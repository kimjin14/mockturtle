module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 , x147 , x148 , x149 , x150 , x151 , x152 , x153 , x154 , x155 , x156 , x157 , x158 , x159 , x160 , x161 , x162 , x163 , x164 , x165 , x166 , x167 , x168 , x169 , x170 , x171 , x172 , x173 , x174 , x175 , x176 , x177 , x178 , x179 , x180 , x181 , x182 , x183 , x184 , x185 , x186 , x187 , x188 , x189 , x190 , x191 , x192 , x193 , x194 , x195 , x196 , x197 , x198 , x199 , x200 , x201 , x202 , x203 , x204 , x205 , x206 , x207 , x208 , x209 , x210 , x211 , x212 , x213 , x214 , x215 , x216 , x217 , x218 , x219 , x220 , x221 , x222 , x223 , x224 , x225 , x226 , x227 , x228 , x229 , x230 , x231 , x232 , x233 , x234 , x235 , x236 , x237 , x238 , x239 , x240 , x241 , x242 , x243 , x244 , x245 , x246 , x247 , x248 , x249 , x250 , x251 , x252 , x253 , x254 , x255 , x256 , x257 , x258 , x259 , x260 , x261 , x262 , x263 , x264 , x265 , x266 , x267 , x268 , x269 , x270 , x271 , x272 , x273 , x274 , x275 , x276 , x277 , x278 , x279 , x280 , x281 , x282 , x283 , x284 , x285 , x286 , x287 , x288 , x289 , x290 , x291 , x292 , x293 , x294 , x295 , x296 , x297 , x298 , x299 , x300 , x301 , x302 , x303 , x304 , x305 , x306 , x307 , x308 , x309 , x310 , x311 , x312 , x313 , x314 , x315 , x316 , x317 , x318 , x319 , x320 , x321 , x322 , x323 , x324 , x325 , x326 , x327 , x328 , x329 , x330 , x331 , x332 , x333 , x334 , x335 , x336 , x337 , x338 , x339 , x340 , x341 , x342 , x343 , x344 , x345 , x346 , x347 , x348 , x349 , x350 , x351 , x352 , x353 , x354 , x355 , x356 , x357 , x358 , x359 , x360 , x361 , x362 , x363 , x364 , x365 , x366 , x367 , x368 , x369 , x370 , x371 , x372 , x373 , x374 , x375 , x376 , x377 , x378 , x379 , x380 , x381 , x382 , x383 , x384 , x385 , x386 , x387 , x388 , x389 , x390 , x391 , x392 , x393 , x394 , x395 , x396 , x397 , x398 , x399 , x400 , x401 , x402 , x403 , x404 , x405 , x406 , x407 , x408 , x409 , x410 , x411 , x412 , x413 , x414 , x415 , x416 , x417 , x418 , x419 , x420 , x421 , x422 , x423 , x424 , x425 , x426 , x427 , x428 , x429 , x430 , x431 , x432 , x433 , x434 , x435 , x436 , x437 , x438 , x439 , x440 , x441 , x442 , x443 , x444 , x445 , x446 , x447 , x448 , x449 , x450 , x451 , x452 , x453 , x454 , x455 , x456 , x457 , x458 , x459 , x460 , x461 , x462 , x463 , x464 , x465 , x466 , x467 , x468 , x469 , x470 , x471 , x472 , x473 , x474 , x475 , x476 , x477 , x478 , x479 , x480 , x481 , x482 , x483 , x484 , x485 , x486 , x487 , x488 , x489 , x490 , x491 , x492 , x493 , x494 , x495 , x496 , x497 , x498 , x499 , x500 , x501 , x502 , x503 , x504 , x505 , x506 , x507 , x508 , x509 , x510 , x511 , x512 , x513 , x514 , x515 , x516 , x517 , x518 , x519 , x520 , x521 , x522 , x523 , x524 , x525 , x526 , x527 , x528 , x529 , x530 , x531 , x532 , x533 , x534 , x535 , x536 , x537 , x538 , x539 , x540 , x541 , x542 , x543 , x544 , x545 , x546 , x547 , x548 , x549 , x550 , x551 , x552 , x553 , x554 , x555 , x556 , x557 , x558 , x559 , x560 , x561 , x562 , x563 , x564 , x565 , x566 , x567 , x568 , x569 , x570 , x571 , x572 , x573 , x574 , x575 , x576 , x577 , x578 , x579 , x580 , x581 , x582 , x583 , x584 , x585 , x586 , x587 , x588 , x589 , x590 , x591 , x592 , x593 , x594 , x595 , x596 , x597 , x598 , x599 , x600 , x601 , x602 , x603 , x604 , x605 , x606 , x607 , x608 , x609 , x610 , x611 , x612 , x613 , x614 , x615 , x616 , x617 , x618 , x619 , x620 , x621 , x622 , x623 , x624 , x625 , x626 , x627 , x628 , x629 , x630 , x631 , x632 , x633 , x634 , x635 , x636 , x637 , x638 , x639 , x640 , x641 , x642 , x643 , x644 , x645 , x646 , x647 , x648 , x649 , x650 , x651 , x652 , x653 , x654 , x655 , x656 , x657 , x658 , x659 , x660 , x661 , x662 , x663 , x664 , x665 , x666 , x667 , x668 , x669 , x670 , x671 , x672 , x673 , x674 , x675 , x676 , x677 , x678 , x679 , x680 , x681 , x682 , x683 , x684 , x685 , x686 , x687 , x688 , x689 , x690 , x691 , x692 , x693 , x694 , x695 , x696 , x697 , x698 , x699 , x700 , x701 , x702 , x703 , x704 , x705 , x706 , x707 , x708 , x709 , x710 , x711 , x712 , x713 , x714 , x715 , x716 , x717 , x718 , x719 , x720 , x721 , x722 , x723 , x724 , x725 , x726 , x727 , x728 , x729 , x730 , x731 , x732 , x733 , x734 , x735 , x736 , x737 , x738 , x739 , x740 , x741 , x742 , x743 , x744 , x745 , x746 , x747 , x748 , x749 , x750 , x751 , x752 , x753 , x754 , x755 , x756 , x757 , x758 , x759 , x760 , x761 , x762 , x763 , x764 , x765 , x766 , x767 , x768 , x769 , x770 , x771 , x772 , x773 , x774 , x775 , x776 , x777 , x778 , x779 , x780 , x781 , x782 , x783 , x784 , x785 , x786 , x787 , x788 , x789 , x790 , x791 , x792 , x793 , x794 , x795 , x796 , x797 , x798 , x799 , x800 , x801 , x802 , x803 , x804 , x805 , x806 , x807 , x808 , x809 , x810 , x811 , x812 , x813 , x814 , x815 , x816 , x817 , x818 , x819 , x820 , x821 , x822 , x823 , x824 , x825 , x826 , x827 , x828 , x829 , x830 , x831 , x832 , x833 , x834 , x835 , x836 , x837 , x838 , x839 , x840 , x841 , x842 , x843 , x844 , x845 , x846 , x847 , x848 , x849 , x850 , x851 , x852 , x853 , x854 , x855 , x856 , x857 , x858 , x859 , x860 , x861 , x862 , x863 , x864 , x865 , x866 , x867 , x868 , x869 , x870 , x871 , x872 , x873 , x874 , x875 , x876 , x877 , x878 , x879 , x880 , x881 , x882 , x883 , x884 , x885 , x886 , x887 , x888 , x889 , x890 , x891 , x892 , x893 , x894 , x895 , x896 , x897 , x898 , x899 , x900 , x901 , x902 , x903 , x904 , x905 , x906 , x907 , x908 , x909 , x910 , x911 , x912 , x913 , x914 , x915 , x916 , x917 , x918 , x919 , x920 , x921 , x922 , x923 , x924 , x925 , x926 , x927 , x928 , x929 , x930 , x931 , x932 , x933 , x934 , x935 , x936 , x937 , x938 , x939 , x940 , x941 , x942 , x943 , x944 , x945 , x946 , x947 , x948 , x949 , x950 , x951 , x952 , x953 , x954 , x955 , x956 , x957 , x958 , x959 , x960 , x961 , x962 , x963 , x964 , x965 , x966 , x967 , x968 , x969 , x970 , x971 , x972 , x973 , x974 , x975 , x976 , x977 , x978 , x979 , x980 , x981 , x982 , x983 , x984 , x985 , x986 , x987 , x988 , x989 , x990 , x991 , x992 , x993 , x994 , x995 , x996 , x997 , x998 , x999 , x1000 , x1001 , x1002 , x1003 , x1004 , x1005 , x1006 , x1007 , x1008 , x1009 , x1010 , x1011 , x1012 , x1013 , x1014 , x1015 , x1016 , x1017 , x1018 , x1019 , x1020 , x1021 , x1022 , x1023 , x1024 , x1025 , x1026 , x1027 , x1028 , x1029 , x1030 , x1031 , x1032 , x1033 , x1034 , x1035 , x1036 , x1037 , x1038 , x1039 , x1040 , x1041 , x1042 , x1043 , x1044 , x1045 , x1046 , x1047 , x1048 , x1049 , x1050 , x1051 , x1052 , x1053 , x1054 , x1055 , x1056 , x1057 , x1058 , x1059 , x1060 , x1061 , x1062 , x1063 , x1064 , x1065 , x1066 , x1067 , x1068 , x1069 , x1070 , x1071 , x1072 , x1073 , x1074 , x1075 , x1076 , x1077 , x1078 , x1079 , x1080 , x1081 , x1082 , x1083 , x1084 , x1085 , x1086 , x1087 , x1088 , x1089 , x1090 , x1091 , x1092 , x1093 , x1094 , x1095 , x1096 , x1097 , x1098 , x1099 , x1100 , x1101 , x1102 , x1103 , x1104 , x1105 , x1106 , x1107 , x1108 , x1109 , x1110 , x1111 , x1112 , x1113 , x1114 , x1115 , x1116 , x1117 , x1118 , x1119 , x1120 , x1121 , x1122 , x1123 , x1124 , x1125 , x1126 , x1127 , x1128 , x1129 , x1130 , x1131 , x1132 , x1133 , x1134 , x1135 , x1136 , x1137 , x1138 , x1139 , x1140 , x1141 , x1142 , x1143 , x1144 , x1145 , x1146 , x1147 , x1148 , x1149 , x1150 , x1151 , x1152 , x1153 , x1154 , x1155 , x1156 , x1157 , x1158 , x1159 , x1160 , x1161 , x1162 , x1163 , x1164 , x1165 , x1166 , x1167 , x1168 , x1169 , x1170 , x1171 , x1172 , x1173 , x1174 , x1175 , x1176 , x1177 , x1178 , x1179 , x1180 , x1181 , x1182 , x1183 , x1184 , x1185 , x1186 , x1187 , x1188 , x1189 , x1190 , x1191 , x1192 , x1193 , x1194 , x1195 , x1196 , x1197 , x1198 , x1199 , x1200 , x1201 , x1202 , x1203 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 , y128 , y129 , y130 , y131 , y132 , y133 , y134 , y135 , y136 , y137 , y138 , y139 , y140 , y141 , y142 , y143 , y144 , y145 , y146 , y147 , y148 , y149 , y150 , y151 , y152 , y153 , y154 , y155 , y156 , y157 , y158 , y159 , y160 , y161 , y162 , y163 , y164 , y165 , y166 , y167 , y168 , y169 , y170 , y171 , y172 , y173 , y174 , y175 , y176 , y177 , y178 , y179 , y180 , y181 , y182 , y183 , y184 , y185 , y186 , y187 , y188 , y189 , y190 , y191 , y192 , y193 , y194 , y195 , y196 , y197 , y198 , y199 , y200 , y201 , y202 , y203 , y204 , y205 , y206 , y207 , y208 , y209 , y210 , y211 , y212 , y213 , y214 , y215 , y216 , y217 , y218 , y219 , y220 , y221 , y222 , y223 , y224 , y225 , y226 , y227 , y228 , y229 , y230 , y231 , y232 , y233 , y234 , y235 , y236 , y237 , y238 , y239 , y240 , y241 , y242 , y243 , y244 , y245 , y246 , y247 , y248 , y249 , y250 , y251 , y252 , y253 , y254 , y255 , y256 , y257 , y258 , y259 , y260 , y261 , y262 , y263 , y264 , y265 , y266 , y267 , y268 , y269 , y270 , y271 , y272 , y273 , y274 , y275 , y276 , y277 , y278 , y279 , y280 , y281 , y282 , y283 , y284 , y285 , y286 , y287 , y288 , y289 , y290 , y291 , y292 , y293 , y294 , y295 , y296 , y297 , y298 , y299 , y300 , y301 , y302 , y303 , y304 , y305 , y306 , y307 , y308 , y309 , y310 , y311 , y312 , y313 , y314 , y315 , y316 , y317 , y318 , y319 , y320 , y321 , y322 , y323 , y324 , y325 , y326 , y327 , y328 , y329 , y330 , y331 , y332 , y333 , y334 , y335 , y336 , y337 , y338 , y339 , y340 , y341 , y342 , y343 , y344 , y345 , y346 , y347 , y348 , y349 , y350 , y351 , y352 , y353 , y354 , y355 , y356 , y357 , y358 , y359 , y360 , y361 , y362 , y363 , y364 , y365 , y366 , y367 , y368 , y369 , y370 , y371 , y372 , y373 , y374 , y375 , y376 , y377 , y378 , y379 , y380 , y381 , y382 , y383 , y384 , y385 , y386 , y387 , y388 , y389 , y390 , y391 , y392 , y393 , y394 , y395 , y396 , y397 , y398 , y399 , y400 , y401 , y402 , y403 , y404 , y405 , y406 , y407 , y408 , y409 , y410 , y411 , y412 , y413 , y414 , y415 , y416 , y417 , y418 , y419 , y420 , y421 , y422 , y423 , y424 , y425 , y426 , y427 , y428 , y429 , y430 , y431 , y432 , y433 , y434 , y435 , y436 , y437 , y438 , y439 , y440 , y441 , y442 , y443 , y444 , y445 , y446 , y447 , y448 , y449 , y450 , y451 , y452 , y453 , y454 , y455 , y456 , y457 , y458 , y459 , y460 , y461 , y462 , y463 , y464 , y465 , y466 , y467 , y468 , y469 , y470 , y471 , y472 , y473 , y474 , y475 , y476 , y477 , y478 , y479 , y480 , y481 , y482 , y483 , y484 , y485 , y486 , y487 , y488 , y489 , y490 , y491 , y492 , y493 , y494 , y495 , y496 , y497 , y498 , y499 , y500 , y501 , y502 , y503 , y504 , y505 , y506 , y507 , y508 , y509 , y510 , y511 , y512 , y513 , y514 , y515 , y516 , y517 , y518 , y519 , y520 , y521 , y522 , y523 , y524 , y525 , y526 , y527 , y528 , y529 , y530 , y531 , y532 , y533 , y534 , y535 , y536 , y537 , y538 , y539 , y540 , y541 , y542 , y543 , y544 , y545 , y546 , y547 , y548 , y549 , y550 , y551 , y552 , y553 , y554 , y555 , y556 , y557 , y558 , y559 , y560 , y561 , y562 , y563 , y564 , y565 , y566 , y567 , y568 , y569 , y570 , y571 , y572 , y573 , y574 , y575 , y576 , y577 , y578 , y579 , y580 , y581 , y582 , y583 , y584 , y585 , y586 , y587 , y588 , y589 , y590 , y591 , y592 , y593 , y594 , y595 , y596 , y597 , y598 , y599 , y600 , y601 , y602 , y603 , y604 , y605 , y606 , y607 , y608 , y609 , y610 , y611 , y612 , y613 , y614 , y615 , y616 , y617 , y618 , y619 , y620 , y621 , y622 , y623 , y624 , y625 , y626 , y627 , y628 , y629 , y630 , y631 , y632 , y633 , y634 , y635 , y636 , y637 , y638 , y639 , y640 , y641 , y642 , y643 , y644 , y645 , y646 , y647 , y648 , y649 , y650 , y651 , y652 , y653 , y654 , y655 , y656 , y657 , y658 , y659 , y660 , y661 , y662 , y663 , y664 , y665 , y666 , y667 , y668 , y669 , y670 , y671 , y672 , y673 , y674 , y675 , y676 , y677 , y678 , y679 , y680 , y681 , y682 , y683 , y684 , y685 , y686 , y687 , y688 , y689 , y690 , y691 , y692 , y693 , y694 , y695 , y696 , y697 , y698 , y699 , y700 , y701 , y702 , y703 , y704 , y705 , y706 , y707 , y708 , y709 , y710 , y711 , y712 , y713 , y714 , y715 , y716 , y717 , y718 , y719 , y720 , y721 , y722 , y723 , y724 , y725 , y726 , y727 , y728 , y729 , y730 , y731 , y732 , y733 , y734 , y735 , y736 , y737 , y738 , y739 , y740 , y741 , y742 , y743 , y744 , y745 , y746 , y747 , y748 , y749 , y750 , y751 , y752 , y753 , y754 , y755 , y756 , y757 , y758 , y759 , y760 , y761 , y762 , y763 , y764 , y765 , y766 , y767 , y768 , y769 , y770 , y771 , y772 , y773 , y774 , y775 , y776 , y777 , y778 , y779 , y780 , y781 , y782 , y783 , y784 , y785 , y786 , y787 , y788 , y789 , y790 , y791 , y792 , y793 , y794 , y795 , y796 , y797 , y798 , y799 , y800 , y801 , y802 , y803 , y804 , y805 , y806 , y807 , y808 , y809 , y810 , y811 , y812 , y813 , y814 , y815 , y816 , y817 , y818 , y819 , y820 , y821 , y822 , y823 , y824 , y825 , y826 , y827 , y828 , y829 , y830 , y831 , y832 , y833 , y834 , y835 , y836 , y837 , y838 , y839 , y840 , y841 , y842 , y843 , y844 , y845 , y846 , y847 , y848 , y849 , y850 , y851 , y852 , y853 , y854 , y855 , y856 , y857 , y858 , y859 , y860 , y861 , y862 , y863 , y864 , y865 , y866 , y867 , y868 , y869 , y870 , y871 , y872 , y873 , y874 , y875 , y876 , y877 , y878 , y879 , y880 , y881 , y882 , y883 , y884 , y885 , y886 , y887 , y888 , y889 , y890 , y891 , y892 , y893 , y894 , y895 , y896 , y897 , y898 , y899 , y900 , y901 , y902 , y903 , y904 , y905 , y906 , y907 , y908 , y909 , y910 , y911 , y912 , y913 , y914 , y915 , y916 , y917 , y918 , y919 , y920 , y921 , y922 , y923 , y924 , y925 , y926 , y927 , y928 , y929 , y930 , y931 , y932 , y933 , y934 , y935 , y936 , y937 , y938 , y939 , y940 , y941 , y942 , y943 , y944 , y945 , y946 , y947 , y948 , y949 , y950 , y951 , y952 , y953 , y954 , y955 , y956 , y957 , y958 , y959 , y960 , y961 , y962 , y963 , y964 , y965 , y966 , y967 , y968 , y969 , y970 , y971 , y972 , y973 , y974 , y975 , y976 , y977 , y978 , y979 , y980 , y981 , y982 , y983 , y984 , y985 , y986 , y987 , y988 , y989 , y990 , y991 , y992 , y993 , y994 , y995 , y996 , y997 , y998 , y999 , y1000 , y1001 , y1002 , y1003 , y1004 , y1005 , y1006 , y1007 , y1008 , y1009 , y1010 , y1011 , y1012 , y1013 , y1014 , y1015 , y1016 , y1017 , y1018 , y1019 , y1020 , y1021 , y1022 , y1023 , y1024 , y1025 , y1026 , y1027 , y1028 , y1029 , y1030 , y1031 , y1032 , y1033 , y1034 , y1035 , y1036 , y1037 , y1038 , y1039 , y1040 , y1041 , y1042 , y1043 , y1044 , y1045 , y1046 , y1047 , y1048 , y1049 , y1050 , y1051 , y1052 , y1053 , y1054 , y1055 , y1056 , y1057 , y1058 , y1059 , y1060 , y1061 , y1062 , y1063 , y1064 , y1065 , y1066 , y1067 , y1068 , y1069 , y1070 , y1071 , y1072 , y1073 , y1074 , y1075 , y1076 , y1077 , y1078 , y1079 , y1080 , y1081 , y1082 , y1083 , y1084 , y1085 , y1086 , y1087 , y1088 , y1089 , y1090 , y1091 , y1092 , y1093 , y1094 , y1095 , y1096 , y1097 , y1098 , y1099 , y1100 , y1101 , y1102 , y1103 , y1104 , y1105 , y1106 , y1107 , y1108 , y1109 , y1110 , y1111 , y1112 , y1113 , y1114 , y1115 , y1116 , y1117 , y1118 , y1119 , y1120 , y1121 , y1122 , y1123 , y1124 , y1125 , y1126 , y1127 , y1128 , y1129 , y1130 , y1131 , y1132 , y1133 , y1134 , y1135 , y1136 , y1137 , y1138 , y1139 , y1140 , y1141 , y1142 , y1143 , y1144 , y1145 , y1146 , y1147 , y1148 , y1149 , y1150 , y1151 , y1152 , y1153 , y1154 , y1155 , y1156 , y1157 , y1158 , y1159 , y1160 , y1161 , y1162 , y1163 , y1164 , y1165 , y1166 , y1167 , y1168 , y1169 , y1170 , y1171 , y1172 , y1173 , y1174 , y1175 , y1176 , y1177 , y1178 , y1179 , y1180 , y1181 , y1182 , y1183 , y1184 , y1185 , y1186 , y1187 , y1188 , y1189 , y1190 , y1191 , y1192 , y1193 , y1194 , y1195 , y1196 , y1197 , y1198 , y1199 , y1200 , y1201 , y1202 , y1203 , y1204 , y1205 , y1206 , y1207 , y1208 , y1209 , y1210 , y1211 , y1212 , y1213 , y1214 , y1215 , y1216 , y1217 , y1218 , y1219 , y1220 , y1221 , y1222 , y1223 , y1224 , y1225 , y1226 , y1227 , y1228 , y1229 , y1230 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 , x147 , x148 , x149 , x150 , x151 , x152 , x153 , x154 , x155 , x156 , x157 , x158 , x159 , x160 , x161 , x162 , x163 , x164 , x165 , x166 , x167 , x168 , x169 , x170 , x171 , x172 , x173 , x174 , x175 , x176 , x177 , x178 , x179 , x180 , x181 , x182 , x183 , x184 , x185 , x186 , x187 , x188 , x189 , x190 , x191 , x192 , x193 , x194 , x195 , x196 , x197 , x198 , x199 , x200 , x201 , x202 , x203 , x204 , x205 , x206 , x207 , x208 , x209 , x210 , x211 , x212 , x213 , x214 , x215 , x216 , x217 , x218 , x219 , x220 , x221 , x222 , x223 , x224 , x225 , x226 , x227 , x228 , x229 , x230 , x231 , x232 , x233 , x234 , x235 , x236 , x237 , x238 , x239 , x240 , x241 , x242 , x243 , x244 , x245 , x246 , x247 , x248 , x249 , x250 , x251 , x252 , x253 , x254 , x255 , x256 , x257 , x258 , x259 , x260 , x261 , x262 , x263 , x264 , x265 , x266 , x267 , x268 , x269 , x270 , x271 , x272 , x273 , x274 , x275 , x276 , x277 , x278 , x279 , x280 , x281 , x282 , x283 , x284 , x285 , x286 , x287 , x288 , x289 , x290 , x291 , x292 , x293 , x294 , x295 , x296 , x297 , x298 , x299 , x300 , x301 , x302 , x303 , x304 , x305 , x306 , x307 , x308 , x309 , x310 , x311 , x312 , x313 , x314 , x315 , x316 , x317 , x318 , x319 , x320 , x321 , x322 , x323 , x324 , x325 , x326 , x327 , x328 , x329 , x330 , x331 , x332 , x333 , x334 , x335 , x336 , x337 , x338 , x339 , x340 , x341 , x342 , x343 , x344 , x345 , x346 , x347 , x348 , x349 , x350 , x351 , x352 , x353 , x354 , x355 , x356 , x357 , x358 , x359 , x360 , x361 , x362 , x363 , x364 , x365 , x366 , x367 , x368 , x369 , x370 , x371 , x372 , x373 , x374 , x375 , x376 , x377 , x378 , x379 , x380 , x381 , x382 , x383 , x384 , x385 , x386 , x387 , x388 , x389 , x390 , x391 , x392 , x393 , x394 , x395 , x396 , x397 , x398 , x399 , x400 , x401 , x402 , x403 , x404 , x405 , x406 , x407 , x408 , x409 , x410 , x411 , x412 , x413 , x414 , x415 , x416 , x417 , x418 , x419 , x420 , x421 , x422 , x423 , x424 , x425 , x426 , x427 , x428 , x429 , x430 , x431 , x432 , x433 , x434 , x435 , x436 , x437 , x438 , x439 , x440 , x441 , x442 , x443 , x444 , x445 , x446 , x447 , x448 , x449 , x450 , x451 , x452 , x453 , x454 , x455 , x456 , x457 , x458 , x459 , x460 , x461 , x462 , x463 , x464 , x465 , x466 , x467 , x468 , x469 , x470 , x471 , x472 , x473 , x474 , x475 , x476 , x477 , x478 , x479 , x480 , x481 , x482 , x483 , x484 , x485 , x486 , x487 , x488 , x489 , x490 , x491 , x492 , x493 , x494 , x495 , x496 , x497 , x498 , x499 , x500 , x501 , x502 , x503 , x504 , x505 , x506 , x507 , x508 , x509 , x510 , x511 , x512 , x513 , x514 , x515 , x516 , x517 , x518 , x519 , x520 , x521 , x522 , x523 , x524 , x525 , x526 , x527 , x528 , x529 , x530 , x531 , x532 , x533 , x534 , x535 , x536 , x537 , x538 , x539 , x540 , x541 , x542 , x543 , x544 , x545 , x546 , x547 , x548 , x549 , x550 , x551 , x552 , x553 , x554 , x555 , x556 , x557 , x558 , x559 , x560 , x561 , x562 , x563 , x564 , x565 , x566 , x567 , x568 , x569 , x570 , x571 , x572 , x573 , x574 , x575 , x576 , x577 , x578 , x579 , x580 , x581 , x582 , x583 , x584 , x585 , x586 , x587 , x588 , x589 , x590 , x591 , x592 , x593 , x594 , x595 , x596 , x597 , x598 , x599 , x600 , x601 , x602 , x603 , x604 , x605 , x606 , x607 , x608 , x609 , x610 , x611 , x612 , x613 , x614 , x615 , x616 , x617 , x618 , x619 , x620 , x621 , x622 , x623 , x624 , x625 , x626 , x627 , x628 , x629 , x630 , x631 , x632 , x633 , x634 , x635 , x636 , x637 , x638 , x639 , x640 , x641 , x642 , x643 , x644 , x645 , x646 , x647 , x648 , x649 , x650 , x651 , x652 , x653 , x654 , x655 , x656 , x657 , x658 , x659 , x660 , x661 , x662 , x663 , x664 , x665 , x666 , x667 , x668 , x669 , x670 , x671 , x672 , x673 , x674 , x675 , x676 , x677 , x678 , x679 , x680 , x681 , x682 , x683 , x684 , x685 , x686 , x687 , x688 , x689 , x690 , x691 , x692 , x693 , x694 , x695 , x696 , x697 , x698 , x699 , x700 , x701 , x702 , x703 , x704 , x705 , x706 , x707 , x708 , x709 , x710 , x711 , x712 , x713 , x714 , x715 , x716 , x717 , x718 , x719 , x720 , x721 , x722 , x723 , x724 , x725 , x726 , x727 , x728 , x729 , x730 , x731 , x732 , x733 , x734 , x735 , x736 , x737 , x738 , x739 , x740 , x741 , x742 , x743 , x744 , x745 , x746 , x747 , x748 , x749 , x750 , x751 , x752 , x753 , x754 , x755 , x756 , x757 , x758 , x759 , x760 , x761 , x762 , x763 , x764 , x765 , x766 , x767 , x768 , x769 , x770 , x771 , x772 , x773 , x774 , x775 , x776 , x777 , x778 , x779 , x780 , x781 , x782 , x783 , x784 , x785 , x786 , x787 , x788 , x789 , x790 , x791 , x792 , x793 , x794 , x795 , x796 , x797 , x798 , x799 , x800 , x801 , x802 , x803 , x804 , x805 , x806 , x807 , x808 , x809 , x810 , x811 , x812 , x813 , x814 , x815 , x816 , x817 , x818 , x819 , x820 , x821 , x822 , x823 , x824 , x825 , x826 , x827 , x828 , x829 , x830 , x831 , x832 , x833 , x834 , x835 , x836 , x837 , x838 , x839 , x840 , x841 , x842 , x843 , x844 , x845 , x846 , x847 , x848 , x849 , x850 , x851 , x852 , x853 , x854 , x855 , x856 , x857 , x858 , x859 , x860 , x861 , x862 , x863 , x864 , x865 , x866 , x867 , x868 , x869 , x870 , x871 , x872 , x873 , x874 , x875 , x876 , x877 , x878 , x879 , x880 , x881 , x882 , x883 , x884 , x885 , x886 , x887 , x888 , x889 , x890 , x891 , x892 , x893 , x894 , x895 , x896 , x897 , x898 , x899 , x900 , x901 , x902 , x903 , x904 , x905 , x906 , x907 , x908 , x909 , x910 , x911 , x912 , x913 , x914 , x915 , x916 , x917 , x918 , x919 , x920 , x921 , x922 , x923 , x924 , x925 , x926 , x927 , x928 , x929 , x930 , x931 , x932 , x933 , x934 , x935 , x936 , x937 , x938 , x939 , x940 , x941 , x942 , x943 , x944 , x945 , x946 , x947 , x948 , x949 , x950 , x951 , x952 , x953 , x954 , x955 , x956 , x957 , x958 , x959 , x960 , x961 , x962 , x963 , x964 , x965 , x966 , x967 , x968 , x969 , x970 , x971 , x972 , x973 , x974 , x975 , x976 , x977 , x978 , x979 , x980 , x981 , x982 , x983 , x984 , x985 , x986 , x987 , x988 , x989 , x990 , x991 , x992 , x993 , x994 , x995 , x996 , x997 , x998 , x999 , x1000 , x1001 , x1002 , x1003 , x1004 , x1005 , x1006 , x1007 , x1008 , x1009 , x1010 , x1011 , x1012 , x1013 , x1014 , x1015 , x1016 , x1017 , x1018 , x1019 , x1020 , x1021 , x1022 , x1023 , x1024 , x1025 , x1026 , x1027 , x1028 , x1029 , x1030 , x1031 , x1032 , x1033 , x1034 , x1035 , x1036 , x1037 , x1038 , x1039 , x1040 , x1041 , x1042 , x1043 , x1044 , x1045 , x1046 , x1047 , x1048 , x1049 , x1050 , x1051 , x1052 , x1053 , x1054 , x1055 , x1056 , x1057 , x1058 , x1059 , x1060 , x1061 , x1062 , x1063 , x1064 , x1065 , x1066 , x1067 , x1068 , x1069 , x1070 , x1071 , x1072 , x1073 , x1074 , x1075 , x1076 , x1077 , x1078 , x1079 , x1080 , x1081 , x1082 , x1083 , x1084 , x1085 , x1086 , x1087 , x1088 , x1089 , x1090 , x1091 , x1092 , x1093 , x1094 , x1095 , x1096 , x1097 , x1098 , x1099 , x1100 , x1101 , x1102 , x1103 , x1104 , x1105 , x1106 , x1107 , x1108 , x1109 , x1110 , x1111 , x1112 , x1113 , x1114 , x1115 , x1116 , x1117 , x1118 , x1119 , x1120 , x1121 , x1122 , x1123 , x1124 , x1125 , x1126 , x1127 , x1128 , x1129 , x1130 , x1131 , x1132 , x1133 , x1134 , x1135 , x1136 , x1137 , x1138 , x1139 , x1140 , x1141 , x1142 , x1143 , x1144 , x1145 , x1146 , x1147 , x1148 , x1149 , x1150 , x1151 , x1152 , x1153 , x1154 , x1155 , x1156 , x1157 , x1158 , x1159 , x1160 , x1161 , x1162 , x1163 , x1164 , x1165 , x1166 , x1167 , x1168 , x1169 , x1170 , x1171 , x1172 , x1173 , x1174 , x1175 , x1176 , x1177 , x1178 , x1179 , x1180 , x1181 , x1182 , x1183 , x1184 , x1185 , x1186 , x1187 , x1188 , x1189 , x1190 , x1191 , x1192 , x1193 , x1194 , x1195 , x1196 , x1197 , x1198 , x1199 , x1200 , x1201 , x1202 , x1203 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 , y128 , y129 , y130 , y131 , y132 , y133 , y134 , y135 , y136 , y137 , y138 , y139 , y140 , y141 , y142 , y143 , y144 , y145 , y146 , y147 , y148 , y149 , y150 , y151 , y152 , y153 , y154 , y155 , y156 , y157 , y158 , y159 , y160 , y161 , y162 , y163 , y164 , y165 , y166 , y167 , y168 , y169 , y170 , y171 , y172 , y173 , y174 , y175 , y176 , y177 , y178 , y179 , y180 , y181 , y182 , y183 , y184 , y185 , y186 , y187 , y188 , y189 , y190 , y191 , y192 , y193 , y194 , y195 , y196 , y197 , y198 , y199 , y200 , y201 , y202 , y203 , y204 , y205 , y206 , y207 , y208 , y209 , y210 , y211 , y212 , y213 , y214 , y215 , y216 , y217 , y218 , y219 , y220 , y221 , y222 , y223 , y224 , y225 , y226 , y227 , y228 , y229 , y230 , y231 , y232 , y233 , y234 , y235 , y236 , y237 , y238 , y239 , y240 , y241 , y242 , y243 , y244 , y245 , y246 , y247 , y248 , y249 , y250 , y251 , y252 , y253 , y254 , y255 , y256 , y257 , y258 , y259 , y260 , y261 , y262 , y263 , y264 , y265 , y266 , y267 , y268 , y269 , y270 , y271 , y272 , y273 , y274 , y275 , y276 , y277 , y278 , y279 , y280 , y281 , y282 , y283 , y284 , y285 , y286 , y287 , y288 , y289 , y290 , y291 , y292 , y293 , y294 , y295 , y296 , y297 , y298 , y299 , y300 , y301 , y302 , y303 , y304 , y305 , y306 , y307 , y308 , y309 , y310 , y311 , y312 , y313 , y314 , y315 , y316 , y317 , y318 , y319 , y320 , y321 , y322 , y323 , y324 , y325 , y326 , y327 , y328 , y329 , y330 , y331 , y332 , y333 , y334 , y335 , y336 , y337 , y338 , y339 , y340 , y341 , y342 , y343 , y344 , y345 , y346 , y347 , y348 , y349 , y350 , y351 , y352 , y353 , y354 , y355 , y356 , y357 , y358 , y359 , y360 , y361 , y362 , y363 , y364 , y365 , y366 , y367 , y368 , y369 , y370 , y371 , y372 , y373 , y374 , y375 , y376 , y377 , y378 , y379 , y380 , y381 , y382 , y383 , y384 , y385 , y386 , y387 , y388 , y389 , y390 , y391 , y392 , y393 , y394 , y395 , y396 , y397 , y398 , y399 , y400 , y401 , y402 , y403 , y404 , y405 , y406 , y407 , y408 , y409 , y410 , y411 , y412 , y413 , y414 , y415 , y416 , y417 , y418 , y419 , y420 , y421 , y422 , y423 , y424 , y425 , y426 , y427 , y428 , y429 , y430 , y431 , y432 , y433 , y434 , y435 , y436 , y437 , y438 , y439 , y440 , y441 , y442 , y443 , y444 , y445 , y446 , y447 , y448 , y449 , y450 , y451 , y452 , y453 , y454 , y455 , y456 , y457 , y458 , y459 , y460 , y461 , y462 , y463 , y464 , y465 , y466 , y467 , y468 , y469 , y470 , y471 , y472 , y473 , y474 , y475 , y476 , y477 , y478 , y479 , y480 , y481 , y482 , y483 , y484 , y485 , y486 , y487 , y488 , y489 , y490 , y491 , y492 , y493 , y494 , y495 , y496 , y497 , y498 , y499 , y500 , y501 , y502 , y503 , y504 , y505 , y506 , y507 , y508 , y509 , y510 , y511 , y512 , y513 , y514 , y515 , y516 , y517 , y518 , y519 , y520 , y521 , y522 , y523 , y524 , y525 , y526 , y527 , y528 , y529 , y530 , y531 , y532 , y533 , y534 , y535 , y536 , y537 , y538 , y539 , y540 , y541 , y542 , y543 , y544 , y545 , y546 , y547 , y548 , y549 , y550 , y551 , y552 , y553 , y554 , y555 , y556 , y557 , y558 , y559 , y560 , y561 , y562 , y563 , y564 , y565 , y566 , y567 , y568 , y569 , y570 , y571 , y572 , y573 , y574 , y575 , y576 , y577 , y578 , y579 , y580 , y581 , y582 , y583 , y584 , y585 , y586 , y587 , y588 , y589 , y590 , y591 , y592 , y593 , y594 , y595 , y596 , y597 , y598 , y599 , y600 , y601 , y602 , y603 , y604 , y605 , y606 , y607 , y608 , y609 , y610 , y611 , y612 , y613 , y614 , y615 , y616 , y617 , y618 , y619 , y620 , y621 , y622 , y623 , y624 , y625 , y626 , y627 , y628 , y629 , y630 , y631 , y632 , y633 , y634 , y635 , y636 , y637 , y638 , y639 , y640 , y641 , y642 , y643 , y644 , y645 , y646 , y647 , y648 , y649 , y650 , y651 , y652 , y653 , y654 , y655 , y656 , y657 , y658 , y659 , y660 , y661 , y662 , y663 , y664 , y665 , y666 , y667 , y668 , y669 , y670 , y671 , y672 , y673 , y674 , y675 , y676 , y677 , y678 , y679 , y680 , y681 , y682 , y683 , y684 , y685 , y686 , y687 , y688 , y689 , y690 , y691 , y692 , y693 , y694 , y695 , y696 , y697 , y698 , y699 , y700 , y701 , y702 , y703 , y704 , y705 , y706 , y707 , y708 , y709 , y710 , y711 , y712 , y713 , y714 , y715 , y716 , y717 , y718 , y719 , y720 , y721 , y722 , y723 , y724 , y725 , y726 , y727 , y728 , y729 , y730 , y731 , y732 , y733 , y734 , y735 , y736 , y737 , y738 , y739 , y740 , y741 , y742 , y743 , y744 , y745 , y746 , y747 , y748 , y749 , y750 , y751 , y752 , y753 , y754 , y755 , y756 , y757 , y758 , y759 , y760 , y761 , y762 , y763 , y764 , y765 , y766 , y767 , y768 , y769 , y770 , y771 , y772 , y773 , y774 , y775 , y776 , y777 , y778 , y779 , y780 , y781 , y782 , y783 , y784 , y785 , y786 , y787 , y788 , y789 , y790 , y791 , y792 , y793 , y794 , y795 , y796 , y797 , y798 , y799 , y800 , y801 , y802 , y803 , y804 , y805 , y806 , y807 , y808 , y809 , y810 , y811 , y812 , y813 , y814 , y815 , y816 , y817 , y818 , y819 , y820 , y821 , y822 , y823 , y824 , y825 , y826 , y827 , y828 , y829 , y830 , y831 , y832 , y833 , y834 , y835 , y836 , y837 , y838 , y839 , y840 , y841 , y842 , y843 , y844 , y845 , y846 , y847 , y848 , y849 , y850 , y851 , y852 , y853 , y854 , y855 , y856 , y857 , y858 , y859 , y860 , y861 , y862 , y863 , y864 , y865 , y866 , y867 , y868 , y869 , y870 , y871 , y872 , y873 , y874 , y875 , y876 , y877 , y878 , y879 , y880 , y881 , y882 , y883 , y884 , y885 , y886 , y887 , y888 , y889 , y890 , y891 , y892 , y893 , y894 , y895 , y896 , y897 , y898 , y899 , y900 , y901 , y902 , y903 , y904 , y905 , y906 , y907 , y908 , y909 , y910 , y911 , y912 , y913 , y914 , y915 , y916 , y917 , y918 , y919 , y920 , y921 , y922 , y923 , y924 , y925 , y926 , y927 , y928 , y929 , y930 , y931 , y932 , y933 , y934 , y935 , y936 , y937 , y938 , y939 , y940 , y941 , y942 , y943 , y944 , y945 , y946 , y947 , y948 , y949 , y950 , y951 , y952 , y953 , y954 , y955 , y956 , y957 , y958 , y959 , y960 , y961 , y962 , y963 , y964 , y965 , y966 , y967 , y968 , y969 , y970 , y971 , y972 , y973 , y974 , y975 , y976 , y977 , y978 , y979 , y980 , y981 , y982 , y983 , y984 , y985 , y986 , y987 , y988 , y989 , y990 , y991 , y992 , y993 , y994 , y995 , y996 , y997 , y998 , y999 , y1000 , y1001 , y1002 , y1003 , y1004 , y1005 , y1006 , y1007 , y1008 , y1009 , y1010 , y1011 , y1012 , y1013 , y1014 , y1015 , y1016 , y1017 , y1018 , y1019 , y1020 , y1021 , y1022 , y1023 , y1024 , y1025 , y1026 , y1027 , y1028 , y1029 , y1030 , y1031 , y1032 , y1033 , y1034 , y1035 , y1036 , y1037 , y1038 , y1039 , y1040 , y1041 , y1042 , y1043 , y1044 , y1045 , y1046 , y1047 , y1048 , y1049 , y1050 , y1051 , y1052 , y1053 , y1054 , y1055 , y1056 , y1057 , y1058 , y1059 , y1060 , y1061 , y1062 , y1063 , y1064 , y1065 , y1066 , y1067 , y1068 , y1069 , y1070 , y1071 , y1072 , y1073 , y1074 , y1075 , y1076 , y1077 , y1078 , y1079 , y1080 , y1081 , y1082 , y1083 , y1084 , y1085 , y1086 , y1087 , y1088 , y1089 , y1090 , y1091 , y1092 , y1093 , y1094 , y1095 , y1096 , y1097 , y1098 , y1099 , y1100 , y1101 , y1102 , y1103 , y1104 , y1105 , y1106 , y1107 , y1108 , y1109 , y1110 , y1111 , y1112 , y1113 , y1114 , y1115 , y1116 , y1117 , y1118 , y1119 , y1120 , y1121 , y1122 , y1123 , y1124 , y1125 , y1126 , y1127 , y1128 , y1129 , y1130 , y1131 , y1132 , y1133 , y1134 , y1135 , y1136 , y1137 , y1138 , y1139 , y1140 , y1141 , y1142 , y1143 , y1144 , y1145 , y1146 , y1147 , y1148 , y1149 , y1150 , y1151 , y1152 , y1153 , y1154 , y1155 , y1156 , y1157 , y1158 , y1159 , y1160 , y1161 , y1162 , y1163 , y1164 , y1165 , y1166 , y1167 , y1168 , y1169 , y1170 , y1171 , y1172 , y1173 , y1174 , y1175 , y1176 , y1177 , y1178 , y1179 , y1180 , y1181 , y1182 , y1183 , y1184 , y1185 , y1186 , y1187 , y1188 , y1189 , y1190 , y1191 , y1192 , y1193 , y1194 , y1195 , y1196 , y1197 , y1198 , y1199 , y1200 , y1201 , y1202 , y1203 , y1204 , y1205 , y1206 , y1207 , y1208 , y1209 , y1210 , y1211 , y1212 , y1213 , y1214 , y1215 , y1216 , y1217 , y1218 , y1219 , y1220 , y1221 , y1222 , y1223 , y1224 , y1225 , y1226 , y1227 , y1228 , y1229 , y1230 ;
  wire n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , n3931 , n3932 , n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , n3940 , n3941 , n3942 , n3943 , n3944 , n3945 , n3946 , n3947 , n3948 , n3949 , n3950 , n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , n3970 , n3971 , n3972 , n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , n3980 , n3981 , n3982 , n3983 , n3984 , n3985 , n3986 , n3987 , n3988 , n3989 , n3990 , n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , n4000 , n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , n4009 , n4010 , n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , n4019 , n4020 , n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , n4029 , n4030 , n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , n4039 , n4040 , n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4049 , n4050 , n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , n4059 , n4060 , n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , n4070 , n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , n4079 , n4080 , n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , n4089 , n4090 , n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , n4097 , n4098 , n4099 , n4100 , n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , n4109 , n4110 , n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , n4119 , n4120 , n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , n4129 , n4130 , n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , n4139 , n4140 , n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , n4150 , n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , n4159 , n4160 , n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , n4169 , n4170 , n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , n4179 , n4180 , n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , n4189 , n4190 , n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , n4197 , n4198 , n4199 , n4200 , n4201 , n4202 , n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , n4209 , n4210 , n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , n4217 , n4218 , n4219 , n4220 , n4221 , n4222 , n4223 , n4224 , n4225 , n4226 , n4227 , n4228 , n4229 , n4230 , n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , n4237 , n4238 , n4239 , n4240 , n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , n4247 , n4248 , n4249 , n4250 , n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , n4259 , n4260 , n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , n4269 , n4270 , n4271 , n4272 , n4273 , n4274 , n4275 , n4276 , n4277 , n4278 , n4279 , n4280 , n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , n4289 , n4290 , n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , n4299 , n4300 , n4301 , n4302 , n4303 , n4304 , n4305 , n4306 , n4307 , n4308 , n4309 , n4310 , n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , n4319 , n4320 , n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , n4329 , n4330 , n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , n4340 , n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , n4349 , n4350 , n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , n4360 , n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , n4370 , n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , n4380 , n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , n4390 , n4391 , n4392 , n4393 , n4394 , n4395 , n4396 , n4397 , n4398 , n4399 , n4400 , n4401 , n4402 , n4403 , n4404 , n4405 , n4406 , n4407 , n4408 , n4409 , n4410 , n4411 , n4412 , n4413 , n4414 , n4415 , n4416 , n4417 , n4418 , n4419 , n4420 , n4421 , n4422 , n4423 , n4424 , n4425 , n4426 , n4427 , n4428 , n4429 , n4430 , n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , n4437 , n4438 , n4439 , n4440 , n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , n4449 , n4450 , n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , n4459 , n4460 , n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , n4469 , n4470 , n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , n4479 , n4480 , n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , n4487 , n4488 , n4489 , n4490 , n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , n4497 , n4498 , n4499 , n4500 , n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , n4509 , n4510 , n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , n4519 , n4520 , n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , n4529 , n4530 , n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , n4537 , n4538 , n4539 , n4540 , n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , n4547 , n4548 , n4549 , n4550 , n4551 , n4552 , n4553 , n4554 , n4555 , n4556 , n4557 , n4558 , n4559 , n4560 , n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , n4567 , n4568 , n4569 , n4570 , n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , n4579 , n4580 , n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , n4589 , n4590 , n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , n4597 , n4598 , n4599 , n4600 , n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , n4607 , n4608 , n4609 , n4610 , n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , n4617 , n4618 , n4619 , n4620 , n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , n4627 , n4628 , n4629 , n4630 , n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , n4637 , n4638 , n4639 , n4640 , n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , n4647 , n4648 , n4649 , n4650 , n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , n4657 , n4658 , n4659 , n4660 , n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , n4669 , n4670 , n4671 , n4672 , n4673 , n4674 , n4675 , n4676 , n4677 , n4678 , n4679 , n4680 , n4681 , n4682 , n4683 , n4684 , n4685 , n4686 , n4687 , n4688 , n4689 , n4690 , n4691 , n4692 , n4693 , n4694 , n4695 , n4696 , n4697 , n4698 , n4699 , n4700 , n4701 , n4702 , n4703 , n4704 , n4705 , n4706 , n4707 , n4708 , n4709 , n4710 , n4711 , n4712 , n4713 , n4714 , n4715 , n4716 , n4717 , n4718 , n4719 , n4720 , n4721 , n4722 , n4723 , n4724 , n4725 , n4726 , n4727 , n4728 , n4729 , n4730 , n4731 , n4732 , n4733 , n4734 , n4735 , n4736 , n4737 , n4738 , n4739 , n4740 , n4741 , n4742 , n4743 , n4744 , n4745 , n4746 , n4747 , n4748 , n4749 , n4750 , n4751 , n4752 , n4753 , n4754 , n4755 , n4756 , n4757 , n4758 , n4759 , n4760 , n4761 , n4762 , n4763 , n4764 , n4765 , n4766 , n4767 , n4768 , n4769 , n4770 , n4771 , n4772 , n4773 , n4774 , n4775 , n4776 , n4777 , n4778 , n4779 , n4780 , n4781 , n4782 , n4783 , n4784 , n4785 , n4786 , n4787 , n4788 , n4789 , n4790 , n4791 , n4792 , n4793 , n4794 , n4795 , n4796 , n4797 , n4798 , n4799 , n4800 , n4801 , n4802 , n4803 , n4804 , n4805 , n4806 , n4807 , n4808 , n4809 , n4810 , n4811 , n4812 , n4813 , n4814 , n4815 , n4816 , n4817 , n4818 , n4819 , n4820 , n4821 , n4822 , n4823 , n4824 , n4825 , n4826 , n4827 , n4828 , n4829 , n4830 , n4831 , n4832 , n4833 , n4834 , n4835 , n4836 , n4837 , n4838 , n4839 , n4840 , n4841 , n4842 , n4843 , n4844 , n4845 , n4846 , n4847 , n4848 , n4849 , n4850 , n4851 , n4852 , n4853 , n4854 , n4855 , n4856 , n4857 , n4858 , n4859 , n4860 , n4861 , n4862 , n4863 , n4864 , n4865 , n4866 , n4867 , n4868 , n4869 , n4870 , n4871 , n4872 , n4873 , n4874 , n4875 , n4876 , n4877 , n4878 , n4879 , n4880 , n4881 , n4882 , n4883 , n4884 , n4885 , n4886 , n4887 , n4888 , n4889 , n4890 , n4891 , n4892 , n4893 , n4894 , n4895 , n4896 , n4897 , n4898 , n4899 , n4900 , n4901 , n4902 , n4903 , n4904 , n4905 , n4906 , n4907 , n4908 , n4909 , n4910 , n4911 , n4912 , n4913 , n4914 , n4915 , n4916 , n4917 , n4918 , n4919 , n4920 , n4921 , n4922 , n4923 , n4924 , n4925 , n4926 , n4927 , n4928 , n4929 , n4930 , n4931 , n4932 , n4933 , n4934 , n4935 , n4936 , n4937 , n4938 , n4939 , n4940 , n4941 , n4942 , n4943 , n4944 , n4945 , n4946 , n4947 , n4948 , n4949 , n4950 , n4951 , n4952 , n4953 , n4954 , n4955 , n4956 , n4957 , n4958 , n4959 , n4960 , n4961 , n4962 , n4963 , n4964 , n4965 , n4966 , n4967 , n4968 , n4969 , n4970 , n4971 , n4972 , n4973 , n4974 , n4975 , n4976 , n4977 , n4978 , n4979 , n4980 , n4981 , n4982 , n4983 , n4984 , n4985 , n4986 , n4987 , n4988 , n4989 , n4990 , n4991 , n4992 , n4993 , n4994 , n4995 , n4996 , n4997 , n4998 , n4999 , n5000 , n5001 , n5002 , n5003 , n5004 , n5005 , n5006 , n5007 , n5008 , n5009 , n5010 , n5011 , n5012 , n5013 , n5014 , n5015 , n5016 , n5017 , n5018 , n5019 , n5020 , n5021 , n5022 , n5023 , n5024 , n5025 , n5026 , n5027 , n5028 , n5029 , n5030 , n5031 , n5032 , n5033 , n5034 , n5035 , n5036 , n5037 , n5038 , n5039 , n5040 , n5041 , n5042 , n5043 , n5044 , n5045 , n5046 , n5047 , n5048 , n5049 , n5050 , n5051 , n5052 , n5053 , n5054 , n5055 , n5056 , n5057 , n5058 , n5059 , n5060 , n5061 , n5062 , n5063 , n5064 , n5065 , n5066 , n5067 , n5068 , n5069 , n5070 , n5071 , n5072 , n5073 , n5074 , n5075 , n5076 , n5077 , n5078 , n5079 , n5080 , n5081 , n5082 , n5083 , n5084 , n5085 , n5086 , n5087 , n5088 , n5089 , n5090 , n5091 , n5092 , n5093 , n5094 , n5095 , n5096 , n5097 , n5098 , n5099 , n5100 , n5101 , n5102 , n5103 , n5104 , n5105 , n5106 , n5107 , n5108 , n5109 , n5110 , n5111 , n5112 , n5113 , n5114 , n5115 , n5116 , n5117 , n5118 , n5119 , n5120 , n5121 , n5122 , n5123 , n5124 , n5125 , n5126 , n5127 , n5128 , n5129 , n5130 , n5131 , n5132 , n5133 , n5134 , n5135 , n5136 , n5137 , n5138 , n5139 , n5140 , n5141 , n5142 , n5143 , n5144 , n5145 , n5146 , n5147 , n5148 , n5149 , n5150 , n5151 , n5152 , n5153 , n5154 , n5155 , n5156 , n5157 , n5158 , n5159 , n5160 , n5161 , n5162 , n5163 , n5164 , n5165 , n5166 , n5167 , n5168 , n5169 , n5170 , n5171 , n5172 , n5173 , n5174 , n5175 , n5176 , n5177 , n5178 , n5179 , n5180 , n5181 , n5182 , n5183 , n5184 , n5185 , n5186 , n5187 , n5188 , n5189 , n5190 , n5191 , n5192 , n5193 , n5194 , n5195 , n5196 , n5197 , n5198 , n5199 , n5200 , n5201 , n5202 , n5203 , n5204 , n5205 , n5206 , n5207 , n5208 , n5209 , n5210 , n5211 , n5212 , n5213 , n5214 , n5215 , n5216 , n5217 , n5218 , n5219 , n5220 , n5221 , n5222 , n5223 , n5224 , n5225 , n5226 , n5227 , n5228 , n5229 , n5230 , n5231 , n5232 , n5233 , n5234 , n5235 , n5236 , n5237 , n5238 , n5239 , n5240 , n5241 , n5242 , n5243 , n5244 , n5245 , n5246 , n5247 , n5248 , n5249 , n5250 , n5251 , n5252 , n5253 , n5254 , n5255 , n5256 , n5257 , n5258 , n5259 , n5260 , n5261 , n5262 , n5263 , n5264 , n5265 , n5266 , n5267 , n5268 , n5269 , n5270 , n5271 , n5272 , n5273 , n5274 , n5275 , n5276 , n5277 , n5278 , n5279 , n5280 , n5281 , n5282 , n5283 , n5284 , n5285 , n5286 , n5287 , n5288 , n5289 , n5290 , n5291 , n5292 , n5293 , n5294 , n5295 , n5296 , n5297 , n5298 , n5299 , n5300 , n5301 , n5302 , n5303 , n5304 , n5305 , n5306 , n5307 , n5308 , n5309 , n5310 , n5311 , n5312 , n5313 , n5314 , n5315 , n5316 , n5317 , n5318 , n5319 , n5320 , n5321 , n5322 , n5323 , n5324 , n5325 , n5326 , n5327 , n5328 , n5329 , n5330 , n5331 , n5332 , n5333 , n5334 , n5335 , n5336 , n5337 , n5338 , n5339 , n5340 , n5341 , n5342 , n5343 , n5344 , n5345 , n5346 , n5347 , n5348 , n5349 , n5350 , n5351 , n5352 , n5353 , n5354 , n5355 , n5356 , n5357 , n5358 , n5359 , n5360 , n5361 , n5362 , n5363 , n5364 , n5365 , n5366 , n5367 , n5368 , n5369 , n5370 , n5371 , n5372 , n5373 , n5374 , n5375 , n5376 , n5377 , n5378 , n5379 , n5380 , n5381 , n5382 , n5383 , n5384 , n5385 , n5386 , n5387 , n5388 , n5389 , n5390 , n5391 , n5392 , n5393 , n5394 , n5395 , n5396 , n5397 , n5398 , n5399 , n5400 , n5401 , n5402 , n5403 , n5404 , n5405 , n5406 , n5407 , n5408 , n5409 , n5410 , n5411 , n5412 , n5413 , n5414 , n5415 , n5416 , n5417 , n5418 , n5419 , n5420 , n5421 , n5422 , n5423 , n5424 , n5425 , n5426 , n5427 , n5428 , n5429 , n5430 , n5431 , n5432 , n5433 , n5434 , n5435 , n5436 , n5437 , n5438 , n5439 , n5440 , n5441 , n5442 , n5443 , n5444 , n5445 , n5446 , n5447 , n5448 , n5449 , n5450 , n5451 , n5452 , n5453 , n5454 , n5455 , n5456 , n5457 , n5458 , n5459 , n5460 , n5461 , n5462 , n5463 , n5464 , n5465 , n5466 , n5467 , n5468 , n5469 , n5470 , n5471 , n5472 , n5473 , n5474 , n5475 , n5476 , n5477 , n5478 , n5479 , n5480 , n5481 , n5482 , n5483 , n5484 , n5485 , n5486 , n5487 , n5488 , n5489 , n5490 , n5491 , n5492 , n5493 , n5494 , n5495 , n5496 , n5497 , n5498 , n5499 , n5500 , n5501 , n5502 , n5503 , n5504 , n5505 , n5506 , n5507 , n5508 , n5509 , n5510 , n5511 , n5512 , n5513 , n5514 , n5515 , n5516 , n5517 , n5518 , n5519 , n5520 , n5521 , n5522 , n5523 , n5524 , n5525 , n5526 , n5527 , n5528 , n5529 , n5530 , n5531 , n5532 , n5533 , n5534 , n5535 , n5536 , n5537 , n5538 , n5539 , n5540 , n5541 , n5542 , n5543 , n5544 , n5545 , n5546 , n5547 , n5548 , n5549 , n5550 , n5551 , n5552 , n5553 , n5554 , n5555 , n5556 , n5557 , n5558 , n5559 , n5560 , n5561 , n5562 , n5563 , n5564 , n5565 , n5566 , n5567 , n5568 , n5569 , n5570 , n5571 , n5572 , n5573 , n5574 , n5575 , n5576 , n5577 , n5578 , n5579 , n5580 , n5581 , n5582 , n5583 , n5584 , n5585 , n5586 , n5587 , n5588 , n5589 , n5590 , n5591 , n5592 , n5593 , n5594 , n5595 , n5596 , n5597 , n5598 , n5599 , n5600 , n5601 , n5602 , n5603 , n5604 , n5605 , n5606 , n5607 , n5608 , n5609 , n5610 , n5611 , n5612 , n5613 , n5614 , n5615 , n5616 , n5617 , n5618 , n5619 , n5620 , n5621 , n5622 , n5623 , n5624 , n5625 , n5626 , n5627 , n5628 , n5629 , n5630 , n5631 , n5632 , n5633 , n5634 , n5635 , n5636 , n5637 , n5638 , n5639 , n5640 , n5641 , n5642 , n5643 , n5644 , n5645 , n5646 , n5647 , n5648 , n5649 , n5650 , n5651 , n5652 , n5653 , n5654 , n5655 , n5656 , n5657 , n5658 , n5659 , n5660 , n5661 , n5662 , n5663 , n5664 , n5665 , n5666 , n5667 , n5668 , n5669 , n5670 , n5671 , n5672 , n5673 , n5674 , n5675 , n5676 , n5677 , n5678 , n5679 , n5680 , n5681 , n5682 , n5683 , n5684 , n5685 , n5686 , n5687 , n5688 , n5689 , n5690 , n5691 , n5692 , n5693 , n5694 , n5695 , n5696 , n5697 , n5698 , n5699 , n5700 , n5701 , n5702 , n5703 , n5704 , n5705 , n5706 , n5707 , n5708 , n5709 , n5710 , n5711 , n5712 , n5713 , n5714 , n5715 , n5716 , n5717 , n5718 , n5719 , n5720 , n5721 , n5722 , n5723 , n5724 , n5725 , n5726 , n5727 , n5728 , n5729 , n5730 , n5731 , n5732 , n5733 , n5734 , n5735 , n5736 , n5737 , n5738 , n5739 , n5740 , n5741 , n5742 , n5743 , n5744 , n5745 , n5746 , n5747 , n5748 , n5749 , n5750 , n5751 , n5752 , n5753 , n5754 , n5755 , n5756 , n5757 , n5758 , n5759 , n5760 , n5761 , n5762 , n5763 , n5764 , n5765 , n5766 , n5767 , n5768 , n5769 , n5770 , n5771 , n5772 , n5773 , n5774 , n5775 , n5776 , n5777 , n5778 , n5779 , n5780 , n5781 , n5782 , n5783 , n5784 , n5785 , n5786 , n5787 , n5788 , n5789 , n5790 , n5791 , n5792 , n5793 , n5794 , n5795 , n5796 , n5797 , n5798 , n5799 , n5800 , n5801 , n5802 , n5803 , n5804 , n5805 , n5806 , n5807 , n5808 , n5809 , n5810 , n5811 , n5812 , n5813 , n5814 , n5815 , n5816 , n5817 , n5818 , n5819 , n5820 , n5821 , n5822 , n5823 , n5824 , n5825 , n5826 , n5827 , n5828 , n5829 , n5830 , n5831 , n5832 , n5833 , n5834 , n5835 , n5836 , n5837 , n5838 , n5839 , n5840 , n5841 , n5842 , n5843 , n5844 , n5845 , n5846 , n5847 , n5848 , n5849 , n5850 , n5851 , n5852 , n5853 , n5854 , n5855 , n5856 , n5857 , n5858 , n5859 , n5860 , n5861 , n5862 , n5863 , n5864 , n5865 , n5866 , n5867 , n5868 , n5869 , n5870 , n5871 , n5872 , n5873 , n5874 , n5875 , n5876 , n5877 , n5878 , n5879 , n5880 , n5881 , n5882 , n5883 , n5884 , n5885 , n5886 , n5887 , n5888 , n5889 , n5890 , n5891 , n5892 , n5893 , n5894 , n5895 , n5896 , n5897 , n5898 , n5899 , n5900 , n5901 , n5902 , n5903 , n5904 , n5905 , n5906 , n5907 , n5908 , n5909 , n5910 , n5911 , n5912 , n5913 , n5914 , n5915 , n5916 , n5917 , n5918 , n5919 , n5920 , n5921 , n5922 , n5923 , n5924 , n5925 , n5926 , n5927 , n5928 , n5929 , n5930 , n5931 , n5932 , n5933 , n5934 , n5935 , n5936 , n5937 , n5938 , n5939 , n5940 , n5941 , n5942 , n5943 , n5944 , n5945 , n5946 , n5947 , n5948 , n5949 , n5950 , n5951 , n5952 , n5953 , n5954 , n5955 , n5956 , n5957 , n5958 , n5959 , n5960 , n5961 , n5962 , n5963 , n5964 , n5965 , n5966 , n5967 , n5968 , n5969 , n5970 , n5971 , n5972 , n5973 , n5974 , n5975 , n5976 , n5977 , n5978 , n5979 , n5980 , n5981 , n5982 , n5983 , n5984 , n5985 , n5986 , n5987 , n5988 , n5989 , n5990 , n5991 , n5992 , n5993 , n5994 , n5995 , n5996 , n5997 , n5998 , n5999 , n6000 , n6001 , n6002 , n6003 , n6004 , n6005 , n6006 , n6007 , n6008 , n6009 , n6010 , n6011 , n6012 , n6013 , n6014 , n6015 , n6016 , n6017 , n6018 , n6019 , n6020 , n6021 , n6022 , n6023 , n6024 , n6025 , n6026 , n6027 , n6028 , n6029 , n6030 , n6031 , n6032 , n6033 , n6034 , n6035 , n6036 , n6037 , n6038 , n6039 , n6040 , n6041 , n6042 , n6043 , n6044 , n6045 , n6046 , n6047 , n6048 , n6049 , n6050 , n6051 , n6052 , n6053 , n6054 , n6055 , n6056 , n6057 , n6058 , n6059 , n6060 , n6061 , n6062 , n6063 , n6064 , n6065 , n6066 , n6067 , n6068 , n6069 , n6070 , n6071 , n6072 , n6073 , n6074 , n6075 , n6076 , n6077 , n6078 , n6079 , n6080 , n6081 , n6082 , n6083 , n6084 , n6085 , n6086 , n6087 , n6088 , n6089 , n6090 , n6091 , n6092 , n6093 , n6094 , n6095 , n6096 , n6097 , n6098 , n6099 , n6100 , n6101 , n6102 , n6103 , n6104 , n6105 , n6106 , n6107 , n6108 , n6109 , n6110 , n6111 , n6112 , n6113 , n6114 , n6115 , n6116 , n6117 , n6118 , n6119 , n6120 , n6121 , n6122 , n6123 , n6124 , n6125 , n6126 , n6127 , n6128 , n6129 , n6130 , n6131 , n6132 , n6133 , n6134 , n6135 , n6136 , n6137 , n6138 , n6139 , n6140 , n6141 , n6142 , n6143 , n6144 , n6145 , n6146 , n6147 , n6148 , n6149 , n6150 , n6151 , n6152 , n6153 , n6154 , n6155 , n6156 , n6157 , n6158 , n6159 , n6160 , n6161 , n6162 , n6163 , n6164 , n6165 , n6166 , n6167 , n6168 , n6169 , n6170 , n6171 , n6172 , n6173 , n6174 , n6175 , n6176 , n6177 , n6178 , n6179 , n6180 , n6181 , n6182 , n6183 , n6184 , n6185 , n6186 , n6187 , n6188 , n6189 , n6190 , n6191 , n6192 , n6193 , n6194 , n6195 , n6196 , n6197 , n6198 , n6199 , n6200 , n6201 , n6202 , n6203 , n6204 , n6205 , n6206 , n6207 , n6208 , n6209 , n6210 , n6211 , n6212 , n6213 , n6214 , n6215 , n6216 , n6217 , n6218 , n6219 , n6220 , n6221 , n6222 , n6223 , n6224 , n6225 , n6226 , n6227 , n6228 , n6229 , n6230 , n6231 , n6232 , n6233 , n6234 , n6235 , n6236 , n6237 , n6238 , n6239 , n6240 , n6241 , n6242 , n6243 , n6244 , n6245 , n6246 , n6247 , n6248 , n6249 , n6250 , n6251 , n6252 , n6253 , n6254 , n6255 , n6256 , n6257 , n6258 , n6259 , n6260 , n6261 , n6262 , n6263 , n6264 , n6265 , n6266 , n6267 , n6268 , n6269 , n6270 , n6271 , n6272 , n6273 , n6274 , n6275 , n6276 , n6277 , n6278 , n6279 , n6280 , n6281 , n6282 , n6283 , n6284 , n6285 , n6286 , n6287 , n6288 , n6289 , n6290 , n6291 , n6292 , n6293 , n6294 , n6295 , n6296 , n6297 , n6298 , n6299 , n6300 , n6301 , n6302 , n6303 , n6304 , n6305 , n6306 , n6307 , n6308 , n6309 , n6310 , n6311 , n6312 , n6313 , n6314 , n6315 , n6316 , n6317 , n6318 , n6319 , n6320 , n6321 , n6322 , n6323 , n6324 , n6325 , n6326 , n6327 , n6328 , n6329 , n6330 , n6331 , n6332 , n6333 , n6334 , n6335 , n6336 , n6337 , n6338 , n6339 , n6340 , n6341 , n6342 , n6343 , n6344 , n6345 , n6346 , n6347 , n6348 , n6349 , n6350 , n6351 , n6352 , n6353 , n6354 , n6355 , n6356 , n6357 , n6358 , n6359 , n6360 , n6361 , n6362 , n6363 , n6364 , n6365 , n6366 , n6367 , n6368 , n6369 , n6370 , n6371 , n6372 , n6373 , n6374 , n6375 , n6376 , n6377 , n6378 , n6379 , n6380 , n6381 , n6382 , n6383 , n6384 , n6385 , n6386 , n6387 , n6388 , n6389 , n6390 , n6391 , n6392 , n6393 , n6394 , n6395 , n6396 , n6397 , n6398 , n6399 , n6400 , n6401 , n6402 , n6403 , n6404 , n6405 , n6406 , n6407 , n6408 , n6409 , n6410 , n6411 , n6412 , n6413 , n6414 , n6415 , n6416 , n6417 , n6418 , n6419 , n6420 , n6421 , n6422 , n6423 , n6424 , n6425 , n6426 , n6427 , n6428 , n6429 , n6430 , n6431 , n6432 , n6433 , n6434 , n6435 , n6436 , n6437 , n6438 , n6439 , n6440 , n6441 , n6442 , n6443 , n6444 , n6445 , n6446 , n6447 , n6448 , n6449 , n6450 , n6451 , n6452 , n6453 , n6454 , n6455 , n6456 , n6457 , n6458 , n6459 , n6460 , n6461 , n6462 , n6463 , n6464 , n6465 , n6466 , n6467 , n6468 , n6469 , n6470 , n6471 , n6472 , n6473 , n6474 , n6475 , n6476 , n6477 , n6478 , n6479 , n6480 , n6481 , n6482 , n6483 , n6484 , n6485 , n6486 , n6487 , n6488 , n6489 , n6490 , n6491 , n6492 , n6493 , n6494 , n6495 , n6496 , n6497 , n6498 , n6499 , n6500 , n6501 , n6502 , n6503 , n6504 , n6505 , n6506 , n6507 , n6508 , n6509 , n6510 , n6511 , n6512 , n6513 , n6514 , n6515 , n6516 , n6517 , n6518 , n6519 , n6520 , n6521 , n6522 , n6523 , n6524 , n6525 , n6526 , n6527 , n6528 , n6529 , n6530 , n6531 , n6532 , n6533 , n6534 , n6535 , n6536 , n6537 , n6538 , n6539 , n6540 , n6541 , n6542 , n6543 , n6544 , n6545 , n6546 , n6547 , n6548 , n6549 , n6550 , n6551 , n6552 , n6553 , n6554 , n6555 , n6556 , n6557 , n6558 , n6559 , n6560 , n6561 , n6562 , n6563 , n6564 , n6565 , n6566 , n6567 , n6568 , n6569 , n6570 , n6571 , n6572 , n6573 , n6574 , n6575 , n6576 , n6577 , n6578 , n6579 , n6580 , n6581 , n6582 , n6583 , n6584 , n6585 , n6586 , n6587 , n6588 , n6589 , n6590 , n6591 , n6592 , n6593 , n6594 , n6595 , n6596 , n6597 , n6598 , n6599 , n6600 , n6601 , n6602 , n6603 , n6604 , n6605 , n6606 , n6607 , n6608 , n6609 , n6610 , n6611 , n6612 , n6613 , n6614 , n6615 , n6616 , n6617 , n6618 , n6619 , n6620 , n6621 , n6622 , n6623 , n6624 , n6625 , n6626 , n6627 , n6628 , n6629 , n6630 , n6631 , n6632 , n6633 , n6634 , n6635 , n6636 , n6637 , n6638 , n6639 , n6640 , n6641 , n6642 , n6643 , n6644 , n6645 , n6646 , n6647 , n6648 , n6649 , n6650 , n6651 , n6652 , n6653 , n6654 , n6655 , n6656 , n6657 , n6658 , n6659 , n6660 , n6661 , n6662 , n6663 , n6664 , n6665 , n6666 , n6667 , n6668 , n6669 , n6670 , n6671 , n6672 , n6673 , n6674 , n6675 , n6676 , n6677 , n6678 , n6679 , n6680 , n6681 , n6682 , n6683 , n6684 , n6685 , n6686 , n6687 , n6688 , n6689 , n6690 , n6691 , n6692 , n6693 , n6694 , n6695 , n6696 , n6697 , n6698 , n6699 , n6700 , n6701 , n6702 , n6703 , n6704 , n6705 , n6706 , n6707 , n6708 , n6709 , n6710 , n6711 , n6712 , n6713 , n6714 , n6715 , n6716 , n6717 , n6718 , n6719 , n6720 , n6721 , n6722 , n6723 , n6724 , n6725 , n6726 , n6727 , n6728 , n6729 , n6730 , n6731 , n6732 , n6733 , n6734 , n6735 , n6736 , n6737 , n6738 , n6739 , n6740 , n6741 , n6742 , n6743 , n6744 , n6745 , n6746 , n6747 , n6748 , n6749 , n6750 , n6751 , n6752 , n6753 , n6754 , n6755 , n6756 , n6757 , n6758 , n6759 , n6760 , n6761 , n6762 , n6763 , n6764 , n6765 , n6766 , n6767 , n6768 , n6769 , n6770 , n6771 , n6772 , n6773 , n6774 , n6775 , n6776 , n6777 , n6778 , n6779 , n6780 , n6781 , n6782 , n6783 , n6784 , n6785 , n6786 , n6787 , n6788 , n6789 , n6790 , n6791 , n6792 , n6793 , n6794 , n6795 , n6796 , n6797 , n6798 , n6799 , n6800 , n6801 , n6802 , n6803 , n6804 , n6805 , n6806 , n6807 , n6808 , n6809 , n6810 , n6811 , n6812 , n6813 , n6814 , n6815 , n6816 , n6817 , n6818 , n6819 , n6820 , n6821 , n6822 , n6823 , n6824 , n6825 , n6826 , n6827 , n6828 , n6829 , n6830 , n6831 , n6832 , n6833 , n6834 , n6835 , n6836 , n6837 , n6838 , n6839 , n6840 , n6841 , n6842 , n6843 , n6844 , n6845 , n6846 , n6847 , n6848 , n6849 , n6850 , n6851 , n6852 , n6853 , n6854 , n6855 , n6856 , n6857 , n6858 , n6859 , n6860 , n6861 , n6862 , n6863 , n6864 , n6865 , n6866 , n6867 , n6868 , n6869 , n6870 , n6871 , n6872 , n6873 , n6874 , n6875 , n6876 , n6877 , n6878 , n6879 , n6880 , n6881 , n6882 , n6883 , n6884 , n6885 , n6886 , n6887 , n6888 , n6889 , n6890 , n6891 , n6892 , n6893 , n6894 , n6895 , n6896 , n6897 , n6898 , n6899 , n6900 , n6901 , n6902 , n6903 , n6904 , n6905 , n6906 , n6907 , n6908 , n6909 , n6910 , n6911 , n6912 , n6913 , n6914 , n6915 , n6916 , n6917 , n6918 , n6919 , n6920 , n6921 , n6922 , n6923 , n6924 , n6925 , n6926 , n6927 , n6928 , n6929 , n6930 , n6931 , n6932 , n6933 , n6934 , n6935 , n6936 , n6937 , n6938 , n6939 , n6940 , n6941 , n6942 , n6943 , n6944 , n6945 , n6946 , n6947 , n6948 , n6949 , n6950 , n6951 , n6952 , n6953 , n6954 , n6955 , n6956 , n6957 , n6958 , n6959 , n6960 , n6961 , n6962 , n6963 , n6964 , n6965 , n6966 , n6967 , n6968 , n6969 , n6970 , n6971 , n6972 , n6973 , n6974 , n6975 , n6976 , n6977 , n6978 , n6979 , n6980 , n6981 , n6982 , n6983 , n6984 , n6985 , n6986 , n6987 , n6988 , n6989 , n6990 , n6991 , n6992 , n6993 , n6994 , n6995 , n6996 , n6997 , n6998 , n6999 , n7000 , n7001 , n7002 , n7003 , n7004 , n7005 , n7006 , n7007 , n7008 , n7009 , n7010 , n7011 , n7012 , n7013 , n7014 , n7015 , n7016 , n7017 , n7018 , n7019 , n7020 , n7021 , n7022 , n7023 , n7024 , n7025 , n7026 , n7027 , n7028 , n7029 , n7030 , n7031 , n7032 , n7033 , n7034 , n7035 , n7036 , n7037 , n7038 , n7039 , n7040 , n7041 , n7042 , n7043 , n7044 , n7045 , n7046 , n7047 , n7048 , n7049 , n7050 , n7051 , n7052 , n7053 , n7054 , n7055 , n7056 , n7057 , n7058 , n7059 , n7060 , n7061 , n7062 , n7063 , n7064 , n7065 , n7066 , n7067 , n7068 , n7069 , n7070 , n7071 , n7072 , n7073 , n7074 , n7075 , n7076 , n7077 , n7078 , n7079 , n7080 , n7081 , n7082 , n7083 , n7084 , n7085 , n7086 , n7087 , n7088 , n7089 , n7090 , n7091 , n7092 , n7093 , n7094 , n7095 , n7096 , n7097 , n7098 , n7099 , n7100 , n7101 , n7102 , n7103 , n7104 , n7105 , n7106 , n7107 , n7108 , n7109 , n7110 , n7111 , n7112 , n7113 , n7114 , n7115 , n7116 , n7117 , n7118 , n7119 , n7120 , n7121 , n7122 , n7123 , n7124 , n7125 , n7126 , n7127 , n7128 , n7129 , n7130 , n7131 , n7132 , n7133 , n7134 , n7135 , n7136 , n7137 , n7138 , n7139 , n7140 , n7141 , n7142 , n7143 , n7144 , n7145 , n7146 , n7147 , n7148 , n7149 , n7150 , n7151 , n7152 , n7153 , n7154 , n7155 , n7156 , n7157 , n7158 , n7159 , n7160 , n7161 , n7162 , n7163 , n7164 , n7165 , n7166 , n7167 , n7168 , n7169 , n7170 , n7171 , n7172 , n7173 , n7174 , n7175 , n7176 , n7177 , n7178 , n7179 , n7180 , n7181 , n7182 , n7183 , n7184 , n7185 , n7186 , n7187 , n7188 , n7189 , n7190 , n7191 , n7192 , n7193 , n7194 , n7195 , n7196 , n7197 , n7198 , n7199 , n7200 , n7201 , n7202 , n7203 , n7204 , n7205 , n7206 , n7207 , n7208 , n7209 , n7210 , n7211 , n7212 , n7213 , n7214 , n7215 , n7216 , n7217 , n7218 , n7219 , n7220 , n7221 , n7222 , n7223 , n7224 , n7225 , n7226 , n7227 , n7228 , n7229 , n7230 , n7231 , n7232 , n7233 , n7234 , n7235 , n7236 , n7237 , n7238 , n7239 , n7240 , n7241 , n7242 , n7243 , n7244 , n7245 , n7246 , n7247 , n7248 , n7249 , n7250 , n7251 , n7252 , n7253 , n7254 , n7255 , n7256 , n7257 , n7258 , n7259 , n7260 , n7261 , n7262 , n7263 , n7264 , n7265 , n7266 , n7267 , n7268 , n7269 , n7270 , n7271 , n7272 , n7273 , n7274 , n7275 , n7276 , n7277 , n7278 , n7279 , n7280 , n7281 , n7282 , n7283 , n7284 , n7285 , n7286 , n7287 , n7288 , n7289 , n7290 , n7291 , n7292 , n7293 , n7294 , n7295 , n7296 , n7297 , n7298 , n7299 , n7300 , n7301 , n7302 , n7303 , n7304 , n7305 , n7306 , n7307 , n7308 , n7309 , n7310 , n7311 , n7312 , n7313 , n7314 , n7315 , n7316 , n7317 , n7318 , n7319 , n7320 , n7321 , n7322 , n7323 , n7324 , n7325 , n7326 , n7327 , n7328 , n7329 , n7330 , n7331 , n7332 , n7333 , n7334 , n7335 , n7336 , n7337 , n7338 , n7339 , n7340 , n7341 , n7342 , n7343 , n7344 , n7345 , n7346 , n7347 , n7348 , n7349 , n7350 , n7351 , n7352 , n7353 , n7354 , n7355 , n7356 , n7357 , n7358 , n7359 , n7360 , n7361 , n7362 , n7363 , n7364 , n7365 , n7366 , n7367 , n7368 , n7369 , n7370 , n7371 , n7372 , n7373 , n7374 , n7375 , n7376 , n7377 , n7378 , n7379 , n7380 , n7381 , n7382 , n7383 , n7384 , n7385 , n7386 , n7387 , n7388 , n7389 , n7390 , n7391 , n7392 , n7393 , n7394 , n7395 , n7396 , n7397 , n7398 , n7399 , n7400 , n7401 , n7402 , n7403 , n7404 , n7405 , n7406 , n7407 , n7408 , n7409 , n7410 , n7411 , n7412 , n7413 , n7414 , n7415 , n7416 , n7417 , n7418 , n7419 , n7420 , n7421 , n7422 , n7423 , n7424 , n7425 , n7426 , n7427 , n7428 , n7429 , n7430 , n7431 , n7432 , n7433 , n7434 , n7435 , n7436 , n7437 , n7438 , n7439 , n7440 , n7441 , n7442 , n7443 , n7444 , n7445 , n7446 , n7447 , n7448 , n7449 , n7450 , n7451 , n7452 , n7453 , n7454 , n7455 , n7456 , n7457 , n7458 , n7459 , n7460 , n7461 , n7462 , n7463 , n7464 , n7465 , n7466 , n7467 , n7468 , n7469 , n7470 , n7471 , n7472 , n7473 , n7474 , n7475 , n7476 , n7477 , n7478 , n7479 , n7480 , n7481 , n7482 , n7483 , n7484 , n7485 , n7486 , n7487 , n7488 , n7489 , n7490 , n7491 , n7492 , n7493 , n7494 , n7495 , n7496 , n7497 , n7498 , n7499 , n7500 , n7501 , n7502 , n7503 , n7504 , n7505 , n7506 , n7507 , n7508 , n7509 , n7510 , n7511 , n7512 , n7513 , n7514 , n7515 , n7516 , n7517 , n7518 , n7519 , n7520 , n7521 , n7522 , n7523 , n7524 , n7525 , n7526 , n7527 , n7528 , n7529 , n7530 , n7531 , n7532 , n7533 , n7534 , n7535 , n7536 , n7537 , n7538 , n7539 , n7540 , n7541 , n7542 , n7543 , n7544 , n7545 , n7546 , n7547 , n7548 , n7549 , n7550 , n7551 , n7552 , n7553 , n7554 , n7555 , n7556 , n7557 , n7558 , n7559 , n7560 , n7561 , n7562 , n7563 , n7564 , n7565 , n7566 , n7567 , n7568 , n7569 , n7570 , n7571 , n7572 , n7573 , n7574 , n7575 , n7576 , n7577 , n7578 , n7579 , n7580 , n7581 , n7582 , n7583 , n7584 , n7585 , n7586 , n7587 , n7588 , n7589 , n7590 , n7591 , n7592 , n7593 , n7594 , n7595 , n7596 , n7597 , n7598 , n7599 , n7600 , n7601 , n7602 , n7603 , n7604 , n7605 , n7606 , n7607 , n7608 , n7609 , n7610 , n7611 , n7612 , n7613 , n7614 , n7615 , n7616 , n7617 , n7618 , n7619 , n7620 , n7621 , n7622 , n7623 , n7624 , n7625 , n7626 , n7627 , n7628 , n7629 , n7630 , n7631 , n7632 , n7633 , n7634 , n7635 , n7636 , n7637 , n7638 , n7639 , n7640 , n7641 , n7642 , n7643 , n7644 , n7645 , n7646 , n7647 , n7648 , n7649 , n7650 , n7651 , n7652 , n7653 , n7654 , n7655 , n7656 , n7657 , n7658 , n7659 , n7660 , n7661 , n7662 , n7663 , n7664 , n7665 , n7666 , n7667 , n7668 , n7669 , n7670 , n7671 , n7672 , n7673 , n7674 , n7675 , n7676 , n7677 , n7678 , n7679 , n7680 , n7681 , n7682 , n7683 , n7684 , n7685 , n7686 , n7687 , n7688 , n7689 , n7690 , n7691 , n7692 , n7693 , n7694 , n7695 , n7696 , n7697 , n7698 , n7699 , n7700 , n7701 , n7702 , n7703 , n7704 , n7705 , n7706 , n7707 , n7708 , n7709 , n7710 , n7711 , n7712 , n7713 , n7714 , n7715 , n7716 , n7717 , n7718 , n7719 , n7720 , n7721 , n7722 , n7723 , n7724 , n7725 , n7726 , n7727 , n7728 , n7729 , n7730 , n7731 , n7732 , n7733 , n7734 , n7735 , n7736 , n7737 , n7738 , n7739 , n7740 , n7741 , n7742 , n7743 , n7744 , n7745 , n7746 , n7747 , n7748 , n7749 , n7750 , n7751 , n7752 , n7753 , n7754 , n7755 , n7756 , n7757 , n7758 , n7759 , n7760 , n7761 , n7762 , n7763 , n7764 , n7765 , n7766 , n7767 , n7768 , n7769 , n7770 , n7771 , n7772 , n7773 , n7774 , n7775 , n7776 , n7777 , n7778 , n7779 , n7780 , n7781 , n7782 , n7783 , n7784 , n7785 , n7786 , n7787 , n7788 , n7789 , n7790 , n7791 , n7792 , n7793 , n7794 , n7795 , n7796 , n7797 , n7798 , n7799 , n7800 , n7801 , n7802 , n7803 , n7804 , n7805 , n7806 , n7807 , n7808 , n7809 , n7810 , n7811 , n7812 , n7813 , n7814 , n7815 , n7816 , n7817 , n7818 , n7819 , n7820 , n7821 , n7822 , n7823 , n7824 , n7825 , n7826 , n7827 , n7828 , n7829 , n7830 , n7831 , n7832 , n7833 , n7834 , n7835 , n7836 , n7837 , n7838 , n7839 , n7840 , n7841 , n7842 , n7843 , n7844 , n7845 , n7846 , n7847 , n7848 , n7849 , n7850 , n7851 , n7852 , n7853 , n7854 , n7855 , n7856 , n7857 , n7858 , n7859 , n7860 , n7861 , n7862 , n7863 , n7864 , n7865 , n7866 , n7867 , n7868 , n7869 , n7870 , n7871 , n7872 , n7873 , n7874 , n7875 , n7876 , n7877 , n7878 , n7879 , n7880 , n7881 , n7882 , n7883 , n7884 , n7885 , n7886 , n7887 , n7888 , n7889 , n7890 , n7891 , n7892 , n7893 , n7894 , n7895 , n7896 , n7897 , n7898 , n7899 , n7900 , n7901 , n7902 , n7903 , n7904 , n7905 , n7906 , n7907 , n7908 , n7909 , n7910 , n7911 , n7912 , n7913 , n7914 , n7915 , n7916 , n7917 , n7918 , n7919 , n7920 , n7921 , n7922 , n7923 , n7924 , n7925 , n7926 , n7927 , n7928 , n7929 , n7930 , n7931 , n7932 , n7933 , n7934 , n7935 , n7936 , n7937 , n7938 , n7939 , n7940 , n7941 , n7942 , n7943 , n7944 , n7945 , n7946 , n7947 , n7948 , n7949 , n7950 , n7951 , n7952 , n7953 , n7954 , n7955 , n7956 , n7957 , n7958 , n7959 , n7960 , n7961 , n7962 , n7963 , n7964 , n7965 , n7966 , n7967 , n7968 , n7969 , n7970 , n7971 , n7972 , n7973 , n7974 , n7975 , n7976 , n7977 , n7978 , n7979 , n7980 , n7981 , n7982 , n7983 , n7984 , n7985 , n7986 , n7987 , n7988 , n7989 , n7990 , n7991 , n7992 , n7993 , n7994 , n7995 , n7996 , n7997 , n7998 , n7999 , n8000 , n8001 , n8002 , n8003 , n8004 , n8005 , n8006 , n8007 , n8008 , n8009 , n8010 , n8011 , n8012 , n8013 , n8014 , n8015 , n8016 , n8017 , n8018 , n8019 , n8020 , n8021 , n8022 , n8023 , n8024 , n8025 , n8026 , n8027 , n8028 , n8029 , n8030 , n8031 , n8032 , n8033 , n8034 , n8035 , n8036 , n8037 , n8038 , n8039 , n8040 , n8041 , n8042 , n8043 , n8044 , n8045 , n8046 , n8047 , n8048 , n8049 , n8050 , n8051 , n8052 , n8053 , n8054 , n8055 , n8056 , n8057 , n8058 , n8059 , n8060 , n8061 , n8062 , n8063 , n8064 , n8065 , n8066 , n8067 , n8068 , n8069 , n8070 , n8071 , n8072 , n8073 , n8074 , n8075 , n8076 , n8077 , n8078 , n8079 , n8080 , n8081 , n8082 , n8083 , n8084 , n8085 , n8086 , n8087 , n8088 , n8089 , n8090 , n8091 , n8092 , n8093 , n8094 , n8095 , n8096 , n8097 , n8098 , n8099 , n8100 , n8101 , n8102 , n8103 , n8104 , n8105 , n8106 , n8107 , n8108 , n8109 , n8110 , n8111 , n8112 , n8113 , n8114 , n8115 , n8116 , n8117 , n8118 , n8119 , n8120 , n8121 , n8122 , n8123 , n8124 , n8125 , n8126 , n8127 , n8128 , n8129 , n8130 , n8131 , n8132 , n8133 , n8134 , n8135 , n8136 , n8137 , n8138 , n8139 , n8140 , n8141 , n8142 , n8143 , n8144 , n8145 , n8146 , n8147 , n8148 , n8149 , n8150 , n8151 , n8152 , n8153 , n8154 , n8155 , n8156 , n8157 , n8158 , n8159 , n8160 , n8161 , n8162 , n8163 , n8164 , n8165 , n8166 , n8167 , n8168 , n8169 , n8170 , n8171 , n8172 , n8173 , n8174 , n8175 , n8176 , n8177 , n8178 , n8179 , n8180 , n8181 , n8182 , n8183 , n8184 , n8185 , n8186 , n8187 , n8188 , n8189 , n8190 , n8191 , n8192 , n8193 , n8194 , n8195 , n8196 , n8197 , n8198 , n8199 , n8200 , n8201 , n8202 , n8203 , n8204 , n8205 , n8206 , n8207 , n8208 , n8209 , n8210 , n8211 , n8212 , n8213 , n8214 , n8215 , n8216 , n8217 , n8218 , n8219 , n8220 , n8221 , n8222 , n8223 , n8224 , n8225 , n8226 , n8227 , n8228 , n8229 , n8230 , n8231 , n8232 , n8233 , n8234 , n8235 , n8236 , n8237 , n8238 , n8239 , n8240 , n8241 , n8242 , n8243 , n8244 , n8245 , n8246 , n8247 , n8248 , n8249 , n8250 , n8251 , n8252 , n8253 , n8254 , n8255 , n8256 , n8257 , n8258 , n8259 , n8260 , n8261 , n8262 , n8263 , n8264 , n8265 , n8266 , n8267 , n8268 , n8269 , n8270 , n8271 , n8272 , n8273 , n8274 , n8275 , n8276 , n8277 , n8278 , n8279 , n8280 , n8281 , n8282 , n8283 , n8284 , n8285 , n8286 , n8287 , n8288 , n8289 , n8290 , n8291 , n8292 , n8293 , n8294 , n8295 , n8296 , n8297 , n8298 , n8299 , n8300 , n8301 , n8302 , n8303 , n8304 , n8305 , n8306 , n8307 , n8308 , n8309 , n8310 , n8311 , n8312 , n8313 , n8314 , n8315 , n8316 , n8317 , n8318 , n8319 , n8320 , n8321 , n8322 , n8323 , n8324 , n8325 , n8326 , n8327 , n8328 , n8329 , n8330 , n8331 , n8332 , n8333 , n8334 , n8335 , n8336 , n8337 , n8338 , n8339 , n8340 , n8341 , n8342 , n8343 , n8344 , n8345 , n8346 , n8347 , n8348 , n8349 , n8350 , n8351 , n8352 , n8353 , n8354 , n8355 , n8356 , n8357 , n8358 , n8359 , n8360 , n8361 , n8362 , n8363 , n8364 , n8365 , n8366 , n8367 , n8368 , n8369 , n8370 , n8371 , n8372 , n8373 , n8374 , n8375 , n8376 , n8377 , n8378 , n8379 , n8380 , n8381 , n8382 , n8383 , n8384 , n8385 , n8386 , n8387 , n8388 , n8389 , n8390 , n8391 , n8392 , n8393 , n8394 , n8395 , n8396 , n8397 , n8398 , n8399 , n8400 , n8401 , n8402 , n8403 , n8404 , n8405 , n8406 , n8407 , n8408 , n8409 , n8410 , n8411 , n8412 , n8413 , n8414 , n8415 , n8416 , n8417 , n8418 , n8419 , n8420 , n8421 , n8422 , n8423 , n8424 , n8425 , n8426 , n8427 , n8428 , n8429 , n8430 , n8431 , n8432 , n8433 , n8434 , n8435 , n8436 , n8437 , n8438 , n8439 , n8440 , n8441 , n8442 , n8443 , n8444 , n8445 , n8446 , n8447 , n8448 , n8449 , n8450 , n8451 , n8452 , n8453 , n8454 , n8455 , n8456 , n8457 , n8458 , n8459 , n8460 , n8461 , n8462 , n8463 , n8464 , n8465 , n8466 , n8467 , n8468 , n8469 , n8470 , n8471 , n8472 , n8473 , n8474 , n8475 , n8476 , n8477 , n8478 , n8479 , n8480 , n8481 , n8482 , n8483 , n8484 , n8485 , n8486 , n8487 , n8488 , n8489 , n8490 , n8491 , n8492 , n8493 , n8494 , n8495 , n8496 , n8497 , n8498 , n8499 , n8500 , n8501 , n8502 , n8503 , n8504 , n8505 , n8506 , n8507 , n8508 , n8509 , n8510 , n8511 , n8512 , n8513 , n8514 , n8515 , n8516 , n8517 , n8518 , n8519 , n8520 , n8521 , n8522 , n8523 , n8524 , n8525 , n8526 , n8527 , n8528 , n8529 , n8530 , n8531 , n8532 , n8533 , n8534 , n8535 , n8536 , n8537 , n8538 , n8539 , n8540 , n8541 , n8542 , n8543 , n8544 , n8545 , n8546 , n8547 , n8548 , n8549 , n8550 , n8551 , n8552 , n8553 , n8554 , n8555 , n8556 , n8557 , n8558 , n8559 , n8560 , n8561 , n8562 , n8563 , n8564 , n8565 , n8566 , n8567 , n8568 , n8569 , n8570 , n8571 , n8572 , n8573 , n8574 , n8575 , n8576 , n8577 , n8578 , n8579 , n8580 , n8581 , n8582 , n8583 , n8584 , n8585 , n8586 , n8587 , n8588 , n8589 , n8590 , n8591 , n8592 , n8593 , n8594 , n8595 , n8596 , n8597 , n8598 , n8599 , n8600 , n8601 , n8602 , n8603 , n8604 , n8605 , n8606 , n8607 , n8608 , n8609 , n8610 , n8611 , n8612 , n8613 , n8614 , n8615 , n8616 , n8617 , n8618 , n8619 , n8620 , n8621 , n8622 , n8623 , n8624 , n8625 , n8626 , n8627 , n8628 , n8629 , n8630 , n8631 , n8632 , n8633 , n8634 , n8635 , n8636 , n8637 , n8638 , n8639 , n8640 , n8641 , n8642 , n8643 , n8644 , n8645 , n8646 , n8647 , n8648 , n8649 , n8650 , n8651 , n8652 , n8653 , n8654 , n8655 , n8656 , n8657 , n8658 , n8659 , n8660 , n8661 , n8662 , n8663 , n8664 , n8665 , n8666 , n8667 , n8668 , n8669 , n8670 , n8671 , n8672 , n8673 , n8674 , n8675 , n8676 , n8677 , n8678 , n8679 , n8680 , n8681 , n8682 , n8683 , n8684 , n8685 , n8686 , n8687 , n8688 , n8689 , n8690 , n8691 , n8692 , n8693 , n8694 , n8695 , n8696 , n8697 , n8698 , n8699 , n8700 , n8701 , n8702 , n8703 , n8704 , n8705 , n8706 , n8707 , n8708 , n8709 , n8710 , n8711 , n8712 , n8713 , n8714 , n8715 , n8716 , n8717 , n8718 , n8719 , n8720 , n8721 , n8722 , n8723 , n8724 , n8725 , n8726 , n8727 , n8728 , n8729 , n8730 , n8731 , n8732 , n8733 , n8734 , n8735 , n8736 , n8737 , n8738 , n8739 , n8740 , n8741 , n8742 , n8743 , n8744 , n8745 , n8746 , n8747 , n8748 , n8749 , n8750 , n8751 , n8752 , n8753 , n8754 , n8755 , n8756 , n8757 , n8758 , n8759 , n8760 , n8761 , n8762 , n8763 , n8764 , n8765 , n8766 , n8767 , n8768 , n8769 , n8770 , n8771 , n8772 , n8773 , n8774 , n8775 , n8776 , n8777 , n8778 , n8779 , n8780 , n8781 , n8782 , n8783 , n8784 , n8785 , n8786 , n8787 , n8788 , n8789 , n8790 , n8791 , n8792 , n8793 , n8794 , n8795 , n8796 , n8797 , n8798 , n8799 , n8800 , n8801 , n8802 , n8803 , n8804 , n8805 , n8806 , n8807 , n8808 , n8809 , n8810 , n8811 , n8812 , n8813 , n8814 , n8815 , n8816 , n8817 , n8818 , n8819 , n8820 , n8821 , n8822 , n8823 , n8824 , n8825 , n8826 , n8827 , n8828 , n8829 , n8830 , n8831 , n8832 , n8833 , n8834 , n8835 , n8836 , n8837 , n8838 , n8839 , n8840 , n8841 , n8842 , n8843 , n8844 , n8845 , n8846 , n8847 , n8848 , n8849 , n8850 , n8851 , n8852 , n8853 , n8854 , n8855 , n8856 , n8857 , n8858 , n8859 , n8860 , n8861 , n8862 , n8863 , n8864 , n8865 , n8866 , n8867 , n8868 , n8869 , n8870 , n8871 , n8872 , n8873 , n8874 , n8875 , n8876 , n8877 , n8878 , n8879 , n8880 , n8881 , n8882 , n8883 , n8884 , n8885 , n8886 , n8887 , n8888 , n8889 , n8890 , n8891 , n8892 , n8893 , n8894 , n8895 , n8896 , n8897 , n8898 , n8899 , n8900 , n8901 , n8902 , n8903 , n8904 , n8905 , n8906 , n8907 , n8908 , n8909 , n8910 , n8911 , n8912 , n8913 , n8914 , n8915 , n8916 , n8917 , n8918 , n8919 , n8920 , n8921 , n8922 , n8923 , n8924 , n8925 , n8926 , n8927 , n8928 , n8929 , n8930 , n8931 , n8932 , n8933 , n8934 , n8935 , n8936 , n8937 , n8938 , n8939 , n8940 , n8941 , n8942 , n8943 , n8944 , n8945 , n8946 , n8947 , n8948 , n8949 , n8950 , n8951 , n8952 , n8953 , n8954 , n8955 , n8956 , n8957 , n8958 , n8959 , n8960 , n8961 , n8962 , n8963 , n8964 , n8965 , n8966 , n8967 , n8968 , n8969 , n8970 , n8971 , n8972 , n8973 , n8974 , n8975 , n8976 , n8977 , n8978 , n8979 , n8980 , n8981 , n8982 , n8983 , n8984 , n8985 , n8986 , n8987 , n8988 , n8989 , n8990 , n8991 , n8992 , n8993 , n8994 , n8995 , n8996 , n8997 , n8998 , n8999 , n9000 , n9001 , n9002 , n9003 , n9004 , n9005 , n9006 , n9007 , n9008 , n9009 , n9010 , n9011 , n9012 , n9013 , n9014 , n9015 , n9016 , n9017 , n9018 , n9019 , n9020 , n9021 , n9022 , n9023 , n9024 , n9025 , n9026 , n9027 , n9028 , n9029 , n9030 , n9031 , n9032 , n9033 , n9034 , n9035 , n9036 , n9037 , n9038 , n9039 , n9040 , n9041 , n9042 , n9043 , n9044 , n9045 , n9046 , n9047 , n9048 , n9049 , n9050 , n9051 , n9052 , n9053 , n9054 , n9055 , n9056 , n9057 , n9058 , n9059 , n9060 , n9061 , n9062 , n9063 , n9064 , n9065 , n9066 , n9067 , n9068 , n9069 , n9070 , n9071 , n9072 , n9073 , n9074 , n9075 , n9076 , n9077 , n9078 , n9079 , n9080 , n9081 , n9082 , n9083 , n9084 , n9085 , n9086 , n9087 , n9088 , n9089 , n9090 , n9091 , n9092 , n9093 , n9094 , n9095 , n9096 , n9097 , n9098 , n9099 , n9100 , n9101 , n9102 , n9103 , n9104 , n9105 , n9106 , n9107 , n9108 , n9109 , n9110 , n9111 , n9112 , n9113 , n9114 , n9115 , n9116 , n9117 , n9118 , n9119 , n9120 , n9121 , n9122 , n9123 , n9124 , n9125 , n9126 , n9127 , n9128 , n9129 , n9130 , n9131 , n9132 , n9133 , n9134 , n9135 , n9136 , n9137 , n9138 , n9139 , n9140 , n9141 , n9142 , n9143 , n9144 , n9145 , n9146 , n9147 , n9148 , n9149 , n9150 , n9151 , n9152 , n9153 , n9154 , n9155 , n9156 , n9157 , n9158 , n9159 , n9160 , n9161 , n9162 , n9163 , n9164 , n9165 , n9166 , n9167 , n9168 , n9169 , n9170 , n9171 , n9172 , n9173 , n9174 , n9175 , n9176 , n9177 , n9178 , n9179 , n9180 , n9181 , n9182 , n9183 , n9184 , n9185 , n9186 , n9187 , n9188 , n9189 , n9190 , n9191 , n9192 , n9193 , n9194 , n9195 , n9196 , n9197 , n9198 , n9199 , n9200 , n9201 , n9202 , n9203 , n9204 , n9205 , n9206 , n9207 , n9208 , n9209 , n9210 , n9211 , n9212 , n9213 , n9214 , n9215 , n9216 , n9217 , n9218 , n9219 , n9220 , n9221 , n9222 , n9223 , n9224 , n9225 , n9226 , n9227 , n9228 , n9229 , n9230 , n9231 , n9232 , n9233 , n9234 , n9235 , n9236 , n9237 , n9238 , n9239 , n9240 , n9241 , n9242 , n9243 , n9244 , n9245 , n9246 , n9247 , n9248 , n9249 , n9250 , n9251 , n9252 , n9253 , n9254 , n9255 , n9256 , n9257 , n9258 , n9259 , n9260 , n9261 , n9262 , n9263 , n9264 , n9265 , n9266 , n9267 , n9268 , n9269 , n9270 , n9271 , n9272 , n9273 , n9274 , n9275 , n9276 , n9277 , n9278 , n9279 , n9280 , n9281 , n9282 , n9283 , n9284 , n9285 , n9286 , n9287 , n9288 , n9289 , n9290 , n9291 , n9292 , n9293 , n9294 , n9295 , n9296 , n9297 , n9298 , n9299 , n9300 , n9301 , n9302 , n9303 , n9304 , n9305 , n9306 , n9307 , n9308 , n9309 , n9310 , n9311 , n9312 , n9313 , n9314 , n9315 , n9316 , n9317 , n9318 , n9319 , n9320 , n9321 , n9322 , n9323 , n9324 , n9325 , n9326 , n9327 , n9328 , n9329 , n9330 , n9331 , n9332 , n9333 , n9334 , n9335 , n9336 , n9337 , n9338 , n9339 , n9340 , n9341 , n9342 , n9343 , n9344 , n9345 , n9346 , n9347 , n9348 , n9349 , n9350 , n9351 , n9352 , n9353 , n9354 , n9355 , n9356 , n9357 , n9358 , n9359 , n9360 , n9361 , n9362 , n9363 , n9364 , n9365 , n9366 , n9367 , n9368 , n9369 , n9370 , n9371 , n9372 , n9373 , n9374 , n9375 , n9376 , n9377 , n9378 , n9379 , n9380 , n9381 , n9382 , n9383 , n9384 , n9385 , n9386 , n9387 , n9388 , n9389 , n9390 , n9391 , n9392 , n9393 , n9394 , n9395 , n9396 , n9397 , n9398 , n9399 , n9400 , n9401 , n9402 , n9403 , n9404 , n9405 , n9406 , n9407 , n9408 , n9409 , n9410 , n9411 , n9412 , n9413 , n9414 , n9415 , n9416 , n9417 , n9418 , n9419 , n9420 , n9421 , n9422 , n9423 , n9424 , n9425 , n9426 , n9427 , n9428 , n9429 , n9430 , n9431 , n9432 , n9433 , n9434 , n9435 , n9436 , n9437 , n9438 , n9439 , n9440 , n9441 , n9442 , n9443 , n9444 , n9445 , n9446 , n9447 , n9448 , n9449 , n9450 , n9451 , n9452 , n9453 , n9454 , n9455 , n9456 , n9457 , n9458 , n9459 , n9460 , n9461 , n9462 , n9463 , n9464 , n9465 , n9466 , n9467 , n9468 , n9469 , n9470 , n9471 , n9472 , n9473 , n9474 , n9475 , n9476 , n9477 , n9478 , n9479 , n9480 , n9481 , n9482 , n9483 , n9484 , n9485 , n9486 , n9487 , n9488 , n9489 , n9490 , n9491 , n9492 , n9493 , n9494 , n9495 , n9496 , n9497 , n9498 , n9499 , n9500 , n9501 , n9502 , n9503 , n9504 , n9505 , n9506 , n9507 , n9508 , n9509 , n9510 , n9511 , n9512 , n9513 , n9514 , n9515 , n9516 , n9517 , n9518 , n9519 , n9520 , n9521 , n9522 , n9523 , n9524 , n9525 , n9526 , n9527 , n9528 , n9529 , n9530 , n9531 , n9532 , n9533 , n9534 , n9535 , n9536 , n9537 , n9538 , n9539 , n9540 , n9541 , n9542 , n9543 , n9544 , n9545 , n9546 , n9547 , n9548 , n9549 , n9550 , n9551 , n9552 , n9553 , n9554 , n9555 , n9556 , n9557 , n9558 , n9559 , n9560 , n9561 , n9562 , n9563 , n9564 , n9565 , n9566 , n9567 , n9568 , n9569 , n9570 , n9571 , n9572 , n9573 , n9574 , n9575 , n9576 , n9577 , n9578 , n9579 , n9580 , n9581 , n9582 , n9583 , n9584 , n9585 , n9586 , n9587 , n9588 , n9589 , n9590 , n9591 , n9592 , n9593 , n9594 , n9595 , n9596 , n9597 , n9598 , n9599 , n9600 , n9601 , n9602 , n9603 , n9604 , n9605 , n9606 , n9607 , n9608 , n9609 , n9610 , n9611 , n9612 , n9613 , n9614 , n9615 , n9616 , n9617 , n9618 , n9619 , n9620 , n9621 , n9622 , n9623 , n9624 , n9625 , n9626 , n9627 , n9628 , n9629 , n9630 , n9631 , n9632 , n9633 , n9634 , n9635 , n9636 , n9637 , n9638 , n9639 , n9640 , n9641 , n9642 , n9643 , n9644 , n9645 , n9646 , n9647 , n9648 , n9649 , n9650 , n9651 , n9652 , n9653 , n9654 , n9655 , n9656 , n9657 , n9658 , n9659 , n9660 , n9661 , n9662 , n9663 , n9664 , n9665 , n9666 , n9667 , n9668 , n9669 , n9670 , n9671 , n9672 , n9673 , n9674 , n9675 , n9676 , n9677 , n9678 , n9679 , n9680 , n9681 , n9682 , n9683 , n9684 , n9685 , n9686 , n9687 , n9688 , n9689 , n9690 , n9691 , n9692 , n9693 , n9694 , n9695 , n9696 , n9697 , n9698 , n9699 , n9700 , n9701 , n9702 , n9703 , n9704 , n9705 , n9706 , n9707 , n9708 , n9709 , n9710 , n9711 , n9712 , n9713 , n9714 , n9715 , n9716 , n9717 , n9718 , n9719 , n9720 , n9721 , n9722 , n9723 , n9724 , n9725 , n9726 , n9727 , n9728 , n9729 , n9730 , n9731 , n9732 , n9733 , n9734 , n9735 , n9736 , n9737 , n9738 , n9739 , n9740 , n9741 , n9742 , n9743 , n9744 , n9745 , n9746 , n9747 , n9748 , n9749 , n9750 , n9751 , n9752 , n9753 , n9754 , n9755 , n9756 , n9757 , n9758 , n9759 , n9760 , n9761 , n9762 , n9763 , n9764 , n9765 , n9766 , n9767 , n9768 , n9769 , n9770 , n9771 , n9772 , n9773 , n9774 , n9775 , n9776 , n9777 , n9778 , n9779 , n9780 , n9781 , n9782 , n9783 , n9784 , n9785 , n9786 , n9787 , n9788 , n9789 , n9790 , n9791 , n9792 , n9793 , n9794 , n9795 , n9796 , n9797 , n9798 , n9799 , n9800 , n9801 , n9802 , n9803 , n9804 , n9805 , n9806 , n9807 , n9808 , n9809 , n9810 , n9811 , n9812 , n9813 , n9814 , n9815 , n9816 , n9817 , n9818 , n9819 , n9820 , n9821 , n9822 , n9823 , n9824 , n9825 , n9826 , n9827 , n9828 , n9829 , n9830 , n9831 , n9832 , n9833 , n9834 , n9835 , n9836 , n9837 , n9838 , n9839 , n9840 , n9841 , n9842 , n9843 , n9844 , n9845 , n9846 , n9847 , n9848 , n9849 , n9850 , n9851 , n9852 , n9853 , n9854 , n9855 , n9856 , n9857 , n9858 , n9859 , n9860 , n9861 , n9862 , n9863 , n9864 , n9865 , n9866 , n9867 , n9868 , n9869 , n9870 , n9871 , n9872 , n9873 , n9874 , n9875 , n9876 , n9877 , n9878 , n9879 , n9880 , n9881 , n9882 , n9883 , n9884 , n9885 , n9886 , n9887 , n9888 , n9889 , n9890 , n9891 , n9892 , n9893 , n9894 , n9895 , n9896 , n9897 , n9898 , n9899 , n9900 , n9901 , n9902 , n9903 , n9904 , n9905 , n9906 , n9907 , n9908 , n9909 , n9910 , n9911 , n9912 , n9913 , n9914 , n9915 , n9916 , n9917 , n9918 , n9919 , n9920 , n9921 , n9922 , n9923 , n9924 , n9925 , n9926 , n9927 , n9928 , n9929 , n9930 , n9931 , n9932 , n9933 , n9934 , n9935 , n9936 , n9937 , n9938 , n9939 , n9940 , n9941 , n9942 , n9943 , n9944 , n9945 , n9946 , n9947 , n9948 , n9949 , n9950 , n9951 , n9952 , n9953 , n9954 , n9955 , n9956 , n9957 , n9958 , n9959 , n9960 , n9961 , n9962 , n9963 , n9964 , n9965 , n9966 , n9967 , n9968 , n9969 , n9970 , n9971 , n9972 , n9973 , n9974 , n9975 , n9976 , n9977 , n9978 , n9979 , n9980 , n9981 , n9982 , n9983 , n9984 , n9985 , n9986 , n9987 , n9988 , n9989 , n9990 , n9991 , n9992 , n9993 , n9994 , n9995 , n9996 , n9997 , n9998 , n9999 , n10000 , n10001 , n10002 , n10003 , n10004 , n10005 , n10006 , n10007 , n10008 , n10009 , n10010 , n10011 , n10012 , n10013 , n10014 , n10015 , n10016 , n10017 , n10018 , n10019 , n10020 , n10021 , n10022 , n10023 , n10024 , n10025 , n10026 , n10027 , n10028 , n10029 , n10030 , n10031 , n10032 , n10033 , n10034 , n10035 , n10036 , n10037 , n10038 , n10039 , n10040 , n10041 , n10042 , n10043 , n10044 , n10045 , n10046 , n10047 , n10048 , n10049 , n10050 , n10051 , n10052 , n10053 , n10054 , n10055 , n10056 , n10057 , n10058 , n10059 , n10060 , n10061 , n10062 , n10063 , n10064 , n10065 , n10066 , n10067 , n10068 , n10069 , n10070 , n10071 , n10072 , n10073 , n10074 , n10075 , n10076 , n10077 , n10078 , n10079 , n10080 , n10081 , n10082 , n10083 , n10084 , n10085 , n10086 , n10087 , n10088 , n10089 , n10090 , n10091 , n10092 , n10093 , n10094 , n10095 , n10096 , n10097 , n10098 , n10099 , n10100 , n10101 , n10102 , n10103 , n10104 , n10105 , n10106 , n10107 , n10108 , n10109 , n10110 , n10111 , n10112 , n10113 , n10114 , n10115 , n10116 , n10117 , n10118 , n10119 , n10120 , n10121 , n10122 , n10123 , n10124 , n10125 , n10126 , n10127 , n10128 , n10129 , n10130 , n10131 , n10132 , n10133 , n10134 , n10135 , n10136 , n10137 , n10138 , n10139 , n10140 , n10141 , n10142 , n10143 , n10144 , n10145 , n10146 , n10147 , n10148 , n10149 , n10150 , n10151 , n10152 , n10153 , n10154 , n10155 , n10156 , n10157 , n10158 , n10159 , n10160 , n10161 , n10162 , n10163 , n10164 , n10165 , n10166 , n10167 , n10168 , n10169 , n10170 , n10171 , n10172 , n10173 , n10174 , n10175 , n10176 , n10177 , n10178 , n10179 , n10180 , n10181 , n10182 , n10183 , n10184 , n10185 , n10186 , n10187 , n10188 , n10189 , n10190 , n10191 , n10192 , n10193 , n10194 , n10195 , n10196 , n10197 , n10198 , n10199 , n10200 , n10201 , n10202 , n10203 , n10204 , n10205 , n10206 , n10207 , n10208 , n10209 , n10210 , n10211 , n10212 , n10213 , n10214 , n10215 , n10216 , n10217 , n10218 , n10219 , n10220 , n10221 , n10222 , n10223 , n10224 , n10225 , n10226 , n10227 , n10228 , n10229 , n10230 , n10231 , n10232 , n10233 , n10234 , n10235 , n10236 , n10237 , n10238 , n10239 , n10240 , n10241 , n10242 , n10243 , n10244 , n10245 , n10246 , n10247 , n10248 , n10249 , n10250 , n10251 , n10252 , n10253 , n10254 , n10255 , n10256 , n10257 , n10258 , n10259 , n10260 , n10261 , n10262 , n10263 , n10264 , n10265 , n10266 , n10267 , n10268 , n10269 , n10270 , n10271 , n10272 , n10273 , n10274 , n10275 , n10276 , n10277 , n10278 , n10279 , n10280 , n10281 , n10282 , n10283 , n10284 , n10285 , n10286 , n10287 , n10288 , n10289 , n10290 , n10291 , n10292 , n10293 , n10294 , n10295 , n10296 , n10297 , n10298 , n10299 , n10300 , n10301 , n10302 , n10303 , n10304 , n10305 , n10306 , n10307 , n10308 , n10309 , n10310 , n10311 , n10312 , n10313 , n10314 , n10315 , n10316 , n10317 , n10318 , n10319 , n10320 , n10321 , n10322 , n10323 , n10324 , n10325 , n10326 , n10327 , n10328 , n10329 , n10330 , n10331 , n10332 , n10333 , n10334 , n10335 , n10336 , n10337 , n10338 , n10339 , n10340 , n10341 , n10342 , n10343 , n10344 , n10345 , n10346 , n10347 , n10348 , n10349 , n10350 , n10351 , n10352 , n10353 , n10354 , n10355 , n10356 , n10357 , n10358 , n10359 , n10360 , n10361 , n10362 , n10363 , n10364 , n10365 , n10366 , n10367 , n10368 , n10369 , n10370 , n10371 , n10372 , n10373 , n10374 , n10375 , n10376 , n10377 , n10378 , n10379 , n10380 , n10381 , n10382 , n10383 , n10384 , n10385 , n10386 , n10387 , n10388 , n10389 , n10390 , n10391 , n10392 , n10393 , n10394 , n10395 , n10396 , n10397 , n10398 , n10399 , n10400 , n10401 , n10402 , n10403 , n10404 , n10405 , n10406 , n10407 , n10408 , n10409 , n10410 , n10411 , n10412 , n10413 , n10414 , n10415 , n10416 , n10417 , n10418 , n10419 , n10420 , n10421 , n10422 , n10423 , n10424 , n10425 , n10426 , n10427 , n10428 , n10429 , n10430 , n10431 , n10432 , n10433 , n10434 , n10435 , n10436 , n10437 , n10438 , n10439 , n10440 , n10441 , n10442 , n10443 , n10444 , n10445 , n10446 , n10447 , n10448 , n10449 , n10450 , n10451 , n10452 , n10453 , n10454 , n10455 , n10456 , n10457 , n10458 , n10459 , n10460 , n10461 , n10462 , n10463 , n10464 , n10465 , n10466 , n10467 , n10468 , n10469 , n10470 , n10471 , n10472 , n10473 , n10474 , n10475 , n10476 , n10477 , n10478 , n10479 , n10480 , n10481 , n10482 , n10483 , n10484 , n10485 , n10486 , n10487 , n10488 , n10489 , n10490 , n10491 , n10492 , n10493 , n10494 , n10495 , n10496 , n10497 , n10498 , n10499 , n10500 , n10501 , n10502 , n10503 , n10504 , n10505 , n10506 , n10507 , n10508 , n10509 , n10510 , n10511 , n10512 , n10513 , n10514 , n10515 , n10516 , n10517 , n10518 , n10519 , n10520 , n10521 , n10522 , n10523 , n10524 , n10525 , n10526 , n10527 , n10528 , n10529 , n10530 , n10531 , n10532 , n10533 , n10534 , n10535 , n10536 , n10537 , n10538 , n10539 , n10540 , n10541 , n10542 , n10543 , n10544 , n10545 , n10546 , n10547 , n10548 , n10549 , n10550 , n10551 , n10552 , n10553 , n10554 , n10555 , n10556 , n10557 , n10558 , n10559 , n10560 , n10561 , n10562 , n10563 , n10564 , n10565 , n10566 , n10567 , n10568 , n10569 , n10570 , n10571 , n10572 , n10573 , n10574 , n10575 , n10576 , n10577 , n10578 , n10579 , n10580 , n10581 , n10582 , n10583 , n10584 , n10585 , n10586 , n10587 , n10588 , n10589 , n10590 , n10591 , n10592 , n10593 , n10594 , n10595 , n10596 , n10597 , n10598 , n10599 , n10600 , n10601 , n10602 , n10603 , n10604 , n10605 , n10606 , n10607 , n10608 , n10609 , n10610 , n10611 , n10612 , n10613 , n10614 , n10615 , n10616 , n10617 , n10618 , n10619 , n10620 , n10621 , n10622 , n10623 , n10624 , n10625 , n10626 , n10627 , n10628 , n10629 , n10630 , n10631 , n10632 , n10633 , n10634 , n10635 , n10636 , n10637 , n10638 , n10639 , n10640 , n10641 , n10642 , n10643 , n10644 , n10645 , n10646 , n10647 , n10648 , n10649 , n10650 , n10651 , n10652 , n10653 , n10654 , n10655 , n10656 , n10657 , n10658 , n10659 , n10660 , n10661 , n10662 , n10663 , n10664 , n10665 , n10666 , n10667 , n10668 , n10669 , n10670 , n10671 , n10672 , n10673 , n10674 , n10675 , n10676 , n10677 , n10678 , n10679 , n10680 , n10681 , n10682 , n10683 , n10684 , n10685 , n10686 , n10687 , n10688 , n10689 , n10690 , n10691 , n10692 , n10693 , n10694 , n10695 , n10696 , n10697 , n10698 , n10699 , n10700 , n10701 , n10702 , n10703 , n10704 , n10705 , n10706 , n10707 , n10708 , n10709 , n10710 , n10711 , n10712 , n10713 , n10714 , n10715 , n10716 , n10717 , n10718 , n10719 , n10720 , n10721 , n10722 , n10723 , n10724 , n10725 , n10726 , n10727 , n10728 , n10729 , n10730 , n10731 , n10732 , n10733 , n10734 , n10735 , n10736 , n10737 , n10738 , n10739 , n10740 , n10741 , n10742 , n10743 , n10744 , n10745 , n10746 , n10747 , n10748 , n10749 , n10750 , n10751 , n10752 , n10753 , n10754 , n10755 , n10756 , n10757 , n10758 , n10759 , n10760 , n10761 , n10762 , n10763 , n10764 , n10765 , n10766 , n10767 , n10768 , n10769 , n10770 , n10771 , n10772 , n10773 , n10774 , n10775 , n10776 , n10777 , n10778 , n10779 , n10780 , n10781 , n10782 , n10783 , n10784 , n10785 , n10786 , n10787 , n10788 , n10789 , n10790 , n10791 , n10792 , n10793 , n10794 , n10795 , n10796 , n10797 , n10798 , n10799 , n10800 , n10801 , n10802 , n10803 , n10804 , n10805 , n10806 , n10807 , n10808 , n10809 , n10810 , n10811 , n10812 , n10813 , n10814 , n10815 , n10816 , n10817 , n10818 , n10819 , n10820 , n10821 , n10822 , n10823 , n10824 , n10825 , n10826 , n10827 , n10828 , n10829 , n10830 , n10831 , n10832 , n10833 , n10834 , n10835 , n10836 , n10837 , n10838 , n10839 , n10840 , n10841 , n10842 , n10843 , n10844 , n10845 , n10846 , n10847 , n10848 , n10849 , n10850 , n10851 , n10852 , n10853 , n10854 , n10855 , n10856 , n10857 , n10858 , n10859 , n10860 , n10861 , n10862 , n10863 , n10864 , n10865 , n10866 , n10867 , n10868 , n10869 , n10870 , n10871 , n10872 , n10873 , n10874 , n10875 , n10876 , n10877 , n10878 , n10879 , n10880 , n10881 , n10882 , n10883 , n10884 , n10885 , n10886 , n10887 , n10888 , n10889 , n10890 , n10891 , n10892 , n10893 , n10894 , n10895 , n10896 , n10897 , n10898 , n10899 , n10900 , n10901 , n10902 , n10903 , n10904 , n10905 , n10906 , n10907 , n10908 , n10909 , n10910 , n10911 , n10912 , n10913 , n10914 , n10915 , n10916 , n10917 , n10918 , n10919 , n10920 , n10921 , n10922 , n10923 , n10924 , n10925 , n10926 , n10927 , n10928 , n10929 , n10930 , n10931 , n10932 , n10933 , n10934 , n10935 , n10936 , n10937 , n10938 , n10939 , n10940 , n10941 , n10942 , n10943 , n10944 , n10945 , n10946 , n10947 , n10948 , n10949 , n10950 , n10951 , n10952 , n10953 , n10954 , n10955 , n10956 , n10957 , n10958 , n10959 , n10960 , n10961 , n10962 , n10963 , n10964 , n10965 , n10966 , n10967 , n10968 , n10969 , n10970 , n10971 , n10972 , n10973 , n10974 , n10975 , n10976 , n10977 , n10978 , n10979 , n10980 , n10981 , n10982 , n10983 , n10984 , n10985 , n10986 , n10987 , n10988 , n10989 , n10990 , n10991 , n10992 , n10993 , n10994 , n10995 , n10996 , n10997 , n10998 , n10999 , n11000 , n11001 , n11002 , n11003 , n11004 , n11005 , n11006 , n11007 , n11008 , n11009 , n11010 , n11011 , n11012 , n11013 , n11014 , n11015 , n11016 , n11017 , n11018 , n11019 , n11020 , n11021 , n11022 , n11023 , n11024 , n11025 , n11026 , n11027 , n11028 , n11029 , n11030 , n11031 , n11032 , n11033 , n11034 , n11035 , n11036 , n11037 , n11038 , n11039 , n11040 , n11041 , n11042 , n11043 , n11044 , n11045 , n11046 , n11047 , n11048 , n11049 , n11050 , n11051 , n11052 , n11053 , n11054 , n11055 , n11056 , n11057 , n11058 , n11059 , n11060 , n11061 , n11062 , n11063 , n11064 , n11065 , n11066 , n11067 , n11068 , n11069 , n11070 , n11071 , n11072 , n11073 , n11074 , n11075 , n11076 , n11077 , n11078 , n11079 , n11080 , n11081 , n11082 , n11083 , n11084 , n11085 , n11086 , n11087 , n11088 , n11089 , n11090 , n11091 , n11092 , n11093 , n11094 , n11095 , n11096 , n11097 , n11098 , n11099 , n11100 , n11101 , n11102 , n11103 , n11104 , n11105 , n11106 , n11107 , n11108 , n11109 , n11110 , n11111 , n11112 , n11113 , n11114 , n11115 , n11116 , n11117 , n11118 , n11119 , n11120 , n11121 , n11122 , n11123 , n11124 , n11125 , n11126 , n11127 , n11128 , n11129 , n11130 , n11131 , n11132 , n11133 , n11134 , n11135 , n11136 , n11137 , n11138 , n11139 , n11140 , n11141 , n11142 , n11143 , n11144 , n11145 , n11146 , n11147 , n11148 , n11149 , n11150 , n11151 , n11152 , n11153 , n11154 , n11155 , n11156 , n11157 , n11158 , n11159 , n11160 , n11161 , n11162 , n11163 , n11164 , n11165 , n11166 , n11167 , n11168 , n11169 , n11170 , n11171 , n11172 , n11173 , n11174 , n11175 , n11176 , n11177 , n11178 , n11179 , n11180 , n11181 , n11182 , n11183 , n11184 , n11185 , n11186 , n11187 , n11188 , n11189 , n11190 , n11191 , n11192 , n11193 , n11194 , n11195 , n11196 , n11197 , n11198 , n11199 , n11200 , n11201 , n11202 , n11203 , n11204 , n11205 , n11206 , n11207 , n11208 , n11209 , n11210 , n11211 , n11212 , n11213 , n11214 , n11215 , n11216 , n11217 , n11218 , n11219 , n11220 , n11221 , n11222 , n11223 , n11224 , n11225 , n11226 , n11227 , n11228 , n11229 , n11230 , n11231 , n11232 , n11233 , n11234 , n11235 , n11236 , n11237 , n11238 , n11239 , n11240 , n11241 , n11242 , n11243 , n11244 , n11245 , n11246 , n11247 , n11248 , n11249 , n11250 , n11251 , n11252 , n11253 , n11254 , n11255 , n11256 , n11257 , n11258 , n11259 , n11260 , n11261 , n11262 , n11263 , n11264 , n11265 , n11266 , n11267 , n11268 , n11269 , n11270 , n11271 , n11272 , n11273 , n11274 , n11275 , n11276 , n11277 , n11278 , n11279 , n11280 , n11281 , n11282 , n11283 , n11284 , n11285 , n11286 , n11287 , n11288 , n11289 , n11290 , n11291 , n11292 , n11293 , n11294 , n11295 , n11296 , n11297 , n11298 , n11299 , n11300 , n11301 , n11302 , n11303 , n11304 , n11305 , n11306 , n11307 , n11308 , n11309 , n11310 , n11311 , n11312 , n11313 , n11314 , n11315 , n11316 , n11317 , n11318 , n11319 , n11320 , n11321 , n11322 , n11323 , n11324 , n11325 , n11326 , n11327 , n11328 , n11329 , n11330 , n11331 , n11332 , n11333 , n11334 , n11335 , n11336 , n11337 , n11338 , n11339 , n11340 , n11341 , n11342 , n11343 , n11344 , n11345 , n11346 , n11347 , n11348 , n11349 , n11350 , n11351 , n11352 , n11353 , n11354 , n11355 , n11356 , n11357 , n11358 , n11359 , n11360 , n11361 , n11362 , n11363 , n11364 , n11365 , n11366 , n11367 , n11368 , n11369 , n11370 , n11371 , n11372 , n11373 , n11374 , n11375 , n11376 , n11377 , n11378 , n11379 , n11380 , n11381 , n11382 , n11383 , n11384 , n11385 , n11386 , n11387 , n11388 , n11389 , n11390 , n11391 , n11392 , n11393 , n11394 , n11395 , n11396 , n11397 , n11398 , n11399 , n11400 , n11401 , n11402 , n11403 , n11404 , n11405 , n11406 , n11407 , n11408 , n11409 , n11410 , n11411 , n11412 , n11413 , n11414 , n11415 , n11416 , n11417 , n11418 , n11419 , n11420 , n11421 , n11422 , n11423 , n11424 , n11425 , n11426 , n11427 , n11428 , n11429 , n11430 , n11431 , n11432 , n11433 , n11434 , n11435 , n11436 , n11437 , n11438 , n11439 , n11440 , n11441 , n11442 , n11443 , n11444 , n11445 , n11446 , n11447 , n11448 , n11449 , n11450 , n11451 , n11452 , n11453 , n11454 , n11455 , n11456 , n11457 , n11458 , n11459 , n11460 , n11461 , n11462 , n11463 , n11464 , n11465 , n11466 , n11467 , n11468 , n11469 , n11470 , n11471 , n11472 , n11473 , n11474 , n11475 , n11476 , n11477 , n11478 , n11479 , n11480 , n11481 , n11482 , n11483 , n11484 , n11485 , n11486 , n11487 , n11488 , n11489 , n11490 , n11491 , n11492 , n11493 , n11494 , n11495 , n11496 , n11497 , n11498 , n11499 , n11500 , n11501 , n11502 , n11503 , n11504 , n11505 , n11506 , n11507 , n11508 , n11509 , n11510 , n11511 , n11512 , n11513 , n11514 , n11515 , n11516 , n11517 , n11518 , n11519 , n11520 , n11521 , n11522 , n11523 , n11524 , n11525 , n11526 , n11527 , n11528 , n11529 , n11530 , n11531 , n11532 , n11533 , n11534 , n11535 , n11536 , n11537 , n11538 , n11539 , n11540 , n11541 , n11542 , n11543 , n11544 , n11545 , n11546 , n11547 , n11548 , n11549 , n11550 , n11551 , n11552 , n11553 , n11554 , n11555 , n11556 , n11557 , n11558 , n11559 , n11560 , n11561 , n11562 , n11563 , n11564 , n11565 , n11566 , n11567 , n11568 , n11569 , n11570 , n11571 , n11572 , n11573 , n11574 , n11575 , n11576 , n11577 , n11578 , n11579 , n11580 , n11581 , n11582 , n11583 , n11584 , n11585 , n11586 , n11587 , n11588 , n11589 , n11590 , n11591 , n11592 , n11593 , n11594 , n11595 , n11596 , n11597 , n11598 , n11599 , n11600 , n11601 , n11602 , n11603 , n11604 , n11605 , n11606 , n11607 , n11608 , n11609 , n11610 , n11611 , n11612 , n11613 , n11614 , n11615 , n11616 , n11617 , n11618 , n11619 , n11620 , n11621 , n11622 , n11623 , n11624 , n11625 , n11626 , n11627 , n11628 , n11629 , n11630 , n11631 , n11632 , n11633 , n11634 , n11635 , n11636 , n11637 , n11638 , n11639 , n11640 , n11641 , n11642 , n11643 , n11644 , n11645 , n11646 , n11647 , n11648 , n11649 , n11650 , n11651 , n11652 , n11653 , n11654 , n11655 , n11656 , n11657 , n11658 , n11659 , n11660 , n11661 , n11662 , n11663 , n11664 , n11665 , n11666 , n11667 , n11668 , n11669 , n11670 , n11671 , n11672 , n11673 , n11674 , n11675 , n11676 , n11677 , n11678 , n11679 , n11680 , n11681 , n11682 , n11683 , n11684 , n11685 , n11686 , n11687 , n11688 , n11689 , n11690 , n11691 , n11692 , n11693 , n11694 , n11695 , n11696 , n11697 , n11698 , n11699 , n11700 , n11701 , n11702 , n11703 , n11704 , n11705 , n11706 , n11707 , n11708 , n11709 , n11710 , n11711 , n11712 , n11713 , n11714 , n11715 , n11716 , n11717 , n11718 , n11719 , n11720 , n11721 , n11722 , n11723 , n11724 , n11725 , n11726 , n11727 , n11728 , n11729 , n11730 , n11731 , n11732 , n11733 , n11734 , n11735 , n11736 , n11737 , n11738 , n11739 , n11740 , n11741 , n11742 , n11743 , n11744 , n11745 , n11746 , n11747 , n11748 , n11749 , n11750 , n11751 , n11752 , n11753 , n11754 , n11755 , n11756 , n11757 , n11758 , n11759 , n11760 , n11761 , n11762 , n11763 , n11764 , n11765 , n11766 , n11767 , n11768 , n11769 , n11770 , n11771 , n11772 , n11773 , n11774 , n11775 , n11776 , n11777 , n11778 , n11779 , n11780 , n11781 , n11782 , n11783 , n11784 , n11785 , n11786 , n11787 , n11788 , n11789 , n11790 , n11791 , n11792 , n11793 , n11794 , n11795 , n11796 , n11797 , n11798 , n11799 , n11800 , n11801 , n11802 , n11803 , n11804 , n11805 , n11806 , n11807 , n11808 , n11809 , n11810 , n11811 , n11812 , n11813 , n11814 , n11815 , n11816 , n11817 , n11818 , n11819 , n11820 , n11821 , n11822 , n11823 , n11824 , n11825 , n11826 , n11827 , n11828 , n11829 , n11830 , n11831 , n11832 , n11833 , n11834 , n11835 , n11836 , n11837 , n11838 , n11839 , n11840 , n11841 , n11842 , n11843 , n11844 , n11845 , n11846 , n11847 , n11848 , n11849 , n11850 , n11851 , n11852 , n11853 , n11854 , n11855 , n11856 , n11857 , n11858 , n11859 , n11860 , n11861 , n11862 , n11863 , n11864 , n11865 , n11866 , n11867 , n11868 , n11869 , n11870 , n11871 , n11872 , n11873 , n11874 , n11875 , n11876 , n11877 , n11878 , n11879 , n11880 , n11881 , n11882 , n11883 , n11884 , n11885 , n11886 , n11887 , n11888 , n11889 , n11890 , n11891 , n11892 , n11893 , n11894 , n11895 , n11896 , n11897 , n11898 , n11899 , n11900 , n11901 , n11902 , n11903 , n11904 , n11905 , n11906 , n11907 , n11908 , n11909 , n11910 , n11911 , n11912 , n11913 , n11914 , n11915 , n11916 , n11917 , n11918 , n11919 , n11920 , n11921 , n11922 , n11923 , n11924 , n11925 , n11926 , n11927 , n11928 , n11929 , n11930 , n11931 , n11932 , n11933 , n11934 , n11935 , n11936 , n11937 , n11938 , n11939 , n11940 , n11941 , n11942 , n11943 , n11944 , n11945 , n11946 , n11947 , n11948 , n11949 , n11950 , n11951 , n11952 , n11953 , n11954 , n11955 , n11956 , n11957 , n11958 , n11959 , n11960 , n11961 , n11962 , n11963 , n11964 , n11965 , n11966 , n11967 , n11968 , n11969 , n11970 , n11971 , n11972 , n11973 , n11974 , n11975 , n11976 , n11977 , n11978 , n11979 , n11980 , n11981 , n11982 , n11983 , n11984 , n11985 , n11986 , n11987 , n11988 , n11989 , n11990 , n11991 , n11992 , n11993 , n11994 , n11995 , n11996 , n11997 , n11998 , n11999 , n12000 , n12001 , n12002 , n12003 , n12004 , n12005 , n12006 , n12007 , n12008 , n12009 , n12010 , n12011 , n12012 , n12013 , n12014 , n12015 , n12016 , n12017 , n12018 , n12019 , n12020 , n12021 , n12022 , n12023 , n12024 , n12025 , n12026 , n12027 , n12028 , n12029 , n12030 , n12031 , n12032 , n12033 , n12034 , n12035 , n12036 , n12037 , n12038 , n12039 , n12040 , n12041 , n12042 , n12043 , n12044 , n12045 , n12046 , n12047 , n12048 , n12049 , n12050 , n12051 , n12052 , n12053 , n12054 , n12055 , n12056 , n12057 , n12058 , n12059 , n12060 , n12061 , n12062 , n12063 , n12064 , n12065 , n12066 , n12067 , n12068 , n12069 , n12070 , n12071 , n12072 , n12073 , n12074 , n12075 , n12076 , n12077 , n12078 , n12079 , n12080 , n12081 , n12082 , n12083 , n12084 , n12085 , n12086 , n12087 , n12088 , n12089 , n12090 , n12091 , n12092 , n12093 , n12094 , n12095 , n12096 , n12097 , n12098 , n12099 , n12100 , n12101 , n12102 , n12103 , n12104 , n12105 , n12106 , n12107 , n12108 , n12109 , n12110 , n12111 , n12112 , n12113 , n12114 , n12115 , n12116 , n12117 , n12118 , n12119 , n12120 , n12121 , n12122 , n12123 , n12124 , n12125 , n12126 , n12127 , n12128 , n12129 , n12130 , n12131 , n12132 , n12133 , n12134 , n12135 , n12136 , n12137 , n12138 , n12139 , n12140 , n12141 , n12142 , n12143 , n12144 , n12145 , n12146 , n12147 , n12148 , n12149 , n12150 , n12151 , n12152 , n12153 , n12154 , n12155 , n12156 , n12157 , n12158 , n12159 , n12160 , n12161 , n12162 , n12163 , n12164 , n12165 , n12166 , n12167 , n12168 , n12169 , n12170 , n12171 , n12172 , n12173 , n12174 , n12175 , n12176 , n12177 , n12178 , n12179 , n12180 , n12181 , n12182 , n12183 , n12184 , n12185 , n12186 , n12187 , n12188 , n12189 , n12190 , n12191 , n12192 , n12193 , n12194 , n12195 , n12196 , n12197 , n12198 , n12199 , n12200 , n12201 , n12202 , n12203 , n12204 , n12205 , n12206 , n12207 , n12208 , n12209 , n12210 , n12211 , n12212 , n12213 , n12214 , n12215 , n12216 , n12217 , n12218 , n12219 , n12220 , n12221 , n12222 , n12223 , n12224 , n12225 , n12226 , n12227 , n12228 , n12229 , n12230 , n12231 , n12232 , n12233 , n12234 , n12235 , n12236 , n12237 , n12238 , n12239 , n12240 , n12241 , n12242 , n12243 , n12244 , n12245 , n12246 , n12247 , n12248 , n12249 , n12250 , n12251 , n12252 , n12253 , n12254 , n12255 , n12256 , n12257 , n12258 , n12259 , n12260 , n12261 , n12262 , n12263 , n12264 , n12265 , n12266 , n12267 , n12268 , n12269 , n12270 , n12271 , n12272 , n12273 , n12274 , n12275 , n12276 , n12277 , n12278 , n12279 , n12280 , n12281 , n12282 , n12283 , n12284 , n12285 , n12286 , n12287 , n12288 , n12289 , n12290 , n12291 , n12292 , n12293 , n12294 , n12295 , n12296 , n12297 , n12298 , n12299 , n12300 , n12301 , n12302 , n12303 , n12304 , n12305 , n12306 , n12307 , n12308 , n12309 , n12310 , n12311 , n12312 , n12313 , n12314 , n12315 , n12316 , n12317 , n12318 , n12319 , n12320 , n12321 , n12322 , n12323 , n12324 , n12325 , n12326 , n12327 , n12328 , n12329 , n12330 , n12331 , n12332 , n12333 , n12334 , n12335 , n12336 , n12337 , n12338 , n12339 , n12340 , n12341 , n12342 , n12343 , n12344 , n12345 , n12346 , n12347 , n12348 , n12349 , n12350 , n12351 , n12352 , n12353 , n12354 , n12355 , n12356 , n12357 , n12358 , n12359 , n12360 , n12361 , n12362 , n12363 , n12364 , n12365 , n12366 , n12367 , n12368 , n12369 , n12370 , n12371 , n12372 , n12373 , n12374 , n12375 , n12376 , n12377 , n12378 , n12379 , n12380 , n12381 , n12382 , n12383 , n12384 , n12385 , n12386 , n12387 , n12388 , n12389 , n12390 , n12391 , n12392 , n12393 , n12394 , n12395 , n12396 , n12397 , n12398 , n12399 , n12400 , n12401 , n12402 , n12403 , n12404 , n12405 , n12406 , n12407 , n12408 , n12409 , n12410 , n12411 , n12412 , n12413 , n12414 , n12415 , n12416 , n12417 , n12418 , n12419 , n12420 , n12421 , n12422 , n12423 , n12424 , n12425 , n12426 , n12427 , n12428 , n12429 , n12430 , n12431 , n12432 , n12433 , n12434 , n12435 , n12436 , n12437 , n12438 , n12439 , n12440 , n12441 , n12442 , n12443 , n12444 , n12445 , n12446 , n12447 , n12448 , n12449 , n12450 , n12451 , n12452 , n12453 , n12454 , n12455 , n12456 , n12457 , n12458 , n12459 , n12460 , n12461 , n12462 , n12463 , n12464 , n12465 , n12466 , n12467 , n12468 , n12469 , n12470 , n12471 , n12472 , n12473 , n12474 , n12475 , n12476 , n12477 , n12478 , n12479 , n12480 , n12481 , n12482 , n12483 , n12484 , n12485 , n12486 , n12487 , n12488 , n12489 , n12490 , n12491 , n12492 , n12493 , n12494 , n12495 , n12496 , n12497 , n12498 , n12499 , n12500 , n12501 , n12502 , n12503 , n12504 , n12505 , n12506 , n12507 , n12508 , n12509 , n12510 , n12511 , n12512 , n12513 , n12514 , n12515 , n12516 , n12517 , n12518 , n12519 , n12520 , n12521 , n12522 , n12523 , n12524 , n12525 , n12526 , n12527 , n12528 , n12529 , n12530 , n12531 , n12532 , n12533 , n12534 , n12535 , n12536 , n12537 , n12538 , n12539 , n12540 , n12541 , n12542 , n12543 , n12544 , n12545 , n12546 , n12547 , n12548 , n12549 , n12550 , n12551 , n12552 , n12553 , n12554 , n12555 , n12556 , n12557 , n12558 , n12559 , n12560 , n12561 , n12562 , n12563 , n12564 , n12565 , n12566 , n12567 , n12568 , n12569 , n12570 , n12571 , n12572 , n12573 , n12574 , n12575 , n12576 , n12577 , n12578 , n12579 , n12580 , n12581 , n12582 , n12583 , n12584 , n12585 , n12586 , n12587 , n12588 , n12589 , n12590 , n12591 , n12592 , n12593 , n12594 , n12595 , n12596 , n12597 , n12598 , n12599 , n12600 , n12601 , n12602 , n12603 , n12604 , n12605 , n12606 , n12607 , n12608 , n12609 , n12610 , n12611 , n12612 , n12613 , n12614 , n12615 , n12616 , n12617 , n12618 , n12619 , n12620 , n12621 , n12622 , n12623 , n12624 , n12625 , n12626 , n12627 , n12628 , n12629 , n12630 , n12631 , n12632 , n12633 , n12634 , n12635 , n12636 , n12637 , n12638 , n12639 , n12640 , n12641 , n12642 , n12643 , n12644 , n12645 , n12646 , n12647 , n12648 , n12649 , n12650 , n12651 , n12652 , n12653 , n12654 , n12655 , n12656 , n12657 , n12658 , n12659 , n12660 , n12661 , n12662 , n12663 , n12664 , n12665 , n12666 , n12667 , n12668 , n12669 , n12670 , n12671 , n12672 , n12673 , n12674 , n12675 , n12676 , n12677 , n12678 , n12679 , n12680 , n12681 , n12682 , n12683 , n12684 , n12685 , n12686 , n12687 , n12688 , n12689 , n12690 , n12691 , n12692 , n12693 , n12694 , n12695 , n12696 , n12697 , n12698 , n12699 , n12700 , n12701 , n12702 , n12703 , n12704 , n12705 , n12706 , n12707 , n12708 , n12709 , n12710 , n12711 , n12712 , n12713 , n12714 , n12715 , n12716 , n12717 , n12718 , n12719 , n12720 , n12721 , n12722 , n12723 , n12724 , n12725 , n12726 , n12727 , n12728 , n12729 , n12730 , n12731 , n12732 , n12733 , n12734 , n12735 , n12736 , n12737 , n12738 , n12739 , n12740 , n12741 , n12742 , n12743 , n12744 , n12745 , n12746 , n12747 , n12748 , n12749 , n12750 , n12751 , n12752 , n12753 , n12754 , n12755 , n12756 , n12757 , n12758 , n12759 , n12760 , n12761 , n12762 , n12763 , n12764 , n12765 , n12766 , n12767 , n12768 , n12769 , n12770 , n12771 , n12772 , n12773 , n12774 , n12775 , n12776 , n12777 , n12778 , n12779 , n12780 , n12781 , n12782 , n12783 , n12784 , n12785 , n12786 , n12787 , n12788 , n12789 , n12790 , n12791 , n12792 , n12793 , n12794 , n12795 , n12796 , n12797 , n12798 , n12799 , n12800 , n12801 , n12802 , n12803 , n12804 , n12805 , n12806 , n12807 , n12808 , n12809 , n12810 , n12811 , n12812 , n12813 , n12814 , n12815 , n12816 , n12817 , n12818 , n12819 , n12820 , n12821 , n12822 , n12823 , n12824 , n12825 , n12826 , n12827 , n12828 , n12829 , n12830 , n12831 , n12832 , n12833 , n12834 , n12835 , n12836 , n12837 , n12838 , n12839 , n12840 , n12841 , n12842 , n12843 , n12844 , n12845 , n12846 , n12847 , n12848 , n12849 , n12850 , n12851 , n12852 , n12853 , n12854 , n12855 , n12856 , n12857 , n12858 , n12859 , n12860 , n12861 , n12862 , n12863 , n12864 , n12865 , n12866 , n12867 , n12868 , n12869 , n12870 , n12871 , n12872 , n12873 , n12874 , n12875 , n12876 , n12877 , n12878 , n12879 , n12880 , n12881 , n12882 , n12883 , n12884 , n12885 , n12886 , n12887 , n12888 , n12889 , n12890 , n12891 , n12892 , n12893 , n12894 , n12895 , n12896 , n12897 , n12898 , n12899 , n12900 , n12901 , n12902 , n12903 , n12904 , n12905 , n12906 , n12907 , n12908 , n12909 , n12910 , n12911 , n12912 , n12913 , n12914 , n12915 , n12916 , n12917 , n12918 , n12919 , n12920 , n12921 , n12922 , n12923 , n12924 , n12925 , n12926 , n12927 , n12928 , n12929 , n12930 , n12931 , n12932 , n12933 , n12934 , n12935 , n12936 , n12937 , n12938 , n12939 , n12940 , n12941 , n12942 , n12943 , n12944 , n12945 , n12946 , n12947 , n12948 , n12949 , n12950 , n12951 , n12952 , n12953 , n12954 , n12955 , n12956 , n12957 , n12958 , n12959 , n12960 , n12961 , n12962 , n12963 , n12964 , n12965 , n12966 , n12967 , n12968 , n12969 , n12970 , n12971 , n12972 , n12973 , n12974 , n12975 , n12976 , n12977 , n12978 , n12979 , n12980 , n12981 , n12982 , n12983 , n12984 , n12985 , n12986 , n12987 , n12988 , n12989 , n12990 , n12991 , n12992 , n12993 , n12994 , n12995 , n12996 , n12997 , n12998 , n12999 , n13000 , n13001 , n13002 , n13003 , n13004 , n13005 , n13006 , n13007 , n13008 , n13009 , n13010 , n13011 , n13012 , n13013 , n13014 , n13015 , n13016 , n13017 , n13018 , n13019 , n13020 , n13021 , n13022 , n13023 , n13024 , n13025 , n13026 , n13027 , n13028 , n13029 , n13030 , n13031 , n13032 , n13033 , n13034 , n13035 , n13036 , n13037 , n13038 , n13039 , n13040 , n13041 , n13042 , n13043 , n13044 , n13045 , n13046 , n13047 , n13048 , n13049 , n13050 , n13051 , n13052 , n13053 , n13054 , n13055 , n13056 , n13057 , n13058 , n13059 , n13060 , n13061 , n13062 , n13063 , n13064 , n13065 , n13066 , n13067 , n13068 , n13069 , n13070 , n13071 , n13072 , n13073 , n13074 , n13075 , n13076 , n13077 , n13078 , n13079 , n13080 , n13081 , n13082 , n13083 , n13084 , n13085 , n13086 , n13087 , n13088 , n13089 , n13090 , n13091 , n13092 , n13093 , n13094 , n13095 , n13096 , n13097 , n13098 , n13099 , n13100 , n13101 , n13102 , n13103 , n13104 , n13105 , n13106 , n13107 , n13108 , n13109 , n13110 , n13111 , n13112 , n13113 , n13114 , n13115 , n13116 , n13117 , n13118 , n13119 , n13120 , n13121 , n13122 , n13123 , n13124 , n13125 , n13126 , n13127 , n13128 , n13129 , n13130 , n13131 , n13132 , n13133 , n13134 , n13135 , n13136 , n13137 , n13138 , n13139 , n13140 , n13141 , n13142 , n13143 , n13144 , n13145 , n13146 , n13147 , n13148 , n13149 , n13150 , n13151 , n13152 , n13153 , n13154 , n13155 , n13156 , n13157 , n13158 , n13159 , n13160 , n13161 , n13162 , n13163 , n13164 , n13165 , n13166 , n13167 , n13168 , n13169 , n13170 , n13171 , n13172 , n13173 , n13174 , n13175 , n13176 , n13177 , n13178 , n13179 , n13180 , n13181 , n13182 , n13183 , n13184 , n13185 , n13186 , n13187 , n13188 , n13189 , n13190 , n13191 , n13192 , n13193 , n13194 , n13195 , n13196 , n13197 , n13198 , n13199 , n13200 , n13201 , n13202 , n13203 , n13204 , n13205 , n13206 , n13207 , n13208 , n13209 , n13210 , n13211 , n13212 , n13213 , n13214 , n13215 , n13216 , n13217 , n13218 , n13219 , n13220 , n13221 , n13222 , n13223 , n13224 , n13225 , n13226 , n13227 , n13228 , n13229 , n13230 , n13231 , n13232 , n13233 , n13234 , n13235 , n13236 , n13237 , n13238 , n13239 , n13240 , n13241 , n13242 , n13243 , n13244 , n13245 , n13246 , n13247 , n13248 , n13249 , n13250 , n13251 , n13252 , n13253 , n13254 , n13255 , n13256 , n13257 , n13258 , n13259 , n13260 , n13261 , n13262 , n13263 , n13264 , n13265 , n13266 , n13267 , n13268 , n13269 , n13270 , n13271 , n13272 , n13273 , n13274 , n13275 , n13276 , n13277 , n13278 , n13279 , n13280 , n13281 , n13282 , n13283 , n13284 , n13285 , n13286 , n13287 , n13288 , n13289 , n13290 , n13291 , n13292 , n13293 , n13294 , n13295 , n13296 , n13297 , n13298 , n13299 , n13300 , n13301 , n13302 , n13303 , n13304 , n13305 , n13306 , n13307 , n13308 , n13309 , n13310 , n13311 , n13312 , n13313 , n13314 , n13315 , n13316 , n13317 , n13318 , n13319 , n13320 , n13321 , n13322 , n13323 , n13324 , n13325 , n13326 , n13327 , n13328 , n13329 , n13330 , n13331 , n13332 , n13333 , n13334 , n13335 , n13336 , n13337 , n13338 , n13339 , n13340 , n13341 , n13342 , n13343 , n13344 , n13345 , n13346 , n13347 , n13348 , n13349 , n13350 , n13351 , n13352 , n13353 , n13354 , n13355 , n13356 , n13357 , n13358 , n13359 , n13360 , n13361 , n13362 , n13363 , n13364 , n13365 , n13366 , n13367 , n13368 , n13369 , n13370 , n13371 , n13372 , n13373 , n13374 , n13375 , n13376 , n13377 , n13378 , n13379 , n13380 , n13381 , n13382 , n13383 , n13384 , n13385 , n13386 , n13387 , n13388 , n13389 , n13390 , n13391 , n13392 , n13393 , n13394 , n13395 , n13396 , n13397 , n13398 , n13399 , n13400 , n13401 , n13402 , n13403 , n13404 , n13405 , n13406 , n13407 , n13408 , n13409 , n13410 , n13411 , n13412 , n13413 , n13414 , n13415 , n13416 , n13417 , n13418 , n13419 , n13420 , n13421 , n13422 , n13423 , n13424 , n13425 , n13426 , n13427 , n13428 , n13429 , n13430 , n13431 , n13432 , n13433 , n13434 , n13435 , n13436 , n13437 , n13438 , n13439 , n13440 , n13441 , n13442 , n13443 , n13444 , n13445 , n13446 , n13447 , n13448 , n13449 , n13450 , n13451 , n13452 , n13453 , n13454 , n13455 , n13456 , n13457 , n13458 , n13459 , n13460 , n13461 , n13462 , n13463 , n13464 , n13465 , n13466 , n13467 , n13468 , n13469 , n13470 , n13471 , n13472 , n13473 , n13474 , n13475 , n13476 , n13477 , n13478 , n13479 , n13480 , n13481 , n13482 , n13483 , n13484 , n13485 , n13486 , n13487 , n13488 , n13489 , n13490 , n13491 , n13492 , n13493 , n13494 , n13495 , n13496 , n13497 , n13498 , n13499 , n13500 , n13501 , n13502 , n13503 , n13504 , n13505 , n13506 , n13507 , n13508 , n13509 , n13510 , n13511 , n13512 , n13513 , n13514 , n13515 , n13516 , n13517 , n13518 , n13519 , n13520 , n13521 , n13522 , n13523 , n13524 , n13525 , n13526 , n13527 , n13528 , n13529 , n13530 , n13531 , n13532 , n13533 , n13534 , n13535 , n13536 , n13537 , n13538 , n13539 , n13540 , n13541 , n13542 , n13543 , n13544 , n13545 , n13546 , n13547 , n13548 , n13549 , n13550 , n13551 , n13552 , n13553 , n13554 , n13555 , n13556 , n13557 , n13558 , n13559 , n13560 , n13561 , n13562 , n13563 , n13564 , n13565 , n13566 , n13567 , n13568 , n13569 , n13570 , n13571 , n13572 , n13573 , n13574 , n13575 , n13576 , n13577 , n13578 , n13579 , n13580 , n13581 , n13582 , n13583 , n13584 , n13585 , n13586 , n13587 , n13588 , n13589 , n13590 , n13591 , n13592 , n13593 , n13594 , n13595 , n13596 , n13597 , n13598 , n13599 , n13600 , n13601 , n13602 , n13603 , n13604 , n13605 , n13606 , n13607 , n13608 , n13609 , n13610 , n13611 , n13612 , n13613 , n13614 , n13615 , n13616 , n13617 , n13618 , n13619 , n13620 , n13621 , n13622 , n13623 , n13624 , n13625 , n13626 , n13627 , n13628 , n13629 , n13630 , n13631 , n13632 , n13633 , n13634 , n13635 , n13636 , n13637 , n13638 , n13639 , n13640 , n13641 , n13642 , n13643 , n13644 , n13645 , n13646 , n13647 , n13648 , n13649 , n13650 , n13651 , n13652 , n13653 , n13654 , n13655 , n13656 , n13657 , n13658 , n13659 , n13660 , n13661 , n13662 , n13663 , n13664 , n13665 , n13666 , n13667 , n13668 , n13669 , n13670 , n13671 , n13672 , n13673 , n13674 , n13675 , n13676 , n13677 , n13678 , n13679 , n13680 , n13681 , n13682 , n13683 , n13684 , n13685 , n13686 , n13687 , n13688 , n13689 , n13690 , n13691 , n13692 , n13693 , n13694 , n13695 , n13696 , n13697 , n13698 , n13699 , n13700 , n13701 , n13702 , n13703 , n13704 , n13705 , n13706 , n13707 , n13708 , n13709 , n13710 , n13711 , n13712 , n13713 , n13714 , n13715 , n13716 , n13717 , n13718 , n13719 , n13720 , n13721 , n13722 , n13723 , n13724 , n13725 , n13726 , n13727 , n13728 , n13729 , n13730 , n13731 , n13732 , n13733 , n13734 , n13735 , n13736 , n13737 , n13738 , n13739 , n13740 , n13741 , n13742 , n13743 , n13744 , n13745 , n13746 , n13747 , n13748 , n13749 , n13750 , n13751 , n13752 , n13753 , n13754 , n13755 , n13756 , n13757 , n13758 , n13759 , n13760 , n13761 , n13762 , n13763 , n13764 , n13765 , n13766 , n13767 , n13768 , n13769 , n13770 , n13771 , n13772 , n13773 , n13774 , n13775 , n13776 , n13777 , n13778 , n13779 , n13780 , n13781 , n13782 , n13783 , n13784 , n13785 , n13786 , n13787 , n13788 , n13789 , n13790 , n13791 , n13792 , n13793 , n13794 , n13795 , n13796 , n13797 , n13798 , n13799 , n13800 , n13801 , n13802 , n13803 , n13804 , n13805 , n13806 , n13807 , n13808 , n13809 , n13810 , n13811 , n13812 , n13813 , n13814 , n13815 , n13816 , n13817 , n13818 , n13819 , n13820 , n13821 , n13822 , n13823 , n13824 , n13825 , n13826 , n13827 , n13828 , n13829 , n13830 , n13831 , n13832 , n13833 , n13834 , n13835 , n13836 , n13837 , n13838 , n13839 , n13840 , n13841 , n13842 , n13843 , n13844 , n13845 , n13846 , n13847 , n13848 , n13849 , n13850 , n13851 , n13852 , n13853 , n13854 , n13855 , n13856 , n13857 , n13858 , n13859 , n13860 , n13861 , n13862 , n13863 , n13864 , n13865 , n13866 , n13867 , n13868 , n13869 , n13870 , n13871 , n13872 , n13873 , n13874 , n13875 , n13876 , n13877 , n13878 , n13879 , n13880 , n13881 , n13882 , n13883 , n13884 , n13885 , n13886 , n13887 , n13888 , n13889 , n13890 , n13891 , n13892 , n13893 , n13894 , n13895 , n13896 , n13897 , n13898 , n13899 , n13900 , n13901 , n13902 , n13903 , n13904 , n13905 , n13906 , n13907 , n13908 , n13909 , n13910 , n13911 , n13912 , n13913 , n13914 , n13915 , n13916 , n13917 , n13918 , n13919 , n13920 , n13921 , n13922 , n13923 , n13924 , n13925 , n13926 , n13927 , n13928 , n13929 , n13930 , n13931 , n13932 , n13933 , n13934 , n13935 , n13936 , n13937 , n13938 , n13939 , n13940 , n13941 , n13942 , n13943 , n13944 , n13945 , n13946 , n13947 , n13948 , n13949 , n13950 , n13951 , n13952 , n13953 , n13954 , n13955 , n13956 , n13957 , n13958 , n13959 , n13960 , n13961 , n13962 , n13963 , n13964 , n13965 , n13966 , n13967 , n13968 , n13969 , n13970 , n13971 , n13972 , n13973 , n13974 , n13975 , n13976 , n13977 , n13978 , n13979 , n13980 , n13981 , n13982 , n13983 , n13984 , n13985 , n13986 , n13987 , n13988 , n13989 , n13990 , n13991 , n13992 , n13993 , n13994 , n13995 , n13996 , n13997 , n13998 , n13999 , n14000 , n14001 , n14002 , n14003 , n14004 , n14005 , n14006 , n14007 , n14008 , n14009 , n14010 , n14011 , n14012 , n14013 , n14014 , n14015 , n14016 , n14017 , n14018 , n14019 , n14020 , n14021 , n14022 , n14023 , n14024 , n14025 , n14026 , n14027 , n14028 , n14029 , n14030 , n14031 , n14032 , n14033 , n14034 , n14035 , n14036 , n14037 , n14038 , n14039 , n14040 , n14041 , n14042 , n14043 , n14044 , n14045 , n14046 , n14047 , n14048 , n14049 , n14050 , n14051 , n14052 , n14053 , n14054 , n14055 , n14056 , n14057 , n14058 , n14059 , n14060 , n14061 , n14062 , n14063 , n14064 , n14065 , n14066 , n14067 , n14068 , n14069 , n14070 , n14071 , n14072 , n14073 , n14074 , n14075 , n14076 , n14077 , n14078 , n14079 , n14080 , n14081 , n14082 , n14083 , n14084 , n14085 , n14086 , n14087 , n14088 , n14089 , n14090 , n14091 , n14092 , n14093 , n14094 , n14095 , n14096 , n14097 , n14098 , n14099 , n14100 , n14101 , n14102 , n14103 , n14104 , n14105 , n14106 , n14107 , n14108 , n14109 , n14110 , n14111 , n14112 , n14113 , n14114 , n14115 , n14116 , n14117 , n14118 , n14119 , n14120 , n14121 , n14122 , n14123 , n14124 , n14125 , n14126 , n14127 , n14128 , n14129 , n14130 , n14131 , n14132 , n14133 , n14134 , n14135 , n14136 , n14137 , n14138 , n14139 , n14140 , n14141 , n14142 , n14143 , n14144 , n14145 , n14146 , n14147 , n14148 , n14149 , n14150 , n14151 , n14152 , n14153 , n14154 , n14155 , n14156 , n14157 , n14158 , n14159 , n14160 , n14161 , n14162 , n14163 , n14164 , n14165 , n14166 , n14167 , n14168 , n14169 , n14170 , n14171 , n14172 , n14173 , n14174 , n14175 , n14176 , n14177 , n14178 , n14179 , n14180 , n14181 , n14182 , n14183 , n14184 , n14185 , n14186 , n14187 , n14188 , n14189 , n14190 , n14191 , n14192 , n14193 , n14194 , n14195 , n14196 , n14197 , n14198 , n14199 , n14200 , n14201 , n14202 , n14203 , n14204 , n14205 , n14206 , n14207 , n14208 , n14209 , n14210 , n14211 , n14212 , n14213 , n14214 , n14215 , n14216 , n14217 , n14218 , n14219 , n14220 , n14221 , n14222 , n14223 , n14224 , n14225 , n14226 , n14227 , n14228 , n14229 , n14230 , n14231 , n14232 , n14233 , n14234 , n14235 , n14236 , n14237 , n14238 , n14239 , n14240 , n14241 , n14242 , n14243 , n14244 , n14245 , n14246 , n14247 , n14248 , n14249 , n14250 , n14251 , n14252 , n14253 , n14254 , n14255 , n14256 , n14257 , n14258 , n14259 , n14260 , n14261 , n14262 , n14263 , n14264 , n14265 , n14266 , n14267 , n14268 , n14269 , n14270 , n14271 , n14272 , n14273 , n14274 , n14275 , n14276 , n14277 , n14278 , n14279 , n14280 , n14281 , n14282 , n14283 , n14284 , n14285 , n14286 , n14287 , n14288 , n14289 , n14290 , n14291 , n14292 , n14293 , n14294 , n14295 , n14296 , n14297 , n14298 , n14299 , n14300 , n14301 , n14302 , n14303 , n14304 , n14305 , n14306 , n14307 , n14308 , n14309 , n14310 , n14311 , n14312 , n14313 , n14314 , n14315 , n14316 , n14317 , n14318 , n14319 , n14320 , n14321 , n14322 , n14323 , n14324 , n14325 , n14326 , n14327 , n14328 , n14329 , n14330 , n14331 , n14332 , n14333 , n14334 , n14335 , n14336 , n14337 , n14338 , n14339 , n14340 , n14341 , n14342 , n14343 , n14344 , n14345 , n14346 , n14347 , n14348 , n14349 , n14350 , n14351 , n14352 , n14353 , n14354 , n14355 , n14356 , n14357 , n14358 , n14359 , n14360 , n14361 , n14362 , n14363 , n14364 , n14365 , n14366 , n14367 , n14368 , n14369 , n14370 , n14371 , n14372 , n14373 , n14374 , n14375 , n14376 , n14377 , n14378 , n14379 , n14380 , n14381 , n14382 , n14383 , n14384 , n14385 , n14386 , n14387 , n14388 , n14389 , n14390 , n14391 , n14392 , n14393 , n14394 , n14395 , n14396 , n14397 , n14398 , n14399 , n14400 , n14401 , n14402 , n14403 , n14404 , n14405 , n14406 , n14407 , n14408 , n14409 , n14410 , n14411 , n14412 , n14413 , n14414 , n14415 , n14416 , n14417 , n14418 , n14419 , n14420 , n14421 , n14422 , n14423 , n14424 , n14425 , n14426 , n14427 , n14428 , n14429 , n14430 , n14431 , n14432 , n14433 , n14434 , n14435 , n14436 , n14437 , n14438 , n14439 , n14440 , n14441 , n14442 , n14443 , n14444 , n14445 , n14446 , n14447 , n14448 , n14449 , n14450 , n14451 , n14452 , n14453 , n14454 , n14455 , n14456 , n14457 , n14458 , n14459 , n14460 , n14461 , n14462 , n14463 , n14464 , n14465 , n14466 , n14467 , n14468 , n14469 , n14470 , n14471 , n14472 , n14473 , n14474 , n14475 , n14476 , n14477 , n14478 , n14479 , n14480 , n14481 , n14482 , n14483 , n14484 , n14485 , n14486 , n14487 , n14488 , n14489 , n14490 , n14491 , n14492 , n14493 , n14494 , n14495 , n14496 , n14497 , n14498 , n14499 , n14500 , n14501 , n14502 , n14503 , n14504 , n14505 , n14506 , n14507 , n14508 , n14509 , n14510 , n14511 , n14512 , n14513 , n14514 , n14515 , n14516 , n14517 , n14518 , n14519 , n14520 , n14521 , n14522 , n14523 , n14524 , n14525 , n14526 , n14527 , n14528 , n14529 , n14530 , n14531 , n14532 , n14533 , n14534 , n14535 , n14536 , n14537 , n14538 , n14539 , n14540 , n14541 , n14542 , n14543 , n14544 , n14545 , n14546 , n14547 , n14548 , n14549 , n14550 , n14551 , n14552 , n14553 , n14554 , n14555 , n14556 , n14557 , n14558 , n14559 , n14560 , n14561 , n14562 , n14563 , n14564 , n14565 , n14566 , n14567 , n14568 , n14569 , n14570 , n14571 , n14572 , n14573 , n14574 , n14575 , n14576 , n14577 , n14578 , n14579 , n14580 , n14581 , n14582 , n14583 , n14584 , n14585 , n14586 , n14587 , n14588 , n14589 , n14590 , n14591 , n14592 , n14593 , n14594 , n14595 , n14596 , n14597 , n14598 , n14599 , n14600 , n14601 , n14602 , n14603 , n14604 , n14605 , n14606 , n14607 , n14608 , n14609 , n14610 , n14611 , n14612 , n14613 , n14614 , n14615 , n14616 , n14617 , n14618 , n14619 , n14620 , n14621 , n14622 , n14623 , n14624 , n14625 , n14626 , n14627 , n14628 , n14629 , n14630 , n14631 , n14632 , n14633 , n14634 , n14635 , n14636 , n14637 , n14638 , n14639 , n14640 , n14641 , n14642 , n14643 , n14644 , n14645 , n14646 , n14647 , n14648 , n14649 , n14650 , n14651 , n14652 , n14653 , n14654 , n14655 , n14656 , n14657 , n14658 , n14659 , n14660 , n14661 , n14662 , n14663 , n14664 , n14665 , n14666 , n14667 , n14668 , n14669 , n14670 , n14671 , n14672 , n14673 , n14674 , n14675 , n14676 , n14677 , n14678 , n14679 , n14680 , n14681 , n14682 , n14683 , n14684 , n14685 , n14686 , n14687 , n14688 , n14689 , n14690 , n14691 , n14692 , n14693 , n14694 , n14695 , n14696 , n14697 , n14698 , n14699 , n14700 , n14701 , n14702 , n14703 , n14704 , n14705 , n14706 , n14707 , n14708 , n14709 , n14710 , n14711 , n14712 , n14713 , n14714 , n14715 , n14716 , n14717 , n14718 , n14719 , n14720 , n14721 , n14722 , n14723 , n14724 , n14725 , n14726 , n14727 , n14728 , n14729 , n14730 , n14731 , n14732 , n14733 , n14734 , n14735 , n14736 , n14737 , n14738 , n14739 , n14740 , n14741 , n14742 , n14743 , n14744 , n14745 , n14746 , n14747 , n14748 , n14749 , n14750 , n14751 , n14752 , n14753 , n14754 , n14755 , n14756 , n14757 , n14758 , n14759 , n14760 , n14761 , n14762 , n14763 , n14764 , n14765 , n14766 , n14767 , n14768 , n14769 , n14770 , n14771 , n14772 , n14773 , n14774 , n14775 , n14776 , n14777 , n14778 , n14779 , n14780 , n14781 , n14782 , n14783 , n14784 , n14785 , n14786 , n14787 , n14788 , n14789 , n14790 , n14791 , n14792 , n14793 , n14794 , n14795 , n14796 , n14797 , n14798 , n14799 , n14800 , n14801 , n14802 , n14803 , n14804 , n14805 , n14806 , n14807 , n14808 , n14809 , n14810 , n14811 , n14812 , n14813 , n14814 , n14815 , n14816 , n14817 , n14818 , n14819 , n14820 , n14821 , n14822 , n14823 , n14824 , n14825 , n14826 , n14827 , n14828 , n14829 , n14830 , n14831 , n14832 , n14833 , n14834 , n14835 , n14836 , n14837 , n14838 , n14839 , n14840 , n14841 , n14842 , n14843 , n14844 , n14845 , n14846 , n14847 , n14848 , n14849 , n14850 , n14851 , n14852 , n14853 , n14854 , n14855 , n14856 , n14857 , n14858 , n14859 , n14860 , n14861 , n14862 , n14863 , n14864 , n14865 , n14866 , n14867 , n14868 , n14869 , n14870 , n14871 , n14872 , n14873 , n14874 , n14875 , n14876 , n14877 , n14878 , n14879 , n14880 , n14881 , n14882 , n14883 , n14884 , n14885 , n14886 , n14887 , n14888 , n14889 , n14890 , n14891 , n14892 , n14893 , n14894 , n14895 , n14896 , n14897 , n14898 , n14899 , n14900 , n14901 , n14902 , n14903 , n14904 , n14905 , n14906 , n14907 , n14908 , n14909 , n14910 , n14911 , n14912 , n14913 , n14914 , n14915 , n14916 , n14917 , n14918 , n14919 , n14920 , n14921 , n14922 , n14923 , n14924 , n14925 , n14926 , n14927 , n14928 , n14929 , n14930 , n14931 , n14932 , n14933 , n14934 , n14935 , n14936 , n14937 , n14938 , n14939 , n14940 , n14941 , n14942 , n14943 , n14944 , n14945 , n14946 , n14947 , n14948 , n14949 , n14950 , n14951 , n14952 , n14953 , n14954 , n14955 , n14956 , n14957 , n14958 , n14959 , n14960 , n14961 , n14962 , n14963 , n14964 , n14965 , n14966 , n14967 , n14968 , n14969 , n14970 , n14971 , n14972 , n14973 , n14974 , n14975 , n14976 , n14977 , n14978 , n14979 , n14980 , n14981 , n14982 , n14983 , n14984 , n14985 , n14986 , n14987 , n14988 , n14989 , n14990 , n14991 , n14992 , n14993 , n14994 , n14995 , n14996 , n14997 , n14998 , n14999 , n15000 , n15001 , n15002 , n15003 , n15004 , n15005 , n15006 , n15007 , n15008 , n15009 , n15010 , n15011 , n15012 , n15013 , n15014 , n15015 , n15016 , n15017 , n15018 , n15019 , n15020 , n15021 , n15022 , n15023 , n15024 , n15025 , n15026 , n15027 , n15028 , n15029 , n15030 , n15031 , n15032 , n15033 , n15034 , n15035 , n15036 , n15037 , n15038 , n15039 , n15040 , n15041 , n15042 , n15043 , n15044 , n15045 , n15046 , n15047 , n15048 , n15049 , n15050 , n15051 , n15052 , n15053 , n15054 , n15055 , n15056 , n15057 , n15058 , n15059 , n15060 , n15061 , n15062 , n15063 , n15064 , n15065 , n15066 , n15067 , n15068 , n15069 , n15070 , n15071 , n15072 , n15073 , n15074 , n15075 , n15076 , n15077 , n15078 , n15079 , n15080 , n15081 , n15082 , n15083 , n15084 , n15085 , n15086 , n15087 , n15088 , n15089 , n15090 , n15091 , n15092 , n15093 , n15094 , n15095 , n15096 , n15097 , n15098 , n15099 , n15100 , n15101 , n15102 , n15103 , n15104 , n15105 , n15106 , n15107 , n15108 , n15109 , n15110 , n15111 , n15112 , n15113 , n15114 , n15115 , n15116 , n15117 , n15118 , n15119 , n15120 , n15121 , n15122 , n15123 , n15124 , n15125 , n15126 , n15127 , n15128 , n15129 , n15130 , n15131 , n15132 , n15133 , n15134 , n15135 , n15136 , n15137 , n15138 , n15139 , n15140 , n15141 , n15142 , n15143 , n15144 , n15145 , n15146 , n15147 , n15148 , n15149 , n15150 , n15151 , n15152 , n15153 , n15154 , n15155 , n15156 , n15157 , n15158 , n15159 , n15160 , n15161 , n15162 , n15163 , n15164 , n15165 , n15166 , n15167 , n15168 , n15169 , n15170 , n15171 , n15172 , n15173 , n15174 , n15175 , n15176 , n15177 , n15178 , n15179 , n15180 , n15181 , n15182 , n15183 , n15184 , n15185 , n15186 , n15187 , n15188 , n15189 , n15190 , n15191 , n15192 , n15193 , n15194 , n15195 , n15196 , n15197 , n15198 , n15199 , n15200 , n15201 , n15202 , n15203 , n15204 , n15205 , n15206 , n15207 , n15208 , n15209 , n15210 , n15211 , n15212 , n15213 , n15214 , n15215 , n15216 , n15217 , n15218 , n15219 , n15220 , n15221 , n15222 , n15223 , n15224 , n15225 , n15226 , n15227 , n15228 , n15229 , n15230 , n15231 , n15232 , n15233 , n15234 , n15235 , n15236 , n15237 , n15238 , n15239 , n15240 , n15241 , n15242 , n15243 , n15244 , n15245 , n15246 , n15247 , n15248 , n15249 , n15250 , n15251 , n15252 , n15253 , n15254 , n15255 , n15256 , n15257 , n15258 , n15259 , n15260 , n15261 , n15262 , n15263 , n15264 , n15265 , n15266 , n15267 , n15268 , n15269 , n15270 , n15271 , n15272 , n15273 , n15274 , n15275 , n15276 , n15277 , n15278 , n15279 , n15280 , n15281 , n15282 , n15283 , n15284 , n15285 , n15286 , n15287 , n15288 , n15289 , n15290 , n15291 , n15292 , n15293 , n15294 , n15295 , n15296 , n15297 , n15298 , n15299 , n15300 , n15301 , n15302 , n15303 , n15304 , n15305 , n15306 , n15307 , n15308 , n15309 , n15310 , n15311 , n15312 , n15313 , n15314 , n15315 , n15316 , n15317 , n15318 , n15319 , n15320 , n15321 , n15322 , n15323 , n15324 , n15325 , n15326 , n15327 , n15328 , n15329 , n15330 , n15331 , n15332 , n15333 , n15334 , n15335 , n15336 , n15337 , n15338 , n15339 , n15340 , n15341 , n15342 , n15343 , n15344 , n15345 , n15346 , n15347 , n15348 , n15349 , n15350 , n15351 , n15352 , n15353 , n15354 , n15355 , n15356 , n15357 , n15358 , n15359 , n15360 , n15361 , n15362 , n15363 , n15364 , n15365 , n15366 , n15367 , n15368 , n15369 , n15370 , n15371 , n15372 , n15373 , n15374 , n15375 , n15376 , n15377 , n15378 , n15379 , n15380 , n15381 , n15382 , n15383 , n15384 , n15385 , n15386 , n15387 , n15388 , n15389 , n15390 , n15391 , n15392 , n15393 , n15394 , n15395 , n15396 , n15397 , n15398 , n15399 , n15400 , n15401 , n15402 , n15403 , n15404 , n15405 , n15406 , n15407 , n15408 , n15409 , n15410 , n15411 , n15412 , n15413 , n15414 , n15415 , n15416 , n15417 , n15418 , n15419 , n15420 , n15421 , n15422 , n15423 , n15424 , n15425 , n15426 , n15427 , n15428 , n15429 , n15430 , n15431 , n15432 , n15433 , n15434 , n15435 , n15436 , n15437 , n15438 , n15439 , n15440 , n15441 , n15442 , n15443 , n15444 , n15445 , n15446 , n15447 , n15448 , n15449 , n15450 , n15451 , n15452 , n15453 , n15454 , n15455 , n15456 , n15457 , n15458 , n15459 , n15460 , n15461 , n15462 , n15463 , n15464 , n15465 , n15466 , n15467 , n15468 , n15469 , n15470 , n15471 , n15472 , n15473 , n15474 , n15475 , n15476 , n15477 , n15478 , n15479 , n15480 , n15481 , n15482 , n15483 , n15484 , n15485 , n15486 , n15487 , n15488 , n15489 , n15490 , n15491 , n15492 , n15493 , n15494 , n15495 , n15496 , n15497 , n15498 , n15499 , n15500 , n15501 , n15502 , n15503 , n15504 , n15505 , n15506 , n15507 , n15508 , n15509 , n15510 , n15511 , n15512 , n15513 , n15514 , n15515 , n15516 , n15517 , n15518 , n15519 , n15520 , n15521 , n15522 , n15523 , n15524 , n15525 , n15526 , n15527 , n15528 , n15529 , n15530 , n15531 , n15532 , n15533 , n15534 , n15535 , n15536 , n15537 , n15538 , n15539 , n15540 , n15541 , n15542 , n15543 , n15544 , n15545 , n15546 , n15547 , n15548 , n15549 , n15550 , n15551 , n15552 , n15553 , n15554 , n15555 , n15556 , n15557 , n15558 , n15559 , n15560 , n15561 , n15562 , n15563 , n15564 , n15565 , n15566 , n15567 , n15568 , n15569 , n15570 , n15571 , n15572 , n15573 , n15574 , n15575 , n15576 , n15577 , n15578 , n15579 , n15580 , n15581 , n15582 , n15583 , n15584 , n15585 , n15586 , n15587 , n15588 , n15589 , n15590 , n15591 , n15592 , n15593 , n15594 , n15595 , n15596 , n15597 , n15598 , n15599 , n15600 , n15601 , n15602 , n15603 , n15604 , n15605 , n15606 , n15607 , n15608 , n15609 , n15610 , n15611 , n15612 , n15613 , n15614 , n15615 , n15616 , n15617 , n15618 , n15619 , n15620 , n15621 , n15622 , n15623 , n15624 , n15625 , n15626 , n15627 , n15628 , n15629 , n15630 , n15631 , n15632 , n15633 , n15634 , n15635 , n15636 , n15637 , n15638 , n15639 , n15640 , n15641 , n15642 , n15643 , n15644 , n15645 , n15646 , n15647 , n15648 , n15649 , n15650 , n15651 , n15652 , n15653 , n15654 , n15655 , n15656 , n15657 , n15658 , n15659 , n15660 , n15661 , n15662 , n15663 , n15664 , n15665 , n15666 , n15667 , n15668 , n15669 , n15670 , n15671 , n15672 , n15673 , n15674 , n15675 , n15676 , n15677 , n15678 , n15679 , n15680 , n15681 , n15682 , n15683 , n15684 , n15685 , n15686 , n15687 , n15688 , n15689 , n15690 , n15691 , n15692 , n15693 , n15694 , n15695 , n15696 , n15697 , n15698 , n15699 , n15700 , n15701 , n15702 , n15703 , n15704 , n15705 , n15706 , n15707 , n15708 , n15709 , n15710 , n15711 , n15712 , n15713 , n15714 , n15715 , n15716 , n15717 , n15718 , n15719 , n15720 , n15721 , n15722 , n15723 , n15724 , n15725 , n15726 , n15727 , n15728 , n15729 , n15730 , n15731 , n15732 , n15733 , n15734 , n15735 , n15736 , n15737 , n15738 , n15739 , n15740 , n15741 , n15742 , n15743 , n15744 , n15745 , n15746 , n15747 , n15748 , n15749 , n15750 , n15751 , n15752 , n15753 , n15754 , n15755 , n15756 , n15757 , n15758 , n15759 , n15760 , n15761 , n15762 , n15763 , n15764 , n15765 , n15766 , n15767 , n15768 , n15769 , n15770 , n15771 , n15772 , n15773 , n15774 , n15775 , n15776 , n15777 , n15778 , n15779 , n15780 , n15781 , n15782 , n15783 , n15784 , n15785 , n15786 , n15787 , n15788 , n15789 , n15790 , n15791 , n15792 , n15793 , n15794 , n15795 , n15796 , n15797 , n15798 , n15799 , n15800 , n15801 , n15802 , n15803 , n15804 , n15805 , n15806 , n15807 , n15808 , n15809 , n15810 , n15811 , n15812 , n15813 , n15814 , n15815 , n15816 , n15817 , n15818 , n15819 , n15820 , n15821 , n15822 , n15823 , n15824 , n15825 , n15826 , n15827 , n15828 , n15829 , n15830 , n15831 , n15832 , n15833 , n15834 , n15835 , n15836 , n15837 , n15838 , n15839 , n15840 , n15841 , n15842 , n15843 , n15844 , n15845 , n15846 , n15847 , n15848 , n15849 , n15850 , n15851 , n15852 , n15853 , n15854 , n15855 , n15856 , n15857 , n15858 , n15859 , n15860 , n15861 , n15862 , n15863 , n15864 , n15865 , n15866 , n15867 , n15868 , n15869 , n15870 , n15871 , n15872 , n15873 , n15874 , n15875 , n15876 , n15877 , n15878 , n15879 , n15880 , n15881 , n15882 , n15883 , n15884 , n15885 , n15886 , n15887 , n15888 , n15889 , n15890 , n15891 , n15892 , n15893 , n15894 , n15895 , n15896 , n15897 , n15898 , n15899 , n15900 , n15901 , n15902 , n15903 , n15904 , n15905 , n15906 , n15907 , n15908 , n15909 , n15910 , n15911 , n15912 , n15913 , n15914 , n15915 , n15916 , n15917 , n15918 , n15919 , n15920 , n15921 , n15922 , n15923 , n15924 , n15925 , n15926 , n15927 , n15928 , n15929 , n15930 , n15931 , n15932 , n15933 , n15934 , n15935 , n15936 , n15937 , n15938 , n15939 , n15940 , n15941 , n15942 , n15943 , n15944 , n15945 , n15946 , n15947 , n15948 , n15949 , n15950 , n15951 , n15952 , n15953 , n15954 , n15955 , n15956 , n15957 , n15958 , n15959 , n15960 , n15961 , n15962 , n15963 , n15964 , n15965 , n15966 , n15967 , n15968 , n15969 , n15970 , n15971 , n15972 , n15973 , n15974 , n15975 , n15976 , n15977 , n15978 , n15979 , n15980 , n15981 , n15982 , n15983 , n15984 , n15985 , n15986 , n15987 , n15988 , n15989 , n15990 , n15991 , n15992 , n15993 , n15994 , n15995 , n15996 , n15997 , n15998 , n15999 , n16000 , n16001 , n16002 , n16003 , n16004 , n16005 , n16006 , n16007 , n16008 , n16009 , n16010 , n16011 , n16012 , n16013 , n16014 , n16015 , n16016 , n16017 , n16018 , n16019 , n16020 , n16021 , n16022 , n16023 , n16024 , n16025 , n16026 , n16027 , n16028 , n16029 , n16030 , n16031 , n16032 , n16033 , n16034 , n16035 , n16036 , n16037 , n16038 , n16039 , n16040 , n16041 , n16042 , n16043 , n16044 , n16045 , n16046 , n16047 , n16048 , n16049 , n16050 , n16051 , n16052 , n16053 , n16054 , n16055 , n16056 , n16057 , n16058 , n16059 , n16060 , n16061 , n16062 , n16063 , n16064 , n16065 , n16066 , n16067 , n16068 , n16069 , n16070 , n16071 , n16072 , n16073 , n16074 , n16075 , n16076 , n16077 , n16078 , n16079 , n16080 , n16081 , n16082 , n16083 , n16084 , n16085 , n16086 , n16087 , n16088 , n16089 , n16090 , n16091 , n16092 , n16093 , n16094 , n16095 , n16096 , n16097 , n16098 , n16099 , n16100 , n16101 , n16102 , n16103 , n16104 , n16105 , n16106 , n16107 , n16108 , n16109 , n16110 , n16111 , n16112 , n16113 , n16114 , n16115 , n16116 , n16117 , n16118 , n16119 , n16120 , n16121 , n16122 , n16123 , n16124 , n16125 , n16126 , n16127 , n16128 , n16129 , n16130 , n16131 , n16132 , n16133 , n16134 , n16135 , n16136 , n16137 , n16138 , n16139 , n16140 , n16141 , n16142 , n16143 , n16144 , n16145 , n16146 , n16147 , n16148 , n16149 , n16150 , n16151 , n16152 , n16153 , n16154 , n16155 , n16156 , n16157 , n16158 , n16159 , n16160 , n16161 , n16162 , n16163 , n16164 , n16165 , n16166 , n16167 , n16168 , n16169 , n16170 , n16171 , n16172 , n16173 , n16174 , n16175 , n16176 , n16177 , n16178 , n16179 , n16180 , n16181 , n16182 , n16183 , n16184 , n16185 , n16186 , n16187 , n16188 , n16189 , n16190 , n16191 , n16192 , n16193 , n16194 , n16195 , n16196 , n16197 , n16198 , n16199 , n16200 , n16201 , n16202 , n16203 , n16204 , n16205 , n16206 , n16207 , n16208 , n16209 , n16210 , n16211 , n16212 , n16213 , n16214 , n16215 , n16216 , n16217 , n16218 , n16219 , n16220 , n16221 , n16222 , n16223 , n16224 , n16225 , n16226 , n16227 , n16228 , n16229 , n16230 , n16231 , n16232 , n16233 , n16234 , n16235 , n16236 , n16237 , n16238 , n16239 , n16240 , n16241 , n16242 , n16243 , n16244 , n16245 , n16246 , n16247 , n16248 , n16249 , n16250 , n16251 , n16252 , n16253 , n16254 , n16255 , n16256 , n16257 , n16258 , n16259 , n16260 , n16261 , n16262 , n16263 , n16264 , n16265 , n16266 , n16267 , n16268 , n16269 , n16270 , n16271 , n16272 , n16273 , n16274 , n16275 , n16276 , n16277 , n16278 , n16279 , n16280 , n16281 , n16282 , n16283 , n16284 , n16285 , n16286 , n16287 , n16288 , n16289 , n16290 , n16291 , n16292 , n16293 , n16294 , n16295 , n16296 , n16297 , n16298 , n16299 , n16300 , n16301 , n16302 , n16303 , n16304 , n16305 , n16306 , n16307 , n16308 , n16309 , n16310 , n16311 , n16312 , n16313 , n16314 , n16315 , n16316 , n16317 , n16318 , n16319 , n16320 , n16321 , n16322 , n16323 , n16324 , n16325 , n16326 , n16327 , n16328 , n16329 , n16330 , n16331 , n16332 , n16333 , n16334 , n16335 , n16336 , n16337 , n16338 , n16339 , n16340 , n16341 , n16342 , n16343 , n16344 , n16345 , n16346 , n16347 , n16348 , n16349 , n16350 , n16351 , n16352 , n16353 , n16354 , n16355 , n16356 , n16357 , n16358 , n16359 , n16360 , n16361 , n16362 , n16363 , n16364 , n16365 , n16366 , n16367 , n16368 , n16369 , n16370 , n16371 , n16372 , n16373 , n16374 , n16375 , n16376 , n16377 , n16378 , n16379 , n16380 , n16381 , n16382 , n16383 , n16384 , n16385 , n16386 , n16387 , n16388 , n16389 , n16390 , n16391 , n16392 , n16393 , n16394 , n16395 , n16396 , n16397 , n16398 , n16399 , n16400 , n16401 , n16402 , n16403 , n16404 , n16405 , n16406 , n16407 , n16408 , n16409 , n16410 , n16411 , n16412 , n16413 , n16414 , n16415 , n16416 , n16417 , n16418 , n16419 , n16420 , n16421 , n16422 , n16423 , n16424 , n16425 , n16426 , n16427 , n16428 , n16429 , n16430 , n16431 , n16432 , n16433 , n16434 , n16435 , n16436 , n16437 , n16438 , n16439 , n16440 , n16441 , n16442 , n16443 , n16444 , n16445 , n16446 , n16447 , n16448 , n16449 , n16450 , n16451 , n16452 , n16453 , n16454 , n16455 , n16456 , n16457 , n16458 , n16459 , n16460 , n16461 , n16462 , n16463 , n16464 , n16465 , n16466 , n16467 , n16468 , n16469 , n16470 , n16471 , n16472 , n16473 , n16474 , n16475 , n16476 , n16477 , n16478 , n16479 , n16480 , n16481 , n16482 , n16483 , n16484 , n16485 , n16486 , n16487 , n16488 , n16489 , n16490 , n16491 , n16492 , n16493 , n16494 , n16495 , n16496 , n16497 , n16498 , n16499 , n16500 , n16501 , n16502 , n16503 , n16504 , n16505 , n16506 , n16507 , n16508 , n16509 , n16510 , n16511 , n16512 , n16513 , n16514 , n16515 , n16516 , n16517 , n16518 , n16519 , n16520 , n16521 , n16522 , n16523 , n16524 , n16525 , n16526 , n16527 , n16528 , n16529 , n16530 , n16531 , n16532 , n16533 , n16534 , n16535 , n16536 , n16537 , n16538 , n16539 , n16540 , n16541 , n16542 , n16543 , n16544 , n16545 , n16546 , n16547 , n16548 , n16549 , n16550 , n16551 , n16552 , n16553 , n16554 , n16555 , n16556 , n16557 , n16558 , n16559 , n16560 , n16561 , n16562 , n16563 , n16564 , n16565 , n16566 , n16567 , n16568 , n16569 , n16570 , n16571 , n16572 , n16573 , n16574 , n16575 , n16576 , n16577 , n16578 , n16579 , n16580 , n16581 , n16582 , n16583 , n16584 , n16585 , n16586 , n16587 , n16588 , n16589 , n16590 , n16591 , n16592 , n16593 , n16594 , n16595 , n16596 , n16597 , n16598 , n16599 , n16600 , n16601 , n16602 , n16603 , n16604 , n16605 , n16606 , n16607 , n16608 , n16609 , n16610 , n16611 , n16612 , n16613 , n16614 , n16615 , n16616 , n16617 , n16618 , n16619 , n16620 , n16621 , n16622 , n16623 , n16624 , n16625 , n16626 , n16627 , n16628 , n16629 , n16630 , n16631 , n16632 , n16633 , n16634 , n16635 , n16636 , n16637 , n16638 , n16639 , n16640 , n16641 , n16642 , n16643 , n16644 , n16645 , n16646 , n16647 , n16648 , n16649 , n16650 , n16651 , n16652 , n16653 , n16654 , n16655 , n16656 , n16657 , n16658 , n16659 , n16660 , n16661 , n16662 , n16663 , n16664 , n16665 , n16666 , n16667 , n16668 , n16669 , n16670 , n16671 , n16672 , n16673 , n16674 , n16675 , n16676 , n16677 , n16678 , n16679 , n16680 , n16681 , n16682 , n16683 , n16684 , n16685 , n16686 , n16687 , n16688 , n16689 , n16690 , n16691 , n16692 , n16693 , n16694 , n16695 , n16696 , n16697 , n16698 , n16699 , n16700 , n16701 , n16702 , n16703 , n16704 , n16705 , n16706 , n16707 , n16708 , n16709 , n16710 , n16711 , n16712 , n16713 , n16714 , n16715 , n16716 , n16717 , n16718 , n16719 , n16720 , n16721 , n16722 , n16723 , n16724 , n16725 , n16726 , n16727 , n16728 , n16729 , n16730 , n16731 , n16732 , n16733 , n16734 , n16735 , n16736 , n16737 , n16738 , n16739 , n16740 , n16741 , n16742 , n16743 , n16744 , n16745 , n16746 , n16747 , n16748 , n16749 , n16750 , n16751 , n16752 , n16753 , n16754 , n16755 , n16756 , n16757 , n16758 , n16759 , n16760 , n16761 , n16762 , n16763 , n16764 , n16765 , n16766 , n16767 , n16768 , n16769 , n16770 , n16771 , n16772 , n16773 , n16774 , n16775 , n16776 , n16777 , n16778 , n16779 , n16780 , n16781 , n16782 , n16783 , n16784 , n16785 , n16786 , n16787 , n16788 , n16789 , n16790 , n16791 , n16792 , n16793 , n16794 , n16795 , n16796 , n16797 , n16798 , n16799 , n16800 , n16801 , n16802 , n16803 , n16804 , n16805 , n16806 , n16807 , n16808 , n16809 , n16810 , n16811 , n16812 , n16813 , n16814 , n16815 , n16816 , n16817 , n16818 , n16819 , n16820 , n16821 , n16822 , n16823 , n16824 , n16825 , n16826 , n16827 , n16828 , n16829 , n16830 , n16831 , n16832 , n16833 , n16834 , n16835 , n16836 , n16837 , n16838 , n16839 , n16840 , n16841 , n16842 , n16843 , n16844 , n16845 , n16846 , n16847 , n16848 , n16849 , n16850 , n16851 , n16852 , n16853 , n16854 , n16855 , n16856 , n16857 , n16858 , n16859 , n16860 , n16861 , n16862 , n16863 , n16864 , n16865 , n16866 , n16867 , n16868 , n16869 , n16870 , n16871 , n16872 , n16873 , n16874 , n16875 , n16876 , n16877 , n16878 , n16879 , n16880 , n16881 , n16882 , n16883 , n16884 , n16885 , n16886 , n16887 , n16888 , n16889 , n16890 , n16891 , n16892 , n16893 , n16894 , n16895 , n16896 , n16897 , n16898 , n16899 , n16900 , n16901 , n16902 , n16903 , n16904 , n16905 , n16906 , n16907 , n16908 , n16909 , n16910 , n16911 , n16912 , n16913 , n16914 , n16915 , n16916 , n16917 , n16918 , n16919 , n16920 , n16921 , n16922 , n16923 , n16924 , n16925 , n16926 , n16927 , n16928 , n16929 , n16930 , n16931 , n16932 , n16933 , n16934 , n16935 , n16936 , n16937 , n16938 , n16939 , n16940 , n16941 , n16942 , n16943 , n16944 , n16945 , n16946 , n16947 , n16948 , n16949 , n16950 , n16951 , n16952 , n16953 , n16954 , n16955 , n16956 , n16957 , n16958 , n16959 , n16960 , n16961 , n16962 , n16963 , n16964 , n16965 , n16966 , n16967 , n16968 , n16969 , n16970 , n16971 , n16972 , n16973 , n16974 , n16975 , n16976 , n16977 , n16978 , n16979 , n16980 , n16981 , n16982 , n16983 , n16984 , n16985 , n16986 , n16987 , n16988 , n16989 , n16990 , n16991 , n16992 , n16993 , n16994 , n16995 , n16996 , n16997 , n16998 , n16999 , n17000 , n17001 , n17002 , n17003 , n17004 , n17005 , n17006 , n17007 , n17008 , n17009 , n17010 , n17011 , n17012 , n17013 , n17014 , n17015 , n17016 , n17017 , n17018 , n17019 , n17020 , n17021 , n17022 , n17023 , n17024 , n17025 , n17026 , n17027 , n17028 , n17029 , n17030 , n17031 , n17032 , n17033 , n17034 , n17035 , n17036 , n17037 , n17038 , n17039 , n17040 , n17041 , n17042 , n17043 , n17044 , n17045 , n17046 , n17047 , n17048 , n17049 , n17050 , n17051 , n17052 , n17053 , n17054 , n17055 , n17056 , n17057 , n17058 , n17059 , n17060 , n17061 , n17062 , n17063 , n17064 , n17065 , n17066 , n17067 , n17068 , n17069 , n17070 , n17071 , n17072 , n17073 , n17074 , n17075 , n17076 , n17077 , n17078 , n17079 , n17080 , n17081 , n17082 , n17083 , n17084 , n17085 , n17086 , n17087 , n17088 , n17089 , n17090 , n17091 , n17092 , n17093 , n17094 , n17095 , n17096 , n17097 , n17098 , n17099 , n17100 , n17101 , n17102 , n17103 , n17104 , n17105 , n17106 , n17107 , n17108 , n17109 , n17110 , n17111 , n17112 , n17113 , n17114 , n17115 , n17116 , n17117 , n17118 , n17119 , n17120 , n17121 , n17122 , n17123 , n17124 , n17125 , n17126 , n17127 , n17128 , n17129 , n17130 , n17131 , n17132 , n17133 , n17134 , n17135 , n17136 , n17137 , n17138 , n17139 , n17140 , n17141 , n17142 , n17143 , n17144 , n17145 , n17146 , n17147 , n17148 , n17149 , n17150 , n17151 , n17152 , n17153 , n17154 , n17155 , n17156 , n17157 , n17158 , n17159 , n17160 , n17161 , n17162 , n17163 , n17164 , n17165 , n17166 , n17167 , n17168 , n17169 , n17170 , n17171 , n17172 , n17173 , n17174 , n17175 , n17176 , n17177 , n17178 , n17179 , n17180 , n17181 , n17182 , n17183 , n17184 , n17185 , n17186 , n17187 , n17188 , n17189 , n17190 , n17191 , n17192 , n17193 , n17194 , n17195 , n17196 , n17197 , n17198 , n17199 , n17200 , n17201 , n17202 , n17203 , n17204 , n17205 , n17206 , n17207 , n17208 , n17209 , n17210 , n17211 , n17212 , n17213 , n17214 , n17215 , n17216 , n17217 , n17218 , n17219 , n17220 , n17221 , n17222 , n17223 , n17224 , n17225 , n17226 , n17227 , n17228 , n17229 , n17230 , n17231 , n17232 , n17233 , n17234 , n17235 , n17236 , n17237 , n17238 , n17239 , n17240 , n17241 , n17242 , n17243 , n17244 , n17245 , n17246 , n17247 , n17248 , n17249 , n17250 , n17251 , n17252 , n17253 , n17254 , n17255 , n17256 , n17257 , n17258 , n17259 , n17260 , n17261 , n17262 , n17263 , n17264 , n17265 , n17266 , n17267 , n17268 , n17269 , n17270 , n17271 , n17272 , n17273 , n17274 , n17275 , n17276 , n17277 , n17278 , n17279 , n17280 , n17281 , n17282 , n17283 , n17284 , n17285 , n17286 , n17287 , n17288 , n17289 , n17290 , n17291 , n17292 , n17293 , n17294 , n17295 , n17296 , n17297 , n17298 , n17299 , n17300 , n17301 , n17302 , n17303 , n17304 , n17305 , n17306 , n17307 , n17308 , n17309 , n17310 , n17311 , n17312 , n17313 , n17314 , n17315 , n17316 , n17317 , n17318 , n17319 , n17320 , n17321 , n17322 , n17323 , n17324 , n17325 , n17326 , n17327 , n17328 , n17329 , n17330 , n17331 , n17332 , n17333 , n17334 , n17335 , n17336 , n17337 , n17338 , n17339 , n17340 , n17341 , n17342 , n17343 , n17344 , n17345 , n17346 , n17347 , n17348 , n17349 , n17350 , n17351 , n17352 , n17353 , n17354 , n17355 , n17356 , n17357 , n17358 , n17359 , n17360 , n17361 , n17362 , n17363 , n17364 , n17365 , n17366 , n17367 , n17368 , n17369 , n17370 , n17371 , n17372 , n17373 , n17374 , n17375 , n17376 , n17377 , n17378 , n17379 , n17380 , n17381 , n17382 , n17383 , n17384 , n17385 , n17386 , n17387 , n17388 , n17389 , n17390 , n17391 , n17392 , n17393 , n17394 , n17395 , n17396 , n17397 , n17398 , n17399 , n17400 , n17401 , n17402 , n17403 , n17404 , n17405 , n17406 , n17407 , n17408 , n17409 , n17410 , n17411 , n17412 , n17413 , n17414 , n17415 , n17416 , n17417 , n17418 , n17419 , n17420 , n17421 , n17422 , n17423 , n17424 , n17425 , n17426 , n17427 , n17428 , n17429 , n17430 , n17431 , n17432 , n17433 , n17434 , n17435 , n17436 , n17437 , n17438 , n17439 , n17440 , n17441 , n17442 , n17443 , n17444 , n17445 , n17446 , n17447 , n17448 , n17449 , n17450 , n17451 , n17452 , n17453 , n17454 , n17455 , n17456 , n17457 , n17458 , n17459 , n17460 , n17461 , n17462 , n17463 , n17464 , n17465 , n17466 , n17467 , n17468 , n17469 , n17470 , n17471 , n17472 , n17473 , n17474 , n17475 , n17476 , n17477 , n17478 , n17479 , n17480 , n17481 , n17482 , n17483 , n17484 , n17485 , n17486 , n17487 , n17488 , n17489 , n17490 , n17491 , n17492 , n17493 , n17494 , n17495 , n17496 , n17497 , n17498 , n17499 , n17500 , n17501 , n17502 , n17503 , n17504 , n17505 , n17506 , n17507 , n17508 , n17509 , n17510 , n17511 , n17512 , n17513 , n17514 , n17515 , n17516 , n17517 , n17518 , n17519 , n17520 , n17521 , n17522 , n17523 , n17524 , n17525 , n17526 , n17527 , n17528 , n17529 , n17530 , n17531 , n17532 , n17533 , n17534 , n17535 , n17536 , n17537 , n17538 , n17539 , n17540 , n17541 , n17542 , n17543 , n17544 , n17545 , n17546 , n17547 , n17548 , n17549 , n17550 , n17551 , n17552 , n17553 , n17554 , n17555 , n17556 , n17557 , n17558 , n17559 , n17560 , n17561 , n17562 , n17563 , n17564 , n17565 , n17566 , n17567 , n17568 , n17569 , n17570 , n17571 , n17572 , n17573 , n17574 , n17575 , n17576 , n17577 , n17578 , n17579 , n17580 , n17581 , n17582 , n17583 , n17584 , n17585 , n17586 , n17587 , n17588 , n17589 , n17590 , n17591 , n17592 , n17593 , n17594 , n17595 , n17596 , n17597 , n17598 , n17599 , n17600 , n17601 , n17602 , n17603 , n17604 , n17605 , n17606 , n17607 , n17608 , n17609 , n17610 , n17611 , n17612 , n17613 , n17614 , n17615 , n17616 , n17617 , n17618 , n17619 , n17620 , n17621 , n17622 , n17623 , n17624 , n17625 , n17626 , n17627 , n17628 , n17629 , n17630 , n17631 , n17632 , n17633 , n17634 , n17635 , n17636 , n17637 , n17638 , n17639 , n17640 , n17641 , n17642 , n17643 , n17644 , n17645 , n17646 , n17647 , n17648 , n17649 , n17650 , n17651 , n17652 , n17653 , n17654 , n17655 , n17656 , n17657 , n17658 , n17659 , n17660 , n17661 , n17662 , n17663 , n17664 , n17665 , n17666 , n17667 , n17668 , n17669 , n17670 , n17671 , n17672 , n17673 , n17674 , n17675 , n17676 , n17677 , n17678 , n17679 , n17680 , n17681 , n17682 , n17683 , n17684 , n17685 , n17686 , n17687 , n17688 , n17689 , n17690 , n17691 , n17692 , n17693 , n17694 , n17695 , n17696 , n17697 , n17698 , n17699 , n17700 , n17701 , n17702 , n17703 , n17704 , n17705 , n17706 , n17707 , n17708 , n17709 , n17710 , n17711 , n17712 , n17713 , n17714 , n17715 , n17716 , n17717 , n17718 , n17719 , n17720 , n17721 , n17722 , n17723 , n17724 , n17725 , n17726 , n17727 , n17728 , n17729 , n17730 , n17731 , n17732 , n17733 , n17734 , n17735 , n17736 , n17737 , n17738 , n17739 , n17740 , n17741 , n17742 , n17743 , n17744 , n17745 , n17746 , n17747 , n17748 , n17749 , n17750 , n17751 , n17752 , n17753 , n17754 , n17755 , n17756 , n17757 , n17758 , n17759 , n17760 , n17761 , n17762 , n17763 , n17764 , n17765 , n17766 , n17767 , n17768 , n17769 , n17770 , n17771 , n17772 , n17773 , n17774 , n17775 , n17776 , n17777 , n17778 , n17779 , n17780 , n17781 , n17782 , n17783 , n17784 , n17785 , n17786 , n17787 , n17788 , n17789 , n17790 , n17791 , n17792 , n17793 , n17794 , n17795 , n17796 , n17797 , n17798 , n17799 , n17800 , n17801 , n17802 , n17803 , n17804 , n17805 , n17806 , n17807 , n17808 , n17809 , n17810 , n17811 , n17812 , n17813 , n17814 , n17815 , n17816 , n17817 , n17818 , n17819 , n17820 , n17821 , n17822 , n17823 , n17824 , n17825 , n17826 , n17827 , n17828 , n17829 , n17830 , n17831 , n17832 , n17833 , n17834 , n17835 , n17836 , n17837 , n17838 , n17839 , n17840 , n17841 , n17842 , n17843 , n17844 , n17845 , n17846 , n17847 , n17848 , n17849 , n17850 , n17851 , n17852 , n17853 , n17854 , n17855 , n17856 , n17857 , n17858 , n17859 , n17860 , n17861 , n17862 , n17863 , n17864 , n17865 , n17866 , n17867 , n17868 , n17869 , n17870 , n17871 , n17872 , n17873 , n17874 , n17875 , n17876 , n17877 , n17878 , n17879 , n17880 , n17881 , n17882 , n17883 , n17884 , n17885 , n17886 , n17887 , n17888 , n17889 , n17890 , n17891 , n17892 , n17893 , n17894 , n17895 , n17896 , n17897 , n17898 , n17899 , n17900 , n17901 , n17902 , n17903 , n17904 , n17905 , n17906 , n17907 , n17908 , n17909 , n17910 , n17911 , n17912 , n17913 , n17914 , n17915 , n17916 , n17917 , n17918 , n17919 , n17920 , n17921 , n17922 , n17923 , n17924 , n17925 , n17926 , n17927 , n17928 , n17929 , n17930 , n17931 , n17932 , n17933 , n17934 , n17935 , n17936 , n17937 , n17938 , n17939 , n17940 , n17941 , n17942 , n17943 , n17944 , n17945 , n17946 , n17947 , n17948 , n17949 , n17950 , n17951 , n17952 , n17953 , n17954 , n17955 , n17956 , n17957 , n17958 , n17959 , n17960 , n17961 , n17962 , n17963 , n17964 , n17965 , n17966 , n17967 , n17968 , n17969 , n17970 , n17971 , n17972 , n17973 , n17974 , n17975 , n17976 , n17977 , n17978 , n17979 , n17980 , n17981 , n17982 , n17983 , n17984 , n17985 , n17986 , n17987 , n17988 , n17989 , n17990 , n17991 , n17992 , n17993 , n17994 , n17995 , n17996 , n17997 , n17998 , n17999 , n18000 , n18001 , n18002 , n18003 , n18004 , n18005 , n18006 , n18007 , n18008 , n18009 , n18010 , n18011 , n18012 , n18013 , n18014 , n18015 , n18016 , n18017 , n18018 , n18019 , n18020 , n18021 , n18022 , n18023 , n18024 , n18025 , n18026 , n18027 , n18028 , n18029 , n18030 , n18031 , n18032 , n18033 , n18034 , n18035 , n18036 , n18037 , n18038 , n18039 , n18040 , n18041 , n18042 , n18043 , n18044 , n18045 , n18046 , n18047 , n18048 , n18049 , n18050 , n18051 , n18052 , n18053 , n18054 , n18055 , n18056 , n18057 , n18058 , n18059 , n18060 , n18061 , n18062 , n18063 , n18064 , n18065 , n18066 , n18067 , n18068 , n18069 , n18070 , n18071 , n18072 , n18073 , n18074 , n18075 , n18076 , n18077 , n18078 , n18079 , n18080 , n18081 , n18082 , n18083 , n18084 , n18085 , n18086 , n18087 , n18088 , n18089 , n18090 , n18091 , n18092 , n18093 , n18094 , n18095 , n18096 , n18097 , n18098 , n18099 , n18100 , n18101 , n18102 , n18103 , n18104 , n18105 , n18106 , n18107 , n18108 , n18109 , n18110 , n18111 , n18112 , n18113 , n18114 , n18115 , n18116 , n18117 , n18118 , n18119 , n18120 , n18121 , n18122 , n18123 , n18124 , n18125 , n18126 , n18127 , n18128 , n18129 , n18130 , n18131 , n18132 , n18133 , n18134 , n18135 , n18136 , n18137 , n18138 , n18139 , n18140 , n18141 , n18142 , n18143 , n18144 , n18145 , n18146 , n18147 , n18148 , n18149 , n18150 , n18151 , n18152 , n18153 , n18154 , n18155 , n18156 , n18157 , n18158 , n18159 , n18160 , n18161 , n18162 , n18163 , n18164 , n18165 , n18166 , n18167 , n18168 , n18169 , n18170 , n18171 , n18172 , n18173 , n18174 , n18175 , n18176 , n18177 , n18178 , n18179 , n18180 , n18181 , n18182 , n18183 , n18184 , n18185 , n18186 , n18187 , n18188 , n18189 , n18190 , n18191 , n18192 , n18193 , n18194 , n18195 , n18196 , n18197 , n18198 , n18199 , n18200 , n18201 , n18202 , n18203 , n18204 , n18205 , n18206 , n18207 , n18208 , n18209 , n18210 , n18211 , n18212 , n18213 , n18214 , n18215 , n18216 , n18217 , n18218 , n18219 , n18220 , n18221 , n18222 , n18223 , n18224 , n18225 , n18226 , n18227 , n18228 , n18229 , n18230 , n18231 , n18232 , n18233 , n18234 , n18235 , n18236 , n18237 , n18238 , n18239 , n18240 , n18241 , n18242 , n18243 , n18244 , n18245 , n18246 , n18247 , n18248 , n18249 , n18250 , n18251 , n18252 , n18253 , n18254 , n18255 , n18256 , n18257 , n18258 , n18259 , n18260 , n18261 , n18262 , n18263 , n18264 , n18265 , n18266 , n18267 , n18268 , n18269 , n18270 , n18271 , n18272 , n18273 , n18274 , n18275 , n18276 , n18277 , n18278 , n18279 , n18280 , n18281 , n18282 , n18283 , n18284 , n18285 , n18286 , n18287 , n18288 , n18289 , n18290 , n18291 , n18292 , n18293 , n18294 , n18295 , n18296 , n18297 , n18298 , n18299 , n18300 , n18301 , n18302 , n18303 , n18304 , n18305 , n18306 , n18307 , n18308 , n18309 , n18310 , n18311 , n18312 , n18313 , n18314 , n18315 , n18316 , n18317 , n18318 , n18319 , n18320 , n18321 , n18322 , n18323 , n18324 , n18325 , n18326 , n18327 , n18328 , n18329 , n18330 , n18331 , n18332 , n18333 , n18334 , n18335 , n18336 , n18337 , n18338 , n18339 , n18340 , n18341 , n18342 , n18343 , n18344 , n18345 , n18346 , n18347 , n18348 , n18349 , n18350 , n18351 , n18352 , n18353 , n18354 , n18355 , n18356 , n18357 , n18358 , n18359 , n18360 , n18361 , n18362 , n18363 , n18364 , n18365 , n18366 , n18367 , n18368 , n18369 , n18370 , n18371 , n18372 , n18373 , n18374 , n18375 , n18376 , n18377 , n18378 , n18379 , n18380 , n18381 , n18382 , n18383 , n18384 , n18385 , n18386 , n18387 , n18388 , n18389 , n18390 , n18391 , n18392 , n18393 , n18394 , n18395 , n18396 , n18397 , n18398 , n18399 , n18400 , n18401 , n18402 , n18403 , n18404 , n18405 , n18406 , n18407 , n18408 , n18409 , n18410 , n18411 , n18412 , n18413 , n18414 , n18415 , n18416 , n18417 , n18418 , n18419 , n18420 , n18421 , n18422 , n18423 , n18424 , n18425 , n18426 , n18427 , n18428 , n18429 , n18430 , n18431 , n18432 , n18433 , n18434 , n18435 , n18436 , n18437 , n18438 , n18439 , n18440 , n18441 , n18442 , n18443 , n18444 , n18445 , n18446 , n18447 , n18448 , n18449 , n18450 , n18451 , n18452 , n18453 , n18454 , n18455 , n18456 , n18457 , n18458 , n18459 , n18460 , n18461 , n18462 , n18463 , n18464 , n18465 , n18466 , n18467 , n18468 , n18469 , n18470 , n18471 , n18472 , n18473 , n18474 , n18475 , n18476 , n18477 , n18478 , n18479 , n18480 , n18481 , n18482 , n18483 , n18484 , n18485 , n18486 , n18487 , n18488 , n18489 , n18490 , n18491 , n18492 , n18493 , n18494 , n18495 , n18496 , n18497 , n18498 , n18499 , n18500 , n18501 , n18502 , n18503 , n18504 , n18505 , n18506 , n18507 , n18508 , n18509 , n18510 , n18511 , n18512 , n18513 , n18514 , n18515 , n18516 , n18517 , n18518 , n18519 , n18520 , n18521 , n18522 , n18523 , n18524 , n18525 , n18526 , n18527 , n18528 , n18529 , n18530 , n18531 , n18532 , n18533 , n18534 , n18535 , n18536 , n18537 , n18538 , n18539 , n18540 , n18541 , n18542 , n18543 , n18544 , n18545 , n18546 , n18547 , n18548 , n18549 , n18550 , n18551 , n18552 , n18553 , n18554 , n18555 , n18556 , n18557 , n18558 , n18559 , n18560 , n18561 , n18562 , n18563 , n18564 , n18565 , n18566 , n18567 , n18568 , n18569 , n18570 , n18571 , n18572 , n18573 , n18574 , n18575 , n18576 , n18577 , n18578 , n18579 , n18580 , n18581 , n18582 , n18583 , n18584 , n18585 , n18586 , n18587 , n18588 , n18589 , n18590 , n18591 , n18592 , n18593 , n18594 , n18595 , n18596 , n18597 , n18598 , n18599 , n18600 , n18601 , n18602 , n18603 , n18604 , n18605 , n18606 , n18607 , n18608 , n18609 , n18610 , n18611 , n18612 , n18613 , n18614 , n18615 , n18616 , n18617 , n18618 , n18619 , n18620 , n18621 , n18622 , n18623 , n18624 , n18625 , n18626 , n18627 , n18628 , n18629 , n18630 , n18631 , n18632 , n18633 , n18634 , n18635 , n18636 , n18637 , n18638 , n18639 , n18640 , n18641 , n18642 , n18643 , n18644 , n18645 , n18646 , n18647 , n18648 , n18649 , n18650 , n18651 , n18652 , n18653 , n18654 , n18655 , n18656 , n18657 , n18658 , n18659 , n18660 , n18661 , n18662 , n18663 , n18664 , n18665 , n18666 , n18667 , n18668 , n18669 , n18670 , n18671 , n18672 , n18673 , n18674 , n18675 , n18676 , n18677 , n18678 , n18679 , n18680 , n18681 , n18682 , n18683 , n18684 , n18685 , n18686 , n18687 , n18688 , n18689 , n18690 , n18691 , n18692 , n18693 , n18694 , n18695 , n18696 , n18697 , n18698 , n18699 , n18700 , n18701 , n18702 , n18703 , n18704 , n18705 , n18706 , n18707 , n18708 , n18709 , n18710 , n18711 , n18712 , n18713 , n18714 , n18715 , n18716 , n18717 , n18718 , n18719 , n18720 , n18721 , n18722 , n18723 , n18724 , n18725 , n18726 , n18727 , n18728 , n18729 , n18730 , n18731 , n18732 , n18733 , n18734 , n18735 , n18736 , n18737 , n18738 , n18739 , n18740 , n18741 , n18742 , n18743 , n18744 , n18745 , n18746 , n18747 , n18748 , n18749 , n18750 , n18751 , n18752 , n18753 , n18754 , n18755 , n18756 , n18757 , n18758 , n18759 , n18760 , n18761 , n18762 , n18763 , n18764 , n18765 , n18766 , n18767 , n18768 , n18769 , n18770 , n18771 , n18772 , n18773 , n18774 , n18775 , n18776 , n18777 , n18778 , n18779 , n18780 , n18781 , n18782 , n18783 , n18784 , n18785 , n18786 , n18787 , n18788 , n18789 , n18790 , n18791 , n18792 , n18793 , n18794 , n18795 , n18796 , n18797 , n18798 , n18799 , n18800 , n18801 , n18802 , n18803 , n18804 , n18805 , n18806 , n18807 , n18808 , n18809 , n18810 , n18811 , n18812 , n18813 , n18814 , n18815 , n18816 , n18817 , n18818 , n18819 , n18820 , n18821 , n18822 , n18823 , n18824 , n18825 , n18826 , n18827 , n18828 , n18829 , n18830 , n18831 , n18832 , n18833 , n18834 , n18835 , n18836 , n18837 , n18838 , n18839 , n18840 , n18841 , n18842 , n18843 , n18844 , n18845 , n18846 , n18847 , n18848 , n18849 , n18850 , n18851 , n18852 , n18853 , n18854 , n18855 , n18856 , n18857 , n18858 , n18859 , n18860 , n18861 , n18862 , n18863 , n18864 , n18865 , n18866 , n18867 , n18868 , n18869 , n18870 , n18871 , n18872 , n18873 , n18874 , n18875 , n18876 , n18877 , n18878 , n18879 , n18880 , n18881 , n18882 , n18883 , n18884 , n18885 , n18886 , n18887 , n18888 , n18889 , n18890 , n18891 , n18892 , n18893 , n18894 , n18895 , n18896 , n18897 , n18898 , n18899 , n18900 , n18901 , n18902 , n18903 , n18904 , n18905 , n18906 , n18907 , n18908 , n18909 , n18910 , n18911 , n18912 , n18913 , n18914 , n18915 , n18916 , n18917 , n18918 , n18919 , n18920 , n18921 , n18922 , n18923 , n18924 , n18925 , n18926 , n18927 , n18928 , n18929 , n18930 , n18931 , n18932 , n18933 , n18934 , n18935 , n18936 , n18937 , n18938 , n18939 , n18940 , n18941 , n18942 , n18943 , n18944 , n18945 , n18946 , n18947 , n18948 , n18949 , n18950 , n18951 , n18952 , n18953 , n18954 , n18955 , n18956 , n18957 , n18958 , n18959 , n18960 , n18961 , n18962 , n18963 , n18964 , n18965 , n18966 , n18967 , n18968 , n18969 , n18970 , n18971 , n18972 , n18973 , n18974 , n18975 , n18976 , n18977 , n18978 , n18979 , n18980 , n18981 , n18982 , n18983 , n18984 , n18985 , n18986 , n18987 , n18988 , n18989 , n18990 , n18991 , n18992 , n18993 , n18994 , n18995 , n18996 , n18997 , n18998 , n18999 , n19000 , n19001 , n19002 , n19003 , n19004 , n19005 , n19006 , n19007 , n19008 , n19009 , n19010 , n19011 , n19012 , n19013 , n19014 , n19015 , n19016 , n19017 , n19018 , n19019 , n19020 , n19021 , n19022 , n19023 , n19024 , n19025 , n19026 , n19027 , n19028 , n19029 , n19030 , n19031 , n19032 , n19033 , n19034 , n19035 , n19036 , n19037 , n19038 , n19039 , n19040 , n19041 , n19042 , n19043 , n19044 , n19045 , n19046 , n19047 , n19048 , n19049 , n19050 , n19051 , n19052 , n19053 , n19054 , n19055 , n19056 , n19057 , n19058 , n19059 , n19060 , n19061 , n19062 , n19063 , n19064 , n19065 , n19066 , n19067 , n19068 , n19069 , n19070 , n19071 , n19072 , n19073 , n19074 , n19075 , n19076 , n19077 , n19078 , n19079 , n19080 , n19081 , n19082 , n19083 , n19084 , n19085 , n19086 , n19087 , n19088 , n19089 , n19090 , n19091 , n19092 , n19093 , n19094 , n19095 , n19096 , n19097 , n19098 , n19099 , n19100 , n19101 , n19102 , n19103 , n19104 , n19105 , n19106 , n19107 , n19108 , n19109 , n19110 , n19111 , n19112 , n19113 , n19114 , n19115 , n19116 , n19117 , n19118 , n19119 , n19120 , n19121 , n19122 , n19123 , n19124 , n19125 , n19126 , n19127 , n19128 , n19129 , n19130 , n19131 , n19132 , n19133 , n19134 , n19135 , n19136 , n19137 , n19138 , n19139 , n19140 , n19141 , n19142 , n19143 , n19144 , n19145 , n19146 , n19147 , n19148 , n19149 , n19150 , n19151 , n19152 , n19153 , n19154 , n19155 , n19156 , n19157 , n19158 , n19159 , n19160 , n19161 , n19162 , n19163 , n19164 , n19165 , n19166 , n19167 , n19168 , n19169 , n19170 , n19171 , n19172 , n19173 , n19174 , n19175 , n19176 , n19177 , n19178 , n19179 , n19180 , n19181 , n19182 , n19183 , n19184 , n19185 , n19186 , n19187 , n19188 , n19189 , n19190 , n19191 , n19192 , n19193 , n19194 , n19195 , n19196 , n19197 , n19198 , n19199 , n19200 , n19201 , n19202 , n19203 , n19204 , n19205 , n19206 , n19207 , n19208 , n19209 , n19210 , n19211 , n19212 , n19213 , n19214 , n19215 , n19216 , n19217 , n19218 , n19219 , n19220 , n19221 , n19222 , n19223 , n19224 , n19225 , n19226 , n19227 , n19228 , n19229 , n19230 , n19231 , n19232 , n19233 , n19234 , n19235 , n19236 , n19237 , n19238 , n19239 , n19240 , n19241 , n19242 , n19243 , n19244 , n19245 , n19246 , n19247 , n19248 , n19249 , n19250 , n19251 , n19252 , n19253 , n19254 , n19255 , n19256 , n19257 , n19258 , n19259 , n19260 , n19261 , n19262 , n19263 , n19264 , n19265 , n19266 , n19267 , n19268 , n19269 , n19270 , n19271 , n19272 , n19273 , n19274 , n19275 , n19276 , n19277 , n19278 , n19279 , n19280 , n19281 , n19282 , n19283 , n19284 , n19285 , n19286 , n19287 , n19288 , n19289 , n19290 , n19291 , n19292 , n19293 , n19294 , n19295 , n19296 , n19297 , n19298 , n19299 , n19300 , n19301 , n19302 , n19303 , n19304 , n19305 , n19306 , n19307 , n19308 , n19309 , n19310 , n19311 , n19312 , n19313 , n19314 , n19315 , n19316 , n19317 , n19318 , n19319 , n19320 , n19321 , n19322 , n19323 , n19324 , n19325 , n19326 , n19327 , n19328 , n19329 , n19330 , n19331 , n19332 , n19333 , n19334 , n19335 , n19336 , n19337 , n19338 , n19339 , n19340 , n19341 , n19342 , n19343 , n19344 , n19345 , n19346 , n19347 , n19348 , n19349 , n19350 , n19351 , n19352 , n19353 , n19354 , n19355 , n19356 , n19357 , n19358 , n19359 , n19360 , n19361 , n19362 , n19363 , n19364 , n19365 , n19366 , n19367 , n19368 , n19369 , n19370 , n19371 , n19372 , n19373 , n19374 , n19375 , n19376 , n19377 , n19378 , n19379 , n19380 , n19381 , n19382 , n19383 , n19384 , n19385 , n19386 , n19387 , n19388 , n19389 , n19390 , n19391 , n19392 , n19393 , n19394 , n19395 , n19396 , n19397 , n19398 , n19399 , n19400 , n19401 , n19402 , n19403 , n19404 , n19405 , n19406 , n19407 , n19408 , n19409 , n19410 , n19411 , n19412 , n19413 , n19414 , n19415 , n19416 , n19417 , n19418 , n19419 , n19420 , n19421 , n19422 , n19423 , n19424 , n19425 , n19426 , n19427 , n19428 , n19429 , n19430 , n19431 , n19432 , n19433 , n19434 , n19435 , n19436 , n19437 , n19438 , n19439 , n19440 , n19441 , n19442 , n19443 , n19444 , n19445 , n19446 , n19447 , n19448 , n19449 , n19450 , n19451 , n19452 , n19453 , n19454 , n19455 , n19456 , n19457 , n19458 , n19459 , n19460 , n19461 , n19462 , n19463 , n19464 , n19465 , n19466 , n19467 , n19468 , n19469 , n19470 , n19471 , n19472 , n19473 , n19474 , n19475 , n19476 , n19477 , n19478 , n19479 , n19480 , n19481 , n19482 , n19483 , n19484 , n19485 , n19486 , n19487 , n19488 , n19489 , n19490 , n19491 , n19492 , n19493 , n19494 , n19495 , n19496 , n19497 , n19498 , n19499 , n19500 , n19501 , n19502 , n19503 , n19504 , n19505 , n19506 , n19507 , n19508 , n19509 , n19510 , n19511 , n19512 , n19513 , n19514 , n19515 , n19516 , n19517 , n19518 , n19519 , n19520 , n19521 , n19522 , n19523 , n19524 , n19525 , n19526 , n19527 , n19528 , n19529 , n19530 , n19531 , n19532 , n19533 , n19534 , n19535 , n19536 , n19537 , n19538 , n19539 , n19540 , n19541 , n19542 , n19543 , n19544 , n19545 , n19546 , n19547 , n19548 , n19549 , n19550 , n19551 , n19552 , n19553 , n19554 , n19555 , n19556 , n19557 , n19558 , n19559 , n19560 , n19561 , n19562 , n19563 , n19564 , n19565 , n19566 , n19567 , n19568 , n19569 , n19570 , n19571 , n19572 , n19573 , n19574 , n19575 , n19576 , n19577 , n19578 , n19579 , n19580 , n19581 , n19582 , n19583 , n19584 , n19585 , n19586 , n19587 , n19588 , n19589 , n19590 , n19591 , n19592 , n19593 , n19594 , n19595 , n19596 , n19597 , n19598 , n19599 , n19600 , n19601 , n19602 , n19603 , n19604 , n19605 , n19606 , n19607 , n19608 , n19609 , n19610 , n19611 , n19612 , n19613 , n19614 , n19615 , n19616 , n19617 , n19618 , n19619 , n19620 , n19621 , n19622 , n19623 , n19624 , n19625 , n19626 , n19627 , n19628 , n19629 , n19630 , n19631 , n19632 , n19633 , n19634 , n19635 , n19636 , n19637 , n19638 , n19639 , n19640 , n19641 , n19642 , n19643 , n19644 , n19645 , n19646 , n19647 , n19648 , n19649 , n19650 , n19651 , n19652 , n19653 , n19654 , n19655 , n19656 , n19657 , n19658 , n19659 , n19660 , n19661 , n19662 , n19663 , n19664 , n19665 , n19666 , n19667 , n19668 , n19669 , n19670 , n19671 , n19672 , n19673 , n19674 , n19675 , n19676 , n19677 , n19678 , n19679 , n19680 , n19681 , n19682 , n19683 , n19684 , n19685 , n19686 , n19687 , n19688 , n19689 , n19690 , n19691 , n19692 , n19693 , n19694 , n19695 , n19696 , n19697 , n19698 , n19699 , n19700 , n19701 , n19702 , n19703 , n19704 , n19705 , n19706 , n19707 , n19708 , n19709 , n19710 , n19711 , n19712 , n19713 , n19714 , n19715 , n19716 , n19717 , n19718 , n19719 , n19720 , n19721 , n19722 , n19723 , n19724 , n19725 , n19726 , n19727 , n19728 , n19729 , n19730 , n19731 , n19732 , n19733 , n19734 , n19735 , n19736 , n19737 , n19738 , n19739 , n19740 , n19741 , n19742 , n19743 , n19744 , n19745 , n19746 , n19747 , n19748 , n19749 , n19750 , n19751 , n19752 , n19753 , n19754 , n19755 , n19756 , n19757 , n19758 , n19759 , n19760 , n19761 , n19762 , n19763 , n19764 , n19765 , n19766 , n19767 , n19768 , n19769 , n19770 , n19771 , n19772 , n19773 , n19774 , n19775 , n19776 , n19777 , n19778 , n19779 , n19780 , n19781 , n19782 , n19783 , n19784 , n19785 , n19786 , n19787 , n19788 , n19789 , n19790 , n19791 , n19792 , n19793 , n19794 , n19795 , n19796 , n19797 , n19798 , n19799 , n19800 , n19801 , n19802 , n19803 , n19804 , n19805 , n19806 , n19807 , n19808 , n19809 , n19810 , n19811 , n19812 , n19813 , n19814 , n19815 , n19816 , n19817 , n19818 , n19819 , n19820 , n19821 , n19822 , n19823 , n19824 , n19825 , n19826 , n19827 , n19828 , n19829 , n19830 , n19831 , n19832 , n19833 , n19834 , n19835 , n19836 , n19837 , n19838 , n19839 , n19840 , n19841 , n19842 , n19843 , n19844 , n19845 , n19846 , n19847 , n19848 , n19849 , n19850 , n19851 , n19852 , n19853 , n19854 , n19855 , n19856 , n19857 , n19858 , n19859 , n19860 , n19861 , n19862 , n19863 , n19864 , n19865 , n19866 , n19867 , n19868 , n19869 , n19870 , n19871 , n19872 , n19873 , n19874 , n19875 , n19876 , n19877 , n19878 , n19879 , n19880 , n19881 , n19882 , n19883 , n19884 , n19885 , n19886 , n19887 , n19888 , n19889 , n19890 , n19891 , n19892 , n19893 , n19894 , n19895 , n19896 , n19897 , n19898 , n19899 , n19900 , n19901 , n19902 , n19903 , n19904 , n19905 , n19906 , n19907 , n19908 , n19909 , n19910 , n19911 , n19912 , n19913 , n19914 , n19915 , n19916 , n19917 , n19918 , n19919 , n19920 , n19921 , n19922 , n19923 , n19924 , n19925 , n19926 , n19927 , n19928 , n19929 , n19930 , n19931 , n19932 , n19933 , n19934 , n19935 , n19936 , n19937 , n19938 , n19939 , n19940 , n19941 , n19942 , n19943 , n19944 , n19945 , n19946 , n19947 , n19948 , n19949 , n19950 , n19951 , n19952 , n19953 , n19954 , n19955 , n19956 , n19957 , n19958 , n19959 , n19960 , n19961 , n19962 , n19963 , n19964 , n19965 , n19966 , n19967 , n19968 , n19969 , n19970 , n19971 , n19972 , n19973 , n19974 , n19975 , n19976 , n19977 , n19978 , n19979 , n19980 , n19981 , n19982 , n19983 , n19984 , n19985 , n19986 , n19987 , n19988 , n19989 , n19990 , n19991 , n19992 , n19993 , n19994 , n19995 , n19996 , n19997 , n19998 , n19999 , n20000 , n20001 , n20002 , n20003 , n20004 , n20005 , n20006 , n20007 , n20008 , n20009 , n20010 , n20011 , n20012 , n20013 , n20014 , n20015 , n20016 , n20017 , n20018 , n20019 , n20020 , n20021 , n20022 , n20023 , n20024 , n20025 , n20026 , n20027 , n20028 , n20029 , n20030 , n20031 , n20032 , n20033 , n20034 , n20035 , n20036 , n20037 , n20038 , n20039 , n20040 , n20041 , n20042 , n20043 , n20044 , n20045 , n20046 , n20047 , n20048 , n20049 , n20050 , n20051 , n20052 , n20053 , n20054 , n20055 , n20056 , n20057 , n20058 , n20059 , n20060 , n20061 , n20062 , n20063 , n20064 , n20065 , n20066 , n20067 , n20068 , n20069 , n20070 , n20071 , n20072 , n20073 , n20074 , n20075 , n20076 , n20077 , n20078 , n20079 , n20080 , n20081 , n20082 , n20083 , n20084 , n20085 , n20086 , n20087 , n20088 , n20089 , n20090 , n20091 , n20092 , n20093 , n20094 , n20095 , n20096 , n20097 , n20098 , n20099 , n20100 , n20101 , n20102 , n20103 , n20104 , n20105 , n20106 , n20107 , n20108 , n20109 , n20110 , n20111 , n20112 , n20113 , n20114 , n20115 , n20116 , n20117 , n20118 , n20119 , n20120 , n20121 , n20122 , n20123 , n20124 , n20125 , n20126 , n20127 , n20128 , n20129 , n20130 , n20131 , n20132 , n20133 , n20134 , n20135 , n20136 , n20137 , n20138 , n20139 , n20140 , n20141 , n20142 , n20143 , n20144 , n20145 , n20146 , n20147 , n20148 , n20149 , n20150 , n20151 , n20152 , n20153 , n20154 , n20155 , n20156 , n20157 , n20158 , n20159 , n20160 , n20161 , n20162 , n20163 , n20164 , n20165 , n20166 , n20167 , n20168 , n20169 , n20170 , n20171 , n20172 , n20173 , n20174 , n20175 , n20176 , n20177 , n20178 , n20179 , n20180 , n20181 , n20182 , n20183 , n20184 , n20185 , n20186 , n20187 , n20188 , n20189 , n20190 , n20191 , n20192 , n20193 , n20194 , n20195 , n20196 , n20197 , n20198 , n20199 , n20200 , n20201 , n20202 , n20203 , n20204 , n20205 , n20206 , n20207 , n20208 , n20209 , n20210 , n20211 , n20212 , n20213 , n20214 , n20215 , n20216 , n20217 , n20218 , n20219 , n20220 , n20221 , n20222 , n20223 , n20224 , n20225 , n20226 , n20227 , n20228 , n20229 , n20230 , n20231 , n20232 , n20233 , n20234 , n20235 , n20236 , n20237 , n20238 , n20239 , n20240 , n20241 , n20242 , n20243 , n20244 , n20245 , n20246 , n20247 , n20248 , n20249 , n20250 , n20251 , n20252 , n20253 , n20254 , n20255 , n20256 , n20257 , n20258 , n20259 , n20260 , n20261 , n20262 , n20263 , n20264 , n20265 , n20266 , n20267 , n20268 , n20269 , n20270 , n20271 , n20272 , n20273 , n20274 , n20275 , n20276 , n20277 , n20278 , n20279 , n20280 , n20281 , n20282 , n20283 , n20284 , n20285 , n20286 , n20287 , n20288 , n20289 , n20290 , n20291 , n20292 , n20293 , n20294 , n20295 , n20296 , n20297 , n20298 , n20299 , n20300 , n20301 , n20302 , n20303 , n20304 , n20305 , n20306 , n20307 , n20308 , n20309 , n20310 , n20311 , n20312 , n20313 , n20314 , n20315 , n20316 , n20317 , n20318 , n20319 , n20320 , n20321 , n20322 , n20323 , n20324 , n20325 , n20326 , n20327 , n20328 , n20329 , n20330 , n20331 , n20332 , n20333 , n20334 , n20335 , n20336 , n20337 , n20338 , n20339 , n20340 , n20341 , n20342 , n20343 , n20344 , n20345 , n20346 , n20347 , n20348 , n20349 , n20350 , n20351 , n20352 , n20353 , n20354 , n20355 , n20356 , n20357 , n20358 , n20359 , n20360 , n20361 , n20362 , n20363 , n20364 , n20365 , n20366 , n20367 , n20368 , n20369 , n20370 , n20371 , n20372 , n20373 , n20374 , n20375 , n20376 , n20377 , n20378 , n20379 , n20380 , n20381 , n20382 , n20383 , n20384 , n20385 , n20386 , n20387 , n20388 , n20389 , n20390 , n20391 , n20392 , n20393 , n20394 , n20395 , n20396 , n20397 , n20398 , n20399 , n20400 , n20401 , n20402 , n20403 , n20404 , n20405 , n20406 , n20407 , n20408 , n20409 , n20410 , n20411 , n20412 , n20413 , n20414 , n20415 , n20416 , n20417 , n20418 , n20419 , n20420 , n20421 , n20422 , n20423 , n20424 , n20425 , n20426 , n20427 , n20428 , n20429 , n20430 , n20431 , n20432 , n20433 , n20434 , n20435 , n20436 , n20437 , n20438 , n20439 , n20440 , n20441 , n20442 , n20443 , n20444 , n20445 , n20446 , n20447 , n20448 , n20449 , n20450 , n20451 , n20452 , n20453 , n20454 , n20455 , n20456 , n20457 , n20458 , n20459 , n20460 , n20461 , n20462 , n20463 , n20464 , n20465 , n20466 , n20467 , n20468 , n20469 , n20470 , n20471 , n20472 , n20473 , n20474 , n20475 , n20476 , n20477 , n20478 , n20479 , n20480 , n20481 , n20482 , n20483 , n20484 , n20485 , n20486 , n20487 , n20488 , n20489 , n20490 , n20491 , n20492 , n20493 , n20494 , n20495 , n20496 , n20497 , n20498 , n20499 , n20500 , n20501 , n20502 , n20503 , n20504 , n20505 , n20506 , n20507 , n20508 , n20509 , n20510 , n20511 , n20512 , n20513 , n20514 , n20515 , n20516 , n20517 , n20518 , n20519 , n20520 , n20521 , n20522 , n20523 , n20524 , n20525 , n20526 , n20527 , n20528 , n20529 , n20530 , n20531 , n20532 , n20533 , n20534 , n20535 , n20536 , n20537 , n20538 , n20539 , n20540 , n20541 , n20542 , n20543 , n20544 , n20545 , n20546 , n20547 , n20548 , n20549 , n20550 , n20551 , n20552 , n20553 , n20554 , n20555 , n20556 , n20557 , n20558 , n20559 , n20560 , n20561 , n20562 , n20563 , n20564 , n20565 , n20566 , n20567 , n20568 , n20569 , n20570 , n20571 , n20572 , n20573 , n20574 , n20575 , n20576 , n20577 , n20578 , n20579 , n20580 , n20581 , n20582 , n20583 , n20584 , n20585 , n20586 , n20587 , n20588 , n20589 , n20590 , n20591 , n20592 , n20593 , n20594 , n20595 , n20596 , n20597 , n20598 , n20599 , n20600 , n20601 , n20602 , n20603 , n20604 , n20605 , n20606 , n20607 , n20608 , n20609 , n20610 , n20611 , n20612 , n20613 , n20614 , n20615 , n20616 , n20617 , n20618 , n20619 , n20620 , n20621 , n20622 , n20623 , n20624 , n20625 , n20626 , n20627 , n20628 , n20629 , n20630 , n20631 , n20632 , n20633 , n20634 , n20635 , n20636 , n20637 , n20638 , n20639 , n20640 , n20641 , n20642 , n20643 , n20644 , n20645 , n20646 , n20647 , n20648 , n20649 , n20650 , n20651 , n20652 , n20653 , n20654 , n20655 , n20656 , n20657 , n20658 , n20659 , n20660 , n20661 , n20662 , n20663 , n20664 , n20665 , n20666 , n20667 , n20668 , n20669 , n20670 , n20671 , n20672 , n20673 , n20674 , n20675 , n20676 , n20677 , n20678 , n20679 , n20680 , n20681 , n20682 , n20683 , n20684 , n20685 , n20686 , n20687 , n20688 , n20689 , n20690 , n20691 , n20692 , n20693 , n20694 , n20695 , n20696 , n20697 , n20698 , n20699 , n20700 , n20701 , n20702 , n20703 , n20704 , n20705 , n20706 , n20707 , n20708 , n20709 , n20710 , n20711 , n20712 , n20713 , n20714 , n20715 , n20716 , n20717 , n20718 , n20719 , n20720 , n20721 , n20722 , n20723 , n20724 , n20725 , n20726 , n20727 , n20728 , n20729 , n20730 , n20731 , n20732 , n20733 , n20734 , n20735 , n20736 , n20737 , n20738 , n20739 , n20740 , n20741 , n20742 , n20743 , n20744 , n20745 , n20746 , n20747 , n20748 , n20749 , n20750 , n20751 , n20752 , n20753 , n20754 , n20755 , n20756 , n20757 , n20758 , n20759 , n20760 , n20761 , n20762 , n20763 , n20764 , n20765 , n20766 , n20767 , n20768 , n20769 , n20770 , n20771 , n20772 , n20773 , n20774 , n20775 , n20776 , n20777 , n20778 , n20779 , n20780 , n20781 , n20782 , n20783 , n20784 , n20785 , n20786 , n20787 , n20788 , n20789 , n20790 , n20791 , n20792 , n20793 , n20794 , n20795 , n20796 , n20797 , n20798 , n20799 , n20800 , n20801 , n20802 , n20803 , n20804 , n20805 , n20806 , n20807 , n20808 , n20809 , n20810 , n20811 , n20812 , n20813 , n20814 , n20815 , n20816 , n20817 , n20818 , n20819 , n20820 , n20821 , n20822 , n20823 , n20824 , n20825 , n20826 , n20827 , n20828 , n20829 , n20830 , n20831 , n20832 , n20833 , n20834 , n20835 , n20836 , n20837 , n20838 , n20839 , n20840 , n20841 , n20842 , n20843 , n20844 , n20845 , n20846 , n20847 , n20848 , n20849 , n20850 , n20851 , n20852 , n20853 , n20854 , n20855 , n20856 , n20857 , n20858 , n20859 , n20860 , n20861 , n20862 , n20863 , n20864 , n20865 , n20866 , n20867 , n20868 , n20869 , n20870 , n20871 , n20872 , n20873 , n20874 , n20875 , n20876 , n20877 , n20878 , n20879 , n20880 , n20881 , n20882 , n20883 , n20884 , n20885 , n20886 , n20887 , n20888 , n20889 , n20890 , n20891 , n20892 , n20893 , n20894 , n20895 , n20896 , n20897 , n20898 , n20899 , n20900 , n20901 , n20902 , n20903 , n20904 , n20905 , n20906 , n20907 , n20908 , n20909 , n20910 , n20911 , n20912 , n20913 , n20914 , n20915 , n20916 , n20917 , n20918 , n20919 , n20920 , n20921 , n20922 , n20923 , n20924 , n20925 , n20926 , n20927 , n20928 , n20929 , n20930 , n20931 , n20932 , n20933 , n20934 , n20935 , n20936 , n20937 , n20938 , n20939 , n20940 , n20941 , n20942 , n20943 , n20944 , n20945 , n20946 , n20947 , n20948 , n20949 , n20950 , n20951 , n20952 , n20953 , n20954 , n20955 , n20956 , n20957 , n20958 , n20959 , n20960 , n20961 , n20962 , n20963 , n20964 , n20965 , n20966 , n20967 , n20968 , n20969 , n20970 , n20971 , n20972 , n20973 , n20974 , n20975 , n20976 , n20977 , n20978 , n20979 , n20980 , n20981 , n20982 , n20983 , n20984 , n20985 , n20986 , n20987 , n20988 , n20989 , n20990 , n20991 , n20992 , n20993 , n20994 , n20995 , n20996 , n20997 , n20998 , n20999 , n21000 , n21001 , n21002 , n21003 , n21004 , n21005 , n21006 , n21007 , n21008 , n21009 , n21010 , n21011 , n21012 , n21013 , n21014 , n21015 , n21016 , n21017 , n21018 , n21019 , n21020 , n21021 , n21022 , n21023 , n21024 , n21025 , n21026 , n21027 , n21028 , n21029 , n21030 , n21031 , n21032 , n21033 , n21034 , n21035 , n21036 , n21037 , n21038 , n21039 , n21040 , n21041 , n21042 , n21043 , n21044 , n21045 , n21046 , n21047 , n21048 , n21049 , n21050 , n21051 , n21052 , n21053 , n21054 , n21055 , n21056 , n21057 , n21058 , n21059 , n21060 , n21061 , n21062 , n21063 , n21064 , n21065 , n21066 , n21067 , n21068 , n21069 , n21070 , n21071 , n21072 , n21073 , n21074 , n21075 , n21076 , n21077 , n21078 , n21079 , n21080 , n21081 , n21082 , n21083 , n21084 , n21085 , n21086 , n21087 , n21088 , n21089 , n21090 , n21091 , n21092 , n21093 , n21094 , n21095 , n21096 , n21097 , n21098 , n21099 , n21100 , n21101 , n21102 , n21103 , n21104 , n21105 , n21106 , n21107 , n21108 , n21109 , n21110 , n21111 , n21112 , n21113 , n21114 , n21115 , n21116 , n21117 , n21118 , n21119 , n21120 , n21121 , n21122 , n21123 , n21124 , n21125 , n21126 , n21127 , n21128 , n21129 , n21130 , n21131 , n21132 , n21133 , n21134 , n21135 , n21136 , n21137 , n21138 , n21139 , n21140 , n21141 , n21142 , n21143 , n21144 , n21145 , n21146 , n21147 , n21148 , n21149 , n21150 , n21151 , n21152 , n21153 , n21154 , n21155 , n21156 , n21157 , n21158 , n21159 , n21160 , n21161 , n21162 , n21163 , n21164 , n21165 , n21166 , n21167 , n21168 , n21169 , n21170 , n21171 , n21172 , n21173 , n21174 , n21175 , n21176 , n21177 , n21178 , n21179 , n21180 , n21181 , n21182 , n21183 , n21184 , n21185 , n21186 , n21187 , n21188 , n21189 , n21190 , n21191 , n21192 , n21193 , n21194 , n21195 , n21196 , n21197 , n21198 , n21199 , n21200 , n21201 , n21202 , n21203 , n21204 , n21205 , n21206 , n21207 , n21208 , n21209 , n21210 , n21211 , n21212 , n21213 , n21214 , n21215 , n21216 , n21217 , n21218 , n21219 , n21220 , n21221 , n21222 , n21223 , n21224 , n21225 , n21226 , n21227 , n21228 , n21229 , n21230 , n21231 , n21232 , n21233 , n21234 , n21235 , n21236 , n21237 , n21238 , n21239 , n21240 , n21241 , n21242 , n21243 , n21244 , n21245 , n21246 , n21247 , n21248 , n21249 , n21250 , n21251 , n21252 , n21253 , n21254 , n21255 , n21256 , n21257 , n21258 , n21259 , n21260 , n21261 , n21262 , n21263 , n21264 , n21265 , n21266 , n21267 , n21268 , n21269 , n21270 , n21271 , n21272 , n21273 , n21274 , n21275 , n21276 , n21277 , n21278 , n21279 , n21280 , n21281 , n21282 , n21283 , n21284 , n21285 , n21286 , n21287 , n21288 , n21289 , n21290 , n21291 , n21292 , n21293 , n21294 , n21295 , n21296 , n21297 , n21298 , n21299 , n21300 , n21301 , n21302 , n21303 , n21304 , n21305 , n21306 , n21307 , n21308 , n21309 , n21310 , n21311 , n21312 , n21313 , n21314 , n21315 , n21316 , n21317 , n21318 , n21319 , n21320 , n21321 , n21322 , n21323 , n21324 , n21325 , n21326 , n21327 , n21328 , n21329 , n21330 , n21331 , n21332 , n21333 , n21334 , n21335 , n21336 , n21337 , n21338 , n21339 , n21340 , n21341 , n21342 , n21343 , n21344 , n21345 , n21346 , n21347 , n21348 , n21349 , n21350 , n21351 , n21352 , n21353 , n21354 , n21355 , n21356 , n21357 , n21358 , n21359 , n21360 , n21361 , n21362 , n21363 , n21364 , n21365 , n21366 , n21367 , n21368 , n21369 , n21370 , n21371 , n21372 , n21373 , n21374 , n21375 , n21376 , n21377 , n21378 , n21379 , n21380 , n21381 , n21382 , n21383 , n21384 , n21385 , n21386 , n21387 , n21388 , n21389 , n21390 , n21391 , n21392 , n21393 , n21394 , n21395 , n21396 , n21397 , n21398 , n21399 , n21400 , n21401 , n21402 , n21403 , n21404 , n21405 , n21406 , n21407 , n21408 , n21409 , n21410 , n21411 , n21412 , n21413 , n21414 , n21415 , n21416 , n21417 , n21418 , n21419 , n21420 , n21421 , n21422 , n21423 , n21424 , n21425 , n21426 , n21427 , n21428 , n21429 , n21430 , n21431 , n21432 , n21433 , n21434 , n21435 , n21436 , n21437 , n21438 , n21439 , n21440 , n21441 , n21442 , n21443 , n21444 , n21445 , n21446 , n21447 , n21448 , n21449 , n21450 , n21451 , n21452 , n21453 , n21454 , n21455 , n21456 , n21457 , n21458 , n21459 , n21460 , n21461 , n21462 , n21463 , n21464 , n21465 , n21466 , n21467 , n21468 , n21469 , n21470 , n21471 , n21472 , n21473 , n21474 , n21475 , n21476 , n21477 , n21478 , n21479 , n21480 , n21481 , n21482 , n21483 , n21484 , n21485 , n21486 , n21487 , n21488 , n21489 , n21490 , n21491 , n21492 , n21493 , n21494 , n21495 , n21496 , n21497 , n21498 , n21499 , n21500 , n21501 , n21502 , n21503 , n21504 , n21505 , n21506 , n21507 , n21508 , n21509 , n21510 , n21511 , n21512 , n21513 , n21514 , n21515 , n21516 , n21517 , n21518 , n21519 , n21520 , n21521 , n21522 , n21523 , n21524 , n21525 , n21526 , n21527 , n21528 , n21529 , n21530 , n21531 , n21532 , n21533 , n21534 , n21535 , n21536 , n21537 , n21538 , n21539 , n21540 , n21541 , n21542 , n21543 , n21544 , n21545 , n21546 , n21547 , n21548 , n21549 , n21550 , n21551 , n21552 , n21553 , n21554 , n21555 , n21556 , n21557 , n21558 , n21559 , n21560 , n21561 , n21562 , n21563 , n21564 , n21565 , n21566 , n21567 , n21568 , n21569 , n21570 , n21571 , n21572 , n21573 , n21574 , n21575 , n21576 , n21577 , n21578 , n21579 , n21580 , n21581 , n21582 , n21583 , n21584 , n21585 , n21586 , n21587 , n21588 , n21589 , n21590 , n21591 , n21592 , n21593 , n21594 , n21595 , n21596 , n21597 , n21598 , n21599 , n21600 , n21601 , n21602 , n21603 , n21604 , n21605 , n21606 , n21607 , n21608 , n21609 , n21610 , n21611 , n21612 , n21613 , n21614 , n21615 , n21616 , n21617 , n21618 , n21619 , n21620 , n21621 , n21622 , n21623 , n21624 , n21625 , n21626 , n21627 , n21628 , n21629 , n21630 , n21631 , n21632 , n21633 , n21634 , n21635 , n21636 , n21637 , n21638 , n21639 , n21640 , n21641 , n21642 , n21643 , n21644 , n21645 , n21646 , n21647 , n21648 , n21649 , n21650 , n21651 , n21652 , n21653 , n21654 , n21655 , n21656 , n21657 , n21658 , n21659 , n21660 , n21661 , n21662 , n21663 , n21664 , n21665 , n21666 , n21667 , n21668 , n21669 , n21670 , n21671 , n21672 , n21673 , n21674 , n21675 , n21676 , n21677 , n21678 , n21679 , n21680 , n21681 , n21682 , n21683 , n21684 , n21685 , n21686 , n21687 , n21688 , n21689 , n21690 , n21691 , n21692 , n21693 , n21694 , n21695 , n21696 , n21697 , n21698 , n21699 , n21700 , n21701 , n21702 , n21703 , n21704 , n21705 , n21706 , n21707 , n21708 , n21709 , n21710 , n21711 , n21712 , n21713 , n21714 , n21715 , n21716 , n21717 , n21718 , n21719 , n21720 , n21721 , n21722 , n21723 , n21724 , n21725 , n21726 , n21727 , n21728 , n21729 , n21730 , n21731 , n21732 , n21733 , n21734 , n21735 , n21736 , n21737 , n21738 , n21739 , n21740 , n21741 , n21742 , n21743 , n21744 , n21745 , n21746 , n21747 , n21748 , n21749 , n21750 , n21751 , n21752 , n21753 , n21754 , n21755 , n21756 , n21757 , n21758 , n21759 , n21760 , n21761 , n21762 , n21763 , n21764 , n21765 , n21766 , n21767 , n21768 , n21769 , n21770 , n21771 , n21772 , n21773 , n21774 , n21775 , n21776 , n21777 , n21778 , n21779 , n21780 , n21781 , n21782 , n21783 , n21784 , n21785 , n21786 , n21787 , n21788 , n21789 , n21790 , n21791 , n21792 , n21793 , n21794 , n21795 , n21796 , n21797 , n21798 , n21799 , n21800 , n21801 , n21802 , n21803 , n21804 , n21805 , n21806 , n21807 , n21808 , n21809 , n21810 , n21811 , n21812 , n21813 , n21814 , n21815 , n21816 , n21817 , n21818 , n21819 , n21820 , n21821 , n21822 , n21823 , n21824 , n21825 , n21826 , n21827 , n21828 , n21829 , n21830 , n21831 , n21832 , n21833 , n21834 , n21835 , n21836 , n21837 , n21838 , n21839 , n21840 , n21841 , n21842 , n21843 , n21844 , n21845 , n21846 , n21847 , n21848 , n21849 , n21850 , n21851 , n21852 , n21853 , n21854 , n21855 , n21856 , n21857 , n21858 , n21859 , n21860 , n21861 , n21862 , n21863 , n21864 , n21865 , n21866 , n21867 , n21868 , n21869 , n21870 , n21871 , n21872 , n21873 , n21874 , n21875 , n21876 , n21877 , n21878 , n21879 , n21880 , n21881 , n21882 , n21883 , n21884 , n21885 , n21886 , n21887 , n21888 , n21889 , n21890 , n21891 , n21892 , n21893 , n21894 , n21895 , n21896 , n21897 , n21898 , n21899 , n21900 , n21901 , n21902 , n21903 , n21904 , n21905 , n21906 , n21907 , n21908 , n21909 , n21910 , n21911 , n21912 , n21913 , n21914 , n21915 , n21916 , n21917 , n21918 , n21919 , n21920 , n21921 , n21922 , n21923 , n21924 , n21925 , n21926 , n21927 , n21928 , n21929 , n21930 , n21931 , n21932 , n21933 , n21934 , n21935 , n21936 , n21937 , n21938 , n21939 , n21940 , n21941 , n21942 , n21943 , n21944 , n21945 , n21946 , n21947 , n21948 , n21949 , n21950 , n21951 , n21952 , n21953 , n21954 , n21955 , n21956 , n21957 , n21958 , n21959 , n21960 , n21961 , n21962 , n21963 , n21964 , n21965 , n21966 , n21967 , n21968 , n21969 , n21970 , n21971 , n21972 , n21973 , n21974 , n21975 , n21976 , n21977 , n21978 , n21979 , n21980 , n21981 , n21982 , n21983 , n21984 , n21985 , n21986 , n21987 , n21988 , n21989 , n21990 , n21991 , n21992 , n21993 , n21994 , n21995 , n21996 , n21997 , n21998 , n21999 , n22000 , n22001 , n22002 , n22003 , n22004 , n22005 , n22006 , n22007 , n22008 , n22009 , n22010 , n22011 , n22012 , n22013 , n22014 , n22015 , n22016 , n22017 , n22018 , n22019 , n22020 , n22021 , n22022 , n22023 , n22024 , n22025 , n22026 , n22027 , n22028 , n22029 , n22030 , n22031 , n22032 , n22033 , n22034 , n22035 , n22036 , n22037 , n22038 , n22039 , n22040 , n22041 , n22042 , n22043 , n22044 , n22045 , n22046 , n22047 , n22048 , n22049 , n22050 , n22051 , n22052 , n22053 , n22054 , n22055 , n22056 , n22057 , n22058 , n22059 , n22060 , n22061 , n22062 , n22063 , n22064 , n22065 , n22066 , n22067 , n22068 , n22069 , n22070 , n22071 , n22072 , n22073 , n22074 , n22075 , n22076 , n22077 , n22078 , n22079 , n22080 , n22081 , n22082 , n22083 , n22084 , n22085 , n22086 , n22087 , n22088 , n22089 , n22090 , n22091 , n22092 , n22093 , n22094 , n22095 , n22096 , n22097 , n22098 , n22099 , n22100 , n22101 , n22102 , n22103 , n22104 , n22105 , n22106 , n22107 , n22108 , n22109 , n22110 , n22111 , n22112 , n22113 , n22114 , n22115 , n22116 , n22117 , n22118 , n22119 , n22120 , n22121 , n22122 , n22123 , n22124 , n22125 , n22126 , n22127 , n22128 , n22129 , n22130 , n22131 , n22132 , n22133 , n22134 , n22135 , n22136 , n22137 , n22138 , n22139 , n22140 , n22141 , n22142 , n22143 , n22144 , n22145 , n22146 , n22147 , n22148 , n22149 , n22150 , n22151 , n22152 , n22153 , n22154 , n22155 , n22156 , n22157 , n22158 , n22159 , n22160 , n22161 , n22162 , n22163 , n22164 , n22165 , n22166 , n22167 , n22168 , n22169 , n22170 , n22171 , n22172 , n22173 , n22174 , n22175 , n22176 , n22177 , n22178 , n22179 , n22180 , n22181 , n22182 , n22183 , n22184 , n22185 , n22186 , n22187 , n22188 , n22189 , n22190 , n22191 , n22192 , n22193 , n22194 , n22195 , n22196 , n22197 , n22198 , n22199 , n22200 , n22201 , n22202 , n22203 , n22204 , n22205 , n22206 , n22207 , n22208 , n22209 , n22210 , n22211 , n22212 , n22213 , n22214 , n22215 , n22216 , n22217 , n22218 , n22219 , n22220 , n22221 , n22222 , n22223 , n22224 , n22225 , n22226 , n22227 , n22228 , n22229 , n22230 , n22231 , n22232 , n22233 , n22234 , n22235 , n22236 , n22237 , n22238 , n22239 , n22240 , n22241 , n22242 , n22243 , n22244 , n22245 , n22246 , n22247 , n22248 , n22249 , n22250 , n22251 , n22252 , n22253 , n22254 , n22255 , n22256 , n22257 , n22258 , n22259 , n22260 , n22261 , n22262 , n22263 , n22264 , n22265 , n22266 , n22267 , n22268 , n22269 , n22270 , n22271 , n22272 , n22273 , n22274 , n22275 , n22276 , n22277 , n22278 , n22279 , n22280 , n22281 , n22282 , n22283 , n22284 , n22285 , n22286 , n22287 , n22288 , n22289 , n22290 , n22291 , n22292 , n22293 , n22294 , n22295 , n22296 , n22297 , n22298 , n22299 , n22300 , n22301 , n22302 , n22303 , n22304 , n22305 , n22306 , n22307 , n22308 , n22309 , n22310 , n22311 , n22312 , n22313 , n22314 , n22315 , n22316 , n22317 , n22318 , n22319 , n22320 , n22321 , n22322 , n22323 , n22324 , n22325 , n22326 , n22327 , n22328 , n22329 , n22330 , n22331 , n22332 , n22333 , n22334 , n22335 , n22336 , n22337 , n22338 , n22339 , n22340 , n22341 , n22342 , n22343 , n22344 , n22345 , n22346 , n22347 , n22348 , n22349 , n22350 , n22351 , n22352 , n22353 , n22354 , n22355 , n22356 , n22357 , n22358 , n22359 , n22360 , n22361 , n22362 , n22363 , n22364 , n22365 , n22366 , n22367 , n22368 , n22369 , n22370 , n22371 , n22372 , n22373 , n22374 , n22375 , n22376 , n22377 , n22378 , n22379 , n22380 , n22381 , n22382 , n22383 , n22384 , n22385 , n22386 , n22387 , n22388 , n22389 , n22390 , n22391 , n22392 , n22393 , n22394 , n22395 , n22396 , n22397 , n22398 , n22399 , n22400 , n22401 , n22402 , n22403 , n22404 , n22405 , n22406 , n22407 , n22408 , n22409 , n22410 , n22411 , n22412 , n22413 , n22414 , n22415 , n22416 , n22417 , n22418 , n22419 , n22420 , n22421 , n22422 , n22423 , n22424 , n22425 , n22426 , n22427 , n22428 , n22429 , n22430 , n22431 , n22432 , n22433 , n22434 , n22435 , n22436 , n22437 , n22438 , n22439 , n22440 , n22441 , n22442 , n22443 , n22444 , n22445 , n22446 , n22447 , n22448 , n22449 , n22450 , n22451 , n22452 , n22453 , n22454 , n22455 , n22456 , n22457 , n22458 , n22459 , n22460 , n22461 , n22462 , n22463 , n22464 , n22465 , n22466 , n22467 , n22468 , n22469 , n22470 , n22471 , n22472 , n22473 , n22474 , n22475 , n22476 , n22477 , n22478 , n22479 , n22480 , n22481 , n22482 , n22483 , n22484 , n22485 , n22486 , n22487 , n22488 , n22489 , n22490 , n22491 , n22492 , n22493 , n22494 , n22495 , n22496 , n22497 , n22498 , n22499 , n22500 , n22501 , n22502 , n22503 , n22504 , n22505 , n22506 , n22507 , n22508 , n22509 , n22510 , n22511 , n22512 , n22513 , n22514 , n22515 , n22516 , n22517 , n22518 , n22519 , n22520 , n22521 , n22522 , n22523 , n22524 , n22525 , n22526 , n22527 , n22528 , n22529 , n22530 , n22531 , n22532 , n22533 , n22534 , n22535 , n22536 , n22537 , n22538 , n22539 , n22540 , n22541 , n22542 , n22543 , n22544 , n22545 , n22546 , n22547 , n22548 , n22549 , n22550 , n22551 , n22552 , n22553 , n22554 , n22555 , n22556 , n22557 , n22558 , n22559 , n22560 , n22561 , n22562 , n22563 , n22564 , n22565 , n22566 , n22567 , n22568 , n22569 , n22570 , n22571 , n22572 , n22573 , n22574 , n22575 , n22576 , n22577 , n22578 , n22579 , n22580 , n22581 , n22582 , n22583 , n22584 , n22585 , n22586 , n22587 , n22588 , n22589 , n22590 , n22591 , n22592 , n22593 , n22594 , n22595 , n22596 , n22597 , n22598 , n22599 , n22600 , n22601 , n22602 , n22603 , n22604 , n22605 , n22606 , n22607 , n22608 , n22609 , n22610 , n22611 , n22612 , n22613 , n22614 , n22615 , n22616 , n22617 , n22618 , n22619 , n22620 , n22621 , n22622 , n22623 , n22624 , n22625 , n22626 , n22627 , n22628 , n22629 , n22630 , n22631 , n22632 , n22633 , n22634 , n22635 , n22636 , n22637 , n22638 , n22639 , n22640 , n22641 , n22642 , n22643 , n22644 , n22645 , n22646 , n22647 , n22648 , n22649 , n22650 , n22651 , n22652 , n22653 , n22654 , n22655 , n22656 , n22657 , n22658 , n22659 , n22660 , n22661 , n22662 , n22663 , n22664 , n22665 , n22666 , n22667 , n22668 , n22669 , n22670 , n22671 , n22672 , n22673 , n22674 , n22675 , n22676 , n22677 , n22678 , n22679 , n22680 , n22681 , n22682 , n22683 , n22684 , n22685 , n22686 , n22687 , n22688 , n22689 , n22690 , n22691 , n22692 , n22693 , n22694 , n22695 , n22696 , n22697 , n22698 , n22699 , n22700 , n22701 , n22702 , n22703 , n22704 , n22705 , n22706 , n22707 , n22708 , n22709 , n22710 , n22711 , n22712 , n22713 , n22714 , n22715 , n22716 , n22717 , n22718 , n22719 , n22720 , n22721 , n22722 , n22723 , n22724 , n22725 , n22726 , n22727 , n22728 , n22729 , n22730 , n22731 , n22732 , n22733 , n22734 , n22735 , n22736 , n22737 , n22738 , n22739 , n22740 , n22741 , n22742 , n22743 , n22744 , n22745 , n22746 , n22747 , n22748 , n22749 , n22750 , n22751 , n22752 , n22753 , n22754 , n22755 , n22756 , n22757 , n22758 , n22759 , n22760 , n22761 , n22762 , n22763 , n22764 , n22765 , n22766 , n22767 , n22768 , n22769 , n22770 , n22771 , n22772 , n22773 , n22774 , n22775 , n22776 , n22777 , n22778 , n22779 , n22780 , n22781 , n22782 , n22783 , n22784 , n22785 , n22786 , n22787 , n22788 , n22789 , n22790 , n22791 , n22792 , n22793 , n22794 , n22795 , n22796 , n22797 , n22798 , n22799 , n22800 , n22801 , n22802 , n22803 , n22804 , n22805 , n22806 , n22807 , n22808 , n22809 , n22810 , n22811 , n22812 , n22813 , n22814 , n22815 , n22816 , n22817 , n22818 , n22819 , n22820 , n22821 , n22822 , n22823 , n22824 , n22825 , n22826 , n22827 , n22828 , n22829 , n22830 , n22831 , n22832 , n22833 , n22834 , n22835 , n22836 , n22837 , n22838 , n22839 , n22840 , n22841 , n22842 , n22843 , n22844 , n22845 , n22846 , n22847 , n22848 , n22849 , n22850 , n22851 , n22852 , n22853 , n22854 , n22855 , n22856 , n22857 , n22858 , n22859 , n22860 , n22861 , n22862 , n22863 , n22864 , n22865 , n22866 , n22867 , n22868 , n22869 , n22870 , n22871 , n22872 , n22873 , n22874 , n22875 , n22876 , n22877 , n22878 , n22879 , n22880 , n22881 , n22882 , n22883 , n22884 , n22885 , n22886 , n22887 , n22888 , n22889 , n22890 , n22891 , n22892 , n22893 , n22894 , n22895 , n22896 , n22897 , n22898 , n22899 , n22900 , n22901 , n22902 , n22903 , n22904 , n22905 , n22906 , n22907 , n22908 , n22909 , n22910 , n22911 , n22912 , n22913 , n22914 , n22915 , n22916 , n22917 , n22918 , n22919 , n22920 , n22921 , n22922 , n22923 , n22924 , n22925 , n22926 , n22927 , n22928 , n22929 , n22930 , n22931 , n22932 , n22933 , n22934 , n22935 , n22936 , n22937 , n22938 , n22939 , n22940 , n22941 , n22942 , n22943 , n22944 , n22945 , n22946 , n22947 , n22948 , n22949 , n22950 , n22951 , n22952 , n22953 , n22954 , n22955 , n22956 , n22957 , n22958 , n22959 , n22960 , n22961 , n22962 , n22963 , n22964 , n22965 , n22966 , n22967 , n22968 , n22969 , n22970 , n22971 , n22972 , n22973 , n22974 , n22975 , n22976 , n22977 , n22978 , n22979 , n22980 , n22981 , n22982 , n22983 , n22984 , n22985 , n22986 , n22987 , n22988 , n22989 , n22990 , n22991 , n22992 , n22993 , n22994 , n22995 , n22996 , n22997 , n22998 , n22999 , n23000 , n23001 , n23002 , n23003 , n23004 , n23005 , n23006 , n23007 , n23008 , n23009 , n23010 , n23011 , n23012 , n23013 , n23014 , n23015 , n23016 , n23017 , n23018 , n23019 , n23020 , n23021 , n23022 , n23023 , n23024 , n23025 , n23026 , n23027 , n23028 , n23029 , n23030 , n23031 , n23032 , n23033 , n23034 , n23035 , n23036 , n23037 , n23038 , n23039 , n23040 , n23041 , n23042 , n23043 , n23044 , n23045 , n23046 , n23047 , n23048 , n23049 , n23050 , n23051 , n23052 , n23053 , n23054 , n23055 , n23056 , n23057 , n23058 , n23059 , n23060 , n23061 , n23062 , n23063 , n23064 , n23065 , n23066 , n23067 , n23068 , n23069 , n23070 , n23071 , n23072 , n23073 , n23074 , n23075 , n23076 , n23077 , n23078 , n23079 , n23080 , n23081 , n23082 , n23083 , n23084 , n23085 , n23086 , n23087 , n23088 , n23089 , n23090 , n23091 , n23092 , n23093 , n23094 , n23095 , n23096 , n23097 , n23098 , n23099 , n23100 , n23101 , n23102 , n23103 , n23104 , n23105 , n23106 , n23107 , n23108 , n23109 , n23110 , n23111 , n23112 , n23113 , n23114 , n23115 , n23116 , n23117 , n23118 , n23119 , n23120 , n23121 , n23122 , n23123 , n23124 , n23125 , n23126 , n23127 , n23128 , n23129 , n23130 , n23131 , n23132 , n23133 , n23134 , n23135 , n23136 , n23137 , n23138 , n23139 , n23140 , n23141 , n23142 , n23143 , n23144 , n23145 , n23146 , n23147 , n23148 , n23149 , n23150 , n23151 , n23152 , n23153 , n23154 , n23155 , n23156 , n23157 , n23158 , n23159 , n23160 , n23161 , n23162 , n23163 , n23164 , n23165 , n23166 , n23167 , n23168 , n23169 , n23170 , n23171 , n23172 , n23173 , n23174 , n23175 , n23176 , n23177 , n23178 , n23179 , n23180 , n23181 , n23182 , n23183 , n23184 , n23185 , n23186 , n23187 , n23188 , n23189 , n23190 , n23191 , n23192 , n23193 , n23194 , n23195 , n23196 , n23197 , n23198 , n23199 , n23200 , n23201 , n23202 , n23203 , n23204 , n23205 , n23206 , n23207 , n23208 , n23209 , n23210 , n23211 , n23212 , n23213 , n23214 , n23215 , n23216 , n23217 , n23218 , n23219 , n23220 , n23221 , n23222 , n23223 , n23224 , n23225 , n23226 , n23227 , n23228 , n23229 , n23230 , n23231 , n23232 , n23233 , n23234 , n23235 , n23236 , n23237 , n23238 , n23239 , n23240 , n23241 , n23242 , n23243 , n23244 , n23245 , n23246 , n23247 , n23248 , n23249 , n23250 , n23251 , n23252 , n23253 , n23254 , n23255 , n23256 , n23257 , n23258 , n23259 , n23260 , n23261 , n23262 , n23263 , n23264 , n23265 , n23266 , n23267 , n23268 , n23269 , n23270 , n23271 , n23272 , n23273 , n23274 , n23275 , n23276 , n23277 , n23278 , n23279 , n23280 , n23281 , n23282 , n23283 , n23284 , n23285 , n23286 , n23287 , n23288 , n23289 , n23290 , n23291 , n23292 , n23293 , n23294 , n23295 , n23296 , n23297 , n23298 , n23299 , n23300 , n23301 , n23302 , n23303 , n23304 , n23305 , n23306 , n23307 , n23308 , n23309 , n23310 , n23311 , n23312 , n23313 , n23314 , n23315 , n23316 , n23317 , n23318 , n23319 , n23320 , n23321 , n23322 , n23323 , n23324 , n23325 , n23326 , n23327 , n23328 , n23329 , n23330 , n23331 , n23332 , n23333 , n23334 , n23335 , n23336 , n23337 , n23338 , n23339 , n23340 , n23341 , n23342 , n23343 , n23344 , n23345 , n23346 , n23347 , n23348 , n23349 , n23350 , n23351 , n23352 , n23353 , n23354 , n23355 , n23356 , n23357 , n23358 , n23359 , n23360 , n23361 , n23362 , n23363 , n23364 , n23365 , n23366 , n23367 , n23368 , n23369 , n23370 , n23371 , n23372 , n23373 , n23374 , n23375 , n23376 , n23377 , n23378 , n23379 , n23380 , n23381 , n23382 , n23383 , n23384 , n23385 , n23386 , n23387 , n23388 , n23389 , n23390 , n23391 , n23392 , n23393 , n23394 , n23395 , n23396 , n23397 , n23398 , n23399 , n23400 , n23401 , n23402 , n23403 , n23404 , n23405 , n23406 , n23407 , n23408 , n23409 , n23410 , n23411 , n23412 , n23413 , n23414 , n23415 , n23416 , n23417 , n23418 , n23419 , n23420 , n23421 , n23422 , n23423 , n23424 , n23425 , n23426 , n23427 , n23428 , n23429 , n23430 , n23431 , n23432 , n23433 , n23434 , n23435 , n23436 , n23437 , n23438 , n23439 , n23440 , n23441 , n23442 , n23443 , n23444 , n23445 , n23446 , n23447 , n23448 , n23449 , n23450 , n23451 , n23452 , n23453 , n23454 , n23455 , n23456 , n23457 , n23458 , n23459 , n23460 , n23461 , n23462 , n23463 , n23464 , n23465 , n23466 , n23467 , n23468 , n23469 , n23470 , n23471 , n23472 , n23473 , n23474 , n23475 , n23476 , n23477 , n23478 , n23479 , n23480 , n23481 , n23482 , n23483 , n23484 , n23485 , n23486 , n23487 , n23488 , n23489 , n23490 , n23491 , n23492 , n23493 , n23494 , n23495 , n23496 , n23497 , n23498 , n23499 , n23500 , n23501 , n23502 , n23503 , n23504 , n23505 , n23506 , n23507 , n23508 , n23509 , n23510 , n23511 , n23512 , n23513 , n23514 , n23515 , n23516 , n23517 , n23518 , n23519 , n23520 , n23521 , n23522 , n23523 , n23524 , n23525 , n23526 , n23527 , n23528 , n23529 , n23530 , n23531 , n23532 , n23533 , n23534 , n23535 , n23536 , n23537 , n23538 , n23539 , n23540 , n23541 , n23542 , n23543 , n23544 , n23545 , n23546 , n23547 , n23548 , n23549 , n23550 , n23551 , n23552 , n23553 , n23554 , n23555 , n23556 , n23557 , n23558 , n23559 , n23560 , n23561 , n23562 , n23563 , n23564 , n23565 , n23566 , n23567 , n23568 , n23569 , n23570 , n23571 , n23572 , n23573 , n23574 , n23575 , n23576 , n23577 , n23578 , n23579 , n23580 , n23581 , n23582 , n23583 , n23584 , n23585 , n23586 , n23587 , n23588 , n23589 , n23590 , n23591 , n23592 , n23593 , n23594 , n23595 , n23596 , n23597 , n23598 , n23599 , n23600 , n23601 , n23602 , n23603 , n23604 , n23605 , n23606 , n23607 , n23608 , n23609 , n23610 , n23611 , n23612 , n23613 , n23614 , n23615 , n23616 , n23617 , n23618 , n23619 , n23620 , n23621 , n23622 , n23623 , n23624 , n23625 , n23626 , n23627 , n23628 , n23629 , n23630 , n23631 , n23632 , n23633 , n23634 , n23635 , n23636 , n23637 , n23638 , n23639 , n23640 , n23641 , n23642 , n23643 , n23644 , n23645 , n23646 , n23647 , n23648 , n23649 , n23650 , n23651 , n23652 , n23653 , n23654 , n23655 , n23656 , n23657 , n23658 , n23659 , n23660 , n23661 , n23662 , n23663 , n23664 , n23665 , n23666 , n23667 , n23668 , n23669 , n23670 , n23671 , n23672 , n23673 , n23674 , n23675 , n23676 , n23677 , n23678 , n23679 , n23680 , n23681 , n23682 , n23683 , n23684 , n23685 , n23686 , n23687 , n23688 , n23689 , n23690 , n23691 , n23692 , n23693 , n23694 , n23695 , n23696 , n23697 , n23698 , n23699 , n23700 , n23701 , n23702 , n23703 , n23704 , n23705 , n23706 , n23707 , n23708 , n23709 , n23710 , n23711 , n23712 , n23713 , n23714 , n23715 , n23716 , n23717 , n23718 , n23719 , n23720 , n23721 , n23722 , n23723 , n23724 , n23725 , n23726 , n23727 , n23728 , n23729 , n23730 , n23731 , n23732 , n23733 , n23734 , n23735 , n23736 , n23737 , n23738 , n23739 , n23740 , n23741 , n23742 , n23743 , n23744 , n23745 , n23746 , n23747 , n23748 , n23749 , n23750 , n23751 , n23752 , n23753 , n23754 , n23755 , n23756 , n23757 , n23758 , n23759 , n23760 , n23761 , n23762 , n23763 , n23764 , n23765 , n23766 , n23767 , n23768 , n23769 , n23770 , n23771 , n23772 , n23773 , n23774 , n23775 , n23776 , n23777 , n23778 , n23779 , n23780 , n23781 , n23782 , n23783 , n23784 , n23785 , n23786 , n23787 , n23788 , n23789 , n23790 , n23791 , n23792 , n23793 , n23794 , n23795 , n23796 , n23797 , n23798 , n23799 , n23800 , n23801 , n23802 , n23803 , n23804 , n23805 , n23806 , n23807 , n23808 , n23809 , n23810 , n23811 , n23812 , n23813 , n23814 , n23815 , n23816 , n23817 , n23818 , n23819 , n23820 , n23821 , n23822 , n23823 , n23824 , n23825 , n23826 , n23827 , n23828 , n23829 , n23830 , n23831 , n23832 , n23833 , n23834 , n23835 , n23836 , n23837 , n23838 , n23839 , n23840 , n23841 , n23842 , n23843 , n23844 , n23845 , n23846 , n23847 , n23848 , n23849 , n23850 , n23851 , n23852 , n23853 , n23854 , n23855 , n23856 , n23857 , n23858 , n23859 , n23860 , n23861 , n23862 , n23863 , n23864 , n23865 , n23866 , n23867 , n23868 , n23869 , n23870 , n23871 , n23872 , n23873 , n23874 , n23875 , n23876 , n23877 , n23878 , n23879 , n23880 , n23881 , n23882 , n23883 , n23884 , n23885 , n23886 , n23887 , n23888 , n23889 , n23890 , n23891 , n23892 , n23893 , n23894 , n23895 , n23896 , n23897 , n23898 , n23899 , n23900 , n23901 , n23902 , n23903 , n23904 , n23905 , n23906 , n23907 , n23908 , n23909 , n23910 , n23911 , n23912 , n23913 , n23914 , n23915 , n23916 , n23917 , n23918 , n23919 , n23920 , n23921 , n23922 , n23923 , n23924 , n23925 , n23926 , n23927 , n23928 , n23929 , n23930 , n23931 , n23932 , n23933 , n23934 , n23935 , n23936 , n23937 , n23938 , n23939 , n23940 , n23941 , n23942 , n23943 , n23944 , n23945 , n23946 , n23947 , n23948 , n23949 , n23950 , n23951 , n23952 , n23953 , n23954 , n23955 , n23956 , n23957 , n23958 , n23959 , n23960 , n23961 , n23962 , n23963 , n23964 , n23965 , n23966 , n23967 , n23968 , n23969 , n23970 , n23971 , n23972 , n23973 , n23974 , n23975 , n23976 , n23977 , n23978 , n23979 , n23980 , n23981 , n23982 , n23983 , n23984 , n23985 , n23986 , n23987 , n23988 , n23989 , n23990 , n23991 , n23992 , n23993 , n23994 , n23995 , n23996 , n23997 , n23998 , n23999 , n24000 , n24001 , n24002 , n24003 , n24004 , n24005 , n24006 , n24007 , n24008 , n24009 , n24010 , n24011 , n24012 , n24013 , n24014 , n24015 , n24016 , n24017 , n24018 , n24019 , n24020 , n24021 , n24022 , n24023 , n24024 , n24025 , n24026 , n24027 , n24028 , n24029 , n24030 , n24031 , n24032 , n24033 , n24034 , n24035 , n24036 , n24037 , n24038 , n24039 , n24040 , n24041 , n24042 , n24043 , n24044 , n24045 , n24046 , n24047 , n24048 , n24049 , n24050 , n24051 , n24052 , n24053 , n24054 , n24055 , n24056 , n24057 , n24058 , n24059 , n24060 , n24061 , n24062 , n24063 , n24064 , n24065 , n24066 , n24067 , n24068 , n24069 , n24070 , n24071 , n24072 , n24073 , n24074 , n24075 , n24076 , n24077 , n24078 , n24079 , n24080 , n24081 , n24082 , n24083 , n24084 , n24085 , n24086 , n24087 , n24088 , n24089 , n24090 , n24091 , n24092 , n24093 , n24094 , n24095 , n24096 , n24097 , n24098 , n24099 , n24100 , n24101 , n24102 , n24103 , n24104 , n24105 , n24106 , n24107 , n24108 , n24109 , n24110 , n24111 , n24112 , n24113 , n24114 , n24115 , n24116 , n24117 , n24118 , n24119 , n24120 , n24121 , n24122 , n24123 , n24124 , n24125 , n24126 , n24127 , n24128 , n24129 , n24130 , n24131 , n24132 , n24133 , n24134 , n24135 , n24136 , n24137 , n24138 , n24139 , n24140 , n24141 , n24142 , n24143 , n24144 , n24145 , n24146 , n24147 , n24148 , n24149 , n24150 , n24151 , n24152 , n24153 , n24154 , n24155 , n24156 , n24157 , n24158 , n24159 , n24160 , n24161 , n24162 , n24163 , n24164 , n24165 , n24166 , n24167 , n24168 , n24169 , n24170 , n24171 , n24172 , n24173 , n24174 , n24175 , n24176 , n24177 , n24178 , n24179 , n24180 , n24181 , n24182 , n24183 , n24184 , n24185 , n24186 , n24187 , n24188 , n24189 , n24190 , n24191 , n24192 , n24193 , n24194 , n24195 , n24196 , n24197 , n24198 , n24199 , n24200 , n24201 , n24202 , n24203 , n24204 , n24205 , n24206 , n24207 , n24208 , n24209 , n24210 , n24211 , n24212 , n24213 , n24214 , n24215 , n24216 , n24217 , n24218 , n24219 , n24220 , n24221 , n24222 , n24223 , n24224 , n24225 , n24226 , n24227 , n24228 , n24229 , n24230 , n24231 , n24232 , n24233 , n24234 , n24235 , n24236 , n24237 , n24238 , n24239 , n24240 , n24241 , n24242 , n24243 , n24244 , n24245 , n24246 , n24247 , n24248 , n24249 , n24250 , n24251 , n24252 , n24253 , n24254 , n24255 , n24256 , n24257 , n24258 , n24259 , n24260 , n24261 , n24262 , n24263 , n24264 , n24265 , n24266 , n24267 , n24268 , n24269 , n24270 , n24271 , n24272 , n24273 , n24274 , n24275 , n24276 , n24277 , n24278 , n24279 , n24280 , n24281 , n24282 , n24283 , n24284 , n24285 , n24286 , n24287 , n24288 , n24289 , n24290 , n24291 , n24292 , n24293 , n24294 , n24295 , n24296 , n24297 , n24298 , n24299 , n24300 , n24301 , n24302 , n24303 , n24304 , n24305 , n24306 , n24307 , n24308 , n24309 , n24310 , n24311 , n24312 , n24313 , n24314 , n24315 , n24316 , n24317 , n24318 , n24319 , n24320 , n24321 , n24322 , n24323 , n24324 , n24325 , n24326 , n24327 , n24328 , n24329 , n24330 , n24331 , n24332 , n24333 , n24334 , n24335 , n24336 , n24337 , n24338 , n24339 , n24340 , n24341 , n24342 , n24343 , n24344 , n24345 , n24346 , n24347 , n24348 , n24349 , n24350 , n24351 , n24352 , n24353 , n24354 , n24355 , n24356 , n24357 , n24358 , n24359 , n24360 , n24361 , n24362 , n24363 , n24364 , n24365 , n24366 , n24367 , n24368 , n24369 , n24370 , n24371 , n24372 , n24373 , n24374 , n24375 , n24376 , n24377 , n24378 , n24379 , n24380 , n24381 , n24382 , n24383 , n24384 , n24385 , n24386 , n24387 , n24388 , n24389 , n24390 , n24391 , n24392 , n24393 , n24394 , n24395 , n24396 , n24397 , n24398 , n24399 , n24400 , n24401 , n24402 , n24403 , n24404 , n24405 , n24406 , n24407 , n24408 , n24409 , n24410 , n24411 , n24412 , n24413 , n24414 , n24415 , n24416 , n24417 , n24418 , n24419 , n24420 , n24421 , n24422 , n24423 , n24424 , n24425 , n24426 , n24427 , n24428 , n24429 , n24430 , n24431 , n24432 , n24433 , n24434 , n24435 , n24436 , n24437 , n24438 , n24439 , n24440 , n24441 , n24442 , n24443 , n24444 , n24445 , n24446 , n24447 , n24448 , n24449 , n24450 , n24451 , n24452 , n24453 , n24454 , n24455 , n24456 , n24457 , n24458 , n24459 , n24460 , n24461 , n24462 , n24463 , n24464 , n24465 , n24466 , n24467 , n24468 , n24469 , n24470 , n24471 , n24472 , n24473 , n24474 , n24475 , n24476 , n24477 , n24478 , n24479 , n24480 , n24481 , n24482 , n24483 , n24484 , n24485 , n24486 , n24487 , n24488 , n24489 , n24490 , n24491 , n24492 , n24493 , n24494 , n24495 , n24496 , n24497 , n24498 , n24499 , n24500 , n24501 , n24502 , n24503 , n24504 , n24505 , n24506 , n24507 , n24508 , n24509 , n24510 , n24511 , n24512 , n24513 , n24514 , n24515 , n24516 , n24517 , n24518 , n24519 , n24520 , n24521 , n24522 , n24523 , n24524 , n24525 , n24526 , n24527 , n24528 , n24529 , n24530 , n24531 , n24532 , n24533 , n24534 , n24535 , n24536 , n24537 , n24538 , n24539 , n24540 , n24541 , n24542 , n24543 , n24544 , n24545 , n24546 , n24547 , n24548 , n24549 , n24550 , n24551 , n24552 , n24553 , n24554 , n24555 , n24556 , n24557 , n24558 , n24559 , n24560 , n24561 , n24562 , n24563 , n24564 , n24565 , n24566 , n24567 , n24568 , n24569 , n24570 , n24571 , n24572 , n24573 , n24574 , n24575 , n24576 , n24577 , n24578 , n24579 , n24580 , n24581 , n24582 , n24583 , n24584 , n24585 , n24586 , n24587 , n24588 , n24589 , n24590 , n24591 , n24592 , n24593 , n24594 , n24595 , n24596 , n24597 , n24598 , n24599 , n24600 , n24601 , n24602 , n24603 , n24604 , n24605 , n24606 , n24607 , n24608 , n24609 , n24610 , n24611 , n24612 , n24613 , n24614 , n24615 , n24616 , n24617 , n24618 , n24619 , n24620 , n24621 , n24622 , n24623 , n24624 , n24625 , n24626 , n24627 , n24628 , n24629 , n24630 , n24631 , n24632 , n24633 , n24634 , n24635 , n24636 , n24637 , n24638 , n24639 , n24640 , n24641 , n24642 , n24643 , n24644 , n24645 , n24646 , n24647 , n24648 , n24649 , n24650 , n24651 , n24652 , n24653 , n24654 , n24655 , n24656 , n24657 , n24658 , n24659 , n24660 , n24661 , n24662 , n24663 , n24664 , n24665 , n24666 , n24667 , n24668 , n24669 , n24670 , n24671 , n24672 , n24673 , n24674 , n24675 , n24676 , n24677 , n24678 , n24679 , n24680 , n24681 , n24682 , n24683 , n24684 , n24685 , n24686 , n24687 , n24688 , n24689 , n24690 , n24691 , n24692 , n24693 , n24694 , n24695 , n24696 , n24697 , n24698 , n24699 , n24700 , n24701 , n24702 , n24703 , n24704 , n24705 , n24706 , n24707 , n24708 , n24709 , n24710 , n24711 , n24712 , n24713 , n24714 , n24715 , n24716 , n24717 , n24718 , n24719 , n24720 , n24721 , n24722 , n24723 , n24724 , n24725 , n24726 , n24727 , n24728 , n24729 , n24730 , n24731 , n24732 , n24733 , n24734 , n24735 , n24736 , n24737 , n24738 , n24739 , n24740 , n24741 , n24742 , n24743 , n24744 , n24745 , n24746 , n24747 , n24748 , n24749 , n24750 , n24751 , n24752 , n24753 , n24754 , n24755 , n24756 , n24757 , n24758 , n24759 , n24760 , n24761 , n24762 , n24763 , n24764 , n24765 , n24766 , n24767 , n24768 , n24769 , n24770 , n24771 , n24772 , n24773 , n24774 , n24775 , n24776 , n24777 , n24778 , n24779 , n24780 , n24781 , n24782 , n24783 , n24784 , n24785 , n24786 , n24787 , n24788 , n24789 , n24790 , n24791 , n24792 , n24793 , n24794 , n24795 , n24796 , n24797 , n24798 , n24799 , n24800 , n24801 , n24802 , n24803 , n24804 , n24805 , n24806 , n24807 , n24808 , n24809 , n24810 , n24811 , n24812 , n24813 , n24814 , n24815 , n24816 , n24817 , n24818 , n24819 , n24820 , n24821 , n24822 , n24823 , n24824 , n24825 , n24826 , n24827 , n24828 , n24829 , n24830 , n24831 , n24832 , n24833 , n24834 , n24835 , n24836 , n24837 , n24838 , n24839 , n24840 , n24841 , n24842 , n24843 , n24844 , n24845 , n24846 , n24847 , n24848 , n24849 , n24850 , n24851 , n24852 , n24853 , n24854 , n24855 , n24856 , n24857 , n24858 , n24859 , n24860 , n24861 , n24862 , n24863 , n24864 , n24865 , n24866 , n24867 , n24868 , n24869 , n24870 , n24871 , n24872 , n24873 , n24874 , n24875 , n24876 , n24877 , n24878 , n24879 , n24880 , n24881 , n24882 , n24883 , n24884 , n24885 , n24886 , n24887 , n24888 , n24889 , n24890 , n24891 , n24892 , n24893 , n24894 , n24895 , n24896 , n24897 , n24898 , n24899 , n24900 , n24901 , n24902 , n24903 , n24904 , n24905 , n24906 , n24907 , n24908 , n24909 , n24910 , n24911 , n24912 , n24913 , n24914 , n24915 , n24916 , n24917 , n24918 , n24919 , n24920 , n24921 , n24922 , n24923 , n24924 , n24925 , n24926 , n24927 , n24928 , n24929 , n24930 , n24931 , n24932 , n24933 , n24934 , n24935 , n24936 , n24937 , n24938 , n24939 , n24940 , n24941 , n24942 , n24943 , n24944 , n24945 , n24946 , n24947 , n24948 , n24949 , n24950 , n24951 , n24952 , n24953 , n24954 , n24955 , n24956 , n24957 , n24958 , n24959 , n24960 , n24961 , n24962 , n24963 , n24964 , n24965 , n24966 , n24967 , n24968 , n24969 , n24970 , n24971 , n24972 , n24973 , n24974 , n24975 , n24976 , n24977 , n24978 , n24979 , n24980 , n24981 , n24982 , n24983 , n24984 , n24985 , n24986 , n24987 , n24988 , n24989 , n24990 , n24991 , n24992 , n24993 , n24994 , n24995 , n24996 , n24997 , n24998 , n24999 , n25000 , n25001 , n25002 , n25003 , n25004 , n25005 , n25006 , n25007 , n25008 , n25009 , n25010 , n25011 , n25012 , n25013 , n25014 , n25015 , n25016 , n25017 , n25018 , n25019 , n25020 , n25021 , n25022 , n25023 , n25024 , n25025 , n25026 , n25027 , n25028 , n25029 , n25030 , n25031 , n25032 , n25033 , n25034 , n25035 , n25036 , n25037 , n25038 , n25039 , n25040 , n25041 , n25042 , n25043 , n25044 , n25045 , n25046 , n25047 , n25048 , n25049 , n25050 , n25051 , n25052 , n25053 , n25054 , n25055 , n25056 , n25057 , n25058 , n25059 , n25060 , n25061 , n25062 , n25063 , n25064 , n25065 , n25066 , n25067 , n25068 , n25069 , n25070 , n25071 , n25072 , n25073 , n25074 , n25075 , n25076 , n25077 , n25078 , n25079 , n25080 , n25081 , n25082 , n25083 , n25084 , n25085 , n25086 , n25087 , n25088 , n25089 , n25090 , n25091 , n25092 , n25093 , n25094 , n25095 , n25096 , n25097 , n25098 , n25099 , n25100 , n25101 , n25102 , n25103 , n25104 , n25105 , n25106 , n25107 , n25108 , n25109 , n25110 , n25111 , n25112 , n25113 , n25114 , n25115 , n25116 , n25117 , n25118 , n25119 , n25120 , n25121 , n25122 , n25123 , n25124 , n25125 , n25126 , n25127 , n25128 , n25129 , n25130 , n25131 , n25132 , n25133 , n25134 , n25135 , n25136 , n25137 , n25138 , n25139 , n25140 , n25141 , n25142 , n25143 , n25144 , n25145 , n25146 , n25147 , n25148 , n25149 , n25150 , n25151 , n25152 , n25153 , n25154 , n25155 , n25156 , n25157 , n25158 , n25159 , n25160 , n25161 , n25162 , n25163 , n25164 , n25165 , n25166 , n25167 , n25168 , n25169 , n25170 , n25171 , n25172 , n25173 , n25174 , n25175 , n25176 , n25177 , n25178 , n25179 , n25180 , n25181 , n25182 , n25183 , n25184 , n25185 , n25186 , n25187 , n25188 , n25189 , n25190 , n25191 , n25192 , n25193 , n25194 , n25195 , n25196 , n25197 , n25198 , n25199 , n25200 , n25201 , n25202 , n25203 , n25204 , n25205 , n25206 , n25207 , n25208 , n25209 , n25210 , n25211 , n25212 , n25213 , n25214 , n25215 , n25216 , n25217 , n25218 , n25219 , n25220 , n25221 , n25222 , n25223 , n25224 , n25225 , n25226 , n25227 , n25228 , n25229 , n25230 , n25231 , n25232 , n25233 , n25234 , n25235 , n25236 , n25237 , n25238 , n25239 , n25240 , n25241 , n25242 , n25243 , n25244 , n25245 , n25246 , n25247 , n25248 , n25249 , n25250 , n25251 , n25252 , n25253 , n25254 , n25255 , n25256 , n25257 , n25258 , n25259 , n25260 , n25261 , n25262 , n25263 , n25264 , n25265 , n25266 , n25267 , n25268 , n25269 , n25270 , n25271 , n25272 , n25273 , n25274 , n25275 , n25276 , n25277 , n25278 , n25279 , n25280 , n25281 , n25282 , n25283 , n25284 , n25285 , n25286 , n25287 , n25288 , n25289 , n25290 , n25291 , n25292 , n25293 , n25294 , n25295 , n25296 , n25297 , n25298 , n25299 , n25300 , n25301 , n25302 , n25303 , n25304 , n25305 , n25306 , n25307 , n25308 , n25309 , n25310 , n25311 , n25312 , n25313 , n25314 , n25315 , n25316 , n25317 , n25318 , n25319 , n25320 , n25321 , n25322 , n25323 , n25324 , n25325 , n25326 , n25327 , n25328 , n25329 , n25330 , n25331 , n25332 , n25333 , n25334 , n25335 , n25336 , n25337 , n25338 , n25339 , n25340 , n25341 , n25342 , n25343 , n25344 , n25345 , n25346 , n25347 , n25348 , n25349 , n25350 , n25351 , n25352 , n25353 , n25354 , n25355 , n25356 , n25357 , n25358 , n25359 , n25360 , n25361 , n25362 , n25363 , n25364 , n25365 , n25366 , n25367 , n25368 , n25369 , n25370 , n25371 , n25372 , n25373 , n25374 , n25375 , n25376 , n25377 , n25378 , n25379 , n25380 , n25381 , n25382 , n25383 , n25384 , n25385 , n25386 , n25387 , n25388 , n25389 , n25390 , n25391 , n25392 , n25393 , n25394 , n25395 , n25396 , n25397 , n25398 , n25399 , n25400 , n25401 , n25402 , n25403 , n25404 , n25405 , n25406 , n25407 , n25408 , n25409 , n25410 , n25411 , n25412 , n25413 , n25414 , n25415 , n25416 , n25417 , n25418 , n25419 , n25420 , n25421 , n25422 , n25423 , n25424 , n25425 , n25426 , n25427 , n25428 , n25429 , n25430 , n25431 , n25432 , n25433 , n25434 , n25435 , n25436 , n25437 , n25438 , n25439 , n25440 , n25441 , n25442 , n25443 , n25444 , n25445 , n25446 , n25447 , n25448 , n25449 , n25450 , n25451 , n25452 , n25453 , n25454 , n25455 , n25456 , n25457 , n25458 , n25459 , n25460 , n25461 , n25462 , n25463 , n25464 , n25465 , n25466 , n25467 , n25468 , n25469 , n25470 , n25471 , n25472 , n25473 , n25474 , n25475 , n25476 , n25477 , n25478 , n25479 , n25480 , n25481 , n25482 , n25483 , n25484 , n25485 , n25486 , n25487 , n25488 , n25489 , n25490 , n25491 , n25492 , n25493 , n25494 , n25495 , n25496 , n25497 , n25498 , n25499 , n25500 , n25501 , n25502 , n25503 , n25504 , n25505 , n25506 , n25507 , n25508 , n25509 , n25510 , n25511 , n25512 , n25513 , n25514 , n25515 , n25516 , n25517 , n25518 , n25519 , n25520 , n25521 , n25522 , n25523 , n25524 , n25525 , n25526 , n25527 , n25528 , n25529 , n25530 , n25531 , n25532 , n25533 , n25534 , n25535 , n25536 , n25537 , n25538 , n25539 , n25540 , n25541 , n25542 , n25543 , n25544 , n25545 , n25546 , n25547 , n25548 , n25549 , n25550 , n25551 , n25552 , n25553 , n25554 , n25555 , n25556 , n25557 , n25558 , n25559 , n25560 , n25561 , n25562 , n25563 , n25564 , n25565 , n25566 , n25567 , n25568 , n25569 , n25570 , n25571 , n25572 , n25573 , n25574 , n25575 , n25576 , n25577 , n25578 , n25579 , n25580 , n25581 , n25582 , n25583 , n25584 , n25585 , n25586 , n25587 , n25588 , n25589 , n25590 , n25591 , n25592 , n25593 , n25594 , n25595 , n25596 , n25597 , n25598 , n25599 , n25600 , n25601 , n25602 , n25603 , n25604 , n25605 , n25606 , n25607 , n25608 , n25609 , n25610 , n25611 , n25612 , n25613 , n25614 , n25615 , n25616 , n25617 , n25618 , n25619 , n25620 , n25621 , n25622 , n25623 , n25624 , n25625 , n25626 , n25627 , n25628 , n25629 , n25630 , n25631 , n25632 , n25633 , n25634 , n25635 , n25636 , n25637 , n25638 , n25639 , n25640 , n25641 , n25642 , n25643 , n25644 , n25645 , n25646 , n25647 , n25648 , n25649 , n25650 , n25651 , n25652 , n25653 , n25654 , n25655 , n25656 , n25657 , n25658 , n25659 , n25660 , n25661 , n25662 , n25663 , n25664 , n25665 , n25666 , n25667 , n25668 , n25669 , n25670 , n25671 , n25672 , n25673 , n25674 , n25675 , n25676 , n25677 , n25678 , n25679 , n25680 , n25681 , n25682 , n25683 , n25684 , n25685 , n25686 , n25687 , n25688 , n25689 , n25690 , n25691 , n25692 , n25693 , n25694 , n25695 , n25696 , n25697 , n25698 , n25699 , n25700 , n25701 , n25702 , n25703 , n25704 , n25705 , n25706 , n25707 , n25708 , n25709 , n25710 , n25711 , n25712 , n25713 , n25714 , n25715 , n25716 , n25717 , n25718 , n25719 , n25720 , n25721 , n25722 , n25723 , n25724 , n25725 , n25726 , n25727 , n25728 , n25729 , n25730 , n25731 , n25732 , n25733 , n25734 , n25735 , n25736 , n25737 , n25738 , n25739 , n25740 , n25741 , n25742 , n25743 , n25744 , n25745 , n25746 , n25747 , n25748 , n25749 , n25750 , n25751 , n25752 , n25753 , n25754 , n25755 , n25756 , n25757 , n25758 , n25759 , n25760 , n25761 , n25762 , n25763 , n25764 , n25765 , n25766 , n25767 , n25768 , n25769 , n25770 , n25771 , n25772 , n25773 , n25774 , n25775 , n25776 , n25777 , n25778 , n25779 , n25780 , n25781 , n25782 , n25783 , n25784 , n25785 , n25786 , n25787 , n25788 , n25789 , n25790 , n25791 , n25792 , n25793 , n25794 , n25795 , n25796 , n25797 , n25798 , n25799 , n25800 , n25801 , n25802 , n25803 , n25804 , n25805 , n25806 , n25807 , n25808 , n25809 , n25810 , n25811 , n25812 , n25813 , n25814 , n25815 , n25816 , n25817 , n25818 , n25819 , n25820 , n25821 , n25822 , n25823 , n25824 , n25825 , n25826 , n25827 , n25828 , n25829 , n25830 , n25831 , n25832 , n25833 , n25834 , n25835 , n25836 , n25837 , n25838 , n25839 , n25840 , n25841 , n25842 , n25843 , n25844 , n25845 , n25846 , n25847 , n25848 , n25849 , n25850 , n25851 , n25852 , n25853 , n25854 , n25855 , n25856 , n25857 , n25858 , n25859 , n25860 , n25861 , n25862 , n25863 , n25864 , n25865 , n25866 , n25867 , n25868 , n25869 , n25870 , n25871 , n25872 , n25873 , n25874 , n25875 , n25876 , n25877 , n25878 , n25879 , n25880 , n25881 , n25882 , n25883 , n25884 , n25885 , n25886 , n25887 , n25888 , n25889 , n25890 , n25891 , n25892 , n25893 , n25894 , n25895 , n25896 , n25897 , n25898 , n25899 , n25900 , n25901 , n25902 , n25903 , n25904 , n25905 , n25906 , n25907 , n25908 , n25909 , n25910 , n25911 , n25912 , n25913 , n25914 , n25915 , n25916 , n25917 , n25918 , n25919 , n25920 , n25921 , n25922 , n25923 , n25924 , n25925 , n25926 , n25927 , n25928 , n25929 , n25930 , n25931 , n25932 , n25933 , n25934 , n25935 , n25936 , n25937 , n25938 , n25939 , n25940 , n25941 , n25942 , n25943 , n25944 , n25945 , n25946 , n25947 , n25948 , n25949 , n25950 , n25951 , n25952 , n25953 , n25954 , n25955 , n25956 , n25957 , n25958 , n25959 , n25960 , n25961 , n25962 , n25963 , n25964 , n25965 , n25966 , n25967 , n25968 , n25969 , n25970 , n25971 , n25972 , n25973 , n25974 , n25975 , n25976 , n25977 , n25978 , n25979 , n25980 , n25981 , n25982 , n25983 , n25984 , n25985 , n25986 , n25987 , n25988 , n25989 , n25990 , n25991 , n25992 , n25993 , n25994 , n25995 , n25996 , n25997 , n25998 , n25999 , n26000 , n26001 , n26002 , n26003 , n26004 , n26005 , n26006 , n26007 , n26008 , n26009 , n26010 , n26011 , n26012 , n26013 , n26014 , n26015 , n26016 , n26017 , n26018 , n26019 , n26020 , n26021 , n26022 , n26023 , n26024 , n26025 , n26026 , n26027 , n26028 , n26029 , n26030 , n26031 , n26032 , n26033 , n26034 , n26035 , n26036 , n26037 , n26038 , n26039 , n26040 , n26041 , n26042 , n26043 , n26044 , n26045 , n26046 , n26047 , n26048 , n26049 , n26050 , n26051 , n26052 , n26053 , n26054 , n26055 , n26056 , n26057 , n26058 , n26059 , n26060 , n26061 , n26062 , n26063 , n26064 , n26065 , n26066 , n26067 , n26068 , n26069 , n26070 , n26071 , n26072 , n26073 , n26074 , n26075 , n26076 , n26077 , n26078 , n26079 , n26080 , n26081 , n26082 , n26083 , n26084 , n26085 , n26086 , n26087 , n26088 , n26089 , n26090 , n26091 , n26092 , n26093 , n26094 , n26095 , n26096 , n26097 , n26098 , n26099 , n26100 , n26101 , n26102 , n26103 , n26104 , n26105 , n26106 , n26107 , n26108 , n26109 , n26110 , n26111 , n26112 , n26113 , n26114 , n26115 , n26116 , n26117 , n26118 , n26119 , n26120 , n26121 , n26122 , n26123 , n26124 , n26125 , n26126 , n26127 , n26128 , n26129 , n26130 , n26131 , n26132 , n26133 , n26134 , n26135 , n26136 , n26137 , n26138 , n26139 , n26140 , n26141 , n26142 , n26143 , n26144 , n26145 , n26146 , n26147 , n26148 , n26149 , n26150 , n26151 , n26152 , n26153 , n26154 , n26155 , n26156 , n26157 , n26158 , n26159 , n26160 , n26161 , n26162 , n26163 , n26164 , n26165 , n26166 , n26167 , n26168 , n26169 , n26170 , n26171 , n26172 , n26173 , n26174 , n26175 , n26176 , n26177 , n26178 , n26179 , n26180 , n26181 , n26182 , n26183 , n26184 , n26185 , n26186 , n26187 , n26188 , n26189 , n26190 , n26191 , n26192 , n26193 , n26194 , n26195 , n26196 , n26197 , n26198 , n26199 , n26200 , n26201 , n26202 , n26203 , n26204 , n26205 , n26206 , n26207 , n26208 , n26209 , n26210 , n26211 , n26212 , n26213 , n26214 , n26215 , n26216 , n26217 , n26218 , n26219 , n26220 , n26221 , n26222 , n26223 , n26224 , n26225 , n26226 , n26227 , n26228 , n26229 , n26230 , n26231 , n26232 , n26233 , n26234 , n26235 , n26236 , n26237 , n26238 , n26239 , n26240 , n26241 , n26242 , n26243 , n26244 , n26245 , n26246 , n26247 , n26248 , n26249 , n26250 , n26251 , n26252 , n26253 , n26254 , n26255 , n26256 , n26257 , n26258 , n26259 , n26260 , n26261 , n26262 , n26263 , n26264 , n26265 , n26266 , n26267 , n26268 , n26269 , n26270 , n26271 , n26272 , n26273 , n26274 , n26275 , n26276 , n26277 , n26278 , n26279 , n26280 , n26281 , n26282 , n26283 , n26284 , n26285 , n26286 , n26287 , n26288 , n26289 , n26290 , n26291 , n26292 , n26293 , n26294 , n26295 , n26296 , n26297 , n26298 , n26299 , n26300 , n26301 , n26302 , n26303 , n26304 , n26305 , n26306 , n26307 , n26308 , n26309 , n26310 , n26311 , n26312 , n26313 , n26314 , n26315 , n26316 , n26317 , n26318 , n26319 , n26320 , n26321 , n26322 , n26323 , n26324 , n26325 , n26326 , n26327 , n26328 , n26329 , n26330 , n26331 , n26332 , n26333 , n26334 , n26335 , n26336 , n26337 , n26338 , n26339 , n26340 , n26341 , n26342 , n26343 , n26344 , n26345 , n26346 , n26347 , n26348 , n26349 , n26350 , n26351 , n26352 , n26353 , n26354 , n26355 , n26356 , n26357 , n26358 , n26359 , n26360 , n26361 , n26362 , n26363 , n26364 , n26365 , n26366 , n26367 , n26368 , n26369 , n26370 , n26371 , n26372 , n26373 , n26374 , n26375 , n26376 , n26377 , n26378 , n26379 , n26380 , n26381 , n26382 , n26383 , n26384 , n26385 , n26386 , n26387 , n26388 , n26389 , n26390 , n26391 , n26392 , n26393 , n26394 , n26395 , n26396 , n26397 , n26398 , n26399 , n26400 , n26401 , n26402 , n26403 , n26404 , n26405 , n26406 , n26407 , n26408 , n26409 , n26410 , n26411 , n26412 , n26413 , n26414 , n26415 , n26416 , n26417 , n26418 , n26419 , n26420 , n26421 , n26422 , n26423 , n26424 , n26425 , n26426 , n26427 , n26428 , n26429 , n26430 , n26431 , n26432 , n26433 , n26434 , n26435 , n26436 , n26437 , n26438 , n26439 , n26440 , n26441 , n26442 , n26443 , n26444 , n26445 , n26446 , n26447 , n26448 , n26449 , n26450 , n26451 , n26452 , n26453 , n26454 , n26455 , n26456 , n26457 , n26458 , n26459 , n26460 , n26461 , n26462 , n26463 , n26464 , n26465 , n26466 , n26467 , n26468 , n26469 , n26470 , n26471 , n26472 , n26473 , n26474 , n26475 , n26476 , n26477 , n26478 , n26479 , n26480 , n26481 , n26482 , n26483 , n26484 , n26485 , n26486 , n26487 , n26488 , n26489 , n26490 , n26491 , n26492 , n26493 , n26494 , n26495 , n26496 , n26497 , n26498 , n26499 , n26500 , n26501 , n26502 , n26503 , n26504 , n26505 , n26506 , n26507 , n26508 , n26509 , n26510 , n26511 , n26512 , n26513 , n26514 , n26515 , n26516 , n26517 , n26518 , n26519 , n26520 , n26521 , n26522 , n26523 , n26524 , n26525 , n26526 , n26527 , n26528 , n26529 , n26530 , n26531 , n26532 , n26533 , n26534 , n26535 , n26536 , n26537 , n26538 , n26539 , n26540 , n26541 , n26542 , n26543 , n26544 , n26545 , n26546 , n26547 , n26548 , n26549 , n26550 , n26551 , n26552 , n26553 , n26554 , n26555 , n26556 , n26557 , n26558 , n26559 , n26560 , n26561 , n26562 , n26563 , n26564 , n26565 , n26566 , n26567 , n26568 , n26569 , n26570 , n26571 , n26572 , n26573 , n26574 , n26575 , n26576 , n26577 , n26578 , n26579 , n26580 , n26581 , n26582 , n26583 , n26584 , n26585 , n26586 , n26587 , n26588 , n26589 , n26590 , n26591 , n26592 , n26593 , n26594 , n26595 , n26596 , n26597 , n26598 , n26599 , n26600 , n26601 , n26602 , n26603 , n26604 , n26605 , n26606 , n26607 , n26608 , n26609 , n26610 , n26611 , n26612 , n26613 , n26614 , n26615 , n26616 , n26617 , n26618 , n26619 , n26620 , n26621 , n26622 , n26623 , n26624 , n26625 , n26626 , n26627 , n26628 , n26629 , n26630 , n26631 , n26632 , n26633 , n26634 , n26635 , n26636 , n26637 , n26638 , n26639 , n26640 , n26641 , n26642 , n26643 , n26644 , n26645 , n26646 , n26647 , n26648 , n26649 , n26650 , n26651 , n26652 , n26653 , n26654 , n26655 , n26656 , n26657 , n26658 , n26659 , n26660 , n26661 , n26662 , n26663 , n26664 , n26665 , n26666 , n26667 , n26668 , n26669 , n26670 , n26671 , n26672 , n26673 , n26674 , n26675 , n26676 , n26677 , n26678 , n26679 , n26680 , n26681 , n26682 , n26683 , n26684 , n26685 , n26686 , n26687 , n26688 , n26689 , n26690 , n26691 , n26692 , n26693 , n26694 , n26695 , n26696 , n26697 , n26698 , n26699 , n26700 , n26701 , n26702 , n26703 , n26704 , n26705 , n26706 , n26707 , n26708 , n26709 , n26710 , n26711 , n26712 , n26713 , n26714 , n26715 , n26716 , n26717 , n26718 , n26719 , n26720 , n26721 , n26722 , n26723 , n26724 , n26725 , n26726 , n26727 , n26728 , n26729 , n26730 , n26731 , n26732 , n26733 , n26734 , n26735 , n26736 , n26737 , n26738 , n26739 , n26740 , n26741 , n26742 , n26743 , n26744 , n26745 , n26746 , n26747 , n26748 , n26749 , n26750 , n26751 , n26752 , n26753 , n26754 , n26755 , n26756 , n26757 , n26758 , n26759 , n26760 , n26761 , n26762 , n26763 , n26764 , n26765 , n26766 , n26767 , n26768 , n26769 , n26770 , n26771 , n26772 , n26773 , n26774 , n26775 , n26776 , n26777 , n26778 , n26779 , n26780 , n26781 , n26782 , n26783 , n26784 , n26785 , n26786 , n26787 , n26788 , n26789 , n26790 , n26791 , n26792 , n26793 , n26794 , n26795 , n26796 , n26797 , n26798 , n26799 , n26800 , n26801 , n26802 , n26803 , n26804 , n26805 , n26806 , n26807 , n26808 , n26809 , n26810 , n26811 , n26812 , n26813 , n26814 , n26815 , n26816 , n26817 , n26818 , n26819 , n26820 , n26821 , n26822 , n26823 , n26824 , n26825 , n26826 , n26827 , n26828 , n26829 , n26830 , n26831 , n26832 , n26833 , n26834 , n26835 , n26836 , n26837 , n26838 , n26839 , n26840 , n26841 , n26842 , n26843 , n26844 , n26845 , n26846 , n26847 , n26848 , n26849 , n26850 , n26851 , n26852 , n26853 , n26854 , n26855 , n26856 , n26857 , n26858 , n26859 , n26860 , n26861 , n26862 , n26863 , n26864 , n26865 , n26866 , n26867 , n26868 , n26869 , n26870 , n26871 , n26872 , n26873 , n26874 , n26875 , n26876 , n26877 , n26878 , n26879 , n26880 , n26881 , n26882 , n26883 , n26884 , n26885 , n26886 , n26887 , n26888 , n26889 , n26890 , n26891 , n26892 , n26893 , n26894 , n26895 , n26896 , n26897 , n26898 , n26899 , n26900 , n26901 , n26902 , n26903 , n26904 , n26905 , n26906 , n26907 , n26908 , n26909 , n26910 , n26911 , n26912 , n26913 , n26914 , n26915 , n26916 , n26917 , n26918 , n26919 , n26920 , n26921 , n26922 , n26923 , n26924 , n26925 , n26926 , n26927 , n26928 , n26929 , n26930 , n26931 , n26932 , n26933 , n26934 , n26935 , n26936 , n26937 , n26938 , n26939 , n26940 , n26941 , n26942 , n26943 , n26944 , n26945 , n26946 , n26947 , n26948 , n26949 , n26950 , n26951 , n26952 , n26953 , n26954 , n26955 , n26956 , n26957 , n26958 , n26959 , n26960 , n26961 , n26962 , n26963 , n26964 , n26965 , n26966 , n26967 , n26968 , n26969 , n26970 , n26971 , n26972 , n26973 , n26974 , n26975 , n26976 , n26977 , n26978 , n26979 , n26980 , n26981 , n26982 , n26983 , n26984 , n26985 , n26986 , n26987 , n26988 , n26989 , n26990 , n26991 , n26992 , n26993 , n26994 , n26995 , n26996 , n26997 , n26998 , n26999 , n27000 , n27001 , n27002 , n27003 , n27004 , n27005 , n27006 , n27007 , n27008 , n27009 , n27010 , n27011 , n27012 , n27013 , n27014 , n27015 , n27016 , n27017 , n27018 , n27019 , n27020 , n27021 , n27022 , n27023 , n27024 , n27025 , n27026 , n27027 , n27028 , n27029 , n27030 , n27031 , n27032 , n27033 , n27034 , n27035 , n27036 , n27037 , n27038 , n27039 , n27040 , n27041 , n27042 , n27043 , n27044 , n27045 , n27046 , n27047 , n27048 , n27049 , n27050 , n27051 , n27052 , n27053 , n27054 , n27055 , n27056 , n27057 , n27058 , n27059 , n27060 , n27061 , n27062 , n27063 , n27064 , n27065 , n27066 , n27067 , n27068 , n27069 , n27070 , n27071 , n27072 , n27073 , n27074 , n27075 , n27076 , n27077 , n27078 , n27079 , n27080 , n27081 , n27082 , n27083 , n27084 , n27085 , n27086 , n27087 , n27088 , n27089 , n27090 , n27091 , n27092 , n27093 , n27094 , n27095 , n27096 , n27097 , n27098 , n27099 , n27100 , n27101 , n27102 , n27103 , n27104 , n27105 , n27106 , n27107 , n27108 , n27109 , n27110 , n27111 , n27112 , n27113 , n27114 , n27115 , n27116 , n27117 , n27118 , n27119 , n27120 , n27121 , n27122 , n27123 , n27124 , n27125 , n27126 , n27127 , n27128 , n27129 , n27130 , n27131 , n27132 , n27133 , n27134 , n27135 , n27136 , n27137 , n27138 , n27139 , n27140 , n27141 , n27142 , n27143 , n27144 , n27145 , n27146 , n27147 , n27148 , n27149 , n27150 , n27151 , n27152 , n27153 , n27154 , n27155 , n27156 , n27157 , n27158 , n27159 , n27160 , n27161 , n27162 , n27163 , n27164 , n27165 , n27166 , n27167 , n27168 , n27169 , n27170 , n27171 , n27172 , n27173 , n27174 , n27175 , n27176 , n27177 , n27178 , n27179 , n27180 , n27181 , n27182 , n27183 , n27184 , n27185 , n27186 , n27187 , n27188 , n27189 , n27190 , n27191 , n27192 , n27193 , n27194 , n27195 , n27196 , n27197 , n27198 , n27199 , n27200 , n27201 , n27202 , n27203 , n27204 , n27205 , n27206 , n27207 , n27208 , n27209 , n27210 , n27211 , n27212 , n27213 , n27214 , n27215 , n27216 , n27217 , n27218 , n27219 , n27220 , n27221 , n27222 , n27223 , n27224 , n27225 , n27226 , n27227 , n27228 , n27229 , n27230 , n27231 , n27232 , n27233 , n27234 , n27235 , n27236 , n27237 , n27238 , n27239 , n27240 , n27241 , n27242 , n27243 , n27244 , n27245 , n27246 , n27247 , n27248 , n27249 , n27250 , n27251 , n27252 , n27253 , n27254 , n27255 , n27256 , n27257 , n27258 , n27259 , n27260 , n27261 , n27262 , n27263 , n27264 , n27265 , n27266 , n27267 , n27268 , n27269 , n27270 , n27271 , n27272 , n27273 , n27274 , n27275 , n27276 , n27277 , n27278 , n27279 , n27280 , n27281 , n27282 , n27283 , n27284 , n27285 , n27286 , n27287 , n27288 , n27289 , n27290 , n27291 , n27292 , n27293 , n27294 , n27295 , n27296 , n27297 , n27298 , n27299 , n27300 , n27301 , n27302 , n27303 , n27304 , n27305 , n27306 , n27307 , n27308 , n27309 , n27310 , n27311 , n27312 , n27313 , n27314 , n27315 , n27316 , n27317 , n27318 , n27319 , n27320 , n27321 , n27322 , n27323 , n27324 , n27325 , n27326 , n27327 , n27328 , n27329 , n27330 , n27331 , n27332 , n27333 , n27334 , n27335 , n27336 , n27337 , n27338 , n27339 , n27340 , n27341 , n27342 , n27343 , n27344 , n27345 , n27346 , n27347 , n27348 , n27349 , n27350 , n27351 , n27352 , n27353 , n27354 , n27355 , n27356 , n27357 , n27358 , n27359 , n27360 , n27361 , n27362 , n27363 , n27364 , n27365 , n27366 , n27367 , n27368 , n27369 , n27370 , n27371 , n27372 , n27373 , n27374 , n27375 , n27376 , n27377 , n27378 , n27379 , n27380 , n27381 , n27382 , n27383 , n27384 , n27385 , n27386 , n27387 , n27388 , n27389 , n27390 , n27391 , n27392 , n27393 , n27394 , n27395 , n27396 , n27397 , n27398 , n27399 , n27400 , n27401 , n27402 , n27403 , n27404 , n27405 , n27406 , n27407 , n27408 , n27409 , n27410 , n27411 , n27412 , n27413 , n27414 , n27415 , n27416 , n27417 , n27418 , n27419 , n27420 , n27421 , n27422 , n27423 , n27424 , n27425 , n27426 , n27427 , n27428 , n27429 , n27430 , n27431 , n27432 , n27433 , n27434 , n27435 , n27436 , n27437 , n27438 , n27439 , n27440 , n27441 , n27442 , n27443 , n27444 , n27445 , n27446 , n27447 , n27448 , n27449 , n27450 , n27451 , n27452 , n27453 , n27454 , n27455 , n27456 , n27457 , n27458 , n27459 , n27460 , n27461 , n27462 , n27463 , n27464 , n27465 , n27466 , n27467 , n27468 , n27469 , n27470 , n27471 , n27472 , n27473 , n27474 , n27475 , n27476 , n27477 , n27478 , n27479 , n27480 , n27481 , n27482 , n27483 , n27484 , n27485 , n27486 , n27487 , n27488 , n27489 , n27490 , n27491 , n27492 , n27493 , n27494 , n27495 , n27496 , n27497 , n27498 , n27499 , n27500 , n27501 , n27502 , n27503 , n27504 , n27505 , n27506 , n27507 , n27508 , n27509 , n27510 , n27511 , n27512 , n27513 , n27514 , n27515 , n27516 , n27517 , n27518 , n27519 , n27520 , n27521 , n27522 , n27523 , n27524 , n27525 , n27526 , n27527 , n27528 , n27529 , n27530 , n27531 , n27532 , n27533 , n27534 , n27535 , n27536 , n27537 , n27538 , n27539 , n27540 , n27541 , n27542 , n27543 , n27544 , n27545 , n27546 , n27547 , n27548 , n27549 , n27550 , n27551 , n27552 , n27553 , n27554 , n27555 , n27556 , n27557 , n27558 , n27559 , n27560 , n27561 , n27562 , n27563 , n27564 , n27565 , n27566 , n27567 , n27568 , n27569 , n27570 , n27571 , n27572 , n27573 , n27574 , n27575 , n27576 , n27577 , n27578 , n27579 , n27580 , n27581 , n27582 , n27583 , n27584 , n27585 , n27586 , n27587 , n27588 , n27589 , n27590 , n27591 , n27592 , n27593 , n27594 , n27595 , n27596 , n27597 , n27598 , n27599 , n27600 , n27601 , n27602 , n27603 , n27604 , n27605 , n27606 , n27607 , n27608 , n27609 , n27610 , n27611 , n27612 , n27613 , n27614 , n27615 , n27616 , n27617 , n27618 , n27619 , n27620 , n27621 , n27622 , n27623 , n27624 , n27625 , n27626 , n27627 , n27628 , n27629 , n27630 , n27631 , n27632 , n27633 , n27634 , n27635 , n27636 , n27637 , n27638 , n27639 , n27640 , n27641 , n27642 , n27643 , n27644 , n27645 , n27646 , n27647 , n27648 , n27649 , n27650 , n27651 , n27652 , n27653 , n27654 , n27655 , n27656 , n27657 , n27658 , n27659 , n27660 , n27661 , n27662 , n27663 , n27664 , n27665 , n27666 , n27667 , n27668 , n27669 , n27670 , n27671 , n27672 , n27673 , n27674 , n27675 , n27676 , n27677 , n27678 , n27679 , n27680 , n27681 , n27682 , n27683 , n27684 , n27685 , n27686 , n27687 , n27688 , n27689 , n27690 , n27691 , n27692 , n27693 , n27694 , n27695 , n27696 , n27697 , n27698 , n27699 , n27700 , n27701 , n27702 , n27703 , n27704 , n27705 , n27706 , n27707 , n27708 , n27709 , n27710 , n27711 , n27712 , n27713 , n27714 , n27715 , n27716 , n27717 , n27718 , n27719 , n27720 , n27721 , n27722 , n27723 , n27724 , n27725 , n27726 , n27727 , n27728 , n27729 , n27730 , n27731 , n27732 , n27733 , n27734 , n27735 , n27736 , n27737 , n27738 , n27739 , n27740 , n27741 , n27742 , n27743 , n27744 , n27745 , n27746 , n27747 , n27748 , n27749 , n27750 , n27751 , n27752 , n27753 , n27754 , n27755 , n27756 , n27757 , n27758 , n27759 , n27760 , n27761 , n27762 , n27763 , n27764 , n27765 , n27766 , n27767 , n27768 , n27769 , n27770 , n27771 , n27772 , n27773 , n27774 , n27775 , n27776 , n27777 , n27778 , n27779 , n27780 , n27781 , n27782 , n27783 , n27784 , n27785 , n27786 , n27787 , n27788 , n27789 , n27790 , n27791 , n27792 , n27793 , n27794 , n27795 , n27796 , n27797 , n27798 , n27799 , n27800 , n27801 , n27802 , n27803 , n27804 , n27805 , n27806 , n27807 , n27808 , n27809 , n27810 , n27811 , n27812 , n27813 , n27814 , n27815 , n27816 , n27817 , n27818 , n27819 , n27820 , n27821 , n27822 , n27823 , n27824 , n27825 , n27826 , n27827 , n27828 , n27829 , n27830 , n27831 , n27832 , n27833 , n27834 , n27835 , n27836 , n27837 , n27838 , n27839 , n27840 , n27841 , n27842 , n27843 , n27844 , n27845 , n27846 , n27847 , n27848 , n27849 , n27850 , n27851 , n27852 , n27853 , n27854 , n27855 , n27856 , n27857 , n27858 , n27859 , n27860 , n27861 , n27862 , n27863 , n27864 , n27865 , n27866 , n27867 , n27868 , n27869 , n27870 , n27871 , n27872 , n27873 , n27874 , n27875 , n27876 , n27877 , n27878 , n27879 , n27880 , n27881 , n27882 , n27883 , n27884 , n27885 , n27886 , n27887 , n27888 , n27889 , n27890 , n27891 , n27892 , n27893 , n27894 , n27895 , n27896 , n27897 , n27898 , n27899 , n27900 , n27901 , n27902 , n27903 , n27904 , n27905 , n27906 , n27907 , n27908 , n27909 , n27910 , n27911 , n27912 , n27913 , n27914 , n27915 , n27916 , n27917 , n27918 , n27919 , n27920 , n27921 , n27922 , n27923 , n27924 , n27925 , n27926 , n27927 , n27928 , n27929 , n27930 , n27931 , n27932 , n27933 , n27934 , n27935 , n27936 , n27937 , n27938 , n27939 , n27940 , n27941 , n27942 , n27943 , n27944 , n27945 , n27946 , n27947 , n27948 , n27949 , n27950 , n27951 , n27952 , n27953 , n27954 , n27955 , n27956 , n27957 , n27958 , n27959 , n27960 , n27961 , n27962 , n27963 , n27964 , n27965 , n27966 , n27967 , n27968 , n27969 , n27970 , n27971 , n27972 , n27973 , n27974 , n27975 , n27976 , n27977 , n27978 , n27979 , n27980 , n27981 , n27982 , n27983 , n27984 , n27985 , n27986 , n27987 , n27988 , n27989 , n27990 , n27991 , n27992 , n27993 , n27994 , n27995 , n27996 , n27997 , n27998 , n27999 , n28000 , n28001 , n28002 , n28003 , n28004 , n28005 , n28006 , n28007 , n28008 , n28009 , n28010 , n28011 , n28012 , n28013 , n28014 , n28015 , n28016 , n28017 , n28018 , n28019 , n28020 , n28021 , n28022 , n28023 , n28024 , n28025 , n28026 , n28027 , n28028 , n28029 , n28030 , n28031 , n28032 , n28033 , n28034 , n28035 , n28036 , n28037 , n28038 , n28039 , n28040 , n28041 , n28042 , n28043 , n28044 , n28045 , n28046 , n28047 , n28048 , n28049 , n28050 , n28051 , n28052 , n28053 , n28054 , n28055 , n28056 , n28057 , n28058 , n28059 , n28060 , n28061 , n28062 , n28063 , n28064 , n28065 , n28066 , n28067 , n28068 , n28069 , n28070 , n28071 , n28072 , n28073 , n28074 , n28075 , n28076 , n28077 , n28078 , n28079 , n28080 , n28081 , n28082 , n28083 , n28084 , n28085 , n28086 , n28087 , n28088 , n28089 , n28090 , n28091 , n28092 , n28093 , n28094 , n28095 , n28096 , n28097 , n28098 , n28099 , n28100 , n28101 , n28102 , n28103 , n28104 , n28105 , n28106 , n28107 , n28108 , n28109 , n28110 , n28111 , n28112 , n28113 , n28114 , n28115 , n28116 , n28117 , n28118 , n28119 , n28120 , n28121 , n28122 , n28123 , n28124 , n28125 , n28126 , n28127 , n28128 , n28129 , n28130 , n28131 , n28132 , n28133 , n28134 , n28135 , n28136 , n28137 , n28138 , n28139 , n28140 , n28141 , n28142 , n28143 , n28144 , n28145 , n28146 , n28147 , n28148 , n28149 , n28150 , n28151 , n28152 , n28153 , n28154 , n28155 , n28156 , n28157 , n28158 , n28159 , n28160 , n28161 , n28162 , n28163 , n28164 , n28165 , n28166 , n28167 , n28168 , n28169 , n28170 , n28171 , n28172 , n28173 , n28174 , n28175 , n28176 , n28177 , n28178 , n28179 , n28180 , n28181 , n28182 , n28183 , n28184 , n28185 , n28186 , n28187 , n28188 , n28189 , n28190 , n28191 , n28192 , n28193 , n28194 , n28195 , n28196 , n28197 , n28198 , n28199 , n28200 , n28201 , n28202 , n28203 , n28204 , n28205 , n28206 , n28207 , n28208 , n28209 , n28210 , n28211 , n28212 , n28213 , n28214 , n28215 , n28216 , n28217 , n28218 , n28219 , n28220 , n28221 , n28222 , n28223 , n28224 , n28225 , n28226 , n28227 , n28228 , n28229 , n28230 , n28231 , n28232 , n28233 , n28234 , n28235 , n28236 , n28237 , n28238 , n28239 , n28240 , n28241 , n28242 , n28243 , n28244 , n28245 , n28246 , n28247 , n28248 , n28249 , n28250 , n28251 , n28252 , n28253 , n28254 , n28255 , n28256 , n28257 , n28258 , n28259 , n28260 , n28261 , n28262 , n28263 , n28264 , n28265 , n28266 , n28267 , n28268 , n28269 , n28270 , n28271 , n28272 , n28273 , n28274 , n28275 , n28276 , n28277 , n28278 , n28279 , n28280 , n28281 , n28282 , n28283 , n28284 , n28285 , n28286 , n28287 , n28288 , n28289 , n28290 , n28291 , n28292 , n28293 , n28294 , n28295 , n28296 , n28297 , n28298 , n28299 , n28300 , n28301 , n28302 , n28303 , n28304 , n28305 , n28306 , n28307 , n28308 , n28309 , n28310 , n28311 , n28312 , n28313 , n28314 , n28315 , n28316 , n28317 , n28318 , n28319 , n28320 , n28321 , n28322 , n28323 , n28324 , n28325 , n28326 , n28327 , n28328 , n28329 , n28330 , n28331 , n28332 , n28333 , n28334 , n28335 , n28336 , n28337 , n28338 , n28339 , n28340 , n28341 , n28342 , n28343 , n28344 , n28345 , n28346 , n28347 , n28348 , n28349 , n28350 , n28351 , n28352 , n28353 , n28354 , n28355 , n28356 , n28357 , n28358 , n28359 , n28360 , n28361 , n28362 , n28363 , n28364 , n28365 , n28366 , n28367 , n28368 , n28369 , n28370 , n28371 , n28372 , n28373 , n28374 , n28375 , n28376 , n28377 , n28378 , n28379 , n28380 , n28381 , n28382 , n28383 , n28384 , n28385 , n28386 , n28387 , n28388 , n28389 , n28390 , n28391 , n28392 , n28393 , n28394 , n28395 , n28396 , n28397 , n28398 , n28399 , n28400 , n28401 , n28402 , n28403 , n28404 , n28405 , n28406 , n28407 , n28408 , n28409 , n28410 , n28411 , n28412 , n28413 , n28414 , n28415 , n28416 , n28417 , n28418 , n28419 , n28420 , n28421 , n28422 , n28423 , n28424 , n28425 , n28426 , n28427 , n28428 , n28429 , n28430 , n28431 , n28432 , n28433 , n28434 , n28435 , n28436 , n28437 , n28438 , n28439 , n28440 , n28441 , n28442 , n28443 , n28444 , n28445 , n28446 , n28447 , n28448 , n28449 , n28450 , n28451 , n28452 , n28453 , n28454 , n28455 , n28456 , n28457 , n28458 , n28459 , n28460 , n28461 , n28462 , n28463 , n28464 , n28465 , n28466 , n28467 , n28468 , n28469 , n28470 , n28471 , n28472 , n28473 , n28474 , n28475 , n28476 , n28477 , n28478 , n28479 , n28480 , n28481 , n28482 , n28483 , n28484 , n28485 , n28486 , n28487 , n28488 , n28489 , n28490 , n28491 , n28492 , n28493 , n28494 , n28495 , n28496 , n28497 , n28498 , n28499 , n28500 , n28501 , n28502 , n28503 , n28504 , n28505 , n28506 , n28507 , n28508 , n28509 , n28510 , n28511 , n28512 , n28513 , n28514 , n28515 , n28516 , n28517 , n28518 , n28519 , n28520 , n28521 , n28522 , n28523 , n28524 , n28525 , n28526 , n28527 , n28528 , n28529 , n28530 , n28531 , n28532 , n28533 , n28534 , n28535 , n28536 , n28537 , n28538 , n28539 , n28540 , n28541 , n28542 , n28543 , n28544 , n28545 , n28546 , n28547 , n28548 , n28549 , n28550 , n28551 , n28552 , n28553 , n28554 , n28555 , n28556 , n28557 , n28558 , n28559 , n28560 , n28561 , n28562 , n28563 , n28564 , n28565 , n28566 , n28567 , n28568 , n28569 , n28570 , n28571 , n28572 , n28573 , n28574 , n28575 , n28576 , n28577 , n28578 , n28579 , n28580 , n28581 , n28582 , n28583 , n28584 , n28585 , n28586 , n28587 , n28588 , n28589 , n28590 , n28591 , n28592 , n28593 , n28594 , n28595 , n28596 , n28597 , n28598 , n28599 , n28600 , n28601 , n28602 , n28603 , n28604 , n28605 , n28606 , n28607 , n28608 , n28609 , n28610 , n28611 , n28612 , n28613 , n28614 , n28615 , n28616 , n28617 , n28618 , n28619 , n28620 , n28621 , n28622 , n28623 , n28624 , n28625 , n28626 , n28627 , n28628 , n28629 , n28630 , n28631 , n28632 , n28633 , n28634 , n28635 , n28636 , n28637 , n28638 , n28639 , n28640 , n28641 , n28642 , n28643 , n28644 , n28645 , n28646 , n28647 , n28648 , n28649 , n28650 , n28651 , n28652 , n28653 , n28654 , n28655 , n28656 , n28657 , n28658 , n28659 , n28660 , n28661 , n28662 , n28663 , n28664 , n28665 , n28666 , n28667 , n28668 , n28669 , n28670 , n28671 , n28672 , n28673 , n28674 , n28675 , n28676 , n28677 , n28678 , n28679 , n28680 , n28681 , n28682 , n28683 , n28684 , n28685 , n28686 , n28687 , n28688 , n28689 , n28690 , n28691 , n28692 , n28693 , n28694 , n28695 , n28696 , n28697 , n28698 , n28699 , n28700 , n28701 , n28702 , n28703 , n28704 , n28705 , n28706 , n28707 , n28708 , n28709 , n28710 , n28711 , n28712 , n28713 , n28714 , n28715 , n28716 , n28717 , n28718 , n28719 , n28720 , n28721 , n28722 , n28723 , n28724 , n28725 , n28726 , n28727 , n28728 , n28729 , n28730 , n28731 , n28732 , n28733 , n28734 , n28735 , n28736 , n28737 , n28738 , n28739 , n28740 , n28741 , n28742 , n28743 , n28744 , n28745 , n28746 , n28747 , n28748 , n28749 , n28750 , n28751 , n28752 , n28753 , n28754 , n28755 , n28756 , n28757 , n28758 , n28759 , n28760 , n28761 , n28762 , n28763 , n28764 , n28765 , n28766 , n28767 , n28768 , n28769 , n28770 , n28771 , n28772 , n28773 , n28774 , n28775 , n28776 , n28777 , n28778 , n28779 , n28780 , n28781 , n28782 , n28783 , n28784 , n28785 , n28786 , n28787 , n28788 , n28789 , n28790 , n28791 , n28792 , n28793 , n28794 , n28795 , n28796 , n28797 , n28798 , n28799 , n28800 , n28801 , n28802 , n28803 , n28804 , n28805 , n28806 , n28807 , n28808 , n28809 , n28810 , n28811 , n28812 , n28813 , n28814 , n28815 , n28816 , n28817 , n28818 , n28819 , n28820 , n28821 , n28822 , n28823 , n28824 , n28825 , n28826 , n28827 , n28828 , n28829 , n28830 , n28831 , n28832 , n28833 , n28834 , n28835 , n28836 , n28837 , n28838 , n28839 , n28840 , n28841 , n28842 , n28843 , n28844 , n28845 , n28846 , n28847 , n28848 , n28849 , n28850 , n28851 , n28852 , n28853 , n28854 , n28855 , n28856 , n28857 , n28858 , n28859 , n28860 , n28861 , n28862 , n28863 , n28864 , n28865 , n28866 , n28867 , n28868 , n28869 , n28870 , n28871 , n28872 , n28873 , n28874 , n28875 , n28876 , n28877 , n28878 , n28879 , n28880 , n28881 , n28882 , n28883 , n28884 , n28885 , n28886 , n28887 , n28888 , n28889 , n28890 , n28891 , n28892 , n28893 , n28894 , n28895 , n28896 , n28897 , n28898 , n28899 , n28900 , n28901 , n28902 , n28903 , n28904 , n28905 , n28906 , n28907 , n28908 , n28909 , n28910 , n28911 , n28912 , n28913 , n28914 , n28915 , n28916 , n28917 , n28918 , n28919 , n28920 , n28921 , n28922 , n28923 , n28924 , n28925 , n28926 , n28927 , n28928 , n28929 , n28930 , n28931 , n28932 , n28933 , n28934 , n28935 , n28936 , n28937 , n28938 , n28939 , n28940 , n28941 , n28942 , n28943 , n28944 , n28945 , n28946 , n28947 , n28948 , n28949 , n28950 , n28951 , n28952 , n28953 , n28954 , n28955 , n28956 , n28957 , n28958 , n28959 , n28960 , n28961 , n28962 , n28963 , n28964 , n28965 , n28966 , n28967 , n28968 , n28969 , n28970 , n28971 , n28972 , n28973 , n28974 , n28975 , n28976 , n28977 , n28978 , n28979 , n28980 , n28981 , n28982 , n28983 , n28984 , n28985 , n28986 , n28987 , n28988 , n28989 , n28990 , n28991 , n28992 , n28993 , n28994 , n28995 , n28996 , n28997 , n28998 , n28999 , n29000 , n29001 , n29002 , n29003 , n29004 , n29005 , n29006 , n29007 , n29008 , n29009 , n29010 , n29011 , n29012 , n29013 , n29014 , n29015 , n29016 , n29017 , n29018 , n29019 , n29020 , n29021 , n29022 , n29023 , n29024 , n29025 , n29026 , n29027 , n29028 , n29029 , n29030 , n29031 , n29032 , n29033 , n29034 , n29035 , n29036 , n29037 , n29038 , n29039 , n29040 , n29041 , n29042 , n29043 , n29044 , n29045 , n29046 , n29047 , n29048 , n29049 , n29050 , n29051 , n29052 , n29053 , n29054 , n29055 , n29056 , n29057 , n29058 , n29059 , n29060 , n29061 , n29062 , n29063 , n29064 , n29065 , n29066 , n29067 , n29068 , n29069 , n29070 , n29071 , n29072 , n29073 , n29074 , n29075 , n29076 , n29077 , n29078 , n29079 , n29080 , n29081 , n29082 , n29083 , n29084 , n29085 , n29086 , n29087 , n29088 , n29089 , n29090 , n29091 , n29092 , n29093 , n29094 , n29095 , n29096 , n29097 , n29098 , n29099 , n29100 , n29101 , n29102 , n29103 , n29104 , n29105 , n29106 , n29107 , n29108 , n29109 , n29110 , n29111 , n29112 , n29113 , n29114 , n29115 , n29116 , n29117 , n29118 , n29119 , n29120 , n29121 , n29122 , n29123 , n29124 , n29125 , n29126 , n29127 , n29128 , n29129 , n29130 , n29131 , n29132 , n29133 , n29134 , n29135 , n29136 , n29137 , n29138 , n29139 , n29140 , n29141 , n29142 , n29143 , n29144 , n29145 , n29146 , n29147 , n29148 , n29149 , n29150 , n29151 , n29152 , n29153 , n29154 , n29155 , n29156 , n29157 , n29158 , n29159 , n29160 , n29161 , n29162 , n29163 , n29164 , n29165 , n29166 , n29167 , n29168 , n29169 , n29170 , n29171 , n29172 , n29173 , n29174 , n29175 , n29176 , n29177 , n29178 , n29179 , n29180 , n29181 , n29182 , n29183 , n29184 , n29185 , n29186 , n29187 , n29188 , n29189 , n29190 , n29191 , n29192 , n29193 , n29194 , n29195 , n29196 , n29197 , n29198 , n29199 , n29200 , n29201 , n29202 , n29203 , n29204 , n29205 , n29206 , n29207 , n29208 , n29209 , n29210 , n29211 , n29212 , n29213 , n29214 , n29215 , n29216 , n29217 , n29218 , n29219 , n29220 , n29221 , n29222 , n29223 , n29224 , n29225 , n29226 , n29227 , n29228 , n29229 , n29230 , n29231 , n29232 , n29233 , n29234 , n29235 , n29236 , n29237 , n29238 , n29239 , n29240 , n29241 , n29242 , n29243 , n29244 , n29245 , n29246 , n29247 , n29248 , n29249 , n29250 , n29251 , n29252 , n29253 , n29254 , n29255 , n29256 , n29257 , n29258 , n29259 , n29260 , n29261 , n29262 , n29263 , n29264 , n29265 , n29266 , n29267 , n29268 , n29269 , n29270 , n29271 , n29272 , n29273 , n29274 , n29275 , n29276 , n29277 , n29278 , n29279 , n29280 , n29281 , n29282 , n29283 , n29284 , n29285 , n29286 , n29287 , n29288 , n29289 , n29290 , n29291 , n29292 , n29293 , n29294 , n29295 , n29296 , n29297 , n29298 , n29299 , n29300 , n29301 , n29302 , n29303 , n29304 , n29305 , n29306 , n29307 , n29308 , n29309 , n29310 , n29311 , n29312 , n29313 , n29314 , n29315 , n29316 , n29317 , n29318 , n29319 , n29320 , n29321 , n29322 , n29323 , n29324 , n29325 , n29326 , n29327 , n29328 , n29329 , n29330 , n29331 , n29332 , n29333 , n29334 , n29335 , n29336 , n29337 , n29338 , n29339 , n29340 , n29341 , n29342 , n29343 , n29344 , n29345 , n29346 , n29347 , n29348 , n29349 , n29350 , n29351 , n29352 , n29353 , n29354 , n29355 , n29356 , n29357 , n29358 , n29359 , n29360 , n29361 , n29362 , n29363 , n29364 , n29365 , n29366 , n29367 , n29368 , n29369 , n29370 , n29371 , n29372 , n29373 , n29374 , n29375 , n29376 , n29377 , n29378 , n29379 , n29380 , n29381 , n29382 , n29383 , n29384 , n29385 , n29386 , n29387 , n29388 , n29389 , n29390 , n29391 , n29392 , n29393 , n29394 , n29395 , n29396 , n29397 , n29398 , n29399 , n29400 , n29401 , n29402 , n29403 , n29404 , n29405 , n29406 , n29407 , n29408 , n29409 , n29410 , n29411 , n29412 , n29413 , n29414 , n29415 , n29416 , n29417 , n29418 , n29419 , n29420 , n29421 , n29422 , n29423 , n29424 , n29425 , n29426 , n29427 , n29428 , n29429 , n29430 , n29431 , n29432 , n29433 , n29434 , n29435 , n29436 , n29437 , n29438 , n29439 , n29440 , n29441 , n29442 , n29443 , n29444 , n29445 , n29446 , n29447 , n29448 , n29449 , n29450 , n29451 , n29452 , n29453 , n29454 , n29455 , n29456 , n29457 , n29458 , n29459 , n29460 , n29461 , n29462 , n29463 , n29464 , n29465 , n29466 , n29467 , n29468 , n29469 , n29470 , n29471 , n29472 , n29473 , n29474 , n29475 , n29476 , n29477 , n29478 , n29479 , n29480 , n29481 , n29482 , n29483 , n29484 , n29485 , n29486 , n29487 , n29488 , n29489 , n29490 , n29491 , n29492 , n29493 , n29494 , n29495 , n29496 , n29497 , n29498 , n29499 , n29500 , n29501 , n29502 , n29503 , n29504 , n29505 , n29506 , n29507 , n29508 , n29509 , n29510 , n29511 , n29512 , n29513 , n29514 , n29515 , n29516 , n29517 , n29518 , n29519 , n29520 , n29521 , n29522 , n29523 , n29524 , n29525 , n29526 , n29527 , n29528 , n29529 , n29530 , n29531 , n29532 , n29533 , n29534 , n29535 , n29536 , n29537 , n29538 , n29539 , n29540 , n29541 , n29542 , n29543 , n29544 , n29545 , n29546 , n29547 , n29548 , n29549 , n29550 , n29551 , n29552 , n29553 , n29554 , n29555 , n29556 , n29557 , n29558 , n29559 , n29560 , n29561 , n29562 , n29563 , n29564 , n29565 , n29566 , n29567 , n29568 , n29569 , n29570 , n29571 , n29572 , n29573 , n29574 , n29575 , n29576 , n29577 , n29578 , n29579 , n29580 , n29581 , n29582 , n29583 , n29584 , n29585 , n29586 , n29587 , n29588 , n29589 , n29590 , n29591 , n29592 , n29593 , n29594 , n29595 , n29596 , n29597 , n29598 , n29599 , n29600 , n29601 , n29602 , n29603 , n29604 , n29605 , n29606 , n29607 , n29608 , n29609 , n29610 , n29611 , n29612 , n29613 , n29614 , n29615 , n29616 , n29617 , n29618 , n29619 , n29620 , n29621 , n29622 , n29623 , n29624 , n29625 , n29626 , n29627 , n29628 , n29629 , n29630 , n29631 , n29632 , n29633 , n29634 , n29635 , n29636 , n29637 , n29638 , n29639 , n29640 , n29641 , n29642 , n29643 , n29644 , n29645 , n29646 , n29647 , n29648 , n29649 , n29650 , n29651 , n29652 , n29653 , n29654 , n29655 , n29656 , n29657 , n29658 , n29659 , n29660 , n29661 , n29662 , n29663 , n29664 , n29665 , n29666 , n29667 , n29668 , n29669 , n29670 , n29671 , n29672 , n29673 , n29674 , n29675 , n29676 , n29677 , n29678 , n29679 , n29680 , n29681 , n29682 , n29683 , n29684 , n29685 , n29686 , n29687 , n29688 , n29689 , n29690 , n29691 , n29692 , n29693 , n29694 , n29695 , n29696 , n29697 , n29698 , n29699 , n29700 , n29701 , n29702 , n29703 , n29704 , n29705 , n29706 , n29707 , n29708 , n29709 , n29710 , n29711 , n29712 , n29713 , n29714 , n29715 , n29716 , n29717 , n29718 , n29719 , n29720 , n29721 , n29722 , n29723 , n29724 , n29725 , n29726 , n29727 , n29728 , n29729 , n29730 , n29731 , n29732 , n29733 , n29734 , n29735 , n29736 , n29737 , n29738 , n29739 , n29740 , n29741 , n29742 , n29743 , n29744 , n29745 , n29746 , n29747 , n29748 , n29749 , n29750 , n29751 , n29752 , n29753 , n29754 , n29755 , n29756 , n29757 , n29758 , n29759 , n29760 , n29761 , n29762 , n29763 , n29764 , n29765 , n29766 , n29767 , n29768 , n29769 , n29770 , n29771 , n29772 , n29773 , n29774 , n29775 , n29776 , n29777 , n29778 , n29779 , n29780 , n29781 , n29782 , n29783 , n29784 , n29785 , n29786 , n29787 , n29788 , n29789 , n29790 , n29791 , n29792 , n29793 , n29794 , n29795 , n29796 , n29797 , n29798 , n29799 , n29800 , n29801 , n29802 , n29803 , n29804 , n29805 , n29806 , n29807 , n29808 , n29809 , n29810 , n29811 , n29812 , n29813 , n29814 , n29815 , n29816 , n29817 , n29818 , n29819 , n29820 , n29821 , n29822 , n29823 , n29824 , n29825 , n29826 , n29827 , n29828 , n29829 , n29830 , n29831 , n29832 , n29833 , n29834 , n29835 , n29836 , n29837 , n29838 , n29839 , n29840 , n29841 , n29842 , n29843 , n29844 , n29845 , n29846 , n29847 , n29848 , n29849 , n29850 , n29851 , n29852 , n29853 , n29854 , n29855 , n29856 , n29857 , n29858 , n29859 , n29860 , n29861 , n29862 , n29863 , n29864 , n29865 , n29866 , n29867 , n29868 , n29869 , n29870 , n29871 , n29872 , n29873 , n29874 , n29875 , n29876 , n29877 , n29878 , n29879 , n29880 , n29881 , n29882 , n29883 , n29884 , n29885 , n29886 , n29887 , n29888 , n29889 , n29890 , n29891 , n29892 , n29893 , n29894 , n29895 , n29896 , n29897 , n29898 , n29899 , n29900 , n29901 , n29902 , n29903 , n29904 , n29905 , n29906 , n29907 , n29908 , n29909 , n29910 , n29911 , n29912 , n29913 , n29914 , n29915 , n29916 , n29917 , n29918 , n29919 , n29920 , n29921 , n29922 , n29923 , n29924 , n29925 , n29926 , n29927 , n29928 , n29929 , n29930 , n29931 , n29932 , n29933 , n29934 , n29935 , n29936 , n29937 , n29938 , n29939 , n29940 , n29941 , n29942 , n29943 , n29944 , n29945 , n29946 , n29947 , n29948 , n29949 , n29950 , n29951 , n29952 , n29953 , n29954 , n29955 , n29956 , n29957 , n29958 , n29959 , n29960 , n29961 , n29962 , n29963 , n29964 , n29965 , n29966 , n29967 , n29968 , n29969 , n29970 , n29971 , n29972 , n29973 , n29974 , n29975 , n29976 , n29977 , n29978 , n29979 , n29980 , n29981 , n29982 , n29983 , n29984 , n29985 , n29986 , n29987 , n29988 , n29989 , n29990 , n29991 , n29992 , n29993 , n29994 , n29995 , n29996 , n29997 , n29998 , n29999 , n30000 , n30001 , n30002 , n30003 , n30004 , n30005 , n30006 , n30007 , n30008 , n30009 , n30010 , n30011 , n30012 , n30013 , n30014 , n30015 , n30016 , n30017 , n30018 , n30019 , n30020 , n30021 , n30022 , n30023 , n30024 , n30025 , n30026 , n30027 , n30028 , n30029 , n30030 , n30031 , n30032 , n30033 , n30034 , n30035 , n30036 , n30037 , n30038 , n30039 , n30040 , n30041 , n30042 , n30043 , n30044 , n30045 , n30046 , n30047 , n30048 , n30049 , n30050 , n30051 , n30052 , n30053 , n30054 , n30055 , n30056 , n30057 , n30058 , n30059 , n30060 , n30061 , n30062 , n30063 , n30064 , n30065 , n30066 , n30067 , n30068 , n30069 , n30070 , n30071 , n30072 , n30073 , n30074 , n30075 , n30076 , n30077 , n30078 , n30079 , n30080 , n30081 , n30082 , n30083 , n30084 , n30085 , n30086 , n30087 , n30088 , n30089 , n30090 , n30091 , n30092 , n30093 , n30094 , n30095 , n30096 , n30097 , n30098 , n30099 , n30100 , n30101 , n30102 , n30103 , n30104 , n30105 , n30106 , n30107 , n30108 , n30109 , n30110 , n30111 , n30112 , n30113 , n30114 , n30115 , n30116 , n30117 , n30118 , n30119 , n30120 , n30121 , n30122 , n30123 , n30124 , n30125 , n30126 , n30127 , n30128 , n30129 , n30130 , n30131 , n30132 , n30133 , n30134 , n30135 , n30136 , n30137 , n30138 , n30139 , n30140 , n30141 , n30142 , n30143 , n30144 , n30145 , n30146 , n30147 , n30148 , n30149 , n30150 , n30151 , n30152 , n30153 , n30154 , n30155 , n30156 , n30157 , n30158 , n30159 , n30160 , n30161 , n30162 , n30163 , n30164 , n30165 , n30166 , n30167 , n30168 , n30169 , n30170 , n30171 , n30172 , n30173 , n30174 , n30175 , n30176 , n30177 , n30178 , n30179 , n30180 , n30181 , n30182 , n30183 , n30184 , n30185 , n30186 , n30187 , n30188 , n30189 , n30190 , n30191 , n30192 , n30193 , n30194 , n30195 , n30196 , n30197 , n30198 , n30199 , n30200 , n30201 , n30202 , n30203 , n30204 , n30205 , n30206 , n30207 , n30208 , n30209 , n30210 , n30211 , n30212 , n30213 , n30214 , n30215 , n30216 , n30217 , n30218 , n30219 , n30220 , n30221 , n30222 , n30223 , n30224 , n30225 , n30226 , n30227 , n30228 , n30229 , n30230 , n30231 , n30232 , n30233 , n30234 , n30235 , n30236 , n30237 , n30238 , n30239 , n30240 , n30241 , n30242 , n30243 , n30244 , n30245 , n30246 , n30247 , n30248 , n30249 , n30250 , n30251 , n30252 , n30253 , n30254 , n30255 , n30256 , n30257 , n30258 , n30259 , n30260 , n30261 , n30262 , n30263 , n30264 , n30265 , n30266 , n30267 , n30268 , n30269 , n30270 , n30271 , n30272 , n30273 , n30274 , n30275 , n30276 , n30277 , n30278 , n30279 , n30280 , n30281 , n30282 , n30283 , n30284 , n30285 , n30286 , n30287 , n30288 , n30289 , n30290 , n30291 , n30292 , n30293 , n30294 , n30295 , n30296 , n30297 , n30298 , n30299 , n30300 , n30301 , n30302 , n30303 , n30304 , n30305 , n30306 , n30307 , n30308 , n30309 , n30310 , n30311 , n30312 , n30313 , n30314 , n30315 , n30316 , n30317 , n30318 , n30319 , n30320 , n30321 , n30322 , n30323 , n30324 , n30325 , n30326 , n30327 , n30328 , n30329 , n30330 , n30331 , n30332 , n30333 , n30334 , n30335 , n30336 , n30337 , n30338 , n30339 , n30340 , n30341 , n30342 , n30343 , n30344 , n30345 , n30346 , n30347 , n30348 , n30349 , n30350 , n30351 , n30352 , n30353 , n30354 , n30355 , n30356 , n30357 , n30358 , n30359 , n30360 , n30361 , n30362 , n30363 , n30364 , n30365 , n30366 , n30367 , n30368 , n30369 , n30370 , n30371 , n30372 , n30373 , n30374 , n30375 , n30376 , n30377 , n30378 , n30379 , n30380 , n30381 , n30382 , n30383 , n30384 , n30385 , n30386 , n30387 , n30388 , n30389 , n30390 , n30391 , n30392 , n30393 , n30394 , n30395 , n30396 , n30397 , n30398 , n30399 , n30400 , n30401 , n30402 , n30403 , n30404 , n30405 , n30406 , n30407 , n30408 , n30409 , n30410 , n30411 , n30412 , n30413 , n30414 , n30415 , n30416 , n30417 , n30418 , n30419 , n30420 , n30421 , n30422 , n30423 , n30424 , n30425 , n30426 , n30427 , n30428 , n30429 , n30430 , n30431 , n30432 , n30433 , n30434 , n30435 , n30436 , n30437 , n30438 , n30439 , n30440 , n30441 , n30442 , n30443 , n30444 , n30445 , n30446 , n30447 , n30448 , n30449 , n30450 , n30451 , n30452 , n30453 , n30454 , n30455 , n30456 , n30457 , n30458 , n30459 , n30460 , n30461 , n30462 , n30463 , n30464 , n30465 , n30466 , n30467 , n30468 , n30469 , n30470 , n30471 , n30472 , n30473 , n30474 , n30475 , n30476 , n30477 , n30478 , n30479 , n30480 , n30481 , n30482 , n30483 , n30484 , n30485 , n30486 , n30487 , n30488 , n30489 , n30490 , n30491 , n30492 , n30493 , n30494 , n30495 , n30496 , n30497 , n30498 , n30499 , n30500 , n30501 , n30502 , n30503 , n30504 , n30505 , n30506 , n30507 , n30508 , n30509 , n30510 , n30511 , n30512 , n30513 , n30514 , n30515 , n30516 , n30517 , n30518 , n30519 , n30520 , n30521 , n30522 , n30523 , n30524 , n30525 , n30526 , n30527 , n30528 , n30529 , n30530 , n30531 , n30532 , n30533 , n30534 , n30535 , n30536 , n30537 , n30538 , n30539 , n30540 , n30541 , n30542 , n30543 , n30544 , n30545 , n30546 , n30547 , n30548 , n30549 , n30550 , n30551 , n30552 , n30553 , n30554 , n30555 , n30556 , n30557 , n30558 , n30559 , n30560 , n30561 , n30562 , n30563 , n30564 , n30565 , n30566 , n30567 , n30568 , n30569 , n30570 , n30571 , n30572 , n30573 , n30574 , n30575 , n30576 , n30577 , n30578 , n30579 , n30580 , n30581 , n30582 , n30583 , n30584 , n30585 , n30586 , n30587 , n30588 , n30589 , n30590 , n30591 , n30592 , n30593 , n30594 , n30595 , n30596 , n30597 , n30598 , n30599 , n30600 , n30601 , n30602 , n30603 , n30604 , n30605 , n30606 , n30607 , n30608 , n30609 , n30610 , n30611 , n30612 , n30613 , n30614 , n30615 , n30616 , n30617 , n30618 , n30619 , n30620 , n30621 , n30622 , n30623 , n30624 , n30625 , n30626 , n30627 , n30628 , n30629 , n30630 , n30631 , n30632 , n30633 , n30634 , n30635 , n30636 , n30637 , n30638 , n30639 , n30640 , n30641 , n30642 , n30643 , n30644 , n30645 , n30646 , n30647 , n30648 , n30649 , n30650 , n30651 , n30652 , n30653 , n30654 , n30655 , n30656 , n30657 , n30658 , n30659 , n30660 , n30661 , n30662 , n30663 , n30664 , n30665 , n30666 , n30667 , n30668 , n30669 , n30670 , n30671 , n30672 , n30673 , n30674 , n30675 , n30676 , n30677 , n30678 , n30679 , n30680 , n30681 , n30682 , n30683 , n30684 , n30685 , n30686 , n30687 , n30688 , n30689 , n30690 , n30691 , n30692 , n30693 , n30694 , n30695 , n30696 , n30697 , n30698 , n30699 , n30700 , n30701 , n30702 , n30703 , n30704 , n30705 , n30706 , n30707 , n30708 , n30709 , n30710 , n30711 , n30712 , n30713 , n30714 , n30715 , n30716 , n30717 , n30718 , n30719 , n30720 , n30721 , n30722 , n30723 , n30724 , n30725 , n30726 , n30727 , n30728 , n30729 , n30730 , n30731 , n30732 , n30733 , n30734 , n30735 , n30736 , n30737 , n30738 , n30739 , n30740 , n30741 , n30742 , n30743 , n30744 , n30745 , n30746 , n30747 , n30748 , n30749 , n30750 , n30751 , n30752 , n30753 , n30754 , n30755 , n30756 , n30757 , n30758 , n30759 , n30760 , n30761 , n30762 , n30763 , n30764 , n30765 , n30766 , n30767 , n30768 , n30769 , n30770 , n30771 , n30772 , n30773 , n30774 , n30775 , n30776 , n30777 , n30778 , n30779 , n30780 , n30781 , n30782 , n30783 , n30784 , n30785 , n30786 , n30787 , n30788 , n30789 , n30790 , n30791 , n30792 , n30793 , n30794 , n30795 , n30796 , n30797 , n30798 , n30799 , n30800 , n30801 , n30802 , n30803 , n30804 , n30805 , n30806 , n30807 , n30808 , n30809 , n30810 , n30811 , n30812 , n30813 , n30814 , n30815 , n30816 , n30817 , n30818 , n30819 , n30820 , n30821 , n30822 , n30823 , n30824 , n30825 , n30826 , n30827 , n30828 , n30829 , n30830 , n30831 , n30832 , n30833 , n30834 , n30835 , n30836 , n30837 , n30838 , n30839 , n30840 , n30841 , n30842 , n30843 , n30844 , n30845 , n30846 , n30847 , n30848 , n30849 , n30850 , n30851 , n30852 , n30853 , n30854 , n30855 , n30856 , n30857 , n30858 , n30859 , n30860 , n30861 , n30862 , n30863 , n30864 , n30865 , n30866 , n30867 , n30868 , n30869 , n30870 , n30871 , n30872 , n30873 , n30874 , n30875 , n30876 , n30877 , n30878 , n30879 , n30880 , n30881 , n30882 , n30883 , n30884 , n30885 , n30886 , n30887 , n30888 , n30889 , n30890 , n30891 , n30892 , n30893 , n30894 , n30895 , n30896 , n30897 , n30898 , n30899 , n30900 , n30901 , n30902 , n30903 , n30904 , n30905 , n30906 , n30907 , n30908 , n30909 , n30910 , n30911 , n30912 , n30913 , n30914 , n30915 , n30916 , n30917 , n30918 , n30919 , n30920 , n30921 , n30922 , n30923 , n30924 , n30925 , n30926 , n30927 , n30928 , n30929 , n30930 , n30931 , n30932 , n30933 , n30934 , n30935 , n30936 , n30937 , n30938 , n30939 , n30940 , n30941 , n30942 , n30943 , n30944 , n30945 , n30946 , n30947 , n30948 , n30949 , n30950 , n30951 , n30952 , n30953 , n30954 , n30955 , n30956 , n30957 , n30958 , n30959 , n30960 , n30961 , n30962 , n30963 , n30964 , n30965 , n30966 , n30967 , n30968 , n30969 , n30970 , n30971 , n30972 , n30973 , n30974 , n30975 , n30976 , n30977 , n30978 , n30979 , n30980 , n30981 , n30982 , n30983 , n30984 , n30985 , n30986 , n30987 , n30988 , n30989 , n30990 , n30991 , n30992 , n30993 , n30994 , n30995 , n30996 , n30997 , n30998 , n30999 , n31000 , n31001 , n31002 , n31003 , n31004 , n31005 , n31006 , n31007 , n31008 , n31009 , n31010 , n31011 , n31012 , n31013 , n31014 , n31015 , n31016 , n31017 , n31018 , n31019 , n31020 , n31021 , n31022 , n31023 , n31024 , n31025 , n31026 , n31027 , n31028 , n31029 , n31030 , n31031 , n31032 , n31033 , n31034 , n31035 , n31036 , n31037 , n31038 , n31039 , n31040 , n31041 , n31042 , n31043 , n31044 , n31045 , n31046 , n31047 , n31048 , n31049 , n31050 , n31051 , n31052 , n31053 , n31054 , n31055 , n31056 , n31057 , n31058 , n31059 , n31060 , n31061 , n31062 , n31063 , n31064 , n31065 , n31066 , n31067 , n31068 , n31069 , n31070 , n31071 , n31072 , n31073 , n31074 , n31075 , n31076 , n31077 , n31078 , n31079 , n31080 , n31081 , n31082 , n31083 , n31084 , n31085 , n31086 , n31087 , n31088 , n31089 , n31090 , n31091 , n31092 , n31093 , n31094 , n31095 , n31096 , n31097 , n31098 , n31099 , n31100 , n31101 , n31102 , n31103 , n31104 , n31105 , n31106 , n31107 , n31108 , n31109 , n31110 , n31111 , n31112 , n31113 , n31114 , n31115 , n31116 , n31117 , n31118 , n31119 , n31120 , n31121 , n31122 , n31123 , n31124 , n31125 , n31126 , n31127 , n31128 , n31129 , n31130 , n31131 , n31132 , n31133 , n31134 , n31135 , n31136 , n31137 , n31138 , n31139 , n31140 , n31141 , n31142 , n31143 , n31144 , n31145 , n31146 , n31147 , n31148 , n31149 , n31150 , n31151 , n31152 , n31153 , n31154 , n31155 , n31156 , n31157 , n31158 , n31159 , n31160 , n31161 , n31162 , n31163 , n31164 , n31165 , n31166 , n31167 , n31168 , n31169 , n31170 , n31171 , n31172 , n31173 , n31174 , n31175 , n31176 , n31177 , n31178 , n31179 , n31180 , n31181 , n31182 , n31183 , n31184 , n31185 , n31186 , n31187 , n31188 , n31189 , n31190 , n31191 , n31192 , n31193 , n31194 , n31195 , n31196 , n31197 , n31198 , n31199 , n31200 , n31201 , n31202 , n31203 , n31204 , n31205 , n31206 , n31207 , n31208 , n31209 , n31210 , n31211 , n31212 , n31213 , n31214 , n31215 , n31216 , n31217 , n31218 , n31219 , n31220 , n31221 , n31222 , n31223 , n31224 , n31225 , n31226 , n31227 , n31228 , n31229 , n31230 , n31231 , n31232 , n31233 , n31234 , n31235 , n31236 , n31237 , n31238 , n31239 , n31240 , n31241 , n31242 , n31243 , n31244 , n31245 , n31246 , n31247 , n31248 , n31249 , n31250 , n31251 , n31252 , n31253 , n31254 , n31255 , n31256 , n31257 , n31258 , n31259 , n31260 , n31261 , n31262 , n31263 , n31264 , n31265 , n31266 , n31267 , n31268 , n31269 , n31270 , n31271 , n31272 , n31273 , n31274 , n31275 , n31276 , n31277 , n31278 , n31279 , n31280 , n31281 , n31282 , n31283 , n31284 , n31285 , n31286 , n31287 , n31288 , n31289 , n31290 , n31291 , n31292 , n31293 , n31294 , n31295 , n31296 , n31297 , n31298 , n31299 , n31300 , n31301 , n31302 , n31303 , n31304 , n31305 , n31306 , n31307 , n31308 , n31309 , n31310 , n31311 , n31312 , n31313 , n31314 , n31315 , n31316 , n31317 , n31318 , n31319 , n31320 , n31321 , n31322 , n31323 , n31324 , n31325 , n31326 , n31327 , n31328 , n31329 , n31330 , n31331 , n31332 , n31333 , n31334 , n31335 , n31336 , n31337 , n31338 , n31339 , n31340 , n31341 , n31342 , n31343 , n31344 , n31345 , n31346 , n31347 , n31348 , n31349 , n31350 , n31351 , n31352 , n31353 , n31354 , n31355 , n31356 , n31357 , n31358 , n31359 , n31360 , n31361 , n31362 , n31363 , n31364 , n31365 , n31366 , n31367 , n31368 , n31369 , n31370 , n31371 , n31372 , n31373 , n31374 , n31375 , n31376 , n31377 , n31378 , n31379 , n31380 , n31381 , n31382 , n31383 , n31384 , n31385 , n31386 , n31387 , n31388 , n31389 , n31390 , n31391 , n31392 , n31393 , n31394 , n31395 , n31396 , n31397 , n31398 , n31399 , n31400 , n31401 , n31402 , n31403 , n31404 , n31405 , n31406 , n31407 , n31408 , n31409 , n31410 , n31411 , n31412 , n31413 , n31414 , n31415 , n31416 , n31417 , n31418 , n31419 , n31420 , n31421 , n31422 , n31423 , n31424 , n31425 , n31426 , n31427 , n31428 , n31429 , n31430 , n31431 , n31432 , n31433 , n31434 , n31435 , n31436 , n31437 , n31438 , n31439 , n31440 , n31441 , n31442 , n31443 , n31444 , n31445 , n31446 , n31447 , n31448 , n31449 , n31450 , n31451 , n31452 , n31453 , n31454 , n31455 , n31456 , n31457 , n31458 , n31459 , n31460 , n31461 , n31462 , n31463 , n31464 , n31465 , n31466 , n31467 , n31468 , n31469 , n31470 , n31471 , n31472 , n31473 , n31474 , n31475 , n31476 , n31477 , n31478 , n31479 , n31480 , n31481 , n31482 , n31483 , n31484 , n31485 , n31486 , n31487 , n31488 , n31489 , n31490 , n31491 , n31492 , n31493 , n31494 , n31495 , n31496 , n31497 , n31498 , n31499 , n31500 , n31501 , n31502 , n31503 , n31504 , n31505 , n31506 , n31507 , n31508 , n31509 , n31510 , n31511 , n31512 , n31513 , n31514 , n31515 , n31516 , n31517 , n31518 , n31519 , n31520 , n31521 , n31522 , n31523 , n31524 , n31525 , n31526 , n31527 , n31528 , n31529 , n31530 , n31531 , n31532 , n31533 , n31534 , n31535 , n31536 , n31537 , n31538 , n31539 , n31540 , n31541 , n31542 , n31543 , n31544 , n31545 , n31546 , n31547 , n31548 , n31549 , n31550 , n31551 , n31552 , n31553 , n31554 , n31555 , n31556 , n31557 , n31558 , n31559 , n31560 , n31561 , n31562 , n31563 , n31564 , n31565 , n31566 , n31567 , n31568 , n31569 , n31570 , n31571 , n31572 , n31573 , n31574 , n31575 , n31576 , n31577 , n31578 , n31579 , n31580 , n31581 , n31582 , n31583 , n31584 , n31585 , n31586 , n31587 , n31588 , n31589 , n31590 , n31591 , n31592 , n31593 , n31594 , n31595 , n31596 , n31597 , n31598 , n31599 , n31600 , n31601 , n31602 , n31603 , n31604 , n31605 , n31606 , n31607 , n31608 , n31609 , n31610 , n31611 , n31612 , n31613 , n31614 , n31615 , n31616 , n31617 , n31618 , n31619 , n31620 , n31621 , n31622 , n31623 , n31624 , n31625 , n31626 , n31627 , n31628 , n31629 , n31630 , n31631 , n31632 , n31633 , n31634 , n31635 , n31636 , n31637 , n31638 , n31639 , n31640 , n31641 , n31642 , n31643 , n31644 , n31645 , n31646 , n31647 , n31648 , n31649 , n31650 , n31651 , n31652 , n31653 , n31654 , n31655 , n31656 , n31657 , n31658 , n31659 , n31660 , n31661 , n31662 , n31663 , n31664 , n31665 , n31666 , n31667 , n31668 , n31669 , n31670 , n31671 , n31672 , n31673 , n31674 , n31675 , n31676 , n31677 , n31678 , n31679 , n31680 , n31681 , n31682 , n31683 , n31684 , n31685 , n31686 , n31687 , n31688 , n31689 , n31690 , n31691 , n31692 , n31693 , n31694 , n31695 , n31696 , n31697 , n31698 , n31699 , n31700 , n31701 , n31702 , n31703 , n31704 , n31705 , n31706 , n31707 , n31708 , n31709 , n31710 , n31711 , n31712 , n31713 , n31714 , n31715 , n31716 , n31717 , n31718 , n31719 , n31720 , n31721 , n31722 , n31723 , n31724 , n31725 , n31726 , n31727 , n31728 , n31729 , n31730 , n31731 , n31732 , n31733 , n31734 , n31735 , n31736 , n31737 , n31738 , n31739 , n31740 , n31741 , n31742 , n31743 , n31744 , n31745 , n31746 , n31747 , n31748 , n31749 , n31750 , n31751 , n31752 , n31753 , n31754 , n31755 , n31756 , n31757 , n31758 , n31759 , n31760 , n31761 , n31762 , n31763 , n31764 , n31765 , n31766 , n31767 , n31768 , n31769 , n31770 , n31771 , n31772 , n31773 , n31774 , n31775 , n31776 , n31777 , n31778 , n31779 , n31780 , n31781 , n31782 , n31783 , n31784 , n31785 , n31786 , n31787 , n31788 , n31789 , n31790 , n31791 , n31792 , n31793 , n31794 , n31795 , n31796 , n31797 , n31798 , n31799 , n31800 , n31801 , n31802 , n31803 , n31804 , n31805 , n31806 , n31807 , n31808 , n31809 , n31810 , n31811 , n31812 , n31813 , n31814 , n31815 , n31816 , n31817 , n31818 , n31819 , n31820 , n31821 , n31822 , n31823 , n31824 , n31825 , n31826 , n31827 , n31828 , n31829 , n31830 , n31831 , n31832 , n31833 , n31834 , n31835 , n31836 , n31837 , n31838 , n31839 , n31840 , n31841 , n31842 , n31843 , n31844 , n31845 , n31846 , n31847 , n31848 , n31849 , n31850 , n31851 , n31852 , n31853 , n31854 , n31855 , n31856 , n31857 , n31858 , n31859 , n31860 , n31861 , n31862 , n31863 , n31864 , n31865 , n31866 , n31867 , n31868 , n31869 , n31870 , n31871 , n31872 , n31873 , n31874 , n31875 , n31876 , n31877 , n31878 , n31879 , n31880 , n31881 , n31882 , n31883 , n31884 , n31885 , n31886 , n31887 , n31888 , n31889 , n31890 , n31891 , n31892 , n31893 , n31894 , n31895 , n31896 , n31897 , n31898 , n31899 , n31900 , n31901 , n31902 , n31903 , n31904 , n31905 , n31906 , n31907 , n31908 , n31909 , n31910 , n31911 , n31912 , n31913 , n31914 , n31915 , n31916 , n31917 , n31918 , n31919 , n31920 , n31921 , n31922 , n31923 , n31924 , n31925 , n31926 , n31927 , n31928 , n31929 , n31930 , n31931 , n31932 , n31933 , n31934 , n31935 , n31936 , n31937 , n31938 , n31939 , n31940 , n31941 , n31942 , n31943 , n31944 , n31945 , n31946 , n31947 , n31948 , n31949 , n31950 , n31951 , n31952 , n31953 , n31954 , n31955 , n31956 , n31957 , n31958 , n31959 , n31960 , n31961 , n31962 , n31963 , n31964 , n31965 , n31966 , n31967 , n31968 , n31969 , n31970 , n31971 , n31972 , n31973 , n31974 , n31975 , n31976 , n31977 , n31978 , n31979 , n31980 , n31981 , n31982 , n31983 , n31984 , n31985 , n31986 , n31987 , n31988 , n31989 , n31990 , n31991 , n31992 , n31993 , n31994 , n31995 , n31996 , n31997 , n31998 , n31999 , n32000 , n32001 , n32002 , n32003 , n32004 , n32005 , n32006 , n32007 , n32008 , n32009 , n32010 , n32011 , n32012 , n32013 , n32014 , n32015 , n32016 , n32017 , n32018 , n32019 , n32020 , n32021 , n32022 , n32023 , n32024 , n32025 , n32026 , n32027 , n32028 , n32029 , n32030 , n32031 , n32032 , n32033 , n32034 , n32035 , n32036 , n32037 , n32038 , n32039 , n32040 , n32041 , n32042 , n32043 , n32044 , n32045 , n32046 , n32047 , n32048 , n32049 , n32050 , n32051 , n32052 , n32053 , n32054 , n32055 , n32056 , n32057 , n32058 , n32059 , n32060 , n32061 , n32062 , n32063 , n32064 , n32065 , n32066 , n32067 , n32068 , n32069 , n32070 , n32071 , n32072 , n32073 , n32074 , n32075 , n32076 , n32077 , n32078 , n32079 , n32080 , n32081 , n32082 , n32083 , n32084 , n32085 , n32086 , n32087 , n32088 , n32089 , n32090 , n32091 , n32092 , n32093 , n32094 , n32095 , n32096 , n32097 , n32098 , n32099 , n32100 , n32101 , n32102 , n32103 , n32104 , n32105 , n32106 , n32107 , n32108 , n32109 , n32110 , n32111 , n32112 , n32113 , n32114 , n32115 , n32116 , n32117 , n32118 , n32119 , n32120 , n32121 , n32122 , n32123 , n32124 , n32125 , n32126 , n32127 , n32128 , n32129 , n32130 , n32131 , n32132 , n32133 , n32134 , n32135 , n32136 , n32137 , n32138 , n32139 , n32140 , n32141 , n32142 , n32143 , n32144 , n32145 , n32146 , n32147 , n32148 , n32149 , n32150 , n32151 , n32152 , n32153 , n32154 , n32155 , n32156 , n32157 , n32158 , n32159 , n32160 , n32161 , n32162 , n32163 , n32164 , n32165 , n32166 , n32167 , n32168 , n32169 , n32170 , n32171 , n32172 , n32173 , n32174 , n32175 , n32176 , n32177 , n32178 , n32179 , n32180 , n32181 , n32182 , n32183 , n32184 , n32185 , n32186 , n32187 , n32188 , n32189 , n32190 , n32191 , n32192 , n32193 , n32194 , n32195 , n32196 , n32197 , n32198 , n32199 , n32200 , n32201 , n32202 , n32203 , n32204 , n32205 , n32206 , n32207 , n32208 , n32209 , n32210 , n32211 , n32212 , n32213 , n32214 , n32215 , n32216 , n32217 , n32218 , n32219 , n32220 , n32221 , n32222 , n32223 , n32224 , n32225 , n32226 , n32227 , n32228 , n32229 , n32230 , n32231 , n32232 , n32233 , n32234 , n32235 , n32236 , n32237 , n32238 , n32239 , n32240 , n32241 , n32242 , n32243 , n32244 , n32245 , n32246 , n32247 , n32248 , n32249 , n32250 , n32251 , n32252 , n32253 , n32254 , n32255 , n32256 , n32257 , n32258 , n32259 , n32260 , n32261 , n32262 , n32263 , n32264 , n32265 , n32266 , n32267 , n32268 , n32269 , n32270 , n32271 , n32272 , n32273 , n32274 , n32275 , n32276 , n32277 , n32278 , n32279 , n32280 , n32281 , n32282 , n32283 , n32284 , n32285 , n32286 , n32287 , n32288 , n32289 , n32290 , n32291 , n32292 , n32293 , n32294 , n32295 , n32296 , n32297 , n32298 , n32299 , n32300 , n32301 , n32302 , n32303 , n32304 , n32305 , n32306 , n32307 , n32308 , n32309 , n32310 , n32311 , n32312 , n32313 , n32314 , n32315 , n32316 , n32317 , n32318 , n32319 , n32320 , n32321 , n32322 , n32323 , n32324 , n32325 , n32326 , n32327 , n32328 , n32329 , n32330 , n32331 , n32332 , n32333 , n32334 , n32335 , n32336 , n32337 , n32338 , n32339 , n32340 , n32341 , n32342 , n32343 , n32344 , n32345 , n32346 , n32347 , n32348 , n32349 , n32350 , n32351 , n32352 , n32353 , n32354 , n32355 , n32356 , n32357 , n32358 , n32359 , n32360 , n32361 , n32362 , n32363 , n32364 , n32365 , n32366 , n32367 , n32368 , n32369 , n32370 , n32371 , n32372 , n32373 , n32374 , n32375 , n32376 , n32377 , n32378 , n32379 , n32380 , n32381 , n32382 , n32383 , n32384 , n32385 , n32386 , n32387 , n32388 , n32389 , n32390 , n32391 , n32392 , n32393 , n32394 , n32395 , n32396 , n32397 , n32398 , n32399 , n32400 , n32401 , n32402 , n32403 , n32404 , n32405 , n32406 , n32407 , n32408 , n32409 , n32410 , n32411 , n32412 , n32413 , n32414 , n32415 , n32416 , n32417 , n32418 , n32419 , n32420 , n32421 , n32422 , n32423 , n32424 , n32425 , n32426 , n32427 , n32428 , n32429 , n32430 , n32431 , n32432 , n32433 , n32434 , n32435 , n32436 , n32437 , n32438 , n32439 , n32440 , n32441 , n32442 , n32443 , n32444 , n32445 , n32446 , n32447 , n32448 , n32449 , n32450 , n32451 , n32452 , n32453 , n32454 , n32455 , n32456 , n32457 , n32458 , n32459 , n32460 , n32461 , n32462 , n32463 , n32464 , n32465 , n32466 , n32467 , n32468 , n32469 , n32470 , n32471 , n32472 , n32473 , n32474 , n32475 , n32476 , n32477 , n32478 , n32479 , n32480 , n32481 , n32482 , n32483 , n32484 , n32485 , n32486 , n32487 , n32488 , n32489 , n32490 , n32491 , n32492 , n32493 , n32494 , n32495 , n32496 , n32497 , n32498 , n32499 , n32500 , n32501 , n32502 , n32503 , n32504 , n32505 , n32506 , n32507 , n32508 , n32509 , n32510 , n32511 , n32512 , n32513 , n32514 , n32515 , n32516 , n32517 , n32518 , n32519 , n32520 , n32521 , n32522 , n32523 , n32524 , n32525 , n32526 , n32527 , n32528 , n32529 , n32530 , n32531 , n32532 , n32533 , n32534 , n32535 , n32536 , n32537 , n32538 , n32539 , n32540 , n32541 , n32542 , n32543 , n32544 , n32545 , n32546 , n32547 , n32548 , n32549 , n32550 , n32551 , n32552 , n32553 , n32554 , n32555 , n32556 , n32557 , n32558 , n32559 , n32560 , n32561 , n32562 , n32563 , n32564 , n32565 , n32566 , n32567 , n32568 , n32569 , n32570 , n32571 , n32572 , n32573 , n32574 , n32575 , n32576 , n32577 , n32578 , n32579 , n32580 , n32581 , n32582 , n32583 , n32584 , n32585 , n32586 , n32587 , n32588 , n32589 , n32590 , n32591 , n32592 , n32593 , n32594 , n32595 , n32596 , n32597 , n32598 , n32599 , n32600 , n32601 , n32602 , n32603 , n32604 , n32605 , n32606 , n32607 , n32608 , n32609 , n32610 , n32611 , n32612 , n32613 , n32614 , n32615 , n32616 , n32617 , n32618 , n32619 , n32620 , n32621 , n32622 , n32623 , n32624 , n32625 , n32626 , n32627 , n32628 , n32629 , n32630 , n32631 , n32632 , n32633 , n32634 , n32635 , n32636 , n32637 , n32638 , n32639 , n32640 , n32641 , n32642 , n32643 , n32644 , n32645 , n32646 , n32647 , n32648 , n32649 , n32650 , n32651 , n32652 , n32653 , n32654 , n32655 , n32656 , n32657 , n32658 , n32659 , n32660 , n32661 , n32662 , n32663 , n32664 , n32665 , n32666 , n32667 , n32668 , n32669 , n32670 , n32671 , n32672 , n32673 , n32674 , n32675 , n32676 , n32677 , n32678 , n32679 , n32680 , n32681 , n32682 , n32683 , n32684 , n32685 , n32686 , n32687 , n32688 , n32689 , n32690 , n32691 , n32692 , n32693 , n32694 , n32695 , n32696 , n32697 , n32698 , n32699 , n32700 , n32701 , n32702 , n32703 , n32704 , n32705 , n32706 , n32707 , n32708 , n32709 , n32710 , n32711 , n32712 , n32713 , n32714 , n32715 , n32716 , n32717 , n32718 , n32719 , n32720 , n32721 , n32722 , n32723 , n32724 , n32725 , n32726 , n32727 , n32728 , n32729 , n32730 , n32731 , n32732 , n32733 , n32734 , n32735 , n32736 , n32737 , n32738 , n32739 , n32740 , n32741 , n32742 , n32743 , n32744 , n32745 , n32746 , n32747 , n32748 , n32749 , n32750 , n32751 , n32752 , n32753 , n32754 , n32755 , n32756 , n32757 , n32758 , n32759 , n32760 , n32761 , n32762 , n32763 , n32764 , n32765 , n32766 , n32767 , n32768 , n32769 , n32770 , n32771 , n32772 , n32773 , n32774 , n32775 , n32776 , n32777 , n32778 , n32779 , n32780 , n32781 , n32782 , n32783 , n32784 , n32785 , n32786 , n32787 , n32788 , n32789 , n32790 , n32791 , n32792 , n32793 , n32794 , n32795 , n32796 , n32797 , n32798 , n32799 , n32800 , n32801 , n32802 , n32803 , n32804 , n32805 , n32806 , n32807 , n32808 , n32809 , n32810 , n32811 , n32812 , n32813 , n32814 , n32815 , n32816 , n32817 , n32818 , n32819 , n32820 , n32821 , n32822 , n32823 , n32824 , n32825 , n32826 , n32827 , n32828 , n32829 , n32830 , n32831 , n32832 , n32833 , n32834 , n32835 , n32836 , n32837 , n32838 , n32839 , n32840 , n32841 , n32842 , n32843 , n32844 , n32845 , n32846 , n32847 , n32848 , n32849 , n32850 , n32851 , n32852 , n32853 , n32854 , n32855 , n32856 , n32857 , n32858 , n32859 , n32860 , n32861 , n32862 , n32863 , n32864 , n32865 , n32866 , n32867 , n32868 , n32869 , n32870 , n32871 , n32872 , n32873 , n32874 , n32875 , n32876 , n32877 , n32878 , n32879 , n32880 , n32881 , n32882 , n32883 , n32884 , n32885 , n32886 , n32887 , n32888 , n32889 , n32890 , n32891 , n32892 , n32893 , n32894 , n32895 , n32896 , n32897 , n32898 , n32899 , n32900 , n32901 , n32902 , n32903 , n32904 , n32905 , n32906 , n32907 , n32908 , n32909 , n32910 , n32911 , n32912 , n32913 , n32914 , n32915 , n32916 , n32917 , n32918 , n32919 , n32920 , n32921 , n32922 , n32923 , n32924 , n32925 , n32926 , n32927 , n32928 , n32929 , n32930 , n32931 , n32932 , n32933 , n32934 , n32935 , n32936 , n32937 , n32938 , n32939 , n32940 , n32941 , n32942 , n32943 , n32944 , n32945 , n32946 , n32947 , n32948 , n32949 , n32950 , n32951 , n32952 , n32953 , n32954 , n32955 , n32956 , n32957 , n32958 , n32959 , n32960 , n32961 , n32962 , n32963 , n32964 , n32965 , n32966 , n32967 , n32968 , n32969 , n32970 , n32971 , n32972 , n32973 , n32974 , n32975 , n32976 , n32977 , n32978 , n32979 , n32980 , n32981 , n32982 , n32983 , n32984 , n32985 , n32986 , n32987 , n32988 , n32989 , n32990 , n32991 , n32992 , n32993 , n32994 , n32995 , n32996 , n32997 , n32998 , n32999 , n33000 , n33001 , n33002 , n33003 , n33004 , n33005 , n33006 , n33007 , n33008 , n33009 , n33010 , n33011 , n33012 , n33013 , n33014 , n33015 , n33016 , n33017 , n33018 , n33019 , n33020 , n33021 , n33022 , n33023 , n33024 , n33025 , n33026 , n33027 , n33028 , n33029 , n33030 , n33031 , n33032 , n33033 , n33034 , n33035 , n33036 , n33037 , n33038 , n33039 , n33040 , n33041 , n33042 , n33043 , n33044 , n33045 , n33046 , n33047 , n33048 , n33049 , n33050 , n33051 , n33052 , n33053 , n33054 , n33055 , n33056 , n33057 , n33058 , n33059 , n33060 , n33061 , n33062 , n33063 , n33064 , n33065 , n33066 , n33067 , n33068 , n33069 , n33070 , n33071 , n33072 , n33073 , n33074 , n33075 , n33076 , n33077 , n33078 , n33079 , n33080 , n33081 , n33082 , n33083 , n33084 , n33085 , n33086 , n33087 , n33088 , n33089 , n33090 , n33091 , n33092 , n33093 , n33094 , n33095 , n33096 , n33097 , n33098 , n33099 , n33100 , n33101 , n33102 , n33103 , n33104 , n33105 , n33106 , n33107 , n33108 , n33109 , n33110 , n33111 , n33112 , n33113 , n33114 , n33115 , n33116 , n33117 , n33118 , n33119 , n33120 , n33121 , n33122 , n33123 , n33124 , n33125 , n33126 , n33127 , n33128 , n33129 , n33130 , n33131 , n33132 , n33133 , n33134 , n33135 , n33136 , n33137 , n33138 , n33139 , n33140 , n33141 , n33142 , n33143 , n33144 , n33145 , n33146 , n33147 , n33148 , n33149 , n33150 , n33151 , n33152 , n33153 , n33154 , n33155 , n33156 , n33157 , n33158 , n33159 , n33160 , n33161 , n33162 , n33163 , n33164 , n33165 , n33166 , n33167 , n33168 , n33169 , n33170 , n33171 , n33172 , n33173 , n33174 , n33175 , n33176 , n33177 , n33178 , n33179 , n33180 , n33181 , n33182 , n33183 , n33184 , n33185 , n33186 , n33187 , n33188 , n33189 , n33190 , n33191 , n33192 , n33193 , n33194 , n33195 , n33196 , n33197 , n33198 , n33199 , n33200 , n33201 , n33202 , n33203 , n33204 , n33205 , n33206 , n33207 , n33208 , n33209 , n33210 , n33211 , n33212 , n33213 , n33214 , n33215 , n33216 , n33217 , n33218 , n33219 , n33220 , n33221 , n33222 , n33223 , n33224 , n33225 , n33226 , n33227 , n33228 , n33229 , n33230 , n33231 , n33232 , n33233 , n33234 , n33235 , n33236 , n33237 , n33238 , n33239 , n33240 , n33241 , n33242 , n33243 , n33244 , n33245 , n33246 , n33247 , n33248 , n33249 , n33250 , n33251 , n33252 , n33253 , n33254 , n33255 , n33256 , n33257 , n33258 , n33259 , n33260 , n33261 , n33262 , n33263 , n33264 , n33265 , n33266 , n33267 , n33268 , n33269 , n33270 , n33271 , n33272 , n33273 , n33274 , n33275 , n33276 , n33277 , n33278 , n33279 , n33280 , n33281 , n33282 , n33283 , n33284 , n33285 , n33286 , n33287 , n33288 , n33289 , n33290 , n33291 , n33292 , n33293 , n33294 , n33295 , n33296 , n33297 , n33298 , n33299 , n33300 , n33301 , n33302 , n33303 , n33304 , n33305 , n33306 , n33307 , n33308 , n33309 , n33310 , n33311 , n33312 , n33313 , n33314 , n33315 , n33316 , n33317 , n33318 , n33319 , n33320 , n33321 , n33322 , n33323 , n33324 , n33325 , n33326 , n33327 , n33328 , n33329 , n33330 , n33331 , n33332 , n33333 , n33334 , n33335 , n33336 , n33337 , n33338 , n33339 , n33340 , n33341 , n33342 , n33343 , n33344 , n33345 , n33346 , n33347 , n33348 , n33349 , n33350 , n33351 , n33352 , n33353 , n33354 , n33355 , n33356 , n33357 , n33358 , n33359 , n33360 , n33361 , n33362 , n33363 , n33364 , n33365 , n33366 , n33367 , n33368 , n33369 , n33370 , n33371 , n33372 , n33373 , n33374 , n33375 , n33376 , n33377 , n33378 , n33379 , n33380 , n33381 , n33382 , n33383 , n33384 , n33385 , n33386 , n33387 , n33388 , n33389 , n33390 , n33391 , n33392 , n33393 , n33394 , n33395 , n33396 , n33397 , n33398 , n33399 , n33400 , n33401 , n33402 , n33403 , n33404 , n33405 , n33406 , n33407 , n33408 , n33409 , n33410 , n33411 , n33412 , n33413 , n33414 , n33415 , n33416 , n33417 , n33418 , n33419 , n33420 , n33421 , n33422 , n33423 , n33424 , n33425 , n33426 , n33427 , n33428 , n33429 , n33430 , n33431 , n33432 , n33433 , n33434 , n33435 , n33436 , n33437 , n33438 , n33439 , n33440 , n33441 , n33442 , n33443 , n33444 , n33445 , n33446 , n33447 , n33448 , n33449 , n33450 , n33451 , n33452 , n33453 , n33454 , n33455 , n33456 , n33457 , n33458 , n33459 , n33460 , n33461 , n33462 , n33463 , n33464 , n33465 , n33466 , n33467 , n33468 , n33469 , n33470 , n33471 , n33472 , n33473 , n33474 , n33475 , n33476 , n33477 , n33478 , n33479 , n33480 , n33481 , n33482 , n33483 , n33484 , n33485 , n33486 , n33487 , n33488 , n33489 , n33490 , n33491 , n33492 , n33493 , n33494 , n33495 , n33496 , n33497 , n33498 , n33499 , n33500 , n33501 , n33502 , n33503 , n33504 , n33505 , n33506 , n33507 , n33508 , n33509 , n33510 , n33511 , n33512 , n33513 , n33514 , n33515 , n33516 , n33517 , n33518 , n33519 , n33520 , n33521 , n33522 , n33523 , n33524 , n33525 , n33526 , n33527 , n33528 , n33529 , n33530 , n33531 , n33532 , n33533 , n33534 , n33535 , n33536 , n33537 , n33538 , n33539 , n33540 , n33541 , n33542 , n33543 , n33544 , n33545 , n33546 , n33547 , n33548 , n33549 , n33550 , n33551 , n33552 , n33553 , n33554 , n33555 , n33556 , n33557 , n33558 , n33559 , n33560 , n33561 , n33562 , n33563 , n33564 , n33565 , n33566 , n33567 , n33568 , n33569 , n33570 , n33571 , n33572 , n33573 , n33574 , n33575 , n33576 , n33577 , n33578 , n33579 , n33580 , n33581 , n33582 , n33583 , n33584 , n33585 , n33586 , n33587 , n33588 , n33589 , n33590 , n33591 , n33592 , n33593 , n33594 , n33595 , n33596 , n33597 , n33598 , n33599 , n33600 , n33601 , n33602 , n33603 , n33604 , n33605 , n33606 , n33607 , n33608 , n33609 , n33610 , n33611 , n33612 , n33613 , n33614 , n33615 , n33616 , n33617 , n33618 , n33619 , n33620 , n33621 , n33622 , n33623 , n33624 , n33625 , n33626 , n33627 , n33628 , n33629 , n33630 , n33631 , n33632 , n33633 , n33634 , n33635 , n33636 , n33637 , n33638 , n33639 , n33640 , n33641 , n33642 , n33643 , n33644 , n33645 , n33646 , n33647 , n33648 , n33649 , n33650 , n33651 , n33652 , n33653 , n33654 , n33655 , n33656 , n33657 , n33658 , n33659 , n33660 , n33661 , n33662 , n33663 , n33664 , n33665 , n33666 , n33667 , n33668 , n33669 , n33670 , n33671 , n33672 , n33673 , n33674 , n33675 , n33676 , n33677 , n33678 , n33679 , n33680 , n33681 , n33682 , n33683 , n33684 , n33685 , n33686 , n33687 , n33688 , n33689 , n33690 , n33691 , n33692 , n33693 , n33694 , n33695 , n33696 , n33697 , n33698 , n33699 , n33700 , n33701 , n33702 , n33703 , n33704 , n33705 , n33706 , n33707 , n33708 , n33709 , n33710 , n33711 , n33712 , n33713 , n33714 , n33715 , n33716 , n33717 , n33718 , n33719 , n33720 , n33721 , n33722 , n33723 , n33724 , n33725 , n33726 , n33727 , n33728 , n33729 , n33730 , n33731 , n33732 , n33733 , n33734 , n33735 , n33736 , n33737 , n33738 , n33739 , n33740 , n33741 , n33742 , n33743 , n33744 , n33745 , n33746 , n33747 , n33748 , n33749 , n33750 , n33751 , n33752 , n33753 , n33754 , n33755 , n33756 , n33757 , n33758 , n33759 , n33760 , n33761 , n33762 , n33763 , n33764 , n33765 , n33766 , n33767 , n33768 , n33769 , n33770 , n33771 , n33772 , n33773 , n33774 , n33775 , n33776 , n33777 , n33778 , n33779 , n33780 , n33781 , n33782 , n33783 , n33784 , n33785 , n33786 , n33787 , n33788 , n33789 , n33790 , n33791 , n33792 , n33793 , n33794 , n33795 , n33796 , n33797 , n33798 , n33799 , n33800 , n33801 , n33802 , n33803 , n33804 , n33805 , n33806 , n33807 , n33808 , n33809 , n33810 , n33811 , n33812 , n33813 , n33814 , n33815 , n33816 , n33817 , n33818 , n33819 , n33820 , n33821 , n33822 , n33823 , n33824 , n33825 , n33826 , n33827 , n33828 , n33829 , n33830 , n33831 , n33832 , n33833 , n33834 , n33835 , n33836 , n33837 , n33838 , n33839 , n33840 , n33841 , n33842 , n33843 , n33844 , n33845 , n33846 , n33847 , n33848 , n33849 , n33850 , n33851 , n33852 , n33853 , n33854 , n33855 , n33856 , n33857 , n33858 , n33859 , n33860 , n33861 , n33862 , n33863 , n33864 , n33865 , n33866 , n33867 , n33868 , n33869 , n33870 , n33871 , n33872 , n33873 , n33874 , n33875 , n33876 , n33877 , n33878 , n33879 , n33880 , n33881 , n33882 , n33883 , n33884 , n33885 , n33886 , n33887 , n33888 , n33889 , n33890 , n33891 , n33892 , n33893 , n33894 , n33895 , n33896 , n33897 , n33898 , n33899 , n33900 , n33901 , n33902 , n33903 , n33904 , n33905 , n33906 , n33907 , n33908 , n33909 , n33910 , n33911 , n33912 , n33913 , n33914 , n33915 , n33916 , n33917 , n33918 , n33919 , n33920 , n33921 , n33922 , n33923 , n33924 , n33925 , n33926 , n33927 , n33928 , n33929 , n33930 , n33931 , n33932 , n33933 , n33934 , n33935 , n33936 , n33937 , n33938 , n33939 , n33940 , n33941 , n33942 , n33943 , n33944 , n33945 , n33946 , n33947 , n33948 , n33949 , n33950 , n33951 , n33952 , n33953 , n33954 , n33955 , n33956 , n33957 , n33958 , n33959 , n33960 , n33961 , n33962 , n33963 , n33964 , n33965 , n33966 , n33967 , n33968 , n33969 , n33970 , n33971 , n33972 , n33973 , n33974 , n33975 , n33976 , n33977 , n33978 , n33979 , n33980 , n33981 , n33982 , n33983 , n33984 , n33985 , n33986 , n33987 , n33988 , n33989 , n33990 , n33991 , n33992 , n33993 , n33994 , n33995 , n33996 , n33997 , n33998 , n33999 , n34000 , n34001 , n34002 , n34003 , n34004 , n34005 , n34006 , n34007 , n34008 , n34009 , n34010 , n34011 , n34012 , n34013 , n34014 , n34015 , n34016 , n34017 , n34018 , n34019 , n34020 , n34021 , n34022 , n34023 , n34024 , n34025 , n34026 , n34027 , n34028 , n34029 , n34030 , n34031 , n34032 , n34033 , n34034 , n34035 , n34036 , n34037 , n34038 , n34039 , n34040 , n34041 , n34042 , n34043 , n34044 , n34045 , n34046 , n34047 , n34048 , n34049 , n34050 , n34051 , n34052 , n34053 , n34054 , n34055 , n34056 , n34057 , n34058 , n34059 , n34060 , n34061 , n34062 , n34063 , n34064 , n34065 , n34066 , n34067 , n34068 , n34069 , n34070 , n34071 , n34072 , n34073 , n34074 , n34075 , n34076 , n34077 , n34078 , n34079 , n34080 , n34081 , n34082 , n34083 , n34084 , n34085 , n34086 , n34087 , n34088 , n34089 , n34090 , n34091 , n34092 , n34093 , n34094 , n34095 , n34096 , n34097 , n34098 , n34099 , n34100 , n34101 , n34102 , n34103 , n34104 , n34105 , n34106 , n34107 , n34108 , n34109 , n34110 , n34111 , n34112 , n34113 , n34114 , n34115 , n34116 , n34117 , n34118 , n34119 , n34120 , n34121 , n34122 , n34123 , n34124 , n34125 , n34126 , n34127 , n34128 , n34129 , n34130 , n34131 , n34132 , n34133 , n34134 , n34135 , n34136 , n34137 , n34138 , n34139 , n34140 , n34141 , n34142 , n34143 , n34144 , n34145 , n34146 , n34147 , n34148 , n34149 , n34150 , n34151 , n34152 , n34153 , n34154 , n34155 , n34156 , n34157 , n34158 , n34159 , n34160 , n34161 , n34162 , n34163 , n34164 , n34165 , n34166 , n34167 , n34168 , n34169 , n34170 , n34171 , n34172 , n34173 , n34174 , n34175 , n34176 , n34177 , n34178 , n34179 , n34180 , n34181 , n34182 , n34183 , n34184 , n34185 , n34186 , n34187 , n34188 , n34189 , n34190 , n34191 , n34192 , n34193 , n34194 , n34195 , n34196 , n34197 , n34198 , n34199 , n34200 , n34201 , n34202 , n34203 , n34204 , n34205 , n34206 , n34207 , n34208 , n34209 , n34210 , n34211 , n34212 , n34213 , n34214 , n34215 , n34216 , n34217 , n34218 , n34219 , n34220 , n34221 , n34222 , n34223 , n34224 , n34225 , n34226 , n34227 , n34228 , n34229 , n34230 , n34231 , n34232 , n34233 , n34234 , n34235 , n34236 , n34237 , n34238 , n34239 , n34240 , n34241 , n34242 , n34243 , n34244 , n34245 , n34246 , n34247 , n34248 , n34249 , n34250 , n34251 , n34252 , n34253 , n34254 , n34255 , n34256 , n34257 , n34258 , n34259 , n34260 , n34261 , n34262 , n34263 , n34264 , n34265 , n34266 , n34267 , n34268 , n34269 , n34270 , n34271 , n34272 , n34273 , n34274 , n34275 , n34276 , n34277 , n34278 , n34279 , n34280 , n34281 , n34282 , n34283 , n34284 , n34285 , n34286 , n34287 , n34288 , n34289 , n34290 , n34291 , n34292 , n34293 , n34294 , n34295 , n34296 , n34297 , n34298 , n34299 , n34300 , n34301 , n34302 , n34303 , n34304 , n34305 , n34306 , n34307 , n34308 , n34309 , n34310 , n34311 , n34312 , n34313 , n34314 , n34315 , n34316 , n34317 , n34318 , n34319 , n34320 , n34321 , n34322 , n34323 , n34324 , n34325 , n34326 , n34327 , n34328 , n34329 , n34330 , n34331 , n34332 , n34333 , n34334 , n34335 , n34336 , n34337 , n34338 , n34339 , n34340 , n34341 , n34342 , n34343 , n34344 , n34345 , n34346 , n34347 , n34348 , n34349 , n34350 , n34351 , n34352 , n34353 , n34354 , n34355 , n34356 , n34357 , n34358 , n34359 , n34360 , n34361 , n34362 , n34363 , n34364 , n34365 , n34366 , n34367 , n34368 , n34369 , n34370 , n34371 , n34372 , n34373 , n34374 , n34375 , n34376 , n34377 , n34378 , n34379 , n34380 , n34381 , n34382 , n34383 , n34384 , n34385 , n34386 , n34387 , n34388 , n34389 , n34390 , n34391 , n34392 , n34393 , n34394 , n34395 , n34396 , n34397 , n34398 , n34399 , n34400 , n34401 , n34402 , n34403 , n34404 , n34405 , n34406 , n34407 , n34408 , n34409 , n34410 , n34411 , n34412 , n34413 , n34414 , n34415 , n34416 , n34417 , n34418 , n34419 , n34420 , n34421 , n34422 , n34423 , n34424 , n34425 , n34426 , n34427 , n34428 , n34429 , n34430 , n34431 , n34432 , n34433 , n34434 , n34435 , n34436 , n34437 , n34438 , n34439 , n34440 , n34441 , n34442 , n34443 , n34444 , n34445 , n34446 , n34447 , n34448 , n34449 , n34450 , n34451 , n34452 , n34453 , n34454 , n34455 , n34456 , n34457 , n34458 , n34459 , n34460 , n34461 , n34462 , n34463 , n34464 , n34465 , n34466 , n34467 , n34468 , n34469 , n34470 , n34471 , n34472 , n34473 , n34474 , n34475 , n34476 , n34477 , n34478 , n34479 , n34480 , n34481 , n34482 , n34483 , n34484 , n34485 , n34486 , n34487 , n34488 , n34489 , n34490 , n34491 , n34492 , n34493 , n34494 , n34495 , n34496 , n34497 , n34498 , n34499 , n34500 , n34501 , n34502 , n34503 , n34504 , n34505 , n34506 , n34507 , n34508 , n34509 , n34510 , n34511 , n34512 , n34513 , n34514 , n34515 , n34516 , n34517 , n34518 , n34519 , n34520 , n34521 , n34522 , n34523 , n34524 , n34525 , n34526 , n34527 , n34528 , n34529 , n34530 , n34531 , n34532 , n34533 , n34534 , n34535 , n34536 , n34537 , n34538 , n34539 , n34540 , n34541 , n34542 , n34543 , n34544 , n34545 , n34546 , n34547 , n34548 , n34549 , n34550 , n34551 , n34552 , n34553 , n34554 , n34555 , n34556 , n34557 , n34558 , n34559 , n34560 , n34561 , n34562 , n34563 , n34564 , n34565 , n34566 , n34567 , n34568 , n34569 , n34570 , n34571 , n34572 , n34573 , n34574 , n34575 , n34576 , n34577 , n34578 , n34579 , n34580 , n34581 , n34582 , n34583 , n34584 , n34585 , n34586 , n34587 , n34588 , n34589 , n34590 , n34591 , n34592 , n34593 , n34594 , n34595 , n34596 , n34597 , n34598 , n34599 , n34600 , n34601 , n34602 , n34603 , n34604 , n34605 , n34606 , n34607 , n34608 , n34609 , n34610 , n34611 , n34612 , n34613 , n34614 , n34615 , n34616 , n34617 , n34618 , n34619 , n34620 , n34621 , n34622 , n34623 , n34624 , n34625 , n34626 , n34627 , n34628 , n34629 , n34630 , n34631 , n34632 , n34633 , n34634 , n34635 , n34636 , n34637 , n34638 , n34639 , n34640 , n34641 , n34642 , n34643 , n34644 , n34645 , n34646 , n34647 , n34648 , n34649 , n34650 , n34651 , n34652 , n34653 , n34654 , n34655 , n34656 , n34657 , n34658 , n34659 , n34660 , n34661 , n34662 , n34663 , n34664 , n34665 , n34666 , n34667 , n34668 , n34669 , n34670 , n34671 , n34672 , n34673 , n34674 , n34675 , n34676 , n34677 , n34678 , n34679 , n34680 , n34681 , n34682 , n34683 , n34684 , n34685 , n34686 , n34687 , n34688 , n34689 , n34690 , n34691 , n34692 , n34693 , n34694 , n34695 , n34696 , n34697 , n34698 , n34699 , n34700 , n34701 , n34702 , n34703 , n34704 , n34705 , n34706 , n34707 , n34708 , n34709 , n34710 , n34711 , n34712 , n34713 , n34714 , n34715 , n34716 , n34717 , n34718 , n34719 , n34720 , n34721 , n34722 , n34723 , n34724 , n34725 , n34726 , n34727 , n34728 , n34729 , n34730 , n34731 , n34732 , n34733 , n34734 , n34735 , n34736 , n34737 , n34738 , n34739 , n34740 , n34741 , n34742 , n34743 , n34744 , n34745 , n34746 , n34747 , n34748 , n34749 , n34750 , n34751 , n34752 , n34753 , n34754 , n34755 , n34756 , n34757 , n34758 , n34759 , n34760 , n34761 , n34762 , n34763 , n34764 , n34765 , n34766 , n34767 , n34768 , n34769 , n34770 , n34771 , n34772 , n34773 , n34774 , n34775 , n34776 , n34777 , n34778 , n34779 , n34780 , n34781 , n34782 , n34783 , n34784 , n34785 , n34786 , n34787 , n34788 , n34789 , n34790 , n34791 , n34792 , n34793 , n34794 , n34795 , n34796 , n34797 , n34798 , n34799 , n34800 , n34801 , n34802 , n34803 , n34804 , n34805 , n34806 , n34807 , n34808 , n34809 , n34810 , n34811 , n34812 , n34813 , n34814 , n34815 , n34816 , n34817 , n34818 , n34819 , n34820 , n34821 , n34822 , n34823 , n34824 , n34825 , n34826 , n34827 , n34828 , n34829 , n34830 , n34831 , n34832 , n34833 , n34834 , n34835 , n34836 , n34837 , n34838 , n34839 , n34840 , n34841 , n34842 , n34843 , n34844 , n34845 , n34846 , n34847 , n34848 , n34849 , n34850 , n34851 , n34852 , n34853 , n34854 , n34855 , n34856 , n34857 , n34858 , n34859 , n34860 , n34861 , n34862 , n34863 , n34864 , n34865 , n34866 , n34867 , n34868 , n34869 , n34870 , n34871 , n34872 , n34873 , n34874 , n34875 , n34876 , n34877 , n34878 , n34879 , n34880 , n34881 , n34882 , n34883 , n34884 , n34885 , n34886 , n34887 , n34888 , n34889 , n34890 , n34891 , n34892 , n34893 , n34894 , n34895 , n34896 , n34897 , n34898 , n34899 , n34900 , n34901 , n34902 , n34903 , n34904 , n34905 , n34906 , n34907 , n34908 , n34909 , n34910 , n34911 , n34912 , n34913 , n34914 , n34915 , n34916 , n34917 , n34918 , n34919 , n34920 , n34921 , n34922 , n34923 , n34924 , n34925 , n34926 , n34927 , n34928 , n34929 , n34930 , n34931 , n34932 , n34933 , n34934 , n34935 , n34936 , n34937 , n34938 , n34939 , n34940 , n34941 , n34942 , n34943 , n34944 , n34945 , n34946 , n34947 , n34948 , n34949 , n34950 , n34951 , n34952 , n34953 , n34954 , n34955 , n34956 , n34957 , n34958 , n34959 , n34960 , n34961 , n34962 , n34963 , n34964 , n34965 , n34966 , n34967 , n34968 , n34969 , n34970 , n34971 , n34972 , n34973 , n34974 , n34975 , n34976 , n34977 , n34978 , n34979 , n34980 , n34981 , n34982 , n34983 , n34984 , n34985 , n34986 , n34987 , n34988 , n34989 , n34990 , n34991 , n34992 , n34993 , n34994 , n34995 , n34996 , n34997 , n34998 , n34999 , n35000 , n35001 , n35002 , n35003 , n35004 , n35005 , n35006 , n35007 , n35008 , n35009 , n35010 , n35011 , n35012 , n35013 , n35014 , n35015 , n35016 , n35017 , n35018 , n35019 , n35020 , n35021 , n35022 , n35023 , n35024 , n35025 , n35026 , n35027 , n35028 , n35029 , n35030 , n35031 , n35032 , n35033 , n35034 , n35035 , n35036 , n35037 , n35038 , n35039 , n35040 , n35041 , n35042 , n35043 , n35044 , n35045 , n35046 , n35047 , n35048 , n35049 , n35050 , n35051 , n35052 , n35053 , n35054 , n35055 , n35056 , n35057 , n35058 , n35059 , n35060 , n35061 , n35062 , n35063 , n35064 , n35065 , n35066 , n35067 , n35068 , n35069 , n35070 , n35071 , n35072 , n35073 , n35074 , n35075 , n35076 , n35077 , n35078 , n35079 , n35080 , n35081 , n35082 , n35083 , n35084 , n35085 , n35086 , n35087 , n35088 , n35089 , n35090 , n35091 , n35092 , n35093 , n35094 , n35095 , n35096 , n35097 , n35098 , n35099 , n35100 , n35101 , n35102 , n35103 , n35104 , n35105 , n35106 , n35107 , n35108 , n35109 , n35110 , n35111 , n35112 , n35113 , n35114 , n35115 , n35116 , n35117 , n35118 , n35119 , n35120 , n35121 , n35122 , n35123 , n35124 , n35125 , n35126 , n35127 , n35128 , n35129 , n35130 , n35131 , n35132 , n35133 , n35134 , n35135 , n35136 , n35137 , n35138 , n35139 , n35140 , n35141 , n35142 , n35143 , n35144 , n35145 , n35146 , n35147 , n35148 , n35149 , n35150 , n35151 , n35152 , n35153 , n35154 , n35155 , n35156 , n35157 , n35158 , n35159 , n35160 , n35161 , n35162 , n35163 , n35164 , n35165 , n35166 , n35167 , n35168 , n35169 , n35170 , n35171 , n35172 , n35173 , n35174 , n35175 , n35176 , n35177 , n35178 , n35179 , n35180 , n35181 , n35182 , n35183 , n35184 , n35185 , n35186 , n35187 , n35188 , n35189 , n35190 , n35191 , n35192 , n35193 , n35194 , n35195 , n35196 , n35197 , n35198 , n35199 , n35200 , n35201 , n35202 , n35203 , n35204 , n35205 , n35206 , n35207 , n35208 , n35209 , n35210 , n35211 , n35212 , n35213 , n35214 , n35215 , n35216 , n35217 , n35218 , n35219 , n35220 , n35221 , n35222 , n35223 , n35224 , n35225 , n35226 , n35227 , n35228 , n35229 , n35230 , n35231 , n35232 , n35233 , n35234 , n35235 , n35236 , n35237 , n35238 , n35239 , n35240 , n35241 , n35242 , n35243 , n35244 , n35245 , n35246 , n35247 , n35248 , n35249 , n35250 , n35251 , n35252 , n35253 , n35254 , n35255 , n35256 , n35257 , n35258 , n35259 , n35260 , n35261 , n35262 , n35263 , n35264 , n35265 , n35266 , n35267 , n35268 , n35269 , n35270 , n35271 , n35272 , n35273 , n35274 , n35275 , n35276 , n35277 , n35278 , n35279 , n35280 , n35281 , n35282 , n35283 , n35284 , n35285 , n35286 , n35287 , n35288 , n35289 , n35290 , n35291 , n35292 , n35293 , n35294 , n35295 , n35296 , n35297 , n35298 , n35299 , n35300 , n35301 , n35302 , n35303 , n35304 , n35305 , n35306 , n35307 , n35308 , n35309 , n35310 , n35311 , n35312 , n35313 , n35314 , n35315 , n35316 , n35317 , n35318 , n35319 , n35320 , n35321 , n35322 , n35323 , n35324 , n35325 , n35326 , n35327 , n35328 , n35329 , n35330 , n35331 , n35332 , n35333 , n35334 , n35335 , n35336 , n35337 , n35338 , n35339 , n35340 , n35341 , n35342 , n35343 , n35344 , n35345 , n35346 , n35347 , n35348 , n35349 , n35350 , n35351 , n35352 , n35353 , n35354 , n35355 , n35356 , n35357 , n35358 , n35359 , n35360 , n35361 , n35362 , n35363 , n35364 , n35365 , n35366 , n35367 , n35368 , n35369 , n35370 , n35371 , n35372 , n35373 , n35374 , n35375 , n35376 , n35377 , n35378 , n35379 , n35380 , n35381 , n35382 , n35383 , n35384 , n35385 , n35386 , n35387 , n35388 , n35389 , n35390 , n35391 , n35392 , n35393 , n35394 , n35395 , n35396 , n35397 , n35398 , n35399 , n35400 , n35401 , n35402 , n35403 , n35404 , n35405 , n35406 , n35407 , n35408 , n35409 , n35410 , n35411 , n35412 , n35413 , n35414 , n35415 , n35416 , n35417 , n35418 , n35419 , n35420 , n35421 , n35422 , n35423 , n35424 , n35425 , n35426 , n35427 , n35428 , n35429 , n35430 , n35431 , n35432 , n35433 , n35434 , n35435 , n35436 , n35437 , n35438 , n35439 , n35440 , n35441 , n35442 , n35443 , n35444 , n35445 , n35446 , n35447 , n35448 , n35449 , n35450 , n35451 , n35452 , n35453 , n35454 , n35455 , n35456 , n35457 , n35458 , n35459 , n35460 , n35461 , n35462 , n35463 , n35464 , n35465 , n35466 , n35467 , n35468 , n35469 , n35470 , n35471 , n35472 , n35473 , n35474 , n35475 , n35476 , n35477 , n35478 , n35479 , n35480 , n35481 , n35482 , n35483 , n35484 , n35485 , n35486 , n35487 , n35488 , n35489 , n35490 , n35491 , n35492 , n35493 , n35494 , n35495 , n35496 , n35497 , n35498 , n35499 , n35500 , n35501 , n35502 , n35503 , n35504 , n35505 , n35506 , n35507 , n35508 , n35509 , n35510 , n35511 , n35512 , n35513 , n35514 , n35515 , n35516 , n35517 , n35518 , n35519 , n35520 , n35521 , n35522 , n35523 , n35524 , n35525 , n35526 , n35527 , n35528 , n35529 , n35530 , n35531 , n35532 , n35533 , n35534 , n35535 , n35536 , n35537 , n35538 , n35539 , n35540 , n35541 , n35542 , n35543 , n35544 , n35545 , n35546 , n35547 , n35548 , n35549 , n35550 , n35551 , n35552 , n35553 , n35554 , n35555 , n35556 , n35557 , n35558 , n35559 , n35560 , n35561 , n35562 , n35563 , n35564 , n35565 , n35566 , n35567 , n35568 , n35569 , n35570 , n35571 , n35572 , n35573 , n35574 , n35575 , n35576 , n35577 , n35578 , n35579 , n35580 , n35581 , n35582 , n35583 , n35584 , n35585 , n35586 , n35587 , n35588 , n35589 , n35590 , n35591 , n35592 , n35593 , n35594 , n35595 , n35596 , n35597 , n35598 , n35599 , n35600 , n35601 , n35602 , n35603 , n35604 , n35605 , n35606 , n35607 , n35608 , n35609 , n35610 , n35611 , n35612 , n35613 , n35614 , n35615 , n35616 , n35617 , n35618 , n35619 , n35620 , n35621 , n35622 , n35623 , n35624 , n35625 , n35626 , n35627 , n35628 , n35629 , n35630 , n35631 , n35632 , n35633 , n35634 , n35635 , n35636 , n35637 , n35638 , n35639 , n35640 , n35641 , n35642 , n35643 , n35644 , n35645 , n35646 , n35647 , n35648 , n35649 , n35650 , n35651 , n35652 , n35653 , n35654 , n35655 , n35656 , n35657 , n35658 , n35659 , n35660 , n35661 , n35662 , n35663 , n35664 , n35665 , n35666 , n35667 , n35668 , n35669 , n35670 , n35671 , n35672 , n35673 , n35674 , n35675 , n35676 , n35677 , n35678 , n35679 , n35680 , n35681 , n35682 , n35683 , n35684 , n35685 , n35686 , n35687 , n35688 , n35689 , n35690 , n35691 , n35692 , n35693 , n35694 , n35695 , n35696 , n35697 , n35698 , n35699 , n35700 , n35701 , n35702 , n35703 , n35704 , n35705 , n35706 , n35707 , n35708 , n35709 , n35710 , n35711 , n35712 , n35713 , n35714 , n35715 , n35716 , n35717 , n35718 , n35719 , n35720 , n35721 , n35722 , n35723 , n35724 , n35725 , n35726 , n35727 , n35728 , n35729 , n35730 , n35731 , n35732 , n35733 , n35734 , n35735 , n35736 , n35737 , n35738 , n35739 , n35740 , n35741 , n35742 , n35743 , n35744 , n35745 , n35746 , n35747 , n35748 , n35749 , n35750 , n35751 , n35752 , n35753 , n35754 , n35755 , n35756 , n35757 , n35758 , n35759 , n35760 , n35761 , n35762 , n35763 , n35764 , n35765 , n35766 , n35767 , n35768 , n35769 , n35770 , n35771 , n35772 , n35773 , n35774 , n35775 , n35776 , n35777 , n35778 , n35779 , n35780 , n35781 , n35782 , n35783 , n35784 , n35785 , n35786 , n35787 , n35788 , n35789 , n35790 , n35791 , n35792 , n35793 , n35794 , n35795 , n35796 , n35797 , n35798 , n35799 , n35800 , n35801 , n35802 , n35803 , n35804 , n35805 , n35806 , n35807 , n35808 , n35809 , n35810 , n35811 , n35812 , n35813 , n35814 , n35815 , n35816 , n35817 , n35818 , n35819 , n35820 , n35821 , n35822 , n35823 , n35824 , n35825 , n35826 , n35827 , n35828 , n35829 , n35830 , n35831 , n35832 , n35833 , n35834 , n35835 , n35836 , n35837 , n35838 , n35839 , n35840 , n35841 , n35842 , n35843 , n35844 , n35845 , n35846 , n35847 , n35848 , n35849 , n35850 , n35851 , n35852 , n35853 , n35854 , n35855 , n35856 , n35857 , n35858 , n35859 , n35860 , n35861 , n35862 , n35863 , n35864 , n35865 , n35866 , n35867 , n35868 , n35869 , n35870 , n35871 , n35872 , n35873 , n35874 , n35875 , n35876 , n35877 , n35878 , n35879 , n35880 , n35881 , n35882 , n35883 , n35884 , n35885 , n35886 , n35887 , n35888 , n35889 , n35890 , n35891 , n35892 , n35893 , n35894 , n35895 , n35896 , n35897 , n35898 , n35899 , n35900 , n35901 , n35902 , n35903 , n35904 , n35905 , n35906 , n35907 , n35908 , n35909 , n35910 , n35911 , n35912 , n35913 , n35914 , n35915 , n35916 , n35917 , n35918 , n35919 , n35920 , n35921 , n35922 , n35923 , n35924 , n35925 , n35926 , n35927 , n35928 , n35929 , n35930 , n35931 , n35932 , n35933 , n35934 , n35935 , n35936 , n35937 , n35938 , n35939 , n35940 , n35941 , n35942 , n35943 , n35944 , n35945 , n35946 , n35947 , n35948 , n35949 , n35950 , n35951 , n35952 , n35953 , n35954 , n35955 , n35956 , n35957 , n35958 , n35959 , n35960 , n35961 , n35962 , n35963 , n35964 , n35965 , n35966 , n35967 , n35968 , n35969 , n35970 , n35971 , n35972 , n35973 , n35974 , n35975 , n35976 , n35977 , n35978 , n35979 , n35980 , n35981 , n35982 , n35983 , n35984 , n35985 , n35986 , n35987 , n35988 , n35989 , n35990 , n35991 , n35992 , n35993 , n35994 , n35995 , n35996 , n35997 , n35998 , n35999 , n36000 , n36001 , n36002 , n36003 , n36004 , n36005 , n36006 , n36007 , n36008 , n36009 , n36010 , n36011 , n36012 , n36013 , n36014 , n36015 , n36016 , n36017 , n36018 , n36019 , n36020 , n36021 , n36022 , n36023 , n36024 , n36025 , n36026 , n36027 , n36028 , n36029 , n36030 , n36031 , n36032 , n36033 , n36034 , n36035 , n36036 , n36037 , n36038 , n36039 , n36040 , n36041 , n36042 , n36043 , n36044 , n36045 , n36046 , n36047 , n36048 , n36049 , n36050 , n36051 , n36052 , n36053 , n36054 , n36055 , n36056 , n36057 , n36058 , n36059 , n36060 , n36061 , n36062 , n36063 , n36064 , n36065 , n36066 , n36067 , n36068 , n36069 , n36070 , n36071 , n36072 , n36073 , n36074 , n36075 , n36076 , n36077 , n36078 , n36079 , n36080 , n36081 , n36082 , n36083 , n36084 , n36085 , n36086 , n36087 , n36088 , n36089 , n36090 , n36091 , n36092 , n36093 , n36094 , n36095 , n36096 , n36097 , n36098 , n36099 , n36100 , n36101 , n36102 , n36103 , n36104 , n36105 , n36106 , n36107 , n36108 , n36109 , n36110 , n36111 , n36112 , n36113 , n36114 , n36115 , n36116 , n36117 , n36118 , n36119 , n36120 , n36121 , n36122 , n36123 , n36124 , n36125 , n36126 , n36127 , n36128 , n36129 , n36130 , n36131 , n36132 , n36133 , n36134 , n36135 , n36136 , n36137 , n36138 , n36139 , n36140 , n36141 , n36142 , n36143 , n36144 , n36145 , n36146 , n36147 , n36148 , n36149 , n36150 , n36151 , n36152 , n36153 , n36154 , n36155 , n36156 , n36157 , n36158 , n36159 , n36160 , n36161 , n36162 , n36163 , n36164 , n36165 , n36166 , n36167 , n36168 , n36169 , n36170 , n36171 , n36172 , n36173 , n36174 , n36175 , n36176 , n36177 , n36178 , n36179 , n36180 , n36181 , n36182 , n36183 , n36184 , n36185 , n36186 , n36187 , n36188 , n36189 , n36190 , n36191 , n36192 , n36193 , n36194 , n36195 , n36196 , n36197 , n36198 , n36199 , n36200 , n36201 , n36202 , n36203 , n36204 , n36205 , n36206 , n36207 , n36208 , n36209 , n36210 , n36211 , n36212 , n36213 , n36214 , n36215 , n36216 , n36217 , n36218 , n36219 , n36220 , n36221 , n36222 , n36223 , n36224 , n36225 , n36226 , n36227 , n36228 , n36229 , n36230 , n36231 , n36232 , n36233 , n36234 , n36235 , n36236 , n36237 , n36238 , n36239 , n36240 , n36241 , n36242 , n36243 , n36244 , n36245 , n36246 , n36247 , n36248 , n36249 , n36250 , n36251 , n36252 , n36253 , n36254 , n36255 , n36256 , n36257 , n36258 , n36259 , n36260 , n36261 , n36262 , n36263 , n36264 , n36265 , n36266 , n36267 , n36268 , n36269 , n36270 , n36271 , n36272 , n36273 , n36274 , n36275 , n36276 , n36277 , n36278 , n36279 , n36280 , n36281 , n36282 , n36283 , n36284 , n36285 , n36286 , n36287 , n36288 , n36289 , n36290 , n36291 , n36292 , n36293 , n36294 , n36295 , n36296 , n36297 , n36298 , n36299 , n36300 , n36301 , n36302 , n36303 , n36304 , n36305 , n36306 , n36307 , n36308 , n36309 , n36310 , n36311 , n36312 , n36313 , n36314 , n36315 , n36316 , n36317 , n36318 , n36319 , n36320 , n36321 , n36322 , n36323 , n36324 , n36325 , n36326 , n36327 , n36328 , n36329 , n36330 , n36331 , n36332 , n36333 , n36334 , n36335 , n36336 , n36337 , n36338 , n36339 , n36340 , n36341 , n36342 , n36343 , n36344 , n36345 , n36346 , n36347 , n36348 , n36349 , n36350 , n36351 , n36352 , n36353 , n36354 , n36355 , n36356 , n36357 , n36358 , n36359 , n36360 , n36361 , n36362 , n36363 , n36364 , n36365 , n36366 , n36367 , n36368 , n36369 , n36370 , n36371 , n36372 , n36373 , n36374 , n36375 , n36376 , n36377 , n36378 , n36379 , n36380 , n36381 , n36382 , n36383 , n36384 , n36385 , n36386 , n36387 , n36388 , n36389 , n36390 , n36391 , n36392 , n36393 , n36394 , n36395 , n36396 , n36397 , n36398 , n36399 , n36400 , n36401 , n36402 , n36403 , n36404 , n36405 , n36406 , n36407 , n36408 , n36409 , n36410 , n36411 , n36412 , n36413 , n36414 , n36415 , n36416 , n36417 , n36418 , n36419 , n36420 , n36421 , n36422 , n36423 , n36424 , n36425 , n36426 , n36427 , n36428 , n36429 , n36430 , n36431 , n36432 , n36433 , n36434 , n36435 , n36436 , n36437 , n36438 , n36439 , n36440 , n36441 , n36442 , n36443 , n36444 , n36445 , n36446 , n36447 , n36448 , n36449 , n36450 , n36451 , n36452 , n36453 , n36454 , n36455 , n36456 , n36457 , n36458 , n36459 , n36460 , n36461 , n36462 , n36463 , n36464 , n36465 , n36466 , n36467 , n36468 , n36469 , n36470 , n36471 , n36472 , n36473 , n36474 , n36475 , n36476 , n36477 , n36478 , n36479 , n36480 , n36481 , n36482 , n36483 , n36484 , n36485 , n36486 , n36487 , n36488 , n36489 , n36490 , n36491 , n36492 , n36493 , n36494 , n36495 , n36496 , n36497 , n36498 , n36499 , n36500 , n36501 , n36502 , n36503 , n36504 , n36505 , n36506 , n36507 , n36508 , n36509 , n36510 , n36511 , n36512 , n36513 , n36514 , n36515 , n36516 , n36517 , n36518 , n36519 , n36520 , n36521 , n36522 , n36523 , n36524 , n36525 , n36526 , n36527 , n36528 , n36529 , n36530 , n36531 , n36532 , n36533 , n36534 , n36535 , n36536 , n36537 , n36538 , n36539 , n36540 , n36541 , n36542 , n36543 , n36544 , n36545 , n36546 , n36547 , n36548 , n36549 , n36550 , n36551 , n36552 , n36553 , n36554 , n36555 , n36556 , n36557 , n36558 , n36559 , n36560 , n36561 , n36562 , n36563 , n36564 , n36565 , n36566 , n36567 , n36568 , n36569 , n36570 , n36571 , n36572 , n36573 , n36574 , n36575 , n36576 , n36577 , n36578 , n36579 , n36580 , n36581 , n36582 , n36583 , n36584 , n36585 , n36586 , n36587 , n36588 , n36589 , n36590 , n36591 , n36592 , n36593 , n36594 , n36595 , n36596 , n36597 , n36598 , n36599 , n36600 , n36601 , n36602 , n36603 , n36604 , n36605 , n36606 , n36607 , n36608 , n36609 , n36610 , n36611 , n36612 , n36613 , n36614 , n36615 , n36616 , n36617 , n36618 , n36619 , n36620 , n36621 , n36622 , n36623 , n36624 , n36625 , n36626 , n36627 , n36628 , n36629 , n36630 , n36631 , n36632 , n36633 , n36634 , n36635 , n36636 , n36637 , n36638 , n36639 , n36640 , n36641 , n36642 , n36643 , n36644 , n36645 , n36646 , n36647 , n36648 , n36649 , n36650 , n36651 , n36652 , n36653 , n36654 , n36655 , n36656 , n36657 , n36658 , n36659 , n36660 , n36661 , n36662 , n36663 , n36664 , n36665 , n36666 , n36667 , n36668 , n36669 , n36670 , n36671 , n36672 , n36673 , n36674 , n36675 , n36676 , n36677 , n36678 , n36679 , n36680 , n36681 , n36682 , n36683 , n36684 , n36685 , n36686 , n36687 , n36688 , n36689 , n36690 , n36691 , n36692 , n36693 , n36694 , n36695 , n36696 , n36697 , n36698 , n36699 , n36700 , n36701 , n36702 , n36703 , n36704 , n36705 , n36706 , n36707 , n36708 , n36709 , n36710 , n36711 , n36712 , n36713 , n36714 , n36715 , n36716 , n36717 , n36718 , n36719 , n36720 , n36721 , n36722 , n36723 , n36724 , n36725 , n36726 , n36727 , n36728 , n36729 , n36730 , n36731 , n36732 , n36733 , n36734 , n36735 , n36736 , n36737 , n36738 , n36739 , n36740 , n36741 , n36742 , n36743 , n36744 , n36745 , n36746 , n36747 , n36748 , n36749 , n36750 , n36751 , n36752 , n36753 , n36754 , n36755 , n36756 , n36757 , n36758 , n36759 , n36760 , n36761 , n36762 , n36763 , n36764 , n36765 , n36766 , n36767 , n36768 , n36769 , n36770 , n36771 , n36772 , n36773 , n36774 , n36775 , n36776 , n36777 , n36778 , n36779 , n36780 , n36781 , n36782 , n36783 , n36784 , n36785 , n36786 , n36787 , n36788 , n36789 , n36790 , n36791 , n36792 , n36793 , n36794 , n36795 , n36796 , n36797 , n36798 , n36799 , n36800 , n36801 , n36802 , n36803 , n36804 , n36805 , n36806 , n36807 , n36808 , n36809 , n36810 , n36811 , n36812 , n36813 , n36814 , n36815 , n36816 , n36817 , n36818 , n36819 , n36820 , n36821 , n36822 , n36823 , n36824 , n36825 , n36826 , n36827 , n36828 , n36829 , n36830 , n36831 , n36832 , n36833 , n36834 , n36835 , n36836 , n36837 , n36838 , n36839 , n36840 , n36841 , n36842 , n36843 , n36844 , n36845 , n36846 , n36847 , n36848 , n36849 , n36850 , n36851 , n36852 , n36853 , n36854 , n36855 , n36856 , n36857 , n36858 , n36859 , n36860 , n36861 , n36862 , n36863 , n36864 , n36865 , n36866 , n36867 , n36868 , n36869 , n36870 , n36871 , n36872 , n36873 , n36874 , n36875 , n36876 , n36877 , n36878 , n36879 , n36880 , n36881 , n36882 , n36883 , n36884 , n36885 , n36886 , n36887 , n36888 , n36889 , n36890 , n36891 , n36892 , n36893 , n36894 , n36895 , n36896 , n36897 , n36898 , n36899 , n36900 , n36901 , n36902 , n36903 , n36904 , n36905 , n36906 , n36907 , n36908 , n36909 , n36910 , n36911 , n36912 , n36913 , n36914 , n36915 , n36916 , n36917 , n36918 , n36919 , n36920 , n36921 , n36922 , n36923 , n36924 , n36925 , n36926 , n36927 , n36928 , n36929 , n36930 , n36931 , n36932 , n36933 , n36934 , n36935 , n36936 , n36937 , n36938 , n36939 , n36940 , n36941 , n36942 , n36943 , n36944 , n36945 , n36946 , n36947 , n36948 , n36949 , n36950 , n36951 , n36952 , n36953 , n36954 , n36955 , n36956 , n36957 , n36958 , n36959 , n36960 , n36961 , n36962 , n36963 , n36964 , n36965 , n36966 , n36967 , n36968 , n36969 , n36970 , n36971 , n36972 , n36973 , n36974 , n36975 , n36976 , n36977 , n36978 , n36979 , n36980 , n36981 , n36982 , n36983 , n36984 , n36985 , n36986 , n36987 , n36988 , n36989 , n36990 , n36991 , n36992 , n36993 , n36994 , n36995 , n36996 , n36997 , n36998 , n36999 , n37000 , n37001 , n37002 , n37003 , n37004 , n37005 , n37006 , n37007 , n37008 , n37009 , n37010 , n37011 , n37012 , n37013 , n37014 , n37015 , n37016 , n37017 , n37018 , n37019 , n37020 , n37021 , n37022 , n37023 , n37024 , n37025 , n37026 , n37027 , n37028 , n37029 , n37030 , n37031 , n37032 , n37033 , n37034 , n37035 , n37036 , n37037 , n37038 , n37039 , n37040 , n37041 , n37042 , n37043 , n37044 , n37045 , n37046 , n37047 , n37048 , n37049 , n37050 , n37051 , n37052 , n37053 , n37054 , n37055 , n37056 , n37057 , n37058 , n37059 , n37060 , n37061 , n37062 , n37063 , n37064 , n37065 , n37066 , n37067 , n37068 , n37069 , n37070 , n37071 , n37072 , n37073 , n37074 , n37075 , n37076 , n37077 , n37078 , n37079 , n37080 , n37081 , n37082 , n37083 , n37084 , n37085 , n37086 , n37087 , n37088 , n37089 , n37090 , n37091 , n37092 , n37093 , n37094 , n37095 , n37096 , n37097 , n37098 , n37099 , n37100 , n37101 , n37102 , n37103 , n37104 , n37105 , n37106 , n37107 , n37108 , n37109 , n37110 , n37111 , n37112 , n37113 , n37114 , n37115 , n37116 , n37117 , n37118 , n37119 , n37120 , n37121 , n37122 , n37123 , n37124 , n37125 , n37126 , n37127 , n37128 , n37129 , n37130 , n37131 , n37132 , n37133 , n37134 , n37135 , n37136 , n37137 , n37138 , n37139 , n37140 , n37141 , n37142 , n37143 , n37144 , n37145 , n37146 , n37147 , n37148 , n37149 , n37150 , n37151 , n37152 , n37153 , n37154 , n37155 , n37156 , n37157 , n37158 , n37159 , n37160 , n37161 , n37162 , n37163 , n37164 , n37165 , n37166 , n37167 , n37168 , n37169 , n37170 , n37171 , n37172 , n37173 , n37174 , n37175 , n37176 , n37177 , n37178 , n37179 , n37180 , n37181 , n37182 , n37183 , n37184 , n37185 , n37186 , n37187 , n37188 , n37189 , n37190 , n37191 , n37192 , n37193 , n37194 , n37195 , n37196 , n37197 , n37198 , n37199 , n37200 , n37201 , n37202 , n37203 , n37204 , n37205 , n37206 , n37207 , n37208 , n37209 , n37210 , n37211 , n37212 , n37213 , n37214 , n37215 , n37216 , n37217 , n37218 , n37219 , n37220 , n37221 , n37222 , n37223 , n37224 , n37225 , n37226 , n37227 , n37228 , n37229 , n37230 , n37231 , n37232 , n37233 , n37234 , n37235 , n37236 , n37237 , n37238 , n37239 , n37240 , n37241 , n37242 , n37243 , n37244 , n37245 , n37246 , n37247 , n37248 , n37249 , n37250 , n37251 , n37252 , n37253 , n37254 , n37255 , n37256 , n37257 , n37258 , n37259 , n37260 , n37261 , n37262 , n37263 , n37264 , n37265 , n37266 , n37267 , n37268 , n37269 , n37270 , n37271 , n37272 , n37273 , n37274 , n37275 , n37276 , n37277 , n37278 , n37279 , n37280 , n37281 , n37282 , n37283 , n37284 , n37285 , n37286 , n37287 , n37288 , n37289 , n37290 , n37291 , n37292 , n37293 , n37294 , n37295 , n37296 , n37297 , n37298 , n37299 , n37300 , n37301 , n37302 , n37303 , n37304 , n37305 , n37306 , n37307 , n37308 , n37309 , n37310 , n37311 , n37312 , n37313 , n37314 , n37315 , n37316 , n37317 , n37318 , n37319 , n37320 , n37321 , n37322 , n37323 , n37324 , n37325 , n37326 , n37327 , n37328 , n37329 , n37330 , n37331 , n37332 , n37333 , n37334 , n37335 , n37336 , n37337 , n37338 , n37339 , n37340 , n37341 , n37342 , n37343 , n37344 , n37345 , n37346 , n37347 , n37348 , n37349 , n37350 , n37351 , n37352 , n37353 , n37354 , n37355 , n37356 , n37357 , n37358 , n37359 , n37360 , n37361 , n37362 , n37363 , n37364 , n37365 , n37366 , n37367 , n37368 , n37369 , n37370 , n37371 , n37372 , n37373 , n37374 , n37375 , n37376 , n37377 , n37378 , n37379 , n37380 , n37381 , n37382 , n37383 , n37384 , n37385 , n37386 , n37387 , n37388 , n37389 , n37390 , n37391 , n37392 , n37393 , n37394 , n37395 , n37396 , n37397 , n37398 , n37399 , n37400 , n37401 , n37402 , n37403 , n37404 , n37405 , n37406 , n37407 , n37408 , n37409 , n37410 , n37411 , n37412 , n37413 , n37414 , n37415 , n37416 , n37417 , n37418 , n37419 , n37420 , n37421 , n37422 , n37423 , n37424 , n37425 , n37426 , n37427 , n37428 , n37429 , n37430 , n37431 , n37432 , n37433 , n37434 , n37435 , n37436 , n37437 , n37438 , n37439 , n37440 , n37441 , n37442 , n37443 , n37444 , n37445 , n37446 , n37447 , n37448 , n37449 , n37450 , n37451 , n37452 , n37453 , n37454 , n37455 , n37456 , n37457 , n37458 , n37459 , n37460 , n37461 , n37462 , n37463 , n37464 , n37465 , n37466 , n37467 , n37468 , n37469 , n37470 , n37471 , n37472 , n37473 , n37474 , n37475 , n37476 , n37477 , n37478 , n37479 , n37480 , n37481 , n37482 , n37483 , n37484 , n37485 , n37486 , n37487 , n37488 , n37489 , n37490 , n37491 , n37492 , n37493 , n37494 , n37495 , n37496 , n37497 , n37498 , n37499 , n37500 , n37501 , n37502 , n37503 , n37504 , n37505 , n37506 , n37507 , n37508 , n37509 , n37510 , n37511 , n37512 , n37513 , n37514 , n37515 , n37516 , n37517 , n37518 , n37519 , n37520 , n37521 , n37522 , n37523 , n37524 , n37525 , n37526 , n37527 , n37528 , n37529 , n37530 , n37531 , n37532 , n37533 , n37534 , n37535 , n37536 , n37537 , n37538 , n37539 , n37540 , n37541 , n37542 , n37543 , n37544 , n37545 , n37546 , n37547 , n37548 , n37549 , n37550 , n37551 , n37552 , n37553 , n37554 , n37555 , n37556 , n37557 , n37558 , n37559 , n37560 , n37561 , n37562 , n37563 , n37564 , n37565 , n37566 , n37567 , n37568 , n37569 , n37570 , n37571 , n37572 , n37573 , n37574 , n37575 , n37576 , n37577 , n37578 , n37579 , n37580 , n37581 , n37582 , n37583 , n37584 , n37585 , n37586 , n37587 , n37588 , n37589 , n37590 , n37591 , n37592 , n37593 , n37594 , n37595 , n37596 , n37597 , n37598 , n37599 , n37600 , n37601 , n37602 , n37603 , n37604 , n37605 , n37606 , n37607 , n37608 , n37609 , n37610 , n37611 , n37612 , n37613 , n37614 , n37615 , n37616 , n37617 , n37618 , n37619 , n37620 , n37621 , n37622 , n37623 , n37624 , n37625 , n37626 , n37627 , n37628 , n37629 , n37630 , n37631 , n37632 , n37633 , n37634 , n37635 , n37636 , n37637 , n37638 , n37639 , n37640 , n37641 , n37642 , n37643 , n37644 , n37645 , n37646 , n37647 , n37648 , n37649 , n37650 , n37651 , n37652 , n37653 , n37654 , n37655 , n37656 , n37657 , n37658 , n37659 , n37660 , n37661 , n37662 , n37663 , n37664 , n37665 , n37666 , n37667 , n37668 , n37669 , n37670 , n37671 , n37672 , n37673 , n37674 , n37675 , n37676 , n37677 , n37678 , n37679 , n37680 , n37681 , n37682 , n37683 , n37684 , n37685 , n37686 , n37687 , n37688 , n37689 , n37690 , n37691 , n37692 , n37693 , n37694 , n37695 , n37696 , n37697 , n37698 , n37699 , n37700 , n37701 , n37702 , n37703 , n37704 , n37705 , n37706 , n37707 , n37708 , n37709 , n37710 , n37711 , n37712 , n37713 , n37714 , n37715 , n37716 , n37717 , n37718 , n37719 , n37720 , n37721 , n37722 , n37723 , n37724 , n37725 , n37726 , n37727 , n37728 , n37729 , n37730 , n37731 , n37732 , n37733 , n37734 , n37735 , n37736 , n37737 , n37738 , n37739 , n37740 , n37741 , n37742 , n37743 , n37744 , n37745 , n37746 , n37747 , n37748 , n37749 , n37750 , n37751 , n37752 , n37753 , n37754 , n37755 , n37756 , n37757 , n37758 , n37759 , n37760 , n37761 , n37762 , n37763 , n37764 , n37765 , n37766 , n37767 , n37768 , n37769 , n37770 , n37771 , n37772 , n37773 , n37774 , n37775 , n37776 , n37777 , n37778 , n37779 , n37780 , n37781 , n37782 , n37783 , n37784 , n37785 , n37786 , n37787 , n37788 , n37789 , n37790 , n37791 , n37792 , n37793 , n37794 , n37795 , n37796 , n37797 , n37798 , n37799 , n37800 , n37801 , n37802 , n37803 , n37804 , n37805 , n37806 , n37807 , n37808 , n37809 , n37810 , n37811 , n37812 , n37813 , n37814 , n37815 , n37816 , n37817 , n37818 , n37819 , n37820 , n37821 , n37822 , n37823 , n37824 , n37825 , n37826 , n37827 , n37828 , n37829 , n37830 , n37831 , n37832 , n37833 , n37834 , n37835 , n37836 , n37837 , n37838 , n37839 , n37840 , n37841 , n37842 , n37843 , n37844 , n37845 , n37846 , n37847 , n37848 , n37849 , n37850 , n37851 , n37852 , n37853 , n37854 , n37855 , n37856 , n37857 , n37858 , n37859 , n37860 , n37861 , n37862 , n37863 , n37864 , n37865 , n37866 , n37867 , n37868 , n37869 , n37870 , n37871 , n37872 , n37873 , n37874 , n37875 , n37876 , n37877 , n37878 , n37879 , n37880 , n37881 , n37882 , n37883 , n37884 , n37885 , n37886 , n37887 , n37888 , n37889 , n37890 , n37891 , n37892 , n37893 , n37894 , n37895 , n37896 , n37897 , n37898 , n37899 , n37900 , n37901 , n37902 , n37903 , n37904 , n37905 , n37906 , n37907 , n37908 , n37909 , n37910 , n37911 , n37912 , n37913 , n37914 , n37915 , n37916 , n37917 , n37918 , n37919 , n37920 , n37921 , n37922 , n37923 , n37924 , n37925 , n37926 , n37927 , n37928 , n37929 , n37930 , n37931 , n37932 , n37933 , n37934 , n37935 , n37936 , n37937 , n37938 , n37939 , n37940 , n37941 , n37942 , n37943 , n37944 , n37945 , n37946 , n37947 , n37948 , n37949 , n37950 , n37951 , n37952 , n37953 , n37954 , n37955 , n37956 , n37957 , n37958 , n37959 , n37960 , n37961 , n37962 , n37963 , n37964 , n37965 , n37966 , n37967 , n37968 , n37969 , n37970 , n37971 , n37972 , n37973 , n37974 , n37975 , n37976 , n37977 , n37978 , n37979 , n37980 , n37981 , n37982 , n37983 , n37984 , n37985 , n37986 , n37987 , n37988 , n37989 , n37990 , n37991 , n37992 , n37993 , n37994 , n37995 , n37996 , n37997 , n37998 , n37999 , n38000 , n38001 , n38002 , n38003 , n38004 , n38005 , n38006 , n38007 , n38008 , n38009 , n38010 , n38011 , n38012 , n38013 , n38014 , n38015 , n38016 , n38017 , n38018 , n38019 , n38020 , n38021 , n38022 , n38023 , n38024 , n38025 , n38026 , n38027 , n38028 , n38029 , n38030 , n38031 , n38032 , n38033 , n38034 , n38035 , n38036 , n38037 , n38038 , n38039 , n38040 , n38041 , n38042 , n38043 , n38044 , n38045 , n38046 , n38047 , n38048 , n38049 , n38050 , n38051 , n38052 , n38053 , n38054 , n38055 , n38056 , n38057 , n38058 , n38059 , n38060 , n38061 , n38062 , n38063 , n38064 , n38065 , n38066 , n38067 , n38068 , n38069 , n38070 , n38071 , n38072 , n38073 , n38074 , n38075 , n38076 , n38077 , n38078 , n38079 , n38080 , n38081 , n38082 , n38083 , n38084 , n38085 , n38086 , n38087 , n38088 , n38089 , n38090 , n38091 , n38092 , n38093 , n38094 , n38095 , n38096 , n38097 , n38098 , n38099 , n38100 , n38101 , n38102 , n38103 , n38104 , n38105 , n38106 , n38107 , n38108 , n38109 , n38110 , n38111 , n38112 , n38113 , n38114 , n38115 , n38116 , n38117 , n38118 , n38119 , n38120 , n38121 , n38122 , n38123 , n38124 , n38125 , n38126 , n38127 , n38128 , n38129 , n38130 , n38131 , n38132 , n38133 , n38134 , n38135 , n38136 , n38137 , n38138 , n38139 , n38140 , n38141 , n38142 , n38143 , n38144 , n38145 , n38146 , n38147 , n38148 , n38149 , n38150 , n38151 , n38152 , n38153 , n38154 , n38155 , n38156 , n38157 , n38158 , n38159 , n38160 , n38161 , n38162 , n38163 , n38164 , n38165 , n38166 , n38167 , n38168 , n38169 , n38170 , n38171 , n38172 , n38173 , n38174 , n38175 , n38176 , n38177 , n38178 , n38179 , n38180 , n38181 , n38182 , n38183 , n38184 , n38185 , n38186 , n38187 , n38188 , n38189 , n38190 , n38191 , n38192 , n38193 , n38194 , n38195 , n38196 , n38197 , n38198 , n38199 , n38200 , n38201 , n38202 , n38203 , n38204 , n38205 , n38206 , n38207 , n38208 , n38209 , n38210 , n38211 , n38212 , n38213 , n38214 , n38215 , n38216 , n38217 , n38218 , n38219 , n38220 , n38221 , n38222 , n38223 , n38224 , n38225 , n38226 , n38227 , n38228 , n38229 , n38230 , n38231 , n38232 , n38233 , n38234 , n38235 , n38236 , n38237 , n38238 , n38239 , n38240 , n38241 , n38242 , n38243 , n38244 , n38245 , n38246 , n38247 , n38248 , n38249 , n38250 , n38251 , n38252 , n38253 , n38254 , n38255 , n38256 , n38257 , n38258 , n38259 , n38260 , n38261 , n38262 , n38263 , n38264 , n38265 , n38266 , n38267 , n38268 , n38269 , n38270 , n38271 , n38272 , n38273 , n38274 , n38275 , n38276 , n38277 , n38278 , n38279 , n38280 , n38281 , n38282 , n38283 , n38284 , n38285 , n38286 , n38287 , n38288 , n38289 , n38290 , n38291 , n38292 , n38293 , n38294 , n38295 , n38296 , n38297 , n38298 , n38299 , n38300 , n38301 , n38302 , n38303 , n38304 , n38305 , n38306 , n38307 , n38308 , n38309 , n38310 , n38311 , n38312 , n38313 , n38314 , n38315 , n38316 , n38317 , n38318 , n38319 , n38320 , n38321 , n38322 , n38323 , n38324 , n38325 , n38326 , n38327 , n38328 , n38329 , n38330 , n38331 , n38332 , n38333 , n38334 , n38335 , n38336 , n38337 , n38338 , n38339 , n38340 , n38341 , n38342 , n38343 , n38344 , n38345 , n38346 , n38347 , n38348 , n38349 , n38350 , n38351 , n38352 , n38353 , n38354 , n38355 , n38356 , n38357 , n38358 , n38359 , n38360 , n38361 , n38362 , n38363 , n38364 , n38365 , n38366 , n38367 , n38368 , n38369 , n38370 , n38371 , n38372 , n38373 , n38374 , n38375 , n38376 , n38377 , n38378 , n38379 , n38380 , n38381 , n38382 , n38383 , n38384 , n38385 , n38386 , n38387 , n38388 , n38389 , n38390 , n38391 , n38392 , n38393 , n38394 , n38395 , n38396 , n38397 , n38398 , n38399 , n38400 , n38401 , n38402 , n38403 , n38404 , n38405 , n38406 , n38407 , n38408 , n38409 , n38410 , n38411 , n38412 , n38413 , n38414 , n38415 , n38416 , n38417 , n38418 , n38419 , n38420 , n38421 , n38422 , n38423 , n38424 , n38425 , n38426 , n38427 , n38428 , n38429 , n38430 , n38431 , n38432 , n38433 , n38434 , n38435 , n38436 , n38437 , n38438 , n38439 , n38440 , n38441 , n38442 , n38443 , n38444 , n38445 , n38446 , n38447 , n38448 , n38449 , n38450 , n38451 , n38452 , n38453 , n38454 , n38455 , n38456 , n38457 , n38458 , n38459 , n38460 , n38461 , n38462 , n38463 , n38464 , n38465 , n38466 , n38467 , n38468 , n38469 , n38470 , n38471 , n38472 , n38473 , n38474 , n38475 , n38476 , n38477 , n38478 , n38479 , n38480 , n38481 , n38482 , n38483 , n38484 , n38485 , n38486 , n38487 , n38488 , n38489 , n38490 , n38491 , n38492 , n38493 , n38494 , n38495 , n38496 , n38497 , n38498 , n38499 , n38500 , n38501 , n38502 , n38503 , n38504 , n38505 , n38506 , n38507 , n38508 , n38509 , n38510 , n38511 , n38512 , n38513 , n38514 , n38515 , n38516 , n38517 , n38518 , n38519 , n38520 , n38521 , n38522 , n38523 , n38524 , n38525 , n38526 , n38527 , n38528 , n38529 , n38530 , n38531 , n38532 , n38533 , n38534 , n38535 , n38536 , n38537 , n38538 , n38539 , n38540 , n38541 , n38542 , n38543 , n38544 , n38545 , n38546 , n38547 , n38548 , n38549 , n38550 , n38551 , n38552 , n38553 , n38554 , n38555 , n38556 , n38557 , n38558 , n38559 , n38560 , n38561 , n38562 , n38563 , n38564 , n38565 , n38566 , n38567 , n38568 , n38569 , n38570 , n38571 , n38572 , n38573 , n38574 , n38575 , n38576 , n38577 , n38578 , n38579 , n38580 , n38581 , n38582 , n38583 , n38584 , n38585 , n38586 , n38587 , n38588 , n38589 , n38590 , n38591 , n38592 , n38593 , n38594 , n38595 , n38596 , n38597 , n38598 , n38599 , n38600 , n38601 , n38602 , n38603 , n38604 , n38605 , n38606 , n38607 , n38608 , n38609 , n38610 , n38611 , n38612 , n38613 , n38614 , n38615 , n38616 , n38617 , n38618 , n38619 , n38620 , n38621 , n38622 , n38623 , n38624 , n38625 , n38626 , n38627 , n38628 , n38629 , n38630 , n38631 , n38632 , n38633 , n38634 , n38635 , n38636 , n38637 , n38638 , n38639 , n38640 , n38641 , n38642 , n38643 , n38644 , n38645 , n38646 , n38647 , n38648 , n38649 , n38650 , n38651 , n38652 , n38653 , n38654 , n38655 , n38656 , n38657 , n38658 , n38659 , n38660 , n38661 , n38662 , n38663 , n38664 , n38665 , n38666 , n38667 , n38668 , n38669 , n38670 , n38671 , n38672 , n38673 , n38674 , n38675 , n38676 , n38677 , n38678 , n38679 , n38680 , n38681 , n38682 , n38683 , n38684 , n38685 , n38686 , n38687 , n38688 , n38689 , n38690 , n38691 , n38692 , n38693 , n38694 , n38695 , n38696 , n38697 , n38698 , n38699 , n38700 , n38701 , n38702 , n38703 , n38704 , n38705 , n38706 , n38707 , n38708 , n38709 , n38710 , n38711 , n38712 , n38713 , n38714 , n38715 , n38716 , n38717 , n38718 , n38719 , n38720 , n38721 , n38722 , n38723 , n38724 , n38725 , n38726 , n38727 , n38728 , n38729 , n38730 , n38731 , n38732 , n38733 , n38734 , n38735 , n38736 , n38737 , n38738 , n38739 , n38740 , n38741 , n38742 , n38743 , n38744 , n38745 , n38746 , n38747 , n38748 , n38749 , n38750 , n38751 , n38752 , n38753 , n38754 , n38755 , n38756 , n38757 , n38758 , n38759 , n38760 , n38761 , n38762 , n38763 , n38764 , n38765 , n38766 , n38767 , n38768 , n38769 , n38770 , n38771 , n38772 , n38773 , n38774 , n38775 , n38776 , n38777 , n38778 , n38779 , n38780 , n38781 , n38782 , n38783 , n38784 , n38785 , n38786 , n38787 , n38788 , n38789 , n38790 , n38791 , n38792 , n38793 , n38794 , n38795 , n38796 , n38797 , n38798 , n38799 , n38800 , n38801 , n38802 , n38803 , n38804 , n38805 , n38806 , n38807 , n38808 , n38809 , n38810 , n38811 , n38812 , n38813 , n38814 , n38815 , n38816 , n38817 , n38818 , n38819 , n38820 , n38821 , n38822 , n38823 , n38824 , n38825 , n38826 , n38827 , n38828 , n38829 , n38830 , n38831 , n38832 , n38833 , n38834 , n38835 , n38836 , n38837 , n38838 , n38839 , n38840 , n38841 , n38842 , n38843 , n38844 , n38845 , n38846 , n38847 , n38848 , n38849 , n38850 , n38851 , n38852 , n38853 , n38854 , n38855 , n38856 , n38857 , n38858 , n38859 , n38860 , n38861 , n38862 , n38863 , n38864 , n38865 , n38866 , n38867 , n38868 , n38869 , n38870 , n38871 , n38872 , n38873 , n38874 , n38875 , n38876 , n38877 , n38878 , n38879 , n38880 , n38881 , n38882 , n38883 , n38884 , n38885 , n38886 , n38887 , n38888 , n38889 , n38890 , n38891 , n38892 , n38893 , n38894 , n38895 , n38896 , n38897 , n38898 , n38899 , n38900 , n38901 , n38902 , n38903 , n38904 , n38905 , n38906 , n38907 , n38908 , n38909 , n38910 , n38911 , n38912 , n38913 , n38914 , n38915 , n38916 , n38917 , n38918 , n38919 , n38920 , n38921 , n38922 , n38923 , n38924 , n38925 , n38926 , n38927 , n38928 , n38929 , n38930 , n38931 , n38932 , n38933 , n38934 , n38935 , n38936 , n38937 , n38938 , n38939 , n38940 , n38941 , n38942 , n38943 , n38944 , n38945 , n38946 , n38947 , n38948 , n38949 , n38950 , n38951 , n38952 , n38953 , n38954 , n38955 , n38956 , n38957 , n38958 , n38959 , n38960 , n38961 , n38962 , n38963 , n38964 , n38965 , n38966 , n38967 , n38968 , n38969 , n38970 , n38971 , n38972 , n38973 , n38974 , n38975 , n38976 , n38977 , n38978 , n38979 , n38980 , n38981 , n38982 , n38983 , n38984 , n38985 , n38986 , n38987 , n38988 , n38989 , n38990 , n38991 , n38992 , n38993 , n38994 , n38995 , n38996 , n38997 , n38998 , n38999 , n39000 , n39001 , n39002 , n39003 , n39004 , n39005 , n39006 , n39007 , n39008 , n39009 , n39010 , n39011 , n39012 , n39013 , n39014 , n39015 , n39016 , n39017 , n39018 , n39019 , n39020 , n39021 , n39022 , n39023 , n39024 , n39025 , n39026 , n39027 , n39028 , n39029 , n39030 , n39031 , n39032 , n39033 , n39034 , n39035 , n39036 , n39037 , n39038 , n39039 , n39040 , n39041 , n39042 , n39043 , n39044 , n39045 , n39046 , n39047 , n39048 , n39049 , n39050 , n39051 , n39052 , n39053 , n39054 , n39055 , n39056 , n39057 , n39058 , n39059 , n39060 , n39061 , n39062 , n39063 , n39064 , n39065 , n39066 , n39067 , n39068 , n39069 , n39070 , n39071 , n39072 , n39073 , n39074 , n39075 , n39076 , n39077 , n39078 , n39079 , n39080 , n39081 , n39082 , n39083 , n39084 , n39085 , n39086 , n39087 , n39088 , n39089 , n39090 , n39091 , n39092 , n39093 , n39094 , n39095 , n39096 , n39097 , n39098 , n39099 , n39100 , n39101 , n39102 , n39103 , n39104 , n39105 , n39106 , n39107 , n39108 , n39109 , n39110 , n39111 , n39112 , n39113 , n39114 , n39115 , n39116 , n39117 , n39118 , n39119 , n39120 , n39121 , n39122 , n39123 , n39124 , n39125 , n39126 , n39127 , n39128 , n39129 , n39130 , n39131 , n39132 , n39133 , n39134 , n39135 , n39136 , n39137 , n39138 , n39139 , n39140 , n39141 , n39142 , n39143 , n39144 , n39145 , n39146 , n39147 , n39148 , n39149 , n39150 , n39151 , n39152 , n39153 , n39154 , n39155 , n39156 , n39157 , n39158 , n39159 , n39160 , n39161 , n39162 , n39163 , n39164 , n39165 , n39166 , n39167 , n39168 , n39169 , n39170 , n39171 , n39172 , n39173 , n39174 , n39175 , n39176 , n39177 , n39178 , n39179 , n39180 , n39181 , n39182 , n39183 , n39184 , n39185 , n39186 , n39187 , n39188 , n39189 , n39190 , n39191 , n39192 , n39193 , n39194 , n39195 , n39196 , n39197 , n39198 , n39199 , n39200 , n39201 , n39202 , n39203 , n39204 , n39205 , n39206 , n39207 , n39208 , n39209 , n39210 , n39211 , n39212 , n39213 , n39214 , n39215 , n39216 , n39217 , n39218 , n39219 , n39220 , n39221 , n39222 , n39223 , n39224 , n39225 , n39226 , n39227 , n39228 , n39229 , n39230 , n39231 , n39232 , n39233 , n39234 , n39235 , n39236 , n39237 , n39238 , n39239 , n39240 , n39241 , n39242 , n39243 , n39244 , n39245 , n39246 , n39247 , n39248 , n39249 , n39250 , n39251 , n39252 , n39253 , n39254 , n39255 , n39256 , n39257 , n39258 , n39259 , n39260 , n39261 , n39262 , n39263 , n39264 , n39265 , n39266 , n39267 , n39268 , n39269 , n39270 , n39271 , n39272 , n39273 , n39274 , n39275 , n39276 , n39277 , n39278 , n39279 , n39280 , n39281 , n39282 , n39283 , n39284 , n39285 , n39286 , n39287 , n39288 , n39289 , n39290 , n39291 , n39292 , n39293 , n39294 , n39295 , n39296 , n39297 , n39298 , n39299 , n39300 , n39301 , n39302 , n39303 , n39304 , n39305 , n39306 , n39307 , n39308 , n39309 , n39310 , n39311 , n39312 , n39313 , n39314 , n39315 , n39316 , n39317 , n39318 , n39319 , n39320 , n39321 , n39322 , n39323 , n39324 , n39325 , n39326 , n39327 , n39328 , n39329 , n39330 , n39331 , n39332 , n39333 , n39334 , n39335 , n39336 , n39337 , n39338 , n39339 , n39340 , n39341 , n39342 , n39343 , n39344 , n39345 , n39346 , n39347 , n39348 , n39349 , n39350 , n39351 , n39352 , n39353 , n39354 , n39355 , n39356 , n39357 , n39358 , n39359 , n39360 , n39361 , n39362 , n39363 , n39364 , n39365 , n39366 , n39367 , n39368 , n39369 , n39370 , n39371 , n39372 , n39373 , n39374 , n39375 , n39376 , n39377 , n39378 , n39379 , n39380 , n39381 , n39382 , n39383 , n39384 , n39385 , n39386 , n39387 , n39388 , n39389 , n39390 , n39391 , n39392 , n39393 , n39394 , n39395 , n39396 , n39397 , n39398 , n39399 , n39400 , n39401 , n39402 , n39403 , n39404 , n39405 , n39406 , n39407 , n39408 , n39409 , n39410 , n39411 , n39412 , n39413 , n39414 , n39415 , n39416 , n39417 , n39418 , n39419 , n39420 , n39421 , n39422 , n39423 , n39424 , n39425 , n39426 , n39427 , n39428 , n39429 , n39430 , n39431 , n39432 , n39433 , n39434 , n39435 , n39436 , n39437 , n39438 , n39439 , n39440 , n39441 , n39442 , n39443 , n39444 , n39445 , n39446 , n39447 , n39448 , n39449 , n39450 , n39451 , n39452 , n39453 , n39454 , n39455 , n39456 , n39457 , n39458 , n39459 , n39460 , n39461 , n39462 , n39463 , n39464 , n39465 , n39466 , n39467 , n39468 , n39469 , n39470 , n39471 , n39472 , n39473 , n39474 , n39475 , n39476 , n39477 , n39478 , n39479 , n39480 , n39481 , n39482 , n39483 , n39484 , n39485 , n39486 , n39487 , n39488 , n39489 , n39490 , n39491 , n39492 , n39493 , n39494 , n39495 , n39496 , n39497 , n39498 , n39499 , n39500 , n39501 , n39502 , n39503 , n39504 , n39505 , n39506 , n39507 , n39508 , n39509 , n39510 , n39511 , n39512 , n39513 , n39514 , n39515 , n39516 , n39517 , n39518 , n39519 , n39520 , n39521 , n39522 , n39523 , n39524 , n39525 , n39526 , n39527 , n39528 , n39529 , n39530 , n39531 , n39532 , n39533 , n39534 , n39535 , n39536 , n39537 , n39538 , n39539 , n39540 , n39541 , n39542 , n39543 , n39544 , n39545 , n39546 , n39547 , n39548 , n39549 , n39550 , n39551 , n39552 , n39553 , n39554 , n39555 , n39556 , n39557 , n39558 , n39559 , n39560 , n39561 , n39562 , n39563 , n39564 , n39565 , n39566 , n39567 , n39568 , n39569 , n39570 , n39571 , n39572 , n39573 , n39574 , n39575 , n39576 , n39577 , n39578 , n39579 , n39580 , n39581 , n39582 , n39583 , n39584 , n39585 , n39586 , n39587 , n39588 , n39589 , n39590 , n39591 , n39592 , n39593 , n39594 , n39595 , n39596 , n39597 , n39598 , n39599 , n39600 , n39601 , n39602 , n39603 , n39604 , n39605 , n39606 , n39607 , n39608 , n39609 , n39610 , n39611 , n39612 , n39613 , n39614 , n39615 , n39616 , n39617 , n39618 , n39619 , n39620 , n39621 , n39622 , n39623 , n39624 , n39625 , n39626 , n39627 , n39628 , n39629 , n39630 , n39631 , n39632 , n39633 , n39634 , n39635 , n39636 , n39637 , n39638 , n39639 , n39640 , n39641 , n39642 , n39643 , n39644 , n39645 , n39646 , n39647 , n39648 , n39649 , n39650 , n39651 , n39652 , n39653 , n39654 , n39655 , n39656 , n39657 , n39658 , n39659 , n39660 , n39661 , n39662 , n39663 , n39664 , n39665 , n39666 , n39667 , n39668 , n39669 , n39670 , n39671 , n39672 , n39673 , n39674 , n39675 , n39676 , n39677 , n39678 , n39679 , n39680 , n39681 , n39682 , n39683 , n39684 , n39685 , n39686 , n39687 , n39688 , n39689 , n39690 , n39691 , n39692 , n39693 , n39694 , n39695 , n39696 , n39697 , n39698 , n39699 , n39700 , n39701 , n39702 , n39703 , n39704 , n39705 , n39706 , n39707 , n39708 , n39709 , n39710 , n39711 , n39712 , n39713 , n39714 , n39715 , n39716 , n39717 , n39718 , n39719 , n39720 , n39721 , n39722 , n39723 , n39724 , n39725 , n39726 , n39727 , n39728 , n39729 , n39730 , n39731 , n39732 , n39733 , n39734 , n39735 , n39736 , n39737 , n39738 , n39739 , n39740 , n39741 , n39742 , n39743 , n39744 , n39745 , n39746 , n39747 , n39748 , n39749 , n39750 , n39751 , n39752 , n39753 , n39754 , n39755 , n39756 , n39757 , n39758 , n39759 , n39760 , n39761 , n39762 , n39763 , n39764 , n39765 , n39766 , n39767 , n39768 , n39769 , n39770 , n39771 , n39772 , n39773 , n39774 , n39775 , n39776 , n39777 , n39778 , n39779 , n39780 , n39781 , n39782 , n39783 , n39784 , n39785 , n39786 , n39787 , n39788 , n39789 , n39790 , n39791 , n39792 , n39793 , n39794 , n39795 , n39796 , n39797 , n39798 , n39799 , n39800 , n39801 , n39802 , n39803 , n39804 , n39805 , n39806 , n39807 , n39808 , n39809 , n39810 , n39811 , n39812 , n39813 , n39814 , n39815 , n39816 , n39817 , n39818 , n39819 , n39820 , n39821 , n39822 , n39823 , n39824 , n39825 , n39826 , n39827 , n39828 , n39829 , n39830 , n39831 , n39832 , n39833 , n39834 , n39835 , n39836 , n39837 , n39838 , n39839 , n39840 , n39841 , n39842 , n39843 , n39844 , n39845 , n39846 , n39847 , n39848 , n39849 , n39850 , n39851 , n39852 , n39853 , n39854 , n39855 , n39856 , n39857 , n39858 , n39859 , n39860 , n39861 , n39862 , n39863 , n39864 , n39865 , n39866 , n39867 , n39868 , n39869 , n39870 , n39871 , n39872 , n39873 , n39874 , n39875 , n39876 , n39877 , n39878 , n39879 , n39880 , n39881 , n39882 , n39883 , n39884 , n39885 , n39886 , n39887 , n39888 , n39889 , n39890 , n39891 , n39892 , n39893 , n39894 , n39895 , n39896 , n39897 , n39898 , n39899 , n39900 , n39901 , n39902 , n39903 , n39904 , n39905 , n39906 , n39907 , n39908 , n39909 , n39910 , n39911 , n39912 , n39913 , n39914 , n39915 , n39916 , n39917 , n39918 , n39919 , n39920 , n39921 , n39922 , n39923 , n39924 , n39925 , n39926 , n39927 , n39928 , n39929 , n39930 , n39931 , n39932 , n39933 , n39934 , n39935 , n39936 , n39937 , n39938 , n39939 , n39940 , n39941 , n39942 , n39943 , n39944 , n39945 , n39946 , n39947 , n39948 , n39949 , n39950 , n39951 , n39952 , n39953 , n39954 , n39955 , n39956 , n39957 , n39958 , n39959 , n39960 , n39961 , n39962 , n39963 , n39964 , n39965 , n39966 , n39967 , n39968 , n39969 , n39970 , n39971 , n39972 , n39973 , n39974 , n39975 , n39976 , n39977 , n39978 , n39979 , n39980 , n39981 , n39982 , n39983 , n39984 , n39985 , n39986 , n39987 , n39988 , n39989 , n39990 , n39991 , n39992 , n39993 , n39994 , n39995 , n39996 , n39997 , n39998 , n39999 , n40000 , n40001 , n40002 , n40003 , n40004 , n40005 , n40006 , n40007 , n40008 , n40009 , n40010 , n40011 , n40012 , n40013 , n40014 , n40015 , n40016 , n40017 , n40018 , n40019 , n40020 , n40021 , n40022 , n40023 , n40024 , n40025 , n40026 , n40027 , n40028 , n40029 , n40030 , n40031 , n40032 , n40033 , n40034 , n40035 , n40036 , n40037 , n40038 , n40039 , n40040 , n40041 , n40042 , n40043 , n40044 , n40045 , n40046 , n40047 , n40048 , n40049 , n40050 , n40051 , n40052 , n40053 , n40054 , n40055 , n40056 , n40057 , n40058 , n40059 , n40060 , n40061 , n40062 , n40063 , n40064 , n40065 , n40066 , n40067 , n40068 , n40069 , n40070 , n40071 , n40072 , n40073 , n40074 , n40075 , n40076 , n40077 , n40078 , n40079 , n40080 , n40081 , n40082 , n40083 , n40084 , n40085 , n40086 , n40087 , n40088 , n40089 , n40090 , n40091 , n40092 , n40093 , n40094 , n40095 , n40096 , n40097 , n40098 , n40099 , n40100 , n40101 , n40102 , n40103 , n40104 , n40105 , n40106 , n40107 , n40108 , n40109 , n40110 , n40111 , n40112 , n40113 , n40114 , n40115 , n40116 , n40117 , n40118 , n40119 , n40120 , n40121 , n40122 , n40123 , n40124 , n40125 , n40126 , n40127 , n40128 , n40129 , n40130 , n40131 , n40132 , n40133 , n40134 , n40135 , n40136 , n40137 , n40138 , n40139 , n40140 , n40141 , n40142 , n40143 , n40144 , n40145 , n40146 , n40147 , n40148 , n40149 , n40150 , n40151 , n40152 , n40153 , n40154 , n40155 , n40156 , n40157 , n40158 , n40159 , n40160 , n40161 , n40162 , n40163 , n40164 , n40165 , n40166 , n40167 , n40168 , n40169 , n40170 , n40171 , n40172 , n40173 , n40174 , n40175 , n40176 , n40177 , n40178 , n40179 , n40180 , n40181 , n40182 , n40183 , n40184 , n40185 , n40186 , n40187 , n40188 , n40189 , n40190 , n40191 , n40192 , n40193 , n40194 , n40195 , n40196 , n40197 , n40198 , n40199 , n40200 , n40201 , n40202 , n40203 , n40204 , n40205 , n40206 , n40207 , n40208 , n40209 , n40210 , n40211 , n40212 , n40213 , n40214 , n40215 , n40216 , n40217 , n40218 , n40219 , n40220 , n40221 , n40222 , n40223 , n40224 , n40225 , n40226 , n40227 , n40228 , n40229 , n40230 , n40231 , n40232 , n40233 , n40234 , n40235 , n40236 , n40237 , n40238 , n40239 , n40240 , n40241 , n40242 , n40243 , n40244 , n40245 , n40246 , n40247 , n40248 , n40249 , n40250 , n40251 , n40252 , n40253 , n40254 , n40255 , n40256 , n40257 , n40258 , n40259 , n40260 , n40261 , n40262 , n40263 , n40264 , n40265 , n40266 , n40267 , n40268 , n40269 , n40270 , n40271 , n40272 , n40273 , n40274 , n40275 , n40276 , n40277 , n40278 , n40279 , n40280 , n40281 , n40282 , n40283 , n40284 , n40285 , n40286 , n40287 , n40288 , n40289 , n40290 , n40291 , n40292 , n40293 , n40294 , n40295 , n40296 , n40297 , n40298 , n40299 , n40300 , n40301 , n40302 , n40303 , n40304 , n40305 , n40306 , n40307 , n40308 , n40309 , n40310 , n40311 , n40312 , n40313 , n40314 , n40315 , n40316 , n40317 , n40318 , n40319 , n40320 , n40321 , n40322 , n40323 , n40324 , n40325 , n40326 , n40327 , n40328 , n40329 , n40330 , n40331 , n40332 , n40333 , n40334 , n40335 , n40336 , n40337 , n40338 , n40339 , n40340 , n40341 , n40342 , n40343 , n40344 , n40345 , n40346 , n40347 , n40348 , n40349 , n40350 , n40351 , n40352 , n40353 , n40354 , n40355 , n40356 , n40357 , n40358 , n40359 , n40360 , n40361 , n40362 , n40363 , n40364 , n40365 , n40366 , n40367 , n40368 , n40369 , n40370 , n40371 , n40372 , n40373 , n40374 , n40375 , n40376 , n40377 , n40378 , n40379 , n40380 , n40381 , n40382 , n40383 , n40384 , n40385 , n40386 , n40387 , n40388 , n40389 , n40390 , n40391 , n40392 , n40393 , n40394 , n40395 , n40396 , n40397 , n40398 , n40399 , n40400 , n40401 , n40402 , n40403 , n40404 , n40405 , n40406 , n40407 , n40408 , n40409 , n40410 , n40411 , n40412 , n40413 , n40414 , n40415 , n40416 , n40417 , n40418 , n40419 , n40420 , n40421 , n40422 , n40423 , n40424 , n40425 , n40426 , n40427 , n40428 , n40429 , n40430 , n40431 , n40432 , n40433 , n40434 , n40435 , n40436 , n40437 , n40438 , n40439 , n40440 , n40441 , n40442 , n40443 , n40444 , n40445 , n40446 , n40447 , n40448 , n40449 , n40450 , n40451 , n40452 , n40453 , n40454 , n40455 , n40456 , n40457 , n40458 , n40459 , n40460 , n40461 , n40462 , n40463 , n40464 , n40465 , n40466 , n40467 , n40468 , n40469 , n40470 , n40471 , n40472 , n40473 , n40474 , n40475 , n40476 , n40477 , n40478 , n40479 , n40480 , n40481 , n40482 , n40483 , n40484 , n40485 , n40486 , n40487 , n40488 , n40489 , n40490 , n40491 , n40492 , n40493 , n40494 , n40495 , n40496 , n40497 , n40498 , n40499 , n40500 , n40501 , n40502 , n40503 , n40504 , n40505 , n40506 , n40507 , n40508 , n40509 , n40510 , n40511 , n40512 , n40513 , n40514 , n40515 , n40516 , n40517 , n40518 , n40519 , n40520 , n40521 , n40522 , n40523 , n40524 , n40525 , n40526 , n40527 , n40528 , n40529 , n40530 , n40531 , n40532 , n40533 , n40534 , n40535 , n40536 , n40537 , n40538 , n40539 , n40540 , n40541 , n40542 , n40543 , n40544 , n40545 , n40546 , n40547 , n40548 , n40549 , n40550 , n40551 , n40552 , n40553 , n40554 , n40555 , n40556 , n40557 , n40558 , n40559 , n40560 , n40561 , n40562 , n40563 , n40564 , n40565 , n40566 , n40567 , n40568 , n40569 , n40570 , n40571 , n40572 , n40573 , n40574 , n40575 , n40576 , n40577 , n40578 , n40579 , n40580 , n40581 , n40582 , n40583 , n40584 , n40585 , n40586 , n40587 , n40588 , n40589 , n40590 , n40591 , n40592 , n40593 , n40594 , n40595 , n40596 , n40597 , n40598 , n40599 , n40600 , n40601 , n40602 , n40603 , n40604 , n40605 , n40606 , n40607 , n40608 , n40609 , n40610 , n40611 , n40612 , n40613 , n40614 , n40615 , n40616 , n40617 , n40618 , n40619 , n40620 , n40621 , n40622 , n40623 , n40624 , n40625 , n40626 , n40627 , n40628 , n40629 , n40630 , n40631 , n40632 , n40633 , n40634 , n40635 , n40636 , n40637 , n40638 , n40639 , n40640 , n40641 , n40642 , n40643 , n40644 , n40645 , n40646 , n40647 , n40648 , n40649 , n40650 , n40651 , n40652 , n40653 , n40654 , n40655 , n40656 , n40657 , n40658 , n40659 , n40660 , n40661 , n40662 , n40663 , n40664 , n40665 , n40666 , n40667 , n40668 , n40669 , n40670 , n40671 , n40672 , n40673 , n40674 , n40675 , n40676 , n40677 , n40678 , n40679 , n40680 , n40681 , n40682 , n40683 , n40684 , n40685 , n40686 , n40687 , n40688 , n40689 , n40690 , n40691 , n40692 , n40693 , n40694 , n40695 , n40696 , n40697 , n40698 , n40699 , n40700 , n40701 , n40702 , n40703 , n40704 , n40705 , n40706 , n40707 , n40708 , n40709 , n40710 , n40711 , n40712 , n40713 , n40714 , n40715 , n40716 , n40717 , n40718 , n40719 , n40720 , n40721 , n40722 , n40723 , n40724 , n40725 , n40726 , n40727 , n40728 , n40729 , n40730 , n40731 , n40732 , n40733 , n40734 , n40735 , n40736 , n40737 , n40738 , n40739 , n40740 , n40741 , n40742 , n40743 , n40744 , n40745 , n40746 , n40747 , n40748 , n40749 , n40750 , n40751 , n40752 , n40753 , n40754 , n40755 , n40756 , n40757 , n40758 , n40759 , n40760 , n40761 , n40762 , n40763 , n40764 , n40765 , n40766 , n40767 , n40768 , n40769 , n40770 , n40771 , n40772 , n40773 , n40774 , n40775 , n40776 , n40777 , n40778 , n40779 , n40780 , n40781 , n40782 , n40783 , n40784 , n40785 , n40786 , n40787 , n40788 , n40789 , n40790 , n40791 , n40792 , n40793 , n40794 , n40795 , n40796 , n40797 , n40798 , n40799 , n40800 , n40801 , n40802 , n40803 , n40804 , n40805 , n40806 , n40807 , n40808 , n40809 , n40810 , n40811 , n40812 , n40813 , n40814 , n40815 , n40816 , n40817 , n40818 , n40819 , n40820 , n40821 , n40822 , n40823 , n40824 , n40825 , n40826 , n40827 , n40828 , n40829 , n40830 , n40831 , n40832 , n40833 , n40834 , n40835 , n40836 , n40837 , n40838 , n40839 , n40840 , n40841 , n40842 , n40843 , n40844 , n40845 , n40846 , n40847 , n40848 , n40849 , n40850 , n40851 , n40852 , n40853 , n40854 , n40855 , n40856 , n40857 , n40858 , n40859 , n40860 , n40861 , n40862 , n40863 , n40864 , n40865 , n40866 , n40867 , n40868 , n40869 , n40870 , n40871 , n40872 , n40873 , n40874 , n40875 , n40876 , n40877 , n40878 , n40879 , n40880 , n40881 , n40882 , n40883 , n40884 , n40885 , n40886 , n40887 , n40888 , n40889 , n40890 , n40891 , n40892 , n40893 , n40894 , n40895 , n40896 , n40897 , n40898 , n40899 , n40900 , n40901 , n40902 , n40903 , n40904 , n40905 , n40906 , n40907 , n40908 , n40909 , n40910 , n40911 , n40912 , n40913 , n40914 , n40915 , n40916 , n40917 , n40918 , n40919 , n40920 , n40921 , n40922 , n40923 , n40924 , n40925 , n40926 , n40927 , n40928 , n40929 , n40930 , n40931 , n40932 , n40933 , n40934 , n40935 , n40936 , n40937 , n40938 , n40939 , n40940 , n40941 , n40942 , n40943 , n40944 , n40945 , n40946 , n40947 , n40948 , n40949 , n40950 , n40951 , n40952 , n40953 , n40954 , n40955 , n40956 , n40957 , n40958 , n40959 , n40960 , n40961 , n40962 , n40963 , n40964 , n40965 , n40966 , n40967 , n40968 , n40969 , n40970 , n40971 , n40972 , n40973 , n40974 , n40975 , n40976 , n40977 , n40978 , n40979 , n40980 , n40981 , n40982 , n40983 , n40984 , n40985 , n40986 , n40987 , n40988 , n40989 , n40990 , n40991 , n40992 , n40993 , n40994 , n40995 , n40996 , n40997 , n40998 , n40999 , n41000 , n41001 , n41002 , n41003 , n41004 , n41005 , n41006 , n41007 , n41008 , n41009 , n41010 , n41011 , n41012 , n41013 , n41014 , n41015 , n41016 , n41017 , n41018 , n41019 , n41020 , n41021 , n41022 , n41023 , n41024 , n41025 , n41026 , n41027 , n41028 , n41029 , n41030 , n41031 , n41032 , n41033 , n41034 , n41035 , n41036 , n41037 , n41038 , n41039 , n41040 , n41041 , n41042 , n41043 , n41044 , n41045 , n41046 , n41047 , n41048 , n41049 , n41050 , n41051 , n41052 , n41053 , n41054 , n41055 , n41056 , n41057 , n41058 , n41059 , n41060 , n41061 , n41062 , n41063 , n41064 , n41065 , n41066 , n41067 , n41068 , n41069 , n41070 , n41071 , n41072 , n41073 , n41074 , n41075 , n41076 , n41077 , n41078 , n41079 , n41080 , n41081 , n41082 , n41083 , n41084 , n41085 , n41086 , n41087 , n41088 , n41089 , n41090 , n41091 , n41092 , n41093 , n41094 , n41095 , n41096 , n41097 , n41098 , n41099 , n41100 , n41101 , n41102 , n41103 , n41104 , n41105 , n41106 , n41107 , n41108 , n41109 , n41110 , n41111 , n41112 , n41113 , n41114 , n41115 , n41116 , n41117 , n41118 , n41119 , n41120 , n41121 , n41122 , n41123 , n41124 , n41125 , n41126 , n41127 , n41128 , n41129 , n41130 , n41131 , n41132 , n41133 , n41134 , n41135 , n41136 , n41137 , n41138 , n41139 , n41140 , n41141 , n41142 , n41143 , n41144 , n41145 , n41146 , n41147 , n41148 , n41149 , n41150 , n41151 , n41152 , n41153 , n41154 , n41155 , n41156 , n41157 , n41158 , n41159 , n41160 , n41161 , n41162 , n41163 , n41164 , n41165 , n41166 , n41167 , n41168 , n41169 , n41170 , n41171 , n41172 , n41173 , n41174 , n41175 , n41176 , n41177 , n41178 , n41179 , n41180 , n41181 , n41182 , n41183 , n41184 , n41185 , n41186 , n41187 , n41188 , n41189 , n41190 , n41191 , n41192 , n41193 , n41194 , n41195 , n41196 , n41197 , n41198 , n41199 , n41200 , n41201 , n41202 , n41203 , n41204 , n41205 , n41206 , n41207 , n41208 , n41209 , n41210 , n41211 , n41212 , n41213 , n41214 , n41215 , n41216 , n41217 , n41218 , n41219 , n41220 , n41221 , n41222 , n41223 , n41224 , n41225 , n41226 , n41227 , n41228 , n41229 , n41230 , n41231 , n41232 , n41233 , n41234 , n41235 , n41236 , n41237 , n41238 , n41239 , n41240 , n41241 , n41242 , n41243 , n41244 , n41245 , n41246 , n41247 , n41248 , n41249 , n41250 , n41251 , n41252 , n41253 , n41254 , n41255 , n41256 , n41257 , n41258 , n41259 , n41260 , n41261 , n41262 , n41263 , n41264 , n41265 , n41266 , n41267 , n41268 , n41269 , n41270 , n41271 , n41272 , n41273 , n41274 , n41275 , n41276 , n41277 , n41278 , n41279 , n41280 , n41281 , n41282 , n41283 , n41284 , n41285 , n41286 , n41287 , n41288 , n41289 , n41290 , n41291 , n41292 , n41293 , n41294 , n41295 , n41296 , n41297 , n41298 , n41299 , n41300 , n41301 , n41302 , n41303 , n41304 , n41305 , n41306 , n41307 , n41308 , n41309 , n41310 , n41311 , n41312 , n41313 , n41314 , n41315 , n41316 , n41317 , n41318 , n41319 , n41320 , n41321 , n41322 , n41323 , n41324 , n41325 , n41326 , n41327 , n41328 , n41329 , n41330 , n41331 , n41332 , n41333 , n41334 , n41335 , n41336 , n41337 , n41338 , n41339 , n41340 , n41341 , n41342 , n41343 , n41344 , n41345 , n41346 , n41347 , n41348 , n41349 , n41350 , n41351 , n41352 , n41353 , n41354 , n41355 , n41356 , n41357 , n41358 , n41359 , n41360 , n41361 , n41362 , n41363 , n41364 , n41365 , n41366 , n41367 , n41368 , n41369 , n41370 , n41371 , n41372 , n41373 , n41374 , n41375 , n41376 , n41377 , n41378 , n41379 , n41380 , n41381 , n41382 , n41383 , n41384 , n41385 , n41386 , n41387 , n41388 , n41389 , n41390 , n41391 , n41392 , n41393 , n41394 , n41395 , n41396 , n41397 , n41398 , n41399 , n41400 , n41401 , n41402 , n41403 , n41404 , n41405 , n41406 , n41407 , n41408 , n41409 , n41410 , n41411 , n41412 , n41413 , n41414 , n41415 , n41416 , n41417 , n41418 , n41419 , n41420 , n41421 , n41422 , n41423 , n41424 , n41425 , n41426 , n41427 , n41428 , n41429 , n41430 , n41431 , n41432 , n41433 , n41434 , n41435 , n41436 , n41437 , n41438 , n41439 , n41440 , n41441 , n41442 , n41443 , n41444 , n41445 , n41446 , n41447 , n41448 , n41449 , n41450 , n41451 , n41452 , n41453 , n41454 , n41455 , n41456 , n41457 , n41458 , n41459 , n41460 , n41461 , n41462 , n41463 , n41464 , n41465 , n41466 , n41467 , n41468 , n41469 , n41470 , n41471 , n41472 , n41473 , n41474 , n41475 , n41476 , n41477 , n41478 , n41479 , n41480 , n41481 , n41482 , n41483 , n41484 , n41485 , n41486 , n41487 , n41488 , n41489 , n41490 , n41491 , n41492 , n41493 , n41494 , n41495 , n41496 , n41497 , n41498 , n41499 , n41500 , n41501 , n41502 , n41503 , n41504 , n41505 , n41506 , n41507 , n41508 , n41509 , n41510 , n41511 , n41512 , n41513 , n41514 , n41515 , n41516 , n41517 , n41518 , n41519 , n41520 , n41521 , n41522 , n41523 , n41524 , n41525 , n41526 , n41527 , n41528 , n41529 , n41530 , n41531 , n41532 , n41533 , n41534 , n41535 , n41536 , n41537 , n41538 , n41539 , n41540 , n41541 , n41542 , n41543 , n41544 , n41545 , n41546 , n41547 , n41548 , n41549 , n41550 , n41551 , n41552 , n41553 , n41554 , n41555 , n41556 , n41557 , n41558 , n41559 , n41560 , n41561 , n41562 , n41563 , n41564 , n41565 , n41566 , n41567 , n41568 , n41569 , n41570 , n41571 , n41572 , n41573 , n41574 , n41575 , n41576 , n41577 , n41578 , n41579 , n41580 , n41581 , n41582 , n41583 , n41584 , n41585 , n41586 , n41587 , n41588 , n41589 , n41590 , n41591 , n41592 , n41593 , n41594 , n41595 , n41596 , n41597 , n41598 , n41599 , n41600 , n41601 , n41602 , n41603 , n41604 , n41605 , n41606 , n41607 , n41608 , n41609 , n41610 , n41611 , n41612 , n41613 , n41614 , n41615 , n41616 , n41617 , n41618 , n41619 , n41620 , n41621 , n41622 , n41623 , n41624 , n41625 , n41626 , n41627 , n41628 , n41629 , n41630 , n41631 , n41632 , n41633 , n41634 , n41635 , n41636 , n41637 , n41638 , n41639 , n41640 , n41641 , n41642 , n41643 , n41644 , n41645 , n41646 , n41647 , n41648 , n41649 , n41650 , n41651 , n41652 , n41653 , n41654 , n41655 , n41656 , n41657 , n41658 , n41659 , n41660 , n41661 , n41662 , n41663 , n41664 , n41665 , n41666 , n41667 , n41668 , n41669 , n41670 , n41671 , n41672 , n41673 , n41674 , n41675 , n41676 , n41677 , n41678 , n41679 , n41680 , n41681 , n41682 , n41683 , n41684 , n41685 , n41686 , n41687 , n41688 , n41689 , n41690 , n41691 , n41692 , n41693 , n41694 , n41695 , n41696 , n41697 , n41698 , n41699 , n41700 , n41701 , n41702 , n41703 , n41704 , n41705 , n41706 , n41707 , n41708 , n41709 , n41710 , n41711 , n41712 , n41713 , n41714 , n41715 , n41716 , n41717 , n41718 , n41719 , n41720 , n41721 , n41722 , n41723 , n41724 , n41725 , n41726 , n41727 , n41728 , n41729 , n41730 , n41731 , n41732 , n41733 , n41734 , n41735 , n41736 , n41737 , n41738 , n41739 , n41740 , n41741 , n41742 , n41743 , n41744 , n41745 , n41746 , n41747 , n41748 , n41749 , n41750 , n41751 , n41752 , n41753 , n41754 , n41755 , n41756 , n41757 , n41758 , n41759 , n41760 , n41761 , n41762 , n41763 , n41764 , n41765 , n41766 , n41767 , n41768 , n41769 , n41770 , n41771 , n41772 , n41773 , n41774 , n41775 , n41776 , n41777 , n41778 , n41779 , n41780 , n41781 , n41782 , n41783 , n41784 , n41785 , n41786 , n41787 , n41788 , n41789 , n41790 , n41791 , n41792 , n41793 , n41794 , n41795 , n41796 , n41797 , n41798 , n41799 , n41800 , n41801 , n41802 , n41803 , n41804 , n41805 , n41806 , n41807 , n41808 , n41809 , n41810 , n41811 , n41812 , n41813 , n41814 , n41815 , n41816 , n41817 , n41818 , n41819 , n41820 , n41821 , n41822 , n41823 , n41824 , n41825 , n41826 , n41827 , n41828 , n41829 , n41830 , n41831 , n41832 , n41833 , n41834 , n41835 , n41836 , n41837 , n41838 , n41839 , n41840 , n41841 , n41842 , n41843 , n41844 , n41845 , n41846 , n41847 , n41848 , n41849 , n41850 , n41851 , n41852 , n41853 , n41854 , n41855 , n41856 , n41857 , n41858 , n41859 , n41860 , n41861 , n41862 , n41863 , n41864 , n41865 , n41866 , n41867 , n41868 , n41869 , n41870 , n41871 , n41872 , n41873 , n41874 , n41875 , n41876 , n41877 , n41878 , n41879 , n41880 , n41881 , n41882 , n41883 , n41884 , n41885 , n41886 , n41887 , n41888 , n41889 , n41890 , n41891 , n41892 , n41893 , n41894 , n41895 , n41896 , n41897 , n41898 , n41899 , n41900 , n41901 , n41902 , n41903 , n41904 , n41905 , n41906 , n41907 , n41908 , n41909 , n41910 , n41911 , n41912 , n41913 , n41914 , n41915 , n41916 , n41917 , n41918 , n41919 , n41920 , n41921 , n41922 , n41923 , n41924 , n41925 , n41926 , n41927 , n41928 , n41929 , n41930 , n41931 , n41932 , n41933 , n41934 , n41935 , n41936 , n41937 , n41938 , n41939 , n41940 , n41941 , n41942 , n41943 , n41944 , n41945 , n41946 , n41947 , n41948 , n41949 , n41950 , n41951 , n41952 , n41953 , n41954 , n41955 , n41956 , n41957 , n41958 , n41959 , n41960 , n41961 , n41962 , n41963 , n41964 , n41965 , n41966 , n41967 , n41968 , n41969 , n41970 , n41971 , n41972 , n41973 , n41974 , n41975 , n41976 , n41977 , n41978 , n41979 , n41980 , n41981 , n41982 , n41983 , n41984 , n41985 , n41986 , n41987 , n41988 , n41989 , n41990 , n41991 , n41992 , n41993 , n41994 , n41995 , n41996 , n41997 , n41998 , n41999 , n42000 , n42001 , n42002 , n42003 , n42004 , n42005 , n42006 , n42007 , n42008 , n42009 , n42010 , n42011 , n42012 , n42013 , n42014 , n42015 , n42016 , n42017 , n42018 , n42019 , n42020 , n42021 , n42022 , n42023 , n42024 , n42025 , n42026 , n42027 , n42028 , n42029 , n42030 , n42031 , n42032 , n42033 , n42034 , n42035 , n42036 , n42037 , n42038 , n42039 , n42040 , n42041 , n42042 , n42043 , n42044 , n42045 , n42046 , n42047 , n42048 , n42049 , n42050 , n42051 , n42052 , n42053 , n42054 , n42055 , n42056 , n42057 , n42058 , n42059 , n42060 , n42061 , n42062 , n42063 , n42064 , n42065 , n42066 , n42067 , n42068 , n42069 , n42070 , n42071 , n42072 , n42073 , n42074 , n42075 , n42076 , n42077 , n42078 , n42079 , n42080 , n42081 , n42082 , n42083 , n42084 , n42085 , n42086 , n42087 , n42088 , n42089 , n42090 , n42091 , n42092 , n42093 , n42094 , n42095 , n42096 , n42097 , n42098 , n42099 , n42100 , n42101 , n42102 , n42103 , n42104 , n42105 , n42106 , n42107 , n42108 , n42109 , n42110 , n42111 , n42112 , n42113 , n42114 , n42115 , n42116 , n42117 , n42118 , n42119 , n42120 , n42121 , n42122 , n42123 , n42124 , n42125 , n42126 , n42127 , n42128 , n42129 , n42130 , n42131 , n42132 , n42133 , n42134 , n42135 , n42136 , n42137 , n42138 , n42139 , n42140 , n42141 , n42142 , n42143 , n42144 , n42145 , n42146 , n42147 , n42148 , n42149 , n42150 , n42151 , n42152 , n42153 , n42154 , n42155 , n42156 , n42157 , n42158 , n42159 , n42160 , n42161 , n42162 , n42163 , n42164 , n42165 , n42166 , n42167 , n42168 , n42169 , n42170 , n42171 , n42172 , n42173 , n42174 , n42175 , n42176 , n42177 , n42178 , n42179 , n42180 , n42181 , n42182 , n42183 , n42184 , n42185 , n42186 , n42187 , n42188 , n42189 , n42190 , n42191 , n42192 , n42193 , n42194 , n42195 , n42196 , n42197 , n42198 , n42199 , n42200 , n42201 , n42202 , n42203 , n42204 , n42205 , n42206 , n42207 , n42208 , n42209 , n42210 , n42211 , n42212 , n42213 , n42214 , n42215 , n42216 , n42217 , n42218 , n42219 , n42220 , n42221 , n42222 , n42223 , n42224 , n42225 , n42226 , n42227 , n42228 , n42229 , n42230 , n42231 , n42232 , n42233 , n42234 , n42235 , n42236 , n42237 , n42238 , n42239 , n42240 , n42241 , n42242 , n42243 , n42244 , n42245 , n42246 , n42247 , n42248 , n42249 , n42250 , n42251 , n42252 , n42253 , n42254 , n42255 , n42256 , n42257 , n42258 , n42259 , n42260 , n42261 , n42262 , n42263 , n42264 , n42265 , n42266 , n42267 , n42268 , n42269 , n42270 , n42271 , n42272 , n42273 , n42274 , n42275 , n42276 , n42277 , n42278 , n42279 , n42280 , n42281 , n42282 , n42283 , n42284 , n42285 , n42286 , n42287 , n42288 , n42289 , n42290 , n42291 , n42292 , n42293 , n42294 , n42295 , n42296 , n42297 , n42298 , n42299 , n42300 , n42301 , n42302 , n42303 , n42304 , n42305 , n42306 , n42307 , n42308 , n42309 , n42310 , n42311 , n42312 , n42313 , n42314 , n42315 , n42316 , n42317 , n42318 , n42319 , n42320 , n42321 , n42322 , n42323 , n42324 , n42325 , n42326 , n42327 , n42328 , n42329 , n42330 , n42331 , n42332 , n42333 , n42334 , n42335 , n42336 , n42337 , n42338 , n42339 , n42340 , n42341 , n42342 , n42343 , n42344 , n42345 , n42346 , n42347 , n42348 , n42349 , n42350 , n42351 , n42352 , n42353 , n42354 , n42355 , n42356 , n42357 , n42358 , n42359 , n42360 , n42361 , n42362 , n42363 , n42364 , n42365 , n42366 , n42367 , n42368 , n42369 , n42370 , n42371 , n42372 , n42373 , n42374 , n42375 , n42376 , n42377 , n42378 , n42379 , n42380 , n42381 , n42382 , n42383 , n42384 , n42385 , n42386 , n42387 , n42388 , n42389 , n42390 , n42391 , n42392 , n42393 , n42394 , n42395 , n42396 , n42397 , n42398 , n42399 , n42400 , n42401 , n42402 , n42403 , n42404 , n42405 , n42406 , n42407 , n42408 , n42409 , n42410 , n42411 , n42412 , n42413 , n42414 , n42415 , n42416 , n42417 , n42418 , n42419 , n42420 , n42421 , n42422 , n42423 , n42424 , n42425 , n42426 , n42427 , n42428 , n42429 , n42430 , n42431 , n42432 , n42433 , n42434 , n42435 , n42436 , n42437 , n42438 , n42439 , n42440 , n42441 , n42442 , n42443 , n42444 , n42445 , n42446 , n42447 , n42448 , n42449 , n42450 , n42451 , n42452 , n42453 , n42454 , n42455 , n42456 , n42457 , n42458 , n42459 , n42460 , n42461 , n42462 , n42463 , n42464 , n42465 , n42466 , n42467 , n42468 , n42469 , n42470 , n42471 , n42472 , n42473 , n42474 , n42475 , n42476 , n42477 , n42478 , n42479 , n42480 , n42481 , n42482 , n42483 , n42484 , n42485 , n42486 , n42487 , n42488 , n42489 , n42490 , n42491 , n42492 , n42493 , n42494 , n42495 , n42496 , n42497 , n42498 , n42499 , n42500 , n42501 , n42502 , n42503 , n42504 , n42505 , n42506 , n42507 , n42508 , n42509 , n42510 , n42511 , n42512 , n42513 , n42514 , n42515 , n42516 , n42517 , n42518 , n42519 , n42520 , n42521 , n42522 , n42523 , n42524 , n42525 , n42526 , n42527 , n42528 , n42529 , n42530 , n42531 , n42532 , n42533 , n42534 , n42535 , n42536 , n42537 , n42538 , n42539 , n42540 , n42541 , n42542 , n42543 , n42544 , n42545 , n42546 , n42547 , n42548 , n42549 , n42550 , n42551 , n42552 , n42553 , n42554 , n42555 , n42556 , n42557 , n42558 , n42559 , n42560 , n42561 , n42562 , n42563 , n42564 , n42565 , n42566 , n42567 , n42568 , n42569 , n42570 , n42571 , n42572 , n42573 , n42574 , n42575 , n42576 , n42577 , n42578 , n42579 , n42580 , n42581 , n42582 , n42583 , n42584 , n42585 , n42586 , n42587 , n42588 , n42589 , n42590 , n42591 , n42592 , n42593 , n42594 , n42595 , n42596 , n42597 , n42598 , n42599 , n42600 , n42601 , n42602 , n42603 , n42604 , n42605 , n42606 , n42607 , n42608 , n42609 , n42610 , n42611 , n42612 , n42613 , n42614 , n42615 , n42616 , n42617 , n42618 , n42619 , n42620 , n42621 , n42622 , n42623 , n42624 , n42625 , n42626 , n42627 , n42628 , n42629 , n42630 , n42631 , n42632 , n42633 , n42634 , n42635 , n42636 , n42637 , n42638 , n42639 , n42640 , n42641 , n42642 , n42643 , n42644 , n42645 , n42646 , n42647 , n42648 , n42649 , n42650 , n42651 , n42652 , n42653 , n42654 , n42655 , n42656 , n42657 , n42658 , n42659 , n42660 , n42661 , n42662 , n42663 , n42664 , n42665 , n42666 , n42667 , n42668 , n42669 , n42670 , n42671 , n42672 , n42673 , n42674 , n42675 , n42676 , n42677 , n42678 , n42679 , n42680 , n42681 , n42682 , n42683 , n42684 , n42685 , n42686 , n42687 , n42688 , n42689 , n42690 , n42691 , n42692 , n42693 , n42694 , n42695 , n42696 , n42697 , n42698 , n42699 , n42700 , n42701 , n42702 , n42703 , n42704 , n42705 , n42706 , n42707 , n42708 , n42709 , n42710 , n42711 , n42712 , n42713 , n42714 , n42715 , n42716 , n42717 , n42718 , n42719 , n42720 , n42721 , n42722 , n42723 , n42724 , n42725 , n42726 , n42727 , n42728 , n42729 , n42730 , n42731 , n42732 , n42733 , n42734 , n42735 , n42736 , n42737 , n42738 , n42739 , n42740 , n42741 , n42742 , n42743 , n42744 , n42745 , n42746 , n42747 , n42748 , n42749 , n42750 , n42751 , n42752 , n42753 , n42754 , n42755 , n42756 , n42757 , n42758 , n42759 , n42760 , n42761 , n42762 , n42763 , n42764 , n42765 , n42766 , n42767 , n42768 , n42769 , n42770 , n42771 , n42772 , n42773 , n42774 , n42775 , n42776 , n42777 , n42778 , n42779 , n42780 , n42781 , n42782 , n42783 , n42784 , n42785 , n42786 , n42787 , n42788 , n42789 , n42790 , n42791 , n42792 , n42793 , n42794 , n42795 , n42796 , n42797 , n42798 , n42799 , n42800 , n42801 , n42802 , n42803 , n42804 , n42805 , n42806 , n42807 , n42808 , n42809 , n42810 , n42811 , n42812 , n42813 , n42814 , n42815 , n42816 , n42817 , n42818 , n42819 , n42820 , n42821 , n42822 , n42823 , n42824 , n42825 , n42826 , n42827 , n42828 , n42829 , n42830 , n42831 , n42832 , n42833 , n42834 , n42835 , n42836 , n42837 , n42838 , n42839 , n42840 , n42841 , n42842 , n42843 , n42844 , n42845 , n42846 , n42847 , n42848 , n42849 , n42850 , n42851 , n42852 , n42853 , n42854 , n42855 , n42856 , n42857 , n42858 , n42859 , n42860 , n42861 , n42862 , n42863 , n42864 , n42865 , n42866 , n42867 , n42868 , n42869 , n42870 , n42871 , n42872 , n42873 , n42874 , n42875 , n42876 , n42877 , n42878 , n42879 , n42880 , n42881 , n42882 , n42883 , n42884 , n42885 , n42886 , n42887 , n42888 , n42889 , n42890 , n42891 , n42892 , n42893 , n42894 , n42895 , n42896 , n42897 , n42898 , n42899 , n42900 , n42901 , n42902 , n42903 , n42904 , n42905 , n42906 , n42907 , n42908 , n42909 , n42910 , n42911 , n42912 , n42913 , n42914 , n42915 , n42916 , n42917 , n42918 , n42919 , n42920 , n42921 , n42922 , n42923 , n42924 , n42925 , n42926 , n42927 , n42928 , n42929 , n42930 , n42931 , n42932 , n42933 , n42934 , n42935 , n42936 , n42937 , n42938 , n42939 , n42940 , n42941 , n42942 , n42943 , n42944 , n42945 , n42946 , n42947 , n42948 , n42949 , n42950 , n42951 , n42952 , n42953 , n42954 , n42955 , n42956 , n42957 , n42958 , n42959 , n42960 , n42961 , n42962 , n42963 , n42964 , n42965 , n42966 , n42967 , n42968 , n42969 , n42970 , n42971 , n42972 , n42973 , n42974 , n42975 , n42976 , n42977 , n42978 , n42979 , n42980 , n42981 , n42982 , n42983 , n42984 , n42985 , n42986 , n42987 , n42988 , n42989 , n42990 , n42991 , n42992 , n42993 , n42994 , n42995 , n42996 , n42997 , n42998 , n42999 , n43000 , n43001 , n43002 , n43003 , n43004 , n43005 , n43006 , n43007 , n43008 , n43009 , n43010 , n43011 , n43012 , n43013 , n43014 , n43015 , n43016 , n43017 , n43018 , n43019 , n43020 , n43021 , n43022 , n43023 , n43024 , n43025 , n43026 , n43027 , n43028 , n43029 , n43030 , n43031 , n43032 , n43033 , n43034 , n43035 , n43036 , n43037 , n43038 , n43039 , n43040 , n43041 , n43042 , n43043 , n43044 , n43045 , n43046 , n43047 , n43048 , n43049 , n43050 , n43051 , n43052 , n43053 , n43054 , n43055 , n43056 , n43057 , n43058 , n43059 , n43060 , n43061 , n43062 , n43063 , n43064 , n43065 , n43066 , n43067 , n43068 , n43069 , n43070 , n43071 , n43072 , n43073 , n43074 , n43075 , n43076 , n43077 , n43078 , n43079 , n43080 , n43081 , n43082 , n43083 , n43084 , n43085 , n43086 , n43087 , n43088 , n43089 , n43090 , n43091 , n43092 , n43093 , n43094 , n43095 , n43096 , n43097 , n43098 , n43099 , n43100 , n43101 , n43102 , n43103 , n43104 , n43105 , n43106 , n43107 , n43108 , n43109 , n43110 , n43111 , n43112 , n43113 , n43114 , n43115 , n43116 , n43117 , n43118 , n43119 , n43120 , n43121 , n43122 , n43123 , n43124 , n43125 , n43126 , n43127 , n43128 , n43129 , n43130 , n43131 , n43132 , n43133 , n43134 , n43135 , n43136 , n43137 , n43138 , n43139 , n43140 , n43141 , n43142 , n43143 , n43144 , n43145 , n43146 , n43147 , n43148 , n43149 , n43150 , n43151 , n43152 , n43153 , n43154 , n43155 , n43156 , n43157 , n43158 , n43159 , n43160 , n43161 , n43162 , n43163 , n43164 , n43165 , n43166 , n43167 , n43168 , n43169 , n43170 , n43171 , n43172 , n43173 , n43174 , n43175 , n43176 , n43177 , n43178 , n43179 , n43180 , n43181 , n43182 , n43183 , n43184 , n43185 , n43186 , n43187 , n43188 , n43189 , n43190 , n43191 , n43192 , n43193 , n43194 , n43195 , n43196 , n43197 , n43198 , n43199 , n43200 , n43201 , n43202 , n43203 , n43204 , n43205 , n43206 , n43207 , n43208 , n43209 , n43210 , n43211 , n43212 , n43213 , n43214 , n43215 , n43216 , n43217 , n43218 , n43219 , n43220 , n43221 , n43222 , n43223 , n43224 , n43225 , n43226 , n43227 , n43228 , n43229 , n43230 , n43231 , n43232 , n43233 , n43234 , n43235 , n43236 , n43237 , n43238 , n43239 , n43240 , n43241 , n43242 , n43243 , n43244 , n43245 , n43246 , n43247 , n43248 , n43249 , n43250 , n43251 , n43252 , n43253 , n43254 , n43255 , n43256 , n43257 , n43258 , n43259 , n43260 , n43261 , n43262 , n43263 , n43264 , n43265 , n43266 , n43267 , n43268 , n43269 , n43270 , n43271 , n43272 , n43273 , n43274 , n43275 , n43276 , n43277 , n43278 , n43279 , n43280 , n43281 , n43282 , n43283 , n43284 , n43285 , n43286 , n43287 , n43288 , n43289 , n43290 , n43291 , n43292 , n43293 , n43294 , n43295 , n43296 , n43297 , n43298 , n43299 , n43300 , n43301 , n43302 , n43303 , n43304 , n43305 , n43306 , n43307 , n43308 , n43309 , n43310 , n43311 , n43312 , n43313 , n43314 , n43315 , n43316 , n43317 , n43318 , n43319 , n43320 , n43321 , n43322 , n43323 , n43324 , n43325 , n43326 , n43327 , n43328 , n43329 , n43330 , n43331 , n43332 , n43333 , n43334 , n43335 , n43336 , n43337 , n43338 , n43339 , n43340 , n43341 , n43342 , n43343 , n43344 , n43345 , n43346 , n43347 , n43348 , n43349 , n43350 , n43351 , n43352 , n43353 , n43354 , n43355 , n43356 , n43357 , n43358 , n43359 , n43360 , n43361 , n43362 , n43363 , n43364 , n43365 , n43366 , n43367 , n43368 , n43369 , n43370 , n43371 , n43372 , n43373 , n43374 , n43375 , n43376 , n43377 , n43378 , n43379 , n43380 , n43381 , n43382 , n43383 , n43384 , n43385 , n43386 , n43387 , n43388 , n43389 , n43390 , n43391 , n43392 , n43393 , n43394 , n43395 , n43396 , n43397 , n43398 , n43399 , n43400 , n43401 , n43402 , n43403 , n43404 , n43405 , n43406 , n43407 , n43408 , n43409 , n43410 , n43411 , n43412 , n43413 , n43414 , n43415 , n43416 , n43417 , n43418 , n43419 , n43420 , n43421 , n43422 , n43423 , n43424 , n43425 , n43426 , n43427 , n43428 , n43429 , n43430 , n43431 , n43432 , n43433 , n43434 , n43435 , n43436 , n43437 , n43438 , n43439 , n43440 , n43441 , n43442 , n43443 , n43444 , n43445 , n43446 , n43447 , n43448 , n43449 , n43450 , n43451 , n43452 , n43453 , n43454 , n43455 , n43456 , n43457 , n43458 , n43459 , n43460 , n43461 , n43462 , n43463 , n43464 , n43465 , n43466 , n43467 , n43468 , n43469 , n43470 , n43471 , n43472 , n43473 , n43474 , n43475 , n43476 , n43477 , n43478 , n43479 , n43480 , n43481 , n43482 , n43483 , n43484 , n43485 , n43486 , n43487 , n43488 , n43489 , n43490 , n43491 , n43492 , n43493 , n43494 , n43495 , n43496 , n43497 , n43498 , n43499 , n43500 , n43501 , n43502 , n43503 , n43504 , n43505 , n43506 , n43507 , n43508 , n43509 , n43510 , n43511 , n43512 , n43513 , n43514 , n43515 , n43516 , n43517 , n43518 , n43519 , n43520 , n43521 , n43522 , n43523 , n43524 , n43525 , n43526 , n43527 , n43528 , n43529 , n43530 , n43531 , n43532 , n43533 , n43534 , n43535 , n43536 , n43537 , n43538 , n43539 , n43540 , n43541 , n43542 , n43543 , n43544 , n43545 , n43546 , n43547 , n43548 , n43549 , n43550 , n43551 , n43552 , n43553 , n43554 , n43555 , n43556 , n43557 , n43558 , n43559 , n43560 , n43561 , n43562 , n43563 , n43564 , n43565 , n43566 , n43567 , n43568 , n43569 , n43570 , n43571 , n43572 , n43573 , n43574 , n43575 , n43576 , n43577 , n43578 , n43579 , n43580 , n43581 , n43582 , n43583 , n43584 , n43585 , n43586 , n43587 , n43588 , n43589 , n43590 , n43591 , n43592 , n43593 , n43594 , n43595 , n43596 , n43597 , n43598 , n43599 , n43600 , n43601 , n43602 , n43603 , n43604 , n43605 , n43606 , n43607 , n43608 , n43609 , n43610 , n43611 , n43612 , n43613 , n43614 , n43615 , n43616 , n43617 , n43618 , n43619 , n43620 , n43621 , n43622 , n43623 , n43624 , n43625 , n43626 , n43627 , n43628 , n43629 , n43630 , n43631 , n43632 , n43633 , n43634 , n43635 , n43636 , n43637 , n43638 , n43639 , n43640 , n43641 , n43642 , n43643 , n43644 , n43645 , n43646 , n43647 , n43648 , n43649 , n43650 , n43651 , n43652 , n43653 , n43654 , n43655 , n43656 , n43657 , n43658 , n43659 , n43660 , n43661 , n43662 , n43663 , n43664 , n43665 , n43666 , n43667 , n43668 , n43669 , n43670 , n43671 , n43672 , n43673 , n43674 , n43675 , n43676 , n43677 , n43678 , n43679 , n43680 , n43681 , n43682 , n43683 , n43684 , n43685 , n43686 , n43687 , n43688 , n43689 , n43690 , n43691 , n43692 , n43693 , n43694 , n43695 , n43696 , n43697 , n43698 , n43699 , n43700 , n43701 , n43702 , n43703 , n43704 , n43705 , n43706 , n43707 , n43708 , n43709 , n43710 , n43711 , n43712 , n43713 , n43714 , n43715 , n43716 , n43717 , n43718 , n43719 , n43720 , n43721 , n43722 , n43723 , n43724 , n43725 , n43726 , n43727 , n43728 , n43729 , n43730 , n43731 , n43732 , n43733 , n43734 , n43735 , n43736 , n43737 , n43738 , n43739 , n43740 , n43741 , n43742 , n43743 , n43744 , n43745 , n43746 , n43747 , n43748 , n43749 , n43750 , n43751 , n43752 , n43753 , n43754 , n43755 , n43756 , n43757 , n43758 , n43759 , n43760 , n43761 , n43762 , n43763 , n43764 , n43765 , n43766 , n43767 , n43768 , n43769 , n43770 , n43771 , n43772 , n43773 , n43774 , n43775 , n43776 , n43777 , n43778 , n43779 , n43780 , n43781 , n43782 , n43783 , n43784 , n43785 , n43786 , n43787 , n43788 , n43789 , n43790 , n43791 , n43792 , n43793 , n43794 , n43795 , n43796 , n43797 , n43798 , n43799 , n43800 , n43801 , n43802 , n43803 , n43804 , n43805 , n43806 , n43807 , n43808 , n43809 , n43810 , n43811 , n43812 , n43813 , n43814 , n43815 , n43816 , n43817 , n43818 , n43819 , n43820 , n43821 , n43822 , n43823 , n43824 , n43825 , n43826 , n43827 , n43828 , n43829 , n43830 , n43831 , n43832 , n43833 , n43834 , n43835 , n43836 , n43837 , n43838 , n43839 , n43840 , n43841 , n43842 , n43843 , n43844 , n43845 , n43846 , n43847 , n43848 , n43849 , n43850 , n43851 , n43852 , n43853 , n43854 , n43855 , n43856 , n43857 , n43858 , n43859 , n43860 , n43861 , n43862 , n43863 , n43864 , n43865 , n43866 , n43867 , n43868 , n43869 , n43870 , n43871 , n43872 , n43873 , n43874 , n43875 , n43876 , n43877 , n43878 , n43879 , n43880 , n43881 , n43882 , n43883 , n43884 , n43885 , n43886 , n43887 , n43888 , n43889 , n43890 , n43891 , n43892 , n43893 , n43894 , n43895 , n43896 , n43897 , n43898 , n43899 , n43900 , n43901 , n43902 , n43903 , n43904 , n43905 , n43906 , n43907 , n43908 , n43909 , n43910 , n43911 , n43912 , n43913 , n43914 , n43915 , n43916 , n43917 , n43918 , n43919 , n43920 , n43921 , n43922 , n43923 , n43924 , n43925 , n43926 , n43927 , n43928 , n43929 , n43930 , n43931 , n43932 , n43933 , n43934 , n43935 , n43936 , n43937 , n43938 , n43939 , n43940 , n43941 , n43942 , n43943 , n43944 , n43945 , n43946 , n43947 , n43948 , n43949 , n43950 , n43951 , n43952 , n43953 , n43954 , n43955 , n43956 , n43957 , n43958 , n43959 , n43960 , n43961 , n43962 , n43963 , n43964 , n43965 , n43966 , n43967 , n43968 , n43969 , n43970 , n43971 , n43972 , n43973 , n43974 , n43975 , n43976 , n43977 , n43978 , n43979 , n43980 , n43981 , n43982 , n43983 , n43984 , n43985 , n43986 , n43987 , n43988 , n43989 , n43990 , n43991 , n43992 , n43993 , n43994 , n43995 , n43996 , n43997 , n43998 , n43999 , n44000 , n44001 , n44002 , n44003 , n44004 , n44005 , n44006 , n44007 , n44008 , n44009 , n44010 , n44011 , n44012 , n44013 , n44014 , n44015 , n44016 , n44017 , n44018 , n44019 , n44020 , n44021 , n44022 , n44023 , n44024 , n44025 , n44026 , n44027 , n44028 , n44029 , n44030 , n44031 , n44032 , n44033 , n44034 , n44035 , n44036 , n44037 , n44038 , n44039 , n44040 , n44041 , n44042 , n44043 , n44044 , n44045 , n44046 , n44047 , n44048 , n44049 , n44050 , n44051 , n44052 , n44053 , n44054 , n44055 , n44056 , n44057 , n44058 , n44059 , n44060 , n44061 , n44062 , n44063 , n44064 , n44065 , n44066 , n44067 , n44068 , n44069 , n44070 , n44071 , n44072 , n44073 , n44074 , n44075 , n44076 , n44077 , n44078 , n44079 , n44080 , n44081 , n44082 , n44083 , n44084 , n44085 , n44086 , n44087 , n44088 , n44089 , n44090 , n44091 , n44092 , n44093 , n44094 , n44095 , n44096 , n44097 , n44098 , n44099 , n44100 , n44101 , n44102 , n44103 , n44104 , n44105 , n44106 , n44107 , n44108 , n44109 , n44110 , n44111 , n44112 , n44113 , n44114 , n44115 , n44116 , n44117 , n44118 , n44119 , n44120 , n44121 , n44122 , n44123 , n44124 , n44125 , n44126 , n44127 , n44128 , n44129 , n44130 , n44131 , n44132 , n44133 , n44134 , n44135 , n44136 , n44137 , n44138 , n44139 , n44140 , n44141 , n44142 , n44143 , n44144 , n44145 , n44146 , n44147 , n44148 , n44149 , n44150 , n44151 , n44152 , n44153 , n44154 , n44155 , n44156 , n44157 , n44158 , n44159 , n44160 , n44161 , n44162 , n44163 , n44164 , n44165 , n44166 , n44167 , n44168 , n44169 , n44170 , n44171 , n44172 , n44173 , n44174 , n44175 , n44176 , n44177 , n44178 , n44179 , n44180 , n44181 , n44182 , n44183 , n44184 , n44185 , n44186 , n44187 , n44188 , n44189 , n44190 , n44191 , n44192 , n44193 , n44194 , n44195 , n44196 , n44197 , n44198 , n44199 , n44200 , n44201 , n44202 , n44203 , n44204 , n44205 , n44206 , n44207 , n44208 , n44209 , n44210 , n44211 , n44212 , n44213 , n44214 , n44215 , n44216 , n44217 , n44218 , n44219 , n44220 , n44221 , n44222 , n44223 , n44224 , n44225 , n44226 , n44227 , n44228 , n44229 , n44230 , n44231 , n44232 , n44233 , n44234 , n44235 , n44236 , n44237 , n44238 , n44239 , n44240 , n44241 , n44242 , n44243 , n44244 , n44245 , n44246 , n44247 , n44248 , n44249 , n44250 , n44251 , n44252 , n44253 , n44254 , n44255 , n44256 , n44257 , n44258 , n44259 , n44260 , n44261 , n44262 , n44263 , n44264 , n44265 , n44266 , n44267 , n44268 , n44269 , n44270 , n44271 , n44272 , n44273 , n44274 , n44275 , n44276 , n44277 , n44278 , n44279 , n44280 , n44281 , n44282 , n44283 , n44284 , n44285 , n44286 , n44287 , n44288 , n44289 , n44290 , n44291 , n44292 , n44293 , n44294 , n44295 , n44296 , n44297 , n44298 , n44299 , n44300 , n44301 , n44302 , n44303 , n44304 , n44305 , n44306 , n44307 , n44308 , n44309 , n44310 , n44311 , n44312 , n44313 , n44314 , n44315 , n44316 , n44317 , n44318 , n44319 , n44320 , n44321 , n44322 , n44323 , n44324 , n44325 , n44326 , n44327 , n44328 , n44329 , n44330 , n44331 , n44332 , n44333 , n44334 , n44335 , n44336 , n44337 , n44338 , n44339 , n44340 , n44341 , n44342 , n44343 , n44344 , n44345 , n44346 , n44347 , n44348 , n44349 , n44350 , n44351 , n44352 , n44353 , n44354 , n44355 , n44356 , n44357 , n44358 , n44359 , n44360 , n44361 , n44362 , n44363 , n44364 , n44365 , n44366 , n44367 , n44368 , n44369 , n44370 , n44371 , n44372 , n44373 , n44374 , n44375 , n44376 , n44377 , n44378 , n44379 , n44380 , n44381 , n44382 , n44383 , n44384 , n44385 , n44386 , n44387 , n44388 , n44389 , n44390 , n44391 , n44392 , n44393 , n44394 , n44395 , n44396 , n44397 , n44398 , n44399 , n44400 , n44401 , n44402 , n44403 , n44404 , n44405 , n44406 , n44407 , n44408 , n44409 , n44410 , n44411 , n44412 , n44413 , n44414 , n44415 , n44416 , n44417 , n44418 , n44419 , n44420 , n44421 , n44422 , n44423 , n44424 , n44425 , n44426 , n44427 , n44428 , n44429 , n44430 , n44431 , n44432 , n44433 , n44434 , n44435 , n44436 , n44437 , n44438 , n44439 , n44440 , n44441 , n44442 , n44443 , n44444 , n44445 , n44446 , n44447 , n44448 , n44449 , n44450 , n44451 , n44452 , n44453 , n44454 , n44455 , n44456 , n44457 , n44458 , n44459 , n44460 , n44461 , n44462 , n44463 , n44464 , n44465 , n44466 , n44467 , n44468 , n44469 , n44470 , n44471 , n44472 , n44473 , n44474 , n44475 , n44476 , n44477 , n44478 , n44479 , n44480 , n44481 , n44482 , n44483 , n44484 , n44485 , n44486 , n44487 , n44488 , n44489 , n44490 , n44491 , n44492 , n44493 , n44494 , n44495 , n44496 , n44497 , n44498 , n44499 , n44500 , n44501 , n44502 , n44503 , n44504 , n44505 , n44506 , n44507 , n44508 , n44509 , n44510 , n44511 , n44512 , n44513 , n44514 , n44515 , n44516 , n44517 , n44518 , n44519 , n44520 , n44521 , n44522 , n44523 , n44524 , n44525 , n44526 , n44527 , n44528 , n44529 , n44530 , n44531 , n44532 , n44533 , n44534 , n44535 , n44536 , n44537 , n44538 , n44539 , n44540 , n44541 , n44542 , n44543 , n44544 , n44545 , n44546 , n44547 , n44548 , n44549 , n44550 , n44551 , n44552 , n44553 , n44554 , n44555 , n44556 , n44557 , n44558 , n44559 , n44560 , n44561 , n44562 , n44563 , n44564 , n44565 , n44566 , n44567 , n44568 , n44569 , n44570 , n44571 , n44572 , n44573 , n44574 , n44575 , n44576 , n44577 , n44578 , n44579 , n44580 , n44581 , n44582 , n44583 , n44584 , n44585 , n44586 , n44587 , n44588 , n44589 , n44590 , n44591 , n44592 , n44593 , n44594 , n44595 , n44596 , n44597 , n44598 , n44599 , n44600 , n44601 , n44602 , n44603 , n44604 , n44605 , n44606 , n44607 , n44608 , n44609 , n44610 , n44611 , n44612 , n44613 , n44614 , n44615 , n44616 , n44617 , n44618 , n44619 , n44620 , n44621 , n44622 , n44623 , n44624 , n44625 , n44626 , n44627 , n44628 , n44629 , n44630 , n44631 , n44632 , n44633 , n44634 , n44635 , n44636 , n44637 , n44638 , n44639 , n44640 , n44641 , n44642 , n44643 , n44644 , n44645 , n44646 , n44647 , n44648 , n44649 , n44650 , n44651 , n44652 , n44653 , n44654 , n44655 , n44656 , n44657 , n44658 , n44659 , n44660 , n44661 , n44662 , n44663 , n44664 , n44665 , n44666 , n44667 , n44668 , n44669 , n44670 , n44671 , n44672 , n44673 , n44674 , n44675 , n44676 , n44677 , n44678 , n44679 , n44680 , n44681 , n44682 , n44683 , n44684 , n44685 , n44686 , n44687 , n44688 , n44689 , n44690 , n44691 , n44692 , n44693 , n44694 , n44695 , n44696 , n44697 , n44698 , n44699 , n44700 , n44701 , n44702 , n44703 , n44704 , n44705 , n44706 , n44707 , n44708 , n44709 , n44710 , n44711 , n44712 , n44713 , n44714 , n44715 , n44716 , n44717 , n44718 , n44719 , n44720 , n44721 , n44722 , n44723 , n44724 , n44725 , n44726 , n44727 , n44728 , n44729 , n44730 , n44731 , n44732 , n44733 , n44734 , n44735 , n44736 , n44737 , n44738 , n44739 , n44740 , n44741 , n44742 , n44743 , n44744 , n44745 , n44746 , n44747 , n44748 , n44749 , n44750 , n44751 , n44752 , n44753 , n44754 , n44755 , n44756 , n44757 , n44758 , n44759 , n44760 , n44761 , n44762 , n44763 , n44764 , n44765 , n44766 , n44767 , n44768 , n44769 , n44770 , n44771 , n44772 , n44773 , n44774 , n44775 , n44776 , n44777 , n44778 , n44779 , n44780 , n44781 , n44782 , n44783 , n44784 , n44785 , n44786 , n44787 , n44788 , n44789 , n44790 , n44791 , n44792 , n44793 , n44794 , n44795 , n44796 , n44797 , n44798 , n44799 , n44800 , n44801 , n44802 , n44803 , n44804 , n44805 , n44806 , n44807 , n44808 , n44809 , n44810 , n44811 , n44812 , n44813 , n44814 , n44815 , n44816 , n44817 , n44818 , n44819 , n44820 , n44821 , n44822 , n44823 , n44824 , n44825 , n44826 , n44827 , n44828 , n44829 , n44830 , n44831 , n44832 , n44833 , n44834 , n44835 , n44836 , n44837 , n44838 , n44839 , n44840 , n44841 , n44842 , n44843 , n44844 , n44845 , n44846 , n44847 , n44848 , n44849 , n44850 , n44851 , n44852 , n44853 , n44854 , n44855 , n44856 , n44857 , n44858 , n44859 , n44860 , n44861 , n44862 , n44863 , n44864 , n44865 , n44866 , n44867 , n44868 , n44869 , n44870 , n44871 , n44872 , n44873 , n44874 , n44875 , n44876 , n44877 , n44878 , n44879 , n44880 , n44881 , n44882 , n44883 , n44884 , n44885 , n44886 , n44887 , n44888 , n44889 , n44890 , n44891 , n44892 , n44893 , n44894 , n44895 , n44896 , n44897 , n44898 , n44899 , n44900 , n44901 , n44902 , n44903 , n44904 , n44905 , n44906 , n44907 , n44908 , n44909 , n44910 , n44911 , n44912 , n44913 , n44914 , n44915 , n44916 , n44917 , n44918 , n44919 , n44920 , n44921 , n44922 , n44923 , n44924 , n44925 , n44926 , n44927 , n44928 , n44929 , n44930 , n44931 , n44932 , n44933 , n44934 , n44935 , n44936 , n44937 , n44938 , n44939 , n44940 , n44941 , n44942 , n44943 , n44944 , n44945 , n44946 , n44947 , n44948 , n44949 , n44950 , n44951 , n44952 , n44953 , n44954 , n44955 , n44956 , n44957 , n44958 , n44959 , n44960 , n44961 , n44962 , n44963 , n44964 , n44965 , n44966 , n44967 , n44968 , n44969 , n44970 , n44971 , n44972 , n44973 , n44974 , n44975 , n44976 , n44977 , n44978 , n44979 , n44980 , n44981 , n44982 , n44983 , n44984 , n44985 , n44986 , n44987 , n44988 , n44989 , n44990 , n44991 , n44992 , n44993 , n44994 , n44995 , n44996 , n44997 , n44998 , n44999 , n45000 , n45001 , n45002 , n45003 , n45004 , n45005 , n45006 , n45007 , n45008 , n45009 , n45010 , n45011 , n45012 , n45013 , n45014 , n45015 , n45016 , n45017 , n45018 , n45019 , n45020 , n45021 , n45022 , n45023 , n45024 , n45025 , n45026 , n45027 , n45028 , n45029 , n45030 , n45031 , n45032 , n45033 , n45034 , n45035 , n45036 , n45037 , n45038 , n45039 , n45040 , n45041 , n45042 , n45043 , n45044 , n45045 , n45046 , n45047 , n45048 , n45049 , n45050 , n45051 , n45052 , n45053 , n45054 , n45055 , n45056 , n45057 , n45058 , n45059 , n45060 , n45061 , n45062 , n45063 , n45064 , n45065 , n45066 , n45067 , n45068 , n45069 , n45070 , n45071 , n45072 , n45073 , n45074 , n45075 , n45076 , n45077 , n45078 , n45079 , n45080 , n45081 , n45082 , n45083 , n45084 , n45085 , n45086 , n45087 , n45088 , n45089 , n45090 , n45091 , n45092 , n45093 , n45094 , n45095 , n45096 , n45097 , n45098 , n45099 , n45100 , n45101 , n45102 , n45103 , n45104 , n45105 , n45106 , n45107 , n45108 , n45109 , n45110 , n45111 , n45112 , n45113 , n45114 , n45115 , n45116 , n45117 , n45118 , n45119 , n45120 , n45121 , n45122 , n45123 , n45124 , n45125 , n45126 , n45127 , n45128 , n45129 , n45130 , n45131 , n45132 , n45133 , n45134 , n45135 , n45136 , n45137 , n45138 , n45139 , n45140 , n45141 , n45142 , n45143 , n45144 , n45145 , n45146 , n45147 , n45148 , n45149 , n45150 , n45151 , n45152 , n45153 , n45154 , n45155 , n45156 , n45157 , n45158 , n45159 , n45160 , n45161 , n45162 , n45163 , n45164 , n45165 , n45166 , n45167 , n45168 , n45169 , n45170 , n45171 , n45172 , n45173 , n45174 , n45175 , n45176 , n45177 , n45178 , n45179 , n45180 , n45181 , n45182 , n45183 , n45184 , n45185 , n45186 , n45187 , n45188 , n45189 , n45190 , n45191 , n45192 , n45193 , n45194 , n45195 , n45196 , n45197 , n45198 , n45199 , n45200 , n45201 , n45202 , n45203 , n45204 , n45205 , n45206 , n45207 , n45208 , n45209 , n45210 , n45211 , n45212 , n45213 , n45214 , n45215 , n45216 , n45217 , n45218 , n45219 , n45220 , n45221 , n45222 , n45223 , n45224 , n45225 , n45226 , n45227 , n45228 , n45229 , n45230 , n45231 , n45232 , n45233 , n45234 , n45235 , n45236 , n45237 , n45238 , n45239 , n45240 , n45241 , n45242 , n45243 , n45244 , n45245 , n45246 , n45247 , n45248 , n45249 , n45250 , n45251 , n45252 , n45253 , n45254 , n45255 , n45256 , n45257 , n45258 , n45259 , n45260 , n45261 , n45262 , n45263 , n45264 , n45265 , n45266 , n45267 , n45268 , n45269 , n45270 , n45271 , n45272 , n45273 ;
  assign n1205 = ~x216 & x833 ;
  assign n1206 = ( x332 & x929 ) | ( x332 & n1205 ) | ( x929 & n1205 ) ;
  assign n1207 = ( x332 & x1144 ) | ( x332 & ~n1205 ) | ( x1144 & ~n1205 ) ;
  assign n1208 = n1206 | n1207 ;
  assign n1209 = x221 & n1208 ;
  assign n1210 = x265 & ~x332 ;
  assign n1211 = x216 & ~n1210 ;
  assign n1212 = x40 | x72 ;
  assign n1213 = x97 | x108 ;
  assign n1214 = x94 | n1213 ;
  assign n1215 = x53 | x60 ;
  assign n1216 = x46 | x86 ;
  assign n1217 = n1215 | n1216 ;
  assign n1218 = n1214 | n1217 ;
  assign n1219 = x61 | x76 ;
  assign n1220 = x85 | x106 ;
  assign n1221 = n1219 | n1220 ;
  assign n1222 = x48 | x89 ;
  assign n1223 = x49 | n1222 ;
  assign n1224 = n1221 | n1223 ;
  assign n1225 = x45 | x104 ;
  assign n1226 = n1224 | n1225 ;
  assign n1227 = x82 | x111 ;
  assign n1228 = x36 | n1227 ;
  assign n1229 = x66 | x73 ;
  assign n1230 = x68 | x84 ;
  assign n1231 = n1229 | n1230 ;
  assign n1232 = n1228 | n1231 ;
  assign n1233 = x83 | x103 ;
  assign n1234 = x67 | x69 ;
  assign n1235 = n1233 | n1234 ;
  assign n1236 = x63 | x107 ;
  assign n1237 = x65 | x71 ;
  assign n1238 = n1236 | n1237 ;
  assign n1239 = n1235 | n1238 ;
  assign n1240 = n1232 | n1239 ;
  assign n1241 = n1226 | n1240 ;
  assign n1242 = x64 | n1241 ;
  assign n1243 = x88 | x98 ;
  assign n1244 = x50 | x77 ;
  assign n1245 = n1243 | n1244 ;
  assign n1246 = x81 | x102 ;
  assign n1247 = n1245 | n1246 ;
  assign n1248 = n1242 | n1247 ;
  assign n1249 = n1218 | n1248 ;
  assign n1250 = x109 | x110 ;
  assign n1251 = x58 | x91 ;
  assign n1252 = x47 | n1251 ;
  assign n1253 = n1250 | n1252 ;
  assign n1254 = n1249 | n1253 ;
  assign n1255 = x90 | x93 ;
  assign n1256 = x70 | x96 ;
  assign n1257 = x35 | x51 ;
  assign n1258 = n1256 | n1257 ;
  assign n1259 = n1255 | n1258 ;
  assign n1260 = n1254 | n1259 ;
  assign n1261 = n1212 | n1260 ;
  assign n1262 = x225 & ~n1261 ;
  assign n1263 = x841 & n1262 ;
  assign n1264 = ( x32 & n1261 ) | ( x32 & n1263 ) | ( n1261 & n1263 ) ;
  assign n1265 = x95 | n1264 ;
  assign n1266 = x47 | x91 ;
  assign n1267 = n1250 | n1266 ;
  assign n1268 = n1218 | n1267 ;
  assign n1269 = x58 | x90 ;
  assign n1270 = n1247 | n1269 ;
  assign n1271 = n1268 | n1270 ;
  assign n1272 = n1242 | n1271 ;
  assign n1273 = x93 | n1272 ;
  assign n1274 = x35 & ~n1273 ;
  assign n1275 = ~x225 & n1274 ;
  assign n1276 = x70 | n1275 ;
  assign n1277 = x51 | x96 ;
  assign n1278 = x35 | x93 ;
  assign n1279 = n1272 | n1278 ;
  assign n1280 = x70 & n1279 ;
  assign n1281 = n1277 | n1280 ;
  assign n1282 = n1212 | n1281 ;
  assign n1283 = n1276 & ~n1282 ;
  assign n1284 = x32 | n1283 ;
  assign n1285 = ~n1265 & n1284 ;
  assign n1286 = x137 & ~n1285 ;
  assign n1287 = ~x833 & x957 ;
  assign n1288 = x1091 & ~n1287 ;
  assign n1289 = x829 & x950 ;
  assign n1290 = x1092 & x1093 ;
  assign n1291 = n1289 & n1290 ;
  assign n1292 = n1288 & n1291 ;
  assign n1293 = x72 | x96 ;
  assign n1294 = x51 | x70 ;
  assign n1295 = n1293 | n1294 ;
  assign n1296 = x40 & ~n1278 ;
  assign n1297 = ~n1295 & n1296 ;
  assign n1298 = ~n1271 & n1297 ;
  assign n1299 = ~n1242 & n1298 ;
  assign n1300 = x32 | n1299 ;
  assign n1301 = x72 & n1260 ;
  assign n1302 = x40 | n1301 ;
  assign n1303 = x51 | n1276 ;
  assign n1304 = x93 & n1272 ;
  assign n1305 = x35 | n1304 ;
  assign n1306 = n1247 | n1268 ;
  assign n1307 = n1242 | n1306 ;
  assign n1308 = x58 & n1307 ;
  assign n1309 = x90 & n1254 ;
  assign n1310 = n1308 | n1309 ;
  assign n1311 = n1218 | n1250 ;
  assign n1312 = x47 | n1311 ;
  assign n1313 = n1248 | n1312 ;
  assign n1314 = x91 & ~n1313 ;
  assign n1315 = n1269 | n1314 ;
  assign n1316 = x109 | n1249 ;
  assign n1317 = x110 & n1316 ;
  assign n1318 = x47 & ~n1246 ;
  assign n1319 = ~n1245 & n1318 ;
  assign n1320 = ~n1311 & n1319 ;
  assign n1321 = ( x91 & n1266 ) | ( x91 & ~n1320 ) | ( n1266 & ~n1320 ) ;
  assign n1322 = x91 | n1266 ;
  assign n1323 = ( n1242 & n1321 ) | ( n1242 & n1322 ) | ( n1321 & n1322 ) ;
  assign n1324 = n1317 | n1323 ;
  assign n1325 = x47 | x110 ;
  assign n1326 = x86 | x94 ;
  assign n1327 = n1215 | n1244 ;
  assign n1328 = n1326 | n1327 ;
  assign n1329 = n1243 | n1246 ;
  assign n1330 = x97 | n1329 ;
  assign n1331 = n1328 | n1330 ;
  assign n1332 = n1242 | n1331 ;
  assign n1333 = x108 & n1332 ;
  assign n1334 = x46 | n1333 ;
  assign n1335 = n1328 | n1329 ;
  assign n1336 = n1242 | n1335 ;
  assign n1337 = x97 & n1336 ;
  assign n1338 = x50 | n1215 ;
  assign n1339 = x77 | n1243 ;
  assign n1340 = n1242 | n1246 ;
  assign n1341 = n1339 | n1340 ;
  assign n1342 = n1338 | n1341 ;
  assign n1343 = ~x86 & x94 ;
  assign n1344 = ~n1342 & n1343 ;
  assign n1345 = x97 | n1344 ;
  assign n1346 = x86 & n1342 ;
  assign n1347 = x94 | n1346 ;
  assign n1348 = n1242 | n1329 ;
  assign n1349 = x77 & ~n1348 ;
  assign n1350 = x50 | n1349 ;
  assign n1351 = x64 & n1241 ;
  assign n1352 = n1226 | n1232 ;
  assign n1353 = n1235 | n1352 ;
  assign n1354 = x71 & n1353 ;
  assign n1355 = x65 | n1354 ;
  assign n1356 = x67 | n1352 ;
  assign n1357 = x69 & n1356 ;
  assign n1358 = n1234 | n1352 ;
  assign n1359 = x83 & n1358 ;
  assign n1360 = x103 | n1359 ;
  assign n1361 = n1357 | n1360 ;
  assign n1362 = x69 | x83 ;
  assign n1363 = x68 | x111 ;
  assign n1364 = n1226 | n1229 ;
  assign n1365 = x84 & n1364 ;
  assign n1366 = n1221 | n1222 ;
  assign n1367 = ( x61 & x85 ) | ( x61 & x106 ) | ( x85 & x106 ) ;
  assign n1368 = x61 | x106 ;
  assign n1369 = ( x76 & x85 ) | ( x76 & n1368 ) | ( x85 & n1368 ) ;
  assign n1370 = n1367 | n1369 ;
  assign n1371 = x48 | n1370 ;
  assign n1372 = n1221 & n1371 ;
  assign n1373 = x48 | n1221 ;
  assign n1374 = x89 & n1373 ;
  assign n1375 = x49 | n1374 ;
  assign n1376 = ( n1366 & n1372 ) | ( n1366 & n1375 ) | ( n1372 & n1375 ) ;
  assign n1377 = x45 | n1376 ;
  assign n1378 = ( x104 & n1224 ) | ( x104 & n1377 ) | ( n1224 & n1377 ) ;
  assign n1379 = n1226 & ~n1378 ;
  assign n1380 = n1229 | n1379 ;
  assign n1381 = ( x66 & x73 ) | ( x66 & n1226 ) | ( x73 & n1226 ) ;
  assign n1382 = n1380 & ~n1381 ;
  assign n1383 = x84 | n1382 ;
  assign n1384 = ~n1365 & n1383 ;
  assign n1385 = n1363 | n1384 ;
  assign n1386 = x84 | n1364 ;
  assign n1387 = x68 | n1386 ;
  assign n1388 = x111 & n1387 ;
  assign n1389 = x82 | n1388 ;
  assign n1390 = x68 & n1386 ;
  assign n1391 = n1389 | n1390 ;
  assign n1392 = n1385 & ~n1391 ;
  assign n1393 = x36 | x67 ;
  assign n1394 = x82 & ~n1363 ;
  assign n1395 = ~n1386 & n1394 ;
  assign n1396 = n1393 | n1395 ;
  assign n1397 = n1392 | n1396 ;
  assign n1398 = x67 & n1352 ;
  assign n1399 = n1227 | n1387 ;
  assign n1400 = x36 & n1399 ;
  assign n1401 = n1398 | n1400 ;
  assign n1402 = n1397 & ~n1401 ;
  assign n1403 = n1362 | n1402 ;
  assign n1404 = ~n1361 & n1403 ;
  assign n1405 = x103 & ~n1362 ;
  assign n1406 = ~n1356 & n1405 ;
  assign n1407 = x71 | n1406 ;
  assign n1408 = n1404 | n1407 ;
  assign n1409 = ~n1355 & n1408 ;
  assign n1410 = x107 | n1409 ;
  assign n1411 = x65 & ~x71 ;
  assign n1412 = ~n1353 & n1411 ;
  assign n1413 = n1410 | n1412 ;
  assign n1414 = n1235 | n1237 ;
  assign n1415 = n1352 | n1414 ;
  assign n1416 = x107 & n1415 ;
  assign n1417 = x63 | n1416 ;
  assign n1418 = n1413 & ~n1417 ;
  assign n1419 = x64 | n1418 ;
  assign n1420 = ~n1351 & n1419 ;
  assign n1421 = n1246 | n1420 ;
  assign n1422 = n1410 & ~n1417 ;
  assign n1423 = x63 & ~x107 ;
  assign n1424 = ~n1415 & n1423 ;
  assign n1425 = x64 | n1424 ;
  assign n1426 = n1422 | n1425 ;
  assign n1427 = ~n1351 & n1426 ;
  assign n1428 = n1421 | n1427 ;
  assign n1429 = ( x81 & x102 ) | ( x81 & n1242 ) | ( x102 & n1242 ) ;
  assign n1430 = n1428 & ~n1429 ;
  assign n1431 = n1243 | n1430 ;
  assign n1432 = x98 & n1340 ;
  assign n1433 = x77 | n1432 ;
  assign n1434 = x88 & x98 ;
  assign n1435 = ( x88 & n1246 ) | ( x88 & n1434 ) | ( n1246 & n1434 ) ;
  assign n1436 = ( x64 & x88 ) | ( x64 & n1435 ) | ( x88 & n1435 ) ;
  assign n1437 = x88 | n1435 ;
  assign n1438 = ( n1241 & n1436 ) | ( n1241 & n1437 ) | ( n1436 & n1437 ) ;
  assign n1439 = n1433 | n1438 ;
  assign n1440 = n1431 & ~n1439 ;
  assign n1441 = n1350 | n1440 ;
  assign n1442 = x50 & n1341 ;
  assign n1443 = x60 | n1442 ;
  assign n1444 = n1441 & ~n1443 ;
  assign n1445 = ~x53 & n1444 ;
  assign n1446 = x86 | n1445 ;
  assign n1447 = ~n1347 & n1446 ;
  assign n1448 = n1345 | n1447 ;
  assign n1449 = ~n1337 & n1448 ;
  assign n1450 = x108 | n1449 ;
  assign n1451 = ~n1334 & n1450 ;
  assign n1452 = x109 | n1451 ;
  assign n1453 = x109 & n1249 ;
  assign n1454 = n1325 | n1453 ;
  assign n1455 = n1452 & ~n1454 ;
  assign n1456 = ( ~n1324 & n1325 ) | ( ~n1324 & n1455 ) | ( n1325 & n1455 ) ;
  assign n1457 = n1315 | n1456 ;
  assign n1458 = ~n1310 & n1457 ;
  assign n1459 = x93 | n1458 ;
  assign n1460 = ~n1305 & n1459 ;
  assign n1461 = n1303 | n1460 ;
  assign n1462 = x70 | n1278 ;
  assign n1463 = n1272 | n1462 ;
  assign n1464 = x51 & n1463 ;
  assign n1465 = x96 | n1464 ;
  assign n1466 = n1280 | n1465 ;
  assign n1467 = n1461 & ~n1466 ;
  assign n1468 = x72 | n1467 ;
  assign n1469 = ~n1302 & n1468 ;
  assign n1470 = n1300 | n1469 ;
  assign n1471 = n1292 | n1470 ;
  assign n1472 = n1292 & ~n1300 ;
  assign n1473 = ~x97 & n1448 ;
  assign n1474 = x108 | n1473 ;
  assign n1475 = ~n1334 & n1474 ;
  assign n1476 = x109 | n1475 ;
  assign n1477 = ~n1454 & n1476 ;
  assign n1478 = ( ~n1324 & n1325 ) | ( ~n1324 & n1477 ) | ( n1325 & n1477 ) ;
  assign n1479 = n1315 | n1478 ;
  assign n1480 = ~n1310 & n1479 ;
  assign n1481 = x93 | n1480 ;
  assign n1482 = ~n1305 & n1481 ;
  assign n1483 = n1303 | n1482 ;
  assign n1484 = ~n1466 & n1483 ;
  assign n1485 = x72 | n1484 ;
  assign n1486 = ~n1302 & n1485 ;
  assign n1487 = n1472 & ~n1486 ;
  assign n1488 = n1264 | n1487 ;
  assign n1489 = n1471 & ~n1488 ;
  assign n1490 = x95 | n1489 ;
  assign n1491 = x95 & ~x479 ;
  assign n1492 = x32 | x40 ;
  assign n1493 = n1278 | n1492 ;
  assign n1494 = n1295 | n1493 ;
  assign n1495 = n1272 | n1494 ;
  assign n1496 = x95 & n1495 ;
  assign n1497 = n1491 | n1496 ;
  assign n1498 = x137 | n1497 ;
  assign n1499 = n1490 & ~n1498 ;
  assign n1500 = ( x137 & ~n1286 ) | ( x137 & n1499 ) | ( ~n1286 & n1499 ) ;
  assign n1501 = x210 | n1500 ;
  assign n1502 = x146 & ~n1501 ;
  assign n1503 = x234 & ~x332 ;
  assign n1504 = x225 | n1261 ;
  assign n1505 = x32 & n1504 ;
  assign n1506 = n1470 & ~n1505 ;
  assign n1507 = x95 | n1506 ;
  assign n1508 = ~n1498 & n1507 ;
  assign n1509 = x95 | n1505 ;
  assign n1510 = x137 & ~n1509 ;
  assign n1511 = n1284 & n1510 ;
  assign n1512 = x210 & ~n1511 ;
  assign n1513 = ~n1508 & n1512 ;
  assign n1514 = n1503 & ~n1513 ;
  assign n1515 = x146 | x210 ;
  assign n1516 = ~n1264 & n1470 ;
  assign n1517 = x95 | n1516 ;
  assign n1518 = ~n1498 & n1517 ;
  assign n1519 = ( x137 & ~n1286 ) | ( x137 & n1518 ) | ( ~n1286 & n1518 ) ;
  assign n1520 = n1515 | n1519 ;
  assign n1521 = n1514 & n1520 ;
  assign n1522 = ~n1502 & n1521 ;
  assign n1523 = x152 | x161 ;
  assign n1524 = x166 | n1523 ;
  assign n1525 = x35 | x70 ;
  assign n1526 = x51 | n1525 ;
  assign n1527 = x93 | n1269 ;
  assign n1528 = x91 | n1527 ;
  assign n1529 = n1526 | n1528 ;
  assign n1530 = n1313 | n1529 ;
  assign n1531 = x96 & ~n1530 ;
  assign n1532 = x72 | n1492 ;
  assign n1533 = n1531 & ~n1532 ;
  assign n1534 = n1284 | n1533 ;
  assign n1535 = ~n1265 & n1534 ;
  assign n1536 = n1491 & ~n1495 ;
  assign n1537 = x137 & ~n1536 ;
  assign n1538 = ~n1535 & n1537 ;
  assign n1539 = x72 | n1531 ;
  assign n1540 = n1467 | n1539 ;
  assign n1541 = ~n1302 & n1540 ;
  assign n1542 = n1300 | n1541 ;
  assign n1543 = n1292 | n1542 ;
  assign n1544 = n1484 | n1539 ;
  assign n1545 = ~n1302 & n1544 ;
  assign n1546 = n1472 & ~n1545 ;
  assign n1547 = n1264 | n1546 ;
  assign n1548 = n1543 & ~n1547 ;
  assign n1549 = x95 | n1548 ;
  assign n1550 = x137 | n1496 ;
  assign n1551 = n1549 & ~n1550 ;
  assign n1552 = ( x137 & ~n1538 ) | ( x137 & n1551 ) | ( ~n1538 & n1551 ) ;
  assign n1553 = x210 | n1552 ;
  assign n1554 = x146 & ~n1553 ;
  assign n1555 = x234 | x332 ;
  assign n1556 = ~n1509 & n1534 ;
  assign n1557 = n1536 | n1556 ;
  assign n1558 = x137 & n1557 ;
  assign n1559 = x210 & ~n1558 ;
  assign n1560 = ~n1509 & n1542 ;
  assign n1561 = ( x95 & ~n1550 ) | ( x95 & n1560 ) | ( ~n1550 & n1560 ) ;
  assign n1562 = n1559 & ~n1561 ;
  assign n1563 = n1555 | n1562 ;
  assign n1564 = ~n1264 & n1542 ;
  assign n1565 = x95 | n1564 ;
  assign n1566 = ~n1550 & n1565 ;
  assign n1567 = ( x137 & ~n1538 ) | ( x137 & n1566 ) | ( ~n1538 & n1566 ) ;
  assign n1568 = n1515 | n1567 ;
  assign n1569 = ~n1563 & n1568 ;
  assign n1570 = ~n1554 & n1569 ;
  assign n1571 = n1524 & ~n1570 ;
  assign n1572 = ~n1522 & n1571 ;
  assign n1573 = n1553 & ~n1563 ;
  assign n1574 = n1501 & n1514 ;
  assign n1575 = n1524 | n1574 ;
  assign n1576 = n1573 | n1575 ;
  assign n1577 = ~x153 & n1576 ;
  assign n1578 = ~n1572 & n1577 ;
  assign n1579 = x153 & ~x332 ;
  assign n1580 = x95 & x479 ;
  assign n1581 = x60 & ~n1248 ;
  assign n1582 = x53 | n1581 ;
  assign n1583 = x60 | n1248 ;
  assign n1584 = x53 & n1583 ;
  assign n1585 = n1326 | n1584 ;
  assign n1586 = n1582 & ~n1585 ;
  assign n1587 = x46 | n1250 ;
  assign n1588 = n1213 | n1266 ;
  assign n1589 = n1587 | n1588 ;
  assign n1590 = x58 | n1589 ;
  assign n1591 = n1255 | n1590 ;
  assign n1592 = n1586 & ~n1591 ;
  assign n1593 = x35 | n1592 ;
  assign n1594 = x35 & n1273 ;
  assign n1595 = n1303 | n1594 ;
  assign n1596 = n1593 & ~n1595 ;
  assign n1597 = x96 | n1596 ;
  assign n1598 = x96 & n1530 ;
  assign n1599 = n1212 | n1598 ;
  assign n1600 = n1597 & ~n1599 ;
  assign n1601 = x32 | n1600 ;
  assign n1602 = x51 | x72 ;
  assign n1603 = x841 & ~n1272 ;
  assign n1604 = ~x93 & n1603 ;
  assign n1605 = ~n1602 & n1604 ;
  assign n1606 = x35 | x40 ;
  assign n1607 = x225 & ~n1606 ;
  assign n1608 = ~n1256 & n1607 ;
  assign n1609 = n1605 & n1608 ;
  assign n1610 = x32 & ~n1609 ;
  assign n1611 = n1601 & ~n1610 ;
  assign n1612 = x95 | n1611 ;
  assign n1613 = ~n1580 & n1612 ;
  assign n1614 = ~n1291 & n1613 ;
  assign n1615 = ~x146 & n1524 ;
  assign n1616 = n1288 & ~n1615 ;
  assign n1617 = ~n1614 & n1616 ;
  assign n1618 = ~n1496 & n1613 ;
  assign n1619 = ~n1617 & n1618 ;
  assign n1620 = ~n1496 & n1616 ;
  assign n1621 = n1291 & ~n1580 ;
  assign n1622 = x97 | n1586 ;
  assign n1623 = x108 | n1337 ;
  assign n1624 = x110 | n1623 ;
  assign n1625 = x46 | x109 ;
  assign n1626 = n1266 | n1625 ;
  assign n1627 = n1527 | n1626 ;
  assign n1628 = n1624 | n1627 ;
  assign n1629 = n1622 & ~n1628 ;
  assign n1630 = x35 | n1629 ;
  assign n1631 = ~n1595 & n1630 ;
  assign n1632 = x96 | n1631 ;
  assign n1633 = ~n1599 & n1632 ;
  assign n1634 = x32 | n1633 ;
  assign n1635 = x95 | n1610 ;
  assign n1636 = n1634 & ~n1635 ;
  assign n1637 = ( x95 & n1621 ) | ( x95 & n1636 ) | ( n1621 & n1636 ) ;
  assign n1638 = n1620 & n1637 ;
  assign n1639 = x137 | n1638 ;
  assign n1640 = n1619 | n1639 ;
  assign n1641 = x40 | n1602 ;
  assign n1642 = n1279 | n1641 ;
  assign n1643 = n1531 & ~n1642 ;
  assign n1644 = ~x51 & x70 ;
  assign n1645 = n1465 | n1644 ;
  assign n1646 = n1275 | n1594 ;
  assign n1647 = x93 & ~n1272 ;
  assign n1648 = x35 | n1647 ;
  assign n1649 = x93 | n1309 ;
  assign n1650 = n1308 | n1649 ;
  assign n1651 = n1444 | n1582 ;
  assign n1652 = ~n1584 & n1651 ;
  assign n1653 = x86 | n1652 ;
  assign n1654 = ~n1347 & n1653 ;
  assign n1655 = n1345 | n1654 ;
  assign n1656 = ~n1337 & n1655 ;
  assign n1657 = x108 | n1656 ;
  assign n1658 = ~n1334 & n1657 ;
  assign n1659 = x109 | n1658 ;
  assign n1660 = ~n1454 & n1659 ;
  assign n1661 = ( ~n1324 & n1325 ) | ( ~n1324 & n1660 ) | ( n1325 & n1660 ) ;
  assign n1662 = n1315 | n1661 ;
  assign n1663 = ~n1650 & n1662 ;
  assign n1664 = n1648 | n1663 ;
  assign n1665 = ~n1646 & n1664 ;
  assign n1666 = x51 | n1665 ;
  assign n1667 = ~n1645 & n1666 ;
  assign n1668 = x72 | n1667 ;
  assign n1669 = ~n1302 & n1668 ;
  assign n1670 = n1300 | n1669 ;
  assign n1671 = n1643 | n1670 ;
  assign n1672 = ~n1610 & n1671 ;
  assign n1673 = x95 | n1672 ;
  assign n1674 = x137 & ~n1496 ;
  assign n1675 = n1673 & n1674 ;
  assign n1676 = ( ~x137 & n1640 ) | ( ~x137 & n1675 ) | ( n1640 & n1675 ) ;
  assign n1677 = x210 | n1676 ;
  assign n1678 = x234 & n1677 ;
  assign n1679 = ~n1635 & n1670 ;
  assign n1680 = ( x95 & ~n1497 ) | ( x95 & n1679 ) | ( ~n1497 & n1679 ) ;
  assign n1681 = x137 & ~n1680 ;
  assign n1682 = x40 | n1293 ;
  assign n1683 = n1596 & ~n1682 ;
  assign n1684 = x32 | n1683 ;
  assign n1685 = ~n1635 & n1684 ;
  assign n1686 = x137 | n1685 ;
  assign n1687 = x210 | x234 ;
  assign n1688 = ( n1615 & ~n1686 ) | ( n1615 & n1687 ) | ( ~n1686 & n1687 ) ;
  assign n1689 = ~n1292 & n1593 ;
  assign n1690 = x1091 & x1093 ;
  assign n1691 = ~n1287 & n1690 ;
  assign n1692 = x950 & x1092 ;
  assign n1693 = x829 & n1692 ;
  assign n1694 = n1691 & n1693 ;
  assign n1695 = n1630 & n1694 ;
  assign n1696 = n1689 | n1695 ;
  assign n1697 = n1595 | n1682 ;
  assign n1698 = n1696 & ~n1697 ;
  assign n1699 = x32 | n1698 ;
  assign n1700 = ~n1635 & n1699 ;
  assign n1701 = x137 | n1700 ;
  assign n1702 = ( n1615 & ~n1687 ) | ( n1615 & n1701 ) | ( ~n1687 & n1701 ) ;
  assign n1703 = ~n1688 & n1702 ;
  assign n1704 = ~n1681 & n1703 ;
  assign n1705 = x32 & ~n1262 ;
  assign n1706 = x95 | n1705 ;
  assign n1707 = n1670 & ~n1706 ;
  assign n1708 = ( x95 & ~n1497 ) | ( x95 & n1707 ) | ( ~n1497 & n1707 ) ;
  assign n1709 = x137 & ~n1708 ;
  assign n1710 = n1684 & ~n1706 ;
  assign n1711 = x137 | n1710 ;
  assign n1712 = x210 & n1711 ;
  assign n1713 = ~n1709 & n1712 ;
  assign n1714 = n1704 | n1713 ;
  assign n1715 = n1678 | n1714 ;
  assign n1716 = n1601 & ~n1706 ;
  assign n1717 = n1491 | n1716 ;
  assign n1718 = ~n1550 & n1717 ;
  assign n1719 = x210 & x234 ;
  assign n1720 = ~n1718 & n1719 ;
  assign n1721 = n1671 & ~n1706 ;
  assign n1722 = ( x95 & n1674 ) | ( x95 & n1721 ) | ( n1674 & n1721 ) ;
  assign n1723 = n1720 & ~n1722 ;
  assign n1724 = n1715 & ~n1723 ;
  assign n1725 = n1579 & ~n1724 ;
  assign n1726 = x228 | n1725 ;
  assign n1727 = n1578 | n1726 ;
  assign n1728 = x137 | n1717 ;
  assign n1729 = x46 & ~n1213 ;
  assign n1730 = ~n1336 & n1729 ;
  assign n1731 = x109 | n1730 ;
  assign n1732 = n1658 | n1731 ;
  assign n1733 = ~n1454 & n1732 ;
  assign n1734 = ( ~n1324 & n1325 ) | ( ~n1324 & n1733 ) | ( n1325 & n1733 ) ;
  assign n1735 = n1315 | n1734 ;
  assign n1736 = ~n1650 & n1735 ;
  assign n1737 = n1648 | n1736 ;
  assign n1738 = ~n1646 & n1737 ;
  assign n1739 = x51 | n1738 ;
  assign n1740 = ~n1645 & n1739 ;
  assign n1741 = x72 | n1740 ;
  assign n1742 = ~n1302 & n1741 ;
  assign n1743 = n1300 | n1742 ;
  assign n1744 = n1643 | n1743 ;
  assign n1745 = ~n1705 & n1744 ;
  assign n1746 = x95 | n1745 ;
  assign n1747 = x479 & n1496 ;
  assign n1748 = n1746 & ~n1747 ;
  assign n1749 = x137 & ~n1748 ;
  assign n1750 = n1728 & ~n1749 ;
  assign n1751 = x210 & ~n1750 ;
  assign n1752 = ~n1610 & n1744 ;
  assign n1753 = x95 | n1752 ;
  assign n1754 = ~n1747 & n1753 ;
  assign n1755 = x137 & ~n1754 ;
  assign n1756 = x137 | n1637 ;
  assign n1757 = n1614 | n1756 ;
  assign n1758 = ( n1288 & n1755 ) | ( n1288 & ~n1757 ) | ( n1755 & ~n1757 ) ;
  assign n1759 = x137 | n1613 ;
  assign n1760 = ( n1288 & ~n1755 ) | ( n1288 & n1759 ) | ( ~n1755 & n1759 ) ;
  assign n1761 = ~n1758 & n1760 ;
  assign n1762 = x210 | n1761 ;
  assign n1763 = ~n1751 & n1762 ;
  assign n1764 = ( x234 & x332 ) | ( x234 & n1763 ) | ( x332 & n1763 ) ;
  assign n1765 = ~n1706 & n1743 ;
  assign n1766 = ( x95 & ~n1497 ) | ( x95 & n1765 ) | ( ~n1497 & n1765 ) ;
  assign n1767 = x137 & ~n1766 ;
  assign n1768 = n1711 & ~n1767 ;
  assign n1769 = x210 & ~n1768 ;
  assign n1770 = ~n1610 & n1743 ;
  assign n1771 = x95 | n1770 ;
  assign n1772 = ~n1497 & n1771 ;
  assign n1773 = x137 & ~n1772 ;
  assign n1774 = n1701 & ~n1773 ;
  assign n1775 = x210 | n1774 ;
  assign n1776 = ~n1769 & n1775 ;
  assign n1777 = ( ~x234 & x332 ) | ( ~x234 & n1776 ) | ( x332 & n1776 ) ;
  assign n1778 = n1764 | n1777 ;
  assign n1779 = ~n1524 & n1778 ;
  assign n1780 = x146 & n1763 ;
  assign n1781 = ~n1755 & n1759 ;
  assign n1782 = x210 | n1781 ;
  assign n1783 = x146 | n1751 ;
  assign n1784 = n1782 & ~n1783 ;
  assign n1785 = n1503 & ~n1784 ;
  assign n1786 = ~n1780 & n1785 ;
  assign n1787 = n1686 & ~n1773 ;
  assign n1788 = x210 | n1787 ;
  assign n1789 = x146 | n1769 ;
  assign n1790 = n1788 & ~n1789 ;
  assign n1791 = x146 & n1776 ;
  assign n1792 = n1555 | n1791 ;
  assign n1793 = n1790 | n1792 ;
  assign n1794 = n1524 & n1793 ;
  assign n1795 = ~n1786 & n1794 ;
  assign n1796 = n1779 | n1795 ;
  assign n1797 = x105 & n1796 ;
  assign n1798 = x105 | n1579 ;
  assign n1799 = x228 & n1798 ;
  assign n1800 = ~n1797 & n1799 ;
  assign n1801 = ( ~x228 & n1727 ) | ( ~x228 & n1800 ) | ( n1727 & n1800 ) ;
  assign n1802 = x216 | n1801 ;
  assign n1803 = ~n1211 & n1802 ;
  assign n1804 = x221 | n1803 ;
  assign n1805 = ~n1209 & n1804 ;
  assign n1806 = x215 | n1805 ;
  assign n1807 = x332 | x1144 ;
  assign n1808 = x215 & n1807 ;
  assign n1809 = x299 & ~n1808 ;
  assign n1810 = n1806 & n1809 ;
  assign n1811 = ~x224 & x833 ;
  assign n1812 = x222 & ~n1811 ;
  assign n1813 = x223 | n1812 ;
  assign n1814 = ~n1807 & n1813 ;
  assign n1815 = x332 | x929 ;
  assign n1816 = n1811 & ~n1815 ;
  assign n1817 = ~x222 & x224 ;
  assign n1818 = ~n1210 & n1817 ;
  assign n1819 = ( x222 & ~n1816 ) | ( x222 & n1818 ) | ( ~n1816 & n1818 ) ;
  assign n1820 = x223 | n1819 ;
  assign n1821 = ~n1814 & n1820 ;
  assign n1822 = x299 | n1821 ;
  assign n1823 = x222 | x224 ;
  assign n1824 = x198 & ~n1750 ;
  assign n1825 = x198 | n1761 ;
  assign n1826 = ~n1824 & n1825 ;
  assign n1827 = x142 & n1826 ;
  assign n1828 = x198 | n1781 ;
  assign n1829 = x142 | n1824 ;
  assign n1830 = n1828 & ~n1829 ;
  assign n1831 = n1503 & ~n1830 ;
  assign n1832 = ~n1827 & n1831 ;
  assign n1833 = x144 | x174 ;
  assign n1834 = x189 | n1833 ;
  assign n1835 = ~x223 & n1834 ;
  assign n1836 = x198 | n1787 ;
  assign n1837 = x198 & ~n1768 ;
  assign n1838 = x142 | n1837 ;
  assign n1839 = n1836 & ~n1838 ;
  assign n1840 = x198 | n1774 ;
  assign n1841 = ~n1837 & n1840 ;
  assign n1842 = x142 & n1841 ;
  assign n1843 = n1555 | n1842 ;
  assign n1844 = n1839 | n1843 ;
  assign n1845 = n1835 & n1844 ;
  assign n1846 = ~n1832 & n1845 ;
  assign n1847 = x223 | n1834 ;
  assign n1848 = ( x234 & x332 ) | ( x234 & n1826 ) | ( x332 & n1826 ) ;
  assign n1849 = ( ~x234 & x332 ) | ( ~x234 & n1841 ) | ( x332 & n1841 ) ;
  assign n1850 = n1848 | n1849 ;
  assign n1851 = ~n1847 & n1850 ;
  assign n1852 = n1846 | n1851 ;
  assign n1853 = ~n1823 & n1852 ;
  assign n1854 = n1822 | n1853 ;
  assign n1855 = ~x39 & n1854 ;
  assign n1856 = ~n1810 & n1855 ;
  assign n1857 = x234 & n1491 ;
  assign n1858 = x332 | n1857 ;
  assign n1859 = x95 | n1494 ;
  assign n1860 = n1272 | n1859 ;
  assign n1861 = ~n1491 & n1860 ;
  assign n1862 = x234 & ~n1861 ;
  assign n1863 = x32 | x95 ;
  assign n1864 = n1212 | n1863 ;
  assign n1865 = n1277 | n1864 ;
  assign n1866 = n1462 | n1865 ;
  assign n1867 = n1271 | n1866 ;
  assign n1868 = n1242 | n1867 ;
  assign n1869 = x234 | n1868 ;
  assign n1870 = ~n1862 & n1869 ;
  assign n1871 = x137 & ~n1870 ;
  assign n1872 = n1858 | n1871 ;
  assign n1873 = x223 | n1823 ;
  assign n1874 = n1872 & ~n1873 ;
  assign n1875 = n1821 | n1874 ;
  assign n1876 = ~x299 & n1875 ;
  assign n1877 = x332 | n1860 ;
  assign n1878 = x137 | x153 ;
  assign n1879 = n1877 | n1878 ;
  assign n1880 = x137 & ~n1868 ;
  assign n1881 = n1579 & ~n1880 ;
  assign n1882 = x228 | n1881 ;
  assign n1883 = n1879 & ~n1882 ;
  assign n1884 = x105 & n1872 ;
  assign n1885 = n1799 & ~n1884 ;
  assign n1886 = ( x228 & n1883 ) | ( x228 & ~n1885 ) | ( n1883 & ~n1885 ) ;
  assign n1887 = ~x216 & n1886 ;
  assign n1888 = n1211 | n1887 ;
  assign n1889 = ~x221 & n1888 ;
  assign n1890 = n1209 | n1889 ;
  assign n1891 = ~x215 & n1890 ;
  assign n1892 = n1808 | n1891 ;
  assign n1893 = x299 & n1892 ;
  assign n1894 = n1876 | n1893 ;
  assign n1895 = x39 & n1894 ;
  assign n1896 = x38 | n1895 ;
  assign n1897 = n1856 | n1896 ;
  assign n1898 = x105 & x228 ;
  assign n1899 = ~n1858 & n1898 ;
  assign n1900 = n1579 & ~n1898 ;
  assign n1901 = x216 | n1900 ;
  assign n1902 = n1899 | n1901 ;
  assign n1903 = ~n1211 & n1902 ;
  assign n1904 = x221 | n1903 ;
  assign n1905 = ~n1209 & n1904 ;
  assign n1906 = x215 | n1905 ;
  assign n1907 = ~n1808 & n1906 ;
  assign n1908 = x215 | x221 ;
  assign n1909 = n1901 | n1908 ;
  assign n1910 = n1872 & ~n1909 ;
  assign n1911 = n1907 & ~n1910 ;
  assign n1912 = x299 & ~n1911 ;
  assign n1913 = n1876 | n1912 ;
  assign n1914 = ~x39 & n1913 ;
  assign n1915 = x299 & n1907 ;
  assign n1916 = n1858 & ~n1873 ;
  assign n1917 = n1822 | n1916 ;
  assign n1918 = ~n1915 & n1917 ;
  assign n1919 = x38 & ~x39 ;
  assign n1920 = ( x38 & ~n1918 ) | ( x38 & n1919 ) | ( ~n1918 & n1919 ) ;
  assign n1921 = ~n1914 & n1920 ;
  assign n1922 = x100 | n1921 ;
  assign n1923 = n1897 & ~n1922 ;
  assign n1924 = x87 | x100 ;
  assign n1925 = x38 | x39 ;
  assign n1926 = ~n1918 & n1925 ;
  assign n1927 = x142 & ~x198 ;
  assign n1928 = ( ~n1870 & n1871 ) | ( ~n1870 & n1927 ) | ( n1871 & n1927 ) ;
  assign n1929 = n1858 | n1928 ;
  assign n1930 = n1835 & n1929 ;
  assign n1931 = ~x137 & x198 ;
  assign n1932 = ~x95 & n1931 ;
  assign n1933 = n1861 | n1932 ;
  assign n1934 = n1503 & n1933 ;
  assign n1935 = n1868 | n1931 ;
  assign n1936 = ~n1555 & n1935 ;
  assign n1937 = n1847 | n1936 ;
  assign n1938 = n1934 | n1937 ;
  assign n1939 = ~n1930 & n1938 ;
  assign n1940 = n1823 | n1939 ;
  assign n1941 = ~n1821 & n1940 ;
  assign n1942 = x299 | n1941 ;
  assign n1943 = ~n1925 & n1942 ;
  assign n1944 = x210 | n1615 ;
  assign n1945 = x95 & x234 ;
  assign n1946 = x137 | n1945 ;
  assign n1947 = n1944 & ~n1946 ;
  assign n1948 = n1870 | n1947 ;
  assign n1949 = ~x332 & n1948 ;
  assign n1950 = x105 & ~n1949 ;
  assign n1951 = n1799 & ~n1950 ;
  assign n1952 = ~x137 & x210 ;
  assign n1953 = x252 | n1952 ;
  assign n1954 = n1615 | n1953 ;
  assign n1955 = n1877 | n1954 ;
  assign n1956 = n1615 & n1880 ;
  assign n1957 = n1579 & ~n1956 ;
  assign n1958 = n1955 & n1957 ;
  assign n1959 = x252 & ~n1615 ;
  assign n1960 = n1944 & ~n1959 ;
  assign n1961 = ~n1879 & n1960 ;
  assign n1962 = n1958 | n1961 ;
  assign n1963 = ~x228 & n1962 ;
  assign n1964 = x216 | n1963 ;
  assign n1965 = n1951 | n1964 ;
  assign n1966 = ~n1211 & n1965 ;
  assign n1967 = x221 | n1966 ;
  assign n1968 = ~n1209 & n1967 ;
  assign n1969 = x215 | n1968 ;
  assign n1970 = n1809 & n1969 ;
  assign n1971 = ( ~x299 & n1943 ) | ( ~x299 & n1970 ) | ( n1943 & n1970 ) ;
  assign n1972 = n1926 | n1971 ;
  assign n1973 = ( x87 & n1924 ) | ( x87 & ~n1972 ) | ( n1924 & ~n1972 ) ;
  assign n1974 = n1923 | n1973 ;
  assign n1975 = x38 | x100 ;
  assign n1976 = x39 | n1975 ;
  assign n1977 = ~n1918 & n1976 ;
  assign n1978 = n1894 | n1976 ;
  assign n1979 = ~n1977 & n1978 ;
  assign n1980 = x87 & ~n1979 ;
  assign n1981 = x75 | n1980 ;
  assign n1982 = n1974 & ~n1981 ;
  assign n1983 = x39 | x87 ;
  assign n1984 = n1975 | n1983 ;
  assign n1985 = ~n1918 & n1984 ;
  assign n1986 = x75 & ~n1985 ;
  assign n1987 = n1942 & ~n1984 ;
  assign n1988 = n1901 | n1951 ;
  assign n1989 = ~n1211 & n1988 ;
  assign n1990 = x221 | n1989 ;
  assign n1991 = ~n1209 & n1990 ;
  assign n1992 = x215 | n1991 ;
  assign n1993 = n1809 & n1992 ;
  assign n1994 = ( ~x299 & n1987 ) | ( ~x299 & n1993 ) | ( n1987 & n1993 ) ;
  assign n1995 = n1986 & ~n1994 ;
  assign n1996 = n1982 | n1995 ;
  assign n1997 = ~x92 & n1996 ;
  assign n1998 = x75 | x87 ;
  assign n1999 = ( x92 & n1918 ) | ( x92 & ~n1998 ) | ( n1918 & ~n1998 ) ;
  assign n2000 = ( x92 & n1979 ) | ( x92 & n1998 ) | ( n1979 & n1998 ) ;
  assign n2001 = n1999 & n2000 ;
  assign n2002 = x54 | n2001 ;
  assign n2003 = n1997 | n2002 ;
  assign n2004 = x75 | x92 ;
  assign n2005 = n1984 | n2004 ;
  assign n2006 = n1918 & n2005 ;
  assign n2007 = x38 | n1924 ;
  assign n2008 = n2004 | n2007 ;
  assign n2009 = n1914 & ~n2008 ;
  assign n2010 = n2006 | n2009 ;
  assign n2011 = x54 & ~n2010 ;
  assign n2012 = x74 | n2011 ;
  assign n2013 = n2003 & ~n2012 ;
  assign n2014 = ( x54 & x74 ) | ( x54 & n2010 ) | ( x74 & n2010 ) ;
  assign n2015 = ( ~x54 & x74 ) | ( ~x54 & n1918 ) | ( x74 & n1918 ) ;
  assign n2016 = n2014 & n2015 ;
  assign n2017 = n2013 | n2016 ;
  assign n2018 = ~x55 & n2017 ;
  assign n2019 = ~x332 & n1870 ;
  assign n2020 = x105 & ~n2019 ;
  assign n2021 = n1799 & ~n2020 ;
  assign n2022 = ~x228 & n1579 ;
  assign n2023 = n1868 & n2022 ;
  assign n2024 = x216 | n2023 ;
  assign n2025 = n2021 | n2024 ;
  assign n2026 = ~n1211 & n2025 ;
  assign n2027 = x221 | n2026 ;
  assign n2028 = ~n1209 & n2027 ;
  assign n2029 = x215 | n2028 ;
  assign n2030 = x54 | x74 ;
  assign n2031 = n2004 | n2030 ;
  assign n2032 = n1924 | n2031 ;
  assign n2033 = n1925 | n2032 ;
  assign n2034 = n1808 | n2033 ;
  assign n2035 = n2029 & ~n2034 ;
  assign n2036 = n1907 & n2033 ;
  assign n2037 = x55 & ~n2036 ;
  assign n2038 = ~n2035 & n2037 ;
  assign n2039 = x56 | n2038 ;
  assign n2040 = n2018 | n2039 ;
  assign n2041 = x100 | n1925 ;
  assign n2042 = x92 | n1998 ;
  assign n2043 = n2030 | n2042 ;
  assign n2044 = x55 | n2043 ;
  assign n2045 = n2041 | n2044 ;
  assign n2046 = n1907 & n2045 ;
  assign n2047 = n1892 | n2045 ;
  assign n2048 = ~n2046 & n2047 ;
  assign n2049 = x56 & ~n2048 ;
  assign n2050 = x62 | n2049 ;
  assign n2051 = n2040 & ~n2050 ;
  assign n2052 = ( x56 & ~x62 ) | ( x56 & n1907 ) | ( ~x62 & n1907 ) ;
  assign n2053 = ( x56 & x62 ) | ( x56 & n2048 ) | ( x62 & n2048 ) ;
  assign n2054 = ~n2052 & n2053 ;
  assign n2055 = x59 | n2054 ;
  assign n2056 = n2051 | n2055 ;
  assign n2057 = x57 | x59 ;
  assign n2058 = x56 | x62 ;
  assign n2059 = n2045 | n2058 ;
  assign n2060 = n1910 & ~n2059 ;
  assign n2061 = n1907 & ~n2060 ;
  assign n2062 = ( x57 & n2057 ) | ( x57 & n2061 ) | ( n2057 & n2061 ) ;
  assign n2063 = n2056 & ~n2062 ;
  assign n2064 = ~x59 & n2060 ;
  assign n2065 = n1907 & ~n2064 ;
  assign n2066 = x57 & ~n2065 ;
  assign n2067 = n2063 | n2066 ;
  assign n2068 = x223 & ~x1146 ;
  assign n2069 = x299 | n2068 ;
  assign n2070 = ( x222 & x939 ) | ( x222 & ~n1811 ) | ( x939 & ~n1811 ) ;
  assign n2071 = ( x222 & x1146 ) | ( x222 & n1811 ) | ( x1146 & n1811 ) ;
  assign n2072 = n2070 & n2071 ;
  assign n2073 = x223 | n2072 ;
  assign n2074 = ( x276 & n1817 ) | ( x276 & n2073 ) | ( n1817 & n2073 ) ;
  assign n2075 = n2073 | n2074 ;
  assign n2076 = ~n2069 & n2075 ;
  assign n2077 = x215 & x1146 ;
  assign n2078 = ( x221 & x939 ) | ( x221 & ~n1205 ) | ( x939 & ~n1205 ) ;
  assign n2079 = ( x221 & x1146 ) | ( x221 & n1205 ) | ( x1146 & n1205 ) ;
  assign n2080 = n2078 & n2079 ;
  assign n2081 = n2077 | n2080 ;
  assign n2082 = x228 | n1868 ;
  assign n2083 = x216 | n2082 ;
  assign n2084 = n2081 | n2083 ;
  assign n2085 = x216 & ~x221 ;
  assign n2086 = x276 & n2085 ;
  assign n2087 = x216 | n1898 ;
  assign n2088 = ~n2086 & n2087 ;
  assign n2089 = x221 | n2088 ;
  assign n2090 = ~n2080 & n2089 ;
  assign n2091 = x215 | n2090 ;
  assign n2092 = ~n2077 & n2091 ;
  assign n2093 = x299 & ~n2092 ;
  assign n2094 = n2084 & n2093 ;
  assign n2095 = n2076 | n2094 ;
  assign n2096 = ~x154 & n2095 ;
  assign n2097 = n2080 | n2086 ;
  assign n2098 = ~x215 & n2097 ;
  assign n2099 = n2077 | n2098 ;
  assign n2100 = x299 & n2099 ;
  assign n2101 = n2076 | n2100 ;
  assign n2102 = x154 & n2101 ;
  assign n2103 = n1976 | n2102 ;
  assign n2104 = n2096 | n2103 ;
  assign n2105 = n1998 | n2104 ;
  assign n2106 = x154 & n2099 ;
  assign n2107 = x154 | n2092 ;
  assign n2108 = ~n2106 & n2107 ;
  assign n2109 = x299 & ~n2108 ;
  assign n2110 = n2076 | n2109 ;
  assign n2111 = n1998 | n2041 ;
  assign n2112 = ~n2110 & n2111 ;
  assign n2113 = x92 & ~n2112 ;
  assign n2114 = n2105 & n2113 ;
  assign n2115 = n2030 | n2114 ;
  assign n2116 = ( x75 & x92 ) | ( x75 & ~n2110 ) | ( x92 & ~n2110 ) ;
  assign n2117 = n1976 & ~n2110 ;
  assign n2118 = n2104 & ~n2117 ;
  assign n2119 = x87 & ~n2118 ;
  assign n2120 = x39 & n1868 ;
  assign n2121 = x70 | n1664 ;
  assign n2122 = n1280 | n1594 ;
  assign n2123 = n2121 & ~n2122 ;
  assign n2124 = x51 | n2123 ;
  assign n2125 = ~n1465 & n2124 ;
  assign n2126 = n1539 | n2125 ;
  assign n2127 = ~n1301 & n2126 ;
  assign n2128 = n1492 | n2127 ;
  assign n2129 = x32 & n1261 ;
  assign n2130 = x40 & n1278 ;
  assign n2131 = ( x40 & n1295 ) | ( x40 & n2130 ) | ( n1295 & n2130 ) ;
  assign n2132 = ( x40 & n1271 ) | ( x40 & n2131 ) | ( n1271 & n2131 ) ;
  assign n2133 = x40 | n2131 ;
  assign n2134 = ( n1242 & n2132 ) | ( n1242 & n2133 ) | ( n2132 & n2133 ) ;
  assign n2135 = n2129 | n2134 ;
  assign n2136 = n2128 & ~n2135 ;
  assign n2137 = x95 | n2136 ;
  assign n2138 = ~n1496 & n2137 ;
  assign n2139 = x39 | n2138 ;
  assign n2140 = ~n2120 & n2139 ;
  assign n2141 = x216 | x228 ;
  assign n2142 = n2081 | n2141 ;
  assign n2143 = n2140 & ~n2142 ;
  assign n2144 = n2093 & ~n2143 ;
  assign n2145 = n2076 | n2144 ;
  assign n2146 = ~x154 & n2145 ;
  assign n2147 = x38 | n2102 ;
  assign n2148 = n2146 | n2147 ;
  assign n2149 = x38 & ~n2110 ;
  assign n2150 = x100 | n2149 ;
  assign n2151 = n2148 & ~n2150 ;
  assign n2152 = ~x146 & n1868 ;
  assign n2153 = x252 | n1868 ;
  assign n2154 = x146 & n2153 ;
  assign n2155 = n2152 | n2154 ;
  assign n2156 = x152 & n2155 ;
  assign n2157 = x161 | x166 ;
  assign n2158 = ( x152 & ~n2155 ) | ( x152 & n2157 ) | ( ~n2155 & n2157 ) ;
  assign n2159 = ( ~x152 & n2153 ) | ( ~x152 & n2157 ) | ( n2153 & n2157 ) ;
  assign n2160 = ~n2158 & n2159 ;
  assign n2161 = n2156 | n2160 ;
  assign n2162 = ~x154 & x299 ;
  assign n2163 = ~x39 & n2162 ;
  assign n2164 = x38 | n2141 ;
  assign n2165 = n2163 & ~n2164 ;
  assign n2166 = ~n2081 & n2165 ;
  assign n2167 = ~n2161 & n2166 ;
  assign n2168 = n2110 & ~n2167 ;
  assign n2169 = ( x87 & n1924 ) | ( x87 & n2168 ) | ( n1924 & n2168 ) ;
  assign n2170 = n2151 | n2169 ;
  assign n2171 = ~n2119 & n2170 ;
  assign n2172 = ( x75 & ~x92 ) | ( x75 & n2171 ) | ( ~x92 & n2171 ) ;
  assign n2173 = ~n2116 & n2172 ;
  assign n2174 = n2115 | n2173 ;
  assign n2175 = n2030 & ~n2110 ;
  assign n2176 = x55 | n2175 ;
  assign n2177 = n2174 & ~n2176 ;
  assign n2178 = n2084 | n2106 ;
  assign n2179 = n2033 | n2178 ;
  assign n2180 = x55 & ~n2108 ;
  assign n2181 = n2179 & n2180 ;
  assign n2182 = x56 | n2181 ;
  assign n2183 = n2177 | n2182 ;
  assign n2184 = x55 | n2033 ;
  assign n2185 = n2108 | n2184 ;
  assign n2186 = n2178 & ~n2185 ;
  assign n2187 = n2045 & ~n2108 ;
  assign n2188 = x56 & ~n2187 ;
  assign n2189 = ~n2186 & n2188 ;
  assign n2190 = x62 | n2189 ;
  assign n2191 = n2183 & ~n2190 ;
  assign n2192 = x56 | n2044 ;
  assign n2193 = n2041 | n2192 ;
  assign n2194 = ~n2108 & n2193 ;
  assign n2195 = n2186 | n2194 ;
  assign n2196 = x62 & n2195 ;
  assign n2197 = n2057 | n2196 ;
  assign n2198 = n2191 | n2197 ;
  assign n2199 = n2057 & n2108 ;
  assign n2200 = x239 | n2199 ;
  assign n2201 = n2198 & ~n2200 ;
  assign n2202 = x100 & n2167 ;
  assign n2203 = x216 | x221 ;
  assign n2204 = x215 | n2203 ;
  assign n2205 = n1491 & n1898 ;
  assign n2206 = ~n2204 & n2205 ;
  assign n2207 = n2099 | n2206 ;
  assign n2208 = x154 & n2207 ;
  assign n2209 = ~x215 & n2207 ;
  assign n2210 = n2107 & ~n2209 ;
  assign n2211 = ~n2208 & n2210 ;
  assign n2212 = x299 & ~n2211 ;
  assign n2213 = x223 | x299 ;
  assign n2214 = n1823 | n2213 ;
  assign n2215 = n1491 & ~n2214 ;
  assign n2216 = n2076 | n2215 ;
  assign n2217 = n2212 | n2216 ;
  assign n2218 = n1975 & n2217 ;
  assign n2219 = ~n2202 & n2218 ;
  assign n2220 = n2084 | n2208 ;
  assign n2221 = ~n2211 & n2220 ;
  assign n2222 = x299 & ~n2221 ;
  assign n2223 = n2217 & ~n2222 ;
  assign n2224 = ( x39 & n1975 ) | ( x39 & ~n2223 ) | ( n1975 & ~n2223 ) ;
  assign n2225 = x299 & ~n2099 ;
  assign n2226 = n1531 & ~n1864 ;
  assign n2227 = n1491 | n2226 ;
  assign n2228 = x105 & n2227 ;
  assign n2229 = x228 & ~n2228 ;
  assign n2230 = ~n1496 & n2227 ;
  assign n2231 = x228 | n2230 ;
  assign n2232 = ~n2229 & n2231 ;
  assign n2233 = ( x154 & n2204 ) | ( x154 & ~n2232 ) | ( n2204 & ~n2232 ) ;
  assign n2234 = x72 | n2125 ;
  assign n2235 = ~n1301 & n2234 ;
  assign n2236 = n1492 | n2235 ;
  assign n2237 = ~n2135 & n2236 ;
  assign n2238 = x95 | n2237 ;
  assign n2239 = ~n1497 & n2238 ;
  assign n2240 = ~x228 & n2239 ;
  assign n2241 = n1898 & ~n2227 ;
  assign n2242 = n2240 | n2241 ;
  assign n2243 = ( ~x154 & n2204 ) | ( ~x154 & n2242 ) | ( n2204 & n2242 ) ;
  assign n2244 = n2233 | n2243 ;
  assign n2245 = n2225 & n2244 ;
  assign n2246 = x224 | n2227 ;
  assign n2247 = x224 & ~x276 ;
  assign n2248 = x222 | n2247 ;
  assign n2249 = n2246 & ~n2248 ;
  assign n2250 = n2073 | n2249 ;
  assign n2251 = ~n2069 & n2250 ;
  assign n2252 = ( x299 & ~n2245 ) | ( x299 & n2251 ) | ( ~n2245 & n2251 ) ;
  assign n2253 = ( x39 & ~n1975 ) | ( x39 & n2252 ) | ( ~n1975 & n2252 ) ;
  assign n2254 = ~n2224 & n2253 ;
  assign n2255 = n2219 | n2254 ;
  assign n2256 = ~x87 & n2255 ;
  assign n2257 = ~n1976 & n2222 ;
  assign n2258 = n2217 & ~n2257 ;
  assign n2259 = ( x75 & n1998 ) | ( x75 & n2258 ) | ( n1998 & n2258 ) ;
  assign n2260 = n2256 | n2259 ;
  assign n2261 = x75 & ~n2217 ;
  assign n2262 = x92 | n2261 ;
  assign n2263 = n2260 & ~n2262 ;
  assign n2264 = ~n2111 & n2222 ;
  assign n2265 = x92 & n2217 ;
  assign n2266 = ~n2264 & n2265 ;
  assign n2267 = n2030 | n2266 ;
  assign n2268 = n2263 | n2267 ;
  assign n2269 = n2030 & ~n2217 ;
  assign n2270 = x55 | n2269 ;
  assign n2271 = n2268 & ~n2270 ;
  assign n2272 = n2033 | n2220 ;
  assign n2273 = x55 & ~n2211 ;
  assign n2274 = n2272 & n2273 ;
  assign n2275 = x56 | n2274 ;
  assign n2276 = n2271 | n2275 ;
  assign n2277 = ~n2184 & n2221 ;
  assign n2278 = n2045 & ~n2211 ;
  assign n2279 = x56 & ~n2278 ;
  assign n2280 = ~n2277 & n2279 ;
  assign n2281 = x62 | n2280 ;
  assign n2282 = n2276 & ~n2281 ;
  assign n2283 = n2193 & ~n2211 ;
  assign n2284 = ~x56 & n2277 ;
  assign n2285 = n2283 | n2284 ;
  assign n2286 = x62 & n2285 ;
  assign n2287 = n2057 | n2286 ;
  assign n2288 = n2282 | n2287 ;
  assign n2289 = n2057 & n2211 ;
  assign n2290 = x239 & ~n2289 ;
  assign n2291 = n2288 & n2290 ;
  assign n2292 = n2201 | n2291 ;
  assign n2293 = x216 & x274 ;
  assign n2294 = x221 | n2293 ;
  assign n2295 = ( x151 & ~x216 ) | ( x151 & n2242 ) | ( ~x216 & n2242 ) ;
  assign n2296 = ( x151 & x216 ) | ( x151 & n2232 ) | ( x216 & n2232 ) ;
  assign n2297 = n2295 & ~n2296 ;
  assign n2298 = n2294 | n2297 ;
  assign n2299 = ( x221 & x927 ) | ( x221 & ~n1205 ) | ( x927 & ~n1205 ) ;
  assign n2300 = ( x221 & x1145 ) | ( x221 & n1205 ) | ( x1145 & n1205 ) ;
  assign n2301 = n2299 & n2300 ;
  assign n2302 = n2298 & ~n2301 ;
  assign n2303 = x215 | n2302 ;
  assign n2304 = x215 & x1145 ;
  assign n2305 = x299 & ~n2304 ;
  assign n2306 = n2303 & n2305 ;
  assign n2307 = x224 & x274 ;
  assign n2308 = x222 | n2307 ;
  assign n2309 = n2246 & ~n2308 ;
  assign n2310 = ( x222 & x927 ) | ( x222 & ~n1811 ) | ( x927 & ~n1811 ) ;
  assign n2311 = ( x222 & x1145 ) | ( x222 & n1811 ) | ( x1145 & n1811 ) ;
  assign n2312 = n2310 & n2311 ;
  assign n2313 = n2309 | n2312 ;
  assign n2314 = ~x223 & n2313 ;
  assign n2315 = x223 & x1145 ;
  assign n2316 = x299 | n2315 ;
  assign n2317 = n2314 | n2316 ;
  assign n2318 = ~x39 & n2317 ;
  assign n2319 = ~n2306 & n2318 ;
  assign n2320 = n1817 & ~n2307 ;
  assign n2321 = n2312 | n2320 ;
  assign n2322 = ~x223 & n2321 ;
  assign n2323 = n2315 | n2322 ;
  assign n2324 = ~x299 & n2323 ;
  assign n2325 = n2215 | n2324 ;
  assign n2326 = x151 | n1898 ;
  assign n2327 = ~n2205 & n2326 ;
  assign n2328 = x151 | n2082 ;
  assign n2329 = ~n2327 & n2328 ;
  assign n2330 = x216 | n2329 ;
  assign n2331 = ~n2294 & n2330 ;
  assign n2332 = n2301 | n2331 ;
  assign n2333 = ~x215 & n2332 ;
  assign n2334 = n2304 | n2333 ;
  assign n2335 = x299 & n2334 ;
  assign n2336 = n2325 | n2335 ;
  assign n2337 = x39 & n2336 ;
  assign n2338 = x38 | n2337 ;
  assign n2339 = n2319 | n2338 ;
  assign n2340 = ~x216 & n2326 ;
  assign n2341 = n2294 | n2340 ;
  assign n2342 = ~n2301 & n2341 ;
  assign n2343 = x215 | n2342 ;
  assign n2344 = ~n2304 & n2343 ;
  assign n2345 = ~n1908 & n2205 ;
  assign n2346 = ~n2293 & n2345 ;
  assign n2347 = n2344 & ~n2346 ;
  assign n2348 = x299 & ~n2347 ;
  assign n2349 = n2325 | n2348 ;
  assign n2350 = x38 & ~n2349 ;
  assign n2351 = x100 | n2350 ;
  assign n2352 = n2339 & ~n2351 ;
  assign n2353 = n1925 | n2325 ;
  assign n2354 = x228 | n2161 ;
  assign n2355 = ~n1491 & n1898 ;
  assign n2356 = n2354 & ~n2355 ;
  assign n2357 = ~x151 & n2356 ;
  assign n2358 = n2330 | n2357 ;
  assign n2359 = ~n2294 & n2358 ;
  assign n2360 = n2301 | n2359 ;
  assign n2361 = ~x215 & n2360 ;
  assign n2362 = n2305 & ~n2361 ;
  assign n2363 = ( x299 & n2353 ) | ( x299 & ~n2362 ) | ( n2353 & ~n2362 ) ;
  assign n2364 = x100 & ~n1925 ;
  assign n2365 = ( x100 & n2349 ) | ( x100 & n2364 ) | ( n2349 & n2364 ) ;
  assign n2366 = n2363 & n2365 ;
  assign n2367 = n2352 | n2366 ;
  assign n2368 = ~x87 & n2367 ;
  assign n2369 = n1976 & ~n2349 ;
  assign n2370 = n1976 | n2336 ;
  assign n2371 = ~n2369 & n2370 ;
  assign n2372 = ( x75 & n1998 ) | ( x75 & n2371 ) | ( n1998 & n2371 ) ;
  assign n2373 = n2368 | n2372 ;
  assign n2374 = x75 & ~n2349 ;
  assign n2375 = x92 | n2374 ;
  assign n2376 = n2373 & ~n2375 ;
  assign n2377 = ( x92 & ~n1998 ) | ( x92 & n2349 ) | ( ~n1998 & n2349 ) ;
  assign n2378 = ( x92 & n1998 ) | ( x92 & n2371 ) | ( n1998 & n2371 ) ;
  assign n2379 = n2377 & n2378 ;
  assign n2380 = n2030 | n2379 ;
  assign n2381 = n2376 | n2380 ;
  assign n2382 = n2030 & ~n2349 ;
  assign n2383 = x55 | n2382 ;
  assign n2384 = n2381 & ~n2383 ;
  assign n2385 = ( x55 & n2033 ) | ( x55 & n2334 ) | ( n2033 & n2334 ) ;
  assign n2386 = ( ~x55 & n2033 ) | ( ~x55 & n2347 ) | ( n2033 & n2347 ) ;
  assign n2387 = n2385 & ~n2386 ;
  assign n2388 = x56 | n2387 ;
  assign n2389 = n2384 | n2388 ;
  assign n2390 = ( x56 & n2045 ) | ( x56 & ~n2334 ) | ( n2045 & ~n2334 ) ;
  assign n2391 = ( x56 & ~n2045 ) | ( x56 & n2347 ) | ( ~n2045 & n2347 ) ;
  assign n2392 = n2390 & n2391 ;
  assign n2393 = x62 | n2392 ;
  assign n2394 = n2389 & ~n2393 ;
  assign n2395 = x235 & ~n2057 ;
  assign n2396 = ( x62 & n2193 ) | ( x62 & n2334 ) | ( n2193 & n2334 ) ;
  assign n2397 = ( ~x62 & n2193 ) | ( ~x62 & n2347 ) | ( n2193 & n2347 ) ;
  assign n2398 = n2396 & ~n2397 ;
  assign n2399 = n2395 & ~n2398 ;
  assign n2400 = ~n2394 & n2399 ;
  assign n2401 = n2301 | n2304 ;
  assign n2402 = n2083 | n2401 ;
  assign n2403 = x299 & ~n2344 ;
  assign n2404 = n2402 & n2403 ;
  assign n2405 = n2041 | n2324 ;
  assign n2406 = n2404 | n2405 ;
  assign n2407 = n1998 | n2406 ;
  assign n2408 = n2324 | n2403 ;
  assign n2409 = n2111 & ~n2408 ;
  assign n2410 = x92 & ~n2409 ;
  assign n2411 = n2407 & n2410 ;
  assign n2412 = n2030 | n2411 ;
  assign n2413 = ( x75 & x92 ) | ( x75 & ~n2408 ) | ( x92 & ~n2408 ) ;
  assign n2414 = n1976 & ~n2408 ;
  assign n2415 = n2406 & ~n2414 ;
  assign n2416 = x87 & ~n2415 ;
  assign n2417 = ~x100 & n2140 ;
  assign n2418 = ~x39 & x100 ;
  assign n2419 = ~n2161 & n2418 ;
  assign n2420 = n2417 | n2419 ;
  assign n2421 = n2164 | n2401 ;
  assign n2422 = n2420 & ~n2421 ;
  assign n2423 = n2403 & ~n2422 ;
  assign n2424 = x87 | n2324 ;
  assign n2425 = n2423 | n2424 ;
  assign n2426 = ~n2416 & n2425 ;
  assign n2427 = ( x75 & ~x92 ) | ( x75 & n2426 ) | ( ~x92 & n2426 ) ;
  assign n2428 = ~n2413 & n2427 ;
  assign n2429 = n2412 | n2428 ;
  assign n2430 = n2030 & ~n2408 ;
  assign n2431 = x55 | n2430 ;
  assign n2432 = n2429 & ~n2431 ;
  assign n2433 = n2033 | n2402 ;
  assign n2434 = x55 & ~n2344 ;
  assign n2435 = n2433 & n2434 ;
  assign n2436 = x56 | n2435 ;
  assign n2437 = n2432 | n2436 ;
  assign n2438 = n2045 | n2402 ;
  assign n2439 = ~n2344 & n2438 ;
  assign n2440 = x56 & ~n2439 ;
  assign n2441 = x62 | n2440 ;
  assign n2442 = n2437 & ~n2441 ;
  assign n2443 = x56 | n2438 ;
  assign n2444 = x62 & ~n2344 ;
  assign n2445 = n2443 & n2444 ;
  assign n2446 = x235 | n2057 ;
  assign n2447 = n2445 | n2446 ;
  assign n2448 = n2442 | n2447 ;
  assign n2449 = x235 & n2346 ;
  assign n2450 = n2057 & ~n2449 ;
  assign n2451 = n2344 & n2450 ;
  assign n2452 = n2448 & ~n2451 ;
  assign n2453 = ~n2400 & n2452 ;
  assign n2454 = x223 & x1143 ;
  assign n2455 = x299 | n2454 ;
  assign n2456 = x224 & x264 ;
  assign n2457 = x222 | n2456 ;
  assign n2458 = x284 | n2227 ;
  assign n2459 = ~x224 & n2458 ;
  assign n2460 = n2457 | n2459 ;
  assign n2461 = ( x222 & x944 ) | ( x222 & ~n1811 ) | ( x944 & ~n1811 ) ;
  assign n2462 = ( x222 & x1143 ) | ( x222 & n1811 ) | ( x1143 & n1811 ) ;
  assign n2463 = n2461 & n2462 ;
  assign n2464 = n2460 & ~n2463 ;
  assign n2465 = n2227 & ~n2457 ;
  assign n2466 = n2464 & ~n2465 ;
  assign n2467 = x223 | n2466 ;
  assign n2468 = ~n2455 & n2467 ;
  assign n2469 = x39 | n2468 ;
  assign n2470 = x215 & x1143 ;
  assign n2471 = x299 & ~n2470 ;
  assign n2472 = x216 & x264 ;
  assign n2473 = x221 | n2472 ;
  assign n2474 = x284 & ~n1491 ;
  assign n2475 = ( ~x105 & x228 ) | ( ~x105 & n2474 ) | ( x228 & n2474 ) ;
  assign n2476 = ( x105 & ~x146 ) | ( x105 & x228 ) | ( ~x146 & x228 ) ;
  assign n2477 = n2475 & n2476 ;
  assign n2478 = ~n2228 & n2477 ;
  assign n2479 = x146 | x284 ;
  assign n2480 = n2138 | n2479 ;
  assign n2481 = ( ~x146 & x284 ) | ( ~x146 & n2239 ) | ( x284 & n2239 ) ;
  assign n2482 = ( x146 & x284 ) | ( x146 & ~n2230 ) | ( x284 & ~n2230 ) ;
  assign n2483 = n2481 & n2482 ;
  assign n2484 = n2480 & ~n2483 ;
  assign n2485 = x228 | n2484 ;
  assign n2486 = ~n2478 & n2485 ;
  assign n2487 = x216 | n2486 ;
  assign n2488 = ~n2473 & n2487 ;
  assign n2489 = ( x221 & x944 ) | ( x221 & ~n1205 ) | ( x944 & ~n1205 ) ;
  assign n2490 = ( x221 & x1143 ) | ( x221 & n1205 ) | ( x1143 & n1205 ) ;
  assign n2491 = n2489 & n2490 ;
  assign n2492 = n2488 | n2491 ;
  assign n2493 = ~x215 & n2492 ;
  assign n2494 = n2471 & ~n2493 ;
  assign n2495 = n2469 | n2494 ;
  assign n2496 = ~x224 & n2474 ;
  assign n2497 = n2457 | n2496 ;
  assign n2498 = ~n2463 & n2497 ;
  assign n2499 = x223 | n2498 ;
  assign n2500 = ~n2454 & n2499 ;
  assign n2501 = x299 | n2500 ;
  assign n2502 = x284 & ~n1868 ;
  assign n2503 = n2152 | n2502 ;
  assign n2504 = ~x228 & n2503 ;
  assign n2505 = n2477 | n2504 ;
  assign n2506 = ~x216 & n2505 ;
  assign n2507 = n2473 | n2506 ;
  assign n2508 = ~n2491 & n2507 ;
  assign n2509 = x215 | n2508 ;
  assign n2510 = ~n2470 & n2509 ;
  assign n2511 = x299 & ~n2510 ;
  assign n2512 = n2501 & ~n2511 ;
  assign n2513 = x39 & ~n2512 ;
  assign n2514 = x38 | n2513 ;
  assign n2515 = n2495 & ~n2514 ;
  assign n2516 = n2205 | n2477 ;
  assign n2517 = x146 | x228 ;
  assign n2518 = ~n2516 & n2517 ;
  assign n2519 = x216 | n2518 ;
  assign n2520 = ~n2473 & n2519 ;
  assign n2521 = n2491 | n2520 ;
  assign n2522 = ~x215 & n2521 ;
  assign n2523 = n2470 | n2522 ;
  assign n2524 = n2345 & ~n2472 ;
  assign n2525 = n2523 | n2524 ;
  assign n2526 = x299 & n2525 ;
  assign n2527 = n2501 & ~n2526 ;
  assign n2528 = x38 & n2527 ;
  assign n2529 = x100 | n2528 ;
  assign n2530 = n2515 | n2529 ;
  assign n2531 = ~n1925 & n2501 ;
  assign n2532 = x252 & ~n1524 ;
  assign n2533 = x284 | n2532 ;
  assign n2534 = n1868 | n2533 ;
  assign n2535 = ~x228 & n2534 ;
  assign n2536 = ~n2154 & n2535 ;
  assign n2537 = n2477 | n2536 ;
  assign n2538 = ~x216 & n2537 ;
  assign n2539 = n2473 | n2538 ;
  assign n2540 = ~n2491 & n2539 ;
  assign n2541 = x215 | n2540 ;
  assign n2542 = n2471 & n2541 ;
  assign n2543 = ( ~x299 & n2531 ) | ( ~x299 & n2542 ) | ( n2531 & n2542 ) ;
  assign n2544 = ( x100 & n2364 ) | ( x100 & ~n2527 ) | ( n2364 & ~n2527 ) ;
  assign n2545 = ~n2543 & n2544 ;
  assign n2546 = n2530 & ~n2545 ;
  assign n2547 = x87 | n2546 ;
  assign n2548 = n1976 & n2527 ;
  assign n2549 = ~n1976 & n2512 ;
  assign n2550 = n2548 | n2549 ;
  assign n2551 = ( x75 & n1998 ) | ( x75 & ~n2550 ) | ( n1998 & ~n2550 ) ;
  assign n2552 = n2547 & ~n2551 ;
  assign n2553 = x75 & n2527 ;
  assign n2554 = x92 | n2553 ;
  assign n2555 = n2552 | n2554 ;
  assign n2556 = ( ~x92 & n1998 ) | ( ~x92 & n2527 ) | ( n1998 & n2527 ) ;
  assign n2557 = ( x92 & n1998 ) | ( x92 & ~n2550 ) | ( n1998 & ~n2550 ) ;
  assign n2558 = ~n2556 & n2557 ;
  assign n2559 = n2030 | n2558 ;
  assign n2560 = n2555 & ~n2559 ;
  assign n2561 = n2030 & n2527 ;
  assign n2562 = x55 | n2561 ;
  assign n2563 = n2560 | n2562 ;
  assign n2564 = ( x55 & n2033 ) | ( x55 & ~n2510 ) | ( n2033 & ~n2510 ) ;
  assign n2565 = ( x55 & ~n2033 ) | ( x55 & n2525 ) | ( ~n2033 & n2525 ) ;
  assign n2566 = n2564 & n2565 ;
  assign n2567 = x56 | n2566 ;
  assign n2568 = n2563 & ~n2567 ;
  assign n2569 = ( x56 & n2045 ) | ( x56 & n2510 ) | ( n2045 & n2510 ) ;
  assign n2570 = ( ~x56 & n2045 ) | ( ~x56 & n2525 ) | ( n2045 & n2525 ) ;
  assign n2571 = n2569 & ~n2570 ;
  assign n2572 = x62 | n2571 ;
  assign n2573 = n2568 | n2572 ;
  assign n2574 = x238 & ~n2057 ;
  assign n2575 = ( x62 & n2193 ) | ( x62 & ~n2510 ) | ( n2193 & ~n2510 ) ;
  assign n2576 = ( x62 & ~n2193 ) | ( x62 & n2525 ) | ( ~n2193 & n2525 ) ;
  assign n2577 = n2575 & n2576 ;
  assign n2578 = n2574 & ~n2577 ;
  assign n2579 = n2573 & n2578 ;
  assign n2580 = x146 | n2239 ;
  assign n2581 = x146 | n2138 ;
  assign n2582 = ( x284 & n2138 ) | ( x284 & ~n2581 ) | ( n2138 & ~n2581 ) ;
  assign n2583 = ~x146 & n2230 ;
  assign n2584 = ( x284 & n2230 ) | ( x284 & n2583 ) | ( n2230 & n2583 ) ;
  assign n2585 = ( n2230 & n2582 ) | ( n2230 & ~n2584 ) | ( n2582 & ~n2584 ) ;
  assign n2586 = n2580 & ~n2585 ;
  assign n2587 = x228 | n2586 ;
  assign n2588 = n1898 & n2227 ;
  assign n2589 = n2477 | n2588 ;
  assign n2590 = n2587 & ~n2589 ;
  assign n2591 = x216 | n2590 ;
  assign n2592 = ~n2473 & n2591 ;
  assign n2593 = n2491 | n2592 ;
  assign n2594 = ~x215 & n2593 ;
  assign n2595 = n2471 & ~n2594 ;
  assign n2596 = ~n2455 & n2464 ;
  assign n2597 = n2469 | n2596 ;
  assign n2598 = n2595 | n2597 ;
  assign n2599 = n1491 & ~n1873 ;
  assign n2600 = n2501 | n2599 ;
  assign n2601 = n2504 | n2516 ;
  assign n2602 = ~x216 & n2601 ;
  assign n2603 = n2473 | n2602 ;
  assign n2604 = ~n2491 & n2603 ;
  assign n2605 = x215 | n2604 ;
  assign n2606 = ~n2470 & n2605 ;
  assign n2607 = x299 & ~n2606 ;
  assign n2608 = n2600 & ~n2607 ;
  assign n2609 = x39 & ~n2608 ;
  assign n2610 = x38 | n2609 ;
  assign n2611 = n2598 & ~n2610 ;
  assign n2612 = x299 & n2523 ;
  assign n2613 = n2600 & ~n2612 ;
  assign n2614 = x38 & n2613 ;
  assign n2615 = x100 | n2614 ;
  assign n2616 = n2611 | n2615 ;
  assign n2617 = ~n1925 & n2600 ;
  assign n2618 = n2516 | n2536 ;
  assign n2619 = ~x216 & n2618 ;
  assign n2620 = n2473 | n2619 ;
  assign n2621 = ~n2491 & n2620 ;
  assign n2622 = x215 | n2621 ;
  assign n2623 = n2471 & n2622 ;
  assign n2624 = ( ~x299 & n2617 ) | ( ~x299 & n2623 ) | ( n2617 & n2623 ) ;
  assign n2625 = ( x100 & n2364 ) | ( x100 & ~n2613 ) | ( n2364 & ~n2613 ) ;
  assign n2626 = ~n2624 & n2625 ;
  assign n2627 = n2616 & ~n2626 ;
  assign n2628 = x87 | n2627 ;
  assign n2629 = n1976 & n2613 ;
  assign n2630 = ~n1976 & n2608 ;
  assign n2631 = n2629 | n2630 ;
  assign n2632 = ( x75 & n1998 ) | ( x75 & ~n2631 ) | ( n1998 & ~n2631 ) ;
  assign n2633 = n2628 & ~n2632 ;
  assign n2634 = x75 & n2613 ;
  assign n2635 = x92 | n2634 ;
  assign n2636 = n2633 | n2635 ;
  assign n2637 = ( ~x92 & n1998 ) | ( ~x92 & n2613 ) | ( n1998 & n2613 ) ;
  assign n2638 = ( x92 & n1998 ) | ( x92 & ~n2631 ) | ( n1998 & ~n2631 ) ;
  assign n2639 = ~n2637 & n2638 ;
  assign n2640 = n2030 | n2639 ;
  assign n2641 = n2636 & ~n2640 ;
  assign n2642 = n2030 & n2613 ;
  assign n2643 = x55 | n2642 ;
  assign n2644 = n2641 | n2643 ;
  assign n2645 = ( x55 & n2033 ) | ( x55 & ~n2606 ) | ( n2033 & ~n2606 ) ;
  assign n2646 = ( x55 & ~n2033 ) | ( x55 & n2523 ) | ( ~n2033 & n2523 ) ;
  assign n2647 = n2645 & n2646 ;
  assign n2648 = x56 | n2647 ;
  assign n2649 = n2644 & ~n2648 ;
  assign n2650 = ( x56 & n2045 ) | ( x56 & n2606 ) | ( n2045 & n2606 ) ;
  assign n2651 = ( ~x56 & n2045 ) | ( ~x56 & n2523 ) | ( n2045 & n2523 ) ;
  assign n2652 = n2650 & ~n2651 ;
  assign n2653 = x62 | n2652 ;
  assign n2654 = n2649 | n2653 ;
  assign n2655 = x238 | n2057 ;
  assign n2656 = ( x62 & n2193 ) | ( x62 & ~n2606 ) | ( n2193 & ~n2606 ) ;
  assign n2657 = ( x62 & ~n2193 ) | ( x62 & n2523 ) | ( ~n2193 & n2523 ) ;
  assign n2658 = n2656 & n2657 ;
  assign n2659 = n2655 | n2658 ;
  assign n2660 = n2654 & ~n2659 ;
  assign n2661 = x238 & n2524 ;
  assign n2662 = n2057 & ~n2661 ;
  assign n2663 = ~n2523 & n2662 ;
  assign n2664 = n2660 | n2663 ;
  assign n2665 = n2579 | n2664 ;
  assign n2666 = x215 & x1142 ;
  assign n2667 = x299 & ~n2666 ;
  assign n2668 = x216 & x277 ;
  assign n2669 = x221 | n2668 ;
  assign n2670 = x262 & n2138 ;
  assign n2671 = x228 | n2670 ;
  assign n2672 = x262 & n2239 ;
  assign n2673 = ( x172 & ~n2239 ) | ( x172 & n2672 ) | ( ~n2239 & n2672 ) ;
  assign n2674 = x262 & n2230 ;
  assign n2675 = ( x172 & n2230 ) | ( x172 & n2674 ) | ( n2230 & n2674 ) ;
  assign n2676 = ( n2230 & n2673 ) | ( n2230 & ~n2675 ) | ( n2673 & ~n2675 ) ;
  assign n2677 = n2671 | n2676 ;
  assign n2678 = x262 & ~n1491 ;
  assign n2679 = x105 & n2678 ;
  assign n2680 = ~n2226 & n2679 ;
  assign n2681 = ~x105 & x172 ;
  assign n2682 = x228 & ~n2681 ;
  assign n2683 = ~n2680 & n2682 ;
  assign n2684 = ~n2228 & n2683 ;
  assign n2685 = x216 | n2684 ;
  assign n2686 = n2677 & ~n2685 ;
  assign n2687 = n2669 | n2686 ;
  assign n2688 = ( x221 & x932 ) | ( x221 & ~n1205 ) | ( x932 & ~n1205 ) ;
  assign n2689 = ( x221 & x1142 ) | ( x221 & n1205 ) | ( x1142 & n1205 ) ;
  assign n2690 = n2688 & n2689 ;
  assign n2691 = n2687 & ~n2690 ;
  assign n2692 = x215 | n2691 ;
  assign n2693 = n2667 & n2692 ;
  assign n2694 = x223 & x1142 ;
  assign n2695 = x299 | n2694 ;
  assign n2696 = x224 & x277 ;
  assign n2697 = x222 | n2696 ;
  assign n2698 = x262 | n2227 ;
  assign n2699 = ~x224 & n2698 ;
  assign n2700 = n2697 | n2699 ;
  assign n2701 = ( x222 & x932 ) | ( x222 & ~n1811 ) | ( x932 & ~n1811 ) ;
  assign n2702 = ( x222 & x1142 ) | ( x222 & n1811 ) | ( x1142 & n1811 ) ;
  assign n2703 = n2701 & n2702 ;
  assign n2704 = n2700 & ~n2703 ;
  assign n2705 = ~n2695 & n2704 ;
  assign n2706 = n2227 & ~n2697 ;
  assign n2707 = n2704 & ~n2706 ;
  assign n2708 = x223 | n2707 ;
  assign n2709 = ~n2695 & n2708 ;
  assign n2710 = x39 | n2709 ;
  assign n2711 = n2705 | n2710 ;
  assign n2712 = n2693 | n2711 ;
  assign n2713 = ~x224 & n2678 ;
  assign n2714 = n2697 | n2713 ;
  assign n2715 = ~n2703 & n2714 ;
  assign n2716 = x223 | n2715 ;
  assign n2717 = ~n2694 & n2716 ;
  assign n2718 = x299 | n2717 ;
  assign n2719 = n2599 | n2718 ;
  assign n2720 = x262 | n1868 ;
  assign n2721 = x172 & ~x228 ;
  assign n2722 = n2082 & ~n2721 ;
  assign n2723 = n2720 & ~n2722 ;
  assign n2724 = n2679 | n2681 ;
  assign n2725 = x228 & n2724 ;
  assign n2726 = n2205 | n2725 ;
  assign n2727 = n2723 | n2726 ;
  assign n2728 = ~x216 & n2727 ;
  assign n2729 = n2669 | n2728 ;
  assign n2730 = ~n2690 & n2729 ;
  assign n2731 = x215 | n2730 ;
  assign n2732 = ~n2666 & n2731 ;
  assign n2733 = x299 & ~n2732 ;
  assign n2734 = n2719 & ~n2733 ;
  assign n2735 = x39 & ~n2734 ;
  assign n2736 = x38 | n2735 ;
  assign n2737 = n2712 & ~n2736 ;
  assign n2738 = n2721 | n2725 ;
  assign n2739 = ~x216 & n2738 ;
  assign n2740 = n2669 | n2739 ;
  assign n2741 = ~n2690 & n2740 ;
  assign n2742 = x215 | n2741 ;
  assign n2743 = ~n2666 & n2742 ;
  assign n2744 = n2206 | n2743 ;
  assign n2745 = x299 & ~n2744 ;
  assign n2746 = n2719 & ~n2745 ;
  assign n2747 = x38 & n2746 ;
  assign n2748 = x100 | n2747 ;
  assign n2749 = n2737 | n2748 ;
  assign n2750 = ~n1925 & n2719 ;
  assign n2751 = x262 | n2161 ;
  assign n2752 = n2354 & ~n2721 ;
  assign n2753 = n2751 & ~n2752 ;
  assign n2754 = n2726 | n2753 ;
  assign n2755 = ~x216 & n2754 ;
  assign n2756 = n2669 | n2755 ;
  assign n2757 = ~n2690 & n2756 ;
  assign n2758 = x215 | n2757 ;
  assign n2759 = n2667 & n2758 ;
  assign n2760 = ( ~x299 & n2750 ) | ( ~x299 & n2759 ) | ( n2750 & n2759 ) ;
  assign n2761 = ( x100 & n2364 ) | ( x100 & ~n2746 ) | ( n2364 & ~n2746 ) ;
  assign n2762 = ~n2760 & n2761 ;
  assign n2763 = n2749 & ~n2762 ;
  assign n2764 = x87 | n2763 ;
  assign n2765 = n1976 & n2746 ;
  assign n2766 = ~n1976 & n2734 ;
  assign n2767 = n2765 | n2766 ;
  assign n2768 = ( x75 & n1998 ) | ( x75 & ~n2767 ) | ( n1998 & ~n2767 ) ;
  assign n2769 = n2764 & ~n2768 ;
  assign n2770 = x75 & n2746 ;
  assign n2771 = x92 | n2770 ;
  assign n2772 = n2769 | n2771 ;
  assign n2773 = ( ~x92 & n1998 ) | ( ~x92 & n2746 ) | ( n1998 & n2746 ) ;
  assign n2774 = ( x92 & n1998 ) | ( x92 & ~n2767 ) | ( n1998 & ~n2767 ) ;
  assign n2775 = ~n2773 & n2774 ;
  assign n2776 = n2030 | n2775 ;
  assign n2777 = n2772 & ~n2776 ;
  assign n2778 = n2030 & n2746 ;
  assign n2779 = x55 | n2778 ;
  assign n2780 = n2777 | n2779 ;
  assign n2781 = ( ~x55 & n2033 ) | ( ~x55 & n2744 ) | ( n2033 & n2744 ) ;
  assign n2782 = ( x55 & n2033 ) | ( x55 & ~n2732 ) | ( n2033 & ~n2732 ) ;
  assign n2783 = ~n2781 & n2782 ;
  assign n2784 = x56 | n2783 ;
  assign n2785 = n2780 & ~n2784 ;
  assign n2786 = ( x56 & ~n2045 ) | ( x56 & n2744 ) | ( ~n2045 & n2744 ) ;
  assign n2787 = ( x56 & n2045 ) | ( x56 & n2732 ) | ( n2045 & n2732 ) ;
  assign n2788 = n2786 & n2787 ;
  assign n2789 = x62 | n2788 ;
  assign n2790 = n2785 | n2789 ;
  assign n2791 = ( ~x62 & n2193 ) | ( ~x62 & n2744 ) | ( n2193 & n2744 ) ;
  assign n2792 = ( x62 & n2193 ) | ( x62 & ~n2732 ) | ( n2193 & ~n2732 ) ;
  assign n2793 = ~n2791 & n2792 ;
  assign n2794 = n2057 | n2793 ;
  assign n2795 = n2790 & ~n2794 ;
  assign n2796 = n2057 & n2744 ;
  assign n2797 = x249 | n2796 ;
  assign n2798 = n2795 | n2797 ;
  assign n2799 = x172 | n2672 ;
  assign n2800 = ( x172 & ~x262 ) | ( x172 & n2230 ) | ( ~x262 & n2230 ) ;
  assign n2801 = ( x172 & x262 ) | ( x172 & n2138 ) | ( x262 & n2138 ) ;
  assign n2802 = n2800 & n2801 ;
  assign n2803 = n2799 & ~n2802 ;
  assign n2804 = x228 | n2803 ;
  assign n2805 = x216 | n2683 ;
  assign n2806 = n2804 & ~n2805 ;
  assign n2807 = n2669 | n2806 ;
  assign n2808 = ~n2690 & n2807 ;
  assign n2809 = x215 | n2808 ;
  assign n2810 = n2667 & n2809 ;
  assign n2811 = n2710 | n2810 ;
  assign n2812 = n2723 | n2725 ;
  assign n2813 = ~x216 & n2812 ;
  assign n2814 = n2669 | n2813 ;
  assign n2815 = ~n2690 & n2814 ;
  assign n2816 = x215 | n2815 ;
  assign n2817 = ~n2666 & n2816 ;
  assign n2818 = x299 & ~n2817 ;
  assign n2819 = n2718 & ~n2818 ;
  assign n2820 = x39 & ~n2819 ;
  assign n2821 = x38 | n2820 ;
  assign n2822 = n2811 & ~n2821 ;
  assign n2823 = x299 & ~n2743 ;
  assign n2824 = n2718 & ~n2823 ;
  assign n2825 = x38 & n2824 ;
  assign n2826 = x100 | n2825 ;
  assign n2827 = n2822 | n2826 ;
  assign n2828 = ~n1925 & n2718 ;
  assign n2829 = n2725 | n2753 ;
  assign n2830 = ~x216 & n2829 ;
  assign n2831 = n2669 | n2830 ;
  assign n2832 = ~n2690 & n2831 ;
  assign n2833 = x215 | n2832 ;
  assign n2834 = n2667 & n2833 ;
  assign n2835 = ( ~x299 & n2828 ) | ( ~x299 & n2834 ) | ( n2828 & n2834 ) ;
  assign n2836 = ( x100 & n2364 ) | ( x100 & ~n2824 ) | ( n2364 & ~n2824 ) ;
  assign n2837 = ~n2835 & n2836 ;
  assign n2838 = n2827 & ~n2837 ;
  assign n2839 = x87 | n2838 ;
  assign n2840 = n1976 & n2824 ;
  assign n2841 = ~n1976 & n2819 ;
  assign n2842 = n2840 | n2841 ;
  assign n2843 = ( x75 & n1998 ) | ( x75 & ~n2842 ) | ( n1998 & ~n2842 ) ;
  assign n2844 = n2839 & ~n2843 ;
  assign n2845 = x75 & n2824 ;
  assign n2846 = x92 | n2845 ;
  assign n2847 = n2844 | n2846 ;
  assign n2848 = ( ~x92 & n1998 ) | ( ~x92 & n2824 ) | ( n1998 & n2824 ) ;
  assign n2849 = ( x92 & n1998 ) | ( x92 & ~n2842 ) | ( n1998 & ~n2842 ) ;
  assign n2850 = ~n2848 & n2849 ;
  assign n2851 = n2030 | n2850 ;
  assign n2852 = n2847 & ~n2851 ;
  assign n2853 = n2030 & n2824 ;
  assign n2854 = x55 | n2853 ;
  assign n2855 = n2852 | n2854 ;
  assign n2856 = ( ~x55 & n2033 ) | ( ~x55 & n2743 ) | ( n2033 & n2743 ) ;
  assign n2857 = ( x55 & n2033 ) | ( x55 & ~n2817 ) | ( n2033 & ~n2817 ) ;
  assign n2858 = ~n2856 & n2857 ;
  assign n2859 = x56 | n2858 ;
  assign n2860 = n2855 & ~n2859 ;
  assign n2861 = ( x56 & ~n2045 ) | ( x56 & n2743 ) | ( ~n2045 & n2743 ) ;
  assign n2862 = ( x56 & n2045 ) | ( x56 & n2817 ) | ( n2045 & n2817 ) ;
  assign n2863 = n2861 & n2862 ;
  assign n2864 = x62 | n2863 ;
  assign n2865 = n2860 | n2864 ;
  assign n2866 = ( ~x62 & n2193 ) | ( ~x62 & n2743 ) | ( n2193 & n2743 ) ;
  assign n2867 = ( x62 & n2193 ) | ( x62 & ~n2817 ) | ( n2193 & ~n2817 ) ;
  assign n2868 = ~n2866 & n2867 ;
  assign n2869 = n2057 | n2868 ;
  assign n2870 = n2865 & ~n2869 ;
  assign n2871 = n2057 & n2743 ;
  assign n2872 = x249 & ~n2871 ;
  assign n2873 = ~n2870 & n2872 ;
  assign n2874 = n2798 & ~n2873 ;
  assign n2875 = x215 & x1141 ;
  assign n2876 = x299 & ~n2875 ;
  assign n2877 = x216 & x270 ;
  assign n2878 = x221 | n2877 ;
  assign n2879 = x861 & n2230 ;
  assign n2880 = x171 | n2879 ;
  assign n2881 = x171 & n2239 ;
  assign n2882 = n2880 & ~n2881 ;
  assign n2883 = n2138 | n2880 ;
  assign n2884 = ( ~x861 & n2882 ) | ( ~x861 & n2883 ) | ( n2882 & n2883 ) ;
  assign n2885 = x228 | n2884 ;
  assign n2886 = x861 & ~n1491 ;
  assign n2887 = ( ~x105 & x228 ) | ( ~x105 & n2886 ) | ( x228 & n2886 ) ;
  assign n2888 = ( x105 & ~x171 ) | ( x105 & x228 ) | ( ~x171 & x228 ) ;
  assign n2889 = n2887 & n2888 ;
  assign n2890 = ~n2228 & n2889 ;
  assign n2891 = x216 | n2890 ;
  assign n2892 = n2885 & ~n2891 ;
  assign n2893 = n2878 | n2892 ;
  assign n2894 = ( x221 & x935 ) | ( x221 & ~n1205 ) | ( x935 & ~n1205 ) ;
  assign n2895 = ( x221 & x1141 ) | ( x221 & n1205 ) | ( x1141 & n1205 ) ;
  assign n2896 = n2894 & n2895 ;
  assign n2897 = n2893 & ~n2896 ;
  assign n2898 = x215 | n2897 ;
  assign n2899 = n2876 & n2898 ;
  assign n2900 = x223 & x1141 ;
  assign n2901 = x299 | n2900 ;
  assign n2902 = x224 & x270 ;
  assign n2903 = x222 | n2902 ;
  assign n2904 = x861 & ~n2227 ;
  assign n2905 = x224 | n2904 ;
  assign n2906 = ~n2903 & n2905 ;
  assign n2907 = ( x222 & x935 ) | ( x222 & ~n1811 ) | ( x935 & ~n1811 ) ;
  assign n2908 = ( x222 & x1141 ) | ( x222 & n1811 ) | ( x1141 & n1811 ) ;
  assign n2909 = n2907 & n2908 ;
  assign n2910 = n2906 | n2909 ;
  assign n2911 = n2901 | n2910 ;
  assign n2912 = n2227 & ~n2903 ;
  assign n2913 = n2910 | n2912 ;
  assign n2914 = ~x223 & n2913 ;
  assign n2915 = n2901 | n2914 ;
  assign n2916 = ~x39 & n2915 ;
  assign n2917 = n2911 & n2916 ;
  assign n2918 = ~n2899 & n2917 ;
  assign n2919 = x224 | n2886 ;
  assign n2920 = ~n2903 & n2919 ;
  assign n2921 = n2909 | n2920 ;
  assign n2922 = ~x223 & n2921 ;
  assign n2923 = n2900 | n2922 ;
  assign n2924 = ~x299 & n2923 ;
  assign n2925 = x216 | n2889 ;
  assign n2926 = x171 & n1868 ;
  assign n2927 = x861 | n1868 ;
  assign n2928 = ~x228 & n2927 ;
  assign n2929 = ~n2926 & n2928 ;
  assign n2930 = n2925 | n2929 ;
  assign n2931 = ~n2878 & n2930 ;
  assign n2932 = n2896 | n2931 ;
  assign n2933 = ~x215 & n2932 ;
  assign n2934 = n2875 | n2933 ;
  assign n2935 = x299 & n2934 ;
  assign n2936 = n2924 | n2935 ;
  assign n2937 = x39 & n2936 ;
  assign n2938 = x38 | n2937 ;
  assign n2939 = n2918 | n2938 ;
  assign n2940 = x171 | x228 ;
  assign n2941 = ~n2925 & n2940 ;
  assign n2942 = n2878 | n2941 ;
  assign n2943 = ~n2896 & n2942 ;
  assign n2944 = x215 | n2943 ;
  assign n2945 = ~n2875 & n2944 ;
  assign n2946 = x299 & ~n2945 ;
  assign n2947 = n2924 | n2946 ;
  assign n2948 = x38 & ~n2947 ;
  assign n2949 = x100 | n2948 ;
  assign n2950 = n2939 & ~n2949 ;
  assign n2951 = n1925 | n2924 ;
  assign n2952 = ( x171 & x228 ) | ( x171 & n2161 ) | ( x228 & n2161 ) ;
  assign n2953 = ( ~x228 & x861 ) | ( ~x228 & n2161 ) | ( x861 & n2161 ) ;
  assign n2954 = ~n2952 & n2953 ;
  assign n2955 = n2925 | n2954 ;
  assign n2956 = ~n2878 & n2955 ;
  assign n2957 = n2896 | n2956 ;
  assign n2958 = ~x215 & n2957 ;
  assign n2959 = n2876 & ~n2958 ;
  assign n2960 = ( x299 & n2951 ) | ( x299 & ~n2959 ) | ( n2951 & ~n2959 ) ;
  assign n2961 = ( x100 & n2364 ) | ( x100 & n2947 ) | ( n2364 & n2947 ) ;
  assign n2962 = n2960 & n2961 ;
  assign n2963 = n2950 | n2962 ;
  assign n2964 = ~x87 & n2963 ;
  assign n2965 = n1976 & ~n2947 ;
  assign n2966 = n1976 | n2936 ;
  assign n2967 = ~n2965 & n2966 ;
  assign n2968 = ( x75 & n1998 ) | ( x75 & n2967 ) | ( n1998 & n2967 ) ;
  assign n2969 = n2964 | n2968 ;
  assign n2970 = x75 & ~n2947 ;
  assign n2971 = x92 | n2970 ;
  assign n2972 = n2969 & ~n2971 ;
  assign n2973 = ( x92 & ~n1998 ) | ( x92 & n2947 ) | ( ~n1998 & n2947 ) ;
  assign n2974 = ( x92 & n1998 ) | ( x92 & n2967 ) | ( n1998 & n2967 ) ;
  assign n2975 = n2973 & n2974 ;
  assign n2976 = n2030 | n2975 ;
  assign n2977 = n2972 | n2976 ;
  assign n2978 = n2030 & ~n2947 ;
  assign n2979 = x55 | n2978 ;
  assign n2980 = n2977 & ~n2979 ;
  assign n2981 = ( x55 & n2033 ) | ( x55 & n2934 ) | ( n2033 & n2934 ) ;
  assign n2982 = ( ~x55 & n2033 ) | ( ~x55 & n2945 ) | ( n2033 & n2945 ) ;
  assign n2983 = n2981 & ~n2982 ;
  assign n2984 = x56 | n2983 ;
  assign n2985 = n2980 | n2984 ;
  assign n2986 = ( x56 & n2045 ) | ( x56 & ~n2934 ) | ( n2045 & ~n2934 ) ;
  assign n2987 = ( x56 & ~n2045 ) | ( x56 & n2945 ) | ( ~n2045 & n2945 ) ;
  assign n2988 = n2986 & n2987 ;
  assign n2989 = x62 | n2988 ;
  assign n2990 = n2985 & ~n2989 ;
  assign n2991 = x241 | n2057 ;
  assign n2992 = ( x62 & n2193 ) | ( x62 & n2934 ) | ( n2193 & n2934 ) ;
  assign n2993 = ( ~x62 & n2193 ) | ( ~x62 & n2945 ) | ( n2193 & n2945 ) ;
  assign n2994 = n2992 & ~n2993 ;
  assign n2995 = n2991 | n2994 ;
  assign n2996 = n2990 | n2995 ;
  assign n2997 = ~x861 & n2239 ;
  assign n2998 = x171 | n2997 ;
  assign n2999 = ( x171 & ~x861 ) | ( x171 & n2138 ) | ( ~x861 & n2138 ) ;
  assign n3000 = ( x171 & x861 ) | ( x171 & n2230 ) | ( x861 & n2230 ) ;
  assign n3001 = n2999 & n3000 ;
  assign n3002 = n2998 & ~n3001 ;
  assign n3003 = x228 | n3002 ;
  assign n3004 = n2588 | n2925 ;
  assign n3005 = n3003 & ~n3004 ;
  assign n3006 = n2878 | n3005 ;
  assign n3007 = ~n2896 & n3006 ;
  assign n3008 = x215 | n3007 ;
  assign n3009 = n2876 & n3008 ;
  assign n3010 = n2916 & ~n3009 ;
  assign n3011 = n2215 | n2924 ;
  assign n3012 = n2205 | n2925 ;
  assign n3013 = n2929 | n3012 ;
  assign n3014 = ~n2878 & n3013 ;
  assign n3015 = n2896 | n3014 ;
  assign n3016 = ~x215 & n3015 ;
  assign n3017 = n2875 | n3016 ;
  assign n3018 = x299 & n3017 ;
  assign n3019 = n3011 | n3018 ;
  assign n3020 = x39 & n3019 ;
  assign n3021 = x38 | n3020 ;
  assign n3022 = n3010 | n3021 ;
  assign n3023 = n2345 & ~n2877 ;
  assign n3024 = n2945 & ~n3023 ;
  assign n3025 = x299 & ~n3024 ;
  assign n3026 = n3011 | n3025 ;
  assign n3027 = x38 & ~n3026 ;
  assign n3028 = x100 | n3027 ;
  assign n3029 = n3022 & ~n3028 ;
  assign n3030 = n1925 | n3011 ;
  assign n3031 = n2954 | n3012 ;
  assign n3032 = ~n2878 & n3031 ;
  assign n3033 = n2896 | n3032 ;
  assign n3034 = ~x215 & n3033 ;
  assign n3035 = n2876 & ~n3034 ;
  assign n3036 = ( x299 & n3030 ) | ( x299 & ~n3035 ) | ( n3030 & ~n3035 ) ;
  assign n3037 = ( x100 & n2364 ) | ( x100 & n3026 ) | ( n2364 & n3026 ) ;
  assign n3038 = n3036 & n3037 ;
  assign n3039 = n3029 | n3038 ;
  assign n3040 = ~x87 & n3039 ;
  assign n3041 = n1976 & ~n3026 ;
  assign n3042 = n1976 | n3019 ;
  assign n3043 = ~n3041 & n3042 ;
  assign n3044 = ( x75 & n1998 ) | ( x75 & n3043 ) | ( n1998 & n3043 ) ;
  assign n3045 = n3040 | n3044 ;
  assign n3046 = x75 & ~n3026 ;
  assign n3047 = x92 | n3046 ;
  assign n3048 = n3045 & ~n3047 ;
  assign n3049 = ( x92 & ~n1998 ) | ( x92 & n3026 ) | ( ~n1998 & n3026 ) ;
  assign n3050 = ( x92 & n1998 ) | ( x92 & n3043 ) | ( n1998 & n3043 ) ;
  assign n3051 = n3049 & n3050 ;
  assign n3052 = n2030 | n3051 ;
  assign n3053 = n3048 | n3052 ;
  assign n3054 = n2030 & ~n3026 ;
  assign n3055 = x55 | n3054 ;
  assign n3056 = n3053 & ~n3055 ;
  assign n3057 = ( x55 & n2033 ) | ( x55 & n3017 ) | ( n2033 & n3017 ) ;
  assign n3058 = ( ~x55 & n2033 ) | ( ~x55 & n3024 ) | ( n2033 & n3024 ) ;
  assign n3059 = n3057 & ~n3058 ;
  assign n3060 = x56 | n3059 ;
  assign n3061 = n3056 | n3060 ;
  assign n3062 = ( x56 & n2045 ) | ( x56 & ~n3017 ) | ( n2045 & ~n3017 ) ;
  assign n3063 = ( x56 & ~n2045 ) | ( x56 & n3024 ) | ( ~n2045 & n3024 ) ;
  assign n3064 = n3062 & n3063 ;
  assign n3065 = x62 | n3064 ;
  assign n3066 = n3061 & ~n3065 ;
  assign n3067 = x241 & ~n2057 ;
  assign n3068 = ( x62 & n2193 ) | ( x62 & n3017 ) | ( n2193 & n3017 ) ;
  assign n3069 = ( ~x62 & n2193 ) | ( ~x62 & n3024 ) | ( n2193 & n3024 ) ;
  assign n3070 = n3068 & ~n3069 ;
  assign n3071 = n3067 & ~n3070 ;
  assign n3072 = ~n3066 & n3071 ;
  assign n3073 = x241 & n3023 ;
  assign n3074 = n2057 & ~n3073 ;
  assign n3075 = n2945 & n3074 ;
  assign n3076 = n3072 | n3075 ;
  assign n3077 = n2996 & ~n3076 ;
  assign n3078 = x215 & x1140 ;
  assign n3079 = x299 & ~n3078 ;
  assign n3080 = x216 & x282 ;
  assign n3081 = x221 | n3080 ;
  assign n3082 = x869 & n2230 ;
  assign n3083 = x170 | n3082 ;
  assign n3084 = x170 & n2239 ;
  assign n3085 = n3083 & ~n3084 ;
  assign n3086 = n2138 | n3083 ;
  assign n3087 = ( ~x869 & n3085 ) | ( ~x869 & n3086 ) | ( n3085 & n3086 ) ;
  assign n3088 = x228 | n3087 ;
  assign n3089 = x869 & ~n1491 ;
  assign n3090 = ( ~x105 & x228 ) | ( ~x105 & n3089 ) | ( x228 & n3089 ) ;
  assign n3091 = ( x105 & ~x170 ) | ( x105 & x228 ) | ( ~x170 & x228 ) ;
  assign n3092 = n3090 & n3091 ;
  assign n3093 = ~n2228 & n3092 ;
  assign n3094 = x216 | n3093 ;
  assign n3095 = n3088 & ~n3094 ;
  assign n3096 = n3081 | n3095 ;
  assign n3097 = ( x221 & x921 ) | ( x221 & ~n1205 ) | ( x921 & ~n1205 ) ;
  assign n3098 = ( x221 & x1140 ) | ( x221 & n1205 ) | ( x1140 & n1205 ) ;
  assign n3099 = n3097 & n3098 ;
  assign n3100 = n3096 & ~n3099 ;
  assign n3101 = x215 | n3100 ;
  assign n3102 = n3079 & n3101 ;
  assign n3103 = x223 & x1140 ;
  assign n3104 = x299 | n3103 ;
  assign n3105 = x224 & x282 ;
  assign n3106 = x222 | n3105 ;
  assign n3107 = x869 & ~n2227 ;
  assign n3108 = x224 | n3107 ;
  assign n3109 = ~n3106 & n3108 ;
  assign n3110 = ( x222 & x921 ) | ( x222 & ~n1811 ) | ( x921 & ~n1811 ) ;
  assign n3111 = ( x222 & x1140 ) | ( x222 & n1811 ) | ( x1140 & n1811 ) ;
  assign n3112 = n3110 & n3111 ;
  assign n3113 = n3109 | n3112 ;
  assign n3114 = n3104 | n3113 ;
  assign n3115 = n2227 & ~n3106 ;
  assign n3116 = n3113 | n3115 ;
  assign n3117 = ~x223 & n3116 ;
  assign n3118 = n3104 | n3117 ;
  assign n3119 = ~x39 & n3118 ;
  assign n3120 = n3114 & n3119 ;
  assign n3121 = ~n3102 & n3120 ;
  assign n3122 = x224 | n3089 ;
  assign n3123 = ~n3106 & n3122 ;
  assign n3124 = n3112 | n3123 ;
  assign n3125 = ~x223 & n3124 ;
  assign n3126 = n3103 | n3125 ;
  assign n3127 = ~x299 & n3126 ;
  assign n3128 = x216 | n3092 ;
  assign n3129 = x170 & n1868 ;
  assign n3130 = x869 | n1868 ;
  assign n3131 = ~x228 & n3130 ;
  assign n3132 = ~n3129 & n3131 ;
  assign n3133 = n3128 | n3132 ;
  assign n3134 = ~n3081 & n3133 ;
  assign n3135 = n3099 | n3134 ;
  assign n3136 = ~x215 & n3135 ;
  assign n3137 = n3078 | n3136 ;
  assign n3138 = x299 & n3137 ;
  assign n3139 = n3127 | n3138 ;
  assign n3140 = x39 & n3139 ;
  assign n3141 = x38 | n3140 ;
  assign n3142 = n3121 | n3141 ;
  assign n3143 = x170 | x228 ;
  assign n3144 = ~n3128 & n3143 ;
  assign n3145 = n3081 | n3144 ;
  assign n3146 = ~n3099 & n3145 ;
  assign n3147 = x215 | n3146 ;
  assign n3148 = ~n3078 & n3147 ;
  assign n3149 = x299 & ~n3148 ;
  assign n3150 = n3127 | n3149 ;
  assign n3151 = x38 & ~n3150 ;
  assign n3152 = x100 | n3151 ;
  assign n3153 = n3142 & ~n3152 ;
  assign n3154 = n1925 | n3127 ;
  assign n3155 = ( x170 & x228 ) | ( x170 & n2161 ) | ( x228 & n2161 ) ;
  assign n3156 = ( ~x228 & x869 ) | ( ~x228 & n2161 ) | ( x869 & n2161 ) ;
  assign n3157 = ~n3155 & n3156 ;
  assign n3158 = n3128 | n3157 ;
  assign n3159 = ~n3081 & n3158 ;
  assign n3160 = n3099 | n3159 ;
  assign n3161 = ~x215 & n3160 ;
  assign n3162 = n3079 & ~n3161 ;
  assign n3163 = ( x299 & n3154 ) | ( x299 & ~n3162 ) | ( n3154 & ~n3162 ) ;
  assign n3164 = ( x100 & n2364 ) | ( x100 & n3150 ) | ( n2364 & n3150 ) ;
  assign n3165 = n3163 & n3164 ;
  assign n3166 = n3153 | n3165 ;
  assign n3167 = ~x87 & n3166 ;
  assign n3168 = n1976 & ~n3150 ;
  assign n3169 = n1976 | n3139 ;
  assign n3170 = ~n3168 & n3169 ;
  assign n3171 = ( x75 & n1998 ) | ( x75 & n3170 ) | ( n1998 & n3170 ) ;
  assign n3172 = n3167 | n3171 ;
  assign n3173 = x75 & ~n3150 ;
  assign n3174 = x92 | n3173 ;
  assign n3175 = n3172 & ~n3174 ;
  assign n3176 = ( x92 & ~n1998 ) | ( x92 & n3150 ) | ( ~n1998 & n3150 ) ;
  assign n3177 = ( x92 & n1998 ) | ( x92 & n3170 ) | ( n1998 & n3170 ) ;
  assign n3178 = n3176 & n3177 ;
  assign n3179 = n2030 | n3178 ;
  assign n3180 = n3175 | n3179 ;
  assign n3181 = n2030 & ~n3150 ;
  assign n3182 = x55 | n3181 ;
  assign n3183 = n3180 & ~n3182 ;
  assign n3184 = ( x55 & n2033 ) | ( x55 & n3137 ) | ( n2033 & n3137 ) ;
  assign n3185 = ( ~x55 & n2033 ) | ( ~x55 & n3148 ) | ( n2033 & n3148 ) ;
  assign n3186 = n3184 & ~n3185 ;
  assign n3187 = x56 | n3186 ;
  assign n3188 = n3183 | n3187 ;
  assign n3189 = ( x56 & n2045 ) | ( x56 & ~n3137 ) | ( n2045 & ~n3137 ) ;
  assign n3190 = ( x56 & ~n2045 ) | ( x56 & n3148 ) | ( ~n2045 & n3148 ) ;
  assign n3191 = n3189 & n3190 ;
  assign n3192 = x62 | n3191 ;
  assign n3193 = n3188 & ~n3192 ;
  assign n3194 = x248 | n2057 ;
  assign n3195 = ( x62 & n2193 ) | ( x62 & n3137 ) | ( n2193 & n3137 ) ;
  assign n3196 = ( ~x62 & n2193 ) | ( ~x62 & n3148 ) | ( n2193 & n3148 ) ;
  assign n3197 = n3195 & ~n3196 ;
  assign n3198 = n3194 | n3197 ;
  assign n3199 = n3193 | n3198 ;
  assign n3200 = ~x869 & n2239 ;
  assign n3201 = x170 | n3200 ;
  assign n3202 = ( x170 & ~x869 ) | ( x170 & n2138 ) | ( ~x869 & n2138 ) ;
  assign n3203 = ( x170 & x869 ) | ( x170 & n2230 ) | ( x869 & n2230 ) ;
  assign n3204 = n3202 & n3203 ;
  assign n3205 = n3201 & ~n3204 ;
  assign n3206 = x228 | n3205 ;
  assign n3207 = n2588 | n3128 ;
  assign n3208 = n3206 & ~n3207 ;
  assign n3209 = n3081 | n3208 ;
  assign n3210 = ~n3099 & n3209 ;
  assign n3211 = x215 | n3210 ;
  assign n3212 = n3079 & n3211 ;
  assign n3213 = n3119 & ~n3212 ;
  assign n3214 = n2215 | n3127 ;
  assign n3215 = n2205 | n3128 ;
  assign n3216 = n3132 | n3215 ;
  assign n3217 = ~n3081 & n3216 ;
  assign n3218 = n3099 | n3217 ;
  assign n3219 = ~x215 & n3218 ;
  assign n3220 = n3078 | n3219 ;
  assign n3221 = x299 & n3220 ;
  assign n3222 = n3214 | n3221 ;
  assign n3223 = x39 & n3222 ;
  assign n3224 = x38 | n3223 ;
  assign n3225 = n3213 | n3224 ;
  assign n3226 = n2345 & ~n3080 ;
  assign n3227 = n3148 & ~n3226 ;
  assign n3228 = x299 & ~n3227 ;
  assign n3229 = n3214 | n3228 ;
  assign n3230 = x38 & ~n3229 ;
  assign n3231 = x100 | n3230 ;
  assign n3232 = n3225 & ~n3231 ;
  assign n3233 = n1925 | n3214 ;
  assign n3234 = n3157 | n3215 ;
  assign n3235 = ~n3081 & n3234 ;
  assign n3236 = n3099 | n3235 ;
  assign n3237 = ~x215 & n3236 ;
  assign n3238 = n3079 & ~n3237 ;
  assign n3239 = ( x299 & n3233 ) | ( x299 & ~n3238 ) | ( n3233 & ~n3238 ) ;
  assign n3240 = ( x100 & n2364 ) | ( x100 & n3229 ) | ( n2364 & n3229 ) ;
  assign n3241 = n3239 & n3240 ;
  assign n3242 = n3232 | n3241 ;
  assign n3243 = ~x87 & n3242 ;
  assign n3244 = n1976 & ~n3229 ;
  assign n3245 = n1976 | n3222 ;
  assign n3246 = ~n3244 & n3245 ;
  assign n3247 = ( x75 & n1998 ) | ( x75 & n3246 ) | ( n1998 & n3246 ) ;
  assign n3248 = n3243 | n3247 ;
  assign n3249 = x75 & ~n3229 ;
  assign n3250 = x92 | n3249 ;
  assign n3251 = n3248 & ~n3250 ;
  assign n3252 = ( x92 & ~n1998 ) | ( x92 & n3229 ) | ( ~n1998 & n3229 ) ;
  assign n3253 = ( x92 & n1998 ) | ( x92 & n3246 ) | ( n1998 & n3246 ) ;
  assign n3254 = n3252 & n3253 ;
  assign n3255 = n2030 | n3254 ;
  assign n3256 = n3251 | n3255 ;
  assign n3257 = n2030 & ~n3229 ;
  assign n3258 = x55 | n3257 ;
  assign n3259 = n3256 & ~n3258 ;
  assign n3260 = ( x55 & n2033 ) | ( x55 & n3220 ) | ( n2033 & n3220 ) ;
  assign n3261 = ( ~x55 & n2033 ) | ( ~x55 & n3227 ) | ( n2033 & n3227 ) ;
  assign n3262 = n3260 & ~n3261 ;
  assign n3263 = x56 | n3262 ;
  assign n3264 = n3259 | n3263 ;
  assign n3265 = ( x56 & n2045 ) | ( x56 & ~n3220 ) | ( n2045 & ~n3220 ) ;
  assign n3266 = ( x56 & ~n2045 ) | ( x56 & n3227 ) | ( ~n2045 & n3227 ) ;
  assign n3267 = n3265 & n3266 ;
  assign n3268 = x62 | n3267 ;
  assign n3269 = n3264 & ~n3268 ;
  assign n3270 = x248 & ~n2057 ;
  assign n3271 = ( x62 & n2193 ) | ( x62 & n3220 ) | ( n2193 & n3220 ) ;
  assign n3272 = ( ~x62 & n2193 ) | ( ~x62 & n3227 ) | ( n2193 & n3227 ) ;
  assign n3273 = n3271 & ~n3272 ;
  assign n3274 = n3270 & ~n3273 ;
  assign n3275 = ~n3269 & n3274 ;
  assign n3276 = x248 & n3226 ;
  assign n3277 = n2057 & ~n3276 ;
  assign n3278 = n3148 & n3277 ;
  assign n3279 = n3275 | n3278 ;
  assign n3280 = n3199 & ~n3279 ;
  assign n3281 = x216 & ~x1139 ;
  assign n3282 = ( x216 & x833 ) | ( x216 & x920 ) | ( x833 & x920 ) ;
  assign n3283 = ( x216 & ~x833 ) | ( x216 & x1139 ) | ( ~x833 & x1139 ) ;
  assign n3284 = n3282 | n3283 ;
  assign n3285 = x221 & n3284 ;
  assign n3286 = ~n3281 & n3285 ;
  assign n3287 = x216 & x281 ;
  assign n3288 = x221 | n3287 ;
  assign n3289 = x216 | x862 ;
  assign n3290 = n2082 & ~n2355 ;
  assign n3291 = n3289 | n3290 ;
  assign n3292 = ~n3288 & n3291 ;
  assign n3293 = n3286 | n3292 ;
  assign n3294 = n2356 & ~n3288 ;
  assign n3295 = n3293 | n3294 ;
  assign n3296 = x148 & ~x215 ;
  assign n3297 = x216 | n3285 ;
  assign n3298 = n2356 & ~n3297 ;
  assign n3299 = n3296 & ~n3298 ;
  assign n3300 = n3295 & n3299 ;
  assign n3301 = x215 & x1139 ;
  assign n3302 = x148 | x215 ;
  assign n3303 = ~n1898 & n2082 ;
  assign n3304 = x862 & ~n2205 ;
  assign n3305 = x216 | n3304 ;
  assign n3306 = n3303 | n3305 ;
  assign n3307 = ~n3288 & n3306 ;
  assign n3308 = n3286 | n3307 ;
  assign n3309 = ~n1898 & n2354 ;
  assign n3310 = ~n3288 & n3309 ;
  assign n3311 = n3308 | n3310 ;
  assign n3312 = ~n3302 & n3311 ;
  assign n3313 = n3301 | n3312 ;
  assign n3314 = n3300 | n3313 ;
  assign n3315 = x299 & n3314 ;
  assign n3316 = x223 & x1139 ;
  assign n3317 = x224 | n3316 ;
  assign n3318 = ( x222 & x920 ) | ( x222 & ~n1811 ) | ( x920 & ~n1811 ) ;
  assign n3319 = ( x222 & x1139 ) | ( x222 & n1811 ) | ( x1139 & n1811 ) ;
  assign n3320 = n3318 & n3319 ;
  assign n3321 = n3317 | n3320 ;
  assign n3322 = n1491 & ~n3321 ;
  assign n3323 = x862 | n3321 ;
  assign n3324 = x281 & n1817 ;
  assign n3325 = ( x222 & ~n3320 ) | ( x222 & n3324 ) | ( ~n3320 & n3324 ) ;
  assign n3326 = x223 | n3325 ;
  assign n3327 = ~n3316 & n3326 ;
  assign n3328 = x299 | n3327 ;
  assign n3329 = n3323 & ~n3328 ;
  assign n3330 = ~n3322 & n3329 ;
  assign n3331 = n1925 | n3330 ;
  assign n3332 = n3315 | n3331 ;
  assign n3333 = n2355 & ~n3289 ;
  assign n3334 = n3288 | n3333 ;
  assign n3335 = ~n3286 & n3334 ;
  assign n3336 = x148 & ~n1898 ;
  assign n3337 = ~n3297 & n3336 ;
  assign n3338 = x215 | n3337 ;
  assign n3339 = n3335 | n3338 ;
  assign n3340 = ~n3301 & n3339 ;
  assign n3341 = n2206 | n3340 ;
  assign n3342 = x299 & ~n3341 ;
  assign n3343 = n3330 | n3342 ;
  assign n3344 = ( x100 & n2364 ) | ( x100 & n3343 ) | ( n2364 & n3343 ) ;
  assign n3345 = n3332 & n3344 ;
  assign n3346 = ( x216 & x862 ) | ( x216 & ~n2232 ) | ( x862 & ~n2232 ) ;
  assign n3347 = ~x228 & n2138 ;
  assign n3348 = n1898 | n3347 ;
  assign n3349 = ( ~x216 & x862 ) | ( ~x216 & n3348 ) | ( x862 & n3348 ) ;
  assign n3350 = ~n3346 & n3349 ;
  assign n3351 = n3288 | n3350 ;
  assign n3352 = ~n3286 & n3351 ;
  assign n3353 = n3302 | n3352 ;
  assign n3354 = n2242 & ~n3289 ;
  assign n3355 = n3288 | n3354 ;
  assign n3356 = ~n3286 & n3355 ;
  assign n3357 = n2242 | n3297 ;
  assign n3358 = n3296 & n3357 ;
  assign n3359 = ~n3356 & n3358 ;
  assign n3360 = x299 & ~n3301 ;
  assign n3361 = ~n3359 & n3360 ;
  assign n3362 = n3353 & n3361 ;
  assign n3363 = n2227 & ~n3321 ;
  assign n3364 = n3323 & ~n3327 ;
  assign n3365 = ~n3363 & n3364 ;
  assign n3366 = x299 | n3365 ;
  assign n3367 = ~x39 & n3366 ;
  assign n3368 = ~n3362 & n3367 ;
  assign n3369 = ~n3302 & n3308 ;
  assign n3370 = n3293 & n3296 ;
  assign n3371 = ( ~n3290 & n3297 ) | ( ~n3290 & n3370 ) | ( n3297 & n3370 ) ;
  assign n3372 = n3370 & n3371 ;
  assign n3373 = n3301 | n3372 ;
  assign n3374 = n3369 | n3373 ;
  assign n3375 = x299 & n3374 ;
  assign n3376 = n3330 | n3375 ;
  assign n3377 = x39 & n3376 ;
  assign n3378 = x38 | n3377 ;
  assign n3379 = n3368 | n3378 ;
  assign n3380 = x38 & ~n3343 ;
  assign n3381 = x100 | n3380 ;
  assign n3382 = n3379 & ~n3381 ;
  assign n3383 = n3345 | n3382 ;
  assign n3384 = ~x87 & n3383 ;
  assign n3385 = n1976 & ~n3343 ;
  assign n3386 = n1976 | n3376 ;
  assign n3387 = ~n3385 & n3386 ;
  assign n3388 = ( x75 & n1998 ) | ( x75 & n3387 ) | ( n1998 & n3387 ) ;
  assign n3389 = n3384 | n3388 ;
  assign n3390 = x75 & ~n3343 ;
  assign n3391 = x92 | n3390 ;
  assign n3392 = n3389 & ~n3391 ;
  assign n3393 = ( x92 & ~n1998 ) | ( x92 & n3343 ) | ( ~n1998 & n3343 ) ;
  assign n3394 = ( x92 & n1998 ) | ( x92 & n3387 ) | ( n1998 & n3387 ) ;
  assign n3395 = n3393 & n3394 ;
  assign n3396 = n2030 | n3395 ;
  assign n3397 = n3392 | n3396 ;
  assign n3398 = n2030 & ~n3343 ;
  assign n3399 = x55 | n3398 ;
  assign n3400 = n3397 & ~n3399 ;
  assign n3401 = ( x55 & n2033 ) | ( x55 & n3374 ) | ( n2033 & n3374 ) ;
  assign n3402 = ( ~x55 & n2033 ) | ( ~x55 & n3341 ) | ( n2033 & n3341 ) ;
  assign n3403 = n3401 & ~n3402 ;
  assign n3404 = x56 | n3403 ;
  assign n3405 = n3400 | n3404 ;
  assign n3406 = ( x56 & n2045 ) | ( x56 & ~n3374 ) | ( n2045 & ~n3374 ) ;
  assign n3407 = ( x56 & ~n2045 ) | ( x56 & n3341 ) | ( ~n2045 & n3341 ) ;
  assign n3408 = n3406 & n3407 ;
  assign n3409 = x62 | n3408 ;
  assign n3410 = n3405 & ~n3409 ;
  assign n3411 = ( x62 & n2193 ) | ( x62 & n3374 ) | ( n2193 & n3374 ) ;
  assign n3412 = ( ~x62 & n2193 ) | ( ~x62 & n3341 ) | ( n2193 & n3341 ) ;
  assign n3413 = n3411 & ~n3412 ;
  assign n3414 = n2057 | n3413 ;
  assign n3415 = n3410 | n3414 ;
  assign n3416 = n2057 & n3341 ;
  assign n3417 = x247 | n3416 ;
  assign n3418 = n3415 & ~n3417 ;
  assign n3419 = n3295 & ~n3302 ;
  assign n3420 = ~n3309 & n3370 ;
  assign n3421 = ( n3297 & n3370 ) | ( n3297 & n3420 ) | ( n3370 & n3420 ) ;
  assign n3422 = n3301 | n3421 ;
  assign n3423 = n3419 | n3422 ;
  assign n3424 = x299 & n3423 ;
  assign n3425 = n2215 | n3329 ;
  assign n3426 = n1925 | n3425 ;
  assign n3427 = n3424 | n3426 ;
  assign n3428 = x299 & ~n3340 ;
  assign n3429 = n3425 | n3428 ;
  assign n3430 = ( x100 & n2364 ) | ( x100 & n3429 ) | ( n2364 & n3429 ) ;
  assign n3431 = n3427 & n3430 ;
  assign n3432 = x38 & ~n3429 ;
  assign n3433 = x100 | n3432 ;
  assign n3434 = n3293 & ~n3338 ;
  assign n3435 = n3373 | n3434 ;
  assign n3436 = x299 & n3435 ;
  assign n3437 = n3425 | n3436 ;
  assign n3438 = ( x38 & x39 ) | ( x38 & n3437 ) | ( x39 & n3437 ) ;
  assign n3439 = ( x216 & x862 ) | ( x216 & n3348 ) | ( x862 & n3348 ) ;
  assign n3440 = ( x216 & ~x862 ) | ( x216 & n2232 ) | ( ~x862 & n2232 ) ;
  assign n3441 = n3439 | n3440 ;
  assign n3442 = ~n3288 & n3441 ;
  assign n3443 = n3286 | n3442 ;
  assign n3444 = n3296 & n3443 ;
  assign n3445 = n3302 | n3356 ;
  assign n3446 = ~n3301 & n3445 ;
  assign n3447 = ~n3444 & n3446 ;
  assign n3448 = x299 & ~n3447 ;
  assign n3449 = ( n2227 & ~n3328 ) | ( n2227 & n3329 ) | ( ~n3328 & n3329 ) ;
  assign n3450 = n3448 | n3449 ;
  assign n3451 = ( x38 & ~x39 ) | ( x38 & n3450 ) | ( ~x39 & n3450 ) ;
  assign n3452 = n3438 | n3451 ;
  assign n3453 = ~n3433 & n3452 ;
  assign n3454 = n3431 | n3453 ;
  assign n3455 = ~x87 & n3454 ;
  assign n3456 = n1976 & ~n3429 ;
  assign n3457 = n1976 | n3437 ;
  assign n3458 = ~n3456 & n3457 ;
  assign n3459 = ( x75 & n1998 ) | ( x75 & n3458 ) | ( n1998 & n3458 ) ;
  assign n3460 = n3455 | n3459 ;
  assign n3461 = x75 & ~n3429 ;
  assign n3462 = x92 | n3461 ;
  assign n3463 = n3460 & ~n3462 ;
  assign n3464 = ( x92 & ~n1998 ) | ( x92 & n3429 ) | ( ~n1998 & n3429 ) ;
  assign n3465 = ( x92 & n1998 ) | ( x92 & n3458 ) | ( n1998 & n3458 ) ;
  assign n3466 = n3464 & n3465 ;
  assign n3467 = n2030 | n3466 ;
  assign n3468 = n3463 | n3467 ;
  assign n3469 = n2030 & ~n3429 ;
  assign n3470 = x55 | n3469 ;
  assign n3471 = n3468 & ~n3470 ;
  assign n3472 = ( x55 & n2033 ) | ( x55 & n3435 ) | ( n2033 & n3435 ) ;
  assign n3473 = ( ~x55 & n2033 ) | ( ~x55 & n3340 ) | ( n2033 & n3340 ) ;
  assign n3474 = n3472 & ~n3473 ;
  assign n3475 = x56 | n3474 ;
  assign n3476 = n3471 | n3475 ;
  assign n3477 = ( x56 & n2045 ) | ( x56 & ~n3435 ) | ( n2045 & ~n3435 ) ;
  assign n3478 = ( x56 & ~n2045 ) | ( x56 & n3340 ) | ( ~n2045 & n3340 ) ;
  assign n3479 = n3477 & n3478 ;
  assign n3480 = x62 | n3479 ;
  assign n3481 = n3476 & ~n3480 ;
  assign n3482 = ( x62 & n2193 ) | ( x62 & n3435 ) | ( n2193 & n3435 ) ;
  assign n3483 = ( ~x62 & n2193 ) | ( ~x62 & n3340 ) | ( n2193 & n3340 ) ;
  assign n3484 = n3482 & ~n3483 ;
  assign n3485 = n2057 | n3484 ;
  assign n3486 = n3481 | n3485 ;
  assign n3487 = n2057 & n3340 ;
  assign n3488 = x247 & ~n3487 ;
  assign n3489 = n3486 & n3488 ;
  assign n3490 = n3418 | n3489 ;
  assign n3491 = x215 & x1138 ;
  assign n3492 = x299 & ~n3491 ;
  assign n3493 = x216 & x269 ;
  assign n3494 = x221 | n3493 ;
  assign n3495 = x877 & n2230 ;
  assign n3496 = x169 | n3495 ;
  assign n3497 = x169 & n2239 ;
  assign n3498 = n3496 & ~n3497 ;
  assign n3499 = n2138 | n3496 ;
  assign n3500 = ( ~x877 & n3498 ) | ( ~x877 & n3499 ) | ( n3498 & n3499 ) ;
  assign n3501 = x228 | n3500 ;
  assign n3502 = x877 & ~n1491 ;
  assign n3503 = ( ~x105 & x228 ) | ( ~x105 & n3502 ) | ( x228 & n3502 ) ;
  assign n3504 = ( x105 & ~x169 ) | ( x105 & x228 ) | ( ~x169 & x228 ) ;
  assign n3505 = n3503 & n3504 ;
  assign n3506 = ~n2228 & n3505 ;
  assign n3507 = x216 | n3506 ;
  assign n3508 = n3501 & ~n3507 ;
  assign n3509 = n3494 | n3508 ;
  assign n3510 = ( x221 & x940 ) | ( x221 & ~n1205 ) | ( x940 & ~n1205 ) ;
  assign n3511 = ( x221 & x1138 ) | ( x221 & n1205 ) | ( x1138 & n1205 ) ;
  assign n3512 = n3510 & n3511 ;
  assign n3513 = n3509 & ~n3512 ;
  assign n3514 = x215 | n3513 ;
  assign n3515 = n3492 & n3514 ;
  assign n3516 = x223 & x1138 ;
  assign n3517 = x299 | n3516 ;
  assign n3518 = x224 & x269 ;
  assign n3519 = x222 | n3518 ;
  assign n3520 = x877 & ~n2227 ;
  assign n3521 = x224 | n3520 ;
  assign n3522 = ~n3519 & n3521 ;
  assign n3523 = ( x222 & x940 ) | ( x222 & ~n1811 ) | ( x940 & ~n1811 ) ;
  assign n3524 = ( x222 & x1138 ) | ( x222 & n1811 ) | ( x1138 & n1811 ) ;
  assign n3525 = n3523 & n3524 ;
  assign n3526 = n3522 | n3525 ;
  assign n3527 = n3517 | n3526 ;
  assign n3528 = n2227 & ~n3519 ;
  assign n3529 = n3526 | n3528 ;
  assign n3530 = ~x223 & n3529 ;
  assign n3531 = n3517 | n3530 ;
  assign n3532 = ~x39 & n3531 ;
  assign n3533 = n3527 & n3532 ;
  assign n3534 = ~n3515 & n3533 ;
  assign n3535 = x224 | n3502 ;
  assign n3536 = ~n3519 & n3535 ;
  assign n3537 = n3525 | n3536 ;
  assign n3538 = ~x223 & n3537 ;
  assign n3539 = n3516 | n3538 ;
  assign n3540 = ~x299 & n3539 ;
  assign n3541 = x216 | n3505 ;
  assign n3542 = ( x169 & x228 ) | ( x169 & n1868 ) | ( x228 & n1868 ) ;
  assign n3543 = ( ~x228 & x877 ) | ( ~x228 & n1868 ) | ( x877 & n1868 ) ;
  assign n3544 = ~n3542 & n3543 ;
  assign n3545 = n3541 | n3544 ;
  assign n3546 = ~n3494 & n3545 ;
  assign n3547 = n3512 | n3546 ;
  assign n3548 = ~x215 & n3547 ;
  assign n3549 = n3491 | n3548 ;
  assign n3550 = x299 & n3549 ;
  assign n3551 = n3540 | n3550 ;
  assign n3552 = x39 & n3551 ;
  assign n3553 = x38 | n3552 ;
  assign n3554 = n3534 | n3553 ;
  assign n3555 = x169 | x228 ;
  assign n3556 = ~n3541 & n3555 ;
  assign n3557 = n3494 | n3556 ;
  assign n3558 = ~n3512 & n3557 ;
  assign n3559 = x215 | n3558 ;
  assign n3560 = ~n3491 & n3559 ;
  assign n3561 = x299 & ~n3560 ;
  assign n3562 = n3540 | n3561 ;
  assign n3563 = x38 & ~n3562 ;
  assign n3564 = x100 | n3563 ;
  assign n3565 = n3554 & ~n3564 ;
  assign n3566 = n1925 | n3540 ;
  assign n3567 = ( x169 & x228 ) | ( x169 & n2161 ) | ( x228 & n2161 ) ;
  assign n3568 = ( ~x228 & x877 ) | ( ~x228 & n2161 ) | ( x877 & n2161 ) ;
  assign n3569 = ~n3567 & n3568 ;
  assign n3570 = n3541 | n3569 ;
  assign n3571 = ~n3494 & n3570 ;
  assign n3572 = n3512 | n3571 ;
  assign n3573 = ~x215 & n3572 ;
  assign n3574 = n3492 & ~n3573 ;
  assign n3575 = ( x299 & n3566 ) | ( x299 & ~n3574 ) | ( n3566 & ~n3574 ) ;
  assign n3576 = ( x100 & n2364 ) | ( x100 & n3562 ) | ( n2364 & n3562 ) ;
  assign n3577 = n3575 & n3576 ;
  assign n3578 = n3565 | n3577 ;
  assign n3579 = ~x87 & n3578 ;
  assign n3580 = n1976 & ~n3562 ;
  assign n3581 = n1976 | n3551 ;
  assign n3582 = ~n3580 & n3581 ;
  assign n3583 = ( x75 & n1998 ) | ( x75 & n3582 ) | ( n1998 & n3582 ) ;
  assign n3584 = n3579 | n3583 ;
  assign n3585 = x75 & ~n3562 ;
  assign n3586 = x92 | n3585 ;
  assign n3587 = n3584 & ~n3586 ;
  assign n3588 = ( x92 & ~n1998 ) | ( x92 & n3562 ) | ( ~n1998 & n3562 ) ;
  assign n3589 = ( x92 & n1998 ) | ( x92 & n3582 ) | ( n1998 & n3582 ) ;
  assign n3590 = n3588 & n3589 ;
  assign n3591 = n2030 | n3590 ;
  assign n3592 = n3587 | n3591 ;
  assign n3593 = n2030 & ~n3562 ;
  assign n3594 = x55 | n3593 ;
  assign n3595 = n3592 & ~n3594 ;
  assign n3596 = ( x55 & n2033 ) | ( x55 & n3549 ) | ( n2033 & n3549 ) ;
  assign n3597 = ( ~x55 & n2033 ) | ( ~x55 & n3560 ) | ( n2033 & n3560 ) ;
  assign n3598 = n3596 & ~n3597 ;
  assign n3599 = x56 | n3598 ;
  assign n3600 = n3595 | n3599 ;
  assign n3601 = ( x56 & n2045 ) | ( x56 & ~n3549 ) | ( n2045 & ~n3549 ) ;
  assign n3602 = ( x56 & ~n2045 ) | ( x56 & n3560 ) | ( ~n2045 & n3560 ) ;
  assign n3603 = n3601 & n3602 ;
  assign n3604 = x62 | n3603 ;
  assign n3605 = n3600 & ~n3604 ;
  assign n3606 = x246 | n2057 ;
  assign n3607 = ( x62 & n2193 ) | ( x62 & n3549 ) | ( n2193 & n3549 ) ;
  assign n3608 = ( ~x62 & n2193 ) | ( ~x62 & n3560 ) | ( n2193 & n3560 ) ;
  assign n3609 = n3607 & ~n3608 ;
  assign n3610 = n3606 | n3609 ;
  assign n3611 = n3605 | n3610 ;
  assign n3612 = ~x877 & n2239 ;
  assign n3613 = x169 | n3612 ;
  assign n3614 = ( x169 & ~x877 ) | ( x169 & n2138 ) | ( ~x877 & n2138 ) ;
  assign n3615 = ( x169 & x877 ) | ( x169 & n2230 ) | ( x877 & n2230 ) ;
  assign n3616 = n3614 & n3615 ;
  assign n3617 = n3613 & ~n3616 ;
  assign n3618 = x228 | n3617 ;
  assign n3619 = n2588 | n3541 ;
  assign n3620 = n3618 & ~n3619 ;
  assign n3621 = n3494 | n3620 ;
  assign n3622 = ~n3512 & n3621 ;
  assign n3623 = x215 | n3622 ;
  assign n3624 = n3492 & n3623 ;
  assign n3625 = n3532 & ~n3624 ;
  assign n3626 = n2215 | n3540 ;
  assign n3627 = n2205 | n3541 ;
  assign n3628 = n3544 | n3627 ;
  assign n3629 = ~n3494 & n3628 ;
  assign n3630 = n3512 | n3629 ;
  assign n3631 = ~x215 & n3630 ;
  assign n3632 = n3491 | n3631 ;
  assign n3633 = x299 & n3632 ;
  assign n3634 = n3626 | n3633 ;
  assign n3635 = x39 & n3634 ;
  assign n3636 = x38 | n3635 ;
  assign n3637 = n3625 | n3636 ;
  assign n3638 = n2345 & ~n3493 ;
  assign n3639 = n3560 & ~n3638 ;
  assign n3640 = x299 & ~n3639 ;
  assign n3641 = n3626 | n3640 ;
  assign n3642 = x38 & ~n3641 ;
  assign n3643 = x100 | n3642 ;
  assign n3644 = n3637 & ~n3643 ;
  assign n3645 = n1925 | n3626 ;
  assign n3646 = n3569 | n3627 ;
  assign n3647 = ~n3494 & n3646 ;
  assign n3648 = n3512 | n3647 ;
  assign n3649 = ~x215 & n3648 ;
  assign n3650 = n3492 & ~n3649 ;
  assign n3651 = ( x299 & n3645 ) | ( x299 & ~n3650 ) | ( n3645 & ~n3650 ) ;
  assign n3652 = ( x100 & n2364 ) | ( x100 & n3641 ) | ( n2364 & n3641 ) ;
  assign n3653 = n3651 & n3652 ;
  assign n3654 = n3644 | n3653 ;
  assign n3655 = ~x87 & n3654 ;
  assign n3656 = n1976 & ~n3641 ;
  assign n3657 = n1976 | n3634 ;
  assign n3658 = ~n3656 & n3657 ;
  assign n3659 = ( x75 & n1998 ) | ( x75 & n3658 ) | ( n1998 & n3658 ) ;
  assign n3660 = n3655 | n3659 ;
  assign n3661 = x75 & ~n3641 ;
  assign n3662 = x92 | n3661 ;
  assign n3663 = n3660 & ~n3662 ;
  assign n3664 = ( x92 & ~n1998 ) | ( x92 & n3641 ) | ( ~n1998 & n3641 ) ;
  assign n3665 = ( x92 & n1998 ) | ( x92 & n3658 ) | ( n1998 & n3658 ) ;
  assign n3666 = n3664 & n3665 ;
  assign n3667 = n2030 | n3666 ;
  assign n3668 = n3663 | n3667 ;
  assign n3669 = n2030 & ~n3641 ;
  assign n3670 = x55 | n3669 ;
  assign n3671 = n3668 & ~n3670 ;
  assign n3672 = ( x55 & n2033 ) | ( x55 & n3632 ) | ( n2033 & n3632 ) ;
  assign n3673 = ( ~x55 & n2033 ) | ( ~x55 & n3639 ) | ( n2033 & n3639 ) ;
  assign n3674 = n3672 & ~n3673 ;
  assign n3675 = x56 | n3674 ;
  assign n3676 = n3671 | n3675 ;
  assign n3677 = ( x56 & n2045 ) | ( x56 & ~n3632 ) | ( n2045 & ~n3632 ) ;
  assign n3678 = ( x56 & ~n2045 ) | ( x56 & n3639 ) | ( ~n2045 & n3639 ) ;
  assign n3679 = n3677 & n3678 ;
  assign n3680 = x62 | n3679 ;
  assign n3681 = n3676 & ~n3680 ;
  assign n3682 = x246 & ~n2057 ;
  assign n3683 = ( x62 & n2193 ) | ( x62 & n3632 ) | ( n2193 & n3632 ) ;
  assign n3684 = ( ~x62 & n2193 ) | ( ~x62 & n3639 ) | ( n2193 & n3639 ) ;
  assign n3685 = n3683 & ~n3684 ;
  assign n3686 = n3682 & ~n3685 ;
  assign n3687 = ~n3681 & n3686 ;
  assign n3688 = x246 & n3638 ;
  assign n3689 = n2057 & ~n3688 ;
  assign n3690 = n3560 & n3689 ;
  assign n3691 = n3687 | n3690 ;
  assign n3692 = n3611 & ~n3691 ;
  assign n3693 = x215 & x1137 ;
  assign n3694 = x299 & ~n3693 ;
  assign n3695 = x216 & x280 ;
  assign n3696 = x221 | n3695 ;
  assign n3697 = x878 & n2230 ;
  assign n3698 = x168 | n3697 ;
  assign n3699 = x168 & n2239 ;
  assign n3700 = n3698 & ~n3699 ;
  assign n3701 = n2138 | n3698 ;
  assign n3702 = ( ~x878 & n3700 ) | ( ~x878 & n3701 ) | ( n3700 & n3701 ) ;
  assign n3703 = x228 | n3702 ;
  assign n3704 = x878 & ~n1491 ;
  assign n3705 = ( ~x105 & x228 ) | ( ~x105 & n3704 ) | ( x228 & n3704 ) ;
  assign n3706 = ( x105 & ~x168 ) | ( x105 & x228 ) | ( ~x168 & x228 ) ;
  assign n3707 = n3705 & n3706 ;
  assign n3708 = ~n2228 & n3707 ;
  assign n3709 = x216 | n3708 ;
  assign n3710 = n3703 & ~n3709 ;
  assign n3711 = n3696 | n3710 ;
  assign n3712 = ( x221 & x933 ) | ( x221 & ~n1205 ) | ( x933 & ~n1205 ) ;
  assign n3713 = ( x221 & x1137 ) | ( x221 & n1205 ) | ( x1137 & n1205 ) ;
  assign n3714 = n3712 & n3713 ;
  assign n3715 = n3711 & ~n3714 ;
  assign n3716 = x215 | n3715 ;
  assign n3717 = n3694 & n3716 ;
  assign n3718 = x223 & x1137 ;
  assign n3719 = x299 | n3718 ;
  assign n3720 = x224 & x280 ;
  assign n3721 = x222 | n3720 ;
  assign n3722 = x878 & ~n2227 ;
  assign n3723 = x224 | n3722 ;
  assign n3724 = ~n3721 & n3723 ;
  assign n3725 = ( x222 & x933 ) | ( x222 & ~n1811 ) | ( x933 & ~n1811 ) ;
  assign n3726 = ( x222 & x1137 ) | ( x222 & n1811 ) | ( x1137 & n1811 ) ;
  assign n3727 = n3725 & n3726 ;
  assign n3728 = n3724 | n3727 ;
  assign n3729 = n3719 | n3728 ;
  assign n3730 = n2227 & ~n3721 ;
  assign n3731 = n3728 | n3730 ;
  assign n3732 = ~x223 & n3731 ;
  assign n3733 = n3719 | n3732 ;
  assign n3734 = ~x39 & n3733 ;
  assign n3735 = n3729 & n3734 ;
  assign n3736 = ~n3717 & n3735 ;
  assign n3737 = x224 | n3704 ;
  assign n3738 = ~n3721 & n3737 ;
  assign n3739 = n3727 | n3738 ;
  assign n3740 = ~x223 & n3739 ;
  assign n3741 = n3718 | n3740 ;
  assign n3742 = ~x299 & n3741 ;
  assign n3743 = x216 | n3707 ;
  assign n3744 = ( x168 & x228 ) | ( x168 & n1868 ) | ( x228 & n1868 ) ;
  assign n3745 = ( ~x228 & x878 ) | ( ~x228 & n1868 ) | ( x878 & n1868 ) ;
  assign n3746 = ~n3744 & n3745 ;
  assign n3747 = n3743 | n3746 ;
  assign n3748 = ~n3696 & n3747 ;
  assign n3749 = n3714 | n3748 ;
  assign n3750 = ~x215 & n3749 ;
  assign n3751 = n3693 | n3750 ;
  assign n3752 = x299 & n3751 ;
  assign n3753 = n3742 | n3752 ;
  assign n3754 = x39 & n3753 ;
  assign n3755 = x38 | n3754 ;
  assign n3756 = n3736 | n3755 ;
  assign n3757 = x168 | x228 ;
  assign n3758 = ~n3743 & n3757 ;
  assign n3759 = n3696 | n3758 ;
  assign n3760 = ~n3714 & n3759 ;
  assign n3761 = x215 | n3760 ;
  assign n3762 = ~n3693 & n3761 ;
  assign n3763 = x299 & ~n3762 ;
  assign n3764 = n3742 | n3763 ;
  assign n3765 = x38 & ~n3764 ;
  assign n3766 = x100 | n3765 ;
  assign n3767 = n3756 & ~n3766 ;
  assign n3768 = n1925 | n3742 ;
  assign n3769 = ( x168 & x228 ) | ( x168 & n2161 ) | ( x228 & n2161 ) ;
  assign n3770 = ( ~x228 & x878 ) | ( ~x228 & n2161 ) | ( x878 & n2161 ) ;
  assign n3771 = ~n3769 & n3770 ;
  assign n3772 = n3743 | n3771 ;
  assign n3773 = ~n3696 & n3772 ;
  assign n3774 = n3714 | n3773 ;
  assign n3775 = ~x215 & n3774 ;
  assign n3776 = n3694 & ~n3775 ;
  assign n3777 = ( x299 & n3768 ) | ( x299 & ~n3776 ) | ( n3768 & ~n3776 ) ;
  assign n3778 = ( x100 & n2364 ) | ( x100 & n3764 ) | ( n2364 & n3764 ) ;
  assign n3779 = n3777 & n3778 ;
  assign n3780 = n3767 | n3779 ;
  assign n3781 = ~x87 & n3780 ;
  assign n3782 = n1976 & ~n3764 ;
  assign n3783 = n1976 | n3753 ;
  assign n3784 = ~n3782 & n3783 ;
  assign n3785 = ( x75 & n1998 ) | ( x75 & n3784 ) | ( n1998 & n3784 ) ;
  assign n3786 = n3781 | n3785 ;
  assign n3787 = x75 & ~n3764 ;
  assign n3788 = x92 | n3787 ;
  assign n3789 = n3786 & ~n3788 ;
  assign n3790 = ( x92 & ~n1998 ) | ( x92 & n3764 ) | ( ~n1998 & n3764 ) ;
  assign n3791 = ( x92 & n1998 ) | ( x92 & n3784 ) | ( n1998 & n3784 ) ;
  assign n3792 = n3790 & n3791 ;
  assign n3793 = n2030 | n3792 ;
  assign n3794 = n3789 | n3793 ;
  assign n3795 = n2030 & ~n3764 ;
  assign n3796 = x55 | n3795 ;
  assign n3797 = n3794 & ~n3796 ;
  assign n3798 = ( x55 & n2033 ) | ( x55 & n3751 ) | ( n2033 & n3751 ) ;
  assign n3799 = ( ~x55 & n2033 ) | ( ~x55 & n3762 ) | ( n2033 & n3762 ) ;
  assign n3800 = n3798 & ~n3799 ;
  assign n3801 = x56 | n3800 ;
  assign n3802 = n3797 | n3801 ;
  assign n3803 = ( x56 & n2045 ) | ( x56 & ~n3751 ) | ( n2045 & ~n3751 ) ;
  assign n3804 = ( x56 & ~n2045 ) | ( x56 & n3762 ) | ( ~n2045 & n3762 ) ;
  assign n3805 = n3803 & n3804 ;
  assign n3806 = x62 | n3805 ;
  assign n3807 = n3802 & ~n3806 ;
  assign n3808 = x240 | n2057 ;
  assign n3809 = ( x62 & n2193 ) | ( x62 & n3751 ) | ( n2193 & n3751 ) ;
  assign n3810 = ( ~x62 & n2193 ) | ( ~x62 & n3762 ) | ( n2193 & n3762 ) ;
  assign n3811 = n3809 & ~n3810 ;
  assign n3812 = n3808 | n3811 ;
  assign n3813 = n3807 | n3812 ;
  assign n3814 = ~x878 & n2239 ;
  assign n3815 = x168 | n3814 ;
  assign n3816 = ( x168 & ~x878 ) | ( x168 & n2138 ) | ( ~x878 & n2138 ) ;
  assign n3817 = ( x168 & x878 ) | ( x168 & n2230 ) | ( x878 & n2230 ) ;
  assign n3818 = n3816 & n3817 ;
  assign n3819 = n3815 & ~n3818 ;
  assign n3820 = x228 | n3819 ;
  assign n3821 = n2588 | n3743 ;
  assign n3822 = n3820 & ~n3821 ;
  assign n3823 = n3696 | n3822 ;
  assign n3824 = ~n3714 & n3823 ;
  assign n3825 = x215 | n3824 ;
  assign n3826 = n3694 & n3825 ;
  assign n3827 = n3734 & ~n3826 ;
  assign n3828 = n2215 | n3742 ;
  assign n3829 = n2205 | n3743 ;
  assign n3830 = n3746 | n3829 ;
  assign n3831 = ~n3696 & n3830 ;
  assign n3832 = n3714 | n3831 ;
  assign n3833 = ~x215 & n3832 ;
  assign n3834 = n3693 | n3833 ;
  assign n3835 = x299 & n3834 ;
  assign n3836 = n3828 | n3835 ;
  assign n3837 = x39 & n3836 ;
  assign n3838 = x38 | n3837 ;
  assign n3839 = n3827 | n3838 ;
  assign n3840 = n2345 & ~n3695 ;
  assign n3841 = n3762 & ~n3840 ;
  assign n3842 = x299 & ~n3841 ;
  assign n3843 = n3828 | n3842 ;
  assign n3844 = x38 & ~n3843 ;
  assign n3845 = x100 | n3844 ;
  assign n3846 = n3839 & ~n3845 ;
  assign n3847 = n1925 | n3828 ;
  assign n3848 = n3771 | n3829 ;
  assign n3849 = ~n3696 & n3848 ;
  assign n3850 = n3714 | n3849 ;
  assign n3851 = ~x215 & n3850 ;
  assign n3852 = n3694 & ~n3851 ;
  assign n3853 = ( x299 & n3847 ) | ( x299 & ~n3852 ) | ( n3847 & ~n3852 ) ;
  assign n3854 = ( x100 & n2364 ) | ( x100 & n3843 ) | ( n2364 & n3843 ) ;
  assign n3855 = n3853 & n3854 ;
  assign n3856 = n3846 | n3855 ;
  assign n3857 = ~x87 & n3856 ;
  assign n3858 = n1976 & ~n3843 ;
  assign n3859 = n1976 | n3836 ;
  assign n3860 = ~n3858 & n3859 ;
  assign n3861 = ( x75 & n1998 ) | ( x75 & n3860 ) | ( n1998 & n3860 ) ;
  assign n3862 = n3857 | n3861 ;
  assign n3863 = x75 & ~n3843 ;
  assign n3864 = x92 | n3863 ;
  assign n3865 = n3862 & ~n3864 ;
  assign n3866 = ( x92 & ~n1998 ) | ( x92 & n3843 ) | ( ~n1998 & n3843 ) ;
  assign n3867 = ( x92 & n1998 ) | ( x92 & n3860 ) | ( n1998 & n3860 ) ;
  assign n3868 = n3866 & n3867 ;
  assign n3869 = n2030 | n3868 ;
  assign n3870 = n3865 | n3869 ;
  assign n3871 = n2030 & ~n3843 ;
  assign n3872 = x55 | n3871 ;
  assign n3873 = n3870 & ~n3872 ;
  assign n3874 = ( x55 & n2033 ) | ( x55 & n3834 ) | ( n2033 & n3834 ) ;
  assign n3875 = ( ~x55 & n2033 ) | ( ~x55 & n3841 ) | ( n2033 & n3841 ) ;
  assign n3876 = n3874 & ~n3875 ;
  assign n3877 = x56 | n3876 ;
  assign n3878 = n3873 | n3877 ;
  assign n3879 = ( x56 & n2045 ) | ( x56 & ~n3834 ) | ( n2045 & ~n3834 ) ;
  assign n3880 = ( x56 & ~n2045 ) | ( x56 & n3841 ) | ( ~n2045 & n3841 ) ;
  assign n3881 = n3879 & n3880 ;
  assign n3882 = x62 | n3881 ;
  assign n3883 = n3878 & ~n3882 ;
  assign n3884 = x240 & ~n2057 ;
  assign n3885 = ( x62 & n2193 ) | ( x62 & n3834 ) | ( n2193 & n3834 ) ;
  assign n3886 = ( ~x62 & n2193 ) | ( ~x62 & n3841 ) | ( n2193 & n3841 ) ;
  assign n3887 = n3885 & ~n3886 ;
  assign n3888 = n3884 & ~n3887 ;
  assign n3889 = ~n3883 & n3888 ;
  assign n3890 = x240 & n3840 ;
  assign n3891 = n2057 & ~n3890 ;
  assign n3892 = n3762 & n3891 ;
  assign n3893 = n3889 | n3892 ;
  assign n3894 = n3813 & ~n3893 ;
  assign n3895 = x216 & x266 ;
  assign n3896 = x875 & ~n1491 ;
  assign n3897 = x105 & ~n3896 ;
  assign n3898 = x105 | x166 ;
  assign n3899 = ~n3897 & n3898 ;
  assign n3900 = n2229 & ~n3899 ;
  assign n3901 = x216 | n3900 ;
  assign n3902 = x166 & ~x875 ;
  assign n3903 = ~n2138 & n3902 ;
  assign n3904 = ( x166 & ~x875 ) | ( x166 & n2230 ) | ( ~x875 & n2230 ) ;
  assign n3905 = ( x166 & x875 ) | ( x166 & n2239 ) | ( x875 & n2239 ) ;
  assign n3906 = ~n3904 & n3905 ;
  assign n3907 = n3903 | n3906 ;
  assign n3908 = ~x228 & n3907 ;
  assign n3909 = n2229 | n3908 ;
  assign n3910 = ~n3901 & n3909 ;
  assign n3911 = n3895 | n3910 ;
  assign n3912 = ~x221 & n3911 ;
  assign n3913 = ( x221 & x928 ) | ( x221 & ~n1205 ) | ( x928 & ~n1205 ) ;
  assign n3914 = ( x221 & x1136 ) | ( x221 & n1205 ) | ( x1136 & n1205 ) ;
  assign n3915 = n3913 & n3914 ;
  assign n3916 = n3912 | n3915 ;
  assign n3917 = ~x215 & n3916 ;
  assign n3918 = x215 & x1136 ;
  assign n3919 = x299 & ~n3918 ;
  assign n3920 = ~n3917 & n3919 ;
  assign n3921 = x224 | x875 ;
  assign n3922 = n1491 | n3921 ;
  assign n3923 = x224 & ~x266 ;
  assign n3924 = x222 | n3923 ;
  assign n3925 = n3922 & ~n3924 ;
  assign n3926 = ~n1823 & n2227 ;
  assign n3927 = n3925 & ~n3926 ;
  assign n3928 = x223 & x1136 ;
  assign n3929 = x299 | n3928 ;
  assign n3930 = ( x222 & x928 ) | ( x222 & ~n1811 ) | ( x928 & ~n1811 ) ;
  assign n3931 = ( x222 & x1136 ) | ( x222 & n1811 ) | ( x1136 & n1811 ) ;
  assign n3932 = n3930 & n3931 ;
  assign n3933 = n3929 | n3932 ;
  assign n3934 = n3927 | n3933 ;
  assign n3935 = n3925 | n3932 ;
  assign n3936 = n3926 | n3935 ;
  assign n3937 = ~x223 & n3936 ;
  assign n3938 = n3929 | n3937 ;
  assign n3939 = ~x39 & n3938 ;
  assign n3940 = n3934 & n3939 ;
  assign n3941 = ~n3920 & n3940 ;
  assign n3942 = ~x223 & n3935 ;
  assign n3943 = n3928 | n3942 ;
  assign n3944 = ~x299 & n3943 ;
  assign n3945 = n1873 | n3896 ;
  assign n3946 = n3944 & n3945 ;
  assign n3947 = x228 & n3899 ;
  assign n3948 = ( ~x166 & x228 ) | ( ~x166 & n1868 ) | ( x228 & n1868 ) ;
  assign n3949 = ( ~x228 & x875 ) | ( ~x228 & n1868 ) | ( x875 & n1868 ) ;
  assign n3950 = ~n3948 & n3949 ;
  assign n3951 = n3947 | n3950 ;
  assign n3952 = ~x216 & n3951 ;
  assign n3953 = n3895 | n3952 ;
  assign n3954 = ~x221 & n3953 ;
  assign n3955 = n3915 | n3954 ;
  assign n3956 = ~x215 & n3955 ;
  assign n3957 = n3918 | n3956 ;
  assign n3958 = x299 & n3957 ;
  assign n3959 = n3946 | n3958 ;
  assign n3960 = x39 & n3959 ;
  assign n3961 = x38 | n3960 ;
  assign n3962 = n3941 | n3961 ;
  assign n3963 = x166 & ~x228 ;
  assign n3964 = n3947 | n3963 ;
  assign n3965 = ~x216 & n3964 ;
  assign n3966 = n3895 | n3965 ;
  assign n3967 = ~x221 & n3966 ;
  assign n3968 = n3915 | n3967 ;
  assign n3969 = ~x215 & n3968 ;
  assign n3970 = n3918 | n3969 ;
  assign n3971 = x299 & n3970 ;
  assign n3972 = n3946 | n3971 ;
  assign n3973 = x38 & ~n3972 ;
  assign n3974 = x100 | n3973 ;
  assign n3975 = n3962 & ~n3974 ;
  assign n3976 = n1925 | n3946 ;
  assign n3977 = ( ~x875 & n1523 ) | ( ~x875 & n2155 ) | ( n1523 & n2155 ) ;
  assign n3978 = ( x875 & n1523 ) | ( x875 & ~n2153 ) | ( n1523 & ~n2153 ) ;
  assign n3979 = ~n3977 & n3978 ;
  assign n3980 = ~n2155 & n3902 ;
  assign n3981 = ( x166 & n3979 ) | ( x166 & ~n3980 ) | ( n3979 & ~n3980 ) ;
  assign n3982 = ~x228 & n3981 ;
  assign n3983 = n3947 | n3982 ;
  assign n3984 = ~x216 & n3983 ;
  assign n3985 = n3895 | n3984 ;
  assign n3986 = ~x221 & n3985 ;
  assign n3987 = n3915 | n3986 ;
  assign n3988 = ~x215 & n3987 ;
  assign n3989 = n3919 & ~n3988 ;
  assign n3990 = ( x299 & n3976 ) | ( x299 & ~n3989 ) | ( n3976 & ~n3989 ) ;
  assign n3991 = ( x100 & n2364 ) | ( x100 & n3972 ) | ( n2364 & n3972 ) ;
  assign n3992 = n3990 & n3991 ;
  assign n3993 = n3975 | n3992 ;
  assign n3994 = ~x87 & n3993 ;
  assign n3995 = n1976 & ~n3972 ;
  assign n3996 = n1976 | n3959 ;
  assign n3997 = ~n3995 & n3996 ;
  assign n3998 = ( x75 & n1998 ) | ( x75 & n3997 ) | ( n1998 & n3997 ) ;
  assign n3999 = n3994 | n3998 ;
  assign n4000 = x75 & ~n3972 ;
  assign n4001 = x92 | n4000 ;
  assign n4002 = n3999 & ~n4001 ;
  assign n4003 = ( x92 & ~n1998 ) | ( x92 & n3972 ) | ( ~n1998 & n3972 ) ;
  assign n4004 = ( x92 & n1998 ) | ( x92 & n3997 ) | ( n1998 & n3997 ) ;
  assign n4005 = n4003 & n4004 ;
  assign n4006 = n2030 | n4005 ;
  assign n4007 = n4002 | n4006 ;
  assign n4008 = n2030 & ~n3972 ;
  assign n4009 = x55 | n4008 ;
  assign n4010 = n4007 & ~n4009 ;
  assign n4011 = ( x55 & ~n2033 ) | ( x55 & n3970 ) | ( ~n2033 & n3970 ) ;
  assign n4012 = ( x55 & n2033 ) | ( x55 & n3957 ) | ( n2033 & n3957 ) ;
  assign n4013 = n4011 & n4012 ;
  assign n4014 = x56 | n4013 ;
  assign n4015 = n4010 | n4014 ;
  assign n4016 = ( ~x56 & n2045 ) | ( ~x56 & n3970 ) | ( n2045 & n3970 ) ;
  assign n4017 = ( x56 & n2045 ) | ( x56 & ~n3957 ) | ( n2045 & ~n3957 ) ;
  assign n4018 = ~n4016 & n4017 ;
  assign n4019 = x62 | n4018 ;
  assign n4020 = n4015 & ~n4019 ;
  assign n4021 = ( x62 & ~n2193 ) | ( x62 & n3970 ) | ( ~n2193 & n3970 ) ;
  assign n4022 = ( x62 & n2193 ) | ( x62 & n3957 ) | ( n2193 & n3957 ) ;
  assign n4023 = n4021 & n4022 ;
  assign n4024 = n2057 | n4023 ;
  assign n4025 = n4020 | n4024 ;
  assign n4026 = n2057 & ~n3970 ;
  assign n4027 = x245 | n4026 ;
  assign n4028 = n4025 & ~n4027 ;
  assign n4029 = x166 | n2138 ;
  assign n4030 = x875 & n4029 ;
  assign n4031 = n3904 & ~n3905 ;
  assign n4032 = x228 | n4031 ;
  assign n4033 = n4030 | n4032 ;
  assign n4034 = ~n3901 & n4033 ;
  assign n4035 = n3895 | n4034 ;
  assign n4036 = ~x221 & n4035 ;
  assign n4037 = n3915 | n4036 ;
  assign n4038 = ~x215 & n4037 ;
  assign n4039 = n3919 & ~n4038 ;
  assign n4040 = n3939 & ~n4039 ;
  assign n4041 = n2205 | n3947 ;
  assign n4042 = n3950 | n4041 ;
  assign n4043 = ~x216 & n4042 ;
  assign n4044 = n3895 | n4043 ;
  assign n4045 = ~x221 & n4044 ;
  assign n4046 = n3915 | n4045 ;
  assign n4047 = ~x215 & n4046 ;
  assign n4048 = n3918 | n4047 ;
  assign n4049 = x299 & n4048 ;
  assign n4050 = n3944 | n4049 ;
  assign n4051 = x39 & n4050 ;
  assign n4052 = x38 | n4051 ;
  assign n4053 = n4040 | n4052 ;
  assign n4054 = n2206 | n3970 ;
  assign n4055 = x299 & n4054 ;
  assign n4056 = n3944 | n4055 ;
  assign n4057 = x38 & ~n4056 ;
  assign n4058 = x100 | n4057 ;
  assign n4059 = n4053 & ~n4058 ;
  assign n4060 = n1925 | n3944 ;
  assign n4061 = n3982 | n4041 ;
  assign n4062 = ~x216 & n4061 ;
  assign n4063 = n3895 | n4062 ;
  assign n4064 = ~x221 & n4063 ;
  assign n4065 = n3915 | n4064 ;
  assign n4066 = ~x215 & n4065 ;
  assign n4067 = n3919 & ~n4066 ;
  assign n4068 = ( x299 & n4060 ) | ( x299 & ~n4067 ) | ( n4060 & ~n4067 ) ;
  assign n4069 = ( x100 & n2364 ) | ( x100 & n4056 ) | ( n2364 & n4056 ) ;
  assign n4070 = n4068 & n4069 ;
  assign n4071 = n4059 | n4070 ;
  assign n4072 = ~x87 & n4071 ;
  assign n4073 = n1976 & ~n4056 ;
  assign n4074 = n1976 | n4050 ;
  assign n4075 = ~n4073 & n4074 ;
  assign n4076 = ( x75 & n1998 ) | ( x75 & n4075 ) | ( n1998 & n4075 ) ;
  assign n4077 = n4072 | n4076 ;
  assign n4078 = x75 & ~n4056 ;
  assign n4079 = x92 | n4078 ;
  assign n4080 = n4077 & ~n4079 ;
  assign n4081 = ( x92 & ~n1998 ) | ( x92 & n4056 ) | ( ~n1998 & n4056 ) ;
  assign n4082 = ( x92 & n1998 ) | ( x92 & n4075 ) | ( n1998 & n4075 ) ;
  assign n4083 = n4081 & n4082 ;
  assign n4084 = n2030 | n4083 ;
  assign n4085 = n4080 | n4084 ;
  assign n4086 = n2030 & ~n4056 ;
  assign n4087 = x55 | n4086 ;
  assign n4088 = n4085 & ~n4087 ;
  assign n4089 = ( x55 & ~n2033 ) | ( x55 & n4054 ) | ( ~n2033 & n4054 ) ;
  assign n4090 = ( x55 & n2033 ) | ( x55 & n4048 ) | ( n2033 & n4048 ) ;
  assign n4091 = n4089 & n4090 ;
  assign n4092 = x56 | n4091 ;
  assign n4093 = n4088 | n4092 ;
  assign n4094 = ( ~x56 & n2045 ) | ( ~x56 & n4054 ) | ( n2045 & n4054 ) ;
  assign n4095 = ( x56 & n2045 ) | ( x56 & ~n4048 ) | ( n2045 & ~n4048 ) ;
  assign n4096 = ~n4094 & n4095 ;
  assign n4097 = x62 | n4096 ;
  assign n4098 = n4093 & ~n4097 ;
  assign n4099 = ( x62 & ~n2193 ) | ( x62 & n4054 ) | ( ~n2193 & n4054 ) ;
  assign n4100 = ( x62 & n2193 ) | ( x62 & n4048 ) | ( n2193 & n4048 ) ;
  assign n4101 = n4099 & n4100 ;
  assign n4102 = n2057 | n4101 ;
  assign n4103 = n4098 | n4102 ;
  assign n4104 = n2057 & ~n4054 ;
  assign n4105 = x245 & ~n4104 ;
  assign n4106 = n4103 & n4105 ;
  assign n4107 = n4028 | n4106 ;
  assign n4108 = x216 & x279 ;
  assign n4109 = x879 & ~n1491 ;
  assign n4110 = x105 & ~n4109 ;
  assign n4111 = x105 | x161 ;
  assign n4112 = ~n4110 & n4111 ;
  assign n4113 = n2229 & ~n4112 ;
  assign n4114 = x216 | n4113 ;
  assign n4115 = x161 & ~x879 ;
  assign n4116 = ~n2138 & n4115 ;
  assign n4117 = ( x161 & ~x879 ) | ( x161 & n2230 ) | ( ~x879 & n2230 ) ;
  assign n4118 = ( x161 & x879 ) | ( x161 & n2239 ) | ( x879 & n2239 ) ;
  assign n4119 = ~n4117 & n4118 ;
  assign n4120 = n4116 | n4119 ;
  assign n4121 = ~x228 & n4120 ;
  assign n4122 = n2229 | n4121 ;
  assign n4123 = ~n4114 & n4122 ;
  assign n4124 = n4108 | n4123 ;
  assign n4125 = ~x221 & n4124 ;
  assign n4126 = ( x221 & x938 ) | ( x221 & ~n1205 ) | ( x938 & ~n1205 ) ;
  assign n4127 = ( x221 & x1135 ) | ( x221 & n1205 ) | ( x1135 & n1205 ) ;
  assign n4128 = n4126 & n4127 ;
  assign n4129 = n4125 | n4128 ;
  assign n4130 = ~x215 & n4129 ;
  assign n4131 = x215 & x1135 ;
  assign n4132 = x299 & ~n4131 ;
  assign n4133 = ~n4130 & n4132 ;
  assign n4134 = x223 & x1135 ;
  assign n4135 = x299 | n4134 ;
  assign n4136 = x224 | x879 ;
  assign n4137 = n1491 | n4136 ;
  assign n4138 = x224 & ~x279 ;
  assign n4139 = x222 | n4138 ;
  assign n4140 = n4137 & ~n4139 ;
  assign n4141 = ( x222 & x938 ) | ( x222 & ~n1811 ) | ( x938 & ~n1811 ) ;
  assign n4142 = ( x222 & x1135 ) | ( x222 & n1811 ) | ( x1135 & n1811 ) ;
  assign n4143 = n4141 & n4142 ;
  assign n4144 = n4140 | n4143 ;
  assign n4145 = ~x223 & n4144 ;
  assign n4146 = n3926 & ~n4143 ;
  assign n4147 = n4145 & ~n4146 ;
  assign n4148 = n4135 | n4147 ;
  assign n4149 = ~x39 & n4148 ;
  assign n4150 = ~n4133 & n4149 ;
  assign n4151 = n4134 | n4145 ;
  assign n4152 = ~x299 & n4151 ;
  assign n4153 = n1873 | n4109 ;
  assign n4154 = n4152 & n4153 ;
  assign n4155 = x228 & n4112 ;
  assign n4156 = x879 | n1868 ;
  assign n4157 = x161 & ~x228 ;
  assign n4158 = n2082 & ~n4157 ;
  assign n4159 = n4156 & ~n4158 ;
  assign n4160 = n4155 | n4159 ;
  assign n4161 = ~x216 & n4160 ;
  assign n4162 = n4108 | n4161 ;
  assign n4163 = ~x221 & n4162 ;
  assign n4164 = n4128 | n4163 ;
  assign n4165 = ~x215 & n4164 ;
  assign n4166 = n4131 | n4165 ;
  assign n4167 = x299 & n4166 ;
  assign n4168 = n4154 | n4167 ;
  assign n4169 = x39 & n4168 ;
  assign n4170 = x38 | n4169 ;
  assign n4171 = n4150 | n4170 ;
  assign n4172 = n4155 | n4157 ;
  assign n4173 = ~x216 & n4172 ;
  assign n4174 = n4108 | n4173 ;
  assign n4175 = ~x221 & n4174 ;
  assign n4176 = n4128 | n4175 ;
  assign n4177 = ~x215 & n4176 ;
  assign n4178 = n4131 | n4177 ;
  assign n4179 = x299 & n4178 ;
  assign n4180 = n4154 | n4179 ;
  assign n4181 = x38 & ~n4180 ;
  assign n4182 = x100 | n4181 ;
  assign n4183 = n4171 & ~n4182 ;
  assign n4184 = n1925 | n4154 ;
  assign n4185 = x152 | x166 ;
  assign n4186 = ( ~x879 & n2155 ) | ( ~x879 & n4185 ) | ( n2155 & n4185 ) ;
  assign n4187 = ( x879 & ~n2153 ) | ( x879 & n4185 ) | ( ~n2153 & n4185 ) ;
  assign n4188 = ~n4186 & n4187 ;
  assign n4189 = ~n2155 & n4115 ;
  assign n4190 = ( x161 & n4188 ) | ( x161 & ~n4189 ) | ( n4188 & ~n4189 ) ;
  assign n4191 = ~x228 & n4190 ;
  assign n4192 = n4155 | n4191 ;
  assign n4193 = ~x216 & n4192 ;
  assign n4194 = n4108 | n4193 ;
  assign n4195 = ~x221 & n4194 ;
  assign n4196 = n4128 | n4195 ;
  assign n4197 = ~x215 & n4196 ;
  assign n4198 = n4132 & ~n4197 ;
  assign n4199 = ( x299 & n4184 ) | ( x299 & ~n4198 ) | ( n4184 & ~n4198 ) ;
  assign n4200 = ( x100 & n2364 ) | ( x100 & n4180 ) | ( n2364 & n4180 ) ;
  assign n4201 = n4199 & n4200 ;
  assign n4202 = n4183 | n4201 ;
  assign n4203 = ~x87 & n4202 ;
  assign n4204 = n1976 & ~n4180 ;
  assign n4205 = n1976 | n4168 ;
  assign n4206 = ~n4204 & n4205 ;
  assign n4207 = ( x75 & n1998 ) | ( x75 & n4206 ) | ( n1998 & n4206 ) ;
  assign n4208 = n4203 | n4207 ;
  assign n4209 = x75 & ~n4180 ;
  assign n4210 = x92 | n4209 ;
  assign n4211 = n4208 & ~n4210 ;
  assign n4212 = ( x92 & ~n1998 ) | ( x92 & n4180 ) | ( ~n1998 & n4180 ) ;
  assign n4213 = ( x92 & n1998 ) | ( x92 & n4206 ) | ( n1998 & n4206 ) ;
  assign n4214 = n4212 & n4213 ;
  assign n4215 = n2030 | n4214 ;
  assign n4216 = n4211 | n4215 ;
  assign n4217 = n2030 & ~n4180 ;
  assign n4218 = x55 | n4217 ;
  assign n4219 = n4216 & ~n4218 ;
  assign n4220 = ( x55 & ~n2033 ) | ( x55 & n4178 ) | ( ~n2033 & n4178 ) ;
  assign n4221 = ( x55 & n2033 ) | ( x55 & n4166 ) | ( n2033 & n4166 ) ;
  assign n4222 = n4220 & n4221 ;
  assign n4223 = x56 | n4222 ;
  assign n4224 = n4219 | n4223 ;
  assign n4225 = ( ~x56 & n2045 ) | ( ~x56 & n4178 ) | ( n2045 & n4178 ) ;
  assign n4226 = ( x56 & n2045 ) | ( x56 & ~n4166 ) | ( n2045 & ~n4166 ) ;
  assign n4227 = ~n4225 & n4226 ;
  assign n4228 = x62 | n4227 ;
  assign n4229 = n4224 & ~n4228 ;
  assign n4230 = ( x62 & ~n2193 ) | ( x62 & n4178 ) | ( ~n2193 & n4178 ) ;
  assign n4231 = ( x62 & n2193 ) | ( x62 & n4166 ) | ( n2193 & n4166 ) ;
  assign n4232 = n4230 & n4231 ;
  assign n4233 = n2057 | n4232 ;
  assign n4234 = n4229 | n4233 ;
  assign n4235 = n2057 & ~n4178 ;
  assign n4236 = x244 | n4235 ;
  assign n4237 = n4234 & ~n4236 ;
  assign n4238 = x161 | n2138 ;
  assign n4239 = x879 & n4238 ;
  assign n4240 = n4117 & ~n4118 ;
  assign n4241 = x228 | n4240 ;
  assign n4242 = n4239 | n4241 ;
  assign n4243 = ~n4114 & n4242 ;
  assign n4244 = n4108 | n4243 ;
  assign n4245 = ~x221 & n4244 ;
  assign n4246 = n4128 | n4245 ;
  assign n4247 = ~x215 & n4246 ;
  assign n4248 = n4132 & ~n4247 ;
  assign n4249 = n3926 | n4144 ;
  assign n4250 = ~x223 & n4249 ;
  assign n4251 = n4135 | n4250 ;
  assign n4252 = ~x39 & n4251 ;
  assign n4253 = ~n4248 & n4252 ;
  assign n4254 = n2205 | n4155 ;
  assign n4255 = n4159 | n4254 ;
  assign n4256 = ~x216 & n4255 ;
  assign n4257 = n4108 | n4256 ;
  assign n4258 = ~x221 & n4257 ;
  assign n4259 = n4128 | n4258 ;
  assign n4260 = ~x215 & n4259 ;
  assign n4261 = n4131 | n4260 ;
  assign n4262 = x299 & n4261 ;
  assign n4263 = n4152 | n4262 ;
  assign n4264 = x39 & n4263 ;
  assign n4265 = x38 | n4264 ;
  assign n4266 = n4253 | n4265 ;
  assign n4267 = n2206 | n4178 ;
  assign n4268 = x299 & n4267 ;
  assign n4269 = n4152 | n4268 ;
  assign n4270 = x38 & ~n4269 ;
  assign n4271 = x100 | n4270 ;
  assign n4272 = n4266 & ~n4271 ;
  assign n4273 = n1925 | n4152 ;
  assign n4274 = n4191 | n4254 ;
  assign n4275 = ~x216 & n4274 ;
  assign n4276 = n4108 | n4275 ;
  assign n4277 = ~x221 & n4276 ;
  assign n4278 = n4128 | n4277 ;
  assign n4279 = ~x215 & n4278 ;
  assign n4280 = n4132 & ~n4279 ;
  assign n4281 = ( x299 & n4273 ) | ( x299 & ~n4280 ) | ( n4273 & ~n4280 ) ;
  assign n4282 = ( x100 & n2364 ) | ( x100 & n4269 ) | ( n2364 & n4269 ) ;
  assign n4283 = n4281 & n4282 ;
  assign n4284 = n4272 | n4283 ;
  assign n4285 = ~x87 & n4284 ;
  assign n4286 = n1976 & ~n4269 ;
  assign n4287 = n1976 | n4263 ;
  assign n4288 = ~n4286 & n4287 ;
  assign n4289 = ( x75 & n1998 ) | ( x75 & n4288 ) | ( n1998 & n4288 ) ;
  assign n4290 = n4285 | n4289 ;
  assign n4291 = x75 & ~n4269 ;
  assign n4292 = x92 | n4291 ;
  assign n4293 = n4290 & ~n4292 ;
  assign n4294 = ( x92 & ~n1998 ) | ( x92 & n4269 ) | ( ~n1998 & n4269 ) ;
  assign n4295 = ( x92 & n1998 ) | ( x92 & n4288 ) | ( n1998 & n4288 ) ;
  assign n4296 = n4294 & n4295 ;
  assign n4297 = n2030 | n4296 ;
  assign n4298 = n4293 | n4297 ;
  assign n4299 = n2030 & ~n4269 ;
  assign n4300 = x55 | n4299 ;
  assign n4301 = n4298 & ~n4300 ;
  assign n4302 = ( x55 & ~n2033 ) | ( x55 & n4267 ) | ( ~n2033 & n4267 ) ;
  assign n4303 = ( x55 & n2033 ) | ( x55 & n4261 ) | ( n2033 & n4261 ) ;
  assign n4304 = n4302 & n4303 ;
  assign n4305 = x56 | n4304 ;
  assign n4306 = n4301 | n4305 ;
  assign n4307 = ( ~x56 & n2045 ) | ( ~x56 & n4267 ) | ( n2045 & n4267 ) ;
  assign n4308 = ( x56 & n2045 ) | ( x56 & ~n4261 ) | ( n2045 & ~n4261 ) ;
  assign n4309 = ~n4307 & n4308 ;
  assign n4310 = x62 | n4309 ;
  assign n4311 = n4306 & ~n4310 ;
  assign n4312 = ( x62 & ~n2193 ) | ( x62 & n4267 ) | ( ~n2193 & n4267 ) ;
  assign n4313 = ( x62 & n2193 ) | ( x62 & n4261 ) | ( n2193 & n4261 ) ;
  assign n4314 = n4312 & n4313 ;
  assign n4315 = n2057 | n4314 ;
  assign n4316 = n4311 | n4315 ;
  assign n4317 = n2057 & ~n4267 ;
  assign n4318 = x244 & ~n4317 ;
  assign n4319 = n4316 & n4318 ;
  assign n4320 = n4237 | n4319 ;
  assign n4321 = x833 & ~x930 ;
  assign n4322 = ~x216 & x221 ;
  assign n4323 = n4321 & n4322 ;
  assign n4324 = x216 & x278 ;
  assign n4325 = x221 | n4324 ;
  assign n4326 = ~x105 & x152 ;
  assign n4327 = x228 & ~n4326 ;
  assign n4328 = x846 | n2227 ;
  assign n4329 = x105 & n4328 ;
  assign n4330 = n4327 & ~n4329 ;
  assign n4331 = x216 | n4330 ;
  assign n4332 = ~x152 & x846 ;
  assign n4333 = ~n2138 & n4332 ;
  assign n4334 = ( ~x152 & x846 ) | ( ~x152 & n2230 ) | ( x846 & n2230 ) ;
  assign n4335 = ( x152 & x846 ) | ( x152 & ~n2239 ) | ( x846 & ~n2239 ) ;
  assign n4336 = n4334 | n4335 ;
  assign n4337 = ~n4333 & n4336 ;
  assign n4338 = x228 | n4337 ;
  assign n4339 = ~n4331 & n4338 ;
  assign n4340 = n4325 | n4339 ;
  assign n4341 = ~n4323 & n4340 ;
  assign n4342 = x221 & ~n1205 ;
  assign n4343 = ~x215 & x299 ;
  assign n4344 = ~n4342 & n4343 ;
  assign n4345 = n4341 & n4344 ;
  assign n4346 = x222 & ~x224 ;
  assign n4347 = n4321 & n4346 ;
  assign n4348 = x224 & x278 ;
  assign n4349 = x222 | n4348 ;
  assign n4350 = ~x224 & n4328 ;
  assign n4351 = n4349 | n4350 ;
  assign n4352 = ~n4347 & n4351 ;
  assign n4353 = n1812 | n2213 ;
  assign n4354 = n4352 & ~n4353 ;
  assign n4355 = x39 | n4354 ;
  assign n4356 = n4345 | n4355 ;
  assign n4357 = x846 & ~n1491 ;
  assign n4358 = ~x224 & n4357 ;
  assign n4359 = n4349 | n4358 ;
  assign n4360 = n1813 | n4347 ;
  assign n4361 = n4359 & ~n4360 ;
  assign n4362 = x299 | n4361 ;
  assign n4363 = n2599 | n4362 ;
  assign n4364 = x215 | n4342 ;
  assign n4365 = n4323 | n4364 ;
  assign n4366 = x105 & n4357 ;
  assign n4367 = n4326 | n4366 ;
  assign n4368 = x228 & n4367 ;
  assign n4369 = n2205 | n4368 ;
  assign n4370 = ( ~x152 & x228 ) | ( ~x152 & n1868 ) | ( x228 & n1868 ) ;
  assign n4371 = ( ~x228 & x846 ) | ( ~x228 & n1868 ) | ( x846 & n1868 ) ;
  assign n4372 = ~n4370 & n4371 ;
  assign n4373 = n4369 | n4372 ;
  assign n4374 = ~x216 & n4373 ;
  assign n4375 = n4325 | n4374 ;
  assign n4376 = ~n4365 & n4375 ;
  assign n4377 = x299 & ~n4376 ;
  assign n4378 = n4363 & ~n4377 ;
  assign n4379 = x39 & ~n4378 ;
  assign n4380 = x38 | n4379 ;
  assign n4381 = n4356 & ~n4380 ;
  assign n4382 = x152 & ~x228 ;
  assign n4383 = n4368 | n4382 ;
  assign n4384 = ~x216 & n4383 ;
  assign n4385 = n4325 | n4384 ;
  assign n4386 = ~n4365 & n4385 ;
  assign n4387 = n2206 | n4386 ;
  assign n4388 = x299 & ~n4387 ;
  assign n4389 = n4363 & ~n4388 ;
  assign n4390 = x38 & n4389 ;
  assign n4391 = x100 | n4390 ;
  assign n4392 = n4381 | n4391 ;
  assign n4393 = x846 & ~n2161 ;
  assign n4394 = ( ~x228 & n2156 ) | ( ~x228 & n4393 ) | ( n2156 & n4393 ) ;
  assign n4395 = n4369 | n4394 ;
  assign n4396 = ~x216 & n4395 ;
  assign n4397 = n4325 | n4396 ;
  assign n4398 = ~n4365 & n4397 ;
  assign n4399 = x299 & ~n4398 ;
  assign n4400 = ~n1925 & n4363 ;
  assign n4401 = ~n4399 & n4400 ;
  assign n4402 = ( x100 & n2364 ) | ( x100 & ~n4389 ) | ( n2364 & ~n4389 ) ;
  assign n4403 = ~n4401 & n4402 ;
  assign n4404 = n4392 & ~n4403 ;
  assign n4405 = x87 | n4404 ;
  assign n4406 = n1976 & n4389 ;
  assign n4407 = ~n1976 & n4378 ;
  assign n4408 = n4406 | n4407 ;
  assign n4409 = ( x75 & n1998 ) | ( x75 & ~n4408 ) | ( n1998 & ~n4408 ) ;
  assign n4410 = n4405 & ~n4409 ;
  assign n4411 = x75 & n4389 ;
  assign n4412 = x92 | n4411 ;
  assign n4413 = n4410 | n4412 ;
  assign n4414 = ( ~x92 & n1998 ) | ( ~x92 & n4389 ) | ( n1998 & n4389 ) ;
  assign n4415 = ( x92 & n1998 ) | ( x92 & ~n4408 ) | ( n1998 & ~n4408 ) ;
  assign n4416 = ~n4414 & n4415 ;
  assign n4417 = n2030 | n4416 ;
  assign n4418 = n4413 & ~n4417 ;
  assign n4419 = n2030 & n4389 ;
  assign n4420 = x55 | n4419 ;
  assign n4421 = n4418 | n4420 ;
  assign n4422 = ( ~x55 & n2033 ) | ( ~x55 & n4387 ) | ( n2033 & n4387 ) ;
  assign n4423 = ( x55 & n2033 ) | ( x55 & ~n4376 ) | ( n2033 & ~n4376 ) ;
  assign n4424 = ~n4422 & n4423 ;
  assign n4425 = x56 | n4424 ;
  assign n4426 = n4421 & ~n4425 ;
  assign n4427 = ( x56 & ~n2045 ) | ( x56 & n4387 ) | ( ~n2045 & n4387 ) ;
  assign n4428 = ( x56 & n2045 ) | ( x56 & n4376 ) | ( n2045 & n4376 ) ;
  assign n4429 = n4427 & n4428 ;
  assign n4430 = x62 | n4429 ;
  assign n4431 = n4426 | n4430 ;
  assign n4432 = ( ~x62 & n2193 ) | ( ~x62 & n4387 ) | ( n2193 & n4387 ) ;
  assign n4433 = ( x62 & n2193 ) | ( x62 & ~n4376 ) | ( n2193 & ~n4376 ) ;
  assign n4434 = ~n4432 & n4433 ;
  assign n4435 = n2057 | n4434 ;
  assign n4436 = n4431 & ~n4435 ;
  assign n4437 = n2057 & n4387 ;
  assign n4438 = x242 & ~n4437 ;
  assign n4439 = ~n4436 & n4438 ;
  assign n4440 = x152 & ~x846 ;
  assign n4441 = ~n2138 & n4440 ;
  assign n4442 = x228 | n4441 ;
  assign n4443 = ( x152 & ~x846 ) | ( x152 & n2230 ) | ( ~x846 & n2230 ) ;
  assign n4444 = ( x152 & x846 ) | ( x152 & n2239 ) | ( x846 & n2239 ) ;
  assign n4445 = ~n4443 & n4444 ;
  assign n4446 = n4442 | n4445 ;
  assign n4447 = n2227 & n4327 ;
  assign n4448 = n4331 | n4447 ;
  assign n4449 = n4446 & ~n4448 ;
  assign n4450 = n4325 | n4449 ;
  assign n4451 = ~n4323 & n4450 ;
  assign n4452 = n4344 & n4451 ;
  assign n4453 = ~n2226 & n4358 ;
  assign n4454 = n4349 | n4453 ;
  assign n4455 = n4347 | n4353 ;
  assign n4456 = n4454 & ~n4455 ;
  assign n4457 = x39 | n4456 ;
  assign n4458 = n4452 | n4457 ;
  assign n4459 = n4368 | n4372 ;
  assign n4460 = ~x216 & n4459 ;
  assign n4461 = n4325 | n4460 ;
  assign n4462 = ~n4365 & n4461 ;
  assign n4463 = x299 & ~n4462 ;
  assign n4464 = n4362 & ~n4463 ;
  assign n4465 = x39 & ~n4464 ;
  assign n4466 = x38 | n4465 ;
  assign n4467 = n4458 & ~n4466 ;
  assign n4468 = x299 & ~n4386 ;
  assign n4469 = n4362 & ~n4468 ;
  assign n4470 = x38 & n4469 ;
  assign n4471 = x100 | n4470 ;
  assign n4472 = n4467 | n4471 ;
  assign n4473 = n4368 | n4394 ;
  assign n4474 = ~x216 & n4473 ;
  assign n4475 = n4325 | n4474 ;
  assign n4476 = ~n4365 & n4475 ;
  assign n4477 = x299 & ~n4476 ;
  assign n4478 = ~n1925 & n4362 ;
  assign n4479 = ~n4477 & n4478 ;
  assign n4480 = ( x100 & n2364 ) | ( x100 & ~n4469 ) | ( n2364 & ~n4469 ) ;
  assign n4481 = ~n4479 & n4480 ;
  assign n4482 = n4472 & ~n4481 ;
  assign n4483 = x87 | n4482 ;
  assign n4484 = n1976 & n4469 ;
  assign n4485 = ~n1976 & n4464 ;
  assign n4486 = n4484 | n4485 ;
  assign n4487 = ( x75 & n1998 ) | ( x75 & ~n4486 ) | ( n1998 & ~n4486 ) ;
  assign n4488 = n4483 & ~n4487 ;
  assign n4489 = x75 & n4469 ;
  assign n4490 = x92 | n4489 ;
  assign n4491 = n4488 | n4490 ;
  assign n4492 = ( ~x92 & n1998 ) | ( ~x92 & n4469 ) | ( n1998 & n4469 ) ;
  assign n4493 = ( x92 & n1998 ) | ( x92 & ~n4486 ) | ( n1998 & ~n4486 ) ;
  assign n4494 = ~n4492 & n4493 ;
  assign n4495 = n2030 | n4494 ;
  assign n4496 = n4491 & ~n4495 ;
  assign n4497 = n2030 & n4469 ;
  assign n4498 = x55 | n4497 ;
  assign n4499 = n4496 | n4498 ;
  assign n4500 = ( ~x55 & n2033 ) | ( ~x55 & n4386 ) | ( n2033 & n4386 ) ;
  assign n4501 = ( x55 & n2033 ) | ( x55 & ~n4462 ) | ( n2033 & ~n4462 ) ;
  assign n4502 = ~n4500 & n4501 ;
  assign n4503 = x56 | n4502 ;
  assign n4504 = n4499 & ~n4503 ;
  assign n4505 = ( x56 & ~n2045 ) | ( x56 & n4386 ) | ( ~n2045 & n4386 ) ;
  assign n4506 = ( x56 & n2045 ) | ( x56 & n4462 ) | ( n2045 & n4462 ) ;
  assign n4507 = n4505 & n4506 ;
  assign n4508 = x62 | n4507 ;
  assign n4509 = n4504 | n4508 ;
  assign n4510 = ( ~x62 & n2193 ) | ( ~x62 & n4386 ) | ( n2193 & n4386 ) ;
  assign n4511 = ( x62 & n2193 ) | ( x62 & ~n4462 ) | ( n2193 & ~n4462 ) ;
  assign n4512 = ~n4510 & n4511 ;
  assign n4513 = n2057 | n4512 ;
  assign n4514 = n4509 & ~n4513 ;
  assign n4515 = n2057 & n4386 ;
  assign n4516 = x242 | n4515 ;
  assign n4517 = n4514 | n4516 ;
  assign n4518 = ~n4439 & n4517 ;
  assign n4519 = x1134 | n4518 ;
  assign n4520 = n2213 | n4352 ;
  assign n4521 = ~x39 & n4520 ;
  assign n4522 = ~n4341 & n4343 ;
  assign n4523 = n4521 & ~n4522 ;
  assign n4524 = n1813 | n4363 ;
  assign n4525 = ~x299 & n4524 ;
  assign n4526 = ~n4323 & n4375 ;
  assign n4527 = x215 | n4526 ;
  assign n4528 = x299 & n4527 ;
  assign n4529 = n4525 | n4528 ;
  assign n4530 = x39 & n4529 ;
  assign n4531 = x38 | n4530 ;
  assign n4532 = n4523 | n4531 ;
  assign n4533 = ~n4323 & n4385 ;
  assign n4534 = x215 | n4533 ;
  assign n4535 = n2206 | n4534 ;
  assign n4536 = x299 & n4535 ;
  assign n4537 = n4525 | n4536 ;
  assign n4538 = x38 & ~n4537 ;
  assign n4539 = x100 | n4538 ;
  assign n4540 = n4532 & ~n4539 ;
  assign n4541 = ~n4323 & n4397 ;
  assign n4542 = x215 | n4541 ;
  assign n4543 = x299 & n4542 ;
  assign n4544 = n1925 | n4525 ;
  assign n4545 = n4543 | n4544 ;
  assign n4546 = ( x100 & n2364 ) | ( x100 & n4537 ) | ( n2364 & n4537 ) ;
  assign n4547 = n4545 & n4546 ;
  assign n4548 = n4540 | n4547 ;
  assign n4549 = ~x87 & n4548 ;
  assign n4550 = n1976 & ~n4537 ;
  assign n4551 = n1976 | n4529 ;
  assign n4552 = ~n4550 & n4551 ;
  assign n4553 = ( x75 & n1998 ) | ( x75 & n4552 ) | ( n1998 & n4552 ) ;
  assign n4554 = n4549 | n4553 ;
  assign n4555 = x75 & ~n4537 ;
  assign n4556 = x92 | n4555 ;
  assign n4557 = n4554 & ~n4556 ;
  assign n4558 = ( x92 & ~n1998 ) | ( x92 & n4537 ) | ( ~n1998 & n4537 ) ;
  assign n4559 = ( x92 & n1998 ) | ( x92 & n4552 ) | ( n1998 & n4552 ) ;
  assign n4560 = n4558 & n4559 ;
  assign n4561 = n2030 | n4560 ;
  assign n4562 = n4557 | n4561 ;
  assign n4563 = n2030 & ~n4537 ;
  assign n4564 = x55 | n4563 ;
  assign n4565 = n4562 & ~n4564 ;
  assign n4566 = ( x55 & ~n2033 ) | ( x55 & n4535 ) | ( ~n2033 & n4535 ) ;
  assign n4567 = ( x55 & n2033 ) | ( x55 & n4527 ) | ( n2033 & n4527 ) ;
  assign n4568 = n4566 & n4567 ;
  assign n4569 = x56 | n4568 ;
  assign n4570 = n4565 | n4569 ;
  assign n4571 = ( ~x56 & n2045 ) | ( ~x56 & n4535 ) | ( n2045 & n4535 ) ;
  assign n4572 = ( x56 & n2045 ) | ( x56 & ~n4527 ) | ( n2045 & ~n4527 ) ;
  assign n4573 = ~n4571 & n4572 ;
  assign n4574 = x62 | n4573 ;
  assign n4575 = n4570 & ~n4574 ;
  assign n4576 = ( x62 & ~n2193 ) | ( x62 & n4535 ) | ( ~n2193 & n4535 ) ;
  assign n4577 = ( x62 & n2193 ) | ( x62 & n4527 ) | ( n2193 & n4527 ) ;
  assign n4578 = n4576 & n4577 ;
  assign n4579 = n2057 | n4578 ;
  assign n4580 = n4575 | n4579 ;
  assign n4581 = n2057 & ~n4535 ;
  assign n4582 = x242 & ~n4581 ;
  assign n4583 = n4580 & n4582 ;
  assign n4584 = n4343 & ~n4451 ;
  assign n4585 = n2213 | n4454 ;
  assign n4586 = n4521 & n4585 ;
  assign n4587 = ~n4584 & n4586 ;
  assign n4588 = x223 | n4359 ;
  assign n4589 = n4525 & n4588 ;
  assign n4590 = ~n4323 & n4461 ;
  assign n4591 = x215 | n4590 ;
  assign n4592 = x299 & n4591 ;
  assign n4593 = n4589 | n4592 ;
  assign n4594 = x39 & n4593 ;
  assign n4595 = x38 | n4594 ;
  assign n4596 = n4587 | n4595 ;
  assign n4597 = x299 & n4534 ;
  assign n4598 = n4589 | n4597 ;
  assign n4599 = x38 & ~n4598 ;
  assign n4600 = x100 | n4599 ;
  assign n4601 = n4596 & ~n4600 ;
  assign n4602 = ~n4323 & n4475 ;
  assign n4603 = x215 | n4602 ;
  assign n4604 = x299 & n4603 ;
  assign n4605 = n1925 | n4589 ;
  assign n4606 = n4604 | n4605 ;
  assign n4607 = ( x100 & n2364 ) | ( x100 & n4598 ) | ( n2364 & n4598 ) ;
  assign n4608 = n4606 & n4607 ;
  assign n4609 = n4601 | n4608 ;
  assign n4610 = ~x87 & n4609 ;
  assign n4611 = n1976 & ~n4598 ;
  assign n4612 = n1976 | n4593 ;
  assign n4613 = ~n4611 & n4612 ;
  assign n4614 = ( x75 & n1998 ) | ( x75 & n4613 ) | ( n1998 & n4613 ) ;
  assign n4615 = n4610 | n4614 ;
  assign n4616 = x75 & ~n4598 ;
  assign n4617 = x92 | n4616 ;
  assign n4618 = n4615 & ~n4617 ;
  assign n4619 = ( x92 & ~n1998 ) | ( x92 & n4598 ) | ( ~n1998 & n4598 ) ;
  assign n4620 = ( x92 & n1998 ) | ( x92 & n4613 ) | ( n1998 & n4613 ) ;
  assign n4621 = n4619 & n4620 ;
  assign n4622 = n2030 | n4621 ;
  assign n4623 = n4618 | n4622 ;
  assign n4624 = n2030 & ~n4598 ;
  assign n4625 = x55 | n4624 ;
  assign n4626 = n4623 & ~n4625 ;
  assign n4627 = ( x55 & ~n2033 ) | ( x55 & n4534 ) | ( ~n2033 & n4534 ) ;
  assign n4628 = ( x55 & n2033 ) | ( x55 & n4591 ) | ( n2033 & n4591 ) ;
  assign n4629 = n4627 & n4628 ;
  assign n4630 = x56 | n4629 ;
  assign n4631 = n4626 | n4630 ;
  assign n4632 = ( ~x56 & n2045 ) | ( ~x56 & n4534 ) | ( n2045 & n4534 ) ;
  assign n4633 = ( x56 & n2045 ) | ( x56 & ~n4591 ) | ( n2045 & ~n4591 ) ;
  assign n4634 = ~n4632 & n4633 ;
  assign n4635 = x62 | n4634 ;
  assign n4636 = n4631 & ~n4635 ;
  assign n4637 = ( x62 & ~n2193 ) | ( x62 & n4534 ) | ( ~n2193 & n4534 ) ;
  assign n4638 = ( x62 & n2193 ) | ( x62 & n4591 ) | ( n2193 & n4591 ) ;
  assign n4639 = n4637 & n4638 ;
  assign n4640 = n2057 | n4639 ;
  assign n4641 = n4636 | n4640 ;
  assign n4642 = n2057 & ~n4534 ;
  assign n4643 = x242 | n4642 ;
  assign n4644 = n4641 & ~n4643 ;
  assign n4645 = x1134 & ~n4644 ;
  assign n4646 = ~n4583 & n4645 ;
  assign n4647 = n4519 & ~n4646 ;
  assign n4648 = n1868 | n2059 ;
  assign n4649 = ( x57 & x59 ) | ( x57 & n4648 ) | ( x59 & n4648 ) ;
  assign n4650 = x57 & n4649 ;
  assign n4651 = n1860 | n1976 ;
  assign n4652 = n2044 | n4651 ;
  assign n4653 = x56 & n4652 ;
  assign n4654 = x54 | n2042 ;
  assign n4655 = n4651 | n4654 ;
  assign n4656 = x74 & n4655 ;
  assign n4657 = x55 | n4656 ;
  assign n4658 = x39 | x95 ;
  assign n4659 = n1494 | n4658 ;
  assign n4660 = n1272 | n4659 ;
  assign n4661 = x38 & n4660 ;
  assign n4662 = x100 | n4661 ;
  assign n4663 = x841 | n1272 ;
  assign n4664 = x93 & n4663 ;
  assign n4665 = x58 & ~n1307 ;
  assign n4666 = x90 | n4665 ;
  assign n4667 = n1326 | n1338 ;
  assign n4668 = n1440 & ~n4667 ;
  assign n4669 = n1345 | n4668 ;
  assign n4670 = ~n1337 & n4669 ;
  assign n4671 = x108 | n4670 ;
  assign n4672 = ~n1334 & n4671 ;
  assign n4673 = x110 | n1731 ;
  assign n4674 = n4672 | n4673 ;
  assign n4675 = n1317 | n1453 ;
  assign n4676 = n4674 & ~n4675 ;
  assign n4677 = x47 | n4676 ;
  assign n4678 = ~n1242 & n1320 ;
  assign n4679 = x47 & ~n4678 ;
  assign n4680 = n1251 | n4679 ;
  assign n4681 = n4677 & ~n4680 ;
  assign n4682 = n4666 | n4681 ;
  assign n4683 = ~n1649 & n4682 ;
  assign n4684 = ( x93 & ~n4664 ) | ( x93 & n4683 ) | ( ~n4664 & n4683 ) ;
  assign n4685 = x35 | n4684 ;
  assign n4686 = ~n1594 & n4685 ;
  assign n4687 = ( x51 & ~n1644 ) | ( x51 & n4686 ) | ( ~n1644 & n4686 ) ;
  assign n4688 = ~n1465 & n4687 ;
  assign n4689 = n1539 | n4688 ;
  assign n4690 = ~n1302 & n4689 ;
  assign n4691 = n1300 | n4690 ;
  assign n4692 = x198 | x299 ;
  assign n4693 = ~x210 & x299 ;
  assign n4694 = n4692 & ~n4693 ;
  assign n4695 = x35 | n1295 ;
  assign n4696 = x40 | n4695 ;
  assign n4697 = n1604 & ~n4696 ;
  assign n4698 = x32 & ~n4697 ;
  assign n4699 = n4694 | n4698 ;
  assign n4700 = ~n2129 & n4694 ;
  assign n4701 = n4699 & ~n4700 ;
  assign n4702 = n4691 & ~n4701 ;
  assign n4703 = x95 | n4702 ;
  assign n4704 = ~n1496 & n4703 ;
  assign n4705 = x39 | n4704 ;
  assign n4706 = x603 & ~x642 ;
  assign n4707 = x614 | x616 ;
  assign n4708 = n4706 & ~n4707 ;
  assign n4709 = ~x662 & x680 ;
  assign n4710 = x661 | x681 ;
  assign n4711 = n4709 & ~n4710 ;
  assign n4712 = n4708 | n4711 ;
  assign n4713 = x332 | x468 ;
  assign n4714 = n4712 & n4713 ;
  assign n4715 = x970 | x972 ;
  assign n4716 = x975 | x978 ;
  assign n4717 = n4715 | n4716 ;
  assign n4718 = x907 | x947 ;
  assign n4719 = x960 | x963 ;
  assign n4720 = n4718 | n4719 ;
  assign n4721 = n4717 | n4720 ;
  assign n4722 = ~n4713 & n4721 ;
  assign n4723 = n4714 | n4722 ;
  assign n4724 = x835 & x950 ;
  assign n4725 = x252 | x1001 ;
  assign n4726 = ~x979 & n4725 ;
  assign n4727 = x835 & x984 ;
  assign n4728 = x287 | n4727 ;
  assign n4729 = n4726 & ~n4728 ;
  assign n4730 = n4724 & n4729 ;
  assign n4731 = n1292 & n4730 ;
  assign n4732 = x216 & x221 ;
  assign n4733 = n4731 & n4732 ;
  assign n4734 = n4723 & n4733 ;
  assign n4735 = n1868 | n4734 ;
  assign n4736 = ~x215 & n4735 ;
  assign n4737 = x299 & ~n4736 ;
  assign n4738 = n1860 | n4713 ;
  assign n4739 = n4712 & ~n4738 ;
  assign n4740 = x1092 & n4730 ;
  assign n4741 = x1093 & ~n1288 ;
  assign n4742 = x829 & ~n4741 ;
  assign n4743 = x1091 & n4741 ;
  assign n4744 = ( x824 & n4742 ) | ( x824 & ~n4743 ) | ( n4742 & ~n4743 ) ;
  assign n4745 = n4740 & n4744 ;
  assign n4746 = n4714 & ~n4745 ;
  assign n4747 = ( n1868 & n4712 ) | ( n1868 & ~n4746 ) | ( n4712 & ~n4746 ) ;
  assign n4748 = ~n4739 & n4747 ;
  assign n4749 = ( x215 & n4721 ) | ( x215 & n4748 ) | ( n4721 & n4748 ) ;
  assign n4750 = ~n4708 & n4713 ;
  assign n4751 = ~n4711 & n4750 ;
  assign n4752 = n4745 & ~n4751 ;
  assign n4753 = n1868 | n4752 ;
  assign n4754 = ( x215 & ~n4721 ) | ( x215 & n4753 ) | ( ~n4721 & n4753 ) ;
  assign n4755 = n4749 & n4754 ;
  assign n4756 = n4737 & ~n4755 ;
  assign n4757 = x39 & x299 ;
  assign n4758 = x969 | x971 ;
  assign n4759 = x974 | x977 ;
  assign n4760 = n4758 | n4759 ;
  assign n4761 = x587 | x602 ;
  assign n4762 = x961 | x967 ;
  assign n4763 = n4761 | n4762 ;
  assign n4764 = n4760 | n4763 ;
  assign n4765 = ~n4713 & n4764 ;
  assign n4766 = n4714 | n4765 ;
  assign n4767 = x222 & x224 ;
  assign n4768 = n4731 & n4767 ;
  assign n4769 = n4766 & n4768 ;
  assign n4770 = n1868 | n4769 ;
  assign n4771 = ~x223 & n4770 ;
  assign n4772 = ( x223 & n4753 ) | ( x223 & ~n4764 ) | ( n4753 & ~n4764 ) ;
  assign n4773 = ( x223 & n4748 ) | ( x223 & n4764 ) | ( n4748 & n4764 ) ;
  assign n4774 = n4772 & n4773 ;
  assign n4775 = n4771 | n4774 ;
  assign n4776 = ( x39 & n4757 ) | ( x39 & n4775 ) | ( n4757 & n4775 ) ;
  assign n4777 = ~n4756 & n4776 ;
  assign n4778 = n4705 & ~n4777 ;
  assign n4779 = x38 | n4778 ;
  assign n4780 = ~n4662 & n4779 ;
  assign n4781 = ~x142 & n1834 ;
  assign n4782 = ~x299 & n4781 ;
  assign n4783 = x299 & n1615 ;
  assign n4784 = n4782 | n4783 ;
  assign n4785 = n2153 & ~n4784 ;
  assign n4786 = x41 | x99 ;
  assign n4787 = x101 | n4786 ;
  assign n4788 = x42 | x43 ;
  assign n4789 = x52 | n4788 ;
  assign n4790 = x113 | x116 ;
  assign n4791 = x114 | x115 ;
  assign n4792 = n4790 | n4791 ;
  assign n4793 = n4789 | n4792 ;
  assign n4794 = n4787 | n4793 ;
  assign n4795 = x44 | n4794 ;
  assign n4796 = ~x683 & n4795 ;
  assign n4797 = x129 & x250 ;
  assign n4798 = x824 | x829 ;
  assign n4799 = n1692 & n4798 ;
  assign n4800 = ~x1093 & n4799 ;
  assign n4801 = x250 | n4800 ;
  assign n4802 = ~n4797 & n4801 ;
  assign n4803 = n4796 | n4802 ;
  assign n4804 = n4784 & n4795 ;
  assign n4805 = ~n4803 & n4804 ;
  assign n4806 = n4785 | n4805 ;
  assign n4807 = ~x38 & x100 ;
  assign n4808 = x39 | n1462 ;
  assign n4809 = n1865 | n4808 ;
  assign n4810 = n1272 | n4809 ;
  assign n4811 = n4807 & ~n4810 ;
  assign n4812 = x87 | n4811 ;
  assign n4813 = ( x87 & ~n4806 ) | ( x87 & n4812 ) | ( ~n4806 & n4812 ) ;
  assign n4814 = n4780 | n4813 ;
  assign n4815 = x87 & n4651 ;
  assign n4816 = x75 | n4815 ;
  assign n4817 = x54 | x92 ;
  assign n4818 = n4816 | n4817 ;
  assign n4819 = n4814 & ~n4818 ;
  assign n4820 = x74 | n4819 ;
  assign n4821 = ~n4657 & n4820 ;
  assign n4822 = x56 | n4821 ;
  assign n4823 = ~n4653 & n4822 ;
  assign n4824 = x62 | n4823 ;
  assign n4825 = n2192 | n4651 ;
  assign n4826 = x62 & n4825 ;
  assign n4827 = x59 | n4826 ;
  assign n4828 = x57 | n4827 ;
  assign n4829 = n4824 & ~n4828 ;
  assign n4830 = ( x57 & ~n4650 ) | ( x57 & n4829 ) | ( ~n4650 & n4829 ) ;
  assign n4831 = x55 | x59 ;
  assign n4832 = n2058 | n4831 ;
  assign n4833 = ~x228 & n4832 ;
  assign n4834 = x57 & ~n4833 ;
  assign n4835 = ~n4711 & n4713 ;
  assign n4836 = x907 | n4713 ;
  assign n4837 = ~n4835 & n4836 ;
  assign n4838 = ~x228 & n2033 ;
  assign n4839 = x30 & x228 ;
  assign n4840 = n2082 & ~n4839 ;
  assign n4841 = n4838 | n4840 ;
  assign n4842 = n4837 & ~n4841 ;
  assign n4843 = n4834 & n4842 ;
  assign n4844 = x602 | n4713 ;
  assign n4845 = ~n4835 & n4844 ;
  assign n4846 = x93 & ~n1603 ;
  assign n4847 = x35 | n4846 ;
  assign n4848 = x91 | x314 ;
  assign n4849 = x67 & ~n1352 ;
  assign n4850 = n1362 | n4849 ;
  assign n4851 = x85 & n1379 ;
  assign n4852 = n1229 | n4851 ;
  assign n4853 = ~n1381 & n4852 ;
  assign n4854 = n1230 | n4853 ;
  assign n4855 = n1365 | n1390 ;
  assign n4856 = n4854 & ~n4855 ;
  assign n4857 = ~n1227 & n4856 ;
  assign n4858 = n1396 | n4857 ;
  assign n4859 = ( ~n1393 & n4850 ) | ( ~n1393 & n4858 ) | ( n4850 & n4858 ) ;
  assign n4860 = ~n1361 & n4859 ;
  assign n4861 = x71 | n4860 ;
  assign n4862 = x64 | n1236 ;
  assign n4863 = n1355 | n4862 ;
  assign n4864 = n4861 & ~n4863 ;
  assign n4865 = x81 | n4864 ;
  assign n4866 = n1406 & ~n4863 ;
  assign n4867 = n4865 | n4866 ;
  assign n4868 = x81 & n1242 ;
  assign n4869 = x102 | n4868 ;
  assign n4870 = n1339 | n4869 ;
  assign n4871 = n4867 & ~n4870 ;
  assign n4872 = n1350 | n4871 ;
  assign n4873 = ~n1443 & n4872 ;
  assign n4874 = n1582 | n4873 ;
  assign n4875 = ~n1584 & n4874 ;
  assign n4876 = x86 | n4875 ;
  assign n4877 = x46 | n1213 ;
  assign n4878 = n1347 | n4877 ;
  assign n4879 = n4876 & ~n4878 ;
  assign n4880 = n1731 | n4879 ;
  assign n4881 = ~n1454 & n4880 ;
  assign n4882 = n4848 | n4881 ;
  assign n4883 = x91 & n1313 ;
  assign n4884 = x58 | n4883 ;
  assign n4885 = ~x91 & x314 ;
  assign n4886 = n4865 & ~n4870 ;
  assign n4887 = n1350 | n4886 ;
  assign n4888 = ~n1443 & n4887 ;
  assign n4889 = n1582 | n4888 ;
  assign n4890 = ~n1584 & n4889 ;
  assign n4891 = x86 | n4890 ;
  assign n4892 = ~n4878 & n4891 ;
  assign n4893 = n1731 | n4892 ;
  assign n4894 = ~n1454 & n4893 ;
  assign n4895 = n4885 & ~n4894 ;
  assign n4896 = n4884 | n4895 ;
  assign n4897 = n4882 & ~n4896 ;
  assign n4898 = x90 | n4897 ;
  assign n4899 = ~n1649 & n4898 ;
  assign n4900 = ( x93 & ~n4847 ) | ( x93 & n4899 ) | ( ~n4847 & n4899 ) ;
  assign n4901 = x70 | n4900 ;
  assign n4902 = ~n1281 & n4901 ;
  assign n4903 = x72 | n4902 ;
  assign n4904 = x95 | n1492 ;
  assign n4905 = n1301 | n4904 ;
  assign n4906 = n4903 & ~n4905 ;
  assign n4907 = n1536 | n4906 ;
  assign n4908 = x93 | x841 ;
  assign n4909 = n1526 | n4908 ;
  assign n4910 = n1682 | n4909 ;
  assign n4911 = n1272 | n4910 ;
  assign n4912 = x32 & ~n4911 ;
  assign n4913 = ~x95 & n4912 ;
  assign n4914 = ~x198 & n4913 ;
  assign n4915 = n4907 | n4914 ;
  assign n4916 = ~x228 & n4915 ;
  assign n4917 = n4839 | n4916 ;
  assign n4918 = n4845 & n4917 ;
  assign n4919 = x299 | n4918 ;
  assign n4920 = x145 & x180 ;
  assign n4921 = x181 & x182 ;
  assign n4922 = n4920 & n4921 ;
  assign n4923 = ~x299 & n4922 ;
  assign n4924 = n4919 & ~n4923 ;
  assign n4925 = n4839 & n4845 ;
  assign n4926 = n4713 & n4915 ;
  assign n4927 = x47 | n1250 ;
  assign n4928 = n1730 | n4879 ;
  assign n4929 = ~n4927 & n4928 ;
  assign n4930 = n4848 | n4929 ;
  assign n4931 = n1730 | n4892 ;
  assign n4932 = ~n4927 & n4931 ;
  assign n4933 = n4885 & ~n4932 ;
  assign n4934 = n4884 | n4933 ;
  assign n4935 = n4930 & ~n4934 ;
  assign n4936 = x90 | n4935 ;
  assign n4937 = ~n1649 & n4936 ;
  assign n4938 = ( x93 & ~n4847 ) | ( x93 & n4937 ) | ( ~n4847 & n4937 ) ;
  assign n4939 = x70 | n4938 ;
  assign n4940 = ~n1281 & n4939 ;
  assign n4941 = x72 | n4940 ;
  assign n4942 = ~n4905 & n4941 ;
  assign n4943 = n1536 | n4942 ;
  assign n4944 = n4914 | n4943 ;
  assign n4945 = ~n4713 & n4944 ;
  assign n4946 = n4926 | n4945 ;
  assign n4947 = ~x228 & n4845 ;
  assign n4948 = n4946 & n4947 ;
  assign n4949 = n4925 | n4948 ;
  assign n4950 = n4922 & n4949 ;
  assign n4951 = n4924 | n4950 ;
  assign n4952 = n4837 & n4839 ;
  assign n4953 = x299 & ~n4952 ;
  assign n4954 = x158 & x159 ;
  assign n4955 = x160 & x197 ;
  assign n4956 = n4954 & n4955 ;
  assign n4957 = ~x210 & n4913 ;
  assign n4958 = n4907 | n4957 ;
  assign n4959 = n4713 & n4958 ;
  assign n4960 = n4943 | n4957 ;
  assign n4961 = ~n4713 & n4960 ;
  assign n4962 = n4959 | n4961 ;
  assign n4963 = n4837 & n4962 ;
  assign n4964 = ( x228 & n4956 ) | ( x228 & ~n4963 ) | ( n4956 & ~n4963 ) ;
  assign n4965 = n4837 & n4958 ;
  assign n4966 = ( ~x228 & n4956 ) | ( ~x228 & n4965 ) | ( n4956 & n4965 ) ;
  assign n4967 = ~n4964 & n4966 ;
  assign n4968 = n4953 & ~n4967 ;
  assign n4969 = x232 & ~n4968 ;
  assign n4970 = n4951 & n4969 ;
  assign n4971 = ~x228 & n4965 ;
  assign n4972 = n4953 & ~n4971 ;
  assign n4973 = x232 | n4972 ;
  assign n4974 = n4919 & ~n4973 ;
  assign n4975 = n4970 | n4974 ;
  assign n4976 = ~x39 & n4975 ;
  assign n4977 = n4726 & ~n4727 ;
  assign n4978 = x835 & n4977 ;
  assign n4979 = x287 | n1462 ;
  assign n4980 = n1865 | n4979 ;
  assign n4981 = n1272 | n4980 ;
  assign n4982 = n4978 & ~n4981 ;
  assign n4983 = x824 & x1093 ;
  assign n4984 = n1692 & n4983 ;
  assign n4985 = n4982 & n4984 ;
  assign n4986 = x829 | n1287 ;
  assign n4987 = x1091 & n4986 ;
  assign n4988 = n4985 & ~n4987 ;
  assign n4989 = x222 & ~x223 ;
  assign n4990 = ( x224 & n4988 ) | ( x224 & n4989 ) | ( n4988 & n4989 ) ;
  assign n4991 = ~x1091 & n4985 ;
  assign n4992 = x1091 & n1287 ;
  assign n4993 = n4984 & ~n4992 ;
  assign n4994 = n1292 | n4993 ;
  assign n4995 = x1091 & n4994 ;
  assign n4996 = n4982 & n4995 ;
  assign n4997 = n4991 | n4996 ;
  assign n4998 = ( ~x224 & n4989 ) | ( ~x224 & n4997 ) | ( n4989 & n4997 ) ;
  assign n4999 = n4990 & n4998 ;
  assign n5000 = ~x228 & n4999 ;
  assign n5001 = n4839 | n5000 ;
  assign n5002 = ~x299 & n4845 ;
  assign n5003 = n5001 & n5002 ;
  assign n5004 = ( x39 & x299 ) | ( x39 & n5003 ) | ( x299 & n5003 ) ;
  assign n5005 = ~x215 & x221 ;
  assign n5006 = x216 & n4997 ;
  assign n5007 = ~x216 & n4988 ;
  assign n5008 = n5006 | n5007 ;
  assign n5009 = ~x228 & n5008 ;
  assign n5010 = n4839 | n5009 ;
  assign n5011 = n5005 & n5010 ;
  assign n5012 = n4839 | n5011 ;
  assign n5013 = x299 & n4837 ;
  assign n5014 = n5012 & n5013 ;
  assign n5015 = ( ~x299 & n5004 ) | ( ~x299 & n5014 ) | ( n5004 & n5014 ) ;
  assign n5016 = x38 | n5015 ;
  assign n5017 = n4976 | n5016 ;
  assign n5018 = n5002 | n5013 ;
  assign n5019 = x39 | n4840 ;
  assign n5020 = n5018 & ~n5019 ;
  assign n5021 = n4839 & n5018 ;
  assign n5022 = x38 & ~n5021 ;
  assign n5023 = ~n5020 & n5022 ;
  assign n5024 = n5017 & ~n5023 ;
  assign n5025 = x100 | n5024 ;
  assign n5026 = n1868 | n4802 ;
  assign n5027 = x683 & n4795 ;
  assign n5028 = ~n5026 & n5027 ;
  assign n5029 = ~n4835 & n5028 ;
  assign n5030 = n4781 & n5029 ;
  assign n5031 = x252 & ~n4781 ;
  assign n5032 = x252 & ~n4738 ;
  assign n5033 = ~n4711 & n5032 ;
  assign n5034 = x252 & ~n1868 ;
  assign n5035 = n4711 & n5034 ;
  assign n5036 = n5033 | n5035 ;
  assign n5037 = n5031 & n5036 ;
  assign n5038 = n5030 | n5037 ;
  assign n5039 = ~x228 & n4844 ;
  assign n5040 = n5038 & n5039 ;
  assign n5041 = x299 | n4925 ;
  assign n5042 = n5040 | n5041 ;
  assign n5043 = ~x228 & n4836 ;
  assign n5044 = ( ~n1615 & n5029 ) | ( ~n1615 & n5043 ) | ( n5029 & n5043 ) ;
  assign n5045 = ( n1615 & n5036 ) | ( n1615 & n5043 ) | ( n5036 & n5043 ) ;
  assign n5046 = n5044 & n5045 ;
  assign n5047 = n4953 & ~n5046 ;
  assign n5048 = n1925 | n5047 ;
  assign n5049 = n5042 & ~n5048 ;
  assign n5050 = n1925 & n5021 ;
  assign n5051 = n5049 | n5050 ;
  assign n5052 = ( x87 & n1924 ) | ( x87 & ~n5051 ) | ( n1924 & ~n5051 ) ;
  assign n5053 = n5025 & ~n5052 ;
  assign n5054 = ( x75 & n1998 ) | ( x75 & n5021 ) | ( n1998 & n5021 ) ;
  assign n5055 = n5053 | n5054 ;
  assign n5056 = n1984 & n5021 ;
  assign n5057 = ~n2007 & n5020 ;
  assign n5058 = n5056 | n5057 ;
  assign n5059 = x75 & ~n5058 ;
  assign n5060 = x92 | n5059 ;
  assign n5061 = n5055 & ~n5060 ;
  assign n5062 = ( x75 & x92 ) | ( x75 & n5058 ) | ( x92 & n5058 ) ;
  assign n5063 = ( ~x75 & x92 ) | ( ~x75 & n5021 ) | ( x92 & n5021 ) ;
  assign n5064 = n5062 & n5063 ;
  assign n5065 = x54 | n5064 ;
  assign n5066 = n5061 | n5065 ;
  assign n5067 = n2004 | n5058 ;
  assign n5068 = n2004 & ~n5021 ;
  assign n5069 = n5067 & ~n5068 ;
  assign n5070 = x54 & ~n5069 ;
  assign n5071 = x74 | n5070 ;
  assign n5072 = n5066 & ~n5071 ;
  assign n5073 = x55 | x74 ;
  assign n5074 = x54 | n5067 ;
  assign n5075 = x54 | n2004 ;
  assign n5076 = ~n5021 & n5075 ;
  assign n5077 = n5074 & ~n5076 ;
  assign n5078 = ( x55 & n5073 ) | ( x55 & n5077 ) | ( n5073 & n5077 ) ;
  assign n5079 = n5072 | n5078 ;
  assign n5080 = x55 & ~n4842 ;
  assign n5081 = n2058 | n5080 ;
  assign n5082 = n5079 & ~n5081 ;
  assign n5083 = n2058 & n4952 ;
  assign n5084 = x59 | n5083 ;
  assign n5085 = n5082 | n5084 ;
  assign n5086 = x55 | n2058 ;
  assign n5087 = ~x228 & n5086 ;
  assign n5088 = n4842 & ~n5087 ;
  assign n5089 = x59 & ~n5088 ;
  assign n5090 = x57 | n5089 ;
  assign n5091 = n5085 & ~n5090 ;
  assign n5092 = n4843 | n5091 ;
  assign n5093 = x947 | n4713 ;
  assign n5094 = ~n4750 & n5093 ;
  assign n5095 = ~n4841 & n5094 ;
  assign n5096 = n4834 & n5095 ;
  assign n5097 = n4839 & n5094 ;
  assign n5098 = x299 & ~n5097 ;
  assign n5099 = n4962 & n5094 ;
  assign n5100 = ( x228 & n4956 ) | ( x228 & ~n5099 ) | ( n4956 & ~n5099 ) ;
  assign n5101 = n4958 & n5094 ;
  assign n5102 = ( ~x228 & n4956 ) | ( ~x228 & n5101 ) | ( n4956 & n5101 ) ;
  assign n5103 = ~n5100 & n5102 ;
  assign n5104 = n5098 & ~n5103 ;
  assign n5105 = x232 & ~n5104 ;
  assign n5106 = x587 | n4713 ;
  assign n5107 = ~n4750 & n5106 ;
  assign n5108 = n4839 & n5107 ;
  assign n5109 = ~x228 & n5107 ;
  assign n5110 = n4946 & n5109 ;
  assign n5111 = n5108 | n5110 ;
  assign n5112 = ( x299 & n4922 ) | ( x299 & n5111 ) | ( n4922 & n5111 ) ;
  assign n5113 = n4917 & n5107 ;
  assign n5114 = ( x299 & ~n4922 ) | ( x299 & n5113 ) | ( ~n4922 & n5113 ) ;
  assign n5115 = n5112 | n5114 ;
  assign n5116 = n5105 & n5115 ;
  assign n5117 = x299 | n5113 ;
  assign n5118 = ~x228 & n5101 ;
  assign n5119 = n5098 & ~n5118 ;
  assign n5120 = x232 | n5119 ;
  assign n5121 = n5117 & ~n5120 ;
  assign n5122 = n5116 | n5121 ;
  assign n5123 = ~x39 & n5122 ;
  assign n5124 = x299 & n5005 ;
  assign n5125 = n5098 | n5124 ;
  assign n5126 = n5011 & n5094 ;
  assign n5127 = n5125 & ~n5126 ;
  assign n5128 = n5001 & n5107 ;
  assign n5129 = x299 | n5128 ;
  assign n5130 = ~n5127 & n5129 ;
  assign n5131 = ( x38 & n1925 ) | ( x38 & n5130 ) | ( n1925 & n5130 ) ;
  assign n5132 = n5123 | n5131 ;
  assign n5133 = x299 & ~n5094 ;
  assign n5134 = x299 | n5107 ;
  assign n5135 = ~n5133 & n5134 ;
  assign n5136 = ~n5019 & n5135 ;
  assign n5137 = n4839 & n5135 ;
  assign n5138 = x38 & ~n5137 ;
  assign n5139 = ~n5136 & n5138 ;
  assign n5140 = n5132 & ~n5139 ;
  assign n5141 = x100 | n5140 ;
  assign n5142 = x228 | n1834 ;
  assign n5143 = n4708 | n5032 ;
  assign n5144 = n4708 & ~n5034 ;
  assign n5145 = n5143 & ~n5144 ;
  assign n5146 = n5106 & n5145 ;
  assign n5147 = n5142 | n5146 ;
  assign n5148 = ~n5108 & n5142 ;
  assign n5149 = ~n4750 & n5028 ;
  assign n5150 = n4708 & n4713 ;
  assign n5151 = x587 | n5150 ;
  assign n5152 = ~x228 & n5151 ;
  assign n5153 = ( x142 & n5149 ) | ( x142 & n5152 ) | ( n5149 & n5152 ) ;
  assign n5154 = ( ~x142 & n5145 ) | ( ~x142 & n5152 ) | ( n5145 & n5152 ) ;
  assign n5155 = n5153 & n5154 ;
  assign n5156 = n5148 & ~n5155 ;
  assign n5157 = n5147 & ~n5156 ;
  assign n5158 = x299 | n5157 ;
  assign n5159 = n1615 & n5093 ;
  assign n5160 = n5149 & n5159 ;
  assign n5161 = x947 | n5150 ;
  assign n5162 = ~n1615 & n5161 ;
  assign n5163 = n5145 & n5162 ;
  assign n5164 = n5160 | n5163 ;
  assign n5165 = ~x228 & n5164 ;
  assign n5166 = n5098 & ~n5165 ;
  assign n5167 = n1925 | n5166 ;
  assign n5168 = n5158 & ~n5167 ;
  assign n5169 = n1925 & n5137 ;
  assign n5170 = n5168 | n5169 ;
  assign n5171 = ( x87 & n1924 ) | ( x87 & ~n5170 ) | ( n1924 & ~n5170 ) ;
  assign n5172 = n5141 & ~n5171 ;
  assign n5173 = ( x75 & n1998 ) | ( x75 & n5137 ) | ( n1998 & n5137 ) ;
  assign n5174 = n5172 | n5173 ;
  assign n5175 = n1984 & n5137 ;
  assign n5176 = ~n2007 & n5136 ;
  assign n5177 = n5175 | n5176 ;
  assign n5178 = x75 & ~n5177 ;
  assign n5179 = x92 | n5178 ;
  assign n5180 = n5174 & ~n5179 ;
  assign n5181 = ( x75 & x92 ) | ( x75 & n5177 ) | ( x92 & n5177 ) ;
  assign n5182 = ( ~x75 & x92 ) | ( ~x75 & n5137 ) | ( x92 & n5137 ) ;
  assign n5183 = n5181 & n5182 ;
  assign n5184 = x54 | n5183 ;
  assign n5185 = n5180 | n5184 ;
  assign n5186 = n2004 | n5177 ;
  assign n5187 = n2004 & ~n5137 ;
  assign n5188 = n5186 & ~n5187 ;
  assign n5189 = x54 & ~n5188 ;
  assign n5190 = x74 | n5189 ;
  assign n5191 = n5185 & ~n5190 ;
  assign n5192 = x54 | n5186 ;
  assign n5193 = n5075 & ~n5137 ;
  assign n5194 = n5192 & ~n5193 ;
  assign n5195 = ( x55 & n5073 ) | ( x55 & n5194 ) | ( n5073 & n5194 ) ;
  assign n5196 = n5191 | n5195 ;
  assign n5197 = x55 & ~n5095 ;
  assign n5198 = n2058 | n5197 ;
  assign n5199 = n5196 & ~n5198 ;
  assign n5200 = n2058 & n5097 ;
  assign n5201 = x59 | n5200 ;
  assign n5202 = n5199 | n5201 ;
  assign n5203 = ~n5087 & n5095 ;
  assign n5204 = x59 & ~n5203 ;
  assign n5205 = x57 | n5204 ;
  assign n5206 = n5202 & ~n5205 ;
  assign n5207 = n5096 | n5206 ;
  assign n5208 = x30 & ~n4713 ;
  assign n5209 = x228 & n5208 ;
  assign n5210 = x970 & n5209 ;
  assign n5211 = ~x228 & x970 ;
  assign n5212 = ~n4738 & n5211 ;
  assign n5213 = ~n2033 & n5212 ;
  assign n5214 = ~n4832 & n5213 ;
  assign n5215 = n5210 | n5214 ;
  assign n5216 = x57 & n5215 ;
  assign n5217 = x299 & ~n5210 ;
  assign n5218 = ~n4713 & n4958 ;
  assign n5219 = n5211 & n5218 ;
  assign n5220 = n5217 & ~n5219 ;
  assign n5221 = x299 & n4954 ;
  assign n5222 = n5220 | n5221 ;
  assign n5223 = n4955 & ~n4961 ;
  assign n5224 = n4955 | n4958 ;
  assign n5225 = ~n5223 & n5224 ;
  assign n5226 = ~n4713 & n5225 ;
  assign n5227 = n5211 & n5226 ;
  assign n5228 = n5210 | n5227 ;
  assign n5229 = n4954 & n5228 ;
  assign n5230 = n5222 & ~n5229 ;
  assign n5231 = ~n4713 & n4917 ;
  assign n5232 = n4922 | n5231 ;
  assign n5233 = ~x228 & n4945 ;
  assign n5234 = n4915 & ~n4922 ;
  assign n5235 = n5209 | n5234 ;
  assign n5236 = n5233 | n5235 ;
  assign n5237 = n5232 & n5236 ;
  assign n5238 = ~x299 & x967 ;
  assign n5239 = n5237 & n5238 ;
  assign n5240 = ( x232 & x299 ) | ( x232 & n5239 ) | ( x299 & n5239 ) ;
  assign n5241 = ~n5230 & n5240 ;
  assign n5242 = x232 | n5220 ;
  assign n5243 = n5231 & n5238 ;
  assign n5244 = ( x299 & ~n5242 ) | ( x299 & n5243 ) | ( ~n5242 & n5243 ) ;
  assign n5245 = n5241 | n5244 ;
  assign n5246 = ~x39 & n5245 ;
  assign n5247 = x299 & x970 ;
  assign n5248 = n5005 & n5008 ;
  assign n5249 = ~n4713 & n5248 ;
  assign n5250 = x228 | n5249 ;
  assign n5251 = n5247 & n5250 ;
  assign n5252 = ~n4713 & n4999 ;
  assign n5253 = x228 | n5252 ;
  assign n5254 = n5238 & n5253 ;
  assign n5255 = n5251 | n5254 ;
  assign n5256 = x228 & ~n5208 ;
  assign n5257 = x39 & ~n5256 ;
  assign n5258 = n5255 & n5257 ;
  assign n5259 = x38 | n5258 ;
  assign n5260 = n5246 | n5259 ;
  assign n5261 = ~n5212 & n5217 ;
  assign n5262 = x39 | n5261 ;
  assign n5263 = ~x228 & n4738 ;
  assign n5264 = n5256 | n5263 ;
  assign n5265 = n5238 & ~n5264 ;
  assign n5266 = ( x299 & ~n5262 ) | ( x299 & n5265 ) | ( ~n5262 & n5265 ) ;
  assign n5267 = n5238 | n5247 ;
  assign n5268 = n5209 & n5267 ;
  assign n5269 = ( x38 & n1919 ) | ( x38 & ~n5268 ) | ( n1919 & ~n5268 ) ;
  assign n5270 = ~n5266 & n5269 ;
  assign n5271 = n5260 & ~n5270 ;
  assign n5272 = x100 | n5271 ;
  assign n5273 = n1925 & n5268 ;
  assign n5274 = ~n4713 & n5028 ;
  assign n5275 = ( x228 & n1615 ) | ( x228 & ~n5274 ) | ( n1615 & ~n5274 ) ;
  assign n5276 = ( ~x228 & n1615 ) | ( ~x228 & n5032 ) | ( n1615 & n5032 ) ;
  assign n5277 = ~n5275 & n5276 ;
  assign n5278 = x970 & n5277 ;
  assign n5279 = n5217 & ~n5278 ;
  assign n5280 = n1925 | n5279 ;
  assign n5281 = ( x228 & n4781 ) | ( x228 & n5274 ) | ( n4781 & n5274 ) ;
  assign n5282 = ( x228 & ~n4781 ) | ( x228 & n5032 ) | ( ~n4781 & n5032 ) ;
  assign n5283 = n5281 | n5282 ;
  assign n5284 = ~n5256 & n5283 ;
  assign n5285 = n5238 & n5284 ;
  assign n5286 = ( x299 & ~n5280 ) | ( x299 & n5285 ) | ( ~n5280 & n5285 ) ;
  assign n5287 = n5273 | n5286 ;
  assign n5288 = ( x87 & n1924 ) | ( x87 & ~n5287 ) | ( n1924 & ~n5287 ) ;
  assign n5289 = n5272 & ~n5288 ;
  assign n5290 = x87 & n5268 ;
  assign n5291 = x75 | n5290 ;
  assign n5292 = n5289 | n5291 ;
  assign n5293 = n1984 & n5268 ;
  assign n5294 = ~n2007 & n5266 ;
  assign n5295 = n5293 | n5294 ;
  assign n5296 = x75 & ~n5295 ;
  assign n5297 = x92 | n5296 ;
  assign n5298 = n5292 & ~n5297 ;
  assign n5299 = ( x75 & x92 ) | ( x75 & n5295 ) | ( x92 & n5295 ) ;
  assign n5300 = ( ~x75 & x92 ) | ( ~x75 & n5268 ) | ( x92 & n5268 ) ;
  assign n5301 = n5299 & n5300 ;
  assign n5302 = x54 | n5301 ;
  assign n5303 = n5298 | n5302 ;
  assign n5304 = n2004 | n5295 ;
  assign n5305 = n2004 & ~n5268 ;
  assign n5306 = n5304 & ~n5305 ;
  assign n5307 = x54 & ~n5306 ;
  assign n5308 = x74 | n5307 ;
  assign n5309 = n5303 & ~n5308 ;
  assign n5310 = x54 | n5304 ;
  assign n5311 = n5075 & ~n5268 ;
  assign n5312 = n5310 & ~n5311 ;
  assign n5313 = ( x55 & n5073 ) | ( x55 & n5312 ) | ( n5073 & n5312 ) ;
  assign n5314 = n5309 | n5313 ;
  assign n5315 = x55 & ~n5210 ;
  assign n5316 = ~n5213 & n5315 ;
  assign n5317 = n2058 | n5316 ;
  assign n5318 = n5314 & ~n5317 ;
  assign n5319 = n2058 & n5210 ;
  assign n5320 = x59 | n5319 ;
  assign n5321 = n5318 | n5320 ;
  assign n5322 = ~n5086 & n5213 ;
  assign n5323 = n5210 | n5322 ;
  assign n5324 = ( x57 & n2057 ) | ( x57 & ~n5323 ) | ( n2057 & ~n5323 ) ;
  assign n5325 = n5321 & ~n5324 ;
  assign n5326 = n5216 | n5325 ;
  assign n5327 = x972 & n5209 ;
  assign n5328 = ~x228 & x972 ;
  assign n5329 = ~n4738 & n5328 ;
  assign n5330 = ~n2033 & n5329 ;
  assign n5331 = ~n4832 & n5330 ;
  assign n5332 = n5327 | n5331 ;
  assign n5333 = x57 & n5332 ;
  assign n5334 = x299 & ~n5327 ;
  assign n5335 = n5218 & n5328 ;
  assign n5336 = n5334 & ~n5335 ;
  assign n5337 = n5221 | n5336 ;
  assign n5338 = n5226 & n5328 ;
  assign n5339 = n5327 | n5338 ;
  assign n5340 = n4954 & n5339 ;
  assign n5341 = n5337 & ~n5340 ;
  assign n5342 = ~x299 & x961 ;
  assign n5343 = n5237 & n5342 ;
  assign n5344 = ( x232 & x299 ) | ( x232 & n5343 ) | ( x299 & n5343 ) ;
  assign n5345 = ~n5341 & n5344 ;
  assign n5346 = x232 | n5336 ;
  assign n5347 = n5231 & n5342 ;
  assign n5348 = ( x299 & ~n5346 ) | ( x299 & n5347 ) | ( ~n5346 & n5347 ) ;
  assign n5349 = n5345 | n5348 ;
  assign n5350 = ~x39 & n5349 ;
  assign n5351 = n5253 & n5342 ;
  assign n5352 = x299 & x972 ;
  assign n5353 = n5250 & n5352 ;
  assign n5354 = n5351 | n5353 ;
  assign n5355 = n5257 & n5354 ;
  assign n5356 = x38 | n5355 ;
  assign n5357 = n5350 | n5356 ;
  assign n5358 = ~n5329 & n5334 ;
  assign n5359 = x39 | n5358 ;
  assign n5360 = ~n5264 & n5342 ;
  assign n5361 = ( x299 & ~n5359 ) | ( x299 & n5360 ) | ( ~n5359 & n5360 ) ;
  assign n5362 = n5342 | n5352 ;
  assign n5363 = n5209 & n5362 ;
  assign n5364 = ( x38 & n1919 ) | ( x38 & ~n5363 ) | ( n1919 & ~n5363 ) ;
  assign n5365 = ~n5361 & n5364 ;
  assign n5366 = n5357 & ~n5365 ;
  assign n5367 = x100 | n5366 ;
  assign n5368 = n1925 & n5363 ;
  assign n5369 = x972 & n5277 ;
  assign n5370 = n5334 & ~n5369 ;
  assign n5371 = n1925 | n5370 ;
  assign n5372 = n5284 & n5342 ;
  assign n5373 = ( x299 & ~n5371 ) | ( x299 & n5372 ) | ( ~n5371 & n5372 ) ;
  assign n5374 = n5368 | n5373 ;
  assign n5375 = ( x87 & n1924 ) | ( x87 & ~n5374 ) | ( n1924 & ~n5374 ) ;
  assign n5376 = n5367 & ~n5375 ;
  assign n5377 = x87 & n5363 ;
  assign n5378 = x75 | n5377 ;
  assign n5379 = n5376 | n5378 ;
  assign n5380 = n1984 & n5363 ;
  assign n5381 = ~n2007 & n5361 ;
  assign n5382 = n5380 | n5381 ;
  assign n5383 = x75 & ~n5382 ;
  assign n5384 = x92 | n5383 ;
  assign n5385 = n5379 & ~n5384 ;
  assign n5386 = ( x75 & x92 ) | ( x75 & n5382 ) | ( x92 & n5382 ) ;
  assign n5387 = ( ~x75 & x92 ) | ( ~x75 & n5363 ) | ( x92 & n5363 ) ;
  assign n5388 = n5386 & n5387 ;
  assign n5389 = x54 | n5388 ;
  assign n5390 = n5385 | n5389 ;
  assign n5391 = n2004 | n5382 ;
  assign n5392 = n2004 & ~n5363 ;
  assign n5393 = n5391 & ~n5392 ;
  assign n5394 = x54 & ~n5393 ;
  assign n5395 = x74 | n5394 ;
  assign n5396 = n5390 & ~n5395 ;
  assign n5397 = x54 | n5391 ;
  assign n5398 = n5075 & ~n5363 ;
  assign n5399 = n5397 & ~n5398 ;
  assign n5400 = ( x55 & n5073 ) | ( x55 & n5399 ) | ( n5073 & n5399 ) ;
  assign n5401 = n5396 | n5400 ;
  assign n5402 = x55 & ~n5327 ;
  assign n5403 = ~n5330 & n5402 ;
  assign n5404 = n2058 | n5403 ;
  assign n5405 = n5401 & ~n5404 ;
  assign n5406 = n2058 & n5327 ;
  assign n5407 = x59 | n5406 ;
  assign n5408 = n5405 | n5407 ;
  assign n5409 = ~n5086 & n5330 ;
  assign n5410 = n5327 | n5409 ;
  assign n5411 = ( x57 & n2057 ) | ( x57 & ~n5410 ) | ( n2057 & ~n5410 ) ;
  assign n5412 = n5408 & ~n5411 ;
  assign n5413 = n5333 | n5412 ;
  assign n5414 = x960 & n5209 ;
  assign n5415 = ~x228 & x960 ;
  assign n5416 = ~n4738 & n5415 ;
  assign n5417 = ~n2033 & n5416 ;
  assign n5418 = ~n4832 & n5417 ;
  assign n5419 = n5414 | n5418 ;
  assign n5420 = x57 & n5419 ;
  assign n5421 = x299 & ~n5414 ;
  assign n5422 = n5218 & n5415 ;
  assign n5423 = n5421 & ~n5422 ;
  assign n5424 = n5221 | n5423 ;
  assign n5425 = n5226 & n5415 ;
  assign n5426 = n5414 | n5425 ;
  assign n5427 = n4954 & n5426 ;
  assign n5428 = n5424 & ~n5427 ;
  assign n5429 = ~x299 & x977 ;
  assign n5430 = n5237 & n5429 ;
  assign n5431 = ( x232 & x299 ) | ( x232 & n5430 ) | ( x299 & n5430 ) ;
  assign n5432 = ~n5428 & n5431 ;
  assign n5433 = x232 | n5423 ;
  assign n5434 = n5231 & n5429 ;
  assign n5435 = ( x299 & ~n5433 ) | ( x299 & n5434 ) | ( ~n5433 & n5434 ) ;
  assign n5436 = n5432 | n5435 ;
  assign n5437 = ~x39 & n5436 ;
  assign n5438 = n5253 & n5429 ;
  assign n5439 = x299 & x960 ;
  assign n5440 = n5250 & n5439 ;
  assign n5441 = n5438 | n5440 ;
  assign n5442 = n5257 & n5441 ;
  assign n5443 = x38 | n5442 ;
  assign n5444 = n5437 | n5443 ;
  assign n5445 = ~n5416 & n5421 ;
  assign n5446 = x39 | n5445 ;
  assign n5447 = ~n5264 & n5429 ;
  assign n5448 = ( x299 & ~n5446 ) | ( x299 & n5447 ) | ( ~n5446 & n5447 ) ;
  assign n5449 = n5429 | n5439 ;
  assign n5450 = n5209 & n5449 ;
  assign n5451 = ( x38 & n1919 ) | ( x38 & ~n5450 ) | ( n1919 & ~n5450 ) ;
  assign n5452 = ~n5448 & n5451 ;
  assign n5453 = n5444 & ~n5452 ;
  assign n5454 = x100 | n5453 ;
  assign n5455 = n1925 & n5450 ;
  assign n5456 = x960 & n5277 ;
  assign n5457 = n5421 & ~n5456 ;
  assign n5458 = n1925 | n5457 ;
  assign n5459 = n5284 & n5429 ;
  assign n5460 = ( x299 & ~n5458 ) | ( x299 & n5459 ) | ( ~n5458 & n5459 ) ;
  assign n5461 = n5455 | n5460 ;
  assign n5462 = ( x87 & n1924 ) | ( x87 & ~n5461 ) | ( n1924 & ~n5461 ) ;
  assign n5463 = n5454 & ~n5462 ;
  assign n5464 = x87 & n5450 ;
  assign n5465 = x75 | n5464 ;
  assign n5466 = n5463 | n5465 ;
  assign n5467 = n1984 & n5450 ;
  assign n5468 = ~n2007 & n5448 ;
  assign n5469 = n5467 | n5468 ;
  assign n5470 = x75 & ~n5469 ;
  assign n5471 = x92 | n5470 ;
  assign n5472 = n5466 & ~n5471 ;
  assign n5473 = ( x75 & x92 ) | ( x75 & n5469 ) | ( x92 & n5469 ) ;
  assign n5474 = ( ~x75 & x92 ) | ( ~x75 & n5450 ) | ( x92 & n5450 ) ;
  assign n5475 = n5473 & n5474 ;
  assign n5476 = x54 | n5475 ;
  assign n5477 = n5472 | n5476 ;
  assign n5478 = n2004 | n5469 ;
  assign n5479 = n2004 & ~n5450 ;
  assign n5480 = n5478 & ~n5479 ;
  assign n5481 = x54 & ~n5480 ;
  assign n5482 = x74 | n5481 ;
  assign n5483 = n5477 & ~n5482 ;
  assign n5484 = x54 | n5478 ;
  assign n5485 = n5075 & ~n5450 ;
  assign n5486 = n5484 & ~n5485 ;
  assign n5487 = ( x55 & n5073 ) | ( x55 & n5486 ) | ( n5073 & n5486 ) ;
  assign n5488 = n5483 | n5487 ;
  assign n5489 = x55 & ~n5414 ;
  assign n5490 = ~n5417 & n5489 ;
  assign n5491 = n2058 | n5490 ;
  assign n5492 = n5488 & ~n5491 ;
  assign n5493 = n2058 & n5414 ;
  assign n5494 = x59 | n5493 ;
  assign n5495 = n5492 | n5494 ;
  assign n5496 = ~n5086 & n5417 ;
  assign n5497 = n5414 | n5496 ;
  assign n5498 = ( x57 & n2057 ) | ( x57 & ~n5497 ) | ( n2057 & ~n5497 ) ;
  assign n5499 = n5495 & ~n5498 ;
  assign n5500 = n5420 | n5499 ;
  assign n5501 = x963 & n5209 ;
  assign n5502 = ~x228 & x963 ;
  assign n5503 = ~n4738 & n5502 ;
  assign n5504 = ~n2033 & n5503 ;
  assign n5505 = ~n4832 & n5504 ;
  assign n5506 = n5501 | n5505 ;
  assign n5507 = x57 & n5506 ;
  assign n5508 = x299 & ~n5501 ;
  assign n5509 = n5218 & n5502 ;
  assign n5510 = n5508 & ~n5509 ;
  assign n5511 = n5221 | n5510 ;
  assign n5512 = n5226 & n5502 ;
  assign n5513 = n5501 | n5512 ;
  assign n5514 = n4954 & n5513 ;
  assign n5515 = n5511 & ~n5514 ;
  assign n5516 = ~x299 & x969 ;
  assign n5517 = n5237 & n5516 ;
  assign n5518 = ( x232 & x299 ) | ( x232 & n5517 ) | ( x299 & n5517 ) ;
  assign n5519 = ~n5515 & n5518 ;
  assign n5520 = x232 | n5510 ;
  assign n5521 = n5231 & n5516 ;
  assign n5522 = ( x299 & ~n5520 ) | ( x299 & n5521 ) | ( ~n5520 & n5521 ) ;
  assign n5523 = n5519 | n5522 ;
  assign n5524 = ~x39 & n5523 ;
  assign n5525 = n5253 & n5516 ;
  assign n5526 = x299 & x963 ;
  assign n5527 = n5250 & n5526 ;
  assign n5528 = n5525 | n5527 ;
  assign n5529 = n5257 & n5528 ;
  assign n5530 = x38 | n5529 ;
  assign n5531 = n5524 | n5530 ;
  assign n5532 = ~n5503 & n5508 ;
  assign n5533 = x39 | n5532 ;
  assign n5534 = ~n5264 & n5516 ;
  assign n5535 = ( x299 & ~n5533 ) | ( x299 & n5534 ) | ( ~n5533 & n5534 ) ;
  assign n5536 = n5516 | n5526 ;
  assign n5537 = n5209 & n5536 ;
  assign n5538 = ( x38 & n1919 ) | ( x38 & ~n5537 ) | ( n1919 & ~n5537 ) ;
  assign n5539 = ~n5535 & n5538 ;
  assign n5540 = n5531 & ~n5539 ;
  assign n5541 = x100 | n5540 ;
  assign n5542 = n1925 & n5537 ;
  assign n5543 = x963 & n5277 ;
  assign n5544 = n5508 & ~n5543 ;
  assign n5545 = n1925 | n5544 ;
  assign n5546 = n5284 & n5516 ;
  assign n5547 = ( x299 & ~n5545 ) | ( x299 & n5546 ) | ( ~n5545 & n5546 ) ;
  assign n5548 = n5542 | n5547 ;
  assign n5549 = ( x87 & n1924 ) | ( x87 & ~n5548 ) | ( n1924 & ~n5548 ) ;
  assign n5550 = n5541 & ~n5549 ;
  assign n5551 = x87 & n5537 ;
  assign n5552 = x75 | n5551 ;
  assign n5553 = n5550 | n5552 ;
  assign n5554 = n1984 & n5537 ;
  assign n5555 = ~n2007 & n5535 ;
  assign n5556 = n5554 | n5555 ;
  assign n5557 = x75 & ~n5556 ;
  assign n5558 = x92 | n5557 ;
  assign n5559 = n5553 & ~n5558 ;
  assign n5560 = ( x75 & x92 ) | ( x75 & n5556 ) | ( x92 & n5556 ) ;
  assign n5561 = ( ~x75 & x92 ) | ( ~x75 & n5537 ) | ( x92 & n5537 ) ;
  assign n5562 = n5560 & n5561 ;
  assign n5563 = x54 | n5562 ;
  assign n5564 = n5559 | n5563 ;
  assign n5565 = n2004 | n5556 ;
  assign n5566 = n2004 & ~n5537 ;
  assign n5567 = n5565 & ~n5566 ;
  assign n5568 = x54 & ~n5567 ;
  assign n5569 = x74 | n5568 ;
  assign n5570 = n5564 & ~n5569 ;
  assign n5571 = x54 | n5565 ;
  assign n5572 = n5075 & ~n5537 ;
  assign n5573 = n5571 & ~n5572 ;
  assign n5574 = ( x55 & n5073 ) | ( x55 & n5573 ) | ( n5073 & n5573 ) ;
  assign n5575 = n5570 | n5574 ;
  assign n5576 = x55 & ~n5501 ;
  assign n5577 = ~n5504 & n5576 ;
  assign n5578 = n2058 | n5577 ;
  assign n5579 = n5575 & ~n5578 ;
  assign n5580 = n2058 & n5501 ;
  assign n5581 = x59 | n5580 ;
  assign n5582 = n5579 | n5581 ;
  assign n5583 = ~n5086 & n5504 ;
  assign n5584 = n5501 | n5583 ;
  assign n5585 = ( x57 & n2057 ) | ( x57 & ~n5584 ) | ( n2057 & ~n5584 ) ;
  assign n5586 = n5582 & ~n5585 ;
  assign n5587 = n5507 | n5586 ;
  assign n5588 = x975 & n5209 ;
  assign n5589 = ~x228 & x975 ;
  assign n5590 = ~n4738 & n5589 ;
  assign n5591 = ~n2033 & n5590 ;
  assign n5592 = ~n4832 & n5591 ;
  assign n5593 = n5588 | n5592 ;
  assign n5594 = x57 & n5593 ;
  assign n5595 = x299 & ~n5588 ;
  assign n5596 = n5218 & n5589 ;
  assign n5597 = n5595 & ~n5596 ;
  assign n5598 = n5221 | n5597 ;
  assign n5599 = n5226 & n5589 ;
  assign n5600 = n5588 | n5599 ;
  assign n5601 = n4954 & n5600 ;
  assign n5602 = n5598 & ~n5601 ;
  assign n5603 = ~x299 & x971 ;
  assign n5604 = n5237 & n5603 ;
  assign n5605 = ( x232 & x299 ) | ( x232 & n5604 ) | ( x299 & n5604 ) ;
  assign n5606 = ~n5602 & n5605 ;
  assign n5607 = x232 | n5597 ;
  assign n5608 = n5231 & n5603 ;
  assign n5609 = ( x299 & ~n5607 ) | ( x299 & n5608 ) | ( ~n5607 & n5608 ) ;
  assign n5610 = n5606 | n5609 ;
  assign n5611 = ~x39 & n5610 ;
  assign n5612 = n5253 & n5603 ;
  assign n5613 = x299 & x975 ;
  assign n5614 = n5250 & n5613 ;
  assign n5615 = n5612 | n5614 ;
  assign n5616 = n5257 & n5615 ;
  assign n5617 = x38 | n5616 ;
  assign n5618 = n5611 | n5617 ;
  assign n5619 = ~n5590 & n5595 ;
  assign n5620 = x39 | n5619 ;
  assign n5621 = ~n5264 & n5603 ;
  assign n5622 = ( x299 & ~n5620 ) | ( x299 & n5621 ) | ( ~n5620 & n5621 ) ;
  assign n5623 = n5603 | n5613 ;
  assign n5624 = n5209 & n5623 ;
  assign n5625 = ( x38 & n1919 ) | ( x38 & ~n5624 ) | ( n1919 & ~n5624 ) ;
  assign n5626 = ~n5622 & n5625 ;
  assign n5627 = n5618 & ~n5626 ;
  assign n5628 = x100 | n5627 ;
  assign n5629 = n1925 & n5624 ;
  assign n5630 = x975 & n5277 ;
  assign n5631 = n5595 & ~n5630 ;
  assign n5632 = n1925 | n5631 ;
  assign n5633 = n5284 & n5603 ;
  assign n5634 = ( x299 & ~n5632 ) | ( x299 & n5633 ) | ( ~n5632 & n5633 ) ;
  assign n5635 = n5629 | n5634 ;
  assign n5636 = ( x87 & n1924 ) | ( x87 & ~n5635 ) | ( n1924 & ~n5635 ) ;
  assign n5637 = n5628 & ~n5636 ;
  assign n5638 = x87 & n5624 ;
  assign n5639 = x75 | n5638 ;
  assign n5640 = n5637 | n5639 ;
  assign n5641 = n1984 & n5624 ;
  assign n5642 = ~n2007 & n5622 ;
  assign n5643 = n5641 | n5642 ;
  assign n5644 = x75 & ~n5643 ;
  assign n5645 = x92 | n5644 ;
  assign n5646 = n5640 & ~n5645 ;
  assign n5647 = ( x75 & x92 ) | ( x75 & n5643 ) | ( x92 & n5643 ) ;
  assign n5648 = ( ~x75 & x92 ) | ( ~x75 & n5624 ) | ( x92 & n5624 ) ;
  assign n5649 = n5647 & n5648 ;
  assign n5650 = x54 | n5649 ;
  assign n5651 = n5646 | n5650 ;
  assign n5652 = n2004 | n5643 ;
  assign n5653 = n2004 & ~n5624 ;
  assign n5654 = n5652 & ~n5653 ;
  assign n5655 = x54 & ~n5654 ;
  assign n5656 = x74 | n5655 ;
  assign n5657 = n5651 & ~n5656 ;
  assign n5658 = x54 | n5652 ;
  assign n5659 = n5075 & ~n5624 ;
  assign n5660 = n5658 & ~n5659 ;
  assign n5661 = ( x55 & n5073 ) | ( x55 & n5660 ) | ( n5073 & n5660 ) ;
  assign n5662 = n5657 | n5661 ;
  assign n5663 = x55 & ~n5588 ;
  assign n5664 = ~n5591 & n5663 ;
  assign n5665 = n2058 | n5664 ;
  assign n5666 = n5662 & ~n5665 ;
  assign n5667 = n2058 & n5588 ;
  assign n5668 = x59 | n5667 ;
  assign n5669 = n5666 | n5668 ;
  assign n5670 = ~n5086 & n5591 ;
  assign n5671 = n5588 | n5670 ;
  assign n5672 = ( x57 & n2057 ) | ( x57 & ~n5671 ) | ( n2057 & ~n5671 ) ;
  assign n5673 = n5669 & ~n5672 ;
  assign n5674 = n5594 | n5673 ;
  assign n5675 = x978 & n5209 ;
  assign n5676 = ~x228 & x978 ;
  assign n5677 = ~n2033 & n5676 ;
  assign n5678 = ~n4738 & n5677 ;
  assign n5679 = ~n4832 & n5678 ;
  assign n5680 = n5675 | n5679 ;
  assign n5681 = x57 & n5680 ;
  assign n5682 = x299 & ~n5675 ;
  assign n5683 = n5218 & n5676 ;
  assign n5684 = n5682 & ~n5683 ;
  assign n5685 = n5221 | n5684 ;
  assign n5686 = n5226 & n5676 ;
  assign n5687 = n5675 | n5686 ;
  assign n5688 = n4954 & n5687 ;
  assign n5689 = n5685 & ~n5688 ;
  assign n5690 = ~x299 & x974 ;
  assign n5691 = n5237 & n5690 ;
  assign n5692 = ( x232 & x299 ) | ( x232 & n5691 ) | ( x299 & n5691 ) ;
  assign n5693 = ~n5689 & n5692 ;
  assign n5694 = x232 | n5684 ;
  assign n5695 = n5231 & n5690 ;
  assign n5696 = ( x299 & ~n5694 ) | ( x299 & n5695 ) | ( ~n5694 & n5695 ) ;
  assign n5697 = n5693 | n5696 ;
  assign n5698 = ~x39 & n5697 ;
  assign n5699 = n5253 & n5690 ;
  assign n5700 = x299 & x978 ;
  assign n5701 = n5250 & n5700 ;
  assign n5702 = n5699 | n5701 ;
  assign n5703 = n5257 & n5702 ;
  assign n5704 = x38 | n5703 ;
  assign n5705 = n5698 | n5704 ;
  assign n5706 = n5690 | n5700 ;
  assign n5707 = n5209 & n5706 ;
  assign n5708 = ( ~x38 & x39 ) | ( ~x38 & n5707 ) | ( x39 & n5707 ) ;
  assign n5709 = ~n5264 & n5706 ;
  assign n5710 = ( x38 & x39 ) | ( x38 & ~n5709 ) | ( x39 & ~n5709 ) ;
  assign n5711 = ~n5708 & n5710 ;
  assign n5712 = n5705 & ~n5711 ;
  assign n5713 = x100 | n5712 ;
  assign n5714 = n1925 & n5707 ;
  assign n5715 = x978 & n5277 ;
  assign n5716 = n5682 & ~n5715 ;
  assign n5717 = n1925 | n5716 ;
  assign n5718 = n5284 & n5690 ;
  assign n5719 = ( x299 & ~n5717 ) | ( x299 & n5718 ) | ( ~n5717 & n5718 ) ;
  assign n5720 = n5714 | n5719 ;
  assign n5721 = ( x87 & n1924 ) | ( x87 & ~n5720 ) | ( n1924 & ~n5720 ) ;
  assign n5722 = n5713 & ~n5721 ;
  assign n5723 = ( x75 & n1998 ) | ( x75 & n5707 ) | ( n1998 & n5707 ) ;
  assign n5724 = n5722 | n5723 ;
  assign n5725 = ~x228 & n1984 ;
  assign n5726 = n5709 & ~n5725 ;
  assign n5727 = x75 & ~n5726 ;
  assign n5728 = x92 | n5727 ;
  assign n5729 = n5724 & ~n5728 ;
  assign n5730 = ( x75 & x92 ) | ( x75 & n5726 ) | ( x92 & n5726 ) ;
  assign n5731 = ( ~x75 & x92 ) | ( ~x75 & n5707 ) | ( x92 & n5707 ) ;
  assign n5732 = n5730 & n5731 ;
  assign n5733 = x54 | n5732 ;
  assign n5734 = n5729 | n5733 ;
  assign n5735 = n2004 | n5726 ;
  assign n5736 = n2004 & ~n5707 ;
  assign n5737 = n5735 & ~n5736 ;
  assign n5738 = x54 & ~n5737 ;
  assign n5739 = x74 | n5738 ;
  assign n5740 = n5734 & ~n5739 ;
  assign n5741 = x54 | n5735 ;
  assign n5742 = n5075 & ~n5707 ;
  assign n5743 = n5741 & ~n5742 ;
  assign n5744 = ( x55 & n5073 ) | ( x55 & n5743 ) | ( n5073 & n5743 ) ;
  assign n5745 = n5740 | n5744 ;
  assign n5746 = x55 & ~n5675 ;
  assign n5747 = ~n5678 & n5746 ;
  assign n5748 = n2058 | n5747 ;
  assign n5749 = n5745 & ~n5748 ;
  assign n5750 = n2058 & n5675 ;
  assign n5751 = x59 | n5750 ;
  assign n5752 = n5749 | n5751 ;
  assign n5753 = ~n5086 & n5678 ;
  assign n5754 = n5675 | n5753 ;
  assign n5755 = ( x57 & n2057 ) | ( x57 & ~n5754 ) | ( n2057 & ~n5754 ) ;
  assign n5756 = n5752 & ~n5755 ;
  assign n5757 = n5681 | n5756 ;
  assign n5758 = n2043 | n4651 ;
  assign n5759 = x55 & n5758 ;
  assign n5760 = x56 | n5759 ;
  assign n5761 = x62 | n5760 ;
  assign n5762 = n2007 | n4810 ;
  assign n5763 = x75 & n5762 ;
  assign n5764 = n1975 | n1998 ;
  assign n5765 = n4810 | n5764 ;
  assign n5766 = x92 & n5765 ;
  assign n5767 = n5763 | n5766 ;
  assign n5768 = x38 | n4810 ;
  assign n5769 = x100 & n5768 ;
  assign n5770 = n4813 | n5769 ;
  assign n5771 = x299 & n4723 ;
  assign n5772 = n5248 & n5771 ;
  assign n5773 = ~x299 & n4766 ;
  assign n5774 = n4999 & n5773 ;
  assign n5775 = x39 & ~n5774 ;
  assign n5776 = ~n5772 & n5775 ;
  assign n5777 = ~n4959 & n5221 ;
  assign n5778 = ~n5225 & n5777 ;
  assign n5779 = n4922 & n4945 ;
  assign n5780 = x299 | n4926 ;
  assign n5781 = n5234 | n5780 ;
  assign n5782 = n5779 | n5781 ;
  assign n5783 = x299 & ~n4958 ;
  assign n5784 = ~n4954 & n5783 ;
  assign n5785 = x232 & ~n5784 ;
  assign n5786 = n5782 & n5785 ;
  assign n5787 = ~n5778 & n5786 ;
  assign n5788 = ~x39 & x232 ;
  assign n5789 = x299 | n4915 ;
  assign n5790 = ~n5783 & n5789 ;
  assign n5791 = ( x39 & ~n5788 ) | ( x39 & n5790 ) | ( ~n5788 & n5790 ) ;
  assign n5792 = n5787 | n5791 ;
  assign n5793 = ~n5776 & n5792 ;
  assign n5794 = x38 | n5793 ;
  assign n5795 = ~n4662 & n5794 ;
  assign n5796 = ( x100 & ~n5770 ) | ( x100 & n5795 ) | ( ~n5770 & n5795 ) ;
  assign n5797 = n2004 | n5796 ;
  assign n5798 = ~n5767 & n5797 ;
  assign n5799 = x54 | n5798 ;
  assign n5800 = x92 | n5765 ;
  assign n5801 = x54 & n5800 ;
  assign n5802 = n5799 & ~n5801 ;
  assign n5803 = x74 | n5802 ;
  assign n5804 = ~n4657 & n5803 ;
  assign n5805 = ( x55 & ~n5761 ) | ( x55 & n5804 ) | ( ~n5761 & n5804 ) ;
  assign n5806 = n2057 | n5805 ;
  assign n5807 = ~n4649 & n5806 ;
  assign n5808 = x954 | n5807 ;
  assign n5809 = x24 & x954 ;
  assign n5810 = n5808 & ~n5809 ;
  assign n5811 = n2041 | n2082 ;
  assign n5812 = n2192 | n5811 ;
  assign n5813 = ~n1898 & n5812 ;
  assign n5814 = x62 & ~n5813 ;
  assign n5815 = x75 & ~n1898 ;
  assign n5816 = x92 | n5815 ;
  assign n5817 = ~x100 & n3347 ;
  assign n5818 = x39 | x100 ;
  assign n5819 = n1868 | n5031 ;
  assign n5820 = ~x299 & n5819 ;
  assign n5821 = x299 & n2161 ;
  assign n5822 = n5820 | n5821 ;
  assign n5823 = n2082 | n5822 ;
  assign n5824 = ( x39 & n5818 ) | ( x39 & ~n5823 ) | ( n5818 & ~n5823 ) ;
  assign n5825 = n5817 | n5824 ;
  assign n5826 = x100 | n2082 ;
  assign n5827 = x39 & n5826 ;
  assign n5828 = x38 | n5827 ;
  assign n5829 = n5825 & ~n5828 ;
  assign n5830 = n1898 | n5829 ;
  assign n5831 = ( x75 & ~x87 ) | ( x75 & n5830 ) | ( ~x87 & n5830 ) ;
  assign n5832 = ~n1898 & n5811 ;
  assign n5833 = ( x75 & x87 ) | ( x75 & ~n5832 ) | ( x87 & ~n5832 ) ;
  assign n5834 = n5831 | n5833 ;
  assign n5835 = ~n5816 & n5834 ;
  assign n5836 = n2082 | n2111 ;
  assign n5837 = ~n1898 & n5836 ;
  assign n5838 = x92 & ~n5837 ;
  assign n5839 = n2030 | n5838 ;
  assign n5840 = n5835 | n5839 ;
  assign n5841 = ~n1898 & n2030 ;
  assign n5842 = x55 | n5841 ;
  assign n5843 = n5840 & ~n5842 ;
  assign n5844 = n2041 | n4654 ;
  assign n5845 = n2082 | n5844 ;
  assign n5846 = x74 | n5845 ;
  assign n5847 = ~n1898 & n5846 ;
  assign n5848 = x55 & ~n5847 ;
  assign n5849 = x56 | n5848 ;
  assign n5850 = n5843 | n5849 ;
  assign n5851 = n2045 | n2082 ;
  assign n5852 = x56 & ~n1898 ;
  assign n5853 = n5851 & n5852 ;
  assign n5854 = x62 | n5853 ;
  assign n5855 = n5850 & ~n5854 ;
  assign n5856 = n5814 | n5855 ;
  assign n5857 = ~n2057 & n5856 ;
  assign n5858 = n1898 & n2057 ;
  assign n5859 = n5857 | n5858 ;
  assign n5860 = x119 & x1056 ;
  assign n5861 = ~x228 & x252 ;
  assign n5862 = x119 | n5861 ;
  assign n5863 = ~x468 & n5862 ;
  assign n5864 = ~n5860 & n5863 ;
  assign n5865 = x119 & x1077 ;
  assign n5866 = n5863 & ~n5865 ;
  assign n5867 = x119 & x1073 ;
  assign n5868 = n5863 & ~n5867 ;
  assign n5869 = x119 & x1041 ;
  assign n5870 = n5863 & ~n5869 ;
  assign n5871 = x352 & ~x353 ;
  assign n5872 = ~x352 & x353 ;
  assign n5873 = n5871 | n5872 ;
  assign n5874 = ( x360 & ~x462 ) | ( x360 & n5873 ) | ( ~x462 & n5873 ) ;
  assign n5875 = ( ~x360 & x462 ) | ( ~x360 & n5874 ) | ( x462 & n5874 ) ;
  assign n5876 = ( ~n5873 & n5874 ) | ( ~n5873 & n5875 ) | ( n5874 & n5875 ) ;
  assign n5877 = x354 & ~n5876 ;
  assign n5878 = ~x354 & n5876 ;
  assign n5879 = n5877 | n5878 ;
  assign n5880 = x74 | n4817 ;
  assign n5881 = ~n1868 & n4800 ;
  assign n5882 = x75 | n2041 ;
  assign n5883 = ( x87 & ~n5881 ) | ( x87 & n5882 ) | ( ~n5881 & n5882 ) ;
  assign n5884 = ~x122 & x829 ;
  assign n5885 = n1525 | n4664 ;
  assign n5886 = x841 | n1254 ;
  assign n5887 = x90 & ~n5886 ;
  assign n5888 = x93 | n5887 ;
  assign n5889 = ~n5885 & n5888 ;
  assign n5890 = x51 | n5889 ;
  assign n5891 = x94 | n1244 ;
  assign n5892 = n1340 | n5891 ;
  assign n5893 = x86 | n1215 ;
  assign n5894 = ~x88 & x98 ;
  assign n5895 = ~n5893 & n5894 ;
  assign n5896 = ~n5892 & n5895 ;
  assign n5897 = x97 | n5896 ;
  assign n5898 = ~n1590 & n5897 ;
  assign n5899 = x35 | n1255 ;
  assign n5900 = x70 | n5899 ;
  assign n5901 = n5898 & ~n5900 ;
  assign n5902 = n5890 | n5901 ;
  assign n5903 = ~n1464 & n5902 ;
  assign n5904 = x96 | n1864 ;
  assign n5905 = n5903 & ~n5904 ;
  assign n5906 = n4799 & n5905 ;
  assign n5907 = ~n5884 & n5906 ;
  assign n5908 = x96 | n5903 ;
  assign n5909 = n1272 | n4909 ;
  assign n5910 = x96 & n5909 ;
  assign n5911 = n1864 | n5910 ;
  assign n5912 = n1692 & n5884 ;
  assign n5913 = ~n5911 & n5912 ;
  assign n5914 = n5908 & n5913 ;
  assign n5915 = n5907 | n5914 ;
  assign n5916 = ~x1093 & n5915 ;
  assign n5917 = ( x87 & ~n5882 ) | ( x87 & n5916 ) | ( ~n5882 & n5916 ) ;
  assign n5918 = ~n5883 & n5917 ;
  assign n5919 = x567 | n5918 ;
  assign n5920 = ~n5880 & n5919 ;
  assign n5921 = ~x299 & n1834 ;
  assign n5922 = x299 & n1524 ;
  assign n5923 = n5921 | n5922 ;
  assign n5924 = x232 & ~n4713 ;
  assign n5925 = ~n5923 & n5924 ;
  assign n5926 = n1984 | n5925 ;
  assign n5927 = ~x24 & n5034 ;
  assign n5928 = ~n1287 & n4795 ;
  assign n5929 = x1091 & n5928 ;
  assign n5930 = n5912 & n5929 ;
  assign n5931 = n5927 & n5930 ;
  assign n5932 = x1093 & n5931 ;
  assign n5933 = ~n5926 & n5932 ;
  assign n5934 = x75 & ~n5933 ;
  assign n5935 = ~n1287 & n1289 ;
  assign n5936 = n4982 & n5935 ;
  assign n5937 = n1290 & n5936 ;
  assign n5938 = x1091 & n5937 ;
  assign n5939 = n4766 & n5938 ;
  assign n5940 = ~x299 & n4989 ;
  assign n5941 = ~x224 & n5940 ;
  assign n5942 = n5939 & n5941 ;
  assign n5943 = n4723 & n5938 ;
  assign n5944 = ~x216 & n5124 ;
  assign n5945 = n5943 & n5944 ;
  assign n5946 = n5942 | n5945 ;
  assign n5947 = ( x38 & n1925 ) | ( x38 & ~n5946 ) | ( n1925 & ~n5946 ) ;
  assign n5948 = x1091 | n5916 ;
  assign n5949 = x1093 & ~n1287 ;
  assign n5950 = x824 & n1692 ;
  assign n5951 = n1464 | n5904 ;
  assign n5952 = n5890 & ~n5951 ;
  assign n5953 = n5950 & n5952 ;
  assign n5954 = ~x829 & n5953 ;
  assign n5955 = n1693 & ~n5911 ;
  assign n5956 = ~x24 & n1314 ;
  assign n5957 = ~x46 & x97 ;
  assign n5958 = ~x108 & n5957 ;
  assign n5959 = ~n4927 & n5958 ;
  assign n5960 = ~n1336 & n5959 ;
  assign n5961 = ~x91 & n5960 ;
  assign n5962 = n5956 | n5961 ;
  assign n5963 = n1269 | n5885 ;
  assign n5964 = n5962 & ~n5963 ;
  assign n5965 = n5890 | n5964 ;
  assign n5966 = ~n1465 & n5965 ;
  assign n5967 = ( x96 & n5955 ) | ( x96 & n5966 ) | ( n5955 & n5966 ) ;
  assign n5968 = n5954 | n5967 ;
  assign n5969 = ~x122 & n5968 ;
  assign n5970 = x122 & n4799 ;
  assign n5971 = n5952 & n5970 ;
  assign n5972 = n5969 | n5971 ;
  assign n5973 = n5949 & n5972 ;
  assign n5974 = x1091 & ~n5973 ;
  assign n5975 = ~n5916 & n5974 ;
  assign n5976 = x39 | n5975 ;
  assign n5977 = n5948 & ~n5976 ;
  assign n5978 = ( x39 & ~n5947 ) | ( x39 & n5977 ) | ( ~n5947 & n5977 ) ;
  assign n5979 = x100 | n5978 ;
  assign n5980 = n4984 & n5952 ;
  assign n5981 = ~n5947 & n5980 ;
  assign n5982 = ~n5974 & n5981 ;
  assign n5983 = n5979 | n5982 ;
  assign n5984 = x1093 & n5912 ;
  assign n5985 = n5928 & n5984 ;
  assign n5986 = ~n1868 & n5985 ;
  assign n5987 = x1091 & n5986 ;
  assign n5988 = x228 & n5987 ;
  assign n5989 = n1925 | n5925 ;
  assign n5990 = n5988 & ~n5989 ;
  assign n5991 = x100 & ~n5990 ;
  assign n5992 = n5983 & ~n5991 ;
  assign n5993 = x87 | n5992 ;
  assign n5994 = ~n1868 & n5950 ;
  assign n5995 = ~x1091 & x1093 ;
  assign n5996 = ~n5994 & n5995 ;
  assign n5997 = x1093 & n1287 ;
  assign n5998 = n4799 & ~n5997 ;
  assign n5999 = ~n1868 & n5998 ;
  assign n6000 = n5995 | n5999 ;
  assign n6001 = ~n1976 & n6000 ;
  assign n6002 = ~n5996 & n6001 ;
  assign n6003 = x87 & ~n6002 ;
  assign n6004 = n5993 & ~n6003 ;
  assign n6005 = x75 | n6004 ;
  assign n6006 = ~n5934 & n6005 ;
  assign n6007 = x567 & ~n6006 ;
  assign n6008 = n5920 & ~n6007 ;
  assign n6009 = x350 & ~x592 ;
  assign n6010 = n6008 | n6009 ;
  assign n6011 = x87 | n5991 ;
  assign n6012 = n5979 & ~n6011 ;
  assign n6013 = x1091 | n5881 ;
  assign n6014 = x1091 & ~n5999 ;
  assign n6015 = x87 & ~x100 ;
  assign n6016 = ~n1925 & n6015 ;
  assign n6017 = ~n6014 & n6016 ;
  assign n6018 = n6013 & n6017 ;
  assign n6019 = x75 | n6018 ;
  assign n6020 = n6012 | n6019 ;
  assign n6021 = ~n5934 & n6020 ;
  assign n6022 = x567 & ~n6021 ;
  assign n6023 = n5920 & ~n6022 ;
  assign n6024 = n6009 & ~n6023 ;
  assign n6025 = ( x316 & ~x348 ) | ( x316 & x349 ) | ( ~x348 & x349 ) ;
  assign n6026 = ( ~x316 & x348 ) | ( ~x316 & n6025 ) | ( x348 & n6025 ) ;
  assign n6027 = ( ~x349 & n6025 ) | ( ~x349 & n6026 ) | ( n6025 & n6026 ) ;
  assign n6028 = ( x315 & ~x322 ) | ( x315 & x359 ) | ( ~x322 & x359 ) ;
  assign n6029 = ( ~x315 & x322 ) | ( ~x315 & n6028 ) | ( x322 & n6028 ) ;
  assign n6030 = ( ~x359 & n6028 ) | ( ~x359 & n6029 ) | ( n6028 & n6029 ) ;
  assign n6031 = ~n6027 & n6030 ;
  assign n6032 = n6027 & ~n6030 ;
  assign n6033 = n6031 | n6032 ;
  assign n6034 = ( x321 & ~x347 ) | ( x321 & n6033 ) | ( ~x347 & n6033 ) ;
  assign n6035 = ( ~x321 & x347 ) | ( ~x321 & n6034 ) | ( x347 & n6034 ) ;
  assign n6036 = ( ~n6033 & n6034 ) | ( ~n6033 & n6035 ) | ( n6034 & n6035 ) ;
  assign n6037 = n6024 | n6036 ;
  assign n6038 = n6010 & ~n6037 ;
  assign n6039 = x452 & ~x455 ;
  assign n6040 = ~x452 & x455 ;
  assign n6041 = n6039 | n6040 ;
  assign n6042 = x355 & ~n6041 ;
  assign n6043 = ~x355 & n6041 ;
  assign n6044 = n6042 | n6043 ;
  assign n6045 = ( x320 & ~x342 ) | ( x320 & x460 ) | ( ~x342 & x460 ) ;
  assign n6046 = ( ~x320 & x342 ) | ( ~x320 & n6045 ) | ( x342 & n6045 ) ;
  assign n6047 = ( ~x460 & n6045 ) | ( ~x460 & n6046 ) | ( n6045 & n6046 ) ;
  assign n6048 = ( x361 & ~x441 ) | ( x361 & n6047 ) | ( ~x441 & n6047 ) ;
  assign n6049 = ( ~x361 & x441 ) | ( ~x361 & n6048 ) | ( x441 & n6048 ) ;
  assign n6050 = ( ~n6047 & n6048 ) | ( ~n6047 & n6049 ) | ( n6048 & n6049 ) ;
  assign n6051 = x458 & ~n6050 ;
  assign n6052 = ~x458 & n6050 ;
  assign n6053 = n6051 | n6052 ;
  assign n6054 = n6044 | n6053 ;
  assign n6055 = n6044 & n6053 ;
  assign n6056 = n6054 & ~n6055 ;
  assign n6057 = x1196 & n6056 ;
  assign n6058 = x350 | x592 ;
  assign n6059 = ~n6008 & n6058 ;
  assign n6060 = n6023 | n6058 ;
  assign n6061 = n6036 & n6060 ;
  assign n6062 = ~n6059 & n6061 ;
  assign n6063 = n6057 | n6062 ;
  assign n6064 = n6038 | n6063 ;
  assign n6065 = x592 | n6023 ;
  assign n6066 = x592 & ~n6008 ;
  assign n6067 = n6065 & ~n6066 ;
  assign n6068 = n6057 & ~n6067 ;
  assign n6069 = x1198 & ~n6068 ;
  assign n6070 = n6064 & n6069 ;
  assign n6071 = x455 | n6067 ;
  assign n6072 = x455 & ~n6008 ;
  assign n6073 = n6071 & ~n6072 ;
  assign n6074 = x452 | n6073 ;
  assign n6075 = x455 & ~n6067 ;
  assign n6076 = x455 | n6008 ;
  assign n6077 = ~n6075 & n6076 ;
  assign n6078 = x452 & ~n6077 ;
  assign n6079 = n6074 & ~n6078 ;
  assign n6080 = x355 | n6079 ;
  assign n6081 = x452 | n6077 ;
  assign n6082 = x452 & ~n6073 ;
  assign n6083 = n6081 & ~n6082 ;
  assign n6084 = x355 & ~n6083 ;
  assign n6085 = n6080 & ~n6084 ;
  assign n6086 = ( x458 & n6050 ) | ( x458 & ~n6085 ) | ( n6050 & ~n6085 ) ;
  assign n6087 = x355 | n6083 ;
  assign n6088 = x355 & ~n6079 ;
  assign n6089 = n6087 & ~n6088 ;
  assign n6090 = ( x458 & ~n6050 ) | ( x458 & n6089 ) | ( ~n6050 & n6089 ) ;
  assign n6091 = ~n6086 & n6090 ;
  assign n6092 = x1196 & ~n6091 ;
  assign n6093 = ( x458 & n6050 ) | ( x458 & n6085 ) | ( n6050 & n6085 ) ;
  assign n6094 = ( ~x458 & n6050 ) | ( ~x458 & n6089 ) | ( n6050 & n6089 ) ;
  assign n6095 = n6093 & n6094 ;
  assign n6096 = n6092 & ~n6095 ;
  assign n6097 = x1196 | n6008 ;
  assign n6098 = ~x1198 & n6097 ;
  assign n6099 = ~n6096 & n6098 ;
  assign n6100 = n6070 | n6099 ;
  assign n6101 = x343 & ~x344 ;
  assign n6102 = ~x343 & x344 ;
  assign n6103 = n6101 | n6102 ;
  assign n6104 = ( x327 & ~x362 ) | ( x327 & n6103 ) | ( ~x362 & n6103 ) ;
  assign n6105 = ( ~x327 & x362 ) | ( ~x327 & n6104 ) | ( x362 & n6104 ) ;
  assign n6106 = ( ~n6103 & n6104 ) | ( ~n6103 & n6105 ) | ( n6104 & n6105 ) ;
  assign n6107 = ( x323 & ~x345 ) | ( x323 & x346 ) | ( ~x345 & x346 ) ;
  assign n6108 = ( ~x323 & x345 ) | ( ~x323 & n6107 ) | ( x345 & n6107 ) ;
  assign n6109 = ( ~x346 & n6107 ) | ( ~x346 & n6108 ) | ( n6107 & n6108 ) ;
  assign n6110 = ( x358 & ~x450 ) | ( x358 & n6109 ) | ( ~x450 & n6109 ) ;
  assign n6111 = ( ~x358 & x450 ) | ( ~x358 & n6110 ) | ( x450 & n6110 ) ;
  assign n6112 = ( ~n6109 & n6110 ) | ( ~n6109 & n6111 ) | ( n6110 & n6111 ) ;
  assign n6113 = ~n6106 & n6112 ;
  assign n6114 = ( x1197 & ~n6112 ) | ( x1197 & n6113 ) | ( ~n6112 & n6113 ) ;
  assign n6115 = ( n6106 & n6113 ) | ( n6106 & n6114 ) | ( n6113 & n6114 ) ;
  assign n6116 = n6100 & ~n6115 ;
  assign n6117 = n6067 & n6115 ;
  assign n6118 = n6116 | n6117 ;
  assign n6119 = ~x351 & x1199 ;
  assign n6120 = n6118 | n6119 ;
  assign n6121 = x1199 & ~n6067 ;
  assign n6122 = ~x351 & n6121 ;
  assign n6123 = n6120 & ~n6122 ;
  assign n6124 = x461 | n6123 ;
  assign n6125 = x351 & x1199 ;
  assign n6126 = n6118 | n6125 ;
  assign n6127 = x351 & n6121 ;
  assign n6128 = n6126 & ~n6127 ;
  assign n6129 = x461 & ~n6128 ;
  assign n6130 = n6124 & ~n6129 ;
  assign n6131 = x357 | n6130 ;
  assign n6132 = x461 | n6128 ;
  assign n6133 = x461 & ~n6123 ;
  assign n6134 = n6132 & ~n6133 ;
  assign n6135 = x357 & ~n6134 ;
  assign n6136 = n6131 & ~n6135 ;
  assign n6137 = ( x356 & n5879 ) | ( x356 & ~n6136 ) | ( n5879 & ~n6136 ) ;
  assign n6138 = x357 | n6134 ;
  assign n6139 = x357 & ~n6130 ;
  assign n6140 = n6138 & ~n6139 ;
  assign n6141 = ( x356 & ~n5879 ) | ( x356 & n6140 ) | ( ~n5879 & n6140 ) ;
  assign n6142 = n6137 & ~n6141 ;
  assign n6143 = x591 | n6142 ;
  assign n6144 = ( x356 & n5879 ) | ( x356 & n6136 ) | ( n5879 & n6136 ) ;
  assign n6145 = ( ~x356 & n5879 ) | ( ~x356 & n6140 ) | ( n5879 & n6140 ) ;
  assign n6146 = n6144 | n6145 ;
  assign n6147 = ~n6143 & n6146 ;
  assign n6148 = x590 & ~x591 ;
  assign n6149 = ( x590 & ~n6008 ) | ( x590 & n6148 ) | ( ~n6008 & n6148 ) ;
  assign n6150 = ~n6147 & n6149 ;
  assign n6151 = x285 | x286 ;
  assign n6152 = x289 | n6151 ;
  assign n6153 = x288 | n6152 ;
  assign n6154 = ( x363 & ~x372 ) | ( x363 & x386 ) | ( ~x372 & x386 ) ;
  assign n6155 = ( ~x363 & x372 ) | ( ~x363 & n6154 ) | ( x372 & n6154 ) ;
  assign n6156 = ( ~x386 & n6154 ) | ( ~x386 & n6155 ) | ( n6154 & n6155 ) ;
  assign n6157 = ( x337 & ~x339 ) | ( x337 & x387 ) | ( ~x339 & x387 ) ;
  assign n6158 = ( ~x337 & x339 ) | ( ~x337 & n6157 ) | ( x339 & n6157 ) ;
  assign n6159 = ( ~x387 & n6157 ) | ( ~x387 & n6158 ) | ( n6157 & n6158 ) ;
  assign n6160 = x380 & n6159 ;
  assign n6161 = x380 | n6159 ;
  assign n6162 = ~n6160 & n6161 ;
  assign n6163 = ( x338 & ~x388 ) | ( x338 & n6162 ) | ( ~x388 & n6162 ) ;
  assign n6164 = ( ~x338 & x388 ) | ( ~x338 & n6163 ) | ( x388 & n6163 ) ;
  assign n6165 = ( ~n6162 & n6163 ) | ( ~n6162 & n6164 ) | ( n6163 & n6164 ) ;
  assign n6166 = ~n6156 & n6165 ;
  assign n6167 = n6156 & ~n6165 ;
  assign n6168 = n6166 | n6167 ;
  assign n6169 = x1196 & n6168 ;
  assign n6170 = x365 & ~x447 ;
  assign n6171 = ~x365 & x447 ;
  assign n6172 = n6170 | n6171 ;
  assign n6173 = x364 & ~x366 ;
  assign n6174 = ~x364 & x366 ;
  assign n6175 = n6173 | n6174 ;
  assign n6176 = ( x336 & ~x383 ) | ( x336 & n6175 ) | ( ~x383 & n6175 ) ;
  assign n6177 = ( ~x336 & x383 ) | ( ~x336 & n6176 ) | ( x383 & n6176 ) ;
  assign n6178 = ( ~n6175 & n6176 ) | ( ~n6175 & n6177 ) | ( n6176 & n6177 ) ;
  assign n6179 = ~n6172 & n6178 ;
  assign n6180 = n6172 & ~n6178 ;
  assign n6181 = n6179 | n6180 ;
  assign n6182 = x367 & n6181 ;
  assign n6183 = x367 | n6181 ;
  assign n6184 = ~n6182 & n6183 ;
  assign n6185 = x368 | x389 ;
  assign n6186 = x368 & x389 ;
  assign n6187 = n6185 & ~n6186 ;
  assign n6188 = ~n6184 & n6187 ;
  assign n6189 = ( x1197 & ~n6187 ) | ( x1197 & n6188 ) | ( ~n6187 & n6188 ) ;
  assign n6190 = ( n6184 & n6188 ) | ( n6184 & n6189 ) | ( n6188 & n6189 ) ;
  assign n6191 = n6169 | n6190 ;
  assign n6192 = x377 & x592 ;
  assign n6193 = n6008 | n6192 ;
  assign n6194 = ~n6023 & n6192 ;
  assign n6195 = ( x376 & ~x381 ) | ( x376 & x439 ) | ( ~x381 & x439 ) ;
  assign n6196 = ( ~x376 & x381 ) | ( ~x376 & n6195 ) | ( x381 & n6195 ) ;
  assign n6197 = ( ~x439 & n6195 ) | ( ~x439 & n6196 ) | ( n6195 & n6196 ) ;
  assign n6198 = ( x317 & ~x378 ) | ( x317 & x385 ) | ( ~x378 & x385 ) ;
  assign n6199 = ( ~x317 & x378 ) | ( ~x317 & n6198 ) | ( x378 & n6198 ) ;
  assign n6200 = ( ~x385 & n6198 ) | ( ~x385 & n6199 ) | ( n6198 & n6199 ) ;
  assign n6201 = ~n6197 & n6200 ;
  assign n6202 = n6197 & ~n6200 ;
  assign n6203 = n6201 | n6202 ;
  assign n6204 = ( x379 & ~x382 ) | ( x379 & n6203 ) | ( ~x382 & n6203 ) ;
  assign n6205 = ( ~x379 & x382 ) | ( ~x379 & n6204 ) | ( x382 & n6204 ) ;
  assign n6206 = ( ~n6203 & n6204 ) | ( ~n6203 & n6205 ) | ( n6204 & n6205 ) ;
  assign n6207 = n6194 | n6206 ;
  assign n6208 = n6193 & ~n6207 ;
  assign n6209 = ~x377 & x592 ;
  assign n6210 = n6008 | n6209 ;
  assign n6211 = ~n6023 & n6209 ;
  assign n6212 = n6206 & ~n6211 ;
  assign n6213 = n6210 & n6212 ;
  assign n6214 = n6208 | n6213 ;
  assign n6215 = ~n6191 & n6214 ;
  assign n6216 = x592 & ~n6023 ;
  assign n6217 = x592 | n6008 ;
  assign n6218 = ~n6216 & n6217 ;
  assign n6219 = n6191 & n6218 ;
  assign n6220 = n6215 | n6219 ;
  assign n6221 = x1199 & ~n6220 ;
  assign n6222 = n6008 & ~n6190 ;
  assign n6223 = x1196 & ~n6218 ;
  assign n6224 = n6190 & n6218 ;
  assign n6225 = ( x1196 & ~n6222 ) | ( x1196 & n6224 ) | ( ~n6222 & n6224 ) ;
  assign n6226 = ( n6222 & ~n6223 ) | ( n6222 & n6225 ) | ( ~n6223 & n6225 ) ;
  assign n6227 = ( x1199 & n6168 ) | ( x1199 & n6226 ) | ( n6168 & n6226 ) ;
  assign n6228 = n6222 | n6224 ;
  assign n6229 = ( x1199 & ~n6168 ) | ( x1199 & n6228 ) | ( ~n6168 & n6228 ) ;
  assign n6230 = n6227 | n6229 ;
  assign n6231 = ~n6221 & n6230 ;
  assign n6232 = x374 | n6231 ;
  assign n6233 = ~x1198 & x1199 ;
  assign n6234 = ~n6220 & n6233 ;
  assign n6235 = ( x1198 & ~n6218 ) | ( x1198 & n6234 ) | ( ~n6218 & n6234 ) ;
  assign n6236 = ( x1198 & n6230 ) | ( x1198 & ~n6234 ) | ( n6230 & ~n6234 ) ;
  assign n6237 = ~n6235 & n6236 ;
  assign n6238 = x374 & ~n6237 ;
  assign n6239 = n6232 & ~n6238 ;
  assign n6240 = x369 & ~n6239 ;
  assign n6241 = x374 | n6237 ;
  assign n6242 = x374 & ~n6231 ;
  assign n6243 = n6241 & ~n6242 ;
  assign n6244 = x369 | n6243 ;
  assign n6245 = ~n6240 & n6244 ;
  assign n6246 = x370 | n6245 ;
  assign n6247 = x369 | n6239 ;
  assign n6248 = x369 & ~n6243 ;
  assign n6249 = n6247 & ~n6248 ;
  assign n6250 = x370 & ~n6249 ;
  assign n6251 = n6246 & ~n6250 ;
  assign n6252 = x371 | n6251 ;
  assign n6253 = x370 | n6249 ;
  assign n6254 = x370 & ~n6245 ;
  assign n6255 = n6253 & ~n6254 ;
  assign n6256 = x371 & ~n6255 ;
  assign n6257 = n6252 & ~n6256 ;
  assign n6258 = x373 | n6257 ;
  assign n6259 = x371 | n6255 ;
  assign n6260 = x371 & ~n6251 ;
  assign n6261 = n6259 & ~n6260 ;
  assign n6262 = x373 & ~n6261 ;
  assign n6263 = n6258 & ~n6262 ;
  assign n6264 = ( x384 & ~x440 ) | ( x384 & x442 ) | ( ~x440 & x442 ) ;
  assign n6265 = ( ~x384 & x440 ) | ( ~x384 & n6264 ) | ( x440 & n6264 ) ;
  assign n6266 = ( ~x442 & n6264 ) | ( ~x442 & n6265 ) | ( n6264 & n6265 ) ;
  assign n6267 = ( x375 & ~n6263 ) | ( x375 & n6266 ) | ( ~n6263 & n6266 ) ;
  assign n6268 = x373 | n6261 ;
  assign n6269 = x373 & ~n6257 ;
  assign n6270 = n6268 & ~n6269 ;
  assign n6271 = ( x375 & ~n6266 ) | ( x375 & n6270 ) | ( ~n6266 & n6270 ) ;
  assign n6272 = n6267 & ~n6271 ;
  assign n6273 = x591 | n6272 ;
  assign n6274 = ( x375 & n6263 ) | ( x375 & n6266 ) | ( n6263 & n6266 ) ;
  assign n6275 = ( ~x375 & n6266 ) | ( ~x375 & n6270 ) | ( n6266 & n6270 ) ;
  assign n6276 = n6274 | n6275 ;
  assign n6277 = ~n6273 & n6276 ;
  assign n6278 = x590 | x591 ;
  assign n6279 = x1197 & ~n6067 ;
  assign n6280 = x394 | x396 ;
  assign n6281 = x394 & x396 ;
  assign n6282 = n6280 & ~n6281 ;
  assign n6283 = ( x328 & ~x408 ) | ( x328 & n6282 ) | ( ~x408 & n6282 ) ;
  assign n6284 = ( ~x328 & x408 ) | ( ~x328 & n6283 ) | ( x408 & n6283 ) ;
  assign n6285 = ( ~n6282 & n6283 ) | ( ~n6282 & n6284 ) | ( n6283 & n6284 ) ;
  assign n6286 = ( x395 & ~x398 ) | ( x395 & x399 ) | ( ~x398 & x399 ) ;
  assign n6287 = ( ~x395 & x398 ) | ( ~x395 & n6286 ) | ( x398 & n6286 ) ;
  assign n6288 = ( ~x399 & n6286 ) | ( ~x399 & n6287 ) | ( n6286 & n6287 ) ;
  assign n6289 = ( x329 & ~x400 ) | ( x329 & n6288 ) | ( ~x400 & n6288 ) ;
  assign n6290 = ( ~x329 & x400 ) | ( ~x329 & n6289 ) | ( x400 & n6289 ) ;
  assign n6291 = ( ~n6288 & n6289 ) | ( ~n6288 & n6290 ) | ( n6289 & n6290 ) ;
  assign n6292 = n6285 & ~n6291 ;
  assign n6293 = ~n6285 & n6291 ;
  assign n6294 = n6292 | n6293 ;
  assign n6295 = x1198 & n6294 ;
  assign n6296 = n6067 & n6295 ;
  assign n6297 = ( x319 & ~x324 ) | ( x319 & x456 ) | ( ~x324 & x456 ) ;
  assign n6298 = ( ~x319 & x324 ) | ( ~x319 & n6297 ) | ( x324 & n6297 ) ;
  assign n6299 = ( ~x456 & n6297 ) | ( ~x456 & n6298 ) | ( n6297 & n6298 ) ;
  assign n6300 = x390 & ~x410 ;
  assign n6301 = ~x390 & x410 ;
  assign n6302 = n6300 | n6301 ;
  assign n6303 = ( x397 & ~x404 ) | ( x397 & x412 ) | ( ~x404 & x412 ) ;
  assign n6304 = ( ~x397 & x404 ) | ( ~x397 & n6303 ) | ( x404 & n6303 ) ;
  assign n6305 = ( ~x412 & n6303 ) | ( ~x412 & n6304 ) | ( n6303 & n6304 ) ;
  assign n6306 = ( n6299 & n6302 ) | ( n6299 & ~n6305 ) | ( n6302 & ~n6305 ) ;
  assign n6307 = ( ~n6302 & n6305 ) | ( ~n6302 & n6306 ) | ( n6305 & n6306 ) ;
  assign n6308 = ( ~n6299 & n6306 ) | ( ~n6299 & n6307 ) | ( n6306 & n6307 ) ;
  assign n6309 = x411 & ~n6308 ;
  assign n6310 = ~x411 & n6308 ;
  assign n6311 = n6309 | n6310 ;
  assign n6312 = ( n5979 & n5983 ) | ( n5979 & ~n6311 ) | ( n5983 & ~n6311 ) ;
  assign n6313 = ~n6011 & n6312 ;
  assign n6314 = n6000 & n6016 ;
  assign n6315 = n5994 & ~n6311 ;
  assign n6316 = n5995 & ~n6315 ;
  assign n6317 = n6314 & ~n6316 ;
  assign n6318 = x75 | x592 ;
  assign n6319 = x1196 & ~n6318 ;
  assign n6320 = ~n6317 & n6319 ;
  assign n6321 = ~n6313 & n6320 ;
  assign n6322 = x1196 | n6005 ;
  assign n6323 = ~n6321 & n6322 ;
  assign n6324 = x1199 | n6323 ;
  assign n6325 = x1196 & n6311 ;
  assign n6326 = ~x75 & n6325 ;
  assign n6327 = ( x401 & ~x402 ) | ( x401 & x406 ) | ( ~x402 & x406 ) ;
  assign n6328 = ( ~x401 & x402 ) | ( ~x401 & n6327 ) | ( x402 & n6327 ) ;
  assign n6329 = ( ~x406 & n6327 ) | ( ~x406 & n6328 ) | ( n6327 & n6328 ) ;
  assign n6330 = x325 & ~x326 ;
  assign n6331 = ~x325 & x326 ;
  assign n6332 = n6330 | n6331 ;
  assign n6333 = ( x403 & ~x405 ) | ( x403 & n6332 ) | ( ~x405 & n6332 ) ;
  assign n6334 = ( ~x403 & x405 ) | ( ~x403 & n6333 ) | ( x405 & n6333 ) ;
  assign n6335 = ( ~n6332 & n6333 ) | ( ~n6332 & n6334 ) | ( n6333 & n6334 ) ;
  assign n6336 = ~n6329 & n6335 ;
  assign n6337 = n6329 & ~n6335 ;
  assign n6338 = n6336 | n6337 ;
  assign n6339 = ( x318 & ~x409 ) | ( x318 & n6338 ) | ( ~x409 & n6338 ) ;
  assign n6340 = ( ~x318 & x409 ) | ( ~x318 & n6339 ) | ( x409 & n6339 ) ;
  assign n6341 = ( ~n6338 & n6339 ) | ( ~n6338 & n6340 ) | ( n6339 & n6340 ) ;
  assign n6342 = n6326 | n6341 ;
  assign n6343 = ( n5979 & n5983 ) | ( n5979 & ~n6342 ) | ( n5983 & ~n6342 ) ;
  assign n6344 = ~n6011 & n6343 ;
  assign n6345 = n5994 & ~n6341 ;
  assign n6346 = n5995 & ~n6345 ;
  assign n6347 = n6314 & ~n6346 ;
  assign n6348 = x1199 & ~n6318 ;
  assign n6349 = n6316 & n6347 ;
  assign n6350 = x1196 & n6349 ;
  assign n6351 = ( ~n6347 & n6348 ) | ( ~n6347 & n6350 ) | ( n6348 & n6350 ) ;
  assign n6352 = ~n6344 & n6351 ;
  assign n6353 = ~n6006 & n6318 ;
  assign n6354 = n6352 | n6353 ;
  assign n6355 = n6324 & ~n6354 ;
  assign n6356 = x567 & ~n6355 ;
  assign n6357 = n5920 & ~n6295 ;
  assign n6358 = ~n6356 & n6357 ;
  assign n6359 = n6296 | n6358 ;
  assign n6360 = x1197 | n6359 ;
  assign n6361 = ~n6279 & n6360 ;
  assign n6362 = x333 & ~n6361 ;
  assign n6363 = x333 | n6359 ;
  assign n6364 = ~n6362 & n6363 ;
  assign n6365 = x391 & ~n6364 ;
  assign n6366 = x333 & n6359 ;
  assign n6367 = ~x333 & n6361 ;
  assign n6368 = n6366 | n6367 ;
  assign n6369 = x391 | n6368 ;
  assign n6370 = ~n6365 & n6369 ;
  assign n6371 = x392 | n6370 ;
  assign n6372 = x391 | n6364 ;
  assign n6373 = x391 & ~n6368 ;
  assign n6374 = n6372 & ~n6373 ;
  assign n6375 = x392 & ~n6374 ;
  assign n6376 = n6371 & ~n6375 ;
  assign n6377 = x393 | n6376 ;
  assign n6378 = x392 | n6374 ;
  assign n6379 = x392 & ~n6370 ;
  assign n6380 = n6378 & ~n6379 ;
  assign n6381 = x393 & ~n6380 ;
  assign n6382 = n6377 & ~n6381 ;
  assign n6383 = x335 & ~x413 ;
  assign n6384 = ~x335 & x413 ;
  assign n6385 = n6383 | n6384 ;
  assign n6386 = ( x407 & ~x463 ) | ( x407 & n6385 ) | ( ~x463 & n6385 ) ;
  assign n6387 = ( ~x407 & x463 ) | ( ~x407 & n6386 ) | ( x463 & n6386 ) ;
  assign n6388 = ( ~n6385 & n6386 ) | ( ~n6385 & n6387 ) | ( n6386 & n6387 ) ;
  assign n6389 = ( x334 & n6382 ) | ( x334 & n6388 ) | ( n6382 & n6388 ) ;
  assign n6390 = x393 | n6380 ;
  assign n6391 = x393 & ~n6376 ;
  assign n6392 = n6390 & ~n6391 ;
  assign n6393 = ( ~x334 & n6388 ) | ( ~x334 & n6392 ) | ( n6388 & n6392 ) ;
  assign n6394 = n6389 | n6393 ;
  assign n6395 = ( x334 & ~n6382 ) | ( x334 & n6388 ) | ( ~n6382 & n6388 ) ;
  assign n6396 = ( x334 & ~n6388 ) | ( x334 & n6392 ) | ( ~n6388 & n6392 ) ;
  assign n6397 = n6395 & ~n6396 ;
  assign n6398 = n6394 & ~n6397 ;
  assign n6399 = ( x590 & n6278 ) | ( x590 & n6398 ) | ( n6278 & n6398 ) ;
  assign n6400 = n6277 | n6399 ;
  assign n6401 = ~n6153 & n6400 ;
  assign n6402 = ~n6150 & n6401 ;
  assign n6403 = n5927 & n5985 ;
  assign n6404 = x1091 & ~n6403 ;
  assign n6405 = n5926 | n6404 ;
  assign n6406 = ~x122 & x1093 ;
  assign n6407 = ~x98 & n5950 ;
  assign n6408 = n6406 & n6407 ;
  assign n6409 = x1091 | n6408 ;
  assign n6410 = ~n6405 & n6409 ;
  assign n6411 = n5950 & n6406 ;
  assign n6412 = ~x1091 & n6411 ;
  assign n6413 = ~x98 & n6412 ;
  assign n6414 = n5926 & n6413 ;
  assign n6415 = x75 & ~n6414 ;
  assign n6416 = ~n6410 & n6415 ;
  assign n6417 = x228 & ~n5925 ;
  assign n6418 = ( ~n1925 & n6413 ) | ( ~n1925 & n6417 ) | ( n6413 & n6417 ) ;
  assign n6419 = x1091 & ~n5986 ;
  assign n6420 = n6409 & ~n6419 ;
  assign n6421 = ( n1925 & n6417 ) | ( n1925 & ~n6420 ) | ( n6417 & ~n6420 ) ;
  assign n6422 = n6418 & ~n6421 ;
  assign n6423 = ( x100 & n2364 ) | ( x100 & ~n6413 ) | ( n2364 & ~n6413 ) ;
  assign n6424 = ~n6422 & n6423 ;
  assign n6425 = x87 | n6424 ;
  assign n6426 = ( x38 & x100 ) | ( x38 & n6413 ) | ( x100 & n6413 ) ;
  assign n6427 = ~x122 & n6407 ;
  assign n6428 = x122 & n5953 ;
  assign n6429 = n6427 | n6428 ;
  assign n6430 = x1093 & n6429 ;
  assign n6431 = n5948 | n6430 ;
  assign n6432 = ~n5976 & n6431 ;
  assign n6433 = ~x216 & n5005 ;
  assign n6434 = n6413 & ~n6433 ;
  assign n6435 = x299 & ~n6434 ;
  assign n6436 = x1091 & ~n5937 ;
  assign n6437 = n6409 & ~n6436 ;
  assign n6438 = n4714 & n6437 ;
  assign n6439 = ~n4714 & n6413 ;
  assign n6440 = n6438 | n6439 ;
  assign n6441 = ( n4721 & n6433 ) | ( n4721 & n6440 ) | ( n6433 & n6440 ) ;
  assign n6442 = ~n4751 & n6437 ;
  assign n6443 = n4751 & n6413 ;
  assign n6444 = n6442 | n6443 ;
  assign n6445 = ( ~n4721 & n6433 ) | ( ~n4721 & n6444 ) | ( n6433 & n6444 ) ;
  assign n6446 = n6441 & n6445 ;
  assign n6447 = n6435 & ~n6446 ;
  assign n6448 = ~x223 & n4346 ;
  assign n6449 = n6413 & ~n6448 ;
  assign n6450 = ( n4764 & n6440 ) | ( n4764 & n6448 ) | ( n6440 & n6448 ) ;
  assign n6451 = ( ~n4764 & n6444 ) | ( ~n4764 & n6448 ) | ( n6444 & n6448 ) ;
  assign n6452 = n6450 & n6451 ;
  assign n6453 = n6449 | n6452 ;
  assign n6454 = ( x39 & n4757 ) | ( x39 & n6453 ) | ( n4757 & n6453 ) ;
  assign n6455 = ~n6447 & n6454 ;
  assign n6456 = n6432 | n6455 ;
  assign n6457 = ( ~x38 & x100 ) | ( ~x38 & n6456 ) | ( x100 & n6456 ) ;
  assign n6458 = n6426 | n6457 ;
  assign n6459 = ~n6425 & n6458 ;
  assign n6460 = x122 & n5994 ;
  assign n6461 = n6427 | n6460 ;
  assign n6462 = x1093 & n6461 ;
  assign n6463 = n6013 | n6462 ;
  assign n6464 = n1976 | n6014 ;
  assign n6465 = n6463 & ~n6464 ;
  assign n6466 = n6413 | n6465 ;
  assign n6467 = x87 & n6466 ;
  assign n6468 = x75 | n6467 ;
  assign n6469 = n6459 | n6468 ;
  assign n6470 = ~n6416 & n6469 ;
  assign n6471 = x567 & ~n6470 ;
  assign n6472 = n5920 & ~n6471 ;
  assign n6473 = x567 & n6413 ;
  assign n6474 = n5880 & n6473 ;
  assign n6475 = n6472 | n6474 ;
  assign n6476 = x592 & ~n6475 ;
  assign n6477 = n6065 & ~n6476 ;
  assign n6478 = n6115 & ~n6477 ;
  assign n6479 = x355 & n6053 ;
  assign n6480 = x355 | n6053 ;
  assign n6481 = ~n6479 & n6480 ;
  assign n6482 = x455 | n6477 ;
  assign n6483 = x455 & ~n6475 ;
  assign n6484 = n6482 & ~n6483 ;
  assign n6485 = ( x452 & n6481 ) | ( x452 & ~n6484 ) | ( n6481 & ~n6484 ) ;
  assign n6486 = x455 & ~n6477 ;
  assign n6487 = x455 | n6475 ;
  assign n6488 = ~n6486 & n6487 ;
  assign n6489 = ( x452 & ~n6481 ) | ( x452 & n6488 ) | ( ~n6481 & n6488 ) ;
  assign n6490 = ~n6485 & n6489 ;
  assign n6491 = x1196 & ~n6490 ;
  assign n6492 = ( x452 & n6481 ) | ( x452 & n6484 ) | ( n6481 & n6484 ) ;
  assign n6493 = ( ~x452 & n6481 ) | ( ~x452 & n6488 ) | ( n6481 & n6488 ) ;
  assign n6494 = n6492 & n6493 ;
  assign n6495 = n6491 & ~n6494 ;
  assign n6496 = x1196 | n6475 ;
  assign n6497 = ~x1198 & n6496 ;
  assign n6498 = ~n6495 & n6497 ;
  assign n6499 = n6058 & ~n6475 ;
  assign n6500 = n6061 & ~n6499 ;
  assign n6501 = n6009 | n6475 ;
  assign n6502 = ~n6037 & n6501 ;
  assign n6503 = n6057 | n6502 ;
  assign n6504 = n6500 | n6503 ;
  assign n6505 = n6057 & ~n6477 ;
  assign n6506 = x1198 & ~n6505 ;
  assign n6507 = n6504 & n6506 ;
  assign n6508 = n6115 | n6507 ;
  assign n6509 = n6498 | n6508 ;
  assign n6510 = ~n6478 & n6509 ;
  assign n6511 = n6119 | n6510 ;
  assign n6512 = x1199 & ~n6477 ;
  assign n6513 = ~x351 & n6512 ;
  assign n6514 = n6511 & ~n6513 ;
  assign n6515 = x461 | n6514 ;
  assign n6516 = n6125 | n6510 ;
  assign n6517 = x351 & n6512 ;
  assign n6518 = n6516 & ~n6517 ;
  assign n6519 = x461 & ~n6518 ;
  assign n6520 = n6515 & ~n6519 ;
  assign n6521 = x357 | n6520 ;
  assign n6522 = x461 | n6518 ;
  assign n6523 = x461 & ~n6514 ;
  assign n6524 = n6522 & ~n6523 ;
  assign n6525 = x357 & ~n6524 ;
  assign n6526 = n6521 & ~n6525 ;
  assign n6527 = ( x356 & n5879 ) | ( x356 & ~n6526 ) | ( n5879 & ~n6526 ) ;
  assign n6528 = x357 | n6524 ;
  assign n6529 = x357 & ~n6520 ;
  assign n6530 = n6528 & ~n6529 ;
  assign n6531 = ( x356 & ~n5879 ) | ( x356 & n6530 ) | ( ~n5879 & n6530 ) ;
  assign n6532 = n6527 & ~n6531 ;
  assign n6533 = x591 | n6532 ;
  assign n6534 = ( x356 & n5879 ) | ( x356 & n6526 ) | ( n5879 & n6526 ) ;
  assign n6535 = ( ~x356 & n5879 ) | ( ~x356 & n6530 ) | ( n5879 & n6530 ) ;
  assign n6536 = n6534 | n6535 ;
  assign n6537 = ~n6533 & n6536 ;
  assign n6538 = x591 & n6475 ;
  assign n6539 = x590 & ~n6538 ;
  assign n6540 = ~n6537 & n6539 ;
  assign n6541 = x592 | n6475 ;
  assign n6542 = ~n6216 & n6541 ;
  assign n6543 = n6191 & n6542 ;
  assign n6544 = n6209 | n6475 ;
  assign n6545 = n6212 & n6544 ;
  assign n6546 = n6192 | n6475 ;
  assign n6547 = ~n6207 & n6546 ;
  assign n6548 = n6545 | n6547 ;
  assign n6549 = ~n6191 & n6548 ;
  assign n6550 = ( x1199 & n6543 ) | ( x1199 & n6549 ) | ( n6543 & n6549 ) ;
  assign n6551 = ~n6191 & n6475 ;
  assign n6552 = ( ~x1199 & n6543 ) | ( ~x1199 & n6551 ) | ( n6543 & n6551 ) ;
  assign n6553 = n6550 | n6552 ;
  assign n6554 = x374 | n6553 ;
  assign n6555 = x1198 | n6553 ;
  assign n6556 = x1198 & ~n6542 ;
  assign n6557 = n6555 & ~n6556 ;
  assign n6558 = x374 & ~n6557 ;
  assign n6559 = n6554 & ~n6558 ;
  assign n6560 = x369 & ~n6559 ;
  assign n6561 = x374 | n6557 ;
  assign n6562 = x374 & ~n6553 ;
  assign n6563 = n6561 & ~n6562 ;
  assign n6564 = x369 | n6563 ;
  assign n6565 = ~n6560 & n6564 ;
  assign n6566 = x370 | n6565 ;
  assign n6567 = x369 | n6559 ;
  assign n6568 = x369 & ~n6563 ;
  assign n6569 = n6567 & ~n6568 ;
  assign n6570 = x370 & ~n6569 ;
  assign n6571 = n6566 & ~n6570 ;
  assign n6572 = ( x373 & ~x375 ) | ( x373 & n6266 ) | ( ~x375 & n6266 ) ;
  assign n6573 = ( ~x373 & x375 ) | ( ~x373 & n6572 ) | ( x375 & n6572 ) ;
  assign n6574 = ( ~n6266 & n6572 ) | ( ~n6266 & n6573 ) | ( n6572 & n6573 ) ;
  assign n6575 = ( x371 & ~n6571 ) | ( x371 & n6574 ) | ( ~n6571 & n6574 ) ;
  assign n6576 = x370 | n6569 ;
  assign n6577 = x370 & ~n6565 ;
  assign n6578 = n6576 & ~n6577 ;
  assign n6579 = ( x371 & ~n6574 ) | ( x371 & n6578 ) | ( ~n6574 & n6578 ) ;
  assign n6580 = n6575 & ~n6579 ;
  assign n6581 = x591 | n6580 ;
  assign n6582 = ( x371 & n6571 ) | ( x371 & n6574 ) | ( n6571 & n6574 ) ;
  assign n6583 = ( ~x371 & n6574 ) | ( ~x371 & n6578 ) | ( n6574 & n6578 ) ;
  assign n6584 = n6582 | n6583 ;
  assign n6585 = ~n6581 & n6584 ;
  assign n6586 = x334 & ~n6388 ;
  assign n6587 = ~x334 & n6388 ;
  assign n6588 = n6586 | n6587 ;
  assign n6589 = x393 & ~n6588 ;
  assign n6590 = ~x393 & n6588 ;
  assign n6591 = n6589 | n6590 ;
  assign n6592 = ~n6311 & n6408 ;
  assign n6593 = ~x1091 & n6592 ;
  assign n6594 = ~n6448 & n6593 ;
  assign n6595 = x299 | n6594 ;
  assign n6596 = ~n6341 & n6408 ;
  assign n6597 = ~x1091 & n6596 ;
  assign n6598 = ~n6448 & n6597 ;
  assign n6599 = x299 | n6598 ;
  assign n6600 = n6595 & n6599 ;
  assign n6601 = ~n6341 & n6593 ;
  assign n6602 = n4714 & n5938 ;
  assign n6603 = n6601 | n6602 ;
  assign n6604 = ( n4764 & n6448 ) | ( n4764 & n6603 ) | ( n6448 & n6603 ) ;
  assign n6605 = ~n4751 & n5938 ;
  assign n6606 = n6601 | n6605 ;
  assign n6607 = ( ~n4764 & n6448 ) | ( ~n4764 & n6606 ) | ( n6448 & n6606 ) ;
  assign n6608 = n6604 & n6607 ;
  assign n6609 = n6600 | n6608 ;
  assign n6610 = ~n6433 & n6593 ;
  assign n6611 = x299 & ~n6610 ;
  assign n6612 = ~n6433 & n6597 ;
  assign n6613 = x299 & ~n6612 ;
  assign n6614 = n6611 | n6613 ;
  assign n6615 = ( n4721 & n6433 ) | ( n4721 & n6603 ) | ( n6433 & n6603 ) ;
  assign n6616 = ( ~n4721 & n6433 ) | ( ~n4721 & n6606 ) | ( n6433 & n6606 ) ;
  assign n6617 = n6615 & n6616 ;
  assign n6618 = n6614 & ~n6617 ;
  assign n6619 = x39 & ~n6618 ;
  assign n6620 = n6609 & n6619 ;
  assign n6621 = ~n5948 & n6311 ;
  assign n6622 = n6432 & ~n6621 ;
  assign n6623 = ~n6341 & n6407 ;
  assign n6624 = x122 | n6623 ;
  assign n6625 = x1093 & n6624 ;
  assign n6626 = ~n6341 & n6428 ;
  assign n6627 = ( ~x122 & n6625 ) | ( ~x122 & n6626 ) | ( n6625 & n6626 ) ;
  assign n6628 = n5948 | n6627 ;
  assign n6629 = n6622 & n6628 ;
  assign n6630 = n6620 | n6629 ;
  assign n6631 = ~x38 & n6630 ;
  assign n6632 = x38 & n6593 ;
  assign n6633 = x100 | n6632 ;
  assign n6634 = x38 & n6597 ;
  assign n6635 = x100 | n6634 ;
  assign n6636 = n6633 & n6635 ;
  assign n6637 = n6631 | n6636 ;
  assign n6638 = n5921 & n5987 ;
  assign n6639 = n4713 | n5922 ;
  assign n6640 = ~n5921 & n6639 ;
  assign n6641 = x1091 | n6601 ;
  assign n6642 = n6640 & n6641 ;
  assign n6643 = ~n6419 & n6642 ;
  assign n6644 = n6638 | n6643 ;
  assign n6645 = x228 & n6644 ;
  assign n6646 = x228 & n6640 ;
  assign n6647 = n6601 & ~n6646 ;
  assign n6648 = x232 & ~n6647 ;
  assign n6649 = ~n6645 & n6648 ;
  assign n6650 = x232 | n6601 ;
  assign n6651 = n5988 | n6650 ;
  assign n6652 = ~n1925 & n6651 ;
  assign n6653 = ~n6649 & n6652 ;
  assign n6654 = ( x100 & n2364 ) | ( x100 & ~n6601 ) | ( n2364 & ~n6601 ) ;
  assign n6655 = ~n6653 & n6654 ;
  assign n6656 = n6637 & ~n6655 ;
  assign n6657 = x87 | n6656 ;
  assign n6658 = n1976 & n6593 ;
  assign n6659 = x87 & ~n6658 ;
  assign n6660 = n1976 & n6597 ;
  assign n6661 = x87 & ~n6660 ;
  assign n6662 = n6659 | n6661 ;
  assign n6663 = ~n6013 & n6311 ;
  assign n6664 = ~n6013 & n6341 ;
  assign n6665 = n6465 & ~n6664 ;
  assign n6666 = ~n6663 & n6665 ;
  assign n6667 = n6662 & ~n6666 ;
  assign n6668 = n6657 & ~n6667 ;
  assign n6669 = x75 | n6668 ;
  assign n6670 = n5926 & n6593 ;
  assign n6671 = x75 & ~n6670 ;
  assign n6672 = n5926 & n6597 ;
  assign n6673 = x75 & ~n6672 ;
  assign n6674 = n6671 | n6673 ;
  assign n6675 = ~n6405 & n6641 ;
  assign n6676 = n6674 & ~n6675 ;
  assign n6677 = n6669 & ~n6676 ;
  assign n6678 = ~x592 & x1196 ;
  assign n6679 = x567 & n6593 ;
  assign n6680 = n5880 & n6679 ;
  assign n6681 = n6678 & ~n6680 ;
  assign n6682 = ( ~n6623 & n6678 ) | ( ~n6623 & n6681 ) | ( n6678 & n6681 ) ;
  assign n6683 = ~n6677 & n6682 ;
  assign n6684 = x567 & n6597 ;
  assign n6685 = n5880 & n6684 ;
  assign n6686 = x592 | x1196 ;
  assign n6687 = n6685 | n6686 ;
  assign n6688 = n6661 & ~n6665 ;
  assign n6689 = n5991 & ~n6597 ;
  assign n6690 = ~n5976 & n6628 ;
  assign n6691 = n6597 | n6605 ;
  assign n6692 = ( ~n4764 & n6448 ) | ( ~n4764 & n6691 ) | ( n6448 & n6691 ) ;
  assign n6693 = n6597 | n6602 ;
  assign n6694 = ( n4764 & n6448 ) | ( n4764 & n6693 ) | ( n6448 & n6693 ) ;
  assign n6695 = n6692 & n6694 ;
  assign n6696 = n6599 | n6695 ;
  assign n6697 = ( ~n4721 & n6433 ) | ( ~n4721 & n6691 ) | ( n6433 & n6691 ) ;
  assign n6698 = ( n4721 & n6433 ) | ( n4721 & n6693 ) | ( n6433 & n6693 ) ;
  assign n6699 = n6697 & n6698 ;
  assign n6700 = n6613 & ~n6699 ;
  assign n6701 = x39 & ~n6700 ;
  assign n6702 = n6696 & n6701 ;
  assign n6703 = n6690 | n6702 ;
  assign n6704 = ~x38 & n6703 ;
  assign n6705 = n6635 | n6704 ;
  assign n6706 = ~n6689 & n6705 ;
  assign n6707 = x87 | n6706 ;
  assign n6708 = ~n6688 & n6707 ;
  assign n6709 = x75 | n6708 ;
  assign n6710 = x1091 | n6596 ;
  assign n6711 = ~n6405 & n6710 ;
  assign n6712 = n6673 & ~n6711 ;
  assign n6713 = n6709 & ~n6712 ;
  assign n6714 = n6687 | n6713 ;
  assign n6715 = ~n6683 & n6714 ;
  assign n6716 = x567 & ~n6715 ;
  assign n6717 = ~n6682 & n6687 ;
  assign n6718 = n5920 | n6717 ;
  assign n6719 = x1199 & n6718 ;
  assign n6720 = ~n6716 & n6719 ;
  assign n6721 = n6593 | n6605 ;
  assign n6722 = ( ~n4764 & n6448 ) | ( ~n4764 & n6721 ) | ( n6448 & n6721 ) ;
  assign n6723 = n6593 | n6602 ;
  assign n6724 = ( n4764 & n6448 ) | ( n4764 & n6723 ) | ( n6448 & n6723 ) ;
  assign n6725 = n6722 & n6724 ;
  assign n6726 = n6595 | n6725 ;
  assign n6727 = ( ~n4721 & n6433 ) | ( ~n4721 & n6721 ) | ( n6433 & n6721 ) ;
  assign n6728 = ( n4721 & n6433 ) | ( n4721 & n6723 ) | ( n6433 & n6723 ) ;
  assign n6729 = n6727 & n6728 ;
  assign n6730 = n6611 & ~n6729 ;
  assign n6731 = x39 & ~n6730 ;
  assign n6732 = n6726 & n6731 ;
  assign n6733 = n6622 | n6732 ;
  assign n6734 = ~x38 & n6733 ;
  assign n6735 = n6633 | n6734 ;
  assign n6736 = n5991 & ~n6593 ;
  assign n6737 = n6735 & ~n6736 ;
  assign n6738 = x87 | n6737 ;
  assign n6739 = n6465 & ~n6663 ;
  assign n6740 = n6659 & ~n6739 ;
  assign n6741 = n6738 & ~n6740 ;
  assign n6742 = x75 | n6741 ;
  assign n6743 = x1091 | n6592 ;
  assign n6744 = ~n6405 & n6743 ;
  assign n6745 = n6671 & ~n6744 ;
  assign n6746 = n6742 & ~n6745 ;
  assign n6747 = x567 & ~n6746 ;
  assign n6748 = n5920 & ~n6747 ;
  assign n6749 = n6681 & ~n6748 ;
  assign n6750 = ~x1199 & n6496 ;
  assign n6751 = ~n6749 & n6750 ;
  assign n6752 = n6295 | n6751 ;
  assign n6753 = n6720 | n6752 ;
  assign n6754 = ~n6065 & n6295 ;
  assign n6755 = n6476 | n6754 ;
  assign n6756 = n6753 & ~n6755 ;
  assign n6757 = x1197 | n6756 ;
  assign n6758 = x1197 & ~n6477 ;
  assign n6759 = n6757 & ~n6758 ;
  assign n6760 = x333 | n6759 ;
  assign n6761 = x333 & ~n6756 ;
  assign n6762 = n6760 & ~n6761 ;
  assign n6763 = x391 | n6762 ;
  assign n6764 = x333 | n6756 ;
  assign n6765 = x333 & ~n6759 ;
  assign n6766 = n6764 & ~n6765 ;
  assign n6767 = x391 & ~n6766 ;
  assign n6768 = n6763 & ~n6767 ;
  assign n6769 = ( x392 & n6591 ) | ( x392 & n6768 ) | ( n6591 & n6768 ) ;
  assign n6770 = x391 | n6766 ;
  assign n6771 = x391 & ~n6762 ;
  assign n6772 = n6770 & ~n6771 ;
  assign n6773 = ( ~x392 & n6591 ) | ( ~x392 & n6772 ) | ( n6591 & n6772 ) ;
  assign n6774 = n6769 | n6773 ;
  assign n6775 = ( x392 & n6591 ) | ( x392 & ~n6768 ) | ( n6591 & ~n6768 ) ;
  assign n6776 = ( x392 & ~n6591 ) | ( x392 & n6772 ) | ( ~n6591 & n6772 ) ;
  assign n6777 = n6775 & ~n6776 ;
  assign n6778 = n6774 & ~n6777 ;
  assign n6779 = ( x590 & n6278 ) | ( x590 & n6778 ) | ( n6278 & n6778 ) ;
  assign n6780 = n6585 | n6779 ;
  assign n6781 = n6153 & n6780 ;
  assign n6782 = ~n6540 & n6781 ;
  assign n6783 = x588 | n6782 ;
  assign n6784 = n6402 | n6783 ;
  assign n6785 = x57 | n4832 ;
  assign n6786 = ( x433 & ~x449 ) | ( x433 & x451 ) | ( ~x449 & x451 ) ;
  assign n6787 = ( ~x433 & x449 ) | ( ~x433 & n6786 ) | ( x449 & n6786 ) ;
  assign n6788 = ( ~x451 & n6786 ) | ( ~x451 & n6787 ) | ( n6786 & n6787 ) ;
  assign n6789 = x448 & n6788 ;
  assign n6790 = x448 | n6788 ;
  assign n6791 = ~n6789 & n6790 ;
  assign n6792 = x432 & ~x459 ;
  assign n6793 = ~x432 & x459 ;
  assign n6794 = n6792 | n6793 ;
  assign n6795 = ( x421 & ~x454 ) | ( x421 & n6794 ) | ( ~x454 & n6794 ) ;
  assign n6796 = ( ~x421 & x454 ) | ( ~x421 & n6795 ) | ( x454 & n6795 ) ;
  assign n6797 = ( ~n6794 & n6795 ) | ( ~n6794 & n6796 ) | ( n6795 & n6796 ) ;
  assign n6798 = x423 & ~x424 ;
  assign n6799 = ~x423 & x424 ;
  assign n6800 = n6798 | n6799 ;
  assign n6801 = ( x419 & ~x420 ) | ( x419 & n6800 ) | ( ~x420 & n6800 ) ;
  assign n6802 = ( ~x419 & x420 ) | ( ~x419 & n6801 ) | ( x420 & n6801 ) ;
  assign n6803 = ( ~n6800 & n6801 ) | ( ~n6800 & n6802 ) | ( n6801 & n6802 ) ;
  assign n6804 = ~n6797 & n6803 ;
  assign n6805 = n6797 & ~n6803 ;
  assign n6806 = n6804 | n6805 ;
  assign n6807 = x425 | n6806 ;
  assign n6808 = x416 & ~x438 ;
  assign n6809 = ~x416 & x438 ;
  assign n6810 = n6808 | n6809 ;
  assign n6811 = ( x415 & ~x431 ) | ( x415 & n6810 ) | ( ~x431 & n6810 ) ;
  assign n6812 = ( ~x415 & x431 ) | ( ~x415 & n6811 ) | ( x431 & n6811 ) ;
  assign n6813 = ( ~n6810 & n6811 ) | ( ~n6810 & n6812 ) | ( n6811 & n6812 ) ;
  assign n6814 = ( x417 & ~x418 ) | ( x417 & x437 ) | ( ~x418 & x437 ) ;
  assign n6815 = ( ~x417 & x418 ) | ( ~x417 & n6814 ) | ( x418 & n6814 ) ;
  assign n6816 = ( ~x437 & n6814 ) | ( ~x437 & n6815 ) | ( n6814 & n6815 ) ;
  assign n6817 = ( x453 & ~x464 ) | ( x453 & n6816 ) | ( ~x464 & n6816 ) ;
  assign n6818 = ( ~x453 & x464 ) | ( ~x453 & n6817 ) | ( x464 & n6817 ) ;
  assign n6819 = ( ~n6816 & n6817 ) | ( ~n6816 & n6818 ) | ( n6817 & n6818 ) ;
  assign n6820 = ~n6813 & n6819 ;
  assign n6821 = ( x1197 & ~n6819 ) | ( x1197 & n6820 ) | ( ~n6819 & n6820 ) ;
  assign n6822 = ( n6813 & n6820 ) | ( n6813 & n6821 ) | ( n6820 & n6821 ) ;
  assign n6823 = ( x425 & ~x1198 ) | ( x425 & n6806 ) | ( ~x1198 & n6806 ) ;
  assign n6824 = ( n6807 & n6822 ) | ( n6807 & ~n6823 ) | ( n6822 & ~n6823 ) ;
  assign n6825 = n6067 & n6824 ;
  assign n6826 = x443 | x592 ;
  assign n6827 = ~n6008 & n6826 ;
  assign n6828 = n6023 | n6826 ;
  assign n6829 = ~n6827 & n6828 ;
  assign n6830 = x444 | n6829 ;
  assign n6831 = x443 & ~x592 ;
  assign n6832 = n6008 | n6831 ;
  assign n6833 = ~n6023 & n6831 ;
  assign n6834 = n6832 & ~n6833 ;
  assign n6835 = x444 & ~n6834 ;
  assign n6836 = n6830 & ~n6835 ;
  assign n6837 = x414 & ~x422 ;
  assign n6838 = ~x414 & x422 ;
  assign n6839 = n6837 | n6838 ;
  assign n6840 = ( x434 & ~x446 ) | ( x434 & n6839 ) | ( ~x446 & n6839 ) ;
  assign n6841 = ( ~x434 & x446 ) | ( ~x434 & n6840 ) | ( x446 & n6840 ) ;
  assign n6842 = ( ~n6839 & n6840 ) | ( ~n6839 & n6841 ) | ( n6840 & n6841 ) ;
  assign n6843 = ( x429 & ~x435 ) | ( x429 & n6842 ) | ( ~x435 & n6842 ) ;
  assign n6844 = ( ~x429 & x435 ) | ( ~x429 & n6843 ) | ( x435 & n6843 ) ;
  assign n6845 = ( ~n6842 & n6843 ) | ( ~n6842 & n6844 ) | ( n6843 & n6844 ) ;
  assign n6846 = ( x436 & n6836 ) | ( x436 & n6845 ) | ( n6836 & n6845 ) ;
  assign n6847 = x444 | n6834 ;
  assign n6848 = x444 & ~n6829 ;
  assign n6849 = n6847 & ~n6848 ;
  assign n6850 = ( ~x436 & n6845 ) | ( ~x436 & n6849 ) | ( n6845 & n6849 ) ;
  assign n6851 = n6846 & n6850 ;
  assign n6852 = x1196 & ~n6851 ;
  assign n6853 = ( x436 & ~n6836 ) | ( x436 & n6845 ) | ( ~n6836 & n6845 ) ;
  assign n6854 = ( x436 & ~n6845 ) | ( x436 & n6849 ) | ( ~n6845 & n6849 ) ;
  assign n6855 = ~n6853 & n6854 ;
  assign n6856 = n6852 & ~n6855 ;
  assign n6857 = n6097 & ~n6824 ;
  assign n6858 = ~n6856 & n6857 ;
  assign n6859 = n6825 | n6858 ;
  assign n6860 = x428 & n6859 ;
  assign n6861 = ~x428 & n6067 ;
  assign n6862 = n6860 | n6861 ;
  assign n6863 = ~x427 & n6862 ;
  assign n6864 = ~x428 & n6859 ;
  assign n6865 = x428 & n6067 ;
  assign n6866 = n6864 | n6865 ;
  assign n6867 = x427 & n6866 ;
  assign n6868 = n6863 | n6867 ;
  assign n6869 = x430 & n6868 ;
  assign n6870 = ~x427 & n6866 ;
  assign n6871 = x427 & n6862 ;
  assign n6872 = n6870 | n6871 ;
  assign n6873 = ~x430 & n6872 ;
  assign n6874 = n6869 | n6873 ;
  assign n6875 = x426 & n6874 ;
  assign n6876 = x430 & n6872 ;
  assign n6877 = ~x430 & n6868 ;
  assign n6878 = n6876 | n6877 ;
  assign n6879 = ~x426 & n6878 ;
  assign n6880 = n6875 | n6879 ;
  assign n6881 = ( x445 & n6791 ) | ( x445 & ~n6880 ) | ( n6791 & ~n6880 ) ;
  assign n6882 = x426 & n6878 ;
  assign n6883 = ~x426 & n6874 ;
  assign n6884 = n6882 | n6883 ;
  assign n6885 = ( x445 & ~n6791 ) | ( x445 & n6884 ) | ( ~n6791 & n6884 ) ;
  assign n6886 = ~n6881 & n6885 ;
  assign n6887 = x1199 & ~n6886 ;
  assign n6888 = ( x445 & n6791 ) | ( x445 & n6880 ) | ( n6791 & n6880 ) ;
  assign n6889 = ( ~x445 & n6791 ) | ( ~x445 & n6884 ) | ( n6791 & n6884 ) ;
  assign n6890 = n6888 & n6889 ;
  assign n6891 = n6887 & ~n6890 ;
  assign n6892 = x1199 | n6859 ;
  assign n6893 = ~n6278 & n6892 ;
  assign n6894 = ~n6891 & n6893 ;
  assign n6895 = n6008 & n6278 ;
  assign n6896 = n6153 | n6895 ;
  assign n6897 = n6894 | n6896 ;
  assign n6898 = n6278 & n6475 ;
  assign n6899 = n6153 & ~n6898 ;
  assign n6900 = n6475 | n6831 ;
  assign n6901 = ~x436 & x444 ;
  assign n6902 = x436 & ~x444 ;
  assign n6903 = n6901 | n6902 ;
  assign n6904 = n6845 & n6903 ;
  assign n6905 = n6845 | n6903 ;
  assign n6906 = ~n6904 & n6905 ;
  assign n6907 = n6833 | n6906 ;
  assign n6908 = n6900 & ~n6907 ;
  assign n6909 = ~n6475 & n6826 ;
  assign n6910 = n6828 & n6906 ;
  assign n6911 = ~n6909 & n6910 ;
  assign n6912 = x1196 & ~n6911 ;
  assign n6913 = ~n6908 & n6912 ;
  assign n6914 = n6496 & ~n6913 ;
  assign n6915 = n6824 | n6914 ;
  assign n6916 = ~n6477 & n6824 ;
  assign n6917 = n6915 & ~n6916 ;
  assign n6918 = ( x1199 & ~n6278 ) | ( x1199 & n6917 ) | ( ~n6278 & n6917 ) ;
  assign n6919 = ( x427 & x428 ) | ( x427 & n6477 ) | ( x428 & n6477 ) ;
  assign n6920 = ( ~x428 & n6917 ) | ( ~x428 & n6919 ) | ( n6917 & n6919 ) ;
  assign n6921 = ( ~x427 & n6919 ) | ( ~x427 & n6920 ) | ( n6919 & n6920 ) ;
  assign n6922 = x430 & ~n6921 ;
  assign n6923 = ~x427 & x428 ;
  assign n6924 = x427 & ~x428 ;
  assign n6925 = n6923 | n6924 ;
  assign n6926 = n6477 & ~n6925 ;
  assign n6927 = n6917 & n6925 ;
  assign n6928 = n6926 | n6927 ;
  assign n6929 = x430 | n6928 ;
  assign n6930 = ~n6922 & n6929 ;
  assign n6931 = x426 | n6930 ;
  assign n6932 = x430 | n6921 ;
  assign n6933 = x430 & ~n6928 ;
  assign n6934 = n6932 & ~n6933 ;
  assign n6935 = x426 & ~n6934 ;
  assign n6936 = n6931 & ~n6935 ;
  assign n6937 = x445 | n6936 ;
  assign n6938 = x426 | n6934 ;
  assign n6939 = x426 & ~n6930 ;
  assign n6940 = n6938 & ~n6939 ;
  assign n6941 = x445 & ~n6940 ;
  assign n6942 = n6937 & ~n6941 ;
  assign n6943 = ( x448 & n6788 ) | ( x448 & n6942 ) | ( n6788 & n6942 ) ;
  assign n6944 = x445 | n6940 ;
  assign n6945 = x445 & ~n6936 ;
  assign n6946 = n6944 & ~n6945 ;
  assign n6947 = ( ~n6788 & n6943 ) | ( ~n6788 & n6946 ) | ( n6943 & n6946 ) ;
  assign n6948 = ( ~x448 & n6943 ) | ( ~x448 & n6947 ) | ( n6943 & n6947 ) ;
  assign n6949 = ( x1199 & n6278 ) | ( x1199 & ~n6948 ) | ( n6278 & ~n6948 ) ;
  assign n6950 = n6918 & ~n6949 ;
  assign n6951 = n6899 & ~n6950 ;
  assign n6952 = n6897 & ~n6951 ;
  assign n6953 = x588 & ~n6952 ;
  assign n6954 = n6785 | n6953 ;
  assign n6955 = n6784 & ~n6954 ;
  assign n6956 = ~x592 & n6056 ;
  assign n6957 = ~n6047 & n6473 ;
  assign n6958 = ~n6956 & n6957 ;
  assign n6959 = ( x361 & ~x458 ) | ( x361 & n6044 ) | ( ~x458 & n6044 ) ;
  assign n6960 = ( ~x361 & x458 ) | ( ~x361 & n6959 ) | ( x458 & n6959 ) ;
  assign n6961 = ( ~n6044 & n6959 ) | ( ~n6044 & n6960 ) | ( n6959 & n6960 ) ;
  assign n6962 = ~x441 & n6961 ;
  assign n6963 = n6047 & n6473 ;
  assign n6964 = ( x441 & x592 ) | ( x441 & ~n6961 ) | ( x592 & ~n6961 ) ;
  assign n6965 = ( n6962 & n6963 ) | ( n6962 & n6964 ) | ( n6963 & n6964 ) ;
  assign n6966 = x1196 & ~n6965 ;
  assign n6967 = ~n6958 & n6966 ;
  assign n6968 = x1198 | n6967 ;
  assign n6969 = ~x592 & n6473 ;
  assign n6970 = x1198 & n6969 ;
  assign n6971 = x350 & n6036 ;
  assign n6972 = ( n6036 & n6057 ) | ( n6036 & ~n6971 ) | ( n6057 & ~n6971 ) ;
  assign n6973 = ( x350 & ~n6971 ) | ( x350 & n6972 ) | ( ~n6971 & n6972 ) ;
  assign n6974 = n6970 & ~n6973 ;
  assign n6975 = n6968 & ~n6974 ;
  assign n6976 = n6115 | n6975 ;
  assign n6977 = ~x592 & n6976 ;
  assign n6978 = n6473 & ~n6977 ;
  assign n6979 = n6119 | n6978 ;
  assign n6980 = x592 & n6473 ;
  assign n6981 = x1199 & ~n6980 ;
  assign n6982 = ~x351 & n6981 ;
  assign n6983 = n6979 & ~n6982 ;
  assign n6984 = x461 | n6983 ;
  assign n6985 = n6125 | n6978 ;
  assign n6986 = x351 & n6981 ;
  assign n6987 = n6985 & ~n6986 ;
  assign n6988 = x461 & ~n6987 ;
  assign n6989 = n6984 & ~n6988 ;
  assign n6990 = x357 | n6989 ;
  assign n6991 = x461 | n6987 ;
  assign n6992 = x461 & ~n6983 ;
  assign n6993 = n6991 & ~n6992 ;
  assign n6994 = x357 & ~n6993 ;
  assign n6995 = n6990 & ~n6994 ;
  assign n6996 = ( x356 & n5879 ) | ( x356 & n6995 ) | ( n5879 & n6995 ) ;
  assign n6997 = x357 | n6993 ;
  assign n6998 = x357 & ~n6989 ;
  assign n6999 = n6997 & ~n6998 ;
  assign n7000 = ( ~n5879 & n6996 ) | ( ~n5879 & n6999 ) | ( n6996 & n6999 ) ;
  assign n7001 = ( ~x356 & n6996 ) | ( ~x356 & n7000 ) | ( n6996 & n7000 ) ;
  assign n7002 = ( x590 & x591 ) | ( x590 & n7001 ) | ( x591 & n7001 ) ;
  assign n7003 = x592 & n6191 ;
  assign n7004 = x377 & n6206 ;
  assign n7005 = ( n6191 & n6206 ) | ( n6191 & ~n7004 ) | ( n6206 & ~n7004 ) ;
  assign n7006 = ( x377 & ~n7004 ) | ( x377 & n7005 ) | ( ~n7004 & n7005 ) ;
  assign n7007 = n6980 & n7006 ;
  assign n7008 = ( x1199 & ~n6473 ) | ( x1199 & n7007 ) | ( ~n6473 & n7007 ) ;
  assign n7009 = n7003 | n7008 ;
  assign n7010 = n6980 & ~n7009 ;
  assign n7011 = ( x369 & ~x370 ) | ( x369 & x374 ) | ( ~x370 & x374 ) ;
  assign n7012 = ( ~x369 & x370 ) | ( ~x369 & n7011 ) | ( x370 & n7011 ) ;
  assign n7013 = ( ~x374 & n7011 ) | ( ~x374 & n7012 ) | ( n7011 & n7012 ) ;
  assign n7014 = ( x371 & ~x373 ) | ( x371 & n7013 ) | ( ~x373 & n7013 ) ;
  assign n7015 = ( ~x371 & x373 ) | ( ~x371 & n7014 ) | ( x373 & n7014 ) ;
  assign n7016 = ( ~n7013 & n7014 ) | ( ~n7013 & n7015 ) | ( n7014 & n7015 ) ;
  assign n7017 = ( x375 & ~n6266 ) | ( x375 & n7016 ) | ( ~n6266 & n7016 ) ;
  assign n7018 = ( ~x375 & n6266 ) | ( ~x375 & n7017 ) | ( n6266 & n7017 ) ;
  assign n7019 = ( ~n7016 & n7017 ) | ( ~n7016 & n7018 ) | ( n7017 & n7018 ) ;
  assign n7020 = x1198 & n7010 ;
  assign n7021 = n7019 & n7020 ;
  assign n7022 = ( n6969 & n7010 ) | ( n6969 & ~n7021 ) | ( n7010 & ~n7021 ) ;
  assign n7023 = ( ~x590 & x591 ) | ( ~x590 & n7022 ) | ( x591 & n7022 ) ;
  assign n7024 = n7002 | n7023 ;
  assign n7025 = x1197 & ~n6980 ;
  assign n7026 = ~x592 & n6684 ;
  assign n7027 = ~n6325 & n7026 ;
  assign n7028 = n6981 & ~n7027 ;
  assign n7029 = ( x1199 & n6678 ) | ( x1199 & n6679 ) | ( n6678 & n6679 ) ;
  assign n7030 = ( x1199 & n6473 ) | ( x1199 & ~n6678 ) | ( n6473 & ~n6678 ) ;
  assign n7031 = n7029 | n7030 ;
  assign n7032 = ~n7028 & n7031 ;
  assign n7033 = x1197 | n7032 ;
  assign n7034 = ~n7025 & n7033 ;
  assign n7035 = x333 | n7034 ;
  assign n7036 = x1198 & ~n6980 ;
  assign n7037 = n7032 & ~n7036 ;
  assign n7038 = n6294 & ~n7037 ;
  assign n7039 = n7032 & ~n7038 ;
  assign n7040 = n7035 & n7039 ;
  assign n7041 = x391 | n7040 ;
  assign n7042 = ( x333 & ~n7034 ) | ( x333 & n7038 ) | ( ~n7034 & n7038 ) ;
  assign n7043 = ( x333 & n7032 ) | ( x333 & ~n7038 ) | ( n7032 & ~n7038 ) ;
  assign n7044 = ~n7042 & n7043 ;
  assign n7045 = x391 & ~n7044 ;
  assign n7046 = n7041 & ~n7045 ;
  assign n7047 = x392 | n7046 ;
  assign n7048 = x391 | n7044 ;
  assign n7049 = x391 & ~n7040 ;
  assign n7050 = n7048 & ~n7049 ;
  assign n7051 = x392 & ~n7050 ;
  assign n7052 = n7047 & ~n7051 ;
  assign n7053 = ( x393 & n6588 ) | ( x393 & n7052 ) | ( n6588 & n7052 ) ;
  assign n7054 = x392 | n7050 ;
  assign n7055 = x392 & ~n7046 ;
  assign n7056 = n7054 & ~n7055 ;
  assign n7057 = ( ~n6588 & n7053 ) | ( ~n6588 & n7056 ) | ( n7053 & n7056 ) ;
  assign n7058 = ( ~x393 & n7053 ) | ( ~x393 & n7057 ) | ( n7053 & n7057 ) ;
  assign n7059 = ( x590 & x591 ) | ( x590 & ~n7058 ) | ( x591 & ~n7058 ) ;
  assign n7060 = ( x590 & ~x591 ) | ( x590 & n6473 ) | ( ~x591 & n6473 ) ;
  assign n7061 = n7059 & ~n7060 ;
  assign n7062 = n7024 & ~n7061 ;
  assign n7063 = x588 | n7062 ;
  assign n7064 = n6153 & n6785 ;
  assign n7065 = ( x436 & ~x443 ) | ( x436 & x444 ) | ( ~x443 & x444 ) ;
  assign n7066 = ( ~x436 & x443 ) | ( ~x436 & n7065 ) | ( x443 & n7065 ) ;
  assign n7067 = ( ~x444 & n7065 ) | ( ~x444 & n7066 ) | ( n7065 & n7066 ) ;
  assign n7068 = n6845 | n7067 ;
  assign n7069 = ( ~n6678 & n6845 ) | ( ~n6678 & n7067 ) | ( n6845 & n7067 ) ;
  assign n7070 = ( n6824 & n7068 ) | ( n6824 & ~n7069 ) | ( n7068 & ~n7069 ) ;
  assign n7071 = n6969 & ~n7070 ;
  assign n7072 = x1199 | n6980 ;
  assign n7073 = n7071 | n7072 ;
  assign n7074 = ~n6278 & n7073 ;
  assign n7075 = ( x426 & ~x430 ) | ( x426 & n6925 ) | ( ~x430 & n6925 ) ;
  assign n7076 = ( ~x426 & x430 ) | ( ~x426 & n7075 ) | ( x430 & n7075 ) ;
  assign n7077 = ( ~n6925 & n7075 ) | ( ~n6925 & n7076 ) | ( n7075 & n7076 ) ;
  assign n7078 = ( x445 & ~x448 ) | ( x445 & n7077 ) | ( ~x448 & n7077 ) ;
  assign n7079 = ( ~x445 & x448 ) | ( ~x445 & n7078 ) | ( x448 & n7078 ) ;
  assign n7080 = ( ~n7077 & n7078 ) | ( ~n7077 & n7079 ) | ( n7078 & n7079 ) ;
  assign n7081 = n7071 & n7080 ;
  assign n7082 = n6980 | n7081 ;
  assign n7083 = ( ~x1199 & n6788 ) | ( ~x1199 & n7082 ) | ( n6788 & n7082 ) ;
  assign n7084 = n7071 & ~n7080 ;
  assign n7085 = n6980 | n7084 ;
  assign n7086 = ( x1199 & n6788 ) | ( x1199 & ~n7085 ) | ( n6788 & ~n7085 ) ;
  assign n7087 = ~n7083 & n7086 ;
  assign n7088 = n7074 & ~n7087 ;
  assign n7089 = n6278 & n6473 ;
  assign n7090 = x588 & ~n7089 ;
  assign n7091 = ~n7088 & n7090 ;
  assign n7092 = n7064 & ~n7091 ;
  assign n7093 = n7063 & n7092 ;
  assign n7094 = x217 | n7093 ;
  assign n7095 = n6955 | n7094 ;
  assign n7096 = n6473 & n7064 ;
  assign n7097 = x217 & ~n7096 ;
  assign n7098 = ( n6153 & ~n6475 ) | ( n6153 & n6785 ) | ( ~n6475 & n6785 ) ;
  assign n7099 = ( n6008 & n6153 ) | ( n6008 & ~n6785 ) | ( n6153 & ~n6785 ) ;
  assign n7100 = ~n7098 & n7099 ;
  assign n7101 = n7097 & ~n7100 ;
  assign n7102 = x1161 | x1162 ;
  assign n7103 = x1163 | n7102 ;
  assign n7104 = n7101 | n7103 ;
  assign n7105 = n7095 & ~n7104 ;
  assign n7106 = x1161 & ~x1163 ;
  assign n7107 = n1290 & n7106 ;
  assign n7108 = ~x31 & x1162 ;
  assign n7109 = n7107 & n7108 ;
  assign n7110 = n7105 | n7109 ;
  assign n7111 = n2057 | n2058 ;
  assign n7112 = n5073 | n7111 ;
  assign n7113 = n4817 | n7112 ;
  assign n7114 = n4784 & ~n4795 ;
  assign n7115 = ~n5026 & n7114 ;
  assign n7116 = ~x137 & n7115 ;
  assign n7117 = x129 & ~n1868 ;
  assign n7118 = ~x137 & x252 ;
  assign n7119 = n4795 & ~n5925 ;
  assign n7120 = n4784 | n7119 ;
  assign n7121 = n7118 & ~n7120 ;
  assign n7122 = n7117 & n7121 ;
  assign n7123 = n7116 | n7122 ;
  assign n7124 = n2364 & n7123 ;
  assign n7125 = x24 | x90 ;
  assign n7126 = n4696 | n7125 ;
  assign n7127 = x50 & ~n1341 ;
  assign n7128 = ~n5893 & n7127 ;
  assign n7129 = n1214 | n1587 ;
  assign n7130 = n1252 | n7129 ;
  assign n7131 = x93 | n7130 ;
  assign n7132 = n7128 & ~n7131 ;
  assign n7133 = ~n7126 & n7132 ;
  assign n7134 = x829 & ~x1093 ;
  assign n7135 = n1692 & n7134 ;
  assign n7136 = n1292 | n7135 ;
  assign n7137 = n6153 & ~n7136 ;
  assign n7138 = x137 | n7137 ;
  assign n7139 = n7133 & n7138 ;
  assign n7140 = x76 & ~x84 ;
  assign n7141 = ~n1227 & n7140 ;
  assign n7142 = x68 | x73 ;
  assign n7143 = x49 | x66 ;
  assign n7144 = n7142 | n7143 ;
  assign n7145 = n7141 & ~n7144 ;
  assign n7146 = x89 | x102 ;
  assign n7147 = n1244 | n7146 ;
  assign n7148 = x64 | x81 ;
  assign n7149 = n1236 | n7148 ;
  assign n7150 = n7147 | n7149 ;
  assign n7151 = n7145 & ~n7150 ;
  assign n7152 = n1243 | n1393 ;
  assign n7153 = x103 | n1220 ;
  assign n7154 = n7152 | n7153 ;
  assign n7155 = n1237 | n1362 ;
  assign n7156 = x45 | x48 ;
  assign n7157 = x61 | x104 ;
  assign n7158 = n7156 | n7157 ;
  assign n7159 = n7155 | n7158 ;
  assign n7160 = n7154 | n7159 ;
  assign n7161 = n7151 & ~n7160 ;
  assign n7162 = ~n5893 & n7161 ;
  assign n7163 = ~n7130 & n7162 ;
  assign n7164 = n1294 | n1682 ;
  assign n7165 = x137 | n5899 ;
  assign n7166 = n7164 | n7165 ;
  assign n7167 = n7137 | n7166 ;
  assign n7168 = ( x24 & ~n7163 ) | ( x24 & n7167 ) | ( ~n7163 & n7167 ) ;
  assign n7169 = n7127 | n7161 ;
  assign n7170 = n1218 | n1253 ;
  assign n7171 = n7169 & ~n7170 ;
  assign n7172 = ( x24 & ~n7167 ) | ( x24 & n7171 ) | ( ~n7167 & n7171 ) ;
  assign n7173 = ~n7168 & n7172 ;
  assign n7174 = n7139 | n7173 ;
  assign n7175 = ~x32 & n7174 ;
  assign n7176 = x24 | x841 ;
  assign n7177 = x32 & n7176 ;
  assign n7178 = ~n1261 & n7177 ;
  assign n7179 = n7175 | n7178 ;
  assign n7180 = ~n4694 & n7179 ;
  assign n7181 = x32 | n7133 ;
  assign n7182 = n4694 & ~n4698 ;
  assign n7183 = n7181 & n7182 ;
  assign n7184 = n7180 | n7183 ;
  assign n7185 = x95 | n2041 ;
  assign n7186 = n7184 & ~n7185 ;
  assign n7187 = n7124 | n7186 ;
  assign n7188 = ~n1998 & n7187 ;
  assign n7189 = x24 | n1279 ;
  assign n7190 = n1256 | n1864 ;
  assign n7191 = x51 | n7190 ;
  assign n7192 = n7189 | n7191 ;
  assign n7193 = n7136 | n7192 ;
  assign n7194 = x252 & ~n7119 ;
  assign n7195 = x87 | n1925 ;
  assign n7196 = x75 & ~x100 ;
  assign n7197 = ~n7195 & n7196 ;
  assign n7198 = ~x137 & n7197 ;
  assign n7199 = ~n4804 & n7198 ;
  assign n7200 = ~n7194 & n7199 ;
  assign n7201 = ~n7193 & n7200 ;
  assign n7202 = n7188 | n7201 ;
  assign n7203 = ~n7113 & n7202 ;
  assign n7204 = x195 | x196 ;
  assign n7205 = x138 | n7204 ;
  assign n7206 = x139 | n7205 ;
  assign n7207 = x118 | n7206 ;
  assign n7208 = x79 | n7207 ;
  assign n7209 = x34 | n7208 ;
  assign n7210 = ~x33 & n7209 ;
  assign n7211 = x149 & x157 ;
  assign n7212 = x149 | x157 ;
  assign n7213 = ~n4713 & n7212 ;
  assign n7214 = ~n7211 & n7213 ;
  assign n7215 = x232 & n7214 ;
  assign n7216 = x75 & ~n7215 ;
  assign n7217 = x100 & ~n7215 ;
  assign n7218 = n7216 | n7217 ;
  assign n7219 = x75 | x100 ;
  assign n7220 = n5924 & ~n7219 ;
  assign n7221 = x169 & n7220 ;
  assign n7222 = n7218 | n7221 ;
  assign n7223 = x74 & n7222 ;
  assign n7224 = x164 & n7220 ;
  assign n7225 = n7218 | n7224 ;
  assign n7226 = ~x74 & n7225 ;
  assign n7227 = n2057 & ~n7226 ;
  assign n7228 = ~n7223 & n7227 ;
  assign n7229 = ( x232 & ~x299 ) | ( x232 & n7214 ) | ( ~x299 & n7214 ) ;
  assign n7230 = x178 & x183 ;
  assign n7231 = x178 | x183 ;
  assign n7232 = ~n4713 & n7231 ;
  assign n7233 = ~n7230 & n7232 ;
  assign n7234 = ( x232 & x299 ) | ( x232 & n7233 ) | ( x299 & n7233 ) ;
  assign n7235 = n7229 & n7234 ;
  assign n7236 = x100 & ~n7235 ;
  assign n7237 = x75 & ~n7235 ;
  assign n7238 = n7236 | n7237 ;
  assign n7239 = x191 & ~x299 ;
  assign n7240 = x169 & x299 ;
  assign n7241 = n7239 | n7240 ;
  assign n7242 = n7220 & n7241 ;
  assign n7243 = n7238 | n7242 ;
  assign n7244 = x74 & n7243 ;
  assign n7245 = x55 | n7244 ;
  assign n7246 = ( x186 & x299 ) | ( x186 & n5924 ) | ( x299 & n5924 ) ;
  assign n7247 = ( x164 & ~x299 ) | ( x164 & n5924 ) | ( ~x299 & n5924 ) ;
  assign n7248 = n7246 & n7247 ;
  assign n7249 = ~n7219 & n7248 ;
  assign n7250 = n7238 | n7249 ;
  assign n7251 = x54 & n7250 ;
  assign n7252 = ~x299 & n5924 ;
  assign n7253 = n4660 & n7252 ;
  assign n7254 = ~x164 & x186 ;
  assign n7255 = n7253 & n7254 ;
  assign n7256 = n4810 & n5924 ;
  assign n7257 = ( x164 & ~x186 ) | ( x164 & n7256 ) | ( ~x186 & n7256 ) ;
  assign n7258 = x299 & n5924 ;
  assign n7259 = n4660 & n7258 ;
  assign n7260 = ( x164 & x186 ) | ( x164 & n7259 ) | ( x186 & n7259 ) ;
  assign n7261 = n7257 & n7260 ;
  assign n7262 = n7255 | n7261 ;
  assign n7263 = x38 & n7262 ;
  assign n7264 = ~x176 & x232 ;
  assign n7265 = x40 | n1236 ;
  assign n7266 = x102 | n7148 ;
  assign n7267 = n1237 | n7266 ;
  assign n7268 = n1245 | n7267 ;
  assign n7269 = n1353 | n7268 ;
  assign n7270 = x60 | n7269 ;
  assign n7271 = n1326 | n1589 ;
  assign n7272 = x53 | n7271 ;
  assign n7273 = n7270 | n7272 ;
  assign n7274 = x58 | n7273 ;
  assign n7275 = n5899 | n7274 ;
  assign n7276 = x32 | n1295 ;
  assign n7277 = n7275 | n7276 ;
  assign n7278 = x95 | n7277 ;
  assign n7279 = n4983 & ~n4987 ;
  assign n7280 = n4740 & n7279 ;
  assign n7281 = n4731 | n7280 ;
  assign n7282 = ~n7278 & n7281 ;
  assign n7283 = n4714 & n7282 ;
  assign n7284 = n7265 | n7283 ;
  assign n7285 = x224 & n4989 ;
  assign n7286 = n7265 | n7285 ;
  assign n7287 = n7284 & n7286 ;
  assign n7288 = ~n7278 & n7280 ;
  assign n7289 = n7265 | n7288 ;
  assign n7290 = ( ~n4713 & n7265 ) | ( ~n4713 & n7289 ) | ( n7265 & n7289 ) ;
  assign n7291 = n4764 & n7290 ;
  assign n7292 = n7286 & n7291 ;
  assign n7293 = x174 & n7292 ;
  assign n7294 = n7287 | n7293 ;
  assign n7295 = ~x299 & n7294 ;
  assign n7296 = x216 & n5005 ;
  assign n7297 = n7265 | n7296 ;
  assign n7298 = x299 & n7297 ;
  assign n7299 = n4731 & ~n7278 ;
  assign n7300 = ~n4751 & n7299 ;
  assign n7301 = n7265 | n7300 ;
  assign n7302 = n4713 | n7301 ;
  assign n7303 = x152 | n7302 ;
  assign n7304 = ~n4713 & n7282 ;
  assign n7305 = n7265 | n7304 ;
  assign n7306 = n4721 & n7305 ;
  assign n7307 = n7284 | n7306 ;
  assign n7308 = ~x154 & n7307 ;
  assign n7309 = n7303 & n7308 ;
  assign n7310 = n4722 & n7289 ;
  assign n7311 = x152 & n7310 ;
  assign n7312 = n7284 | n7311 ;
  assign n7313 = x154 & n7312 ;
  assign n7314 = n7296 & ~n7313 ;
  assign n7315 = ~n7309 & n7314 ;
  assign n7316 = n7298 & ~n7315 ;
  assign n7317 = n7295 | n7316 ;
  assign n7318 = n4765 & n7299 ;
  assign n7319 = ~n7265 & n7285 ;
  assign n7320 = ~n7318 & n7319 ;
  assign n7321 = n7286 & ~n7320 ;
  assign n7322 = ~x299 & n7321 ;
  assign n7323 = n7317 | n7322 ;
  assign n7324 = n7264 & n7323 ;
  assign n7325 = x176 & x232 ;
  assign n7326 = n7317 & n7325 ;
  assign n7327 = n7298 & n7307 ;
  assign n7328 = n4764 & n7305 ;
  assign n7329 = n7286 & n7328 ;
  assign n7330 = n7287 | n7329 ;
  assign n7331 = ~x299 & n7330 ;
  assign n7332 = n7327 | n7331 ;
  assign n7333 = ~x232 & n7332 ;
  assign n7334 = x39 & ~n7333 ;
  assign n7335 = ~n7326 & n7334 ;
  assign n7336 = ~n7324 & n7335 ;
  assign n7337 = x95 & n7265 ;
  assign n7338 = n1491 | n7337 ;
  assign n7339 = x40 | x479 ;
  assign n7340 = ~n1236 & n7277 ;
  assign n7341 = ~n7339 & n7340 ;
  assign n7342 = n7338 & ~n7341 ;
  assign n7343 = x32 & n7265 ;
  assign n7344 = ~n1236 & n7275 ;
  assign n7345 = x70 & ~n7344 ;
  assign n7346 = ~n1236 & n7273 ;
  assign n7347 = x58 & ~n7346 ;
  assign n7348 = x53 & n7270 ;
  assign n7349 = ~x60 & n7127 ;
  assign n7350 = n1582 | n7349 ;
  assign n7351 = ~n7348 & n7350 ;
  assign n7352 = x111 | n1233 ;
  assign n7353 = x68 | n1234 ;
  assign n7354 = x36 | n7353 ;
  assign n7355 = n7352 | n7354 ;
  assign n7356 = x66 | x84 ;
  assign n7357 = x73 & ~x82 ;
  assign n7358 = ~n7356 & n7357 ;
  assign n7359 = ~n7355 & n7358 ;
  assign n7360 = ~n7268 & n7359 ;
  assign n7361 = ~n1226 & n7360 ;
  assign n7362 = ~n1215 & n7361 ;
  assign n7363 = n1236 | n7362 ;
  assign n7364 = n7351 | n7363 ;
  assign n7365 = ~n1326 & n7364 ;
  assign n7366 = n1236 & n1326 ;
  assign n7367 = n1589 | n7366 ;
  assign n7368 = n7365 | n7367 ;
  assign n7369 = ~n1236 & n1589 ;
  assign n7370 = x58 | n7369 ;
  assign n7371 = n7368 & ~n7370 ;
  assign n7372 = n7347 | n7371 ;
  assign n7373 = ~x90 & n7372 ;
  assign n7374 = x841 | n7274 ;
  assign n7375 = ~n1236 & n7374 ;
  assign n7376 = x90 & ~n7375 ;
  assign n7377 = n1278 | n7376 ;
  assign n7378 = n7373 | n7377 ;
  assign n7379 = ~n1236 & n1278 ;
  assign n7380 = x70 | n7379 ;
  assign n7381 = n7378 & ~n7380 ;
  assign n7382 = n7345 | n7381 ;
  assign n7383 = ~x51 & n7382 ;
  assign n7384 = x51 & n1236 ;
  assign n7385 = n1293 | n7384 ;
  assign n7386 = n7383 | n7385 ;
  assign n7387 = ~n1236 & n1293 ;
  assign n7388 = x40 | n7387 ;
  assign n7389 = n7386 & ~n7388 ;
  assign n7390 = ( ~x32 & x40 ) | ( ~x32 & n7389 ) | ( x40 & n7389 ) ;
  assign n7391 = n7343 | n7390 ;
  assign n7392 = ~x95 & n7391 ;
  assign n7393 = n7342 | n7392 ;
  assign n7394 = x72 | x93 ;
  assign n7395 = x90 | n7394 ;
  assign n7396 = n1258 | n7395 ;
  assign n7397 = n7374 | n7396 ;
  assign n7398 = ~n7265 & n7397 ;
  assign n7399 = x32 & ~n7398 ;
  assign n7400 = n7390 | n7399 ;
  assign n7401 = ~x95 & n7400 ;
  assign n7402 = ~x198 & n7401 ;
  assign n7403 = n7393 | n7402 ;
  assign n7404 = n4713 & ~n7403 ;
  assign n7405 = ~n7271 & n7351 ;
  assign n7406 = n1236 | n7405 ;
  assign n7407 = ~x58 & n7406 ;
  assign n7408 = n7347 | n7407 ;
  assign n7409 = ~x90 & n7408 ;
  assign n7410 = n7377 | n7409 ;
  assign n7411 = ~n7380 & n7410 ;
  assign n7412 = n7345 | n7411 ;
  assign n7413 = ~x51 & n7412 ;
  assign n7414 = n7385 | n7413 ;
  assign n7415 = ~n7387 & n7414 ;
  assign n7416 = x40 | n7415 ;
  assign n7417 = ~x32 & n7416 ;
  assign n7418 = n7399 | n7417 ;
  assign n7419 = ~x95 & n7418 ;
  assign n7420 = ~x198 & n7419 ;
  assign n7421 = n4713 | n7337 ;
  assign n7422 = n7343 | n7417 ;
  assign n7423 = ~x95 & n7422 ;
  assign n7424 = n7421 | n7423 ;
  assign n7425 = n7420 | n7424 ;
  assign n7426 = ~n7404 & n7425 ;
  assign n7427 = x183 | n7426 ;
  assign n7428 = x40 | n7343 ;
  assign n7429 = ~n1236 & n4695 ;
  assign n7430 = x32 | n7429 ;
  assign n7431 = x93 & n1236 ;
  assign n7432 = n4695 | n7431 ;
  assign n7433 = n1236 | n7347 ;
  assign n7434 = ~x90 & n7433 ;
  assign n7435 = n7376 | n7434 ;
  assign n7436 = ~x93 & n7435 ;
  assign n7437 = n7432 | n7436 ;
  assign n7438 = ~n7430 & n7437 ;
  assign n7439 = n7428 | n7438 ;
  assign n7440 = ~x95 & n7439 ;
  assign n7441 = n7421 | n7440 ;
  assign n7442 = ~n7404 & n7441 ;
  assign n7443 = x183 & ~n7442 ;
  assign n7444 = n7427 & ~n7443 ;
  assign n7445 = ~x95 & n7444 ;
  assign n7446 = x174 | n7342 ;
  assign n7447 = n7445 | n7446 ;
  assign n7448 = x183 & ~n4713 ;
  assign n7449 = n7403 & ~n7448 ;
  assign n7450 = ~n7170 & n7361 ;
  assign n7451 = ~x90 & n7450 ;
  assign n7452 = n7435 | n7451 ;
  assign n7453 = ~x93 & n7452 ;
  assign n7454 = n7432 | n7453 ;
  assign n7455 = ~n7430 & n7454 ;
  assign n7456 = n7428 | n7455 ;
  assign n7457 = ~x95 & n7456 ;
  assign n7458 = n7342 | n7457 ;
  assign n7459 = ~n4713 & n7458 ;
  assign n7460 = x183 & n7459 ;
  assign n7461 = x174 & ~n7460 ;
  assign n7462 = ~n7449 & n7461 ;
  assign n7463 = x180 | n7462 ;
  assign n7464 = n7447 & ~n7463 ;
  assign n7465 = x174 | n7444 ;
  assign n7466 = x180 & n7465 ;
  assign n7467 = n7421 | n7457 ;
  assign n7468 = ~n7404 & n7467 ;
  assign n7469 = ( ~x174 & x183 ) | ( ~x174 & n7468 ) | ( x183 & n7468 ) ;
  assign n7470 = x40 | n4713 ;
  assign n7471 = n7337 | n7392 ;
  assign n7472 = n7402 | n7471 ;
  assign n7473 = n7470 | n7472 ;
  assign n7474 = ~n7404 & n7473 ;
  assign n7475 = ( x174 & x183 ) | ( x174 & ~n7474 ) | ( x183 & ~n7474 ) ;
  assign n7476 = ~n7469 & n7475 ;
  assign n7477 = n7466 & ~n7476 ;
  assign n7478 = n7464 | n7477 ;
  assign n7479 = ~x193 & n7478 ;
  assign n7480 = ~x40 & n1236 ;
  assign n7481 = x95 & ~n7480 ;
  assign n7482 = x32 & ~n7480 ;
  assign n7483 = n1269 | n1278 ;
  assign n7484 = n1236 & n7483 ;
  assign n7485 = ~n5899 & n7407 ;
  assign n7486 = n7484 | n7485 ;
  assign n7487 = ~x70 & n7486 ;
  assign n7488 = n7345 | n7487 ;
  assign n7489 = ~x51 & n7488 ;
  assign n7490 = n7385 | n7489 ;
  assign n7491 = ~n7387 & n7490 ;
  assign n7492 = ~x40 & n7491 ;
  assign n7493 = x32 | n7492 ;
  assign n7494 = ~n7482 & n7493 ;
  assign n7495 = x95 | n7494 ;
  assign n7496 = ~n7481 & n7495 ;
  assign n7497 = x198 & ~n7496 ;
  assign n7498 = ( x32 & x40 ) | ( x32 & n7398 ) | ( x40 & n7398 ) ;
  assign n7499 = n7493 & ~n7498 ;
  assign n7500 = x95 | n7499 ;
  assign n7501 = ~n7481 & n7500 ;
  assign n7502 = x198 | n7501 ;
  assign n7503 = ~n7497 & n7502 ;
  assign n7504 = n7470 | n7503 ;
  assign n7505 = ~n7404 & n7504 ;
  assign n7506 = x183 | n7505 ;
  assign n7507 = ~n4713 & n7265 ;
  assign n7508 = n4713 & n7403 ;
  assign n7509 = n7507 | n7508 ;
  assign n7510 = x174 | x183 ;
  assign n7511 = ( x174 & ~n7509 ) | ( x174 & n7510 ) | ( ~n7509 & n7510 ) ;
  assign n7512 = n7506 & ~n7511 ;
  assign n7513 = n1295 | n5899 ;
  assign n7514 = n7170 | n7513 ;
  assign n7515 = x32 | n7514 ;
  assign n7516 = n7361 & ~n7515 ;
  assign n7517 = n7265 | n7516 ;
  assign n7518 = ~x95 & n7517 ;
  assign n7519 = n7421 | n7518 ;
  assign n7520 = ~n7404 & n7519 ;
  assign n7521 = ( x174 & ~x183 ) | ( x174 & n7520 ) | ( ~x183 & n7520 ) ;
  assign n7522 = ~n5899 & n7371 ;
  assign n7523 = n7484 | n7522 ;
  assign n7524 = ~x70 & n7523 ;
  assign n7525 = n7345 | n7524 ;
  assign n7526 = ~x51 & n7525 ;
  assign n7527 = n7385 | n7526 ;
  assign n7528 = ~n7388 & n7527 ;
  assign n7529 = x32 | n7528 ;
  assign n7530 = ~n7482 & n7529 ;
  assign n7531 = n1682 & n7265 ;
  assign n7532 = n7530 | n7531 ;
  assign n7533 = ~x95 & n7532 ;
  assign n7534 = n7337 | n7533 ;
  assign n7535 = ~n7498 & n7529 ;
  assign n7536 = x95 | n7535 ;
  assign n7537 = ~n7481 & n7536 ;
  assign n7538 = n7534 | n7537 ;
  assign n7539 = ~x198 & n7538 ;
  assign n7540 = n4713 | n7539 ;
  assign n7541 = n7534 | n7540 ;
  assign n7542 = ~n7404 & n7541 ;
  assign n7543 = ( x174 & x183 ) | ( x174 & n7542 ) | ( x183 & n7542 ) ;
  assign n7544 = n7521 & n7543 ;
  assign n7545 = x180 & ~n7544 ;
  assign n7546 = ~n7512 & n7545 ;
  assign n7547 = ~x95 & n7265 ;
  assign n7548 = n7342 | n7547 ;
  assign n7549 = n4713 | n7548 ;
  assign n7550 = ~n7404 & n7549 ;
  assign n7551 = ( x174 & x183 ) | ( x174 & ~n7550 ) | ( x183 & ~n7550 ) ;
  assign n7552 = x40 | n7491 ;
  assign n7553 = ~x32 & n7552 ;
  assign n7554 = n7343 | n7553 ;
  assign n7555 = ~x95 & n7554 ;
  assign n7556 = n7342 | n7555 ;
  assign n7557 = n7399 | n7553 ;
  assign n7558 = ~x95 & n7557 ;
  assign n7559 = ~x198 & n7558 ;
  assign n7560 = n7556 | n7559 ;
  assign n7561 = ~n4713 & n7560 ;
  assign n7562 = n7508 | n7561 ;
  assign n7563 = ( ~x174 & x183 ) | ( ~x174 & n7562 ) | ( x183 & n7562 ) ;
  assign n7564 = ~n7551 & n7563 ;
  assign n7565 = x180 | n7564 ;
  assign n7566 = n4713 | n7518 ;
  assign n7567 = n7342 | n7566 ;
  assign n7568 = ~n7404 & n7567 ;
  assign n7569 = ( x174 & ~x183 ) | ( x174 & n7568 ) | ( ~x183 & n7568 ) ;
  assign n7570 = n7342 | n7533 ;
  assign n7571 = ~n7507 & n7540 ;
  assign n7572 = n7570 | n7571 ;
  assign n7573 = ~n7404 & n7572 ;
  assign n7574 = ( x174 & x183 ) | ( x174 & n7573 ) | ( x183 & n7573 ) ;
  assign n7575 = n7569 & n7574 ;
  assign n7576 = n7565 | n7575 ;
  assign n7577 = x193 & n7576 ;
  assign n7578 = ~n7546 & n7577 ;
  assign n7579 = n7479 | n7578 ;
  assign n7580 = ~x299 & n7579 ;
  assign n7581 = x158 & x299 ;
  assign n7582 = ~x210 & n7401 ;
  assign n7583 = n7393 | n7582 ;
  assign n7584 = n4713 & n7583 ;
  assign n7585 = n7471 | n7582 ;
  assign n7586 = ~n4713 & n7585 ;
  assign n7587 = n7584 | n7586 ;
  assign n7588 = ( x152 & x172 ) | ( x152 & ~n7587 ) | ( x172 & ~n7587 ) ;
  assign n7589 = n4713 & ~n7583 ;
  assign n7590 = ~x210 & n7419 ;
  assign n7591 = n7424 | n7590 ;
  assign n7592 = ~n7589 & n7591 ;
  assign n7593 = ( x152 & ~x172 ) | ( x152 & n7592 ) | ( ~x172 & n7592 ) ;
  assign n7594 = ~n7588 & n7593 ;
  assign n7595 = n7337 | n7558 ;
  assign n7596 = ~x210 & n7595 ;
  assign n7597 = n4713 | n7596 ;
  assign n7598 = n7337 | n7555 ;
  assign n7599 = n7597 | n7598 ;
  assign n7600 = ~n7589 & n7599 ;
  assign n7601 = ( x152 & x172 ) | ( x152 & n7600 ) | ( x172 & n7600 ) ;
  assign n7602 = ~x210 & n7538 ;
  assign n7603 = n4713 | n7602 ;
  assign n7604 = n7534 | n7603 ;
  assign n7605 = ~n7589 & n7604 ;
  assign n7606 = ( ~x152 & x172 ) | ( ~x152 & n7605 ) | ( x172 & n7605 ) ;
  assign n7607 = n7601 & n7606 ;
  assign n7608 = n7594 | n7607 ;
  assign n7609 = n7581 & n7608 ;
  assign n7610 = ~x158 & x299 ;
  assign n7611 = ~n7589 & n7610 ;
  assign n7612 = ( x152 & x172 ) | ( x152 & n7583 ) | ( x172 & n7583 ) ;
  assign n7613 = n7342 | n7423 ;
  assign n7614 = n7590 | n7613 ;
  assign n7615 = n4713 | n7614 ;
  assign n7616 = ( ~x152 & x172 ) | ( ~x152 & n7615 ) | ( x172 & n7615 ) ;
  assign n7617 = n7612 | n7616 ;
  assign n7618 = n7611 & n7617 ;
  assign n7619 = ~n7507 & n7597 ;
  assign n7620 = n7556 | n7619 ;
  assign n7621 = ( x152 & x172 ) | ( x152 & ~n7620 ) | ( x172 & ~n7620 ) ;
  assign n7622 = ~n7507 & n7603 ;
  assign n7623 = n7570 | n7622 ;
  assign n7624 = ( x152 & ~x172 ) | ( x152 & n7623 ) | ( ~x172 & n7623 ) ;
  assign n7625 = n7621 & ~n7624 ;
  assign n7626 = n7618 & ~n7625 ;
  assign n7627 = x149 | n7626 ;
  assign n7628 = n7609 | n7627 ;
  assign n7629 = n7549 & ~n7589 ;
  assign n7630 = ( x152 & x172 ) | ( x152 & n7629 ) | ( x172 & n7629 ) ;
  assign n7631 = n7567 & ~n7589 ;
  assign n7632 = ( ~x152 & x172 ) | ( ~x152 & n7631 ) | ( x172 & n7631 ) ;
  assign n7633 = n7630 & n7632 ;
  assign n7634 = n7459 | n7584 ;
  assign n7635 = ( x152 & x172 ) | ( x152 & ~n7634 ) | ( x172 & ~n7634 ) ;
  assign n7636 = n7342 | n7440 ;
  assign n7637 = ~n4713 & n7636 ;
  assign n7638 = n7584 | n7637 ;
  assign n7639 = ( x152 & ~x172 ) | ( x152 & n7638 ) | ( ~x172 & n7638 ) ;
  assign n7640 = ~n7635 & n7639 ;
  assign n7641 = n7633 | n7640 ;
  assign n7642 = n7610 & n7641 ;
  assign n7643 = n7467 & ~n7589 ;
  assign n7644 = ( x152 & x172 ) | ( x152 & ~n7643 ) | ( x172 & ~n7643 ) ;
  assign n7645 = n7441 & ~n7589 ;
  assign n7646 = ( x152 & ~x172 ) | ( x152 & n7645 ) | ( ~x172 & n7645 ) ;
  assign n7647 = ~n7644 & n7646 ;
  assign n7648 = n7507 | n7584 ;
  assign n7649 = ( x152 & x172 ) | ( x152 & n7648 ) | ( x172 & n7648 ) ;
  assign n7650 = n7519 & ~n7589 ;
  assign n7651 = ( ~x152 & x172 ) | ( ~x152 & n7650 ) | ( x172 & n7650 ) ;
  assign n7652 = n7649 & n7651 ;
  assign n7653 = n7647 | n7652 ;
  assign n7654 = n7581 & n7653 ;
  assign n7655 = x149 & ~n7654 ;
  assign n7656 = ~n7642 & n7655 ;
  assign n7657 = n7628 & ~n7656 ;
  assign n7658 = n7580 | n7657 ;
  assign n7659 = x232 & n7658 ;
  assign n7660 = ~n4694 & n7401 ;
  assign n7661 = n7393 | n7660 ;
  assign n7662 = ~x232 & n7661 ;
  assign n7663 = x39 | n7662 ;
  assign n7664 = n7659 | n7663 ;
  assign n7665 = ~n7336 & n7664 ;
  assign n7666 = x38 | n7665 ;
  assign n7667 = ~n7263 & n7666 ;
  assign n7668 = x100 | n7667 ;
  assign n7669 = x87 | n7236 ;
  assign n7670 = n7668 & ~n7669 ;
  assign n7671 = x38 & n7248 ;
  assign n7672 = ~x100 & n7671 ;
  assign n7673 = n7236 | n7672 ;
  assign n7674 = n1975 | n7265 ;
  assign n7675 = x87 & n7674 ;
  assign n7676 = ~n7673 & n7675 ;
  assign n7677 = n2004 | n7676 ;
  assign n7678 = n7670 | n7677 ;
  assign n7679 = ~x75 & x92 ;
  assign n7680 = x232 & ~n2162 ;
  assign n7681 = x176 | x299 ;
  assign n7682 = ~n4713 & n7681 ;
  assign n7683 = n7680 & n7682 ;
  assign n7684 = n1983 | n7278 ;
  assign n7685 = n7683 | n7684 ;
  assign n7686 = ~n7674 & n7685 ;
  assign n7687 = n7673 | n7686 ;
  assign n7688 = n7679 & n7687 ;
  assign n7689 = n7237 | n7688 ;
  assign n7690 = n7678 & ~n7689 ;
  assign n7691 = x54 | n7690 ;
  assign n7692 = ~n7251 & n7691 ;
  assign n7693 = x74 | n7692 ;
  assign n7694 = ~n7245 & n7693 ;
  assign n7695 = x55 & ~n7223 ;
  assign n7696 = x54 & n7225 ;
  assign n7697 = x92 | n7216 ;
  assign n7698 = x164 & n5924 ;
  assign n7699 = x38 & ~n7698 ;
  assign n7700 = ~x38 & n7265 ;
  assign n7701 = x100 | n7700 ;
  assign n7702 = n7699 | n7701 ;
  assign n7703 = x87 & ~n7702 ;
  assign n7704 = n7217 | n7703 ;
  assign n7705 = n1924 | n7699 ;
  assign n7706 = x149 & n5924 ;
  assign n7707 = x39 | n7706 ;
  assign n7708 = n7278 | n7707 ;
  assign n7709 = x38 | n7265 ;
  assign n7710 = n7708 & ~n7709 ;
  assign n7711 = ( x38 & ~n7705 ) | ( x38 & n7710 ) | ( ~n7705 & n7710 ) ;
  assign n7712 = n7704 | n7711 ;
  assign n7713 = ~x75 & n7712 ;
  assign n7714 = n7697 | n7713 ;
  assign n7715 = x75 | n7702 ;
  assign n7716 = ~n7218 & n7715 ;
  assign n7717 = ( x54 & n4817 ) | ( x54 & n7716 ) | ( n4817 & n7716 ) ;
  assign n7718 = n7714 & ~n7717 ;
  assign n7719 = n7696 | n7718 ;
  assign n7720 = ~x74 & n7719 ;
  assign n7721 = n7695 & ~n7720 ;
  assign n7722 = n2058 | n7721 ;
  assign n7723 = n7694 | n7722 ;
  assign n7724 = x38 & n7698 ;
  assign n7725 = ~n7219 & n7724 ;
  assign n7726 = n7218 | n7725 ;
  assign n7727 = n7696 | n7726 ;
  assign n7728 = ~x74 & n7727 ;
  assign n7729 = n7223 | n7728 ;
  assign n7730 = n2058 & n7729 ;
  assign n7731 = n2057 | n7730 ;
  assign n7732 = n7219 | n7709 ;
  assign n7733 = n2030 | n7732 ;
  assign n7734 = n2058 & ~n7733 ;
  assign n7735 = n7731 | n7734 ;
  assign n7736 = n7723 & ~n7735 ;
  assign n7737 = n7228 | n7736 ;
  assign n7738 = ( x954 & ~n7210 ) | ( x954 & n7737 ) | ( ~n7210 & n7737 ) ;
  assign n7739 = n4765 & n4988 ;
  assign n7740 = n7285 & n7739 ;
  assign n7741 = ~x174 & n7740 ;
  assign n7742 = x299 | n7741 ;
  assign n7743 = n7264 & n7742 ;
  assign n7744 = n4765 & n7285 ;
  assign n7745 = n5938 & n7744 ;
  assign n7746 = ( x174 & x299 ) | ( x174 & n7745 ) | ( x299 & n7745 ) ;
  assign n7747 = n4997 & n7285 ;
  assign n7748 = n4765 & n7747 ;
  assign n7749 = ( ~x174 & x299 ) | ( ~x174 & n7748 ) | ( x299 & n7748 ) ;
  assign n7750 = n7746 | n7749 ;
  assign n7751 = n7325 & n7750 ;
  assign n7752 = n7743 | n7751 ;
  assign n7753 = ~n4713 & n5938 ;
  assign n7754 = n4721 & n7753 ;
  assign n7755 = x152 & x154 ;
  assign n7756 = n7754 & n7755 ;
  assign n7757 = n4722 & n4997 ;
  assign n7758 = ( x152 & x154 ) | ( x152 & ~n7757 ) | ( x154 & ~n7757 ) ;
  assign n7759 = n4722 & n4988 ;
  assign n7760 = ( ~x152 & x154 ) | ( ~x152 & n7759 ) | ( x154 & n7759 ) ;
  assign n7761 = ~n7758 & n7760 ;
  assign n7762 = n7756 | n7761 ;
  assign n7763 = n7296 & n7762 ;
  assign n7764 = x299 & ~n7763 ;
  assign n7765 = x39 & ~n7764 ;
  assign n7766 = n7752 & n7765 ;
  assign n7767 = x90 & n5886 ;
  assign n7768 = ~n1278 & n4666 ;
  assign n7769 = ~n7767 & n7768 ;
  assign n7770 = x90 | n1590 ;
  assign n7771 = n1278 | n7770 ;
  assign n7772 = n1585 | n7771 ;
  assign n7773 = n1236 | n7772 ;
  assign n7774 = n7365 & ~n7773 ;
  assign n7775 = x70 | n7774 ;
  assign n7776 = n7769 | n7775 ;
  assign n7777 = n1281 | n1864 ;
  assign n7778 = n7776 & ~n7777 ;
  assign n7779 = n7775 & ~n7777 ;
  assign n7780 = n4913 | n7779 ;
  assign n7781 = ~x198 & n7780 ;
  assign n7782 = n7778 | n7781 ;
  assign n7783 = n7448 & n7782 ;
  assign n7784 = n1258 | n7394 ;
  assign n7785 = n7767 | n7784 ;
  assign n7786 = ~n1236 & n7450 ;
  assign n7787 = n4666 | n7786 ;
  assign n7788 = ~n7785 & n7787 ;
  assign n7789 = n1863 | n4713 ;
  assign n7790 = x40 | n7789 ;
  assign n7791 = n7788 & ~n7790 ;
  assign n7792 = ~x183 & n7791 ;
  assign n7793 = x174 | n7792 ;
  assign n7794 = n7783 | n7793 ;
  assign n7795 = n7350 & ~n7772 ;
  assign n7796 = x70 | n7795 ;
  assign n7797 = n7769 | n7796 ;
  assign n7798 = ~n7777 & n7797 ;
  assign n7799 = n4914 | n7798 ;
  assign n7800 = ~n4713 & n7799 ;
  assign n7801 = ( ~x174 & x183 ) | ( ~x174 & n7800 ) | ( x183 & n7800 ) ;
  assign n7802 = n4666 & ~n7785 ;
  assign n7803 = ~n7790 & n7802 ;
  assign n7804 = ( x174 & x183 ) | ( x174 & ~n7803 ) | ( x183 & ~n7803 ) ;
  assign n7805 = ~n7801 & n7804 ;
  assign n7806 = n7794 & ~n7805 ;
  assign n7807 = x193 & ~n7806 ;
  assign n7808 = ~n7396 & n7786 ;
  assign n7809 = ~n1863 & n7808 ;
  assign n7810 = ~n7470 & n7809 ;
  assign n7811 = ~n7510 & n7810 ;
  assign n7812 = x193 | n7811 ;
  assign n7813 = ~n7777 & n7796 ;
  assign n7814 = n4914 | n7813 ;
  assign n7815 = ( ~x174 & n7448 ) | ( ~x174 & n7814 ) | ( n7448 & n7814 ) ;
  assign n7816 = n4914 | n7779 ;
  assign n7817 = ( x174 & n7448 ) | ( x174 & n7816 ) | ( n7448 & n7816 ) ;
  assign n7818 = n7815 & n7817 ;
  assign n7819 = n7812 | n7818 ;
  assign n7820 = ~n7807 & n7819 ;
  assign n7821 = n1536 & ~n4713 ;
  assign n7822 = x180 & n7821 ;
  assign n7823 = x299 | n7822 ;
  assign n7824 = n7820 | n7823 ;
  assign n7825 = x172 & n7778 ;
  assign n7826 = n4957 | n7779 ;
  assign n7827 = x152 | n7826 ;
  assign n7828 = n7825 | n7827 ;
  assign n7829 = n4957 | n7813 ;
  assign n7830 = x172 & n7798 ;
  assign n7831 = x152 & ~n7830 ;
  assign n7832 = ~n7829 & n7831 ;
  assign n7833 = x149 & ~n4713 ;
  assign n7834 = ~n7832 & n7833 ;
  assign n7835 = n7828 & n7834 ;
  assign n7836 = ~x152 & n7791 ;
  assign n7837 = n7803 | n7836 ;
  assign n7838 = x172 & n7837 ;
  assign n7839 = x152 | x172 ;
  assign n7840 = n7810 & ~n7839 ;
  assign n7841 = n7838 | n7840 ;
  assign n7842 = ~x149 & n7841 ;
  assign n7843 = x158 & n7821 ;
  assign n7844 = x299 & ~n7843 ;
  assign n7845 = ~n7842 & n7844 ;
  assign n7846 = ~n7835 & n7845 ;
  assign n7847 = n5788 & ~n7846 ;
  assign n7848 = n7824 & n7847 ;
  assign n7849 = n7766 | n7848 ;
  assign n7850 = ~x38 & n7849 ;
  assign n7851 = x87 | n7263 ;
  assign n7852 = n7850 | n7851 ;
  assign n7853 = x87 & ~n7671 ;
  assign n7854 = x100 | n7853 ;
  assign n7855 = n7852 & ~n7854 ;
  assign n7856 = n7236 | n7855 ;
  assign n7857 = ~n2004 & n7856 ;
  assign n7858 = x38 | x87 ;
  assign n7859 = x100 | n7858 ;
  assign n7860 = n7683 & ~n7859 ;
  assign n7861 = ~n4660 & n7860 ;
  assign n7862 = n7673 | n7861 ;
  assign n7863 = n7679 & n7862 ;
  assign n7864 = n7237 | n7863 ;
  assign n7865 = n7857 | n7864 ;
  assign n7866 = ~x54 & n7865 ;
  assign n7867 = n7251 | n7866 ;
  assign n7868 = ~x74 & n7867 ;
  assign n7869 = n7245 | n7868 ;
  assign n7870 = ~n4660 & n7706 ;
  assign n7871 = x38 | n7870 ;
  assign n7872 = ~n7705 & n7871 ;
  assign n7873 = n6015 & n7724 ;
  assign n7874 = n7217 | n7873 ;
  assign n7875 = n7872 | n7874 ;
  assign n7876 = ~x75 & n7875 ;
  assign n7877 = n7697 | n7876 ;
  assign n7878 = ( x54 & n4817 ) | ( x54 & ~n7726 ) | ( n4817 & ~n7726 ) ;
  assign n7879 = n7877 & ~n7878 ;
  assign n7880 = n7696 | n7879 ;
  assign n7881 = ~x74 & n7880 ;
  assign n7882 = n7695 & ~n7881 ;
  assign n7883 = n2058 | n7882 ;
  assign n7884 = n7869 & ~n7883 ;
  assign n7885 = n7731 | n7884 ;
  assign n7886 = ~n7228 & n7885 ;
  assign n7887 = ( x954 & n7210 ) | ( x954 & ~n7886 ) | ( n7210 & ~n7886 ) ;
  assign n7888 = n7738 | n7887 ;
  assign n7889 = ( ~x33 & x954 ) | ( ~x33 & n7886 ) | ( x954 & n7886 ) ;
  assign n7890 = ( x33 & x954 ) | ( x33 & ~n7737 ) | ( x954 & ~n7737 ) ;
  assign n7891 = n7889 & n7890 ;
  assign n7892 = n7888 & ~n7891 ;
  assign n7893 = ( x162 & x197 ) | ( x162 & ~n7212 ) | ( x197 & ~n7212 ) ;
  assign n7894 = ( x162 & x197 ) | ( x162 & n7212 ) | ( x197 & n7212 ) ;
  assign n7895 = ( n7212 & n7893 ) | ( n7212 & ~n7894 ) | ( n7893 & ~n7894 ) ;
  assign n7896 = ~n4713 & n7895 ;
  assign n7897 = x232 & n7896 ;
  assign n7898 = n7219 & n7897 ;
  assign n7899 = x167 & n5924 ;
  assign n7900 = ~n7219 & n7899 ;
  assign n7901 = n7898 | n7900 ;
  assign n7902 = x74 | n7901 ;
  assign n7903 = x148 & n7220 ;
  assign n7904 = x74 & ~n7903 ;
  assign n7905 = ~n7898 & n7904 ;
  assign n7906 = n7902 & ~n7905 ;
  assign n7907 = n2057 & n7906 ;
  assign n7908 = x54 | n7898 ;
  assign n7909 = x38 & n7900 ;
  assign n7910 = n7908 | n7909 ;
  assign n7911 = x74 | n7910 ;
  assign n7912 = n7906 & n7911 ;
  assign n7913 = n2058 & ~n7912 ;
  assign n7914 = n2057 | n7913 ;
  assign n7915 = x299 & ~n7896 ;
  assign n7916 = x232 & x299 ;
  assign n7917 = x140 & x145 ;
  assign n7918 = x140 | x145 ;
  assign n7919 = ~n7917 & n7918 ;
  assign n7920 = n7232 & ~n7919 ;
  assign n7921 = n7231 | n7917 ;
  assign n7922 = ~n4713 & n7918 ;
  assign n7923 = ~n7921 & n7922 ;
  assign n7924 = n7920 | n7923 ;
  assign n7925 = ( x232 & n7916 ) | ( x232 & n7924 ) | ( n7916 & n7924 ) ;
  assign n7926 = ~n7915 & n7925 ;
  assign n7927 = x100 & ~n7926 ;
  assign n7928 = x75 & ~n7926 ;
  assign n7929 = n7927 | n7928 ;
  assign n7930 = x141 & ~x299 ;
  assign n7931 = x148 & x299 ;
  assign n7932 = n7930 | n7931 ;
  assign n7933 = n5924 & n7932 ;
  assign n7934 = n7219 | n7933 ;
  assign n7935 = ~n7929 & n7934 ;
  assign n7936 = x74 & ~n7935 ;
  assign n7937 = x55 | n7936 ;
  assign n7938 = x188 & ~x299 ;
  assign n7939 = x167 & x299 ;
  assign n7940 = n7938 | n7939 ;
  assign n7941 = n5924 & n7940 ;
  assign n7942 = x100 | n7941 ;
  assign n7943 = x75 | n7942 ;
  assign n7944 = ~n7929 & n7943 ;
  assign n7945 = x54 & ~n7944 ;
  assign n7946 = x181 & n7821 ;
  assign n7947 = x299 | n7946 ;
  assign n7948 = x140 & n4713 ;
  assign n7949 = ~x142 & n7803 ;
  assign n7950 = x140 | n7949 ;
  assign n7951 = ~x142 & n7798 ;
  assign n7952 = x140 & ~n7951 ;
  assign n7953 = ~n7814 & n7952 ;
  assign n7954 = n7950 & ~n7953 ;
  assign n7955 = ( x144 & n7948 ) | ( x144 & ~n7954 ) | ( n7948 & ~n7954 ) ;
  assign n7956 = ~x142 & n7778 ;
  assign n7957 = x140 & ~n7816 ;
  assign n7958 = ~n7956 & n7957 ;
  assign n7959 = ( x140 & x142 ) | ( x140 & n7810 ) | ( x142 & n7810 ) ;
  assign n7960 = ( x140 & ~x142 ) | ( x140 & n7791 ) | ( ~x142 & n7791 ) ;
  assign n7961 = n7959 | n7960 ;
  assign n7962 = ~n7958 & n7961 ;
  assign n7963 = ( x144 & ~n7948 ) | ( x144 & n7962 ) | ( ~n7948 & n7962 ) ;
  assign n7964 = ~n7955 & n7963 ;
  assign n7965 = n7947 | n7964 ;
  assign n7966 = ~x146 & x161 ;
  assign n7967 = n7803 & n7966 ;
  assign n7968 = ( x146 & x161 ) | ( x146 & ~n7810 ) | ( x161 & ~n7810 ) ;
  assign n7969 = ( x146 & ~x161 ) | ( x146 & n7791 ) | ( ~x161 & n7791 ) ;
  assign n7970 = ~n7968 & n7969 ;
  assign n7971 = n7967 | n7970 ;
  assign n7972 = ~x162 & n7971 ;
  assign n7973 = x162 & ~n4713 ;
  assign n7974 = ~x159 & x299 ;
  assign n7975 = x159 & x299 ;
  assign n7976 = ~x162 & n7821 ;
  assign n7977 = n7975 & ~n7976 ;
  assign n7978 = n7974 | n7977 ;
  assign n7979 = ~n7973 & n7978 ;
  assign n7980 = ~x146 & n7798 ;
  assign n7981 = n7829 | n7980 ;
  assign n7982 = x159 & n1536 ;
  assign n7983 = x299 & ~n7982 ;
  assign n7984 = ( x161 & n7981 ) | ( x161 & ~n7983 ) | ( n7981 & ~n7983 ) ;
  assign n7985 = ~x146 & n7778 ;
  assign n7986 = n7826 | n7985 ;
  assign n7987 = ( x161 & n7983 ) | ( x161 & ~n7986 ) | ( n7983 & ~n7986 ) ;
  assign n7988 = ~n7984 & n7987 ;
  assign n7989 = n7979 | n7988 ;
  assign n7990 = ~n7972 & n7989 ;
  assign n7991 = x232 & ~n7990 ;
  assign n7992 = n7965 & n7991 ;
  assign n7993 = n1925 | n7992 ;
  assign n7994 = x188 & n7253 ;
  assign n7995 = x167 | n7994 ;
  assign n7996 = x188 | n7259 ;
  assign n7997 = x167 & x188 ;
  assign n7998 = ~n7256 & n7997 ;
  assign n7999 = n7996 & ~n7998 ;
  assign n8000 = n7995 & n7999 ;
  assign n8001 = x38 & ~n8000 ;
  assign n8002 = ~x38 & x155 ;
  assign n8003 = ( x161 & n7296 ) | ( x161 & n7757 ) | ( n7296 & n7757 ) ;
  assign n8004 = ( ~x161 & n7296 ) | ( ~x161 & n7754 ) | ( n7296 & n7754 ) ;
  assign n8005 = n8003 & n8004 ;
  assign n8006 = n8002 & ~n8005 ;
  assign n8007 = x38 | x155 ;
  assign n8008 = ~x161 & n7296 ;
  assign n8009 = n7759 & n8008 ;
  assign n8010 = n8007 | n8009 ;
  assign n8011 = ~n8006 & n8010 ;
  assign n8012 = x299 & ~n8011 ;
  assign n8013 = x177 | x299 ;
  assign n8014 = ~x144 & n7740 ;
  assign n8015 = n8013 | n8014 ;
  assign n8016 = x232 & n8015 ;
  assign n8017 = x177 & ~x299 ;
  assign n8018 = ( x144 & n7745 ) | ( x144 & ~n8017 ) | ( n7745 & ~n8017 ) ;
  assign n8019 = ( x144 & ~n7748 ) | ( x144 & n8017 ) | ( ~n7748 & n8017 ) ;
  assign n8020 = ~n8018 & n8019 ;
  assign n8021 = n8016 & ~n8020 ;
  assign n8022 = x38 | n8021 ;
  assign n8023 = ~n8012 & n8022 ;
  assign n8024 = x39 & ~n8023 ;
  assign n8025 = n8001 | n8024 ;
  assign n8026 = n7993 & ~n8025 ;
  assign n8027 = x100 | n8026 ;
  assign n8028 = ~n7927 & n8027 ;
  assign n8029 = x87 | n8028 ;
  assign n8030 = n1975 & n7942 ;
  assign n8031 = ~n7927 & n8030 ;
  assign n8032 = x87 & ~n8031 ;
  assign n8033 = n8029 & ~n8032 ;
  assign n8034 = n2004 | n8033 ;
  assign n8035 = x38 & n7940 ;
  assign n8036 = x155 & x299 ;
  assign n8037 = n8017 | n8036 ;
  assign n8038 = ~n1925 & n8037 ;
  assign n8039 = ~n1860 & n8038 ;
  assign n8040 = n8035 | n8039 ;
  assign n8041 = n5924 & n8040 ;
  assign n8042 = x100 | n8041 ;
  assign n8043 = ~n7927 & n8042 ;
  assign n8044 = x87 | n8043 ;
  assign n8045 = ~n8032 & n8044 ;
  assign n8046 = n7679 & ~n8045 ;
  assign n8047 = n7928 | n8046 ;
  assign n8048 = n8034 & ~n8047 ;
  assign n8049 = x54 | n8048 ;
  assign n8050 = ~n7945 & n8049 ;
  assign n8051 = x74 | n8050 ;
  assign n8052 = ~n7937 & n8051 ;
  assign n8053 = x55 & ~n7905 ;
  assign n8054 = x54 & ~n7901 ;
  assign n8055 = x38 & n7899 ;
  assign n8056 = ~x92 & x162 ;
  assign n8057 = n5788 & n8056 ;
  assign n8058 = ~n7858 & n8057 ;
  assign n8059 = ~n4738 & n8058 ;
  assign n8060 = n8055 | n8059 ;
  assign n8061 = ~n7219 & n8060 ;
  assign n8062 = n7908 | n8061 ;
  assign n8063 = ~n8054 & n8062 ;
  assign n8064 = x74 | n8063 ;
  assign n8065 = n8053 & n8064 ;
  assign n8066 = n2058 | n8065 ;
  assign n8067 = n8052 | n8066 ;
  assign n8068 = ~n7914 & n8067 ;
  assign n8069 = n7907 | n8068 ;
  assign n8070 = x33 | x954 ;
  assign n8071 = ( ~x34 & n8069 ) | ( ~x34 & n8070 ) | ( n8069 & n8070 ) ;
  assign n8072 = n2058 & n7733 ;
  assign n8073 = n2057 | n8072 ;
  assign n8074 = n7914 & n8073 ;
  assign n8075 = ( x140 & x142 ) | ( x140 & ~n7426 ) | ( x142 & ~n7426 ) ;
  assign n8076 = ( ~x140 & x142 ) | ( ~x140 & n7505 ) | ( x142 & n7505 ) ;
  assign n8077 = ~n8075 & n8076 ;
  assign n8078 = ( x140 & ~x142 ) | ( x140 & n7442 ) | ( ~x142 & n7442 ) ;
  assign n8079 = ( x140 & x142 ) | ( x140 & n7509 ) | ( x142 & n7509 ) ;
  assign n8080 = n8078 & n8079 ;
  assign n8081 = n8077 | n8080 ;
  assign n8082 = ( x144 & x181 ) | ( x144 & n8081 ) | ( x181 & n8081 ) ;
  assign n8083 = x142 | n7562 ;
  assign n8084 = n7420 | n7613 ;
  assign n8085 = ~n4713 & n8084 ;
  assign n8086 = x142 & ~n8085 ;
  assign n8087 = ~n7508 & n8086 ;
  assign n8088 = x140 | n8087 ;
  assign n8089 = n8083 & ~n8088 ;
  assign n8090 = x142 | n7550 ;
  assign n8091 = x142 & ~n7637 ;
  assign n8092 = ~n7508 & n8091 ;
  assign n8093 = x140 & ~n8092 ;
  assign n8094 = n8090 & n8093 ;
  assign n8095 = n8089 | n8094 ;
  assign n8096 = ( x144 & ~x181 ) | ( x144 & n8095 ) | ( ~x181 & n8095 ) ;
  assign n8097 = n8082 | n8096 ;
  assign n8098 = ~x299 & n8097 ;
  assign n8099 = ( x140 & x142 ) | ( x140 & ~n7474 ) | ( x142 & ~n7474 ) ;
  assign n8100 = ( ~x140 & x142 ) | ( ~x140 & n7542 ) | ( x142 & n7542 ) ;
  assign n8101 = ~n8099 & n8100 ;
  assign n8102 = ( x140 & ~x142 ) | ( x140 & n7468 ) | ( ~x142 & n7468 ) ;
  assign n8103 = ( x140 & x142 ) | ( x140 & n7520 ) | ( x142 & n7520 ) ;
  assign n8104 = n8102 & n8103 ;
  assign n8105 = n8101 | n8104 ;
  assign n8106 = ( ~x144 & x181 ) | ( ~x144 & n8105 ) | ( x181 & n8105 ) ;
  assign n8107 = x142 | n7568 ;
  assign n8108 = x142 & ~n7459 ;
  assign n8109 = ~n7508 & n8108 ;
  assign n8110 = x140 & ~n8109 ;
  assign n8111 = n8107 & n8110 ;
  assign n8112 = ( x140 & x142 ) | ( x140 & ~n7403 ) | ( x142 & ~n7403 ) ;
  assign n8113 = ( ~x140 & x142 ) | ( ~x140 & n7573 ) | ( x142 & n7573 ) ;
  assign n8114 = ~n8112 & n8113 ;
  assign n8115 = n8111 | n8114 ;
  assign n8116 = ( x144 & x181 ) | ( x144 & ~n8115 ) | ( x181 & ~n8115 ) ;
  assign n8117 = ~n8106 & n8116 ;
  assign n8118 = n8098 & ~n8117 ;
  assign n8119 = ( x146 & x161 ) | ( x146 & ~n7638 ) | ( x161 & ~n7638 ) ;
  assign n8120 = ( x146 & ~x161 ) | ( x146 & n7629 ) | ( ~x161 & n7629 ) ;
  assign n8121 = ~n8119 & n8120 ;
  assign n8122 = ( x146 & x161 ) | ( x146 & n7631 ) | ( x161 & n7631 ) ;
  assign n8123 = ( ~x146 & x161 ) | ( ~x146 & n7634 ) | ( x161 & n7634 ) ;
  assign n8124 = n8122 & n8123 ;
  assign n8125 = n8121 | n8124 ;
  assign n8126 = x162 & n8125 ;
  assign n8127 = x162 | n7589 ;
  assign n8128 = ( ~x146 & x161 ) | ( ~x146 & n7583 ) | ( x161 & n7583 ) ;
  assign n8129 = ( x146 & x161 ) | ( x146 & ~n7615 ) | ( x161 & ~n7615 ) ;
  assign n8130 = ~n8128 & n8129 ;
  assign n8131 = n8127 | n8130 ;
  assign n8132 = ( x146 & x161 ) | ( x146 & n7623 ) | ( x161 & n7623 ) ;
  assign n8133 = ( x146 & ~x161 ) | ( x146 & n7620 ) | ( ~x161 & n7620 ) ;
  assign n8134 = n8132 | n8133 ;
  assign n8135 = ~n8131 & n8134 ;
  assign n8136 = n8126 | n8135 ;
  assign n8137 = n7974 & n8136 ;
  assign n8138 = ( x146 & x161 ) | ( x146 & ~n7645 ) | ( x161 & ~n7645 ) ;
  assign n8139 = ( x146 & ~x161 ) | ( x146 & n7648 ) | ( ~x161 & n7648 ) ;
  assign n8140 = ~n8138 & n8139 ;
  assign n8141 = x162 & ~n8140 ;
  assign n8142 = ( x146 & x161 ) | ( x146 & n7650 ) | ( x161 & n7650 ) ;
  assign n8143 = ( ~x146 & x161 ) | ( ~x146 & n7643 ) | ( x161 & n7643 ) ;
  assign n8144 = n8142 & n8143 ;
  assign n8145 = n8141 & ~n8144 ;
  assign n8146 = ( x146 & x161 ) | ( x146 & n7605 ) | ( x161 & n7605 ) ;
  assign n8147 = ( ~x146 & x161 ) | ( ~x146 & n7587 ) | ( x161 & n7587 ) ;
  assign n8148 = n8146 & n8147 ;
  assign n8149 = x162 | n8148 ;
  assign n8150 = ( x146 & x161 ) | ( x146 & ~n7592 ) | ( x161 & ~n7592 ) ;
  assign n8151 = ( x146 & ~x161 ) | ( x146 & n7600 ) | ( ~x161 & n7600 ) ;
  assign n8152 = ~n8150 & n8151 ;
  assign n8153 = n8149 | n8152 ;
  assign n8154 = n7975 & n8153 ;
  assign n8155 = ~n8145 & n8154 ;
  assign n8156 = n8137 | n8155 ;
  assign n8157 = n8118 | n8156 ;
  assign n8158 = x232 & n8157 ;
  assign n8159 = n7662 | n8158 ;
  assign n8160 = ~n1925 & n8159 ;
  assign n8161 = x144 & ~n7330 ;
  assign n8162 = x144 | n7287 ;
  assign n8163 = n7321 | n8162 ;
  assign n8164 = ~n8013 & n8163 ;
  assign n8165 = ~n8161 & n8164 ;
  assign n8166 = n7287 | n7292 ;
  assign n8167 = n8017 & n8162 ;
  assign n8168 = n8166 & n8167 ;
  assign n8169 = n8165 | n8168 ;
  assign n8170 = x232 & n8169 ;
  assign n8171 = n7333 | n8170 ;
  assign n8172 = ~x38 & n8171 ;
  assign n8173 = x161 | n7302 ;
  assign n8174 = n7307 & n8173 ;
  assign n8175 = n7296 & ~n8174 ;
  assign n8176 = n7298 & ~n8007 ;
  assign n8177 = ~n8175 & n8176 ;
  assign n8178 = x161 & n7310 ;
  assign n8179 = ~n7284 & n7296 ;
  assign n8180 = ~n8178 & n8179 ;
  assign n8181 = n7298 & n8002 ;
  assign n8182 = ~n8180 & n8181 ;
  assign n8183 = n8177 | n8182 ;
  assign n8184 = x232 & n8183 ;
  assign n8185 = n8172 | n8184 ;
  assign n8186 = x39 & n8185 ;
  assign n8187 = x87 | n8001 ;
  assign n8188 = n8186 | n8187 ;
  assign n8189 = n8160 | n8188 ;
  assign n8190 = x38 & ~n7941 ;
  assign n8191 = n7700 | n8190 ;
  assign n8192 = x87 & ~n8191 ;
  assign n8193 = x100 | n8192 ;
  assign n8194 = n8189 & ~n8193 ;
  assign n8195 = n7927 | n8194 ;
  assign n8196 = ~n2004 & n8195 ;
  assign n8197 = x38 | n8037 ;
  assign n8198 = n5924 & n8197 ;
  assign n8199 = n7684 | n8198 ;
  assign n8200 = ~n8191 & n8199 ;
  assign n8201 = x100 | n8200 ;
  assign n8202 = ~n7927 & n8201 ;
  assign n8203 = n7679 & ~n8202 ;
  assign n8204 = n7928 | n8203 ;
  assign n8205 = n8196 | n8204 ;
  assign n8206 = ~x54 & n8205 ;
  assign n8207 = n7945 | n8206 ;
  assign n8208 = ~x74 & n8207 ;
  assign n8209 = n7937 | n8208 ;
  assign n8210 = n7732 & ~n7910 ;
  assign n8211 = n4817 & ~n8210 ;
  assign n8212 = ( x75 & x92 ) | ( x75 & ~n7897 ) | ( x92 & ~n7897 ) ;
  assign n8213 = x100 & ~n7897 ;
  assign n8214 = n7684 | n7973 ;
  assign n8215 = ~n7709 & n8214 ;
  assign n8216 = x100 | n8215 ;
  assign n8217 = x232 | n7684 ;
  assign n8218 = n8216 & n8217 ;
  assign n8219 = n8055 | n8218 ;
  assign n8220 = ~n8213 & n8219 ;
  assign n8221 = ( x75 & ~x92 ) | ( x75 & n8220 ) | ( ~x92 & n8220 ) ;
  assign n8222 = ~n8212 & n8221 ;
  assign n8223 = n8211 | n8222 ;
  assign n8224 = ~n8054 & n8223 ;
  assign n8225 = x74 | n8224 ;
  assign n8226 = n8053 & n8225 ;
  assign n8227 = n2058 | n8226 ;
  assign n8228 = n8209 & ~n8227 ;
  assign n8229 = n8074 | n8228 ;
  assign n8230 = ~n7907 & n8229 ;
  assign n8231 = ( x34 & n8070 ) | ( x34 & ~n8230 ) | ( n8070 & ~n8230 ) ;
  assign n8232 = n8071 & n8231 ;
  assign n8233 = ~x34 & n7208 ;
  assign n8234 = ( ~n8069 & n8070 ) | ( ~n8069 & n8233 ) | ( n8070 & n8233 ) ;
  assign n8235 = ( n8070 & n8230 ) | ( n8070 & ~n8233 ) | ( n8230 & ~n8233 ) ;
  assign n8236 = n8234 | n8235 ;
  assign n8237 = ~n8232 & n8236 ;
  assign n8238 = x24 | n5800 ;
  assign n8239 = x54 & n8238 ;
  assign n8240 = n2058 | n5073 ;
  assign n8241 = n8239 | n8240 ;
  assign n8242 = x137 & n7115 ;
  assign n8243 = n1287 & n1690 ;
  assign n8244 = n5950 & ~n8243 ;
  assign n8245 = x683 & n8244 ;
  assign n8246 = x252 & n4795 ;
  assign n8247 = ~n8245 & n8246 ;
  assign n8248 = ~n5924 & n8247 ;
  assign n8249 = x146 & n5922 ;
  assign n8250 = x142 & n5921 ;
  assign n8251 = n8249 | n8250 ;
  assign n8252 = ~n8247 & n8251 ;
  assign n8253 = ( n5923 & n8248 ) | ( n5923 & ~n8252 ) | ( n8248 & ~n8252 ) ;
  assign n8254 = n7118 | n8253 ;
  assign n8255 = ~n4784 & n7120 ;
  assign n8256 = ~n8247 & n8255 ;
  assign n8257 = n8254 & ~n8256 ;
  assign n8258 = n7117 & ~n8257 ;
  assign n8259 = n8242 | n8258 ;
  assign n8260 = n2364 & n8259 ;
  assign n8261 = ~x90 & n4665 ;
  assign n8262 = x93 | n8261 ;
  assign n8263 = ~n4664 & n8262 ;
  assign n8264 = x35 | n8263 ;
  assign n8265 = x35 & ~n1604 ;
  assign n8266 = n7164 | n8265 ;
  assign n8267 = n8264 & ~n8266 ;
  assign n8268 = ~x32 & n8267 ;
  assign n8269 = x32 & ~x93 ;
  assign n8270 = ~n7126 & n8269 ;
  assign n8271 = ~n5886 & n8270 ;
  assign n8272 = n8268 | n8271 ;
  assign n8273 = x95 | n4694 ;
  assign n8274 = n8272 & ~n8273 ;
  assign n8275 = n1299 | n8267 ;
  assign n8276 = x1082 & ~n1863 ;
  assign n8277 = n8275 & n8276 ;
  assign n8278 = n4694 & n8264 ;
  assign n8279 = x137 | n4694 ;
  assign n8280 = x122 | n4800 ;
  assign n8281 = ( n6153 & n8279 ) | ( n6153 & ~n8280 ) | ( n8279 & ~n8280 ) ;
  assign n8282 = n1288 & n5984 ;
  assign n8283 = ( ~n6153 & n8279 ) | ( ~n6153 & n8282 ) | ( n8279 & n8282 ) ;
  assign n8284 = n8281 & n8283 ;
  assign n8285 = n8278 | n8284 ;
  assign n8286 = ~n1255 & n7163 ;
  assign n8287 = n8264 | n8286 ;
  assign n8288 = n1863 | n8266 ;
  assign n8289 = n8287 & ~n8288 ;
  assign n8290 = n8285 & n8289 ;
  assign n8291 = x38 | n8290 ;
  assign n8292 = n8277 | n8291 ;
  assign n8293 = n8274 | n8292 ;
  assign n8294 = x38 & n7192 ;
  assign n8295 = n5818 | n8294 ;
  assign n8296 = n8293 & ~n8295 ;
  assign n8297 = n8260 | n8296 ;
  assign n8298 = ~n1998 & n8297 ;
  assign n8299 = x137 & ~n7136 ;
  assign n8300 = ~n4804 & n8299 ;
  assign n8301 = n7194 | n8300 ;
  assign n8302 = n7197 & n8301 ;
  assign n8303 = ~n7192 & n8302 ;
  assign n8304 = n8298 | n8303 ;
  assign n8305 = ~n4817 & n8304 ;
  assign n8306 = ( x54 & ~n8241 ) | ( x54 & n8305 ) | ( ~n8241 & n8305 ) ;
  assign n8307 = ( ~x57 & x59 ) | ( ~x57 & n8306 ) | ( x59 & n8306 ) ;
  assign n8308 = n2033 | n2058 ;
  assign n8309 = n7192 | n8308 ;
  assign n8310 = x55 | n8309 ;
  assign n8311 = ( x57 & x59 ) | ( x57 & n8310 ) | ( x59 & n8310 ) ;
  assign n8312 = n8307 & ~n8311 ;
  assign n8313 = n1328 | n1590 ;
  assign n8314 = x83 | n1399 ;
  assign n8315 = x65 | n1243 ;
  assign n8316 = n1236 | n8315 ;
  assign n8317 = n7266 | n8316 ;
  assign n8318 = x69 | n8317 ;
  assign n8319 = x67 | x71 ;
  assign n8320 = x36 & ~x103 ;
  assign n8321 = ~n8319 & n8320 ;
  assign n8322 = ~n8318 & n8321 ;
  assign n8323 = ~n8314 & n8322 ;
  assign n8324 = ~n8313 & n8323 ;
  assign n8325 = ~x58 & n5956 ;
  assign n8326 = n8324 | n8325 ;
  assign n8327 = n1255 | n4904 ;
  assign n8328 = n4695 | n8327 ;
  assign n8329 = n2030 | n6785 ;
  assign n8330 = n2111 | n8329 ;
  assign n8331 = x92 | n8330 ;
  assign n8332 = n8328 | n8331 ;
  assign n8333 = n4800 & ~n8332 ;
  assign n8334 = n8326 & n8333 ;
  assign n8335 = x81 | n1351 ;
  assign n8336 = n4904 | n7483 ;
  assign n8337 = n1268 | n8336 ;
  assign n8338 = n1295 | n8337 ;
  assign n8339 = x71 | n1236 ;
  assign n8340 = x104 | n1221 ;
  assign n8341 = n8339 | n8340 ;
  assign n8342 = x45 | x73 ;
  assign n8343 = n7143 | n8342 ;
  assign n8344 = x48 | x65 ;
  assign n8345 = x82 | x84 ;
  assign n8346 = x89 & ~n8345 ;
  assign n8347 = ~n8344 & n8346 ;
  assign n8348 = ~n8343 & n8347 ;
  assign n8349 = ~n7355 & n8348 ;
  assign n8350 = ~n8341 & n8349 ;
  assign n8351 = x332 & n8350 ;
  assign n8352 = x64 | n8351 ;
  assign n8353 = x102 | n1245 ;
  assign n8354 = x39 | x841 ;
  assign n8355 = n8353 | n8354 ;
  assign n8356 = n8352 & ~n8355 ;
  assign n8357 = ~n8338 & n8356 ;
  assign n8358 = ~n8335 & n8357 ;
  assign n8359 = n2032 | n6785 ;
  assign n8360 = ( x38 & n8358 ) | ( x38 & ~n8359 ) | ( n8358 & ~n8359 ) ;
  assign n8361 = x39 | n1864 ;
  assign n8362 = x24 & ~n8361 ;
  assign n8363 = ~n1260 & n8362 ;
  assign n8364 = ( x38 & n8359 ) | ( x38 & ~n8363 ) | ( n8359 & ~n8363 ) ;
  assign n8365 = n8360 & ~n8364 ;
  assign n8366 = x38 | n8359 ;
  assign n8367 = ( x835 & n1692 ) | ( x835 & n4727 ) | ( n1692 & n4727 ) ;
  assign n8368 = n4726 & ~n8367 ;
  assign n8369 = n4744 & ~n8368 ;
  assign n8370 = x1093 & n8369 ;
  assign n8371 = n4977 & ~n4981 ;
  assign n8372 = ~n8370 & n8371 ;
  assign n8373 = ~x215 & n8372 ;
  assign n8374 = ~n4751 & n8369 ;
  assign n8375 = n8371 & ~n8374 ;
  assign n8376 = ( ~x299 & n4721 ) | ( ~x299 & n8375 ) | ( n4721 & n8375 ) ;
  assign n8377 = n4714 & n8369 ;
  assign n8378 = n8371 & ~n8377 ;
  assign n8379 = ( x299 & n4721 ) | ( x299 & ~n8378 ) | ( n4721 & ~n8378 ) ;
  assign n8380 = ~n8376 & n8379 ;
  assign n8381 = ~n8373 & n8380 ;
  assign n8382 = x786 & ~x1082 ;
  assign n8383 = ~x223 & n8372 ;
  assign n8384 = ( x299 & n4764 ) | ( x299 & n8375 ) | ( n4764 & n8375 ) ;
  assign n8385 = ( x299 & ~n4764 ) | ( x299 & n8378 ) | ( ~n4764 & n8378 ) ;
  assign n8386 = n8384 | n8385 ;
  assign n8387 = n8383 | n8386 ;
  assign n8388 = ~n8382 & n8387 ;
  assign n8389 = ~n8381 & n8388 ;
  assign n8390 = n4343 & n4723 ;
  assign n8391 = ~n2213 & n4766 ;
  assign n8392 = n8390 | n8391 ;
  assign n8393 = n4800 & n8382 ;
  assign n8394 = n8392 & n8393 ;
  assign n8395 = n4982 & n8394 ;
  assign n8396 = n8389 | n8395 ;
  assign n8397 = x39 & n8396 ;
  assign n8398 = n4694 & n4912 ;
  assign n8399 = x35 & n4908 ;
  assign n8400 = n1295 | n8399 ;
  assign n8401 = ( n1271 & n4695 ) | ( n1271 & n8400 ) | ( n4695 & n8400 ) ;
  assign n8402 = n4695 | n8400 ;
  assign n8403 = ( n1242 & n8401 ) | ( n1242 & n8402 ) | ( n8401 & n8402 ) ;
  assign n8404 = n1492 | n8403 ;
  assign n8405 = n1333 | n1587 ;
  assign n8406 = n7147 | n7152 ;
  assign n8407 = n7352 | n8406 ;
  assign n8408 = n7148 | n7356 ;
  assign n8409 = x65 | x69 ;
  assign n8410 = n8408 | n8409 ;
  assign n8411 = x48 & ~x49 ;
  assign n8412 = x68 | x82 ;
  assign n8413 = n8411 & ~n8412 ;
  assign n8414 = ~n8342 & n8413 ;
  assign n8415 = ~n8410 & n8414 ;
  assign n8416 = ~n8407 & n8415 ;
  assign n8417 = ~n8341 & n8416 ;
  assign n8418 = x841 | n1215 ;
  assign n8419 = n1326 | n8418 ;
  assign n8420 = x97 | n8419 ;
  assign n8421 = n8417 & ~n8420 ;
  assign n8422 = ~n8405 & n8421 ;
  assign n8423 = ~x46 & x108 ;
  assign n8424 = ~n1250 & n8423 ;
  assign n8425 = ~n1331 & n8424 ;
  assign n8426 = ~n1242 & n8425 ;
  assign n8427 = x47 | n8426 ;
  assign n8428 = n8422 | n8427 ;
  assign n8429 = x986 | n4800 ;
  assign n8430 = x252 & n8429 ;
  assign n8431 = x314 & ~n8430 ;
  assign n8432 = ~n4680 & n8431 ;
  assign n8433 = n8428 & n8432 ;
  assign n8434 = x47 | x841 ;
  assign n8435 = n8417 & ~n8434 ;
  assign n8436 = ~n1242 & n1319 ;
  assign n8437 = n8435 | n8436 ;
  assign n8438 = n1251 | n1311 ;
  assign n8439 = n8431 | n8438 ;
  assign n8440 = n8437 & ~n8439 ;
  assign n8441 = n8433 | n8440 ;
  assign n8442 = ~n5899 & n8441 ;
  assign n8443 = ( x35 & ~n8404 ) | ( x35 & n8442 ) | ( ~n8404 & n8442 ) ;
  assign n8444 = n8398 | n8443 ;
  assign n8445 = ~n4658 & n8444 ;
  assign n8446 = n8397 | n8445 ;
  assign n8447 = ~n8366 & n8446 ;
  assign n8448 = x81 | n1242 ;
  assign n8449 = ~x93 & x102 ;
  assign n8450 = ~n1269 & n8449 ;
  assign n8451 = ~n1245 & n8450 ;
  assign n8452 = ~n4695 & n8451 ;
  assign n8453 = ~n1268 & n8452 ;
  assign n8454 = ~n8448 & n8453 ;
  assign n8455 = ~n4904 & n8454 ;
  assign n8456 = ( x1082 & n8331 ) | ( x1082 & ~n8455 ) | ( n8331 & ~n8455 ) ;
  assign n8457 = x40 | n8454 ;
  assign n8458 = n1863 | n2131 ;
  assign n8459 = x40 | n1863 ;
  assign n8460 = ( n1271 & n8458 ) | ( n1271 & n8459 ) | ( n8458 & n8459 ) ;
  assign n8461 = n8458 | n8459 ;
  assign n8462 = ( n1242 & n8460 ) | ( n1242 & n8461 ) | ( n8460 & n8461 ) ;
  assign n8463 = n8457 & ~n8462 ;
  assign n8464 = ( x1082 & ~n8331 ) | ( x1082 & n8463 ) | ( ~n8331 & n8463 ) ;
  assign n8465 = ~n8456 & n8464 ;
  assign n8466 = x166 | n4713 ;
  assign n8467 = x161 & ~n8466 ;
  assign n8468 = ~x152 & n8467 ;
  assign n8469 = x39 & x232 ;
  assign n8470 = n8468 & n8469 ;
  assign n8471 = x41 | x72 ;
  assign n8472 = ~x39 & n8471 ;
  assign n8473 = x72 | n8472 ;
  assign n8474 = n6785 & ~n8473 ;
  assign n8475 = ~n8470 & n8474 ;
  assign n8476 = n5921 | n8468 ;
  assign n8477 = x189 | n4713 ;
  assign n8478 = x144 & ~n8477 ;
  assign n8479 = ~x174 & n8478 ;
  assign n8480 = x299 | n8479 ;
  assign n8481 = x232 & n8480 ;
  assign n8482 = n8476 & n8481 ;
  assign n8483 = x72 | n8482 ;
  assign n8484 = x39 & n8483 ;
  assign n8485 = n8472 | n8484 ;
  assign n8486 = ( n5880 & n6785 ) | ( n5880 & n8485 ) | ( n6785 & n8485 ) ;
  assign n8487 = ~n6417 & n8471 ;
  assign n8488 = x44 | n1868 ;
  assign n8489 = x101 | n8488 ;
  assign n8490 = n5984 & ~n8489 ;
  assign n8491 = n5927 & n8490 ;
  assign n8492 = x41 & ~n8491 ;
  assign n8493 = ~x41 & x72 ;
  assign n8494 = n1288 & ~n8493 ;
  assign n8495 = x99 | n4793 ;
  assign n8496 = ~x72 & x101 ;
  assign n8497 = x41 | n8496 ;
  assign n8498 = x24 | n1260 ;
  assign n8499 = x252 & ~n4904 ;
  assign n8500 = n5984 & n8499 ;
  assign n8501 = ~n8498 & n8500 ;
  assign n8502 = ~x44 & n8501 ;
  assign n8503 = ~n8497 & n8502 ;
  assign n8504 = n8495 & n8503 ;
  assign n8505 = n8494 & ~n8504 ;
  assign n8506 = ~n8492 & n8505 ;
  assign n8507 = n1288 & n6417 ;
  assign n8508 = ( n6417 & n8471 ) | ( n6417 & n8507 ) | ( n8471 & n8507 ) ;
  assign n8509 = ~n8506 & n8508 ;
  assign n8510 = n8487 | n8509 ;
  assign n8511 = ~x39 & n8510 ;
  assign n8512 = n2007 | n8484 ;
  assign n8513 = n8511 | n8512 ;
  assign n8514 = n2007 & ~n8485 ;
  assign n8515 = x75 & ~n8514 ;
  assign n8516 = n8513 & n8515 ;
  assign n8517 = n5905 & ~n5912 ;
  assign n8518 = x1093 | n5914 ;
  assign n8519 = n8517 | n8518 ;
  assign n8520 = ~x44 & n8519 ;
  assign n8521 = ~n1626 & n5897 ;
  assign n8522 = ~n1624 & n8521 ;
  assign n8523 = n5956 | n8522 ;
  assign n8524 = ~n1269 & n8523 ;
  assign n8525 = n5888 | n8524 ;
  assign n8526 = ~n5885 & n8525 ;
  assign n8527 = x51 | n8526 ;
  assign n8528 = ~n1464 & n8527 ;
  assign n8529 = x96 | n8528 ;
  assign n8530 = n4904 | n5910 ;
  assign n8531 = ~x72 & n5912 ;
  assign n8532 = ~n8530 & n8531 ;
  assign n8533 = n8529 & n8532 ;
  assign n8534 = n8517 | n8533 ;
  assign n8535 = x1093 & ~n8534 ;
  assign n8536 = n8520 & ~n8535 ;
  assign n8537 = ~x101 & n8536 ;
  assign n8538 = x41 & ~n8537 ;
  assign n8539 = x44 & x72 ;
  assign n8540 = x72 | n5905 ;
  assign n8541 = n5912 | n8540 ;
  assign n8542 = ~x1093 & n8541 ;
  assign n8543 = n5908 & n8532 ;
  assign n8544 = ( ~n8531 & n8542 ) | ( ~n8531 & n8543 ) | ( n8542 & n8543 ) ;
  assign n8545 = ~x72 & n8535 ;
  assign n8546 = ( x1093 & n8544 ) | ( x1093 & ~n8545 ) | ( n8544 & ~n8545 ) ;
  assign n8547 = ~x44 & n8546 ;
  assign n8548 = n8539 | n8547 ;
  assign n8549 = x101 | n8548 ;
  assign n8550 = ~n8497 & n8549 ;
  assign n8551 = n1288 & ~n8550 ;
  assign n8552 = ~n8538 & n8551 ;
  assign n8553 = n8540 | n8544 ;
  assign n8554 = ~x44 & n8553 ;
  assign n8555 = n8539 | n8554 ;
  assign n8556 = x101 | n8555 ;
  assign n8557 = ~n8497 & n8556 ;
  assign n8558 = n1288 | n8557 ;
  assign n8559 = x1093 & ~n5905 ;
  assign n8560 = n8520 & ~n8559 ;
  assign n8561 = ~x101 & n8560 ;
  assign n8562 = ( x41 & n8558 ) | ( x41 & ~n8561 ) | ( n8558 & ~n8561 ) ;
  assign n8563 = n8558 | n8562 ;
  assign n8564 = x228 & n8563 ;
  assign n8565 = ~n8552 & n8564 ;
  assign n8566 = x109 | n4877 ;
  assign n8567 = n1344 & ~n8566 ;
  assign n8568 = x110 | n8567 ;
  assign n8569 = n1251 | n1317 ;
  assign n8570 = ~x480 & x949 ;
  assign n8571 = ~n1259 & n8570 ;
  assign n8572 = ~x47 & n8571 ;
  assign n8573 = ~n8569 & n8572 ;
  assign n8574 = n8568 & n8573 ;
  assign n8575 = x901 & ~x959 ;
  assign n8576 = n1344 & ~n1590 ;
  assign n8577 = ~n1259 & n8576 ;
  assign n8578 = ~n8570 & n8577 ;
  assign n8579 = n8575 & ~n8578 ;
  assign n8580 = ~n8574 & n8579 ;
  assign n8581 = n1252 | n1316 ;
  assign n8582 = x110 & ~n8581 ;
  assign n8583 = n8571 & n8582 ;
  assign n8584 = n8575 | n8583 ;
  assign n8585 = ~x250 & x252 ;
  assign n8586 = ~n4904 & n8585 ;
  assign n8587 = n8584 & n8586 ;
  assign n8588 = ~n8580 & n8587 ;
  assign n8589 = ~x72 & n8588 ;
  assign n8590 = ~n8328 & n8582 ;
  assign n8591 = n8570 & ~n8585 ;
  assign n8592 = n8590 & n8591 ;
  assign n8593 = n8589 | n8592 ;
  assign n8594 = ~x44 & n8593 ;
  assign n8595 = ~x101 & n8594 ;
  assign n8596 = x41 & ~n8595 ;
  assign n8597 = n4904 | n8585 ;
  assign n8598 = n8583 & ~n8597 ;
  assign n8599 = x72 | n8598 ;
  assign n8600 = n8588 | n8599 ;
  assign n8601 = ~x44 & n8600 ;
  assign n8602 = n8539 | n8601 ;
  assign n8603 = x101 | n8602 ;
  assign n8604 = ~n8497 & n8603 ;
  assign n8605 = n8596 | n8604 ;
  assign n8606 = ~x228 & n8605 ;
  assign n8607 = x39 | n8606 ;
  assign n8608 = n8565 | n8607 ;
  assign n8609 = x287 & ~n1868 ;
  assign n8610 = n8482 & n8609 ;
  assign n8611 = n8483 & ~n8610 ;
  assign n8612 = x39 & ~n8611 ;
  assign n8613 = n1975 | n8612 ;
  assign n8614 = n8608 & ~n8613 ;
  assign n8615 = n1260 | n4904 ;
  assign n8616 = x44 | n8615 ;
  assign n8617 = n8497 | n8616 ;
  assign n8618 = ~n8493 & n8617 ;
  assign n8619 = x72 | n5984 ;
  assign n8620 = ~n8618 & n8619 ;
  assign n8621 = n8495 & n8620 ;
  assign n8622 = x41 & ~n8490 ;
  assign n8623 = n1288 & n8495 ;
  assign n8624 = n8494 | n8623 ;
  assign n8625 = ~n8622 & n8624 ;
  assign n8626 = ~n8621 & n8625 ;
  assign n8627 = n8508 & ~n8626 ;
  assign n8628 = n8487 | n8627 ;
  assign n8629 = ~x39 & n8628 ;
  assign n8630 = n8484 | n8629 ;
  assign n8631 = n4807 & n8630 ;
  assign n8632 = x38 & n8485 ;
  assign n8633 = x87 | n8632 ;
  assign n8634 = n8631 | n8633 ;
  assign n8635 = n8614 | n8634 ;
  assign n8636 = x41 & n8489 ;
  assign n8637 = x228 & n8618 ;
  assign n8638 = ~n8636 & n8637 ;
  assign n8639 = x228 | n8471 ;
  assign n8640 = ~n1976 & n8639 ;
  assign n8641 = ~n8638 & n8640 ;
  assign n8642 = n1975 & n8472 ;
  assign n8643 = x87 & ~n8642 ;
  assign n8644 = ~n8484 & n8643 ;
  assign n8645 = ~n8641 & n8644 ;
  assign n8646 = x75 | n8645 ;
  assign n8647 = n8635 & ~n8646 ;
  assign n8648 = n8516 | n8647 ;
  assign n8649 = ( ~n5880 & n6785 ) | ( ~n5880 & n8648 ) | ( n6785 & n8648 ) ;
  assign n8650 = n8486 | n8649 ;
  assign n8651 = ~n8475 & n8650 ;
  assign n8652 = x211 & x214 ;
  assign n8653 = x212 & n8652 ;
  assign n8654 = x219 | n8653 ;
  assign n8655 = ~x115 & n1288 ;
  assign n8656 = x42 & ~x114 ;
  assign n8657 = x72 & x116 ;
  assign n8658 = ~x99 & n8550 ;
  assign n8659 = ~x72 & x113 ;
  assign n8660 = x72 & n4786 ;
  assign n8661 = ( x113 & ~n8658 ) | ( x113 & n8660 ) | ( ~n8658 & n8660 ) ;
  assign n8662 = ( n8658 & ~n8659 ) | ( n8658 & n8661 ) | ( ~n8659 & n8661 ) ;
  assign n8663 = ~x116 & n8662 ;
  assign n8664 = n8657 | n8663 ;
  assign n8665 = n8656 & n8664 ;
  assign n8666 = x42 & ~x72 ;
  assign n8667 = x114 & ~n8666 ;
  assign n8668 = ~n4786 & n8537 ;
  assign n8669 = ~n4790 & n8668 ;
  assign n8670 = x42 | n8669 ;
  assign n8671 = ~n8667 & n8670 ;
  assign n8672 = ~n8665 & n8671 ;
  assign n8673 = n8655 & ~n8672 ;
  assign n8674 = x115 | n1288 ;
  assign n8675 = ~n4786 & n8561 ;
  assign n8676 = ~n4790 & n8675 ;
  assign n8677 = ( ~x42 & x114 ) | ( ~x42 & n8676 ) | ( x114 & n8676 ) ;
  assign n8678 = x72 & x113 ;
  assign n8679 = ~x99 & n8557 ;
  assign n8680 = n8660 | n8679 ;
  assign n8681 = ~x113 & n8680 ;
  assign n8682 = n8678 | n8681 ;
  assign n8683 = ~x116 & n8682 ;
  assign n8684 = n8657 | n8683 ;
  assign n8685 = ( x42 & x114 ) | ( x42 & ~n8684 ) | ( x114 & ~n8684 ) ;
  assign n8686 = n8677 | n8685 ;
  assign n8687 = ~n8667 & n8686 ;
  assign n8688 = n8674 | n8687 ;
  assign n8689 = x115 & ~n8666 ;
  assign n8690 = x228 & ~n8689 ;
  assign n8691 = n8688 & n8690 ;
  assign n8692 = ~n8673 & n8691 ;
  assign n8693 = ~x39 & x228 ;
  assign n8694 = ~x99 & n8604 ;
  assign n8695 = n8660 | n8694 ;
  assign n8696 = ~x113 & n8695 ;
  assign n8697 = n8678 | n8696 ;
  assign n8698 = ~x116 & n8697 ;
  assign n8699 = n8657 | n8698 ;
  assign n8700 = n8656 & n8699 ;
  assign n8701 = ~n4786 & n8595 ;
  assign n8702 = ~x113 & n8701 ;
  assign n8703 = ~x116 & n8702 ;
  assign n8704 = x42 | n8703 ;
  assign n8705 = ~n8667 & n8704 ;
  assign n8706 = ~n8700 & n8705 ;
  assign n8707 = x115 | n8706 ;
  assign n8708 = ~n8689 & n8707 ;
  assign n8709 = ( x39 & ~n8693 ) | ( x39 & n8708 ) | ( ~n8693 & n8708 ) ;
  assign n8710 = n8692 | n8709 ;
  assign n8711 = ~x72 & x199 ;
  assign n8712 = x232 | n8711 ;
  assign n8713 = ~x299 & n8712 ;
  assign n8714 = ~x72 & n8477 ;
  assign n8715 = ~n4713 & n8609 ;
  assign n8716 = ~x189 & n8715 ;
  assign n8717 = n8714 | n8716 ;
  assign n8718 = x199 & n8717 ;
  assign n8719 = x232 & ~n8718 ;
  assign n8720 = n8713 & ~n8719 ;
  assign n8721 = x39 & ~n8720 ;
  assign n8722 = n8710 & ~n8721 ;
  assign n8723 = n1975 | n8722 ;
  assign n8724 = n6417 | n8666 ;
  assign n8725 = n8655 & ~n8667 ;
  assign n8726 = n4786 | n8489 ;
  assign n8727 = n4790 | n8726 ;
  assign n8728 = n5984 & ~n8727 ;
  assign n8729 = ~x114 & n4789 ;
  assign n8730 = n8728 & n8729 ;
  assign n8731 = ( ~x42 & x114 ) | ( ~x42 & n8730 ) | ( x114 & n8730 ) ;
  assign n8732 = n4787 | n8616 ;
  assign n8733 = n4790 | n8732 ;
  assign n8734 = ~x72 & n8733 ;
  assign n8735 = n8619 & ~n8734 ;
  assign n8736 = ( x42 & x114 ) | ( x42 & ~n8735 ) | ( x114 & ~n8735 ) ;
  assign n8737 = n8731 | n8736 ;
  assign n8738 = n8725 & n8737 ;
  assign n8739 = n6417 & n8655 ;
  assign n8740 = ( n6417 & ~n8666 ) | ( n6417 & n8739 ) | ( ~n8666 & n8739 ) ;
  assign n8741 = ~n8738 & n8740 ;
  assign n8742 = n8724 & ~n8741 ;
  assign n8743 = x39 | n8742 ;
  assign n8744 = x199 & n8714 ;
  assign n8745 = x232 & ~n8744 ;
  assign n8746 = n8713 & ~n8745 ;
  assign n8747 = x39 & ~n8746 ;
  assign n8748 = n8743 & ~n8747 ;
  assign n8749 = n4807 & ~n8748 ;
  assign n8750 = x39 | n8666 ;
  assign n8751 = ~n8747 & n8750 ;
  assign n8752 = x38 & ~n8751 ;
  assign n8753 = x87 | n8752 ;
  assign n8754 = n8749 | n8753 ;
  assign n8755 = n8723 & ~n8754 ;
  assign n8756 = x228 & ~n8727 ;
  assign n8757 = ~x115 & n8756 ;
  assign n8758 = ~x114 & n8757 ;
  assign n8759 = ~x42 & n8758 ;
  assign n8760 = x228 & ~n8732 ;
  assign n8761 = ~n4792 & n8760 ;
  assign n8762 = n8666 & ~n8761 ;
  assign n8763 = n1976 | n8762 ;
  assign n8764 = n8759 | n8763 ;
  assign n8765 = n1975 & ~n8750 ;
  assign n8766 = x87 & ~n8765 ;
  assign n8767 = n8764 & n8766 ;
  assign n8768 = ~n8747 & n8767 ;
  assign n8769 = x75 | n8768 ;
  assign n8770 = n8755 | n8769 ;
  assign n8771 = n5927 & n8730 ;
  assign n8772 = ~x42 & n8771 ;
  assign n8773 = ~n4787 & n8502 ;
  assign n8774 = ~x113 & n8773 ;
  assign n8775 = ~x116 & n8774 ;
  assign n8776 = n8666 & ~n8775 ;
  assign n8777 = x114 | n8776 ;
  assign n8778 = n8772 | n8777 ;
  assign n8779 = n8725 & n8778 ;
  assign n8780 = n8740 & ~n8779 ;
  assign n8781 = ~n2007 & n8724 ;
  assign n8782 = ~n8780 & n8781 ;
  assign n8783 = n2007 & n8666 ;
  assign n8784 = x39 | n8783 ;
  assign n8785 = n8782 | n8784 ;
  assign n8786 = ~n8747 & n8785 ;
  assign n8787 = x75 & ~n8786 ;
  assign n8788 = n5880 | n8787 ;
  assign n8789 = n8770 & ~n8788 ;
  assign n8790 = x207 & x208 ;
  assign n8791 = n5880 & n8751 ;
  assign n8792 = n8790 | n8791 ;
  assign n8793 = n8789 | n8792 ;
  assign n8794 = ~x72 & x200 ;
  assign n8795 = x232 | n8794 ;
  assign n8796 = ~x299 & n8795 ;
  assign n8797 = x200 & n8714 ;
  assign n8798 = x232 & ~n8797 ;
  assign n8799 = n8796 & ~n8798 ;
  assign n8800 = x39 & ~n8799 ;
  assign n8801 = ~n8746 & n8800 ;
  assign n8802 = n8750 & ~n8801 ;
  assign n8803 = n5880 & n8802 ;
  assign n8804 = n8790 & ~n8803 ;
  assign n8805 = x200 & n8717 ;
  assign n8806 = n8719 & ~n8805 ;
  assign n8807 = n8713 | n8796 ;
  assign n8808 = ~n8806 & n8807 ;
  assign n8809 = x39 & ~n8808 ;
  assign n8810 = n8710 & ~n8809 ;
  assign n8811 = n1975 | n8810 ;
  assign n8812 = x38 & ~n8802 ;
  assign n8813 = x87 | n8812 ;
  assign n8814 = n8743 & ~n8801 ;
  assign n8815 = n4807 & ~n8814 ;
  assign n8816 = n8813 | n8815 ;
  assign n8817 = n8811 & ~n8816 ;
  assign n8818 = n8767 & ~n8801 ;
  assign n8819 = x75 | n8818 ;
  assign n8820 = n8817 | n8819 ;
  assign n8821 = n8785 & ~n8801 ;
  assign n8822 = x75 & ~n8821 ;
  assign n8823 = n5880 | n8822 ;
  assign n8824 = n8820 & ~n8823 ;
  assign n8825 = n8804 & ~n8824 ;
  assign n8826 = n8793 & ~n8825 ;
  assign n8827 = n8654 | n8826 ;
  assign n8828 = x232 & ~x299 ;
  assign n8829 = ~n8718 & n8828 ;
  assign n8830 = ~n8466 & n8609 ;
  assign n8831 = ~x166 & n5924 ;
  assign n8832 = x72 | n8831 ;
  assign n8833 = n7916 & n8832 ;
  assign n8834 = ~n8830 & n8833 ;
  assign n8835 = x72 & ~x232 ;
  assign n8836 = x299 & ~n8835 ;
  assign n8837 = n8712 | n8836 ;
  assign n8838 = ~n8834 & n8837 ;
  assign n8839 = ~n8829 & n8838 ;
  assign n8840 = x39 & ~n8839 ;
  assign n8841 = n8710 & ~n8840 ;
  assign n8842 = n1975 | n8841 ;
  assign n8843 = x299 & ~n8832 ;
  assign n8844 = x39 & ~n8843 ;
  assign n8845 = ~n8746 & n8844 ;
  assign n8846 = n8743 & ~n8845 ;
  assign n8847 = n4807 & ~n8846 ;
  assign n8848 = n8750 & ~n8845 ;
  assign n8849 = x38 & ~n8848 ;
  assign n8850 = x87 | n8849 ;
  assign n8851 = n8847 | n8850 ;
  assign n8852 = n8842 & ~n8851 ;
  assign n8853 = n8767 & ~n8845 ;
  assign n8854 = x75 | n8853 ;
  assign n8855 = n8852 | n8854 ;
  assign n8856 = n8785 & ~n8845 ;
  assign n8857 = x75 & ~n8856 ;
  assign n8858 = n5880 | n8857 ;
  assign n8859 = n8855 & ~n8858 ;
  assign n8860 = n8790 | n8859 ;
  assign n8861 = ~x299 & n8806 ;
  assign n8862 = n8794 | n8837 ;
  assign n8863 = ~n8834 & n8862 ;
  assign n8864 = ~n8861 & n8863 ;
  assign n8865 = x39 & ~n8864 ;
  assign n8866 = n8710 & ~n8865 ;
  assign n8867 = n1975 | n8866 ;
  assign n8868 = n8800 & n8845 ;
  assign n8869 = n8743 & ~n8868 ;
  assign n8870 = n4807 & ~n8869 ;
  assign n8871 = n8813 & n8850 ;
  assign n8872 = n8870 | n8871 ;
  assign n8873 = n8867 & ~n8872 ;
  assign n8874 = n8766 & ~n8868 ;
  assign n8875 = n8764 & n8874 ;
  assign n8876 = x75 | n8875 ;
  assign n8877 = n8873 | n8876 ;
  assign n8878 = n8785 & ~n8868 ;
  assign n8879 = x75 & ~n8878 ;
  assign n8880 = n5880 | n8879 ;
  assign n8881 = n8877 & ~n8880 ;
  assign n8882 = n8804 & ~n8881 ;
  assign n8883 = n8860 & ~n8882 ;
  assign n8884 = n5880 & n8848 ;
  assign n8885 = n8654 & ~n8884 ;
  assign n8886 = ~n8883 & n8885 ;
  assign n8887 = n6785 | n8886 ;
  assign n8888 = n8827 & ~n8887 ;
  assign n8889 = n8654 & ~n8832 ;
  assign n8890 = x39 & ~n8889 ;
  assign n8891 = n6785 & n8750 ;
  assign n8892 = ~n8890 & n8891 ;
  assign n8893 = n8888 | n8892 ;
  assign n8894 = x212 & x214 ;
  assign n8895 = x211 | x219 ;
  assign n8896 = n8894 & n8895 ;
  assign n8897 = x211 | n8894 ;
  assign n8898 = ~n8896 & n8897 ;
  assign n8899 = ~n8832 & n8898 ;
  assign n8900 = x39 & ~n8899 ;
  assign n8901 = x43 & ~x72 ;
  assign n8902 = x39 | n8901 ;
  assign n8903 = n6785 & n8902 ;
  assign n8904 = ~n8900 & n8903 ;
  assign n8905 = ~x228 & n8699 ;
  assign n8906 = ( x228 & ~n1288 ) | ( x228 & n8664 ) | ( ~n1288 & n8664 ) ;
  assign n8907 = ( x228 & n1288 ) | ( x228 & n8684 ) | ( n1288 & n8684 ) ;
  assign n8908 = n8906 & n8907 ;
  assign n8909 = n8905 | n8908 ;
  assign n8910 = x42 | n4791 ;
  assign n8911 = x43 & ~n8910 ;
  assign n8912 = n8909 & n8911 ;
  assign n8913 = x228 | n8703 ;
  assign n8914 = n1288 | n8675 ;
  assign n8915 = n1288 & ~n8668 ;
  assign n8916 = n8914 & ~n8915 ;
  assign n8917 = ~n4790 & n8916 ;
  assign n8918 = x228 & ~n8917 ;
  assign n8919 = n8913 & ~n8918 ;
  assign n8920 = x43 | n8919 ;
  assign n8921 = ~n8901 & n8910 ;
  assign n8922 = n8920 & ~n8921 ;
  assign n8923 = ~n8912 & n8922 ;
  assign n8924 = x39 | n8923 ;
  assign n8925 = x232 & ~n8805 ;
  assign n8926 = n8796 & ~n8925 ;
  assign n8927 = x39 & ~n8926 ;
  assign n8928 = n8924 & ~n8927 ;
  assign n8929 = n1975 | n8928 ;
  assign n8930 = n6417 | n8901 ;
  assign n8931 = n1288 & ~n8910 ;
  assign n8932 = n8901 & ~n8931 ;
  assign n8933 = n6417 & ~n8932 ;
  assign n8934 = ~x43 & x52 ;
  assign n8935 = n8728 & n8934 ;
  assign n8936 = x43 & ~n8735 ;
  assign n8937 = n8935 | n8936 ;
  assign n8938 = n8931 & n8937 ;
  assign n8939 = n8933 & ~n8938 ;
  assign n8940 = n8930 & ~n8939 ;
  assign n8941 = x39 | n8940 ;
  assign n8942 = ~n8800 & n8941 ;
  assign n8943 = n4807 & ~n8942 ;
  assign n8944 = ~n8800 & n8902 ;
  assign n8945 = x38 & ~n8944 ;
  assign n8946 = x87 | n8945 ;
  assign n8947 = n8943 | n8946 ;
  assign n8948 = n8929 & ~n8947 ;
  assign n8949 = x228 & ~n8910 ;
  assign n8950 = n8901 & ~n8949 ;
  assign n8951 = n1976 | n8950 ;
  assign n8952 = ( ~x43 & n8734 ) | ( ~x43 & n8949 ) | ( n8734 & n8949 ) ;
  assign n8953 = ( x43 & ~n8727 ) | ( x43 & n8949 ) | ( ~n8727 & n8949 ) ;
  assign n8954 = n8952 & n8953 ;
  assign n8955 = n8951 | n8954 ;
  assign n8956 = n1975 & ~n8902 ;
  assign n8957 = x87 & ~n8956 ;
  assign n8958 = n8955 & n8957 ;
  assign n8959 = ~n8800 & n8958 ;
  assign n8960 = x75 | n8959 ;
  assign n8961 = n8948 | n8960 ;
  assign n8962 = x72 | n8775 ;
  assign n8963 = x43 & ~n8962 ;
  assign n8964 = n5927 & n8728 ;
  assign n8965 = n8934 & n8964 ;
  assign n8966 = n8963 | n8965 ;
  assign n8967 = n8931 & n8966 ;
  assign n8968 = n8933 & ~n8967 ;
  assign n8969 = n8930 & ~n8968 ;
  assign n8970 = ( x39 & ~n2007 ) | ( x39 & n8969 ) | ( ~n2007 & n8969 ) ;
  assign n8971 = ( x39 & n2007 ) | ( x39 & n8901 ) | ( n2007 & n8901 ) ;
  assign n8972 = n8970 | n8971 ;
  assign n8973 = ~n8800 & n8972 ;
  assign n8974 = x75 & ~n8973 ;
  assign n8975 = n5880 | n8974 ;
  assign n8976 = n8961 & ~n8975 ;
  assign n8977 = n5880 & n8944 ;
  assign n8978 = n8790 | n8977 ;
  assign n8979 = n8976 | n8978 ;
  assign n8980 = x199 | x200 ;
  assign n8981 = ~x299 & n8980 ;
  assign n8982 = x72 | n8981 ;
  assign n8983 = ~x232 & n8982 ;
  assign n8984 = x299 | n8983 ;
  assign n8985 = n8717 & ~n8980 ;
  assign n8986 = x232 & ~n8985 ;
  assign n8987 = n8984 | n8986 ;
  assign n8988 = x39 & n8987 ;
  assign n8989 = n8924 & ~n8988 ;
  assign n8990 = n1975 | n8989 ;
  assign n8991 = n8714 & ~n8980 ;
  assign n8992 = x232 & ~n8991 ;
  assign n8993 = n8984 | n8992 ;
  assign n8994 = x39 & n8993 ;
  assign n8995 = n8941 & ~n8994 ;
  assign n8996 = n4807 & ~n8995 ;
  assign n8997 = n8902 & ~n8994 ;
  assign n8998 = x38 & ~n8997 ;
  assign n8999 = x87 | n8998 ;
  assign n9000 = n8996 | n8999 ;
  assign n9001 = n8990 & ~n9000 ;
  assign n9002 = n2041 & ~n8997 ;
  assign n9003 = n8958 & ~n9002 ;
  assign n9004 = x75 | n9003 ;
  assign n9005 = n9001 | n9004 ;
  assign n9006 = n8972 & ~n8994 ;
  assign n9007 = x75 & ~n9006 ;
  assign n9008 = n5880 | n9007 ;
  assign n9009 = n9005 & ~n9008 ;
  assign n9010 = n5880 & n8997 ;
  assign n9011 = n8790 & ~n9010 ;
  assign n9012 = ~n9009 & n9011 ;
  assign n9013 = n8979 & ~n9012 ;
  assign n9014 = ( ~n6785 & n8898 ) | ( ~n6785 & n9013 ) | ( n8898 & n9013 ) ;
  assign n9015 = ~n8805 & n8828 ;
  assign n9016 = ~n8834 & n8836 ;
  assign n9017 = ( n8795 & ~n8834 ) | ( n8795 & n9016 ) | ( ~n8834 & n9016 ) ;
  assign n9018 = ~n9015 & n9017 ;
  assign n9019 = x39 & ~n9018 ;
  assign n9020 = n8924 & ~n9019 ;
  assign n9021 = n1975 | n9020 ;
  assign n9022 = ~n8799 & n8844 ;
  assign n9023 = n8941 & ~n9022 ;
  assign n9024 = n4807 & ~n9023 ;
  assign n9025 = n8902 & ~n9022 ;
  assign n9026 = x38 & ~n9025 ;
  assign n9027 = x87 | n9026 ;
  assign n9028 = n9024 | n9027 ;
  assign n9029 = n9021 & ~n9028 ;
  assign n9030 = n8958 & ~n9022 ;
  assign n9031 = x75 | n9030 ;
  assign n9032 = n9029 | n9031 ;
  assign n9033 = n8972 & ~n9022 ;
  assign n9034 = x75 & ~n9033 ;
  assign n9035 = n5880 | n9034 ;
  assign n9036 = n9032 & ~n9035 ;
  assign n9037 = n5880 & n9025 ;
  assign n9038 = n8790 | n9037 ;
  assign n9039 = n9036 | n9038 ;
  assign n9040 = n8828 & ~n8985 ;
  assign n9041 = n8834 | n8983 ;
  assign n9042 = n9040 | n9041 ;
  assign n9043 = x39 & n9042 ;
  assign n9044 = n8924 & ~n9043 ;
  assign n9045 = n1975 | n9044 ;
  assign n9046 = ~n8843 & n8994 ;
  assign n9047 = n8941 & ~n9046 ;
  assign n9048 = n4807 & ~n9047 ;
  assign n9049 = n8902 & ~n9046 ;
  assign n9050 = x38 & ~n9049 ;
  assign n9051 = x87 | n9050 ;
  assign n9052 = n9048 | n9051 ;
  assign n9053 = n9045 & ~n9052 ;
  assign n9054 = n8958 & ~n9046 ;
  assign n9055 = x75 | n9054 ;
  assign n9056 = n9053 | n9055 ;
  assign n9057 = n8972 & ~n9046 ;
  assign n9058 = x75 & ~n9057 ;
  assign n9059 = n5880 | n9058 ;
  assign n9060 = n9056 & ~n9059 ;
  assign n9061 = n5880 & n9049 ;
  assign n9062 = n8790 & ~n9061 ;
  assign n9063 = ~n9060 & n9062 ;
  assign n9064 = n9039 & ~n9063 ;
  assign n9065 = ( n6785 & n8898 ) | ( n6785 & ~n9064 ) | ( n8898 & ~n9064 ) ;
  assign n9066 = n9014 & ~n9065 ;
  assign n9067 = n8904 | n9066 ;
  assign n9068 = ~n1524 & n5924 ;
  assign n9069 = ~x72 & n9068 ;
  assign n9070 = x39 & ~n9069 ;
  assign n9071 = x44 & ~x72 ;
  assign n9072 = x39 | n9071 ;
  assign n9073 = n6785 & n9072 ;
  assign n9074 = ~n9070 & n9073 ;
  assign n9075 = ~x72 & n5925 ;
  assign n9076 = x39 & ~n9075 ;
  assign n9077 = n9072 & ~n9076 ;
  assign n9078 = ( n5880 & n6785 ) | ( n5880 & ~n9077 ) | ( n6785 & ~n9077 ) ;
  assign n9079 = x44 & ~n8546 ;
  assign n9080 = n1288 & ~n8536 ;
  assign n9081 = ~n9079 & n9080 ;
  assign n9082 = x44 & ~n8553 ;
  assign n9083 = n1288 | n8560 ;
  assign n9084 = n9082 | n9083 ;
  assign n9085 = ~n9081 & n9084 ;
  assign n9086 = x228 & ~n9085 ;
  assign n9087 = x44 & ~n8600 ;
  assign n9088 = n8594 | n9087 ;
  assign n9089 = ( ~x39 & n8693 ) | ( ~x39 & n9088 ) | ( n8693 & n9088 ) ;
  assign n9090 = ~n9086 & n9089 ;
  assign n9091 = x39 & n5925 ;
  assign n9092 = x287 & ~n8615 ;
  assign n9093 = x72 | n9092 ;
  assign n9094 = n9091 & ~n9093 ;
  assign n9095 = n1975 | n9094 ;
  assign n9096 = n9090 | n9095 ;
  assign n9097 = n6417 | n9071 ;
  assign n9098 = ~x39 & n9097 ;
  assign n9099 = n5929 & ~n8539 ;
  assign n9100 = n5984 & ~n8488 ;
  assign n9101 = n5984 & ~n8615 ;
  assign n9102 = x44 & ~n9101 ;
  assign n9103 = n9100 | n9102 ;
  assign n9104 = n9099 & n9103 ;
  assign n9105 = ( n6417 & n8507 ) | ( n6417 & ~n9071 ) | ( n8507 & ~n9071 ) ;
  assign n9106 = ~n9104 & n9105 ;
  assign n9107 = n9098 & ~n9106 ;
  assign n9108 = ~x72 & n9091 ;
  assign n9109 = n4807 & ~n9108 ;
  assign n9110 = ~n9107 & n9109 ;
  assign n9111 = x38 & ~n9077 ;
  assign n9112 = x87 | n9111 ;
  assign n9113 = n9110 | n9112 ;
  assign n9114 = n9096 & ~n9113 ;
  assign n9115 = x228 & ~n1975 ;
  assign n9116 = ~n8488 & n9115 ;
  assign n9117 = ~n8615 & n9115 ;
  assign n9118 = n9071 & ~n9117 ;
  assign n9119 = x39 | n9118 ;
  assign n9120 = n9116 | n9119 ;
  assign n9121 = ~n9076 & n9120 ;
  assign n9122 = ( x75 & n1998 ) | ( x75 & n9121 ) | ( n1998 & n9121 ) ;
  assign n9123 = n9114 | n9122 ;
  assign n9124 = ( ~x75 & n2007 ) | ( ~x75 & n9077 ) | ( n2007 & n9077 ) ;
  assign n9125 = n5927 & n9100 ;
  assign n9126 = x44 & ~n8501 ;
  assign n9127 = n9125 | n9126 ;
  assign n9128 = n9099 & n9127 ;
  assign n9129 = n9105 & ~n9128 ;
  assign n9130 = n9098 & ~n9129 ;
  assign n9131 = n9108 | n9130 ;
  assign n9132 = ( x75 & n2007 ) | ( x75 & ~n9131 ) | ( n2007 & ~n9131 ) ;
  assign n9133 = ~n9124 & n9132 ;
  assign n9134 = n9123 & ~n9133 ;
  assign n9135 = ( n5880 & ~n6785 ) | ( n5880 & n9134 ) | ( ~n6785 & n9134 ) ;
  assign n9136 = ~n9078 & n9135 ;
  assign n9137 = n9074 | n9136 ;
  assign n9138 = ~x38 & x39 ;
  assign n9139 = ~n8359 & n9138 ;
  assign n9140 = x979 & n9139 ;
  assign n9141 = ~n4981 & n9140 ;
  assign n9142 = x49 | x76 ;
  assign n9143 = n7142 | n9142 ;
  assign n9144 = x102 | x104 ;
  assign n9145 = x111 | n9144 ;
  assign n9146 = n8339 | n9145 ;
  assign n9147 = n9143 | n9146 ;
  assign n9148 = x61 & ~x82 ;
  assign n9149 = x83 | x89 ;
  assign n9150 = n9148 & ~n9149 ;
  assign n9151 = n1244 | n7156 ;
  assign n9152 = n9150 & ~n9151 ;
  assign n9153 = ~n7154 & n9152 ;
  assign n9154 = ~n8410 & n9153 ;
  assign n9155 = ~n9147 & n9154 ;
  assign n9156 = ~n7170 & n9155 ;
  assign n9157 = ~x841 & n9156 ;
  assign n9158 = ~n1253 & n1730 ;
  assign n9159 = x24 & n9158 ;
  assign n9160 = n9157 | n9159 ;
  assign n9161 = ~n8332 & n9160 ;
  assign n9162 = x82 | n1366 ;
  assign n9163 = ~x84 & x104 ;
  assign n9164 = ~n1363 & n9163 ;
  assign n9165 = ~n8343 & n9164 ;
  assign n9166 = ~n9162 & n9165 ;
  assign n9167 = x36 | n9166 ;
  assign n9168 = n7155 | n7266 ;
  assign n9169 = x67 | x103 ;
  assign n9170 = n1236 | n9169 ;
  assign n9171 = x98 | n9170 ;
  assign n9172 = n9168 | n9171 ;
  assign n9173 = n9167 & ~n9172 ;
  assign n9174 = ~n1400 & n9173 ;
  assign n9175 = x88 | n9174 ;
  assign n9176 = ~n1312 & n9175 ;
  assign n9177 = n1244 | n1437 ;
  assign n9178 = n1244 | n1436 ;
  assign n9179 = ( n1241 & n9177 ) | ( n1241 & n9178 ) | ( n9177 & n9178 ) ;
  assign n9180 = n9176 & ~n9179 ;
  assign n9181 = ~n1251 & n9180 ;
  assign n9182 = n8325 | n9181 ;
  assign n9183 = ~n8328 & n9182 ;
  assign n9184 = n5997 & ~n9183 ;
  assign n9185 = ~n1692 & n9183 ;
  assign n9186 = ~x36 & n9173 ;
  assign n9187 = x88 | n9186 ;
  assign n9188 = ~n9179 & n9187 ;
  assign n9189 = ~n8338 & n9188 ;
  assign n9190 = ~x824 & n1692 ;
  assign n9191 = n9189 & n9190 ;
  assign n9192 = x829 & ~n9191 ;
  assign n9193 = ~n9185 & n9192 ;
  assign n9194 = ~n1287 & n9193 ;
  assign n9195 = n9184 | n9194 ;
  assign n9196 = x1091 & n9195 ;
  assign n9197 = ~n5950 & n9183 ;
  assign n9198 = x829 | n9197 ;
  assign n9199 = ~n9193 & n9198 ;
  assign n9200 = x1093 | n9199 ;
  assign n9201 = n5950 & ~n8328 ;
  assign n9202 = n8326 & n9201 ;
  assign n9203 = n4986 & ~n5995 ;
  assign n9204 = n9202 | n9203 ;
  assign n9205 = n9197 | n9204 ;
  assign n9206 = ~n8331 & n9205 ;
  assign n9207 = n9200 & n9206 ;
  assign n9208 = ~n9196 & n9207 ;
  assign n9209 = ~x72 & x841 ;
  assign n9210 = ~n1256 & n9209 ;
  assign n9211 = ~x51 & n9210 ;
  assign n9212 = n8417 & n9211 ;
  assign n9213 = ~n8331 & n9212 ;
  assign n9214 = ~n8337 & n9213 ;
  assign n9215 = x103 | n1393 ;
  assign n9216 = n8408 | n9215 ;
  assign n9217 = n7142 | n7155 ;
  assign n9218 = n9216 | n9217 ;
  assign n9219 = n1236 | n1245 ;
  assign n9220 = ~x45 & x49 ;
  assign n9221 = ~n9145 & n9220 ;
  assign n9222 = ~n9219 & n9221 ;
  assign n9223 = ~n9218 & n9222 ;
  assign n9224 = ~n9162 & n9223 ;
  assign n9225 = n1257 | n7170 ;
  assign n9226 = n9224 & ~n9225 ;
  assign n9227 = ~n8327 & n9210 ;
  assign n9228 = n9226 & n9227 ;
  assign n9229 = n5844 | n6785 ;
  assign n9230 = ( x74 & n9228 ) | ( x74 & ~n9229 ) | ( n9228 & ~n9229 ) ;
  assign n9231 = ( x74 & n7192 ) | ( x74 & n9229 ) | ( n7192 & n9229 ) ;
  assign n9232 = n9230 & ~n9231 ;
  assign n9233 = x24 & ~n7130 ;
  assign n9234 = n8576 | n9233 ;
  assign n9235 = x24 & ~x94 ;
  assign n9236 = ~n7128 & n9235 ;
  assign n9237 = x252 | n7119 ;
  assign n9238 = x252 & ~n7136 ;
  assign n9239 = n9237 & ~n9238 ;
  assign n9240 = ~n8328 & n9239 ;
  assign n9241 = ~n9236 & n9240 ;
  assign n9242 = n9234 & n9241 ;
  assign n9243 = n1526 | n5904 ;
  assign n9244 = x24 & ~x90 ;
  assign n9245 = ~n9243 & n9244 ;
  assign n9246 = ~n9239 & n9245 ;
  assign n9247 = n7132 & n9246 ;
  assign n9248 = n9242 | n9247 ;
  assign n9249 = ~x100 & n9248 ;
  assign n9250 = x100 & n4784 ;
  assign n9251 = n5028 & n9250 ;
  assign n9252 = n9249 | n9251 ;
  assign n9253 = n1925 | n1998 ;
  assign n9254 = n9252 & ~n9253 ;
  assign n9255 = n4804 & n7197 ;
  assign n9256 = ~n7193 & n9255 ;
  assign n9257 = n9254 | n9256 ;
  assign n9258 = ~n7113 & n9257 ;
  assign n9259 = n1251 | n8332 ;
  assign n9260 = n1312 | n9259 ;
  assign n9261 = n7267 | n9219 ;
  assign n9262 = n1233 | n9261 ;
  assign n9263 = x69 | n9262 ;
  assign n9264 = n1393 | n9263 ;
  assign n9265 = n1395 & ~n9264 ;
  assign n9266 = ~n9260 & n9265 ;
  assign n9267 = x219 | n8897 ;
  assign n9268 = x52 & ~x72 ;
  assign n9269 = ~x39 & n9268 ;
  assign n9270 = n5880 & ~n9269 ;
  assign n9271 = n8790 & ~n9270 ;
  assign n9272 = x114 | n4788 ;
  assign n9273 = n8739 & ~n9272 ;
  assign n9274 = n8775 & n9273 ;
  assign n9275 = ~n2007 & n9274 ;
  assign n9276 = n9269 & ~n9275 ;
  assign n9277 = ( x75 & n5880 ) | ( x75 & n9276 ) | ( n5880 & n9276 ) ;
  assign n9278 = n5984 & n9273 ;
  assign n9279 = ~n8733 & n9278 ;
  assign n9280 = n9268 & ~n9279 ;
  assign n9281 = ( x39 & x100 ) | ( x39 & ~n9280 ) | ( x100 & ~n9280 ) ;
  assign n9282 = ( x52 & n8655 ) | ( x52 & ~n8669 ) | ( n8655 & ~n8669 ) ;
  assign n9283 = ( ~x52 & n8655 ) | ( ~x52 & n8664 ) | ( n8655 & n8664 ) ;
  assign n9284 = n9282 & n9283 ;
  assign n9285 = ( ~x52 & n8674 ) | ( ~x52 & n8676 ) | ( n8674 & n8676 ) ;
  assign n9286 = ( x52 & n8674 ) | ( x52 & ~n8684 ) | ( n8674 & ~n8684 ) ;
  assign n9287 = n9285 | n9286 ;
  assign n9288 = ~n9284 & n9287 ;
  assign n9289 = n9272 | n9288 ;
  assign n9290 = n4788 | n4791 ;
  assign n9291 = ~n9268 & n9290 ;
  assign n9292 = x228 & ~n9291 ;
  assign n9293 = n9289 & n9292 ;
  assign n9294 = ( ~x52 & n8703 ) | ( ~x52 & n9290 ) | ( n8703 & n9290 ) ;
  assign n9295 = ( x52 & ~n8699 ) | ( x52 & n9290 ) | ( ~n8699 & n9290 ) ;
  assign n9296 = n9294 | n9295 ;
  assign n9297 = ~n9291 & n9296 ;
  assign n9298 = ( x39 & ~n8693 ) | ( x39 & n9297 ) | ( ~n8693 & n9297 ) ;
  assign n9299 = n9293 | n9298 ;
  assign n9300 = ( ~x39 & x100 ) | ( ~x39 & n9299 ) | ( x100 & n9299 ) ;
  assign n9301 = ~n9281 & n9300 ;
  assign n9302 = x38 | n9301 ;
  assign n9303 = x38 & ~n9269 ;
  assign n9304 = x87 | n9303 ;
  assign n9305 = n9302 & ~n9304 ;
  assign n9306 = ~x100 & n9138 ;
  assign n9307 = x87 & ~n9306 ;
  assign n9308 = ( ~x100 & n9269 ) | ( ~x100 & n9307 ) | ( n9269 & n9307 ) ;
  assign n9309 = x228 & ~n9290 ;
  assign n9310 = n9268 & ~n9309 ;
  assign n9311 = ( ~x52 & n8734 ) | ( ~x52 & n9309 ) | ( n8734 & n9309 ) ;
  assign n9312 = ( x52 & ~n8727 ) | ( x52 & n9309 ) | ( ~n8727 & n9309 ) ;
  assign n9313 = n9311 & n9312 ;
  assign n9314 = n9310 | n9313 ;
  assign n9315 = x38 | n9314 ;
  assign n9316 = ~n9303 & n9315 ;
  assign n9317 = ( x100 & n9307 ) | ( x100 & n9316 ) | ( n9307 & n9316 ) ;
  assign n9318 = n9308 & n9317 ;
  assign n9319 = n9305 | n9318 ;
  assign n9320 = ( ~x75 & n5880 ) | ( ~x75 & n9319 ) | ( n5880 & n9319 ) ;
  assign n9321 = n9277 | n9320 ;
  assign n9322 = n9271 & n9321 ;
  assign n9323 = ~n8988 & n9299 ;
  assign n9324 = n1975 | n9323 ;
  assign n9325 = x39 | n9280 ;
  assign n9326 = ~n8994 & n9325 ;
  assign n9327 = n4807 & ~n9326 ;
  assign n9328 = x39 | n9268 ;
  assign n9329 = ~n8994 & n9328 ;
  assign n9330 = x38 & ~n9329 ;
  assign n9331 = x87 | n9330 ;
  assign n9332 = n9327 | n9331 ;
  assign n9333 = n9324 & ~n9332 ;
  assign n9334 = n1975 & n9329 ;
  assign n9335 = x39 | n9314 ;
  assign n9336 = n1975 | n8994 ;
  assign n9337 = n9335 & ~n9336 ;
  assign n9338 = n9334 | n9337 ;
  assign n9339 = x87 & n9338 ;
  assign n9340 = x75 | n9339 ;
  assign n9341 = n9333 | n9340 ;
  assign n9342 = n2007 & n9329 ;
  assign n9343 = x75 & ~n9342 ;
  assign n9344 = n2007 | n8994 ;
  assign n9345 = n9269 & ~n9274 ;
  assign n9346 = ( x39 & ~n9344 ) | ( x39 & n9345 ) | ( ~n9344 & n9345 ) ;
  assign n9347 = n9343 & ~n9346 ;
  assign n9348 = n5880 | n8790 ;
  assign n9349 = n9347 | n9348 ;
  assign n9350 = n9341 & ~n9349 ;
  assign n9351 = n9322 | n9350 ;
  assign n9352 = n9267 & n9351 ;
  assign n9353 = x39 & ~n9016 ;
  assign n9354 = n9299 & ~n9353 ;
  assign n9355 = n1975 | n9354 ;
  assign n9356 = ~n8844 & n9328 ;
  assign n9357 = x38 & ~n9356 ;
  assign n9358 = ~n8844 & n9325 ;
  assign n9359 = n4807 & ~n9358 ;
  assign n9360 = n9357 | n9359 ;
  assign n9361 = n9355 & ~n9360 ;
  assign n9362 = x87 | n9361 ;
  assign n9363 = n1975 & n9356 ;
  assign n9364 = x87 & ~n9363 ;
  assign n9365 = n1975 | n8844 ;
  assign n9366 = n9335 & ~n9365 ;
  assign n9367 = n9364 & ~n9366 ;
  assign n9368 = n8790 & ~n9367 ;
  assign n9369 = n9362 & n9368 ;
  assign n9370 = ~n9043 & n9299 ;
  assign n9371 = n1975 | n9370 ;
  assign n9372 = ~n9046 & n9325 ;
  assign n9373 = n4807 & ~n9372 ;
  assign n9374 = n9330 & ~n9356 ;
  assign n9375 = n9373 | n9374 ;
  assign n9376 = n9371 & ~n9375 ;
  assign n9377 = x87 | n9376 ;
  assign n9378 = n1975 | n9046 ;
  assign n9379 = n9335 & ~n9378 ;
  assign n9380 = ~n9334 & n9364 ;
  assign n9381 = ~n9379 & n9380 ;
  assign n9382 = n8790 | n9381 ;
  assign n9383 = n9377 & ~n9382 ;
  assign n9384 = n9369 | n9383 ;
  assign n9385 = ~x75 & n9384 ;
  assign n9386 = ( ~x75 & n8790 ) | ( ~x75 & n8844 ) | ( n8790 & n8844 ) ;
  assign n9387 = ( x75 & n8790 ) | ( x75 & ~n9046 ) | ( n8790 & ~n9046 ) ;
  assign n9388 = ~n9386 & n9387 ;
  assign n9389 = ( x39 & n9276 ) | ( x39 & n9388 ) | ( n9276 & n9388 ) ;
  assign n9390 = n5880 | n9389 ;
  assign n9391 = n9385 | n9390 ;
  assign n9392 = n5880 & ~n9356 ;
  assign n9393 = n9267 | n9392 ;
  assign n9394 = n9391 & ~n9393 ;
  assign n9395 = n5880 & ~n8790 ;
  assign n9396 = n9329 & n9395 ;
  assign n9397 = n6785 | n9396 ;
  assign n9398 = n9394 | n9397 ;
  assign n9399 = n9352 | n9398 ;
  assign n9400 = x39 & ~n9267 ;
  assign n9401 = ~n8832 & n9400 ;
  assign n9402 = n6785 & ~n9269 ;
  assign n9403 = ~n9401 & n9402 ;
  assign n9404 = n9399 & ~n9403 ;
  assign n9405 = x287 | x979 ;
  assign n9406 = n4727 & ~n9405 ;
  assign n9407 = x39 & ~n9406 ;
  assign n9408 = n8366 | n9407 ;
  assign n9409 = x53 & ~n1326 ;
  assign n9410 = ~n1590 & n9409 ;
  assign n9411 = ~n1583 & n9410 ;
  assign n9412 = x24 & ~n8328 ;
  assign n9413 = ~x39 & n9412 ;
  assign n9414 = n9411 & n9413 ;
  assign n9415 = ( x39 & ~n9408 ) | ( x39 & n9414 ) | ( ~n9408 & n9414 ) ;
  assign n9416 = ~n2120 & n9415 ;
  assign n9417 = n7130 | n7272 ;
  assign n9418 = x60 | x85 ;
  assign n9419 = x106 & ~n9418 ;
  assign n9420 = n1227 | n7146 ;
  assign n9421 = n9419 & ~n9420 ;
  assign n9422 = ~n9143 & n9421 ;
  assign n9423 = n7159 | n9216 ;
  assign n9424 = n9422 & ~n9423 ;
  assign n9425 = ~n9219 & n9424 ;
  assign n9426 = ~n9417 & n9425 ;
  assign n9427 = x841 | n1255 ;
  assign n9428 = n7190 | n9427 ;
  assign n9429 = n1257 | n2005 ;
  assign n9430 = n9428 | n9429 ;
  assign n9431 = n9426 & ~n9430 ;
  assign n9432 = ( x54 & ~n7112 ) | ( x54 & n9431 ) | ( ~n7112 & n9431 ) ;
  assign n9433 = ~n2008 & n8363 ;
  assign n9434 = ( x54 & n7112 ) | ( x54 & ~n9433 ) | ( n7112 & ~n9433 ) ;
  assign n9435 = n9432 & ~n9434 ;
  assign n9436 = x104 | n1224 ;
  assign n9437 = x45 & ~n1227 ;
  assign n9438 = ~n1236 & n9437 ;
  assign n9439 = ~n9218 & n9438 ;
  assign n9440 = ~n9436 & n9439 ;
  assign n9441 = n4904 | n7514 ;
  assign n9442 = n2033 | n8353 ;
  assign n9443 = n9441 | n9442 ;
  assign n9444 = n9440 & ~n9443 ;
  assign n9445 = ( x55 & ~n7111 ) | ( x55 & n9444 ) | ( ~n7111 & n9444 ) ;
  assign n9446 = ~x54 & n9433 ;
  assign n9447 = ~x74 & n9446 ;
  assign n9448 = ( x55 & n7111 ) | ( x55 & ~n9447 ) | ( n7111 & ~n9447 ) ;
  assign n9449 = n9445 & ~n9448 ;
  assign n9450 = x56 & ~x62 ;
  assign n9451 = x55 & ~n8309 ;
  assign n9452 = n9450 | n9451 ;
  assign n9453 = n1863 | n2045 ;
  assign n9454 = n4697 & ~n9453 ;
  assign n9455 = x56 & ~n9454 ;
  assign n9456 = n2057 | n9455 ;
  assign n9457 = n9452 & ~n9456 ;
  assign n9458 = ~n5086 & n9447 ;
  assign n9459 = ( x57 & x59 ) | ( x57 & ~n9458 ) | ( x59 & ~n9458 ) ;
  assign n9460 = n4911 | n9453 ;
  assign n9461 = ~x56 & x62 ;
  assign n9462 = ~x924 & n9461 ;
  assign n9463 = n9450 | n9462 ;
  assign n9464 = ~n9460 & n9463 ;
  assign n9465 = ( x57 & ~x59 ) | ( x57 & n9464 ) | ( ~x59 & n9464 ) ;
  assign n9466 = ~n9459 & n9465 ;
  assign n9467 = x93 | n9243 ;
  assign n9468 = n8331 | n9467 ;
  assign n9469 = n5887 & ~n9468 ;
  assign n9470 = x924 & n9461 ;
  assign n9471 = ~n9460 & n9470 ;
  assign n9472 = ( ~x57 & x59 ) | ( ~x57 & n9471 ) | ( x59 & n9471 ) ;
  assign n9473 = ~n9459 & n9472 ;
  assign n9474 = x39 & ~x979 ;
  assign n9475 = ~n4727 & n9474 ;
  assign n9476 = ~n4725 & n9475 ;
  assign n9477 = ~n4981 & n9476 ;
  assign n9478 = n9413 & ~n9417 ;
  assign n9479 = n1581 & n9478 ;
  assign n9480 = n9477 | n9479 ;
  assign n9481 = ~n8366 & n9480 ;
  assign n9482 = x841 & n9156 ;
  assign n9483 = x24 | n9417 ;
  assign n9484 = n1581 & ~n9483 ;
  assign n9485 = n9482 | n9484 ;
  assign n9486 = ~n8332 & n9485 ;
  assign n9487 = n9454 & n9461 ;
  assign n9488 = ( x57 & ~x59 ) | ( x57 & n9487 ) | ( ~x59 & n9487 ) ;
  assign n9489 = ~n8311 & n9488 ;
  assign n9490 = n1423 & ~n7170 ;
  assign n9491 = ~n7269 & n9490 ;
  assign n9492 = x999 & n9491 ;
  assign n9493 = ~x24 & n9158 ;
  assign n9494 = n9492 | n9493 ;
  assign n9495 = ~n8332 & n9494 ;
  assign n9496 = ~x63 & x107 ;
  assign n9497 = ~n7269 & n9496 ;
  assign n9498 = ( x841 & ~n9260 ) | ( x841 & n9497 ) | ( ~n9260 & n9497 ) ;
  assign n9499 = ~n1415 & n9496 ;
  assign n9500 = x64 | n9499 ;
  assign n9501 = ~n8353 & n9500 ;
  assign n9502 = ~n8335 & n9501 ;
  assign n9503 = ( x841 & n9260 ) | ( x841 & ~n9502 ) | ( n9260 & ~n9502 ) ;
  assign n9504 = n9498 & ~n9503 ;
  assign n9505 = x39 & n8382 ;
  assign n9506 = ~n8366 & n9505 ;
  assign n9507 = n8386 & n9506 ;
  assign n9508 = ~n8380 & n9507 ;
  assign n9509 = x314 & ~n1245 ;
  assign n9510 = ~n9441 & n9509 ;
  assign n9511 = x81 & ~x102 ;
  assign n9512 = n9510 & n9511 ;
  assign n9513 = ~n1242 & n9512 ;
  assign n9514 = n1975 | n2031 ;
  assign n9515 = x199 & ~x299 ;
  assign n9516 = ~n1983 & n9515 ;
  assign n9517 = ~n9514 & n9516 ;
  assign n9518 = n9513 & n9517 ;
  assign n9519 = ( x219 & ~n6785 ) | ( x219 & n9518 ) | ( ~n6785 & n9518 ) ;
  assign n9520 = x199 | x299 ;
  assign n9521 = ~n2033 & n9513 ;
  assign n9522 = n9520 & n9521 ;
  assign n9523 = ( x219 & n6785 ) | ( x219 & ~n9522 ) | ( n6785 & ~n9522 ) ;
  assign n9524 = n9519 & ~n9523 ;
  assign n9525 = x83 & ~x103 ;
  assign n9526 = ~n9261 & n9525 ;
  assign n9527 = ~n8331 & n9526 ;
  assign n9528 = n9510 & n9527 ;
  assign n9529 = ~n1358 & n9528 ;
  assign n9530 = n4723 & n4988 ;
  assign n9531 = n2085 & n4343 ;
  assign n9532 = n9530 & n9531 ;
  assign n9533 = n4766 & n4988 ;
  assign n9534 = n1817 & ~n2213 ;
  assign n9535 = n9533 & n9534 ;
  assign n9536 = n9532 | n9535 ;
  assign n9537 = n9139 & n9536 ;
  assign n9538 = x69 & ~n9215 ;
  assign n9539 = ~n8314 & n9538 ;
  assign n9540 = x71 | n9539 ;
  assign n9541 = x81 | x314 ;
  assign n9542 = n8353 | n9541 ;
  assign n9543 = n4863 | n9542 ;
  assign n9544 = n9540 & ~n9543 ;
  assign n9545 = x71 & x314 ;
  assign n9546 = ~n1244 & n9545 ;
  assign n9547 = ~n8317 & n9546 ;
  assign n9548 = ~n1353 & n9547 ;
  assign n9549 = n9544 | n9548 ;
  assign n9550 = ~n9260 & n9549 ;
  assign n9551 = ~n1279 & n1644 ;
  assign n9552 = ~x96 & n9551 ;
  assign n9553 = n8362 & n9552 ;
  assign n9554 = x198 & x589 ;
  assign n9555 = ~n2214 & n4766 ;
  assign n9556 = n9554 & n9555 ;
  assign n9557 = x210 & x589 ;
  assign n9558 = ~x221 & n4343 ;
  assign n9559 = ~x216 & n9558 ;
  assign n9560 = n4723 & n9559 ;
  assign n9561 = n9557 & n9560 ;
  assign n9562 = n9556 | n9561 ;
  assign n9563 = ~x593 & n4978 ;
  assign n9564 = n4994 & n9563 ;
  assign n9565 = n9562 & n9564 ;
  assign n9566 = x287 | n9565 ;
  assign n9567 = x39 & n9566 ;
  assign n9568 = ~n1868 & n9567 ;
  assign n9569 = n9553 | n9568 ;
  assign n9570 = ~n8366 & n9569 ;
  assign n9571 = x50 | n7170 ;
  assign n9572 = n4870 | n9571 ;
  assign n9573 = ~n1232 & n4851 ;
  assign n9574 = ~n9170 & n9573 ;
  assign n9575 = x64 | n7155 ;
  assign n9576 = n9574 & ~n9575 ;
  assign n9577 = x81 | n9576 ;
  assign n9578 = ~x199 & x200 ;
  assign n9579 = ~x299 & n9578 ;
  assign n9580 = x211 & ~x219 ;
  assign n9581 = x299 & n9580 ;
  assign n9582 = n9579 | n9581 ;
  assign n9583 = x314 & n9582 ;
  assign n9584 = ~n8328 & n9583 ;
  assign n9585 = n9577 & n9584 ;
  assign n9586 = ~n9572 & n9585 ;
  assign n9587 = n9168 | n9582 ;
  assign n9588 = n9510 & ~n9587 ;
  assign n9589 = n9574 & n9588 ;
  assign n9590 = n9586 | n9589 ;
  assign n9591 = ~n8331 & n9590 ;
  assign n9592 = x24 & ~n1260 ;
  assign n9593 = x72 & n9592 ;
  assign n9594 = x88 & ~n8313 ;
  assign n9595 = n4993 & ~n7396 ;
  assign n9596 = n9594 & n9595 ;
  assign n9597 = x98 | n1246 ;
  assign n9598 = n1242 | n9597 ;
  assign n9599 = n9596 & ~n9598 ;
  assign n9600 = n9593 | n9599 ;
  assign n9601 = ~n4904 & n9600 ;
  assign n9602 = x39 | n9601 ;
  assign n9603 = n5941 & n9533 ;
  assign n9604 = n5944 & n9530 ;
  assign n9605 = x39 & ~n9604 ;
  assign n9606 = ~n9603 & n9605 ;
  assign n9607 = n8366 | n9606 ;
  assign n9608 = n9602 & ~n9607 ;
  assign n9609 = ~x314 & x1050 ;
  assign n9610 = n7786 & ~n8328 ;
  assign n9611 = n9609 & n9610 ;
  assign n9612 = ( x39 & ~n8366 ) | ( x39 & n9611 ) | ( ~n8366 & n9611 ) ;
  assign n9613 = n7285 & n9533 ;
  assign n9614 = x299 | n9613 ;
  assign n9615 = n7296 & n9530 ;
  assign n9616 = x299 & ~n9615 ;
  assign n9617 = n9614 & ~n9616 ;
  assign n9618 = ( x39 & n8366 ) | ( x39 & ~n9617 ) | ( n8366 & ~n9617 ) ;
  assign n9619 = n9612 & ~n9618 ;
  assign n9620 = x74 & n9446 ;
  assign n9621 = ~n1529 & n5960 ;
  assign n9622 = x96 | n9621 ;
  assign n9623 = x96 | x1093 ;
  assign n9624 = n5950 & ~n9623 ;
  assign n9625 = n2111 | n5880 ;
  assign n9626 = n9624 | n9625 ;
  assign n9627 = x96 | n4694 ;
  assign n9628 = x479 & n9627 ;
  assign n9629 = n7136 | n9628 ;
  assign n9630 = n9626 | n9629 ;
  assign n9631 = n9622 & ~n9630 ;
  assign n9632 = ~n5911 & n9631 ;
  assign n9633 = n9620 | n9632 ;
  assign n9634 = ~n6785 & n9633 ;
  assign n9635 = ~n2007 & n8363 ;
  assign n9636 = ( x75 & n7113 ) | ( x75 & ~n9635 ) | ( n7113 & ~n9635 ) ;
  assign n9637 = x96 & ~x1093 ;
  assign n9638 = n1691 & n9622 ;
  assign n9639 = n9637 | n9638 ;
  assign n9640 = ~n1984 & n9639 ;
  assign n9641 = n5955 & n9640 ;
  assign n9642 = ( x75 & ~n7113 ) | ( x75 & n9641 ) | ( ~n7113 & n9641 ) ;
  assign n9643 = ~n9636 & n9642 ;
  assign n9644 = ~n1864 & n8577 ;
  assign n9645 = x252 & n1693 ;
  assign n9646 = n9644 & ~n9645 ;
  assign n9647 = ~x137 & n9646 ;
  assign n9648 = ~x137 & n1288 ;
  assign n9649 = n7130 & ~n8576 ;
  assign n9650 = x94 | n7162 ;
  assign n9651 = ~n8328 & n9650 ;
  assign n9652 = ~n9649 & n9651 ;
  assign n9653 = n1693 | n9652 ;
  assign n9654 = n7161 & ~n8338 ;
  assign n9655 = ( x252 & ~n1693 ) | ( x252 & n9654 ) | ( ~n1693 & n9654 ) ;
  assign n9656 = ( x252 & n1693 ) | ( x252 & ~n9652 ) | ( n1693 & ~n9652 ) ;
  assign n9657 = ~n9655 & n9656 ;
  assign n9658 = n9653 & ~n9657 ;
  assign n9659 = x122 & ~n9658 ;
  assign n9660 = n5950 & ~n9653 ;
  assign n9661 = n4799 | n9644 ;
  assign n9662 = ~n9657 & n9661 ;
  assign n9663 = ~n9660 & n9662 ;
  assign n9664 = x122 | n9663 ;
  assign n9665 = ~n9659 & n9664 ;
  assign n9666 = x1093 | n9665 ;
  assign n9667 = x122 | n9646 ;
  assign n9668 = ~n9659 & n9667 ;
  assign n9669 = x1093 & ~n9668 ;
  assign n9670 = n9666 & ~n9669 ;
  assign n9671 = n1288 & ~n9670 ;
  assign n9672 = n9648 | n9671 ;
  assign n9673 = ~n9647 & n9672 ;
  assign n9674 = ~x122 & n9644 ;
  assign n9675 = x1093 & ~n9652 ;
  assign n9676 = n6406 | n9675 ;
  assign n9677 = ~n9674 & n9676 ;
  assign n9678 = n9666 & ~n9677 ;
  assign n9679 = n1288 | n9678 ;
  assign n9680 = x137 | n1288 ;
  assign n9681 = n9679 & n9680 ;
  assign n9682 = x252 & x1092 ;
  assign n9683 = ~x1093 & n9682 ;
  assign n9684 = n1289 & n9683 ;
  assign n9685 = x137 | n9684 ;
  assign n9686 = n9644 & ~n9685 ;
  assign n9687 = n9681 | n9686 ;
  assign n9688 = ~n9673 & n9687 ;
  assign n9689 = n4795 | n9688 ;
  assign n9690 = n8280 & n9654 ;
  assign n9691 = n4795 & ~n9690 ;
  assign n9692 = ~x137 & n4795 ;
  assign n9693 = n9691 | n9692 ;
  assign n9694 = n9689 & ~n9693 ;
  assign n9695 = x210 | n9694 ;
  assign n9696 = ~n9671 & n9679 ;
  assign n9697 = n4795 | n9696 ;
  assign n9698 = ~n9691 & n9697 ;
  assign n9699 = x210 & ~n9698 ;
  assign n9700 = n9695 & ~n9699 ;
  assign n9701 = n1523 | n8466 ;
  assign n9702 = ~n9700 & n9701 ;
  assign n9703 = ( x210 & n9696 ) | ( x210 & n9701 ) | ( n9696 & n9701 ) ;
  assign n9704 = ( ~x210 & n9688 ) | ( ~x210 & n9701 ) | ( n9688 & n9701 ) ;
  assign n9705 = n9703 | n9704 ;
  assign n9706 = x299 & n9705 ;
  assign n9707 = ~n9702 & n9706 ;
  assign n9708 = x198 | n9694 ;
  assign n9709 = x198 & ~n9698 ;
  assign n9710 = n9708 & ~n9709 ;
  assign n9711 = n1834 | n4713 ;
  assign n9712 = ~n9710 & n9711 ;
  assign n9713 = ( x198 & n9696 ) | ( x198 & n9711 ) | ( n9696 & n9711 ) ;
  assign n9714 = ( ~x198 & n9688 ) | ( ~x198 & n9711 ) | ( n9688 & n9711 ) ;
  assign n9715 = n9713 | n9714 ;
  assign n9716 = ~x299 & n9715 ;
  assign n9717 = ~n9712 & n9716 ;
  assign n9718 = n9707 | n9717 ;
  assign n9719 = x232 & n9718 ;
  assign n9720 = ( x232 & x299 ) | ( x232 & ~n9700 ) | ( x299 & ~n9700 ) ;
  assign n9721 = ( ~x232 & x299 ) | ( ~x232 & n9710 ) | ( x299 & n9710 ) ;
  assign n9722 = ~n9720 & n9721 ;
  assign n9723 = n9719 | n9722 ;
  assign n9724 = ~n6153 & n9723 ;
  assign n9725 = x1093 | n9658 ;
  assign n9726 = ( n1288 & ~n9675 ) | ( n1288 & n9725 ) | ( ~n9675 & n9725 ) ;
  assign n9727 = n1693 & ~n9644 ;
  assign n9728 = ~n9645 & n9653 ;
  assign n9729 = ~n9727 & n9728 ;
  assign n9730 = n6406 & ~n9729 ;
  assign n9731 = n9659 | n9730 ;
  assign n9732 = ( n1288 & ~n9725 ) | ( n1288 & n9731 ) | ( ~n9725 & n9731 ) ;
  assign n9733 = n9726 & ~n9732 ;
  assign n9734 = ~n4795 & n9733 ;
  assign n9735 = n4795 & n9654 ;
  assign n9736 = ~n8282 & n9735 ;
  assign n9737 = n9734 | n9736 ;
  assign n9738 = x210 & n9737 ;
  assign n9739 = x137 | n9729 ;
  assign n9740 = x1093 | n9739 ;
  assign n9741 = x137 & ~n9725 ;
  assign n9742 = n9675 | n9741 ;
  assign n9743 = n9740 & ~n9742 ;
  assign n9744 = ~n4795 & n9743 ;
  assign n9745 = n9735 | n9744 ;
  assign n9746 = n7135 & n9692 ;
  assign n9747 = n1288 | n9746 ;
  assign n9748 = n9745 & ~n9747 ;
  assign n9749 = x137 & n9731 ;
  assign n9750 = n9739 & ~n9741 ;
  assign n9751 = ~n9749 & n9750 ;
  assign n9752 = n4795 | n9751 ;
  assign n9753 = x137 & ~n6406 ;
  assign n9754 = n1693 & ~n9753 ;
  assign n9755 = n9735 & ~n9754 ;
  assign n9756 = ( n1288 & ~n4795 ) | ( n1288 & n9755 ) | ( ~n4795 & n9755 ) ;
  assign n9757 = n9752 & n9756 ;
  assign n9758 = n9748 | n9757 ;
  assign n9759 = ~x210 & n9758 ;
  assign n9760 = n9738 | n9759 ;
  assign n9761 = n9701 & n9760 ;
  assign n9762 = ( x210 & n9701 ) | ( x210 & ~n9733 ) | ( n9701 & ~n9733 ) ;
  assign n9763 = ~n1288 & n9743 ;
  assign n9764 = n1288 & n9751 ;
  assign n9765 = n9763 | n9764 ;
  assign n9766 = ( x210 & ~n9701 ) | ( x210 & n9765 ) | ( ~n9701 & n9765 ) ;
  assign n9767 = ~n9762 & n9766 ;
  assign n9768 = x299 & ~n9767 ;
  assign n9769 = ~n9761 & n9768 ;
  assign n9770 = x198 & n9737 ;
  assign n9771 = ~x198 & n9758 ;
  assign n9772 = n9770 | n9771 ;
  assign n9773 = n9711 & n9772 ;
  assign n9774 = ( x198 & n9711 ) | ( x198 & ~n9733 ) | ( n9711 & ~n9733 ) ;
  assign n9775 = ( x198 & ~n9711 ) | ( x198 & n9765 ) | ( ~n9711 & n9765 ) ;
  assign n9776 = ~n9774 & n9775 ;
  assign n9777 = x299 | n9776 ;
  assign n9778 = n9773 | n9777 ;
  assign n9779 = ~n9769 & n9778 ;
  assign n9780 = x232 & ~n9779 ;
  assign n9781 = ( x232 & x299 ) | ( x232 & n9760 ) | ( x299 & n9760 ) ;
  assign n9782 = ( x232 & ~x299 ) | ( x232 & n9772 ) | ( ~x299 & n9772 ) ;
  assign n9783 = n9781 | n9782 ;
  assign n9784 = n6153 & n9783 ;
  assign n9785 = ~n9780 & n9784 ;
  assign n9786 = n9724 | n9785 ;
  assign n9787 = ~n8331 & n9786 ;
  assign n9788 = x86 & ~n7130 ;
  assign n9789 = ~n1342 & n9788 ;
  assign n9790 = ( x314 & n8332 ) | ( x314 & ~n9789 ) | ( n8332 & ~n9789 ) ;
  assign n9791 = ~n1338 & n1349 ;
  assign n9792 = x86 | n9791 ;
  assign n9793 = ~n4878 & n9792 ;
  assign n9794 = ~n1253 & n9793 ;
  assign n9795 = ( x314 & ~n8332 ) | ( x314 & n9794 ) | ( ~n8332 & n9794 ) ;
  assign n9796 = ~n9790 & n9795 ;
  assign n9797 = x119 & x232 ;
  assign n9798 = ~x468 & n9797 ;
  assign n9799 = x197 & ~n7212 ;
  assign n9800 = n7973 & n9799 ;
  assign n9801 = x162 | x197 ;
  assign n9802 = n7213 & n9801 ;
  assign n9803 = n4713 | n9802 ;
  assign n9804 = n9800 | n9803 ;
  assign n9805 = x163 & n9804 ;
  assign n9806 = x163 | n9800 ;
  assign n9807 = n9802 | n9806 ;
  assign n9808 = ~n9805 & n9807 ;
  assign n9809 = x232 & n9808 ;
  assign n9810 = x75 & ~n9809 ;
  assign n9811 = x100 & ~n9809 ;
  assign n9812 = n9810 | n9811 ;
  assign n9813 = x147 & n5924 ;
  assign n9814 = ~n7219 & n9813 ;
  assign n9815 = n9812 | n9814 ;
  assign n9816 = n7219 & n9809 ;
  assign n9817 = x74 & ~n9816 ;
  assign n9818 = n2057 & ~n9817 ;
  assign n9819 = ~n9815 & n9818 ;
  assign n9820 = x54 & n9815 ;
  assign n9821 = x38 | x40 ;
  assign n9822 = x38 & ~n9813 ;
  assign n9823 = x100 | n9822 ;
  assign n9824 = n9821 & ~n9823 ;
  assign n9825 = n9811 | n9824 ;
  assign n9826 = ~x75 & n9825 ;
  assign n9827 = n9810 | n9826 ;
  assign n9828 = ~x54 & n9827 ;
  assign n9829 = n9820 | n9828 ;
  assign n9830 = ~x74 & n9829 ;
  assign n9831 = n9817 | n9830 ;
  assign n9832 = n2058 & n9831 ;
  assign n9833 = n2057 | n9832 ;
  assign n9834 = x299 & ~n9808 ;
  assign n9835 = n7921 & n7922 ;
  assign n9836 = x184 | n9835 ;
  assign n9837 = ( n4713 & n9835 ) | ( n4713 & n9836 ) | ( n9835 & n9836 ) ;
  assign n9838 = ( x299 & n9836 ) | ( x299 & ~n9837 ) | ( n9836 & ~n9837 ) ;
  assign n9839 = ( ~x184 & n9836 ) | ( ~x184 & n9838 ) | ( n9836 & n9838 ) ;
  assign n9840 = x232 & n9839 ;
  assign n9841 = ~n9834 & n9840 ;
  assign n9842 = n7219 & n9841 ;
  assign n9843 = x74 & ~n9842 ;
  assign n9844 = x55 | n9843 ;
  assign n9845 = ( x187 & x299 ) | ( x187 & n5924 ) | ( x299 & n5924 ) ;
  assign n9846 = ( x147 & ~x299 ) | ( x147 & n5924 ) | ( ~x299 & n5924 ) ;
  assign n9847 = n9845 & n9846 ;
  assign n9848 = n7219 | n9847 ;
  assign n9849 = x54 & n9848 ;
  assign n9850 = ~n9842 & n9849 ;
  assign n9851 = ~x147 & x187 ;
  assign n9852 = n7253 & n9851 ;
  assign n9853 = ( x147 & ~x187 ) | ( x147 & n7256 ) | ( ~x187 & n7256 ) ;
  assign n9854 = ( x147 & x187 ) | ( x147 & n7259 ) | ( x187 & n7259 ) ;
  assign n9855 = n9853 & n9854 ;
  assign n9856 = n9852 | n9855 ;
  assign n9857 = x38 & n9856 ;
  assign n9858 = ~x32 & x95 ;
  assign n9859 = ~x479 & n9858 ;
  assign n9860 = n1278 | n1295 ;
  assign n9861 = n1272 | n9860 ;
  assign n9862 = n9859 & ~n9861 ;
  assign n9863 = x40 | n9862 ;
  assign n9864 = n7826 | n9863 ;
  assign n9865 = ~n8466 & n9864 ;
  assign n9866 = x166 & ~n4713 ;
  assign n9867 = n7829 | n9863 ;
  assign n9868 = n9866 & n9867 ;
  assign n9869 = x153 | n9868 ;
  assign n9870 = n9865 | n9869 ;
  assign n9871 = ~x210 & n7780 ;
  assign n9872 = n7778 | n9863 ;
  assign n9873 = n9871 | n9872 ;
  assign n9874 = ~n8466 & n9873 ;
  assign n9875 = n7798 | n9867 ;
  assign n9876 = n9866 & n9875 ;
  assign n9877 = x153 & ~n9876 ;
  assign n9878 = ~n9874 & n9877 ;
  assign n9879 = n9870 & ~n9878 ;
  assign n9880 = x40 & n4713 ;
  assign n9881 = x163 & ~n9880 ;
  assign n9882 = ~n9879 & n9881 ;
  assign n9883 = x160 & ~n9882 ;
  assign n9884 = x153 & n7778 ;
  assign n9885 = n7826 | n9884 ;
  assign n9886 = ~n8466 & n9885 ;
  assign n9887 = x153 & n7798 ;
  assign n9888 = n7829 | n9887 ;
  assign n9889 = n9866 & n9888 ;
  assign n9890 = ~x40 & x163 ;
  assign n9891 = ~n9889 & n9890 ;
  assign n9892 = ~n9886 & n9891 ;
  assign n9893 = x153 & ~n7789 ;
  assign n9894 = n7802 & n9893 ;
  assign n9895 = n7809 & ~n8466 ;
  assign n9896 = x40 | x163 ;
  assign n9897 = n9895 | n9896 ;
  assign n9898 = n9894 | n9897 ;
  assign n9899 = ~x160 & n9898 ;
  assign n9900 = ~n9892 & n9899 ;
  assign n9901 = n9883 | n9900 ;
  assign n9902 = ~n4713 & n9862 ;
  assign n9903 = n9898 | n9902 ;
  assign n9904 = x299 & n9903 ;
  assign n9905 = n9901 & n9904 ;
  assign n9906 = x182 & n9862 ;
  assign n9907 = ( x189 & n1863 ) | ( x189 & ~n7802 ) | ( n1863 & ~n7802 ) ;
  assign n9908 = ( x189 & ~n1863 ) | ( x189 & n7788 ) | ( ~n1863 & n7788 ) ;
  assign n9909 = ~n9907 & n9908 ;
  assign n9910 = n9906 | n9909 ;
  assign n9911 = ~n4713 & n9910 ;
  assign n9912 = x184 | n9911 ;
  assign n9913 = n7782 & ~n8477 ;
  assign n9914 = x189 & n7800 ;
  assign n9915 = ~x182 & x184 ;
  assign n9916 = ~n9914 & n9915 ;
  assign n9917 = ~n9913 & n9916 ;
  assign n9918 = n9912 & ~n9917 ;
  assign n9919 = x40 | n9918 ;
  assign n9920 = x175 & ~x299 ;
  assign n9921 = n7781 | n9872 ;
  assign n9922 = ~n8477 & n9921 ;
  assign n9923 = x189 & ~n4713 ;
  assign n9924 = n7799 | n9863 ;
  assign n9925 = n9923 & n9924 ;
  assign n9926 = x182 & x184 ;
  assign n9927 = ~n9880 & n9926 ;
  assign n9928 = ~n9925 & n9927 ;
  assign n9929 = ~n9922 & n9928 ;
  assign n9930 = n9920 & ~n9929 ;
  assign n9931 = n9919 & n9930 ;
  assign n9932 = x175 | x299 ;
  assign n9933 = x184 & x189 ;
  assign n9934 = n7814 & n9933 ;
  assign n9935 = n9906 | n9934 ;
  assign n9936 = ( x184 & x189 ) | ( x184 & ~n7816 ) | ( x189 & ~n7816 ) ;
  assign n9937 = ( x184 & ~x189 ) | ( x184 & n7809 ) | ( ~x189 & n7809 ) ;
  assign n9938 = ~n9936 & n9937 ;
  assign n9939 = n9935 | n9938 ;
  assign n9940 = ~n7470 & n9939 ;
  assign n9941 = ( x40 & ~n9932 ) | ( x40 & n9940 ) | ( ~n9932 & n9940 ) ;
  assign n9942 = n9931 | n9941 ;
  assign n9943 = n9905 | n9942 ;
  assign n9944 = ~x39 & n9943 ;
  assign n9945 = n7789 | n9861 ;
  assign n9946 = ~x189 & n7280 ;
  assign n9947 = x179 & n4731 ;
  assign n9948 = n9946 | n9947 ;
  assign n9949 = n4764 & n7285 ;
  assign n9950 = n9948 & n9949 ;
  assign n9951 = ~n9945 & n9950 ;
  assign n9952 = x40 | x299 ;
  assign n9953 = n9951 | n9952 ;
  assign n9954 = n4721 & n7296 ;
  assign n9955 = x156 & n4731 ;
  assign n9956 = ~x166 & n7280 ;
  assign n9957 = n9955 | n9956 ;
  assign n9958 = n9954 & n9957 ;
  assign n9959 = ~n9945 & n9958 ;
  assign n9960 = ~x40 & x299 ;
  assign n9961 = ~n9959 & n9960 ;
  assign n9962 = x39 & ~n9961 ;
  assign n9963 = n9953 & n9962 ;
  assign n9964 = x232 & ~n9963 ;
  assign n9965 = ~n9944 & n9964 ;
  assign n9966 = x40 | x232 ;
  assign n9967 = ~x38 & n9966 ;
  assign n9968 = ~n9965 & n9967 ;
  assign n9969 = n9857 | n9968 ;
  assign n9970 = ~n1924 & n9969 ;
  assign n9971 = x100 & ~n9841 ;
  assign n9972 = x38 & ~n9847 ;
  assign n9973 = x100 | n9972 ;
  assign n9974 = x87 & n9821 ;
  assign n9975 = ~n9973 & n9974 ;
  assign n9976 = n9971 | n9975 ;
  assign n9977 = n9970 | n9976 ;
  assign n9978 = ~n2004 & n9977 ;
  assign n9979 = x75 & ~n9841 ;
  assign n9980 = n1863 | n1983 ;
  assign n9981 = ( x179 & x299 ) | ( x179 & n5924 ) | ( x299 & n5924 ) ;
  assign n9982 = ( x156 & ~x299 ) | ( x156 & n5924 ) | ( ~x299 & n5924 ) ;
  assign n9983 = n9981 & n9982 ;
  assign n9984 = ~n9980 & n9983 ;
  assign n9985 = ~n9861 & n9984 ;
  assign n9986 = n9821 | n9985 ;
  assign n9987 = ~n9973 & n9986 ;
  assign n9988 = n9971 | n9987 ;
  assign n9989 = n7679 & n9988 ;
  assign n9990 = n9979 | n9989 ;
  assign n9991 = n9978 | n9990 ;
  assign n9992 = ~x54 & n9991 ;
  assign n9993 = n9850 | n9992 ;
  assign n9994 = ~x74 & n9993 ;
  assign n9995 = n9844 | n9994 ;
  assign n9996 = x55 & ~n9817 ;
  assign n9997 = x163 & x232 ;
  assign n9998 = x92 | n1983 ;
  assign n9999 = n9997 & ~n9998 ;
  assign n10000 = ~n9945 & n9999 ;
  assign n10001 = n9821 | n10000 ;
  assign n10002 = x75 | n9823 ;
  assign n10003 = n10001 & ~n10002 ;
  assign n10004 = n9812 | n10003 ;
  assign n10005 = ~x54 & n10004 ;
  assign n10006 = n9820 | n10005 ;
  assign n10007 = ~x74 & n10006 ;
  assign n10008 = n9996 & ~n10007 ;
  assign n10009 = n2058 | n10008 ;
  assign n10010 = n9995 & ~n10009 ;
  assign n10011 = n9833 | n10010 ;
  assign n10012 = ~n9819 & n10011 ;
  assign n10013 = x34 | n8070 ;
  assign n10014 = ( x79 & n10012 ) | ( x79 & ~n10013 ) | ( n10012 & ~n10013 ) ;
  assign n10015 = ~x40 & n7439 ;
  assign n10016 = x95 | n10015 ;
  assign n10017 = ~x40 & n7456 ;
  assign n10018 = x166 & n10017 ;
  assign n10019 = n10016 | n10018 ;
  assign n10020 = n4713 | n7481 ;
  assign n10021 = n10019 & ~n10020 ;
  assign n10022 = x153 | n10021 ;
  assign n10023 = ~x40 & n7517 ;
  assign n10024 = x95 | n10023 ;
  assign n10025 = x166 & n10024 ;
  assign n10026 = ~n10020 & n10025 ;
  assign n10027 = n7480 & ~n8466 ;
  assign n10028 = x153 & ~n10027 ;
  assign n10029 = ~n10026 & n10028 ;
  assign n10030 = x160 & ~n10029 ;
  assign n10031 = n10022 & n10030 ;
  assign n10032 = x153 | n10019 ;
  assign n10033 = n1491 | n7481 ;
  assign n10034 = n7339 | n7340 ;
  assign n10035 = n10033 & n10034 ;
  assign n10036 = ~n9610 & n10024 ;
  assign n10037 = x153 & ~n10025 ;
  assign n10038 = ~n10036 & n10037 ;
  assign n10039 = x160 | n4713 ;
  assign n10040 = n10038 | n10039 ;
  assign n10041 = n10035 | n10040 ;
  assign n10042 = n10032 & ~n10041 ;
  assign n10043 = x163 & ~n10042 ;
  assign n10044 = ~n10031 & n10043 ;
  assign n10045 = ~x40 & n7585 ;
  assign n10046 = x95 | n10045 ;
  assign n10047 = ~n10035 & n10046 ;
  assign n10048 = x166 & n10047 ;
  assign n10049 = ~x40 & n7415 ;
  assign n10050 = x32 | n10049 ;
  assign n10051 = ~n7482 & n10050 ;
  assign n10052 = x95 | n10051 ;
  assign n10053 = ~n10035 & n10052 ;
  assign n10054 = ( x210 & n8466 ) | ( x210 & ~n10053 ) | ( n8466 & ~n10053 ) ;
  assign n10055 = ~n7498 & n10050 ;
  assign n10056 = x95 | n10055 ;
  assign n10057 = ~n10035 & n10056 ;
  assign n10058 = ( x210 & ~n8466 ) | ( x210 & n10057 ) | ( ~n8466 & n10057 ) ;
  assign n10059 = ~n10054 & n10058 ;
  assign n10060 = x153 | n10059 ;
  assign n10061 = n10048 | n10060 ;
  assign n10062 = x95 | n7530 ;
  assign n10063 = ~n10035 & n10062 ;
  assign n10064 = ( ~x210 & n9866 ) | ( ~x210 & n10063 ) | ( n9866 & n10063 ) ;
  assign n10065 = n7536 & ~n10035 ;
  assign n10066 = ( x210 & n9866 ) | ( x210 & n10065 ) | ( n9866 & n10065 ) ;
  assign n10067 = n10064 & n10066 ;
  assign n10068 = x153 & ~n10067 ;
  assign n10069 = n7500 & ~n10035 ;
  assign n10070 = ( x210 & ~n8466 ) | ( x210 & n10069 ) | ( ~n8466 & n10069 ) ;
  assign n10071 = n7495 & ~n10035 ;
  assign n10072 = ( x210 & n8466 ) | ( x210 & ~n10071 ) | ( n8466 & ~n10071 ) ;
  assign n10073 = n10070 & ~n10072 ;
  assign n10074 = n10068 & ~n10073 ;
  assign n10075 = x160 | n10074 ;
  assign n10076 = n10061 & ~n10075 ;
  assign n10077 = n9866 & n10045 ;
  assign n10078 = ~n7481 & n10056 ;
  assign n10079 = ( x210 & ~n8466 ) | ( x210 & n10078 ) | ( ~n8466 & n10078 ) ;
  assign n10080 = ~n7481 & n10052 ;
  assign n10081 = ( x210 & n8466 ) | ( x210 & ~n10080 ) | ( n8466 & ~n10080 ) ;
  assign n10082 = n10079 & ~n10081 ;
  assign n10083 = x153 | n10082 ;
  assign n10084 = n10077 | n10083 ;
  assign n10085 = ( x210 & ~n7496 ) | ( x210 & n8466 ) | ( ~n7496 & n8466 ) ;
  assign n10086 = ( x210 & n7501 ) | ( x210 & ~n8466 ) | ( n7501 & ~n8466 ) ;
  assign n10087 = ~n10085 & n10086 ;
  assign n10088 = x153 & ~n10087 ;
  assign n10089 = ( x210 & n7537 ) | ( x210 & n9866 ) | ( n7537 & n9866 ) ;
  assign n10090 = ~n7481 & n10062 ;
  assign n10091 = ( ~x210 & n9866 ) | ( ~x210 & n10090 ) | ( n9866 & n10090 ) ;
  assign n10092 = n10089 & n10091 ;
  assign n10093 = n10088 & ~n10092 ;
  assign n10094 = x160 & ~n10093 ;
  assign n10095 = n10084 & n10094 ;
  assign n10096 = x163 | n10095 ;
  assign n10097 = n10076 | n10096 ;
  assign n10098 = ~n10044 & n10097 ;
  assign n10099 = n4713 & n10047 ;
  assign n10100 = x299 & ~n10099 ;
  assign n10101 = ~n10098 & n10100 ;
  assign n10102 = ~x40 & n7472 ;
  assign n10103 = x95 | n10102 ;
  assign n10104 = ~n10035 & n10103 ;
  assign n10105 = n4713 & n10104 ;
  assign n10106 = x189 & n10017 ;
  assign n10107 = n10016 | n10106 ;
  assign n10108 = ~x182 & n10035 ;
  assign n10109 = x182 & n7481 ;
  assign n10110 = n4713 | n10109 ;
  assign n10111 = n10108 | n10110 ;
  assign n10112 = n10107 & ~n10111 ;
  assign n10113 = x184 & ~n10112 ;
  assign n10114 = n9923 & n10102 ;
  assign n10115 = x182 & ~x184 ;
  assign n10116 = ( x198 & ~n8477 ) | ( x198 & n10078 ) | ( ~n8477 & n10078 ) ;
  assign n10117 = ( x198 & n8477 ) | ( x198 & ~n10080 ) | ( n8477 & ~n10080 ) ;
  assign n10118 = n10116 & ~n10117 ;
  assign n10119 = n10115 & ~n10118 ;
  assign n10120 = ~n10114 & n10119 ;
  assign n10121 = n10113 | n10120 ;
  assign n10122 = ~n9932 & n10121 ;
  assign n10123 = n7503 & ~n8477 ;
  assign n10124 = x182 & ~n10123 ;
  assign n10125 = ( x198 & n7537 ) | ( x198 & n9923 ) | ( n7537 & n9923 ) ;
  assign n10126 = ( ~x198 & n9923 ) | ( ~x198 & n10090 ) | ( n9923 & n10090 ) ;
  assign n10127 = n10125 & n10126 ;
  assign n10128 = n10124 & ~n10127 ;
  assign n10129 = ( x198 & n9923 ) | ( x198 & n10065 ) | ( n9923 & n10065 ) ;
  assign n10130 = ( ~x198 & n9923 ) | ( ~x198 & n10063 ) | ( n9923 & n10063 ) ;
  assign n10131 = n10129 & n10130 ;
  assign n10132 = x182 | n10131 ;
  assign n10133 = ~n10128 & n10132 ;
  assign n10134 = x95 & ~x182 ;
  assign n10135 = n7503 | n10134 ;
  assign n10136 = n8477 | n10035 ;
  assign n10137 = n10135 & ~n10136 ;
  assign n10138 = n10133 | n10137 ;
  assign n10139 = ~x184 & n10138 ;
  assign n10140 = x184 & ~n4713 ;
  assign n10141 = ~x95 & x189 ;
  assign n10142 = n1236 | n10141 ;
  assign n10143 = n10023 & n10142 ;
  assign n10144 = n10134 | n10143 ;
  assign n10145 = n10140 & n10144 ;
  assign n10146 = ~n10108 & n10145 ;
  assign n10147 = n9920 & ~n10146 ;
  assign n10148 = ~n10139 & n10147 ;
  assign n10149 = n10122 | n10148 ;
  assign n10150 = ~n10105 & n10149 ;
  assign n10151 = n8477 & n10104 ;
  assign n10152 = x182 | x184 ;
  assign n10153 = n9932 | n10152 ;
  assign n10154 = ( x198 & n8477 ) | ( x198 & ~n10053 ) | ( n8477 & ~n10053 ) ;
  assign n10155 = ( x198 & ~n8477 ) | ( x198 & n10057 ) | ( ~n8477 & n10057 ) ;
  assign n10156 = ~n10154 & n10155 ;
  assign n10157 = n10153 | n10156 ;
  assign n10158 = n10151 | n10157 ;
  assign n10159 = ~n10150 & n10158 ;
  assign n10160 = ~n10101 & n10159 ;
  assign n10161 = x232 & ~n10160 ;
  assign n10162 = ( x232 & x299 ) | ( x232 & n10047 ) | ( x299 & n10047 ) ;
  assign n10163 = ( x232 & ~x299 ) | ( x232 & n10104 ) | ( ~x299 & n10104 ) ;
  assign n10164 = n10162 | n10163 ;
  assign n10165 = ~x39 & n10164 ;
  assign n10166 = ~n10161 & n10165 ;
  assign n10167 = n7285 | n7480 ;
  assign n10168 = ~x40 & n7284 ;
  assign n10169 = x189 | n10168 ;
  assign n10170 = n1236 | n7288 ;
  assign n10171 = ~n7470 & n10170 ;
  assign n10172 = n4751 & n7480 ;
  assign n10173 = n1236 | n7282 ;
  assign n10174 = ~x40 & n10173 ;
  assign n10175 = n4714 & n10174 ;
  assign n10176 = n10172 | n10175 ;
  assign n10177 = n10171 | n10176 ;
  assign n10178 = x189 & n4764 ;
  assign n10179 = ~n10177 & n10178 ;
  assign n10180 = n10169 & ~n10179 ;
  assign n10181 = x179 & ~n10180 ;
  assign n10182 = n4764 | n10168 ;
  assign n10183 = ~n4751 & n10174 ;
  assign n10184 = n10172 | n10183 ;
  assign n10185 = ~x179 & n4764 ;
  assign n10186 = ( x189 & n10184 ) | ( x189 & ~n10185 ) | ( n10184 & ~n10185 ) ;
  assign n10187 = n1236 | n7299 ;
  assign n10188 = ~n7470 & n10187 ;
  assign n10189 = n10176 | n10188 ;
  assign n10190 = ( x189 & n10185 ) | ( x189 & ~n10189 ) | ( n10185 & ~n10189 ) ;
  assign n10191 = ~n10186 & n10190 ;
  assign n10192 = n10182 & ~n10191 ;
  assign n10193 = ~n10181 & n10192 ;
  assign n10194 = n7285 & ~n10193 ;
  assign n10195 = n10167 & ~n10194 ;
  assign n10196 = x299 | n10195 ;
  assign n10197 = ~n7296 & n7480 ;
  assign n10198 = x299 & ~n10197 ;
  assign n10199 = x166 & n4721 ;
  assign n10200 = ( n7296 & n10168 ) | ( n7296 & n10199 ) | ( n10168 & n10199 ) ;
  assign n10201 = ( n7296 & n10177 ) | ( n7296 & ~n10199 ) | ( n10177 & ~n10199 ) ;
  assign n10202 = n10200 & n10201 ;
  assign n10203 = n10198 & ~n10202 ;
  assign n10204 = n10196 & ~n10203 ;
  assign n10205 = x156 & x232 ;
  assign n10206 = ~n10204 & n10205 ;
  assign n10207 = ~x166 & n4721 ;
  assign n10208 = ( n7296 & n10189 ) | ( n7296 & ~n10207 ) | ( n10189 & ~n10207 ) ;
  assign n10209 = n4721 | n10168 ;
  assign n10210 = n4721 & ~n10184 ;
  assign n10211 = n10209 & ~n10210 ;
  assign n10212 = ( n7296 & n10207 ) | ( n7296 & n10211 ) | ( n10207 & n10211 ) ;
  assign n10213 = n10208 & n10212 ;
  assign n10214 = n10198 & ~n10213 ;
  assign n10215 = n10196 & ~n10214 ;
  assign n10216 = ~x156 & x232 ;
  assign n10217 = ~n10215 & n10216 ;
  assign n10218 = n4764 & ~n10184 ;
  assign n10219 = n10182 & ~n10218 ;
  assign n10220 = n7285 & ~n10219 ;
  assign n10221 = ~x299 & n10167 ;
  assign n10222 = ~n10220 & n10221 ;
  assign n10223 = n7298 & n10211 ;
  assign n10224 = n10222 | n10223 ;
  assign n10225 = ( x39 & n8469 ) | ( x39 & n10224 ) | ( n8469 & n10224 ) ;
  assign n10226 = ~n10217 & n10225 ;
  assign n10227 = ~n10206 & n10226 ;
  assign n10228 = x38 | n10227 ;
  assign n10229 = n10166 | n10228 ;
  assign n10230 = ~n9857 & n10229 ;
  assign n10231 = n1924 | n10230 ;
  assign n10232 = x87 & n1236 ;
  assign n10233 = ~n9821 & n10232 ;
  assign n10234 = n9973 | n10233 ;
  assign n10235 = x87 & ~n10234 ;
  assign n10236 = n9971 | n10235 ;
  assign n10237 = n10231 & ~n10236 ;
  assign n10238 = n2004 | n10237 ;
  assign n10239 = x39 & ~n7480 ;
  assign n10240 = n7858 | n10239 ;
  assign n10241 = ~n1236 & n7278 ;
  assign n10242 = x40 | n10241 ;
  assign n10243 = ~n1236 & n9983 ;
  assign n10244 = n10242 | n10243 ;
  assign n10245 = ~x39 & n10244 ;
  assign n10246 = n10240 | n10245 ;
  assign n10247 = ~n10234 & n10246 ;
  assign n10248 = n9971 | n10247 ;
  assign n10249 = n7679 & n10248 ;
  assign n10250 = n9979 | n10249 ;
  assign n10251 = n10238 & ~n10250 ;
  assign n10252 = x54 | n10251 ;
  assign n10253 = ~n9850 & n10252 ;
  assign n10254 = x74 | n10253 ;
  assign n10255 = ~n9844 & n10254 ;
  assign n10256 = n4713 & ~n7278 ;
  assign n10257 = n7265 | n10256 ;
  assign n10258 = n9997 & ~n10257 ;
  assign n10259 = n10242 | n10258 ;
  assign n10260 = ~x39 & n10259 ;
  assign n10261 = n10240 | n10260 ;
  assign n10262 = n9823 | n10233 ;
  assign n10263 = n10261 & ~n10262 ;
  assign n10264 = n9811 | n10263 ;
  assign n10265 = ~n2004 & n10264 ;
  assign n10266 = n7674 & ~n9825 ;
  assign n10267 = n7679 & ~n10266 ;
  assign n10268 = n9810 | n10267 ;
  assign n10269 = n10265 | n10268 ;
  assign n10270 = ~x54 & n10269 ;
  assign n10271 = n9820 | n10270 ;
  assign n10272 = ~x74 & n10271 ;
  assign n10273 = n9996 & ~n10272 ;
  assign n10274 = n2058 | n10273 ;
  assign n10275 = n10255 | n10274 ;
  assign n10276 = n7734 | n9833 ;
  assign n10277 = n10275 & ~n10276 ;
  assign n10278 = n9819 | n10277 ;
  assign n10279 = ( x79 & n10013 ) | ( x79 & n10278 ) | ( n10013 & n10278 ) ;
  assign n10280 = ~n10014 & n10279 ;
  assign n10281 = ~x79 & n7207 ;
  assign n10282 = ( n10012 & n10013 ) | ( n10012 & n10281 ) | ( n10013 & n10281 ) ;
  assign n10283 = ( ~n10013 & n10278 ) | ( ~n10013 & n10281 ) | ( n10278 & n10281 ) ;
  assign n10284 = ~n10282 & n10283 ;
  assign n10285 = n10280 | n10284 ;
  assign n10286 = x98 & x1092 ;
  assign n10287 = x1093 & n10286 ;
  assign n10288 = ~x567 & n1290 ;
  assign n10289 = n10287 | n10288 ;
  assign n10290 = n6278 & ~n10289 ;
  assign n10291 = x588 & ~n10290 ;
  assign n10292 = x592 & n10289 ;
  assign n10293 = n5880 & ~n10289 ;
  assign n10294 = n5880 | n10288 ;
  assign n10295 = x75 & n10287 ;
  assign n10296 = x1091 & n10287 ;
  assign n10297 = x110 | n1252 ;
  assign n10298 = x86 | x88 ;
  assign n10299 = n1215 | n10298 ;
  assign n10300 = n8566 | n10299 ;
  assign n10301 = n10297 | n10300 ;
  assign n10302 = n5892 | n10301 ;
  assign n10303 = n5900 | n10302 ;
  assign n10304 = x51 & ~n10303 ;
  assign n10305 = ( x90 & x93 ) | ( x90 & x841 ) | ( x93 & x841 ) ;
  assign n10306 = ( x90 & x93 ) | ( x90 & ~n1526 ) | ( x93 & ~n1526 ) ;
  assign n10307 = ~n10305 & n10306 ;
  assign n10308 = ~n10302 & n10307 ;
  assign n10309 = n10304 | n10308 ;
  assign n10310 = x824 & x950 ;
  assign n10311 = ~n5904 & n10310 ;
  assign n10312 = n10309 & n10311 ;
  assign n10313 = x98 | n10312 ;
  assign n10314 = x1092 & n10313 ;
  assign n10315 = n10296 | n10314 ;
  assign n10316 = n5995 | n10296 ;
  assign n10317 = ~n1984 & n10316 ;
  assign n10318 = n10315 & n10317 ;
  assign n10319 = ~n1865 & n10310 ;
  assign n10320 = ~n10303 & n10319 ;
  assign n10321 = x98 | n10320 ;
  assign n10322 = x1092 & n10321 ;
  assign n10323 = n10296 | n10322 ;
  assign n10324 = n6016 & n10316 ;
  assign n10325 = n10323 & n10324 ;
  assign n10326 = n1976 & n10287 ;
  assign n10327 = n10325 | n10326 ;
  assign n10328 = n10318 | n10327 ;
  assign n10329 = ~x75 & n10328 ;
  assign n10330 = n10295 | n10329 ;
  assign n10331 = x567 & n10330 ;
  assign n10332 = n10294 | n10331 ;
  assign n10333 = ~n10293 & n10332 ;
  assign n10334 = ~x592 & n10333 ;
  assign n10335 = n10292 | n10334 ;
  assign n10336 = n6824 & ~n10335 ;
  assign n10337 = ~x1196 & n10289 ;
  assign n10338 = n6824 | n10337 ;
  assign n10339 = ~x443 & n10289 ;
  assign n10340 = x443 & n10335 ;
  assign n10341 = n10339 | n10340 ;
  assign n10342 = n6903 | n10341 ;
  assign n10343 = x443 & n10289 ;
  assign n10344 = ~x443 & n10335 ;
  assign n10345 = n10343 | n10344 ;
  assign n10346 = n6903 & ~n10345 ;
  assign n10347 = n10342 & ~n10346 ;
  assign n10348 = x435 & ~n10347 ;
  assign n10349 = ( x436 & x444 ) | ( x436 & n10341 ) | ( x444 & n10341 ) ;
  assign n10350 = ( ~x444 & n10345 ) | ( ~x444 & n10349 ) | ( n10345 & n10349 ) ;
  assign n10351 = ( ~x436 & n10349 ) | ( ~x436 & n10350 ) | ( n10349 & n10350 ) ;
  assign n10352 = x435 | n10351 ;
  assign n10353 = ~n10348 & n10352 ;
  assign n10354 = ( x429 & n6842 ) | ( x429 & ~n10353 ) | ( n6842 & ~n10353 ) ;
  assign n10355 = x435 | n10347 ;
  assign n10356 = x435 & ~n10351 ;
  assign n10357 = n10355 & ~n10356 ;
  assign n10358 = ( x429 & ~n6842 ) | ( x429 & n10357 ) | ( ~n6842 & n10357 ) ;
  assign n10359 = n10354 & ~n10358 ;
  assign n10360 = x1196 & ~n10359 ;
  assign n10361 = ( x429 & n6842 ) | ( x429 & n10353 ) | ( n6842 & n10353 ) ;
  assign n10362 = ( ~x429 & n6842 ) | ( ~x429 & n10357 ) | ( n6842 & n10357 ) ;
  assign n10363 = n10361 | n10362 ;
  assign n10364 = n10360 & n10363 ;
  assign n10365 = n10338 | n10364 ;
  assign n10366 = ~n10336 & n10365 ;
  assign n10367 = x428 | n10366 ;
  assign n10368 = x428 & ~n10335 ;
  assign n10369 = n10367 & ~n10368 ;
  assign n10370 = x427 | n10369 ;
  assign n10371 = x428 & ~n10366 ;
  assign n10372 = x428 | n10335 ;
  assign n10373 = ~n10371 & n10372 ;
  assign n10374 = x427 & ~n10373 ;
  assign n10375 = n10370 & ~n10374 ;
  assign n10376 = x430 & ~n10375 ;
  assign n10377 = x427 | n10373 ;
  assign n10378 = x427 & ~n10369 ;
  assign n10379 = n10377 & ~n10378 ;
  assign n10380 = x430 | n10379 ;
  assign n10381 = ~n10376 & n10380 ;
  assign n10382 = x426 & ~n10381 ;
  assign n10383 = x430 & ~n10379 ;
  assign n10384 = x430 | n10375 ;
  assign n10385 = ~n10383 & n10384 ;
  assign n10386 = x426 | n10385 ;
  assign n10387 = ~n10382 & n10386 ;
  assign n10388 = x445 & ~n10387 ;
  assign n10389 = x426 & ~n10385 ;
  assign n10390 = x426 | n10381 ;
  assign n10391 = ~n10389 & n10390 ;
  assign n10392 = x445 | n10391 ;
  assign n10393 = ~n10388 & n10392 ;
  assign n10394 = ( x448 & n6788 ) | ( x448 & n10393 ) | ( n6788 & n10393 ) ;
  assign n10395 = x445 & ~n10391 ;
  assign n10396 = x445 | n10387 ;
  assign n10397 = ~n10395 & n10396 ;
  assign n10398 = ( ~x448 & n6788 ) | ( ~x448 & n10397 ) | ( n6788 & n10397 ) ;
  assign n10399 = n10394 | n10398 ;
  assign n10400 = x1199 & n10399 ;
  assign n10401 = ( x448 & n6788 ) | ( x448 & ~n10393 ) | ( n6788 & ~n10393 ) ;
  assign n10402 = ( x448 & ~n6788 ) | ( x448 & n10397 ) | ( ~n6788 & n10397 ) ;
  assign n10403 = n10401 & ~n10402 ;
  assign n10404 = n10400 & ~n10403 ;
  assign n10405 = ~x1199 & n10366 ;
  assign n10406 = n6278 | n10405 ;
  assign n10407 = n10404 | n10406 ;
  assign n10408 = n10291 & n10407 ;
  assign n10409 = x591 & n10289 ;
  assign n10410 = x590 & ~n10409 ;
  assign n10411 = n6973 | n10289 ;
  assign n10412 = n6973 & ~n10335 ;
  assign n10413 = n10411 & ~n10412 ;
  assign n10414 = x1198 & ~n10413 ;
  assign n10415 = x1198 | n10337 ;
  assign n10416 = n6041 | n10289 ;
  assign n10417 = n6041 & ~n10335 ;
  assign n10418 = n10416 & ~n10417 ;
  assign n10419 = x355 & ~n10418 ;
  assign n10420 = ( x452 & x455 ) | ( x452 & n10289 ) | ( x455 & n10289 ) ;
  assign n10421 = ( ~x455 & n10335 ) | ( ~x455 & n10420 ) | ( n10335 & n10420 ) ;
  assign n10422 = ( ~x452 & n10420 ) | ( ~x452 & n10421 ) | ( n10420 & n10421 ) ;
  assign n10423 = x355 | n10422 ;
  assign n10424 = ~n10419 & n10423 ;
  assign n10425 = ( x458 & n6050 ) | ( x458 & ~n10424 ) | ( n6050 & ~n10424 ) ;
  assign n10426 = x355 | n10418 ;
  assign n10427 = x355 & ~n10422 ;
  assign n10428 = n10426 & ~n10427 ;
  assign n10429 = ( x458 & ~n6050 ) | ( x458 & n10428 ) | ( ~n6050 & n10428 ) ;
  assign n10430 = n10425 & ~n10429 ;
  assign n10431 = x1196 & ~n10430 ;
  assign n10432 = ( ~x458 & n6050 ) | ( ~x458 & n10428 ) | ( n6050 & n10428 ) ;
  assign n10433 = ( x458 & n6050 ) | ( x458 & n10424 ) | ( n6050 & n10424 ) ;
  assign n10434 = n10432 | n10433 ;
  assign n10435 = n10431 & n10434 ;
  assign n10436 = n10415 | n10435 ;
  assign n10437 = ~n10414 & n10436 ;
  assign n10438 = n6115 | n10437 ;
  assign n10439 = n6115 & ~n10335 ;
  assign n10440 = n10438 & ~n10439 ;
  assign n10441 = ~n6119 & n10440 ;
  assign n10442 = x1199 & n10335 ;
  assign n10443 = ~x351 & n10442 ;
  assign n10444 = n10441 | n10443 ;
  assign n10445 = ~x461 & n10444 ;
  assign n10446 = ~n6125 & n10440 ;
  assign n10447 = x351 & n10442 ;
  assign n10448 = n10446 | n10447 ;
  assign n10449 = x461 & n10448 ;
  assign n10450 = n10445 | n10449 ;
  assign n10451 = ~x357 & n10450 ;
  assign n10452 = ~x461 & n10448 ;
  assign n10453 = x461 & n10444 ;
  assign n10454 = n10452 | n10453 ;
  assign n10455 = x357 & n10454 ;
  assign n10456 = n10451 | n10455 ;
  assign n10457 = ~x356 & n10456 ;
  assign n10458 = ~x357 & n10454 ;
  assign n10459 = x357 & n10450 ;
  assign n10460 = n10458 | n10459 ;
  assign n10461 = x356 & n10460 ;
  assign n10462 = n10457 | n10461 ;
  assign n10463 = ( x354 & n5876 ) | ( x354 & n10462 ) | ( n5876 & n10462 ) ;
  assign n10464 = ~x356 & n10460 ;
  assign n10465 = x356 & n10456 ;
  assign n10466 = n10464 | n10465 ;
  assign n10467 = ( ~x354 & n5876 ) | ( ~x354 & n10466 ) | ( n5876 & n10466 ) ;
  assign n10468 = n10463 | n10467 ;
  assign n10469 = ~x591 & n10468 ;
  assign n10470 = ( x354 & n5876 ) | ( x354 & ~n10462 ) | ( n5876 & ~n10462 ) ;
  assign n10471 = ( x354 & ~n5876 ) | ( x354 & n10466 ) | ( ~n5876 & n10466 ) ;
  assign n10472 = n10470 & ~n10471 ;
  assign n10473 = n10469 & ~n10472 ;
  assign n10474 = n10410 & ~n10473 ;
  assign n10475 = x1197 | n6295 ;
  assign n10476 = n10335 & n10475 ;
  assign n10477 = n6678 & ~n10293 ;
  assign n10478 = ~x411 & n10286 ;
  assign n10479 = n6308 | n10478 ;
  assign n10480 = x411 & n10314 ;
  assign n10481 = n10479 | n10480 ;
  assign n10482 = n6308 & ~n10286 ;
  assign n10483 = n6310 | n10482 ;
  assign n10484 = ~x411 & n10314 ;
  assign n10485 = n10483 & ~n10484 ;
  assign n10486 = n10481 & ~n10485 ;
  assign n10487 = n10296 | n10486 ;
  assign n10488 = n10317 & n10487 ;
  assign n10489 = x411 & ~n10483 ;
  assign n10490 = ( x411 & ~n10322 ) | ( x411 & n10483 ) | ( ~n10322 & n10483 ) ;
  assign n10491 = ( n10479 & n10489 ) | ( n10479 & ~n10490 ) | ( n10489 & ~n10490 ) ;
  assign n10492 = n10296 | n10491 ;
  assign n10493 = n10324 & n10492 ;
  assign n10494 = n10326 | n10493 ;
  assign n10495 = n10488 | n10494 ;
  assign n10496 = ~x75 & n10495 ;
  assign n10497 = n10295 | n10496 ;
  assign n10498 = x567 & n10497 ;
  assign n10499 = n10294 | n10498 ;
  assign n10500 = n10477 & n10499 ;
  assign n10501 = n10292 | n10337 ;
  assign n10502 = x1199 | n10501 ;
  assign n10503 = n10500 | n10502 ;
  assign n10504 = n6341 & n10325 ;
  assign n10505 = n6341 & n10314 ;
  assign n10506 = ~n6341 & n10286 ;
  assign n10507 = n10505 | n10506 ;
  assign n10508 = n10318 & n10507 ;
  assign n10509 = n10504 | n10508 ;
  assign n10510 = n10495 | n10509 ;
  assign n10511 = n10477 & n10510 ;
  assign n10512 = n6341 & n10322 ;
  assign n10513 = n10506 | n10512 ;
  assign n10514 = n10325 & n10513 ;
  assign n10515 = n10326 | n10514 ;
  assign n10516 = n10508 | n10515 ;
  assign n10517 = n6686 | n10293 ;
  assign n10518 = n10516 & ~n10517 ;
  assign n10519 = n10511 | n10518 ;
  assign n10520 = ~x75 & x567 ;
  assign n10521 = n10519 & n10520 ;
  assign n10522 = n6318 | n10294 ;
  assign n10523 = n10289 & n10522 ;
  assign n10524 = x1199 & ~n10523 ;
  assign n10525 = ~n10521 & n10524 ;
  assign n10526 = n6295 | n10525 ;
  assign n10527 = n10503 & ~n10526 ;
  assign n10528 = ~x1197 & n10527 ;
  assign n10529 = n10476 | n10528 ;
  assign n10530 = ~x333 & n10529 ;
  assign n10531 = n6295 & n10335 ;
  assign n10532 = n10527 | n10531 ;
  assign n10533 = x333 & n10532 ;
  assign n10534 = n10530 | n10533 ;
  assign n10535 = ~x391 & n10534 ;
  assign n10536 = x333 & n10529 ;
  assign n10537 = ~x333 & n10532 ;
  assign n10538 = n10536 | n10537 ;
  assign n10539 = x391 & n10538 ;
  assign n10540 = n10535 | n10539 ;
  assign n10541 = ~x392 & n10540 ;
  assign n10542 = ~x391 & n10538 ;
  assign n10543 = x391 & n10534 ;
  assign n10544 = n10542 | n10543 ;
  assign n10545 = x392 & n10544 ;
  assign n10546 = n10541 | n10545 ;
  assign n10547 = ( x393 & n6588 ) | ( x393 & ~n10546 ) | ( n6588 & ~n10546 ) ;
  assign n10548 = ~x392 & n10544 ;
  assign n10549 = x392 & n10540 ;
  assign n10550 = n10548 | n10549 ;
  assign n10551 = ( x393 & ~n6588 ) | ( x393 & n10550 ) | ( ~n6588 & n10550 ) ;
  assign n10552 = n10547 & ~n10551 ;
  assign n10553 = x591 & ~n10552 ;
  assign n10554 = ( ~x393 & n6588 ) | ( ~x393 & n10550 ) | ( n6588 & n10550 ) ;
  assign n10555 = ( x393 & n6588 ) | ( x393 & n10546 ) | ( n6588 & n10546 ) ;
  assign n10556 = n10554 | n10555 ;
  assign n10557 = n10553 & n10556 ;
  assign n10558 = ~x590 & x591 ;
  assign n10559 = ~x592 & n10289 ;
  assign n10560 = x592 & n10333 ;
  assign n10561 = n10559 | n10560 ;
  assign n10562 = n7006 & ~n10561 ;
  assign n10563 = n7006 | n10289 ;
  assign n10564 = x1199 & n10563 ;
  assign n10565 = ~n10562 & n10564 ;
  assign n10566 = ~x1197 & n10289 ;
  assign n10567 = n6169 | n10566 ;
  assign n10568 = ( x367 & n6181 ) | ( x367 & ~n6187 ) | ( n6181 & ~n6187 ) ;
  assign n10569 = ( ~x367 & n6187 ) | ( ~x367 & n10568 ) | ( n6187 & n10568 ) ;
  assign n10570 = ( ~n6181 & n10568 ) | ( ~n6181 & n10569 ) | ( n10568 & n10569 ) ;
  assign n10571 = ( x1197 & n10561 ) | ( x1197 & ~n10570 ) | ( n10561 & ~n10570 ) ;
  assign n10572 = ( x1197 & n10289 ) | ( x1197 & n10570 ) | ( n10289 & n10570 ) ;
  assign n10573 = n10571 & n10572 ;
  assign n10574 = n10567 | n10573 ;
  assign n10575 = n6169 & ~n10561 ;
  assign n10576 = x1199 | n10575 ;
  assign n10577 = n10574 & ~n10576 ;
  assign n10578 = n10565 | n10577 ;
  assign n10579 = ~x374 & n10578 ;
  assign n10580 = ~x1198 & n10578 ;
  assign n10581 = x1198 & n10561 ;
  assign n10582 = n10580 | n10581 ;
  assign n10583 = x374 & n10582 ;
  assign n10584 = n10579 | n10583 ;
  assign n10585 = ( x370 & ~x371 ) | ( x370 & n6574 ) | ( ~x371 & n6574 ) ;
  assign n10586 = ( ~x370 & x371 ) | ( ~x370 & n10585 ) | ( x371 & n10585 ) ;
  assign n10587 = ( ~n6574 & n10585 ) | ( ~n6574 & n10586 ) | ( n10585 & n10586 ) ;
  assign n10588 = ( x369 & n10584 ) | ( x369 & ~n10587 ) | ( n10584 & ~n10587 ) ;
  assign n10589 = ~x374 & n10582 ;
  assign n10590 = x374 & n10578 ;
  assign n10591 = n10589 | n10590 ;
  assign n10592 = ( x369 & n10587 ) | ( x369 & ~n10591 ) | ( n10587 & ~n10591 ) ;
  assign n10593 = ~n10588 & n10592 ;
  assign n10594 = ( x369 & n10587 ) | ( x369 & n10591 ) | ( n10587 & n10591 ) ;
  assign n10595 = ( ~x369 & n10584 ) | ( ~x369 & n10587 ) | ( n10584 & n10587 ) ;
  assign n10596 = n10594 | n10595 ;
  assign n10597 = ~n10593 & n10596 ;
  assign n10598 = ( x590 & ~n10558 ) | ( x590 & n10597 ) | ( ~n10558 & n10597 ) ;
  assign n10599 = n10557 | n10598 ;
  assign n10600 = ~x588 & n10599 ;
  assign n10601 = ~n10474 & n10600 ;
  assign n10602 = n6153 | n10601 ;
  assign n10603 = n10408 | n10602 ;
  assign n10604 = n6412 | n10287 ;
  assign n10605 = x122 | n10604 ;
  assign n10606 = n5995 & n10605 ;
  assign n10607 = n1976 | n10296 ;
  assign n10608 = n10606 | n10607 ;
  assign n10609 = x87 | n10607 ;
  assign n10610 = n10314 | n10609 ;
  assign n10611 = x87 & ~n10607 ;
  assign n10612 = ~n10322 & n10611 ;
  assign n10613 = n10610 & ~n10612 ;
  assign n10614 = x122 & ~n10613 ;
  assign n10615 = n10608 & ~n10614 ;
  assign n10616 = x75 | n10615 ;
  assign n10617 = x567 & ~n5880 ;
  assign n10618 = n5882 & ~n10604 ;
  assign n10619 = n10617 & ~n10618 ;
  assign n10620 = n10616 & n10619 ;
  assign n10621 = n5880 & n10604 ;
  assign n10622 = n10288 | n10621 ;
  assign n10623 = n10620 | n10622 ;
  assign n10624 = ~x592 & n10623 ;
  assign n10625 = n10292 | n10624 ;
  assign n10626 = n6824 & ~n10625 ;
  assign n10627 = x443 & n10625 ;
  assign n10628 = n10339 | n10627 ;
  assign n10629 = n6903 | n10628 ;
  assign n10630 = ~x443 & n10625 ;
  assign n10631 = n10343 | n10630 ;
  assign n10632 = n6903 & ~n10631 ;
  assign n10633 = n10629 & ~n10632 ;
  assign n10634 = x435 & ~n10633 ;
  assign n10635 = ( x436 & x444 ) | ( x436 & n10628 ) | ( x444 & n10628 ) ;
  assign n10636 = ( ~x444 & n10631 ) | ( ~x444 & n10635 ) | ( n10631 & n10635 ) ;
  assign n10637 = ( ~x436 & n10635 ) | ( ~x436 & n10636 ) | ( n10635 & n10636 ) ;
  assign n10638 = x435 | n10637 ;
  assign n10639 = ~n10634 & n10638 ;
  assign n10640 = ( x429 & n6842 ) | ( x429 & ~n10639 ) | ( n6842 & ~n10639 ) ;
  assign n10641 = x435 | n10633 ;
  assign n10642 = x435 & ~n10637 ;
  assign n10643 = n10641 & ~n10642 ;
  assign n10644 = ( x429 & ~n6842 ) | ( x429 & n10643 ) | ( ~n6842 & n10643 ) ;
  assign n10645 = n10640 & ~n10644 ;
  assign n10646 = x1196 & ~n10645 ;
  assign n10647 = ( x429 & n6842 ) | ( x429 & n10639 ) | ( n6842 & n10639 ) ;
  assign n10648 = ( ~x429 & n6842 ) | ( ~x429 & n10643 ) | ( n6842 & n10643 ) ;
  assign n10649 = n10647 | n10648 ;
  assign n10650 = n10646 & n10649 ;
  assign n10651 = n10338 | n10650 ;
  assign n10652 = ~n10626 & n10651 ;
  assign n10653 = x428 | n10652 ;
  assign n10654 = x428 & ~n10625 ;
  assign n10655 = n10653 & ~n10654 ;
  assign n10656 = x427 | n10655 ;
  assign n10657 = x428 & ~n10652 ;
  assign n10658 = x428 | n10625 ;
  assign n10659 = ~n10657 & n10658 ;
  assign n10660 = x427 & ~n10659 ;
  assign n10661 = n10656 & ~n10660 ;
  assign n10662 = x430 & ~n10661 ;
  assign n10663 = x427 | n10659 ;
  assign n10664 = x427 & ~n10655 ;
  assign n10665 = n10663 & ~n10664 ;
  assign n10666 = x430 | n10665 ;
  assign n10667 = ~n10662 & n10666 ;
  assign n10668 = x426 & ~n10667 ;
  assign n10669 = x430 & ~n10665 ;
  assign n10670 = x430 | n10661 ;
  assign n10671 = ~n10669 & n10670 ;
  assign n10672 = x426 | n10671 ;
  assign n10673 = ~n10668 & n10672 ;
  assign n10674 = x445 & ~n10673 ;
  assign n10675 = x426 & ~n10671 ;
  assign n10676 = x426 | n10667 ;
  assign n10677 = ~n10675 & n10676 ;
  assign n10678 = x445 | n10677 ;
  assign n10679 = ~n10674 & n10678 ;
  assign n10680 = ( x448 & n6788 ) | ( x448 & ~n10679 ) | ( n6788 & ~n10679 ) ;
  assign n10681 = x445 & ~n10677 ;
  assign n10682 = x445 | n10673 ;
  assign n10683 = ~n10681 & n10682 ;
  assign n10684 = ( x448 & ~n6788 ) | ( x448 & n10683 ) | ( ~n6788 & n10683 ) ;
  assign n10685 = n10680 & ~n10684 ;
  assign n10686 = x1199 & ~n10685 ;
  assign n10687 = ( ~x448 & n6788 ) | ( ~x448 & n10683 ) | ( n6788 & n10683 ) ;
  assign n10688 = ( x448 & n6788 ) | ( x448 & n10679 ) | ( n6788 & n10679 ) ;
  assign n10689 = n10687 | n10688 ;
  assign n10690 = n10686 & n10689 ;
  assign n10691 = ~x1199 & n10652 ;
  assign n10692 = n6278 | n10691 ;
  assign n10693 = n10690 | n10692 ;
  assign n10694 = n10291 & n10693 ;
  assign n10695 = n6973 & ~n10625 ;
  assign n10696 = n10411 & ~n10695 ;
  assign n10697 = x1198 & ~n10696 ;
  assign n10698 = n6041 & ~n10625 ;
  assign n10699 = n10416 & ~n10698 ;
  assign n10700 = x355 | n10699 ;
  assign n10701 = x455 & n10289 ;
  assign n10702 = ~x455 & n10625 ;
  assign n10703 = n10701 | n10702 ;
  assign n10704 = ~x452 & n10703 ;
  assign n10705 = ~x455 & n10289 ;
  assign n10706 = x455 & n10625 ;
  assign n10707 = n10705 | n10706 ;
  assign n10708 = x452 & n10707 ;
  assign n10709 = n10704 | n10708 ;
  assign n10710 = x355 & ~n10709 ;
  assign n10711 = n10700 & ~n10710 ;
  assign n10712 = ( ~x458 & n6050 ) | ( ~x458 & n10711 ) | ( n6050 & n10711 ) ;
  assign n10713 = x355 & ~n10699 ;
  assign n10714 = x355 | n10709 ;
  assign n10715 = ~n10713 & n10714 ;
  assign n10716 = ( x458 & n6050 ) | ( x458 & n10715 ) | ( n6050 & n10715 ) ;
  assign n10717 = n10712 | n10716 ;
  assign n10718 = x1196 & n10717 ;
  assign n10719 = ( x458 & n6050 ) | ( x458 & ~n10715 ) | ( n6050 & ~n10715 ) ;
  assign n10720 = ( x458 & ~n6050 ) | ( x458 & n10711 ) | ( ~n6050 & n10711 ) ;
  assign n10721 = n10719 & ~n10720 ;
  assign n10722 = n10718 & ~n10721 ;
  assign n10723 = n10415 | n10722 ;
  assign n10724 = ~n10697 & n10723 ;
  assign n10725 = n6115 | n10724 ;
  assign n10726 = n6115 & ~n10625 ;
  assign n10727 = n10725 & ~n10726 ;
  assign n10728 = ~n6119 & n10727 ;
  assign n10729 = x1199 & n10625 ;
  assign n10730 = ~x351 & n10729 ;
  assign n10731 = n10728 | n10730 ;
  assign n10732 = ~x461 & n10731 ;
  assign n10733 = ~n6125 & n10727 ;
  assign n10734 = x351 & n10729 ;
  assign n10735 = n10733 | n10734 ;
  assign n10736 = x461 & n10735 ;
  assign n10737 = n10732 | n10736 ;
  assign n10738 = ~x357 & n10737 ;
  assign n10739 = ~x461 & n10735 ;
  assign n10740 = x461 & n10731 ;
  assign n10741 = n10739 | n10740 ;
  assign n10742 = x357 & n10741 ;
  assign n10743 = n10738 | n10742 ;
  assign n10744 = ~x356 & n10743 ;
  assign n10745 = ~x357 & n10741 ;
  assign n10746 = x357 & n10737 ;
  assign n10747 = n10745 | n10746 ;
  assign n10748 = x356 & n10747 ;
  assign n10749 = n10744 | n10748 ;
  assign n10750 = ( x354 & n5876 ) | ( x354 & n10749 ) | ( n5876 & n10749 ) ;
  assign n10751 = ~x356 & n10747 ;
  assign n10752 = x356 & n10743 ;
  assign n10753 = n10751 | n10752 ;
  assign n10754 = ( ~x354 & n5876 ) | ( ~x354 & n10753 ) | ( n5876 & n10753 ) ;
  assign n10755 = n10750 | n10754 ;
  assign n10756 = ~x591 & n10755 ;
  assign n10757 = ( x354 & n5876 ) | ( x354 & ~n10749 ) | ( n5876 & ~n10749 ) ;
  assign n10758 = ( x354 & ~n5876 ) | ( x354 & n10753 ) | ( ~n5876 & n10753 ) ;
  assign n10759 = n10757 & ~n10758 ;
  assign n10760 = n10756 & ~n10759 ;
  assign n10761 = n10410 & ~n10760 ;
  assign n10762 = x367 & n10289 ;
  assign n10763 = x592 & n10623 ;
  assign n10764 = n10559 | n10763 ;
  assign n10765 = ~x367 & n10764 ;
  assign n10766 = n10762 | n10765 ;
  assign n10767 = n6187 | n10766 ;
  assign n10768 = ~x367 & n10289 ;
  assign n10769 = x367 & n10764 ;
  assign n10770 = n10768 | n10769 ;
  assign n10771 = n6187 & ~n10770 ;
  assign n10772 = n10767 & ~n10771 ;
  assign n10773 = ( n6172 & n6178 ) | ( n6172 & n10772 ) | ( n6178 & n10772 ) ;
  assign n10774 = n6187 & n10766 ;
  assign n10775 = ~n6187 & n10770 ;
  assign n10776 = n10774 | n10775 ;
  assign n10777 = ( ~n6172 & n6178 ) | ( ~n6172 & n10776 ) | ( n6178 & n10776 ) ;
  assign n10778 = n10773 | n10777 ;
  assign n10779 = x1197 & n10778 ;
  assign n10780 = ( n6172 & n6178 ) | ( n6172 & ~n10772 ) | ( n6178 & ~n10772 ) ;
  assign n10781 = ( n6172 & ~n6178 ) | ( n6172 & n10776 ) | ( ~n6178 & n10776 ) ;
  assign n10782 = n10780 & ~n10781 ;
  assign n10783 = n10779 & ~n10782 ;
  assign n10784 = n10567 | n10783 ;
  assign n10785 = n6169 & ~n10764 ;
  assign n10786 = x1199 | n10785 ;
  assign n10787 = n10784 & ~n10786 ;
  assign n10788 = n7006 & ~n10764 ;
  assign n10789 = n10563 & ~n10788 ;
  assign n10790 = x1199 & n10789 ;
  assign n10791 = n10787 | n10790 ;
  assign n10792 = ~x374 & n10791 ;
  assign n10793 = n6233 & n10789 ;
  assign n10794 = ( x1198 & n10764 ) | ( x1198 & n10793 ) | ( n10764 & n10793 ) ;
  assign n10795 = ( ~x1198 & n10787 ) | ( ~x1198 & n10793 ) | ( n10787 & n10793 ) ;
  assign n10796 = n10794 | n10795 ;
  assign n10797 = x374 & n10796 ;
  assign n10798 = n10792 | n10797 ;
  assign n10799 = ( x369 & ~n10587 ) | ( x369 & n10798 ) | ( ~n10587 & n10798 ) ;
  assign n10800 = ~x374 & n10796 ;
  assign n10801 = x374 & n10791 ;
  assign n10802 = n10800 | n10801 ;
  assign n10803 = ( x369 & n10587 ) | ( x369 & ~n10802 ) | ( n10587 & ~n10802 ) ;
  assign n10804 = ~n10799 & n10803 ;
  assign n10805 = x591 | n10804 ;
  assign n10806 = ( x369 & n10587 ) | ( x369 & n10802 ) | ( n10587 & n10802 ) ;
  assign n10807 = ( ~x369 & n10587 ) | ( ~x369 & n10798 ) | ( n10587 & n10798 ) ;
  assign n10808 = n10806 | n10807 ;
  assign n10809 = ~n10805 & n10808 ;
  assign n10810 = n10475 & ~n10625 ;
  assign n10811 = ( x397 & ~x404 ) | ( x397 & x411 ) | ( ~x404 & x411 ) ;
  assign n10812 = ( ~x397 & x404 ) | ( ~x397 & n10811 ) | ( x404 & n10811 ) ;
  assign n10813 = ( ~x411 & n10811 ) | ( ~x411 & n10812 ) | ( n10811 & n10812 ) ;
  assign n10814 = n6302 & n10813 ;
  assign n10815 = n6302 | n10813 ;
  assign n10816 = ~n10814 & n10815 ;
  assign n10817 = n5950 & ~n10816 ;
  assign n10818 = n10286 | n10817 ;
  assign n10819 = ( x412 & n6299 ) | ( x412 & ~n10818 ) | ( n6299 & ~n10818 ) ;
  assign n10820 = n5950 & n10816 ;
  assign n10821 = n10286 | n10820 ;
  assign n10822 = ( x412 & ~n6299 ) | ( x412 & n10821 ) | ( ~n6299 & n10821 ) ;
  assign n10823 = n10819 & ~n10822 ;
  assign n10824 = x122 | n10823 ;
  assign n10825 = ( x412 & n6299 ) | ( x412 & n10818 ) | ( n6299 & n10818 ) ;
  assign n10826 = ( ~x412 & n6299 ) | ( ~x412 & n10821 ) | ( n6299 & n10821 ) ;
  assign n10827 = n10825 | n10826 ;
  assign n10828 = ~n10824 & n10827 ;
  assign n10829 = n10286 | n10828 ;
  assign n10830 = n5995 & n10829 ;
  assign n10831 = n10296 | n10830 ;
  assign n10832 = x567 & n10831 ;
  assign n10833 = ~x122 & n5950 ;
  assign n10834 = n10286 | n10833 ;
  assign n10835 = n5950 & n6341 ;
  assign n10836 = x122 | n10286 ;
  assign n10837 = n10835 | n10836 ;
  assign n10838 = n10316 & n10837 ;
  assign n10839 = n10834 & n10838 ;
  assign n10840 = x567 & n10839 ;
  assign n10841 = n10288 | n10840 ;
  assign n10842 = n10832 | n10841 ;
  assign n10843 = n10294 & n10842 ;
  assign n10844 = n1976 | n10838 ;
  assign n10845 = n10830 | n10844 ;
  assign n10846 = n10507 | n10609 ;
  assign n10847 = n6308 & ~n10484 ;
  assign n10848 = n10481 & ~n10847 ;
  assign n10849 = n10846 | n10848 ;
  assign n10850 = ~n10512 & n10611 ;
  assign n10851 = ~n10491 & n10850 ;
  assign n10852 = n10849 & ~n10851 ;
  assign n10853 = ~x122 & n10835 ;
  assign n10854 = n10828 | n10853 ;
  assign n10855 = n10852 | n10854 ;
  assign n10856 = n10845 & n10855 ;
  assign n10857 = x75 | n10856 ;
  assign n10858 = n5882 & ~n10839 ;
  assign n10859 = ~n10830 & n10858 ;
  assign n10860 = n10617 & ~n10859 ;
  assign n10861 = n10857 & n10860 ;
  assign n10862 = n10843 | n10861 ;
  assign n10863 = n6678 & n10862 ;
  assign n10864 = n10294 & n10841 ;
  assign n10865 = ~n10513 & n10611 ;
  assign n10866 = n10846 & ~n10865 ;
  assign n10867 = x122 & ~n10866 ;
  assign n10868 = n10844 & ~n10867 ;
  assign n10869 = x75 | n10868 ;
  assign n10870 = n10617 & ~n10858 ;
  assign n10871 = n10869 & n10870 ;
  assign n10872 = n10864 | n10871 ;
  assign n10873 = ~n6686 & n10872 ;
  assign n10874 = n10863 | n10873 ;
  assign n10875 = ( x1199 & n10292 ) | ( x1199 & n10874 ) | ( n10292 & n10874 ) ;
  assign n10876 = n10288 | n10832 ;
  assign n10877 = n10294 & n10876 ;
  assign n10878 = ( ~x75 & n10617 ) | ( ~x75 & n10831 ) | ( n10617 & n10831 ) ;
  assign n10879 = x122 & n10486 ;
  assign n10880 = n10828 | n10879 ;
  assign n10881 = n5995 & n10880 ;
  assign n10882 = n10609 | n10881 ;
  assign n10883 = x122 & n10491 ;
  assign n10884 = n10828 | n10883 ;
  assign n10885 = n5995 & n10884 ;
  assign n10886 = n10611 & ~n10885 ;
  assign n10887 = n1976 & ~n10831 ;
  assign n10888 = n10886 | n10887 ;
  assign n10889 = n10882 & ~n10888 ;
  assign n10890 = ( x75 & n10617 ) | ( x75 & n10889 ) | ( n10617 & n10889 ) ;
  assign n10891 = n10878 & n10890 ;
  assign n10892 = n10877 | n10891 ;
  assign n10893 = n6678 & n10892 ;
  assign n10894 = n10337 | n10893 ;
  assign n10895 = ( ~x1199 & n10292 ) | ( ~x1199 & n10894 ) | ( n10292 & n10894 ) ;
  assign n10896 = n10875 | n10895 ;
  assign n10897 = n10475 | n10896 ;
  assign n10898 = ~n10810 & n10897 ;
  assign n10899 = x333 & ~n10898 ;
  assign n10900 = n6295 & n10625 ;
  assign n10901 = ~n6295 & n10896 ;
  assign n10902 = n10900 | n10901 ;
  assign n10903 = x333 | n10902 ;
  assign n10904 = ~n10899 & n10903 ;
  assign n10905 = x391 & ~n10904 ;
  assign n10906 = x333 & n10902 ;
  assign n10907 = ~x333 & n10898 ;
  assign n10908 = n10906 | n10907 ;
  assign n10909 = x391 | n10908 ;
  assign n10910 = ~n10905 & n10909 ;
  assign n10911 = x392 | n10910 ;
  assign n10912 = ~x391 & n10904 ;
  assign n10913 = x391 & n10908 ;
  assign n10914 = n10912 | n10913 ;
  assign n10915 = x392 & ~n10914 ;
  assign n10916 = n10911 & ~n10915 ;
  assign n10917 = ( x393 & n6588 ) | ( x393 & n10916 ) | ( n6588 & n10916 ) ;
  assign n10918 = x392 & ~n10910 ;
  assign n10919 = x392 | n10914 ;
  assign n10920 = ~n10918 & n10919 ;
  assign n10921 = ( ~x393 & n6588 ) | ( ~x393 & n10920 ) | ( n6588 & n10920 ) ;
  assign n10922 = n10917 | n10921 ;
  assign n10923 = ( x393 & n6588 ) | ( x393 & ~n10916 ) | ( n6588 & ~n10916 ) ;
  assign n10924 = ( x393 & ~n6588 ) | ( x393 & n10920 ) | ( ~n6588 & n10920 ) ;
  assign n10925 = n10923 & ~n10924 ;
  assign n10926 = n10922 & ~n10925 ;
  assign n10927 = ( x590 & n6278 ) | ( x590 & n10926 ) | ( n6278 & n10926 ) ;
  assign n10928 = n10809 | n10927 ;
  assign n10929 = ~x588 & n10928 ;
  assign n10930 = ~n10761 & n10929 ;
  assign n10931 = n6153 & ~n10930 ;
  assign n10932 = ~n10694 & n10931 ;
  assign n10933 = x80 | n6785 ;
  assign n10934 = n10932 | n10933 ;
  assign n10935 = n10603 & ~n10934 ;
  assign n10936 = x392 & ~n6591 ;
  assign n10937 = ~x392 & n6591 ;
  assign n10938 = n10936 | n10937 ;
  assign n10939 = n6969 | n10289 ;
  assign n10940 = n10475 & n10939 ;
  assign n10941 = n6678 & n10842 ;
  assign n10942 = ~n6686 & n10841 ;
  assign n10943 = n10292 | n10942 ;
  assign n10944 = n10941 | n10943 ;
  assign n10945 = x1199 & n10944 ;
  assign n10946 = n6678 & n10876 ;
  assign n10947 = n10502 | n10946 ;
  assign n10948 = ( ~x1199 & n10945 ) | ( ~x1199 & n10947 ) | ( n10945 & n10947 ) ;
  assign n10949 = ~n10475 & n10948 ;
  assign n10950 = n10940 | n10949 ;
  assign n10951 = ~x333 & n10950 ;
  assign n10952 = n6295 & n10939 ;
  assign n10953 = ~n6295 & n10948 ;
  assign n10954 = n10952 | n10953 ;
  assign n10955 = x333 & n10954 ;
  assign n10956 = n10951 | n10955 ;
  assign n10957 = ( x391 & n10938 ) | ( x391 & ~n10956 ) | ( n10938 & ~n10956 ) ;
  assign n10958 = x333 & n10950 ;
  assign n10959 = ~x333 & n10954 ;
  assign n10960 = n10958 | n10959 ;
  assign n10961 = ( x391 & ~n10938 ) | ( x391 & n10960 ) | ( ~n10938 & n10960 ) ;
  assign n10962 = n10957 & ~n10961 ;
  assign n10963 = x591 & ~n10962 ;
  assign n10964 = ( x391 & n10938 ) | ( x391 & n10956 ) | ( n10938 & n10956 ) ;
  assign n10965 = ( ~x391 & n10938 ) | ( ~x391 & n10960 ) | ( n10938 & n10960 ) ;
  assign n10966 = n10964 | n10965 ;
  assign n10967 = n10963 & n10966 ;
  assign n10968 = ~n6969 & n7022 ;
  assign n10969 = n6473 & n7009 ;
  assign n10970 = x1198 | n10969 ;
  assign n10971 = ~n7036 & n10970 ;
  assign n10972 = ~n10968 & n10971 ;
  assign n10973 = n10289 | n10972 ;
  assign n10974 = ~x591 & n10973 ;
  assign n10975 = x590 | n10974 ;
  assign n10976 = n10967 | n10975 ;
  assign n10977 = n6980 | n10289 ;
  assign n10978 = n6976 | n10977 ;
  assign n10979 = n6125 | n10978 ;
  assign n10980 = n10939 & n10979 ;
  assign n10981 = x461 & ~n10980 ;
  assign n10982 = n6119 | n10978 ;
  assign n10983 = n10939 & n10982 ;
  assign n10984 = x461 | n10983 ;
  assign n10985 = ~n10981 & n10984 ;
  assign n10986 = x357 & ~n10985 ;
  assign n10987 = x461 & ~n10983 ;
  assign n10988 = x461 | n10980 ;
  assign n10989 = ~n10987 & n10988 ;
  assign n10990 = x357 | n10989 ;
  assign n10991 = ~n10986 & n10990 ;
  assign n10992 = x356 & ~n10991 ;
  assign n10993 = x357 & ~n10989 ;
  assign n10994 = x357 | n10985 ;
  assign n10995 = ~n10993 & n10994 ;
  assign n10996 = x356 | n10995 ;
  assign n10997 = ~n10992 & n10996 ;
  assign n10998 = ( x354 & n5876 ) | ( x354 & n10997 ) | ( n5876 & n10997 ) ;
  assign n10999 = x356 & ~n10995 ;
  assign n11000 = x356 | n10991 ;
  assign n11001 = ~n10999 & n11000 ;
  assign n11002 = ( ~x354 & n5876 ) | ( ~x354 & n11001 ) | ( n5876 & n11001 ) ;
  assign n11003 = n10998 | n11002 ;
  assign n11004 = ~x591 & n11003 ;
  assign n11005 = ( x354 & ~n5876 ) | ( x354 & n11001 ) | ( ~n5876 & n11001 ) ;
  assign n11006 = ( x354 & n5876 ) | ( x354 & ~n10997 ) | ( n5876 & ~n10997 ) ;
  assign n11007 = ~n11005 & n11006 ;
  assign n11008 = n11004 & ~n11007 ;
  assign n11009 = n10410 & ~n11008 ;
  assign n11010 = x588 | n11009 ;
  assign n11011 = n10976 & ~n11010 ;
  assign n11012 = x592 & n6824 ;
  assign n11013 = n6473 & n7070 ;
  assign n11014 = ~n11012 & n11013 ;
  assign n11015 = n10289 | n11014 ;
  assign n11016 = x428 & n11015 ;
  assign n11017 = ~x428 & n10939 ;
  assign n11018 = n11016 | n11017 ;
  assign n11019 = ~x427 & n11018 ;
  assign n11020 = ~x428 & n11015 ;
  assign n11021 = x428 & n10939 ;
  assign n11022 = n11020 | n11021 ;
  assign n11023 = x427 & n11022 ;
  assign n11024 = n11019 | n11023 ;
  assign n11025 = ~x430 & n11024 ;
  assign n11026 = ~x427 & n11022 ;
  assign n11027 = x427 & n11018 ;
  assign n11028 = n11026 | n11027 ;
  assign n11029 = x430 & n11028 ;
  assign n11030 = n11025 | n11029 ;
  assign n11031 = ~x426 & n11030 ;
  assign n11032 = ~x430 & n11028 ;
  assign n11033 = x430 & n11024 ;
  assign n11034 = n11032 | n11033 ;
  assign n11035 = x426 & n11034 ;
  assign n11036 = n11031 | n11035 ;
  assign n11037 = ~x445 & n11036 ;
  assign n11038 = ~x426 & n11034 ;
  assign n11039 = x426 & n11030 ;
  assign n11040 = n11038 | n11039 ;
  assign n11041 = x445 & n11040 ;
  assign n11042 = n11037 | n11041 ;
  assign n11043 = ( x448 & n6788 ) | ( x448 & n11042 ) | ( n6788 & n11042 ) ;
  assign n11044 = ~x445 & n11040 ;
  assign n11045 = x445 & n11036 ;
  assign n11046 = n11044 | n11045 ;
  assign n11047 = ( ~x448 & n6788 ) | ( ~x448 & n11046 ) | ( n6788 & n11046 ) ;
  assign n11048 = n11043 | n11047 ;
  assign n11049 = x1199 & n11048 ;
  assign n11050 = ( x448 & n6788 ) | ( x448 & ~n11042 ) | ( n6788 & ~n11042 ) ;
  assign n11051 = ( x448 & ~n6788 ) | ( x448 & n11046 ) | ( ~n6788 & n11046 ) ;
  assign n11052 = n11050 & ~n11051 ;
  assign n11053 = n11049 & ~n11052 ;
  assign n11054 = ~x1199 & n11015 ;
  assign n11055 = n6278 | n11054 ;
  assign n11056 = n11053 | n11055 ;
  assign n11057 = n10291 & n11056 ;
  assign n11058 = n6153 & ~n11057 ;
  assign n11059 = ~n11011 & n11058 ;
  assign n11060 = n6153 | n10289 ;
  assign n11061 = ~x80 & n6785 ;
  assign n11062 = n11060 & n11061 ;
  assign n11063 = ~n11059 & n11062 ;
  assign n11064 = x217 | n11063 ;
  assign n11065 = n10935 | n11064 ;
  assign n11066 = ~x80 & n10289 ;
  assign n11067 = x217 & ~n11066 ;
  assign n11068 = n7103 | n11067 ;
  assign n11069 = n11065 & ~n11068 ;
  assign n11070 = n6785 | n9443 ;
  assign n11071 = x81 & ~x314 ;
  assign n11072 = ~n1242 & n11071 ;
  assign n11073 = x68 & ~x81 ;
  assign n11074 = ~n1228 & n11073 ;
  assign n11075 = ~n9170 & n11074 ;
  assign n11076 = ~n9575 & n11075 ;
  assign n11077 = ~n1386 & n11076 ;
  assign n11078 = n11072 | n11077 ;
  assign n11079 = ~n11070 & n11078 ;
  assign n11080 = x69 & x314 ;
  assign n11081 = ~n1356 & n11080 ;
  assign n11082 = n1228 | n1230 ;
  assign n11083 = n1226 | n11082 ;
  assign n11084 = x66 & ~x73 ;
  assign n11085 = ~n1234 & n11084 ;
  assign n11086 = ~n11083 & n11085 ;
  assign n11087 = n11081 | n11086 ;
  assign n11088 = n9260 | n9262 ;
  assign n11089 = n11087 & ~n11088 ;
  assign n11090 = n1218 | n9261 ;
  assign n11091 = n1253 | n11090 ;
  assign n11092 = n1228 | n1364 ;
  assign n11093 = x84 & ~n7353 ;
  assign n11094 = ~n11092 & n11093 ;
  assign n11095 = ~n1233 & n11094 ;
  assign n11096 = ~n11091 & n11095 ;
  assign n11097 = ( x314 & n8332 ) | ( x314 & ~n11096 ) | ( n8332 & ~n11096 ) ;
  assign n11098 = x83 | n11094 ;
  assign n11099 = ~n11091 & n11098 ;
  assign n11100 = ~n1360 & n11099 ;
  assign n11101 = ( x314 & ~n8332 ) | ( x314 & n11100 ) | ( ~n8332 & n11100 ) ;
  assign n11102 = ~n11097 & n11101 ;
  assign n11103 = x211 & x299 ;
  assign n11104 = x219 & x299 ;
  assign n11105 = n11103 | n11104 ;
  assign n11106 = n8981 | n11105 ;
  assign n11107 = n6785 | n11106 ;
  assign n11108 = n9521 & ~n11107 ;
  assign n11109 = n4849 & ~n9263 ;
  assign n11110 = x314 | n9264 ;
  assign n11111 = n9573 & ~n11110 ;
  assign n11112 = n11109 | n11111 ;
  assign n11113 = ~n9260 & n11112 ;
  assign n11114 = n5943 & n9531 ;
  assign n11115 = n5939 & n9534 ;
  assign n11116 = n11114 | n11115 ;
  assign n11117 = n9139 & n11116 ;
  assign n11118 = n1406 & ~n11090 ;
  assign n11119 = x314 & ~n8332 ;
  assign n11120 = ~n1253 & n11119 ;
  assign n11121 = n11118 & n11120 ;
  assign n11122 = ~n1259 & n5950 ;
  assign n11123 = x1093 | n1864 ;
  assign n11124 = n2033 | n11123 ;
  assign n11125 = n11122 & ~n11124 ;
  assign n11126 = n9594 & n11125 ;
  assign n11127 = ~n9598 & n11126 ;
  assign n11128 = ( n6153 & n6785 ) | ( n6153 & ~n11127 ) | ( n6785 & ~n11127 ) ;
  assign n11129 = n5891 | n10300 ;
  assign n11130 = n9186 & ~n11129 ;
  assign n11131 = n9201 & ~n10297 ;
  assign n11132 = n11130 & n11131 ;
  assign n11133 = n2033 | n8243 ;
  assign n11134 = ( x1093 & ~n11132 ) | ( x1093 & n11133 ) | ( ~n11132 & n11133 ) ;
  assign n11135 = n5950 & n9189 ;
  assign n11136 = ( x1093 & ~n11133 ) | ( x1093 & n11135 ) | ( ~n11133 & n11135 ) ;
  assign n11137 = ~n11134 & n11136 ;
  assign n11138 = ( n6153 & ~n6785 ) | ( n6153 & n11137 ) | ( ~n6785 & n11137 ) ;
  assign n11139 = ~n11128 & n11138 ;
  assign n11140 = x70 & n7189 ;
  assign n11141 = n1865 | n8331 ;
  assign n11142 = x70 | x841 ;
  assign n11143 = n7148 | n8353 ;
  assign n11144 = n7170 | n11143 ;
  assign n11145 = n8350 & ~n11144 ;
  assign n11146 = ~n5899 & n11145 ;
  assign n11147 = ( x70 & n11142 ) | ( x70 & n11146 ) | ( n11142 & n11146 ) ;
  assign n11148 = ~n11141 & n11147 ;
  assign n11149 = ~n11140 & n11148 ;
  assign n11150 = ~x1050 & n7786 ;
  assign n11151 = x90 | n11150 ;
  assign n11152 = ~n9468 & n11151 ;
  assign n11153 = ~n1309 & n11152 ;
  assign n11154 = ~n5887 & n11153 ;
  assign n11155 = ~x58 & n1314 ;
  assign n11156 = n8324 | n11155 ;
  assign n11157 = n1292 & ~n8328 ;
  assign n11158 = n11156 & n11157 ;
  assign n11159 = x24 & ~n1527 ;
  assign n11160 = ~n1292 & n11159 ;
  assign n11161 = ~n9243 & n11160 ;
  assign n11162 = n1314 & n11161 ;
  assign n11163 = x39 | n11162 ;
  assign n11164 = n11158 | n11163 ;
  assign n11165 = ~n8359 & n11164 ;
  assign n11166 = ~n5947 & n11165 ;
  assign n11167 = x92 & ~n1868 ;
  assign n11168 = ~n2111 & n9609 ;
  assign n11169 = n11167 & n11168 ;
  assign n11170 = n4343 & n4732 ;
  assign n11171 = n5943 & n11170 ;
  assign n11172 = ~n2213 & n4767 ;
  assign n11173 = n5939 & n11172 ;
  assign n11174 = n11171 | n11173 ;
  assign n11175 = ~n2042 & n9306 ;
  assign n11176 = n11174 & n11175 ;
  assign n11177 = n11169 | n11176 ;
  assign n11178 = ~n8329 & n11177 ;
  assign n11179 = x93 & ~n9243 ;
  assign n11180 = n1603 & n11179 ;
  assign n11181 = ( x92 & ~n8330 ) | ( x92 & n11180 ) | ( ~n8330 & n11180 ) ;
  assign n11182 = x1050 | n1868 ;
  assign n11183 = ( x92 & n8330 ) | ( x92 & n11182 ) | ( n8330 & n11182 ) ;
  assign n11184 = n11181 & ~n11183 ;
  assign n11185 = n9226 & ~n9428 ;
  assign n11186 = ( n7119 & ~n8331 ) | ( n7119 & n11185 ) | ( ~n8331 & n11185 ) ;
  assign n11187 = ( x1093 & n4741 ) | ( x1093 & ~n11185 ) | ( n4741 & ~n11185 ) ;
  assign n11188 = n1693 & ~n11187 ;
  assign n11189 = ~n8419 & n9224 ;
  assign n11190 = n1344 | n11189 ;
  assign n11191 = n1590 | n8328 ;
  assign n11192 = x252 & ~n11191 ;
  assign n11193 = n11190 & n11192 ;
  assign n11194 = n11188 | n11193 ;
  assign n11195 = n7136 & ~n11185 ;
  assign n11196 = ~x252 & n11185 ;
  assign n11197 = ( n11194 & ~n11195 ) | ( n11194 & n11196 ) | ( ~n11195 & n11196 ) ;
  assign n11198 = ( n7119 & n8331 ) | ( n7119 & ~n11197 ) | ( n8331 & ~n11197 ) ;
  assign n11199 = n11186 & ~n11198 ;
  assign n11200 = n4766 & n4997 ;
  assign n11201 = n2214 | n9554 ;
  assign n11202 = n11200 & ~n11201 ;
  assign n11203 = ~n9557 & n9560 ;
  assign n11204 = n4997 & n11203 ;
  assign n11205 = x39 & ~n11204 ;
  assign n11206 = ~n11202 & n11205 ;
  assign n11207 = ~n1212 & n9858 ;
  assign n11208 = n9592 & n11207 ;
  assign n11209 = x332 | n8328 ;
  assign n11210 = n9427 | n11209 ;
  assign n11211 = n11145 & ~n11210 ;
  assign n11212 = x39 | n11211 ;
  assign n11213 = n11208 | n11212 ;
  assign n11214 = ~n8366 & n11213 ;
  assign n11215 = ~n11206 & n11214 ;
  assign n11216 = ~n8498 & n11207 ;
  assign n11217 = x479 & ~n7136 ;
  assign n11218 = n1533 & n11217 ;
  assign n11219 = x96 & ~n1492 ;
  assign n11220 = ~n1525 & n11219 ;
  assign n11221 = ~n11217 & n11220 ;
  assign n11222 = n1605 & n11221 ;
  assign n11223 = n11218 | n11222 ;
  assign n11224 = ~x95 & n11223 ;
  assign n11225 = n11216 | n11224 ;
  assign n11226 = ~n8331 & n11225 ;
  assign n11227 = x39 & x593 ;
  assign n11228 = n9562 & n11227 ;
  assign n11229 = n4997 & n11228 ;
  assign n11230 = n4694 & n11217 ;
  assign n11231 = n4800 | n11230 ;
  assign n11232 = x96 | n8361 ;
  assign n11233 = n11231 & ~n11232 ;
  assign n11234 = n9621 & n11233 ;
  assign n11235 = n11229 | n11234 ;
  assign n11236 = ~n8366 & n11235 ;
  assign n11237 = ~x92 & n9610 ;
  assign n11238 = n11167 | n11237 ;
  assign n11239 = x314 & x1050 ;
  assign n11240 = ~n8330 & n11239 ;
  assign n11241 = n11238 & n11240 ;
  assign n11242 = ~x72 & x152 ;
  assign n11243 = n8467 & n11242 ;
  assign n11244 = x299 & n11243 ;
  assign n11245 = ~x72 & x174 ;
  assign n11246 = ~x299 & n11245 ;
  assign n11247 = n8478 & n11246 ;
  assign n11248 = n11244 | n11247 ;
  assign n11249 = x232 & n11248 ;
  assign n11250 = x39 & ~n11249 ;
  assign n11251 = ~x72 & x99 ;
  assign n11252 = x39 | n11251 ;
  assign n11253 = ~n11250 & n11252 ;
  assign n11254 = ( n5880 & n6785 ) | ( n5880 & ~n11253 ) | ( n6785 & ~n11253 ) ;
  assign n11255 = n6417 | n11251 ;
  assign n11256 = ~n8503 & n11251 ;
  assign n11257 = ~n4787 & n9125 ;
  assign n11258 = n11256 | n11257 ;
  assign n11259 = n8623 & n11258 ;
  assign n11260 = ( n6417 & n8507 ) | ( n6417 & ~n11251 ) | ( n8507 & ~n11251 ) ;
  assign n11261 = ~n11259 & n11260 ;
  assign n11262 = n11255 & ~n11261 ;
  assign n11263 = x39 | n11262 ;
  assign n11264 = n2007 | n11250 ;
  assign n11265 = n11263 & ~n11264 ;
  assign n11266 = n2007 & n11253 ;
  assign n11267 = x75 & ~n11266 ;
  assign n11268 = ~n11265 & n11267 ;
  assign n11269 = x41 & x72 ;
  assign n11270 = x99 & ~n11269 ;
  assign n11271 = ~n8550 & n11270 ;
  assign n11272 = n8915 & ~n11271 ;
  assign n11273 = ~n8557 & n11270 ;
  assign n11274 = n8914 | n11273 ;
  assign n11275 = ~n11272 & n11274 ;
  assign n11276 = x228 & ~n11275 ;
  assign n11277 = ~n8604 & n11270 ;
  assign n11278 = n8701 | n11277 ;
  assign n11279 = ( ~x39 & n8693 ) | ( ~x39 & n11278 ) | ( n8693 & n11278 ) ;
  assign n11280 = ~n11276 & n11279 ;
  assign n11281 = n8469 & n11248 ;
  assign n11282 = ~n9092 & n11281 ;
  assign n11283 = n1975 | n11282 ;
  assign n11284 = n11280 | n11283 ;
  assign n11285 = ~n8620 & n11251 ;
  assign n11286 = ~n4786 & n8490 ;
  assign n11287 = n11285 | n11286 ;
  assign n11288 = n8623 & n11287 ;
  assign n11289 = n11260 & ~n11288 ;
  assign n11290 = n11255 & ~n11289 ;
  assign n11291 = x39 | n11290 ;
  assign n11292 = ~n11250 & n11291 ;
  assign n11293 = n4807 & ~n11292 ;
  assign n11294 = x38 & ~n11253 ;
  assign n11295 = x87 | n11294 ;
  assign n11296 = n11293 | n11295 ;
  assign n11297 = n11284 & ~n11296 ;
  assign n11298 = x228 & ~n8726 ;
  assign n11299 = x228 & ~n8617 ;
  assign n11300 = n11251 & ~n11299 ;
  assign n11301 = n2041 | n11300 ;
  assign n11302 = n11298 | n11301 ;
  assign n11303 = n2041 & ~n11253 ;
  assign n11304 = n11302 & ~n11303 ;
  assign n11305 = ( x75 & n1998 ) | ( x75 & n11304 ) | ( n1998 & n11304 ) ;
  assign n11306 = n11297 | n11305 ;
  assign n11307 = ~n11268 & n11306 ;
  assign n11308 = ( n5880 & ~n6785 ) | ( n5880 & n11307 ) | ( ~n6785 & n11307 ) ;
  assign n11309 = ~n11254 & n11308 ;
  assign n11310 = n6785 & n11252 ;
  assign n11311 = n8469 & n11243 ;
  assign n11312 = ( ~x39 & n11310 ) | ( ~x39 & n11311 ) | ( n11310 & n11311 ) ;
  assign n11313 = n11309 | n11312 ;
  assign n11314 = x129 & ~n8248 ;
  assign n11315 = n5923 | n11314 ;
  assign n11316 = n4784 & n4803 ;
  assign n11317 = x129 & ~n8247 ;
  assign n11318 = n8251 & ~n11317 ;
  assign n11319 = n11316 | n11318 ;
  assign n11320 = n11315 & ~n11319 ;
  assign n11321 = x75 | n1983 ;
  assign n11322 = n4807 & ~n11321 ;
  assign n11323 = ~n11320 & n11322 ;
  assign n11324 = ~x24 & n7197 ;
  assign n11325 = n7136 & n11324 ;
  assign n11326 = ~n7194 & n11325 ;
  assign n11327 = n11323 | n11326 ;
  assign n11328 = ~n7113 & n11327 ;
  assign n11329 = ~n1868 & n11328 ;
  assign n11330 = x152 & ~n2157 ;
  assign n11331 = ~n4713 & n11330 ;
  assign n11332 = ~x72 & n11331 ;
  assign n11333 = ( x232 & ~x299 ) | ( x232 & n11332 ) | ( ~x299 & n11332 ) ;
  assign n11334 = ~x144 & x174 ;
  assign n11335 = ~n8477 & n11334 ;
  assign n11336 = ~x72 & n11335 ;
  assign n11337 = ( x232 & x299 ) | ( x232 & n11336 ) | ( x299 & n11336 ) ;
  assign n11338 = n11333 & n11337 ;
  assign n11339 = x39 & ~n11338 ;
  assign n11340 = x39 | n8496 ;
  assign n11341 = ~n11339 & n11340 ;
  assign n11342 = ( n5880 & n6785 ) | ( n5880 & ~n11341 ) | ( n6785 & ~n11341 ) ;
  assign n11343 = n6417 | n8496 ;
  assign n11344 = n1288 & n4794 ;
  assign n11345 = n8496 & ~n8502 ;
  assign n11346 = n8491 | n11345 ;
  assign n11347 = n11344 & n11346 ;
  assign n11348 = ( n6417 & ~n8496 ) | ( n6417 & n8507 ) | ( ~n8496 & n8507 ) ;
  assign n11349 = ~n11347 & n11348 ;
  assign n11350 = n11343 & ~n11349 ;
  assign n11351 = x39 | n11350 ;
  assign n11352 = n2007 | n11339 ;
  assign n11353 = n11351 & ~n11352 ;
  assign n11354 = n2007 & n11341 ;
  assign n11355 = x75 & ~n11354 ;
  assign n11356 = ~n11353 & n11355 ;
  assign n11357 = x101 & ~n8548 ;
  assign n11358 = n1288 & ~n8537 ;
  assign n11359 = ~n11357 & n11358 ;
  assign n11360 = x101 & ~n8555 ;
  assign n11361 = n1288 | n8561 ;
  assign n11362 = n11360 | n11361 ;
  assign n11363 = ~n11359 & n11362 ;
  assign n11364 = x228 & ~n11363 ;
  assign n11365 = x101 & ~n8602 ;
  assign n11366 = n8595 | n11365 ;
  assign n11367 = ( ~x39 & n8693 ) | ( ~x39 & n11366 ) | ( n8693 & n11366 ) ;
  assign n11368 = ~n11364 & n11367 ;
  assign n11369 = ~n9093 & n11331 ;
  assign n11370 = ( ~x299 & n8469 ) | ( ~x299 & n11369 ) | ( n8469 & n11369 ) ;
  assign n11371 = ~n9093 & n11335 ;
  assign n11372 = ( x299 & n8469 ) | ( x299 & n11371 ) | ( n8469 & n11371 ) ;
  assign n11373 = n11370 & n11372 ;
  assign n11374 = n1975 | n11373 ;
  assign n11375 = n11368 | n11374 ;
  assign n11376 = ~x44 & n9101 ;
  assign n11377 = n8496 & ~n11376 ;
  assign n11378 = n8490 | n11377 ;
  assign n11379 = n11344 & n11378 ;
  assign n11380 = n11348 & ~n11379 ;
  assign n11381 = n11343 & ~n11380 ;
  assign n11382 = x39 | n11381 ;
  assign n11383 = ~n11339 & n11382 ;
  assign n11384 = n4807 & ~n11383 ;
  assign n11385 = x38 & ~n11341 ;
  assign n11386 = x87 | n11385 ;
  assign n11387 = n11384 | n11386 ;
  assign n11388 = n11375 & ~n11387 ;
  assign n11389 = ~x101 & n9116 ;
  assign n11390 = ~n8616 & n9115 ;
  assign n11391 = n8496 & ~n11390 ;
  assign n11392 = x39 | n11391 ;
  assign n11393 = n11389 | n11392 ;
  assign n11394 = ~n11339 & n11393 ;
  assign n11395 = ( x75 & n1998 ) | ( x75 & n11394 ) | ( n1998 & n11394 ) ;
  assign n11396 = n11388 | n11395 ;
  assign n11397 = ~n11356 & n11396 ;
  assign n11398 = ( n5880 & ~n6785 ) | ( n5880 & n11397 ) | ( ~n6785 & n11397 ) ;
  assign n11399 = ~n11342 & n11398 ;
  assign n11400 = n6785 & n11340 ;
  assign n11401 = n8469 & n11332 ;
  assign n11402 = ( ~x39 & n11400 ) | ( ~x39 & n11401 ) | ( n11400 & n11401 ) ;
  assign n11403 = n11399 | n11402 ;
  assign n11404 = n1412 & ~n7149 ;
  assign n11405 = ~n11070 & n11404 ;
  assign n11406 = x109 & ~n1325 ;
  assign n11407 = ~n1249 & n11406 ;
  assign n11408 = ( x314 & n9259 ) | ( x314 & ~n11407 ) | ( n9259 & ~n11407 ) ;
  assign n11409 = x109 | n11118 ;
  assign n11410 = ~n1454 & n11409 ;
  assign n11411 = ( x314 & ~n9259 ) | ( x314 & n11410 ) | ( ~n9259 & n11410 ) ;
  assign n11412 = ~n11408 & n11411 ;
  assign n11413 = n7119 & n8244 ;
  assign n11414 = ( n6153 & n8244 ) | ( n6153 & n11413 ) | ( n8244 & n11413 ) ;
  assign n11415 = n8590 & ~n11414 ;
  assign n11416 = x110 | n11130 ;
  assign n11417 = ~x47 & n9201 ;
  assign n11418 = n11416 & n11417 ;
  assign n11419 = ~n8569 & n11418 ;
  assign n11420 = n5925 & ~n8243 ;
  assign n11421 = n11419 & n11420 ;
  assign n11422 = n5925 | n8243 ;
  assign n11423 = ( n4795 & ~n11132 ) | ( n4795 & n11422 ) | ( ~n11132 & n11422 ) ;
  assign n11424 = ( n4795 & n11419 ) | ( n4795 & ~n11422 ) | ( n11419 & ~n11422 ) ;
  assign n11425 = ~n11423 & n11424 ;
  assign n11426 = n11421 | n11425 ;
  assign n11427 = n6153 & n11426 ;
  assign n11428 = n11415 | n11427 ;
  assign n11429 = ~n8331 & n11428 ;
  assign n11430 = x24 & n9426 ;
  assign n11431 = x53 | n9425 ;
  assign n11432 = ~n1585 & n11431 ;
  assign n11433 = x24 | n1590 ;
  assign n11434 = n11432 & ~n11433 ;
  assign n11435 = n11430 | n11434 ;
  assign n11436 = x841 & n11435 ;
  assign n11437 = ~n7176 & n9411 ;
  assign n11438 = n11436 | n11437 ;
  assign n11439 = ~n8332 & n11438 ;
  assign n11440 = x999 | n8332 ;
  assign n11441 = n9491 & ~n11440 ;
  assign n11442 = ~x97 & n5896 ;
  assign n11443 = x108 | n11442 ;
  assign n11444 = ~n1252 & n11443 ;
  assign n11445 = ~n8405 & n11444 ;
  assign n11446 = ~n5900 & n8430 ;
  assign n11447 = n11445 & n11446 ;
  assign n11448 = x51 | n11447 ;
  assign n11449 = n5900 | n8430 ;
  assign n11450 = ( x314 & ~n5898 ) | ( x314 & n11449 ) | ( ~n5898 & n11449 ) ;
  assign n11451 = ( x314 & n11445 ) | ( x314 & ~n11449 ) | ( n11445 & ~n11449 ) ;
  assign n11452 = ~n11450 & n11451 ;
  assign n11453 = n11448 | n11452 ;
  assign n11454 = n1976 | n5951 ;
  assign n11455 = n11453 & ~n11454 ;
  assign n11456 = x87 | n11455 ;
  assign n11457 = n4816 | n7113 ;
  assign n11458 = n11456 & ~n11457 ;
  assign n11459 = n1349 & ~n9571 ;
  assign n11460 = n11119 & n11459 ;
  assign n11461 = x82 | x109 ;
  assign n11462 = x111 & ~n11461 ;
  assign n11463 = ~n10297 & n11462 ;
  assign n11464 = ~n1218 & n11463 ;
  assign n11465 = ~n9264 & n11464 ;
  assign n11466 = ~n1387 & n11465 ;
  assign n11467 = x314 & n11466 ;
  assign n11468 = n8582 & n11413 ;
  assign n11469 = n11467 | n11468 ;
  assign n11470 = ~n8332 & n11469 ;
  assign n11471 = x72 & ~n8498 ;
  assign n11472 = ~x314 & n11466 ;
  assign n11473 = ~n7396 & n11472 ;
  assign n11474 = n11471 | n11473 ;
  assign n11475 = n4904 | n8331 ;
  assign n11476 = n11474 & ~n11475 ;
  assign n11477 = x124 & ~x468 ;
  assign n11478 = ~x99 & n8558 ;
  assign n11479 = ~n8551 & n11478 ;
  assign n11480 = x113 & ~n8660 ;
  assign n11481 = ~n11479 & n11480 ;
  assign n11482 = ~x113 & n8916 ;
  assign n11483 = x228 & ~n11482 ;
  assign n11484 = ~n11481 & n11483 ;
  assign n11485 = x113 & ~n8695 ;
  assign n11486 = n8702 | n11485 ;
  assign n11487 = ( ~x39 & n8693 ) | ( ~x39 & n11486 ) | ( n8693 & n11486 ) ;
  assign n11488 = ~n11484 & n11487 ;
  assign n11489 = n1975 | n11488 ;
  assign n11490 = ~x39 & n8659 ;
  assign n11491 = x38 & ~n11490 ;
  assign n11492 = n4793 & n8507 ;
  assign n11493 = ~x113 & n11492 ;
  assign n11494 = n11286 & n11493 ;
  assign n11495 = n5984 & ~n8732 ;
  assign n11496 = n11492 & ~n11495 ;
  assign n11497 = ( ~n8507 & n8659 ) | ( ~n8507 & n11496 ) | ( n8659 & n11496 ) ;
  assign n11498 = n11494 | n11497 ;
  assign n11499 = ~x39 & n11498 ;
  assign n11500 = n4807 & ~n11499 ;
  assign n11501 = n11491 | n11500 ;
  assign n11502 = n11489 & ~n11501 ;
  assign n11503 = x87 | n11502 ;
  assign n11504 = n8659 & ~n8760 ;
  assign n11505 = ~x113 & n11298 ;
  assign n11506 = n11504 | n11505 ;
  assign n11507 = ~n2041 & n11506 ;
  assign n11508 = n1975 & n11490 ;
  assign n11509 = x87 & ~n11508 ;
  assign n11510 = ~n11507 & n11509 ;
  assign n11511 = n11503 & ~n11510 ;
  assign n11512 = x75 | n11511 ;
  assign n11513 = n5927 & n11494 ;
  assign n11514 = n4793 & ~n8773 ;
  assign n11515 = n8507 & ~n11514 ;
  assign n11516 = n8659 & ~n11515 ;
  assign n11517 = n11513 | n11516 ;
  assign n11518 = ~n1984 & n11517 ;
  assign n11519 = n2007 & n11490 ;
  assign n11520 = x75 & ~n11519 ;
  assign n11521 = ~n11518 & n11520 ;
  assign n11522 = n11512 & ~n11521 ;
  assign n11523 = n7113 | n11522 ;
  assign n11524 = n7113 & ~n11490 ;
  assign n11525 = n11523 & ~n11524 ;
  assign n11526 = x114 & ~n8962 ;
  assign n11527 = n8739 & ~n11526 ;
  assign n11528 = ~n8771 & n11527 ;
  assign n11529 = ~x72 & x114 ;
  assign n11530 = n8739 | n11529 ;
  assign n11531 = ~n1984 & n11530 ;
  assign n11532 = ~n11528 & n11531 ;
  assign n11533 = ~x39 & n11529 ;
  assign n11534 = n2007 & n11533 ;
  assign n11535 = x75 & ~n11534 ;
  assign n11536 = ~n11532 & n11535 ;
  assign n11537 = x115 & ~n11529 ;
  assign n11538 = x39 | n11537 ;
  assign n11539 = ( ~x114 & x115 ) | ( ~x114 & n8919 ) | ( x115 & n8919 ) ;
  assign n11540 = ( x114 & x115 ) | ( x114 & ~n8909 ) | ( x115 & ~n8909 ) ;
  assign n11541 = n11539 | n11540 ;
  assign n11542 = ~n11538 & n11541 ;
  assign n11543 = n1975 | n11542 ;
  assign n11544 = x114 & ~n8735 ;
  assign n11545 = n8739 & ~n11544 ;
  assign n11546 = ~n8730 & n11545 ;
  assign n11547 = ~x39 & n11530 ;
  assign n11548 = ~n11546 & n11547 ;
  assign n11549 = n4807 & ~n11548 ;
  assign n11550 = x38 & ~n11533 ;
  assign n11551 = x87 | n11550 ;
  assign n11552 = n11549 | n11551 ;
  assign n11553 = n11543 & ~n11552 ;
  assign n11554 = x228 & ~n8733 ;
  assign n11555 = ~x115 & n11554 ;
  assign n11556 = n11529 & ~n11555 ;
  assign n11557 = n1975 | n11556 ;
  assign n11558 = n8758 | n11557 ;
  assign n11559 = n1975 & ~n11533 ;
  assign n11560 = n9307 & ~n11559 ;
  assign n11561 = n11558 & n11560 ;
  assign n11562 = x75 | n11561 ;
  assign n11563 = n11553 | n11562 ;
  assign n11564 = ~n11536 & n11563 ;
  assign n11565 = n7113 | n11564 ;
  assign n11566 = n7113 & ~n11533 ;
  assign n11567 = n11565 & ~n11566 ;
  assign n11568 = x52 | n9272 ;
  assign n11569 = ~x115 & n11568 ;
  assign n11570 = n8728 & n11569 ;
  assign n11571 = n5927 & n11570 ;
  assign n11572 = x115 & ~n8962 ;
  assign n11573 = n8507 & ~n11572 ;
  assign n11574 = ~n11571 & n11573 ;
  assign n11575 = ~x72 & x115 ;
  assign n11576 = n8507 | n11575 ;
  assign n11577 = ~n1984 & n11576 ;
  assign n11578 = ~n11574 & n11577 ;
  assign n11579 = ~x39 & n11575 ;
  assign n11580 = n2007 & n11579 ;
  assign n11581 = x75 & ~n11580 ;
  assign n11582 = ~n11578 & n11581 ;
  assign n11583 = ( ~x39 & x115 ) | ( ~x39 & n8919 ) | ( x115 & n8919 ) ;
  assign n11584 = ( x39 & x115 ) | ( x39 & n8909 ) | ( x115 & n8909 ) ;
  assign n11585 = n11583 & ~n11584 ;
  assign n11586 = n1975 | n11585 ;
  assign n11587 = x115 & ~n8735 ;
  assign n11588 = n8507 & ~n11587 ;
  assign n11589 = ~n11570 & n11588 ;
  assign n11590 = ~x39 & n11576 ;
  assign n11591 = ~n11589 & n11590 ;
  assign n11592 = n4807 & ~n11591 ;
  assign n11593 = x38 & ~n11579 ;
  assign n11594 = x87 | n11593 ;
  assign n11595 = n11592 | n11594 ;
  assign n11596 = n11586 & ~n11595 ;
  assign n11597 = ~n11554 & n11575 ;
  assign n11598 = n1975 | n11597 ;
  assign n11599 = n8757 | n11598 ;
  assign n11600 = n1975 & ~n11579 ;
  assign n11601 = n9307 & ~n11600 ;
  assign n11602 = n11599 & n11601 ;
  assign n11603 = x75 | n11602 ;
  assign n11604 = n11596 | n11603 ;
  assign n11605 = ~n11582 & n11604 ;
  assign n11606 = n7113 | n11605 ;
  assign n11607 = n7113 & ~n11579 ;
  assign n11608 = n11606 & ~n11607 ;
  assign n11609 = x116 & ~n8682 ;
  assign n11610 = n1288 | n11609 ;
  assign n11611 = n1288 & n8662 ;
  assign n11612 = x116 & ~n11611 ;
  assign n11613 = n8669 | n11612 ;
  assign n11614 = n11610 & n11613 ;
  assign n11615 = ~n1288 & n8676 ;
  assign n11616 = x228 & ~n11615 ;
  assign n11617 = ~n11614 & n11616 ;
  assign n11618 = x116 & ~n8697 ;
  assign n11619 = n8913 | n11618 ;
  assign n11620 = ~x39 & n11619 ;
  assign n11621 = ~n11617 & n11620 ;
  assign n11622 = n1975 | n11621 ;
  assign n11623 = ~x72 & x116 ;
  assign n11624 = ~n8507 & n11623 ;
  assign n11625 = ~x113 & n11495 ;
  assign n11626 = n11623 & ~n11625 ;
  assign n11627 = n8728 | n11626 ;
  assign n11628 = n11492 & n11627 ;
  assign n11629 = n11624 | n11628 ;
  assign n11630 = ~x39 & n11629 ;
  assign n11631 = n4807 & ~n11630 ;
  assign n11632 = ~x39 & n11623 ;
  assign n11633 = x38 & ~n11632 ;
  assign n11634 = x87 | n11633 ;
  assign n11635 = n11631 | n11634 ;
  assign n11636 = n11622 & ~n11635 ;
  assign n11637 = ( ~x100 & n9307 ) | ( ~x100 & n11632 ) | ( n9307 & n11632 ) ;
  assign n11638 = ~x113 & n8760 ;
  assign n11639 = n11623 & ~n11638 ;
  assign n11640 = x38 | n11639 ;
  assign n11641 = n8756 | n11640 ;
  assign n11642 = ~n11633 & n11641 ;
  assign n11643 = ( x100 & n9307 ) | ( x100 & n11642 ) | ( n9307 & n11642 ) ;
  assign n11644 = n11637 & n11643 ;
  assign n11645 = x75 | n11644 ;
  assign n11646 = n11636 | n11645 ;
  assign n11647 = ~n8774 & n11623 ;
  assign n11648 = n8964 | n11647 ;
  assign n11649 = n11492 & n11648 ;
  assign n11650 = n11624 | n11649 ;
  assign n11651 = ~n1984 & n11650 ;
  assign n11652 = n2007 & n11632 ;
  assign n11653 = x75 & ~n11652 ;
  assign n11654 = ~n11651 & n11653 ;
  assign n11655 = n11646 & ~n11654 ;
  assign n11656 = n7113 | n11655 ;
  assign n11657 = n7113 & ~n11632 ;
  assign n11658 = n11656 & ~n11657 ;
  assign n11659 = n2418 & ~n5822 ;
  assign n11660 = n2417 | n11659 ;
  assign n11661 = ~x38 & n11660 ;
  assign n11662 = x87 | n11661 ;
  assign n11663 = ~n4816 & n11662 ;
  assign n11664 = x92 | n11663 ;
  assign n11665 = x54 | n5766 ;
  assign n11666 = x74 | n11665 ;
  assign n11667 = n11664 & ~n11666 ;
  assign n11668 = x55 | n11667 ;
  assign n11669 = ~n5759 & n11668 ;
  assign n11670 = x56 | n11669 ;
  assign n11671 = ~n4653 & n11670 ;
  assign n11672 = x62 | n11671 ;
  assign n11673 = ~n4828 & n11672 ;
  assign n11674 = x163 & ~n4713 ;
  assign n11675 = n9808 | n11674 ;
  assign n11676 = ~x150 & n11675 ;
  assign n11677 = x150 & ~n9803 ;
  assign n11678 = ~n9806 & n11677 ;
  assign n11679 = n11676 | n11678 ;
  assign n11680 = x232 & n11679 ;
  assign n11681 = n7219 & n11680 ;
  assign n11682 = x74 & ~n11681 ;
  assign n11683 = x165 & n5924 ;
  assign n11684 = x38 | x54 ;
  assign n11685 = ~n11683 & n11684 ;
  assign n11686 = ~n7219 & n11685 ;
  assign n11687 = x74 | n11681 ;
  assign n11688 = n11686 | n11687 ;
  assign n11689 = ~n11682 & n11688 ;
  assign n11690 = n2058 & ~n11689 ;
  assign n11691 = n2057 | n11690 ;
  assign n11692 = n8073 & n11691 ;
  assign n11693 = ( x232 & ~x299 ) | ( x232 & n11679 ) | ( ~x299 & n11679 ) ;
  assign n11694 = ~x185 & n9836 ;
  assign n11695 = ( n4713 & n9836 ) | ( n4713 & ~n11694 ) | ( n9836 & ~n11694 ) ;
  assign n11696 = ( x185 & n11694 ) | ( x185 & ~n11695 ) | ( n11694 & ~n11695 ) ;
  assign n11697 = ( x232 & x299 ) | ( x232 & n11696 ) | ( x299 & n11696 ) ;
  assign n11698 = n11693 & n11697 ;
  assign n11699 = n7219 & n11698 ;
  assign n11700 = x74 & ~n11699 ;
  assign n11701 = x55 | n11700 ;
  assign n11702 = ( x143 & x299 ) | ( x143 & n5924 ) | ( x299 & n5924 ) ;
  assign n11703 = ( x165 & ~x299 ) | ( x165 & n5924 ) | ( ~x299 & n5924 ) ;
  assign n11704 = n11702 & n11703 ;
  assign n11705 = n7219 | n11704 ;
  assign n11706 = x54 & n11705 ;
  assign n11707 = ~n11699 & n11706 ;
  assign n11708 = x143 & ~x165 ;
  assign n11709 = n7253 & n11708 ;
  assign n11710 = x38 & ~n11709 ;
  assign n11711 = ( x143 & x165 ) | ( x143 & n7259 ) | ( x165 & n7259 ) ;
  assign n11712 = ( ~x143 & x165 ) | ( ~x143 & n7256 ) | ( x165 & n7256 ) ;
  assign n11713 = n11711 & n11712 ;
  assign n11714 = n11710 & ~n11713 ;
  assign n11715 = n1924 | n11714 ;
  assign n11716 = n4713 & ~n7548 ;
  assign n11717 = x151 & ~x168 ;
  assign n11718 = n7615 & n11717 ;
  assign n11719 = ( x151 & x168 ) | ( x151 & ~n7623 ) | ( x168 & ~n7623 ) ;
  assign n11720 = ( ~x151 & x168 ) | ( ~x151 & n7620 ) | ( x168 & n7620 ) ;
  assign n11721 = ~n11719 & n11720 ;
  assign n11722 = n11718 | n11721 ;
  assign n11723 = ~n11716 & n11722 ;
  assign n11724 = n4713 & n7548 ;
  assign n11725 = ~n4713 & n7583 ;
  assign n11726 = n11724 | n11725 ;
  assign n11727 = x151 & x168 ;
  assign n11728 = n11726 & n11727 ;
  assign n11729 = x150 & ~n11728 ;
  assign n11730 = ~n11723 & n11729 ;
  assign n11731 = n7459 | n11724 ;
  assign n11732 = x168 & ~n11731 ;
  assign n11733 = n7637 | n11724 ;
  assign n11734 = ( x151 & n11727 ) | ( x151 & n11733 ) | ( n11727 & n11733 ) ;
  assign n11735 = ~n11732 & n11734 ;
  assign n11736 = x168 & ~n7567 ;
  assign n11737 = x168 & ~n4713 ;
  assign n11738 = n7548 | n11737 ;
  assign n11739 = ~x151 & n11738 ;
  assign n11740 = ~n11736 & n11739 ;
  assign n11741 = x150 | n11740 ;
  assign n11742 = n11735 | n11741 ;
  assign n11743 = x299 & n11742 ;
  assign n11744 = ~n11730 & n11743 ;
  assign n11745 = n7572 & ~n11716 ;
  assign n11746 = x173 | n11745 ;
  assign n11747 = ~n4713 & n7403 ;
  assign n11748 = x173 & ~n11724 ;
  assign n11749 = ~n11747 & n11748 ;
  assign n11750 = x185 & ~n11749 ;
  assign n11751 = n11746 & n11750 ;
  assign n11752 = ( x173 & x185 ) | ( x173 & ~n11731 ) | ( x185 & ~n11731 ) ;
  assign n11753 = n7567 & ~n11716 ;
  assign n11754 = ( x173 & ~x185 ) | ( x173 & n11753 ) | ( ~x185 & n11753 ) ;
  assign n11755 = ~n11752 & n11754 ;
  assign n11756 = x190 & ~n11755 ;
  assign n11757 = ~n11751 & n11756 ;
  assign n11758 = x185 & ~n11716 ;
  assign n11759 = ( ~x173 & n4713 ) | ( ~x173 & n7560 ) | ( n4713 & n7560 ) ;
  assign n11760 = ( x173 & n4713 ) | ( x173 & n8084 ) | ( n4713 & n8084 ) ;
  assign n11761 = n11759 | n11760 ;
  assign n11762 = n11758 & n11761 ;
  assign n11763 = ( x173 & x185 ) | ( x173 & ~n11733 ) | ( x185 & ~n11733 ) ;
  assign n11764 = ( x173 & ~x185 ) | ( x173 & n7548 ) | ( ~x185 & n7548 ) ;
  assign n11765 = ~n11763 & n11764 ;
  assign n11766 = x190 | n11765 ;
  assign n11767 = n11762 | n11766 ;
  assign n11768 = ~n11757 & n11767 ;
  assign n11769 = ( x232 & n7916 ) | ( x232 & ~n11768 ) | ( n7916 & ~n11768 ) ;
  assign n11770 = ~n11744 & n11769 ;
  assign n11771 = ( ~x39 & n5788 ) | ( ~x39 & n7548 ) | ( n5788 & n7548 ) ;
  assign n11772 = ~n11770 & n11771 ;
  assign n11773 = x178 | x299 ;
  assign n11774 = x168 & n7288 ;
  assign n11775 = x157 & n7299 ;
  assign n11776 = n11774 | n11775 ;
  assign n11777 = ~n4713 & n9954 ;
  assign n11778 = n11776 & n11777 ;
  assign n11779 = x299 & ~n11778 ;
  assign n11780 = n11773 & ~n11779 ;
  assign n11781 = n7265 | n11780 ;
  assign n11782 = x178 & ~n7321 ;
  assign n11783 = x190 | n11782 ;
  assign n11784 = ~x299 & n11783 ;
  assign n11785 = n11781 & ~n11784 ;
  assign n11786 = ( n4764 & n7285 ) | ( n4764 & n7319 ) | ( n7285 & n7319 ) ;
  assign n11787 = x178 & n11786 ;
  assign n11788 = ~n7328 & n11787 ;
  assign n11789 = ~x178 & n11786 ;
  assign n11790 = ~n7291 & n11789 ;
  assign n11791 = ~x299 & n7286 ;
  assign n11792 = x190 & n11791 ;
  assign n11793 = ~n11790 & n11792 ;
  assign n11794 = ~n11788 & n11793 ;
  assign n11795 = x232 & ~n11794 ;
  assign n11796 = ~n11785 & n11795 ;
  assign n11797 = x232 | n7265 ;
  assign n11798 = ~n11796 & n11797 ;
  assign n11799 = ( x38 & n1925 ) | ( x38 & n11798 ) | ( n1925 & n11798 ) ;
  assign n11800 = n11772 | n11799 ;
  assign n11801 = ~n11715 & n11800 ;
  assign n11802 = x100 & ~n11698 ;
  assign n11803 = x38 & ~n11704 ;
  assign n11804 = n6015 & ~n11803 ;
  assign n11805 = n7709 & n11804 ;
  assign n11806 = n11802 | n11805 ;
  assign n11807 = n11801 | n11806 ;
  assign n11808 = ~n2004 & n11807 ;
  assign n11809 = x75 & ~n11698 ;
  assign n11810 = x100 | n11803 ;
  assign n11811 = ~x157 & x299 ;
  assign n11812 = n11773 & ~n11811 ;
  assign n11813 = n5924 & n11812 ;
  assign n11814 = ~n7684 & n11813 ;
  assign n11815 = n7709 | n11814 ;
  assign n11816 = ~n11810 & n11815 ;
  assign n11817 = n11802 | n11816 ;
  assign n11818 = n7679 & n11817 ;
  assign n11819 = n11809 | n11818 ;
  assign n11820 = n11808 | n11819 ;
  assign n11821 = ~x54 & n11820 ;
  assign n11822 = n11707 | n11821 ;
  assign n11823 = ~x74 & n11822 ;
  assign n11824 = n11701 | n11823 ;
  assign n11825 = x55 & ~n11682 ;
  assign n11826 = x150 & n5924 ;
  assign n11827 = x92 | n7684 ;
  assign n11828 = n11826 & ~n11827 ;
  assign n11829 = n7265 | n11684 ;
  assign n11830 = n11828 | n11829 ;
  assign n11831 = ~n11685 & n11830 ;
  assign n11832 = n7219 | n11831 ;
  assign n11833 = ~n11687 & n11832 ;
  assign n11834 = n11825 & ~n11833 ;
  assign n11835 = n2058 | n11834 ;
  assign n11836 = n11824 & ~n11835 ;
  assign n11837 = n11692 | n11836 ;
  assign n11838 = ( n2057 & n7219 ) | ( n2057 & ~n11683 ) | ( n7219 & ~n11683 ) ;
  assign n11839 = ( n2057 & ~n7219 ) | ( n2057 & n11680 ) | ( ~n7219 & n11680 ) ;
  assign n11840 = n11838 & n11839 ;
  assign n11841 = ~n11682 & n11840 ;
  assign n11842 = n11837 & ~n11841 ;
  assign n11843 = x79 | n10013 ;
  assign n11844 = ( x118 & n11842 ) | ( x118 & ~n11843 ) | ( n11842 & ~n11843 ) ;
  assign n11845 = n4714 & n4997 ;
  assign n11846 = ~x157 & n7754 ;
  assign n11847 = x168 & ~n11846 ;
  assign n11848 = x157 & ~n7759 ;
  assign n11849 = x157 | x168 ;
  assign n11850 = n7757 | n11849 ;
  assign n11851 = ~n11848 & n11850 ;
  assign n11852 = ~n11847 & n11851 ;
  assign n11853 = n11845 | n11852 ;
  assign n11854 = n11170 & n11853 ;
  assign n11855 = ~x178 & n4764 ;
  assign n11856 = n7753 & n11855 ;
  assign n11857 = n11845 | n11856 ;
  assign n11858 = x190 & n11857 ;
  assign n11859 = x178 | n11200 ;
  assign n11860 = x178 & ~n7739 ;
  assign n11861 = ~n11845 & n11860 ;
  assign n11862 = x190 | n11861 ;
  assign n11863 = n11859 & ~n11862 ;
  assign n11864 = n11858 | n11863 ;
  assign n11865 = n11172 & n11864 ;
  assign n11866 = x232 & ~n11865 ;
  assign n11867 = ~n11854 & n11866 ;
  assign n11868 = n5773 & n7747 ;
  assign n11869 = n4723 & n11170 ;
  assign n11870 = n4997 & n11869 ;
  assign n11871 = n11868 | n11870 ;
  assign n11872 = ( x39 & n8469 ) | ( x39 & n11871 ) | ( n8469 & n11871 ) ;
  assign n11873 = ~n11867 & n11872 ;
  assign n11874 = n7808 & n11717 ;
  assign n11875 = ( x151 & x168 ) | ( x151 & ~n7802 ) | ( x168 & ~n7802 ) ;
  assign n11876 = ( ~x151 & x168 ) | ( ~x151 & n7788 ) | ( x168 & n7788 ) ;
  assign n11877 = ~n11875 & n11876 ;
  assign n11878 = n11874 | n11877 ;
  assign n11879 = ~n7790 & n11878 ;
  assign n11880 = x150 & ~n11879 ;
  assign n11881 = ~x151 & n7778 ;
  assign n11882 = n7826 | n11881 ;
  assign n11883 = ~x168 & n11882 ;
  assign n11884 = ~x151 & n7798 ;
  assign n11885 = n7829 | n11884 ;
  assign n11886 = n11737 & n11885 ;
  assign n11887 = x150 | n11886 ;
  assign n11888 = n11883 | n11887 ;
  assign n11889 = ~n11880 & n11888 ;
  assign n11890 = n7778 | n9871 ;
  assign n11891 = n4713 & n11890 ;
  assign n11892 = x299 & ~n11891 ;
  assign n11893 = ~n11889 & n11892 ;
  assign n11894 = x190 | n4713 ;
  assign n11895 = ( x173 & n4904 ) | ( x173 & ~n7808 ) | ( n4904 & ~n7808 ) ;
  assign n11896 = ( x173 & ~n4904 ) | ( x173 & n7788 ) | ( ~n4904 & n7788 ) ;
  assign n11897 = ~n11895 & n11896 ;
  assign n11898 = ~n11894 & n11897 ;
  assign n11899 = ~x173 & x190 ;
  assign n11900 = n7803 & n11899 ;
  assign n11901 = x185 & ~n11900 ;
  assign n11902 = ~n11898 & n11901 ;
  assign n11903 = ~x173 & n7778 ;
  assign n11904 = n7816 | n11903 ;
  assign n11905 = ~x190 & n11904 ;
  assign n11906 = x173 & ~n7814 ;
  assign n11907 = x190 & n7800 ;
  assign n11908 = ~n11906 & n11907 ;
  assign n11909 = x185 | n11908 ;
  assign n11910 = n11905 | n11909 ;
  assign n11911 = ~n11902 & n11910 ;
  assign n11912 = n4713 & n7782 ;
  assign n11913 = x299 | n11912 ;
  assign n11914 = n11911 | n11913 ;
  assign n11915 = ~n11893 & n11914 ;
  assign n11916 = x232 & ~n11915 ;
  assign n11917 = ~n4694 & n7780 ;
  assign n11918 = n7778 | n11917 ;
  assign n11919 = ( ~x39 & n5788 ) | ( ~x39 & n11918 ) | ( n5788 & n11918 ) ;
  assign n11920 = ~n11916 & n11919 ;
  assign n11921 = n11873 | n11920 ;
  assign n11922 = ~x38 & n11921 ;
  assign n11923 = n11715 | n11922 ;
  assign n11924 = n11802 | n11804 ;
  assign n11925 = n11923 & ~n11924 ;
  assign n11926 = n2004 | n11925 ;
  assign n11927 = n7195 | n11813 ;
  assign n11928 = n1868 | n11927 ;
  assign n11929 = ~n11810 & n11928 ;
  assign n11930 = n11802 | n11929 ;
  assign n11931 = n7679 & n11930 ;
  assign n11932 = n11809 | n11931 ;
  assign n11933 = n11926 & ~n11932 ;
  assign n11934 = x54 | n11933 ;
  assign n11935 = ~n11707 & n11934 ;
  assign n11936 = x74 | n11935 ;
  assign n11937 = ~n11701 & n11936 ;
  assign n11938 = x54 & n11683 ;
  assign n11939 = x92 | n7219 ;
  assign n11940 = n7195 | n11939 ;
  assign n11941 = n11826 | n11940 ;
  assign n11942 = n11938 | n11941 ;
  assign n11943 = n1868 | n11942 ;
  assign n11944 = ~n11688 & n11943 ;
  assign n11945 = n11825 & ~n11944 ;
  assign n11946 = n2058 | n11945 ;
  assign n11947 = n11937 | n11946 ;
  assign n11948 = ~n11691 & n11947 ;
  assign n11949 = n11841 | n11948 ;
  assign n11950 = ( x118 & n11843 ) | ( x118 & n11949 ) | ( n11843 & n11949 ) ;
  assign n11951 = ~n11844 & n11950 ;
  assign n11952 = ~x118 & n7206 ;
  assign n11953 = ( ~n11843 & n11949 ) | ( ~n11843 & n11952 ) | ( n11949 & n11952 ) ;
  assign n11954 = ( n11842 & n11843 ) | ( n11842 & n11952 ) | ( n11843 & n11952 ) ;
  assign n11955 = n11953 & ~n11954 ;
  assign n11956 = n11951 | n11955 ;
  assign n11957 = x128 & x228 ;
  assign n11958 = n8329 & n11957 ;
  assign n11959 = x87 & ~n11957 ;
  assign n11960 = x75 | n11959 ;
  assign n11961 = n1823 & ~n2213 ;
  assign n11962 = n5939 & n11961 ;
  assign n11963 = n2203 & n4343 ;
  assign n11964 = n5943 & n11963 ;
  assign n11965 = n11962 | n11964 ;
  assign n11966 = x39 & n11965 ;
  assign n11967 = x299 & n4956 ;
  assign n11968 = n4923 | n11967 ;
  assign n11969 = n5924 & n11968 ;
  assign n11970 = ~n1327 & n8323 ;
  assign n11971 = n9792 | n11970 ;
  assign n11972 = ~n1347 & n11971 ;
  assign n11973 = x97 | n11972 ;
  assign n11974 = ~x46 & n1292 ;
  assign n11975 = ~n1623 & n11974 ;
  assign n11976 = n11973 & n11975 ;
  assign n11977 = x109 & ~n11969 ;
  assign n11978 = ~n1292 & n9793 ;
  assign n11979 = n11977 | n11978 ;
  assign n11980 = n11976 | n11979 ;
  assign n11981 = ( ~n1454 & n11969 ) | ( ~n1454 & n11980 ) | ( n11969 & n11980 ) ;
  assign n11982 = ( n4927 & n11969 ) | ( n4927 & ~n11980 ) | ( n11969 & ~n11980 ) ;
  assign n11983 = n11981 & ~n11982 ;
  assign n11984 = x91 | n11983 ;
  assign n11985 = n1527 | n4883 ;
  assign n11986 = n11984 & ~n11985 ;
  assign n11987 = n1647 | n11986 ;
  assign n11988 = x39 | n9243 ;
  assign n11989 = n11987 & ~n11988 ;
  assign n11990 = n11966 | n11989 ;
  assign n11991 = ~x38 & n11990 ;
  assign n11992 = ~x228 & n11991 ;
  assign n11993 = n11957 | n11992 ;
  assign n11994 = ( x87 & ~x100 ) | ( x87 & n11993 ) | ( ~x100 & n11993 ) ;
  assign n11995 = n1925 | n2082 ;
  assign n11996 = ~n11957 & n11995 ;
  assign n11997 = ( x87 & x100 ) | ( x87 & ~n11996 ) | ( x100 & ~n11996 ) ;
  assign n11998 = n11994 | n11997 ;
  assign n11999 = ~n11960 & n11998 ;
  assign n12000 = n5826 | n7195 ;
  assign n12001 = ~n11957 & n12000 ;
  assign n12002 = x75 & ~n12001 ;
  assign n12003 = x92 | n12002 ;
  assign n12004 = n11999 | n12003 ;
  assign n12005 = x92 & ~n11957 ;
  assign n12006 = n5836 & n12005 ;
  assign n12007 = n8329 | n12006 ;
  assign n12008 = n12004 & ~n12007 ;
  assign n12009 = n11958 | n12008 ;
  assign n12010 = x31 | x80 ;
  assign n12011 = x818 & ~n12010 ;
  assign n12012 = n5880 & n6412 ;
  assign n12013 = n6153 & ~n12012 ;
  assign n12014 = ~x120 & n5880 ;
  assign n12015 = ~x1093 & n12014 ;
  assign n12016 = n12013 & ~n12015 ;
  assign n12017 = ~n1925 & n6417 ;
  assign n12018 = ~n1868 & n5930 ;
  assign n12019 = x120 & ~n6412 ;
  assign n12020 = ~n5987 & n12019 ;
  assign n12021 = ~x120 & x1093 ;
  assign n12022 = n5987 & ~n12021 ;
  assign n12023 = ( n12018 & ~n12020 ) | ( n12018 & n12022 ) | ( ~n12020 & n12022 ) ;
  assign n12024 = n12017 & n12023 ;
  assign n12025 = ~x1091 & n10833 ;
  assign n12026 = n12021 & ~n12025 ;
  assign n12027 = n12019 | n12026 ;
  assign n12028 = x100 & n12027 ;
  assign n12029 = ~n12024 & n12028 ;
  assign n12030 = x1093 | n5915 ;
  assign n12031 = x120 & ~n12030 ;
  assign n12032 = x39 | n12031 ;
  assign n12033 = n5955 & n8529 ;
  assign n12034 = n5905 & n5950 ;
  assign n12035 = ( x122 & ~n5884 ) | ( x122 & n12034 ) | ( ~n5884 & n12034 ) ;
  assign n12036 = n12033 | n12035 ;
  assign n12037 = x122 & ~n5906 ;
  assign n12038 = n1287 | n12037 ;
  assign n12039 = n12036 & ~n12038 ;
  assign n12040 = n1690 & ~n12039 ;
  assign n12041 = n5995 & ~n12034 ;
  assign n12042 = ~n10833 & n12041 ;
  assign n12043 = n12040 | n12042 ;
  assign n12044 = n12032 | n12043 ;
  assign n12045 = n6448 | n12027 ;
  assign n12046 = ~x299 & n12045 ;
  assign n12047 = n4714 | n12027 ;
  assign n12048 = ~n5938 & n12019 ;
  assign n12049 = x1091 & x1092 ;
  assign n12050 = n5936 & n12049 ;
  assign n12051 = n12026 & ~n12050 ;
  assign n12052 = n12048 | n12051 ;
  assign n12053 = n4714 & ~n12052 ;
  assign n12054 = n12047 & ~n12053 ;
  assign n12055 = ( n4764 & n6448 ) | ( n4764 & ~n12054 ) | ( n6448 & ~n12054 ) ;
  assign n12056 = n4751 & n12027 ;
  assign n12057 = ~n4751 & n12052 ;
  assign n12058 = n12056 | n12057 ;
  assign n12059 = ( n4764 & ~n6448 ) | ( n4764 & n12058 ) | ( ~n6448 & n12058 ) ;
  assign n12060 = n12055 & ~n12059 ;
  assign n12061 = n12046 & ~n12060 ;
  assign n12062 = n6433 | n12027 ;
  assign n12063 = x299 & n12062 ;
  assign n12064 = ( n4721 & n6433 ) | ( n4721 & ~n12054 ) | ( n6433 & ~n12054 ) ;
  assign n12065 = ( n4721 & ~n6433 ) | ( n4721 & n12058 ) | ( ~n6433 & n12058 ) ;
  assign n12066 = n12064 & ~n12065 ;
  assign n12067 = n12063 & ~n12066 ;
  assign n12068 = x39 & ~n12067 ;
  assign n12069 = ~n12061 & n12068 ;
  assign n12070 = n12044 & ~n12069 ;
  assign n12071 = x38 | n12070 ;
  assign n12072 = x38 & n6412 ;
  assign n12073 = x120 | x1093 ;
  assign n12074 = x38 & ~n12073 ;
  assign n12075 = x100 | n12074 ;
  assign n12076 = n12072 | n12075 ;
  assign n12077 = n12071 & ~n12076 ;
  assign n12078 = n12029 | n12077 ;
  assign n12079 = ~x87 & n12078 ;
  assign n12080 = n6003 & n12073 ;
  assign n12081 = n5995 & ~n10833 ;
  assign n12082 = ~n6460 & n12081 ;
  assign n12083 = n6001 & ~n12082 ;
  assign n12084 = n1976 & n6412 ;
  assign n12085 = x87 & ~n12084 ;
  assign n12086 = ~n12083 & n12085 ;
  assign n12087 = n12080 & n12086 ;
  assign n12088 = n12079 | n12087 ;
  assign n12089 = ~x75 & n12088 ;
  assign n12090 = ( x75 & ~n1984 ) | ( x75 & n12027 ) | ( ~n1984 & n12027 ) ;
  assign n12091 = n5925 & ~n12027 ;
  assign n12092 = ~n5931 & n12026 ;
  assign n12093 = x1091 | n6411 ;
  assign n12094 = ~n6404 & n12093 ;
  assign n12095 = x120 & ~n12094 ;
  assign n12096 = n5925 | n12095 ;
  assign n12097 = n12092 | n12096 ;
  assign n12098 = ~n12091 & n12097 ;
  assign n12099 = ( x75 & n1984 ) | ( x75 & n12098 ) | ( n1984 & n12098 ) ;
  assign n12100 = n12090 & n12099 ;
  assign n12101 = n5880 | n12100 ;
  assign n12102 = n12089 | n12101 ;
  assign n12103 = n12016 & n12102 ;
  assign n12104 = n12040 | n12041 ;
  assign n12105 = n12032 | n12104 ;
  assign n12106 = ( n4751 & n4764 ) | ( n4751 & ~n6448 ) | ( n4764 & ~n6448 ) ;
  assign n12107 = x1093 & ~n4714 ;
  assign n12108 = ( n4764 & n6448 ) | ( n4764 & ~n12107 ) | ( n6448 & ~n12107 ) ;
  assign n12109 = ~n12106 & n12108 ;
  assign n12110 = n5938 & n12109 ;
  assign n12111 = ~x299 & n12073 ;
  assign n12112 = ~n12110 & n12111 ;
  assign n12113 = ( n4721 & n4751 ) | ( n4721 & ~n6433 ) | ( n4751 & ~n6433 ) ;
  assign n12114 = ( n4721 & n6433 ) | ( n4721 & ~n12107 ) | ( n6433 & ~n12107 ) ;
  assign n12115 = ~n12113 & n12114 ;
  assign n12116 = n5938 & n12115 ;
  assign n12117 = x299 & n12073 ;
  assign n12118 = ~n12116 & n12117 ;
  assign n12119 = x39 & ~n12118 ;
  assign n12120 = ~n12112 & n12119 ;
  assign n12121 = n12105 & ~n12120 ;
  assign n12122 = x38 | n12121 ;
  assign n12123 = ~n12075 & n12122 ;
  assign n12124 = x120 & n5987 ;
  assign n12125 = ~x120 & n12018 ;
  assign n12126 = n12124 | n12125 ;
  assign n12127 = n12017 & n12126 ;
  assign n12128 = x100 & n12073 ;
  assign n12129 = ~n12127 & n12128 ;
  assign n12130 = n12123 | n12129 ;
  assign n12131 = ~x87 & n12130 ;
  assign n12132 = n12080 | n12131 ;
  assign n12133 = ~x75 & n12132 ;
  assign n12134 = n5934 & n12073 ;
  assign n12135 = n5880 | n12134 ;
  assign n12136 = n12133 | n12135 ;
  assign n12137 = n6153 | n12015 ;
  assign n12138 = n12136 & ~n12137 ;
  assign n12139 = n12103 | n12138 ;
  assign n12140 = n12011 & n12139 ;
  assign n12141 = n6785 | n12140 ;
  assign n12142 = n6153 & ~n12027 ;
  assign n12143 = x120 & ~n12142 ;
  assign n12144 = n12011 & n12073 ;
  assign n12145 = ~n12142 & n12144 ;
  assign n12146 = n6785 & ~n12145 ;
  assign n12147 = ~n12143 & n12146 ;
  assign n12148 = n7103 & ~n12147 ;
  assign n12149 = x951 & x982 ;
  assign n12150 = x1092 & n12149 ;
  assign n12151 = x1093 & n12150 ;
  assign n12152 = x120 | n12151 ;
  assign n12153 = ~n12142 & n12152 ;
  assign n12154 = n12146 & ~n12153 ;
  assign n12155 = n7103 | n12154 ;
  assign n12156 = ~n12148 & n12155 ;
  assign n12157 = n12141 & ~n12156 ;
  assign n12158 = x120 & n5932 ;
  assign n12159 = ~x1091 & n12151 ;
  assign n12160 = x120 | n12159 ;
  assign n12161 = n1690 & n12150 ;
  assign n12162 = x93 | x122 ;
  assign n12163 = n1293 | n12162 ;
  assign n12164 = n1289 & ~n7125 ;
  assign n12165 = ~n12163 & n12164 ;
  assign n12166 = ~n1526 & n12165 ;
  assign n12167 = n8499 & n12166 ;
  assign n12168 = n5928 & n12167 ;
  assign n12169 = ~n1254 & n12168 ;
  assign n12170 = n12161 & ~n12169 ;
  assign n12171 = n12160 | n12170 ;
  assign n12172 = ~n12158 & n12171 ;
  assign n12173 = n5925 | n12172 ;
  assign n12174 = ( n1984 & n5926 ) | ( n1984 & ~n12152 ) | ( n5926 & ~n12152 ) ;
  assign n12175 = n12173 & ~n12174 ;
  assign n12176 = n1984 & n12152 ;
  assign n12177 = x75 & ~n12176 ;
  assign n12178 = ~n12175 & n12177 ;
  assign n12179 = n6448 | n12152 ;
  assign n12180 = ~x299 & n12179 ;
  assign n12181 = ~n6605 & n12152 ;
  assign n12182 = ( n4764 & ~n6448 ) | ( n4764 & n12181 ) | ( ~n6448 & n12181 ) ;
  assign n12183 = ~n6602 & n12152 ;
  assign n12184 = ( n4764 & n6448 ) | ( n4764 & ~n12183 ) | ( n6448 & ~n12183 ) ;
  assign n12185 = ~n12182 & n12184 ;
  assign n12186 = n12180 & ~n12185 ;
  assign n12187 = n6433 | n12152 ;
  assign n12188 = x299 & n12187 ;
  assign n12189 = ( n4721 & ~n6433 ) | ( n4721 & n12181 ) | ( ~n6433 & n12181 ) ;
  assign n12190 = ( n4721 & n6433 ) | ( n4721 & ~n12183 ) | ( n6433 & ~n12183 ) ;
  assign n12191 = ~n12189 & n12190 ;
  assign n12192 = n12188 & ~n12191 ;
  assign n12193 = n12186 | n12192 ;
  assign n12194 = x39 & n12193 ;
  assign n12195 = n12030 & ~n12104 ;
  assign n12196 = x120 & n12195 ;
  assign n12197 = n5884 & n12150 ;
  assign n12198 = ~x72 & x950 ;
  assign n12199 = ~n8530 & n12198 ;
  assign n12200 = ~n1328 & n5894 ;
  assign n12201 = ~n1340 & n12200 ;
  assign n12202 = x97 | n12201 ;
  assign n12203 = ~n1626 & n12202 ;
  assign n12204 = ~n1624 & n12203 ;
  assign n12205 = n5956 | n12204 ;
  assign n12206 = ~n1269 & n12205 ;
  assign n12207 = n5888 | n12206 ;
  assign n12208 = ~n5885 & n12207 ;
  assign n12209 = x51 | n12208 ;
  assign n12210 = ~n1465 & n12209 ;
  assign n12211 = ( x96 & n12199 ) | ( x96 & n12210 ) | ( n12199 & n12210 ) ;
  assign n12212 = n12197 & ~n12211 ;
  assign n12213 = ~n7770 & n12201 ;
  assign n12214 = ~n5885 & n12213 ;
  assign n12215 = n5890 | n12214 ;
  assign n12216 = x950 & ~n5951 ;
  assign n12217 = n12215 & n12216 ;
  assign n12218 = x824 & n12217 ;
  assign n12219 = n12150 & ~n12218 ;
  assign n12220 = ~x829 & n12219 ;
  assign n12221 = x829 & x1092 ;
  assign n12222 = x122 & n12149 ;
  assign n12223 = n12221 & n12222 ;
  assign n12224 = ~n12217 & n12223 ;
  assign n12225 = n12220 | n12224 ;
  assign n12226 = n12212 | n12225 ;
  assign n12227 = n5949 & n12226 ;
  assign n12228 = n1287 & n12151 ;
  assign n12229 = n12227 | n12228 ;
  assign n12230 = x1091 & n12229 ;
  assign n12231 = n12159 & ~n12218 ;
  assign n12232 = x120 | n12231 ;
  assign n12233 = n12230 | n12232 ;
  assign n12234 = ~x39 & n12233 ;
  assign n12235 = ~n12196 & n12234 ;
  assign n12236 = n12194 | n12235 ;
  assign n12237 = ~n1975 & n12236 ;
  assign n12238 = n12017 | n12152 ;
  assign n12239 = x950 & ~n1868 ;
  assign n12240 = n5884 & n5928 ;
  assign n12241 = n12239 & n12240 ;
  assign n12242 = n12161 & ~n12241 ;
  assign n12243 = n12160 | n12242 ;
  assign n12244 = ~n12124 & n12243 ;
  assign n12245 = ~x39 & n6417 ;
  assign n12246 = ~n12244 & n12245 ;
  assign n12247 = n4807 & ~n12246 ;
  assign n12248 = ( x38 & n12238 ) | ( x38 & n12247 ) | ( n12238 & n12247 ) ;
  assign n12249 = n12237 | n12248 ;
  assign n12250 = ~x87 & n12249 ;
  assign n12251 = n1976 & ~n12152 ;
  assign n12252 = x87 & ~n12251 ;
  assign n12253 = ~n1287 & n4798 ;
  assign n12254 = n12239 & n12253 ;
  assign n12255 = n12161 & ~n12254 ;
  assign n12256 = x824 & n12239 ;
  assign n12257 = n12159 & ~n12256 ;
  assign n12258 = n12255 | n12257 ;
  assign n12259 = ~x120 & n12258 ;
  assign n12260 = ~n5996 & n6000 ;
  assign n12261 = x120 & ~n12260 ;
  assign n12262 = n1976 | n12261 ;
  assign n12263 = n12259 | n12262 ;
  assign n12264 = n12252 & n12263 ;
  assign n12265 = x75 | n12264 ;
  assign n12266 = n12250 | n12265 ;
  assign n12267 = ~n12178 & n12266 ;
  assign n12268 = n5880 | n12267 ;
  assign n12269 = ~n6153 & n12268 ;
  assign n12270 = ~n10833 & n12159 ;
  assign n12271 = n12242 | n12270 ;
  assign n12272 = ~x120 & n12271 ;
  assign n12273 = n12020 | n12272 ;
  assign n12274 = n6417 & n12273 ;
  assign n12275 = n12027 & n12152 ;
  assign n12276 = ( n1925 & ~n12017 ) | ( n1925 & n12275 ) | ( ~n12017 & n12275 ) ;
  assign n12277 = n12274 | n12276 ;
  assign n12278 = n1925 & ~n12275 ;
  assign n12279 = x100 & ~n12278 ;
  assign n12280 = n12277 & n12279 ;
  assign n12281 = ( x38 & x100 ) | ( x38 & ~n12275 ) | ( x100 & ~n12275 ) ;
  assign n12282 = n12030 & ~n12043 ;
  assign n12283 = x120 & n12282 ;
  assign n12284 = n12081 & n12219 ;
  assign n12285 = x120 | n12284 ;
  assign n12286 = n12230 | n12285 ;
  assign n12287 = ~n12283 & n12286 ;
  assign n12288 = x39 | n12287 ;
  assign n12289 = n6412 & ~n6433 ;
  assign n12290 = n12188 & ~n12289 ;
  assign n12291 = ~n5936 & n12161 ;
  assign n12292 = n12270 | n12291 ;
  assign n12293 = ~x120 & n12292 ;
  assign n12294 = n12048 | n12293 ;
  assign n12295 = n4714 & n12294 ;
  assign n12296 = ~n4714 & n12275 ;
  assign n12297 = n12295 | n12296 ;
  assign n12298 = ( n4721 & n6433 ) | ( n4721 & ~n12297 ) | ( n6433 & ~n12297 ) ;
  assign n12299 = ~n4751 & n12294 ;
  assign n12300 = n4751 & n12275 ;
  assign n12301 = n12299 | n12300 ;
  assign n12302 = ( n4721 & ~n6433 ) | ( n4721 & n12301 ) | ( ~n6433 & n12301 ) ;
  assign n12303 = n12298 & ~n12302 ;
  assign n12304 = n12290 & ~n12303 ;
  assign n12305 = n12045 & n12180 ;
  assign n12306 = ( n4764 & n6448 ) | ( n4764 & ~n12297 ) | ( n6448 & ~n12297 ) ;
  assign n12307 = ( n4764 & ~n6448 ) | ( n4764 & n12301 ) | ( ~n6448 & n12301 ) ;
  assign n12308 = n12306 & ~n12307 ;
  assign n12309 = n12305 & ~n12308 ;
  assign n12310 = x39 & ~n12309 ;
  assign n12311 = ~n12304 & n12310 ;
  assign n12312 = n12288 & ~n12311 ;
  assign n12313 = ( x38 & ~x100 ) | ( x38 & n12312 ) | ( ~x100 & n12312 ) ;
  assign n12314 = ~n12281 & n12313 ;
  assign n12315 = n12280 | n12314 ;
  assign n12316 = ~x87 & n12315 ;
  assign n12317 = ~n12083 & n12262 ;
  assign n12318 = n12255 | n12270 ;
  assign n12319 = n12259 & n12318 ;
  assign n12320 = n12317 | n12319 ;
  assign n12321 = ~n12084 & n12252 ;
  assign n12322 = n12320 & n12321 ;
  assign n12323 = n12316 | n12322 ;
  assign n12324 = ~x75 & n12323 ;
  assign n12325 = ( x75 & ~n1984 ) | ( x75 & n12275 ) | ( ~n1984 & n12275 ) ;
  assign n12326 = n5925 & ~n12275 ;
  assign n12327 = n12170 | n12270 ;
  assign n12328 = ~x120 & n12327 ;
  assign n12329 = n12096 | n12328 ;
  assign n12330 = ~n12326 & n12329 ;
  assign n12331 = ( x75 & n1984 ) | ( x75 & n12330 ) | ( n1984 & n12330 ) ;
  assign n12332 = n12325 & n12331 ;
  assign n12333 = n5880 | n12332 ;
  assign n12334 = n12324 | n12333 ;
  assign n12335 = n12016 & n12334 ;
  assign n12336 = n12269 | n12335 ;
  assign n12337 = n12014 & ~n12151 ;
  assign n12338 = n12155 | n12337 ;
  assign n12339 = n12336 & ~n12338 ;
  assign n12340 = x39 | n12195 ;
  assign n12341 = ~n5947 & n12340 ;
  assign n12342 = x100 | n12341 ;
  assign n12343 = ~n6011 & n12342 ;
  assign n12344 = ( x87 & ~n6003 ) | ( x87 & n12343 ) | ( ~n6003 & n12343 ) ;
  assign n12345 = x75 | n12344 ;
  assign n12346 = ~n5934 & n12345 ;
  assign n12347 = n6153 | n12014 ;
  assign n12348 = n12346 | n12347 ;
  assign n12349 = n5991 & ~n6412 ;
  assign n12350 = x100 | n12072 ;
  assign n12351 = n6412 & ~n6448 ;
  assign n12352 = x299 | n12351 ;
  assign n12353 = ~n6436 & n12093 ;
  assign n12354 = n4714 & ~n12353 ;
  assign n12355 = n4714 | n6412 ;
  assign n12356 = ~n12354 & n12355 ;
  assign n12357 = ( n4764 & n6448 ) | ( n4764 & n12356 ) | ( n6448 & n12356 ) ;
  assign n12358 = n4751 | n12353 ;
  assign n12359 = n4751 & ~n6412 ;
  assign n12360 = n12358 & ~n12359 ;
  assign n12361 = ( ~n4764 & n6448 ) | ( ~n4764 & n12360 ) | ( n6448 & n12360 ) ;
  assign n12362 = n12357 & n12361 ;
  assign n12363 = n12352 | n12362 ;
  assign n12364 = x299 & ~n12289 ;
  assign n12365 = ( n4721 & n6433 ) | ( n4721 & n12356 ) | ( n6433 & n12356 ) ;
  assign n12366 = ( ~n4721 & n6433 ) | ( ~n4721 & n12360 ) | ( n6433 & n12360 ) ;
  assign n12367 = n12365 & n12366 ;
  assign n12368 = n12364 & ~n12367 ;
  assign n12369 = n12363 & ~n12368 ;
  assign n12370 = ( x38 & x39 ) | ( x38 & ~n12369 ) | ( x39 & ~n12369 ) ;
  assign n12371 = ( ~x38 & x39 ) | ( ~x38 & n12282 ) | ( x39 & n12282 ) ;
  assign n12372 = ~n12370 & n12371 ;
  assign n12373 = n12350 | n12372 ;
  assign n12374 = ~n12349 & n12373 ;
  assign n12375 = x87 | n12374 ;
  assign n12376 = ~n12086 & n12375 ;
  assign n12377 = x75 | n12376 ;
  assign n12378 = ( ~x75 & n5926 ) | ( ~x75 & n6412 ) | ( n5926 & n6412 ) ;
  assign n12379 = ( x75 & n5926 ) | ( x75 & ~n12094 ) | ( n5926 & ~n12094 ) ;
  assign n12380 = ~n12378 & n12379 ;
  assign n12381 = n12377 & ~n12380 ;
  assign n12382 = n12013 & ~n12381 ;
  assign n12383 = n5880 & ~n12142 ;
  assign n12384 = n12382 | n12383 ;
  assign n12385 = n12348 & ~n12384 ;
  assign n12386 = x120 & n12148 ;
  assign n12387 = ~n12385 & n12386 ;
  assign n12388 = n12339 | n12387 ;
  assign n12389 = ~n12011 & n12388 ;
  assign n12390 = n12157 | n12389 ;
  assign n12391 = x134 | x135 ;
  assign n12392 = x136 | n12391 ;
  assign n12393 = x130 | n12392 ;
  assign n12394 = x132 | n12393 ;
  assign n12395 = x126 | n12394 ;
  assign n12396 = x121 | n12395 ;
  assign n12397 = x125 | x133 ;
  assign n12398 = x121 & n12397 ;
  assign n12399 = x121 | n12397 ;
  assign n12400 = ~n12398 & n12399 ;
  assign n12401 = n12396 & ~n12400 ;
  assign n12402 = n1230 | n8319 ;
  assign n12403 = x51 | n12402 ;
  assign n12404 = x87 | n12403 ;
  assign n12405 = n12401 | n12404 ;
  assign n12406 = n6785 & n12405 ;
  assign n12407 = ~n4713 & n12403 ;
  assign n12408 = x51 & x146 ;
  assign n12409 = x51 & ~n4713 ;
  assign n12410 = ~x146 & n12409 ;
  assign n12411 = x161 & ~n12410 ;
  assign n12412 = n12408 | n12411 ;
  assign n12413 = n12407 & ~n12412 ;
  assign n12414 = ( x87 & x232 ) | ( x87 & n12413 ) | ( x232 & n12413 ) ;
  assign n12415 = ( ~x87 & x232 ) | ( ~x87 & n11674 ) | ( x232 & n11674 ) ;
  assign n12416 = n12414 & n12415 ;
  assign n12417 = n12406 & ~n12416 ;
  assign n12418 = x299 & ~n12413 ;
  assign n12419 = ~x142 & n12409 ;
  assign n12420 = x144 & ~n12419 ;
  assign n12421 = x51 & x142 ;
  assign n12422 = n12407 & ~n12421 ;
  assign n12423 = ~n12420 & n12422 ;
  assign n12424 = x299 | n12423 ;
  assign n12425 = x232 & n12424 ;
  assign n12426 = ~n12418 & n12425 ;
  assign n12427 = x38 & ~n12426 ;
  assign n12428 = x100 | n12427 ;
  assign n12429 = x38 & n12403 ;
  assign n12430 = x100 | n12429 ;
  assign n12431 = n12428 & n12430 ;
  assign n12432 = n1233 | n8318 ;
  assign n12433 = n11092 | n12432 ;
  assign n12434 = ~x50 & x77 ;
  assign n12435 = ~n5893 & n12434 ;
  assign n12436 = ~n12433 & n12435 ;
  assign n12437 = n1256 | n5899 ;
  assign n12438 = ~x24 & x314 ;
  assign n12439 = ~n12437 & n12438 ;
  assign n12440 = ~n7130 & n12439 ;
  assign n12441 = n12436 & n12440 ;
  assign n12442 = ~n1864 & n12441 ;
  assign n12443 = n1327 | n12433 ;
  assign n12444 = x58 | n12437 ;
  assign n12445 = n7271 | n12444 ;
  assign n12446 = n12443 | n12445 ;
  assign n12447 = x72 & ~n4904 ;
  assign n12448 = ~n12446 & n12447 ;
  assign n12449 = ~n12402 & n12437 ;
  assign n12450 = x51 | n12449 ;
  assign n12451 = x86 & ~n12443 ;
  assign n12452 = n12436 | n12451 ;
  assign n12453 = n9233 & n12452 ;
  assign n12454 = ~x24 & n9788 ;
  assign n12455 = ~n12443 & n12454 ;
  assign n12456 = n12402 | n12455 ;
  assign n12457 = n12453 | n12456 ;
  assign n12458 = ~n12450 & n12457 ;
  assign n12459 = ~n1864 & n12458 ;
  assign n12460 = n12403 | n12442 ;
  assign n12461 = n12459 | n12460 ;
  assign n12462 = n4713 & n12461 ;
  assign n12463 = n12407 | n12462 ;
  assign n12464 = n12448 | n12463 ;
  assign n12465 = n12442 | n12464 ;
  assign n12466 = n12420 & n12465 ;
  assign n12467 = x180 | n12466 ;
  assign n12468 = n12403 | n12459 ;
  assign n12469 = n12448 | n12468 ;
  assign n12470 = n12442 | n12469 ;
  assign n12471 = n4713 & n12470 ;
  assign n12472 = x72 & ~n8615 ;
  assign n12473 = n12409 | n12472 ;
  assign n12474 = ~n4713 & n12473 ;
  assign n12475 = n12471 | n12474 ;
  assign n12476 = ~x51 & n12439 ;
  assign n12477 = n11459 & n12476 ;
  assign n12478 = n1864 | n4713 ;
  assign n12479 = n12477 & ~n12478 ;
  assign n12480 = n12475 | n12479 ;
  assign n12481 = ( x142 & x144 ) | ( x142 & ~n12480 ) | ( x144 & ~n12480 ) ;
  assign n12482 = n4713 & ~n12470 ;
  assign n12483 = x72 | n12477 ;
  assign n12484 = ~n4905 & n12483 ;
  assign n12485 = n4713 | n12484 ;
  assign n12486 = ~n12482 & n12485 ;
  assign n12487 = ( x142 & ~x144 ) | ( x142 & n12486 ) | ( ~x144 & n12486 ) ;
  assign n12488 = ~n12481 & n12487 ;
  assign n12489 = n12467 | n12488 ;
  assign n12490 = ( x144 & n12419 ) | ( x144 & ~n12464 ) | ( n12419 & ~n12464 ) ;
  assign n12491 = ( x144 & ~n12419 ) | ( x144 & n12475 ) | ( ~n12419 & n12475 ) ;
  assign n12492 = ~n12490 & n12491 ;
  assign n12493 = x180 & ~n12492 ;
  assign n12494 = x179 & ~n12493 ;
  assign n12495 = n12489 & n12494 ;
  assign n12496 = n12420 & n12470 ;
  assign n12497 = x180 | n12496 ;
  assign n12498 = x24 | n9789 ;
  assign n12499 = x24 & ~n9794 ;
  assign n12500 = n12498 & ~n12499 ;
  assign n12501 = x314 | n12500 ;
  assign n12502 = x314 & ~n9794 ;
  assign n12503 = n12501 & ~n12502 ;
  assign n12504 = n5899 | n7190 ;
  assign n12505 = n12503 & ~n12504 ;
  assign n12506 = x51 | n12505 ;
  assign n12507 = n12472 | n12506 ;
  assign n12508 = ~n4713 & n12507 ;
  assign n12509 = n12471 | n12508 ;
  assign n12510 = ( x142 & x144 ) | ( x142 & ~n12509 ) | ( x144 & ~n12509 ) ;
  assign n12511 = ~n1259 & n12503 ;
  assign n12512 = x72 | n12511 ;
  assign n12513 = ~n4905 & n12512 ;
  assign n12514 = n4713 | n12513 ;
  assign n12515 = ~n12482 & n12514 ;
  assign n12516 = ( x142 & ~x144 ) | ( x142 & n12515 ) | ( ~x144 & n12515 ) ;
  assign n12517 = ~n12510 & n12516 ;
  assign n12518 = n12497 | n12517 ;
  assign n12519 = x51 | n4713 ;
  assign n12520 = n12469 & ~n12519 ;
  assign n12521 = n12471 | n12520 ;
  assign n12522 = ~n4713 & n12468 ;
  assign n12523 = x142 | n12522 ;
  assign n12524 = ~x51 & n12402 ;
  assign n12525 = ~n4713 & n12524 ;
  assign n12526 = n12478 & ~n12525 ;
  assign n12527 = n1864 | n12458 ;
  assign n12528 = ~n12526 & n12527 ;
  assign n12529 = x142 & ~n12528 ;
  assign n12530 = n12523 & ~n12529 ;
  assign n12531 = n12463 & ~n12530 ;
  assign n12532 = n12521 | n12531 ;
  assign n12533 = x144 & n12532 ;
  assign n12534 = x180 & ~n12533 ;
  assign n12535 = ~n1259 & n12500 ;
  assign n12536 = ~n12478 & n12535 ;
  assign n12537 = n12474 | n12536 ;
  assign n12538 = n12471 | n12537 ;
  assign n12539 = ( x142 & x144 ) | ( x142 & ~n12538 ) | ( x144 & ~n12538 ) ;
  assign n12540 = x72 | n12535 ;
  assign n12541 = ~n4905 & n12540 ;
  assign n12542 = n4713 | n12541 ;
  assign n12543 = ~n12482 & n12542 ;
  assign n12544 = ( x142 & ~x144 ) | ( x142 & n12543 ) | ( ~x144 & n12543 ) ;
  assign n12545 = ~n12539 & n12544 ;
  assign n12546 = n12534 & ~n12545 ;
  assign n12547 = x179 | n12546 ;
  assign n12548 = n12518 & ~n12547 ;
  assign n12549 = n12495 | n12548 ;
  assign n12550 = ~x299 & n12549 ;
  assign n12551 = x161 | n12410 ;
  assign n12552 = n12475 & ~n12551 ;
  assign n12553 = n12402 | n12448 ;
  assign n12554 = ~n12519 & n12553 ;
  assign n12555 = x146 | n12554 ;
  assign n12556 = n12471 | n12555 ;
  assign n12557 = x146 & ~n12464 ;
  assign n12558 = x161 & ~n12557 ;
  assign n12559 = n12556 & n12558 ;
  assign n12560 = n12552 | n12559 ;
  assign n12561 = n7581 & n12560 ;
  assign n12562 = n12519 | n12553 ;
  assign n12563 = n12442 | n12562 ;
  assign n12564 = ~n12409 & n12563 ;
  assign n12565 = x146 & n12403 ;
  assign n12566 = n12564 | n12565 ;
  assign n12567 = x161 & n12566 ;
  assign n12568 = ~n12482 & n12567 ;
  assign n12569 = ( x146 & x161 ) | ( x146 & ~n12480 ) | ( x161 & ~n12480 ) ;
  assign n12570 = ( x146 & ~x161 ) | ( x146 & n12486 ) | ( ~x161 & n12486 ) ;
  assign n12571 = ~n12569 & n12570 ;
  assign n12572 = n12568 | n12571 ;
  assign n12573 = n7610 & n12572 ;
  assign n12574 = n12561 | n12573 ;
  assign n12575 = x156 & n12574 ;
  assign n12576 = ( ~x146 & n7581 ) | ( ~x146 & n12538 ) | ( n7581 & n12538 ) ;
  assign n12577 = ( x146 & n7581 ) | ( x146 & n12543 ) | ( n7581 & n12543 ) ;
  assign n12578 = n12576 & n12577 ;
  assign n12579 = x161 | n12578 ;
  assign n12580 = ( x146 & n7610 ) | ( x146 & n12515 ) | ( n7610 & n12515 ) ;
  assign n12581 = ( ~x146 & n7610 ) | ( ~x146 & n12509 ) | ( n7610 & n12509 ) ;
  assign n12582 = n12580 & n12581 ;
  assign n12583 = n12579 | n12582 ;
  assign n12584 = x146 | n12522 ;
  assign n12585 = x146 & ~n12528 ;
  assign n12586 = n12584 & ~n12585 ;
  assign n12587 = n12463 & ~n12586 ;
  assign n12588 = n12521 | n12587 ;
  assign n12589 = n7581 & n12588 ;
  assign n12590 = n7610 & ~n12410 ;
  assign n12591 = n12470 & n12590 ;
  assign n12592 = x161 & ~n12591 ;
  assign n12593 = ~n12589 & n12592 ;
  assign n12594 = x156 | n12593 ;
  assign n12595 = n12583 & ~n12594 ;
  assign n12596 = n12575 | n12595 ;
  assign n12597 = n12550 | n12596 ;
  assign n12598 = n5788 & n12597 ;
  assign n12599 = n1864 | n12446 ;
  assign n12600 = ~n12403 & n12599 ;
  assign n12601 = n4713 & ~n12600 ;
  assign n12602 = n1463 | n5904 ;
  assign n12603 = ~x51 & n12602 ;
  assign n12604 = n4713 | n12603 ;
  assign n12605 = ~n12601 & n12604 ;
  assign n12606 = ( x146 & x161 ) | ( x146 & ~n12605 ) | ( x161 & ~n12605 ) ;
  assign n12607 = n4738 & ~n12601 ;
  assign n12608 = ( x146 & ~x161 ) | ( x146 & n12607 ) | ( ~x161 & n12607 ) ;
  assign n12609 = ~n12606 & n12608 ;
  assign n12610 = n12411 & ~n12600 ;
  assign n12611 = ( x161 & n12609 ) | ( x161 & ~n12610 ) | ( n12609 & ~n12610 ) ;
  assign n12612 = n5005 & n12611 ;
  assign n12613 = n7296 | n12612 ;
  assign n12614 = x287 | n4713 ;
  assign n12615 = x51 | n12614 ;
  assign n12616 = ~n12605 & n12615 ;
  assign n12617 = ~n12551 & n12616 ;
  assign n12618 = ~n12599 & n12614 ;
  assign n12619 = n12403 | n12618 ;
  assign n12620 = n12411 & n12619 ;
  assign n12621 = n12617 | n12620 ;
  assign n12622 = x216 & n12621 ;
  assign n12623 = n12613 & ~n12622 ;
  assign n12624 = ( n5005 & n12403 ) | ( n5005 & ~n12413 ) | ( n12403 & ~n12413 ) ;
  assign n12625 = n7975 & n12624 ;
  assign n12626 = ~n12623 & n12625 ;
  assign n12627 = ( x142 & n4989 ) | ( x142 & n12607 ) | ( n4989 & n12607 ) ;
  assign n12628 = ( ~x142 & n4989 ) | ( ~x142 & n12605 ) | ( n4989 & n12605 ) ;
  assign n12629 = n12627 & n12628 ;
  assign n12630 = n7285 | n12629 ;
  assign n12631 = x224 & ~n12419 ;
  assign n12632 = n12616 & n12631 ;
  assign n12633 = n12630 & ~n12632 ;
  assign n12634 = n12403 & ~n12419 ;
  assign n12635 = n4989 | n12634 ;
  assign n12636 = x144 & n12635 ;
  assign n12637 = ~n4989 & n12525 ;
  assign n12638 = n12635 & ~n12637 ;
  assign n12639 = ~n12636 & n12638 ;
  assign n12640 = ~n12633 & n12639 ;
  assign n12641 = x51 | n12600 ;
  assign n12642 = ~x287 & n12641 ;
  assign n12643 = ~n12525 & n12614 ;
  assign n12644 = n12642 | n12643 ;
  assign n12645 = ~n12422 & n12644 ;
  assign n12646 = n7285 & ~n12645 ;
  assign n12647 = ~n12402 & n12646 ;
  assign n12648 = x51 & n4713 ;
  assign n12649 = n12641 & ~n12648 ;
  assign n12650 = n4989 & ~n12421 ;
  assign n12651 = n12649 & n12650 ;
  assign n12652 = n12636 & ~n12651 ;
  assign n12653 = ~n12647 & n12652 ;
  assign n12654 = x181 & ~n12653 ;
  assign n12655 = ~n12640 & n12654 ;
  assign n12656 = ~n12629 & n12639 ;
  assign n12657 = x181 | n12652 ;
  assign n12658 = n12656 | n12657 ;
  assign n12659 = ~x299 & n12658 ;
  assign n12660 = ~n12655 & n12659 ;
  assign n12661 = n7974 & n12624 ;
  assign n12662 = ~n12612 & n12661 ;
  assign n12663 = x232 & ~n12662 ;
  assign n12664 = ~n12660 & n12663 ;
  assign n12665 = ~n12626 & n12664 ;
  assign n12666 = n5124 | n5940 ;
  assign n12667 = ~n12599 & n12666 ;
  assign n12668 = n12403 | n12667 ;
  assign n12669 = ( x39 & n8469 ) | ( x39 & n12668 ) | ( n8469 & n12668 ) ;
  assign n12670 = ~n12665 & n12669 ;
  assign n12671 = x39 | x232 ;
  assign n12672 = n12470 & ~n12671 ;
  assign n12673 = n12670 | n12672 ;
  assign n12674 = n12598 | n12673 ;
  assign n12675 = ~x38 & n12674 ;
  assign n12676 = n12431 | n12675 ;
  assign n12677 = x100 & ~n12403 ;
  assign n12678 = n2043 | n12677 ;
  assign n12679 = x100 & n12426 ;
  assign n12680 = n12678 | n12679 ;
  assign n12681 = n12676 & ~n12680 ;
  assign n12682 = ~x87 & n2031 ;
  assign n12683 = n12403 & n12682 ;
  assign n12684 = ~n12426 & n12683 ;
  assign n12685 = x184 | x299 ;
  assign n12686 = ~x163 & x299 ;
  assign n12687 = n12685 & ~n12686 ;
  assign n12688 = n5924 & n12687 ;
  assign n12689 = x87 & ~n12688 ;
  assign n12690 = n12401 | n12689 ;
  assign n12691 = n12684 | n12690 ;
  assign n12692 = n12681 | n12691 ;
  assign n12693 = ~n4713 & n12506 ;
  assign n12694 = ~n12421 & n12693 ;
  assign n12695 = x144 & ~n12694 ;
  assign n12696 = n12402 | n12441 ;
  assign n12697 = n12437 | n12696 ;
  assign n12698 = ( ~n12450 & n12458 ) | ( ~n12450 & n12697 ) | ( n12458 & n12697 ) ;
  assign n12699 = n1864 | n12698 ;
  assign n12700 = ~n12526 & n12699 ;
  assign n12701 = ( x142 & x144 ) | ( x142 & n12700 ) | ( x144 & n12700 ) ;
  assign n12702 = ~n4713 & n12461 ;
  assign n12703 = ( ~x142 & x144 ) | ( ~x142 & n12702 ) | ( x144 & n12702 ) ;
  assign n12704 = n12701 | n12703 ;
  assign n12705 = x180 & n12704 ;
  assign n12706 = ~n12695 & n12705 ;
  assign n12707 = n12420 & ~n12536 ;
  assign n12708 = x144 | n12530 ;
  assign n12709 = ~x180 & n12708 ;
  assign n12710 = ~n12707 & n12709 ;
  assign n12711 = x179 & ~n12710 ;
  assign n12712 = ~n12706 & n12711 ;
  assign n12713 = n12420 & ~n12479 ;
  assign n12714 = ~x51 & n12696 ;
  assign n12715 = n1864 | n12714 ;
  assign n12716 = ~n12526 & n12715 ;
  assign n12717 = ( x142 & x144 ) | ( x142 & n12716 ) | ( x144 & n12716 ) ;
  assign n12718 = ~n4713 & n12460 ;
  assign n12719 = ( ~x142 & x144 ) | ( ~x142 & n12718 ) | ( x144 & n12718 ) ;
  assign n12720 = n12717 | n12719 ;
  assign n12721 = x180 & n12720 ;
  assign n12722 = ~n12713 & n12721 ;
  assign n12723 = ~x180 & n12423 ;
  assign n12724 = x179 | n12723 ;
  assign n12725 = n12722 | n12724 ;
  assign n12726 = ~n12712 & n12725 ;
  assign n12727 = x299 | n12726 ;
  assign n12728 = ~n12408 & n12693 ;
  assign n12729 = x161 & ~n12728 ;
  assign n12730 = ( x146 & x161 ) | ( x146 & n12700 ) | ( x161 & n12700 ) ;
  assign n12731 = ( ~x146 & x161 ) | ( ~x146 & n12702 ) | ( x161 & n12702 ) ;
  assign n12732 = n12730 | n12731 ;
  assign n12733 = ~n12729 & n12732 ;
  assign n12734 = n7581 & ~n12733 ;
  assign n12735 = n12411 & ~n12536 ;
  assign n12736 = x161 | n12586 ;
  assign n12737 = ~n12735 & n12736 ;
  assign n12738 = n7610 & ~n12737 ;
  assign n12739 = x232 & ~n12738 ;
  assign n12740 = ~n12734 & n12739 ;
  assign n12741 = x156 & ~n12740 ;
  assign n12742 = x39 | n12741 ;
  assign n12743 = n12727 & ~n12742 ;
  assign n12744 = n7285 & ~n12614 ;
  assign n12745 = ( x142 & n1868 ) | ( x142 & ~n12744 ) | ( n1868 & ~n12744 ) ;
  assign n12746 = ( x142 & ~n12602 ) | ( x142 & n12744 ) | ( ~n12602 & n12744 ) ;
  assign n12747 = ~n12745 & n12746 ;
  assign n12748 = n12420 & ~n12747 ;
  assign n12749 = x144 | n12422 ;
  assign n12750 = n12646 | n12749 ;
  assign n12751 = x181 & n12750 ;
  assign n12752 = ~n12748 & n12751 ;
  assign n12753 = ~x181 & n12423 ;
  assign n12754 = x299 | n12753 ;
  assign n12755 = n12752 | n12754 ;
  assign n12756 = n4713 | n4981 ;
  assign n12757 = n12411 & n12756 ;
  assign n12758 = ~n12551 & n12644 ;
  assign n12759 = n7296 & ~n12758 ;
  assign n12760 = ~n12757 & n12759 ;
  assign n12761 = ~n7296 & n12413 ;
  assign n12762 = n7975 & ~n12761 ;
  assign n12763 = ~n12760 & n12762 ;
  assign n12764 = ~x159 & n12418 ;
  assign n12765 = n8469 & ~n12764 ;
  assign n12766 = ~n12763 & n12765 ;
  assign n12767 = n12755 & n12766 ;
  assign n12768 = x38 | n12767 ;
  assign n12769 = n12743 | n12768 ;
  assign n12770 = n12411 & ~n12479 ;
  assign n12771 = ( x146 & x161 ) | ( x146 & n12716 ) | ( x161 & n12716 ) ;
  assign n12772 = ( ~x146 & x161 ) | ( ~x146 & n12718 ) | ( x161 & n12718 ) ;
  assign n12773 = n12771 | n12772 ;
  assign n12774 = ~n12770 & n12773 ;
  assign n12775 = n7581 & ~n12774 ;
  assign n12776 = ~x158 & n12418 ;
  assign n12777 = x232 & ~n12776 ;
  assign n12778 = ~n12775 & n12777 ;
  assign n12779 = x156 | n1925 ;
  assign n12780 = n12778 | n12779 ;
  assign n12781 = ~n12428 & n12780 ;
  assign n12782 = n12769 & n12781 ;
  assign n12783 = n2043 | n12679 ;
  assign n12784 = n12782 | n12783 ;
  assign n12785 = ~n12426 & n12682 ;
  assign n12786 = n12401 & ~n12689 ;
  assign n12787 = ~n12785 & n12786 ;
  assign n12788 = n12784 & n12787 ;
  assign n12789 = n6785 | n12788 ;
  assign n12790 = n12692 & ~n12789 ;
  assign n12791 = n12417 | n12790 ;
  assign n12792 = n6412 & n7064 ;
  assign n12793 = ~n5880 & n12346 ;
  assign n12794 = n6153 | n12793 ;
  assign n12795 = ( n5880 & n12013 ) | ( n5880 & n12382 ) | ( n12013 & n12382 ) ;
  assign n12796 = n6785 | n12795 ;
  assign n12797 = n12794 & ~n12796 ;
  assign n12798 = n12792 | n12797 ;
  assign n12799 = x110 & n8244 ;
  assign n12800 = ~n9068 & n12799 ;
  assign n12801 = n4795 & n12800 ;
  assign n12802 = ( x39 & n6785 ) | ( x39 & n12801 ) | ( n6785 & n12801 ) ;
  assign n12803 = ~x110 & n7280 ;
  assign n12804 = n4723 & n5005 ;
  assign n12805 = n12803 & n12804 ;
  assign n12806 = ( ~x39 & n6785 ) | ( ~x39 & n12805 ) | ( n6785 & n12805 ) ;
  assign n12807 = n12802 & n12806 ;
  assign n12808 = x38 | n2032 ;
  assign n12809 = x299 & n12805 ;
  assign n12810 = n4766 & n5940 ;
  assign n12811 = n12803 & n12810 ;
  assign n12812 = x39 & ~n12811 ;
  assign n12813 = ~n12809 & n12812 ;
  assign n12814 = x110 & n11413 ;
  assign n12815 = x39 | n12814 ;
  assign n12816 = ~n12813 & n12815 ;
  assign n12817 = ( n6785 & n12808 ) | ( n6785 & ~n12816 ) | ( n12808 & ~n12816 ) ;
  assign n12818 = x111 | n4856 ;
  assign n12819 = x36 | n1389 ;
  assign n12820 = n12818 & ~n12819 ;
  assign n12821 = n1234 | n12820 ;
  assign n12822 = n1357 | n1398 ;
  assign n12823 = n12821 & ~n12822 ;
  assign n12824 = x83 | n12823 ;
  assign n12825 = ~n1360 & n12824 ;
  assign n12826 = x71 | n12825 ;
  assign n12827 = ~n4863 & n12826 ;
  assign n12828 = x81 | n12827 ;
  assign n12829 = ~n9572 & n12828 ;
  assign n12830 = x90 | n12829 ;
  assign n12831 = ~n1258 & n12830 ;
  assign n12832 = x90 & n8581 ;
  assign n12833 = n7394 | n12832 ;
  assign n12834 = n12831 & ~n12833 ;
  assign n12835 = x72 & ~n1259 ;
  assign n12836 = ~n8581 & n12835 ;
  assign n12837 = n12834 | n12836 ;
  assign n12838 = ~n4904 & n12837 ;
  assign n12839 = x110 | n12838 ;
  assign n12840 = n11413 & n12839 ;
  assign n12841 = ~n1649 & n12831 ;
  assign n12842 = x72 | n12841 ;
  assign n12843 = n4905 | n11413 ;
  assign n12844 = n12842 & ~n12843 ;
  assign n12845 = x39 | n12844 ;
  assign n12846 = n12840 | n12845 ;
  assign n12847 = ~n12813 & n12846 ;
  assign n12848 = ( ~n6785 & n12808 ) | ( ~n6785 & n12847 ) | ( n12808 & n12847 ) ;
  assign n12849 = ~n12817 & n12848 ;
  assign n12850 = n12807 | n12849 ;
  assign n12851 = x125 | n12396 ;
  assign n12852 = ( x133 & ~n12397 ) | ( x133 & n12851 ) | ( ~n12397 & n12851 ) ;
  assign n12853 = ( x125 & ~n12397 ) | ( x125 & n12852 ) | ( ~n12397 & n12852 ) ;
  assign n12854 = n12403 | n12853 ;
  assign n12855 = x172 & n12409 ;
  assign n12856 = ~x152 & n12525 ;
  assign n12857 = n12855 | n12856 ;
  assign n12858 = x232 & n12857 ;
  assign n12859 = n12854 & ~n12858 ;
  assign n12860 = x87 | n12859 ;
  assign n12861 = x87 & n5924 ;
  assign n12862 = x162 & n12861 ;
  assign n12863 = n6785 & ~n12862 ;
  assign n12864 = n12860 & n12863 ;
  assign n12865 = x152 | n4713 ;
  assign n12866 = n12472 & n12865 ;
  assign n12867 = ~x152 & n12554 ;
  assign n12868 = x197 | n12867 ;
  assign n12869 = n12866 | n12868 ;
  assign n12870 = n4713 & n12472 ;
  assign n12871 = n12519 & ~n12870 ;
  assign n12872 = n12563 & ~n12871 ;
  assign n12873 = ~x152 & x197 ;
  assign n12874 = ~n12872 & n12873 ;
  assign n12875 = n12869 & ~n12874 ;
  assign n12876 = n12855 | n12875 ;
  assign n12877 = n12409 | n12479 ;
  assign n12878 = n12472 | n12877 ;
  assign n12879 = x152 & x197 ;
  assign n12880 = ( x172 & n12878 ) | ( x172 & ~n12879 ) | ( n12878 & ~n12879 ) ;
  assign n12881 = n4713 & ~n12472 ;
  assign n12882 = n12485 & ~n12881 ;
  assign n12883 = ( x172 & n12879 ) | ( x172 & ~n12882 ) | ( n12879 & ~n12882 ) ;
  assign n12884 = ~n12880 & n12883 ;
  assign n12885 = n12876 & ~n12884 ;
  assign n12886 = n8007 | n12885 ;
  assign n12887 = n4713 | n12470 ;
  assign n12888 = ~n12871 & n12887 ;
  assign n12889 = x152 | n12855 ;
  assign n12890 = n12888 | n12889 ;
  assign n12891 = x197 & n12890 ;
  assign n12892 = n12507 & ~n12881 ;
  assign n12893 = ( ~x152 & x172 ) | ( ~x152 & n12892 ) | ( x172 & n12892 ) ;
  assign n12894 = n12514 & ~n12881 ;
  assign n12895 = ( x152 & x172 ) | ( x152 & ~n12894 ) | ( x172 & ~n12894 ) ;
  assign n12896 = ~n12893 & n12895 ;
  assign n12897 = n12891 & ~n12896 ;
  assign n12898 = n12469 | n12562 ;
  assign n12899 = ~n12881 & n12898 ;
  assign n12900 = ( x152 & x172 ) | ( x152 & ~n12899 ) | ( x172 & ~n12899 ) ;
  assign n12901 = n12473 | n12536 ;
  assign n12902 = ( x152 & ~x172 ) | ( x152 & n12901 ) | ( ~x172 & n12901 ) ;
  assign n12903 = n12900 & ~n12902 ;
  assign n12904 = x197 | n12903 ;
  assign n12905 = n12542 & ~n12881 ;
  assign n12906 = ( x152 & x172 ) | ( x152 & n12905 ) | ( x172 & n12905 ) ;
  assign n12907 = n12520 | n12870 ;
  assign n12908 = ( ~x152 & x172 ) | ( ~x152 & n12907 ) | ( x172 & n12907 ) ;
  assign n12909 = n12906 | n12908 ;
  assign n12910 = ~n12904 & n12909 ;
  assign n12911 = n8002 & ~n12910 ;
  assign n12912 = ~n12897 & n12911 ;
  assign n12913 = n12886 & ~n12912 ;
  assign n12914 = x299 & ~n12913 ;
  assign n12915 = ( x145 & x174 ) | ( x145 & ~n12472 ) | ( x174 & ~n12472 ) ;
  assign n12916 = ( x145 & ~x174 ) | ( x145 & n12882 ) | ( ~x174 & n12882 ) ;
  assign n12917 = n12915 & ~n12916 ;
  assign n12918 = ( x145 & x174 ) | ( x145 & n12872 ) | ( x174 & n12872 ) ;
  assign n12919 = n12554 | n12870 ;
  assign n12920 = ( ~x145 & x174 ) | ( ~x145 & n12919 ) | ( x174 & n12919 ) ;
  assign n12921 = n12918 | n12920 ;
  assign n12922 = ~n12917 & n12921 ;
  assign n12923 = x193 | n12922 ;
  assign n12924 = ~x145 & n12479 ;
  assign n12925 = n12877 & ~n12924 ;
  assign n12926 = n12472 | n12925 ;
  assign n12927 = x174 & n12926 ;
  assign n12928 = n12409 | n12442 ;
  assign n12929 = x145 & n12928 ;
  assign n12930 = n12562 | n12929 ;
  assign n12931 = ~x174 & n12930 ;
  assign n12932 = ~n12881 & n12931 ;
  assign n12933 = x193 & ~n12932 ;
  assign n12934 = ~n12927 & n12933 ;
  assign n12935 = n12923 & ~n12934 ;
  assign n12936 = n8013 | n12935 ;
  assign n12937 = ( x145 & x193 ) | ( x145 & ~n12901 ) | ( x193 & ~n12901 ) ;
  assign n12938 = ( x145 & ~x193 ) | ( x145 & n12892 ) | ( ~x193 & n12892 ) ;
  assign n12939 = n12937 & ~n12938 ;
  assign n12940 = x174 & ~n12939 ;
  assign n12941 = ( x145 & x193 ) | ( x145 & n12894 ) | ( x193 & n12894 ) ;
  assign n12942 = ( ~x145 & x193 ) | ( ~x145 & n12905 ) | ( x193 & n12905 ) ;
  assign n12943 = n12941 | n12942 ;
  assign n12944 = n12940 & n12943 ;
  assign n12945 = x193 & n12409 ;
  assign n12946 = x145 & ~n12945 ;
  assign n12947 = ~n12888 & n12946 ;
  assign n12948 = x174 | n12947 ;
  assign n12949 = ( x145 & x193 ) | ( x145 & n12899 ) | ( x193 & n12899 ) ;
  assign n12950 = ( x145 & ~x193 ) | ( x145 & n12907 ) | ( ~x193 & n12907 ) ;
  assign n12951 = n12949 | n12950 ;
  assign n12952 = ~n12948 & n12951 ;
  assign n12953 = n8017 & ~n12952 ;
  assign n12954 = ~n12944 & n12953 ;
  assign n12955 = n12936 & ~n12954 ;
  assign n12956 = x38 | n12955 ;
  assign n12957 = ~n12914 & n12956 ;
  assign n12958 = n5788 & ~n12957 ;
  assign n12959 = x299 | n6448 ;
  assign n12960 = x299 & ~n6433 ;
  assign n12961 = n12959 & ~n12960 ;
  assign n12962 = ~n1868 & n12961 ;
  assign n12963 = x232 | n12962 ;
  assign n12964 = x39 & n12963 ;
  assign n12965 = n6448 | n12744 ;
  assign n12966 = ~n1868 & n12965 ;
  assign n12967 = ( x174 & x193 ) | ( x174 & n12966 ) | ( x193 & n12966 ) ;
  assign n12968 = ( x224 & ~n4989 ) | ( x224 & n12644 ) | ( ~n4989 & n12644 ) ;
  assign n12969 = ~n1868 & n4713 ;
  assign n12970 = n4713 | n12641 ;
  assign n12971 = ~n12969 & n12970 ;
  assign n12972 = ( x224 & n4989 ) | ( x224 & ~n12971 ) | ( n4989 & ~n12971 ) ;
  assign n12973 = ~n12968 & n12972 ;
  assign n12974 = n12637 | n12973 ;
  assign n12975 = ( ~x174 & x193 ) | ( ~x174 & n12974 ) | ( x193 & n12974 ) ;
  assign n12976 = n12967 | n12975 ;
  assign n12977 = x180 & n12976 ;
  assign n12978 = n4713 | n12600 ;
  assign n12979 = ~n12969 & n12978 ;
  assign n12980 = n6448 & n12979 ;
  assign n12981 = n12599 | n12614 ;
  assign n12982 = x224 & n12981 ;
  assign n12983 = n4989 & ~n12982 ;
  assign n12984 = n12407 | n12983 ;
  assign n12985 = ~n12980 & n12984 ;
  assign n12986 = ( x174 & x193 ) | ( x174 & ~n12985 ) | ( x193 & ~n12985 ) ;
  assign n12987 = n12602 | n12614 ;
  assign n12988 = ~n12409 & n12987 ;
  assign n12989 = x224 & n12988 ;
  assign n12990 = n4989 & ~n12989 ;
  assign n12991 = n12604 & ~n12969 ;
  assign n12992 = n6448 & n12991 ;
  assign n12993 = n12990 & ~n12992 ;
  assign n12994 = n12409 | n12993 ;
  assign n12995 = ( x174 & ~x193 ) | ( x174 & n12994 ) | ( ~x193 & n12994 ) ;
  assign n12996 = n12986 & ~n12995 ;
  assign n12997 = n12977 & ~n12996 ;
  assign n12998 = ~n1868 & n6448 ;
  assign n12999 = ( x174 & n12945 ) | ( x174 & n12998 ) | ( n12945 & n12998 ) ;
  assign n13000 = n6448 | n12407 ;
  assign n13001 = ~n12971 & n13000 ;
  assign n13002 = ( ~x174 & n12945 ) | ( ~x174 & n13001 ) | ( n12945 & n13001 ) ;
  assign n13003 = n12999 | n13002 ;
  assign n13004 = ~x180 & n13003 ;
  assign n13005 = x299 | n13004 ;
  assign n13006 = n12997 | n13005 ;
  assign n13007 = n6433 | n12857 ;
  assign n13008 = x51 & ~x172 ;
  assign n13009 = ( x152 & n12991 ) | ( x152 & n13008 ) | ( n12991 & n13008 ) ;
  assign n13010 = ( ~x152 & n12979 ) | ( ~x152 & n13008 ) | ( n12979 & n13008 ) ;
  assign n13011 = n13009 | n13010 ;
  assign n13012 = ~x216 & n13011 ;
  assign n13013 = n5005 & n13012 ;
  assign n13014 = n13007 & ~n13013 ;
  assign n13015 = n7610 & ~n13014 ;
  assign n13016 = ~n12407 & n12981 ;
  assign n13017 = ( x152 & x172 ) | ( x152 & ~n13016 ) | ( x172 & ~n13016 ) ;
  assign n13018 = ( x152 & ~x172 ) | ( x152 & n12988 ) | ( ~x172 & n12988 ) ;
  assign n13019 = n13017 & ~n13018 ;
  assign n13020 = x216 & ~n13019 ;
  assign n13021 = ( x152 & x172 ) | ( x152 & n12756 ) | ( x172 & n12756 ) ;
  assign n13022 = ( ~x152 & x172 ) | ( ~x152 & n12644 ) | ( x172 & n12644 ) ;
  assign n13023 = n13021 | n13022 ;
  assign n13024 = n13020 & n13023 ;
  assign n13025 = n5005 & ~n13024 ;
  assign n13026 = ~n13012 & n13025 ;
  assign n13027 = ~n5005 & n12857 ;
  assign n13028 = n7581 & ~n13027 ;
  assign n13029 = ~n13026 & n13028 ;
  assign n13030 = n13015 | n13029 ;
  assign n13031 = n13006 & ~n13030 ;
  assign n13032 = x232 & ~n13031 ;
  assign n13033 = n12964 & ~n13032 ;
  assign n13034 = x232 | n12472 ;
  assign n13035 = ~x39 & n13034 ;
  assign n13036 = x38 | n13035 ;
  assign n13037 = n13033 | n13036 ;
  assign n13038 = x299 & ~n12857 ;
  assign n13039 = ~x174 & n12525 ;
  assign n13040 = n12945 | n13039 ;
  assign n13041 = ( x232 & n7916 ) | ( x232 & n13040 ) | ( n7916 & n13040 ) ;
  assign n13042 = ~n13038 & n13041 ;
  assign n13043 = x38 & ~n13042 ;
  assign n13044 = x100 | n13043 ;
  assign n13045 = n13037 & ~n13044 ;
  assign n13046 = ~n12958 & n13045 ;
  assign n13047 = x100 & n13042 ;
  assign n13048 = n2043 | n13047 ;
  assign n13049 = n13046 | n13048 ;
  assign n13050 = n12682 & ~n13042 ;
  assign n13051 = x140 & ~x299 ;
  assign n13052 = x162 & x299 ;
  assign n13053 = n13051 | n13052 ;
  assign n13054 = n5924 & n13053 ;
  assign n13055 = x87 & ~n13054 ;
  assign n13056 = n12853 & ~n13055 ;
  assign n13057 = ~n13050 & n13056 ;
  assign n13058 = n13049 & n13057 ;
  assign n13059 = x145 | n12462 ;
  assign n13060 = n12693 | n13059 ;
  assign n13061 = n12462 | n12536 ;
  assign n13062 = x145 & ~n13061 ;
  assign n13063 = ~x51 & n13062 ;
  assign n13064 = x174 | n13063 ;
  assign n13065 = n13060 & ~n13064 ;
  assign n13066 = ~x145 & n12460 ;
  assign n13067 = n4713 & n12460 ;
  assign n13068 = n12407 | n13067 ;
  assign n13069 = n12459 | n13068 ;
  assign n13070 = n13066 | n13069 ;
  assign n13071 = x174 & n13070 ;
  assign n13072 = x193 | n13071 ;
  assign n13073 = n13065 | n13072 ;
  assign n13074 = ~n12478 & n12511 ;
  assign n13075 = n12462 | n13074 ;
  assign n13076 = x145 | n13075 ;
  assign n13077 = x174 | n13062 ;
  assign n13078 = n13076 & ~n13077 ;
  assign n13079 = n1864 | n13070 ;
  assign n13080 = n12462 | n12700 ;
  assign n13081 = x174 & n13080 ;
  assign n13082 = n13079 & n13081 ;
  assign n13083 = x193 & ~n13082 ;
  assign n13084 = ~n13078 & n13083 ;
  assign n13085 = n8013 | n13084 ;
  assign n13086 = n13073 & ~n13085 ;
  assign n13087 = n12409 | n12462 ;
  assign n13088 = x174 | n12924 ;
  assign n13089 = x145 & ~n12402 ;
  assign n13090 = n13088 & ~n13089 ;
  assign n13091 = n13087 | n13090 ;
  assign n13092 = n12462 | n12718 ;
  assign n13093 = x174 & ~n13092 ;
  assign n13094 = n13091 & ~n13093 ;
  assign n13095 = x193 | n13094 ;
  assign n13096 = x145 & ~n12525 ;
  assign n13097 = ~x145 & x174 ;
  assign n13098 = ~n12716 & n13097 ;
  assign n13099 = n13096 | n13098 ;
  assign n13100 = n13088 & ~n13099 ;
  assign n13101 = x193 & ~n12462 ;
  assign n13102 = ~n13100 & n13101 ;
  assign n13103 = n8017 & ~n13102 ;
  assign n13104 = n13095 & n13103 ;
  assign n13105 = n13086 | n13104 ;
  assign n13106 = ~x38 & n13105 ;
  assign n13107 = ~x152 & n12693 ;
  assign n13108 = n12461 & n12865 ;
  assign n13109 = x172 | n13108 ;
  assign n13110 = n13107 | n13109 ;
  assign n13111 = ( x152 & x172 ) | ( x152 & ~n13075 ) | ( x172 & ~n13075 ) ;
  assign n13112 = ( x152 & ~x172 ) | ( x152 & n13080 ) | ( ~x172 & n13080 ) ;
  assign n13113 = n13111 & ~n13112 ;
  assign n13114 = n13110 & ~n13113 ;
  assign n13115 = x197 | n13114 ;
  assign n13116 = ~x152 & n13061 ;
  assign n13117 = ~x172 & n12409 ;
  assign n13118 = x197 & ~n13117 ;
  assign n13119 = n12462 | n12528 ;
  assign n13120 = ( x152 & ~x172 ) | ( x152 & n13119 ) | ( ~x172 & n13119 ) ;
  assign n13121 = ( x152 & x172 ) | ( x152 & n13069 ) | ( x172 & n13069 ) ;
  assign n13122 = n13120 & n13121 ;
  assign n13123 = n13118 & ~n13122 ;
  assign n13124 = ~n13116 & n13123 ;
  assign n13125 = x299 & ~n8007 ;
  assign n13126 = ~n13124 & n13125 ;
  assign n13127 = n13115 & n13126 ;
  assign n13128 = n12462 | n12479 ;
  assign n13129 = x152 | n13128 ;
  assign n13130 = n12409 | n13129 ;
  assign n13131 = x152 & ~n13092 ;
  assign n13132 = x172 | n13131 ;
  assign n13133 = n13130 & ~n13132 ;
  assign n13134 = n12462 | n12716 ;
  assign n13135 = x152 & ~n13134 ;
  assign n13136 = x172 & ~n13135 ;
  assign n13137 = n13129 & n13136 ;
  assign n13138 = x197 | n13137 ;
  assign n13139 = n13133 | n13138 ;
  assign n13140 = x172 | n12856 ;
  assign n13141 = n12463 & ~n13140 ;
  assign n13142 = x152 & n12525 ;
  assign n13143 = n12462 | n13142 ;
  assign n13144 = x172 & n13143 ;
  assign n13145 = x197 & ~n13144 ;
  assign n13146 = ~n13141 & n13145 ;
  assign n13147 = x299 & n8002 ;
  assign n13148 = ~n13146 & n13147 ;
  assign n13149 = n13139 & n13148 ;
  assign n13150 = n13127 | n13149 ;
  assign n13151 = n13106 | n13150 ;
  assign n13152 = n5788 & n13151 ;
  assign n13153 = n12430 & n13044 ;
  assign n13154 = n12403 & ~n12857 ;
  assign n13155 = n7296 | n13154 ;
  assign n13156 = ~n12600 & n12865 ;
  assign n13157 = x152 | n12604 ;
  assign n13158 = ~n13156 & n13157 ;
  assign n13159 = x172 | n13158 ;
  assign n13160 = n7296 & n13159 ;
  assign n13161 = ( x152 & x172 ) | ( x152 & ~n12607 ) | ( x172 & ~n12607 ) ;
  assign n13162 = ( x152 & ~x172 ) | ( x152 & n12649 ) | ( ~x172 & n12649 ) ;
  assign n13163 = n13161 & ~n13162 ;
  assign n13164 = n13160 & ~n13163 ;
  assign n13165 = n7610 & ~n13164 ;
  assign n13166 = n12616 & ~n12889 ;
  assign n13167 = x152 & ~n12855 ;
  assign n13168 = n12619 & n13167 ;
  assign n13169 = n7296 & ~n13168 ;
  assign n13170 = ~n13166 & n13169 ;
  assign n13171 = n7581 & ~n13170 ;
  assign n13172 = n13165 | n13171 ;
  assign n13173 = n13155 & n13172 ;
  assign n13174 = n4713 & n12402 ;
  assign n13175 = n7285 | n13174 ;
  assign n13176 = n12648 | n13175 ;
  assign n13177 = n7285 & ~n12601 ;
  assign n13178 = ~n8715 & n13177 ;
  assign n13179 = n13176 & ~n13178 ;
  assign n13180 = ( x174 & x180 ) | ( x174 & n13179 ) | ( x180 & n13179 ) ;
  assign n13181 = ~x51 & n12619 ;
  assign n13182 = n4713 | n13181 ;
  assign n13183 = ( n7285 & n12403 ) | ( n7285 & ~n12600 ) | ( n12403 & ~n12600 ) ;
  assign n13184 = n13182 & n13183 ;
  assign n13185 = ( ~x174 & x180 ) | ( ~x174 & n13184 ) | ( x180 & n13184 ) ;
  assign n13186 = n13180 & n13185 ;
  assign n13187 = x193 & ~n13186 ;
  assign n13188 = ~n12409 & n13183 ;
  assign n13189 = ( x174 & x180 ) | ( x174 & ~n13188 ) | ( x180 & ~n13188 ) ;
  assign n13190 = n7285 & n12607 ;
  assign n13191 = n13176 & ~n13190 ;
  assign n13192 = ( x174 & ~x180 ) | ( x174 & n13191 ) | ( ~x180 & n13191 ) ;
  assign n13193 = ~n13189 & n13192 ;
  assign n13194 = n13187 & ~n13193 ;
  assign n13195 = n7285 & n12605 ;
  assign n13196 = x51 | n13175 ;
  assign n13197 = ~n13195 & n13196 ;
  assign n13198 = x180 & ~n12615 ;
  assign n13199 = x174 | n13198 ;
  assign n13200 = n13197 & ~n13199 ;
  assign n13201 = x180 & ~n12619 ;
  assign n13202 = x174 & n13183 ;
  assign n13203 = ~n13201 & n13202 ;
  assign n13204 = x193 | n13203 ;
  assign n13205 = n13200 | n13204 ;
  assign n13206 = ~x299 & n13205 ;
  assign n13207 = ~n13194 & n13206 ;
  assign n13208 = n13173 | n13207 ;
  assign n13209 = x232 & n13208 ;
  assign n13210 = ~x299 & n13183 ;
  assign n13211 = n7296 & ~n12599 ;
  assign n13212 = n12403 | n13211 ;
  assign n13213 = x299 & n13212 ;
  assign n13214 = n13210 | n13213 ;
  assign n13215 = ~x232 & n13214 ;
  assign n13216 = x39 & ~n13215 ;
  assign n13217 = ~n13209 & n13216 ;
  assign n13218 = ~x232 & n12461 ;
  assign n13219 = x39 | n13218 ;
  assign n13220 = ~x38 & n13219 ;
  assign n13221 = ~n13217 & n13220 ;
  assign n13222 = n13153 | n13221 ;
  assign n13223 = n13152 | n13222 ;
  assign n13224 = n12678 | n13047 ;
  assign n13225 = n13223 & ~n13224 ;
  assign n13226 = n12683 & ~n13042 ;
  assign n13227 = n12853 | n13055 ;
  assign n13228 = n13226 | n13227 ;
  assign n13229 = n13225 | n13228 ;
  assign n13230 = ~n6785 & n13229 ;
  assign n13231 = ~n13058 & n13230 ;
  assign n13232 = n12864 | n13231 ;
  assign n13233 = x189 & ~n12882 ;
  assign n13234 = x189 | n12872 ;
  assign n13235 = ~x178 & n13234 ;
  assign n13236 = ~n13233 & n13235 ;
  assign n13237 = x189 & n12894 ;
  assign n13238 = ~x189 & n12888 ;
  assign n13239 = x178 & ~n13238 ;
  assign n13240 = ~n13237 & n13239 ;
  assign n13241 = ( x178 & n13236 ) | ( x178 & ~n13240 ) | ( n13236 & ~n13240 ) ;
  assign n13242 = x181 & n13241 ;
  assign n13243 = ~x189 & n12919 ;
  assign n13244 = x189 & n12472 ;
  assign n13245 = x178 | n13244 ;
  assign n13246 = n12409 | n13245 ;
  assign n13247 = n13243 | n13246 ;
  assign n13248 = ~x181 & n13247 ;
  assign n13249 = n12919 | n13245 ;
  assign n13250 = n13248 & n13249 ;
  assign n13251 = ( ~x178 & x189 ) | ( ~x178 & n12905 ) | ( x189 & n12905 ) ;
  assign n13252 = ( x178 & x189 ) | ( x178 & ~n12907 ) | ( x189 & ~n12907 ) ;
  assign n13253 = ~n13251 & n13252 ;
  assign n13254 = n13250 & ~n13253 ;
  assign n13255 = n9932 | n13254 ;
  assign n13256 = n13242 | n13255 ;
  assign n13257 = ( x153 & x157 ) | ( x153 & ~n12894 ) | ( x157 & ~n12894 ) ;
  assign n13258 = ( x153 & ~x157 ) | ( x153 & n12892 ) | ( ~x157 & n12892 ) ;
  assign n13259 = n13257 & ~n13258 ;
  assign n13260 = ( x153 & x157 ) | ( x153 & n12878 ) | ( x157 & n12878 ) ;
  assign n13261 = ( ~x153 & x157 ) | ( ~x153 & n12882 ) | ( x157 & n12882 ) ;
  assign n13262 = n13260 | n13261 ;
  assign n13263 = ~n13259 & n13262 ;
  assign n13264 = x166 & ~n13263 ;
  assign n13265 = x153 & n12409 ;
  assign n13266 = x166 | n13265 ;
  assign n13267 = ( x157 & n12888 ) | ( x157 & n13266 ) | ( n12888 & n13266 ) ;
  assign n13268 = ( ~x157 & n12872 ) | ( ~x157 & n13266 ) | ( n12872 & n13266 ) ;
  assign n13269 = n13267 | n13268 ;
  assign n13270 = ~n13264 & n13269 ;
  assign n13271 = n7975 & ~n13270 ;
  assign n13272 = x166 & n12901 ;
  assign n13273 = x153 & x166 ;
  assign n13274 = ( x153 & ~n12899 ) | ( x153 & n13273 ) | ( ~n12899 & n13273 ) ;
  assign n13275 = ~n13272 & n13274 ;
  assign n13276 = ( x153 & x166 ) | ( x153 & n12905 ) | ( x166 & n12905 ) ;
  assign n13277 = ( x153 & ~x166 ) | ( x153 & n12907 ) | ( ~x166 & n12907 ) ;
  assign n13278 = n13276 | n13277 ;
  assign n13279 = ~n13275 & n13278 ;
  assign n13280 = x157 & ~n13279 ;
  assign n13281 = x157 | n13265 ;
  assign n13282 = ( x166 & n12472 ) | ( x166 & n13281 ) | ( n12472 & n13281 ) ;
  assign n13283 = ( ~x166 & n12919 ) | ( ~x166 & n13281 ) | ( n12919 & n13281 ) ;
  assign n13284 = n13282 | n13283 ;
  assign n13285 = ~n13280 & n13284 ;
  assign n13286 = n7974 & ~n13285 ;
  assign n13287 = x189 | n13087 ;
  assign n13288 = n12892 & n13287 ;
  assign n13289 = n13239 & ~n13288 ;
  assign n13290 = x189 & ~n12878 ;
  assign n13291 = n12409 | n13234 ;
  assign n13292 = ~n13290 & n13291 ;
  assign n13293 = x178 | n13292 ;
  assign n13294 = x181 & n13293 ;
  assign n13295 = ~n13289 & n13294 ;
  assign n13296 = ( ~x178 & x189 ) | ( ~x178 & n12901 ) | ( x189 & n12901 ) ;
  assign n13297 = ( x178 & x189 ) | ( x178 & ~n12899 ) | ( x189 & ~n12899 ) ;
  assign n13298 = ~n13296 & n13297 ;
  assign n13299 = n13248 & ~n13298 ;
  assign n13300 = n9920 & ~n13299 ;
  assign n13301 = ~n13295 & n13300 ;
  assign n13302 = n13286 | n13301 ;
  assign n13303 = n13271 | n13302 ;
  assign n13304 = n13256 & ~n13303 ;
  assign n13305 = x232 & ~n13304 ;
  assign n13306 = n13035 & ~n13305 ;
  assign n13307 = x126 | n12399 ;
  assign n13308 = x126 & n12399 ;
  assign n13309 = n13307 & ~n13308 ;
  assign n13310 = n12395 & ~n13309 ;
  assign n13311 = x51 | n12525 ;
  assign n13312 = n8466 & n12402 ;
  assign n13313 = x51 | n13312 ;
  assign n13314 = ~n13265 & n13313 ;
  assign n13315 = n13311 & ~n13314 ;
  assign n13316 = ~x160 & n7296 ;
  assign n13317 = ( ~n5005 & n13315 ) | ( ~n5005 & n13316 ) | ( n13315 & n13316 ) ;
  assign n13318 = x299 & ~n13317 ;
  assign n13319 = ( x153 & x166 ) | ( x153 & ~n12756 ) | ( x166 & ~n12756 ) ;
  assign n13320 = ( ~x153 & x166 ) | ( ~x153 & n12644 ) | ( x166 & n12644 ) ;
  assign n13321 = ~n13319 & n13320 ;
  assign n13322 = x160 & ~n13321 ;
  assign n13323 = ( x153 & ~x166 ) | ( x153 & n12988 ) | ( ~x166 & n12988 ) ;
  assign n13324 = ( x153 & x166 ) | ( x153 & n13016 ) | ( x166 & n13016 ) ;
  assign n13325 = n13323 & n13324 ;
  assign n13326 = n13322 & ~n13325 ;
  assign n13327 = ( ~x216 & n5005 ) | ( ~x216 & n13326 ) | ( n5005 & n13326 ) ;
  assign n13328 = x51 & ~x153 ;
  assign n13329 = ( x166 & n12991 ) | ( x166 & n13328 ) | ( n12991 & n13328 ) ;
  assign n13330 = ( ~x166 & n12979 ) | ( ~x166 & n13328 ) | ( n12979 & n13328 ) ;
  assign n13331 = n13329 | n13330 ;
  assign n13332 = ( x216 & n5005 ) | ( x216 & ~n13331 ) | ( n5005 & ~n13331 ) ;
  assign n13333 = n13327 & n13332 ;
  assign n13334 = n13318 & ~n13333 ;
  assign n13335 = ( x182 & x189 ) | ( x182 & n12998 ) | ( x189 & n12998 ) ;
  assign n13336 = ( x182 & ~x189 ) | ( x182 & n13001 ) | ( ~x189 & n13001 ) ;
  assign n13337 = n13335 | n13336 ;
  assign n13338 = n12409 | n13337 ;
  assign n13339 = ( ~x182 & x189 ) | ( ~x182 & n12994 ) | ( x189 & n12994 ) ;
  assign n13340 = ( x182 & x189 ) | ( x182 & ~n12985 ) | ( x189 & ~n12985 ) ;
  assign n13341 = ~n13339 & n13340 ;
  assign n13342 = n13338 & ~n13341 ;
  assign n13343 = n9920 & ~n13342 ;
  assign n13344 = ( ~x182 & x189 ) | ( ~x182 & n12966 ) | ( x189 & n12966 ) ;
  assign n13345 = ( x182 & x189 ) | ( x182 & ~n12974 ) | ( x189 & ~n12974 ) ;
  assign n13346 = ~n13344 & n13345 ;
  assign n13347 = n13337 & ~n13346 ;
  assign n13348 = n9932 | n13347 ;
  assign n13349 = ~n13343 & n13348 ;
  assign n13350 = ~n13334 & n13349 ;
  assign n13351 = x232 & ~n13350 ;
  assign n13352 = n12964 & ~n13351 ;
  assign n13353 = n13310 & ~n13352 ;
  assign n13354 = ~n13306 & n13353 ;
  assign n13355 = ~x166 & n12693 ;
  assign n13356 = n8466 & n12461 ;
  assign n13357 = x153 | n13356 ;
  assign n13358 = n13355 | n13357 ;
  assign n13359 = ( ~x153 & x166 ) | ( ~x153 & n13080 ) | ( x166 & n13080 ) ;
  assign n13360 = ( x153 & x166 ) | ( x153 & ~n13075 ) | ( x166 & ~n13075 ) ;
  assign n13361 = ~n13359 & n13360 ;
  assign n13362 = n13358 & ~n13361 ;
  assign n13363 = x157 | n13362 ;
  assign n13364 = x51 & ~n8466 ;
  assign n13365 = x166 & n13092 ;
  assign n13366 = n13364 | n13365 ;
  assign n13367 = ~x153 & n13366 ;
  assign n13368 = ~x166 & n13128 ;
  assign n13369 = n13134 & n13273 ;
  assign n13370 = x157 & ~n13369 ;
  assign n13371 = ~n13368 & n13370 ;
  assign n13372 = ~n13367 & n13371 ;
  assign n13373 = n7974 & ~n13372 ;
  assign n13374 = n13363 & n13373 ;
  assign n13375 = n8477 & n12461 ;
  assign n13376 = ~x189 & n12693 ;
  assign n13377 = n13375 | n13376 ;
  assign n13378 = ~x178 & n13377 ;
  assign n13379 = x189 & ~n13092 ;
  assign n13380 = x178 & n13287 ;
  assign n13381 = x189 | n13128 ;
  assign n13382 = x178 & n13381 ;
  assign n13383 = n13380 | n13382 ;
  assign n13384 = ~n13379 & n13383 ;
  assign n13385 = x181 | n13384 ;
  assign n13386 = n13378 | n13385 ;
  assign n13387 = n12536 | n13287 ;
  assign n13388 = x189 & ~n13069 ;
  assign n13389 = x178 | n13388 ;
  assign n13390 = n13387 & ~n13389 ;
  assign n13391 = x189 & ~n12463 ;
  assign n13392 = n13380 & ~n13391 ;
  assign n13393 = x181 & ~n13392 ;
  assign n13394 = ~n13390 & n13393 ;
  assign n13395 = n9932 | n13394 ;
  assign n13396 = n13386 & ~n13395 ;
  assign n13397 = x189 & ~n13134 ;
  assign n13398 = n13382 & ~n13397 ;
  assign n13399 = x181 | n13398 ;
  assign n13400 = ( x178 & x189 ) | ( x178 & ~n13080 ) | ( x189 & ~n13080 ) ;
  assign n13401 = ( ~x178 & x189 ) | ( ~x178 & n13075 ) | ( x189 & n13075 ) ;
  assign n13402 = ~n13400 & n13401 ;
  assign n13403 = n13399 | n13402 ;
  assign n13404 = x178 & n9923 ;
  assign n13405 = n12524 & n13404 ;
  assign n13406 = x181 & ~n13405 ;
  assign n13407 = ~n12462 & n13406 ;
  assign n13408 = ( x178 & x189 ) | ( x178 & ~n12528 ) | ( x189 & ~n12528 ) ;
  assign n13409 = ( ~x178 & x189 ) | ( ~x178 & n12536 ) | ( x189 & n12536 ) ;
  assign n13410 = ~n13408 & n13409 ;
  assign n13411 = n13407 & ~n13410 ;
  assign n13412 = n9920 & ~n13411 ;
  assign n13413 = n13403 & n13412 ;
  assign n13414 = ~x166 & n13061 ;
  assign n13415 = x166 & n13069 ;
  assign n13416 = n13364 | n13415 ;
  assign n13417 = ~x153 & n13416 ;
  assign n13418 = n13119 & n13273 ;
  assign n13419 = x157 | n13418 ;
  assign n13420 = n13417 | n13419 ;
  assign n13421 = n13414 | n13420 ;
  assign n13422 = x153 | n13315 ;
  assign n13423 = n12463 & ~n13422 ;
  assign n13424 = x166 & n12525 ;
  assign n13425 = n12462 | n13424 ;
  assign n13426 = x153 & n13425 ;
  assign n13427 = x157 & ~n13426 ;
  assign n13428 = ~n13423 & n13427 ;
  assign n13429 = n7975 & ~n13428 ;
  assign n13430 = n13421 & n13429 ;
  assign n13431 = n13413 | n13430 ;
  assign n13432 = n13396 | n13431 ;
  assign n13433 = n13374 | n13432 ;
  assign n13434 = x232 & n13433 ;
  assign n13435 = n13219 | n13434 ;
  assign n13436 = n8466 & ~n12600 ;
  assign n13437 = x166 | n12604 ;
  assign n13438 = ~n13436 & n13437 ;
  assign n13439 = x153 | n13438 ;
  assign n13440 = ( ~x153 & x166 ) | ( ~x153 & n12649 ) | ( x166 & n12649 ) ;
  assign n13441 = ( x153 & x166 ) | ( x153 & ~n12607 ) | ( x166 & ~n12607 ) ;
  assign n13442 = ~n13440 & n13441 ;
  assign n13443 = n13439 & ~n13442 ;
  assign n13444 = x160 | n13443 ;
  assign n13445 = x160 & ~n13265 ;
  assign n13446 = ( x166 & n12616 ) | ( x166 & n13445 ) | ( n12616 & n13445 ) ;
  assign n13447 = ( ~x166 & n12619 ) | ( ~x166 & n13445 ) | ( n12619 & n13445 ) ;
  assign n13448 = n13446 & n13447 ;
  assign n13449 = n7296 & ~n13448 ;
  assign n13450 = n13444 & n13449 ;
  assign n13451 = n7296 | n13314 ;
  assign n13452 = x299 & n13451 ;
  assign n13453 = ~n13450 & n13452 ;
  assign n13454 = x182 & ~n12619 ;
  assign n13455 = x189 & n13183 ;
  assign n13456 = ~n13454 & n13455 ;
  assign n13457 = x182 & ~n12615 ;
  assign n13458 = x189 | n13457 ;
  assign n13459 = n13197 & ~n13458 ;
  assign n13460 = n13456 | n13459 ;
  assign n13461 = ~n9932 & n13460 ;
  assign n13462 = ( x182 & x189 ) | ( x182 & ~n13188 ) | ( x189 & ~n13188 ) ;
  assign n13463 = ( ~x182 & x189 ) | ( ~x182 & n13191 ) | ( x189 & n13191 ) ;
  assign n13464 = ~n13462 & n13463 ;
  assign n13465 = ( x182 & ~x189 ) | ( x182 & n13184 ) | ( ~x189 & n13184 ) ;
  assign n13466 = ( x182 & x189 ) | ( x182 & n13179 ) | ( x189 & n13179 ) ;
  assign n13467 = n13465 & n13466 ;
  assign n13468 = n13464 | n13467 ;
  assign n13469 = n9920 & n13468 ;
  assign n13470 = n13461 | n13469 ;
  assign n13471 = n13453 | n13470 ;
  assign n13472 = x232 & n13471 ;
  assign n13473 = n13216 & ~n13472 ;
  assign n13474 = n13310 | n13473 ;
  assign n13475 = n13435 & ~n13474 ;
  assign n13476 = n1975 | n13475 ;
  assign n13477 = n13354 | n13476 ;
  assign n13478 = x299 & ~n13315 ;
  assign n13479 = ~x189 & n12525 ;
  assign n13480 = x175 & n12409 ;
  assign n13481 = n13479 | n13480 ;
  assign n13482 = ( x232 & n7916 ) | ( x232 & n13481 ) | ( n7916 & n13481 ) ;
  assign n13483 = ~n13478 & n13482 ;
  assign n13484 = n1975 & n13483 ;
  assign n13485 = n1975 & ~n12403 ;
  assign n13486 = ~n13310 & n13485 ;
  assign n13487 = n2043 | n13486 ;
  assign n13488 = n13484 | n13487 ;
  assign n13489 = n13477 & ~n13488 ;
  assign n13490 = n12404 | n13310 ;
  assign n13491 = n12682 & ~n13483 ;
  assign n13492 = ~x150 & x299 ;
  assign n13493 = x185 | x299 ;
  assign n13494 = ~n13492 & n13493 ;
  assign n13495 = n12861 & n13494 ;
  assign n13496 = ( x87 & n13491 ) | ( x87 & ~n13495 ) | ( n13491 & ~n13495 ) ;
  assign n13497 = n13490 & n13496 ;
  assign n13498 = n6785 | n13497 ;
  assign n13499 = n13489 | n13498 ;
  assign n13500 = ( ~x87 & n6785 ) | ( ~x87 & n11826 ) | ( n6785 & n11826 ) ;
  assign n13501 = x232 & n13311 ;
  assign n13502 = n13310 & ~n13501 ;
  assign n13503 = ~x232 & n12403 ;
  assign n13504 = n13314 | n13503 ;
  assign n13505 = n13502 | n13504 ;
  assign n13506 = ( x87 & n6785 ) | ( x87 & ~n13505 ) | ( n6785 & ~n13505 ) ;
  assign n13507 = n13500 & n13506 ;
  assign n13508 = n13499 & ~n13507 ;
  assign n13509 = x57 & x59 ;
  assign n13510 = ~n2045 & n7117 ;
  assign n13511 = ~n2058 & n13510 ;
  assign n13512 = ( n2057 & n13509 ) | ( n2057 & ~n13511 ) | ( n13509 & ~n13511 ) ;
  assign n13513 = n2058 & ~n13510 ;
  assign n13514 = x129 & ~n5762 ;
  assign n13515 = x75 & n13514 ;
  assign n13516 = x92 | n13515 ;
  assign n13517 = n1976 & n7195 ;
  assign n13518 = n7117 & ~n13517 ;
  assign n13519 = ( x75 & n1924 ) | ( x75 & ~n13518 ) | ( n1924 & ~n13518 ) ;
  assign n13520 = x129 & ~n4660 ;
  assign n13521 = x38 & ~n13520 ;
  assign n13522 = n1304 | n1594 ;
  assign n13523 = x250 & ~n5925 ;
  assign n13524 = n8246 & n13523 ;
  assign n13525 = n1421 & ~n1429 ;
  assign n13526 = n1243 | n13525 ;
  assign n13527 = ~n1439 & n13526 ;
  assign n13528 = n1350 | n13527 ;
  assign n13529 = ~n1443 & n13528 ;
  assign n13530 = n1582 | n13529 ;
  assign n13531 = ~n1584 & n13530 ;
  assign n13532 = x86 | n13531 ;
  assign n13533 = ~n1347 & n13532 ;
  assign n13534 = x97 | n13533 ;
  assign n13535 = ~n1337 & n13534 ;
  assign n13536 = x108 | n13535 ;
  assign n13537 = ~n1334 & n13536 ;
  assign n13538 = n1731 | n13537 ;
  assign n13539 = ~n1454 & n13538 ;
  assign n13540 = ( ~n1324 & n1325 ) | ( ~n1324 & n13539 ) | ( n1325 & n13539 ) ;
  assign n13541 = ( n4800 & ~n13524 ) | ( n4800 & n13540 ) | ( ~n13524 & n13540 ) ;
  assign n13542 = n1345 | n13533 ;
  assign n13543 = ~n1337 & n13542 ;
  assign n13544 = x108 | n13543 ;
  assign n13545 = ~n1334 & n13544 ;
  assign n13546 = n1731 | n13545 ;
  assign n13547 = ~n1454 & n13546 ;
  assign n13548 = ( ~n1324 & n1325 ) | ( ~n1324 & n13547 ) | ( n1325 & n13547 ) ;
  assign n13549 = ( n4800 & n13524 ) | ( n4800 & ~n13548 ) | ( n13524 & ~n13548 ) ;
  assign n13550 = ~n13541 & n13549 ;
  assign n13551 = ( x127 & n13524 ) | ( x127 & n13548 ) | ( n13524 & n13548 ) ;
  assign n13552 = ( ~x127 & n13524 ) | ( ~x127 & n13540 ) | ( n13524 & n13540 ) ;
  assign n13553 = n13551 | n13552 ;
  assign n13554 = ~n13550 & n13553 ;
  assign n13555 = n1315 | n13554 ;
  assign n13556 = ~n1310 & n13555 ;
  assign n13557 = n1278 | n13556 ;
  assign n13558 = ~n13522 & n13557 ;
  assign n13559 = x70 | n13558 ;
  assign n13560 = ~n1280 & n13559 ;
  assign n13561 = x51 | n13560 ;
  assign n13562 = ~n1465 & n13561 ;
  assign n13563 = n1539 | n13562 ;
  assign n13564 = ~n1301 & n13563 ;
  assign n13565 = n1492 | n13564 ;
  assign n13566 = ~n2135 & n13565 ;
  assign n13567 = x95 | n13566 ;
  assign n13568 = ~x39 & x129 ;
  assign n13569 = ~n1496 & n13568 ;
  assign n13570 = n13567 & n13569 ;
  assign n13571 = ( x38 & n1925 ) | ( x38 & n7117 ) | ( n1925 & n7117 ) ;
  assign n13572 = n13570 | n13571 ;
  assign n13573 = ~n13521 & n13572 ;
  assign n13574 = ( ~x75 & n1924 ) | ( ~x75 & n13573 ) | ( n1924 & n13573 ) ;
  assign n13575 = ~n13519 & n13574 ;
  assign n13576 = n13516 | n13575 ;
  assign n13577 = x92 & ~x129 ;
  assign n13578 = n11665 | n13577 ;
  assign n13579 = n13576 & ~n13578 ;
  assign n13580 = x54 & ~n2005 ;
  assign n13581 = n7117 & n13580 ;
  assign n13582 = x74 | n13581 ;
  assign n13583 = n13579 | n13582 ;
  assign n13584 = ~n5075 & n13514 ;
  assign n13585 = x74 & ~n13584 ;
  assign n13586 = x55 | n13585 ;
  assign n13587 = n13583 & ~n13586 ;
  assign n13588 = x55 & ~n2031 ;
  assign n13589 = n13514 & n13588 ;
  assign n13590 = n13587 | n13589 ;
  assign n13591 = ( x62 & ~n9450 ) | ( x62 & n13590 ) | ( ~n9450 & n13590 ) ;
  assign n13592 = ( n9450 & ~n13513 ) | ( n9450 & n13591 ) | ( ~n13513 & n13591 ) ;
  assign n13593 = ( ~x56 & n9450 ) | ( ~x56 & n13592 ) | ( n9450 & n13592 ) ;
  assign n13594 = ( n2057 & ~n13509 ) | ( n2057 & n13593 ) | ( ~n13509 & n13593 ) ;
  assign n13595 = ~n13512 & n13594 ;
  assign n13596 = n4656 | n5759 ;
  assign n13597 = x38 | n2140 ;
  assign n13598 = ~n4662 & n13597 ;
  assign n13599 = ~n4802 & n4811 ;
  assign n13600 = x87 | n13599 ;
  assign n13601 = n13598 | n13600 ;
  assign n13602 = ~n4816 & n13601 ;
  assign n13603 = n7119 & n8585 ;
  assign n13604 = ( n4800 & ~n7197 ) | ( n4800 & n13603 ) | ( ~n7197 & n13603 ) ;
  assign n13605 = ( x129 & n7197 ) | ( x129 & n13603 ) | ( n7197 & n13603 ) ;
  assign n13606 = ~n13604 & n13605 ;
  assign n13607 = ~n1868 & n13606 ;
  assign n13608 = n4817 | n13607 ;
  assign n13609 = n13602 | n13608 ;
  assign n13610 = n5766 | n5801 ;
  assign n13611 = n13609 & ~n13610 ;
  assign n13612 = n5073 | n13611 ;
  assign n13613 = ~n13596 & n13612 ;
  assign n13614 = x56 | n13613 ;
  assign n13615 = ~n4653 & n13614 ;
  assign n13616 = x62 | n13615 ;
  assign n13617 = ~n4826 & n13616 ;
  assign n13618 = n2057 | n13617 ;
  assign n13619 = ~n4649 & n13618 ;
  assign n13620 = ~x51 & n13214 ;
  assign n13621 = x232 | n13620 ;
  assign n13622 = n9138 & n13621 ;
  assign n13623 = x169 & ~n4713 ;
  assign n13624 = ~n7296 & n12524 ;
  assign n13625 = ~n13623 & n13624 ;
  assign n13626 = x299 & ~n13625 ;
  assign n13627 = ~x162 & n7296 ;
  assign n13628 = ( ~n12641 & n13623 ) | ( ~n12641 & n13627 ) | ( n13623 & n13627 ) ;
  assign n13629 = ( n1868 & n13623 ) | ( n1868 & ~n13627 ) | ( n13623 & ~n13627 ) ;
  assign n13630 = n13628 & ~n13629 ;
  assign n13631 = n13626 & ~n13630 ;
  assign n13632 = x162 & n7296 ;
  assign n13633 = ( x169 & n13181 ) | ( x169 & n13632 ) | ( n13181 & n13632 ) ;
  assign n13634 = x51 | n12605 ;
  assign n13635 = n12614 & ~n13634 ;
  assign n13636 = ( ~x169 & n13632 ) | ( ~x169 & n13635 ) | ( n13632 & n13635 ) ;
  assign n13637 = n13633 & n13636 ;
  assign n13638 = n13631 & ~n13637 ;
  assign n13639 = x191 | x299 ;
  assign n13640 = ~x51 & n13183 ;
  assign n13641 = x140 & ~n13182 ;
  assign n13642 = n13640 & ~n13641 ;
  assign n13643 = n13639 | n13642 ;
  assign n13644 = ~x51 & n13197 ;
  assign n13645 = x140 & ~n12614 ;
  assign n13646 = n13644 & ~n13645 ;
  assign n13647 = n7239 & ~n13646 ;
  assign n13648 = n13643 & ~n13647 ;
  assign n13649 = ~n13638 & n13648 ;
  assign n13650 = x232 & ~n13649 ;
  assign n13651 = n13622 & ~n13650 ;
  assign n13652 = n5924 & n7241 ;
  assign n13653 = n12524 & ~n13652 ;
  assign n13654 = ( x100 & ~n9306 ) | ( x100 & n13653 ) | ( ~n9306 & n13653 ) ;
  assign n13655 = n13651 | n13654 ;
  assign n13656 = n13311 & ~n13653 ;
  assign n13657 = x100 & n13656 ;
  assign n13658 = n2043 | n13657 ;
  assign n13659 = n12677 | n13658 ;
  assign n13660 = n13655 & ~n13659 ;
  assign n13661 = x87 & ~n7941 ;
  assign n13662 = n12682 & ~n13656 ;
  assign n13663 = n13661 | n13662 ;
  assign n13664 = n12404 & n13663 ;
  assign n13665 = x132 | n13307 ;
  assign n13666 = x130 & n13665 ;
  assign n13667 = x130 | n13665 ;
  assign n13668 = ~n13666 & n13667 ;
  assign n13669 = n12393 & ~n13668 ;
  assign n13670 = n13664 | n13669 ;
  assign n13671 = n13660 | n13670 ;
  assign n13672 = ( x38 & x100 ) | ( x38 & ~n13656 ) | ( x100 & ~n13656 ) ;
  assign n13673 = n12603 | n13623 ;
  assign n13674 = x169 & ~n12978 ;
  assign n13675 = n13673 & ~n13674 ;
  assign n13676 = x216 | n13675 ;
  assign n13677 = ~n12648 & n13016 ;
  assign n13678 = x162 & x216 ;
  assign n13679 = ( x169 & n13677 ) | ( x169 & ~n13678 ) | ( n13677 & ~n13678 ) ;
  assign n13680 = ~x51 & n12987 ;
  assign n13681 = ( x169 & n13678 ) | ( x169 & ~n13680 ) | ( n13678 & ~n13680 ) ;
  assign n13682 = ~n13679 & n13681 ;
  assign n13683 = n13676 & ~n13682 ;
  assign n13684 = n5005 & ~n13683 ;
  assign n13685 = x169 & n12525 ;
  assign n13686 = x51 | n13685 ;
  assign n13687 = ( ~n5005 & n13627 ) | ( ~n5005 & n13686 ) | ( n13627 & n13686 ) ;
  assign n13688 = n13684 | n13687 ;
  assign n13689 = x299 & n13688 ;
  assign n13690 = n6448 & ~n12602 ;
  assign n13691 = x51 | n13690 ;
  assign n13692 = ( x140 & ~n13639 ) | ( x140 & n13691 ) | ( ~n13639 & n13691 ) ;
  assign n13693 = ~n12602 & n12990 ;
  assign n13694 = x51 | n13693 ;
  assign n13695 = ( x140 & n13639 ) | ( x140 & ~n13694 ) | ( n13639 & ~n13694 ) ;
  assign n13696 = n13692 & ~n13695 ;
  assign n13697 = n13689 | n13696 ;
  assign n13698 = n4713 & ~n12603 ;
  assign n13699 = n12978 & ~n13698 ;
  assign n13700 = n6448 & ~n13699 ;
  assign n13701 = ~n6448 & n13311 ;
  assign n13702 = n13700 | n13701 ;
  assign n13703 = ( x140 & n7239 ) | ( x140 & n13702 ) | ( n7239 & n13702 ) ;
  assign n13704 = ~n4989 & n13311 ;
  assign n13705 = ( x224 & n4989 ) | ( x224 & ~n13699 ) | ( n4989 & ~n13699 ) ;
  assign n13706 = ( x224 & ~n4989 ) | ( x224 & n13677 ) | ( ~n4989 & n13677 ) ;
  assign n13707 = n13705 & ~n13706 ;
  assign n13708 = n13704 | n13707 ;
  assign n13709 = ( ~x140 & n7239 ) | ( ~x140 & n13708 ) | ( n7239 & n13708 ) ;
  assign n13710 = n13703 & n13709 ;
  assign n13711 = n13697 | n13710 ;
  assign n13712 = x232 & n13711 ;
  assign n13713 = ( x51 & ~n12603 ) | ( x51 & n12961 ) | ( ~n12603 & n12961 ) ;
  assign n13714 = ~x232 & n13713 ;
  assign n13715 = x39 & ~n13714 ;
  assign n13716 = ~n13712 & n13715 ;
  assign n13717 = ~x232 & n12507 ;
  assign n13718 = x39 | n13717 ;
  assign n13719 = n4713 & ~n12507 ;
  assign n13720 = n12887 & ~n13719 ;
  assign n13721 = ( x232 & ~n7241 ) | ( x232 & n13720 ) | ( ~n7241 & n13720 ) ;
  assign n13722 = ( x232 & n7241 ) | ( x232 & n12507 ) | ( n7241 & n12507 ) ;
  assign n13723 = n13721 & n13722 ;
  assign n13724 = n13718 | n13723 ;
  assign n13725 = ~n13716 & n13724 ;
  assign n13726 = ( x38 & ~x100 ) | ( x38 & n13725 ) | ( ~x100 & n13725 ) ;
  assign n13727 = ~n13672 & n13726 ;
  assign n13728 = n13658 | n13727 ;
  assign n13729 = ~n13663 & n13669 ;
  assign n13730 = n13728 & n13729 ;
  assign n13731 = n13671 & ~n13730 ;
  assign n13732 = n6785 | n13731 ;
  assign n13733 = x51 | x87 ;
  assign n13734 = n13685 | n13733 ;
  assign n13735 = n13669 & ~n13734 ;
  assign n13736 = x169 & n5924 ;
  assign n13737 = ~x87 & n12524 ;
  assign n13738 = ~n13736 & n13737 ;
  assign n13739 = x87 & ~n7899 ;
  assign n13740 = n6785 & ~n13739 ;
  assign n13741 = ~n13738 & n13740 ;
  assign n13742 = ~n13735 & n13741 ;
  assign n13743 = n13732 & ~n13742 ;
  assign n13744 = x100 | n11991 ;
  assign n13745 = x87 | n5769 ;
  assign n13746 = n13744 & ~n13745 ;
  assign n13747 = x75 | n13746 ;
  assign n13748 = ~n5763 & n13747 ;
  assign n13749 = x92 | n13748 ;
  assign n13750 = n7112 | n11665 ;
  assign n13751 = n13749 & ~n13750 ;
  assign n13752 = x51 & ~x151 ;
  assign n13753 = n11737 | n12409 ;
  assign n13754 = ~n13752 & n13753 ;
  assign n13755 = n12407 & n13754 ;
  assign n13756 = x232 & n13755 ;
  assign n13757 = x132 & n13307 ;
  assign n13758 = n13665 & ~n13757 ;
  assign n13759 = n12394 & ~n13758 ;
  assign n13760 = n12403 | n13759 ;
  assign n13761 = ~n13756 & n13760 ;
  assign n13762 = x87 | n13761 ;
  assign n13763 = x164 & n12861 ;
  assign n13764 = n6785 & ~n13763 ;
  assign n13765 = n13762 & n13764 ;
  assign n13766 = x190 | x299 ;
  assign n13767 = n4713 & ~n12541 ;
  assign n13768 = x182 & ~n13767 ;
  assign n13769 = n12514 & n13768 ;
  assign n13770 = ~x182 & n12541 ;
  assign n13771 = x173 | n13770 ;
  assign n13772 = n13769 | n13771 ;
  assign n13773 = n4713 & n12541 ;
  assign n13774 = n12508 | n13773 ;
  assign n13775 = ( ~x173 & x182 ) | ( ~x173 & n13774 ) | ( x182 & n13774 ) ;
  assign n13776 = n12537 | n13773 ;
  assign n13777 = ( x173 & x182 ) | ( x173 & ~n13776 ) | ( x182 & ~n13776 ) ;
  assign n13778 = ~n13775 & n13777 ;
  assign n13779 = n13772 & ~n13778 ;
  assign n13780 = n13766 | n13779 ;
  assign n13781 = ( x151 & x168 ) | ( x151 & ~n12507 ) | ( x168 & ~n12507 ) ;
  assign n13782 = ( x151 & ~x168 ) | ( x151 & n12513 ) | ( ~x168 & n12513 ) ;
  assign n13783 = ~n13781 & n13782 ;
  assign n13784 = x168 & ~n13752 ;
  assign n13785 = ( n4713 & n12887 ) | ( n4713 & n13784 ) | ( n12887 & n13784 ) ;
  assign n13786 = n13783 | n13785 ;
  assign n13787 = x160 & ~n13767 ;
  assign n13788 = n13786 & n13787 ;
  assign n13789 = ~x168 & n13776 ;
  assign n13790 = n12898 & ~n13767 ;
  assign n13791 = ( x151 & n11717 ) | ( x151 & ~n13790 ) | ( n11717 & ~n13790 ) ;
  assign n13792 = ~n13789 & n13791 ;
  assign n13793 = ~n11737 & n12541 ;
  assign n13794 = x168 & n12520 ;
  assign n13795 = x151 | n13794 ;
  assign n13796 = n13793 | n13795 ;
  assign n13797 = ~x160 & n13796 ;
  assign n13798 = ~n13792 & n13797 ;
  assign n13799 = x299 & ~n13798 ;
  assign n13800 = ~n13788 & n13799 ;
  assign n13801 = x190 & ~x299 ;
  assign n13802 = x182 & n12442 ;
  assign n13803 = n12469 | n13802 ;
  assign n13804 = x51 & ~x173 ;
  assign n13805 = n4713 | n13804 ;
  assign n13806 = n13803 & ~n13805 ;
  assign n13807 = n13801 & ~n13806 ;
  assign n13808 = ~n13773 & n13807 ;
  assign n13809 = x232 & ~n13808 ;
  assign n13810 = ~n13800 & n13809 ;
  assign n13811 = n13780 & n13810 ;
  assign n13812 = ~x232 & n12541 ;
  assign n13813 = n13811 | n13812 ;
  assign n13814 = ~x39 & n13813 ;
  assign n13815 = ~x149 & n7296 ;
  assign n13816 = ( ~n5005 & n13755 ) | ( ~n5005 & n13815 ) | ( n13755 & n13815 ) ;
  assign n13817 = x299 & ~n13816 ;
  assign n13818 = ( x151 & x168 ) | ( x151 & ~n12644 ) | ( x168 & ~n12644 ) ;
  assign n13819 = ( ~x151 & x168 ) | ( ~x151 & n12756 ) | ( x168 & n12756 ) ;
  assign n13820 = ~n13818 & n13819 ;
  assign n13821 = x149 & ~n13820 ;
  assign n13822 = ( x151 & ~x168 ) | ( x151 & n13016 ) | ( ~x168 & n13016 ) ;
  assign n13823 = ( x151 & x168 ) | ( x151 & n12988 ) | ( x168 & n12988 ) ;
  assign n13824 = n13822 & n13823 ;
  assign n13825 = n13821 & ~n13824 ;
  assign n13826 = ( ~x216 & n5005 ) | ( ~x216 & n13825 ) | ( n5005 & n13825 ) ;
  assign n13827 = ( x168 & n12979 ) | ( x168 & n13752 ) | ( n12979 & n13752 ) ;
  assign n13828 = ( ~x168 & n12991 ) | ( ~x168 & n13752 ) | ( n12991 & n13752 ) ;
  assign n13829 = n13827 | n13828 ;
  assign n13830 = ( x216 & n5005 ) | ( x216 & ~n13829 ) | ( n5005 & ~n13829 ) ;
  assign n13831 = n13826 & n13830 ;
  assign n13832 = n13817 & ~n13831 ;
  assign n13833 = x183 | n13000 ;
  assign n13834 = x183 | n12980 ;
  assign n13835 = x173 & ~n12985 ;
  assign n13836 = n13834 & n13835 ;
  assign n13837 = n13833 & ~n13836 ;
  assign n13838 = ( ~x173 & x183 ) | ( ~x173 & n12971 ) | ( x183 & n12971 ) ;
  assign n13839 = ( x173 & x183 ) | ( x173 & n12974 ) | ( x183 & n12974 ) ;
  assign n13840 = n13838 & ~n13839 ;
  assign n13841 = n13837 & ~n13840 ;
  assign n13842 = n13801 & ~n13841 ;
  assign n13843 = x183 & ~n12994 ;
  assign n13844 = x183 | n12409 ;
  assign n13845 = n12998 | n13844 ;
  assign n13846 = x173 & n13845 ;
  assign n13847 = ~n13843 & n13846 ;
  assign n13848 = x183 | n6448 ;
  assign n13849 = ~x173 & n13848 ;
  assign n13850 = n12966 & n13849 ;
  assign n13851 = n13766 | n13850 ;
  assign n13852 = n13847 | n13851 ;
  assign n13853 = ~n13842 & n13852 ;
  assign n13854 = ~n13832 & n13853 ;
  assign n13855 = x232 & ~n13854 ;
  assign n13856 = n12964 & ~n13855 ;
  assign n13857 = n13814 | n13856 ;
  assign n13858 = ~n1975 & n13857 ;
  assign n13859 = x299 & ~n13755 ;
  assign n13860 = x190 & n12525 ;
  assign n13861 = x173 & n12409 ;
  assign n13862 = n13860 | n13861 ;
  assign n13863 = ( x232 & n7916 ) | ( x232 & n13862 ) | ( n7916 & n13862 ) ;
  assign n13864 = ~n13859 & n13863 ;
  assign n13865 = n1975 & n13864 ;
  assign n13866 = n2043 | n13865 ;
  assign n13867 = n13858 | n13866 ;
  assign n13868 = n12682 & ~n13864 ;
  assign n13869 = x87 & ~n7248 ;
  assign n13870 = n13759 & ~n13869 ;
  assign n13871 = ~n13868 & n13870 ;
  assign n13872 = n13867 & n13871 ;
  assign n13873 = n2043 | n13485 ;
  assign n13874 = n13865 | n13873 ;
  assign n13875 = ~x151 & n12409 ;
  assign n13876 = x168 & ~n13875 ;
  assign n13877 = ~n12479 & n13876 ;
  assign n13878 = ( x151 & x168 ) | ( x151 & n12716 ) | ( x168 & n12716 ) ;
  assign n13879 = ( ~x151 & x168 ) | ( ~x151 & n12460 ) | ( x168 & n12460 ) ;
  assign n13880 = n13878 | n13879 ;
  assign n13881 = ~n13877 & n13880 ;
  assign n13882 = x160 | n13067 ;
  assign n13883 = n13881 | n13882 ;
  assign n13884 = x151 | n13755 ;
  assign n13885 = n13068 & ~n13884 ;
  assign n13886 = ~x168 & n12525 ;
  assign n13887 = n13067 | n13886 ;
  assign n13888 = x151 & n13887 ;
  assign n13889 = x160 & ~n13888 ;
  assign n13890 = ~n13885 & n13889 ;
  assign n13891 = x299 & ~n13890 ;
  assign n13892 = n13883 & n13891 ;
  assign n13893 = ~x182 & n12479 ;
  assign n13894 = n13067 | n13804 ;
  assign n13895 = n13893 | n13894 ;
  assign n13896 = n13801 & n13895 ;
  assign n13897 = x182 & ~n13068 ;
  assign n13898 = n13766 | n13861 ;
  assign n13899 = n12460 & ~n13898 ;
  assign n13900 = ~n13897 & n13899 ;
  assign n13901 = x232 & ~n13900 ;
  assign n13902 = ~n13896 & n13901 ;
  assign n13903 = ~n13892 & n13902 ;
  assign n13904 = ( ~x39 & n5788 ) | ( ~x39 & n12460 ) | ( n5788 & n12460 ) ;
  assign n13905 = ~n13903 & n13904 ;
  assign n13906 = n1975 | n13905 ;
  assign n13907 = x183 & ~n12615 ;
  assign n13908 = x173 | n13907 ;
  assign n13909 = n13197 & ~n13908 ;
  assign n13910 = ( x173 & ~x183 ) | ( x173 & n13179 ) | ( ~x183 & n13179 ) ;
  assign n13911 = ( x173 & x183 ) | ( x173 & n13191 ) | ( x183 & n13191 ) ;
  assign n13912 = n13910 & n13911 ;
  assign n13913 = n13909 | n13912 ;
  assign n13914 = n13801 & n13913 ;
  assign n13915 = n12403 & n13859 ;
  assign n13916 = n11170 | n13915 ;
  assign n13917 = x168 & ~n12604 ;
  assign n13918 = n11737 | n12600 ;
  assign n13919 = ~x151 & n13918 ;
  assign n13920 = ~n13917 & n13919 ;
  assign n13921 = x149 | n13920 ;
  assign n13922 = ( x151 & ~x168 ) | ( x151 & n12607 ) | ( ~x168 & n12607 ) ;
  assign n13923 = ( x151 & x168 ) | ( x151 & n12649 ) | ( x168 & n12649 ) ;
  assign n13924 = n13922 & n13923 ;
  assign n13925 = n13921 | n13924 ;
  assign n13926 = n7296 & n13925 ;
  assign n13927 = n12988 | n13752 ;
  assign n13928 = ~n12605 & n13927 ;
  assign n13929 = ( x149 & ~x168 ) | ( x149 & n13928 ) | ( ~x168 & n13928 ) ;
  assign n13930 = n12619 & ~n13754 ;
  assign n13931 = ( x149 & x168 ) | ( x149 & n13930 ) | ( x168 & n13930 ) ;
  assign n13932 = n13929 & n13931 ;
  assign n13933 = n13926 & ~n13932 ;
  assign n13934 = n13916 & ~n13933 ;
  assign n13935 = x183 & ~n12619 ;
  assign n13936 = n13183 & ~n13898 ;
  assign n13937 = ~n13935 & n13936 ;
  assign n13938 = n13934 | n13937 ;
  assign n13939 = n13914 | n13938 ;
  assign n13940 = x232 & n13939 ;
  assign n13941 = n13216 & ~n13940 ;
  assign n13942 = ( x39 & n13906 ) | ( x39 & ~n13941 ) | ( n13906 & ~n13941 ) ;
  assign n13943 = ~n13874 & n13942 ;
  assign n13944 = n12683 & ~n13864 ;
  assign n13945 = n13759 | n13869 ;
  assign n13946 = n13944 | n13945 ;
  assign n13947 = n13943 | n13946 ;
  assign n13948 = ~n6785 & n13947 ;
  assign n13949 = ~n13872 & n13948 ;
  assign n13950 = n13765 | n13949 ;
  assign n13951 = x197 & ~n12614 ;
  assign n13952 = n4322 | n13951 ;
  assign n13953 = n5124 & n13952 ;
  assign n13954 = x145 | n6448 ;
  assign n13955 = ~x299 & n13954 ;
  assign n13956 = n12965 & n13955 ;
  assign n13957 = n13953 | n13956 ;
  assign n13958 = ~n1868 & n13957 ;
  assign n13959 = x232 & ~n13958 ;
  assign n13960 = n12963 & ~n13959 ;
  assign n13961 = x39 & ~n13960 ;
  assign n13962 = n9514 | n13961 ;
  assign n13963 = ~x39 & x176 ;
  assign n13964 = ( n7680 & ~n12484 ) | ( n7680 & n13963 ) | ( ~n12484 & n13963 ) ;
  assign n13965 = n4713 & ~n12484 ;
  assign n13966 = n12514 & ~n13965 ;
  assign n13967 = ( n7680 & ~n13963 ) | ( n7680 & n13966 ) | ( ~n13963 & n13966 ) ;
  assign n13968 = n13964 & ~n13967 ;
  assign n13969 = n13962 | n13968 ;
  assign n13970 = x39 | x176 ;
  assign n13971 = x154 & n7916 ;
  assign n13972 = ( n12484 & n13970 ) | ( n12484 & ~n13971 ) | ( n13970 & ~n13971 ) ;
  assign n13973 = ( n13966 & n13970 ) | ( n13966 & n13971 ) | ( n13970 & n13971 ) ;
  assign n13974 = n13972 | n13973 ;
  assign n13975 = ~n13969 & n13974 ;
  assign n13976 = ~x133 & n12851 ;
  assign n13977 = ~x87 & n13976 ;
  assign n13978 = ~n13975 & n13977 ;
  assign n13979 = x145 & ~n12619 ;
  assign n13980 = n13210 & ~n13979 ;
  assign n13981 = n13211 & ~n13951 ;
  assign n13982 = n12403 | n13981 ;
  assign n13983 = x299 & n13982 ;
  assign n13984 = n13980 | n13983 ;
  assign n13985 = x232 & n13984 ;
  assign n13986 = n13216 & ~n13985 ;
  assign n13987 = ~n7683 & n12459 ;
  assign n13988 = n12403 | n13987 ;
  assign n13989 = ( ~x38 & n9138 ) | ( ~x38 & n13988 ) | ( n9138 & n13988 ) ;
  assign n13990 = ~n13986 & n13989 ;
  assign n13991 = n12430 | n13990 ;
  assign n13992 = ~n12678 & n13991 ;
  assign n13993 = n12683 | n13992 ;
  assign n13994 = ~n13976 & n13993 ;
  assign n13995 = x183 | x299 ;
  assign n13996 = ~x149 & x299 ;
  assign n13997 = n13995 & ~n13996 ;
  assign n13998 = n12861 & n13997 ;
  assign n13999 = ( x87 & n13994 ) | ( x87 & ~n13998 ) | ( n13994 & ~n13998 ) ;
  assign n14000 = n13978 | n13999 ;
  assign n14001 = ~n6785 & n14000 ;
  assign n14002 = n12404 | n13976 ;
  assign n14003 = x149 & n12861 ;
  assign n14004 = n6785 & ~n14003 ;
  assign n14005 = n14002 & n14004 ;
  assign n14006 = n14001 | n14005 ;
  assign n14007 = x136 | n13667 ;
  assign n14008 = x135 | n14007 ;
  assign n14009 = x134 & n14008 ;
  assign n14010 = n12402 | n14009 ;
  assign n14011 = n6785 & ~n13733 ;
  assign n14012 = x171 & ~n4713 ;
  assign n14013 = n12402 & n14012 ;
  assign n14014 = x232 & n14013 ;
  assign n14015 = n14011 & ~n14014 ;
  assign n14016 = n14010 & n14015 ;
  assign n14017 = x39 & x186 ;
  assign n14018 = x192 & ~x299 ;
  assign n14019 = n12614 & n13644 ;
  assign n14020 = n14018 & ~n14019 ;
  assign n14021 = x192 | x299 ;
  assign n14022 = n13182 & n13640 ;
  assign n14023 = n14021 | n14022 ;
  assign n14024 = ~n14020 & n14023 ;
  assign n14025 = n13624 & ~n14012 ;
  assign n14026 = x299 & ~n14025 ;
  assign n14027 = ( x171 & n7296 ) | ( x171 & n13181 ) | ( n7296 & n13181 ) ;
  assign n14028 = ( ~x171 & n7296 ) | ( ~x171 & n13635 ) | ( n7296 & n13635 ) ;
  assign n14029 = n14027 & n14028 ;
  assign n14030 = n14026 & ~n14029 ;
  assign n14031 = n14024 & ~n14030 ;
  assign n14032 = x232 & ~n14031 ;
  assign n14033 = n13621 & ~n14032 ;
  assign n14034 = n14017 & ~n14033 ;
  assign n14035 = x39 & ~x186 ;
  assign n14036 = ~n13644 & n14018 ;
  assign n14037 = n13640 | n14021 ;
  assign n14038 = ~n14036 & n14037 ;
  assign n14039 = ~n14030 & n14038 ;
  assign n14040 = x232 & ~n14039 ;
  assign n14041 = n13621 & ~n14040 ;
  assign n14042 = n14035 & ~n14041 ;
  assign n14043 = x171 & x299 ;
  assign n14044 = n14018 | n14043 ;
  assign n14045 = n5924 & n14044 ;
  assign n14046 = n12524 & ~n14045 ;
  assign n14047 = x39 | n14046 ;
  assign n14048 = x164 & n14047 ;
  assign n14049 = ~n14042 & n14048 ;
  assign n14050 = ~n14034 & n14049 ;
  assign n14051 = n2926 & ~n4713 ;
  assign n14052 = n12641 & ~n14012 ;
  assign n14053 = n7296 & ~n14052 ;
  assign n14054 = ~n14051 & n14053 ;
  assign n14055 = n14026 & ~n14054 ;
  assign n14056 = n14024 & ~n14055 ;
  assign n14057 = x232 & ~n14056 ;
  assign n14058 = n13621 & ~n14057 ;
  assign n14059 = n14017 & ~n14058 ;
  assign n14060 = n14038 & ~n14055 ;
  assign n14061 = x232 & ~n14060 ;
  assign n14062 = n13621 & ~n14061 ;
  assign n14063 = n14035 & ~n14062 ;
  assign n14064 = ~x164 & n14047 ;
  assign n14065 = ~n14063 & n14064 ;
  assign n14066 = ~n14059 & n14065 ;
  assign n14067 = n1975 | n14066 ;
  assign n14068 = n14050 | n14067 ;
  assign n14069 = n13311 & ~n14046 ;
  assign n14070 = n1975 & n14069 ;
  assign n14071 = n2043 | n14070 ;
  assign n14072 = n13485 | n14071 ;
  assign n14073 = n14068 & ~n14072 ;
  assign n14074 = n12682 & n14046 ;
  assign n14075 = n14009 | n14074 ;
  assign n14076 = n14073 | n14075 ;
  assign n14077 = n12603 | n14012 ;
  assign n14078 = x171 & ~n12978 ;
  assign n14079 = n14077 & ~n14078 ;
  assign n14080 = x216 | n14079 ;
  assign n14081 = x164 & x216 ;
  assign n14082 = ( x171 & n13677 ) | ( x171 & ~n14081 ) | ( n13677 & ~n14081 ) ;
  assign n14083 = ( x171 & ~n13680 ) | ( x171 & n14081 ) | ( ~n13680 & n14081 ) ;
  assign n14084 = ~n14082 & n14083 ;
  assign n14085 = n14080 & ~n14084 ;
  assign n14086 = n5005 & ~n14085 ;
  assign n14087 = x51 | n14013 ;
  assign n14088 = ~x164 & n7296 ;
  assign n14089 = ( ~n5005 & n14087 ) | ( ~n5005 & n14088 ) | ( n14087 & n14088 ) ;
  assign n14090 = n14086 | n14089 ;
  assign n14091 = x299 & n14090 ;
  assign n14092 = n13702 & n14018 ;
  assign n14093 = n13691 & ~n14021 ;
  assign n14094 = n14017 | n14093 ;
  assign n14095 = n14092 | n14094 ;
  assign n14096 = n13708 & n14018 ;
  assign n14097 = n13694 & ~n14021 ;
  assign n14098 = x186 & ~n14097 ;
  assign n14099 = ~n14096 & n14098 ;
  assign n14100 = n14095 & ~n14099 ;
  assign n14101 = n14091 | n14100 ;
  assign n14102 = x232 & n14101 ;
  assign n14103 = n13715 & ~n14102 ;
  assign n14104 = n1975 | n14103 ;
  assign n14105 = x232 & n14044 ;
  assign n14106 = ( x39 & n13720 ) | ( x39 & n14105 ) | ( n13720 & n14105 ) ;
  assign n14107 = ( x39 & n12507 ) | ( x39 & ~n14105 ) | ( n12507 & ~n14105 ) ;
  assign n14108 = n14106 | n14107 ;
  assign n14109 = ~n14104 & n14108 ;
  assign n14110 = n14071 | n14109 ;
  assign n14111 = n12682 & ~n14069 ;
  assign n14112 = n14009 & ~n14111 ;
  assign n14113 = n14110 & n14112 ;
  assign n14114 = n6785 | n14113 ;
  assign n14115 = n14076 & ~n14114 ;
  assign n14116 = n14016 | n14115 ;
  assign n14117 = x170 & ~n4713 ;
  assign n14118 = n7916 & n14117 ;
  assign n14119 = n12524 & ~n14118 ;
  assign n14120 = x194 & n7252 ;
  assign n14121 = n14119 & ~n14120 ;
  assign n14122 = n13311 & ~n14121 ;
  assign n14123 = x100 & n14122 ;
  assign n14124 = n2043 | n14123 ;
  assign n14125 = n13311 & ~n14119 ;
  assign n14126 = ( x38 & x194 ) | ( x38 & ~n14125 ) | ( x194 & ~n14125 ) ;
  assign n14127 = n12603 | n14117 ;
  assign n14128 = x170 & ~n12978 ;
  assign n14129 = n6433 & ~n14128 ;
  assign n14130 = n14127 & n14129 ;
  assign n14131 = n7296 | n14130 ;
  assign n14132 = ( x170 & x216 ) | ( x170 & ~n13680 ) | ( x216 & ~n13680 ) ;
  assign n14133 = ( x170 & ~x216 ) | ( x170 & n13677 ) | ( ~x216 & n13677 ) ;
  assign n14134 = n14132 & ~n14133 ;
  assign n14135 = n14131 & ~n14134 ;
  assign n14136 = x150 & x299 ;
  assign n14137 = n12402 & n14117 ;
  assign n14138 = x51 | n14137 ;
  assign n14139 = n5005 | n14138 ;
  assign n14140 = n14136 & n14139 ;
  assign n14141 = ~n14135 & n14140 ;
  assign n14142 = n6433 | n14138 ;
  assign n14143 = n13492 & n14142 ;
  assign n14144 = ~n14130 & n14143 ;
  assign n14145 = n14141 | n14144 ;
  assign n14146 = ( x185 & x299 ) | ( x185 & ~n13694 ) | ( x299 & ~n13694 ) ;
  assign n14147 = ( x185 & ~x299 ) | ( x185 & n13691 ) | ( ~x299 & n13691 ) ;
  assign n14148 = ~n14146 & n14147 ;
  assign n14149 = n14145 | n14148 ;
  assign n14150 = x232 & n14149 ;
  assign n14151 = n13715 & ~n14150 ;
  assign n14152 = ~x299 & n12507 ;
  assign n14153 = ( x170 & n7916 ) | ( x170 & n12507 ) | ( n7916 & n12507 ) ;
  assign n14154 = ( ~x170 & n7916 ) | ( ~x170 & n13720 ) | ( n7916 & n13720 ) ;
  assign n14155 = n14153 & n14154 ;
  assign n14156 = n13718 | n14155 ;
  assign n14157 = n14152 | n14156 ;
  assign n14158 = ~n14151 & n14157 ;
  assign n14159 = ( x38 & ~x194 ) | ( x38 & n14158 ) | ( ~x194 & n14158 ) ;
  assign n14160 = ~n14126 & n14159 ;
  assign n14161 = ( x185 & x299 ) | ( x185 & ~n13708 ) | ( x299 & ~n13708 ) ;
  assign n14162 = ( x185 & ~x299 ) | ( x185 & n13702 ) | ( ~x299 & n13702 ) ;
  assign n14163 = ~n14161 & n14162 ;
  assign n14164 = n14145 | n14163 ;
  assign n14165 = x232 & n14164 ;
  assign n14166 = n13715 & ~n14165 ;
  assign n14167 = n8828 & n13720 ;
  assign n14168 = n14156 | n14167 ;
  assign n14169 = ~n14166 & n14168 ;
  assign n14170 = ( x38 & x194 ) | ( x38 & n14169 ) | ( x194 & n14169 ) ;
  assign n14171 = x170 & n5924 ;
  assign n14172 = n7252 | n14171 ;
  assign n14173 = n12524 & ~n14172 ;
  assign n14174 = n13311 & ~n14173 ;
  assign n14175 = ( ~x38 & x194 ) | ( ~x38 & n14174 ) | ( x194 & n14174 ) ;
  assign n14176 = n14170 & n14175 ;
  assign n14177 = n14160 | n14176 ;
  assign n14178 = ~x100 & n14177 ;
  assign n14179 = n14124 | n14178 ;
  assign n14180 = x135 & n14007 ;
  assign n14181 = x134 & ~n14008 ;
  assign n14182 = n14180 | n14181 ;
  assign n14183 = n12682 & ~n14122 ;
  assign n14184 = n14182 & ~n14183 ;
  assign n14185 = n14179 & n14184 ;
  assign n14186 = x185 & ~n13182 ;
  assign n14187 = n13640 & ~n14186 ;
  assign n14188 = ~n9138 & n14119 ;
  assign n14189 = x194 | n14188 ;
  assign n14190 = n14187 | n14189 ;
  assign n14191 = ~x185 & n13644 ;
  assign n14192 = ~n9138 & n14173 ;
  assign n14193 = x194 & ~n14192 ;
  assign n14194 = ~n14019 & n14193 ;
  assign n14195 = ~n14191 & n14194 ;
  assign n14196 = n14190 & ~n14195 ;
  assign n14197 = x299 | n14196 ;
  assign n14198 = ( x170 & n7296 ) | ( x170 & n13181 ) | ( n7296 & n13181 ) ;
  assign n14199 = ( ~x170 & n7296 ) | ( ~x170 & n13635 ) | ( n7296 & n13635 ) ;
  assign n14200 = n14198 & n14199 ;
  assign n14201 = n14136 & ~n14200 ;
  assign n14202 = n3129 & ~n4713 ;
  assign n14203 = n12641 & ~n14117 ;
  assign n14204 = n7296 & ~n14203 ;
  assign n14205 = ~n14202 & n14204 ;
  assign n14206 = n13492 & ~n14205 ;
  assign n14207 = n14201 | n14206 ;
  assign n14208 = n13624 & ~n14117 ;
  assign n14209 = n14189 & ~n14193 ;
  assign n14210 = n14208 | n14209 ;
  assign n14211 = n14207 & ~n14210 ;
  assign n14212 = n14197 & ~n14211 ;
  assign n14213 = x232 & ~n14212 ;
  assign n14214 = n13622 | n14209 ;
  assign n14215 = ~n14213 & n14214 ;
  assign n14216 = x100 | n14215 ;
  assign n14217 = n12677 | n14124 ;
  assign n14218 = n14216 & ~n14217 ;
  assign n14219 = n12682 & n14121 ;
  assign n14220 = n14182 | n14219 ;
  assign n14221 = n14218 | n14220 ;
  assign n14222 = ~n6785 & n14221 ;
  assign n14223 = ~n14185 & n14222 ;
  assign n14224 = ( n12402 & ~n14011 ) | ( n12402 & n14171 ) | ( ~n14011 & n14171 ) ;
  assign n14225 = ( n12402 & n14011 ) | ( n12402 & n14182 ) | ( n14011 & n14182 ) ;
  assign n14226 = ~n14224 & n14225 ;
  assign n14227 = n14223 | n14226 ;
  assign n14228 = x136 & n13667 ;
  assign n14229 = n14007 & ~n14228 ;
  assign n14230 = n12392 & ~n14229 ;
  assign n14231 = ~n12524 & n14230 ;
  assign n14232 = x148 & n5924 ;
  assign n14233 = n12402 & ~n14232 ;
  assign n14234 = n14231 | n14233 ;
  assign n14235 = n14011 & n14234 ;
  assign n14236 = ( x232 & ~n7932 ) | ( x232 & n13720 ) | ( ~n7932 & n13720 ) ;
  assign n14237 = ( x232 & n7932 ) | ( x232 & n12507 ) | ( n7932 & n12507 ) ;
  assign n14238 = n14236 & n14237 ;
  assign n14239 = n13718 | n14238 ;
  assign n14240 = n6433 & ~n13699 ;
  assign n14241 = x163 & n5005 ;
  assign n14242 = n13677 & n14241 ;
  assign n14243 = n5005 | n13311 ;
  assign n14244 = ~n6433 & n13311 ;
  assign n14245 = ( x163 & n14243 ) | ( x163 & n14244 ) | ( n14243 & n14244 ) ;
  assign n14246 = ~n14242 & n14245 ;
  assign n14247 = x148 & ~n14246 ;
  assign n14248 = ~n14240 & n14247 ;
  assign n14249 = ~x287 & n11674 ;
  assign n14250 = x216 & ~n14249 ;
  assign n14251 = n5005 & ~n14250 ;
  assign n14252 = ~n12602 & n14251 ;
  assign n14253 = x51 | x148 ;
  assign n14254 = n14252 | n14253 ;
  assign n14255 = x299 & n14254 ;
  assign n14256 = ~n14248 & n14255 ;
  assign n14257 = x141 | x299 ;
  assign n14258 = ( x184 & n13691 ) | ( x184 & ~n14257 ) | ( n13691 & ~n14257 ) ;
  assign n14259 = ( x184 & ~n13694 ) | ( x184 & n14257 ) | ( ~n13694 & n14257 ) ;
  assign n14260 = n14258 & ~n14259 ;
  assign n14261 = n14256 | n14260 ;
  assign n14262 = ( x184 & n7930 ) | ( x184 & n13702 ) | ( n7930 & n13702 ) ;
  assign n14263 = ( ~x184 & n7930 ) | ( ~x184 & n13708 ) | ( n7930 & n13708 ) ;
  assign n14264 = n14262 & n14263 ;
  assign n14265 = n14261 | n14264 ;
  assign n14266 = x232 & n14265 ;
  assign n14267 = n13715 & ~n14266 ;
  assign n14268 = n1975 | n14267 ;
  assign n14269 = n14239 & ~n14268 ;
  assign n14270 = n7933 & n12402 ;
  assign n14271 = x51 | n14270 ;
  assign n14272 = n1975 & n14271 ;
  assign n14273 = n2043 | n14272 ;
  assign n14274 = n14269 | n14273 ;
  assign n14275 = n12682 & ~n14271 ;
  assign n14276 = n14230 & ~n14275 ;
  assign n14277 = n14274 & n14276 ;
  assign n14278 = ~n9306 & n12402 ;
  assign n14279 = ~n14271 & n14278 ;
  assign n14280 = n7296 & ~n13634 ;
  assign n14281 = x148 & ~n4713 ;
  assign n14282 = ( x148 & ~n13624 ) | ( x148 & n14281 ) | ( ~n13624 & n14281 ) ;
  assign n14283 = ~n14280 & n14282 ;
  assign n14284 = ~x51 & n13211 ;
  assign n14285 = x148 | n14284 ;
  assign n14286 = ~n14249 & n14285 ;
  assign n14287 = ~x148 & n12524 ;
  assign n14288 = n14286 | n14287 ;
  assign n14289 = ~n14283 & n14288 ;
  assign n14290 = x299 & ~n14289 ;
  assign n14291 = x184 & ~n13182 ;
  assign n14292 = n13640 & ~n14291 ;
  assign n14293 = n14257 | n14292 ;
  assign n14294 = x184 & ~n12614 ;
  assign n14295 = n13644 & ~n14294 ;
  assign n14296 = n7930 & ~n14295 ;
  assign n14297 = n14293 & ~n14296 ;
  assign n14298 = ~n14290 & n14297 ;
  assign n14299 = x232 & ~n14298 ;
  assign n14300 = ~x100 & n13622 ;
  assign n14301 = ~n14299 & n14300 ;
  assign n14302 = n14279 | n14301 ;
  assign n14303 = ~n2043 & n14302 ;
  assign n14304 = n12402 & n14275 ;
  assign n14305 = n14230 | n14304 ;
  assign n14306 = n14303 | n14305 ;
  assign n14307 = ~n6785 & n14306 ;
  assign n14308 = ~n14277 & n14307 ;
  assign n14309 = n14235 | n14308 ;
  assign n14310 = ~x39 & x137 ;
  assign n14311 = n8609 & ~n12808 ;
  assign n14312 = n4693 & ~n9701 ;
  assign n14313 = x299 | n6785 ;
  assign n14314 = x198 | n9711 ;
  assign n14315 = n14313 | n14314 ;
  assign n14316 = ~n14312 & n14315 ;
  assign n14317 = n14311 | n14316 ;
  assign n14318 = x210 | n9701 ;
  assign n14319 = n6785 & ~n14318 ;
  assign n14320 = n14317 & ~n14319 ;
  assign n14321 = n8469 & ~n14320 ;
  assign n14322 = n14310 | n14321 ;
  assign n14323 = n7684 & ~n7732 ;
  assign n14324 = x92 & ~n14323 ;
  assign n14325 = n2030 | n14324 ;
  assign n14326 = x75 | n7675 ;
  assign n14327 = n7614 & ~n14281 ;
  assign n14328 = x148 & n11725 ;
  assign n14329 = n14327 | n14328 ;
  assign n14330 = x299 & n14329 ;
  assign n14331 = ~x299 & n8084 ;
  assign n14332 = ( x141 & x232 ) | ( x141 & ~n14331 ) | ( x232 & ~n14331 ) ;
  assign n14333 = n4713 & n8084 ;
  assign n14334 = n11747 | n14333 ;
  assign n14335 = ~x299 & n14334 ;
  assign n14336 = ( x141 & ~x232 ) | ( x141 & n14335 ) | ( ~x232 & n14335 ) ;
  assign n14337 = n14332 & ~n14336 ;
  assign n14338 = ~n14330 & n14337 ;
  assign n14339 = x299 & n7614 ;
  assign n14340 = n14331 | n14339 ;
  assign n14341 = ( ~x39 & n5788 ) | ( ~x39 & n14340 ) | ( n5788 & n14340 ) ;
  assign n14342 = ~n14338 & n14341 ;
  assign n14343 = n7301 & n10257 ;
  assign n14344 = n7320 & ~n14343 ;
  assign n14345 = n11791 & ~n14344 ;
  assign n14346 = n4721 & n7301 ;
  assign n14347 = n7296 & ~n14343 ;
  assign n14348 = ~n14346 & n14347 ;
  assign n14349 = n7298 & ~n14348 ;
  assign n14350 = n14345 | n14349 ;
  assign n14351 = ~x232 & n14350 ;
  assign n14352 = n7306 | n14343 ;
  assign n14353 = n7297 & n14352 ;
  assign n14354 = x148 & ~n14353 ;
  assign n14355 = n7931 | n14349 ;
  assign n14356 = ~n14354 & n14355 ;
  assign n14357 = ~n7328 & n14344 ;
  assign n14358 = n11791 & ~n14357 ;
  assign n14359 = ( x141 & n14356 ) | ( x141 & n14358 ) | ( n14356 & n14358 ) ;
  assign n14360 = ( ~x141 & n14345 ) | ( ~x141 & n14356 ) | ( n14345 & n14356 ) ;
  assign n14361 = n14359 | n14360 ;
  assign n14362 = x232 & n14361 ;
  assign n14363 = n14351 | n14362 ;
  assign n14364 = x39 & n14363 ;
  assign n14365 = n1975 | n14364 ;
  assign n14366 = n14342 | n14365 ;
  assign n14367 = ~x87 & n14366 ;
  assign n14368 = n14326 | n14367 ;
  assign n14369 = ~x92 & n14368 ;
  assign n14370 = n14325 | n14369 ;
  assign n14371 = ~x55 & n14370 ;
  assign n14372 = ~n7733 & n11827 ;
  assign n14373 = x55 & ~n14372 ;
  assign n14374 = n14371 | n14373 ;
  assign n14375 = ~n2058 & n14374 ;
  assign n14376 = n8073 | n14375 ;
  assign n14377 = x118 | n11843 ;
  assign n14378 = x139 | n14377 ;
  assign n14379 = ( ~x138 & n14376 ) | ( ~x138 & n14378 ) | ( n14376 & n14378 ) ;
  assign n14380 = ~n4904 & n7808 ;
  assign n14381 = ~n7933 & n14380 ;
  assign n14382 = ( x39 & ~n8366 ) | ( x39 & n14381 ) | ( ~n8366 & n14381 ) ;
  assign n14383 = x232 | n9617 ;
  assign n14384 = n4714 & n4988 ;
  assign n14385 = n7285 & n14384 ;
  assign n14386 = ~n4714 & n7931 ;
  assign n14387 = ( n7930 & ~n14385 ) | ( n7930 & n14386 ) | ( ~n14385 & n14386 ) ;
  assign n14388 = ( n7930 & n9617 ) | ( n7930 & ~n14386 ) | ( n9617 & ~n14386 ) ;
  assign n14389 = ~n14387 & n14388 ;
  assign n14390 = x232 & ~n14389 ;
  assign n14391 = n14383 & ~n14390 ;
  assign n14392 = ( x39 & n8366 ) | ( x39 & ~n14391 ) | ( n8366 & ~n14391 ) ;
  assign n14393 = n14382 & ~n14392 ;
  assign n14394 = ( x138 & n14378 ) | ( x138 & ~n14393 ) | ( n14378 & ~n14393 ) ;
  assign n14395 = n14379 & n14394 ;
  assign n14396 = ~x138 & n7204 ;
  assign n14397 = ( n14378 & n14393 ) | ( n14378 & ~n14396 ) | ( n14393 & ~n14396 ) ;
  assign n14398 = ( ~n14376 & n14378 ) | ( ~n14376 & n14396 ) | ( n14378 & n14396 ) ;
  assign n14399 = n14397 | n14398 ;
  assign n14400 = ~n14395 & n14399 ;
  assign n14401 = n7614 & ~n13623 ;
  assign n14402 = x169 & n11725 ;
  assign n14403 = n14401 | n14402 ;
  assign n14404 = x299 & n14403 ;
  assign n14405 = ( x191 & x232 ) | ( x191 & ~n14331 ) | ( x232 & ~n14331 ) ;
  assign n14406 = ( x191 & ~x232 ) | ( x191 & n14335 ) | ( ~x232 & n14335 ) ;
  assign n14407 = n14405 & ~n14406 ;
  assign n14408 = ~n14404 & n14407 ;
  assign n14409 = n14341 & ~n14408 ;
  assign n14410 = x169 | n7301 ;
  assign n14411 = n14352 & n14410 ;
  assign n14412 = n7296 & ~n14411 ;
  assign n14413 = n7298 & ~n14412 ;
  assign n14414 = ( x191 & n14358 ) | ( x191 & n14413 ) | ( n14358 & n14413 ) ;
  assign n14415 = ( ~x191 & n14345 ) | ( ~x191 & n14413 ) | ( n14345 & n14413 ) ;
  assign n14416 = n14414 | n14415 ;
  assign n14417 = x232 & n14416 ;
  assign n14418 = n14351 | n14417 ;
  assign n14419 = x39 & n14418 ;
  assign n14420 = n1975 | n14419 ;
  assign n14421 = n14409 | n14420 ;
  assign n14422 = ~x87 & n14421 ;
  assign n14423 = n14326 | n14422 ;
  assign n14424 = ~x92 & n14423 ;
  assign n14425 = n14325 | n14424 ;
  assign n14426 = ~x55 & n14425 ;
  assign n14427 = n14373 | n14426 ;
  assign n14428 = ~n2058 & n14427 ;
  assign n14429 = n8073 | n14428 ;
  assign n14430 = ( ~x139 & n14377 ) | ( ~x139 & n14429 ) | ( n14377 & n14429 ) ;
  assign n14431 = ~n13652 & n14380 ;
  assign n14432 = ( x39 & ~n8366 ) | ( x39 & n14431 ) | ( ~n8366 & n14431 ) ;
  assign n14433 = ~n4714 & n7240 ;
  assign n14434 = n9616 | n14433 ;
  assign n14435 = n9613 | n13639 ;
  assign n14436 = n7239 & ~n14385 ;
  assign n14437 = n14435 & ~n14436 ;
  assign n14438 = ~n14434 & n14437 ;
  assign n14439 = x232 & ~n14438 ;
  assign n14440 = n14383 & ~n14439 ;
  assign n14441 = ( x39 & n8366 ) | ( x39 & ~n14440 ) | ( n8366 & ~n14440 ) ;
  assign n14442 = n14432 & ~n14441 ;
  assign n14443 = ( x139 & n14377 ) | ( x139 & ~n14442 ) | ( n14377 & ~n14442 ) ;
  assign n14444 = n14430 & n14443 ;
  assign n14445 = ~x139 & n7205 ;
  assign n14446 = ( n14377 & n14442 ) | ( n14377 & ~n14445 ) | ( n14442 & ~n14445 ) ;
  assign n14447 = ( n14377 & ~n14429 ) | ( n14377 & n14445 ) | ( ~n14429 & n14445 ) ;
  assign n14448 = n14446 | n14447 ;
  assign n14449 = ~n14444 & n14448 ;
  assign n14450 = n4717 | n4719 ;
  assign n14451 = n1290 & ~n4977 ;
  assign n14452 = ~n4980 & n14451 ;
  assign n14453 = ~n1271 & n14452 ;
  assign n14454 = ~n1242 & n14453 ;
  assign n14455 = x120 | n14454 ;
  assign n14456 = n1290 & ~n1462 ;
  assign n14457 = ~n1865 & n14456 ;
  assign n14458 = ~n12253 & n14457 ;
  assign n14459 = x120 & ~n14457 ;
  assign n14460 = x120 & n4730 ;
  assign n14461 = ( ~n14458 & n14459 ) | ( ~n14458 & n14460 ) | ( n14459 & n14460 ) ;
  assign n14462 = x1091 & ~n14461 ;
  assign n14463 = ~x120 & x1091 ;
  assign n14464 = ( ~n1272 & n14462 ) | ( ~n1272 & n14463 ) | ( n14462 & n14463 ) ;
  assign n14465 = n14455 & n14464 ;
  assign n14466 = ( x120 & n1271 ) | ( x120 & n14459 ) | ( n1271 & n14459 ) ;
  assign n14467 = x120 | n14459 ;
  assign n14468 = ( n1242 & n14466 ) | ( n1242 & n14467 ) | ( n14466 & n14467 ) ;
  assign n14469 = x1091 | n14468 ;
  assign n14470 = x120 & x824 ;
  assign n14471 = x1091 | n14470 ;
  assign n14472 = n14468 | n14471 ;
  assign n14473 = ( n4730 & n14469 ) | ( n4730 & n14472 ) | ( n14469 & n14472 ) ;
  assign n14474 = n14455 & ~n14473 ;
  assign n14475 = n14465 | n14474 ;
  assign n14476 = n4977 | n4980 ;
  assign n14477 = n1271 | n14476 ;
  assign n14478 = n1242 | n14477 ;
  assign n14479 = ~x120 & n14478 ;
  assign n14480 = x120 & n1868 ;
  assign n14481 = n14479 | n14480 ;
  assign n14482 = n1290 | n4713 ;
  assign n14483 = ~n4713 & n14482 ;
  assign n14484 = ~n14481 & n14483 ;
  assign n14485 = n1290 | n4706 ;
  assign n14486 = ( n4706 & ~n14481 ) | ( n4706 & n14485 ) | ( ~n14481 & n14485 ) ;
  assign n14487 = ~n4706 & n14485 ;
  assign n14488 = ~n14481 & n14487 ;
  assign n14489 = ( n14484 & n14486 ) | ( n14484 & n14488 ) | ( n14486 & n14488 ) ;
  assign n14490 = ( n4713 & ~n14481 ) | ( n4713 & n14482 ) | ( ~n14481 & n14482 ) ;
  assign n14491 = ( n14486 & n14488 ) | ( n14486 & n14490 ) | ( n14488 & n14490 ) ;
  assign n14492 = ( n14475 & n14489 ) | ( n14475 & n14491 ) | ( n14489 & n14491 ) ;
  assign n14493 = x616 & ~n1290 ;
  assign n14494 = ( x616 & n14481 ) | ( x616 & n14493 ) | ( n14481 & n14493 ) ;
  assign n14495 = x614 & ~x616 ;
  assign n14496 = x614 & ~n1290 ;
  assign n14497 = ~x616 & n14496 ;
  assign n14498 = ( n14481 & n14495 ) | ( n14481 & n14497 ) | ( n14495 & n14497 ) ;
  assign n14499 = n14494 | n14498 ;
  assign n14500 = x616 & ~n14493 ;
  assign n14501 = ~n14481 & n14500 ;
  assign n14502 = ( x614 & ~n14499 ) | ( x614 & n14501 ) | ( ~n14499 & n14501 ) ;
  assign n14503 = n14499 & ~n14501 ;
  assign n14504 = ( n14492 & n14502 ) | ( n14492 & ~n14503 ) | ( n14502 & ~n14503 ) ;
  assign n14505 = n4709 | n14504 ;
  assign n14506 = n4709 & ~n14465 ;
  assign n14507 = ~n14474 & n14506 ;
  assign n14508 = n4713 & ~n14507 ;
  assign n14509 = ~n4713 & n14465 ;
  assign n14510 = ( ~n4713 & n14474 ) | ( ~n4713 & n14509 ) | ( n14474 & n14509 ) ;
  assign n14511 = n14508 | n14510 ;
  assign n14512 = ~x661 & n14511 ;
  assign n14513 = ~x661 & n14510 ;
  assign n14514 = ( n14505 & n14512 ) | ( n14505 & n14513 ) | ( n14512 & n14513 ) ;
  assign n14515 = x614 | n14492 ;
  assign n14516 = n1290 & n4713 ;
  assign n14517 = ~n14481 & n14516 ;
  assign n14518 = x616 & n14517 ;
  assign n14519 = ( x616 & n14510 ) | ( x616 & n14518 ) | ( n14510 & n14518 ) ;
  assign n14520 = x681 & ~n14519 ;
  assign n14521 = n14510 | n14517 ;
  assign n14522 = x681 & ~n14521 ;
  assign n14523 = ( ~n14515 & n14520 ) | ( ~n14515 & n14522 ) | ( n14520 & n14522 ) ;
  assign n14524 = ( x681 & n4710 ) | ( x681 & n14519 ) | ( n4710 & n14519 ) ;
  assign n14525 = ( x681 & n4710 ) | ( x681 & n14521 ) | ( n4710 & n14521 ) ;
  assign n14526 = ( n14515 & n14524 ) | ( n14515 & n14525 ) | ( n14524 & n14525 ) ;
  assign n14527 = ~n14523 & n14526 ;
  assign n14528 = ( n14514 & ~n14523 ) | ( n14514 & n14527 ) | ( ~n14523 & n14527 ) ;
  assign n14529 = n14450 & ~n14528 ;
  assign n14530 = x680 & ~n14484 ;
  assign n14531 = x680 & ~n14482 ;
  assign n14532 = x680 & ~n4713 ;
  assign n14533 = ( n14481 & n14531 ) | ( n14481 & n14532 ) | ( n14531 & n14532 ) ;
  assign n14534 = ( ~n14475 & n14530 ) | ( ~n14475 & n14533 ) | ( n14530 & n14533 ) ;
  assign n14535 = x616 | x662 ;
  assign n14536 = n4710 | n14535 ;
  assign n14537 = n14534 | n14536 ;
  assign n14538 = ~x616 & n14498 ;
  assign n14539 = ~x680 & n14538 ;
  assign n14540 = ( x614 & x616 ) | ( x614 & ~n14498 ) | ( x616 & ~n14498 ) ;
  assign n14541 = x680 | n14540 ;
  assign n14542 = ( n14492 & ~n14539 ) | ( n14492 & n14541 ) | ( ~n14539 & n14541 ) ;
  assign n14543 = ~n14537 & n14542 ;
  assign n14544 = x680 | n1290 ;
  assign n14545 = x616 & ~x662 ;
  assign n14546 = ~n4710 & n14545 ;
  assign n14547 = n14544 & n14546 ;
  assign n14548 = x680 & n14546 ;
  assign n14549 = ( ~n14481 & n14547 ) | ( ~n14481 & n14548 ) | ( n14547 & n14548 ) ;
  assign n14550 = ~n14484 & n14549 ;
  assign n14551 = ~n14490 & n14549 ;
  assign n14552 = ( ~n14475 & n14550 ) | ( ~n14475 & n14551 ) | ( n14550 & n14551 ) ;
  assign n14553 = x662 | n4710 ;
  assign n14554 = x616 & n1290 ;
  assign n14555 = n14553 & n14554 ;
  assign n14556 = ~n14481 & n14555 ;
  assign n14557 = n14549 | n14556 ;
  assign n14558 = x681 | n14557 ;
  assign n14559 = ( ~x680 & n14549 ) | ( ~x680 & n14556 ) | ( n14549 & n14556 ) ;
  assign n14560 = x681 | n14559 ;
  assign n14561 = ( ~n14552 & n14558 ) | ( ~n14552 & n14560 ) | ( n14558 & n14560 ) ;
  assign n14562 = ~x616 & x662 ;
  assign n14563 = ( ~x616 & n4710 ) | ( ~x616 & n14562 ) | ( n4710 & n14562 ) ;
  assign n14564 = ~n14496 & n14563 ;
  assign n14565 = ~x614 & n14563 ;
  assign n14566 = ( ~n14481 & n14564 ) | ( ~n14481 & n14565 ) | ( n14564 & n14565 ) ;
  assign n14567 = x614 & n14566 ;
  assign n14568 = ( n14492 & n14566 ) | ( n14492 & n14567 ) | ( n14566 & n14567 ) ;
  assign n14569 = n14561 | n14568 ;
  assign n14570 = n14543 | n14569 ;
  assign n14571 = x681 & ~n14504 ;
  assign n14572 = n14450 | n14571 ;
  assign n14573 = n14570 & ~n14572 ;
  assign n14574 = ( ~n4718 & n14450 ) | ( ~n4718 & n14573 ) | ( n14450 & n14573 ) ;
  assign n14575 = ~n14529 & n14574 ;
  assign n14576 = x215 & ~n4718 ;
  assign n14577 = ( x215 & ~n14528 ) | ( x215 & n14576 ) | ( ~n14528 & n14576 ) ;
  assign n14578 = x299 & n14577 ;
  assign n14579 = ~n14575 & n14578 ;
  assign n14580 = ~x661 & n4709 ;
  assign n14581 = n1287 & n14454 ;
  assign n14582 = n4980 | n8368 ;
  assign n14583 = n1271 | n14582 ;
  assign n14584 = n1242 | n14583 ;
  assign n14585 = x1092 | n9190 ;
  assign n14586 = ( n9190 & ~n14584 ) | ( n9190 & n14585 ) | ( ~n14584 & n14585 ) ;
  assign n14587 = ~n4798 & n14478 ;
  assign n14588 = ( x829 & n14586 ) | ( x829 & ~n14587 ) | ( n14586 & ~n14587 ) ;
  assign n14589 = ~x829 & x1093 ;
  assign n14590 = ~n1287 & n14589 ;
  assign n14591 = ( x1092 & n5949 ) | ( x1092 & n14590 ) | ( n5949 & n14590 ) ;
  assign n14592 = n5949 & n14590 ;
  assign n14593 = ( ~n14584 & n14591 ) | ( ~n14584 & n14592 ) | ( n14591 & n14592 ) ;
  assign n14594 = n14581 | n14593 ;
  assign n14595 = ( n14581 & n14588 ) | ( n14581 & n14594 ) | ( n14588 & n14594 ) ;
  assign n14596 = x120 | x1091 ;
  assign n14597 = ~n14468 & n14596 ;
  assign n14598 = x120 & ~n14468 ;
  assign n14599 = ( n14595 & n14597 ) | ( n14595 & n14598 ) | ( n14597 & n14598 ) ;
  assign n14600 = ( x1093 & n4983 ) | ( x1093 & ~n14478 ) | ( n4983 & ~n14478 ) ;
  assign n14601 = n14586 & n14600 ;
  assign n14602 = x120 & ~x1091 ;
  assign n14603 = ~n14468 & n14602 ;
  assign n14604 = ( ~n14469 & n14601 ) | ( ~n14469 & n14603 ) | ( n14601 & n14603 ) ;
  assign n14605 = n14580 & n14604 ;
  assign n14606 = ( n14580 & n14599 ) | ( n14580 & n14605 ) | ( n14599 & n14605 ) ;
  assign n14607 = x681 | n14606 ;
  assign n14608 = ~n4713 & n14604 ;
  assign n14609 = ( ~n4713 & n14599 ) | ( ~n4713 & n14608 ) | ( n14599 & n14608 ) ;
  assign n14610 = n4708 | n14517 ;
  assign n14611 = n14609 | n14610 ;
  assign n14612 = n4708 & ~n14604 ;
  assign n14613 = ~n14599 & n14612 ;
  assign n14614 = n14611 & ~n14613 ;
  assign n14615 = ~x681 & n14580 ;
  assign n14616 = ~n14606 & n14615 ;
  assign n14617 = ( n14607 & n14614 ) | ( n14607 & ~n14616 ) | ( n14614 & ~n14616 ) ;
  assign n14618 = x681 & n14613 ;
  assign n14619 = ( x681 & ~n14611 ) | ( x681 & n14618 ) | ( ~n14611 & n14618 ) ;
  assign n14620 = n14450 & n14619 ;
  assign n14621 = ( n14450 & ~n14617 ) | ( n14450 & n14620 ) | ( ~n14617 & n14620 ) ;
  assign n14622 = n4718 | n14621 ;
  assign n14623 = n4713 & ~n14604 ;
  assign n14624 = ~n14599 & n14623 ;
  assign n14625 = x614 & n1290 ;
  assign n14626 = n14553 & n14625 ;
  assign n14627 = ~n14481 & n14626 ;
  assign n14628 = x614 & ~x662 ;
  assign n14629 = ~n4710 & n14628 ;
  assign n14630 = n14544 & n14629 ;
  assign n14631 = x680 & n14629 ;
  assign n14632 = ( ~n14481 & n14630 ) | ( ~n14481 & n14631 ) | ( n14630 & n14631 ) ;
  assign n14633 = ~n14533 & n14632 ;
  assign n14634 = n14627 | n14633 ;
  assign n14635 = ~x680 & n14631 ;
  assign n14636 = ~x680 & n14630 ;
  assign n14637 = ( ~n14481 & n14635 ) | ( ~n14481 & n14636 ) | ( n14635 & n14636 ) ;
  assign n14638 = n14627 | n14637 ;
  assign n14639 = ( ~n14624 & n14634 ) | ( ~n14624 & n14638 ) | ( n14634 & n14638 ) ;
  assign n14640 = x681 | n14639 ;
  assign n14641 = n14490 & ~n14624 ;
  assign n14642 = x603 | n1290 ;
  assign n14643 = ( x603 & ~n14481 ) | ( x603 & n14642 ) | ( ~n14481 & n14642 ) ;
  assign n14644 = x603 & ~n14482 ;
  assign n14645 = x603 & ~n4713 ;
  assign n14646 = ( n14481 & n14644 ) | ( n14481 & n14645 ) | ( n14644 & n14645 ) ;
  assign n14647 = n14643 & ~n14646 ;
  assign n14648 = x642 | n14647 ;
  assign n14649 = ~x603 & n14642 ;
  assign n14650 = ~n14481 & n14649 ;
  assign n14651 = x642 | n14650 ;
  assign n14652 = ( ~n14624 & n14648 ) | ( ~n14624 & n14651 ) | ( n14648 & n14651 ) ;
  assign n14653 = x614 | n4711 ;
  assign n14654 = ( x616 & ~n14554 ) | ( x616 & n14653 ) | ( ~n14554 & n14653 ) ;
  assign n14655 = x616 | n14653 ;
  assign n14656 = ( n14481 & n14654 ) | ( n14481 & n14655 ) | ( n14654 & n14655 ) ;
  assign n14657 = ~x616 & n14486 ;
  assign n14658 = ( x616 & ~n14656 ) | ( x616 & n14657 ) | ( ~n14656 & n14657 ) ;
  assign n14659 = x616 & ~n14656 ;
  assign n14660 = ( n14652 & n14658 ) | ( n14652 & n14659 ) | ( n14658 & n14659 ) ;
  assign n14661 = ~x614 & n4711 ;
  assign n14662 = n14658 | n14661 ;
  assign n14663 = n14659 | n14661 ;
  assign n14664 = ( n14652 & n14662 ) | ( n14652 & n14663 ) | ( n14662 & n14663 ) ;
  assign n14665 = ( n14641 & n14660 ) | ( n14641 & n14664 ) | ( n14660 & n14664 ) ;
  assign n14666 = n14640 | n14665 ;
  assign n14667 = ( x614 & n14481 ) | ( x614 & n14496 ) | ( n14481 & n14496 ) ;
  assign n14668 = x614 | n14485 ;
  assign n14669 = x614 | n4706 ;
  assign n14670 = ( ~n14481 & n14668 ) | ( ~n14481 & n14669 ) | ( n14668 & n14669 ) ;
  assign n14671 = ~n14667 & n14670 ;
  assign n14672 = x616 | n14671 ;
  assign n14673 = ~n14494 & n14672 ;
  assign n14674 = x614 & ~n14496 ;
  assign n14675 = x616 | n14674 ;
  assign n14676 = ( x616 & ~n14481 ) | ( x616 & n14675 ) | ( ~n14481 & n14675 ) ;
  assign n14677 = ~n14494 & n14676 ;
  assign n14678 = ( n14652 & n14673 ) | ( n14652 & n14677 ) | ( n14673 & n14677 ) ;
  assign n14679 = x681 & ~n14678 ;
  assign n14680 = ~n14450 & n14679 ;
  assign n14681 = ( n14450 & n14666 ) | ( n14450 & ~n14680 ) | ( n14666 & ~n14680 ) ;
  assign n14682 = ~n14622 & n14681 ;
  assign n14683 = n4718 & ~n14619 ;
  assign n14684 = n14617 & n14683 ;
  assign n14685 = n1290 & ~n2203 ;
  assign n14686 = x215 | n14685 ;
  assign n14687 = ( x215 & ~n14481 ) | ( x215 & n14686 ) | ( ~n14481 & n14686 ) ;
  assign n14688 = n2203 | n14687 ;
  assign n14689 = ( n14684 & n14687 ) | ( n14684 & n14688 ) | ( n14687 & n14688 ) ;
  assign n14690 = n2203 | n14689 ;
  assign n14691 = ( n14682 & n14689 ) | ( n14682 & n14690 ) | ( n14689 & n14690 ) ;
  assign n14692 = ( x299 & n14579 ) | ( x299 & ~n14691 ) | ( n14579 & ~n14691 ) ;
  assign n14693 = ~n4764 & n14679 ;
  assign n14694 = ( n4764 & n14666 ) | ( n4764 & ~n14693 ) | ( n14666 & ~n14693 ) ;
  assign n14695 = n4764 & n14619 ;
  assign n14696 = ( n4764 & ~n14617 ) | ( n4764 & n14695 ) | ( ~n14617 & n14695 ) ;
  assign n14697 = n1823 & ~n14696 ;
  assign n14698 = n14694 & n14697 ;
  assign n14699 = n1290 & ~n1823 ;
  assign n14700 = x223 | n14699 ;
  assign n14701 = ( x223 & ~n14481 ) | ( x223 & n14700 ) | ( ~n14481 & n14700 ) ;
  assign n14702 = n14698 | n14701 ;
  assign n14703 = n4764 & ~n14528 ;
  assign n14704 = ~n4764 & n14571 ;
  assign n14705 = ( n4764 & n14570 ) | ( n4764 & ~n14704 ) | ( n14570 & ~n14704 ) ;
  assign n14706 = x223 & ~n14705 ;
  assign n14707 = ( x223 & n14703 ) | ( x223 & n14706 ) | ( n14703 & n14706 ) ;
  assign n14708 = ~x299 & n14707 ;
  assign n14709 = ( x299 & n14702 ) | ( x299 & ~n14708 ) | ( n14702 & ~n14708 ) ;
  assign n14710 = ~n14692 & n14709 ;
  assign n14711 = n1323 | n1527 ;
  assign n14712 = x314 & n8425 ;
  assign n14713 = ~n1242 & n14712 ;
  assign n14714 = ~n14711 & n14713 ;
  assign n14715 = x40 | n8403 ;
  assign n14716 = n1244 | n10299 ;
  assign n14717 = ~x102 & n9436 ;
  assign n14718 = ( x102 & n9439 ) | ( x102 & ~n14717 ) | ( n9439 & ~n14717 ) ;
  assign n14719 = ~n14716 & n14718 ;
  assign n14720 = ~x47 & n7129 ;
  assign n14721 = x81 & x102 ;
  assign n14722 = x102 | n14721 ;
  assign n14723 = x98 | n14722 ;
  assign n14724 = ( x64 & x102 ) | ( x64 & n14721 ) | ( x102 & n14721 ) ;
  assign n14725 = x98 | n14724 ;
  assign n14726 = ( n1241 & n14723 ) | ( n1241 & n14725 ) | ( n14723 & n14725 ) ;
  assign n14727 = ( ~x47 & n14720 ) | ( ~x47 & n14726 ) | ( n14720 & n14726 ) ;
  assign n14728 = x47 & ~n14720 ;
  assign n14729 = ( n14719 & ~n14727 ) | ( n14719 & n14728 ) | ( ~n14727 & n14728 ) ;
  assign n14730 = n14715 | n14729 ;
  assign n14731 = n14711 & ~n14715 ;
  assign n14732 = ( n14714 & n14730 ) | ( n14714 & ~n14731 ) | ( n14730 & ~n14731 ) ;
  assign n14733 = x252 & ~n1299 ;
  assign n14734 = ( ~x35 & n14715 ) | ( ~x35 & n14733 ) | ( n14715 & n14733 ) ;
  assign n14735 = n14715 & n14733 ;
  assign n14736 = ( ~n14732 & n14734 ) | ( ~n14732 & n14735 ) | ( n14734 & n14735 ) ;
  assign n14737 = ~x252 & n8462 ;
  assign n14738 = ~x40 & n7396 ;
  assign n14739 = ( ~x40 & n7130 ) | ( ~x40 & n14738 ) | ( n7130 & n14738 ) ;
  assign n14740 = ( ~x40 & n14726 ) | ( ~x40 & n14739 ) | ( n14726 & n14739 ) ;
  assign n14741 = x40 & ~n14739 ;
  assign n14742 = ( n14719 & ~n14740 ) | ( n14719 & n14741 ) | ( ~n14740 & n14741 ) ;
  assign n14743 = ( x252 & ~n14737 ) | ( x252 & n14742 ) | ( ~n14737 & n14742 ) ;
  assign n14744 = ~n1863 & n14743 ;
  assign n14745 = x1092 & n1690 ;
  assign n14746 = n1287 & n14745 ;
  assign n14747 = n1288 | n14746 ;
  assign n14748 = ( n1288 & n14744 ) | ( n1288 & n14747 ) | ( n14744 & n14747 ) ;
  assign n14749 = n1288 & n14747 ;
  assign n14750 = ( ~n14736 & n14748 ) | ( ~n14736 & n14749 ) | ( n14748 & n14749 ) ;
  assign n14751 = n1287 & n14750 ;
  assign n14752 = n5950 & ~n8462 ;
  assign n14753 = x88 | n14718 ;
  assign n14754 = ( x88 & ~n14726 ) | ( x88 & n14753 ) | ( ~n14726 & n14753 ) ;
  assign n14755 = x252 | n7513 ;
  assign n14756 = n7170 | n14755 ;
  assign n14757 = n9179 | n14756 ;
  assign n14758 = ~x40 & n14757 ;
  assign n14759 = ( x40 & n14754 ) | ( x40 & ~n14758 ) | ( n14754 & ~n14758 ) ;
  assign n14760 = n14752 & n14759 ;
  assign n14761 = x47 | n14713 ;
  assign n14762 = ~n14711 & n14761 ;
  assign n14763 = x252 & ~n8403 ;
  assign n14764 = n1311 | n9178 ;
  assign n14765 = n1311 | n9177 ;
  assign n14766 = ( n1241 & n14764 ) | ( n1241 & n14765 ) | ( n14764 & n14765 ) ;
  assign n14767 = n14726 | n14766 ;
  assign n14768 = x88 & ~n14766 ;
  assign n14769 = ( n14753 & ~n14767 ) | ( n14753 & n14768 ) | ( ~n14767 & n14768 ) ;
  assign n14770 = x35 & x252 ;
  assign n14771 = ~n8403 & n14770 ;
  assign n14772 = ( n14763 & n14769 ) | ( n14763 & n14771 ) | ( n14769 & n14771 ) ;
  assign n14773 = ( ~n14711 & n14763 ) | ( ~n14711 & n14771 ) | ( n14763 & n14771 ) ;
  assign n14774 = ( n14762 & n14772 ) | ( n14762 & n14773 ) | ( n14772 & n14773 ) ;
  assign n14775 = ( n14752 & n14760 ) | ( n14752 & n14774 ) | ( n14760 & n14774 ) ;
  assign n14776 = x1093 & n14775 ;
  assign n14777 = x1092 & ~n10310 ;
  assign n14778 = n14744 & n14777 ;
  assign n14779 = ~n14736 & n14778 ;
  assign n14780 = ( x1093 & n14776 ) | ( x1093 & n14779 ) | ( n14776 & n14779 ) ;
  assign n14781 = ( n14750 & n14751 ) | ( n14750 & n14780 ) | ( n14751 & n14780 ) ;
  assign n14782 = ~x1091 & n14780 ;
  assign n14783 = n14781 | n14782 ;
  assign n14784 = x210 | n14783 ;
  assign n14785 = ~n2134 & n14759 ;
  assign n14786 = ( ~n2134 & n14774 ) | ( ~n2134 & n14785 ) | ( n14774 & n14785 ) ;
  assign n14787 = x32 & ~n1271 ;
  assign n14788 = ~n1242 & n14787 ;
  assign n14789 = ~x95 & n1692 ;
  assign n14790 = ( x32 & n4910 ) | ( x32 & ~n14789 ) | ( n4910 & ~n14789 ) ;
  assign n14791 = x32 & ~n14790 ;
  assign n14792 = ~x32 & n14789 ;
  assign n14793 = x32 & n14792 ;
  assign n14794 = ( n14788 & n14791 ) | ( n14788 & n14793 ) | ( n14791 & n14793 ) ;
  assign n14795 = x824 & n14794 ;
  assign n14796 = ( n14788 & ~n14790 ) | ( n14788 & n14792 ) | ( ~n14790 & n14792 ) ;
  assign n14797 = x824 & n14796 ;
  assign n14798 = ( n14786 & n14795 ) | ( n14786 & n14797 ) | ( n14795 & n14797 ) ;
  assign n14799 = n14779 | n14798 ;
  assign n14800 = x32 | n14743 ;
  assign n14801 = ~x824 & x829 ;
  assign n14802 = ~n14790 & n14801 ;
  assign n14803 = n14792 & n14801 ;
  assign n14804 = ( n14788 & n14802 ) | ( n14788 & n14803 ) | ( n14802 & n14803 ) ;
  assign n14805 = n14800 & n14804 ;
  assign n14806 = x32 & n14804 ;
  assign n14807 = ( ~n14736 & n14805 ) | ( ~n14736 & n14806 ) | ( n14805 & n14806 ) ;
  assign n14808 = x1093 & n14807 ;
  assign n14809 = ( x1093 & n14799 ) | ( x1093 & n14808 ) | ( n14799 & n14808 ) ;
  assign n14810 = ( n14750 & n14751 ) | ( n14750 & n14809 ) | ( n14751 & n14809 ) ;
  assign n14811 = x210 & ~n5995 ;
  assign n14812 = ( x210 & ~n14799 ) | ( x210 & n14811 ) | ( ~n14799 & n14811 ) ;
  assign n14813 = ~n14810 & n14812 ;
  assign n14814 = n14784 & ~n14813 ;
  assign n14815 = x299 & ~n14814 ;
  assign n14816 = x198 | n14783 ;
  assign n14817 = x198 & ~n5995 ;
  assign n14818 = ( x198 & ~n14799 ) | ( x198 & n14817 ) | ( ~n14799 & n14817 ) ;
  assign n14819 = ~n14810 & n14818 ;
  assign n14820 = n14816 & ~n14819 ;
  assign n14821 = x299 | n14820 ;
  assign n14822 = ~n14815 & n14821 ;
  assign n14823 = ~x39 & n14822 ;
  assign n14824 = n1290 & ~n4658 ;
  assign n14825 = ~n1494 & n14824 ;
  assign n14826 = ~n1271 & n14825 ;
  assign n14827 = ~n1242 & n14826 ;
  assign n14828 = ( n2032 & n12808 ) | ( n2032 & ~n14827 ) | ( n12808 & ~n14827 ) ;
  assign n14829 = x38 & ~n2032 ;
  assign n14830 = n14827 & n14829 ;
  assign n14831 = ( n14823 & ~n14828 ) | ( n14823 & n14830 ) | ( ~n14828 & n14830 ) ;
  assign n14832 = x39 | n14822 ;
  assign n14833 = ( ~n14828 & n14830 ) | ( ~n14828 & n14832 ) | ( n14830 & n14832 ) ;
  assign n14834 = ( n14710 & n14831 ) | ( n14710 & n14833 ) | ( n14831 & n14833 ) ;
  assign n14835 = x140 | n14834 ;
  assign n14836 = ( x626 & x1158 ) | ( x626 & ~n14835 ) | ( x1158 & ~n14835 ) ;
  assign n14837 = x140 & n2032 ;
  assign n14838 = x621 & x1091 ;
  assign n14839 = x603 & ~n14838 ;
  assign n14840 = n1290 & n14839 ;
  assign n14841 = ~x215 & n2203 ;
  assign n14842 = ( x215 & n14840 ) | ( x215 & ~n14841 ) | ( n14840 & ~n14841 ) ;
  assign n14843 = x215 & ~n14841 ;
  assign n14844 = ( ~n14481 & n14842 ) | ( ~n14481 & n14843 ) | ( n14842 & n14843 ) ;
  assign n14845 = ~n4711 & n14613 ;
  assign n14846 = ( n4711 & n14611 ) | ( n4711 & ~n14845 ) | ( n14611 & ~n14845 ) ;
  assign n14847 = n4711 & ~n14604 ;
  assign n14848 = ~n14599 & n14847 ;
  assign n14849 = n14839 & ~n14848 ;
  assign n14850 = n4721 & ~n14849 ;
  assign n14851 = ( n4721 & ~n14846 ) | ( n4721 & n14850 ) | ( ~n14846 & n14850 ) ;
  assign n14852 = ~n14844 & n14851 ;
  assign n14853 = n2203 & n4721 ;
  assign n14854 = x614 | x642 ;
  assign n14855 = x616 | n14854 ;
  assign n14856 = n14840 & n14855 ;
  assign n14857 = ~n14481 & n14856 ;
  assign n14858 = n4713 & n14839 ;
  assign n14859 = ~n14855 & n14858 ;
  assign n14860 = n14482 & n14839 ;
  assign n14861 = ~n14855 & n14860 ;
  assign n14862 = ( ~n14481 & n14859 ) | ( ~n14481 & n14861 ) | ( n14859 & n14861 ) ;
  assign n14863 = n14857 | n14862 ;
  assign n14864 = ~n4711 & n14863 ;
  assign n14865 = ~n4711 & n14857 ;
  assign n14866 = ( ~n14624 & n14864 ) | ( ~n14624 & n14865 ) | ( n14864 & n14865 ) ;
  assign n14867 = ( ~n14481 & n14858 ) | ( ~n14481 & n14860 ) | ( n14858 & n14860 ) ;
  assign n14868 = n4711 & n14867 ;
  assign n14869 = ~n14624 & n14868 ;
  assign n14870 = n14866 | n14869 ;
  assign n14871 = ( n2203 & n14853 ) | ( n2203 & n14870 ) | ( n14853 & n14870 ) ;
  assign n14872 = n4721 & ~n14517 ;
  assign n14873 = ~n14510 & n14872 ;
  assign n14874 = ~n14481 & n14840 ;
  assign n14875 = n14517 & n14874 ;
  assign n14876 = ( n14510 & n14874 ) | ( n14510 & n14875 ) | ( n14874 & n14875 ) ;
  assign n14877 = n4713 & ~n14855 ;
  assign n14878 = ~n14465 & n14877 ;
  assign n14879 = ~n14474 & n14878 ;
  assign n14880 = n4711 | n14879 ;
  assign n14881 = n14876 & ~n14880 ;
  assign n14882 = ~n4713 & n14840 ;
  assign n14883 = ~n14481 & n14882 ;
  assign n14884 = ( n14475 & n14874 ) | ( n14475 & n14883 ) | ( n14874 & n14883 ) ;
  assign n14885 = ~n14873 & n14884 ;
  assign n14886 = ( ~n14873 & n14881 ) | ( ~n14873 & n14885 ) | ( n14881 & n14885 ) ;
  assign n14887 = ( x299 & n4343 ) | ( x299 & n14886 ) | ( n4343 & n14886 ) ;
  assign n14888 = n14871 & n14887 ;
  assign n14889 = n14844 & n14887 ;
  assign n14890 = ( ~n14852 & n14888 ) | ( ~n14852 & n14889 ) | ( n14888 & n14889 ) ;
  assign n14891 = n14699 & n14839 ;
  assign n14892 = x223 | n14891 ;
  assign n14893 = ( x223 & ~n14481 ) | ( x223 & n14892 ) | ( ~n14481 & n14892 ) ;
  assign n14894 = n4764 & ~n14849 ;
  assign n14895 = ( n4764 & ~n14846 ) | ( n4764 & n14894 ) | ( ~n14846 & n14894 ) ;
  assign n14896 = ~n14893 & n14895 ;
  assign n14897 = n1823 & n4764 ;
  assign n14898 = ( n1823 & n14870 ) | ( n1823 & n14897 ) | ( n14870 & n14897 ) ;
  assign n14899 = n4764 & ~n14517 ;
  assign n14900 = ~n14510 & n14899 ;
  assign n14901 = n14884 & ~n14900 ;
  assign n14902 = ( n14881 & ~n14900 ) | ( n14881 & n14901 ) | ( ~n14900 & n14901 ) ;
  assign n14903 = ( x299 & n2213 ) | ( x299 & ~n14902 ) | ( n2213 & ~n14902 ) ;
  assign n14904 = n14898 & ~n14903 ;
  assign n14905 = n14893 & ~n14903 ;
  assign n14906 = ( ~n14896 & n14904 ) | ( ~n14896 & n14905 ) | ( n14904 & n14905 ) ;
  assign n14907 = n14890 | n14906 ;
  assign n14908 = x39 & ~n14907 ;
  assign n14910 = x621 & ~n5995 ;
  assign n14911 = ( x621 & ~n14799 ) | ( x621 & n14910 ) | ( ~n14799 & n14910 ) ;
  assign n14909 = n5995 & n14799 ;
  assign n14912 = n14909 & ~n14911 ;
  assign n14913 = ( n14810 & ~n14911 ) | ( n14810 & n14912 ) | ( ~n14911 & n14912 ) ;
  assign n14914 = x210 & ~n14913 ;
  assign n14915 = ~x210 & n14838 ;
  assign n14916 = ~x210 & x621 ;
  assign n14917 = ( ~n14780 & n14915 ) | ( ~n14780 & n14916 ) | ( n14915 & n14916 ) ;
  assign n14918 = ( x210 & n14783 ) | ( x210 & ~n14917 ) | ( n14783 & ~n14917 ) ;
  assign n14919 = x603 & n14918 ;
  assign n14920 = ~n14914 & n14919 ;
  assign n14921 = x299 & ~n14920 ;
  assign n14922 = x198 & n14913 ;
  assign n14923 = x198 | x621 ;
  assign n14924 = x198 | n14838 ;
  assign n14925 = ( ~n14780 & n14923 ) | ( ~n14780 & n14924 ) | ( n14923 & n14924 ) ;
  assign n14926 = x603 & ~n14925 ;
  assign n14927 = n14783 & n14926 ;
  assign n14928 = x299 | n14927 ;
  assign n14929 = x299 | x603 ;
  assign n14930 = ( n14922 & n14928 ) | ( n14922 & n14929 ) | ( n14928 & n14929 ) ;
  assign n14931 = x39 | n14930 ;
  assign n14932 = ( x39 & ~n14921 ) | ( x39 & n14931 ) | ( ~n14921 & n14931 ) ;
  assign n14933 = ~n14908 & n14932 ;
  assign n14934 = x140 & ~x761 ;
  assign n14935 = n14933 & n14934 ;
  assign n14936 = ( n14710 & n14823 ) | ( n14710 & n14832 ) | ( n14823 & n14832 ) ;
  assign n14937 = ( x140 & x761 ) | ( x140 & n14936 ) | ( x761 & n14936 ) ;
  assign n14938 = x621 & n14751 ;
  assign n14939 = x621 & n14750 ;
  assign n14940 = ( n14809 & n14938 ) | ( n14809 & n14939 ) | ( n14938 & n14939 ) ;
  assign n14941 = x210 & ~n14940 ;
  assign n14942 = x210 | x621 ;
  assign n14943 = ( x210 & n14781 ) | ( x210 & n14942 ) | ( n14781 & n14942 ) ;
  assign n14944 = x603 & ~n14943 ;
  assign n14945 = ( x603 & n14941 ) | ( x603 & n14944 ) | ( n14941 & n14944 ) ;
  assign n14946 = n14814 & ~n14945 ;
  assign n14947 = x299 & ~n14946 ;
  assign n14948 = x603 | n14925 ;
  assign n14949 = n14783 & ~n14948 ;
  assign n14950 = ( ~x603 & n14922 ) | ( ~x603 & n14949 ) | ( n14922 & n14949 ) ;
  assign n14951 = x198 & ~n14940 ;
  assign n14952 = ( x198 & n14781 ) | ( x198 & n14923 ) | ( n14781 & n14923 ) ;
  assign n14953 = ~n14951 & n14952 ;
  assign n14954 = x299 | n14953 ;
  assign n14955 = n14950 | n14954 ;
  assign n14956 = ~n14947 & n14955 ;
  assign n14957 = x39 | n14956 ;
  assign n14958 = x215 & ~n4721 ;
  assign n14959 = n1290 & ~n14839 ;
  assign n14960 = n14517 & n14959 ;
  assign n14961 = ( n14510 & n14959 ) | ( n14510 & n14960 ) | ( n14959 & n14960 ) ;
  assign n14962 = ( ~n4708 & n14465 ) | ( ~n4708 & n14961 ) | ( n14465 & n14961 ) ;
  assign n14963 = n14465 & n14959 ;
  assign n14964 = ( n14474 & n14959 ) | ( n14474 & n14963 ) | ( n14959 & n14963 ) ;
  assign n14965 = n4711 & ~n14964 ;
  assign n14966 = n4711 & n14964 ;
  assign n14967 = ( n14961 & ~n14965 ) | ( n14961 & n14966 ) | ( ~n14965 & n14966 ) ;
  assign n14968 = ~n14965 & n14966 ;
  assign n14969 = ( n14962 & n14967 ) | ( n14962 & n14968 ) | ( n14967 & n14968 ) ;
  assign n14970 = ( x215 & n14958 ) | ( x215 & n14969 ) | ( n14958 & n14969 ) ;
  assign n14971 = n1290 & n14838 ;
  assign n14972 = n4713 | n14971 ;
  assign n14973 = x603 & ~n14972 ;
  assign n14974 = ( n14481 & n14645 ) | ( n14481 & n14973 ) | ( n14645 & n14973 ) ;
  assign n14975 = ~x621 & n4713 ;
  assign n14976 = ( n4713 & ~n14465 ) | ( n4713 & n14975 ) | ( ~n14465 & n14975 ) ;
  assign n14977 = ( x603 & n14974 ) | ( x603 & n14976 ) | ( n14974 & n14976 ) ;
  assign n14978 = n4711 & n14484 ;
  assign n14979 = n4711 & n14490 ;
  assign n14980 = ( n14475 & n14978 ) | ( n14475 & n14979 ) | ( n14978 & n14979 ) ;
  assign n14981 = ~n14977 & n14980 ;
  assign n14982 = n14855 & n14959 ;
  assign n14983 = ~n14481 & n14982 ;
  assign n14984 = n14642 & ~n14855 ;
  assign n14985 = x603 & ~n14855 ;
  assign n14986 = ( ~n14481 & n14984 ) | ( ~n14481 & n14985 ) | ( n14984 & n14985 ) ;
  assign n14987 = n14983 | n14986 ;
  assign n14988 = ( ~n14977 & n14983 ) | ( ~n14977 & n14987 ) | ( n14983 & n14987 ) ;
  assign n14989 = ~n4711 & n14988 ;
  assign n14990 = n14981 | n14989 ;
  assign n14991 = n4721 | n14990 ;
  assign n14992 = n14970 & n14991 ;
  assign n14993 = x215 & ~n14992 ;
  assign n14994 = ~n2203 & n14959 ;
  assign n14995 = ~n14481 & n14994 ;
  assign n14996 = ( n14992 & ~n14993 ) | ( n14992 & n14995 ) | ( ~n14993 & n14995 ) ;
  assign n14997 = n14846 & ~n14848 ;
  assign n14998 = ( x603 & ~n14516 ) | ( x603 & n14839 ) | ( ~n14516 & n14839 ) ;
  assign n14999 = ( x603 & n14481 ) | ( x603 & n14998 ) | ( n14481 & n14998 ) ;
  assign n15000 = x120 & n14838 ;
  assign n15001 = ~n14468 & n15000 ;
  assign n15002 = ~n4713 & n15001 ;
  assign n15003 = n14596 & n14838 ;
  assign n15004 = ~n14468 & n15003 ;
  assign n15005 = ~n4713 & n15004 ;
  assign n15006 = ( n14595 & n15002 ) | ( n14595 & n15005 ) | ( n15002 & n15005 ) ;
  assign n15007 = n14999 & ~n15006 ;
  assign n15008 = x603 | n14517 ;
  assign n15009 = n14609 | n15008 ;
  assign n15010 = ~n15007 & n15009 ;
  assign n15011 = ( n14595 & n15001 ) | ( n14595 & n15004 ) | ( n15001 & n15004 ) ;
  assign n15012 = x603 & ~n15001 ;
  assign n15013 = x603 & ~n15004 ;
  assign n15014 = ( ~n14595 & n15012 ) | ( ~n14595 & n15013 ) | ( n15012 & n15013 ) ;
  assign n15015 = x621 & ~n14603 ;
  assign n15016 = x621 & n14469 ;
  assign n15017 = ( ~n14601 & n15015 ) | ( ~n14601 & n15016 ) | ( n15015 & n15016 ) ;
  assign n15018 = n14604 & ~n15017 ;
  assign n15019 = ( n14599 & ~n15017 ) | ( n14599 & n15018 ) | ( ~n15017 & n15018 ) ;
  assign n15020 = ( n15011 & ~n15014 ) | ( n15011 & n15019 ) | ( ~n15014 & n15019 ) ;
  assign n15021 = n15010 | n15020 ;
  assign n15022 = n14997 & n15021 ;
  assign n15023 = n2203 & ~n4721 ;
  assign n15024 = n4713 & ~n15001 ;
  assign n15025 = n4713 & ~n15004 ;
  assign n15026 = ( ~n14595 & n15024 ) | ( ~n14595 & n15025 ) | ( n15024 & n15025 ) ;
  assign n15027 = ( x603 & n14974 ) | ( x603 & n15026 ) | ( n14974 & n15026 ) ;
  assign n15028 = n4711 & n15027 ;
  assign n15029 = ( n4711 & ~n14641 ) | ( n4711 & n15028 ) | ( ~n14641 & n15028 ) ;
  assign n15030 = n4711 | n14982 ;
  assign n15031 = ( n4711 & ~n14481 ) | ( n4711 & n15030 ) | ( ~n14481 & n15030 ) ;
  assign n15032 = ~n14974 & n14986 ;
  assign n15033 = ~x603 & n14986 ;
  assign n15034 = ( ~n15026 & n15032 ) | ( ~n15026 & n15033 ) | ( n15032 & n15033 ) ;
  assign n15035 = n15031 | n15034 ;
  assign n15036 = n4721 | n15035 ;
  assign n15037 = ( n4721 & ~n15029 ) | ( n4721 & n15036 ) | ( ~n15029 & n15036 ) ;
  assign n15038 = n15023 & n15037 ;
  assign n15039 = n2203 & n15037 ;
  assign n15040 = ( n15022 & n15038 ) | ( n15022 & n15039 ) | ( n15038 & n15039 ) ;
  assign n15041 = x299 & n15040 ;
  assign n15042 = x299 & ~n14993 ;
  assign n15043 = ( n14996 & n15041 ) | ( n14996 & n15042 ) | ( n15041 & n15042 ) ;
  assign n15044 = x223 & ~n4764 ;
  assign n15045 = ( x223 & n14969 ) | ( x223 & n15044 ) | ( n14969 & n15044 ) ;
  assign n15046 = n4764 | n14990 ;
  assign n15047 = n15045 & n15046 ;
  assign n15048 = x223 & ~n15047 ;
  assign n15049 = ~n1823 & n14959 ;
  assign n15050 = ~n14481 & n15049 ;
  assign n15051 = ( n15047 & ~n15048 ) | ( n15047 & n15050 ) | ( ~n15048 & n15050 ) ;
  assign n15052 = n1823 & ~n4764 ;
  assign n15053 = n4764 | n15035 ;
  assign n15054 = ( n4764 & ~n15029 ) | ( n4764 & n15053 ) | ( ~n15029 & n15053 ) ;
  assign n15055 = n15052 & n15054 ;
  assign n15056 = n1823 & n15054 ;
  assign n15057 = ( n15022 & n15055 ) | ( n15022 & n15056 ) | ( n15055 & n15056 ) ;
  assign n15058 = ~x299 & n15057 ;
  assign n15059 = x299 | n15048 ;
  assign n15060 = ( n15051 & n15058 ) | ( n15051 & ~n15059 ) | ( n15058 & ~n15059 ) ;
  assign n15061 = n15043 | n15060 ;
  assign n15062 = x39 & ~n15061 ;
  assign n15063 = n14957 & ~n15062 ;
  assign n15064 = ( x140 & ~x761 ) | ( x140 & n15063 ) | ( ~x761 & n15063 ) ;
  assign n15065 = n14937 | n15064 ;
  assign n15066 = ~n14935 & n15065 ;
  assign n15067 = x38 | n15066 ;
  assign n15068 = n1290 & ~n4809 ;
  assign n15069 = ~n1271 & n15068 ;
  assign n15070 = ~n1242 & n15069 ;
  assign n15071 = x140 | n15070 ;
  assign n15072 = ~n4810 & n14840 ;
  assign n15073 = ~x761 & n15072 ;
  assign n15074 = n15071 & ~n15073 ;
  assign n15075 = x38 & ~n15074 ;
  assign n15076 = n15067 & ~n15075 ;
  assign n15077 = ~n2032 & n15076 ;
  assign n15078 = n14837 | n15077 ;
  assign n15079 = ~x608 & x1153 ;
  assign n15080 = x608 & ~x1153 ;
  assign n15081 = n15079 | n15080 ;
  assign n15082 = x778 & n15081 ;
  assign n15083 = n15078 & ~n15082 ;
  assign n15084 = n14835 & n15082 ;
  assign n15085 = n15083 | n15084 ;
  assign n15086 = ~x785 & n15085 ;
  assign n15087 = x609 & ~x778 ;
  assign n15088 = ( x609 & ~n15081 ) | ( x609 & n15087 ) | ( ~n15081 & n15087 ) ;
  assign n15089 = n14835 & ~n15088 ;
  assign n15090 = x609 & n15083 ;
  assign n15091 = n15089 | n15090 ;
  assign n15092 = x1155 & n15091 ;
  assign n15093 = x609 | x778 ;
  assign n15094 = ( x609 & n15081 ) | ( x609 & n15093 ) | ( n15081 & n15093 ) ;
  assign n15095 = n14835 & n15094 ;
  assign n15096 = ~x609 & n15083 ;
  assign n15097 = n15095 | n15096 ;
  assign n15098 = ~x1155 & n15097 ;
  assign n15099 = n15092 | n15098 ;
  assign n15100 = x785 & n15099 ;
  assign n15101 = n15086 | n15100 ;
  assign n15102 = ~x781 & n15101 ;
  assign n15103 = ( x618 & x1154 ) | ( x618 & n14835 ) | ( x1154 & n14835 ) ;
  assign n15104 = ( ~x618 & x1154 ) | ( ~x618 & n15101 ) | ( x1154 & n15101 ) ;
  assign n15105 = n15103 & n15104 ;
  assign n15106 = ( x618 & x1154 ) | ( x618 & ~n14835 ) | ( x1154 & ~n14835 ) ;
  assign n15107 = ( x618 & ~x1154 ) | ( x618 & n15101 ) | ( ~x1154 & n15101 ) ;
  assign n15108 = ~n15106 & n15107 ;
  assign n15109 = n15105 | n15108 ;
  assign n15110 = x781 & n15109 ;
  assign n15111 = n15102 | n15110 ;
  assign n15112 = ~x789 & n15111 ;
  assign n15113 = ( x619 & x1159 ) | ( x619 & n14835 ) | ( x1159 & n14835 ) ;
  assign n15114 = ( ~x619 & x1159 ) | ( ~x619 & n15111 ) | ( x1159 & n15111 ) ;
  assign n15115 = n15113 & n15114 ;
  assign n15116 = ( x619 & x1159 ) | ( x619 & ~n14835 ) | ( x1159 & ~n14835 ) ;
  assign n15117 = ( x619 & ~x1159 ) | ( x619 & n15111 ) | ( ~x1159 & n15111 ) ;
  assign n15118 = ~n15116 & n15117 ;
  assign n15119 = n15115 | n15118 ;
  assign n15120 = x789 & n15119 ;
  assign n15121 = n15112 | n15120 ;
  assign n15122 = ( x626 & ~x1158 ) | ( x626 & n15121 ) | ( ~x1158 & n15121 ) ;
  assign n15123 = ~n14836 & n15122 ;
  assign n15124 = ( x626 & x1158 ) | ( x626 & n14835 ) | ( x1158 & n14835 ) ;
  assign n15125 = ( ~x626 & x1158 ) | ( ~x626 & n15121 ) | ( x1158 & n15121 ) ;
  assign n15126 = n15124 & n15125 ;
  assign n15127 = n15123 | n15126 ;
  assign n15128 = x788 & n15127 ;
  assign n15129 = ~x788 & n15121 ;
  assign n15130 = n15128 | n15129 ;
  assign n15131 = ~x629 & x1156 ;
  assign n15132 = x629 & ~x1156 ;
  assign n15133 = n15131 | n15132 ;
  assign n15134 = x792 & n15133 ;
  assign n15135 = n15130 | n15134 ;
  assign n15136 = ~n14835 & n15134 ;
  assign n15137 = n15135 & ~n15136 ;
  assign n15138 = ~x630 & x1157 ;
  assign n15139 = x630 & ~x1157 ;
  assign n15140 = n15138 | n15139 ;
  assign n15141 = x787 & n15140 ;
  assign n15142 = n15137 & ~n15141 ;
  assign n15143 = n14835 & n15141 ;
  assign n15144 = n15142 | n15143 ;
  assign n15145 = ( x644 & x715 ) | ( x644 & n15144 ) | ( x715 & n15144 ) ;
  assign n15146 = ( ~x644 & x715 ) | ( ~x644 & n14835 ) | ( x715 & n14835 ) ;
  assign n15147 = n15145 & n15146 ;
  assign n15148 = x1160 | n15147 ;
  assign n15149 = x665 & x1091 ;
  assign n15150 = n1290 & ~n15149 ;
  assign n15151 = ~n14481 & n15150 ;
  assign n15152 = x665 & ~n14603 ;
  assign n15153 = x665 & n14469 ;
  assign n15154 = ( ~n14601 & n15152 ) | ( ~n14601 & n15153 ) | ( n15152 & n15153 ) ;
  assign n15155 = n14604 & ~n15154 ;
  assign n15156 = ( n14599 & ~n15154 ) | ( n14599 & n15155 ) | ( ~n15154 & n15155 ) ;
  assign n15157 = n15151 | n15156 ;
  assign n15158 = n14641 & n15157 ;
  assign n15159 = x662 & x680 ;
  assign n15160 = ( x680 & n4710 ) | ( x680 & n15159 ) | ( n4710 & n15159 ) ;
  assign n15161 = ( x680 & n15158 ) | ( x680 & n15160 ) | ( n15158 & n15160 ) ;
  assign n15162 = ~n4708 & n15150 ;
  assign n15163 = n4708 | n15162 ;
  assign n15164 = ( n4708 & ~n14481 ) | ( n4708 & n15163 ) | ( ~n14481 & n15163 ) ;
  assign n15165 = n14553 & ~n15164 ;
  assign n15166 = ~n14481 & n15162 ;
  assign n15167 = n14553 & ~n15166 ;
  assign n15168 = ( ~n15158 & n15165 ) | ( ~n15158 & n15167 ) | ( n15165 & n15167 ) ;
  assign n15169 = n15161 & ~n15168 ;
  assign n15170 = ( n1823 & n14897 ) | ( n1823 & n15169 ) | ( n14897 & n15169 ) ;
  assign n15171 = x680 & ~n15149 ;
  assign n15172 = n14699 & n15171 ;
  assign n15173 = ~n14481 & n15172 ;
  assign n15174 = ~n14613 & n15171 ;
  assign n15175 = n14611 & n15174 ;
  assign n15176 = n4711 | n14553 ;
  assign n15177 = ( n14553 & n15156 ) | ( n14553 & n15176 ) | ( n15156 & n15176 ) ;
  assign n15178 = n4764 & ~n15177 ;
  assign n15179 = n4711 & n15156 ;
  assign n15180 = n4764 & ~n15179 ;
  assign n15181 = ( ~n15175 & n15178 ) | ( ~n15175 & n15180 ) | ( n15178 & n15180 ) ;
  assign n15182 = ~n15173 & n15181 ;
  assign n15183 = ~n4713 & n15150 ;
  assign n15184 = ~n14481 & n15183 ;
  assign n15185 = n15166 | n15184 ;
  assign n15186 = n15151 | n15166 ;
  assign n15187 = ( n14475 & n15185 ) | ( n14475 & n15186 ) | ( n15185 & n15186 ) ;
  assign n15188 = x680 & n15187 ;
  assign n15189 = x223 & x662 ;
  assign n15190 = ( x223 & n4710 ) | ( x223 & n15189 ) | ( n4710 & n15189 ) ;
  assign n15191 = ( x223 & n15184 ) | ( x223 & n15190 ) | ( n15184 & n15190 ) ;
  assign n15192 = ( x223 & n15151 ) | ( x223 & n15190 ) | ( n15151 & n15190 ) ;
  assign n15193 = ( n14475 & n15191 ) | ( n14475 & n15192 ) | ( n15191 & n15192 ) ;
  assign n15194 = ~n14900 & n15193 ;
  assign n15195 = n15188 & n15194 ;
  assign n15196 = x223 & ~n15195 ;
  assign n15197 = ( n15182 & ~n15195 ) | ( n15182 & n15196 ) | ( ~n15195 & n15196 ) ;
  assign n15198 = ( n15173 & n15195 ) | ( n15173 & ~n15196 ) | ( n15195 & ~n15196 ) ;
  assign n15199 = ( n15170 & ~n15197 ) | ( n15170 & n15198 ) | ( ~n15197 & n15198 ) ;
  assign n15200 = ~x299 & n15199 ;
  assign n15201 = n4721 | n15169 ;
  assign n15202 = n1290 & n15171 ;
  assign n15203 = ~n2203 & n15202 ;
  assign n15204 = ~n14481 & n15203 ;
  assign n15205 = ( n2203 & n15023 ) | ( n2203 & n15177 ) | ( n15023 & n15177 ) ;
  assign n15206 = ( n2203 & n15023 ) | ( n2203 & n15179 ) | ( n15023 & n15179 ) ;
  assign n15207 = ( n15175 & n15205 ) | ( n15175 & n15206 ) | ( n15205 & n15206 ) ;
  assign n15208 = n15204 | n15207 ;
  assign n15209 = x215 & x662 ;
  assign n15210 = ( x215 & n4710 ) | ( x215 & n15209 ) | ( n4710 & n15209 ) ;
  assign n15211 = ( x215 & n15184 ) | ( x215 & n15210 ) | ( n15184 & n15210 ) ;
  assign n15212 = ( x215 & n15151 ) | ( x215 & n15210 ) | ( n15151 & n15210 ) ;
  assign n15213 = ( n14475 & n15211 ) | ( n14475 & n15212 ) | ( n15211 & n15212 ) ;
  assign n15214 = ~n14873 & n15213 ;
  assign n15215 = n15188 & n15214 ;
  assign n15216 = x215 & ~n15215 ;
  assign n15217 = ( n15208 & n15215 ) | ( n15208 & ~n15216 ) | ( n15215 & ~n15216 ) ;
  assign n15218 = ( n15204 & n15215 ) | ( n15204 & ~n15216 ) | ( n15215 & ~n15216 ) ;
  assign n15219 = ( n15201 & n15217 ) | ( n15201 & n15218 ) | ( n15217 & n15218 ) ;
  assign n15220 = x299 & n15219 ;
  assign n15221 = n15200 | n15220 ;
  assign n15222 = x140 & n15221 ;
  assign n15223 = x39 & x140 ;
  assign n15224 = n1290 & n15149 ;
  assign n15225 = ~n4708 & n15224 ;
  assign n15226 = x680 & ~n15225 ;
  assign n15227 = ( x680 & n14481 ) | ( x680 & n15226 ) | ( n14481 & n15226 ) ;
  assign n15228 = n4713 | n15224 ;
  assign n15229 = ( n4713 & ~n14481 ) | ( n4713 & n15228 ) | ( ~n14481 & n15228 ) ;
  assign n15230 = n15227 & ~n15229 ;
  assign n15231 = ( ~n4708 & n15227 ) | ( ~n4708 & n15230 ) | ( n15227 & n15230 ) ;
  assign n15232 = x680 & ~n15227 ;
  assign n15233 = n14596 & n15149 ;
  assign n15234 = ~n14468 & n15233 ;
  assign n15235 = n4713 & ~n15234 ;
  assign n15236 = x680 & ~n15235 ;
  assign n15237 = x120 & n15149 ;
  assign n15238 = ~n14468 & n15237 ;
  assign n15239 = n4713 & ~n15238 ;
  assign n15240 = x680 & ~n15239 ;
  assign n15241 = ( n14595 & n15236 ) | ( n14595 & n15240 ) | ( n15236 & n15240 ) ;
  assign n15242 = ( ~n15231 & n15232 ) | ( ~n15231 & n15241 ) | ( n15232 & n15241 ) ;
  assign n15243 = n14553 & n15242 ;
  assign n15244 = ( ~n14595 & n15235 ) | ( ~n14595 & n15239 ) | ( n15235 & n15239 ) ;
  assign n15245 = ( n15227 & n15231 ) | ( n15227 & n15244 ) | ( n15231 & n15244 ) ;
  assign n15246 = n14553 & ~n15245 ;
  assign n15247 = ( n14678 & n15243 ) | ( n14678 & n15246 ) | ( n15243 & n15246 ) ;
  assign n15248 = ( x680 & n14553 ) | ( x680 & ~n15229 ) | ( n14553 & ~n15229 ) ;
  assign n15249 = x680 | n14553 ;
  assign n15250 = ( ~n15241 & n15248 ) | ( ~n15241 & n15249 ) | ( n15248 & n15249 ) ;
  assign n15251 = x680 & ~n15250 ;
  assign n15252 = ( n14678 & ~n15250 ) | ( n14678 & n15251 ) | ( ~n15250 & n15251 ) ;
  assign n15253 = n15247 | n15252 ;
  assign n15254 = n4764 | n15253 ;
  assign n15255 = ~x665 & x680 ;
  assign n15256 = ( x680 & ~n14465 ) | ( x680 & n15255 ) | ( ~n14465 & n15255 ) ;
  assign n15257 = n14516 & n15149 ;
  assign n15258 = ~n4708 & n15257 ;
  assign n15259 = ~n14481 & n15258 ;
  assign n15260 = n15256 & ~n15259 ;
  assign n15261 = x680 & ~n15260 ;
  assign n15262 = ( n14519 & ~n15260 ) | ( n14519 & n15261 ) | ( ~n15260 & n15261 ) ;
  assign n15263 = ( n14521 & ~n15260 ) | ( n14521 & n15261 ) | ( ~n15260 & n15261 ) ;
  assign n15264 = ( n14515 & n15262 ) | ( n14515 & n15263 ) | ( n15262 & n15263 ) ;
  assign n15265 = n4711 & ~n15228 ;
  assign n15266 = n4711 & ~n4713 ;
  assign n15267 = ( n14481 & n15265 ) | ( n14481 & n15266 ) | ( n15265 & n15266 ) ;
  assign n15268 = ~x665 & n4713 ;
  assign n15269 = ( n4713 & ~n14465 ) | ( n4713 & n15268 ) | ( ~n14465 & n15268 ) ;
  assign n15270 = ( n4711 & n15267 ) | ( n4711 & n15269 ) | ( n15267 & n15269 ) ;
  assign n15271 = ( n15227 & n15230 ) | ( n15227 & n15269 ) | ( n15230 & n15269 ) ;
  assign n15272 = n15270 | n15271 ;
  assign n15273 = n4764 & ~n15272 ;
  assign n15274 = n15264 & n15273 ;
  assign n15275 = x680 | n14504 ;
  assign n15276 = x223 & n4764 ;
  assign n15277 = ( x223 & n15272 ) | ( x223 & n15276 ) | ( n15272 & n15276 ) ;
  assign n15278 = x223 | n15276 ;
  assign n15279 = ( ~n15275 & n15277 ) | ( ~n15275 & n15278 ) | ( n15277 & n15278 ) ;
  assign n15280 = ~n15274 & n15279 ;
  assign n15281 = n14699 & ~n15171 ;
  assign n15282 = x223 | n15281 ;
  assign n15283 = ( x223 & ~n14481 ) | ( x223 & n15282 ) | ( ~n14481 & n15282 ) ;
  assign n15284 = ~x680 & n14613 ;
  assign n15285 = ( x680 & n14611 ) | ( x680 & ~n15284 ) | ( n14611 & ~n15284 ) ;
  assign n15286 = ~n14553 & n15234 ;
  assign n15287 = x680 & ~n15286 ;
  assign n15288 = ~n14553 & n15238 ;
  assign n15289 = x680 & ~n15288 ;
  assign n15290 = ( ~n14595 & n15287 ) | ( ~n14595 & n15289 ) | ( n15287 & n15289 ) ;
  assign n15291 = ~n4750 & n15238 ;
  assign n15292 = ~n4750 & n15234 ;
  assign n15293 = ( n14595 & n15291 ) | ( n14595 & n15292 ) | ( n15291 & n15292 ) ;
  assign n15294 = n14553 & n15259 ;
  assign n15295 = ( n14553 & n15293 ) | ( n14553 & n15294 ) | ( n15293 & n15294 ) ;
  assign n15296 = n15290 & ~n15295 ;
  assign n15297 = n4764 & n15296 ;
  assign n15298 = ( n4764 & ~n15285 ) | ( n4764 & n15297 ) | ( ~n15285 & n15297 ) ;
  assign n15299 = n1823 | n15283 ;
  assign n15300 = ( n15283 & ~n15298 ) | ( n15283 & n15299 ) | ( ~n15298 & n15299 ) ;
  assign n15301 = ~n15280 & n15300 ;
  assign n15302 = ~n15280 & n15283 ;
  assign n15303 = ( n15254 & n15301 ) | ( n15254 & n15302 ) | ( n15301 & n15302 ) ;
  assign n15304 = x299 | n15303 ;
  assign n15305 = n4721 | n15253 ;
  assign n15306 = n4721 & ~n15272 ;
  assign n15307 = n15264 & n15306 ;
  assign n15308 = x215 & n4721 ;
  assign n15309 = ( x215 & n15272 ) | ( x215 & n15308 ) | ( n15272 & n15308 ) ;
  assign n15310 = x215 | n15308 ;
  assign n15311 = ( ~n15275 & n15309 ) | ( ~n15275 & n15310 ) | ( n15309 & n15310 ) ;
  assign n15312 = ~n15307 & n15311 ;
  assign n15313 = n1290 & ~n15171 ;
  assign n15314 = ( x215 & ~n14841 ) | ( x215 & n15313 ) | ( ~n14841 & n15313 ) ;
  assign n15315 = ( ~n14481 & n14843 ) | ( ~n14481 & n15314 ) | ( n14843 & n15314 ) ;
  assign n15316 = n4721 & n15296 ;
  assign n15317 = ( n4721 & ~n15285 ) | ( n4721 & n15316 ) | ( ~n15285 & n15316 ) ;
  assign n15318 = n2203 | n15315 ;
  assign n15319 = ( n15315 & ~n15317 ) | ( n15315 & n15318 ) | ( ~n15317 & n15318 ) ;
  assign n15320 = ~n15312 & n15319 ;
  assign n15321 = ~n15312 & n15315 ;
  assign n15322 = ( n15305 & n15320 ) | ( n15305 & n15321 ) | ( n15320 & n15321 ) ;
  assign n15323 = x299 & ~n15322 ;
  assign n15324 = n15304 & ~n15323 ;
  assign n15325 = x39 & n15324 ;
  assign n15326 = n15223 | n15325 ;
  assign n15327 = ~n15222 & n15326 ;
  assign n15328 = x665 & n14751 ;
  assign n15329 = x665 & n14750 ;
  assign n15330 = ( n14809 & n15328 ) | ( n14809 & n15329 ) | ( n15328 & n15329 ) ;
  assign n15331 = x198 & ~n15330 ;
  assign n15332 = x198 | x665 ;
  assign n15333 = ( x198 & n14781 ) | ( x198 & n15332 ) | ( n14781 & n15332 ) ;
  assign n15334 = x680 & ~n15333 ;
  assign n15335 = ( x680 & n15331 ) | ( x680 & n15334 ) | ( n15331 & n15334 ) ;
  assign n15336 = n14820 & ~n15335 ;
  assign n15337 = x299 | n15336 ;
  assign n15338 = x210 & ~n15330 ;
  assign n15339 = x210 | x665 ;
  assign n15340 = ( x210 & n14781 ) | ( x210 & n15339 ) | ( n14781 & n15339 ) ;
  assign n15341 = x680 & ~n15340 ;
  assign n15342 = ( x680 & n15338 ) | ( x680 & n15341 ) | ( n15338 & n15341 ) ;
  assign n15343 = n14814 & ~n15342 ;
  assign n15344 = x299 & ~n15343 ;
  assign n15345 = n15337 & ~n15344 ;
  assign n15346 = ( ~x39 & x140 ) | ( ~x39 & n15345 ) | ( x140 & n15345 ) ;
  assign n15347 = ~x198 & n15149 ;
  assign n15348 = ~x198 & x665 ;
  assign n15349 = ( ~n14780 & n15347 ) | ( ~n14780 & n15348 ) | ( n15347 & n15348 ) ;
  assign n15350 = ( x198 & n14783 ) | ( x198 & ~n15349 ) | ( n14783 & ~n15349 ) ;
  assign n15351 = x665 & ~n5995 ;
  assign n15352 = ( x665 & ~n14799 ) | ( x665 & n15351 ) | ( ~n14799 & n15351 ) ;
  assign n15353 = x198 & n15352 ;
  assign n15354 = x198 & ~n14909 ;
  assign n15355 = ( ~n14810 & n15353 ) | ( ~n14810 & n15354 ) | ( n15353 & n15354 ) ;
  assign n15356 = n15350 & ~n15355 ;
  assign n15357 = x299 | x680 ;
  assign n15358 = ( x299 & n15356 ) | ( x299 & n15357 ) | ( n15356 & n15357 ) ;
  assign n15359 = ~x210 & n15149 ;
  assign n15360 = ~x210 & x665 ;
  assign n15361 = ( ~n14780 & n15359 ) | ( ~n14780 & n15360 ) | ( n15359 & n15360 ) ;
  assign n15362 = ( x210 & n14783 ) | ( x210 & ~n15361 ) | ( n14783 & ~n15361 ) ;
  assign n15363 = x210 & n15352 ;
  assign n15364 = x210 & ~n14909 ;
  assign n15365 = ( ~n14810 & n15363 ) | ( ~n14810 & n15364 ) | ( n15363 & n15364 ) ;
  assign n15366 = n15362 & ~n15365 ;
  assign n15367 = x299 & ~x680 ;
  assign n15368 = ( x299 & ~n15366 ) | ( x299 & n15367 ) | ( ~n15366 & n15367 ) ;
  assign n15369 = n15358 & ~n15368 ;
  assign n15370 = ( x39 & x140 ) | ( x39 & n15369 ) | ( x140 & n15369 ) ;
  assign n15371 = n15346 & ~n15370 ;
  assign n15372 = n15327 | n15371 ;
  assign n15373 = ~x38 & n15372 ;
  assign n15374 = ~n4810 & n15202 ;
  assign n15375 = x38 & ~n15374 ;
  assign n15376 = n15071 & n15375 ;
  assign n15377 = x738 | n15376 ;
  assign n15378 = n15373 | n15377 ;
  assign n15379 = ~x140 & x738 ;
  assign n15380 = x38 & ~n14827 ;
  assign n15381 = x38 & n14827 ;
  assign n15382 = ( n14936 & ~n15380 ) | ( n14936 & n15381 ) | ( ~n15380 & n15381 ) ;
  assign n15383 = n15379 & ~n15382 ;
  assign n15384 = n2032 | n15383 ;
  assign n15385 = n15378 & ~n15384 ;
  assign n15386 = n14837 | n15385 ;
  assign n15387 = ~x778 & n15386 ;
  assign n15388 = ( x625 & x1153 ) | ( x625 & n14835 ) | ( x1153 & n14835 ) ;
  assign n15389 = ( ~x625 & x1153 ) | ( ~x625 & n15386 ) | ( x1153 & n15386 ) ;
  assign n15390 = n15388 & n15389 ;
  assign n15391 = ( x625 & x1153 ) | ( x625 & ~n14835 ) | ( x1153 & ~n14835 ) ;
  assign n15392 = ( x625 & ~x1153 ) | ( x625 & n15386 ) | ( ~x1153 & n15386 ) ;
  assign n15393 = ~n15391 & n15392 ;
  assign n15394 = n15390 | n15393 ;
  assign n15395 = x778 & n15394 ;
  assign n15396 = n15387 | n15395 ;
  assign n15397 = x660 | x1155 ;
  assign n15398 = x660 & x1155 ;
  assign n15399 = x785 & ~n15398 ;
  assign n15400 = n15397 & n15399 ;
  assign n15401 = n15396 & ~n15400 ;
  assign n15402 = n14835 & n15400 ;
  assign n15403 = n15401 | n15402 ;
  assign n15404 = x627 | x1154 ;
  assign n15405 = x627 & x1154 ;
  assign n15406 = x781 & ~n15405 ;
  assign n15407 = n15404 & n15406 ;
  assign n15408 = n15403 | n15407 ;
  assign n15409 = ~n14835 & n15407 ;
  assign n15410 = n15408 & ~n15409 ;
  assign n15411 = ~x648 & x1159 ;
  assign n15412 = x648 & ~x1159 ;
  assign n15413 = n15411 | n15412 ;
  assign n15414 = x789 & n15413 ;
  assign n15415 = n15410 & ~n15414 ;
  assign n15416 = n14835 & n15414 ;
  assign n15417 = n15415 | n15416 ;
  assign n15418 = ~x641 & x1158 ;
  assign n15419 = x641 & ~x1158 ;
  assign n15420 = n15418 | n15419 ;
  assign n15421 = x788 & n15420 ;
  assign n15422 = n15417 | n15421 ;
  assign n15423 = ~n14835 & n15421 ;
  assign n15424 = n15422 & ~n15423 ;
  assign n15425 = ~x792 & n15424 ;
  assign n15426 = ( x628 & x1156 ) | ( x628 & n14835 ) | ( x1156 & n14835 ) ;
  assign n15427 = ( ~x628 & x1156 ) | ( ~x628 & n15424 ) | ( x1156 & n15424 ) ;
  assign n15428 = n15426 & n15427 ;
  assign n15429 = ( x628 & x1156 ) | ( x628 & ~n14835 ) | ( x1156 & ~n14835 ) ;
  assign n15430 = ( x628 & ~x1156 ) | ( x628 & n15424 ) | ( ~x1156 & n15424 ) ;
  assign n15431 = ~n15429 & n15430 ;
  assign n15432 = n15428 | n15431 ;
  assign n15433 = x792 & n15432 ;
  assign n15434 = n15425 | n15433 ;
  assign n15435 = ~x787 & n15434 ;
  assign n15436 = ( x647 & x1157 ) | ( x647 & n14835 ) | ( x1157 & n14835 ) ;
  assign n15437 = ( ~x647 & x1157 ) | ( ~x647 & n15434 ) | ( x1157 & n15434 ) ;
  assign n15438 = n15436 & n15437 ;
  assign n15439 = ( x647 & x1157 ) | ( x647 & ~n14835 ) | ( x1157 & ~n14835 ) ;
  assign n15440 = ( x647 & ~x1157 ) | ( x647 & n15434 ) | ( ~x1157 & n15434 ) ;
  assign n15441 = ~n15439 & n15440 ;
  assign n15442 = n15438 | n15441 ;
  assign n15443 = x787 & n15442 ;
  assign n15444 = n15435 | n15443 ;
  assign n15445 = ( x644 & x715 ) | ( x644 & ~n15444 ) | ( x715 & ~n15444 ) ;
  assign n15446 = x630 | n15438 ;
  assign n15447 = ( x647 & x1157 ) | ( x647 & ~n15137 ) | ( x1157 & ~n15137 ) ;
  assign n15448 = x629 | n15428 ;
  assign n15449 = ( x628 & x1156 ) | ( x628 & ~n15130 ) | ( x1156 & ~n15130 ) ;
  assign n15450 = x648 | n15115 ;
  assign n15451 = ( x619 & x1159 ) | ( x619 & ~n15410 ) | ( x1159 & ~n15410 ) ;
  assign n15452 = x627 | n15105 ;
  assign n15453 = ( x618 & x1154 ) | ( x618 & ~n15403 ) | ( x1154 & ~n15403 ) ;
  assign n15454 = x660 | n15092 ;
  assign n15455 = ( x609 & x1155 ) | ( x609 & ~n15396 ) | ( x1155 & ~n15396 ) ;
  assign n15456 = x608 | n15390 ;
  assign n15457 = ( x625 & x1153 ) | ( x625 & ~n15078 ) | ( x1153 & ~n15078 ) ;
  assign n15458 = ( x738 & n2032 ) | ( x738 & ~n15076 ) | ( n2032 & ~n15076 ) ;
  assign n15459 = x603 & x665 ;
  assign n15460 = x603 & ~n15459 ;
  assign n15461 = ( n15150 & ~n15459 ) | ( n15150 & n15460 ) | ( ~n15459 & n15460 ) ;
  assign n15462 = n14959 & n15461 ;
  assign n15463 = x603 & ~x665 ;
  assign n15464 = n14959 & n15463 ;
  assign n15465 = ( ~n14481 & n15462 ) | ( ~n14481 & n15464 ) | ( n15462 & n15464 ) ;
  assign n15466 = n14517 & n15465 ;
  assign n15467 = ( n14510 & n15465 ) | ( n14510 & n15466 ) | ( n15465 & n15466 ) ;
  assign n15468 = ( ~n14481 & n15461 ) | ( ~n14481 & n15463 ) | ( n15461 & n15463 ) ;
  assign n15469 = x642 | n15468 ;
  assign n15470 = ( x642 & ~n14977 ) | ( x642 & n15469 ) | ( ~n14977 & n15469 ) ;
  assign n15471 = n15467 & n15470 ;
  assign n15472 = n4707 | n15471 ;
  assign n15473 = n14495 & ~n15467 ;
  assign n15474 = n14553 & ~n15473 ;
  assign n15475 = n15472 & n15474 ;
  assign n15476 = x616 & ~n15467 ;
  assign n15477 = ~n14839 & n15171 ;
  assign n15478 = n15160 | n15477 ;
  assign n15479 = ( n14465 & n15160 ) | ( n14465 & n15478 ) | ( n15160 & n15478 ) ;
  assign n15480 = n15160 | n15478 ;
  assign n15481 = ( n14474 & n15479 ) | ( n14474 & n15480 ) | ( n15479 & n15480 ) ;
  assign n15482 = ( n14553 & n15476 ) | ( n14553 & ~n15481 ) | ( n15476 & ~n15481 ) ;
  assign n15483 = n4764 & n15482 ;
  assign n15484 = ~n14553 & n15481 ;
  assign n15485 = n4764 & ~n15484 ;
  assign n15486 = ( ~n15475 & n15483 ) | ( ~n15475 & n15485 ) | ( n15483 & n15485 ) ;
  assign n15487 = ~n14977 & n15468 ;
  assign n15488 = n14980 & n15487 ;
  assign n15489 = ~x616 & n15149 ;
  assign n15490 = ~n14839 & n15150 ;
  assign n15491 = x616 & n15490 ;
  assign n15492 = ( ~x616 & n15160 ) | ( ~x616 & n15491 ) | ( n15160 & n15491 ) ;
  assign n15493 = ~x616 & n15160 ;
  assign n15494 = ( ~n14481 & n15492 ) | ( ~n14481 & n15493 ) | ( n15492 & n15493 ) ;
  assign n15495 = ~n15489 & n15494 ;
  assign n15496 = x616 & n15494 ;
  assign n15497 = ( n14988 & n15495 ) | ( n14988 & n15496 ) | ( n15495 & n15496 ) ;
  assign n15498 = n15488 | n15497 ;
  assign n15499 = x299 | n15276 ;
  assign n15500 = ( n2213 & n15498 ) | ( n2213 & n15499 ) | ( n15498 & n15499 ) ;
  assign n15501 = ( x299 & ~n15486 ) | ( x299 & n15500 ) | ( ~n15486 & n15500 ) ;
  assign n15502 = n15010 & n15157 ;
  assign n15503 = n14517 | n14609 ;
  assign n15504 = n15157 & n15503 ;
  assign n15505 = ~x665 & n15004 ;
  assign n15506 = x603 & ~n15505 ;
  assign n15507 = ~x665 & n15001 ;
  assign n15508 = x603 & ~n15507 ;
  assign n15509 = ( ~n14595 & n15506 ) | ( ~n14595 & n15508 ) | ( n15506 & n15508 ) ;
  assign n15510 = x603 & ~n15509 ;
  assign n15511 = n14855 | n15510 ;
  assign n15512 = ~n14855 & n15509 ;
  assign n15513 = ( n15504 & n15511 ) | ( n15504 & ~n15512 ) | ( n15511 & ~n15512 ) ;
  assign n15514 = n15502 & n15513 ;
  assign n15515 = ~n14854 & n15510 ;
  assign n15516 = x616 | n15515 ;
  assign n15517 = n14854 | n15509 ;
  assign n15518 = ~x616 & n15517 ;
  assign n15519 = ( n15504 & n15516 ) | ( n15504 & ~n15518 ) | ( n15516 & ~n15518 ) ;
  assign n15520 = n15514 | n15519 ;
  assign n15521 = ~n15160 & n15509 ;
  assign n15522 = ( n15160 & n15179 ) | ( n15160 & ~n15521 ) | ( n15179 & ~n15521 ) ;
  assign n15523 = x616 & ~n15157 ;
  assign n15524 = ( x616 & ~n15010 ) | ( x616 & n15523 ) | ( ~n15010 & n15523 ) ;
  assign n15525 = n14553 & ~n15524 ;
  assign n15526 = ( ~n14553 & n15522 ) | ( ~n14553 & n15525 ) | ( n15522 & n15525 ) ;
  assign n15527 = ~n14553 & n15522 ;
  assign n15528 = ( n15520 & n15526 ) | ( n15520 & n15527 ) | ( n15526 & n15527 ) ;
  assign n15529 = ~n14839 & n15202 ;
  assign n15530 = n1290 & n14840 ;
  assign n15531 = ( n1290 & n15529 ) | ( n1290 & n15530 ) | ( n15529 & n15530 ) ;
  assign n15532 = n1823 | n15531 ;
  assign n15533 = ( n1823 & ~n14481 ) | ( n1823 & n15532 ) | ( ~n14481 & n15532 ) ;
  assign n15534 = ~n14893 & n15533 ;
  assign n15535 = n14838 & n15463 ;
  assign n15536 = n14644 | n15535 ;
  assign n15537 = n14645 | n15535 ;
  assign n15538 = ( n14481 & n15536 ) | ( n14481 & n15537 ) | ( n15536 & n15537 ) ;
  assign n15539 = ( x603 & n14624 ) | ( x603 & n15538 ) | ( n14624 & n15538 ) ;
  assign n15540 = x603 | n15228 ;
  assign n15541 = x603 | n4713 ;
  assign n15542 = ( ~n14481 & n15540 ) | ( ~n14481 & n15541 ) | ( n15540 & n15541 ) ;
  assign n15543 = n4711 & ~n15542 ;
  assign n15544 = ~x603 & n4711 ;
  assign n15545 = ( n15244 & n15543 ) | ( n15244 & n15544 ) | ( n15543 & n15544 ) ;
  assign n15546 = ( n4711 & n15539 ) | ( n4711 & n15545 ) | ( n15539 & n15545 ) ;
  assign n15547 = ~n14974 & n15468 ;
  assign n15548 = ~x603 & n15468 ;
  assign n15549 = ( ~n15026 & n15547 ) | ( ~n15026 & n15548 ) | ( n15547 & n15548 ) ;
  assign n15550 = ( x616 & n14855 ) | ( x616 & n15490 ) | ( n14855 & n15490 ) ;
  assign n15551 = n14854 & ~n15550 ;
  assign n15552 = ~x616 & n14854 ;
  assign n15553 = ( n14481 & n15551 ) | ( n14481 & n15552 ) | ( n15551 & n15552 ) ;
  assign n15554 = n15494 & ~n15553 ;
  assign n15555 = ( x616 & ~n14481 ) | ( x616 & n15550 ) | ( ~n14481 & n15550 ) ;
  assign n15556 = n15494 & n15555 ;
  assign n15557 = ( n15549 & n15554 ) | ( n15549 & n15556 ) | ( n15554 & n15556 ) ;
  assign n15558 = n14641 | n15557 ;
  assign n15559 = ( n15546 & n15557 ) | ( n15546 & n15558 ) | ( n15557 & n15558 ) ;
  assign n15560 = ( n1823 & n14897 ) | ( n1823 & ~n15559 ) | ( n14897 & ~n15559 ) ;
  assign n15561 = n4764 & n15560 ;
  assign n15562 = ( n15534 & ~n15560 ) | ( n15534 & n15561 ) | ( ~n15560 & n15561 ) ;
  assign n15563 = n15534 & ~n15560 ;
  assign n15564 = ( n15528 & n15562 ) | ( n15528 & n15563 ) | ( n15562 & n15563 ) ;
  assign n15565 = n15501 | n15564 ;
  assign n15566 = ( x215 & n14686 ) | ( x215 & n15477 ) | ( n14686 & n15477 ) ;
  assign n15567 = ( x215 & ~n14481 ) | ( x215 & n15566 ) | ( ~n14481 & n15566 ) ;
  assign n15568 = n2203 | n15567 ;
  assign n15569 = ( ~n4721 & n15567 ) | ( ~n4721 & n15568 ) | ( n15567 & n15568 ) ;
  assign n15570 = n14853 | n15567 ;
  assign n15571 = ( ~n4721 & n15567 ) | ( ~n4721 & n15570 ) | ( n15567 & n15570 ) ;
  assign n15572 = ( n15559 & n15569 ) | ( n15559 & n15571 ) | ( n15569 & n15571 ) ;
  assign n15573 = n4721 & ~n15482 ;
  assign n15574 = n4721 & n15484 ;
  assign n15575 = ( n15475 & n15573 ) | ( n15475 & n15574 ) | ( n15573 & n15574 ) ;
  assign n15576 = ( x215 & n15308 ) | ( x215 & ~n15498 ) | ( n15308 & ~n15498 ) ;
  assign n15577 = x299 & n15576 ;
  assign n15578 = ~n15575 & n15577 ;
  assign n15579 = ( x299 & ~n15572 ) | ( x299 & n15578 ) | ( ~n15572 & n15578 ) ;
  assign n15580 = ( n15559 & n15568 ) | ( n15559 & n15570 ) | ( n15568 & n15570 ) ;
  assign n15581 = ( x299 & n15578 ) | ( x299 & ~n15580 ) | ( n15578 & ~n15580 ) ;
  assign n15582 = ( ~n15528 & n15579 ) | ( ~n15528 & n15581 ) | ( n15579 & n15581 ) ;
  assign n15583 = n15565 & ~n15582 ;
  assign n15584 = ( x140 & ~x761 ) | ( x140 & n15583 ) | ( ~x761 & n15583 ) ;
  assign n15585 = n14839 | n15149 ;
  assign n15586 = ~n14613 & n15585 ;
  assign n15587 = n14611 & n15586 ;
  assign n15588 = n15160 & ~n15587 ;
  assign n15589 = x603 & ~x621 ;
  assign n15590 = n15234 & ~n15589 ;
  assign n15591 = n4711 & ~n15590 ;
  assign n15592 = n15238 & ~n15589 ;
  assign n15593 = n4711 & ~n15592 ;
  assign n15594 = ( ~n14595 & n15591 ) | ( ~n14595 & n15593 ) | ( n15591 & n15593 ) ;
  assign n15595 = ~x603 & n15594 ;
  assign n15596 = ( ~n15019 & n15594 ) | ( ~n15019 & n15595 ) | ( n15594 & n15595 ) ;
  assign n15597 = n15285 & ~n15596 ;
  assign n15598 = ~n15588 & n15597 ;
  assign n15599 = ( n1823 & n15052 ) | ( n1823 & ~n15598 ) | ( n15052 & ~n15598 ) ;
  assign n15600 = x680 | n14678 ;
  assign n15601 = n14647 & n15585 ;
  assign n15602 = n14650 & n15585 ;
  assign n15603 = ( ~n14624 & n15601 ) | ( ~n14624 & n15602 ) | ( n15601 & n15602 ) ;
  assign n15604 = ( n1290 & n14839 ) | ( n1290 & n15224 ) | ( n14839 & n15224 ) ;
  assign n15605 = x614 & ~n15604 ;
  assign n15606 = ( x614 & n14481 ) | ( x614 & n15605 ) | ( n14481 & n15605 ) ;
  assign n15607 = x642 & ~n15604 ;
  assign n15608 = x642 & ~n15607 ;
  assign n15609 = x614 | n15608 ;
  assign n15610 = ( x614 & ~n14481 ) | ( x614 & n15609 ) | ( ~n14481 & n15609 ) ;
  assign n15611 = ~n15606 & n15610 ;
  assign n15612 = x616 | n15611 ;
  assign n15613 = x616 & ~n15604 ;
  assign n15614 = n15160 & n15613 ;
  assign n15615 = x616 & n15160 ;
  assign n15616 = ( n14481 & n15614 ) | ( n14481 & n15615 ) | ( n15614 & n15615 ) ;
  assign n15617 = ( n15160 & ~n15612 ) | ( n15160 & n15616 ) | ( ~n15612 & n15616 ) ;
  assign n15618 = ~x614 & n15607 ;
  assign n15619 = ~x614 & x642 ;
  assign n15620 = ( n14481 & n15618 ) | ( n14481 & n15619 ) | ( n15618 & n15619 ) ;
  assign n15621 = n15606 | n15620 ;
  assign n15622 = ~x616 & n15621 ;
  assign n15623 = ( n15160 & n15616 ) | ( n15160 & n15622 ) | ( n15616 & n15622 ) ;
  assign n15624 = ( ~n15603 & n15617 ) | ( ~n15603 & n15623 ) | ( n15617 & n15623 ) ;
  assign n15625 = n15546 | n15624 ;
  assign n15626 = n15600 & ~n15625 ;
  assign n15627 = ~n4764 & n15626 ;
  assign n15628 = n15599 & ~n15627 ;
  assign n15629 = ~x223 & n1823 ;
  assign n15630 = n1290 & ~n15477 ;
  assign n15631 = ~n1823 & n15630 ;
  assign n15632 = ( ~x223 & n1823 ) | ( ~x223 & n15631 ) | ( n1823 & n15631 ) ;
  assign n15633 = ( ~n14481 & n15629 ) | ( ~n14481 & n15632 ) | ( n15629 & n15632 ) ;
  assign n15634 = ~n15628 & n15633 ;
  assign n15635 = n14475 & n14874 ;
  assign n15636 = x665 & n14465 ;
  assign n15637 = ~x603 & n15257 ;
  assign n15638 = ~n14481 & n15637 ;
  assign n15639 = n15636 | n15638 ;
  assign n15640 = n14855 | n15639 ;
  assign n15641 = n15635 | n15640 ;
  assign n15642 = ~n14481 & n15257 ;
  assign n15643 = n15636 | n15642 ;
  assign n15644 = n14855 & ~n15643 ;
  assign n15645 = ~n14876 & n15644 ;
  assign n15646 = n15641 & ~n15645 ;
  assign n15647 = ~x665 & n4711 ;
  assign n15648 = ( n4711 & ~n14465 ) | ( n4711 & n15647 ) | ( ~n14465 & n15647 ) ;
  assign n15649 = ~n14874 & n15648 ;
  assign n15650 = ( ~n14475 & n15648 ) | ( ~n14475 & n15649 ) | ( n15648 & n15649 ) ;
  assign n15651 = n15160 | n15650 ;
  assign n15652 = ( ~n15646 & n15650 ) | ( ~n15646 & n15651 ) | ( n15650 & n15651 ) ;
  assign n15653 = x680 | n14519 ;
  assign n15654 = x680 | n14521 ;
  assign n15655 = ( n14515 & n15653 ) | ( n14515 & n15654 ) | ( n15653 & n15654 ) ;
  assign n15656 = n4764 & ~n15655 ;
  assign n15657 = ( n4764 & n15652 ) | ( n4764 & n15656 ) | ( n15652 & n15656 ) ;
  assign n15658 = x223 & ~n15657 ;
  assign n15659 = ~n14884 & n15270 ;
  assign n15660 = n15275 & ~n15659 ;
  assign n15661 = n15635 | n15639 ;
  assign n15662 = x642 | n15228 ;
  assign n15663 = x642 | n4713 ;
  assign n15664 = ( ~n14481 & n15662 ) | ( ~n14481 & n15663 ) | ( n15662 & n15663 ) ;
  assign n15665 = ( x642 & ~n15269 ) | ( x642 & n15664 ) | ( ~n15269 & n15664 ) ;
  assign n15666 = n14884 | n15665 ;
  assign n15667 = n15661 | n15666 ;
  assign n15668 = ( x616 & n14481 ) | ( x616 & n15613 ) | ( n14481 & n15613 ) ;
  assign n15669 = n15622 | n15668 ;
  assign n15670 = n15160 & n15669 ;
  assign n15671 = x614 & ~n15605 ;
  assign n15672 = x616 | n15671 ;
  assign n15673 = ( x616 & ~n14481 ) | ( x616 & n15672 ) | ( ~n14481 & n15672 ) ;
  assign n15674 = ~n15668 & n15673 ;
  assign n15675 = n15160 & ~n15674 ;
  assign n15676 = ( ~n15667 & n15670 ) | ( ~n15667 & n15675 ) | ( n15670 & n15675 ) ;
  assign n15677 = n15660 & ~n15676 ;
  assign n15678 = n4764 | n15677 ;
  assign n15679 = n15658 & n15678 ;
  assign n15680 = ~x299 & n15679 ;
  assign n15681 = ( ~x299 & n15634 ) | ( ~x299 & n15680 ) | ( n15634 & n15680 ) ;
  assign n15682 = n4721 & ~n15598 ;
  assign n15683 = n4721 | n15626 ;
  assign n15684 = ~n15682 & n15683 ;
  assign n15685 = ~n2203 & n15630 ;
  assign n15686 = ( ~x215 & n2203 ) | ( ~x215 & n15685 ) | ( n2203 & n15685 ) ;
  assign n15687 = ( ~n14481 & n14841 ) | ( ~n14481 & n15686 ) | ( n14841 & n15686 ) ;
  assign n15688 = ~n2203 & n15686 ;
  assign n15689 = ~n2203 & n14841 ;
  assign n15690 = ( ~n14481 & n15688 ) | ( ~n14481 & n15689 ) | ( n15688 & n15689 ) ;
  assign n15691 = ( n15684 & n15687 ) | ( n15684 & n15690 ) | ( n15687 & n15690 ) ;
  assign n15692 = n4721 & ~n15655 ;
  assign n15693 = ( n4721 & n15652 ) | ( n4721 & n15692 ) | ( n15652 & n15692 ) ;
  assign n15694 = x215 & ~n15693 ;
  assign n15695 = n4721 | n15677 ;
  assign n15696 = n15694 & n15695 ;
  assign n15697 = x299 & n15696 ;
  assign n15698 = ( x299 & n15691 ) | ( x299 & n15697 ) | ( n15691 & n15697 ) ;
  assign n15699 = n15681 | n15698 ;
  assign n15700 = ( x140 & x761 ) | ( x140 & n15699 ) | ( x761 & n15699 ) ;
  assign n15701 = ~n15584 & n15700 ;
  assign n15702 = x680 | n14982 ;
  assign n15703 = ( x680 & ~n14481 ) | ( x680 & n15702 ) | ( ~n14481 & n15702 ) ;
  assign n15704 = n15034 | n15703 ;
  assign n15705 = n15149 & ~n15589 ;
  assign n15706 = n15228 & n15705 ;
  assign n15707 = n4711 & ~n15706 ;
  assign n15708 = n4713 & n15705 ;
  assign n15709 = n4711 & ~n15708 ;
  assign n15710 = ( n14481 & n15707 ) | ( n14481 & n15709 ) | ( n15707 & n15709 ) ;
  assign n15711 = ( n4711 & n15244 ) | ( n4711 & n15710 ) | ( n15244 & n15710 ) ;
  assign n15712 = n15704 & ~n15711 ;
  assign n15713 = n15224 & ~n15589 ;
  assign n15714 = ~n14855 & n15160 ;
  assign n15715 = ( n15160 & ~n15713 ) | ( n15160 & n15714 ) | ( ~n15713 & n15714 ) ;
  assign n15716 = n15160 | n15714 ;
  assign n15717 = ( n14481 & n15715 ) | ( n14481 & n15716 ) | ( n15715 & n15716 ) ;
  assign n15718 = ~n15149 & n15716 ;
  assign n15719 = ~n15149 & n15715 ;
  assign n15720 = ( n14481 & n15718 ) | ( n14481 & n15719 ) | ( n15718 & n15719 ) ;
  assign n15721 = ( ~n15034 & n15717 ) | ( ~n15034 & n15720 ) | ( n15717 & n15720 ) ;
  assign n15722 = n4764 | n15721 ;
  assign n15723 = n15712 & ~n15722 ;
  assign n15724 = n1823 & n15723 ;
  assign n15725 = n14613 | n14839 ;
  assign n15726 = n14611 & ~n15725 ;
  assign n15727 = ~n15292 & n15705 ;
  assign n15728 = ~n15291 & n15705 ;
  assign n15729 = ( ~n14595 & n15727 ) | ( ~n14595 & n15728 ) | ( n15727 & n15728 ) ;
  assign n15730 = ( ~n15160 & n15259 ) | ( ~n15160 & n15705 ) | ( n15259 & n15705 ) ;
  assign n15731 = n15160 & ~n15705 ;
  assign n15732 = ( n15729 & ~n15730 ) | ( n15729 & n15731 ) | ( ~n15730 & n15731 ) ;
  assign n15733 = x680 & ~n15594 ;
  assign n15734 = ~n15732 & n15733 ;
  assign n15735 = n4764 & n15734 ;
  assign n15736 = n15594 | n15732 ;
  assign n15737 = n4764 & ~n15736 ;
  assign n15738 = ( n15726 & n15735 ) | ( n15726 & n15737 ) | ( n15735 & n15737 ) ;
  assign n15739 = ( n1823 & n15724 ) | ( n1823 & n15738 ) | ( n15724 & n15738 ) ;
  assign n15740 = n15255 | n15589 ;
  assign n15741 = n4711 & n15740 ;
  assign n15742 = x680 | n15589 ;
  assign n15743 = n4711 & n15742 ;
  assign n15744 = ( ~n14465 & n15741 ) | ( ~n14465 & n15743 ) | ( n15741 & n15743 ) ;
  assign n15745 = x680 & ~n15743 ;
  assign n15746 = x680 & ~n15741 ;
  assign n15747 = ( n14465 & n15745 ) | ( n14465 & n15746 ) | ( n15745 & n15746 ) ;
  assign n15748 = ( n14961 & ~n15744 ) | ( n14961 & n15747 ) | ( ~n15744 & n15747 ) ;
  assign n15749 = ~n15744 & n15747 ;
  assign n15750 = ( n14962 & n15748 ) | ( n14962 & n15749 ) | ( n15748 & n15749 ) ;
  assign n15751 = n15160 & ~n15643 ;
  assign n15752 = ( ~n14988 & n15160 ) | ( ~n14988 & n15751 ) | ( n15160 & n15751 ) ;
  assign n15753 = n4764 & ~n15752 ;
  assign n15754 = n15750 & n15753 ;
  assign n15755 = ~n1271 & n14457 ;
  assign n15756 = ~n1242 & n15755 ;
  assign n15757 = ( n14839 & n15171 ) | ( n14839 & n15756 ) | ( n15171 & n15756 ) ;
  assign n15758 = n15756 & ~n15757 ;
  assign n15759 = ( ~x223 & n14479 ) | ( ~x223 & n15629 ) | ( n14479 & n15629 ) ;
  assign n15760 = x223 & ~n15629 ;
  assign n15761 = ( n15758 & ~n15759 ) | ( n15758 & n15760 ) | ( ~n15759 & n15760 ) ;
  assign n15762 = n4711 & ~n15589 ;
  assign n15763 = n15228 & n15762 ;
  assign n15764 = n4713 & n15762 ;
  assign n15765 = ( ~n14481 & n15763 ) | ( ~n14481 & n15764 ) | ( n15763 & n15764 ) ;
  assign n15766 = ~n15269 & n15765 ;
  assign n15767 = n15171 & ~n15766 ;
  assign n15768 = ( x223 & n15276 ) | ( x223 & n15767 ) | ( n15276 & n15767 ) ;
  assign n15769 = ( x223 & n15276 ) | ( x223 & ~n15766 ) | ( n15276 & ~n15766 ) ;
  assign n15770 = ( ~n14989 & n15768 ) | ( ~n14989 & n15769 ) | ( n15768 & n15769 ) ;
  assign n15771 = n15761 & ~n15770 ;
  assign n15772 = ( n15754 & n15761 ) | ( n15754 & n15771 ) | ( n15761 & n15771 ) ;
  assign n15773 = x299 | n15772 ;
  assign n15774 = ~n15754 & n15770 ;
  assign n15775 = ~x299 & n15774 ;
  assign n15776 = ( n15739 & n15773 ) | ( n15739 & ~n15775 ) | ( n15773 & ~n15775 ) ;
  assign n15777 = n4721 | n15721 ;
  assign n15778 = n15712 & ~n15777 ;
  assign n15779 = n2203 & n15778 ;
  assign n15780 = n4721 & n15734 ;
  assign n15781 = n4721 & ~n15736 ;
  assign n15782 = ( n15726 & n15780 ) | ( n15726 & n15781 ) | ( n15780 & n15781 ) ;
  assign n15783 = ( n2203 & n15779 ) | ( n2203 & n15782 ) | ( n15779 & n15782 ) ;
  assign n15784 = n4721 & ~n15752 ;
  assign n15785 = n15750 & n15784 ;
  assign n15786 = ( ~x215 & n14479 ) | ( ~x215 & n14841 ) | ( n14479 & n14841 ) ;
  assign n15787 = ( n14843 & n15758 ) | ( n14843 & ~n15786 ) | ( n15758 & ~n15786 ) ;
  assign n15788 = ( x215 & n15308 ) | ( x215 & n15767 ) | ( n15308 & n15767 ) ;
  assign n15789 = ( x215 & n15308 ) | ( x215 & ~n15766 ) | ( n15308 & ~n15766 ) ;
  assign n15790 = ( ~n14989 & n15788 ) | ( ~n14989 & n15789 ) | ( n15788 & n15789 ) ;
  assign n15791 = n15787 & ~n15790 ;
  assign n15792 = ( n15785 & n15787 ) | ( n15785 & n15791 ) | ( n15787 & n15791 ) ;
  assign n15793 = x299 & ~n15792 ;
  assign n15794 = ~n15785 & n15790 ;
  assign n15795 = x299 & n15794 ;
  assign n15796 = ( ~n15783 & n15793 ) | ( ~n15783 & n15795 ) | ( n15793 & n15795 ) ;
  assign n15797 = n15776 & ~n15796 ;
  assign n15798 = ( x140 & ~x761 ) | ( x140 & n15797 ) | ( ~x761 & n15797 ) ;
  assign n15799 = ~n14624 & n14867 ;
  assign n15800 = ~n14855 & n15549 ;
  assign n15801 = ( ~n14855 & n15799 ) | ( ~n14855 & n15800 ) | ( n15799 & n15800 ) ;
  assign n15802 = n1290 & ~n15705 ;
  assign n15803 = ( n15160 & n15714 ) | ( n15160 & ~n15802 ) | ( n15714 & ~n15802 ) ;
  assign n15804 = ( n14481 & n15716 ) | ( n14481 & n15803 ) | ( n15716 & n15803 ) ;
  assign n15805 = ~n15801 & n15804 ;
  assign n15806 = x680 | n14863 ;
  assign n15807 = x680 | n14857 ;
  assign n15808 = ( ~n14624 & n15806 ) | ( ~n14624 & n15807 ) | ( n15806 & n15807 ) ;
  assign n15809 = n4711 & ~n14867 ;
  assign n15810 = ( n4711 & n14624 ) | ( n4711 & n15809 ) | ( n14624 & n15809 ) ;
  assign n15811 = n15808 & ~n15810 ;
  assign n15812 = ( n15158 & n15808 ) | ( n15158 & n15811 ) | ( n15808 & n15811 ) ;
  assign n15813 = ~n15805 & n15812 ;
  assign n15814 = ( n1823 & n14897 ) | ( n1823 & ~n15813 ) | ( n14897 & ~n15813 ) ;
  assign n15815 = x603 & n15019 ;
  assign n15816 = ( x603 & ~n15509 ) | ( x603 & n15815 ) | ( ~n15509 & n15815 ) ;
  assign n15817 = n15509 & ~n15815 ;
  assign n15818 = ( n15504 & n15816 ) | ( n15504 & ~n15817 ) | ( n15816 & ~n15817 ) ;
  assign n15819 = ~n14855 & n15818 ;
  assign n15820 = n14517 & n14839 ;
  assign n15821 = ( n14609 & n14839 ) | ( n14609 & n15820 ) | ( n14839 & n15820 ) ;
  assign n15822 = n14855 & n15821 ;
  assign n15823 = ( n14855 & n15504 ) | ( n14855 & n15822 ) | ( n15504 & n15822 ) ;
  assign n15824 = n15160 & ~n15823 ;
  assign n15825 = ~n15819 & n15824 ;
  assign n15826 = n4711 | n15160 ;
  assign n15827 = ( n15156 & n15160 ) | ( n15156 & n15826 ) | ( n15160 & n15826 ) ;
  assign n15828 = n14849 | n15827 ;
  assign n15829 = ( n14846 & n15827 ) | ( n14846 & n15828 ) | ( n15827 & n15828 ) ;
  assign n15830 = n4764 & n15829 ;
  assign n15831 = ~n15825 & n15830 ;
  assign n15832 = n15814 & ~n15831 ;
  assign n15833 = ~n14855 & n14883 ;
  assign n15834 = ~n14855 & n14874 ;
  assign n15835 = ( n14475 & n15833 ) | ( n14475 & n15834 ) | ( n15833 & n15834 ) ;
  assign n15836 = ( ~n14855 & n15187 ) | ( ~n14855 & n15835 ) | ( n15187 & n15835 ) ;
  assign n15837 = n15804 & ~n15836 ;
  assign n15838 = ( x680 & n15160 ) | ( x680 & n15184 ) | ( n15160 & n15184 ) ;
  assign n15839 = ( x680 & n15151 ) | ( x680 & n15160 ) | ( n15151 & n15160 ) ;
  assign n15840 = ( n14475 & n15838 ) | ( n14475 & n15839 ) | ( n15838 & n15839 ) ;
  assign n15841 = n14884 | n15840 ;
  assign n15842 = n14881 | n15841 ;
  assign n15843 = ~n15837 & n15842 ;
  assign n15844 = n4764 | n15843 ;
  assign n15845 = n14881 | n15635 ;
  assign n15846 = n15187 & n15840 ;
  assign n15847 = n14517 & n15151 ;
  assign n15848 = ( n14510 & n15151 ) | ( n14510 & n15847 ) | ( n15151 & n15847 ) ;
  assign n15849 = n15846 & n15848 ;
  assign n15850 = n15845 | n15849 ;
  assign n15851 = ( x223 & n15044 ) | ( x223 & n15850 ) | ( n15044 & n15850 ) ;
  assign n15852 = n15844 & n15851 ;
  assign n15853 = x299 | n15852 ;
  assign n15854 = ( ~x223 & n15531 ) | ( ~x223 & n15629 ) | ( n15531 & n15629 ) ;
  assign n15855 = ( ~n14481 & n15629 ) | ( ~n14481 & n15854 ) | ( n15629 & n15854 ) ;
  assign n15856 = x299 | n15855 ;
  assign n15857 = n15852 | n15856 ;
  assign n15858 = ( ~n15832 & n15853 ) | ( ~n15832 & n15857 ) | ( n15853 & n15857 ) ;
  assign n15859 = n15023 & n15813 ;
  assign n15860 = n4721 & n15829 ;
  assign n15861 = ~n15825 & n15860 ;
  assign n15862 = ( n2203 & n15859 ) | ( n2203 & n15861 ) | ( n15859 & n15861 ) ;
  assign n15863 = ~n4721 & n15843 ;
  assign n15864 = ( x215 & n14958 ) | ( x215 & ~n15850 ) | ( n14958 & ~n15850 ) ;
  assign n15865 = ~n15863 & n15864 ;
  assign n15866 = ( x215 & ~n14841 ) | ( x215 & n15531 ) | ( ~n14841 & n15531 ) ;
  assign n15867 = ( ~n14481 & n14843 ) | ( ~n14481 & n15866 ) | ( n14843 & n15866 ) ;
  assign n15868 = n15865 | n15867 ;
  assign n15869 = ( x299 & n15865 ) | ( x299 & ~n15868 ) | ( n15865 & ~n15868 ) ;
  assign n15870 = x299 & n15865 ;
  assign n15871 = ( ~n15862 & n15869 ) | ( ~n15862 & n15870 ) | ( n15869 & n15870 ) ;
  assign n15872 = n15858 & ~n15871 ;
  assign n15873 = ( x140 & x761 ) | ( x140 & n15872 ) | ( x761 & n15872 ) ;
  assign n15874 = n15798 & ~n15873 ;
  assign n15875 = n15701 | n15874 ;
  assign n15876 = x39 & n15875 ;
  assign n15877 = x603 & ~n14952 ;
  assign n15878 = ( x603 & n14951 ) | ( x603 & n15877 ) | ( n14951 & n15877 ) ;
  assign n15879 = n15459 | n15878 ;
  assign n15880 = x603 | n15356 ;
  assign n15881 = ~n15879 & n15880 ;
  assign n15882 = ( x299 & x680 ) | ( x299 & n15881 ) | ( x680 & n15881 ) ;
  assign n15883 = n14945 | n15459 ;
  assign n15884 = x603 | n15366 ;
  assign n15885 = ~n15883 & n15884 ;
  assign n15886 = ( ~x299 & x680 ) | ( ~x299 & n15885 ) | ( x680 & n15885 ) ;
  assign n15887 = n15882 & n15886 ;
  assign n15888 = ( ~x140 & x761 ) | ( ~x140 & n15887 ) | ( x761 & n15887 ) ;
  assign n15889 = x680 & n14930 ;
  assign n15890 = ~n14921 & n15889 ;
  assign n15891 = n15345 | n15890 ;
  assign n15892 = ( x140 & x761 ) | ( x140 & ~n15891 ) | ( x761 & ~n15891 ) ;
  assign n15893 = n15888 & n15892 ;
  assign n15894 = n14956 & n15345 ;
  assign n15895 = ( ~x140 & x761 ) | ( ~x140 & n15894 ) | ( x761 & n15894 ) ;
  assign n15896 = ~n14921 & n14930 ;
  assign n15897 = n15369 | n15896 ;
  assign n15898 = ( x140 & x761 ) | ( x140 & ~n15897 ) | ( x761 & ~n15897 ) ;
  assign n15899 = n15895 | n15898 ;
  assign n15900 = ~n15893 & n15899 ;
  assign n15901 = ( x38 & ~n9138 ) | ( x38 & n15900 ) | ( ~n9138 & n15900 ) ;
  assign n15902 = n15876 | n15901 ;
  assign n15903 = x140 | n15758 ;
  assign n15904 = n14840 | n15529 ;
  assign n15905 = x140 & n15904 ;
  assign n15906 = ~n1868 & n15905 ;
  assign n15907 = x761 | n15906 ;
  assign n15908 = n15903 & ~n15907 ;
  assign n15909 = x140 | n15756 ;
  assign n15910 = x761 & n15909 ;
  assign n15911 = n14457 & n15477 ;
  assign n15912 = ~n1271 & n15911 ;
  assign n15913 = ~n1242 & n15912 ;
  assign n15914 = n15910 & ~n15913 ;
  assign n15915 = n15908 | n15914 ;
  assign n15916 = ~x39 & n15915 ;
  assign n15917 = x38 & ~n15223 ;
  assign n15918 = ~n15916 & n15917 ;
  assign n15919 = n15902 & ~n15918 ;
  assign n15920 = ( x738 & ~n2032 ) | ( x738 & n15919 ) | ( ~n2032 & n15919 ) ;
  assign n15921 = ~n15458 & n15920 ;
  assign n15922 = n14837 | n15921 ;
  assign n15923 = ( x625 & ~x1153 ) | ( x625 & n15922 ) | ( ~x1153 & n15922 ) ;
  assign n15924 = ~n15457 & n15923 ;
  assign n15925 = n15456 | n15924 ;
  assign n15926 = x608 & ~n15393 ;
  assign n15927 = ( x625 & x1153 ) | ( x625 & n15078 ) | ( x1153 & n15078 ) ;
  assign n15928 = ( ~x625 & x1153 ) | ( ~x625 & n15922 ) | ( x1153 & n15922 ) ;
  assign n15929 = n15927 & n15928 ;
  assign n15930 = n15926 & ~n15929 ;
  assign n15931 = n15925 & ~n15930 ;
  assign n15932 = x778 & ~n15931 ;
  assign n15933 = x778 | n15922 ;
  assign n15934 = ~n15932 & n15933 ;
  assign n15935 = ( x609 & ~x1155 ) | ( x609 & n15934 ) | ( ~x1155 & n15934 ) ;
  assign n15936 = ~n15455 & n15935 ;
  assign n15937 = n15454 | n15936 ;
  assign n15938 = x660 & ~n15098 ;
  assign n15939 = ( x609 & x1155 ) | ( x609 & n15396 ) | ( x1155 & n15396 ) ;
  assign n15940 = ( ~x609 & x1155 ) | ( ~x609 & n15934 ) | ( x1155 & n15934 ) ;
  assign n15941 = n15939 & n15940 ;
  assign n15942 = n15938 & ~n15941 ;
  assign n15943 = n15937 & ~n15942 ;
  assign n15944 = x785 & ~n15943 ;
  assign n15945 = x785 | n15934 ;
  assign n15946 = ~n15944 & n15945 ;
  assign n15947 = ( x618 & ~x1154 ) | ( x618 & n15946 ) | ( ~x1154 & n15946 ) ;
  assign n15948 = ~n15453 & n15947 ;
  assign n15949 = n15452 | n15948 ;
  assign n15950 = x627 & ~n15108 ;
  assign n15951 = ( x618 & x1154 ) | ( x618 & n15403 ) | ( x1154 & n15403 ) ;
  assign n15952 = ( ~x618 & x1154 ) | ( ~x618 & n15946 ) | ( x1154 & n15946 ) ;
  assign n15953 = n15951 & n15952 ;
  assign n15954 = n15950 & ~n15953 ;
  assign n15955 = n15949 & ~n15954 ;
  assign n15956 = x781 & ~n15955 ;
  assign n15957 = x781 | n15946 ;
  assign n15958 = ~n15956 & n15957 ;
  assign n15959 = ( x619 & ~x1159 ) | ( x619 & n15958 ) | ( ~x1159 & n15958 ) ;
  assign n15960 = ~n15451 & n15959 ;
  assign n15961 = n15450 | n15960 ;
  assign n15962 = x648 & ~n15118 ;
  assign n15963 = ( x619 & x1159 ) | ( x619 & n15410 ) | ( x1159 & n15410 ) ;
  assign n15964 = ( ~x619 & x1159 ) | ( ~x619 & n15958 ) | ( x1159 & n15958 ) ;
  assign n15965 = n15963 & n15964 ;
  assign n15966 = n15962 & ~n15965 ;
  assign n15967 = n15961 & ~n15966 ;
  assign n15968 = x789 & ~n15967 ;
  assign n15969 = x789 | n15958 ;
  assign n15970 = ~n15968 & n15969 ;
  assign n15971 = ~x788 & n15970 ;
  assign n15972 = x641 | x1158 ;
  assign n15973 = ~n15123 & n15972 ;
  assign n15974 = ( x626 & x641 ) | ( x626 & n15417 ) | ( x641 & n15417 ) ;
  assign n15975 = ( ~x626 & x641 ) | ( ~x626 & n15970 ) | ( x641 & n15970 ) ;
  assign n15976 = n15974 | n15975 ;
  assign n15977 = ~n15973 & n15976 ;
  assign n15978 = x641 & x1158 ;
  assign n15979 = n15126 | n15978 ;
  assign n15980 = ( x626 & x641 ) | ( x626 & ~n15417 ) | ( x641 & ~n15417 ) ;
  assign n15981 = ( x626 & ~x641 ) | ( x626 & n15970 ) | ( ~x641 & n15970 ) ;
  assign n15982 = n15980 & ~n15981 ;
  assign n15983 = n15979 & ~n15982 ;
  assign n15984 = n15977 | n15983 ;
  assign n15985 = x788 & n15984 ;
  assign n15986 = n15971 | n15985 ;
  assign n15987 = ( x628 & ~x1156 ) | ( x628 & n15986 ) | ( ~x1156 & n15986 ) ;
  assign n15988 = ~n15449 & n15987 ;
  assign n15989 = n15448 | n15988 ;
  assign n15990 = x629 & ~n15431 ;
  assign n15991 = ( x628 & x1156 ) | ( x628 & n15130 ) | ( x1156 & n15130 ) ;
  assign n15992 = ( ~x628 & x1156 ) | ( ~x628 & n15986 ) | ( x1156 & n15986 ) ;
  assign n15993 = n15991 & n15992 ;
  assign n15994 = n15990 & ~n15993 ;
  assign n15995 = n15989 & ~n15994 ;
  assign n15996 = x792 & ~n15995 ;
  assign n15997 = x792 | n15986 ;
  assign n15998 = ~n15996 & n15997 ;
  assign n15999 = ( x647 & ~x1157 ) | ( x647 & n15998 ) | ( ~x1157 & n15998 ) ;
  assign n16000 = ~n15447 & n15999 ;
  assign n16001 = n15446 | n16000 ;
  assign n16002 = x630 & ~n15441 ;
  assign n16003 = ( x647 & x1157 ) | ( x647 & n15137 ) | ( x1157 & n15137 ) ;
  assign n16004 = ( ~x647 & x1157 ) | ( ~x647 & n15998 ) | ( x1157 & n15998 ) ;
  assign n16005 = n16003 & n16004 ;
  assign n16006 = n16002 & ~n16005 ;
  assign n16007 = n16001 & ~n16006 ;
  assign n16008 = x787 & ~n16007 ;
  assign n16009 = x787 | n15998 ;
  assign n16010 = ~n16008 & n16009 ;
  assign n16011 = ( x644 & ~x715 ) | ( x644 & n16010 ) | ( ~x715 & n16010 ) ;
  assign n16012 = ~n15445 & n16011 ;
  assign n16013 = n15148 | n16012 ;
  assign n16014 = ( x644 & x715 ) | ( x644 & ~n15144 ) | ( x715 & ~n15144 ) ;
  assign n16015 = ( x644 & ~x715 ) | ( x644 & n14835 ) | ( ~x715 & n14835 ) ;
  assign n16016 = ~n16014 & n16015 ;
  assign n16017 = x1160 & ~n16016 ;
  assign n16018 = ( x644 & x715 ) | ( x644 & n15444 ) | ( x715 & n15444 ) ;
  assign n16019 = ( ~x644 & x715 ) | ( ~x644 & n16010 ) | ( x715 & n16010 ) ;
  assign n16020 = n16018 & n16019 ;
  assign n16021 = n16017 & ~n16020 ;
  assign n16022 = x790 & ~n16021 ;
  assign n16023 = n16013 & n16022 ;
  assign n16024 = ~x790 & n16010 ;
  assign n16025 = n6785 | n16024 ;
  assign n16026 = n16023 | n16025 ;
  assign n16027 = ~x140 & n6785 ;
  assign n16028 = x832 | n16027 ;
  assign n16029 = n16026 & ~n16028 ;
  assign n16030 = x140 | n1290 ;
  assign n16031 = ( x647 & x1157 ) | ( x647 & n16030 ) | ( x1157 & n16030 ) ;
  assign n16032 = ~x738 & n15202 ;
  assign n16033 = n16030 & ~n16032 ;
  assign n16034 = ~x778 & n16033 ;
  assign n16035 = ~x625 & n16032 ;
  assign n16036 = n16033 | n16035 ;
  assign n16037 = x1153 & n16036 ;
  assign n16038 = ~x1153 & n16030 ;
  assign n16039 = ~n16035 & n16038 ;
  assign n16040 = n16037 | n16039 ;
  assign n16041 = x778 & n16040 ;
  assign n16042 = n16034 | n16041 ;
  assign n16043 = n1290 & n15400 ;
  assign n16044 = n16042 | n16043 ;
  assign n16045 = n1290 & n15407 ;
  assign n16046 = n16044 | n16045 ;
  assign n16047 = n1290 & n15414 ;
  assign n16048 = n16046 | n16047 ;
  assign n16049 = n1290 & n15421 ;
  assign n16050 = n16048 | n16049 ;
  assign n16051 = ~x628 & x1156 ;
  assign n16052 = x628 & ~x1156 ;
  assign n16053 = n16051 | n16052 ;
  assign n16054 = x792 & n16053 ;
  assign n16055 = n1290 & n16054 ;
  assign n16056 = n16050 | n16055 ;
  assign n16057 = ( ~x647 & x1157 ) | ( ~x647 & n16056 ) | ( x1157 & n16056 ) ;
  assign n16058 = n16031 & n16057 ;
  assign n16059 = x630 | n16058 ;
  assign n16060 = n1290 & n15082 ;
  assign n16061 = ~x761 & n14840 ;
  assign n16062 = n16030 & ~n16061 ;
  assign n16063 = n16060 | n16062 ;
  assign n16064 = ~x785 & n16063 ;
  assign n16065 = n1290 & ~n15088 ;
  assign n16066 = n16062 | n16065 ;
  assign n16067 = x1155 & n16066 ;
  assign n16068 = x609 & n1290 ;
  assign n16069 = n16063 | n16068 ;
  assign n16070 = ~x1155 & n16069 ;
  assign n16071 = n16067 | n16070 ;
  assign n16072 = x785 & n16071 ;
  assign n16073 = n16064 | n16072 ;
  assign n16074 = ~x781 & n16073 ;
  assign n16075 = ~x618 & n1290 ;
  assign n16076 = n16073 | n16075 ;
  assign n16077 = x1154 & n16076 ;
  assign n16078 = x618 & n1290 ;
  assign n16079 = n16073 | n16078 ;
  assign n16080 = ~x1154 & n16079 ;
  assign n16081 = n16077 | n16080 ;
  assign n16082 = x781 & n16081 ;
  assign n16083 = n16074 | n16082 ;
  assign n16084 = ~x789 & n16083 ;
  assign n16085 = ( x619 & x1159 ) | ( x619 & n16030 ) | ( x1159 & n16030 ) ;
  assign n16086 = ( ~x619 & x1159 ) | ( ~x619 & n16083 ) | ( x1159 & n16083 ) ;
  assign n16087 = n16085 & n16086 ;
  assign n16088 = ( x619 & x1159 ) | ( x619 & ~n16030 ) | ( x1159 & ~n16030 ) ;
  assign n16089 = ( x619 & ~x1159 ) | ( x619 & n16083 ) | ( ~x1159 & n16083 ) ;
  assign n16090 = ~n16088 & n16089 ;
  assign n16091 = n16087 | n16090 ;
  assign n16092 = x789 & n16091 ;
  assign n16093 = n16084 | n16092 ;
  assign n16094 = ~x788 & n16093 ;
  assign n16095 = ( x626 & x1158 ) | ( x626 & n16030 ) | ( x1158 & n16030 ) ;
  assign n16096 = ( ~x1158 & n16093 ) | ( ~x1158 & n16095 ) | ( n16093 & n16095 ) ;
  assign n16097 = ( ~x626 & n16095 ) | ( ~x626 & n16096 ) | ( n16095 & n16096 ) ;
  assign n16098 = x788 & n16097 ;
  assign n16099 = n16094 | n16098 ;
  assign n16100 = n15134 | n16099 ;
  assign n16101 = n15134 & ~n16030 ;
  assign n16102 = n16100 & ~n16101 ;
  assign n16103 = ( x647 & x1157 ) | ( x647 & ~n16102 ) | ( x1157 & ~n16102 ) ;
  assign n16104 = ~x628 & n1290 ;
  assign n16105 = n16050 | n16104 ;
  assign n16106 = x1156 & n16105 ;
  assign n16107 = x629 | n16106 ;
  assign n16108 = ( x628 & x1156 ) | ( x628 & ~n16099 ) | ( x1156 & ~n16099 ) ;
  assign n16109 = ~x626 & x1158 ;
  assign n16110 = x626 & ~x1158 ;
  assign n16111 = n16109 | n16110 ;
  assign n16112 = ~x626 & x641 ;
  assign n16113 = x626 & ~x641 ;
  assign n16114 = n16112 | n16113 ;
  assign n16115 = n16111 & n16114 ;
  assign n16116 = ~n16048 & n16115 ;
  assign n16117 = n15420 & ~n16097 ;
  assign n16118 = n16116 | n16117 ;
  assign n16119 = x788 & n16118 ;
  assign n16120 = x648 & ~n16090 ;
  assign n16121 = ( x619 & x1159 ) | ( x619 & n16046 ) | ( x1159 & n16046 ) ;
  assign n16122 = x627 | n16077 ;
  assign n16123 = ( x618 & x1154 ) | ( x618 & ~n16044 ) | ( x1154 & ~n16044 ) ;
  assign n16124 = x660 | n16067 ;
  assign n16125 = ( x609 & x1155 ) | ( x609 & ~n16042 ) | ( x1155 & ~n16042 ) ;
  assign n16126 = n14839 | n16033 ;
  assign n16127 = x625 & ~n16126 ;
  assign n16128 = n16062 & n16126 ;
  assign n16129 = n16127 | n16128 ;
  assign n16130 = n16038 & n16129 ;
  assign n16131 = x608 | n16037 ;
  assign n16132 = n16130 | n16131 ;
  assign n16133 = x1153 & n16062 ;
  assign n16134 = ~n16127 & n16133 ;
  assign n16135 = x608 & ~n16039 ;
  assign n16136 = ~n16134 & n16135 ;
  assign n16137 = n16132 & ~n16136 ;
  assign n16138 = x778 & ~n16137 ;
  assign n16139 = x778 | n16128 ;
  assign n16140 = ~n16138 & n16139 ;
  assign n16141 = ( x609 & ~x1155 ) | ( x609 & n16140 ) | ( ~x1155 & n16140 ) ;
  assign n16142 = ~n16125 & n16141 ;
  assign n16143 = n16124 | n16142 ;
  assign n16144 = x660 & ~n16070 ;
  assign n16145 = ( x609 & x1155 ) | ( x609 & n16042 ) | ( x1155 & n16042 ) ;
  assign n16146 = ( ~x609 & x1155 ) | ( ~x609 & n16140 ) | ( x1155 & n16140 ) ;
  assign n16147 = n16145 & n16146 ;
  assign n16148 = n16144 & ~n16147 ;
  assign n16149 = n16143 & ~n16148 ;
  assign n16150 = x785 & ~n16149 ;
  assign n16151 = x785 | n16140 ;
  assign n16152 = ~n16150 & n16151 ;
  assign n16153 = ( x618 & ~x1154 ) | ( x618 & n16152 ) | ( ~x1154 & n16152 ) ;
  assign n16154 = ~n16123 & n16153 ;
  assign n16155 = n16122 | n16154 ;
  assign n16156 = x627 & ~n16080 ;
  assign n16157 = ( x618 & x1154 ) | ( x618 & n16044 ) | ( x1154 & n16044 ) ;
  assign n16158 = ( ~x618 & x1154 ) | ( ~x618 & n16152 ) | ( x1154 & n16152 ) ;
  assign n16159 = n16157 & n16158 ;
  assign n16160 = n16156 & ~n16159 ;
  assign n16161 = n16155 & ~n16160 ;
  assign n16162 = x781 & ~n16161 ;
  assign n16163 = x781 | n16152 ;
  assign n16164 = ~n16162 & n16163 ;
  assign n16165 = ( ~x619 & x1159 ) | ( ~x619 & n16164 ) | ( x1159 & n16164 ) ;
  assign n16166 = n16121 & n16165 ;
  assign n16167 = n16120 & ~n16166 ;
  assign n16168 = x648 | n16087 ;
  assign n16169 = ( x619 & x1159 ) | ( x619 & ~n16046 ) | ( x1159 & ~n16046 ) ;
  assign n16170 = ( x619 & ~x1159 ) | ( x619 & n16164 ) | ( ~x1159 & n16164 ) ;
  assign n16171 = ~n16169 & n16170 ;
  assign n16172 = n16168 | n16171 ;
  assign n16173 = x789 & n16172 ;
  assign n16174 = ~n16167 & n16173 ;
  assign n16175 = ~x789 & n16164 ;
  assign n16176 = x788 & n16111 ;
  assign n16177 = n15421 | n16176 ;
  assign n16178 = n16175 | n16177 ;
  assign n16179 = n16174 | n16178 ;
  assign n16180 = ~n16119 & n16179 ;
  assign n16181 = ( x628 & ~x1156 ) | ( x628 & n16180 ) | ( ~x1156 & n16180 ) ;
  assign n16182 = ~n16108 & n16181 ;
  assign n16183 = n16107 | n16182 ;
  assign n16184 = x628 & n1290 ;
  assign n16185 = n16050 | n16184 ;
  assign n16186 = ~x1156 & n16185 ;
  assign n16187 = x629 & ~n16186 ;
  assign n16188 = ( x628 & x1156 ) | ( x628 & n16099 ) | ( x1156 & n16099 ) ;
  assign n16189 = ( ~x628 & x1156 ) | ( ~x628 & n16180 ) | ( x1156 & n16180 ) ;
  assign n16190 = n16188 & n16189 ;
  assign n16191 = n16187 & ~n16190 ;
  assign n16192 = n16183 & ~n16191 ;
  assign n16193 = x792 & ~n16192 ;
  assign n16194 = x792 | n16180 ;
  assign n16195 = ~n16193 & n16194 ;
  assign n16196 = ( x647 & ~x1157 ) | ( x647 & n16195 ) | ( ~x1157 & n16195 ) ;
  assign n16197 = ~n16103 & n16196 ;
  assign n16198 = n16059 | n16197 ;
  assign n16199 = ( x647 & x1157 ) | ( x647 & ~n16030 ) | ( x1157 & ~n16030 ) ;
  assign n16200 = ( x647 & ~x1157 ) | ( x647 & n16056 ) | ( ~x1157 & n16056 ) ;
  assign n16201 = ~n16199 & n16200 ;
  assign n16202 = x630 & ~n16201 ;
  assign n16203 = ( x647 & x1157 ) | ( x647 & n16102 ) | ( x1157 & n16102 ) ;
  assign n16204 = ( ~x647 & x1157 ) | ( ~x647 & n16195 ) | ( x1157 & n16195 ) ;
  assign n16205 = n16203 & n16204 ;
  assign n16206 = n16202 & ~n16205 ;
  assign n16207 = n16198 & ~n16206 ;
  assign n16208 = x787 & ~n16207 ;
  assign n16209 = x787 | n16195 ;
  assign n16210 = ~n16208 & n16209 ;
  assign n16211 = ( x790 & x832 ) | ( x790 & n16210 ) | ( x832 & n16210 ) ;
  assign n16212 = n15141 & n16030 ;
  assign n16213 = ~n15141 & n16102 ;
  assign n16214 = n16212 | n16213 ;
  assign n16215 = ( x644 & x715 ) | ( x644 & ~n16214 ) | ( x715 & ~n16214 ) ;
  assign n16216 = ( x644 & ~x715 ) | ( x644 & n16030 ) | ( ~x715 & n16030 ) ;
  assign n16217 = ~n16215 & n16216 ;
  assign n16218 = x1160 & ~n16217 ;
  assign n16219 = ~x787 & n16056 ;
  assign n16220 = n16058 | n16201 ;
  assign n16221 = x787 & n16220 ;
  assign n16222 = n16219 | n16221 ;
  assign n16223 = ( x644 & x715 ) | ( x644 & n16222 ) | ( x715 & n16222 ) ;
  assign n16224 = ( ~x644 & x715 ) | ( ~x644 & n16210 ) | ( x715 & n16210 ) ;
  assign n16225 = n16223 & n16224 ;
  assign n16226 = n16218 & ~n16225 ;
  assign n16227 = ( x644 & x715 ) | ( x644 & n16214 ) | ( x715 & n16214 ) ;
  assign n16228 = ( ~x644 & x715 ) | ( ~x644 & n16030 ) | ( x715 & n16030 ) ;
  assign n16229 = n16227 & n16228 ;
  assign n16230 = x1160 | n16229 ;
  assign n16231 = ( x644 & x715 ) | ( x644 & ~n16222 ) | ( x715 & ~n16222 ) ;
  assign n16232 = ( x644 & ~x715 ) | ( x644 & n16210 ) | ( ~x715 & n16210 ) ;
  assign n16233 = ~n16231 & n16232 ;
  assign n16234 = n16230 | n16233 ;
  assign n16235 = ~n16226 & n16234 ;
  assign n16236 = ( ~x790 & x832 ) | ( ~x790 & n16235 ) | ( x832 & n16235 ) ;
  assign n16237 = n16211 & n16236 ;
  assign n16238 = n16029 | n16237 ;
  assign n16239 = x141 | n14834 ;
  assign n16240 = n15141 & n16239 ;
  assign n16241 = ( x626 & x1158 ) | ( x626 & ~n16239 ) | ( x1158 & ~n16239 ) ;
  assign n16242 = x141 & n2032 ;
  assign n16243 = x141 | n15070 ;
  assign n16244 = x749 & n15072 ;
  assign n16245 = n16243 & ~n16244 ;
  assign n16246 = x38 & ~n16245 ;
  assign n16247 = ~x749 & n14710 ;
  assign n16248 = x141 & ~n14907 ;
  assign n16249 = n16247 | n16248 ;
  assign n16250 = x39 & n16249 ;
  assign n16251 = x141 | x749 ;
  assign n16252 = n14823 | n16251 ;
  assign n16253 = ( ~x141 & x749 ) | ( ~x141 & n14932 ) | ( x749 & n14932 ) ;
  assign n16254 = ( x141 & x749 ) | ( x141 & ~n15063 ) | ( x749 & ~n15063 ) ;
  assign n16255 = n16253 & n16254 ;
  assign n16256 = n16252 & ~n16255 ;
  assign n16257 = x38 | n16256 ;
  assign n16258 = n16250 | n16257 ;
  assign n16259 = ~n16246 & n16258 ;
  assign n16260 = ~n2032 & n16259 ;
  assign n16261 = n16242 | n16260 ;
  assign n16262 = ~n15082 & n16261 ;
  assign n16263 = n15082 & n16239 ;
  assign n16264 = n16262 | n16263 ;
  assign n16265 = ~x785 & n16264 ;
  assign n16266 = ~n15088 & n16239 ;
  assign n16267 = x609 & n16262 ;
  assign n16268 = n16266 | n16267 ;
  assign n16269 = x1155 & n16268 ;
  assign n16270 = n15094 & n16239 ;
  assign n16271 = ~x609 & n16262 ;
  assign n16272 = n16270 | n16271 ;
  assign n16273 = ~x1155 & n16272 ;
  assign n16274 = n16269 | n16273 ;
  assign n16275 = x785 & n16274 ;
  assign n16276 = n16265 | n16275 ;
  assign n16277 = ~x781 & n16276 ;
  assign n16278 = ( x618 & x1154 ) | ( x618 & n16239 ) | ( x1154 & n16239 ) ;
  assign n16279 = ( ~x618 & x1154 ) | ( ~x618 & n16276 ) | ( x1154 & n16276 ) ;
  assign n16280 = n16278 & n16279 ;
  assign n16281 = ( x618 & x1154 ) | ( x618 & ~n16239 ) | ( x1154 & ~n16239 ) ;
  assign n16282 = ( x618 & ~x1154 ) | ( x618 & n16276 ) | ( ~x1154 & n16276 ) ;
  assign n16283 = ~n16281 & n16282 ;
  assign n16284 = n16280 | n16283 ;
  assign n16285 = x781 & n16284 ;
  assign n16286 = n16277 | n16285 ;
  assign n16287 = ~x789 & n16286 ;
  assign n16288 = ( x619 & x1159 ) | ( x619 & n16239 ) | ( x1159 & n16239 ) ;
  assign n16289 = ( ~x619 & x1159 ) | ( ~x619 & n16286 ) | ( x1159 & n16286 ) ;
  assign n16290 = n16288 & n16289 ;
  assign n16291 = ( x619 & x1159 ) | ( x619 & ~n16239 ) | ( x1159 & ~n16239 ) ;
  assign n16292 = ( x619 & ~x1159 ) | ( x619 & n16286 ) | ( ~x1159 & n16286 ) ;
  assign n16293 = ~n16291 & n16292 ;
  assign n16294 = n16290 | n16293 ;
  assign n16295 = x789 & n16294 ;
  assign n16296 = n16287 | n16295 ;
  assign n16297 = ( x626 & ~x1158 ) | ( x626 & n16296 ) | ( ~x1158 & n16296 ) ;
  assign n16298 = ~n16241 & n16297 ;
  assign n16299 = ( x626 & x1158 ) | ( x626 & n16239 ) | ( x1158 & n16239 ) ;
  assign n16300 = ( ~x626 & x1158 ) | ( ~x626 & n16296 ) | ( x1158 & n16296 ) ;
  assign n16301 = n16299 & n16300 ;
  assign n16302 = n16298 | n16301 ;
  assign n16303 = x788 & n16302 ;
  assign n16304 = ~x788 & n16296 ;
  assign n16305 = n16303 | n16304 ;
  assign n16306 = n15134 | n16305 ;
  assign n16307 = n15134 & ~n16239 ;
  assign n16308 = n16306 & ~n16307 ;
  assign n16309 = ~n15141 & n16308 ;
  assign n16310 = n16240 | n16309 ;
  assign n16311 = ( x644 & x715 ) | ( x644 & n16310 ) | ( x715 & n16310 ) ;
  assign n16312 = ( ~x644 & x715 ) | ( ~x644 & n16239 ) | ( x715 & n16239 ) ;
  assign n16313 = n16311 & n16312 ;
  assign n16314 = x1160 | n16313 ;
  assign n16315 = n15414 & n16239 ;
  assign n16316 = n15375 & n16243 ;
  assign n16317 = x706 & ~n16316 ;
  assign n16318 = ~x39 & n15345 ;
  assign n16319 = n15325 | n16318 ;
  assign n16320 = ( ~x38 & x141 ) | ( ~x38 & n16319 ) | ( x141 & n16319 ) ;
  assign n16321 = x39 & n15221 ;
  assign n16322 = ~x39 & n15369 ;
  assign n16323 = n16321 | n16322 ;
  assign n16324 = ( x38 & x141 ) | ( x38 & n16323 ) | ( x141 & n16323 ) ;
  assign n16325 = n16320 & ~n16324 ;
  assign n16326 = n16317 & ~n16325 ;
  assign n16327 = x141 | x706 ;
  assign n16328 = n15382 | n16327 ;
  assign n16329 = ~n2032 & n16328 ;
  assign n16330 = ~n16326 & n16329 ;
  assign n16331 = n16242 | n16330 ;
  assign n16332 = ~x778 & n16331 ;
  assign n16333 = ( x625 & x1153 ) | ( x625 & n16239 ) | ( x1153 & n16239 ) ;
  assign n16334 = ( ~x625 & x1153 ) | ( ~x625 & n16331 ) | ( x1153 & n16331 ) ;
  assign n16335 = n16333 & n16334 ;
  assign n16336 = ( x625 & x1153 ) | ( x625 & ~n16239 ) | ( x1153 & ~n16239 ) ;
  assign n16337 = ( x625 & ~x1153 ) | ( x625 & n16331 ) | ( ~x1153 & n16331 ) ;
  assign n16338 = ~n16336 & n16337 ;
  assign n16339 = n16335 | n16338 ;
  assign n16340 = x778 & n16339 ;
  assign n16341 = n16332 | n16340 ;
  assign n16342 = ~n15400 & n16341 ;
  assign n16343 = n15400 & n16239 ;
  assign n16344 = n16342 | n16343 ;
  assign n16345 = n15407 | n16344 ;
  assign n16346 = n15407 & ~n16239 ;
  assign n16347 = n16345 & ~n16346 ;
  assign n16348 = ~n15414 & n16347 ;
  assign n16349 = n16315 | n16348 ;
  assign n16350 = n15421 | n16349 ;
  assign n16351 = n15421 & ~n16239 ;
  assign n16352 = n16350 & ~n16351 ;
  assign n16353 = ~x792 & n16352 ;
  assign n16354 = ( x628 & x1156 ) | ( x628 & n16239 ) | ( x1156 & n16239 ) ;
  assign n16355 = ( ~x628 & x1156 ) | ( ~x628 & n16352 ) | ( x1156 & n16352 ) ;
  assign n16356 = n16354 & n16355 ;
  assign n16357 = ( x628 & x1156 ) | ( x628 & ~n16239 ) | ( x1156 & ~n16239 ) ;
  assign n16358 = ( x628 & ~x1156 ) | ( x628 & n16352 ) | ( ~x1156 & n16352 ) ;
  assign n16359 = ~n16357 & n16358 ;
  assign n16360 = n16356 | n16359 ;
  assign n16361 = x792 & n16360 ;
  assign n16362 = n16353 | n16361 ;
  assign n16363 = ~x787 & n16362 ;
  assign n16364 = ( x647 & x1157 ) | ( x647 & n16239 ) | ( x1157 & n16239 ) ;
  assign n16365 = ( ~x647 & x1157 ) | ( ~x647 & n16362 ) | ( x1157 & n16362 ) ;
  assign n16366 = n16364 & n16365 ;
  assign n16367 = ( x647 & x1157 ) | ( x647 & ~n16239 ) | ( x1157 & ~n16239 ) ;
  assign n16368 = ( x647 & ~x1157 ) | ( x647 & n16362 ) | ( ~x1157 & n16362 ) ;
  assign n16369 = ~n16367 & n16368 ;
  assign n16370 = n16366 | n16369 ;
  assign n16371 = x787 & n16370 ;
  assign n16372 = n16363 | n16371 ;
  assign n16373 = ( x644 & x715 ) | ( x644 & ~n16372 ) | ( x715 & ~n16372 ) ;
  assign n16374 = x630 | n16366 ;
  assign n16375 = ( x647 & x1157 ) | ( x647 & ~n16308 ) | ( x1157 & ~n16308 ) ;
  assign n16376 = x629 | n16356 ;
  assign n16377 = ( x628 & x1156 ) | ( x628 & ~n16305 ) | ( x1156 & ~n16305 ) ;
  assign n16378 = x648 | n16290 ;
  assign n16379 = ( x619 & x1159 ) | ( x619 & ~n16347 ) | ( x1159 & ~n16347 ) ;
  assign n16380 = x627 | n16280 ;
  assign n16381 = ( x618 & x1154 ) | ( x618 & ~n16344 ) | ( x1154 & ~n16344 ) ;
  assign n16382 = x660 | n16269 ;
  assign n16383 = ( x609 & x1155 ) | ( x609 & ~n16341 ) | ( x1155 & ~n16341 ) ;
  assign n16384 = x608 | n16335 ;
  assign n16385 = ( x625 & x1153 ) | ( x625 & ~n16261 ) | ( x1153 & ~n16261 ) ;
  assign n16386 = ( x141 & ~x749 ) | ( x141 & n15872 ) | ( ~x749 & n15872 ) ;
  assign n16387 = ( x141 & x749 ) | ( x141 & n15797 ) | ( x749 & n15797 ) ;
  assign n16388 = ~n16386 & n16387 ;
  assign n16389 = x39 & ~n16388 ;
  assign n16390 = ( x141 & ~x749 ) | ( x141 & n15699 ) | ( ~x749 & n15699 ) ;
  assign n16391 = ( x141 & x749 ) | ( x141 & n15583 ) | ( x749 & n15583 ) ;
  assign n16392 = n16390 & ~n16391 ;
  assign n16393 = n16389 & ~n16392 ;
  assign n16394 = ( x141 & ~x749 ) | ( x141 & n15891 ) | ( ~x749 & n15891 ) ;
  assign n16395 = ( x141 & x749 ) | ( x141 & n15887 ) | ( x749 & n15887 ) ;
  assign n16396 = n16394 & ~n16395 ;
  assign n16397 = ( x141 & ~x749 ) | ( x141 & n15897 ) | ( ~x749 & n15897 ) ;
  assign n16398 = ( x141 & x749 ) | ( x141 & n15894 ) | ( x749 & n15894 ) ;
  assign n16399 = ~n16397 & n16398 ;
  assign n16400 = n16396 | n16399 ;
  assign n16401 = ( ~x38 & n9138 ) | ( ~x38 & n16400 ) | ( n9138 & n16400 ) ;
  assign n16402 = ~n16393 & n16401 ;
  assign n16403 = ~x39 & n15913 ;
  assign n16404 = x38 & ~n16403 ;
  assign n16405 = n16245 & n16404 ;
  assign n16406 = x706 & ~n16405 ;
  assign n16407 = ~n16402 & n16406 ;
  assign n16408 = x706 | n16259 ;
  assign n16409 = ~n2032 & n16408 ;
  assign n16410 = ~n16407 & n16409 ;
  assign n16411 = n16242 | n16410 ;
  assign n16412 = ( x625 & ~x1153 ) | ( x625 & n16411 ) | ( ~x1153 & n16411 ) ;
  assign n16413 = ~n16385 & n16412 ;
  assign n16414 = n16384 | n16413 ;
  assign n16415 = x608 & ~n16338 ;
  assign n16416 = ( x625 & x1153 ) | ( x625 & n16261 ) | ( x1153 & n16261 ) ;
  assign n16417 = ( ~x625 & x1153 ) | ( ~x625 & n16411 ) | ( x1153 & n16411 ) ;
  assign n16418 = n16416 & n16417 ;
  assign n16419 = n16415 & ~n16418 ;
  assign n16420 = n16414 & ~n16419 ;
  assign n16421 = x778 & ~n16420 ;
  assign n16422 = x778 | n16411 ;
  assign n16423 = ~n16421 & n16422 ;
  assign n16424 = ( x609 & ~x1155 ) | ( x609 & n16423 ) | ( ~x1155 & n16423 ) ;
  assign n16425 = ~n16383 & n16424 ;
  assign n16426 = n16382 | n16425 ;
  assign n16427 = x660 & ~n16273 ;
  assign n16428 = ( x609 & x1155 ) | ( x609 & n16341 ) | ( x1155 & n16341 ) ;
  assign n16429 = ( ~x609 & x1155 ) | ( ~x609 & n16423 ) | ( x1155 & n16423 ) ;
  assign n16430 = n16428 & n16429 ;
  assign n16431 = n16427 & ~n16430 ;
  assign n16432 = n16426 & ~n16431 ;
  assign n16433 = x785 & ~n16432 ;
  assign n16434 = x785 | n16423 ;
  assign n16435 = ~n16433 & n16434 ;
  assign n16436 = ( x618 & ~x1154 ) | ( x618 & n16435 ) | ( ~x1154 & n16435 ) ;
  assign n16437 = ~n16381 & n16436 ;
  assign n16438 = n16380 | n16437 ;
  assign n16439 = x627 & ~n16283 ;
  assign n16440 = ( x618 & x1154 ) | ( x618 & n16344 ) | ( x1154 & n16344 ) ;
  assign n16441 = ( ~x618 & x1154 ) | ( ~x618 & n16435 ) | ( x1154 & n16435 ) ;
  assign n16442 = n16440 & n16441 ;
  assign n16443 = n16439 & ~n16442 ;
  assign n16444 = n16438 & ~n16443 ;
  assign n16445 = x781 & ~n16444 ;
  assign n16446 = x781 | n16435 ;
  assign n16447 = ~n16445 & n16446 ;
  assign n16448 = ( x619 & ~x1159 ) | ( x619 & n16447 ) | ( ~x1159 & n16447 ) ;
  assign n16449 = ~n16379 & n16448 ;
  assign n16450 = n16378 | n16449 ;
  assign n16451 = x648 & ~n16293 ;
  assign n16452 = ( x619 & x1159 ) | ( x619 & n16347 ) | ( x1159 & n16347 ) ;
  assign n16453 = ( ~x619 & x1159 ) | ( ~x619 & n16447 ) | ( x1159 & n16447 ) ;
  assign n16454 = n16452 & n16453 ;
  assign n16455 = n16451 & ~n16454 ;
  assign n16456 = n16450 & ~n16455 ;
  assign n16457 = x789 & ~n16456 ;
  assign n16458 = x789 | n16447 ;
  assign n16459 = ~n16457 & n16458 ;
  assign n16460 = ~x788 & n16459 ;
  assign n16461 = n15972 & ~n16298 ;
  assign n16462 = ( x626 & x641 ) | ( x626 & n16349 ) | ( x641 & n16349 ) ;
  assign n16463 = ( ~x626 & x641 ) | ( ~x626 & n16459 ) | ( x641 & n16459 ) ;
  assign n16464 = n16462 | n16463 ;
  assign n16465 = ~n16461 & n16464 ;
  assign n16466 = n15978 | n16301 ;
  assign n16467 = ( x626 & x641 ) | ( x626 & ~n16349 ) | ( x641 & ~n16349 ) ;
  assign n16468 = ( x626 & ~x641 ) | ( x626 & n16459 ) | ( ~x641 & n16459 ) ;
  assign n16469 = n16467 & ~n16468 ;
  assign n16470 = n16466 & ~n16469 ;
  assign n16471 = n16465 | n16470 ;
  assign n16472 = x788 & n16471 ;
  assign n16473 = n16460 | n16472 ;
  assign n16474 = ( x628 & ~x1156 ) | ( x628 & n16473 ) | ( ~x1156 & n16473 ) ;
  assign n16475 = ~n16377 & n16474 ;
  assign n16476 = n16376 | n16475 ;
  assign n16477 = x629 & ~n16359 ;
  assign n16478 = ( x628 & x1156 ) | ( x628 & n16305 ) | ( x1156 & n16305 ) ;
  assign n16479 = ( ~x628 & x1156 ) | ( ~x628 & n16473 ) | ( x1156 & n16473 ) ;
  assign n16480 = n16478 & n16479 ;
  assign n16481 = n16477 & ~n16480 ;
  assign n16482 = n16476 & ~n16481 ;
  assign n16483 = x792 & ~n16482 ;
  assign n16484 = x792 | n16473 ;
  assign n16485 = ~n16483 & n16484 ;
  assign n16486 = ( x647 & ~x1157 ) | ( x647 & n16485 ) | ( ~x1157 & n16485 ) ;
  assign n16487 = ~n16375 & n16486 ;
  assign n16488 = n16374 | n16487 ;
  assign n16489 = x630 & ~n16369 ;
  assign n16490 = ( x647 & x1157 ) | ( x647 & n16308 ) | ( x1157 & n16308 ) ;
  assign n16491 = ( ~x647 & x1157 ) | ( ~x647 & n16485 ) | ( x1157 & n16485 ) ;
  assign n16492 = n16490 & n16491 ;
  assign n16493 = n16489 & ~n16492 ;
  assign n16494 = n16488 & ~n16493 ;
  assign n16495 = x787 & ~n16494 ;
  assign n16496 = x787 | n16485 ;
  assign n16497 = ~n16495 & n16496 ;
  assign n16498 = ( x644 & ~x715 ) | ( x644 & n16497 ) | ( ~x715 & n16497 ) ;
  assign n16499 = ~n16373 & n16498 ;
  assign n16500 = n16314 | n16499 ;
  assign n16501 = ( x644 & x715 ) | ( x644 & ~n16310 ) | ( x715 & ~n16310 ) ;
  assign n16502 = ( x644 & ~x715 ) | ( x644 & n16239 ) | ( ~x715 & n16239 ) ;
  assign n16503 = ~n16501 & n16502 ;
  assign n16504 = x1160 & ~n16503 ;
  assign n16505 = ( x644 & x715 ) | ( x644 & n16372 ) | ( x715 & n16372 ) ;
  assign n16506 = ( ~x644 & x715 ) | ( ~x644 & n16497 ) | ( x715 & n16497 ) ;
  assign n16507 = n16505 & n16506 ;
  assign n16508 = n16504 & ~n16507 ;
  assign n16509 = x790 & ~n16508 ;
  assign n16510 = n16500 & n16509 ;
  assign n16511 = ~x790 & n16497 ;
  assign n16512 = n6785 | n16511 ;
  assign n16513 = n16510 | n16512 ;
  assign n16514 = ~x141 & n6785 ;
  assign n16515 = x832 | n16514 ;
  assign n16516 = n16513 & ~n16515 ;
  assign n16517 = x141 | n1290 ;
  assign n16518 = ( x647 & x1157 ) | ( x647 & n16517 ) | ( x1157 & n16517 ) ;
  assign n16519 = x706 & n15202 ;
  assign n16520 = n16517 & ~n16519 ;
  assign n16521 = ~x778 & n16520 ;
  assign n16522 = ~x625 & n16519 ;
  assign n16523 = n16520 | n16522 ;
  assign n16524 = x1153 & n16523 ;
  assign n16525 = ~x1153 & n16517 ;
  assign n16526 = ~n16522 & n16525 ;
  assign n16527 = n16524 | n16526 ;
  assign n16528 = x778 & n16527 ;
  assign n16529 = n16521 | n16528 ;
  assign n16530 = n16043 | n16529 ;
  assign n16531 = n16045 | n16530 ;
  assign n16532 = n16047 | n16531 ;
  assign n16533 = n16049 | n16532 ;
  assign n16534 = n16055 | n16533 ;
  assign n16535 = ( ~x647 & x1157 ) | ( ~x647 & n16534 ) | ( x1157 & n16534 ) ;
  assign n16536 = n16518 & n16535 ;
  assign n16537 = x630 | n16536 ;
  assign n16538 = x749 & n14840 ;
  assign n16539 = n16517 & ~n16538 ;
  assign n16540 = n16060 | n16539 ;
  assign n16541 = ~x785 & n16540 ;
  assign n16542 = n16065 | n16539 ;
  assign n16543 = x1155 & n16542 ;
  assign n16544 = n16068 | n16540 ;
  assign n16545 = ~x1155 & n16544 ;
  assign n16546 = n16543 | n16545 ;
  assign n16547 = x785 & n16546 ;
  assign n16548 = n16541 | n16547 ;
  assign n16549 = ~x781 & n16548 ;
  assign n16550 = n16075 | n16548 ;
  assign n16551 = x1154 & n16550 ;
  assign n16552 = n16078 | n16548 ;
  assign n16553 = ~x1154 & n16552 ;
  assign n16554 = n16551 | n16553 ;
  assign n16555 = x781 & n16554 ;
  assign n16556 = n16549 | n16555 ;
  assign n16557 = ~x789 & n16556 ;
  assign n16558 = ( x619 & x1159 ) | ( x619 & n16517 ) | ( x1159 & n16517 ) ;
  assign n16559 = ( ~x619 & x1159 ) | ( ~x619 & n16556 ) | ( x1159 & n16556 ) ;
  assign n16560 = n16558 & n16559 ;
  assign n16561 = ( x619 & x1159 ) | ( x619 & ~n16517 ) | ( x1159 & ~n16517 ) ;
  assign n16562 = ( x619 & ~x1159 ) | ( x619 & n16556 ) | ( ~x1159 & n16556 ) ;
  assign n16563 = ~n16561 & n16562 ;
  assign n16564 = n16560 | n16563 ;
  assign n16565 = x789 & n16564 ;
  assign n16566 = n16557 | n16565 ;
  assign n16567 = ~x788 & n16566 ;
  assign n16568 = ( x626 & x1158 ) | ( x626 & n16517 ) | ( x1158 & n16517 ) ;
  assign n16569 = ( ~x1158 & n16566 ) | ( ~x1158 & n16568 ) | ( n16566 & n16568 ) ;
  assign n16570 = ( ~x626 & n16568 ) | ( ~x626 & n16569 ) | ( n16568 & n16569 ) ;
  assign n16571 = x788 & n16570 ;
  assign n16572 = n16567 | n16571 ;
  assign n16573 = n15134 | n16572 ;
  assign n16574 = n15134 & ~n16517 ;
  assign n16575 = n16573 & ~n16574 ;
  assign n16576 = ( x647 & x1157 ) | ( x647 & ~n16575 ) | ( x1157 & ~n16575 ) ;
  assign n16577 = ( x628 & x1156 ) | ( x628 & ~n16572 ) | ( x1156 & ~n16572 ) ;
  assign n16578 = n16115 & ~n16532 ;
  assign n16579 = n15420 & ~n16570 ;
  assign n16580 = n16578 | n16579 ;
  assign n16581 = x788 & n16580 ;
  assign n16582 = x648 & ~n16563 ;
  assign n16583 = ( x619 & x1159 ) | ( x619 & n16531 ) | ( x1159 & n16531 ) ;
  assign n16584 = x627 | n16551 ;
  assign n16585 = ( x618 & x1154 ) | ( x618 & ~n16530 ) | ( x1154 & ~n16530 ) ;
  assign n16586 = x660 | n16543 ;
  assign n16587 = ( x609 & x1155 ) | ( x609 & ~n16529 ) | ( x1155 & ~n16529 ) ;
  assign n16588 = n14839 | n16520 ;
  assign n16589 = x625 & ~n16588 ;
  assign n16590 = n16539 & n16588 ;
  assign n16591 = n16589 | n16590 ;
  assign n16592 = n16525 & n16591 ;
  assign n16593 = x608 | n16524 ;
  assign n16594 = n16592 | n16593 ;
  assign n16595 = x1153 & n16539 ;
  assign n16596 = ~n16589 & n16595 ;
  assign n16597 = x608 & ~n16526 ;
  assign n16598 = ~n16596 & n16597 ;
  assign n16599 = n16594 & ~n16598 ;
  assign n16600 = x778 & ~n16599 ;
  assign n16601 = x778 | n16590 ;
  assign n16602 = ~n16600 & n16601 ;
  assign n16603 = ( x609 & ~x1155 ) | ( x609 & n16602 ) | ( ~x1155 & n16602 ) ;
  assign n16604 = ~n16587 & n16603 ;
  assign n16605 = n16586 | n16604 ;
  assign n16606 = x660 & ~n16545 ;
  assign n16607 = ( x609 & x1155 ) | ( x609 & n16529 ) | ( x1155 & n16529 ) ;
  assign n16608 = ( ~x609 & x1155 ) | ( ~x609 & n16602 ) | ( x1155 & n16602 ) ;
  assign n16609 = n16607 & n16608 ;
  assign n16610 = n16606 & ~n16609 ;
  assign n16611 = n16605 & ~n16610 ;
  assign n16612 = x785 & ~n16611 ;
  assign n16613 = x785 | n16602 ;
  assign n16614 = ~n16612 & n16613 ;
  assign n16615 = ( x618 & ~x1154 ) | ( x618 & n16614 ) | ( ~x1154 & n16614 ) ;
  assign n16616 = ~n16585 & n16615 ;
  assign n16617 = n16584 | n16616 ;
  assign n16618 = x627 & ~n16553 ;
  assign n16619 = ( x618 & x1154 ) | ( x618 & n16530 ) | ( x1154 & n16530 ) ;
  assign n16620 = ( ~x618 & x1154 ) | ( ~x618 & n16614 ) | ( x1154 & n16614 ) ;
  assign n16621 = n16619 & n16620 ;
  assign n16622 = n16618 & ~n16621 ;
  assign n16623 = n16617 & ~n16622 ;
  assign n16624 = x781 & ~n16623 ;
  assign n16625 = x781 | n16614 ;
  assign n16626 = ~n16624 & n16625 ;
  assign n16627 = ( ~x619 & x1159 ) | ( ~x619 & n16626 ) | ( x1159 & n16626 ) ;
  assign n16628 = n16583 & n16627 ;
  assign n16629 = n16582 & ~n16628 ;
  assign n16630 = x648 | n16560 ;
  assign n16631 = ( x619 & x1159 ) | ( x619 & ~n16531 ) | ( x1159 & ~n16531 ) ;
  assign n16632 = ( x619 & ~x1159 ) | ( x619 & n16626 ) | ( ~x1159 & n16626 ) ;
  assign n16633 = ~n16631 & n16632 ;
  assign n16634 = n16630 | n16633 ;
  assign n16635 = x789 & n16634 ;
  assign n16636 = ~n16629 & n16635 ;
  assign n16637 = ~x789 & n16626 ;
  assign n16638 = n16177 | n16637 ;
  assign n16639 = n16636 | n16638 ;
  assign n16640 = ~n16581 & n16639 ;
  assign n16641 = ( x628 & ~x1156 ) | ( x628 & n16640 ) | ( ~x1156 & n16640 ) ;
  assign n16642 = ~n16577 & n16641 ;
  assign n16643 = x1156 & ~n16104 ;
  assign n16644 = ~n16533 & n16643 ;
  assign n16645 = ( x629 & x1156 ) | ( x629 & ~n16644 ) | ( x1156 & ~n16644 ) ;
  assign n16646 = n16642 | n16645 ;
  assign n16647 = ( x628 & x1156 ) | ( x628 & n16572 ) | ( x1156 & n16572 ) ;
  assign n16648 = ( ~x628 & x1156 ) | ( ~x628 & n16640 ) | ( x1156 & n16640 ) ;
  assign n16649 = n16647 & n16648 ;
  assign n16650 = x1156 | n16184 ;
  assign n16651 = n16533 | n16650 ;
  assign n16652 = ( x629 & x1156 ) | ( x629 & ~n16651 ) | ( x1156 & ~n16651 ) ;
  assign n16653 = ~n16649 & n16652 ;
  assign n16654 = n16646 & ~n16653 ;
  assign n16655 = x792 & ~n16654 ;
  assign n16656 = x792 | n16640 ;
  assign n16657 = ~n16655 & n16656 ;
  assign n16658 = ( x647 & ~x1157 ) | ( x647 & n16657 ) | ( ~x1157 & n16657 ) ;
  assign n16659 = ~n16576 & n16658 ;
  assign n16660 = n16537 | n16659 ;
  assign n16661 = ( x647 & x1157 ) | ( x647 & ~n16517 ) | ( x1157 & ~n16517 ) ;
  assign n16662 = ( x647 & ~x1157 ) | ( x647 & n16534 ) | ( ~x1157 & n16534 ) ;
  assign n16663 = ~n16661 & n16662 ;
  assign n16664 = x630 & ~n16663 ;
  assign n16665 = ( x647 & x1157 ) | ( x647 & n16575 ) | ( x1157 & n16575 ) ;
  assign n16666 = ( ~x647 & x1157 ) | ( ~x647 & n16657 ) | ( x1157 & n16657 ) ;
  assign n16667 = n16665 & n16666 ;
  assign n16668 = n16664 & ~n16667 ;
  assign n16669 = n16660 & ~n16668 ;
  assign n16670 = x787 & ~n16669 ;
  assign n16671 = x787 | n16657 ;
  assign n16672 = ~n16670 & n16671 ;
  assign n16673 = ( x790 & x832 ) | ( x790 & n16672 ) | ( x832 & n16672 ) ;
  assign n16674 = n15141 & n16517 ;
  assign n16675 = ~n15141 & n16575 ;
  assign n16676 = n16674 | n16675 ;
  assign n16677 = ( x644 & x715 ) | ( x644 & ~n16676 ) | ( x715 & ~n16676 ) ;
  assign n16678 = ( x644 & ~x715 ) | ( x644 & n16517 ) | ( ~x715 & n16517 ) ;
  assign n16679 = ~n16677 & n16678 ;
  assign n16680 = x1160 & ~n16679 ;
  assign n16681 = ~x787 & n16534 ;
  assign n16682 = n16536 | n16663 ;
  assign n16683 = x787 & n16682 ;
  assign n16684 = n16681 | n16683 ;
  assign n16685 = ( x644 & x715 ) | ( x644 & n16684 ) | ( x715 & n16684 ) ;
  assign n16686 = ( ~x644 & x715 ) | ( ~x644 & n16672 ) | ( x715 & n16672 ) ;
  assign n16687 = n16685 & n16686 ;
  assign n16688 = n16680 & ~n16687 ;
  assign n16689 = ( x644 & x715 ) | ( x644 & n16676 ) | ( x715 & n16676 ) ;
  assign n16690 = ( ~x644 & x715 ) | ( ~x644 & n16517 ) | ( x715 & n16517 ) ;
  assign n16691 = n16689 & n16690 ;
  assign n16692 = x1160 | n16691 ;
  assign n16693 = ( x644 & x715 ) | ( x644 & ~n16684 ) | ( x715 & ~n16684 ) ;
  assign n16694 = ( x644 & ~x715 ) | ( x644 & n16672 ) | ( ~x715 & n16672 ) ;
  assign n16695 = ~n16693 & n16694 ;
  assign n16696 = n16692 | n16695 ;
  assign n16697 = ~n16688 & n16696 ;
  assign n16698 = ( ~x790 & x832 ) | ( ~x790 & n16697 ) | ( x832 & n16697 ) ;
  assign n16699 = n16673 & n16698 ;
  assign n16700 = n16516 | n16699 ;
  assign n16701 = x142 & n14828 ;
  assign n16702 = x39 & n14709 ;
  assign n16703 = x142 & ~n14823 ;
  assign n16704 = ~n16702 & n16703 ;
  assign n16705 = n1290 & ~n14481 ;
  assign n16706 = x142 & ~n16705 ;
  assign n16707 = n2203 | n16706 ;
  assign n16708 = ~x215 & n16707 ;
  assign n16709 = n14617 & ~n14619 ;
  assign n16710 = x142 & ~n16709 ;
  assign n16711 = ( ~n2203 & n4721 ) | ( ~n2203 & n16710 ) | ( n4721 & n16710 ) ;
  assign n16712 = n14666 & ~n14679 ;
  assign n16713 = x142 & ~n16712 ;
  assign n16714 = ( n2203 & n4721 ) | ( n2203 & ~n16713 ) | ( n4721 & ~n16713 ) ;
  assign n16715 = ~n16711 & n16714 ;
  assign n16716 = n16708 & ~n16715 ;
  assign n16717 = x142 & ~n14528 ;
  assign n16718 = ( x215 & ~n4721 ) | ( x215 & n16717 ) | ( ~n4721 & n16717 ) ;
  assign n16719 = n14570 & ~n14571 ;
  assign n16720 = x142 & ~n16719 ;
  assign n16721 = ( x215 & n4721 ) | ( x215 & n16720 ) | ( n4721 & n16720 ) ;
  assign n16722 = n16718 & n16721 ;
  assign n16723 = n16716 | n16722 ;
  assign n16724 = n4757 & n16723 ;
  assign n16725 = n16704 | n16724 ;
  assign n16726 = ~n12808 & n16725 ;
  assign n16727 = n16701 | n16726 ;
  assign n16728 = n15141 & n16727 ;
  assign n16729 = ( x626 & x1158 ) | ( x626 & ~n16727 ) | ( x1158 & ~n16727 ) ;
  assign n16730 = x142 & n2032 ;
  assign n16731 = x743 & n14874 ;
  assign n16732 = n16706 | n16731 ;
  assign n16733 = ~n2203 & n16732 ;
  assign n16734 = x215 | n16733 ;
  assign n16735 = x743 | n16710 ;
  assign n16736 = x142 & ~n15022 ;
  assign n16737 = n14846 & n14849 ;
  assign n16738 = x743 & ~n16737 ;
  assign n16739 = ~n16736 & n16738 ;
  assign n16740 = n16735 & ~n16739 ;
  assign n16741 = ( n2203 & ~n4721 ) | ( n2203 & n16740 ) | ( ~n4721 & n16740 ) ;
  assign n16742 = x743 | n16713 ;
  assign n16743 = ~n15029 & n15035 ;
  assign n16744 = ( ~x142 & x743 ) | ( ~x142 & n16743 ) | ( x743 & n16743 ) ;
  assign n16745 = ( x142 & x743 ) | ( x142 & ~n14870 ) | ( x743 & ~n14870 ) ;
  assign n16746 = n16744 & n16745 ;
  assign n16747 = n16742 & ~n16746 ;
  assign n16748 = ( n2203 & n4721 ) | ( n2203 & n16747 ) | ( n4721 & n16747 ) ;
  assign n16749 = n16741 & n16748 ;
  assign n16750 = n16734 | n16749 ;
  assign n16751 = x743 | n16717 ;
  assign n16752 = x142 & ~n14969 ;
  assign n16753 = x743 & ~n15845 ;
  assign n16754 = ~n16752 & n16753 ;
  assign n16755 = n16751 & ~n16754 ;
  assign n16756 = n4721 & n16755 ;
  assign n16757 = x743 | n16720 ;
  assign n16758 = x142 & ~n14990 ;
  assign n16759 = n14881 | n14884 ;
  assign n16760 = x743 & ~n16759 ;
  assign n16761 = ~n16758 & n16760 ;
  assign n16762 = n16757 & ~n16761 ;
  assign n16763 = ( x215 & n15308 ) | ( x215 & ~n16762 ) | ( n15308 & ~n16762 ) ;
  assign n16764 = ~n16756 & n16763 ;
  assign n16765 = n16750 & ~n16764 ;
  assign n16766 = x299 & ~n16765 ;
  assign n16767 = ~n4764 & n16747 ;
  assign n16768 = ( n1823 & n15052 ) | ( n1823 & ~n16740 ) | ( n15052 & ~n16740 ) ;
  assign n16769 = ~n16767 & n16768 ;
  assign n16770 = n1823 | n16732 ;
  assign n16771 = ~x223 & n16770 ;
  assign n16772 = ~n16769 & n16771 ;
  assign n16773 = ( x223 & ~n4764 ) | ( x223 & n16755 ) | ( ~n4764 & n16755 ) ;
  assign n16774 = ( x223 & n4764 ) | ( x223 & n16762 ) | ( n4764 & n16762 ) ;
  assign n16775 = n16773 & n16774 ;
  assign n16776 = n16772 | n16775 ;
  assign n16777 = ( x39 & n4757 ) | ( x39 & n16776 ) | ( n4757 & n16776 ) ;
  assign n16778 = ~n16766 & n16777 ;
  assign n16779 = n14950 | n14953 ;
  assign n16780 = x142 & n16779 ;
  assign n16781 = ( x603 & n14922 ) | ( x603 & n14927 ) | ( n14922 & n14927 ) ;
  assign n16782 = x142 | n16781 ;
  assign n16783 = x743 & n16782 ;
  assign n16784 = ~n16780 & n16783 ;
  assign n16785 = x142 & ~x743 ;
  assign n16786 = ~n14820 & n16785 ;
  assign n16787 = x299 | n16786 ;
  assign n16788 = n16784 | n16787 ;
  assign n16789 = x142 & n14946 ;
  assign n16790 = x142 | n14920 ;
  assign n16791 = x142 & ~n14814 ;
  assign n16792 = ( x743 & n16790 ) | ( x743 & n16791 ) | ( n16790 & n16791 ) ;
  assign n16793 = ~n16789 & n16792 ;
  assign n16794 = x299 & ~n16793 ;
  assign n16795 = n16788 & ~n16794 ;
  assign n16796 = ( x38 & ~n9138 ) | ( x38 & n16795 ) | ( ~n9138 & n16795 ) ;
  assign n16797 = n16778 | n16796 ;
  assign n16798 = x39 & x142 ;
  assign n16799 = x38 & ~n16798 ;
  assign n16800 = x142 & ~n15756 ;
  assign n16801 = x743 & n14840 ;
  assign n16802 = ~n1868 & n16801 ;
  assign n16803 = n16800 | n16802 ;
  assign n16804 = ~x39 & n16803 ;
  assign n16805 = n16799 & ~n16804 ;
  assign n16806 = n2032 | n16805 ;
  assign n16807 = n16797 & ~n16806 ;
  assign n16808 = n16730 | n16807 ;
  assign n16809 = ~n15082 & n16808 ;
  assign n16810 = n15082 & n16727 ;
  assign n16811 = n16809 | n16810 ;
  assign n16812 = ~x785 & n16811 ;
  assign n16813 = ~n15088 & n16727 ;
  assign n16814 = x609 & n16809 ;
  assign n16815 = n16813 | n16814 ;
  assign n16816 = x1155 & n16815 ;
  assign n16817 = n15094 & n16727 ;
  assign n16818 = ~x609 & n16809 ;
  assign n16819 = n16817 | n16818 ;
  assign n16820 = ~x1155 & n16819 ;
  assign n16821 = n16816 | n16820 ;
  assign n16822 = x785 & n16821 ;
  assign n16823 = n16812 | n16822 ;
  assign n16824 = ~x781 & n16823 ;
  assign n16825 = ( x618 & x1154 ) | ( x618 & n16727 ) | ( x1154 & n16727 ) ;
  assign n16826 = ( ~x618 & x1154 ) | ( ~x618 & n16823 ) | ( x1154 & n16823 ) ;
  assign n16827 = n16825 & n16826 ;
  assign n16828 = ( x618 & x1154 ) | ( x618 & ~n16727 ) | ( x1154 & ~n16727 ) ;
  assign n16829 = ( x618 & ~x1154 ) | ( x618 & n16823 ) | ( ~x1154 & n16823 ) ;
  assign n16830 = ~n16828 & n16829 ;
  assign n16831 = n16827 | n16830 ;
  assign n16832 = x781 & n16831 ;
  assign n16833 = n16824 | n16832 ;
  assign n16834 = ~x789 & n16833 ;
  assign n16835 = ( x619 & x1159 ) | ( x619 & n16727 ) | ( x1159 & n16727 ) ;
  assign n16836 = ( ~x619 & x1159 ) | ( ~x619 & n16833 ) | ( x1159 & n16833 ) ;
  assign n16837 = n16835 & n16836 ;
  assign n16838 = ( x619 & x1159 ) | ( x619 & ~n16727 ) | ( x1159 & ~n16727 ) ;
  assign n16839 = ( x619 & ~x1159 ) | ( x619 & n16833 ) | ( ~x1159 & n16833 ) ;
  assign n16840 = ~n16838 & n16839 ;
  assign n16841 = n16837 | n16840 ;
  assign n16842 = x789 & n16841 ;
  assign n16843 = n16834 | n16842 ;
  assign n16844 = ( x626 & ~x1158 ) | ( x626 & n16843 ) | ( ~x1158 & n16843 ) ;
  assign n16845 = ~n16729 & n16844 ;
  assign n16846 = ( x626 & x1158 ) | ( x626 & n16727 ) | ( x1158 & n16727 ) ;
  assign n16847 = ( ~x626 & x1158 ) | ( ~x626 & n16843 ) | ( x1158 & n16843 ) ;
  assign n16848 = n16846 & n16847 ;
  assign n16849 = n16845 | n16848 ;
  assign n16850 = x788 & n16849 ;
  assign n16851 = ~x788 & n16843 ;
  assign n16852 = n16850 | n16851 ;
  assign n16853 = n15134 | n16852 ;
  assign n16854 = n15134 & ~n16727 ;
  assign n16855 = n16853 & ~n16854 ;
  assign n16856 = ~n15141 & n16855 ;
  assign n16857 = n16728 | n16856 ;
  assign n16858 = ( x644 & x715 ) | ( x644 & n16857 ) | ( x715 & n16857 ) ;
  assign n16859 = ( ~x644 & x715 ) | ( ~x644 & n16727 ) | ( x715 & n16727 ) ;
  assign n16860 = n16858 & n16859 ;
  assign n16861 = x1160 | n16860 ;
  assign n16862 = n15407 & n16727 ;
  assign n16863 = x735 | n16710 ;
  assign n16864 = n15285 & ~n15296 ;
  assign n16865 = ( ~x142 & x735 ) | ( ~x142 & n16864 ) | ( x735 & n16864 ) ;
  assign n16866 = ( n15175 & n15177 ) | ( n15175 & n15179 ) | ( n15177 & n15179 ) ;
  assign n16867 = ( x142 & x735 ) | ( x142 & ~n16866 ) | ( x735 & ~n16866 ) ;
  assign n16868 = n16865 & n16867 ;
  assign n16869 = n16863 & ~n16868 ;
  assign n16870 = ( ~n1823 & n4764 ) | ( ~n1823 & n16869 ) | ( n4764 & n16869 ) ;
  assign n16871 = x735 | n16713 ;
  assign n16872 = ( ~x142 & x735 ) | ( ~x142 & n15253 ) | ( x735 & n15253 ) ;
  assign n16873 = ( x142 & x735 ) | ( x142 & ~n15169 ) | ( x735 & ~n15169 ) ;
  assign n16874 = n16872 & n16873 ;
  assign n16875 = n16871 & ~n16874 ;
  assign n16876 = ( n1823 & n4764 ) | ( n1823 & ~n16875 ) | ( n4764 & ~n16875 ) ;
  assign n16877 = ~n16870 & n16876 ;
  assign n16878 = x735 & n15202 ;
  assign n16879 = ~n14481 & n16878 ;
  assign n16880 = n16706 | n16879 ;
  assign n16881 = ( ~x223 & n15629 ) | ( ~x223 & n16880 ) | ( n15629 & n16880 ) ;
  assign n16882 = ~n16877 & n16881 ;
  assign n16883 = x735 | n16717 ;
  assign n16884 = n15264 & ~n15272 ;
  assign n16885 = x142 & ~n16884 ;
  assign n16886 = ~x142 & n15846 ;
  assign n16887 = n15848 & n16886 ;
  assign n16888 = x735 & ~n16887 ;
  assign n16889 = ~n16885 & n16888 ;
  assign n16890 = n16883 & ~n16889 ;
  assign n16891 = ( x223 & ~n4764 ) | ( x223 & n16890 ) | ( ~n4764 & n16890 ) ;
  assign n16892 = x735 | n16720 ;
  assign n16893 = ~n15272 & n15275 ;
  assign n16894 = x142 & ~n16893 ;
  assign n16895 = x735 & ~n16886 ;
  assign n16896 = ~n16894 & n16895 ;
  assign n16897 = n16892 & ~n16896 ;
  assign n16898 = ( x223 & n4764 ) | ( x223 & n16897 ) | ( n4764 & n16897 ) ;
  assign n16899 = n16891 & n16898 ;
  assign n16900 = x299 | n16899 ;
  assign n16901 = n16882 | n16900 ;
  assign n16902 = n2203 | n16880 ;
  assign n16903 = ~x215 & n16902 ;
  assign n16904 = ( ~n2203 & n4721 ) | ( ~n2203 & n16869 ) | ( n4721 & n16869 ) ;
  assign n16905 = ( n2203 & n4721 ) | ( n2203 & ~n16875 ) | ( n4721 & ~n16875 ) ;
  assign n16906 = ~n16904 & n16905 ;
  assign n16907 = n16903 & ~n16906 ;
  assign n16908 = ( x215 & ~n4721 ) | ( x215 & n16890 ) | ( ~n4721 & n16890 ) ;
  assign n16909 = ( x215 & n4721 ) | ( x215 & n16897 ) | ( n4721 & n16897 ) ;
  assign n16910 = n16908 & n16909 ;
  assign n16911 = x299 & ~n16910 ;
  assign n16912 = ~n16907 & n16911 ;
  assign n16913 = x39 & ~n16912 ;
  assign n16914 = n16901 & n16913 ;
  assign n16915 = x142 & ~x735 ;
  assign n16916 = ~n14822 & n16915 ;
  assign n16917 = ( x142 & ~x735 ) | ( x142 & n15345 ) | ( ~x735 & n15345 ) ;
  assign n16918 = ( x142 & x735 ) | ( x142 & n15369 ) | ( x735 & n15369 ) ;
  assign n16919 = ~n16917 & n16918 ;
  assign n16920 = n16916 | n16919 ;
  assign n16921 = ~x39 & n16920 ;
  assign n16922 = x38 | n16921 ;
  assign n16923 = n16914 | n16922 ;
  assign n16924 = ~n1868 & n16878 ;
  assign n16925 = n16800 | n16924 ;
  assign n16926 = ~x39 & n16925 ;
  assign n16927 = n16799 & ~n16926 ;
  assign n16928 = n2032 | n16927 ;
  assign n16929 = n16923 & ~n16928 ;
  assign n16930 = n16730 | n16929 ;
  assign n16931 = ~x778 & n16930 ;
  assign n16932 = ( x625 & x1153 ) | ( x625 & ~n16727 ) | ( x1153 & ~n16727 ) ;
  assign n16933 = ( x625 & ~x1153 ) | ( x625 & n16930 ) | ( ~x1153 & n16930 ) ;
  assign n16934 = ~n16932 & n16933 ;
  assign n16935 = ( x625 & x1153 ) | ( x625 & n16727 ) | ( x1153 & n16727 ) ;
  assign n16936 = ( ~x625 & x1153 ) | ( ~x625 & n16930 ) | ( x1153 & n16930 ) ;
  assign n16937 = n16935 & n16936 ;
  assign n16938 = n16934 | n16937 ;
  assign n16939 = x778 & n16938 ;
  assign n16940 = n16931 | n16939 ;
  assign n16941 = n15400 | n16940 ;
  assign n16942 = n15400 & ~n16727 ;
  assign n16943 = n16941 & ~n16942 ;
  assign n16944 = ~n15407 & n16943 ;
  assign n16945 = n16862 | n16944 ;
  assign n16946 = n15414 | n16945 ;
  assign n16947 = n15414 & ~n16727 ;
  assign n16948 = n16946 & ~n16947 ;
  assign n16949 = n15421 | n16948 ;
  assign n16950 = n15421 & ~n16727 ;
  assign n16951 = n16949 & ~n16950 ;
  assign n16952 = ~x792 & n16951 ;
  assign n16953 = ( x628 & x1156 ) | ( x628 & n16727 ) | ( x1156 & n16727 ) ;
  assign n16954 = ( ~x628 & x1156 ) | ( ~x628 & n16951 ) | ( x1156 & n16951 ) ;
  assign n16955 = n16953 & n16954 ;
  assign n16956 = ( x628 & x1156 ) | ( x628 & ~n16727 ) | ( x1156 & ~n16727 ) ;
  assign n16957 = ( x628 & ~x1156 ) | ( x628 & n16951 ) | ( ~x1156 & n16951 ) ;
  assign n16958 = ~n16956 & n16957 ;
  assign n16959 = n16955 | n16958 ;
  assign n16960 = x792 & n16959 ;
  assign n16961 = n16952 | n16960 ;
  assign n16962 = ~x787 & n16961 ;
  assign n16963 = ( x647 & x1157 ) | ( x647 & n16727 ) | ( x1157 & n16727 ) ;
  assign n16964 = ( ~x647 & x1157 ) | ( ~x647 & n16961 ) | ( x1157 & n16961 ) ;
  assign n16965 = n16963 & n16964 ;
  assign n16966 = ( x647 & x1157 ) | ( x647 & ~n16727 ) | ( x1157 & ~n16727 ) ;
  assign n16967 = ( x647 & ~x1157 ) | ( x647 & n16961 ) | ( ~x1157 & n16961 ) ;
  assign n16968 = ~n16966 & n16967 ;
  assign n16969 = n16965 | n16968 ;
  assign n16970 = x787 & n16969 ;
  assign n16971 = n16962 | n16970 ;
  assign n16972 = ( x644 & x715 ) | ( x644 & ~n16971 ) | ( x715 & ~n16971 ) ;
  assign n16973 = x630 | n16965 ;
  assign n16974 = ( x647 & x1157 ) | ( x647 & ~n16855 ) | ( x1157 & ~n16855 ) ;
  assign n16975 = x629 | n16955 ;
  assign n16976 = ( x628 & x1156 ) | ( x628 & ~n16852 ) | ( x1156 & ~n16852 ) ;
  assign n16977 = x648 | n16837 ;
  assign n16978 = ( x619 & x1159 ) | ( x619 & ~n16945 ) | ( x1159 & ~n16945 ) ;
  assign n16979 = x627 | n16827 ;
  assign n16980 = ( x618 & x1154 ) | ( x618 & ~n16943 ) | ( x1154 & ~n16943 ) ;
  assign n16981 = x660 | n16816 ;
  assign n16982 = ( x609 & x1155 ) | ( x609 & ~n16940 ) | ( x1155 & ~n16940 ) ;
  assign n16983 = x608 & ~n16934 ;
  assign n16984 = ( x625 & x1153 ) | ( x625 & n16808 ) | ( x1153 & n16808 ) ;
  assign n16985 = n15336 & n16780 ;
  assign n16986 = x680 & n15356 ;
  assign n16987 = n16782 | n16986 ;
  assign n16988 = ~n16985 & n16987 ;
  assign n16989 = x743 & ~n16988 ;
  assign n16990 = x680 & n15881 ;
  assign n16991 = ~x142 & n16990 ;
  assign n16992 = x142 & ~n15336 ;
  assign n16993 = ~n16781 & n16992 ;
  assign n16994 = x743 | n16993 ;
  assign n16995 = n16991 | n16994 ;
  assign n16996 = ~x299 & n16995 ;
  assign n16997 = ~n16989 & n16996 ;
  assign n16998 = x680 & n15885 ;
  assign n16999 = ~x142 & n16998 ;
  assign n17000 = x142 & ~n15343 ;
  assign n17001 = ~n14920 & n17000 ;
  assign n17002 = x743 | n17001 ;
  assign n17003 = n16999 | n17002 ;
  assign n17004 = x680 & n15366 ;
  assign n17005 = n16790 | n17004 ;
  assign n17006 = ~n15342 & n16789 ;
  assign n17007 = n17005 & ~n17006 ;
  assign n17008 = x743 & ~n17007 ;
  assign n17009 = x299 & ~n17008 ;
  assign n17010 = n17003 & n17009 ;
  assign n17011 = n16997 | n17010 ;
  assign n17012 = ( x39 & x735 ) | ( x39 & n17011 ) | ( x735 & n17011 ) ;
  assign n17013 = ( x39 & ~x735 ) | ( x39 & n16795 ) | ( ~x735 & n16795 ) ;
  assign n17014 = n17012 | n17013 ;
  assign n17015 = n15913 | n16803 ;
  assign n17016 = ~n14479 & n17015 ;
  assign n17017 = ( x735 & n16706 ) | ( x735 & n17016 ) | ( n16706 & n17016 ) ;
  assign n17018 = ( ~x735 & n16706 ) | ( ~x735 & n16731 ) | ( n16706 & n16731 ) ;
  assign n17019 = n17017 | n17018 ;
  assign n17020 = n2203 | n17019 ;
  assign n17021 = ~x215 & n17020 ;
  assign n17022 = ( n15726 & n15734 ) | ( n15726 & ~n15736 ) | ( n15734 & ~n15736 ) ;
  assign n17023 = ( x142 & ~x743 ) | ( x142 & n17022 ) | ( ~x743 & n17022 ) ;
  assign n17024 = ~n15825 & n15829 ;
  assign n17025 = ( x142 & x743 ) | ( x142 & n17024 ) | ( x743 & n17024 ) ;
  assign n17026 = ~n17023 & n17025 ;
  assign n17027 = ( x142 & ~x743 ) | ( x142 & n15528 ) | ( ~x743 & n15528 ) ;
  assign n17028 = ( x142 & x743 ) | ( x142 & n15598 ) | ( x743 & n15598 ) ;
  assign n17029 = n17027 & ~n17028 ;
  assign n17030 = n17026 | n17029 ;
  assign n17031 = x735 & n17030 ;
  assign n17032 = ~x735 & n16740 ;
  assign n17033 = n17031 | n17032 ;
  assign n17034 = ( ~n2203 & n4721 ) | ( ~n2203 & n17033 ) | ( n4721 & n17033 ) ;
  assign n17035 = n15712 & ~n15721 ;
  assign n17036 = ( x142 & ~x743 ) | ( x142 & n17035 ) | ( ~x743 & n17035 ) ;
  assign n17037 = ( x142 & x743 ) | ( x142 & n15813 ) | ( x743 & n15813 ) ;
  assign n17038 = ~n17036 & n17037 ;
  assign n17039 = ( x142 & ~x743 ) | ( x142 & n15559 ) | ( ~x743 & n15559 ) ;
  assign n17040 = ( x142 & x743 ) | ( x142 & n15626 ) | ( x743 & n15626 ) ;
  assign n17041 = n17039 & ~n17040 ;
  assign n17042 = n17038 | n17041 ;
  assign n17043 = x735 & n17042 ;
  assign n17044 = ~x735 & n16747 ;
  assign n17045 = n17043 | n17044 ;
  assign n17046 = ( n2203 & n4721 ) | ( n2203 & ~n17045 ) | ( n4721 & ~n17045 ) ;
  assign n17047 = ~n17034 & n17046 ;
  assign n17048 = n17021 & ~n17047 ;
  assign n17049 = n15750 & ~n15752 ;
  assign n17050 = ( x142 & ~x743 ) | ( x142 & n17049 ) | ( ~x743 & n17049 ) ;
  assign n17051 = ( x142 & x743 ) | ( x142 & n15850 ) | ( x743 & n15850 ) ;
  assign n17052 = ~n17050 & n17051 ;
  assign n17053 = ( n15475 & ~n15482 ) | ( n15475 & n15484 ) | ( ~n15482 & n15484 ) ;
  assign n17054 = ( x142 & ~x743 ) | ( x142 & n17053 ) | ( ~x743 & n17053 ) ;
  assign n17055 = ~n15652 & n15655 ;
  assign n17056 = ( x142 & x743 ) | ( x142 & n17055 ) | ( x743 & n17055 ) ;
  assign n17057 = n17054 & ~n17056 ;
  assign n17058 = n17052 | n17057 ;
  assign n17059 = x735 & n17058 ;
  assign n17060 = ~x735 & n16755 ;
  assign n17061 = n17059 | n17060 ;
  assign n17062 = ( x215 & ~n4721 ) | ( x215 & n17061 ) | ( ~n4721 & n17061 ) ;
  assign n17063 = ( n14989 & n15766 ) | ( n14989 & ~n15767 ) | ( n15766 & ~n15767 ) ;
  assign n17064 = ( x142 & ~x743 ) | ( x142 & n17063 ) | ( ~x743 & n17063 ) ;
  assign n17065 = ( x142 & x743 ) | ( x142 & n15843 ) | ( x743 & n15843 ) ;
  assign n17066 = ~n17064 & n17065 ;
  assign n17067 = ( x142 & ~x743 ) | ( x142 & n15498 ) | ( ~x743 & n15498 ) ;
  assign n17068 = ( x142 & x743 ) | ( x142 & n15677 ) | ( x743 & n15677 ) ;
  assign n17069 = n17067 & ~n17068 ;
  assign n17070 = n17066 | n17069 ;
  assign n17071 = x735 & n17070 ;
  assign n17072 = ~x735 & n16762 ;
  assign n17073 = n17071 | n17072 ;
  assign n17074 = ( x215 & n4721 ) | ( x215 & n17073 ) | ( n4721 & n17073 ) ;
  assign n17075 = n17062 & n17074 ;
  assign n17076 = n17048 | n17075 ;
  assign n17077 = ( ~x39 & x299 ) | ( ~x39 & n17076 ) | ( x299 & n17076 ) ;
  assign n17078 = n1823 | n17019 ;
  assign n17079 = ~x223 & n17078 ;
  assign n17080 = ( ~n1823 & n4764 ) | ( ~n1823 & n17033 ) | ( n4764 & n17033 ) ;
  assign n17081 = ( n1823 & n4764 ) | ( n1823 & ~n17045 ) | ( n4764 & ~n17045 ) ;
  assign n17082 = ~n17080 & n17081 ;
  assign n17083 = n17079 & ~n17082 ;
  assign n17084 = ( x223 & ~n4764 ) | ( x223 & n17061 ) | ( ~n4764 & n17061 ) ;
  assign n17085 = ( x223 & n4764 ) | ( x223 & n17073 ) | ( n4764 & n17073 ) ;
  assign n17086 = n17084 & n17085 ;
  assign n17087 = n17083 | n17086 ;
  assign n17088 = ( x39 & x299 ) | ( x39 & ~n17087 ) | ( x299 & ~n17087 ) ;
  assign n17089 = ~n17077 & n17088 ;
  assign n17090 = n17014 & ~n17089 ;
  assign n17091 = x38 | n17090 ;
  assign n17092 = x735 & n15913 ;
  assign n17093 = n16803 | n17092 ;
  assign n17094 = ~x39 & n17093 ;
  assign n17095 = n16799 & ~n17094 ;
  assign n17096 = n2032 | n17095 ;
  assign n17097 = n17091 & ~n17096 ;
  assign n17098 = n16730 | n17097 ;
  assign n17099 = ( ~x625 & x1153 ) | ( ~x625 & n17098 ) | ( x1153 & n17098 ) ;
  assign n17100 = n16984 & n17099 ;
  assign n17101 = n16983 & ~n17100 ;
  assign n17102 = x608 | n16937 ;
  assign n17103 = ( x625 & x1153 ) | ( x625 & ~n16808 ) | ( x1153 & ~n16808 ) ;
  assign n17104 = ( x625 & ~x1153 ) | ( x625 & n17098 ) | ( ~x1153 & n17098 ) ;
  assign n17105 = ~n17103 & n17104 ;
  assign n17106 = n17102 | n17105 ;
  assign n17107 = ~n17101 & n17106 ;
  assign n17108 = x778 & ~n17107 ;
  assign n17109 = x778 | n17098 ;
  assign n17110 = ~n17108 & n17109 ;
  assign n17111 = ( x609 & ~x1155 ) | ( x609 & n17110 ) | ( ~x1155 & n17110 ) ;
  assign n17112 = ~n16982 & n17111 ;
  assign n17113 = n16981 | n17112 ;
  assign n17114 = x660 & ~n16820 ;
  assign n17115 = ( x609 & x1155 ) | ( x609 & n16940 ) | ( x1155 & n16940 ) ;
  assign n17116 = ( ~x609 & x1155 ) | ( ~x609 & n17110 ) | ( x1155 & n17110 ) ;
  assign n17117 = n17115 & n17116 ;
  assign n17118 = n17114 & ~n17117 ;
  assign n17119 = n17113 & ~n17118 ;
  assign n17120 = x785 & ~n17119 ;
  assign n17121 = x785 | n17110 ;
  assign n17122 = ~n17120 & n17121 ;
  assign n17123 = ( x618 & ~x1154 ) | ( x618 & n17122 ) | ( ~x1154 & n17122 ) ;
  assign n17124 = ~n16980 & n17123 ;
  assign n17125 = n16979 | n17124 ;
  assign n17126 = x627 & ~n16830 ;
  assign n17127 = ( x618 & x1154 ) | ( x618 & n16943 ) | ( x1154 & n16943 ) ;
  assign n17128 = ( ~x618 & x1154 ) | ( ~x618 & n17122 ) | ( x1154 & n17122 ) ;
  assign n17129 = n17127 & n17128 ;
  assign n17130 = n17126 & ~n17129 ;
  assign n17131 = n17125 & ~n17130 ;
  assign n17132 = x781 & ~n17131 ;
  assign n17133 = x781 | n17122 ;
  assign n17134 = ~n17132 & n17133 ;
  assign n17135 = ( x619 & ~x1159 ) | ( x619 & n17134 ) | ( ~x1159 & n17134 ) ;
  assign n17136 = ~n16978 & n17135 ;
  assign n17137 = n16977 | n17136 ;
  assign n17138 = x648 & ~n16840 ;
  assign n17139 = ( x619 & x1159 ) | ( x619 & n16945 ) | ( x1159 & n16945 ) ;
  assign n17140 = ( ~x619 & x1159 ) | ( ~x619 & n17134 ) | ( x1159 & n17134 ) ;
  assign n17141 = n17139 & n17140 ;
  assign n17142 = n17138 & ~n17141 ;
  assign n17143 = n17137 & ~n17142 ;
  assign n17144 = x789 & ~n17143 ;
  assign n17145 = x789 | n17134 ;
  assign n17146 = ~n17144 & n17145 ;
  assign n17147 = ~x788 & n17146 ;
  assign n17148 = n15972 & ~n16845 ;
  assign n17149 = ( x626 & x641 ) | ( x626 & n16948 ) | ( x641 & n16948 ) ;
  assign n17150 = ( ~x626 & x641 ) | ( ~x626 & n17146 ) | ( x641 & n17146 ) ;
  assign n17151 = n17149 | n17150 ;
  assign n17152 = ~n17148 & n17151 ;
  assign n17153 = n15978 | n16848 ;
  assign n17154 = ( x626 & x641 ) | ( x626 & ~n16948 ) | ( x641 & ~n16948 ) ;
  assign n17155 = ( x626 & ~x641 ) | ( x626 & n17146 ) | ( ~x641 & n17146 ) ;
  assign n17156 = n17154 & ~n17155 ;
  assign n17157 = n17153 & ~n17156 ;
  assign n17158 = n17152 | n17157 ;
  assign n17159 = x788 & n17158 ;
  assign n17160 = n17147 | n17159 ;
  assign n17161 = ( x628 & ~x1156 ) | ( x628 & n17160 ) | ( ~x1156 & n17160 ) ;
  assign n17162 = ~n16976 & n17161 ;
  assign n17163 = n16975 | n17162 ;
  assign n17164 = x629 & ~n16958 ;
  assign n17165 = ( x628 & x1156 ) | ( x628 & n16852 ) | ( x1156 & n16852 ) ;
  assign n17166 = ( ~x628 & x1156 ) | ( ~x628 & n17160 ) | ( x1156 & n17160 ) ;
  assign n17167 = n17165 & n17166 ;
  assign n17168 = n17164 & ~n17167 ;
  assign n17169 = n17163 & ~n17168 ;
  assign n17170 = x792 & ~n17169 ;
  assign n17171 = x792 | n17160 ;
  assign n17172 = ~n17170 & n17171 ;
  assign n17173 = ( x647 & ~x1157 ) | ( x647 & n17172 ) | ( ~x1157 & n17172 ) ;
  assign n17174 = ~n16974 & n17173 ;
  assign n17175 = n16973 | n17174 ;
  assign n17176 = x630 & ~n16968 ;
  assign n17177 = ( x647 & x1157 ) | ( x647 & n16855 ) | ( x1157 & n16855 ) ;
  assign n17178 = ( ~x647 & x1157 ) | ( ~x647 & n17172 ) | ( x1157 & n17172 ) ;
  assign n17179 = n17177 & n17178 ;
  assign n17180 = n17176 & ~n17179 ;
  assign n17181 = n17175 & ~n17180 ;
  assign n17182 = x787 & ~n17181 ;
  assign n17183 = x787 | n17172 ;
  assign n17184 = ~n17182 & n17183 ;
  assign n17185 = ( x644 & ~x715 ) | ( x644 & n17184 ) | ( ~x715 & n17184 ) ;
  assign n17186 = ~n16972 & n17185 ;
  assign n17187 = n16861 | n17186 ;
  assign n17188 = ( x644 & x715 ) | ( x644 & ~n16857 ) | ( x715 & ~n16857 ) ;
  assign n17189 = ( x644 & ~x715 ) | ( x644 & n16727 ) | ( ~x715 & n16727 ) ;
  assign n17190 = ~n17188 & n17189 ;
  assign n17191 = x1160 & ~n17190 ;
  assign n17192 = ( x644 & x715 ) | ( x644 & n16971 ) | ( x715 & n16971 ) ;
  assign n17193 = ( ~x644 & x715 ) | ( ~x644 & n17184 ) | ( x715 & n17184 ) ;
  assign n17194 = n17192 & n17193 ;
  assign n17195 = n17191 & ~n17194 ;
  assign n17196 = x790 & ~n17195 ;
  assign n17197 = n17187 & n17196 ;
  assign n17198 = ~x790 & n17184 ;
  assign n17199 = n4832 | n17198 ;
  assign n17200 = n17197 | n17199 ;
  assign n17201 = ~x142 & n4832 ;
  assign n17202 = x57 | n17201 ;
  assign n17203 = n17200 & ~n17202 ;
  assign n17204 = x57 & x142 ;
  assign n17205 = x832 | n17204 ;
  assign n17206 = n17203 | n17205 ;
  assign n17207 = x142 & ~n1290 ;
  assign n17208 = ~x625 & x1153 ;
  assign n17209 = ( x778 & ~x1153 ) | ( x778 & n17208 ) | ( ~x1153 & n17208 ) ;
  assign n17210 = ( x625 & n17208 ) | ( x625 & n17209 ) | ( n17208 & n17209 ) ;
  assign n17211 = n16878 & ~n17210 ;
  assign n17212 = n17207 | n17211 ;
  assign n17213 = n15414 | n15421 ;
  assign n17214 = n15400 | n15407 ;
  assign n17215 = n17213 | n17214 ;
  assign n17216 = n17212 & ~n17215 ;
  assign n17217 = x628 | x1156 ;
  assign n17218 = x628 & x1156 ;
  assign n17219 = x792 & ~n17218 ;
  assign n17220 = n17217 & n17219 ;
  assign n17221 = n17216 & ~n17220 ;
  assign n17222 = x647 & n17221 ;
  assign n17223 = x1157 & ~n17207 ;
  assign n17224 = ~n17222 & n17223 ;
  assign n17225 = x630 | n17224 ;
  assign n17226 = ~n15082 & n16801 ;
  assign n17227 = x609 & n17226 ;
  assign n17228 = x1155 & ~n17207 ;
  assign n17229 = ~n17227 & n17228 ;
  assign n17230 = ~x609 & n17226 ;
  assign n17231 = x1155 | n17207 ;
  assign n17232 = n17230 | n17231 ;
  assign n17233 = ~n17229 & n17232 ;
  assign n17234 = x785 & ~n17233 ;
  assign n17235 = x785 | n17207 ;
  assign n17236 = n17226 | n17235 ;
  assign n17237 = ~n17234 & n17236 ;
  assign n17238 = x781 | n17237 ;
  assign n17239 = ( x618 & x1154 ) | ( x618 & ~n17207 ) | ( x1154 & ~n17207 ) ;
  assign n17240 = ( x618 & ~x1154 ) | ( x618 & n17237 ) | ( ~x1154 & n17237 ) ;
  assign n17241 = n17239 & ~n17240 ;
  assign n17242 = ( x618 & x1154 ) | ( x618 & n17207 ) | ( x1154 & n17207 ) ;
  assign n17243 = ( ~x618 & x1154 ) | ( ~x618 & n17237 ) | ( x1154 & n17237 ) ;
  assign n17244 = n17242 | n17243 ;
  assign n17245 = ~n17241 & n17244 ;
  assign n17246 = x781 & ~n17245 ;
  assign n17247 = n17238 & ~n17246 ;
  assign n17248 = x789 | n17247 ;
  assign n17249 = ( x619 & x1159 ) | ( x619 & ~n17207 ) | ( x1159 & ~n17207 ) ;
  assign n17250 = ( x619 & ~x1159 ) | ( x619 & n17247 ) | ( ~x1159 & n17247 ) ;
  assign n17251 = n17249 & ~n17250 ;
  assign n17252 = ( x619 & x1159 ) | ( x619 & n17207 ) | ( x1159 & n17207 ) ;
  assign n17253 = ( ~x619 & x1159 ) | ( ~x619 & n17247 ) | ( x1159 & n17247 ) ;
  assign n17254 = n17252 | n17253 ;
  assign n17255 = ~n17251 & n17254 ;
  assign n17256 = x789 & ~n17255 ;
  assign n17257 = n17248 & ~n17256 ;
  assign n17258 = x788 | n17257 ;
  assign n17259 = ( x626 & x1158 ) | ( x626 & n17207 ) | ( x1158 & n17207 ) ;
  assign n17260 = ( ~x1158 & n17257 ) | ( ~x1158 & n17259 ) | ( n17257 & n17259 ) ;
  assign n17261 = ( ~x626 & n17259 ) | ( ~x626 & n17260 ) | ( n17259 & n17260 ) ;
  assign n17262 = x788 & ~n17261 ;
  assign n17263 = n17258 & ~n17262 ;
  assign n17264 = ~n15134 & n17263 ;
  assign n17265 = n15134 & n17207 ;
  assign n17266 = n17264 | n17265 ;
  assign n17267 = ( x647 & x1157 ) | ( x647 & n17266 ) | ( x1157 & n17266 ) ;
  assign n17268 = x628 & n17216 ;
  assign n17269 = n17207 | n17268 ;
  assign n17270 = x1156 & n17269 ;
  assign n17271 = x629 | n17270 ;
  assign n17272 = ( x628 & x1156 ) | ( x628 & ~n17263 ) | ( x1156 & ~n17263 ) ;
  assign n17273 = n15420 & n17261 ;
  assign n17274 = n15414 & ~n17207 ;
  assign n17275 = n16115 & ~n17274 ;
  assign n17276 = ( n17207 & n17212 ) | ( n17207 & ~n17214 ) | ( n17212 & ~n17214 ) ;
  assign n17277 = n17275 & n17276 ;
  assign n17278 = n17273 | n17277 ;
  assign n17279 = x788 & n17278 ;
  assign n17280 = x648 & n17254 ;
  assign n17281 = ( x619 & x1159 ) | ( x619 & ~n17276 ) | ( x1159 & ~n17276 ) ;
  assign n17282 = x627 | n17241 ;
  assign n17283 = ~n15400 & n17212 ;
  assign n17284 = n17207 | n17283 ;
  assign n17285 = ( x618 & x1154 ) | ( x618 & n17284 ) | ( x1154 & n17284 ) ;
  assign n17286 = x660 | n17229 ;
  assign n17287 = ( x609 & x1155 ) | ( x609 & n17212 ) | ( x1155 & n17212 ) ;
  assign n17288 = x735 & n15529 ;
  assign n17289 = x625 & n17288 ;
  assign n17290 = n16801 | n17207 ;
  assign n17291 = n17288 | n17290 ;
  assign n17292 = ~n17289 & n17291 ;
  assign n17293 = x1153 | n17292 ;
  assign n17294 = x625 & n16878 ;
  assign n17295 = x1153 & ~n17207 ;
  assign n17296 = ~n17294 & n17295 ;
  assign n17297 = x608 | n17296 ;
  assign n17298 = n17293 & ~n17297 ;
  assign n17299 = n16801 | n17289 ;
  assign n17300 = x1153 & n17299 ;
  assign n17301 = x625 | x1153 ;
  assign n17302 = n16878 & ~n17301 ;
  assign n17303 = n17207 | n17302 ;
  assign n17304 = n17300 | n17303 ;
  assign n17305 = x608 & n17304 ;
  assign n17306 = n17298 | n17305 ;
  assign n17307 = x778 & n17306 ;
  assign n17308 = ~x778 & n17291 ;
  assign n17309 = n17307 | n17308 ;
  assign n17310 = ( ~x609 & x1155 ) | ( ~x609 & n17309 ) | ( x1155 & n17309 ) ;
  assign n17311 = n17287 | n17310 ;
  assign n17312 = ~n17286 & n17311 ;
  assign n17313 = x660 & n17232 ;
  assign n17314 = ( x609 & x1155 ) | ( x609 & ~n17212 ) | ( x1155 & ~n17212 ) ;
  assign n17315 = ( x609 & ~x1155 ) | ( x609 & n17309 ) | ( ~x1155 & n17309 ) ;
  assign n17316 = n17314 & ~n17315 ;
  assign n17317 = n17313 & ~n17316 ;
  assign n17318 = n17312 | n17317 ;
  assign n17319 = x785 & n17318 ;
  assign n17320 = ~x785 & n17309 ;
  assign n17321 = n17319 | n17320 ;
  assign n17322 = ( ~x618 & x1154 ) | ( ~x618 & n17321 ) | ( x1154 & n17321 ) ;
  assign n17323 = n17285 | n17322 ;
  assign n17324 = ~n17282 & n17323 ;
  assign n17325 = x627 & n17244 ;
  assign n17326 = ( x618 & x1154 ) | ( x618 & ~n17284 ) | ( x1154 & ~n17284 ) ;
  assign n17327 = ( x618 & ~x1154 ) | ( x618 & n17321 ) | ( ~x1154 & n17321 ) ;
  assign n17328 = n17326 & ~n17327 ;
  assign n17329 = n17325 & ~n17328 ;
  assign n17330 = n17324 | n17329 ;
  assign n17331 = x781 & n17330 ;
  assign n17332 = ~x781 & n17321 ;
  assign n17333 = n17331 | n17332 ;
  assign n17334 = ( x619 & ~x1159 ) | ( x619 & n17333 ) | ( ~x1159 & n17333 ) ;
  assign n17335 = n17281 & ~n17334 ;
  assign n17336 = n17280 & ~n17335 ;
  assign n17337 = x648 | n17251 ;
  assign n17338 = ( x619 & x1159 ) | ( x619 & n17276 ) | ( x1159 & n17276 ) ;
  assign n17339 = ( ~x619 & x1159 ) | ( ~x619 & n17333 ) | ( x1159 & n17333 ) ;
  assign n17340 = n17338 | n17339 ;
  assign n17341 = ~n17337 & n17340 ;
  assign n17342 = x789 & ~n17341 ;
  assign n17343 = ~n17336 & n17342 ;
  assign n17344 = x789 | n17333 ;
  assign n17345 = ~n16177 & n17344 ;
  assign n17346 = ~n17343 & n17345 ;
  assign n17347 = n17279 | n17346 ;
  assign n17348 = ( x628 & ~x1156 ) | ( x628 & n17347 ) | ( ~x1156 & n17347 ) ;
  assign n17349 = ~n17272 & n17348 ;
  assign n17350 = n17271 | n17349 ;
  assign n17351 = ~x628 & n17216 ;
  assign n17352 = n17207 | n17351 ;
  assign n17353 = ~x1156 & n17352 ;
  assign n17354 = x629 & ~n17353 ;
  assign n17355 = ( x628 & x1156 ) | ( x628 & n17263 ) | ( x1156 & n17263 ) ;
  assign n17356 = ( ~x628 & x1156 ) | ( ~x628 & n17347 ) | ( x1156 & n17347 ) ;
  assign n17357 = n17355 & n17356 ;
  assign n17358 = n17354 & ~n17357 ;
  assign n17359 = n17350 & ~n17358 ;
  assign n17360 = x792 & ~n17359 ;
  assign n17361 = x792 | n17347 ;
  assign n17362 = ~n17360 & n17361 ;
  assign n17363 = ( ~x647 & x1157 ) | ( ~x647 & n17362 ) | ( x1157 & n17362 ) ;
  assign n17364 = n17267 | n17363 ;
  assign n17365 = ~n17225 & n17364 ;
  assign n17366 = ~x647 & n17221 ;
  assign n17367 = x1157 | n17207 ;
  assign n17368 = n17366 | n17367 ;
  assign n17369 = x630 & n17368 ;
  assign n17370 = ( x647 & x1157 ) | ( x647 & ~n17266 ) | ( x1157 & ~n17266 ) ;
  assign n17371 = ( x647 & ~x1157 ) | ( x647 & n17362 ) | ( ~x1157 & n17362 ) ;
  assign n17372 = n17370 & ~n17371 ;
  assign n17373 = n17369 & ~n17372 ;
  assign n17374 = n17365 | n17373 ;
  assign n17375 = x787 & n17374 ;
  assign n17376 = ~x787 & n17362 ;
  assign n17377 = n17375 | n17376 ;
  assign n17378 = ( x790 & x832 ) | ( x790 & ~n17377 ) | ( x832 & ~n17377 ) ;
  assign n17379 = n15141 & ~n17207 ;
  assign n17380 = n15141 | n17266 ;
  assign n17381 = ~n17379 & n17380 ;
  assign n17382 = ( x644 & x715 ) | ( x644 & n17381 ) | ( x715 & n17381 ) ;
  assign n17383 = ( ~x644 & x715 ) | ( ~x644 & n17207 ) | ( x715 & n17207 ) ;
  assign n17384 = n17382 | n17383 ;
  assign n17385 = x1160 & n17384 ;
  assign n17386 = ~x647 & x1157 ;
  assign n17387 = x647 & ~x1157 ;
  assign n17388 = n17386 | n17387 ;
  assign n17389 = x787 & n17388 ;
  assign n17390 = n17221 & ~n17389 ;
  assign n17391 = n17207 | n17390 ;
  assign n17392 = ( x644 & x715 ) | ( x644 & ~n17391 ) | ( x715 & ~n17391 ) ;
  assign n17393 = ( x644 & ~x715 ) | ( x644 & n17377 ) | ( ~x715 & n17377 ) ;
  assign n17394 = n17392 & ~n17393 ;
  assign n17395 = n17385 & ~n17394 ;
  assign n17396 = ( x644 & x715 ) | ( x644 & ~n17381 ) | ( x715 & ~n17381 ) ;
  assign n17397 = ( x644 & ~x715 ) | ( x644 & n17207 ) | ( ~x715 & n17207 ) ;
  assign n17398 = n17396 & ~n17397 ;
  assign n17399 = x1160 | n17398 ;
  assign n17400 = ( x644 & x715 ) | ( x644 & n17391 ) | ( x715 & n17391 ) ;
  assign n17401 = ( ~x644 & x715 ) | ( ~x644 & n17377 ) | ( x715 & n17377 ) ;
  assign n17402 = n17400 | n17401 ;
  assign n17403 = ~n17399 & n17402 ;
  assign n17404 = n17395 | n17403 ;
  assign n17405 = ( x790 & ~x832 ) | ( x790 & n17404 ) | ( ~x832 & n17404 ) ;
  assign n17406 = n17378 & ~n17405 ;
  assign n17407 = n17206 & ~n17406 ;
  assign n17408 = x143 | n14834 ;
  assign n17409 = n15141 & n17408 ;
  assign n17410 = ( x626 & x1158 ) | ( x626 & ~n17408 ) | ( x1158 & ~n17408 ) ;
  assign n17411 = x143 & n2032 ;
  assign n17412 = x143 | n15382 ;
  assign n17413 = x774 & n17412 ;
  assign n17414 = ~n4660 & n14840 ;
  assign n17415 = x38 & n17414 ;
  assign n17416 = ~x38 & n14933 ;
  assign n17417 = x143 & ~n17416 ;
  assign n17418 = x38 | n15063 ;
  assign n17419 = ~n4810 & n14959 ;
  assign n17420 = x38 & ~n17419 ;
  assign n17421 = n17418 & ~n17420 ;
  assign n17422 = x143 | x774 ;
  assign n17423 = n17421 & ~n17422 ;
  assign n17424 = n17417 | n17423 ;
  assign n17425 = ~n17415 & n17424 ;
  assign n17426 = n17413 | n17425 ;
  assign n17427 = ~n2032 & n17426 ;
  assign n17428 = n17411 | n17427 ;
  assign n17429 = ~n15082 & n17428 ;
  assign n17430 = n15082 & n17408 ;
  assign n17431 = n17429 | n17430 ;
  assign n17432 = ~x785 & n17431 ;
  assign n17433 = ~n15088 & n17408 ;
  assign n17434 = x609 & n17429 ;
  assign n17435 = n17433 | n17434 ;
  assign n17436 = x1155 & n17435 ;
  assign n17437 = n15094 & n17408 ;
  assign n17438 = ~x609 & n17429 ;
  assign n17439 = n17437 | n17438 ;
  assign n17440 = ~x1155 & n17439 ;
  assign n17441 = n17436 | n17440 ;
  assign n17442 = x785 & n17441 ;
  assign n17443 = n17432 | n17442 ;
  assign n17444 = ~x781 & n17443 ;
  assign n17445 = ( x618 & x1154 ) | ( x618 & n17408 ) | ( x1154 & n17408 ) ;
  assign n17446 = ( ~x618 & x1154 ) | ( ~x618 & n17443 ) | ( x1154 & n17443 ) ;
  assign n17447 = n17445 & n17446 ;
  assign n17448 = ( x618 & x1154 ) | ( x618 & ~n17408 ) | ( x1154 & ~n17408 ) ;
  assign n17449 = ( x618 & ~x1154 ) | ( x618 & n17443 ) | ( ~x1154 & n17443 ) ;
  assign n17450 = ~n17448 & n17449 ;
  assign n17451 = n17447 | n17450 ;
  assign n17452 = x781 & n17451 ;
  assign n17453 = n17444 | n17452 ;
  assign n17454 = ~x789 & n17453 ;
  assign n17455 = ( x619 & x1159 ) | ( x619 & n17408 ) | ( x1159 & n17408 ) ;
  assign n17456 = ( ~x619 & x1159 ) | ( ~x619 & n17453 ) | ( x1159 & n17453 ) ;
  assign n17457 = n17455 & n17456 ;
  assign n17458 = ( x619 & x1159 ) | ( x619 & ~n17408 ) | ( x1159 & ~n17408 ) ;
  assign n17459 = ( x619 & ~x1159 ) | ( x619 & n17453 ) | ( ~x1159 & n17453 ) ;
  assign n17460 = ~n17458 & n17459 ;
  assign n17461 = n17457 | n17460 ;
  assign n17462 = x789 & n17461 ;
  assign n17463 = n17454 | n17462 ;
  assign n17464 = ( x626 & ~x1158 ) | ( x626 & n17463 ) | ( ~x1158 & n17463 ) ;
  assign n17465 = ~n17410 & n17464 ;
  assign n17466 = ( x626 & x1158 ) | ( x626 & n17408 ) | ( x1158 & n17408 ) ;
  assign n17467 = ( ~x626 & x1158 ) | ( ~x626 & n17463 ) | ( x1158 & n17463 ) ;
  assign n17468 = n17466 & n17467 ;
  assign n17469 = n17465 | n17468 ;
  assign n17470 = x788 & n17469 ;
  assign n17471 = ~x788 & n17463 ;
  assign n17472 = n17470 | n17471 ;
  assign n17473 = n15134 | n17472 ;
  assign n17474 = n15134 & ~n17408 ;
  assign n17475 = n17473 & ~n17474 ;
  assign n17476 = ~n15141 & n17475 ;
  assign n17477 = n17409 | n17476 ;
  assign n17478 = ( x644 & x715 ) | ( x644 & n17477 ) | ( x715 & n17477 ) ;
  assign n17479 = ( ~x644 & x715 ) | ( ~x644 & n17408 ) | ( x715 & n17408 ) ;
  assign n17480 = n17478 & n17479 ;
  assign n17481 = x1160 | n17480 ;
  assign n17482 = n15414 & n17408 ;
  assign n17483 = x143 | n15070 ;
  assign n17484 = n15375 & n17483 ;
  assign n17485 = x687 & ~n17484 ;
  assign n17486 = ( ~x38 & x143 ) | ( ~x38 & n16319 ) | ( x143 & n16319 ) ;
  assign n17487 = ( x38 & x143 ) | ( x38 & n16323 ) | ( x143 & n16323 ) ;
  assign n17488 = n17486 & ~n17487 ;
  assign n17489 = n17485 & ~n17488 ;
  assign n17490 = x687 | n17412 ;
  assign n17491 = ~n2032 & n17490 ;
  assign n17492 = ~n17489 & n17491 ;
  assign n17493 = n17411 | n17492 ;
  assign n17494 = ~x778 & n17493 ;
  assign n17495 = ( x625 & x1153 ) | ( x625 & n17408 ) | ( x1153 & n17408 ) ;
  assign n17496 = ( ~x625 & x1153 ) | ( ~x625 & n17493 ) | ( x1153 & n17493 ) ;
  assign n17497 = n17495 & n17496 ;
  assign n17498 = ( x625 & x1153 ) | ( x625 & ~n17408 ) | ( x1153 & ~n17408 ) ;
  assign n17499 = ( x625 & ~x1153 ) | ( x625 & n17493 ) | ( ~x1153 & n17493 ) ;
  assign n17500 = ~n17498 & n17499 ;
  assign n17501 = n17497 | n17500 ;
  assign n17502 = x778 & n17501 ;
  assign n17503 = n17494 | n17502 ;
  assign n17504 = ~n15400 & n17503 ;
  assign n17505 = n15400 & n17408 ;
  assign n17506 = n17504 | n17505 ;
  assign n17507 = n15407 | n17506 ;
  assign n17508 = n15407 & ~n17408 ;
  assign n17509 = n17507 & ~n17508 ;
  assign n17510 = ~n15414 & n17509 ;
  assign n17511 = n17482 | n17510 ;
  assign n17512 = n15421 | n17511 ;
  assign n17513 = n15421 & ~n17408 ;
  assign n17514 = n17512 & ~n17513 ;
  assign n17515 = ~x792 & n17514 ;
  assign n17516 = ( x628 & x1156 ) | ( x628 & n17408 ) | ( x1156 & n17408 ) ;
  assign n17517 = ( ~x628 & x1156 ) | ( ~x628 & n17514 ) | ( x1156 & n17514 ) ;
  assign n17518 = n17516 & n17517 ;
  assign n17519 = ( x628 & x1156 ) | ( x628 & ~n17408 ) | ( x1156 & ~n17408 ) ;
  assign n17520 = ( x628 & ~x1156 ) | ( x628 & n17514 ) | ( ~x1156 & n17514 ) ;
  assign n17521 = ~n17519 & n17520 ;
  assign n17522 = n17518 | n17521 ;
  assign n17523 = x792 & n17522 ;
  assign n17524 = n17515 | n17523 ;
  assign n17525 = ~x787 & n17524 ;
  assign n17526 = ( x647 & x1157 ) | ( x647 & n17408 ) | ( x1157 & n17408 ) ;
  assign n17527 = ( ~x647 & x1157 ) | ( ~x647 & n17524 ) | ( x1157 & n17524 ) ;
  assign n17528 = n17526 & n17527 ;
  assign n17529 = ( x647 & x1157 ) | ( x647 & ~n17408 ) | ( x1157 & ~n17408 ) ;
  assign n17530 = ( x647 & ~x1157 ) | ( x647 & n17524 ) | ( ~x1157 & n17524 ) ;
  assign n17531 = ~n17529 & n17530 ;
  assign n17532 = n17528 | n17531 ;
  assign n17533 = x787 & n17532 ;
  assign n17534 = n17525 | n17533 ;
  assign n17535 = ( x644 & x715 ) | ( x644 & ~n17534 ) | ( x715 & ~n17534 ) ;
  assign n17536 = x630 | n17528 ;
  assign n17537 = ( x647 & x1157 ) | ( x647 & ~n17475 ) | ( x1157 & ~n17475 ) ;
  assign n17538 = x629 | n17518 ;
  assign n17539 = ( x628 & x1156 ) | ( x628 & ~n17472 ) | ( x1156 & ~n17472 ) ;
  assign n17540 = x648 | n17457 ;
  assign n17541 = ( x619 & x1159 ) | ( x619 & ~n17509 ) | ( x1159 & ~n17509 ) ;
  assign n17542 = x627 | n17447 ;
  assign n17543 = ( x618 & x1154 ) | ( x618 & ~n17506 ) | ( x1154 & ~n17506 ) ;
  assign n17544 = x660 | n17436 ;
  assign n17545 = ( x609 & x1155 ) | ( x609 & ~n17503 ) | ( x1155 & ~n17503 ) ;
  assign n17546 = x608 | n17497 ;
  assign n17547 = ( x625 & x1153 ) | ( x625 & ~n17428 ) | ( x1153 & ~n17428 ) ;
  assign n17548 = x687 | n17426 ;
  assign n17549 = x39 & ~n15797 ;
  assign n17550 = ~x39 & n15758 ;
  assign n17551 = ( x38 & n17549 ) | ( x38 & ~n17550 ) | ( n17549 & ~n17550 ) ;
  assign n17552 = x39 | n15894 ;
  assign n17553 = ( x38 & ~n17549 ) | ( x38 & n17552 ) | ( ~n17549 & n17552 ) ;
  assign n17554 = ~n17551 & n17553 ;
  assign n17555 = ( x143 & ~x774 ) | ( x143 & n17554 ) | ( ~x774 & n17554 ) ;
  assign n17556 = ~n4810 & n15904 ;
  assign n17557 = x38 & ~n17556 ;
  assign n17558 = x39 & ~n15872 ;
  assign n17559 = n14932 | n15369 ;
  assign n17560 = ~n17558 & n17559 ;
  assign n17561 = x38 | n17560 ;
  assign n17562 = ~n17557 & n17561 ;
  assign n17563 = ( x143 & x774 ) | ( x143 & n17562 ) | ( x774 & n17562 ) ;
  assign n17564 = n17555 & ~n17563 ;
  assign n17565 = x687 & ~n17564 ;
  assign n17566 = x39 | n15887 ;
  assign n17567 = x39 & ~n15583 ;
  assign n17568 = n17566 & ~n17567 ;
  assign n17569 = ~x38 & n17568 ;
  assign n17570 = n1919 & n15913 ;
  assign n17571 = x774 & ~n17570 ;
  assign n17572 = ( x143 & n17569 ) | ( x143 & ~n17571 ) | ( n17569 & ~n17571 ) ;
  assign n17573 = n15070 & ~n15477 ;
  assign n17574 = x38 & n17573 ;
  assign n17575 = x39 & n15699 ;
  assign n17576 = ~x39 & n15891 ;
  assign n17577 = n17575 | n17576 ;
  assign n17578 = ~x38 & n17577 ;
  assign n17579 = n17574 | n17578 ;
  assign n17580 = ( x143 & n17571 ) | ( x143 & n17579 ) | ( n17571 & n17579 ) ;
  assign n17581 = ~n17572 & n17580 ;
  assign n17582 = n17565 & ~n17581 ;
  assign n17583 = n2032 | n17582 ;
  assign n17584 = n17548 & ~n17583 ;
  assign n17585 = n17411 | n17584 ;
  assign n17586 = ( x625 & ~x1153 ) | ( x625 & n17585 ) | ( ~x1153 & n17585 ) ;
  assign n17587 = ~n17547 & n17586 ;
  assign n17588 = n17546 | n17587 ;
  assign n17589 = x608 & ~n17500 ;
  assign n17590 = ( x625 & x1153 ) | ( x625 & n17428 ) | ( x1153 & n17428 ) ;
  assign n17591 = ( ~x625 & x1153 ) | ( ~x625 & n17585 ) | ( x1153 & n17585 ) ;
  assign n17592 = n17590 & n17591 ;
  assign n17593 = n17589 & ~n17592 ;
  assign n17594 = n17588 & ~n17593 ;
  assign n17595 = x778 & ~n17594 ;
  assign n17596 = x778 | n17585 ;
  assign n17597 = ~n17595 & n17596 ;
  assign n17598 = ( x609 & ~x1155 ) | ( x609 & n17597 ) | ( ~x1155 & n17597 ) ;
  assign n17599 = ~n17545 & n17598 ;
  assign n17600 = n17544 | n17599 ;
  assign n17601 = x660 & ~n17440 ;
  assign n17602 = ( x609 & x1155 ) | ( x609 & n17503 ) | ( x1155 & n17503 ) ;
  assign n17603 = ( ~x609 & x1155 ) | ( ~x609 & n17597 ) | ( x1155 & n17597 ) ;
  assign n17604 = n17602 & n17603 ;
  assign n17605 = n17601 & ~n17604 ;
  assign n17606 = n17600 & ~n17605 ;
  assign n17607 = x785 & ~n17606 ;
  assign n17608 = x785 | n17597 ;
  assign n17609 = ~n17607 & n17608 ;
  assign n17610 = ( x618 & ~x1154 ) | ( x618 & n17609 ) | ( ~x1154 & n17609 ) ;
  assign n17611 = ~n17543 & n17610 ;
  assign n17612 = n17542 | n17611 ;
  assign n17613 = x627 & ~n17450 ;
  assign n17614 = ( x618 & x1154 ) | ( x618 & n17506 ) | ( x1154 & n17506 ) ;
  assign n17615 = ( ~x618 & x1154 ) | ( ~x618 & n17609 ) | ( x1154 & n17609 ) ;
  assign n17616 = n17614 & n17615 ;
  assign n17617 = n17613 & ~n17616 ;
  assign n17618 = n17612 & ~n17617 ;
  assign n17619 = x781 & ~n17618 ;
  assign n17620 = x781 | n17609 ;
  assign n17621 = ~n17619 & n17620 ;
  assign n17622 = ( x619 & ~x1159 ) | ( x619 & n17621 ) | ( ~x1159 & n17621 ) ;
  assign n17623 = ~n17541 & n17622 ;
  assign n17624 = n17540 | n17623 ;
  assign n17625 = x648 & ~n17460 ;
  assign n17626 = ( x619 & x1159 ) | ( x619 & n17509 ) | ( x1159 & n17509 ) ;
  assign n17627 = ( ~x619 & x1159 ) | ( ~x619 & n17621 ) | ( x1159 & n17621 ) ;
  assign n17628 = n17626 & n17627 ;
  assign n17629 = n17625 & ~n17628 ;
  assign n17630 = n17624 & ~n17629 ;
  assign n17631 = x789 & ~n17630 ;
  assign n17632 = x789 | n17621 ;
  assign n17633 = ~n17631 & n17632 ;
  assign n17634 = ~x788 & n17633 ;
  assign n17635 = n15972 & ~n17465 ;
  assign n17636 = ( x626 & x641 ) | ( x626 & n17511 ) | ( x641 & n17511 ) ;
  assign n17637 = ( ~x626 & x641 ) | ( ~x626 & n17633 ) | ( x641 & n17633 ) ;
  assign n17638 = n17636 | n17637 ;
  assign n17639 = ~n17635 & n17638 ;
  assign n17640 = n15978 | n17468 ;
  assign n17641 = ( x626 & x641 ) | ( x626 & ~n17511 ) | ( x641 & ~n17511 ) ;
  assign n17642 = ( x626 & ~x641 ) | ( x626 & n17633 ) | ( ~x641 & n17633 ) ;
  assign n17643 = n17641 & ~n17642 ;
  assign n17644 = n17640 & ~n17643 ;
  assign n17645 = n17639 | n17644 ;
  assign n17646 = x788 & n17645 ;
  assign n17647 = n17634 | n17646 ;
  assign n17648 = ( x628 & ~x1156 ) | ( x628 & n17647 ) | ( ~x1156 & n17647 ) ;
  assign n17649 = ~n17539 & n17648 ;
  assign n17650 = n17538 | n17649 ;
  assign n17651 = x629 & ~n17521 ;
  assign n17652 = ( x628 & x1156 ) | ( x628 & n17472 ) | ( x1156 & n17472 ) ;
  assign n17653 = ( ~x628 & x1156 ) | ( ~x628 & n17647 ) | ( x1156 & n17647 ) ;
  assign n17654 = n17652 & n17653 ;
  assign n17655 = n17651 & ~n17654 ;
  assign n17656 = n17650 & ~n17655 ;
  assign n17657 = x792 & ~n17656 ;
  assign n17658 = x792 | n17647 ;
  assign n17659 = ~n17657 & n17658 ;
  assign n17660 = ( x647 & ~x1157 ) | ( x647 & n17659 ) | ( ~x1157 & n17659 ) ;
  assign n17661 = ~n17537 & n17660 ;
  assign n17662 = n17536 | n17661 ;
  assign n17663 = x630 & ~n17531 ;
  assign n17664 = ( x647 & x1157 ) | ( x647 & n17475 ) | ( x1157 & n17475 ) ;
  assign n17665 = ( ~x647 & x1157 ) | ( ~x647 & n17659 ) | ( x1157 & n17659 ) ;
  assign n17666 = n17664 & n17665 ;
  assign n17667 = n17663 & ~n17666 ;
  assign n17668 = n17662 & ~n17667 ;
  assign n17669 = x787 & ~n17668 ;
  assign n17670 = x787 | n17659 ;
  assign n17671 = ~n17669 & n17670 ;
  assign n17672 = ( x644 & ~x715 ) | ( x644 & n17671 ) | ( ~x715 & n17671 ) ;
  assign n17673 = ~n17535 & n17672 ;
  assign n17674 = n17481 | n17673 ;
  assign n17675 = ( x644 & x715 ) | ( x644 & ~n17477 ) | ( x715 & ~n17477 ) ;
  assign n17676 = ( x644 & ~x715 ) | ( x644 & n17408 ) | ( ~x715 & n17408 ) ;
  assign n17677 = ~n17675 & n17676 ;
  assign n17678 = x1160 & ~n17677 ;
  assign n17679 = ( x644 & x715 ) | ( x644 & n17534 ) | ( x715 & n17534 ) ;
  assign n17680 = ( ~x644 & x715 ) | ( ~x644 & n17671 ) | ( x715 & n17671 ) ;
  assign n17681 = n17679 & n17680 ;
  assign n17682 = n17678 & ~n17681 ;
  assign n17683 = x790 & ~n17682 ;
  assign n17684 = n17674 & n17683 ;
  assign n17685 = ~x790 & n17671 ;
  assign n17686 = n6785 | n17685 ;
  assign n17687 = n17684 | n17686 ;
  assign n17688 = ~x143 & n6785 ;
  assign n17689 = x832 | n17688 ;
  assign n17690 = n17687 & ~n17689 ;
  assign n17691 = x143 | n1290 ;
  assign n17692 = ( x647 & x1157 ) | ( x647 & n17691 ) | ( x1157 & n17691 ) ;
  assign n17693 = x687 & n15202 ;
  assign n17694 = n17691 & ~n17693 ;
  assign n17695 = ~x778 & n17694 ;
  assign n17696 = ~x625 & n17693 ;
  assign n17697 = n17694 | n17696 ;
  assign n17698 = x1153 & n17697 ;
  assign n17699 = ~x1153 & n17691 ;
  assign n17700 = ~n17696 & n17699 ;
  assign n17701 = n17698 | n17700 ;
  assign n17702 = x778 & n17701 ;
  assign n17703 = n17695 | n17702 ;
  assign n17704 = n16043 | n17703 ;
  assign n17705 = n16045 | n17704 ;
  assign n17706 = n16047 | n17705 ;
  assign n17707 = n16049 | n17706 ;
  assign n17708 = n16055 | n17707 ;
  assign n17709 = ( ~x647 & x1157 ) | ( ~x647 & n17708 ) | ( x1157 & n17708 ) ;
  assign n17710 = n17692 & n17709 ;
  assign n17711 = x630 | n17710 ;
  assign n17712 = ~x774 & n14840 ;
  assign n17713 = n17691 & ~n17712 ;
  assign n17714 = n16060 | n17713 ;
  assign n17715 = ~x785 & n17714 ;
  assign n17716 = n16065 | n17713 ;
  assign n17717 = x1155 & n17716 ;
  assign n17718 = n16068 | n17714 ;
  assign n17719 = ~x1155 & n17718 ;
  assign n17720 = n17717 | n17719 ;
  assign n17721 = x785 & n17720 ;
  assign n17722 = n17715 | n17721 ;
  assign n17723 = ~x781 & n17722 ;
  assign n17724 = n16075 | n17722 ;
  assign n17725 = x1154 & n17724 ;
  assign n17726 = n16078 | n17722 ;
  assign n17727 = ~x1154 & n17726 ;
  assign n17728 = n17725 | n17727 ;
  assign n17729 = x781 & n17728 ;
  assign n17730 = n17723 | n17729 ;
  assign n17731 = ~x789 & n17730 ;
  assign n17732 = ( x619 & x1159 ) | ( x619 & n17691 ) | ( x1159 & n17691 ) ;
  assign n17733 = ( ~x619 & x1159 ) | ( ~x619 & n17730 ) | ( x1159 & n17730 ) ;
  assign n17734 = n17732 & n17733 ;
  assign n17735 = ( x619 & x1159 ) | ( x619 & ~n17691 ) | ( x1159 & ~n17691 ) ;
  assign n17736 = ( x619 & ~x1159 ) | ( x619 & n17730 ) | ( ~x1159 & n17730 ) ;
  assign n17737 = ~n17735 & n17736 ;
  assign n17738 = n17734 | n17737 ;
  assign n17739 = x789 & n17738 ;
  assign n17740 = n17731 | n17739 ;
  assign n17741 = ~x788 & n17740 ;
  assign n17742 = ( x626 & x1158 ) | ( x626 & n17691 ) | ( x1158 & n17691 ) ;
  assign n17743 = ( ~x1158 & n17740 ) | ( ~x1158 & n17742 ) | ( n17740 & n17742 ) ;
  assign n17744 = ( ~x626 & n17742 ) | ( ~x626 & n17743 ) | ( n17742 & n17743 ) ;
  assign n17745 = x788 & n17744 ;
  assign n17746 = n17741 | n17745 ;
  assign n17747 = n15134 | n17746 ;
  assign n17748 = n15134 & ~n17691 ;
  assign n17749 = n17747 & ~n17748 ;
  assign n17750 = ( x647 & x1157 ) | ( x647 & ~n17749 ) | ( x1157 & ~n17749 ) ;
  assign n17751 = ( x628 & x1156 ) | ( x628 & ~n17746 ) | ( x1156 & ~n17746 ) ;
  assign n17752 = n16115 & ~n17706 ;
  assign n17753 = n15420 & ~n17744 ;
  assign n17754 = n17752 | n17753 ;
  assign n17755 = x788 & n17754 ;
  assign n17756 = x648 & ~n17737 ;
  assign n17757 = ( x619 & x1159 ) | ( x619 & n17705 ) | ( x1159 & n17705 ) ;
  assign n17758 = x627 | n17725 ;
  assign n17759 = ( x618 & x1154 ) | ( x618 & ~n17704 ) | ( x1154 & ~n17704 ) ;
  assign n17760 = x660 | n17717 ;
  assign n17761 = ( x609 & x1155 ) | ( x609 & ~n17703 ) | ( x1155 & ~n17703 ) ;
  assign n17762 = n14839 | n17694 ;
  assign n17763 = x625 & ~n17762 ;
  assign n17764 = n17713 & n17762 ;
  assign n17765 = n17763 | n17764 ;
  assign n17766 = n17699 & n17765 ;
  assign n17767 = x608 | n17698 ;
  assign n17768 = n17766 | n17767 ;
  assign n17769 = x1153 & n17713 ;
  assign n17770 = ~n17763 & n17769 ;
  assign n17771 = x608 & ~n17700 ;
  assign n17772 = ~n17770 & n17771 ;
  assign n17773 = n17768 & ~n17772 ;
  assign n17774 = x778 & ~n17773 ;
  assign n17775 = x778 | n17764 ;
  assign n17776 = ~n17774 & n17775 ;
  assign n17777 = ( x609 & ~x1155 ) | ( x609 & n17776 ) | ( ~x1155 & n17776 ) ;
  assign n17778 = ~n17761 & n17777 ;
  assign n17779 = n17760 | n17778 ;
  assign n17780 = x660 & ~n17719 ;
  assign n17781 = ( x609 & x1155 ) | ( x609 & n17703 ) | ( x1155 & n17703 ) ;
  assign n17782 = ( ~x609 & x1155 ) | ( ~x609 & n17776 ) | ( x1155 & n17776 ) ;
  assign n17783 = n17781 & n17782 ;
  assign n17784 = n17780 & ~n17783 ;
  assign n17785 = n17779 & ~n17784 ;
  assign n17786 = x785 & ~n17785 ;
  assign n17787 = x785 | n17776 ;
  assign n17788 = ~n17786 & n17787 ;
  assign n17789 = ( x618 & ~x1154 ) | ( x618 & n17788 ) | ( ~x1154 & n17788 ) ;
  assign n17790 = ~n17759 & n17789 ;
  assign n17791 = n17758 | n17790 ;
  assign n17792 = x627 & ~n17727 ;
  assign n17793 = ( x618 & x1154 ) | ( x618 & n17704 ) | ( x1154 & n17704 ) ;
  assign n17794 = ( ~x618 & x1154 ) | ( ~x618 & n17788 ) | ( x1154 & n17788 ) ;
  assign n17795 = n17793 & n17794 ;
  assign n17796 = n17792 & ~n17795 ;
  assign n17797 = n17791 & ~n17796 ;
  assign n17798 = x781 & ~n17797 ;
  assign n17799 = x781 | n17788 ;
  assign n17800 = ~n17798 & n17799 ;
  assign n17801 = ( ~x619 & x1159 ) | ( ~x619 & n17800 ) | ( x1159 & n17800 ) ;
  assign n17802 = n17757 & n17801 ;
  assign n17803 = n17756 & ~n17802 ;
  assign n17804 = x648 | n17734 ;
  assign n17805 = ( x619 & x1159 ) | ( x619 & ~n17705 ) | ( x1159 & ~n17705 ) ;
  assign n17806 = ( x619 & ~x1159 ) | ( x619 & n17800 ) | ( ~x1159 & n17800 ) ;
  assign n17807 = ~n17805 & n17806 ;
  assign n17808 = n17804 | n17807 ;
  assign n17809 = x789 & n17808 ;
  assign n17810 = ~n17803 & n17809 ;
  assign n17811 = ~x789 & n17800 ;
  assign n17812 = n16177 | n17811 ;
  assign n17813 = n17810 | n17812 ;
  assign n17814 = ~n17755 & n17813 ;
  assign n17815 = ( x628 & ~x1156 ) | ( x628 & n17814 ) | ( ~x1156 & n17814 ) ;
  assign n17816 = ~n17751 & n17815 ;
  assign n17817 = n16643 & ~n17707 ;
  assign n17818 = ( x629 & x1156 ) | ( x629 & ~n17817 ) | ( x1156 & ~n17817 ) ;
  assign n17819 = n17816 | n17818 ;
  assign n17820 = ( x628 & x1156 ) | ( x628 & n17746 ) | ( x1156 & n17746 ) ;
  assign n17821 = ( ~x628 & x1156 ) | ( ~x628 & n17814 ) | ( x1156 & n17814 ) ;
  assign n17822 = n17820 & n17821 ;
  assign n17823 = n16650 | n17707 ;
  assign n17824 = ( x629 & x1156 ) | ( x629 & ~n17823 ) | ( x1156 & ~n17823 ) ;
  assign n17825 = ~n17822 & n17824 ;
  assign n17826 = n17819 & ~n17825 ;
  assign n17827 = x792 & ~n17826 ;
  assign n17828 = x792 | n17814 ;
  assign n17829 = ~n17827 & n17828 ;
  assign n17830 = ( x647 & ~x1157 ) | ( x647 & n17829 ) | ( ~x1157 & n17829 ) ;
  assign n17831 = ~n17750 & n17830 ;
  assign n17832 = n17711 | n17831 ;
  assign n17833 = ( x647 & x1157 ) | ( x647 & ~n17691 ) | ( x1157 & ~n17691 ) ;
  assign n17834 = ( x647 & ~x1157 ) | ( x647 & n17708 ) | ( ~x1157 & n17708 ) ;
  assign n17835 = ~n17833 & n17834 ;
  assign n17836 = x630 & ~n17835 ;
  assign n17837 = ( x647 & x1157 ) | ( x647 & n17749 ) | ( x1157 & n17749 ) ;
  assign n17838 = ( ~x647 & x1157 ) | ( ~x647 & n17829 ) | ( x1157 & n17829 ) ;
  assign n17839 = n17837 & n17838 ;
  assign n17840 = n17836 & ~n17839 ;
  assign n17841 = n17832 & ~n17840 ;
  assign n17842 = x787 & ~n17841 ;
  assign n17843 = x787 | n17829 ;
  assign n17844 = ~n17842 & n17843 ;
  assign n17845 = ( x790 & x832 ) | ( x790 & n17844 ) | ( x832 & n17844 ) ;
  assign n17846 = n15141 & n17691 ;
  assign n17847 = ~n15141 & n17749 ;
  assign n17848 = n17846 | n17847 ;
  assign n17849 = ( x644 & x715 ) | ( x644 & ~n17848 ) | ( x715 & ~n17848 ) ;
  assign n17850 = ( x644 & ~x715 ) | ( x644 & n17691 ) | ( ~x715 & n17691 ) ;
  assign n17851 = ~n17849 & n17850 ;
  assign n17852 = x1160 & ~n17851 ;
  assign n17853 = ~x787 & n17708 ;
  assign n17854 = n17710 | n17835 ;
  assign n17855 = x787 & n17854 ;
  assign n17856 = n17853 | n17855 ;
  assign n17857 = ( x644 & x715 ) | ( x644 & n17856 ) | ( x715 & n17856 ) ;
  assign n17858 = ( ~x644 & x715 ) | ( ~x644 & n17844 ) | ( x715 & n17844 ) ;
  assign n17859 = n17857 & n17858 ;
  assign n17860 = n17852 & ~n17859 ;
  assign n17861 = ( x644 & x715 ) | ( x644 & n17848 ) | ( x715 & n17848 ) ;
  assign n17862 = ( ~x644 & x715 ) | ( ~x644 & n17691 ) | ( x715 & n17691 ) ;
  assign n17863 = n17861 & n17862 ;
  assign n17864 = x1160 | n17863 ;
  assign n17865 = ( x644 & x715 ) | ( x644 & ~n17856 ) | ( x715 & ~n17856 ) ;
  assign n17866 = ( x644 & ~x715 ) | ( x644 & n17844 ) | ( ~x715 & n17844 ) ;
  assign n17867 = ~n17865 & n17866 ;
  assign n17868 = n17864 | n17867 ;
  assign n17869 = ~n17860 & n17868 ;
  assign n17870 = ( ~x790 & x832 ) | ( ~x790 & n17869 ) | ( x832 & n17869 ) ;
  assign n17871 = n17845 & n17870 ;
  assign n17872 = n17690 | n17871 ;
  assign n17873 = x144 & ~n14830 ;
  assign n17874 = x144 & n14828 ;
  assign n17875 = ( ~n14936 & n17873 ) | ( ~n14936 & n17874 ) | ( n17873 & n17874 ) ;
  assign n17876 = n15421 & n17875 ;
  assign n17877 = n15421 & ~n17876 ;
  assign n17878 = x628 & n17877 ;
  assign n17879 = x628 | n17873 ;
  assign n17880 = x628 | n17874 ;
  assign n17881 = ( ~n14936 & n17879 ) | ( ~n14936 & n17880 ) | ( n17879 & n17880 ) ;
  assign n17882 = x1156 & n17881 ;
  assign n17883 = ~n17878 & n17882 ;
  assign n17884 = x628 & ~n17876 ;
  assign n17885 = n17882 & ~n17884 ;
  assign n17886 = n15414 & ~n17875 ;
  assign n17887 = x736 & ~n2032 ;
  assign n17888 = n17875 | n17887 ;
  assign n17889 = ~n4809 & n15313 ;
  assign n17890 = ~n1271 & n17889 ;
  assign n17891 = ~n1242 & n17890 ;
  assign n17892 = x38 & ~n17891 ;
  assign n17893 = x144 | n15070 ;
  assign n17894 = n17887 & ~n17893 ;
  assign n17895 = ( n17887 & ~n17892 ) | ( n17887 & n17894 ) | ( ~n17892 & n17894 ) ;
  assign n17896 = n17888 & ~n17895 ;
  assign n17897 = ( ~x38 & x144 ) | ( ~x38 & n16323 ) | ( x144 & n16323 ) ;
  assign n17898 = ( x38 & x144 ) | ( x38 & n16319 ) | ( x144 & n16319 ) ;
  assign n17899 = n17897 & ~n17898 ;
  assign n17900 = ( n17888 & n17896 ) | ( n17888 & n17899 ) | ( n17896 & n17899 ) ;
  assign n17901 = ~x778 & n17900 ;
  assign n17902 = x625 | n17873 ;
  assign n17903 = x625 | n17874 ;
  assign n17904 = ( ~n14936 & n17902 ) | ( ~n14936 & n17903 ) | ( n17902 & n17903 ) ;
  assign n17905 = x1153 & n17904 ;
  assign n17906 = ~x625 & n17905 ;
  assign n17907 = ( n17900 & n17905 ) | ( n17900 & n17906 ) | ( n17905 & n17906 ) ;
  assign n17908 = x625 & ~n17873 ;
  assign n17909 = x625 & ~n17874 ;
  assign n17910 = ( n14936 & n17908 ) | ( n14936 & n17909 ) | ( n17908 & n17909 ) ;
  assign n17911 = x1153 | n17910 ;
  assign n17912 = x625 & ~n17911 ;
  assign n17913 = ( n17900 & ~n17911 ) | ( n17900 & n17912 ) | ( ~n17911 & n17912 ) ;
  assign n17914 = n17907 | n17913 ;
  assign n17915 = x778 | n17901 ;
  assign n17916 = ( n17901 & n17914 ) | ( n17901 & n17915 ) | ( n17914 & n17915 ) ;
  assign n17917 = n15400 & ~n17875 ;
  assign n17918 = n15400 & ~n17917 ;
  assign n17919 = ~n15407 & n17918 ;
  assign n17920 = n15407 & n17875 ;
  assign n17921 = n17919 | n17920 ;
  assign n17922 = n15414 | n17921 ;
  assign n17923 = n15407 | n17917 ;
  assign n17924 = ~n17920 & n17923 ;
  assign n17925 = ~n15414 & n17924 ;
  assign n17926 = ( n17916 & n17922 ) | ( n17916 & ~n17925 ) | ( n17922 & ~n17925 ) ;
  assign n17927 = ~n17886 & n17926 ;
  assign n17928 = ( n17883 & n17885 ) | ( n17883 & n17927 ) | ( n17885 & n17927 ) ;
  assign n17929 = ~x628 & n17877 ;
  assign n17930 = x628 & ~n17873 ;
  assign n17931 = x628 & ~n17874 ;
  assign n17932 = ( n14936 & n17930 ) | ( n14936 & n17931 ) | ( n17930 & n17931 ) ;
  assign n17933 = x1156 | n17932 ;
  assign n17934 = n17929 | n17933 ;
  assign n17935 = x628 | n17876 ;
  assign n17936 = ~n17933 & n17935 ;
  assign n17937 = ( n17927 & ~n17934 ) | ( n17927 & n17936 ) | ( ~n17934 & n17936 ) ;
  assign n17938 = n17928 | n17937 ;
  assign n17939 = ( n17876 & ~n17877 ) | ( n17876 & n17927 ) | ( ~n17877 & n17927 ) ;
  assign n17940 = ~x792 & n17939 ;
  assign n17941 = x792 | n17940 ;
  assign n17942 = ( n17938 & n17940 ) | ( n17938 & n17941 ) | ( n17940 & n17941 ) ;
  assign n17943 = ~x787 & n17942 ;
  assign n17944 = x647 | n17873 ;
  assign n17945 = x647 | n17874 ;
  assign n17946 = ( ~n14936 & n17944 ) | ( ~n14936 & n17945 ) | ( n17944 & n17945 ) ;
  assign n17947 = x1157 & n17946 ;
  assign n17948 = ~x647 & n17947 ;
  assign n17949 = ( n17942 & n17947 ) | ( n17942 & n17948 ) | ( n17947 & n17948 ) ;
  assign n17950 = x647 & ~n17873 ;
  assign n17951 = x647 & ~n17874 ;
  assign n17952 = ( n14936 & n17950 ) | ( n14936 & n17951 ) | ( n17950 & n17951 ) ;
  assign n17953 = x1157 | n17952 ;
  assign n17954 = x647 & ~n17953 ;
  assign n17955 = ( n17942 & ~n17953 ) | ( n17942 & n17954 ) | ( ~n17953 & n17954 ) ;
  assign n17956 = n17949 | n17955 ;
  assign n17957 = x787 | n17943 ;
  assign n17958 = ( n17943 & n17956 ) | ( n17943 & n17957 ) | ( n17956 & n17957 ) ;
  assign n17959 = x644 | x715 ;
  assign n17960 = ( x715 & ~n17958 ) | ( x715 & n17959 ) | ( ~n17958 & n17959 ) ;
  assign n17961 = n15134 & n17875 ;
  assign n17962 = n15141 | n17961 ;
  assign n17963 = n15141 & ~n17875 ;
  assign n17964 = n17962 & ~n17963 ;
  assign n17965 = x644 | n17964 ;
  assign n17966 = x644 & ~n17873 ;
  assign n17967 = x644 & ~n17874 ;
  assign n17968 = ( n14936 & n17966 ) | ( n14936 & n17967 ) | ( n17966 & n17967 ) ;
  assign n17969 = x715 & ~n17968 ;
  assign n17970 = n17965 & n17969 ;
  assign n17971 = ~x644 & n17963 ;
  assign n17972 = n17969 & ~n17971 ;
  assign n17973 = x144 & n2032 ;
  assign n17974 = n15082 | n17973 ;
  assign n17975 = n15082 & ~n17875 ;
  assign n17976 = n17974 & ~n17975 ;
  assign n17977 = n2032 & ~n17973 ;
  assign n17978 = ~n15082 & n17977 ;
  assign n17979 = n17975 | n17978 ;
  assign n17980 = x38 & n17893 ;
  assign n17981 = x603 & x758 ;
  assign n17982 = ( n14838 & n15070 ) | ( n14838 & ~n17981 ) | ( n15070 & ~n17981 ) ;
  assign n17983 = n15070 & n17982 ;
  assign n17984 = n17980 & ~n17983 ;
  assign n17985 = x758 & ~n15061 ;
  assign n17986 = x758 | n14710 ;
  assign n17987 = ~n17985 & n17986 ;
  assign n17988 = x39 & ~n17987 ;
  assign n17989 = ( x39 & x758 ) | ( x39 & n14956 ) | ( x758 & n14956 ) ;
  assign n17990 = ( x39 & ~x758 ) | ( x39 & n14822 ) | ( ~x758 & n14822 ) ;
  assign n17991 = n17989 | n17990 ;
  assign n17992 = x144 & ~n17991 ;
  assign n17993 = ( x144 & n17988 ) | ( x144 & n17992 ) | ( n17988 & n17992 ) ;
  assign n17994 = ~x144 & x758 ;
  assign n17995 = ~n14908 & n17994 ;
  assign n17996 = n14932 & n17995 ;
  assign n17997 = x38 | n17996 ;
  assign n17998 = n17993 | n17997 ;
  assign n17999 = ( ~x38 & n17984 ) | ( ~x38 & n17998 ) | ( n17984 & n17998 ) ;
  assign n18000 = ( n17976 & ~n17979 ) | ( n17976 & n17999 ) | ( ~n17979 & n17999 ) ;
  assign n18001 = x609 & ~n18000 ;
  assign n18002 = x609 | n17873 ;
  assign n18003 = x609 | n17874 ;
  assign n18004 = ( ~n14936 & n18002 ) | ( ~n14936 & n18003 ) | ( n18002 & n18003 ) ;
  assign n18005 = x1155 & n18004 ;
  assign n18006 = ~n18001 & n18005 ;
  assign n18007 = x609 | n18000 ;
  assign n18008 = x609 & ~n17873 ;
  assign n18009 = x609 & ~n17874 ;
  assign n18010 = ( n14936 & n18008 ) | ( n14936 & n18009 ) | ( n18008 & n18009 ) ;
  assign n18011 = x1155 | n18010 ;
  assign n18012 = n18007 & ~n18011 ;
  assign n18013 = n18006 | n18012 ;
  assign n18014 = ~x785 & n18000 ;
  assign n18015 = x785 | n18014 ;
  assign n18016 = ( n18013 & n18014 ) | ( n18013 & n18015 ) | ( n18014 & n18015 ) ;
  assign n18017 = x618 & ~n18016 ;
  assign n18018 = x618 | n17873 ;
  assign n18019 = x618 | n17874 ;
  assign n18020 = ( ~n14936 & n18018 ) | ( ~n14936 & n18019 ) | ( n18018 & n18019 ) ;
  assign n18021 = x1154 & n18020 ;
  assign n18022 = ~n18017 & n18021 ;
  assign n18023 = x618 | n18016 ;
  assign n18024 = x618 & ~n17873 ;
  assign n18025 = x618 & ~n17874 ;
  assign n18026 = ( n14936 & n18024 ) | ( n14936 & n18025 ) | ( n18024 & n18025 ) ;
  assign n18027 = x1154 | n18026 ;
  assign n18028 = n18023 & ~n18027 ;
  assign n18029 = n18022 | n18028 ;
  assign n18030 = ~x781 & n18016 ;
  assign n18031 = x781 | n18030 ;
  assign n18032 = ( n18029 & n18030 ) | ( n18029 & n18031 ) | ( n18030 & n18031 ) ;
  assign n18033 = x619 & ~n18032 ;
  assign n18034 = x619 | n17873 ;
  assign n18035 = x619 | n17874 ;
  assign n18036 = ( ~n14936 & n18034 ) | ( ~n14936 & n18035 ) | ( n18034 & n18035 ) ;
  assign n18037 = x1159 & n18036 ;
  assign n18038 = ~n18033 & n18037 ;
  assign n18039 = x619 | n18032 ;
  assign n18040 = x619 & ~n17873 ;
  assign n18041 = x619 & ~n17874 ;
  assign n18042 = ( n14936 & n18040 ) | ( n14936 & n18041 ) | ( n18040 & n18041 ) ;
  assign n18043 = x1159 | n18042 ;
  assign n18044 = n18039 & ~n18043 ;
  assign n18045 = n18038 | n18044 ;
  assign n18046 = ~x789 & n18032 ;
  assign n18047 = x789 | n18046 ;
  assign n18048 = ( n18045 & n18046 ) | ( n18045 & n18047 ) | ( n18046 & n18047 ) ;
  assign n18049 = x626 | n18048 ;
  assign n18050 = x626 & ~n17873 ;
  assign n18051 = x626 & ~n17874 ;
  assign n18052 = ( n14936 & n18050 ) | ( n14936 & n18051 ) | ( n18050 & n18051 ) ;
  assign n18053 = x1158 | n18052 ;
  assign n18054 = n18049 & ~n18053 ;
  assign n18055 = x626 & ~n18048 ;
  assign n18056 = x626 | n17873 ;
  assign n18057 = x626 | n17874 ;
  assign n18058 = ( ~n14936 & n18056 ) | ( ~n14936 & n18057 ) | ( n18056 & n18057 ) ;
  assign n18059 = x1158 & n18058 ;
  assign n18060 = ~n18055 & n18059 ;
  assign n18061 = n18054 | n18060 ;
  assign n18062 = ~x788 & n18048 ;
  assign n18063 = x788 | n18062 ;
  assign n18064 = ( n18061 & n18062 ) | ( n18061 & n18063 ) | ( n18062 & n18063 ) ;
  assign n18065 = ~n15134 & n18064 ;
  assign n18066 = ( n17970 & n17972 ) | ( n17970 & n18065 ) | ( n17972 & n18065 ) ;
  assign n18067 = x1160 | n18066 ;
  assign n18068 = x647 & ~n17961 ;
  assign n18069 = x1157 | n18068 ;
  assign n18070 = ( x1157 & ~n18065 ) | ( x1157 & n18069 ) | ( ~n18065 & n18069 ) ;
  assign n18071 = x630 | n17949 ;
  assign n18072 = x628 & ~n18064 ;
  assign n18073 = x1156 | n18072 ;
  assign n18074 = x629 | n17928 ;
  assign n18075 = x619 & ~n17921 ;
  assign n18076 = x619 & n17924 ;
  assign n18077 = ( ~n17916 & n18075 ) | ( ~n17916 & n18076 ) | ( n18075 & n18076 ) ;
  assign n18078 = x1159 | n18077 ;
  assign n18079 = x648 | n18038 ;
  assign n18080 = x618 & ~n17918 ;
  assign n18081 = x618 & n17917 ;
  assign n18082 = ( ~n17916 & n18080 ) | ( ~n17916 & n18081 ) | ( n18080 & n18081 ) ;
  assign n18083 = x1154 | n18082 ;
  assign n18084 = x627 | n18022 ;
  assign n18085 = x609 | x1155 ;
  assign n18086 = ( x1155 & ~n17916 ) | ( x1155 & n18085 ) | ( ~n17916 & n18085 ) ;
  assign n18087 = x660 | n18006 ;
  assign n18088 = x625 & n17977 ;
  assign n18089 = x625 & ~n17973 ;
  assign n18090 = ( ~n17999 & n18088 ) | ( ~n17999 & n18089 ) | ( n18088 & n18089 ) ;
  assign n18091 = x1153 | n18090 ;
  assign n18092 = x608 | n17907 ;
  assign n18093 = x736 & ~n17570 ;
  assign n18094 = ~n17984 & n18093 ;
  assign n18095 = x144 & n15699 ;
  assign n18096 = x144 & ~x758 ;
  assign n18097 = ( ~x758 & n15583 ) | ( ~x758 & n18096 ) | ( n15583 & n18096 ) ;
  assign n18098 = ~n18095 & n18097 ;
  assign n18099 = x144 | n15872 ;
  assign n18100 = ( x758 & ~n15797 ) | ( x758 & n17994 ) | ( ~n15797 & n17994 ) ;
  assign n18101 = x39 & ~n18100 ;
  assign n18102 = ( x39 & ~n18099 ) | ( x39 & n18101 ) | ( ~n18099 & n18101 ) ;
  assign n18103 = ~n18098 & n18102 ;
  assign n18104 = n18094 & n18103 ;
  assign n18105 = ( ~x758 & n15887 ) | ( ~x758 & n18096 ) | ( n15887 & n18096 ) ;
  assign n18106 = x144 & n15891 ;
  assign n18107 = n18105 & ~n18106 ;
  assign n18108 = ( x144 & ~x758 ) | ( x144 & n15894 ) | ( ~x758 & n15894 ) ;
  assign n18109 = ( x144 & x758 ) | ( x144 & n15897 ) | ( x758 & n15897 ) ;
  assign n18110 = ~n18108 & n18109 ;
  assign n18111 = n18107 | n18110 ;
  assign n18112 = ( ~x38 & n9138 ) | ( ~x38 & n18111 ) | ( n9138 & n18111 ) ;
  assign n18113 = ( n18094 & n18104 ) | ( n18094 & ~n18112 ) | ( n18104 & ~n18112 ) ;
  assign n18114 = n2032 | n18113 ;
  assign n18115 = x736 | n17999 ;
  assign n18116 = n17973 | n18115 ;
  assign n18117 = ( n17973 & ~n18114 ) | ( n17973 & n18116 ) | ( ~n18114 & n18116 ) ;
  assign n18118 = n18091 | n18117 ;
  assign n18119 = x625 | n18118 ;
  assign n18120 = ( ~n18091 & n18092 ) | ( ~n18091 & n18119 ) | ( n18092 & n18119 ) ;
  assign n18121 = ~x625 & n17977 ;
  assign n18122 = x625 | n17973 ;
  assign n18123 = ( n17999 & ~n18121 ) | ( n17999 & n18122 ) | ( ~n18121 & n18122 ) ;
  assign n18124 = x1153 & n18123 ;
  assign n18125 = x608 & ~n17913 ;
  assign n18126 = ~n18117 & n18124 ;
  assign n18127 = x625 & n18126 ;
  assign n18128 = ( ~n18124 & n18125 ) | ( ~n18124 & n18127 ) | ( n18125 & n18127 ) ;
  assign n18129 = n18120 & ~n18128 ;
  assign n18130 = x778 | n18117 ;
  assign n18131 = ~x778 & n18130 ;
  assign n18132 = ( n18129 & n18130 ) | ( n18129 & n18131 ) | ( n18130 & n18131 ) ;
  assign n18133 = n18086 | n18132 ;
  assign n18134 = x609 | n18133 ;
  assign n18135 = ( ~n18086 & n18087 ) | ( ~n18086 & n18134 ) | ( n18087 & n18134 ) ;
  assign n18136 = x609 & x1155 ;
  assign n18137 = ( x1155 & n17916 ) | ( x1155 & n18136 ) | ( n17916 & n18136 ) ;
  assign n18138 = x660 & ~n18012 ;
  assign n18139 = ~n18132 & n18137 ;
  assign n18140 = x609 & n18139 ;
  assign n18141 = ( ~n18137 & n18138 ) | ( ~n18137 & n18140 ) | ( n18138 & n18140 ) ;
  assign n18142 = n18135 & ~n18141 ;
  assign n18143 = x785 | n18132 ;
  assign n18144 = ~x785 & n18143 ;
  assign n18145 = ( n18142 & n18143 ) | ( n18142 & n18144 ) | ( n18143 & n18144 ) ;
  assign n18146 = n18083 | n18145 ;
  assign n18147 = x618 | n18146 ;
  assign n18148 = ( ~n18083 & n18084 ) | ( ~n18083 & n18147 ) | ( n18084 & n18147 ) ;
  assign n18149 = x618 | n17918 ;
  assign n18150 = ~x618 & n17917 ;
  assign n18151 = ( n17916 & n18149 ) | ( n17916 & ~n18150 ) | ( n18149 & ~n18150 ) ;
  assign n18152 = x1154 & n18151 ;
  assign n18153 = x627 & ~n18028 ;
  assign n18154 = ~n18145 & n18152 ;
  assign n18155 = x618 & n18154 ;
  assign n18156 = ( ~n18152 & n18153 ) | ( ~n18152 & n18155 ) | ( n18153 & n18155 ) ;
  assign n18157 = n18148 & ~n18156 ;
  assign n18158 = x781 | n18145 ;
  assign n18159 = ~x781 & n18158 ;
  assign n18160 = ( n18157 & n18158 ) | ( n18157 & n18159 ) | ( n18158 & n18159 ) ;
  assign n18161 = n18078 | n18160 ;
  assign n18162 = x619 | n18161 ;
  assign n18163 = ( ~n18078 & n18079 ) | ( ~n18078 & n18162 ) | ( n18079 & n18162 ) ;
  assign n18164 = x619 | n17921 ;
  assign n18165 = ~x619 & n17924 ;
  assign n18166 = ( n17916 & n18164 ) | ( n17916 & ~n18165 ) | ( n18164 & ~n18165 ) ;
  assign n18167 = x1159 & n18166 ;
  assign n18168 = x648 & ~n18044 ;
  assign n18169 = ~n18160 & n18167 ;
  assign n18170 = x619 & n18169 ;
  assign n18171 = ( ~n18167 & n18168 ) | ( ~n18167 & n18170 ) | ( n18168 & n18170 ) ;
  assign n18172 = n18163 & ~n18171 ;
  assign n18173 = x789 | n18160 ;
  assign n18174 = ~x789 & n18173 ;
  assign n18175 = ( n18172 & n18173 ) | ( n18172 & n18174 ) | ( n18173 & n18174 ) ;
  assign n18176 = ~x788 & n18175 ;
  assign n18177 = x626 | x641 ;
  assign n18178 = ( x641 & n17927 ) | ( x641 & n18177 ) | ( n17927 & n18177 ) ;
  assign n18179 = n15972 & ~n18054 ;
  assign n18180 = n18175 & ~n18178 ;
  assign n18181 = ~x626 & n18180 ;
  assign n18182 = ( n18178 & ~n18179 ) | ( n18178 & n18181 ) | ( ~n18179 & n18181 ) ;
  assign n18183 = x626 & x641 ;
  assign n18184 = ( x641 & ~n17927 ) | ( x641 & n18183 ) | ( ~n17927 & n18183 ) ;
  assign n18185 = n15978 | n18060 ;
  assign n18186 = n18175 & n18184 ;
  assign n18187 = x626 & n18186 ;
  assign n18188 = ( ~n18184 & n18185 ) | ( ~n18184 & n18187 ) | ( n18185 & n18187 ) ;
  assign n18189 = n18182 | n18188 ;
  assign n18190 = x788 | n18176 ;
  assign n18191 = ( n18176 & n18189 ) | ( n18176 & n18190 ) | ( n18189 & n18190 ) ;
  assign n18192 = n18073 | n18191 ;
  assign n18193 = x628 | n18192 ;
  assign n18194 = ( ~n18073 & n18074 ) | ( ~n18073 & n18193 ) | ( n18074 & n18193 ) ;
  assign n18195 = x628 | n18064 ;
  assign n18196 = x1156 & n18195 ;
  assign n18197 = x629 & ~n17937 ;
  assign n18198 = ~n18191 & n18196 ;
  assign n18199 = x628 & n18198 ;
  assign n18200 = ( ~n18196 & n18197 ) | ( ~n18196 & n18199 ) | ( n18197 & n18199 ) ;
  assign n18201 = n18194 & ~n18200 ;
  assign n18202 = x792 | n18191 ;
  assign n18203 = ~x792 & n18202 ;
  assign n18204 = ( n18201 & n18202 ) | ( n18201 & n18203 ) | ( n18202 & n18203 ) ;
  assign n18205 = n18070 | n18204 ;
  assign n18206 = x647 | n18205 ;
  assign n18207 = ( ~n18070 & n18071 ) | ( ~n18070 & n18206 ) | ( n18071 & n18206 ) ;
  assign n18208 = x647 | n17961 ;
  assign n18209 = x1157 & n18208 ;
  assign n18210 = ( x1157 & n18065 ) | ( x1157 & n18209 ) | ( n18065 & n18209 ) ;
  assign n18211 = x630 & ~n17955 ;
  assign n18212 = ~n18204 & n18210 ;
  assign n18213 = x647 & n18212 ;
  assign n18214 = ( ~n18210 & n18211 ) | ( ~n18210 & n18213 ) | ( n18211 & n18213 ) ;
  assign n18215 = n18207 & ~n18214 ;
  assign n18216 = x787 | n18204 ;
  assign n18217 = ~x787 & n18216 ;
  assign n18218 = ( n18215 & n18216 ) | ( n18215 & n18217 ) | ( n18216 & n18217 ) ;
  assign n18219 = n17960 | n18218 ;
  assign n18220 = x644 | n18219 ;
  assign n18221 = ( ~n17960 & n18067 ) | ( ~n17960 & n18220 ) | ( n18067 & n18220 ) ;
  assign n18222 = x644 & x715 ;
  assign n18223 = ( x715 & n17958 ) | ( x715 & n18222 ) | ( n17958 & n18222 ) ;
  assign n18224 = x644 & ~n17964 ;
  assign n18225 = x644 | n17873 ;
  assign n18226 = x644 | n17874 ;
  assign n18227 = ( ~n14936 & n18225 ) | ( ~n14936 & n18226 ) | ( n18225 & n18226 ) ;
  assign n18228 = ~x715 & n18227 ;
  assign n18229 = ~n18224 & n18228 ;
  assign n18230 = x644 & n17963 ;
  assign n18231 = n18228 & ~n18230 ;
  assign n18232 = ( n18065 & n18229 ) | ( n18065 & n18231 ) | ( n18229 & n18231 ) ;
  assign n18233 = x1160 & ~n18232 ;
  assign n18234 = ~n18223 & n18233 ;
  assign n18235 = ~x644 & n18223 ;
  assign n18236 = n18233 & ~n18235 ;
  assign n18237 = ( ~n18218 & n18234 ) | ( ~n18218 & n18236 ) | ( n18234 & n18236 ) ;
  assign n18238 = x790 & ~n18237 ;
  assign n18239 = n18221 & n18238 ;
  assign n18240 = ~x57 & x144 ;
  assign n18241 = ( x57 & n4832 ) | ( x57 & ~n18240 ) | ( n4832 & ~n18240 ) ;
  assign n18242 = x790 & ~n4832 ;
  assign n18243 = ( n4832 & n18218 ) | ( n4832 & ~n18242 ) | ( n18218 & ~n18242 ) ;
  assign n18244 = ~n18241 & n18243 ;
  assign n18245 = ( n18239 & ~n18241 ) | ( n18239 & n18244 ) | ( ~n18241 & n18244 ) ;
  assign n18246 = x618 & x1154 ;
  assign n18247 = x618 | x1154 ;
  assign n18248 = x781 & n18247 ;
  assign n18249 = ~n18246 & n18248 ;
  assign n18250 = ~x619 & x1159 ;
  assign n18251 = x619 & ~x1159 ;
  assign n18252 = n18250 | n18251 ;
  assign n18253 = x789 & n18252 ;
  assign n18254 = n15082 | n18253 ;
  assign n18255 = n18249 | n18254 ;
  assign n18256 = x785 & n18085 ;
  assign n18257 = ~n18136 & n18256 ;
  assign n18258 = x758 & n14840 ;
  assign n18259 = ~n18257 & n18258 ;
  assign n18260 = ~n16176 & n18259 ;
  assign n18261 = ~n18255 & n18260 ;
  assign n18262 = x144 & ~n1290 ;
  assign n18263 = x715 | n18262 ;
  assign n18264 = n15134 | n15141 ;
  assign n18265 = x644 & ~n18264 ;
  assign n18266 = n18263 | n18265 ;
  assign n18267 = ( n18261 & n18263 ) | ( n18261 & n18266 ) | ( n18263 & n18266 ) ;
  assign n18268 = x1160 & n18267 ;
  assign n18269 = x626 & n18259 ;
  assign n18270 = ~n18255 & n18269 ;
  assign n18271 = ( x641 & n15972 ) | ( x641 & n18262 ) | ( n15972 & n18262 ) ;
  assign n18272 = ( n15972 & n18270 ) | ( n15972 & n18271 ) | ( n18270 & n18271 ) ;
  assign n18273 = n15414 & ~n18262 ;
  assign n18274 = n18262 & ~n18273 ;
  assign n18275 = n15407 & ~n18262 ;
  assign n18276 = n18273 | n18275 ;
  assign n18277 = x736 & n15202 ;
  assign n18278 = n18262 | n18277 ;
  assign n18279 = x625 & n18277 ;
  assign n18280 = n18278 & ~n18279 ;
  assign n18281 = x1153 & ~n18262 ;
  assign n18282 = ~n18279 & n18281 ;
  assign n18283 = x1153 & ~n18282 ;
  assign n18284 = ( n18280 & ~n18282 ) | ( n18280 & n18283 ) | ( ~n18282 & n18283 ) ;
  assign n18285 = x778 | n18278 ;
  assign n18286 = ~x778 & n18285 ;
  assign n18287 = ( n18284 & n18285 ) | ( n18284 & n18286 ) | ( n18285 & n18286 ) ;
  assign n18288 = ~n15400 & n18287 ;
  assign n18289 = ( n18274 & ~n18276 ) | ( n18274 & n18288 ) | ( ~n18276 & n18288 ) ;
  assign n18290 = n16110 & n18289 ;
  assign n18291 = n18272 | n18290 ;
  assign n18292 = ~x626 & n18259 ;
  assign n18293 = ~n18255 & n18292 ;
  assign n18294 = ~x1158 & n18262 ;
  assign n18295 = x641 & ~n18294 ;
  assign n18296 = ( n15978 & ~n18293 ) | ( n15978 & n18295 ) | ( ~n18293 & n18295 ) ;
  assign n18297 = x788 & ~n18296 ;
  assign n18298 = n16109 & n18289 ;
  assign n18299 = ( x788 & n18297 ) | ( x788 & n18298 ) | ( n18297 & n18298 ) ;
  assign n18300 = n18291 & n18299 ;
  assign n18301 = x619 | x778 ;
  assign n18302 = ( x619 & n15081 ) | ( x619 & n18301 ) | ( n15081 & n18301 ) ;
  assign n18303 = n18249 | n18302 ;
  assign n18304 = n18259 & ~n18303 ;
  assign n18305 = x1159 | n18262 ;
  assign n18306 = x648 & n18305 ;
  assign n18307 = ( x648 & n18304 ) | ( x648 & n18306 ) | ( n18304 & n18306 ) ;
  assign n18308 = x619 | n18275 ;
  assign n18309 = ~x619 & n18262 ;
  assign n18310 = ( n18288 & ~n18308 ) | ( n18288 & n18309 ) | ( ~n18308 & n18309 ) ;
  assign n18311 = x1159 & ~n18310 ;
  assign n18312 = n18307 & ~n18311 ;
  assign n18313 = x1154 & ~n18262 ;
  assign n18314 = x618 & ~x778 ;
  assign n18315 = ( x618 & ~n15081 ) | ( x618 & n18314 ) | ( ~n15081 & n18314 ) ;
  assign n18316 = n18313 & ~n18315 ;
  assign n18317 = ( ~n18259 & n18313 ) | ( ~n18259 & n18316 ) | ( n18313 & n18316 ) ;
  assign n18318 = x627 | n18317 ;
  assign n18319 = x618 & n18262 ;
  assign n18320 = x1154 | n18319 ;
  assign n18321 = ( n18247 & n18288 ) | ( n18247 & n18320 ) | ( n18288 & n18320 ) ;
  assign n18322 = ~n18318 & n18321 ;
  assign n18323 = n15088 & n18258 ;
  assign n18324 = x1155 & ~n18262 ;
  assign n18325 = x660 | n18324 ;
  assign n18326 = ( x660 & ~n18323 ) | ( x660 & n18325 ) | ( ~n18323 & n18325 ) ;
  assign n18327 = x609 & n18287 ;
  assign n18328 = x1155 | n18327 ;
  assign n18329 = ~n18326 & n18328 ;
  assign n18330 = x736 & n15529 ;
  assign n18331 = x625 & n18330 ;
  assign n18332 = n18258 | n18262 ;
  assign n18333 = x1153 & ~n18332 ;
  assign n18334 = ~n18331 & n18333 ;
  assign n18335 = x608 & x1153 ;
  assign n18336 = ( x608 & n18280 ) | ( x608 & n18335 ) | ( n18280 & n18335 ) ;
  assign n18337 = ~n18334 & n18336 ;
  assign n18338 = n18330 | n18332 ;
  assign n18339 = ~n18331 & n18338 ;
  assign n18340 = x608 | n18282 ;
  assign n18341 = x1153 & ~n18340 ;
  assign n18342 = ( n18339 & ~n18340 ) | ( n18339 & n18341 ) | ( ~n18340 & n18341 ) ;
  assign n18343 = n18337 | n18342 ;
  assign n18344 = ~x778 & n18338 ;
  assign n18345 = x778 | n18344 ;
  assign n18346 = ( n18343 & n18344 ) | ( n18343 & n18345 ) | ( n18344 & n18345 ) ;
  assign n18347 = ~x609 & n18346 ;
  assign n18348 = ( ~n18326 & n18329 ) | ( ~n18326 & n18347 ) | ( n18329 & n18347 ) ;
  assign n18349 = ~n15094 & n18258 ;
  assign n18350 = x1155 | n18262 ;
  assign n18351 = x660 & n18350 ;
  assign n18352 = ( x660 & n18349 ) | ( x660 & n18351 ) | ( n18349 & n18351 ) ;
  assign n18353 = ~x609 & n18287 ;
  assign n18354 = x1155 & ~n18353 ;
  assign n18355 = n18352 & ~n18354 ;
  assign n18356 = x609 & n18346 ;
  assign n18357 = ( n18352 & n18355 ) | ( n18352 & n18356 ) | ( n18355 & n18356 ) ;
  assign n18358 = n18348 | n18357 ;
  assign n18359 = ~x785 & n18346 ;
  assign n18360 = x785 | n18359 ;
  assign n18361 = ( n18358 & n18359 ) | ( n18358 & n18360 ) | ( n18359 & n18360 ) ;
  assign n18362 = ~x618 & n18361 ;
  assign n18363 = ( ~n18318 & n18322 ) | ( ~n18318 & n18362 ) | ( n18322 & n18362 ) ;
  assign n18364 = x1154 | n18262 ;
  assign n18365 = x618 | x778 ;
  assign n18366 = ( x618 & n15081 ) | ( x618 & n18365 ) | ( n15081 & n18365 ) ;
  assign n18367 = ~n18364 & n18366 ;
  assign n18368 = ( n18259 & n18364 ) | ( n18259 & ~n18367 ) | ( n18364 & ~n18367 ) ;
  assign n18369 = x627 & n18368 ;
  assign n18370 = ~x618 & n18262 ;
  assign n18371 = x1154 & ~n18370 ;
  assign n18372 = ( n18246 & ~n18288 ) | ( n18246 & n18371 ) | ( ~n18288 & n18371 ) ;
  assign n18373 = n18369 & ~n18372 ;
  assign n18374 = x618 & n18361 ;
  assign n18375 = ( n18369 & n18373 ) | ( n18369 & n18374 ) | ( n18373 & n18374 ) ;
  assign n18376 = n18363 | n18375 ;
  assign n18377 = ~x781 & n18361 ;
  assign n18378 = x781 | n18377 ;
  assign n18379 = ( n18376 & n18377 ) | ( n18376 & n18378 ) | ( n18377 & n18378 ) ;
  assign n18380 = x619 & n18379 ;
  assign n18381 = ( n18307 & n18312 ) | ( n18307 & n18380 ) | ( n18312 & n18380 ) ;
  assign n18382 = x619 & ~x778 ;
  assign n18383 = ( x619 & ~n15081 ) | ( x619 & n18382 ) | ( ~n15081 & n18382 ) ;
  assign n18384 = ~n18249 & n18383 ;
  assign n18385 = n18259 & n18384 ;
  assign n18386 = x1159 & ~n18262 ;
  assign n18387 = x648 | n18386 ;
  assign n18388 = ( x648 & ~n18385 ) | ( x648 & n18387 ) | ( ~n18385 & n18387 ) ;
  assign n18389 = x619 & ~n18275 ;
  assign n18390 = x619 & n18262 ;
  assign n18391 = ( n18288 & n18389 ) | ( n18288 & n18390 ) | ( n18389 & n18390 ) ;
  assign n18392 = x1159 | n18391 ;
  assign n18393 = ~x619 & n18379 ;
  assign n18394 = n18388 | n18393 ;
  assign n18395 = n18392 | n18394 ;
  assign n18396 = ( x789 & n18388 ) | ( x789 & ~n18395 ) | ( n18388 & ~n18395 ) ;
  assign n18397 = ~n18381 & n18396 ;
  assign n18398 = x789 | n18379 ;
  assign n18399 = ~n16177 & n18398 ;
  assign n18400 = n18300 | n18399 ;
  assign n18401 = ( n18300 & ~n18397 ) | ( n18300 & n18400 ) | ( ~n18397 & n18400 ) ;
  assign n18402 = x630 & ~n15134 ;
  assign n18403 = x1157 & ~n18402 ;
  assign n18404 = ( x1157 & ~n18261 ) | ( x1157 & n18403 ) | ( ~n18261 & n18403 ) ;
  assign n18405 = ~n17215 & n18287 ;
  assign n18406 = ~x630 & n18405 ;
  assign n18407 = ~n17220 & n18406 ;
  assign n18408 = ( x630 & x647 ) | ( x630 & n18407 ) | ( x647 & n18407 ) ;
  assign n18409 = n18404 & ~n18408 ;
  assign n18410 = x630 & n17220 ;
  assign n18411 = ( x630 & ~n18405 ) | ( x630 & n18410 ) | ( ~n18405 & n18410 ) ;
  assign n18412 = x630 | n15134 ;
  assign n18413 = ( n17387 & ~n18261 ) | ( n17387 & n18412 ) | ( ~n18261 & n18412 ) ;
  assign n18414 = n17387 & n18413 ;
  assign n18415 = ( ~x1157 & n18411 ) | ( ~x1157 & n18414 ) | ( n18411 & n18414 ) ;
  assign n18416 = n18409 | n18415 ;
  assign n18417 = x787 & ~n18262 ;
  assign n18418 = n18416 & n18417 ;
  assign n18419 = x628 & n18405 ;
  assign n18420 = x628 & x629 ;
  assign n18421 = x1156 & ~n18420 ;
  assign n18422 = ( n15131 & ~n18261 ) | ( n15131 & n18421 ) | ( ~n18261 & n18421 ) ;
  assign n18423 = ~n18419 & n18422 ;
  assign n18424 = ( x629 & ~n18405 ) | ( x629 & n18420 ) | ( ~n18405 & n18420 ) ;
  assign n18425 = x628 & ~n18261 ;
  assign n18426 = ~x1156 & n18425 ;
  assign n18427 = ( ~x1156 & n18424 ) | ( ~x1156 & n18426 ) | ( n18424 & n18426 ) ;
  assign n18428 = n18423 | n18427 ;
  assign n18429 = x792 & ~n18262 ;
  assign n18430 = n18428 & n18429 ;
  assign n18431 = ( x787 & n15141 ) | ( x787 & n17388 ) | ( n15141 & n17388 ) ;
  assign n18432 = ( x629 & ~x792 ) | ( x629 & n17218 ) | ( ~x792 & n17218 ) ;
  assign n18433 = ( x629 & x792 ) | ( x629 & n17217 ) | ( x792 & n17217 ) ;
  assign n18434 = ~n18432 & n18433 ;
  assign n18435 = n18428 & n18434 ;
  assign n18436 = ~n18262 & n18435 ;
  assign n18437 = ( n18431 & n18434 ) | ( n18431 & ~n18436 ) | ( n18434 & ~n18436 ) ;
  assign n18438 = ~n18418 & n18437 ;
  assign n18439 = ( n18418 & n18430 ) | ( n18418 & ~n18438 ) | ( n18430 & ~n18438 ) ;
  assign n18440 = x644 & ~n18439 ;
  assign n18441 = n17220 | n17389 ;
  assign n18442 = ~n18262 & n18441 ;
  assign n18443 = x644 | n18442 ;
  assign n18444 = ~x644 & n18262 ;
  assign n18445 = ( n18405 & ~n18443 ) | ( n18405 & n18444 ) | ( ~n18443 & n18444 ) ;
  assign n18446 = x715 & ~n18445 ;
  assign n18447 = ~n18440 & n18446 ;
  assign n18448 = x644 & n18438 ;
  assign n18449 = n18446 & ~n18448 ;
  assign n18450 = ( ~n18401 & n18447 ) | ( ~n18401 & n18449 ) | ( n18447 & n18449 ) ;
  assign n18451 = n18268 & ~n18450 ;
  assign n18452 = x715 & ~n18262 ;
  assign n18453 = x644 | n18264 ;
  assign n18454 = n18452 & n18453 ;
  assign n18455 = ( ~n18261 & n18452 ) | ( ~n18261 & n18454 ) | ( n18452 & n18454 ) ;
  assign n18456 = x1160 | n18455 ;
  assign n18457 = x644 | n18439 ;
  assign n18458 = x644 & ~n18442 ;
  assign n18459 = x644 & n18262 ;
  assign n18460 = ( n18405 & n18458 ) | ( n18405 & n18459 ) | ( n18458 & n18459 ) ;
  assign n18461 = x715 | n18460 ;
  assign n18462 = n18457 & ~n18461 ;
  assign n18463 = ~x644 & n18438 ;
  assign n18464 = n18461 | n18463 ;
  assign n18465 = ( n18401 & ~n18462 ) | ( n18401 & n18464 ) | ( ~n18462 & n18464 ) ;
  assign n18466 = ~n18456 & n18465 ;
  assign n18467 = n18451 | n18466 ;
  assign n18468 = x790 | n18439 ;
  assign n18469 = ~x790 & n18438 ;
  assign n18470 = ( n18401 & ~n18468 ) | ( n18401 & n18469 ) | ( ~n18468 & n18469 ) ;
  assign n18471 = x832 & ~n18470 ;
  assign n18472 = ~x790 & n18471 ;
  assign n18473 = ( ~n18467 & n18471 ) | ( ~n18467 & n18472 ) | ( n18471 & n18472 ) ;
  assign n18474 = x57 & x144 ;
  assign n18475 = x832 | n18474 ;
  assign n18476 = ~n18473 & n18475 ;
  assign n18477 = ( n18245 & ~n18473 ) | ( n18245 & n18476 ) | ( ~n18473 & n18476 ) ;
  assign n18478 = x145 | n14834 ;
  assign n18479 = n15414 & n18478 ;
  assign n18480 = x698 | n2032 ;
  assign n18481 = ~n18478 & n18480 ;
  assign n18482 = x145 & n16323 ;
  assign n18483 = x38 | n18482 ;
  assign n18484 = ~n2032 & n18483 ;
  assign n18485 = x145 | n16319 ;
  assign n18486 = ~n18484 & n18485 ;
  assign n18487 = x145 | n15070 ;
  assign n18488 = n15375 & n18487 ;
  assign n18489 = x698 | n18488 ;
  assign n18490 = n18486 | n18489 ;
  assign n18491 = ~n18481 & n18490 ;
  assign n18492 = ~x778 & n18491 ;
  assign n18493 = ( x625 & x1153 ) | ( x625 & n18478 ) | ( x1153 & n18478 ) ;
  assign n18494 = ( ~x625 & x1153 ) | ( ~x625 & n18491 ) | ( x1153 & n18491 ) ;
  assign n18495 = n18493 & n18494 ;
  assign n18496 = ( x625 & x1153 ) | ( x625 & ~n18478 ) | ( x1153 & ~n18478 ) ;
  assign n18497 = ( x625 & ~x1153 ) | ( x625 & n18491 ) | ( ~x1153 & n18491 ) ;
  assign n18498 = ~n18496 & n18497 ;
  assign n18499 = n18495 | n18498 ;
  assign n18500 = x778 & n18499 ;
  assign n18501 = n18492 | n18500 ;
  assign n18502 = ~n15400 & n18501 ;
  assign n18503 = n15400 & n18478 ;
  assign n18504 = n18502 | n18503 ;
  assign n18505 = n15407 | n18504 ;
  assign n18506 = n15407 & ~n18478 ;
  assign n18507 = n18505 & ~n18506 ;
  assign n18508 = ~n15414 & n18507 ;
  assign n18509 = n18479 | n18508 ;
  assign n18510 = n15421 | n18509 ;
  assign n18511 = n15421 & ~n18478 ;
  assign n18512 = n18510 & ~n18511 ;
  assign n18513 = ~x792 & n18512 ;
  assign n18514 = ( x628 & x1156 ) | ( x628 & n18478 ) | ( x1156 & n18478 ) ;
  assign n18515 = ( ~x628 & x1156 ) | ( ~x628 & n18512 ) | ( x1156 & n18512 ) ;
  assign n18516 = n18514 & n18515 ;
  assign n18517 = ( x628 & x1156 ) | ( x628 & ~n18478 ) | ( x1156 & ~n18478 ) ;
  assign n18518 = ( x628 & ~x1156 ) | ( x628 & n18512 ) | ( ~x1156 & n18512 ) ;
  assign n18519 = ~n18517 & n18518 ;
  assign n18520 = n18516 | n18519 ;
  assign n18521 = x792 & n18520 ;
  assign n18522 = n18513 | n18521 ;
  assign n18523 = x787 | n18522 ;
  assign n18524 = x647 & n18522 ;
  assign n18525 = ~x647 & n18478 ;
  assign n18526 = n18524 | n18525 ;
  assign n18527 = ( ~x787 & x1157 ) | ( ~x787 & n18526 ) | ( x1157 & n18526 ) ;
  assign n18528 = ~x647 & n18522 ;
  assign n18529 = x647 & n18478 ;
  assign n18530 = n18528 | n18529 ;
  assign n18531 = ( x787 & x1157 ) | ( x787 & ~n18530 ) | ( x1157 & ~n18530 ) ;
  assign n18532 = ~n18527 & n18531 ;
  assign n18533 = n18523 & ~n18532 ;
  assign n18534 = x644 | n18533 ;
  assign n18535 = x715 & n18534 ;
  assign n18536 = x145 & n2032 ;
  assign n18537 = x145 | n14936 ;
  assign n18538 = x767 & n18537 ;
  assign n18539 = x145 & ~n14933 ;
  assign n18540 = x145 | x767 ;
  assign n18541 = n15063 & ~n18540 ;
  assign n18542 = n18539 | n18541 ;
  assign n18543 = n18538 | n18542 ;
  assign n18544 = ~x38 & n18543 ;
  assign n18545 = ~x767 & n15072 ;
  assign n18546 = x38 & n18487 ;
  assign n18547 = ~n18545 & n18546 ;
  assign n18548 = n18544 | n18547 ;
  assign n18549 = ~n2032 & n18548 ;
  assign n18550 = n18536 | n18549 ;
  assign n18551 = ~n15082 & n18550 ;
  assign n18552 = n15082 & n18478 ;
  assign n18553 = n18551 | n18552 ;
  assign n18554 = ~x785 & n18553 ;
  assign n18555 = ~n15088 & n18478 ;
  assign n18556 = x609 & n18551 ;
  assign n18557 = n18555 | n18556 ;
  assign n18558 = x1155 & n18557 ;
  assign n18559 = n15094 & n18478 ;
  assign n18560 = ~x609 & n18551 ;
  assign n18561 = n18559 | n18560 ;
  assign n18562 = ~x1155 & n18561 ;
  assign n18563 = n18558 | n18562 ;
  assign n18564 = x785 & n18563 ;
  assign n18565 = n18554 | n18564 ;
  assign n18566 = ~x781 & n18565 ;
  assign n18567 = ( x618 & x1154 ) | ( x618 & n18478 ) | ( x1154 & n18478 ) ;
  assign n18568 = ( ~x618 & x1154 ) | ( ~x618 & n18565 ) | ( x1154 & n18565 ) ;
  assign n18569 = n18567 & n18568 ;
  assign n18570 = ( x618 & x1154 ) | ( x618 & ~n18478 ) | ( x1154 & ~n18478 ) ;
  assign n18571 = ( x618 & ~x1154 ) | ( x618 & n18565 ) | ( ~x1154 & n18565 ) ;
  assign n18572 = ~n18570 & n18571 ;
  assign n18573 = n18569 | n18572 ;
  assign n18574 = x781 & n18573 ;
  assign n18575 = n18566 | n18574 ;
  assign n18576 = ~x789 & n18575 ;
  assign n18577 = ( x619 & x1159 ) | ( x619 & n18478 ) | ( x1159 & n18478 ) ;
  assign n18578 = ( ~x619 & x1159 ) | ( ~x619 & n18575 ) | ( x1159 & n18575 ) ;
  assign n18579 = n18577 & n18578 ;
  assign n18580 = ( x619 & x1159 ) | ( x619 & ~n18478 ) | ( x1159 & ~n18478 ) ;
  assign n18581 = ( x619 & ~x1159 ) | ( x619 & n18575 ) | ( ~x1159 & n18575 ) ;
  assign n18582 = ~n18580 & n18581 ;
  assign n18583 = n18579 | n18582 ;
  assign n18584 = x789 & n18583 ;
  assign n18585 = n18576 | n18584 ;
  assign n18586 = ~x788 & n18585 ;
  assign n18587 = ( x626 & x1158 ) | ( x626 & n18478 ) | ( x1158 & n18478 ) ;
  assign n18588 = ( ~x1158 & n18585 ) | ( ~x1158 & n18587 ) | ( n18585 & n18587 ) ;
  assign n18589 = ( ~x626 & n18587 ) | ( ~x626 & n18588 ) | ( n18587 & n18588 ) ;
  assign n18590 = x788 & n18589 ;
  assign n18591 = n18586 | n18590 ;
  assign n18592 = n15134 | n18591 ;
  assign n18593 = n15134 & ~n18478 ;
  assign n18594 = n18592 & ~n18593 ;
  assign n18595 = n15141 | n18594 ;
  assign n18596 = n15141 & ~n18478 ;
  assign n18597 = n18595 & ~n18596 ;
  assign n18598 = ( x644 & x715 ) | ( x644 & ~n18597 ) | ( x715 & ~n18597 ) ;
  assign n18599 = ( x644 & ~x715 ) | ( x644 & n18478 ) | ( ~x715 & n18478 ) ;
  assign n18600 = ~n18598 & n18599 ;
  assign n18601 = x1160 & ~n18600 ;
  assign n18602 = ~n18535 & n18601 ;
  assign n18603 = ( x644 & x715 ) | ( x644 & n18597 ) | ( x715 & n18597 ) ;
  assign n18604 = ( ~x644 & x715 ) | ( ~x644 & n18478 ) | ( x715 & n18478 ) ;
  assign n18605 = n18603 & n18604 ;
  assign n18606 = x1160 | n18605 ;
  assign n18607 = ( x644 & x715 ) | ( x644 & ~n18533 ) | ( x715 & ~n18533 ) ;
  assign n18608 = x630 & n17386 ;
  assign n18609 = ~x630 & n17387 ;
  assign n18610 = n18608 | n18609 ;
  assign n18611 = n18594 & n18610 ;
  assign n18612 = n15139 & n18530 ;
  assign n18613 = n15138 & n18526 ;
  assign n18614 = n18612 | n18613 ;
  assign n18615 = n18611 | n18614 ;
  assign n18616 = x787 & n18615 ;
  assign n18617 = ~x628 & x629 ;
  assign n18618 = x1156 & n18617 ;
  assign n18619 = x628 & ~x629 ;
  assign n18620 = ~x1156 & n18619 ;
  assign n18621 = n18618 | n18620 ;
  assign n18622 = n18591 & n18621 ;
  assign n18623 = ( x629 & n18519 ) | ( x629 & n18622 ) | ( n18519 & n18622 ) ;
  assign n18624 = ( ~x629 & n18516 ) | ( ~x629 & n18622 ) | ( n18516 & n18622 ) ;
  assign n18625 = n18623 | n18624 ;
  assign n18626 = x792 & n18625 ;
  assign n18627 = x648 & ~n18582 ;
  assign n18628 = ( x619 & x1159 ) | ( x619 & n18507 ) | ( x1159 & n18507 ) ;
  assign n18629 = x627 | n18569 ;
  assign n18630 = ( x618 & x1154 ) | ( x618 & ~n18504 ) | ( x1154 & ~n18504 ) ;
  assign n18631 = x660 | n18558 ;
  assign n18632 = ( x609 & x1155 ) | ( x609 & ~n18501 ) | ( x1155 & ~n18501 ) ;
  assign n18633 = x608 | n18495 ;
  assign n18634 = ( x625 & x1153 ) | ( x625 & ~n18550 ) | ( x1153 & ~n18550 ) ;
  assign n18635 = x698 & ~n18548 ;
  assign n18636 = ( x145 & ~x767 ) | ( x145 & n15797 ) | ( ~x767 & n15797 ) ;
  assign n18637 = ( x145 & x767 ) | ( x145 & n15872 ) | ( x767 & n15872 ) ;
  assign n18638 = n18636 & ~n18637 ;
  assign n18639 = x39 & ~n18638 ;
  assign n18640 = ( x145 & ~x767 ) | ( x145 & n15583 ) | ( ~x767 & n15583 ) ;
  assign n18641 = ( x145 & x767 ) | ( x145 & n15699 ) | ( x767 & n15699 ) ;
  assign n18642 = ~n18640 & n18641 ;
  assign n18643 = n18639 & ~n18642 ;
  assign n18644 = ( ~x145 & x767 ) | ( ~x145 & n15887 ) | ( x767 & n15887 ) ;
  assign n18645 = ( x145 & x767 ) | ( x145 & ~n15891 ) | ( x767 & ~n15891 ) ;
  assign n18646 = n18644 & n18645 ;
  assign n18647 = ( ~x145 & x767 ) | ( ~x145 & n15894 ) | ( x767 & n15894 ) ;
  assign n18648 = ( x145 & x767 ) | ( x145 & ~n15897 ) | ( x767 & ~n15897 ) ;
  assign n18649 = n18647 | n18648 ;
  assign n18650 = ~n18646 & n18649 ;
  assign n18651 = x39 | n18650 ;
  assign n18652 = ~x38 & n18651 ;
  assign n18653 = ~n18643 & n18652 ;
  assign n18654 = x767 | n15758 ;
  assign n18655 = n17573 & n18654 ;
  assign n18656 = x145 | n18655 ;
  assign n18657 = ~x767 & n14840 ;
  assign n18658 = n15529 | n18657 ;
  assign n18659 = x145 & n18658 ;
  assign n18660 = ~n4810 & n18659 ;
  assign n18661 = x38 & ~n18660 ;
  assign n18662 = n18656 & n18661 ;
  assign n18663 = x698 | n18662 ;
  assign n18664 = n18653 | n18663 ;
  assign n18665 = ~n2032 & n18664 ;
  assign n18666 = ~n18635 & n18665 ;
  assign n18667 = n18536 | n18666 ;
  assign n18668 = ( x625 & ~x1153 ) | ( x625 & n18667 ) | ( ~x1153 & n18667 ) ;
  assign n18669 = ~n18634 & n18668 ;
  assign n18670 = n18633 | n18669 ;
  assign n18671 = x608 & ~n18498 ;
  assign n18672 = ( x625 & x1153 ) | ( x625 & n18550 ) | ( x1153 & n18550 ) ;
  assign n18673 = ( ~x625 & x1153 ) | ( ~x625 & n18667 ) | ( x1153 & n18667 ) ;
  assign n18674 = n18672 & n18673 ;
  assign n18675 = n18671 & ~n18674 ;
  assign n18676 = n18670 & ~n18675 ;
  assign n18677 = x778 & ~n18676 ;
  assign n18678 = x778 | n18667 ;
  assign n18679 = ~n18677 & n18678 ;
  assign n18680 = ( x609 & ~x1155 ) | ( x609 & n18679 ) | ( ~x1155 & n18679 ) ;
  assign n18681 = ~n18632 & n18680 ;
  assign n18682 = n18631 | n18681 ;
  assign n18683 = x660 & ~n18562 ;
  assign n18684 = ( x609 & x1155 ) | ( x609 & n18501 ) | ( x1155 & n18501 ) ;
  assign n18685 = ( ~x609 & x1155 ) | ( ~x609 & n18679 ) | ( x1155 & n18679 ) ;
  assign n18686 = n18684 & n18685 ;
  assign n18687 = n18683 & ~n18686 ;
  assign n18688 = n18682 & ~n18687 ;
  assign n18689 = x785 & ~n18688 ;
  assign n18690 = x785 | n18679 ;
  assign n18691 = ~n18689 & n18690 ;
  assign n18692 = ( x618 & ~x1154 ) | ( x618 & n18691 ) | ( ~x1154 & n18691 ) ;
  assign n18693 = ~n18630 & n18692 ;
  assign n18694 = n18629 | n18693 ;
  assign n18695 = x627 & ~n18572 ;
  assign n18696 = ( x618 & x1154 ) | ( x618 & n18504 ) | ( x1154 & n18504 ) ;
  assign n18697 = ( ~x618 & x1154 ) | ( ~x618 & n18691 ) | ( x1154 & n18691 ) ;
  assign n18698 = n18696 & n18697 ;
  assign n18699 = n18695 & ~n18698 ;
  assign n18700 = n18694 & ~n18699 ;
  assign n18701 = x781 & ~n18700 ;
  assign n18702 = x781 | n18691 ;
  assign n18703 = ~n18701 & n18702 ;
  assign n18704 = ( ~x619 & x1159 ) | ( ~x619 & n18703 ) | ( x1159 & n18703 ) ;
  assign n18705 = n18628 & n18704 ;
  assign n18706 = n18627 & ~n18705 ;
  assign n18707 = x648 | n18579 ;
  assign n18708 = ( x619 & x1159 ) | ( x619 & ~n18507 ) | ( x1159 & ~n18507 ) ;
  assign n18709 = ( x619 & ~x1159 ) | ( x619 & n18703 ) | ( ~x1159 & n18703 ) ;
  assign n18710 = ~n18708 & n18709 ;
  assign n18711 = n18707 | n18710 ;
  assign n18712 = x789 & n18711 ;
  assign n18713 = ~n18706 & n18712 ;
  assign n18714 = ~x789 & n18703 ;
  assign n18715 = n16177 | n18714 ;
  assign n18716 = n18713 | n18715 ;
  assign n18717 = n16115 & ~n18509 ;
  assign n18718 = n15420 & ~n18589 ;
  assign n18719 = n18717 | n18718 ;
  assign n18720 = x788 & n18719 ;
  assign n18721 = n18434 | n18720 ;
  assign n18722 = n18716 & ~n18721 ;
  assign n18723 = n18626 | n18722 ;
  assign n18724 = ~n18431 & n18723 ;
  assign n18725 = n18616 | n18724 ;
  assign n18726 = ( x644 & ~x715 ) | ( x644 & n18725 ) | ( ~x715 & n18725 ) ;
  assign n18727 = ~n18607 & n18726 ;
  assign n18728 = n18606 | n18727 ;
  assign n18729 = ~n18602 & n18728 ;
  assign n18730 = x790 & ~n18729 ;
  assign n18731 = x644 & n18601 ;
  assign n18732 = x790 & ~n18731 ;
  assign n18733 = n18725 | n18732 ;
  assign n18734 = ~n18730 & n18733 ;
  assign n18735 = ( ~x832 & n6785 ) | ( ~x832 & n18734 ) | ( n6785 & n18734 ) ;
  assign n18736 = ( ~x145 & x832 ) | ( ~x145 & n6785 ) | ( x832 & n6785 ) ;
  assign n18737 = n18735 & ~n18736 ;
  assign n18738 = x145 | n1290 ;
  assign n18739 = ~n18657 & n18738 ;
  assign n18740 = n16060 | n18739 ;
  assign n18741 = ~x785 & n18740 ;
  assign n18742 = n16065 | n18739 ;
  assign n18743 = x1155 & n18742 ;
  assign n18744 = n16068 | n18740 ;
  assign n18745 = ~x1155 & n18744 ;
  assign n18746 = n18743 | n18745 ;
  assign n18747 = x785 & n18746 ;
  assign n18748 = n18741 | n18747 ;
  assign n18749 = ~x781 & n18748 ;
  assign n18750 = n16075 | n18748 ;
  assign n18751 = x1154 & n18750 ;
  assign n18752 = n16078 | n18748 ;
  assign n18753 = ~x1154 & n18752 ;
  assign n18754 = n18751 | n18753 ;
  assign n18755 = x781 & n18754 ;
  assign n18756 = n18749 | n18755 ;
  assign n18757 = ~x789 & n18756 ;
  assign n18758 = ( x619 & x1159 ) | ( x619 & n18738 ) | ( x1159 & n18738 ) ;
  assign n18759 = ( ~x619 & x1159 ) | ( ~x619 & n18756 ) | ( x1159 & n18756 ) ;
  assign n18760 = n18758 & n18759 ;
  assign n18761 = ( x619 & x1159 ) | ( x619 & ~n18738 ) | ( x1159 & ~n18738 ) ;
  assign n18762 = ( x619 & ~x1159 ) | ( x619 & n18756 ) | ( ~x1159 & n18756 ) ;
  assign n18763 = ~n18761 & n18762 ;
  assign n18764 = n18760 | n18763 ;
  assign n18765 = x789 & n18764 ;
  assign n18766 = n18757 | n18765 ;
  assign n18767 = ~x788 & n18766 ;
  assign n18768 = ( x626 & x1158 ) | ( x626 & n18738 ) | ( x1158 & n18738 ) ;
  assign n18769 = ( ~x1158 & n18766 ) | ( ~x1158 & n18768 ) | ( n18766 & n18768 ) ;
  assign n18770 = ( ~x626 & n18768 ) | ( ~x626 & n18769 ) | ( n18768 & n18769 ) ;
  assign n18771 = x788 & n18770 ;
  assign n18772 = n18767 | n18771 ;
  assign n18773 = n15134 | n18772 ;
  assign n18774 = n15134 & ~n18738 ;
  assign n18775 = n18773 & ~n18774 ;
  assign n18776 = n18610 & n18775 ;
  assign n18777 = ( x647 & x1157 ) | ( x647 & ~n18738 ) | ( x1157 & ~n18738 ) ;
  assign n18778 = ~x698 & n15202 ;
  assign n18779 = n18738 & ~n18778 ;
  assign n18780 = ~x778 & n18779 ;
  assign n18781 = ~x625 & n18778 ;
  assign n18782 = n18779 | n18781 ;
  assign n18783 = x1153 & n18782 ;
  assign n18784 = ~x1153 & n18738 ;
  assign n18785 = ~n18781 & n18784 ;
  assign n18786 = n18783 | n18785 ;
  assign n18787 = x778 & n18786 ;
  assign n18788 = n18780 | n18787 ;
  assign n18789 = n16043 | n18788 ;
  assign n18790 = n16045 | n18789 ;
  assign n18791 = n16047 | n18790 ;
  assign n18792 = n16049 | n18791 ;
  assign n18793 = n16055 | n18792 ;
  assign n18794 = ( x647 & ~x1157 ) | ( x647 & n18793 ) | ( ~x1157 & n18793 ) ;
  assign n18795 = ~n18777 & n18794 ;
  assign n18796 = x630 & n18795 ;
  assign n18797 = x647 & n18793 ;
  assign n18798 = ~x647 & n18738 ;
  assign n18799 = n18797 | n18798 ;
  assign n18800 = n15138 & n18799 ;
  assign n18801 = n18796 | n18800 ;
  assign n18802 = n18776 | n18801 ;
  assign n18803 = x787 & n18802 ;
  assign n18804 = n16115 & ~n18791 ;
  assign n18805 = n15420 & ~n18770 ;
  assign n18806 = n18804 | n18805 ;
  assign n18807 = x788 & n18806 ;
  assign n18808 = x648 & ~n18763 ;
  assign n18809 = ( x619 & x1159 ) | ( x619 & n18790 ) | ( x1159 & n18790 ) ;
  assign n18810 = x627 | n18751 ;
  assign n18811 = ( x618 & x1154 ) | ( x618 & ~n18789 ) | ( x1154 & ~n18789 ) ;
  assign n18812 = x660 | n18743 ;
  assign n18813 = ( x609 & x1155 ) | ( x609 & ~n18788 ) | ( x1155 & ~n18788 ) ;
  assign n18814 = n14839 | n18779 ;
  assign n18815 = x625 & ~n18814 ;
  assign n18816 = n18739 & n18814 ;
  assign n18817 = n18815 | n18816 ;
  assign n18818 = n18784 & n18817 ;
  assign n18819 = x608 | n18783 ;
  assign n18820 = n18818 | n18819 ;
  assign n18821 = x1153 & n18739 ;
  assign n18822 = ~n18815 & n18821 ;
  assign n18823 = x608 & ~n18785 ;
  assign n18824 = ~n18822 & n18823 ;
  assign n18825 = n18820 & ~n18824 ;
  assign n18826 = x778 & ~n18825 ;
  assign n18827 = x778 | n18816 ;
  assign n18828 = ~n18826 & n18827 ;
  assign n18829 = ( x609 & ~x1155 ) | ( x609 & n18828 ) | ( ~x1155 & n18828 ) ;
  assign n18830 = ~n18813 & n18829 ;
  assign n18831 = n18812 | n18830 ;
  assign n18832 = x660 & ~n18745 ;
  assign n18833 = ( x609 & x1155 ) | ( x609 & n18788 ) | ( x1155 & n18788 ) ;
  assign n18834 = ( ~x609 & x1155 ) | ( ~x609 & n18828 ) | ( x1155 & n18828 ) ;
  assign n18835 = n18833 & n18834 ;
  assign n18836 = n18832 & ~n18835 ;
  assign n18837 = n18831 & ~n18836 ;
  assign n18838 = x785 & ~n18837 ;
  assign n18839 = x785 | n18828 ;
  assign n18840 = ~n18838 & n18839 ;
  assign n18841 = ( x618 & ~x1154 ) | ( x618 & n18840 ) | ( ~x1154 & n18840 ) ;
  assign n18842 = ~n18811 & n18841 ;
  assign n18843 = n18810 | n18842 ;
  assign n18844 = x627 & ~n18753 ;
  assign n18845 = ( x618 & x1154 ) | ( x618 & n18789 ) | ( x1154 & n18789 ) ;
  assign n18846 = ( ~x618 & x1154 ) | ( ~x618 & n18840 ) | ( x1154 & n18840 ) ;
  assign n18847 = n18845 & n18846 ;
  assign n18848 = n18844 & ~n18847 ;
  assign n18849 = n18843 & ~n18848 ;
  assign n18850 = x781 & ~n18849 ;
  assign n18851 = x781 | n18840 ;
  assign n18852 = ~n18850 & n18851 ;
  assign n18853 = ( ~x619 & x1159 ) | ( ~x619 & n18852 ) | ( x1159 & n18852 ) ;
  assign n18854 = n18809 & n18853 ;
  assign n18855 = n18808 & ~n18854 ;
  assign n18856 = x648 | n18760 ;
  assign n18857 = ( x619 & x1159 ) | ( x619 & ~n18790 ) | ( x1159 & ~n18790 ) ;
  assign n18858 = ( x619 & ~x1159 ) | ( x619 & n18852 ) | ( ~x1159 & n18852 ) ;
  assign n18859 = ~n18857 & n18858 ;
  assign n18860 = n18856 | n18859 ;
  assign n18861 = x789 & n18860 ;
  assign n18862 = ~n18855 & n18861 ;
  assign n18863 = ~x789 & n18852 ;
  assign n18864 = n16177 | n18863 ;
  assign n18865 = n18862 | n18864 ;
  assign n18866 = ~n18807 & n18865 ;
  assign n18867 = n18434 | n18866 ;
  assign n18868 = n16650 | n18792 ;
  assign n18869 = n16051 & ~n18772 ;
  assign n18870 = n18868 & ~n18869 ;
  assign n18871 = ( x629 & ~x792 ) | ( x629 & n18870 ) | ( ~x792 & n18870 ) ;
  assign n18872 = n16052 & ~n18772 ;
  assign n18873 = n16643 & ~n18792 ;
  assign n18874 = n18872 | n18873 ;
  assign n18875 = ( x629 & x792 ) | ( x629 & n18874 ) | ( x792 & n18874 ) ;
  assign n18876 = ~n18871 & n18875 ;
  assign n18877 = n18431 | n18876 ;
  assign n18878 = n18867 & ~n18877 ;
  assign n18879 = n18803 | n18878 ;
  assign n18880 = ( x790 & x832 ) | ( x790 & n18879 ) | ( x832 & n18879 ) ;
  assign n18881 = n15141 | n18775 ;
  assign n18882 = n15141 & ~n18738 ;
  assign n18883 = n18881 & ~n18882 ;
  assign n18884 = ( x644 & x715 ) | ( x644 & ~n18883 ) | ( x715 & ~n18883 ) ;
  assign n18885 = ( x644 & ~x715 ) | ( x644 & n18738 ) | ( ~x715 & n18738 ) ;
  assign n18886 = ~n18884 & n18885 ;
  assign n18887 = x1160 & ~n18886 ;
  assign n18888 = ~x787 & n18793 ;
  assign n18889 = x1157 & n18799 ;
  assign n18890 = n18795 | n18889 ;
  assign n18891 = x787 & n18890 ;
  assign n18892 = n18888 | n18891 ;
  assign n18893 = ( x644 & x715 ) | ( x644 & n18892 ) | ( x715 & n18892 ) ;
  assign n18894 = ( ~x644 & x715 ) | ( ~x644 & n18879 ) | ( x715 & n18879 ) ;
  assign n18895 = n18893 & n18894 ;
  assign n18896 = n18887 & ~n18895 ;
  assign n18897 = ( x644 & x715 ) | ( x644 & n18883 ) | ( x715 & n18883 ) ;
  assign n18898 = ( ~x644 & x715 ) | ( ~x644 & n18738 ) | ( x715 & n18738 ) ;
  assign n18899 = n18897 & n18898 ;
  assign n18900 = x1160 | n18899 ;
  assign n18901 = ( x644 & x715 ) | ( x644 & ~n18892 ) | ( x715 & ~n18892 ) ;
  assign n18902 = ( x644 & ~x715 ) | ( x644 & n18879 ) | ( ~x715 & n18879 ) ;
  assign n18903 = ~n18901 & n18902 ;
  assign n18904 = n18900 | n18903 ;
  assign n18905 = ~n18896 & n18904 ;
  assign n18906 = ( ~x790 & x832 ) | ( ~x790 & n18905 ) | ( x832 & n18905 ) ;
  assign n18907 = n18880 & n18906 ;
  assign n18908 = n18737 | n18907 ;
  assign n18909 = n4718 & n14528 ;
  assign n18910 = n14575 | n18909 ;
  assign n18911 = x146 & ~n18910 ;
  assign n18912 = x743 & x947 ;
  assign n18913 = x907 & ~x947 ;
  assign n18914 = x735 & n18913 ;
  assign n18915 = n18912 | n18914 ;
  assign n18916 = n14528 & n18915 ;
  assign n18917 = x215 & ~n18916 ;
  assign n18918 = ~n18911 & n18917 ;
  assign n18919 = x907 | n14450 ;
  assign n18920 = x146 & ~n16709 ;
  assign n18921 = n18919 & n18920 ;
  assign n18922 = x146 & ~n16712 ;
  assign n18923 = ~n18919 & n18922 ;
  assign n18924 = x735 & x907 ;
  assign n18925 = x947 | n16709 ;
  assign n18926 = ( x947 & n18924 ) | ( x947 & n18925 ) | ( n18924 & n18925 ) ;
  assign n18927 = n18923 | n18926 ;
  assign n18928 = x743 & n16709 ;
  assign n18929 = x947 & ~n18920 ;
  assign n18930 = ~n18928 & n18929 ;
  assign n18931 = n18927 & ~n18930 ;
  assign n18932 = n18921 | n18931 ;
  assign n18933 = ( x215 & n2203 ) | ( x215 & n18932 ) | ( n2203 & n18932 ) ;
  assign n18934 = n16705 & n18915 ;
  assign n18935 = x146 & ~n16705 ;
  assign n18936 = n18934 | n18935 ;
  assign n18937 = ( x215 & ~n2203 ) | ( x215 & n18936 ) | ( ~n2203 & n18936 ) ;
  assign n18938 = n18933 | n18937 ;
  assign n18939 = ~n18918 & n18938 ;
  assign n18940 = x299 & ~n18939 ;
  assign n18941 = n16709 & n18915 ;
  assign n18942 = n4764 & ~n18920 ;
  assign n18943 = ~n18941 & n18942 ;
  assign n18944 = n16712 & n18915 ;
  assign n18945 = n4764 | n18922 ;
  assign n18946 = n18944 | n18945 ;
  assign n18947 = ~n18943 & n18946 ;
  assign n18948 = n1823 & ~n18947 ;
  assign n18949 = ( ~x223 & n15629 ) | ( ~x223 & n18936 ) | ( n15629 & n18936 ) ;
  assign n18950 = ~n18948 & n18949 ;
  assign n18951 = x146 & ~n14528 ;
  assign n18952 = n18916 | n18951 ;
  assign n18953 = n4764 & n18952 ;
  assign n18954 = ( x146 & ~n4764 ) | ( x146 & n16719 ) | ( ~n4764 & n16719 ) ;
  assign n18955 = ( n4764 & n16719 ) | ( n4764 & ~n18915 ) | ( n16719 & ~n18915 ) ;
  assign n18956 = n18954 & ~n18955 ;
  assign n18957 = n18953 | n18956 ;
  assign n18958 = x223 & n18957 ;
  assign n18959 = x299 | n18958 ;
  assign n18960 = n18950 | n18959 ;
  assign n18961 = ~n18940 & n18960 ;
  assign n18962 = x39 & ~n18961 ;
  assign n18963 = ( x146 & ~x299 ) | ( x146 & n14820 ) | ( ~x299 & n14820 ) ;
  assign n18964 = ( x299 & n14820 ) | ( x299 & ~n18915 ) | ( n14820 & ~n18915 ) ;
  assign n18965 = n18963 & ~n18964 ;
  assign n18966 = ( x146 & x299 ) | ( x146 & n14814 ) | ( x299 & n14814 ) ;
  assign n18967 = ( x299 & ~n14814 ) | ( x299 & n18915 ) | ( ~n14814 & n18915 ) ;
  assign n18968 = n18966 & n18967 ;
  assign n18969 = n18965 | n18968 ;
  assign n18970 = ( ~x38 & n9138 ) | ( ~x38 & n18969 ) | ( n9138 & n18969 ) ;
  assign n18971 = ~n18962 & n18970 ;
  assign n18972 = x146 | n15070 ;
  assign n18973 = n1290 & ~n18915 ;
  assign n18974 = ~n4810 & n18973 ;
  assign n18975 = x38 & ~n18974 ;
  assign n18976 = n18972 & n18975 ;
  assign n18977 = n8359 | n18976 ;
  assign n18978 = n18971 | n18977 ;
  assign n18979 = ~x146 & n8359 ;
  assign n18980 = x832 | n18979 ;
  assign n18981 = n18978 & ~n18980 ;
  assign n18982 = x146 | n1290 ;
  assign n18983 = x832 & n18982 ;
  assign n18984 = ~n18973 & n18983 ;
  assign n18985 = n18981 | n18984 ;
  assign n18986 = ~x947 & n14822 ;
  assign n18987 = x39 | n18986 ;
  assign n18988 = n14702 & ~n14707 ;
  assign n18989 = ~x299 & n18988 ;
  assign n18990 = x947 & n18989 ;
  assign n18991 = ~n14481 & n14685 ;
  assign n18992 = ~x947 & n18991 ;
  assign n18993 = n16709 & n18913 ;
  assign n18994 = n14682 | n18993 ;
  assign n18995 = n2203 & n18994 ;
  assign n18996 = x215 | n18995 ;
  assign n18997 = n18992 | n18996 ;
  assign n18998 = x215 & ~n14575 ;
  assign n18999 = n14528 & n18913 ;
  assign n19000 = n18998 & ~n18999 ;
  assign n19001 = n18997 & ~n19000 ;
  assign n19002 = x299 & ~n19001 ;
  assign n19003 = n14709 & ~n19002 ;
  assign n19004 = ~n18990 & n19003 ;
  assign n19005 = x39 & ~n19004 ;
  assign n19006 = n18987 & ~n19005 ;
  assign n19007 = ~x38 & n19006 ;
  assign n19008 = x38 & ~x947 ;
  assign n19009 = n14827 & n19008 ;
  assign n19010 = n19007 | n19009 ;
  assign n19011 = x770 | n19010 ;
  assign n19012 = x770 & ~n15382 ;
  assign n19013 = n19011 & ~n19012 ;
  assign n19014 = x147 | n19013 ;
  assign n19015 = n15380 | n19009 ;
  assign n19016 = x947 & n14822 ;
  assign n19017 = x39 | n19016 ;
  assign n19018 = x947 & n18988 ;
  assign n19019 = x299 | n19018 ;
  assign n19020 = x215 & x947 ;
  assign n19021 = n14528 & n19020 ;
  assign n19022 = x299 & ~n19021 ;
  assign n19023 = x947 & n16709 ;
  assign n19024 = n2203 & ~n19023 ;
  assign n19025 = x947 & n16705 ;
  assign n19026 = n2203 | n19025 ;
  assign n19027 = ~x215 & n19026 ;
  assign n19028 = ~n19024 & n19027 ;
  assign n19029 = n19022 & ~n19028 ;
  assign n19030 = n19019 & ~n19029 ;
  assign n19031 = x39 & ~n19030 ;
  assign n19032 = n19017 & ~n19031 ;
  assign n19033 = x38 | n19032 ;
  assign n19034 = ~n19015 & n19033 ;
  assign n19035 = x147 & ~x770 ;
  assign n19036 = n19034 & n19035 ;
  assign n19037 = x726 | n19036 ;
  assign n19038 = n19014 & ~n19037 ;
  assign n19039 = x147 | n15070 ;
  assign n19040 = n15070 & n18913 ;
  assign n19041 = x38 & ~n19040 ;
  assign n19042 = n19039 & n19041 ;
  assign n19043 = x770 & ~n19042 ;
  assign n19044 = ~n18913 & n18991 ;
  assign n19045 = n14682 | n19023 ;
  assign n19046 = n2203 & n19045 ;
  assign n19047 = x215 | n19046 ;
  assign n19048 = n19044 | n19047 ;
  assign n19049 = ~n18998 & n19048 ;
  assign n19050 = n19021 | n19049 ;
  assign n19051 = x299 & n19050 ;
  assign n19052 = ~n18913 & n18989 ;
  assign n19053 = n19051 | n19052 ;
  assign n19054 = x39 & n19053 ;
  assign n19055 = n14822 & ~n18913 ;
  assign n19056 = ~x39 & n19055 ;
  assign n19057 = n19054 | n19056 ;
  assign n19058 = ( ~x38 & x147 ) | ( ~x38 & n19057 ) | ( x147 & n19057 ) ;
  assign n19059 = x215 & ~n18999 ;
  assign n19060 = n2203 & ~n18993 ;
  assign n19061 = x907 & n16705 ;
  assign n19062 = ~x947 & n19061 ;
  assign n19063 = n2203 | n19062 ;
  assign n19064 = ~n19060 & n19063 ;
  assign n19065 = x215 | n19064 ;
  assign n19066 = ~n19059 & n19065 ;
  assign n19067 = x299 & ~n19066 ;
  assign n19068 = n18913 & n18988 ;
  assign n19069 = x299 | n19068 ;
  assign n19070 = ~n19067 & n19069 ;
  assign n19071 = x39 & ~n19070 ;
  assign n19072 = n14822 & n18913 ;
  assign n19073 = x39 | n19072 ;
  assign n19074 = ~n19071 & n19073 ;
  assign n19075 = ( x38 & x147 ) | ( x38 & n19074 ) | ( x147 & n19074 ) ;
  assign n19076 = n19058 & ~n19075 ;
  assign n19077 = n19043 & ~n19076 ;
  assign n19078 = ~n4718 & n14827 ;
  assign n19079 = x147 | n19078 ;
  assign n19080 = n4718 & n15070 ;
  assign n19081 = x38 & ~n19080 ;
  assign n19082 = n19079 & n19081 ;
  assign n19083 = x770 | n19082 ;
  assign n19084 = ~n14481 & n14699 ;
  assign n19085 = ~n1868 & n19084 ;
  assign n19086 = n14698 | n19085 ;
  assign n19087 = ~n4718 & n19086 ;
  assign n19088 = x223 | n19087 ;
  assign n19089 = ~n14703 & n14705 ;
  assign n19090 = ~x947 & n19089 ;
  assign n19091 = x223 & ~n19090 ;
  assign n19092 = ~n18913 & n19089 ;
  assign n19093 = x223 & ~n19092 ;
  assign n19094 = n19091 | n19093 ;
  assign n19095 = n19088 & ~n19094 ;
  assign n19096 = x299 | n19095 ;
  assign n19097 = x299 & x947 ;
  assign n19098 = ( x299 & ~n19049 ) | ( x299 & n19097 ) | ( ~n19049 & n19097 ) ;
  assign n19099 = n19096 & ~n19098 ;
  assign n19100 = x39 & n19099 ;
  assign n19101 = n4718 & n14822 ;
  assign n19102 = x39 | n19101 ;
  assign n19103 = n14822 & ~n19102 ;
  assign n19104 = n19100 | n19103 ;
  assign n19105 = ( ~x38 & x147 ) | ( ~x38 & n19104 ) | ( x147 & n19104 ) ;
  assign n19106 = n4718 & n18988 ;
  assign n19107 = ~x299 & n19106 ;
  assign n19108 = n2203 & n14684 ;
  assign n19109 = n4718 & n16705 ;
  assign n19110 = ( x215 & ~n14841 ) | ( x215 & n19109 ) | ( ~n14841 & n19109 ) ;
  assign n19111 = n19108 | n19110 ;
  assign n19112 = x299 & ~n14577 ;
  assign n19113 = n19111 & n19112 ;
  assign n19114 = n19107 | n19113 ;
  assign n19115 = x39 & ~n19114 ;
  assign n19116 = n19102 & ~n19115 ;
  assign n19117 = ( x38 & x147 ) | ( x38 & n19116 ) | ( x147 & n19116 ) ;
  assign n19118 = n19105 & ~n19117 ;
  assign n19119 = n19083 | n19118 ;
  assign n19120 = x726 & n19119 ;
  assign n19121 = ~n19077 & n19120 ;
  assign n19122 = n8359 | n19121 ;
  assign n19123 = n19038 | n19122 ;
  assign n19124 = ~x147 & n8359 ;
  assign n19125 = x832 | n19124 ;
  assign n19126 = n19123 & ~n19125 ;
  assign n19127 = ~x770 & x947 ;
  assign n19128 = x726 & n18913 ;
  assign n19129 = n19127 | n19128 ;
  assign n19130 = ( ~x832 & n1290 ) | ( ~x832 & n19129 ) | ( n1290 & n19129 ) ;
  assign n19131 = ( x147 & x832 ) | ( x147 & n1290 ) | ( x832 & n1290 ) ;
  assign n19132 = ~n19130 & n19131 ;
  assign n19133 = n19126 | n19132 ;
  assign n19134 = ~n7931 & n19053 ;
  assign n19135 = n14709 & ~n19067 ;
  assign n19136 = x148 & ~n19135 ;
  assign n19137 = x749 | n19136 ;
  assign n19138 = n19134 | n19137 ;
  assign n19139 = x39 & n19138 ;
  assign n19140 = ( ~x148 & x749 ) | ( ~x148 & n19114 ) | ( x749 & n19114 ) ;
  assign n19141 = ( x148 & x749 ) | ( x148 & ~n19099 ) | ( x749 & ~n19099 ) ;
  assign n19142 = n19140 & n19141 ;
  assign n19143 = n19139 & ~n19142 ;
  assign n19144 = x148 | n14822 ;
  assign n19145 = ~x39 & n19144 ;
  assign n19146 = ~x749 & x947 ;
  assign n19147 = n19101 & ~n19146 ;
  assign n19148 = n19145 & ~n19147 ;
  assign n19149 = x38 | n19148 ;
  assign n19150 = n19143 | n19149 ;
  assign n19151 = n19080 & ~n19146 ;
  assign n19152 = x148 | n15070 ;
  assign n19153 = ~n19151 & n19152 ;
  assign n19154 = x38 & ~n19153 ;
  assign n19155 = x706 & ~n19154 ;
  assign n19156 = n19150 & n19155 ;
  assign n19157 = n2032 | n4832 ;
  assign n19158 = x148 | n18988 ;
  assign n19159 = ~n19019 & n19158 ;
  assign n19160 = x749 & ~n19159 ;
  assign n19161 = n19021 | n19028 ;
  assign n19162 = ( x148 & ~x299 ) | ( x148 & n19161 ) | ( ~x299 & n19161 ) ;
  assign n19163 = ( x148 & x299 ) | ( x148 & n19001 ) | ( x299 & n19001 ) ;
  assign n19164 = ~n19162 & n19163 ;
  assign n19165 = n19160 & ~n19164 ;
  assign n19166 = x148 | x749 ;
  assign n19167 = n14710 | n19166 ;
  assign n19168 = x39 & n19167 ;
  assign n19169 = ~n19165 & n19168 ;
  assign n19170 = x749 & x947 ;
  assign n19171 = n14822 & n19170 ;
  assign n19172 = n19145 & ~n19171 ;
  assign n19173 = x38 | n19172 ;
  assign n19174 = n19169 | n19173 ;
  assign n19175 = x148 & ~n14827 ;
  assign n19176 = n15070 & ~n19170 ;
  assign n19177 = x38 & ~n19176 ;
  assign n19178 = ~n19175 & n19177 ;
  assign n19179 = x706 | n19178 ;
  assign n19180 = n19174 & ~n19179 ;
  assign n19181 = n19157 | n19180 ;
  assign n19182 = n19156 | n19181 ;
  assign n19183 = ~x148 & n19157 ;
  assign n19184 = x57 | n19183 ;
  assign n19185 = n19182 & ~n19184 ;
  assign n19186 = x57 & x148 ;
  assign n19187 = x832 | n19186 ;
  assign n19188 = n19185 | n19187 ;
  assign n19189 = x706 & n18913 ;
  assign n19190 = n1290 & ~n19170 ;
  assign n19191 = ~n19189 & n19190 ;
  assign n19192 = x148 & ~n1290 ;
  assign n19193 = x832 & ~n19192 ;
  assign n19194 = ~n19191 & n19193 ;
  assign n19195 = n19188 & ~n19194 ;
  assign n19196 = ~x755 & x947 ;
  assign n19197 = ~x725 & n18913 ;
  assign n19198 = n19196 | n19197 ;
  assign n19199 = ( ~x832 & n1290 ) | ( ~x832 & n19198 ) | ( n1290 & n19198 ) ;
  assign n19200 = ( x149 & x832 ) | ( x149 & n1290 ) | ( x832 & n1290 ) ;
  assign n19201 = ~n19199 & n19200 ;
  assign n19202 = x149 & ~n14827 ;
  assign n19203 = n15070 & ~n19196 ;
  assign n19204 = x38 & ~n19203 ;
  assign n19205 = ~n19202 & n19204 ;
  assign n19206 = x149 | n19001 ;
  assign n19207 = n13996 | n19029 ;
  assign n19208 = n19206 & n19207 ;
  assign n19209 = x149 | n18988 ;
  assign n19210 = ~n19019 & n19209 ;
  assign n19211 = x755 | n19210 ;
  assign n19212 = n19208 | n19211 ;
  assign n19213 = ~x149 & x755 ;
  assign n19214 = ~n14710 & n19213 ;
  assign n19215 = x39 & ~n19214 ;
  assign n19216 = n19212 & n19215 ;
  assign n19217 = ( x39 & n14822 ) | ( x39 & n19196 ) | ( n14822 & n19196 ) ;
  assign n19218 = ( ~x39 & x149 ) | ( ~x39 & n14822 ) | ( x149 & n14822 ) ;
  assign n19219 = ~n19217 & n19218 ;
  assign n19220 = x38 | n19219 ;
  assign n19221 = n19216 | n19220 ;
  assign n19222 = ~n19205 & n19221 ;
  assign n19223 = x725 & ~n19222 ;
  assign n19224 = ~n19072 & n19219 ;
  assign n19225 = x755 & ~n19052 ;
  assign n19226 = ( ~x149 & n19135 ) | ( ~x149 & n19225 ) | ( n19135 & n19225 ) ;
  assign n19227 = ( x149 & ~n19051 ) | ( x149 & n19225 ) | ( ~n19051 & n19225 ) ;
  assign n19228 = n19226 & n19227 ;
  assign n19229 = x39 & ~n19228 ;
  assign n19230 = ( ~x149 & x755 ) | ( ~x149 & n19099 ) | ( x755 & n19099 ) ;
  assign n19231 = ( x149 & x755 ) | ( x149 & ~n19114 ) | ( x755 & ~n19114 ) ;
  assign n19232 = n19230 | n19231 ;
  assign n19233 = n19229 & n19232 ;
  assign n19234 = n19224 | n19233 ;
  assign n19235 = ~x38 & n19234 ;
  assign n19236 = n4718 & n15756 ;
  assign n19237 = x755 & x947 ;
  assign n19238 = x39 | n19237 ;
  assign n19239 = n19236 & ~n19238 ;
  assign n19240 = x149 | n15070 ;
  assign n19241 = x38 & n19240 ;
  assign n19242 = ~n19239 & n19241 ;
  assign n19243 = x725 | n19242 ;
  assign n19244 = n19235 | n19243 ;
  assign n19245 = ~n19223 & n19244 ;
  assign n19246 = ( ~x832 & n8359 ) | ( ~x832 & n19245 ) | ( n8359 & n19245 ) ;
  assign n19247 = ( ~x149 & x832 ) | ( ~x149 & n8359 ) | ( x832 & n8359 ) ;
  assign n19248 = n19246 & ~n19247 ;
  assign n19249 = n19201 | n19248 ;
  assign n19250 = ~x150 & x751 ;
  assign n19251 = ~n14710 & n19250 ;
  assign n19252 = ( ~x150 & x751 ) | ( ~x150 & n19004 ) | ( x751 & n19004 ) ;
  assign n19253 = ( x150 & x751 ) | ( x150 & ~n19030 ) | ( x751 & ~n19030 ) ;
  assign n19254 = n19252 | n19253 ;
  assign n19255 = ~n19251 & n19254 ;
  assign n19256 = x39 & ~n19255 ;
  assign n19257 = x150 & ~n14822 ;
  assign n19258 = x751 & n14822 ;
  assign n19259 = n19257 | n19258 ;
  assign n19260 = n18987 | n19259 ;
  assign n19261 = ~x38 & n19260 ;
  assign n19262 = ~n19256 & n19261 ;
  assign n19263 = x150 & ~n14827 ;
  assign n19264 = ~x751 & x947 ;
  assign n19265 = n15070 & ~n19264 ;
  assign n19266 = n19263 | n19265 ;
  assign n19267 = x38 & n19266 ;
  assign n19268 = x701 & ~n19267 ;
  assign n19269 = ~n19262 & n19268 ;
  assign n19270 = ( ~x150 & x751 ) | ( ~x150 & n19070 ) | ( x751 & n19070 ) ;
  assign n19271 = ( x150 & x751 ) | ( x150 & ~n19053 ) | ( x751 & ~n19053 ) ;
  assign n19272 = n19270 & n19271 ;
  assign n19273 = ( ~x150 & x751 ) | ( ~x150 & n19099 ) | ( x751 & n19099 ) ;
  assign n19274 = ( x150 & x751 ) | ( x150 & ~n19114 ) | ( x751 & ~n19114 ) ;
  assign n19275 = n19273 | n19274 ;
  assign n19276 = ~n19272 & n19275 ;
  assign n19277 = x39 & ~n19276 ;
  assign n19278 = n19055 & ~n19264 ;
  assign n19279 = n19257 | n19278 ;
  assign n19280 = ( ~x38 & n9138 ) | ( ~x38 & n19279 ) | ( n9138 & n19279 ) ;
  assign n19281 = ~n19277 & n19280 ;
  assign n19282 = x751 & x947 ;
  assign n19283 = x39 | n19282 ;
  assign n19284 = n19236 & ~n19283 ;
  assign n19285 = x150 | n15070 ;
  assign n19286 = x38 & n19285 ;
  assign n19287 = ~n19284 & n19286 ;
  assign n19288 = x701 | n19287 ;
  assign n19289 = n19281 | n19288 ;
  assign n19290 = ~n19269 & n19289 ;
  assign n19291 = ( ~x832 & n8359 ) | ( ~x832 & n19290 ) | ( n8359 & n19290 ) ;
  assign n19292 = ( ~x150 & x832 ) | ( ~x150 & n8359 ) | ( x832 & n8359 ) ;
  assign n19293 = n19291 & ~n19292 ;
  assign n19294 = ~x701 & n18913 ;
  assign n19295 = n19264 | n19294 ;
  assign n19296 = ( ~x832 & n1290 ) | ( ~x832 & n19295 ) | ( n1290 & n19295 ) ;
  assign n19297 = ( x150 & x832 ) | ( x150 & n1290 ) | ( x832 & n1290 ) ;
  assign n19298 = ~n19296 & n19297 ;
  assign n19299 = n19293 | n19298 ;
  assign n19300 = ~x745 & x947 ;
  assign n19301 = ~x723 & n18913 ;
  assign n19302 = n19300 | n19301 ;
  assign n19303 = ( ~x832 & n1290 ) | ( ~x832 & n19302 ) | ( n1290 & n19302 ) ;
  assign n19304 = ( x151 & x832 ) | ( x151 & n1290 ) | ( x832 & n1290 ) ;
  assign n19305 = ~n19303 & n19304 ;
  assign n19306 = x151 | n14822 ;
  assign n19307 = ~x745 & n19016 ;
  assign n19308 = n19306 & ~n19307 ;
  assign n19309 = ~n19073 & n19308 ;
  assign n19310 = n14575 | n18999 ;
  assign n19311 = x151 | n19310 ;
  assign n19312 = ~n18909 & n19311 ;
  assign n19313 = x215 & ~n19312 ;
  assign n19314 = n2203 & n14682 ;
  assign n19315 = x151 & n2203 ;
  assign n19316 = ~n14684 & n19315 ;
  assign n19317 = n19314 | n19316 ;
  assign n19318 = x151 | n16705 ;
  assign n19319 = ~n19063 & n19318 ;
  assign n19320 = ~n19109 & n19319 ;
  assign n19321 = x215 | n19320 ;
  assign n19322 = n19317 | n19321 ;
  assign n19323 = ~n19313 & n19322 ;
  assign n19324 = x299 & ~n19323 ;
  assign n19325 = x151 & ~n19106 ;
  assign n19326 = n19096 | n19325 ;
  assign n19327 = ~n19324 & n19326 ;
  assign n19328 = x745 | n19327 ;
  assign n19329 = x151 | n18988 ;
  assign n19330 = ~n19069 & n19329 ;
  assign n19331 = x745 & ~n19330 ;
  assign n19332 = n19317 | n19319 ;
  assign n19333 = n19047 | n19332 ;
  assign n19334 = ~n19313 & n19333 ;
  assign n19335 = n19022 & ~n19334 ;
  assign n19336 = ( ~x299 & n19331 ) | ( ~x299 & n19335 ) | ( n19331 & n19335 ) ;
  assign n19337 = x39 & ~n19336 ;
  assign n19338 = n19328 & n19337 ;
  assign n19339 = n19309 | n19338 ;
  assign n19340 = ~x38 & n19339 ;
  assign n19341 = x745 & x947 ;
  assign n19342 = x39 | n19341 ;
  assign n19343 = n19236 & ~n19342 ;
  assign n19344 = x151 | n15070 ;
  assign n19345 = x38 & n19344 ;
  assign n19346 = ~n19343 & n19345 ;
  assign n19347 = x723 | n19346 ;
  assign n19348 = n19340 | n19347 ;
  assign n19349 = x151 & ~n14827 ;
  assign n19350 = n15070 & ~n19300 ;
  assign n19351 = n19349 | n19350 ;
  assign n19352 = x38 & n19351 ;
  assign n19353 = x723 & ~n19352 ;
  assign n19354 = ~x745 & n14709 ;
  assign n19355 = x151 | n14710 ;
  assign n19356 = n19354 | n19355 ;
  assign n19357 = ~n19026 & n19318 ;
  assign n19358 = n19317 | n19357 ;
  assign n19359 = n18996 | n19358 ;
  assign n19360 = n19059 & ~n19312 ;
  assign n19361 = x299 & ~n19360 ;
  assign n19362 = n19359 & n19361 ;
  assign n19363 = ~x745 & n19019 ;
  assign n19364 = ~n19362 & n19363 ;
  assign n19365 = n19356 & ~n19364 ;
  assign n19366 = ( x38 & x39 ) | ( x38 & ~n19365 ) | ( x39 & ~n19365 ) ;
  assign n19367 = ( ~x38 & x39 ) | ( ~x38 & n19308 ) | ( x39 & n19308 ) ;
  assign n19368 = ~n19366 & n19367 ;
  assign n19369 = n19353 & ~n19368 ;
  assign n19370 = n19348 & ~n19369 ;
  assign n19371 = ( ~x832 & n8359 ) | ( ~x832 & n19370 ) | ( n8359 & n19370 ) ;
  assign n19372 = ( ~x151 & x832 ) | ( ~x151 & n8359 ) | ( x832 & n8359 ) ;
  assign n19373 = n19371 & ~n19372 ;
  assign n19374 = n19305 | n19373 ;
  assign n19375 = x696 & n18913 ;
  assign n19376 = x759 & x947 ;
  assign n19377 = n1290 & ~n19376 ;
  assign n19378 = ~n19375 & n19377 ;
  assign n19379 = x152 | n1290 ;
  assign n19380 = x832 & n19379 ;
  assign n19381 = ~n19378 & n19380 ;
  assign n19382 = n14694 & ~n14696 ;
  assign n19383 = x152 | n19382 ;
  assign n19384 = ~x947 & n19382 ;
  assign n19385 = n1823 & ~n19384 ;
  assign n19386 = n19383 & n19385 ;
  assign n19387 = n4718 & n19382 ;
  assign n19388 = n1823 & ~n19387 ;
  assign n19389 = ~n19386 & n19388 ;
  assign n19390 = x152 & ~n16705 ;
  assign n19391 = n19109 | n19390 ;
  assign n19392 = ( ~x223 & n15629 ) | ( ~x223 & n19391 ) | ( n15629 & n19391 ) ;
  assign n19393 = ~n19389 & n19392 ;
  assign n19394 = x152 | n19089 ;
  assign n19395 = n19093 & n19394 ;
  assign n19396 = n19091 & n19394 ;
  assign n19397 = x299 | n19396 ;
  assign n19398 = n19395 | n19397 ;
  assign n19399 = n19393 | n19398 ;
  assign n19400 = n2203 | n19391 ;
  assign n19401 = ~x215 & n19400 ;
  assign n19402 = x152 & ~n19045 ;
  assign n19403 = n19060 & ~n19402 ;
  assign n19404 = ~n14684 & n19403 ;
  assign n19405 = n19401 & ~n19404 ;
  assign n19406 = x152 | n18909 ;
  assign n19407 = n18998 & n19406 ;
  assign n19408 = x299 & ~n19407 ;
  assign n19409 = ~n19405 & n19408 ;
  assign n19410 = x759 & ~n19409 ;
  assign n19411 = n19399 & n19410 ;
  assign n19412 = n19062 | n19390 ;
  assign n19413 = ~n1823 & n19412 ;
  assign n19414 = ~n18913 & n19382 ;
  assign n19415 = n1823 & ~n19414 ;
  assign n19416 = n19383 & n19415 ;
  assign n19417 = n19413 | n19416 ;
  assign n19418 = ~x223 & n19417 ;
  assign n19419 = x299 | n19395 ;
  assign n19420 = n19418 | n19419 ;
  assign n19421 = ~n19044 & n19401 ;
  assign n19422 = ~n19403 & n19421 ;
  assign n19423 = n14577 | n18913 ;
  assign n19424 = n19407 & n19423 ;
  assign n19425 = x299 & ~n19424 ;
  assign n19426 = ~n19422 & n19425 ;
  assign n19427 = x759 | n19426 ;
  assign n19428 = n19420 & ~n19427 ;
  assign n19429 = x39 & ~n19428 ;
  assign n19430 = ~n19411 & n19429 ;
  assign n19431 = x152 & ~n14822 ;
  assign n19432 = x39 | n19376 ;
  assign n19433 = n14832 & n19432 ;
  assign n19434 = n19431 | n19433 ;
  assign n19435 = n19072 | n19434 ;
  assign n19436 = ~x38 & n19435 ;
  assign n19437 = ~n19430 & n19436 ;
  assign n19438 = n15756 & ~n18913 ;
  assign n19439 = ~n19432 & n19438 ;
  assign n19440 = x152 | n15070 ;
  assign n19441 = x38 & n19440 ;
  assign n19442 = ~n19439 & n19441 ;
  assign n19443 = x696 & ~n19442 ;
  assign n19444 = ~n19437 & n19443 ;
  assign n19445 = n18995 | n19403 ;
  assign n19446 = ~n19023 & n19445 ;
  assign n19447 = n19025 | n19390 ;
  assign n19448 = ( ~x215 & n14841 ) | ( ~x215 & n19447 ) | ( n14841 & n19447 ) ;
  assign n19449 = ~n19446 & n19448 ;
  assign n19450 = x152 & n19000 ;
  assign n19451 = n19022 & ~n19450 ;
  assign n19452 = ~n19449 & n19451 ;
  assign n19453 = ~n1823 & n19447 ;
  assign n19454 = n19386 | n19453 ;
  assign n19455 = ~x223 & n19454 ;
  assign n19456 = n19397 | n19455 ;
  assign n19457 = x759 & n19456 ;
  assign n19458 = ~n19452 & n19457 ;
  assign n19459 = x759 | n14710 ;
  assign n19460 = x152 & ~n19459 ;
  assign n19461 = x39 & ~n19460 ;
  assign n19462 = ~n19458 & n19461 ;
  assign n19463 = ~x38 & n19434 ;
  assign n19464 = ~n19462 & n19463 ;
  assign n19465 = x152 | n14827 ;
  assign n19466 = n15070 & ~n19376 ;
  assign n19467 = x38 & ~n19466 ;
  assign n19468 = n19465 & n19467 ;
  assign n19469 = x696 | n19468 ;
  assign n19470 = n19464 | n19469 ;
  assign n19471 = ~n19444 & n19470 ;
  assign n19472 = ( ~x832 & n8359 ) | ( ~x832 & n19471 ) | ( n8359 & n19471 ) ;
  assign n19473 = ( ~x152 & x832 ) | ( ~x152 & n8359 ) | ( x832 & n8359 ) ;
  assign n19474 = n19472 & ~n19473 ;
  assign n19475 = n19381 | n19474 ;
  assign n19476 = x766 & x947 ;
  assign n19477 = n1290 & ~n19476 ;
  assign n19478 = x700 & n18913 ;
  assign n19479 = n19477 & ~n19478 ;
  assign n19480 = x153 & ~n1290 ;
  assign n19481 = x832 & ~n19480 ;
  assign n19482 = ~n19479 & n19481 ;
  assign n19483 = x153 | n14822 ;
  assign n19484 = ~x766 & n14823 ;
  assign n19485 = n19017 & ~n19484 ;
  assign n19486 = n19483 & ~n19485 ;
  assign n19487 = ~n19072 & n19486 ;
  assign n19488 = x153 & ~n18909 ;
  assign n19489 = n18998 & ~n19488 ;
  assign n19490 = x153 & n2203 ;
  assign n19491 = ~n14684 & n19490 ;
  assign n19492 = n19314 | n19491 ;
  assign n19493 = x153 | n16705 ;
  assign n19494 = ~n19026 & n19493 ;
  assign n19495 = ~n19061 & n19494 ;
  assign n19496 = x215 | n19495 ;
  assign n19497 = n19492 | n19496 ;
  assign n19498 = ~n19489 & n19497 ;
  assign n19499 = x299 & ~n19498 ;
  assign n19500 = x153 & ~n19106 ;
  assign n19501 = n19096 | n19500 ;
  assign n19502 = ~n19499 & n19501 ;
  assign n19503 = x766 & ~n19502 ;
  assign n19504 = ~n19063 & n19493 ;
  assign n19505 = n19046 | n19504 ;
  assign n19506 = n19492 | n19505 ;
  assign n19507 = ~x215 & n19506 ;
  assign n19508 = n14577 & ~n19489 ;
  assign n19509 = n19021 | n19508 ;
  assign n19510 = n19507 | n19509 ;
  assign n19511 = x299 & n19510 ;
  assign n19512 = x153 | n18988 ;
  assign n19513 = ~n19069 & n19512 ;
  assign n19514 = x766 | n19513 ;
  assign n19515 = n19511 | n19514 ;
  assign n19516 = x39 & n19515 ;
  assign n19517 = ~n19503 & n19516 ;
  assign n19518 = n19487 | n19517 ;
  assign n19519 = ~x38 & n19518 ;
  assign n19520 = ~x766 & x947 ;
  assign n19521 = x39 | n19520 ;
  assign n19522 = n19236 & ~n19521 ;
  assign n19523 = x153 | n15070 ;
  assign n19524 = x38 & n19523 ;
  assign n19525 = ~n19522 & n19524 ;
  assign n19526 = n19519 | n19525 ;
  assign n19527 = x700 & n19526 ;
  assign n19528 = ~n19019 & n19512 ;
  assign n19529 = n19492 | n19494 ;
  assign n19530 = n18996 | n19529 ;
  assign n19531 = n19000 & ~n19488 ;
  assign n19532 = x299 & ~n19531 ;
  assign n19533 = n19530 & n19532 ;
  assign n19534 = x766 & ~n19533 ;
  assign n19535 = ~n19528 & n19534 ;
  assign n19536 = x153 | x766 ;
  assign n19537 = n14710 | n19536 ;
  assign n19538 = x39 & n19537 ;
  assign n19539 = ~n19535 & n19538 ;
  assign n19540 = x38 | n19486 ;
  assign n19541 = n19539 | n19540 ;
  assign n19542 = x153 & ~n14827 ;
  assign n19543 = ~n4810 & n19477 ;
  assign n19544 = x38 & ~n19543 ;
  assign n19545 = ~n19542 & n19544 ;
  assign n19546 = x700 | n19545 ;
  assign n19547 = n19541 & ~n19546 ;
  assign n19548 = n19157 | n19547 ;
  assign n19549 = n19527 | n19548 ;
  assign n19550 = ~x153 & n19157 ;
  assign n19551 = x57 | n19550 ;
  assign n19552 = n19549 & ~n19551 ;
  assign n19553 = x57 & x153 ;
  assign n19554 = x832 | n19553 ;
  assign n19555 = n19552 | n19554 ;
  assign n19556 = ~n19482 & n19555 ;
  assign n19557 = x154 | n14822 ;
  assign n19558 = ~n19073 & n19557 ;
  assign n19559 = ~n19101 & n19558 ;
  assign n19560 = ( x39 & x154 ) | ( x39 & n19099 ) | ( x154 & n19099 ) ;
  assign n19561 = ( ~x39 & x154 ) | ( ~x39 & n19114 ) | ( x154 & n19114 ) ;
  assign n19562 = n19560 & ~n19561 ;
  assign n19563 = n19559 | n19562 ;
  assign n19564 = ~x38 & n19563 ;
  assign n19565 = x154 | n15070 ;
  assign n19566 = n19081 & n19565 ;
  assign n19567 = x742 | n19566 ;
  assign n19568 = n19564 | n19567 ;
  assign n19569 = ( x39 & x154 ) | ( x39 & n19053 ) | ( x154 & n19053 ) ;
  assign n19570 = ( ~x39 & x154 ) | ( ~x39 & n19070 ) | ( x154 & n19070 ) ;
  assign n19571 = n19569 & ~n19570 ;
  assign n19572 = n19558 | n19571 ;
  assign n19573 = ~x38 & n19572 ;
  assign n19574 = n19041 & n19565 ;
  assign n19575 = x742 & ~n19574 ;
  assign n19576 = ~n19573 & n19575 ;
  assign n19577 = x704 | n19576 ;
  assign n19578 = n19568 & ~n19577 ;
  assign n19579 = ~n19017 & n19557 ;
  assign n19580 = ( x39 & x154 ) | ( x39 & n19004 ) | ( x154 & n19004 ) ;
  assign n19581 = ( ~x39 & x154 ) | ( ~x39 & n19030 ) | ( x154 & n19030 ) ;
  assign n19582 = n19580 & ~n19581 ;
  assign n19583 = n19579 | n19582 ;
  assign n19584 = ~x38 & n19583 ;
  assign n19585 = x154 | n14827 ;
  assign n19586 = n19015 & n19585 ;
  assign n19587 = x742 | n19586 ;
  assign n19588 = n19584 | n19587 ;
  assign n19589 = ~x154 & x742 ;
  assign n19590 = ~n15382 & n19589 ;
  assign n19591 = x704 & ~n19590 ;
  assign n19592 = n19588 & n19591 ;
  assign n19593 = n8359 | n19592 ;
  assign n19594 = n19578 | n19593 ;
  assign n19595 = ~x154 & n8359 ;
  assign n19596 = x832 | n19595 ;
  assign n19597 = n19594 & ~n19596 ;
  assign n19598 = ~x742 & x947 ;
  assign n19599 = ~x704 & n18913 ;
  assign n19600 = n19598 | n19599 ;
  assign n19601 = ( ~x832 & n1290 ) | ( ~x832 & n19600 ) | ( n1290 & n19600 ) ;
  assign n19602 = ( x154 & x832 ) | ( x154 & n1290 ) | ( x832 & n1290 ) ;
  assign n19603 = ~n19601 & n19602 ;
  assign n19604 = n19597 | n19603 ;
  assign n19605 = ~x757 & n19034 ;
  assign n19606 = x686 & ~n19605 ;
  assign n19607 = n8359 | n19606 ;
  assign n19608 = x38 | n19074 ;
  assign n19609 = ~n19041 & n19608 ;
  assign n19610 = ( x686 & x757 ) | ( x686 & n19609 ) | ( x757 & n19609 ) ;
  assign n19611 = x38 | n19116 ;
  assign n19612 = ~n19081 & n19611 ;
  assign n19613 = ( x686 & ~x757 ) | ( x686 & n19612 ) | ( ~x757 & n19612 ) ;
  assign n19614 = n19610 | n19613 ;
  assign n19615 = ~n19607 & n19614 ;
  assign n19616 = x155 & ~n19615 ;
  assign n19617 = x757 | n19010 ;
  assign n19618 = x757 & ~n15382 ;
  assign n19619 = x686 & ~n19618 ;
  assign n19620 = n19617 & n19619 ;
  assign n19621 = ~x38 & n19057 ;
  assign n19622 = n15070 & n19041 ;
  assign n19623 = n19621 | n19622 ;
  assign n19624 = ( x686 & x757 ) | ( x686 & ~n19623 ) | ( x757 & ~n19623 ) ;
  assign n19625 = ~x38 & n19104 ;
  assign n19626 = x38 & n19078 ;
  assign n19627 = n19625 | n19626 ;
  assign n19628 = ( ~x686 & x757 ) | ( ~x686 & n19627 ) | ( x757 & n19627 ) ;
  assign n19629 = ~n19624 & n19628 ;
  assign n19630 = n19620 | n19629 ;
  assign n19631 = x155 | n8359 ;
  assign n19632 = n19630 & ~n19631 ;
  assign n19633 = n19616 | n19632 ;
  assign n19634 = ~x832 & n19633 ;
  assign n19635 = ~x757 & x947 ;
  assign n19636 = ~x686 & n18913 ;
  assign n19637 = n19635 | n19636 ;
  assign n19638 = ( ~x832 & n1290 ) | ( ~x832 & n19637 ) | ( n1290 & n19637 ) ;
  assign n19639 = ( x155 & x832 ) | ( x155 & n1290 ) | ( x832 & n1290 ) ;
  assign n19640 = ~n19638 & n19639 ;
  assign n19641 = n19634 | n19640 ;
  assign n19642 = ~x741 & n19010 ;
  assign n19643 = x741 & n15382 ;
  assign n19644 = x724 & ~n19643 ;
  assign n19645 = ~n19642 & n19644 ;
  assign n19646 = n8359 | n19645 ;
  assign n19647 = ( x724 & x741 ) | ( x724 & n19623 ) | ( x741 & n19623 ) ;
  assign n19648 = ( x724 & ~x741 ) | ( x724 & n19627 ) | ( ~x741 & n19627 ) ;
  assign n19649 = n19647 | n19648 ;
  assign n19650 = ~n19646 & n19649 ;
  assign n19651 = x156 | n19650 ;
  assign n19652 = x724 & ~x741 ;
  assign n19653 = n19034 & n19652 ;
  assign n19654 = ( x724 & x741 ) | ( x724 & ~n19609 ) | ( x741 & ~n19609 ) ;
  assign n19655 = ( ~x724 & x741 ) | ( ~x724 & n19612 ) | ( x741 & n19612 ) ;
  assign n19656 = ~n19654 & n19655 ;
  assign n19657 = n19653 | n19656 ;
  assign n19658 = x156 & ~n8359 ;
  assign n19659 = n19657 & n19658 ;
  assign n19660 = x832 | n19659 ;
  assign n19661 = n19651 & ~n19660 ;
  assign n19662 = ~x741 & x947 ;
  assign n19663 = ~x724 & n18913 ;
  assign n19664 = n19662 | n19663 ;
  assign n19665 = ( ~x832 & n1290 ) | ( ~x832 & n19664 ) | ( n1290 & n19664 ) ;
  assign n19666 = ( x156 & x832 ) | ( x156 & n1290 ) | ( x832 & n1290 ) ;
  assign n19667 = ~n19665 & n19666 ;
  assign n19668 = n19661 | n19667 ;
  assign n19669 = ~x760 & x947 ;
  assign n19670 = ~x688 & n18913 ;
  assign n19671 = n19669 | n19670 ;
  assign n19672 = ( ~x832 & n1290 ) | ( ~x832 & n19671 ) | ( n1290 & n19671 ) ;
  assign n19673 = ( x157 & x832 ) | ( x157 & n1290 ) | ( x832 & n1290 ) ;
  assign n19674 = ~n19672 & n19673 ;
  assign n19675 = x157 & ~n14827 ;
  assign n19676 = n15070 & ~n19669 ;
  assign n19677 = x38 & ~n19676 ;
  assign n19678 = ~n19675 & n19677 ;
  assign n19679 = x157 | n19001 ;
  assign n19680 = n11811 | n19029 ;
  assign n19681 = n19679 & n19680 ;
  assign n19682 = x157 | n18988 ;
  assign n19683 = ~n19019 & n19682 ;
  assign n19684 = x760 | n19683 ;
  assign n19685 = n19681 | n19684 ;
  assign n19686 = ~x157 & x760 ;
  assign n19687 = ~n14710 & n19686 ;
  assign n19688 = x39 & ~n19687 ;
  assign n19689 = n19685 & n19688 ;
  assign n19690 = ( x39 & n14822 ) | ( x39 & n19669 ) | ( n14822 & n19669 ) ;
  assign n19691 = ( ~x39 & x157 ) | ( ~x39 & n14822 ) | ( x157 & n14822 ) ;
  assign n19692 = ~n19690 & n19691 ;
  assign n19693 = x38 | n19692 ;
  assign n19694 = n19689 | n19693 ;
  assign n19695 = ~n19678 & n19694 ;
  assign n19696 = x688 & ~n19695 ;
  assign n19697 = ~n19072 & n19692 ;
  assign n19698 = ( x157 & ~x760 ) | ( x157 & n19070 ) | ( ~x760 & n19070 ) ;
  assign n19699 = ( x157 & x760 ) | ( x157 & n19114 ) | ( x760 & n19114 ) ;
  assign n19700 = n19698 & n19699 ;
  assign n19701 = x39 & ~n19700 ;
  assign n19702 = ( x157 & x760 ) | ( x157 & n19053 ) | ( x760 & n19053 ) ;
  assign n19703 = ( x157 & ~x760 ) | ( x157 & n19099 ) | ( ~x760 & n19099 ) ;
  assign n19704 = n19702 | n19703 ;
  assign n19705 = n19701 & n19704 ;
  assign n19706 = n19697 | n19705 ;
  assign n19707 = ~x38 & n19706 ;
  assign n19708 = x760 & x947 ;
  assign n19709 = x39 | n19708 ;
  assign n19710 = n19236 & ~n19709 ;
  assign n19711 = x157 | n15070 ;
  assign n19712 = x38 & n19711 ;
  assign n19713 = ~n19710 & n19712 ;
  assign n19714 = x688 | n19713 ;
  assign n19715 = n19707 | n19714 ;
  assign n19716 = ~n19696 & n19715 ;
  assign n19717 = ( ~x832 & n8359 ) | ( ~x832 & n19716 ) | ( n8359 & n19716 ) ;
  assign n19718 = ( ~x157 & x832 ) | ( ~x157 & n8359 ) | ( x832 & n8359 ) ;
  assign n19719 = n19717 & ~n19718 ;
  assign n19720 = n19674 | n19719 ;
  assign n19721 = ~x158 & x753 ;
  assign n19722 = ~n14710 & n19721 ;
  assign n19723 = ( ~x158 & x753 ) | ( ~x158 & n19004 ) | ( x753 & n19004 ) ;
  assign n19724 = ( x158 & x753 ) | ( x158 & ~n19030 ) | ( x753 & ~n19030 ) ;
  assign n19725 = n19723 | n19724 ;
  assign n19726 = ~n19722 & n19725 ;
  assign n19727 = x39 & ~n19726 ;
  assign n19728 = x158 & ~n14822 ;
  assign n19729 = x753 & n14822 ;
  assign n19730 = n19728 | n19729 ;
  assign n19731 = n18987 | n19730 ;
  assign n19732 = ~x38 & n19731 ;
  assign n19733 = ~n19727 & n19732 ;
  assign n19734 = x158 & ~n14827 ;
  assign n19735 = ~x753 & x947 ;
  assign n19736 = n15070 & ~n19735 ;
  assign n19737 = n19734 | n19736 ;
  assign n19738 = x38 & n19737 ;
  assign n19739 = x702 & ~n19738 ;
  assign n19740 = ~n19733 & n19739 ;
  assign n19741 = ( ~x158 & x753 ) | ( ~x158 & n19070 ) | ( x753 & n19070 ) ;
  assign n19742 = ( x158 & x753 ) | ( x158 & ~n19053 ) | ( x753 & ~n19053 ) ;
  assign n19743 = n19741 & n19742 ;
  assign n19744 = ( ~x158 & x753 ) | ( ~x158 & n19099 ) | ( x753 & n19099 ) ;
  assign n19745 = ( x158 & x753 ) | ( x158 & ~n19114 ) | ( x753 & ~n19114 ) ;
  assign n19746 = n19744 | n19745 ;
  assign n19747 = ~n19743 & n19746 ;
  assign n19748 = x39 & ~n19747 ;
  assign n19749 = n19055 & ~n19735 ;
  assign n19750 = n19728 | n19749 ;
  assign n19751 = ( ~x38 & n9138 ) | ( ~x38 & n19750 ) | ( n9138 & n19750 ) ;
  assign n19752 = ~n19748 & n19751 ;
  assign n19753 = x753 & x947 ;
  assign n19754 = x39 | n19753 ;
  assign n19755 = n19236 & ~n19754 ;
  assign n19756 = x158 | n15070 ;
  assign n19757 = x38 & n19756 ;
  assign n19758 = ~n19755 & n19757 ;
  assign n19759 = x702 | n19758 ;
  assign n19760 = n19752 | n19759 ;
  assign n19761 = ~n19740 & n19760 ;
  assign n19762 = ( ~x832 & n8359 ) | ( ~x832 & n19761 ) | ( n8359 & n19761 ) ;
  assign n19763 = ( ~x158 & x832 ) | ( ~x158 & n8359 ) | ( x832 & n8359 ) ;
  assign n19764 = n19762 & ~n19763 ;
  assign n19765 = ~x702 & n18913 ;
  assign n19766 = n19735 | n19765 ;
  assign n19767 = ( ~x832 & n1290 ) | ( ~x832 & n19766 ) | ( n1290 & n19766 ) ;
  assign n19768 = ( x158 & x832 ) | ( x158 & n1290 ) | ( x832 & n1290 ) ;
  assign n19769 = ~n19767 & n19768 ;
  assign n19770 = n19764 | n19769 ;
  assign n19771 = ~x159 & x754 ;
  assign n19772 = ~n14710 & n19771 ;
  assign n19773 = ( ~x159 & x754 ) | ( ~x159 & n19004 ) | ( x754 & n19004 ) ;
  assign n19774 = ( x159 & x754 ) | ( x159 & ~n19030 ) | ( x754 & ~n19030 ) ;
  assign n19775 = n19773 | n19774 ;
  assign n19776 = ~n19772 & n19775 ;
  assign n19777 = x39 & ~n19776 ;
  assign n19778 = x159 & ~n14822 ;
  assign n19779 = x754 & n14822 ;
  assign n19780 = n19778 | n19779 ;
  assign n19781 = n18987 | n19780 ;
  assign n19782 = ~x38 & n19781 ;
  assign n19783 = ~n19777 & n19782 ;
  assign n19784 = x159 & ~n14827 ;
  assign n19785 = ~x754 & x947 ;
  assign n19786 = n15070 & ~n19785 ;
  assign n19787 = n19784 | n19786 ;
  assign n19788 = x38 & n19787 ;
  assign n19789 = x709 & ~n19788 ;
  assign n19790 = ~n19783 & n19789 ;
  assign n19791 = ( ~x159 & x754 ) | ( ~x159 & n19070 ) | ( x754 & n19070 ) ;
  assign n19792 = ( x159 & x754 ) | ( x159 & ~n19053 ) | ( x754 & ~n19053 ) ;
  assign n19793 = n19791 & n19792 ;
  assign n19794 = ( ~x159 & x754 ) | ( ~x159 & n19099 ) | ( x754 & n19099 ) ;
  assign n19795 = ( x159 & x754 ) | ( x159 & ~n19114 ) | ( x754 & ~n19114 ) ;
  assign n19796 = n19794 | n19795 ;
  assign n19797 = ~n19793 & n19796 ;
  assign n19798 = x39 & ~n19797 ;
  assign n19799 = n19055 & ~n19785 ;
  assign n19800 = n19778 | n19799 ;
  assign n19801 = ( ~x38 & n9138 ) | ( ~x38 & n19800 ) | ( n9138 & n19800 ) ;
  assign n19802 = ~n19798 & n19801 ;
  assign n19803 = x754 & x947 ;
  assign n19804 = x39 | n19803 ;
  assign n19805 = n19236 & ~n19804 ;
  assign n19806 = x159 | n15070 ;
  assign n19807 = x38 & n19806 ;
  assign n19808 = ~n19805 & n19807 ;
  assign n19809 = x709 | n19808 ;
  assign n19810 = n19802 | n19809 ;
  assign n19811 = ~n19790 & n19810 ;
  assign n19812 = ( ~x832 & n8359 ) | ( ~x832 & n19811 ) | ( n8359 & n19811 ) ;
  assign n19813 = ( ~x159 & x832 ) | ( ~x159 & n8359 ) | ( x832 & n8359 ) ;
  assign n19814 = n19812 & ~n19813 ;
  assign n19815 = ~x709 & n18913 ;
  assign n19816 = n19785 | n19815 ;
  assign n19817 = ( ~x832 & n1290 ) | ( ~x832 & n19816 ) | ( n1290 & n19816 ) ;
  assign n19818 = ( x159 & x832 ) | ( x159 & n1290 ) | ( x832 & n1290 ) ;
  assign n19819 = ~n19817 & n19818 ;
  assign n19820 = n19814 | n19819 ;
  assign n19821 = ~x756 & x947 ;
  assign n19822 = ~x734 & n18913 ;
  assign n19823 = n19821 | n19822 ;
  assign n19824 = ( ~x832 & n1290 ) | ( ~x832 & n19823 ) | ( n1290 & n19823 ) ;
  assign n19825 = ( x160 & x832 ) | ( x160 & n1290 ) | ( x832 & n1290 ) ;
  assign n19826 = ~n19824 & n19825 ;
  assign n19827 = x160 & ~n14827 ;
  assign n19828 = n15070 & ~n19821 ;
  assign n19829 = x38 & ~n19828 ;
  assign n19830 = ~n19827 & n19829 ;
  assign n19831 = x160 | n18988 ;
  assign n19832 = ~n19019 & n19831 ;
  assign n19833 = x756 | n19832 ;
  assign n19834 = ( x160 & ~x299 ) | ( x160 & n19161 ) | ( ~x299 & n19161 ) ;
  assign n19835 = ( x160 & x299 ) | ( x160 & n19001 ) | ( x299 & n19001 ) ;
  assign n19836 = ~n19834 & n19835 ;
  assign n19837 = n19833 | n19836 ;
  assign n19838 = ~x160 & x756 ;
  assign n19839 = ~n14710 & n19838 ;
  assign n19840 = x39 & ~n19839 ;
  assign n19841 = n19837 & n19840 ;
  assign n19842 = ( x39 & n14822 ) | ( x39 & n19821 ) | ( n14822 & n19821 ) ;
  assign n19843 = ( ~x39 & x160 ) | ( ~x39 & n14822 ) | ( x160 & n14822 ) ;
  assign n19844 = ~n19842 & n19843 ;
  assign n19845 = x38 | n19844 ;
  assign n19846 = n19841 | n19845 ;
  assign n19847 = ~n19830 & n19846 ;
  assign n19848 = x734 & ~n19847 ;
  assign n19849 = ~n19072 & n19844 ;
  assign n19850 = x756 & ~n19052 ;
  assign n19851 = ( ~x160 & n19135 ) | ( ~x160 & n19850 ) | ( n19135 & n19850 ) ;
  assign n19852 = ( x160 & ~n19051 ) | ( x160 & n19850 ) | ( ~n19051 & n19850 ) ;
  assign n19853 = n19851 & n19852 ;
  assign n19854 = x39 & ~n19853 ;
  assign n19855 = ( ~x160 & x756 ) | ( ~x160 & n19099 ) | ( x756 & n19099 ) ;
  assign n19856 = ( x160 & x756 ) | ( x160 & ~n19114 ) | ( x756 & ~n19114 ) ;
  assign n19857 = n19855 | n19856 ;
  assign n19858 = n19854 & n19857 ;
  assign n19859 = n19849 | n19858 ;
  assign n19860 = ~x38 & n19859 ;
  assign n19861 = x756 & x947 ;
  assign n19862 = x39 | n19861 ;
  assign n19863 = n19236 & ~n19862 ;
  assign n19864 = x160 | n15070 ;
  assign n19865 = x38 & n19864 ;
  assign n19866 = ~n19863 & n19865 ;
  assign n19867 = x734 | n19866 ;
  assign n19868 = n19860 | n19867 ;
  assign n19869 = ~n19848 & n19868 ;
  assign n19870 = ( ~x832 & n8359 ) | ( ~x832 & n19869 ) | ( n8359 & n19869 ) ;
  assign n19871 = ( ~x160 & x832 ) | ( ~x160 & n8359 ) | ( x832 & n8359 ) ;
  assign n19872 = n19870 & ~n19871 ;
  assign n19873 = n19826 | n19872 ;
  assign n19874 = x736 & n18913 ;
  assign n19875 = x758 & x947 ;
  assign n19876 = n1290 & ~n19875 ;
  assign n19877 = ~n19874 & n19876 ;
  assign n19878 = x161 | n1290 ;
  assign n19879 = x832 & n19878 ;
  assign n19880 = ~n19877 & n19879 ;
  assign n19881 = x161 | n19382 ;
  assign n19882 = n19385 & n19881 ;
  assign n19883 = n19388 & ~n19882 ;
  assign n19884 = x161 & ~n16705 ;
  assign n19885 = n19109 | n19884 ;
  assign n19886 = ( ~x223 & n15629 ) | ( ~x223 & n19885 ) | ( n15629 & n19885 ) ;
  assign n19887 = ~n19883 & n19886 ;
  assign n19888 = x161 | n19089 ;
  assign n19889 = n19093 & n19888 ;
  assign n19890 = n19091 & n19888 ;
  assign n19891 = x299 | n19890 ;
  assign n19892 = n19889 | n19891 ;
  assign n19893 = n19887 | n19892 ;
  assign n19894 = n2203 | n19885 ;
  assign n19895 = ~x215 & n19894 ;
  assign n19896 = x161 & ~n19045 ;
  assign n19897 = n19060 & ~n19896 ;
  assign n19898 = ~n14684 & n19897 ;
  assign n19899 = n19895 & ~n19898 ;
  assign n19900 = x161 | n18909 ;
  assign n19901 = n18998 & n19900 ;
  assign n19902 = x299 & ~n19901 ;
  assign n19903 = ~n19899 & n19902 ;
  assign n19904 = x758 & ~n19903 ;
  assign n19905 = n19893 & n19904 ;
  assign n19906 = n19062 | n19884 ;
  assign n19907 = ~n1823 & n19906 ;
  assign n19908 = n19415 & n19881 ;
  assign n19909 = n19907 | n19908 ;
  assign n19910 = ~x223 & n19909 ;
  assign n19911 = x299 | n19889 ;
  assign n19912 = n19910 | n19911 ;
  assign n19913 = ~n19044 & n19895 ;
  assign n19914 = ~n19897 & n19913 ;
  assign n19915 = n19423 & n19901 ;
  assign n19916 = x299 & ~n19915 ;
  assign n19917 = ~n19914 & n19916 ;
  assign n19918 = x758 | n19917 ;
  assign n19919 = n19912 & ~n19918 ;
  assign n19920 = x39 & ~n19919 ;
  assign n19921 = ~n19905 & n19920 ;
  assign n19922 = ( x39 & n14822 ) | ( x39 & n19875 ) | ( n14822 & n19875 ) ;
  assign n19923 = ( x39 & x161 ) | ( x39 & ~n14822 ) | ( x161 & ~n14822 ) ;
  assign n19924 = n19922 | n19923 ;
  assign n19925 = n19072 | n19924 ;
  assign n19926 = ~x38 & n19925 ;
  assign n19927 = ~n19921 & n19926 ;
  assign n19928 = x39 | n19875 ;
  assign n19929 = n19438 & ~n19928 ;
  assign n19930 = x161 | n15070 ;
  assign n19931 = x38 & n19930 ;
  assign n19932 = ~n19929 & n19931 ;
  assign n19933 = x736 & ~n19932 ;
  assign n19934 = ~n19927 & n19933 ;
  assign n19935 = n18995 | n19897 ;
  assign n19936 = ~n19023 & n19935 ;
  assign n19937 = n19025 | n19884 ;
  assign n19938 = ( ~x215 & n14841 ) | ( ~x215 & n19937 ) | ( n14841 & n19937 ) ;
  assign n19939 = ~n19936 & n19938 ;
  assign n19940 = x161 & n19000 ;
  assign n19941 = n19022 & ~n19940 ;
  assign n19942 = ~n19939 & n19941 ;
  assign n19943 = ~n1823 & n19937 ;
  assign n19944 = n19882 | n19943 ;
  assign n19945 = ~x223 & n19944 ;
  assign n19946 = n19891 | n19945 ;
  assign n19947 = x758 & n19946 ;
  assign n19948 = ~n19942 & n19947 ;
  assign n19949 = x161 & ~n17986 ;
  assign n19950 = x39 & ~n19949 ;
  assign n19951 = ~n19948 & n19950 ;
  assign n19952 = ~x38 & n19924 ;
  assign n19953 = ~n19951 & n19952 ;
  assign n19954 = x161 | n14827 ;
  assign n19955 = n15070 & ~n19875 ;
  assign n19956 = x38 & ~n19955 ;
  assign n19957 = n19954 & n19956 ;
  assign n19958 = x736 | n19957 ;
  assign n19959 = n19953 | n19958 ;
  assign n19960 = ~n19934 & n19959 ;
  assign n19961 = ( ~x832 & n8359 ) | ( ~x832 & n19960 ) | ( n8359 & n19960 ) ;
  assign n19962 = ( ~x161 & x832 ) | ( ~x161 & n8359 ) | ( x832 & n8359 ) ;
  assign n19963 = n19961 & ~n19962 ;
  assign n19964 = n19880 | n19963 ;
  assign n19965 = x162 & ~n14827 ;
  assign n19966 = ~x761 & x947 ;
  assign n19967 = n15070 & ~n19966 ;
  assign n19968 = x38 & ~n19967 ;
  assign n19969 = ~n19965 & n19968 ;
  assign n19970 = n13052 & n19161 ;
  assign n19971 = n18990 | n19970 ;
  assign n19972 = ~x761 & n19971 ;
  assign n19973 = x39 & ~n19972 ;
  assign n19974 = ( x162 & x761 ) | ( x162 & n14710 ) | ( x761 & n14710 ) ;
  assign n19975 = ( x162 & ~x761 ) | ( x162 & n19003 ) | ( ~x761 & n19003 ) ;
  assign n19976 = n19974 | n19975 ;
  assign n19977 = n19973 & n19976 ;
  assign n19978 = ( x39 & n14822 ) | ( x39 & n19966 ) | ( n14822 & n19966 ) ;
  assign n19979 = ( ~x39 & x162 ) | ( ~x39 & n14822 ) | ( x162 & n14822 ) ;
  assign n19980 = ~n19978 & n19979 ;
  assign n19981 = x38 | n19980 ;
  assign n19982 = n19977 | n19981 ;
  assign n19983 = ~n19969 & n19982 ;
  assign n19984 = x738 & ~n19983 ;
  assign n19985 = ~n19072 & n19980 ;
  assign n19986 = ~n13052 & n19053 ;
  assign n19987 = x162 & ~n19135 ;
  assign n19988 = x761 & ~n19987 ;
  assign n19989 = ~n19986 & n19988 ;
  assign n19990 = x39 & ~n19989 ;
  assign n19991 = ( ~x162 & x761 ) | ( ~x162 & n19099 ) | ( x761 & n19099 ) ;
  assign n19992 = ( x162 & x761 ) | ( x162 & ~n19114 ) | ( x761 & ~n19114 ) ;
  assign n19993 = n19991 | n19992 ;
  assign n19994 = n19990 & n19993 ;
  assign n19995 = n19985 | n19994 ;
  assign n19996 = ~x38 & n19995 ;
  assign n19997 = x761 & x947 ;
  assign n19998 = x39 | n19997 ;
  assign n19999 = n19236 & ~n19998 ;
  assign n20000 = x162 | n15070 ;
  assign n20001 = x38 & n20000 ;
  assign n20002 = ~n19999 & n20001 ;
  assign n20003 = x738 | n20002 ;
  assign n20004 = n19996 | n20003 ;
  assign n20005 = ~n19984 & n20004 ;
  assign n20006 = ( ~x832 & n8359 ) | ( ~x832 & n20005 ) | ( n8359 & n20005 ) ;
  assign n20007 = ( ~x162 & x832 ) | ( ~x162 & n8359 ) | ( x832 & n8359 ) ;
  assign n20008 = n20006 & ~n20007 ;
  assign n20009 = ~x738 & n18913 ;
  assign n20010 = n19966 | n20009 ;
  assign n20011 = ( ~x832 & n1290 ) | ( ~x832 & n20010 ) | ( n1290 & n20010 ) ;
  assign n20012 = ( x162 & x832 ) | ( x162 & n1290 ) | ( x832 & n1290 ) ;
  assign n20013 = ~n20011 & n20012 ;
  assign n20014 = n20008 | n20013 ;
  assign n20015 = ~x777 & x947 ;
  assign n20016 = ~x737 & n18913 ;
  assign n20017 = n20015 | n20016 ;
  assign n20018 = ( ~x832 & n1290 ) | ( ~x832 & n20017 ) | ( n1290 & n20017 ) ;
  assign n20019 = ( x163 & x832 ) | ( x163 & n1290 ) | ( x832 & n1290 ) ;
  assign n20020 = ~n20018 & n20019 ;
  assign n20021 = x163 & ~n14827 ;
  assign n20022 = n15070 & ~n20015 ;
  assign n20023 = x38 & ~n20022 ;
  assign n20024 = ~n20021 & n20023 ;
  assign n20025 = x163 | n19001 ;
  assign n20026 = n12686 | n19029 ;
  assign n20027 = n20025 & n20026 ;
  assign n20028 = x163 | n18988 ;
  assign n20029 = ~n19019 & n20028 ;
  assign n20030 = x777 | n20029 ;
  assign n20031 = n20027 | n20030 ;
  assign n20032 = ~x163 & x777 ;
  assign n20033 = ~n14710 & n20032 ;
  assign n20034 = x39 & ~n20033 ;
  assign n20035 = n20031 & n20034 ;
  assign n20036 = ( x39 & n14822 ) | ( x39 & n20015 ) | ( n14822 & n20015 ) ;
  assign n20037 = ( ~x39 & x163 ) | ( ~x39 & n14822 ) | ( x163 & n14822 ) ;
  assign n20038 = ~n20036 & n20037 ;
  assign n20039 = x38 | n20038 ;
  assign n20040 = n20035 | n20039 ;
  assign n20041 = ~n20024 & n20040 ;
  assign n20042 = x737 & ~n20041 ;
  assign n20043 = ~n19072 & n20038 ;
  assign n20044 = x777 & ~n19052 ;
  assign n20045 = ( ~x163 & n19135 ) | ( ~x163 & n20044 ) | ( n19135 & n20044 ) ;
  assign n20046 = ( x163 & ~n19051 ) | ( x163 & n20044 ) | ( ~n19051 & n20044 ) ;
  assign n20047 = n20045 & n20046 ;
  assign n20048 = x39 & ~n20047 ;
  assign n20049 = ( ~x163 & x777 ) | ( ~x163 & n19099 ) | ( x777 & n19099 ) ;
  assign n20050 = ( x163 & x777 ) | ( x163 & ~n19114 ) | ( x777 & ~n19114 ) ;
  assign n20051 = n20049 | n20050 ;
  assign n20052 = n20048 & n20051 ;
  assign n20053 = n20043 | n20052 ;
  assign n20054 = ~x38 & n20053 ;
  assign n20055 = x777 & x947 ;
  assign n20056 = x39 | n20055 ;
  assign n20057 = n19236 & ~n20056 ;
  assign n20058 = x163 | n15070 ;
  assign n20059 = x38 & n20058 ;
  assign n20060 = ~n20057 & n20059 ;
  assign n20061 = x737 | n20060 ;
  assign n20062 = n20054 | n20061 ;
  assign n20063 = ~n20042 & n20062 ;
  assign n20064 = ( ~x832 & n8359 ) | ( ~x832 & n20063 ) | ( n8359 & n20063 ) ;
  assign n20065 = ( ~x163 & x832 ) | ( ~x163 & n8359 ) | ( x832 & n8359 ) ;
  assign n20066 = n20064 & ~n20065 ;
  assign n20067 = n20020 | n20066 ;
  assign n20068 = ~x752 & x947 ;
  assign n20069 = x703 & n18913 ;
  assign n20070 = n20068 | n20069 ;
  assign n20071 = ( ~x832 & n1290 ) | ( ~x832 & n20070 ) | ( n1290 & n20070 ) ;
  assign n20072 = ( x164 & x832 ) | ( x164 & n1290 ) | ( x832 & n1290 ) ;
  assign n20073 = ~n20071 & n20072 ;
  assign n20074 = x164 | n19078 ;
  assign n20075 = n19081 & n20074 ;
  assign n20076 = x752 | n20075 ;
  assign n20077 = ( ~x38 & x164 ) | ( ~x38 & n19104 ) | ( x164 & n19104 ) ;
  assign n20078 = ( x38 & x164 ) | ( x38 & n19116 ) | ( x164 & n19116 ) ;
  assign n20079 = n20077 & ~n20078 ;
  assign n20080 = n20076 | n20079 ;
  assign n20081 = x164 | n15070 ;
  assign n20082 = n19041 & n20081 ;
  assign n20083 = x752 & ~n20082 ;
  assign n20084 = ( ~x38 & x164 ) | ( ~x38 & n19057 ) | ( x164 & n19057 ) ;
  assign n20085 = ( x38 & x164 ) | ( x38 & n19074 ) | ( x164 & n19074 ) ;
  assign n20086 = n20084 & ~n20085 ;
  assign n20087 = n20083 & ~n20086 ;
  assign n20088 = n20080 & ~n20087 ;
  assign n20089 = x703 & ~n20088 ;
  assign n20090 = x164 & ~n19009 ;
  assign n20091 = x752 | n20090 ;
  assign n20092 = n19010 & ~n20091 ;
  assign n20093 = ~x752 & n19034 ;
  assign n20094 = x164 & ~n20093 ;
  assign n20095 = x752 & n15382 ;
  assign n20096 = x703 | n20095 ;
  assign n20097 = n20094 | n20096 ;
  assign n20098 = n20092 | n20097 ;
  assign n20099 = ~n20089 & n20098 ;
  assign n20100 = ( ~x832 & n8359 ) | ( ~x832 & n20099 ) | ( n8359 & n20099 ) ;
  assign n20101 = ( ~x164 & x832 ) | ( ~x164 & n8359 ) | ( x832 & n8359 ) ;
  assign n20102 = n20100 & ~n20101 ;
  assign n20103 = n20073 | n20102 ;
  assign n20104 = ~x774 & x947 ;
  assign n20105 = x687 & n18913 ;
  assign n20106 = n20104 | n20105 ;
  assign n20107 = ( ~x832 & n1290 ) | ( ~x832 & n20106 ) | ( n1290 & n20106 ) ;
  assign n20108 = ( x165 & x832 ) | ( x165 & n1290 ) | ( x832 & n1290 ) ;
  assign n20109 = ~n20107 & n20108 ;
  assign n20110 = x165 | n19078 ;
  assign n20111 = n19081 & n20110 ;
  assign n20112 = x774 | n20111 ;
  assign n20113 = ( ~x38 & x165 ) | ( ~x38 & n19104 ) | ( x165 & n19104 ) ;
  assign n20114 = ( x38 & x165 ) | ( x38 & n19116 ) | ( x165 & n19116 ) ;
  assign n20115 = n20113 & ~n20114 ;
  assign n20116 = n20112 | n20115 ;
  assign n20117 = x165 | n15070 ;
  assign n20118 = n19041 & n20117 ;
  assign n20119 = x774 & ~n20118 ;
  assign n20120 = ( ~x38 & x165 ) | ( ~x38 & n19057 ) | ( x165 & n19057 ) ;
  assign n20121 = ( x38 & x165 ) | ( x38 & n19074 ) | ( x165 & n19074 ) ;
  assign n20122 = n20120 & ~n20121 ;
  assign n20123 = n20119 & ~n20122 ;
  assign n20124 = n20116 & ~n20123 ;
  assign n20125 = x687 & ~n20124 ;
  assign n20126 = x165 & ~n19009 ;
  assign n20127 = x774 | n20126 ;
  assign n20128 = n19010 & ~n20127 ;
  assign n20129 = ~x774 & n19034 ;
  assign n20130 = x165 & ~n20129 ;
  assign n20131 = x774 & n15382 ;
  assign n20132 = x687 | n20131 ;
  assign n20133 = n20130 | n20132 ;
  assign n20134 = n20128 | n20133 ;
  assign n20135 = ~n20125 & n20134 ;
  assign n20136 = ( ~x832 & n8359 ) | ( ~x832 & n20135 ) | ( n8359 & n20135 ) ;
  assign n20137 = ( ~x165 & x832 ) | ( ~x165 & n8359 ) | ( x832 & n8359 ) ;
  assign n20138 = n20136 & ~n20137 ;
  assign n20139 = n20109 | n20138 ;
  assign n20140 = x727 & n18913 ;
  assign n20141 = x772 & x947 ;
  assign n20142 = n1290 & ~n20141 ;
  assign n20143 = ~n20140 & n20142 ;
  assign n20144 = x166 | n1290 ;
  assign n20145 = x832 & n20144 ;
  assign n20146 = ~n20143 & n20145 ;
  assign n20147 = x166 & ~n19045 ;
  assign n20148 = n19060 & ~n20147 ;
  assign n20149 = n18995 | n20148 ;
  assign n20150 = ~n19023 & n20149 ;
  assign n20151 = x166 & ~n16705 ;
  assign n20152 = n19025 | n20151 ;
  assign n20153 = ( ~x215 & n14841 ) | ( ~x215 & n20152 ) | ( n14841 & n20152 ) ;
  assign n20154 = ~n20150 & n20153 ;
  assign n20155 = x166 & n19000 ;
  assign n20156 = n19022 & ~n20155 ;
  assign n20157 = ~n20154 & n20156 ;
  assign n20158 = x166 | n19089 ;
  assign n20159 = n19091 & n20158 ;
  assign n20160 = x299 | n20159 ;
  assign n20161 = ~n1823 & n20152 ;
  assign n20162 = x166 | n19382 ;
  assign n20163 = n19385 & n20162 ;
  assign n20164 = n20161 | n20163 ;
  assign n20165 = ~x223 & n20164 ;
  assign n20166 = n20160 | n20165 ;
  assign n20167 = x772 & n20166 ;
  assign n20168 = ~n20157 & n20167 ;
  assign n20169 = x772 | n14710 ;
  assign n20170 = x166 & ~n20169 ;
  assign n20171 = x39 & ~n20170 ;
  assign n20172 = ~n20168 & n20171 ;
  assign n20173 = x166 & ~n14822 ;
  assign n20174 = x39 | n20141 ;
  assign n20175 = n14832 & n20174 ;
  assign n20176 = n20173 | n20175 ;
  assign n20177 = ~x38 & n20176 ;
  assign n20178 = ~n20172 & n20177 ;
  assign n20179 = x166 | n14827 ;
  assign n20180 = n15070 & ~n20141 ;
  assign n20181 = x38 & ~n20180 ;
  assign n20182 = n20179 & n20181 ;
  assign n20183 = x727 | n20182 ;
  assign n20184 = n20178 | n20183 ;
  assign n20185 = n19109 | n20151 ;
  assign n20186 = ( ~x215 & n14841 ) | ( ~x215 & n20185 ) | ( n14841 & n20185 ) ;
  assign n20187 = ~n19044 & n20186 ;
  assign n20188 = ~n20148 & n20187 ;
  assign n20189 = x166 | n18909 ;
  assign n20190 = n18998 & n20189 ;
  assign n20191 = n19423 & n20190 ;
  assign n20192 = x299 & ~n20191 ;
  assign n20193 = ~n20188 & n20192 ;
  assign n20194 = n4718 & n19089 ;
  assign n20195 = x166 | n20194 ;
  assign n20196 = n19093 & n20195 ;
  assign n20197 = x299 | n20196 ;
  assign n20198 = n1823 | n20185 ;
  assign n20199 = ~x223 & n20198 ;
  assign n20200 = ( n1823 & ~n19025 ) | ( n1823 & n20199 ) | ( ~n19025 & n20199 ) ;
  assign n20201 = ~n19414 & n20162 ;
  assign n20202 = ( ~n1823 & n20199 ) | ( ~n1823 & n20201 ) | ( n20199 & n20201 ) ;
  assign n20203 = n20200 & n20202 ;
  assign n20204 = n20197 | n20203 ;
  assign n20205 = ~x772 & n20204 ;
  assign n20206 = ~n20193 & n20205 ;
  assign n20207 = ~n14684 & n20148 ;
  assign n20208 = n20186 & ~n20207 ;
  assign n20209 = x299 & ~n20190 ;
  assign n20210 = ~n20208 & n20209 ;
  assign n20211 = n19388 & ~n20201 ;
  assign n20212 = n20199 & ~n20211 ;
  assign n20213 = n20160 | n20196 ;
  assign n20214 = n20212 | n20213 ;
  assign n20215 = x772 & n20214 ;
  assign n20216 = ~n20210 & n20215 ;
  assign n20217 = x39 & ~n20216 ;
  assign n20218 = ~n20206 & n20217 ;
  assign n20219 = n19072 | n20176 ;
  assign n20220 = ~x38 & n20219 ;
  assign n20221 = ~n20218 & n20220 ;
  assign n20222 = x166 | n15070 ;
  assign n20223 = n19438 & ~n20174 ;
  assign n20224 = x38 & ~n20223 ;
  assign n20225 = n20222 & n20224 ;
  assign n20226 = x727 & ~n20225 ;
  assign n20227 = ~n20221 & n20226 ;
  assign n20228 = n20184 & ~n20227 ;
  assign n20229 = ( ~x832 & n8359 ) | ( ~x832 & n20228 ) | ( n8359 & n20228 ) ;
  assign n20230 = ( ~x166 & x832 ) | ( ~x166 & n8359 ) | ( x832 & n8359 ) ;
  assign n20231 = n20229 & ~n20230 ;
  assign n20232 = n20146 | n20231 ;
  assign n20233 = x167 | n19078 ;
  assign n20234 = n19081 & n20233 ;
  assign n20235 = x768 | n20234 ;
  assign n20236 = ( ~x38 & x167 ) | ( ~x38 & n19104 ) | ( x167 & n19104 ) ;
  assign n20237 = ( x38 & x167 ) | ( x38 & n19116 ) | ( x167 & n19116 ) ;
  assign n20238 = n20236 & ~n20237 ;
  assign n20239 = n20235 | n20238 ;
  assign n20240 = x167 | n15070 ;
  assign n20241 = n19041 & n20240 ;
  assign n20242 = x768 & ~n20241 ;
  assign n20243 = ( ~x38 & x167 ) | ( ~x38 & n19057 ) | ( x167 & n19057 ) ;
  assign n20244 = ( x38 & x167 ) | ( x38 & n19074 ) | ( x167 & n19074 ) ;
  assign n20245 = n20243 & ~n20244 ;
  assign n20246 = n20242 & ~n20245 ;
  assign n20247 = x705 & ~n20246 ;
  assign n20248 = n20239 & n20247 ;
  assign n20249 = x167 | n14827 ;
  assign n20250 = n19015 & n20249 ;
  assign n20251 = x768 | n20250 ;
  assign n20252 = ( ~x38 & x167 ) | ( ~x38 & n19006 ) | ( x167 & n19006 ) ;
  assign n20253 = ( x38 & x167 ) | ( x38 & n19032 ) | ( x167 & n19032 ) ;
  assign n20254 = n20252 & ~n20253 ;
  assign n20255 = n20251 | n20254 ;
  assign n20256 = x768 & ~n15382 ;
  assign n20257 = ~x167 & n20256 ;
  assign n20258 = x705 | n20257 ;
  assign n20259 = n20255 & ~n20258 ;
  assign n20260 = n8359 | n20259 ;
  assign n20261 = n20248 | n20260 ;
  assign n20262 = ~x167 & n8359 ;
  assign n20263 = x832 | n20262 ;
  assign n20264 = n20261 & ~n20263 ;
  assign n20265 = ~x768 & x947 ;
  assign n20266 = x705 & n18913 ;
  assign n20267 = n20265 | n20266 ;
  assign n20268 = ( ~x832 & n1290 ) | ( ~x832 & n20267 ) | ( n1290 & n20267 ) ;
  assign n20269 = ( x167 & x832 ) | ( x167 & n1290 ) | ( x832 & n1290 ) ;
  assign n20270 = ~n20268 & n20269 ;
  assign n20271 = n20264 | n20270 ;
  assign n20272 = x763 & x947 ;
  assign n20273 = n1290 & ~n20272 ;
  assign n20274 = x699 & n18913 ;
  assign n20275 = n20273 & ~n20274 ;
  assign n20276 = x168 & ~n1290 ;
  assign n20277 = x832 & ~n20276 ;
  assign n20278 = ~n20275 & n20277 ;
  assign n20279 = x168 | n14822 ;
  assign n20280 = ~x763 & n14823 ;
  assign n20281 = n19017 & ~n20280 ;
  assign n20282 = n20279 & ~n20281 ;
  assign n20283 = ~n19072 & n20282 ;
  assign n20284 = x168 & ~n18909 ;
  assign n20285 = n18998 & ~n20284 ;
  assign n20286 = x168 & n2203 ;
  assign n20287 = ~n14684 & n20286 ;
  assign n20288 = n19314 | n20287 ;
  assign n20289 = x168 | n16705 ;
  assign n20290 = ~n19026 & n20289 ;
  assign n20291 = ~n19061 & n20290 ;
  assign n20292 = x215 | n20291 ;
  assign n20293 = n20288 | n20292 ;
  assign n20294 = ~n20285 & n20293 ;
  assign n20295 = x299 & ~n20294 ;
  assign n20296 = x168 & ~n19106 ;
  assign n20297 = n19096 | n20296 ;
  assign n20298 = ~n20295 & n20297 ;
  assign n20299 = x763 & ~n20298 ;
  assign n20300 = ~n19063 & n20289 ;
  assign n20301 = n19046 | n20300 ;
  assign n20302 = n20288 | n20301 ;
  assign n20303 = ~x215 & n20302 ;
  assign n20304 = n14577 & ~n20285 ;
  assign n20305 = n19021 | n20304 ;
  assign n20306 = n20303 | n20305 ;
  assign n20307 = x299 & n20306 ;
  assign n20308 = x168 | n18988 ;
  assign n20309 = ~n19069 & n20308 ;
  assign n20310 = x763 | n20309 ;
  assign n20311 = n20307 | n20310 ;
  assign n20312 = x39 & n20311 ;
  assign n20313 = ~n20299 & n20312 ;
  assign n20314 = n20283 | n20313 ;
  assign n20315 = ~x38 & n20314 ;
  assign n20316 = ~x763 & x947 ;
  assign n20317 = x39 | n20316 ;
  assign n20318 = n19236 & ~n20317 ;
  assign n20319 = x168 | n15070 ;
  assign n20320 = x38 & n20319 ;
  assign n20321 = ~n20318 & n20320 ;
  assign n20322 = n20315 | n20321 ;
  assign n20323 = x699 & n20322 ;
  assign n20324 = ~n19019 & n20308 ;
  assign n20325 = n20288 | n20290 ;
  assign n20326 = n18996 | n20325 ;
  assign n20327 = n19000 & ~n20284 ;
  assign n20328 = x299 & ~n20327 ;
  assign n20329 = n20326 & n20328 ;
  assign n20330 = x763 & ~n20329 ;
  assign n20331 = ~n20324 & n20330 ;
  assign n20332 = x168 | x763 ;
  assign n20333 = n14710 | n20332 ;
  assign n20334 = x39 & n20333 ;
  assign n20335 = ~n20331 & n20334 ;
  assign n20336 = x38 | n20282 ;
  assign n20337 = n20335 | n20336 ;
  assign n20338 = x168 & ~n14827 ;
  assign n20339 = ~n4810 & n20273 ;
  assign n20340 = x38 & ~n20339 ;
  assign n20341 = ~n20338 & n20340 ;
  assign n20342 = x699 | n20341 ;
  assign n20343 = n20337 & ~n20342 ;
  assign n20344 = n19157 | n20343 ;
  assign n20345 = n20323 | n20344 ;
  assign n20346 = ~x168 & n19157 ;
  assign n20347 = x57 | n20346 ;
  assign n20348 = n20345 & ~n20347 ;
  assign n20349 = x57 & x168 ;
  assign n20350 = x832 | n20349 ;
  assign n20351 = n20348 | n20350 ;
  assign n20352 = ~n20278 & n20351 ;
  assign n20353 = x746 & x947 ;
  assign n20354 = n1290 & ~n20353 ;
  assign n20355 = x729 & n18913 ;
  assign n20356 = n20354 & ~n20355 ;
  assign n20357 = x169 & ~n1290 ;
  assign n20358 = x832 & ~n20357 ;
  assign n20359 = ~n20356 & n20358 ;
  assign n20360 = x169 | n14822 ;
  assign n20361 = ~x746 & n14823 ;
  assign n20362 = n19017 & ~n20361 ;
  assign n20363 = n20360 & ~n20362 ;
  assign n20364 = ~n19072 & n20363 ;
  assign n20365 = x169 & ~n18909 ;
  assign n20366 = n18998 & ~n20365 ;
  assign n20367 = x169 & n2203 ;
  assign n20368 = ~n14684 & n20367 ;
  assign n20369 = n19314 | n20368 ;
  assign n20370 = x169 | n16705 ;
  assign n20371 = ~n19026 & n20370 ;
  assign n20372 = ~n19061 & n20371 ;
  assign n20373 = x215 | n20372 ;
  assign n20374 = n20369 | n20373 ;
  assign n20375 = ~n20366 & n20374 ;
  assign n20376 = x299 & ~n20375 ;
  assign n20377 = x169 & ~n19106 ;
  assign n20378 = n19096 | n20377 ;
  assign n20379 = ~n20376 & n20378 ;
  assign n20380 = x746 & ~n20379 ;
  assign n20381 = ~n19063 & n20370 ;
  assign n20382 = n19046 | n20381 ;
  assign n20383 = n20369 | n20382 ;
  assign n20384 = ~x215 & n20383 ;
  assign n20385 = n14577 & ~n20366 ;
  assign n20386 = n19021 | n20385 ;
  assign n20387 = n20384 | n20386 ;
  assign n20388 = x299 & n20387 ;
  assign n20389 = x169 | n18988 ;
  assign n20390 = ~n19069 & n20389 ;
  assign n20391 = x746 | n20390 ;
  assign n20392 = n20388 | n20391 ;
  assign n20393 = x39 & n20392 ;
  assign n20394 = ~n20380 & n20393 ;
  assign n20395 = n20364 | n20394 ;
  assign n20396 = ~x38 & n20395 ;
  assign n20397 = ~x746 & x947 ;
  assign n20398 = x39 | n20397 ;
  assign n20399 = n19236 & ~n20398 ;
  assign n20400 = x169 | n15070 ;
  assign n20401 = x38 & n20400 ;
  assign n20402 = ~n20399 & n20401 ;
  assign n20403 = n20396 | n20402 ;
  assign n20404 = x729 & n20403 ;
  assign n20405 = ~n19019 & n20389 ;
  assign n20406 = n20369 | n20371 ;
  assign n20407 = n18996 | n20406 ;
  assign n20408 = n19000 & ~n20365 ;
  assign n20409 = x299 & ~n20408 ;
  assign n20410 = n20407 & n20409 ;
  assign n20411 = x746 & ~n20410 ;
  assign n20412 = ~n20405 & n20411 ;
  assign n20413 = x169 | x746 ;
  assign n20414 = n14710 | n20413 ;
  assign n20415 = x39 & n20414 ;
  assign n20416 = ~n20412 & n20415 ;
  assign n20417 = x38 | n20363 ;
  assign n20418 = n20416 | n20417 ;
  assign n20419 = x169 & ~n14827 ;
  assign n20420 = ~n4810 & n20354 ;
  assign n20421 = x38 & ~n20420 ;
  assign n20422 = ~n20419 & n20421 ;
  assign n20423 = x729 | n20422 ;
  assign n20424 = n20418 & ~n20423 ;
  assign n20425 = n19157 | n20424 ;
  assign n20426 = n20404 | n20425 ;
  assign n20427 = ~x169 & n19157 ;
  assign n20428 = x57 | n20427 ;
  assign n20429 = n20426 & ~n20428 ;
  assign n20430 = x57 & x169 ;
  assign n20431 = x832 | n20430 ;
  assign n20432 = n20429 | n20431 ;
  assign n20433 = ~n20359 & n20432 ;
  assign n20434 = x730 & n18913 ;
  assign n20435 = x748 & x947 ;
  assign n20436 = n1290 & ~n20435 ;
  assign n20437 = ~n20434 & n20436 ;
  assign n20438 = x170 & ~n1290 ;
  assign n20439 = x832 & ~n20438 ;
  assign n20440 = ~n20437 & n20439 ;
  assign n20441 = x170 & n2203 ;
  assign n20442 = ~n14684 & n20441 ;
  assign n20443 = n19314 | n20442 ;
  assign n20444 = x170 | n16705 ;
  assign n20445 = ~n19063 & n20444 ;
  assign n20446 = n19046 | n20445 ;
  assign n20447 = n20443 | n20446 ;
  assign n20448 = ~x215 & n20447 ;
  assign n20449 = x170 & ~n18909 ;
  assign n20450 = n18998 & ~n20449 ;
  assign n20451 = n14577 & ~n20450 ;
  assign n20452 = n19021 | n20451 ;
  assign n20453 = n20448 | n20452 ;
  assign n20454 = x299 & n20453 ;
  assign n20455 = x170 | n18988 ;
  assign n20456 = ~x299 & n20455 ;
  assign n20457 = ~n19068 & n20456 ;
  assign n20458 = n20454 | n20457 ;
  assign n20459 = x39 & n20458 ;
  assign n20460 = x170 | n14822 ;
  assign n20461 = ~n19073 & n20460 ;
  assign n20462 = n20459 | n20461 ;
  assign n20463 = ~x38 & n20462 ;
  assign n20464 = x170 | n15070 ;
  assign n20465 = n19041 & n20464 ;
  assign n20466 = x748 | n20465 ;
  assign n20467 = n20463 | n20466 ;
  assign n20468 = ~n19102 & n20460 ;
  assign n20469 = x170 & ~n19106 ;
  assign n20470 = n19096 | n20469 ;
  assign n20471 = ~n19026 & n20444 ;
  assign n20472 = ~n19061 & n20471 ;
  assign n20473 = x215 | n20472 ;
  assign n20474 = n20443 | n20473 ;
  assign n20475 = ~n20450 & n20474 ;
  assign n20476 = x299 & ~n20475 ;
  assign n20477 = x39 & ~n20476 ;
  assign n20478 = n20470 & n20477 ;
  assign n20479 = n20468 | n20478 ;
  assign n20480 = ~x38 & n20479 ;
  assign n20481 = n19081 & n20464 ;
  assign n20482 = x748 & ~n20481 ;
  assign n20483 = ~n20480 & n20482 ;
  assign n20484 = x730 & ~n20483 ;
  assign n20485 = n20467 & n20484 ;
  assign n20486 = ~n19017 & n20460 ;
  assign n20487 = n20443 | n20471 ;
  assign n20488 = n18996 | n20487 ;
  assign n20489 = n19000 & ~n20449 ;
  assign n20490 = x299 & ~n20489 ;
  assign n20491 = n20488 & n20490 ;
  assign n20492 = ~n19018 & n20456 ;
  assign n20493 = n20491 | n20492 ;
  assign n20494 = x39 & n20493 ;
  assign n20495 = n20486 | n20494 ;
  assign n20496 = ~x38 & n20495 ;
  assign n20497 = x170 | n14827 ;
  assign n20498 = n19015 & n20497 ;
  assign n20499 = x748 & ~n20498 ;
  assign n20500 = ~n20496 & n20499 ;
  assign n20501 = x170 | x748 ;
  assign n20502 = n15382 | n20501 ;
  assign n20503 = ~x730 & n20502 ;
  assign n20504 = ~n20500 & n20503 ;
  assign n20505 = n19157 | n20504 ;
  assign n20506 = n20485 | n20505 ;
  assign n20507 = ~x170 & n19157 ;
  assign n20508 = x57 | n20507 ;
  assign n20509 = n20506 & ~n20508 ;
  assign n20510 = x57 & x170 ;
  assign n20511 = x832 | n20510 ;
  assign n20512 = n20509 | n20511 ;
  assign n20513 = ~n20440 & n20512 ;
  assign n20514 = x764 & x947 ;
  assign n20515 = n1290 & ~n20514 ;
  assign n20516 = x691 & n18913 ;
  assign n20517 = n20515 & ~n20516 ;
  assign n20518 = x171 & ~n1290 ;
  assign n20519 = x832 & ~n20518 ;
  assign n20520 = ~n20517 & n20519 ;
  assign n20521 = x171 | n14822 ;
  assign n20522 = ~x764 & n14823 ;
  assign n20523 = n19017 & ~n20522 ;
  assign n20524 = n20521 & ~n20523 ;
  assign n20525 = ~n19072 & n20524 ;
  assign n20526 = x171 & ~n18909 ;
  assign n20527 = n18998 & ~n20526 ;
  assign n20528 = x171 & n2203 ;
  assign n20529 = ~n14684 & n20528 ;
  assign n20530 = n19314 | n20529 ;
  assign n20531 = x171 | n16705 ;
  assign n20532 = ~n19026 & n20531 ;
  assign n20533 = ~n19061 & n20532 ;
  assign n20534 = x215 | n20533 ;
  assign n20535 = n20530 | n20534 ;
  assign n20536 = ~n20527 & n20535 ;
  assign n20537 = x299 & ~n20536 ;
  assign n20538 = x171 & ~n19106 ;
  assign n20539 = n19096 | n20538 ;
  assign n20540 = ~n20537 & n20539 ;
  assign n20541 = x764 & ~n20540 ;
  assign n20542 = ~n19063 & n20531 ;
  assign n20543 = n19046 | n20542 ;
  assign n20544 = n20530 | n20543 ;
  assign n20545 = ~x215 & n20544 ;
  assign n20546 = n14577 & ~n20527 ;
  assign n20547 = n19021 | n20546 ;
  assign n20548 = n20545 | n20547 ;
  assign n20549 = x299 & n20548 ;
  assign n20550 = x171 | n18988 ;
  assign n20551 = ~n19069 & n20550 ;
  assign n20552 = x764 | n20551 ;
  assign n20553 = n20549 | n20552 ;
  assign n20554 = x39 & n20553 ;
  assign n20555 = ~n20541 & n20554 ;
  assign n20556 = n20525 | n20555 ;
  assign n20557 = ~x38 & n20556 ;
  assign n20558 = ~x764 & x947 ;
  assign n20559 = x39 | n20558 ;
  assign n20560 = n19236 & ~n20559 ;
  assign n20561 = x171 | n15070 ;
  assign n20562 = x38 & n20561 ;
  assign n20563 = ~n20560 & n20562 ;
  assign n20564 = n20557 | n20563 ;
  assign n20565 = x691 & n20564 ;
  assign n20566 = ~n19019 & n20550 ;
  assign n20567 = n20530 | n20532 ;
  assign n20568 = n18996 | n20567 ;
  assign n20569 = n19000 & ~n20526 ;
  assign n20570 = x299 & ~n20569 ;
  assign n20571 = n20568 & n20570 ;
  assign n20572 = x764 & ~n20571 ;
  assign n20573 = ~n20566 & n20572 ;
  assign n20574 = x171 | x764 ;
  assign n20575 = n14710 | n20574 ;
  assign n20576 = x39 & n20575 ;
  assign n20577 = ~n20573 & n20576 ;
  assign n20578 = x38 | n20524 ;
  assign n20579 = n20577 | n20578 ;
  assign n20580 = x171 & ~n14827 ;
  assign n20581 = ~n4810 & n20515 ;
  assign n20582 = x38 & ~n20581 ;
  assign n20583 = ~n20580 & n20582 ;
  assign n20584 = x691 | n20583 ;
  assign n20585 = n20579 & ~n20584 ;
  assign n20586 = n19157 | n20585 ;
  assign n20587 = n20565 | n20586 ;
  assign n20588 = ~x171 & n19157 ;
  assign n20589 = x57 | n20588 ;
  assign n20590 = n20587 & ~n20589 ;
  assign n20591 = x57 & x171 ;
  assign n20592 = x832 | n20591 ;
  assign n20593 = n20590 | n20592 ;
  assign n20594 = ~n20520 & n20593 ;
  assign n20595 = x739 & x947 ;
  assign n20596 = n1290 & ~n20595 ;
  assign n20597 = x690 & n18913 ;
  assign n20598 = n20596 & ~n20597 ;
  assign n20599 = x172 & ~n1290 ;
  assign n20600 = x832 & ~n20599 ;
  assign n20601 = ~n20598 & n20600 ;
  assign n20602 = ( x39 & n14822 ) | ( x39 & n20595 ) | ( n14822 & n20595 ) ;
  assign n20603 = ( ~x39 & x172 ) | ( ~x39 & n14822 ) | ( x172 & n14822 ) ;
  assign n20604 = ~n20602 & n20603 ;
  assign n20605 = ~n19072 & n20604 ;
  assign n20606 = x172 & ~n18909 ;
  assign n20607 = n18998 & ~n20606 ;
  assign n20608 = x172 & n2203 ;
  assign n20609 = ~n14684 & n20608 ;
  assign n20610 = n19314 | n20609 ;
  assign n20611 = x172 | n16705 ;
  assign n20612 = ~n19026 & n20611 ;
  assign n20613 = ~n19061 & n20612 ;
  assign n20614 = x215 | n20613 ;
  assign n20615 = n20610 | n20614 ;
  assign n20616 = ~n20607 & n20615 ;
  assign n20617 = x299 & ~n20616 ;
  assign n20618 = x172 & ~n19106 ;
  assign n20619 = n19096 | n20618 ;
  assign n20620 = ~n20617 & n20619 ;
  assign n20621 = x739 & ~n20620 ;
  assign n20622 = ~n19063 & n20611 ;
  assign n20623 = n19046 | n20622 ;
  assign n20624 = n20610 | n20623 ;
  assign n20625 = ~x215 & n20624 ;
  assign n20626 = n14577 & ~n20607 ;
  assign n20627 = n19021 | n20626 ;
  assign n20628 = n20625 | n20627 ;
  assign n20629 = x299 & n20628 ;
  assign n20630 = x172 | n18988 ;
  assign n20631 = ~n19069 & n20630 ;
  assign n20632 = x739 | n20631 ;
  assign n20633 = n20629 | n20632 ;
  assign n20634 = x39 & n20633 ;
  assign n20635 = ~n20621 & n20634 ;
  assign n20636 = n20605 | n20635 ;
  assign n20637 = ~x38 & n20636 ;
  assign n20638 = ~x739 & x947 ;
  assign n20639 = x39 | n20638 ;
  assign n20640 = n19236 & ~n20639 ;
  assign n20641 = x172 | n15070 ;
  assign n20642 = x38 & n20641 ;
  assign n20643 = ~n20640 & n20642 ;
  assign n20644 = n20637 | n20643 ;
  assign n20645 = x690 & n20644 ;
  assign n20646 = ~n19019 & n20630 ;
  assign n20647 = n20610 | n20612 ;
  assign n20648 = n18996 | n20647 ;
  assign n20649 = n19000 & ~n20606 ;
  assign n20650 = x299 & ~n20649 ;
  assign n20651 = n20648 & n20650 ;
  assign n20652 = x739 & ~n20651 ;
  assign n20653 = ~n20646 & n20652 ;
  assign n20654 = x172 | x739 ;
  assign n20655 = n14710 | n20654 ;
  assign n20656 = x39 & n20655 ;
  assign n20657 = ~n20653 & n20656 ;
  assign n20658 = x38 | n20604 ;
  assign n20659 = n20657 | n20658 ;
  assign n20660 = x172 & ~n14827 ;
  assign n20661 = ~n4810 & n20596 ;
  assign n20662 = x38 & ~n20661 ;
  assign n20663 = ~n20660 & n20662 ;
  assign n20664 = x690 | n20663 ;
  assign n20665 = n20659 & ~n20664 ;
  assign n20666 = n19157 | n20665 ;
  assign n20667 = n20645 | n20666 ;
  assign n20668 = ~x172 & n19157 ;
  assign n20669 = x57 | n20668 ;
  assign n20670 = n20667 & ~n20669 ;
  assign n20671 = x57 & x172 ;
  assign n20672 = x832 | n20671 ;
  assign n20673 = n20670 | n20672 ;
  assign n20674 = ~n20601 & n20673 ;
  assign n20675 = x173 | n14834 ;
  assign n20676 = n15414 & n20675 ;
  assign n20677 = x723 | n2032 ;
  assign n20678 = ~n20675 & n20677 ;
  assign n20679 = x173 & n16323 ;
  assign n20680 = x38 | n20679 ;
  assign n20681 = ~n2032 & n20680 ;
  assign n20682 = x173 | n16319 ;
  assign n20683 = ~n20681 & n20682 ;
  assign n20684 = x173 | n15070 ;
  assign n20685 = n15375 & n20684 ;
  assign n20686 = x723 | n20685 ;
  assign n20687 = n20683 | n20686 ;
  assign n20688 = ~n20678 & n20687 ;
  assign n20689 = ~x778 & n20688 ;
  assign n20690 = ( x625 & x1153 ) | ( x625 & n20675 ) | ( x1153 & n20675 ) ;
  assign n20691 = ( ~x625 & x1153 ) | ( ~x625 & n20688 ) | ( x1153 & n20688 ) ;
  assign n20692 = n20690 & n20691 ;
  assign n20693 = ( x625 & x1153 ) | ( x625 & ~n20675 ) | ( x1153 & ~n20675 ) ;
  assign n20694 = ( x625 & ~x1153 ) | ( x625 & n20688 ) | ( ~x1153 & n20688 ) ;
  assign n20695 = ~n20693 & n20694 ;
  assign n20696 = n20692 | n20695 ;
  assign n20697 = x778 & n20696 ;
  assign n20698 = n20689 | n20697 ;
  assign n20699 = ~n15400 & n20698 ;
  assign n20700 = n15400 & n20675 ;
  assign n20701 = n20699 | n20700 ;
  assign n20702 = n15407 | n20701 ;
  assign n20703 = n15407 & ~n20675 ;
  assign n20704 = n20702 & ~n20703 ;
  assign n20705 = ~n15414 & n20704 ;
  assign n20706 = n20676 | n20705 ;
  assign n20707 = n15421 | n20706 ;
  assign n20708 = n15421 & ~n20675 ;
  assign n20709 = n20707 & ~n20708 ;
  assign n20710 = ~x792 & n20709 ;
  assign n20711 = ( x628 & x1156 ) | ( x628 & n20675 ) | ( x1156 & n20675 ) ;
  assign n20712 = ( ~x628 & x1156 ) | ( ~x628 & n20709 ) | ( x1156 & n20709 ) ;
  assign n20713 = n20711 & n20712 ;
  assign n20714 = ( x628 & x1156 ) | ( x628 & ~n20675 ) | ( x1156 & ~n20675 ) ;
  assign n20715 = ( x628 & ~x1156 ) | ( x628 & n20709 ) | ( ~x1156 & n20709 ) ;
  assign n20716 = ~n20714 & n20715 ;
  assign n20717 = n20713 | n20716 ;
  assign n20718 = x792 & n20717 ;
  assign n20719 = n20710 | n20718 ;
  assign n20720 = x787 | n20719 ;
  assign n20721 = x647 & n20719 ;
  assign n20722 = ~x647 & n20675 ;
  assign n20723 = n20721 | n20722 ;
  assign n20724 = ( ~x787 & x1157 ) | ( ~x787 & n20723 ) | ( x1157 & n20723 ) ;
  assign n20725 = ~x647 & n20719 ;
  assign n20726 = x647 & n20675 ;
  assign n20727 = n20725 | n20726 ;
  assign n20728 = ( x787 & x1157 ) | ( x787 & ~n20727 ) | ( x1157 & ~n20727 ) ;
  assign n20729 = ~n20724 & n20728 ;
  assign n20730 = n20720 & ~n20729 ;
  assign n20731 = x644 | n20730 ;
  assign n20732 = x715 & n20731 ;
  assign n20733 = x173 & n2032 ;
  assign n20734 = x173 | n14936 ;
  assign n20735 = x745 & n20734 ;
  assign n20736 = x173 & ~n14933 ;
  assign n20737 = x173 | x745 ;
  assign n20738 = n15063 & ~n20737 ;
  assign n20739 = n20736 | n20738 ;
  assign n20740 = n20735 | n20739 ;
  assign n20741 = ~x38 & n20740 ;
  assign n20742 = ~x745 & n15072 ;
  assign n20743 = x38 & n20684 ;
  assign n20744 = ~n20742 & n20743 ;
  assign n20745 = n20741 | n20744 ;
  assign n20746 = ~n2032 & n20745 ;
  assign n20747 = n20733 | n20746 ;
  assign n20748 = ~n15082 & n20747 ;
  assign n20749 = n15082 & n20675 ;
  assign n20750 = n20748 | n20749 ;
  assign n20751 = ~x785 & n20750 ;
  assign n20752 = ~n15088 & n20675 ;
  assign n20753 = x609 & n20748 ;
  assign n20754 = n20752 | n20753 ;
  assign n20755 = x1155 & n20754 ;
  assign n20756 = n15094 & n20675 ;
  assign n20757 = ~x609 & n20748 ;
  assign n20758 = n20756 | n20757 ;
  assign n20759 = ~x1155 & n20758 ;
  assign n20760 = n20755 | n20759 ;
  assign n20761 = x785 & n20760 ;
  assign n20762 = n20751 | n20761 ;
  assign n20763 = ~x781 & n20762 ;
  assign n20764 = ( x618 & x1154 ) | ( x618 & n20675 ) | ( x1154 & n20675 ) ;
  assign n20765 = ( ~x618 & x1154 ) | ( ~x618 & n20762 ) | ( x1154 & n20762 ) ;
  assign n20766 = n20764 & n20765 ;
  assign n20767 = ( x618 & x1154 ) | ( x618 & ~n20675 ) | ( x1154 & ~n20675 ) ;
  assign n20768 = ( x618 & ~x1154 ) | ( x618 & n20762 ) | ( ~x1154 & n20762 ) ;
  assign n20769 = ~n20767 & n20768 ;
  assign n20770 = n20766 | n20769 ;
  assign n20771 = x781 & n20770 ;
  assign n20772 = n20763 | n20771 ;
  assign n20773 = ~x789 & n20772 ;
  assign n20774 = ( x619 & x1159 ) | ( x619 & n20675 ) | ( x1159 & n20675 ) ;
  assign n20775 = ( ~x619 & x1159 ) | ( ~x619 & n20772 ) | ( x1159 & n20772 ) ;
  assign n20776 = n20774 & n20775 ;
  assign n20777 = ( x619 & x1159 ) | ( x619 & ~n20675 ) | ( x1159 & ~n20675 ) ;
  assign n20778 = ( x619 & ~x1159 ) | ( x619 & n20772 ) | ( ~x1159 & n20772 ) ;
  assign n20779 = ~n20777 & n20778 ;
  assign n20780 = n20776 | n20779 ;
  assign n20781 = x789 & n20780 ;
  assign n20782 = n20773 | n20781 ;
  assign n20783 = ~x788 & n20782 ;
  assign n20784 = ( x626 & x1158 ) | ( x626 & n20675 ) | ( x1158 & n20675 ) ;
  assign n20785 = ( ~x1158 & n20782 ) | ( ~x1158 & n20784 ) | ( n20782 & n20784 ) ;
  assign n20786 = ( ~x626 & n20784 ) | ( ~x626 & n20785 ) | ( n20784 & n20785 ) ;
  assign n20787 = x788 & n20786 ;
  assign n20788 = n20783 | n20787 ;
  assign n20789 = n15134 | n20788 ;
  assign n20790 = n15134 & ~n20675 ;
  assign n20791 = n20789 & ~n20790 ;
  assign n20792 = n15141 | n20791 ;
  assign n20793 = n15141 & ~n20675 ;
  assign n20794 = n20792 & ~n20793 ;
  assign n20795 = ( x644 & x715 ) | ( x644 & ~n20794 ) | ( x715 & ~n20794 ) ;
  assign n20796 = ( x644 & ~x715 ) | ( x644 & n20675 ) | ( ~x715 & n20675 ) ;
  assign n20797 = ~n20795 & n20796 ;
  assign n20798 = x1160 & ~n20797 ;
  assign n20799 = ~n20732 & n20798 ;
  assign n20800 = ( x644 & x715 ) | ( x644 & n20794 ) | ( x715 & n20794 ) ;
  assign n20801 = ( ~x644 & x715 ) | ( ~x644 & n20675 ) | ( x715 & n20675 ) ;
  assign n20802 = n20800 & n20801 ;
  assign n20803 = x1160 | n20802 ;
  assign n20804 = ( x644 & x715 ) | ( x644 & ~n20730 ) | ( x715 & ~n20730 ) ;
  assign n20805 = n18610 & n20791 ;
  assign n20806 = n15139 & n20727 ;
  assign n20807 = n15138 & n20723 ;
  assign n20808 = n20806 | n20807 ;
  assign n20809 = n20805 | n20808 ;
  assign n20810 = x787 & n20809 ;
  assign n20811 = n18621 & n20788 ;
  assign n20812 = ( x629 & n20716 ) | ( x629 & n20811 ) | ( n20716 & n20811 ) ;
  assign n20813 = ( ~x629 & n20713 ) | ( ~x629 & n20811 ) | ( n20713 & n20811 ) ;
  assign n20814 = n20812 | n20813 ;
  assign n20815 = x792 & n20814 ;
  assign n20816 = x648 & ~n20779 ;
  assign n20817 = ( x619 & x1159 ) | ( x619 & n20704 ) | ( x1159 & n20704 ) ;
  assign n20818 = x627 | n20766 ;
  assign n20819 = ( x618 & x1154 ) | ( x618 & ~n20701 ) | ( x1154 & ~n20701 ) ;
  assign n20820 = x660 | n20755 ;
  assign n20821 = ( x609 & x1155 ) | ( x609 & ~n20698 ) | ( x1155 & ~n20698 ) ;
  assign n20822 = x608 | n20692 ;
  assign n20823 = ( x625 & x1153 ) | ( x625 & ~n20747 ) | ( x1153 & ~n20747 ) ;
  assign n20824 = x723 & ~n20745 ;
  assign n20825 = ( x173 & ~x745 ) | ( x173 & n15797 ) | ( ~x745 & n15797 ) ;
  assign n20826 = ( x173 & x745 ) | ( x173 & n15872 ) | ( x745 & n15872 ) ;
  assign n20827 = n20825 & ~n20826 ;
  assign n20828 = x39 & ~n20827 ;
  assign n20829 = ( x173 & ~x745 ) | ( x173 & n15583 ) | ( ~x745 & n15583 ) ;
  assign n20830 = ( x173 & x745 ) | ( x173 & n15699 ) | ( x745 & n15699 ) ;
  assign n20831 = ~n20829 & n20830 ;
  assign n20832 = n20828 & ~n20831 ;
  assign n20833 = ( ~x173 & x745 ) | ( ~x173 & n15887 ) | ( x745 & n15887 ) ;
  assign n20834 = ( x173 & x745 ) | ( x173 & ~n15891 ) | ( x745 & ~n15891 ) ;
  assign n20835 = n20833 & n20834 ;
  assign n20836 = ( ~x173 & x745 ) | ( ~x173 & n15894 ) | ( x745 & n15894 ) ;
  assign n20837 = ( x173 & x745 ) | ( x173 & ~n15897 ) | ( x745 & ~n15897 ) ;
  assign n20838 = n20836 | n20837 ;
  assign n20839 = ~n20835 & n20838 ;
  assign n20840 = x39 | n20839 ;
  assign n20841 = ~x38 & n20840 ;
  assign n20842 = ~n20832 & n20841 ;
  assign n20843 = x745 | n15758 ;
  assign n20844 = n17573 & n20843 ;
  assign n20845 = x173 | n20844 ;
  assign n20846 = ~x745 & n14840 ;
  assign n20847 = n15529 | n20846 ;
  assign n20848 = x173 & n20847 ;
  assign n20849 = ~n4810 & n20848 ;
  assign n20850 = x38 & ~n20849 ;
  assign n20851 = n20845 & n20850 ;
  assign n20852 = x723 | n20851 ;
  assign n20853 = n20842 | n20852 ;
  assign n20854 = ~n2032 & n20853 ;
  assign n20855 = ~n20824 & n20854 ;
  assign n20856 = n20733 | n20855 ;
  assign n20857 = ( x625 & ~x1153 ) | ( x625 & n20856 ) | ( ~x1153 & n20856 ) ;
  assign n20858 = ~n20823 & n20857 ;
  assign n20859 = n20822 | n20858 ;
  assign n20860 = x608 & ~n20695 ;
  assign n20861 = ( x625 & x1153 ) | ( x625 & n20747 ) | ( x1153 & n20747 ) ;
  assign n20862 = ( ~x625 & x1153 ) | ( ~x625 & n20856 ) | ( x1153 & n20856 ) ;
  assign n20863 = n20861 & n20862 ;
  assign n20864 = n20860 & ~n20863 ;
  assign n20865 = n20859 & ~n20864 ;
  assign n20866 = x778 & ~n20865 ;
  assign n20867 = x778 | n20856 ;
  assign n20868 = ~n20866 & n20867 ;
  assign n20869 = ( x609 & ~x1155 ) | ( x609 & n20868 ) | ( ~x1155 & n20868 ) ;
  assign n20870 = ~n20821 & n20869 ;
  assign n20871 = n20820 | n20870 ;
  assign n20872 = x660 & ~n20759 ;
  assign n20873 = ( x609 & x1155 ) | ( x609 & n20698 ) | ( x1155 & n20698 ) ;
  assign n20874 = ( ~x609 & x1155 ) | ( ~x609 & n20868 ) | ( x1155 & n20868 ) ;
  assign n20875 = n20873 & n20874 ;
  assign n20876 = n20872 & ~n20875 ;
  assign n20877 = n20871 & ~n20876 ;
  assign n20878 = x785 & ~n20877 ;
  assign n20879 = x785 | n20868 ;
  assign n20880 = ~n20878 & n20879 ;
  assign n20881 = ( x618 & ~x1154 ) | ( x618 & n20880 ) | ( ~x1154 & n20880 ) ;
  assign n20882 = ~n20819 & n20881 ;
  assign n20883 = n20818 | n20882 ;
  assign n20884 = x627 & ~n20769 ;
  assign n20885 = ( x618 & x1154 ) | ( x618 & n20701 ) | ( x1154 & n20701 ) ;
  assign n20886 = ( ~x618 & x1154 ) | ( ~x618 & n20880 ) | ( x1154 & n20880 ) ;
  assign n20887 = n20885 & n20886 ;
  assign n20888 = n20884 & ~n20887 ;
  assign n20889 = n20883 & ~n20888 ;
  assign n20890 = x781 & ~n20889 ;
  assign n20891 = x781 | n20880 ;
  assign n20892 = ~n20890 & n20891 ;
  assign n20893 = ( ~x619 & x1159 ) | ( ~x619 & n20892 ) | ( x1159 & n20892 ) ;
  assign n20894 = n20817 & n20893 ;
  assign n20895 = n20816 & ~n20894 ;
  assign n20896 = x648 | n20776 ;
  assign n20897 = ( x619 & x1159 ) | ( x619 & ~n20704 ) | ( x1159 & ~n20704 ) ;
  assign n20898 = ( x619 & ~x1159 ) | ( x619 & n20892 ) | ( ~x1159 & n20892 ) ;
  assign n20899 = ~n20897 & n20898 ;
  assign n20900 = n20896 | n20899 ;
  assign n20901 = x789 & n20900 ;
  assign n20902 = ~n20895 & n20901 ;
  assign n20903 = ~x789 & n20892 ;
  assign n20904 = n16177 | n20903 ;
  assign n20905 = n20902 | n20904 ;
  assign n20906 = n16115 & ~n20706 ;
  assign n20907 = n15420 & ~n20786 ;
  assign n20908 = n20906 | n20907 ;
  assign n20909 = x788 & n20908 ;
  assign n20910 = n18434 | n20909 ;
  assign n20911 = n20905 & ~n20910 ;
  assign n20912 = n20815 | n20911 ;
  assign n20913 = ~n18431 & n20912 ;
  assign n20914 = n20810 | n20913 ;
  assign n20915 = ( x644 & ~x715 ) | ( x644 & n20914 ) | ( ~x715 & n20914 ) ;
  assign n20916 = ~n20804 & n20915 ;
  assign n20917 = n20803 | n20916 ;
  assign n20918 = ~n20799 & n20917 ;
  assign n20919 = x790 & ~n20918 ;
  assign n20920 = x644 & n20798 ;
  assign n20921 = x790 & ~n20920 ;
  assign n20922 = n20914 | n20921 ;
  assign n20923 = ~n20919 & n20922 ;
  assign n20924 = ( ~x832 & n6785 ) | ( ~x832 & n20923 ) | ( n6785 & n20923 ) ;
  assign n20925 = ( ~x173 & x832 ) | ( ~x173 & n6785 ) | ( x832 & n6785 ) ;
  assign n20926 = n20924 & ~n20925 ;
  assign n20927 = x173 | n1290 ;
  assign n20928 = ~n20846 & n20927 ;
  assign n20929 = n16060 | n20928 ;
  assign n20930 = ~x785 & n20929 ;
  assign n20931 = ~n15094 & n20846 ;
  assign n20932 = n20929 | n20931 ;
  assign n20933 = x1155 & n20932 ;
  assign n20934 = ~x1155 & n20927 ;
  assign n20935 = ~n20931 & n20934 ;
  assign n20936 = n20933 | n20935 ;
  assign n20937 = x785 & n20936 ;
  assign n20938 = n20930 | n20937 ;
  assign n20939 = ~x781 & n20938 ;
  assign n20940 = n16075 | n20938 ;
  assign n20941 = x1154 & n20940 ;
  assign n20942 = n16078 | n20938 ;
  assign n20943 = ~x1154 & n20942 ;
  assign n20944 = n20941 | n20943 ;
  assign n20945 = x781 & n20944 ;
  assign n20946 = n20939 | n20945 ;
  assign n20947 = ~x789 & n20946 ;
  assign n20948 = ~x619 & n1290 ;
  assign n20949 = n20946 | n20948 ;
  assign n20950 = x1159 & n20949 ;
  assign n20951 = x619 & n1290 ;
  assign n20952 = n20946 | n20951 ;
  assign n20953 = ~x1159 & n20952 ;
  assign n20954 = n20950 | n20953 ;
  assign n20955 = x789 & n20954 ;
  assign n20956 = n20947 | n20955 ;
  assign n20957 = ~x788 & n20956 ;
  assign n20958 = ( x626 & x1158 ) | ( x626 & n20927 ) | ( x1158 & n20927 ) ;
  assign n20959 = ( ~x1158 & n20956 ) | ( ~x1158 & n20958 ) | ( n20956 & n20958 ) ;
  assign n20960 = ( ~x626 & n20958 ) | ( ~x626 & n20959 ) | ( n20958 & n20959 ) ;
  assign n20961 = x788 & n20960 ;
  assign n20962 = n20957 | n20961 ;
  assign n20963 = n15134 | n20962 ;
  assign n20964 = n15134 & ~n20927 ;
  assign n20965 = n20963 & ~n20964 ;
  assign n20966 = n18610 & n20965 ;
  assign n20967 = ( x647 & x1157 ) | ( x647 & ~n20927 ) | ( x1157 & ~n20927 ) ;
  assign n20968 = ~x723 & n15202 ;
  assign n20969 = n20927 & ~n20968 ;
  assign n20970 = x778 | n20969 ;
  assign n20971 = ~x625 & n20968 ;
  assign n20972 = n20969 | n20971 ;
  assign n20973 = x1153 & n20972 ;
  assign n20974 = ~x1153 & n20927 ;
  assign n20975 = ~n20971 & n20974 ;
  assign n20976 = x778 & ~n20975 ;
  assign n20977 = ~n20973 & n20976 ;
  assign n20978 = n20970 & ~n20977 ;
  assign n20979 = n16043 | n20978 ;
  assign n20980 = n16045 | n20979 ;
  assign n20981 = n16047 | n20980 ;
  assign n20982 = n16049 | n20981 ;
  assign n20983 = n16055 | n20982 ;
  assign n20984 = ( x647 & ~x1157 ) | ( x647 & n20983 ) | ( ~x1157 & n20983 ) ;
  assign n20985 = ~n20967 & n20984 ;
  assign n20986 = x630 & n20985 ;
  assign n20987 = x647 & n20983 ;
  assign n20988 = ~x647 & n20927 ;
  assign n20989 = n20987 | n20988 ;
  assign n20990 = n15138 & n20989 ;
  assign n20991 = n20986 | n20990 ;
  assign n20992 = n20966 | n20991 ;
  assign n20993 = x787 & n20992 ;
  assign n20994 = n16115 & ~n20981 ;
  assign n20995 = n15420 & ~n20960 ;
  assign n20996 = n20994 | n20995 ;
  assign n20997 = x788 & n20996 ;
  assign n20998 = x648 & ~n20953 ;
  assign n20999 = ( x619 & x1159 ) | ( x619 & n20980 ) | ( x1159 & n20980 ) ;
  assign n21000 = x627 | n20941 ;
  assign n21001 = ( x618 & x1154 ) | ( x618 & ~n20979 ) | ( x1154 & ~n20979 ) ;
  assign n21002 = x660 | n20933 ;
  assign n21003 = ( x609 & x1155 ) | ( x609 & ~n20978 ) | ( x1155 & ~n20978 ) ;
  assign n21004 = n14839 | n20969 ;
  assign n21005 = x625 & ~n21004 ;
  assign n21006 = n20928 & n21004 ;
  assign n21007 = n21005 | n21006 ;
  assign n21008 = n20974 & n21007 ;
  assign n21009 = x608 | n20973 ;
  assign n21010 = n21008 | n21009 ;
  assign n21011 = x1153 & n20928 ;
  assign n21012 = ~n21005 & n21011 ;
  assign n21013 = x608 & ~n20975 ;
  assign n21014 = ~n21012 & n21013 ;
  assign n21015 = n21010 & ~n21014 ;
  assign n21016 = x778 & ~n21015 ;
  assign n21017 = x778 | n21006 ;
  assign n21018 = ~n21016 & n21017 ;
  assign n21019 = ( x609 & ~x1155 ) | ( x609 & n21018 ) | ( ~x1155 & n21018 ) ;
  assign n21020 = ~n21003 & n21019 ;
  assign n21021 = n21002 | n21020 ;
  assign n21022 = x660 & ~n20935 ;
  assign n21023 = ( x609 & x1155 ) | ( x609 & n20978 ) | ( x1155 & n20978 ) ;
  assign n21024 = ( ~x609 & x1155 ) | ( ~x609 & n21018 ) | ( x1155 & n21018 ) ;
  assign n21025 = n21023 & n21024 ;
  assign n21026 = n21022 & ~n21025 ;
  assign n21027 = n21021 & ~n21026 ;
  assign n21028 = x785 & ~n21027 ;
  assign n21029 = x785 | n21018 ;
  assign n21030 = ~n21028 & n21029 ;
  assign n21031 = ( x618 & ~x1154 ) | ( x618 & n21030 ) | ( ~x1154 & n21030 ) ;
  assign n21032 = ~n21001 & n21031 ;
  assign n21033 = n21000 | n21032 ;
  assign n21034 = x627 & ~n20943 ;
  assign n21035 = ( x618 & x1154 ) | ( x618 & n20979 ) | ( x1154 & n20979 ) ;
  assign n21036 = ( ~x618 & x1154 ) | ( ~x618 & n21030 ) | ( x1154 & n21030 ) ;
  assign n21037 = n21035 & n21036 ;
  assign n21038 = n21034 & ~n21037 ;
  assign n21039 = n21033 & ~n21038 ;
  assign n21040 = x781 & ~n21039 ;
  assign n21041 = x781 | n21030 ;
  assign n21042 = ~n21040 & n21041 ;
  assign n21043 = ( ~x619 & x1159 ) | ( ~x619 & n21042 ) | ( x1159 & n21042 ) ;
  assign n21044 = n20999 & n21043 ;
  assign n21045 = n20998 & ~n21044 ;
  assign n21046 = x648 | n20950 ;
  assign n21047 = ( x619 & x1159 ) | ( x619 & ~n20980 ) | ( x1159 & ~n20980 ) ;
  assign n21048 = ( x619 & ~x1159 ) | ( x619 & n21042 ) | ( ~x1159 & n21042 ) ;
  assign n21049 = ~n21047 & n21048 ;
  assign n21050 = n21046 | n21049 ;
  assign n21051 = x789 & n21050 ;
  assign n21052 = ~n21045 & n21051 ;
  assign n21053 = ~x789 & n21042 ;
  assign n21054 = n16177 | n21053 ;
  assign n21055 = n21052 | n21054 ;
  assign n21056 = ~n20997 & n21055 ;
  assign n21057 = n18434 | n21056 ;
  assign n21058 = n16650 | n20982 ;
  assign n21059 = n16051 & ~n20962 ;
  assign n21060 = n21058 & ~n21059 ;
  assign n21061 = ( x629 & ~x792 ) | ( x629 & n21060 ) | ( ~x792 & n21060 ) ;
  assign n21062 = n16052 & ~n20962 ;
  assign n21063 = n16643 & ~n20982 ;
  assign n21064 = n21062 | n21063 ;
  assign n21065 = ( x629 & x792 ) | ( x629 & n21064 ) | ( x792 & n21064 ) ;
  assign n21066 = ~n21061 & n21065 ;
  assign n21067 = n18431 | n21066 ;
  assign n21068 = n21057 & ~n21067 ;
  assign n21069 = n20993 | n21068 ;
  assign n21070 = ( x790 & x832 ) | ( x790 & n21069 ) | ( x832 & n21069 ) ;
  assign n21071 = n15141 | n20965 ;
  assign n21072 = n15141 & ~n20927 ;
  assign n21073 = n21071 & ~n21072 ;
  assign n21074 = ( x644 & x715 ) | ( x644 & ~n21073 ) | ( x715 & ~n21073 ) ;
  assign n21075 = ( x644 & ~x715 ) | ( x644 & n20927 ) | ( ~x715 & n20927 ) ;
  assign n21076 = ~n21074 & n21075 ;
  assign n21077 = x1160 & ~n21076 ;
  assign n21078 = ~x787 & n20983 ;
  assign n21079 = x1157 & n20989 ;
  assign n21080 = n20985 | n21079 ;
  assign n21081 = x787 & n21080 ;
  assign n21082 = n21078 | n21081 ;
  assign n21083 = ( x644 & x715 ) | ( x644 & n21082 ) | ( x715 & n21082 ) ;
  assign n21084 = ( ~x644 & x715 ) | ( ~x644 & n21069 ) | ( x715 & n21069 ) ;
  assign n21085 = n21083 & n21084 ;
  assign n21086 = n21077 & ~n21085 ;
  assign n21087 = ( x644 & x715 ) | ( x644 & n21073 ) | ( x715 & n21073 ) ;
  assign n21088 = ( ~x644 & x715 ) | ( ~x644 & n20927 ) | ( x715 & n20927 ) ;
  assign n21089 = n21087 & n21088 ;
  assign n21090 = x1160 | n21089 ;
  assign n21091 = ( x644 & x715 ) | ( x644 & ~n21082 ) | ( x715 & ~n21082 ) ;
  assign n21092 = ( x644 & ~x715 ) | ( x644 & n21069 ) | ( ~x715 & n21069 ) ;
  assign n21093 = ~n21091 & n21092 ;
  assign n21094 = n21090 | n21093 ;
  assign n21095 = ~n21086 & n21094 ;
  assign n21096 = ( ~x790 & x832 ) | ( ~x790 & n21095 ) | ( x832 & n21095 ) ;
  assign n21097 = n21070 & n21096 ;
  assign n21098 = n20926 | n21097 ;
  assign n21099 = ( x174 & x619 ) | ( x174 & x1159 ) | ( x619 & x1159 ) ;
  assign n21100 = x619 & x1159 ;
  assign n21101 = ( ~n14834 & n21099 ) | ( ~n14834 & n21100 ) | ( n21099 & n21100 ) ;
  assign n21102 = ( x174 & x618 ) | ( x174 & x1154 ) | ( x618 & x1154 ) ;
  assign n21103 = ( ~n14834 & n18246 ) | ( ~n14834 & n21102 ) | ( n18246 & n21102 ) ;
  assign n21104 = ( x174 & x609 ) | ( x174 & x1155 ) | ( x609 & x1155 ) ;
  assign n21105 = ( ~n14834 & n18136 ) | ( ~n14834 & n21104 ) | ( n18136 & n21104 ) ;
  assign n21106 = x759 & ~n15061 ;
  assign n21107 = x39 & n21106 ;
  assign n21108 = ( x39 & ~n19459 ) | ( x39 & n21107 ) | ( ~n19459 & n21107 ) ;
  assign n21109 = ( x39 & x759 ) | ( x39 & n14956 ) | ( x759 & n14956 ) ;
  assign n21110 = ( x39 & ~x759 ) | ( x39 & n14822 ) | ( ~x759 & n14822 ) ;
  assign n21111 = n21109 | n21110 ;
  assign n21112 = x174 & ~n21111 ;
  assign n21113 = ( x174 & n21108 ) | ( x174 & n21112 ) | ( n21108 & n21112 ) ;
  assign n21114 = x603 & x759 ;
  assign n21115 = ~n14838 & n21114 ;
  assign n21116 = n15070 & ~n21115 ;
  assign n21117 = x38 & x174 ;
  assign n21118 = ( x38 & n15070 ) | ( x38 & n21117 ) | ( n15070 & n21117 ) ;
  assign n21119 = ~n21116 & n21118 ;
  assign n21120 = ~x174 & x759 ;
  assign n21121 = ~n14908 & n21120 ;
  assign n21122 = n14932 & n21121 ;
  assign n21123 = ~x38 & n21122 ;
  assign n21124 = n21119 | n21123 ;
  assign n21125 = ~n2032 & n21124 ;
  assign n21126 = x38 & ~n21119 ;
  assign n21127 = n2032 | n21126 ;
  assign n21128 = ( n21113 & n21125 ) | ( n21113 & ~n21127 ) | ( n21125 & ~n21127 ) ;
  assign n21129 = ~x174 & n15082 ;
  assign n21130 = ( n14834 & n15082 ) | ( n14834 & n21129 ) | ( n15082 & n21129 ) ;
  assign n21131 = x174 & n1924 ;
  assign n21132 = ( x174 & n2031 ) | ( x174 & n21131 ) | ( n2031 & n21131 ) ;
  assign n21133 = n15082 | n21132 ;
  assign n21134 = ~n21130 & n21133 ;
  assign n21135 = ( ~x609 & x1155 ) | ( ~x609 & n21134 ) | ( x1155 & n21134 ) ;
  assign n21136 = ( x609 & ~x1155 ) | ( x609 & n21130 ) | ( ~x1155 & n21130 ) ;
  assign n21137 = ( n21128 & n21135 ) | ( n21128 & ~n21136 ) | ( n21135 & ~n21136 ) ;
  assign n21138 = n21105 & n21137 ;
  assign n21139 = ( ~x174 & x609 ) | ( ~x174 & x1155 ) | ( x609 & x1155 ) ;
  assign n21140 = ( n14834 & n18085 ) | ( n14834 & n21139 ) | ( n18085 & n21139 ) ;
  assign n21141 = ( x609 & ~x1155 ) | ( x609 & n21134 ) | ( ~x1155 & n21134 ) ;
  assign n21142 = ( ~x609 & x1155 ) | ( ~x609 & n21130 ) | ( x1155 & n21130 ) ;
  assign n21143 = ( n21128 & n21141 ) | ( n21128 & ~n21142 ) | ( n21141 & ~n21142 ) ;
  assign n21144 = ~n21140 & n21143 ;
  assign n21145 = n21138 | n21144 ;
  assign n21146 = ~x785 & n21134 ;
  assign n21147 = x785 | n21130 ;
  assign n21148 = ( n21128 & n21146 ) | ( n21128 & ~n21147 ) | ( n21146 & ~n21147 ) ;
  assign n21149 = x785 | n21148 ;
  assign n21150 = ( ~x618 & x1154 ) | ( ~x618 & n21149 ) | ( x1154 & n21149 ) ;
  assign n21151 = ( ~x618 & x1154 ) | ( ~x618 & n21148 ) | ( x1154 & n21148 ) ;
  assign n21152 = ( n21145 & n21150 ) | ( n21145 & n21151 ) | ( n21150 & n21151 ) ;
  assign n21153 = n21103 & n21152 ;
  assign n21154 = ( ~x174 & x618 ) | ( ~x174 & x1154 ) | ( x618 & x1154 ) ;
  assign n21155 = ( n14834 & n18247 ) | ( n14834 & n21154 ) | ( n18247 & n21154 ) ;
  assign n21156 = ( x618 & ~x1154 ) | ( x618 & n21149 ) | ( ~x1154 & n21149 ) ;
  assign n21157 = ( x618 & ~x1154 ) | ( x618 & n21148 ) | ( ~x1154 & n21148 ) ;
  assign n21158 = ( n21145 & n21156 ) | ( n21145 & n21157 ) | ( n21156 & n21157 ) ;
  assign n21159 = ~n21155 & n21158 ;
  assign n21160 = n21153 | n21159 ;
  assign n21161 = ~x781 & n21149 ;
  assign n21162 = ~x781 & n21148 ;
  assign n21163 = ( n21145 & n21161 ) | ( n21145 & n21162 ) | ( n21161 & n21162 ) ;
  assign n21164 = x781 | n21163 ;
  assign n21165 = ( ~x619 & x1159 ) | ( ~x619 & n21164 ) | ( x1159 & n21164 ) ;
  assign n21166 = ( ~x619 & x1159 ) | ( ~x619 & n21163 ) | ( x1159 & n21163 ) ;
  assign n21167 = ( n21160 & n21165 ) | ( n21160 & n21166 ) | ( n21165 & n21166 ) ;
  assign n21168 = n21101 & n21167 ;
  assign n21169 = ( ~x174 & x619 ) | ( ~x174 & x1159 ) | ( x619 & x1159 ) ;
  assign n21170 = x619 | x1159 ;
  assign n21171 = ( n14834 & n21169 ) | ( n14834 & n21170 ) | ( n21169 & n21170 ) ;
  assign n21172 = ( x619 & ~x1159 ) | ( x619 & n21164 ) | ( ~x1159 & n21164 ) ;
  assign n21173 = ( x619 & ~x1159 ) | ( x619 & n21163 ) | ( ~x1159 & n21163 ) ;
  assign n21174 = ( n21160 & n21172 ) | ( n21160 & n21173 ) | ( n21172 & n21173 ) ;
  assign n21175 = ~n21171 & n21174 ;
  assign n21176 = n21168 | n21175 ;
  assign n21177 = ~x789 & n21164 ;
  assign n21178 = ~x789 & n21163 ;
  assign n21179 = ( n21160 & n21177 ) | ( n21160 & n21178 ) | ( n21177 & n21178 ) ;
  assign n21180 = x789 | n21179 ;
  assign n21181 = ~n16176 & n21180 ;
  assign n21182 = ~n16176 & n21179 ;
  assign n21183 = ( n21176 & n21181 ) | ( n21176 & n21182 ) | ( n21181 & n21182 ) ;
  assign n21184 = ~x174 & n15141 ;
  assign n21185 = ( n14834 & n15141 ) | ( n14834 & n21184 ) | ( n15141 & n21184 ) ;
  assign n21186 = x174 & n16176 ;
  assign n21187 = ~n14834 & n21186 ;
  assign n21188 = ~n15134 & n21187 ;
  assign n21189 = x174 & n15134 ;
  assign n21190 = ~n14834 & n21189 ;
  assign n21191 = n21188 | n21190 ;
  assign n21192 = n15141 | n21191 ;
  assign n21193 = ~n21185 & n21192 ;
  assign n21194 = ( x644 & x715 ) | ( x644 & n21193 ) | ( x715 & n21193 ) ;
  assign n21195 = ~x644 & x715 ;
  assign n21196 = ( x174 & ~x644 ) | ( x174 & x715 ) | ( ~x644 & x715 ) ;
  assign n21197 = ( ~n14834 & n21195 ) | ( ~n14834 & n21196 ) | ( n21195 & n21196 ) ;
  assign n21198 = n21194 & n21197 ;
  assign n21199 = x1160 | n21198 ;
  assign n21200 = n15134 & ~n21190 ;
  assign n21201 = ~n15141 & n21200 ;
  assign n21202 = n21185 | n21201 ;
  assign n21203 = ( x644 & x715 ) | ( x644 & ~n21202 ) | ( x715 & ~n21202 ) ;
  assign n21204 = n21197 & n21203 ;
  assign n21205 = x1160 | n21204 ;
  assign n21206 = ( n21183 & n21199 ) | ( n21183 & n21205 ) | ( n21199 & n21205 ) ;
  assign n21207 = ( x174 & x625 ) | ( x174 & x1153 ) | ( x625 & x1153 ) ;
  assign n21208 = x625 & x1153 ;
  assign n21209 = ( ~n14834 & n21207 ) | ( ~n14834 & n21208 ) | ( n21207 & n21208 ) ;
  assign n21210 = x174 | n15070 ;
  assign n21211 = n17892 & n21210 ;
  assign n21212 = x696 & ~n1924 ;
  assign n21213 = ~n2031 & n21212 ;
  assign n21214 = ~n21211 & n21213 ;
  assign n21215 = ( x38 & x174 ) | ( x38 & n16319 ) | ( x174 & n16319 ) ;
  assign n21216 = ( ~x38 & x174 ) | ( ~x38 & n16322 ) | ( x174 & n16322 ) ;
  assign n21217 = x38 & ~x174 ;
  assign n21218 = ( n16321 & n21216 ) | ( n16321 & ~n21217 ) | ( n21216 & ~n21217 ) ;
  assign n21219 = n21214 & ~n21218 ;
  assign n21220 = ( n21214 & n21215 ) | ( n21214 & n21219 ) | ( n21215 & n21219 ) ;
  assign n21221 = x174 | n21213 ;
  assign n21222 = ( ~n14834 & n21213 ) | ( ~n14834 & n21221 ) | ( n21213 & n21221 ) ;
  assign n21223 = ( ~x625 & x1153 ) | ( ~x625 & n21222 ) | ( x1153 & n21222 ) ;
  assign n21224 = ( n17208 & ~n21220 ) | ( n17208 & n21223 ) | ( ~n21220 & n21223 ) ;
  assign n21225 = n21209 & n21224 ;
  assign n21226 = ( ~x174 & x625 ) | ( ~x174 & x1153 ) | ( x625 & x1153 ) ;
  assign n21227 = ( n14834 & n17301 ) | ( n14834 & n21226 ) | ( n17301 & n21226 ) ;
  assign n21228 = ( x625 & ~x1153 ) | ( x625 & n21222 ) | ( ~x1153 & n21222 ) ;
  assign n21229 = x625 & ~x1153 ;
  assign n21230 = ( ~n21220 & n21228 ) | ( ~n21220 & n21229 ) | ( n21228 & n21229 ) ;
  assign n21231 = ~n21227 & n21230 ;
  assign n21232 = n21225 | n21231 ;
  assign n21233 = ~x778 & n21222 ;
  assign n21234 = ~n21220 & n21233 ;
  assign n21235 = x778 | n21234 ;
  assign n21236 = n15400 | n21235 ;
  assign n21237 = n15400 | n21234 ;
  assign n21238 = ( n21232 & n21236 ) | ( n21232 & n21237 ) | ( n21236 & n21237 ) ;
  assign n21239 = ~x174 & n15414 ;
  assign n21240 = ( n14834 & n15414 ) | ( n14834 & n21239 ) | ( n15414 & n21239 ) ;
  assign n21241 = ~x174 & n15400 ;
  assign n21242 = ( n14834 & n15400 ) | ( n14834 & n21241 ) | ( n15400 & n21241 ) ;
  assign n21243 = n15407 | n21242 ;
  assign n21244 = x174 & n15407 ;
  assign n21245 = ~n14834 & n21244 ;
  assign n21246 = n21243 & ~n21245 ;
  assign n21247 = ~n15414 & n21246 ;
  assign n21248 = n21240 | n21247 ;
  assign n21249 = n15421 | n21248 ;
  assign n21250 = n15414 | n21245 ;
  assign n21251 = ~n21240 & n21250 ;
  assign n21252 = ~n15421 & n21251 ;
  assign n21253 = ( n21238 & ~n21249 ) | ( n21238 & n21252 ) | ( ~n21249 & n21252 ) ;
  assign n21254 = ( x174 & x628 ) | ( x174 & x1156 ) | ( x628 & x1156 ) ;
  assign n21255 = ( ~n14834 & n17218 ) | ( ~n14834 & n21254 ) | ( n17218 & n21254 ) ;
  assign n21256 = x174 & n15421 ;
  assign n21257 = ~n14834 & n21256 ;
  assign n21258 = ( ~x628 & x1156 ) | ( ~x628 & n21257 ) | ( x1156 & n21257 ) ;
  assign n21259 = n21255 & n21258 ;
  assign n21260 = ~n16052 & n21255 ;
  assign n21261 = ( n21253 & n21259 ) | ( n21253 & n21260 ) | ( n21259 & n21260 ) ;
  assign n21262 = ( ~x174 & x628 ) | ( ~x174 & x1156 ) | ( x628 & x1156 ) ;
  assign n21263 = ( n14834 & n17217 ) | ( n14834 & n21262 ) | ( n17217 & n21262 ) ;
  assign n21264 = ( x628 & ~x1156 ) | ( x628 & n21257 ) | ( ~x1156 & n21257 ) ;
  assign n21265 = ~n21263 & n21264 ;
  assign n21266 = n16051 | n21263 ;
  assign n21267 = ( n21253 & n21265 ) | ( n21253 & ~n21266 ) | ( n21265 & ~n21266 ) ;
  assign n21268 = n21261 | n21267 ;
  assign n21269 = ~x792 & n21257 ;
  assign n21270 = ( ~x792 & n21253 ) | ( ~x792 & n21269 ) | ( n21253 & n21269 ) ;
  assign n21271 = x792 | n21270 ;
  assign n21272 = ( n21268 & n21270 ) | ( n21268 & n21271 ) | ( n21270 & n21271 ) ;
  assign n21273 = ( x174 & x647 ) | ( x174 & x1157 ) | ( x647 & x1157 ) ;
  assign n21274 = x647 & x1157 ;
  assign n21275 = ( ~n14834 & n21273 ) | ( ~n14834 & n21274 ) | ( n21273 & n21274 ) ;
  assign n21276 = ~x647 & n21275 ;
  assign n21277 = x630 | n21276 ;
  assign n21278 = x1157 & n21275 ;
  assign n21279 = x630 | n21278 ;
  assign n21280 = ( n21272 & n21277 ) | ( n21272 & n21279 ) | ( n21277 & n21279 ) ;
  assign n21281 = x629 | n21259 ;
  assign n21282 = x629 | n21260 ;
  assign n21283 = ( n21253 & n21281 ) | ( n21253 & n21282 ) | ( n21281 & n21282 ) ;
  assign n21284 = ( x626 & x641 ) | ( x626 & ~n21180 ) | ( x641 & ~n21180 ) ;
  assign n21285 = ( x626 & x641 ) | ( x626 & ~n21179 ) | ( x641 & ~n21179 ) ;
  assign n21286 = ( ~n21176 & n21284 ) | ( ~n21176 & n21285 ) | ( n21284 & n21285 ) ;
  assign n21287 = ( x174 & x626 ) | ( x174 & ~x641 ) | ( x626 & ~x641 ) ;
  assign n21288 = ( ~n14834 & n16113 ) | ( ~n14834 & n21287 ) | ( n16113 & n21287 ) ;
  assign n21289 = ~x1158 & n21288 ;
  assign n21290 = ( x1158 & n21286 ) | ( x1158 & ~n21289 ) | ( n21286 & ~n21289 ) ;
  assign n21291 = x648 | n21101 ;
  assign n21292 = ( x648 & n21167 ) | ( x648 & n21291 ) | ( n21167 & n21291 ) ;
  assign n21293 = x627 | n21103 ;
  assign n21294 = ( x627 & n21152 ) | ( x627 & n21293 ) | ( n21152 & n21293 ) ;
  assign n21295 = x660 | n21105 ;
  assign n21296 = ( x660 & n21137 ) | ( x660 & n21295 ) | ( n21137 & n21295 ) ;
  assign n21297 = x608 | n21209 ;
  assign n21298 = ( x608 & n21224 ) | ( x608 & n21297 ) | ( n21224 & n21297 ) ;
  assign n21299 = ( x174 & ~x759 ) | ( x174 & n15887 ) | ( ~x759 & n15887 ) ;
  assign n21300 = ( x174 & x759 ) | ( x174 & n15891 ) | ( x759 & n15891 ) ;
  assign n21301 = n21299 & ~n21300 ;
  assign n21302 = ( x174 & ~x759 ) | ( x174 & n15894 ) | ( ~x759 & n15894 ) ;
  assign n21303 = ( x174 & x759 ) | ( x174 & n15369 ) | ( x759 & n15369 ) ;
  assign n21304 = x174 | x759 ;
  assign n21305 = ( n15896 & n21303 ) | ( n15896 & n21304 ) | ( n21303 & n21304 ) ;
  assign n21306 = ~n21302 & n21305 ;
  assign n21307 = n21301 | n21306 ;
  assign n21308 = ( ~x38 & n9138 ) | ( ~x38 & n21307 ) | ( n9138 & n21307 ) ;
  assign n21309 = x696 & ~n1919 ;
  assign n21310 = ( x696 & ~n15913 ) | ( x696 & n21309 ) | ( ~n15913 & n21309 ) ;
  assign n21311 = ~n21119 & n21310 ;
  assign n21312 = ( x174 & ~x759 ) | ( x174 & n15797 ) | ( ~x759 & n15797 ) ;
  assign n21313 = x759 & ~n21312 ;
  assign n21314 = x174 & ~n21312 ;
  assign n21315 = ( n15872 & n21313 ) | ( n15872 & n21314 ) | ( n21313 & n21314 ) ;
  assign n21316 = x39 & ~n21315 ;
  assign n21317 = ( x174 & x759 ) | ( x174 & n15699 ) | ( x759 & n15699 ) ;
  assign n21318 = ( ~x174 & x759 ) | ( ~x174 & n15582 ) | ( x759 & n15582 ) ;
  assign n21319 = x174 & ~x759 ;
  assign n21320 = ( n15565 & ~n21318 ) | ( n15565 & n21319 ) | ( ~n21318 & n21319 ) ;
  assign n21321 = ~n21317 & n21320 ;
  assign n21322 = n21316 & ~n21321 ;
  assign n21323 = n21311 & n21322 ;
  assign n21324 = ( ~n21308 & n21311 ) | ( ~n21308 & n21323 ) | ( n21311 & n21323 ) ;
  assign n21325 = x696 | n21124 ;
  assign n21326 = ~x696 & n21126 ;
  assign n21327 = ( n21113 & n21325 ) | ( n21113 & ~n21326 ) | ( n21325 & ~n21326 ) ;
  assign n21328 = ~n2032 & n21327 ;
  assign n21329 = ~n21324 & n21328 ;
  assign n21330 = ( x625 & x1153 ) | ( x625 & ~n21132 ) | ( x1153 & ~n21132 ) ;
  assign n21331 = ( ~n21128 & n21208 ) | ( ~n21128 & n21330 ) | ( n21208 & n21330 ) ;
  assign n21332 = ( x625 & ~x1153 ) | ( x625 & n21132 ) | ( ~x1153 & n21132 ) ;
  assign n21333 = ~n21331 & n21332 ;
  assign n21334 = n17208 | n21331 ;
  assign n21335 = ( n21329 & n21333 ) | ( n21329 & ~n21334 ) | ( n21333 & ~n21334 ) ;
  assign n21336 = n21298 | n21335 ;
  assign n21337 = x608 & n21227 ;
  assign n21338 = ( x608 & ~n21230 ) | ( x608 & n21337 ) | ( ~n21230 & n21337 ) ;
  assign n21339 = ( x625 & x1153 ) | ( x625 & n21132 ) | ( x1153 & n21132 ) ;
  assign n21340 = ( n17301 & n21128 ) | ( n17301 & n21339 ) | ( n21128 & n21339 ) ;
  assign n21341 = ( ~x625 & x1153 ) | ( ~x625 & n21132 ) | ( x1153 & n21132 ) ;
  assign n21342 = n21340 & n21341 ;
  assign n21343 = ~n21229 & n21340 ;
  assign n21344 = ( n21329 & n21342 ) | ( n21329 & n21343 ) | ( n21342 & n21343 ) ;
  assign n21345 = n21338 & ~n21344 ;
  assign n21346 = n21336 & ~n21345 ;
  assign n21347 = x778 | n21132 ;
  assign n21348 = n21329 | n21347 ;
  assign n21349 = ~x778 & n21348 ;
  assign n21350 = ( x609 & ~x1155 ) | ( x609 & n21349 ) | ( ~x1155 & n21349 ) ;
  assign n21351 = ( x609 & ~x1155 ) | ( x609 & n21348 ) | ( ~x1155 & n21348 ) ;
  assign n21352 = ( n21346 & n21350 ) | ( n21346 & n21351 ) | ( n21350 & n21351 ) ;
  assign n21353 = ( x609 & x1155 ) | ( x609 & ~n21235 ) | ( x1155 & ~n21235 ) ;
  assign n21354 = ( x609 & x1155 ) | ( x609 & ~n21234 ) | ( x1155 & ~n21234 ) ;
  assign n21355 = ( ~n21232 & n21353 ) | ( ~n21232 & n21354 ) | ( n21353 & n21354 ) ;
  assign n21356 = ~n21296 & n21355 ;
  assign n21357 = ( n21296 & n21352 ) | ( n21296 & ~n21356 ) | ( n21352 & ~n21356 ) ;
  assign n21358 = x660 & n21140 ;
  assign n21359 = ( x660 & ~n21143 ) | ( x660 & n21358 ) | ( ~n21143 & n21358 ) ;
  assign n21360 = ( ~x609 & x1155 ) | ( ~x609 & n21349 ) | ( x1155 & n21349 ) ;
  assign n21361 = ( ~x609 & x1155 ) | ( ~x609 & n21348 ) | ( x1155 & n21348 ) ;
  assign n21362 = ( n21346 & n21360 ) | ( n21346 & n21361 ) | ( n21360 & n21361 ) ;
  assign n21363 = ( x609 & x1155 ) | ( x609 & n21235 ) | ( x1155 & n21235 ) ;
  assign n21364 = ( x609 & x1155 ) | ( x609 & n21234 ) | ( x1155 & n21234 ) ;
  assign n21365 = ( n21232 & n21363 ) | ( n21232 & n21364 ) | ( n21363 & n21364 ) ;
  assign n21366 = n21359 & ~n21365 ;
  assign n21367 = ( n21359 & ~n21362 ) | ( n21359 & n21366 ) | ( ~n21362 & n21366 ) ;
  assign n21368 = n21357 & ~n21367 ;
  assign n21369 = x785 | n21349 ;
  assign n21370 = x785 | n21348 ;
  assign n21371 = ( n21346 & n21369 ) | ( n21346 & n21370 ) | ( n21369 & n21370 ) ;
  assign n21372 = ~x785 & n21371 ;
  assign n21373 = ( x618 & ~x1154 ) | ( x618 & n21372 ) | ( ~x1154 & n21372 ) ;
  assign n21374 = ( x618 & ~x1154 ) | ( x618 & n21371 ) | ( ~x1154 & n21371 ) ;
  assign n21375 = ( n21368 & n21373 ) | ( n21368 & n21374 ) | ( n21373 & n21374 ) ;
  assign n21376 = ( x618 & x1154 ) | ( x618 & n21242 ) | ( x1154 & n21242 ) ;
  assign n21377 = ( n18247 & ~n21238 ) | ( n18247 & n21376 ) | ( ~n21238 & n21376 ) ;
  assign n21378 = ~n21294 & n21377 ;
  assign n21379 = ( n21294 & n21375 ) | ( n21294 & ~n21378 ) | ( n21375 & ~n21378 ) ;
  assign n21380 = x627 & n21155 ;
  assign n21381 = ( x627 & ~n21158 ) | ( x627 & n21380 ) | ( ~n21158 & n21380 ) ;
  assign n21382 = ( ~x618 & x1154 ) | ( ~x618 & n21372 ) | ( x1154 & n21372 ) ;
  assign n21383 = ( ~x618 & x1154 ) | ( ~x618 & n21371 ) | ( x1154 & n21371 ) ;
  assign n21384 = ( n21368 & n21382 ) | ( n21368 & n21383 ) | ( n21382 & n21383 ) ;
  assign n21385 = ( x618 & x1154 ) | ( x618 & ~n21242 ) | ( x1154 & ~n21242 ) ;
  assign n21386 = ( n18246 & n21238 ) | ( n18246 & n21385 ) | ( n21238 & n21385 ) ;
  assign n21387 = n21381 & ~n21386 ;
  assign n21388 = ( n21381 & ~n21384 ) | ( n21381 & n21387 ) | ( ~n21384 & n21387 ) ;
  assign n21389 = n21379 & ~n21388 ;
  assign n21390 = x781 | n21372 ;
  assign n21391 = x781 | n21371 ;
  assign n21392 = ( n21368 & n21390 ) | ( n21368 & n21391 ) | ( n21390 & n21391 ) ;
  assign n21393 = ~x781 & n21392 ;
  assign n21394 = ( x619 & ~x1159 ) | ( x619 & n21393 ) | ( ~x1159 & n21393 ) ;
  assign n21395 = ( x619 & ~x1159 ) | ( x619 & n21392 ) | ( ~x1159 & n21392 ) ;
  assign n21396 = ( n21389 & n21394 ) | ( n21389 & n21395 ) | ( n21394 & n21395 ) ;
  assign n21397 = ( x619 & x1159 ) | ( x619 & n21246 ) | ( x1159 & n21246 ) ;
  assign n21398 = ( x619 & x1159 ) | ( x619 & ~n21245 ) | ( x1159 & ~n21245 ) ;
  assign n21399 = ( ~n21238 & n21397 ) | ( ~n21238 & n21398 ) | ( n21397 & n21398 ) ;
  assign n21400 = ~n21292 & n21399 ;
  assign n21401 = ( n21292 & n21396 ) | ( n21292 & ~n21400 ) | ( n21396 & ~n21400 ) ;
  assign n21402 = x648 & n21171 ;
  assign n21403 = ( x648 & ~n21174 ) | ( x648 & n21402 ) | ( ~n21174 & n21402 ) ;
  assign n21404 = ( ~x619 & x1159 ) | ( ~x619 & n21393 ) | ( x1159 & n21393 ) ;
  assign n21405 = ( ~x619 & x1159 ) | ( ~x619 & n21392 ) | ( x1159 & n21392 ) ;
  assign n21406 = ( n21389 & n21404 ) | ( n21389 & n21405 ) | ( n21404 & n21405 ) ;
  assign n21407 = ( x619 & x1159 ) | ( x619 & ~n21246 ) | ( x1159 & ~n21246 ) ;
  assign n21408 = ( x619 & x1159 ) | ( x619 & n21245 ) | ( x1159 & n21245 ) ;
  assign n21409 = ( n21238 & n21407 ) | ( n21238 & n21408 ) | ( n21407 & n21408 ) ;
  assign n21410 = n21403 & ~n21409 ;
  assign n21411 = ( n21403 & ~n21406 ) | ( n21403 & n21410 ) | ( ~n21406 & n21410 ) ;
  assign n21412 = n21401 & ~n21411 ;
  assign n21413 = x789 | n21393 ;
  assign n21414 = x789 | n21392 ;
  assign n21415 = ( n21389 & n21413 ) | ( n21389 & n21414 ) | ( n21413 & n21414 ) ;
  assign n21416 = ~x789 & n21415 ;
  assign n21417 = ( ~x626 & x641 ) | ( ~x626 & n21416 ) | ( x641 & n21416 ) ;
  assign n21418 = ( ~x626 & x641 ) | ( ~x626 & n21415 ) | ( x641 & n21415 ) ;
  assign n21419 = ( n21412 & n21417 ) | ( n21412 & n21418 ) | ( n21417 & n21418 ) ;
  assign n21420 = ( x626 & x641 ) | ( x626 & ~n21248 ) | ( x641 & ~n21248 ) ;
  assign n21421 = ( x626 & x641 ) | ( x626 & n21251 ) | ( x641 & n21251 ) ;
  assign n21422 = ( n21238 & n21420 ) | ( n21238 & n21421 ) | ( n21420 & n21421 ) ;
  assign n21423 = ~n21290 & n21422 ;
  assign n21424 = ( ~n21290 & n21419 ) | ( ~n21290 & n21423 ) | ( n21419 & n21423 ) ;
  assign n21425 = ( x626 & x641 ) | ( x626 & n21180 ) | ( x641 & n21180 ) ;
  assign n21426 = ( x626 & x641 ) | ( x626 & n21179 ) | ( x641 & n21179 ) ;
  assign n21427 = ( n21176 & n21425 ) | ( n21176 & n21426 ) | ( n21425 & n21426 ) ;
  assign n21428 = ( x174 & ~x626 ) | ( x174 & x641 ) | ( ~x626 & x641 ) ;
  assign n21429 = ( ~n14834 & n16112 ) | ( ~n14834 & n21428 ) | ( n16112 & n21428 ) ;
  assign n21430 = x1158 & n21429 ;
  assign n21431 = ( x1158 & n21427 ) | ( x1158 & n21430 ) | ( n21427 & n21430 ) ;
  assign n21432 = ( x626 & ~x641 ) | ( x626 & n21416 ) | ( ~x641 & n21416 ) ;
  assign n21433 = ( x626 & ~x641 ) | ( x626 & n21415 ) | ( ~x641 & n21415 ) ;
  assign n21434 = ( n21412 & n21432 ) | ( n21412 & n21433 ) | ( n21432 & n21433 ) ;
  assign n21435 = ( x626 & x641 ) | ( x626 & n21248 ) | ( x641 & n21248 ) ;
  assign n21436 = ( x626 & x641 ) | ( x626 & ~n21251 ) | ( x641 & ~n21251 ) ;
  assign n21437 = ( ~n21238 & n21435 ) | ( ~n21238 & n21436 ) | ( n21435 & n21436 ) ;
  assign n21438 = n21431 & ~n21437 ;
  assign n21439 = ( n21431 & n21434 ) | ( n21431 & n21438 ) | ( n21434 & n21438 ) ;
  assign n21440 = n21424 | n21439 ;
  assign n21441 = ~x788 & n21416 ;
  assign n21442 = ~x788 & n21415 ;
  assign n21443 = ( n21412 & n21441 ) | ( n21412 & n21442 ) | ( n21441 & n21442 ) ;
  assign n21444 = x788 | n21443 ;
  assign n21445 = ( x628 & ~x1156 ) | ( x628 & n21444 ) | ( ~x1156 & n21444 ) ;
  assign n21446 = ( x628 & ~x1156 ) | ( x628 & n21443 ) | ( ~x1156 & n21443 ) ;
  assign n21447 = ( n21440 & n21445 ) | ( n21440 & n21446 ) | ( n21445 & n21446 ) ;
  assign n21448 = ( x628 & x1156 ) | ( x628 & ~n21187 ) | ( x1156 & ~n21187 ) ;
  assign n21449 = ( n17218 & ~n21183 ) | ( n17218 & n21448 ) | ( ~n21183 & n21448 ) ;
  assign n21450 = ~n21283 & n21449 ;
  assign n21451 = ( n21283 & n21447 ) | ( n21283 & ~n21450 ) | ( n21447 & ~n21450 ) ;
  assign n21452 = x629 & ~n21265 ;
  assign n21453 = x629 & n21266 ;
  assign n21454 = ( ~n21253 & n21452 ) | ( ~n21253 & n21453 ) | ( n21452 & n21453 ) ;
  assign n21455 = ( ~x628 & x1156 ) | ( ~x628 & n21444 ) | ( x1156 & n21444 ) ;
  assign n21456 = ( ~x628 & x1156 ) | ( ~x628 & n21443 ) | ( x1156 & n21443 ) ;
  assign n21457 = ( n21440 & n21455 ) | ( n21440 & n21456 ) | ( n21455 & n21456 ) ;
  assign n21458 = ( x628 & x1156 ) | ( x628 & n21187 ) | ( x1156 & n21187 ) ;
  assign n21459 = ( n17217 & n21183 ) | ( n17217 & n21458 ) | ( n21183 & n21458 ) ;
  assign n21460 = n21454 & ~n21459 ;
  assign n21461 = ( n21454 & ~n21457 ) | ( n21454 & n21460 ) | ( ~n21457 & n21460 ) ;
  assign n21462 = n21451 & ~n21461 ;
  assign n21463 = x792 | n21444 ;
  assign n21464 = x792 | n21443 ;
  assign n21465 = ( n21440 & n21463 ) | ( n21440 & n21464 ) | ( n21463 & n21464 ) ;
  assign n21466 = ~x792 & n21465 ;
  assign n21467 = ( x647 & ~x1157 ) | ( x647 & n21466 ) | ( ~x1157 & n21466 ) ;
  assign n21468 = ( x647 & ~x1157 ) | ( x647 & n21465 ) | ( ~x1157 & n21465 ) ;
  assign n21469 = ( n21462 & n21467 ) | ( n21462 & n21468 ) | ( n21467 & n21468 ) ;
  assign n21470 = ( x647 & x1157 ) | ( x647 & ~n21191 ) | ( x1157 & ~n21191 ) ;
  assign n21471 = ( x647 & x1157 ) | ( x647 & n21200 ) | ( x1157 & n21200 ) ;
  assign n21472 = ( ~n21183 & n21470 ) | ( ~n21183 & n21471 ) | ( n21470 & n21471 ) ;
  assign n21473 = ~n21280 & n21472 ;
  assign n21474 = ( n21280 & n21469 ) | ( n21280 & ~n21473 ) | ( n21469 & ~n21473 ) ;
  assign n21475 = ( ~x174 & x647 ) | ( ~x174 & x1157 ) | ( x647 & x1157 ) ;
  assign n21476 = x647 | x1157 ;
  assign n21477 = ( n14834 & n21475 ) | ( n14834 & n21476 ) | ( n21475 & n21476 ) ;
  assign n21478 = x647 & ~n21477 ;
  assign n21479 = x630 & ~n21478 ;
  assign n21480 = x1157 | n21477 ;
  assign n21481 = x630 & n21480 ;
  assign n21482 = ( ~n21272 & n21479 ) | ( ~n21272 & n21481 ) | ( n21479 & n21481 ) ;
  assign n21483 = ( ~x647 & x1157 ) | ( ~x647 & n21466 ) | ( x1157 & n21466 ) ;
  assign n21484 = ( ~x647 & x1157 ) | ( ~x647 & n21465 ) | ( x1157 & n21465 ) ;
  assign n21485 = ( n21462 & n21483 ) | ( n21462 & n21484 ) | ( n21483 & n21484 ) ;
  assign n21486 = ( x647 & x1157 ) | ( x647 & n21191 ) | ( x1157 & n21191 ) ;
  assign n21487 = ( x647 & x1157 ) | ( x647 & ~n21200 ) | ( x1157 & ~n21200 ) ;
  assign n21488 = ( n21183 & n21486 ) | ( n21183 & n21487 ) | ( n21486 & n21487 ) ;
  assign n21489 = n21482 & ~n21488 ;
  assign n21490 = ( n21482 & ~n21485 ) | ( n21482 & n21489 ) | ( ~n21485 & n21489 ) ;
  assign n21491 = n21474 & ~n21490 ;
  assign n21492 = x787 | n21466 ;
  assign n21493 = x787 | n21465 ;
  assign n21494 = ( n21462 & n21492 ) | ( n21462 & n21493 ) | ( n21492 & n21493 ) ;
  assign n21495 = ~x787 & n21494 ;
  assign n21496 = ( x644 & ~x715 ) | ( x644 & n21495 ) | ( ~x715 & n21495 ) ;
  assign n21497 = ( x644 & ~x715 ) | ( x644 & n21494 ) | ( ~x715 & n21494 ) ;
  assign n21498 = ( n21491 & n21496 ) | ( n21491 & n21497 ) | ( n21496 & n21497 ) ;
  assign n21499 = ~x787 & n21272 ;
  assign n21500 = ( n21272 & n21276 ) | ( n21272 & n21278 ) | ( n21276 & n21278 ) ;
  assign n21501 = ( n21272 & n21478 ) | ( n21272 & ~n21480 ) | ( n21478 & ~n21480 ) ;
  assign n21502 = n21500 | n21501 ;
  assign n21503 = x787 | n21499 ;
  assign n21504 = ( n21499 & n21502 ) | ( n21499 & n21503 ) | ( n21502 & n21503 ) ;
  assign n21505 = ( x644 & x715 ) | ( x644 & ~n21504 ) | ( x715 & ~n21504 ) ;
  assign n21506 = ~n21206 & n21505 ;
  assign n21507 = ( n21206 & n21498 ) | ( n21206 & ~n21506 ) | ( n21498 & ~n21506 ) ;
  assign n21508 = ( ~x644 & x715 ) | ( ~x644 & n21495 ) | ( x715 & n21495 ) ;
  assign n21509 = ( ~x644 & x715 ) | ( ~x644 & n21494 ) | ( x715 & n21494 ) ;
  assign n21510 = ( n21491 & n21508 ) | ( n21491 & n21509 ) | ( n21508 & n21509 ) ;
  assign n21511 = ( x644 & x715 ) | ( x644 & n21504 ) | ( x715 & n21504 ) ;
  assign n21512 = ( x644 & x715 ) | ( x644 & ~n21193 ) | ( x715 & ~n21193 ) ;
  assign n21513 = x644 & ~x715 ;
  assign n21514 = ( x174 & x644 ) | ( x174 & ~x715 ) | ( x644 & ~x715 ) ;
  assign n21515 = ( ~n14834 & n21513 ) | ( ~n14834 & n21514 ) | ( n21513 & n21514 ) ;
  assign n21516 = ~n21512 & n21515 ;
  assign n21517 = x1160 & ~n21516 ;
  assign n21518 = ( x644 & x715 ) | ( x644 & n21202 ) | ( x715 & n21202 ) ;
  assign n21519 = n21515 & ~n21518 ;
  assign n21520 = x1160 & ~n21519 ;
  assign n21521 = ( ~n21183 & n21517 ) | ( ~n21183 & n21520 ) | ( n21517 & n21520 ) ;
  assign n21522 = ~n21511 & n21521 ;
  assign n21523 = x790 & ~n21522 ;
  assign n21524 = x790 & ~n21521 ;
  assign n21525 = ( n21510 & n21523 ) | ( n21510 & n21524 ) | ( n21523 & n21524 ) ;
  assign n21526 = n21507 & n21525 ;
  assign n21527 = ~x57 & x174 ;
  assign n21528 = ( x57 & n4832 ) | ( x57 & ~n21527 ) | ( n4832 & ~n21527 ) ;
  assign n21529 = ~x790 & n21495 ;
  assign n21530 = ~x790 & n21494 ;
  assign n21531 = ( n21491 & n21529 ) | ( n21491 & n21530 ) | ( n21529 & n21530 ) ;
  assign n21532 = n4832 | n21531 ;
  assign n21533 = ~n21528 & n21532 ;
  assign n21534 = ( n21526 & ~n21528 ) | ( n21526 & n21533 ) | ( ~n21528 & n21533 ) ;
  assign n21535 = x759 & n1290 ;
  assign n21536 = n14839 & n21535 ;
  assign n21537 = ~n18257 & n21536 ;
  assign n21538 = ~n16176 & n21537 ;
  assign n21539 = ~n18255 & n21538 ;
  assign n21540 = x174 | x715 ;
  assign n21541 = ( x715 & ~n1290 ) | ( x715 & n21540 ) | ( ~n1290 & n21540 ) ;
  assign n21542 = n18265 | n21541 ;
  assign n21543 = ( n21539 & n21541 ) | ( n21539 & n21542 ) | ( n21541 & n21542 ) ;
  assign n21544 = x1160 & n21543 ;
  assign n21545 = x174 & ~n1290 ;
  assign n21546 = n18315 | n21545 ;
  assign n21547 = ( n21537 & n21545 ) | ( n21537 & n21546 ) | ( n21545 & n21546 ) ;
  assign n21548 = ( x627 & n15404 ) | ( x627 & ~n21547 ) | ( n15404 & ~n21547 ) ;
  assign n21549 = x696 & ~n14839 ;
  assign n21550 = n15202 & n21549 ;
  assign n21551 = x625 & n21550 ;
  assign n21552 = x1153 & ~n21545 ;
  assign n21553 = ~n21536 & n21552 ;
  assign n21554 = ~n21551 & n21553 ;
  assign n21555 = x696 & n1290 ;
  assign n21556 = n15171 & n21555 ;
  assign n21557 = n21545 | n21556 ;
  assign n21558 = x625 & n21556 ;
  assign n21559 = n21557 & ~n21558 ;
  assign n21560 = ( x608 & n18335 ) | ( x608 & n21559 ) | ( n18335 & n21559 ) ;
  assign n21561 = ~n21554 & n21560 ;
  assign n21562 = n21536 | n21545 ;
  assign n21563 = n21550 | n21562 ;
  assign n21564 = ~n21551 & n21563 ;
  assign n21565 = ~x174 & x1153 ;
  assign n21566 = ( x1153 & n1290 ) | ( x1153 & n21565 ) | ( n1290 & n21565 ) ;
  assign n21567 = ~x625 & n21566 ;
  assign n21568 = ( ~n21556 & n21566 ) | ( ~n21556 & n21567 ) | ( n21566 & n21567 ) ;
  assign n21569 = x608 | n21568 ;
  assign n21570 = x1153 & ~n21569 ;
  assign n21571 = ( n21564 & ~n21569 ) | ( n21564 & n21570 ) | ( ~n21569 & n21570 ) ;
  assign n21572 = n21561 | n21571 ;
  assign n21573 = ~x778 & n21563 ;
  assign n21574 = x778 | n21573 ;
  assign n21575 = ( ~x609 & x1155 ) | ( ~x609 & n21574 ) | ( x1155 & n21574 ) ;
  assign n21576 = ( ~x609 & x1155 ) | ( ~x609 & n21573 ) | ( x1155 & n21573 ) ;
  assign n21577 = ( n21572 & n21575 ) | ( n21572 & n21576 ) | ( n21575 & n21576 ) ;
  assign n21578 = n15088 & n21536 ;
  assign n21579 = ( x660 & n15397 ) | ( x660 & ~n21545 ) | ( n15397 & ~n21545 ) ;
  assign n21580 = x660 & n15397 ;
  assign n21581 = ( ~n21578 & n21579 ) | ( ~n21578 & n21580 ) | ( n21579 & n21580 ) ;
  assign n21582 = x1153 & ~n21568 ;
  assign n21583 = ( n21559 & ~n21568 ) | ( n21559 & n21582 ) | ( ~n21568 & n21582 ) ;
  assign n21584 = x778 | n21545 ;
  assign n21585 = n21556 | n21584 ;
  assign n21586 = ~x778 & n21585 ;
  assign n21587 = ( x609 & x1155 ) | ( x609 & n21586 ) | ( x1155 & n21586 ) ;
  assign n21588 = ( x609 & x1155 ) | ( x609 & n21585 ) | ( x1155 & n21585 ) ;
  assign n21589 = ( n21583 & n21587 ) | ( n21583 & n21588 ) | ( n21587 & n21588 ) ;
  assign n21590 = ~n21581 & n21589 ;
  assign n21591 = ( n21577 & ~n21581 ) | ( n21577 & n21590 ) | ( ~n21581 & n21590 ) ;
  assign n21592 = ( x609 & ~x1155 ) | ( x609 & n21574 ) | ( ~x1155 & n21574 ) ;
  assign n21593 = ( x609 & ~x1155 ) | ( x609 & n21573 ) | ( ~x1155 & n21573 ) ;
  assign n21594 = ( n21572 & n21592 ) | ( n21572 & n21593 ) | ( n21592 & n21593 ) ;
  assign n21595 = ~n15094 & n21536 ;
  assign n21596 = ( x660 & n15398 ) | ( x660 & n21545 ) | ( n15398 & n21545 ) ;
  assign n21597 = x660 | n15398 ;
  assign n21598 = ( n21595 & n21596 ) | ( n21595 & n21597 ) | ( n21596 & n21597 ) ;
  assign n21599 = ( x609 & x1155 ) | ( x609 & ~n21586 ) | ( x1155 & ~n21586 ) ;
  assign n21600 = ( x609 & x1155 ) | ( x609 & ~n21585 ) | ( x1155 & ~n21585 ) ;
  assign n21601 = ( ~n21583 & n21599 ) | ( ~n21583 & n21600 ) | ( n21599 & n21600 ) ;
  assign n21602 = n21598 & ~n21601 ;
  assign n21603 = ( n21594 & n21598 ) | ( n21594 & n21602 ) | ( n21598 & n21602 ) ;
  assign n21604 = n21591 | n21603 ;
  assign n21605 = ~x785 & n21574 ;
  assign n21606 = ~x785 & n21573 ;
  assign n21607 = ( n21572 & n21605 ) | ( n21572 & n21606 ) | ( n21605 & n21606 ) ;
  assign n21608 = x785 | n21607 ;
  assign n21609 = ( ~x618 & x1154 ) | ( ~x618 & n21608 ) | ( x1154 & n21608 ) ;
  assign n21610 = ( ~x618 & x1154 ) | ( ~x618 & n21607 ) | ( x1154 & n21607 ) ;
  assign n21611 = ( n21604 & n21609 ) | ( n21604 & n21610 ) | ( n21609 & n21610 ) ;
  assign n21612 = ~n15400 & n21586 ;
  assign n21613 = ~n15400 & n21585 ;
  assign n21614 = ( n21583 & n21612 ) | ( n21583 & n21613 ) | ( n21612 & n21613 ) ;
  assign n21615 = ( x618 & x1154 ) | ( x618 & n21545 ) | ( x1154 & n21545 ) ;
  assign n21616 = ( n18247 & n21614 ) | ( n18247 & n21615 ) | ( n21614 & n21615 ) ;
  assign n21617 = ~n21548 & n21616 ;
  assign n21618 = ( ~n21548 & n21611 ) | ( ~n21548 & n21617 ) | ( n21611 & n21617 ) ;
  assign n21619 = n18366 & ~n21545 ;
  assign n21620 = ( n21537 & n21545 ) | ( n21537 & ~n21619 ) | ( n21545 & ~n21619 ) ;
  assign n21621 = ( x627 & n15405 ) | ( x627 & n21620 ) | ( n15405 & n21620 ) ;
  assign n21622 = ( x618 & ~x1154 ) | ( x618 & n21608 ) | ( ~x1154 & n21608 ) ;
  assign n21623 = ( x618 & ~x1154 ) | ( x618 & n21607 ) | ( ~x1154 & n21607 ) ;
  assign n21624 = ( n21604 & n21622 ) | ( n21604 & n21623 ) | ( n21622 & n21623 ) ;
  assign n21625 = ( x618 & x1154 ) | ( x618 & ~n21545 ) | ( x1154 & ~n21545 ) ;
  assign n21626 = ( n18246 & ~n21614 ) | ( n18246 & n21625 ) | ( ~n21614 & n21625 ) ;
  assign n21627 = n21621 & ~n21626 ;
  assign n21628 = ( n21621 & n21624 ) | ( n21621 & n21627 ) | ( n21624 & n21627 ) ;
  assign n21629 = n21618 | n21628 ;
  assign n21630 = x648 & n18250 ;
  assign n21631 = ~x648 & n18251 ;
  assign n21632 = n21630 | n21631 ;
  assign n21633 = ~n17214 & n21586 ;
  assign n21634 = ~n17214 & n21585 ;
  assign n21635 = ( n21583 & n21633 ) | ( n21583 & n21634 ) | ( n21633 & n21634 ) ;
  assign n21636 = n21632 & ~n21635 ;
  assign n21637 = ~x174 & x789 ;
  assign n21638 = ( x789 & n1290 ) | ( x789 & n21637 ) | ( n1290 & n21637 ) ;
  assign n21639 = ~n18303 & n21537 ;
  assign n21640 = n15412 & ~n21639 ;
  assign n21641 = n18384 & n21537 ;
  assign n21642 = n15411 & ~n21641 ;
  assign n21643 = n21640 | n21642 ;
  assign n21644 = n21638 & n21643 ;
  assign n21645 = ( n21636 & n21638 ) | ( n21636 & n21644 ) | ( n21638 & n21644 ) ;
  assign n21646 = n16177 | n21645 ;
  assign n21647 = ( x789 & n15414 ) | ( x789 & n21632 ) | ( n15414 & n21632 ) ;
  assign n21648 = ( ~x781 & n21608 ) | ( ~x781 & n21647 ) | ( n21608 & n21647 ) ;
  assign n21649 = ( ~x781 & n21607 ) | ( ~x781 & n21647 ) | ( n21607 & n21647 ) ;
  assign n21650 = ( n21604 & n21648 ) | ( n21604 & n21649 ) | ( n21648 & n21649 ) ;
  assign n21651 = x781 | n21650 ;
  assign n21652 = ~n21646 & n21651 ;
  assign n21653 = n21647 | n21650 ;
  assign n21654 = ~n21646 & n21653 ;
  assign n21655 = ( n21629 & n21652 ) | ( n21629 & n21654 ) | ( n21652 & n21654 ) ;
  assign n21656 = ~n17215 & n21586 ;
  assign n21657 = ~n17215 & n21585 ;
  assign n21658 = ( n21583 & n21656 ) | ( n21583 & n21657 ) | ( n21656 & n21657 ) ;
  assign n21659 = ~x630 & n17220 ;
  assign n21660 = x647 & ~n21659 ;
  assign n21661 = x630 & x647 ;
  assign n21662 = ( n21658 & n21660 ) | ( n21658 & n21661 ) | ( n21660 & n21661 ) ;
  assign n21663 = ( x1157 & n18403 ) | ( x1157 & ~n21539 ) | ( n18403 & ~n21539 ) ;
  assign n21664 = ~n21662 & n21663 ;
  assign n21665 = ( x630 & n18410 ) | ( x630 & ~n21658 ) | ( n18410 & ~n21658 ) ;
  assign n21666 = ~n18412 & n21539 ;
  assign n21667 = x1157 | n21666 ;
  assign n21668 = ( n17387 & n21665 ) | ( n17387 & ~n21667 ) | ( n21665 & ~n21667 ) ;
  assign n21669 = n21664 | n21668 ;
  assign n21670 = ~x174 & x787 ;
  assign n21671 = ( x787 & n1290 ) | ( x787 & n21670 ) | ( n1290 & n21670 ) ;
  assign n21672 = n21669 & n21671 ;
  assign n21673 = n15414 & ~n21545 ;
  assign n21674 = n16110 & ~n21673 ;
  assign n21675 = n16110 & n21545 ;
  assign n21676 = ( n21635 & n21674 ) | ( n21635 & n21675 ) | ( n21674 & n21675 ) ;
  assign n21677 = x626 & n21537 ;
  assign n21678 = ~n18255 & n21677 ;
  assign n21679 = x1158 & n21545 ;
  assign n21680 = x641 | n21679 ;
  assign n21681 = ( n15972 & n21678 ) | ( n15972 & n21680 ) | ( n21678 & n21680 ) ;
  assign n21682 = n21676 | n21681 ;
  assign n21683 = n16109 & ~n21673 ;
  assign n21684 = n16109 & n21545 ;
  assign n21685 = ( n21635 & n21683 ) | ( n21635 & n21684 ) | ( n21683 & n21684 ) ;
  assign n21686 = ~x626 & n21537 ;
  assign n21687 = ~n18255 & n21686 ;
  assign n21688 = ~x1158 & n21545 ;
  assign n21689 = x641 & ~n21688 ;
  assign n21690 = ( n15978 & ~n21687 ) | ( n15978 & n21689 ) | ( ~n21687 & n21689 ) ;
  assign n21691 = x788 & ~n21690 ;
  assign n21692 = ( x788 & n21685 ) | ( x788 & n21691 ) | ( n21685 & n21691 ) ;
  assign n21693 = n21682 & n21692 ;
  assign n21694 = n18434 | n21693 ;
  assign n21695 = x628 & n21658 ;
  assign n21696 = ( n15131 & n18421 ) | ( n15131 & ~n21539 ) | ( n18421 & ~n21539 ) ;
  assign n21697 = ~n21695 & n21696 ;
  assign n21698 = x629 & ~n21658 ;
  assign n21699 = ( x628 & n18420 ) | ( x628 & ~n21539 ) | ( n18420 & ~n21539 ) ;
  assign n21700 = ~x1156 & n21699 ;
  assign n21701 = ( ~x1156 & n21698 ) | ( ~x1156 & n21700 ) | ( n21698 & n21700 ) ;
  assign n21702 = n21697 | n21701 ;
  assign n21703 = ~x174 & x792 ;
  assign n21704 = ( x792 & n1290 ) | ( x792 & n21703 ) | ( n1290 & n21703 ) ;
  assign n21705 = n21702 & n21704 ;
  assign n21706 = n21694 & ~n21705 ;
  assign n21707 = n18431 | n21706 ;
  assign n21708 = ~n21672 & n21707 ;
  assign n21709 = ( x644 & ~x715 ) | ( x644 & n21708 ) | ( ~x715 & n21708 ) ;
  assign n21710 = ~n18431 & n21705 ;
  assign n21711 = n21672 | n21710 ;
  assign n21712 = ( ~x644 & x715 ) | ( ~x644 & n21711 ) | ( x715 & n21711 ) ;
  assign n21713 = ( n21655 & n21709 ) | ( n21655 & ~n21712 ) | ( n21709 & ~n21712 ) ;
  assign n21714 = n18441 & ~n21545 ;
  assign n21715 = ( x644 & x715 ) | ( x644 & n21714 ) | ( x715 & n21714 ) ;
  assign n21716 = ( x644 & x715 ) | ( x644 & ~n21545 ) | ( x715 & ~n21545 ) ;
  assign n21717 = ( ~n21658 & n21715 ) | ( ~n21658 & n21716 ) | ( n21715 & n21716 ) ;
  assign n21718 = n21544 & ~n21717 ;
  assign n21719 = ( n21544 & n21713 ) | ( n21544 & n21718 ) | ( n21713 & n21718 ) ;
  assign n21720 = ~x174 & x715 ;
  assign n21721 = ( x715 & n1290 ) | ( x715 & n21720 ) | ( n1290 & n21720 ) ;
  assign n21722 = n18453 & n21721 ;
  assign n21723 = ( ~n21539 & n21721 ) | ( ~n21539 & n21722 ) | ( n21721 & n21722 ) ;
  assign n21724 = x1160 | n21723 ;
  assign n21725 = ( ~x644 & x715 ) | ( ~x644 & n21708 ) | ( x715 & n21708 ) ;
  assign n21726 = ( x644 & ~x715 ) | ( x644 & n21711 ) | ( ~x715 & n21711 ) ;
  assign n21727 = ( n21655 & n21725 ) | ( n21655 & ~n21726 ) | ( n21725 & ~n21726 ) ;
  assign n21728 = ( x644 & x715 ) | ( x644 & ~n21714 ) | ( x715 & ~n21714 ) ;
  assign n21729 = ( x644 & x715 ) | ( x644 & n21545 ) | ( x715 & n21545 ) ;
  assign n21730 = ( n21658 & n21728 ) | ( n21658 & n21729 ) | ( n21728 & n21729 ) ;
  assign n21731 = ~n21724 & n21730 ;
  assign n21732 = ( ~n21724 & n21727 ) | ( ~n21724 & n21731 ) | ( n21727 & n21731 ) ;
  assign n21733 = n21719 | n21732 ;
  assign n21734 = ( x790 & x832 ) | ( x790 & ~n21708 ) | ( x832 & ~n21708 ) ;
  assign n21735 = ( x790 & x832 ) | ( x790 & n21711 ) | ( x832 & n21711 ) ;
  assign n21736 = ( ~n21655 & n21734 ) | ( ~n21655 & n21735 ) | ( n21734 & n21735 ) ;
  assign n21737 = x832 & n21736 ;
  assign n21738 = ~x790 & n21736 ;
  assign n21739 = ( ~n21733 & n21737 ) | ( ~n21733 & n21738 ) | ( n21737 & n21738 ) ;
  assign n21740 = x57 & x174 ;
  assign n21741 = x832 | n21740 ;
  assign n21742 = ~n21739 & n21741 ;
  assign n21743 = ( n21534 & ~n21739 ) | ( n21534 & n21742 ) | ( ~n21739 & n21742 ) ;
  assign n21744 = x175 | n1290 ;
  assign n21745 = x766 & n14840 ;
  assign n21746 = n21744 & ~n21745 ;
  assign n21747 = n16060 | n21746 ;
  assign n21748 = ~x785 & n21747 ;
  assign n21749 = ~n15094 & n21745 ;
  assign n21750 = n21747 | n21749 ;
  assign n21751 = x1155 & n21750 ;
  assign n21752 = ~x1155 & n21744 ;
  assign n21753 = ~n21749 & n21752 ;
  assign n21754 = n21751 | n21753 ;
  assign n21755 = x785 & n21754 ;
  assign n21756 = n21748 | n21755 ;
  assign n21757 = ~x781 & n21756 ;
  assign n21758 = n16075 | n21756 ;
  assign n21759 = x1154 & n21758 ;
  assign n21760 = n16078 | n21756 ;
  assign n21761 = ~x1154 & n21760 ;
  assign n21762 = n21759 | n21761 ;
  assign n21763 = x781 & n21762 ;
  assign n21764 = n21757 | n21763 ;
  assign n21765 = ~x789 & n21764 ;
  assign n21766 = n20948 | n21764 ;
  assign n21767 = x1159 & n21766 ;
  assign n21768 = n20951 | n21764 ;
  assign n21769 = ~x1159 & n21768 ;
  assign n21770 = n21767 | n21769 ;
  assign n21771 = x789 & n21770 ;
  assign n21772 = n21765 | n21771 ;
  assign n21773 = n16176 | n21772 ;
  assign n21774 = n16176 & ~n21744 ;
  assign n21775 = n21773 & ~n21774 ;
  assign n21776 = n15134 | n21775 ;
  assign n21777 = n15134 & ~n21744 ;
  assign n21778 = n21776 & ~n21777 ;
  assign n21779 = n18610 & n21778 ;
  assign n21780 = ( x647 & x1157 ) | ( x647 & ~n21744 ) | ( x1157 & ~n21744 ) ;
  assign n21781 = x700 & n15202 ;
  assign n21782 = n21744 & ~n21781 ;
  assign n21783 = x778 | n21782 ;
  assign n21784 = ~x625 & n21781 ;
  assign n21785 = n21782 | n21784 ;
  assign n21786 = x1153 & n21785 ;
  assign n21787 = ~x1153 & n21744 ;
  assign n21788 = ~n21784 & n21787 ;
  assign n21789 = x778 & ~n21788 ;
  assign n21790 = ~n21786 & n21789 ;
  assign n21791 = n21783 & ~n21790 ;
  assign n21792 = n16043 | n21791 ;
  assign n21793 = n16045 | n21792 ;
  assign n21794 = n16047 | n21793 ;
  assign n21795 = n16049 | n21794 ;
  assign n21796 = n16055 | n21795 ;
  assign n21797 = ( x647 & ~x1157 ) | ( x647 & n21796 ) | ( ~x1157 & n21796 ) ;
  assign n21798 = ~n21780 & n21797 ;
  assign n21799 = x630 & n21798 ;
  assign n21800 = x647 & n21796 ;
  assign n21801 = ~x647 & n21744 ;
  assign n21802 = n21800 | n21801 ;
  assign n21803 = n15138 & n21802 ;
  assign n21804 = n21799 | n21803 ;
  assign n21805 = n21779 | n21804 ;
  assign n21806 = x787 & n21805 ;
  assign n21807 = n16115 & ~n21794 ;
  assign n21808 = ( x626 & ~n15419 ) | ( x626 & n21744 ) | ( ~n15419 & n21744 ) ;
  assign n21809 = ( x626 & n15419 ) | ( x626 & ~n21772 ) | ( n15419 & ~n21772 ) ;
  assign n21810 = ~n21808 & n21809 ;
  assign n21811 = n21807 | n21810 ;
  assign n21812 = ( x626 & n15418 ) | ( x626 & ~n21744 ) | ( n15418 & ~n21744 ) ;
  assign n21813 = ( x626 & ~n15418 ) | ( x626 & n21772 ) | ( ~n15418 & n21772 ) ;
  assign n21814 = n21812 & ~n21813 ;
  assign n21815 = n21811 | n21814 ;
  assign n21816 = x788 & n21815 ;
  assign n21817 = x648 & ~n21769 ;
  assign n21818 = ( x619 & x1159 ) | ( x619 & n21793 ) | ( x1159 & n21793 ) ;
  assign n21819 = x627 | n21759 ;
  assign n21820 = ( x618 & x1154 ) | ( x618 & ~n21792 ) | ( x1154 & ~n21792 ) ;
  assign n21821 = x660 | n21751 ;
  assign n21822 = ( x609 & x1155 ) | ( x609 & ~n21791 ) | ( x1155 & ~n21791 ) ;
  assign n21823 = n14839 | n21782 ;
  assign n21824 = x625 & ~n21823 ;
  assign n21825 = n21746 & n21823 ;
  assign n21826 = n21824 | n21825 ;
  assign n21827 = n21787 & n21826 ;
  assign n21828 = x608 | n21786 ;
  assign n21829 = n21827 | n21828 ;
  assign n21830 = x1153 & n21746 ;
  assign n21831 = ~n21824 & n21830 ;
  assign n21832 = x608 & ~n21788 ;
  assign n21833 = ~n21831 & n21832 ;
  assign n21834 = n21829 & ~n21833 ;
  assign n21835 = x778 & ~n21834 ;
  assign n21836 = x778 | n21825 ;
  assign n21837 = ~n21835 & n21836 ;
  assign n21838 = ( x609 & ~x1155 ) | ( x609 & n21837 ) | ( ~x1155 & n21837 ) ;
  assign n21839 = ~n21822 & n21838 ;
  assign n21840 = n21821 | n21839 ;
  assign n21841 = x660 & ~n21753 ;
  assign n21842 = ( x609 & x1155 ) | ( x609 & n21791 ) | ( x1155 & n21791 ) ;
  assign n21843 = ( ~x609 & x1155 ) | ( ~x609 & n21837 ) | ( x1155 & n21837 ) ;
  assign n21844 = n21842 & n21843 ;
  assign n21845 = n21841 & ~n21844 ;
  assign n21846 = n21840 & ~n21845 ;
  assign n21847 = x785 & ~n21846 ;
  assign n21848 = x785 | n21837 ;
  assign n21849 = ~n21847 & n21848 ;
  assign n21850 = ( x618 & ~x1154 ) | ( x618 & n21849 ) | ( ~x1154 & n21849 ) ;
  assign n21851 = ~n21820 & n21850 ;
  assign n21852 = n21819 | n21851 ;
  assign n21853 = x627 & ~n21761 ;
  assign n21854 = ( x618 & x1154 ) | ( x618 & n21792 ) | ( x1154 & n21792 ) ;
  assign n21855 = ( ~x618 & x1154 ) | ( ~x618 & n21849 ) | ( x1154 & n21849 ) ;
  assign n21856 = n21854 & n21855 ;
  assign n21857 = n21853 & ~n21856 ;
  assign n21858 = n21852 & ~n21857 ;
  assign n21859 = x781 & ~n21858 ;
  assign n21860 = x781 | n21849 ;
  assign n21861 = ~n21859 & n21860 ;
  assign n21862 = ( ~x619 & x1159 ) | ( ~x619 & n21861 ) | ( x1159 & n21861 ) ;
  assign n21863 = n21818 & n21862 ;
  assign n21864 = n21817 & ~n21863 ;
  assign n21865 = x648 | n21767 ;
  assign n21866 = ( x619 & x1159 ) | ( x619 & ~n21793 ) | ( x1159 & ~n21793 ) ;
  assign n21867 = ( x619 & ~x1159 ) | ( x619 & n21861 ) | ( ~x1159 & n21861 ) ;
  assign n21868 = ~n21866 & n21867 ;
  assign n21869 = n21865 | n21868 ;
  assign n21870 = x789 & n21869 ;
  assign n21871 = ~n21864 & n21870 ;
  assign n21872 = ~x789 & n21861 ;
  assign n21873 = n16177 | n21872 ;
  assign n21874 = n21871 | n21873 ;
  assign n21875 = ~n21816 & n21874 ;
  assign n21876 = n18434 | n21875 ;
  assign n21877 = n16650 | n21795 ;
  assign n21878 = n16051 & ~n21775 ;
  assign n21879 = n21877 & ~n21878 ;
  assign n21880 = ( x629 & ~x792 ) | ( x629 & n21879 ) | ( ~x792 & n21879 ) ;
  assign n21881 = n16052 & ~n21775 ;
  assign n21882 = n16643 & ~n21795 ;
  assign n21883 = n21881 | n21882 ;
  assign n21884 = ( x629 & x792 ) | ( x629 & n21883 ) | ( x792 & n21883 ) ;
  assign n21885 = ~n21880 & n21884 ;
  assign n21886 = n18431 | n21885 ;
  assign n21887 = n21876 & ~n21886 ;
  assign n21888 = n21806 | n21887 ;
  assign n21889 = ( x790 & x832 ) | ( x790 & n21888 ) | ( x832 & n21888 ) ;
  assign n21890 = n15141 | n21778 ;
  assign n21891 = n15141 & ~n21744 ;
  assign n21892 = n21890 & ~n21891 ;
  assign n21893 = ( x644 & x715 ) | ( x644 & ~n21892 ) | ( x715 & ~n21892 ) ;
  assign n21894 = ( x644 & ~x715 ) | ( x644 & n21744 ) | ( ~x715 & n21744 ) ;
  assign n21895 = ~n21893 & n21894 ;
  assign n21896 = x1160 & ~n21895 ;
  assign n21897 = ~x787 & n21796 ;
  assign n21898 = x1157 & n21802 ;
  assign n21899 = n21798 | n21898 ;
  assign n21900 = x787 & n21899 ;
  assign n21901 = n21897 | n21900 ;
  assign n21902 = ( x644 & x715 ) | ( x644 & n21901 ) | ( x715 & n21901 ) ;
  assign n21903 = ( ~x644 & x715 ) | ( ~x644 & n21888 ) | ( x715 & n21888 ) ;
  assign n21904 = n21902 & n21903 ;
  assign n21905 = n21896 & ~n21904 ;
  assign n21906 = ( x644 & x715 ) | ( x644 & n21892 ) | ( x715 & n21892 ) ;
  assign n21907 = ( ~x644 & x715 ) | ( ~x644 & n21744 ) | ( x715 & n21744 ) ;
  assign n21908 = n21906 & n21907 ;
  assign n21909 = x1160 | n21908 ;
  assign n21910 = ( x644 & x715 ) | ( x644 & ~n21901 ) | ( x715 & ~n21901 ) ;
  assign n21911 = ( x644 & ~x715 ) | ( x644 & n21888 ) | ( ~x715 & n21888 ) ;
  assign n21912 = ~n21910 & n21911 ;
  assign n21913 = n21909 | n21912 ;
  assign n21914 = ~n21905 & n21913 ;
  assign n21915 = ( ~x790 & x832 ) | ( ~x790 & n21914 ) | ( x832 & n21914 ) ;
  assign n21916 = n21889 & n21915 ;
  assign n21917 = x175 | n14834 ;
  assign n21918 = n15414 & n21917 ;
  assign n21919 = x175 & n2032 ;
  assign n21920 = x175 | n15070 ;
  assign n21921 = n15375 & n21920 ;
  assign n21922 = x700 & ~n21921 ;
  assign n21923 = ( ~x38 & x175 ) | ( ~x38 & n16319 ) | ( x175 & n16319 ) ;
  assign n21924 = ( x38 & x175 ) | ( x38 & n16323 ) | ( x175 & n16323 ) ;
  assign n21925 = n21923 & ~n21924 ;
  assign n21926 = n21922 & ~n21925 ;
  assign n21927 = x175 | x700 ;
  assign n21928 = n15382 | n21927 ;
  assign n21929 = ~n2032 & n21928 ;
  assign n21930 = ~n21926 & n21929 ;
  assign n21931 = n21919 | n21930 ;
  assign n21932 = ~x778 & n21931 ;
  assign n21933 = ( x625 & x1153 ) | ( x625 & n21917 ) | ( x1153 & n21917 ) ;
  assign n21934 = ( ~x625 & x1153 ) | ( ~x625 & n21931 ) | ( x1153 & n21931 ) ;
  assign n21935 = n21933 & n21934 ;
  assign n21936 = ( x625 & x1153 ) | ( x625 & ~n21917 ) | ( x1153 & ~n21917 ) ;
  assign n21937 = ( x625 & ~x1153 ) | ( x625 & n21931 ) | ( ~x1153 & n21931 ) ;
  assign n21938 = ~n21936 & n21937 ;
  assign n21939 = n21935 | n21938 ;
  assign n21940 = x778 & n21939 ;
  assign n21941 = n21932 | n21940 ;
  assign n21942 = ~n15400 & n21941 ;
  assign n21943 = n15400 & n21917 ;
  assign n21944 = n21942 | n21943 ;
  assign n21945 = n15407 | n21944 ;
  assign n21946 = n15407 & ~n21917 ;
  assign n21947 = n21945 & ~n21946 ;
  assign n21948 = ~n15414 & n21947 ;
  assign n21949 = n21918 | n21948 ;
  assign n21950 = n15421 | n21949 ;
  assign n21951 = n15421 & ~n21917 ;
  assign n21952 = n21950 & ~n21951 ;
  assign n21953 = x792 | n21952 ;
  assign n21954 = x628 & ~n21952 ;
  assign n21955 = x628 | n21917 ;
  assign n21956 = ~n21954 & n21955 ;
  assign n21957 = ( ~x792 & x1156 ) | ( ~x792 & n21956 ) | ( x1156 & n21956 ) ;
  assign n21958 = x628 | n21952 ;
  assign n21959 = x628 & ~n21917 ;
  assign n21960 = n21958 & ~n21959 ;
  assign n21961 = ( x792 & x1156 ) | ( x792 & ~n21960 ) | ( x1156 & ~n21960 ) ;
  assign n21962 = ~n21957 & n21961 ;
  assign n21963 = n21953 & ~n21962 ;
  assign n21964 = x787 | n21963 ;
  assign n21965 = x647 & ~n21963 ;
  assign n21966 = x647 | n21917 ;
  assign n21967 = ~n21965 & n21966 ;
  assign n21968 = ( ~x787 & x1157 ) | ( ~x787 & n21967 ) | ( x1157 & n21967 ) ;
  assign n21969 = x647 | n21963 ;
  assign n21970 = x647 & ~n21917 ;
  assign n21971 = n21969 & ~n21970 ;
  assign n21972 = ( x787 & x1157 ) | ( x787 & ~n21971 ) | ( x1157 & ~n21971 ) ;
  assign n21973 = ~n21968 & n21972 ;
  assign n21974 = n21964 & ~n21973 ;
  assign n21975 = x644 | n21974 ;
  assign n21976 = x715 & n21975 ;
  assign n21977 = ~x766 & n14710 ;
  assign n21978 = x175 & ~n14907 ;
  assign n21979 = n21977 | n21978 ;
  assign n21980 = x39 & n21979 ;
  assign n21981 = ~x175 & x766 ;
  assign n21982 = n15063 & n21981 ;
  assign n21983 = x766 & n14932 ;
  assign n21984 = x175 & ~n21983 ;
  assign n21985 = n19484 | n21984 ;
  assign n21986 = n21982 | n21985 ;
  assign n21987 = n21980 | n21986 ;
  assign n21988 = ~x38 & n21987 ;
  assign n21989 = x766 & n15072 ;
  assign n21990 = x38 & n21920 ;
  assign n21991 = ~n21989 & n21990 ;
  assign n21992 = n21988 | n21991 ;
  assign n21993 = ~n2032 & n21992 ;
  assign n21994 = n21919 | n21993 ;
  assign n21995 = ~n15082 & n21994 ;
  assign n21996 = n15082 & n21917 ;
  assign n21997 = n21995 | n21996 ;
  assign n21998 = ~x785 & n21997 ;
  assign n21999 = ~n15088 & n21917 ;
  assign n22000 = x609 & n21995 ;
  assign n22001 = n21999 | n22000 ;
  assign n22002 = x1155 & n22001 ;
  assign n22003 = n15094 & n21917 ;
  assign n22004 = ~x609 & n21995 ;
  assign n22005 = n22003 | n22004 ;
  assign n22006 = ~x1155 & n22005 ;
  assign n22007 = n22002 | n22006 ;
  assign n22008 = x785 & n22007 ;
  assign n22009 = n21998 | n22008 ;
  assign n22010 = ~x781 & n22009 ;
  assign n22011 = ( x618 & x1154 ) | ( x618 & n21917 ) | ( x1154 & n21917 ) ;
  assign n22012 = ( ~x618 & x1154 ) | ( ~x618 & n22009 ) | ( x1154 & n22009 ) ;
  assign n22013 = n22011 & n22012 ;
  assign n22014 = ( x618 & x1154 ) | ( x618 & ~n21917 ) | ( x1154 & ~n21917 ) ;
  assign n22015 = ( x618 & ~x1154 ) | ( x618 & n22009 ) | ( ~x1154 & n22009 ) ;
  assign n22016 = ~n22014 & n22015 ;
  assign n22017 = n22013 | n22016 ;
  assign n22018 = x781 & n22017 ;
  assign n22019 = n22010 | n22018 ;
  assign n22020 = ~x789 & n22019 ;
  assign n22021 = ( x619 & x1159 ) | ( x619 & n21917 ) | ( x1159 & n21917 ) ;
  assign n22022 = ( ~x619 & x1159 ) | ( ~x619 & n22019 ) | ( x1159 & n22019 ) ;
  assign n22023 = n22021 & n22022 ;
  assign n22024 = ( x619 & x1159 ) | ( x619 & ~n21917 ) | ( x1159 & ~n21917 ) ;
  assign n22025 = ( x619 & ~x1159 ) | ( x619 & n22019 ) | ( ~x1159 & n22019 ) ;
  assign n22026 = ~n22024 & n22025 ;
  assign n22027 = n22023 | n22026 ;
  assign n22028 = x789 & n22027 ;
  assign n22029 = n22020 | n22028 ;
  assign n22030 = n16176 | n22029 ;
  assign n22031 = n16176 & ~n21917 ;
  assign n22032 = n22030 & ~n22031 ;
  assign n22033 = n15134 | n22032 ;
  assign n22034 = n15134 & ~n21917 ;
  assign n22035 = n22033 & ~n22034 ;
  assign n22036 = n15141 | n22035 ;
  assign n22037 = n15141 & ~n21917 ;
  assign n22038 = n22036 & ~n22037 ;
  assign n22039 = ( x644 & x715 ) | ( x644 & ~n22038 ) | ( x715 & ~n22038 ) ;
  assign n22040 = ( x644 & ~x715 ) | ( x644 & n21917 ) | ( ~x715 & n21917 ) ;
  assign n22041 = ~n22039 & n22040 ;
  assign n22042 = x1160 & ~n22041 ;
  assign n22043 = ~n21976 & n22042 ;
  assign n22044 = x644 & ~n21974 ;
  assign n22045 = x715 | n22044 ;
  assign n22046 = ( x644 & x715 ) | ( x644 & n22038 ) | ( x715 & n22038 ) ;
  assign n22047 = ( ~x644 & x715 ) | ( ~x644 & n21917 ) | ( x715 & n21917 ) ;
  assign n22048 = n22046 & n22047 ;
  assign n22049 = x1160 | n22048 ;
  assign n22050 = n22045 & ~n22049 ;
  assign n22051 = n22043 | n22050 ;
  assign n22052 = x790 & n22051 ;
  assign n22053 = n18621 & n22032 ;
  assign n22054 = n15132 & n21960 ;
  assign n22055 = n15131 & n21956 ;
  assign n22056 = n22054 | n22055 ;
  assign n22057 = n22053 | n22056 ;
  assign n22058 = x792 & n22057 ;
  assign n22059 = x648 & ~n22026 ;
  assign n22060 = ( x619 & x1159 ) | ( x619 & n21947 ) | ( x1159 & n21947 ) ;
  assign n22061 = x627 | n22013 ;
  assign n22062 = ( x618 & x1154 ) | ( x618 & ~n21944 ) | ( x1154 & ~n21944 ) ;
  assign n22063 = x660 | n22002 ;
  assign n22064 = ( x609 & x1155 ) | ( x609 & ~n21941 ) | ( x1155 & ~n21941 ) ;
  assign n22065 = x608 | n21935 ;
  assign n22066 = ( x625 & x1153 ) | ( x625 & ~n21994 ) | ( x1153 & ~n21994 ) ;
  assign n22067 = x700 | n21992 ;
  assign n22068 = ( x175 & ~x766 ) | ( x175 & n15872 ) | ( ~x766 & n15872 ) ;
  assign n22069 = ( x175 & x766 ) | ( x175 & n15797 ) | ( x766 & n15797 ) ;
  assign n22070 = ~n22068 & n22069 ;
  assign n22071 = x39 & ~n22070 ;
  assign n22072 = ( x175 & ~x766 ) | ( x175 & n15699 ) | ( ~x766 & n15699 ) ;
  assign n22073 = ( x175 & x766 ) | ( x175 & n15583 ) | ( x766 & n15583 ) ;
  assign n22074 = n22072 & ~n22073 ;
  assign n22075 = n22071 & ~n22074 ;
  assign n22076 = ( x175 & ~x766 ) | ( x175 & n15891 ) | ( ~x766 & n15891 ) ;
  assign n22077 = ( x175 & x766 ) | ( x175 & n15887 ) | ( x766 & n15887 ) ;
  assign n22078 = n22076 & ~n22077 ;
  assign n22079 = ( x175 & ~x766 ) | ( x175 & n15897 ) | ( ~x766 & n15897 ) ;
  assign n22080 = ( x175 & x766 ) | ( x175 & n15894 ) | ( x766 & n15894 ) ;
  assign n22081 = ~n22079 & n22080 ;
  assign n22082 = n22078 | n22081 ;
  assign n22083 = ( ~x38 & n9138 ) | ( ~x38 & n22082 ) | ( n9138 & n22082 ) ;
  assign n22084 = ~n22075 & n22083 ;
  assign n22085 = n15585 & n15756 ;
  assign n22086 = ~x766 & n22085 ;
  assign n22087 = n15758 | n22086 ;
  assign n22088 = ~x39 & n22087 ;
  assign n22089 = x175 | n22088 ;
  assign n22090 = n15529 | n21745 ;
  assign n22091 = x175 & n22090 ;
  assign n22092 = ~n4810 & n22091 ;
  assign n22093 = x38 & ~n22092 ;
  assign n22094 = n22089 & n22093 ;
  assign n22095 = x700 & ~n22094 ;
  assign n22096 = ~n22084 & n22095 ;
  assign n22097 = n2032 | n22096 ;
  assign n22098 = n22067 & ~n22097 ;
  assign n22099 = n21919 | n22098 ;
  assign n22100 = ( x625 & ~x1153 ) | ( x625 & n22099 ) | ( ~x1153 & n22099 ) ;
  assign n22101 = ~n22066 & n22100 ;
  assign n22102 = n22065 | n22101 ;
  assign n22103 = x608 & ~n21938 ;
  assign n22104 = ( x625 & x1153 ) | ( x625 & n21994 ) | ( x1153 & n21994 ) ;
  assign n22105 = ( ~x625 & x1153 ) | ( ~x625 & n22099 ) | ( x1153 & n22099 ) ;
  assign n22106 = n22104 & n22105 ;
  assign n22107 = n22103 & ~n22106 ;
  assign n22108 = n22102 & ~n22107 ;
  assign n22109 = x778 & ~n22108 ;
  assign n22110 = x778 | n22099 ;
  assign n22111 = ~n22109 & n22110 ;
  assign n22112 = ( x609 & ~x1155 ) | ( x609 & n22111 ) | ( ~x1155 & n22111 ) ;
  assign n22113 = ~n22064 & n22112 ;
  assign n22114 = n22063 | n22113 ;
  assign n22115 = x660 & ~n22006 ;
  assign n22116 = ( x609 & x1155 ) | ( x609 & n21941 ) | ( x1155 & n21941 ) ;
  assign n22117 = ( ~x609 & x1155 ) | ( ~x609 & n22111 ) | ( x1155 & n22111 ) ;
  assign n22118 = n22116 & n22117 ;
  assign n22119 = n22115 & ~n22118 ;
  assign n22120 = n22114 & ~n22119 ;
  assign n22121 = x785 & ~n22120 ;
  assign n22122 = x785 | n22111 ;
  assign n22123 = ~n22121 & n22122 ;
  assign n22124 = ( x618 & ~x1154 ) | ( x618 & n22123 ) | ( ~x1154 & n22123 ) ;
  assign n22125 = ~n22062 & n22124 ;
  assign n22126 = n22061 | n22125 ;
  assign n22127 = x627 & ~n22016 ;
  assign n22128 = ( x618 & x1154 ) | ( x618 & n21944 ) | ( x1154 & n21944 ) ;
  assign n22129 = ( ~x618 & x1154 ) | ( ~x618 & n22123 ) | ( x1154 & n22123 ) ;
  assign n22130 = n22128 & n22129 ;
  assign n22131 = n22127 & ~n22130 ;
  assign n22132 = n22126 & ~n22131 ;
  assign n22133 = x781 & ~n22132 ;
  assign n22134 = x781 | n22123 ;
  assign n22135 = ~n22133 & n22134 ;
  assign n22136 = ( ~x619 & x1159 ) | ( ~x619 & n22135 ) | ( x1159 & n22135 ) ;
  assign n22137 = n22060 & n22136 ;
  assign n22138 = n22059 & ~n22137 ;
  assign n22139 = x648 | n22023 ;
  assign n22140 = ( x619 & x1159 ) | ( x619 & ~n21947 ) | ( x1159 & ~n21947 ) ;
  assign n22141 = ( x619 & ~x1159 ) | ( x619 & n22135 ) | ( ~x1159 & n22135 ) ;
  assign n22142 = ~n22140 & n22141 ;
  assign n22143 = n22139 | n22142 ;
  assign n22144 = x789 & n22143 ;
  assign n22145 = ~n22138 & n22144 ;
  assign n22146 = ~x789 & n22135 ;
  assign n22147 = n16177 | n22146 ;
  assign n22148 = n22145 | n22147 ;
  assign n22149 = n16115 & ~n21949 ;
  assign n22150 = ( x626 & ~n15419 ) | ( x626 & n21917 ) | ( ~n15419 & n21917 ) ;
  assign n22151 = ( x626 & n15419 ) | ( x626 & ~n22029 ) | ( n15419 & ~n22029 ) ;
  assign n22152 = ~n22150 & n22151 ;
  assign n22153 = n22149 | n22152 ;
  assign n22154 = ( x626 & n15418 ) | ( x626 & ~n21917 ) | ( n15418 & ~n21917 ) ;
  assign n22155 = ( x626 & ~n15418 ) | ( x626 & n22029 ) | ( ~n15418 & n22029 ) ;
  assign n22156 = n22154 & ~n22155 ;
  assign n22157 = n22153 | n22156 ;
  assign n22158 = x788 & n22157 ;
  assign n22159 = n18434 | n22158 ;
  assign n22160 = n22148 & ~n22159 ;
  assign n22161 = n22058 | n22160 ;
  assign n22162 = ~n18431 & n22161 ;
  assign n22163 = n15138 & n21967 ;
  assign n22164 = n15139 & n21971 ;
  assign n22165 = n18610 & n22035 ;
  assign n22166 = n22164 | n22165 ;
  assign n22167 = n22163 | n22166 ;
  assign n22168 = x787 & n22167 ;
  assign n22169 = n22162 | n22168 ;
  assign n22170 = ( x644 & ~x790 ) | ( x644 & n22042 ) | ( ~x790 & n22042 ) ;
  assign n22171 = ( x644 & x790 ) | ( x644 & n22049 ) | ( x790 & n22049 ) ;
  assign n22172 = ~n22170 & n22171 ;
  assign n22173 = n22169 | n22172 ;
  assign n22174 = ~n22052 & n22173 ;
  assign n22175 = ( ~x832 & n6785 ) | ( ~x832 & n22174 ) | ( n6785 & n22174 ) ;
  assign n22176 = ( ~x175 & x832 ) | ( ~x175 & n6785 ) | ( x832 & n6785 ) ;
  assign n22177 = n22175 & ~n22176 ;
  assign n22178 = n21916 | n22177 ;
  assign n22179 = x176 | n1290 ;
  assign n22180 = ~x742 & n14840 ;
  assign n22181 = n22179 & ~n22180 ;
  assign n22182 = n16060 | n22181 ;
  assign n22183 = ~x785 & n22182 ;
  assign n22184 = n16065 | n22181 ;
  assign n22185 = x1155 & n22184 ;
  assign n22186 = n16068 | n22182 ;
  assign n22187 = ~x1155 & n22186 ;
  assign n22188 = n22185 | n22187 ;
  assign n22189 = x785 & n22188 ;
  assign n22190 = n22183 | n22189 ;
  assign n22191 = ~x781 & n22190 ;
  assign n22192 = n16075 | n22190 ;
  assign n22193 = x1154 & n22192 ;
  assign n22194 = n16078 | n22190 ;
  assign n22195 = ~x1154 & n22194 ;
  assign n22196 = n22193 | n22195 ;
  assign n22197 = x781 & n22196 ;
  assign n22198 = n22191 | n22197 ;
  assign n22199 = ~x789 & n22198 ;
  assign n22200 = ( x619 & x1159 ) | ( x619 & n22179 ) | ( x1159 & n22179 ) ;
  assign n22201 = ( ~x619 & x1159 ) | ( ~x619 & n22198 ) | ( x1159 & n22198 ) ;
  assign n22202 = n22200 & n22201 ;
  assign n22203 = ( x619 & x1159 ) | ( x619 & ~n22179 ) | ( x1159 & ~n22179 ) ;
  assign n22204 = ( x619 & ~x1159 ) | ( x619 & n22198 ) | ( ~x1159 & n22198 ) ;
  assign n22205 = ~n22203 & n22204 ;
  assign n22206 = n22202 | n22205 ;
  assign n22207 = x789 & n22206 ;
  assign n22208 = n22199 | n22207 ;
  assign n22209 = n16176 | n22208 ;
  assign n22210 = n16176 & ~n22179 ;
  assign n22211 = n22209 & ~n22210 ;
  assign n22212 = n15134 | n22211 ;
  assign n22213 = n15134 & ~n22179 ;
  assign n22214 = n22212 & ~n22213 ;
  assign n22215 = n18610 & n22214 ;
  assign n22216 = ( x647 & x1157 ) | ( x647 & ~n22179 ) | ( x1157 & ~n22179 ) ;
  assign n22217 = ~x704 & n15202 ;
  assign n22218 = n22179 & ~n22217 ;
  assign n22219 = ~x778 & n22218 ;
  assign n22220 = ~x625 & n22217 ;
  assign n22221 = n22218 | n22220 ;
  assign n22222 = x1153 & n22221 ;
  assign n22223 = ~x1153 & n22179 ;
  assign n22224 = ~n22220 & n22223 ;
  assign n22225 = n22222 | n22224 ;
  assign n22226 = x778 & n22225 ;
  assign n22227 = n22219 | n22226 ;
  assign n22228 = n16043 | n22227 ;
  assign n22229 = n16045 | n22228 ;
  assign n22230 = n16047 | n22229 ;
  assign n22231 = n16049 | n22230 ;
  assign n22232 = n16055 | n22231 ;
  assign n22233 = ( x647 & ~x1157 ) | ( x647 & n22232 ) | ( ~x1157 & n22232 ) ;
  assign n22234 = ~n22216 & n22233 ;
  assign n22235 = x630 & n22234 ;
  assign n22236 = x647 & n22232 ;
  assign n22237 = ~x647 & n22179 ;
  assign n22238 = n22236 | n22237 ;
  assign n22239 = n15138 & n22238 ;
  assign n22240 = n22235 | n22239 ;
  assign n22241 = n22215 | n22240 ;
  assign n22242 = x787 & n22241 ;
  assign n22243 = n16115 & ~n22230 ;
  assign n22244 = ( x626 & ~n15419 ) | ( x626 & n22179 ) | ( ~n15419 & n22179 ) ;
  assign n22245 = ( x626 & n15419 ) | ( x626 & ~n22208 ) | ( n15419 & ~n22208 ) ;
  assign n22246 = ~n22244 & n22245 ;
  assign n22247 = n22243 | n22246 ;
  assign n22248 = ( x626 & n15418 ) | ( x626 & ~n22179 ) | ( n15418 & ~n22179 ) ;
  assign n22249 = ( x626 & ~n15418 ) | ( x626 & n22208 ) | ( ~n15418 & n22208 ) ;
  assign n22250 = n22248 & ~n22249 ;
  assign n22251 = n22247 | n22250 ;
  assign n22252 = x788 & n22251 ;
  assign n22253 = x648 & ~n22205 ;
  assign n22254 = ( x619 & x1159 ) | ( x619 & n22229 ) | ( x1159 & n22229 ) ;
  assign n22255 = x627 | n22193 ;
  assign n22256 = ( x618 & x1154 ) | ( x618 & ~n22228 ) | ( x1154 & ~n22228 ) ;
  assign n22257 = x660 | n22185 ;
  assign n22258 = ( x609 & x1155 ) | ( x609 & ~n22227 ) | ( x1155 & ~n22227 ) ;
  assign n22259 = n14839 | n22218 ;
  assign n22260 = x625 & ~n22259 ;
  assign n22261 = n22181 & n22259 ;
  assign n22262 = n22260 | n22261 ;
  assign n22263 = n22223 & n22262 ;
  assign n22264 = x608 | n22222 ;
  assign n22265 = n22263 | n22264 ;
  assign n22266 = x1153 & n22181 ;
  assign n22267 = ~n22260 & n22266 ;
  assign n22268 = x608 & ~n22224 ;
  assign n22269 = ~n22267 & n22268 ;
  assign n22270 = n22265 & ~n22269 ;
  assign n22271 = x778 & ~n22270 ;
  assign n22272 = x778 | n22261 ;
  assign n22273 = ~n22271 & n22272 ;
  assign n22274 = ( x609 & ~x1155 ) | ( x609 & n22273 ) | ( ~x1155 & n22273 ) ;
  assign n22275 = ~n22258 & n22274 ;
  assign n22276 = n22257 | n22275 ;
  assign n22277 = x660 & ~n22187 ;
  assign n22278 = ( x609 & x1155 ) | ( x609 & n22227 ) | ( x1155 & n22227 ) ;
  assign n22279 = ( ~x609 & x1155 ) | ( ~x609 & n22273 ) | ( x1155 & n22273 ) ;
  assign n22280 = n22278 & n22279 ;
  assign n22281 = n22277 & ~n22280 ;
  assign n22282 = n22276 & ~n22281 ;
  assign n22283 = x785 & ~n22282 ;
  assign n22284 = x785 | n22273 ;
  assign n22285 = ~n22283 & n22284 ;
  assign n22286 = ( x618 & ~x1154 ) | ( x618 & n22285 ) | ( ~x1154 & n22285 ) ;
  assign n22287 = ~n22256 & n22286 ;
  assign n22288 = n22255 | n22287 ;
  assign n22289 = x627 & ~n22195 ;
  assign n22290 = ( x618 & x1154 ) | ( x618 & n22228 ) | ( x1154 & n22228 ) ;
  assign n22291 = ( ~x618 & x1154 ) | ( ~x618 & n22285 ) | ( x1154 & n22285 ) ;
  assign n22292 = n22290 & n22291 ;
  assign n22293 = n22289 & ~n22292 ;
  assign n22294 = n22288 & ~n22293 ;
  assign n22295 = x781 & ~n22294 ;
  assign n22296 = x781 | n22285 ;
  assign n22297 = ~n22295 & n22296 ;
  assign n22298 = ( ~x619 & x1159 ) | ( ~x619 & n22297 ) | ( x1159 & n22297 ) ;
  assign n22299 = n22254 & n22298 ;
  assign n22300 = n22253 & ~n22299 ;
  assign n22301 = x648 | n22202 ;
  assign n22302 = ( x619 & x1159 ) | ( x619 & ~n22229 ) | ( x1159 & ~n22229 ) ;
  assign n22303 = ( x619 & ~x1159 ) | ( x619 & n22297 ) | ( ~x1159 & n22297 ) ;
  assign n22304 = ~n22302 & n22303 ;
  assign n22305 = n22301 | n22304 ;
  assign n22306 = x789 & n22305 ;
  assign n22307 = ~n22300 & n22306 ;
  assign n22308 = ~x789 & n22297 ;
  assign n22309 = n16177 | n22308 ;
  assign n22310 = n22307 | n22309 ;
  assign n22311 = ~n22252 & n22310 ;
  assign n22312 = n18434 | n22311 ;
  assign n22313 = n16650 | n22231 ;
  assign n22314 = n16051 & ~n22211 ;
  assign n22315 = n22313 & ~n22314 ;
  assign n22316 = ( x629 & ~x792 ) | ( x629 & n22315 ) | ( ~x792 & n22315 ) ;
  assign n22317 = n16052 & ~n22211 ;
  assign n22318 = n16643 & ~n22231 ;
  assign n22319 = n22317 | n22318 ;
  assign n22320 = ( x629 & x792 ) | ( x629 & n22319 ) | ( x792 & n22319 ) ;
  assign n22321 = ~n22316 & n22320 ;
  assign n22322 = n18431 | n22321 ;
  assign n22323 = n22312 & ~n22322 ;
  assign n22324 = n22242 | n22323 ;
  assign n22325 = ( x790 & x832 ) | ( x790 & n22324 ) | ( x832 & n22324 ) ;
  assign n22326 = n15141 | n22214 ;
  assign n22327 = n15141 & ~n22179 ;
  assign n22328 = n22326 & ~n22327 ;
  assign n22329 = ( x644 & x715 ) | ( x644 & ~n22328 ) | ( x715 & ~n22328 ) ;
  assign n22330 = ( x644 & ~x715 ) | ( x644 & n22179 ) | ( ~x715 & n22179 ) ;
  assign n22331 = ~n22329 & n22330 ;
  assign n22332 = x1160 & ~n22331 ;
  assign n22333 = ~x787 & n22232 ;
  assign n22334 = x1157 & n22238 ;
  assign n22335 = n22234 | n22334 ;
  assign n22336 = x787 & n22335 ;
  assign n22337 = n22333 | n22336 ;
  assign n22338 = ( x644 & x715 ) | ( x644 & n22337 ) | ( x715 & n22337 ) ;
  assign n22339 = ( ~x644 & x715 ) | ( ~x644 & n22324 ) | ( x715 & n22324 ) ;
  assign n22340 = n22338 & n22339 ;
  assign n22341 = n22332 & ~n22340 ;
  assign n22342 = ( x644 & x715 ) | ( x644 & n22328 ) | ( x715 & n22328 ) ;
  assign n22343 = ( ~x644 & x715 ) | ( ~x644 & n22179 ) | ( x715 & n22179 ) ;
  assign n22344 = n22342 & n22343 ;
  assign n22345 = x1160 | n22344 ;
  assign n22346 = ( x644 & x715 ) | ( x644 & ~n22337 ) | ( x715 & ~n22337 ) ;
  assign n22347 = ( x644 & ~x715 ) | ( x644 & n22324 ) | ( ~x715 & n22324 ) ;
  assign n22348 = ~n22346 & n22347 ;
  assign n22349 = n22345 | n22348 ;
  assign n22350 = ~n22341 & n22349 ;
  assign n22351 = ( ~x790 & x832 ) | ( ~x790 & n22350 ) | ( x832 & n22350 ) ;
  assign n22352 = n22325 & n22351 ;
  assign n22353 = x176 | n14834 ;
  assign n22354 = n15414 & n22353 ;
  assign n22355 = x38 | n16323 ;
  assign n22356 = n2032 | n15375 ;
  assign n22357 = n22355 & ~n22356 ;
  assign n22358 = x176 & ~n22357 ;
  assign n22359 = x176 | n15382 ;
  assign n22360 = ( x704 & n2032 ) | ( x704 & ~n22359 ) | ( n2032 & ~n22359 ) ;
  assign n22361 = x38 | n16319 ;
  assign n22362 = ~n17892 & n22361 ;
  assign n22363 = ~x176 & n22362 ;
  assign n22364 = ( x704 & ~n2032 ) | ( x704 & n22363 ) | ( ~n2032 & n22363 ) ;
  assign n22365 = ~n22360 & n22364 ;
  assign n22366 = n22358 | n22365 ;
  assign n22367 = ~x778 & n22366 ;
  assign n22368 = ( x625 & x1153 ) | ( x625 & n22353 ) | ( x1153 & n22353 ) ;
  assign n22369 = ( ~x625 & x1153 ) | ( ~x625 & n22366 ) | ( x1153 & n22366 ) ;
  assign n22370 = n22368 & n22369 ;
  assign n22371 = ( x625 & x1153 ) | ( x625 & ~n22353 ) | ( x1153 & ~n22353 ) ;
  assign n22372 = ( x625 & ~x1153 ) | ( x625 & n22366 ) | ( ~x1153 & n22366 ) ;
  assign n22373 = ~n22371 & n22372 ;
  assign n22374 = n22370 | n22373 ;
  assign n22375 = x778 & n22374 ;
  assign n22376 = n22367 | n22375 ;
  assign n22377 = ~n15400 & n22376 ;
  assign n22378 = n15400 & n22353 ;
  assign n22379 = n22377 | n22378 ;
  assign n22380 = n15407 | n22379 ;
  assign n22381 = n15407 & ~n22353 ;
  assign n22382 = n22380 & ~n22381 ;
  assign n22383 = ~n15414 & n22382 ;
  assign n22384 = n22354 | n22383 ;
  assign n22385 = n15421 | n22384 ;
  assign n22386 = n15421 & ~n22353 ;
  assign n22387 = n22385 & ~n22386 ;
  assign n22388 = x792 | n22387 ;
  assign n22389 = x628 & ~n22387 ;
  assign n22390 = x628 | n22353 ;
  assign n22391 = ~n22389 & n22390 ;
  assign n22392 = ( ~x792 & x1156 ) | ( ~x792 & n22391 ) | ( x1156 & n22391 ) ;
  assign n22393 = x628 | n22387 ;
  assign n22394 = x628 & ~n22353 ;
  assign n22395 = n22393 & ~n22394 ;
  assign n22396 = ( x792 & x1156 ) | ( x792 & ~n22395 ) | ( x1156 & ~n22395 ) ;
  assign n22397 = ~n22392 & n22396 ;
  assign n22398 = n22388 & ~n22397 ;
  assign n22399 = x787 | n22398 ;
  assign n22400 = x647 & ~n22398 ;
  assign n22401 = x647 | n22353 ;
  assign n22402 = ~n22400 & n22401 ;
  assign n22403 = ( ~x787 & x1157 ) | ( ~x787 & n22402 ) | ( x1157 & n22402 ) ;
  assign n22404 = x647 | n22398 ;
  assign n22405 = x647 & ~n22353 ;
  assign n22406 = n22404 & ~n22405 ;
  assign n22407 = ( x787 & x1157 ) | ( x787 & ~n22406 ) | ( x1157 & ~n22406 ) ;
  assign n22408 = ~n22403 & n22407 ;
  assign n22409 = n22399 & ~n22408 ;
  assign n22410 = x644 | n22409 ;
  assign n22411 = x715 & n22410 ;
  assign n22412 = x176 & n2032 ;
  assign n22413 = x742 & n22359 ;
  assign n22414 = ( x176 & ~x742 ) | ( x176 & n17421 ) | ( ~x742 & n17421 ) ;
  assign n22415 = n17415 | n17416 ;
  assign n22416 = ( x176 & x742 ) | ( x176 & n22415 ) | ( x742 & n22415 ) ;
  assign n22417 = n22414 & ~n22416 ;
  assign n22418 = n22413 | n22417 ;
  assign n22419 = ~n2032 & n22418 ;
  assign n22420 = n22412 | n22419 ;
  assign n22421 = ~n15082 & n22420 ;
  assign n22422 = n15082 & n22353 ;
  assign n22423 = n22421 | n22422 ;
  assign n22424 = ~x785 & n22423 ;
  assign n22425 = ~n15088 & n22353 ;
  assign n22426 = x609 & n22421 ;
  assign n22427 = n22425 | n22426 ;
  assign n22428 = x1155 & n22427 ;
  assign n22429 = n15094 & n22353 ;
  assign n22430 = ~x609 & n22421 ;
  assign n22431 = n22429 | n22430 ;
  assign n22432 = ~x1155 & n22431 ;
  assign n22433 = n22428 | n22432 ;
  assign n22434 = x785 & n22433 ;
  assign n22435 = n22424 | n22434 ;
  assign n22436 = ~x781 & n22435 ;
  assign n22437 = ( x618 & x1154 ) | ( x618 & n22353 ) | ( x1154 & n22353 ) ;
  assign n22438 = ( ~x618 & x1154 ) | ( ~x618 & n22435 ) | ( x1154 & n22435 ) ;
  assign n22439 = n22437 & n22438 ;
  assign n22440 = ( x618 & x1154 ) | ( x618 & ~n22353 ) | ( x1154 & ~n22353 ) ;
  assign n22441 = ( x618 & ~x1154 ) | ( x618 & n22435 ) | ( ~x1154 & n22435 ) ;
  assign n22442 = ~n22440 & n22441 ;
  assign n22443 = n22439 | n22442 ;
  assign n22444 = x781 & n22443 ;
  assign n22445 = n22436 | n22444 ;
  assign n22446 = ~x789 & n22445 ;
  assign n22447 = ( x619 & x1159 ) | ( x619 & n22353 ) | ( x1159 & n22353 ) ;
  assign n22448 = ( ~x619 & x1159 ) | ( ~x619 & n22445 ) | ( x1159 & n22445 ) ;
  assign n22449 = n22447 & n22448 ;
  assign n22450 = ( x619 & x1159 ) | ( x619 & ~n22353 ) | ( x1159 & ~n22353 ) ;
  assign n22451 = ( x619 & ~x1159 ) | ( x619 & n22445 ) | ( ~x1159 & n22445 ) ;
  assign n22452 = ~n22450 & n22451 ;
  assign n22453 = n22449 | n22452 ;
  assign n22454 = x789 & n22453 ;
  assign n22455 = n22446 | n22454 ;
  assign n22456 = n16176 | n22455 ;
  assign n22457 = n16176 & ~n22353 ;
  assign n22458 = n22456 & ~n22457 ;
  assign n22459 = n15134 | n22458 ;
  assign n22460 = n15134 & ~n22353 ;
  assign n22461 = n22459 & ~n22460 ;
  assign n22462 = n15141 | n22461 ;
  assign n22463 = n15141 & ~n22353 ;
  assign n22464 = n22462 & ~n22463 ;
  assign n22465 = ( x644 & x715 ) | ( x644 & ~n22464 ) | ( x715 & ~n22464 ) ;
  assign n22466 = ( x644 & ~x715 ) | ( x644 & n22353 ) | ( ~x715 & n22353 ) ;
  assign n22467 = ~n22465 & n22466 ;
  assign n22468 = x1160 & ~n22467 ;
  assign n22469 = ~n22411 & n22468 ;
  assign n22470 = x644 & ~n22409 ;
  assign n22471 = x715 | n22470 ;
  assign n22472 = ( x644 & x715 ) | ( x644 & n22464 ) | ( x715 & n22464 ) ;
  assign n22473 = ( ~x644 & x715 ) | ( ~x644 & n22353 ) | ( x715 & n22353 ) ;
  assign n22474 = n22472 & n22473 ;
  assign n22475 = x1160 | n22474 ;
  assign n22476 = n22471 & ~n22475 ;
  assign n22477 = n22469 | n22476 ;
  assign n22478 = x790 & n22477 ;
  assign n22479 = n15138 & n22402 ;
  assign n22480 = n15139 & n22406 ;
  assign n22481 = n18610 & n22461 ;
  assign n22482 = n22480 | n22481 ;
  assign n22483 = n22479 | n22482 ;
  assign n22484 = x787 & n22483 ;
  assign n22485 = n18621 & n22458 ;
  assign n22486 = n15132 & n22395 ;
  assign n22487 = n15131 & n22391 ;
  assign n22488 = n22486 | n22487 ;
  assign n22489 = n22485 | n22488 ;
  assign n22490 = x792 & n22489 ;
  assign n22491 = n16115 & ~n22384 ;
  assign n22492 = ( x626 & ~n15419 ) | ( x626 & n22353 ) | ( ~n15419 & n22353 ) ;
  assign n22493 = ( x626 & n15419 ) | ( x626 & ~n22455 ) | ( n15419 & ~n22455 ) ;
  assign n22494 = ~n22492 & n22493 ;
  assign n22495 = n22491 | n22494 ;
  assign n22496 = ( x626 & n15418 ) | ( x626 & ~n22353 ) | ( n15418 & ~n22353 ) ;
  assign n22497 = ( x626 & ~n15418 ) | ( x626 & n22455 ) | ( ~n15418 & n22455 ) ;
  assign n22498 = n22496 & ~n22497 ;
  assign n22499 = n22495 | n22498 ;
  assign n22500 = x788 & n22499 ;
  assign n22501 = x648 & ~n22452 ;
  assign n22502 = ( x619 & x1159 ) | ( x619 & n22382 ) | ( x1159 & n22382 ) ;
  assign n22503 = x627 | n22439 ;
  assign n22504 = ( x618 & x1154 ) | ( x618 & ~n22379 ) | ( x1154 & ~n22379 ) ;
  assign n22505 = x660 | n22428 ;
  assign n22506 = ( x609 & x1155 ) | ( x609 & ~n22376 ) | ( x1155 & ~n22376 ) ;
  assign n22507 = x608 | n22370 ;
  assign n22508 = ( x625 & x1153 ) | ( x625 & ~n22420 ) | ( x1153 & ~n22420 ) ;
  assign n22509 = x704 & ~n22418 ;
  assign n22510 = ( x176 & ~x742 ) | ( x176 & n17554 ) | ( ~x742 & n17554 ) ;
  assign n22511 = ( x176 & x742 ) | ( x176 & n17562 ) | ( x742 & n17562 ) ;
  assign n22512 = n22510 & ~n22511 ;
  assign n22513 = x704 | n22512 ;
  assign n22514 = n17569 | n17570 ;
  assign n22515 = ( x176 & ~x742 ) | ( x176 & n22514 ) | ( ~x742 & n22514 ) ;
  assign n22516 = ( x176 & x742 ) | ( x176 & n17579 ) | ( x742 & n17579 ) ;
  assign n22517 = ~n22515 & n22516 ;
  assign n22518 = n22513 | n22517 ;
  assign n22519 = ~n2032 & n22518 ;
  assign n22520 = ~n22509 & n22519 ;
  assign n22521 = n22412 | n22520 ;
  assign n22522 = ( x625 & ~x1153 ) | ( x625 & n22521 ) | ( ~x1153 & n22521 ) ;
  assign n22523 = ~n22508 & n22522 ;
  assign n22524 = n22507 | n22523 ;
  assign n22525 = x608 & ~n22373 ;
  assign n22526 = ( x625 & x1153 ) | ( x625 & n22420 ) | ( x1153 & n22420 ) ;
  assign n22527 = ( ~x625 & x1153 ) | ( ~x625 & n22521 ) | ( x1153 & n22521 ) ;
  assign n22528 = n22526 & n22527 ;
  assign n22529 = n22525 & ~n22528 ;
  assign n22530 = n22524 & ~n22529 ;
  assign n22531 = x778 & ~n22530 ;
  assign n22532 = x778 | n22521 ;
  assign n22533 = ~n22531 & n22532 ;
  assign n22534 = ( x609 & ~x1155 ) | ( x609 & n22533 ) | ( ~x1155 & n22533 ) ;
  assign n22535 = ~n22506 & n22534 ;
  assign n22536 = n22505 | n22535 ;
  assign n22537 = x660 & ~n22432 ;
  assign n22538 = ( x609 & x1155 ) | ( x609 & n22376 ) | ( x1155 & n22376 ) ;
  assign n22539 = ( ~x609 & x1155 ) | ( ~x609 & n22533 ) | ( x1155 & n22533 ) ;
  assign n22540 = n22538 & n22539 ;
  assign n22541 = n22537 & ~n22540 ;
  assign n22542 = n22536 & ~n22541 ;
  assign n22543 = x785 & ~n22542 ;
  assign n22544 = x785 | n22533 ;
  assign n22545 = ~n22543 & n22544 ;
  assign n22546 = ( x618 & ~x1154 ) | ( x618 & n22545 ) | ( ~x1154 & n22545 ) ;
  assign n22547 = ~n22504 & n22546 ;
  assign n22548 = n22503 | n22547 ;
  assign n22549 = x627 & ~n22442 ;
  assign n22550 = ( x618 & x1154 ) | ( x618 & n22379 ) | ( x1154 & n22379 ) ;
  assign n22551 = ( ~x618 & x1154 ) | ( ~x618 & n22545 ) | ( x1154 & n22545 ) ;
  assign n22552 = n22550 & n22551 ;
  assign n22553 = n22549 & ~n22552 ;
  assign n22554 = n22548 & ~n22553 ;
  assign n22555 = x781 & ~n22554 ;
  assign n22556 = x781 | n22545 ;
  assign n22557 = ~n22555 & n22556 ;
  assign n22558 = ( ~x619 & x1159 ) | ( ~x619 & n22557 ) | ( x1159 & n22557 ) ;
  assign n22559 = n22502 & n22558 ;
  assign n22560 = n22501 & ~n22559 ;
  assign n22561 = x648 | n22449 ;
  assign n22562 = ( x619 & x1159 ) | ( x619 & ~n22382 ) | ( x1159 & ~n22382 ) ;
  assign n22563 = ( x619 & ~x1159 ) | ( x619 & n22557 ) | ( ~x1159 & n22557 ) ;
  assign n22564 = ~n22562 & n22563 ;
  assign n22565 = n22561 | n22564 ;
  assign n22566 = x789 & n22565 ;
  assign n22567 = ~n22560 & n22566 ;
  assign n22568 = ~x789 & n22557 ;
  assign n22569 = n16177 | n22568 ;
  assign n22570 = n22567 | n22569 ;
  assign n22571 = ~n22500 & n22570 ;
  assign n22572 = n22490 | n22571 ;
  assign n22573 = n18431 | n18434 ;
  assign n22574 = ( n18431 & ~n22489 ) | ( n18431 & n22573 ) | ( ~n22489 & n22573 ) ;
  assign n22575 = n22572 & ~n22574 ;
  assign n22576 = n22484 | n22575 ;
  assign n22577 = ( x644 & ~x790 ) | ( x644 & n22468 ) | ( ~x790 & n22468 ) ;
  assign n22578 = ( x644 & x790 ) | ( x644 & n22475 ) | ( x790 & n22475 ) ;
  assign n22579 = ~n22577 & n22578 ;
  assign n22580 = n22576 | n22579 ;
  assign n22581 = ~n22478 & n22580 ;
  assign n22582 = ( ~x832 & n6785 ) | ( ~x832 & n22581 ) | ( n6785 & n22581 ) ;
  assign n22583 = ( ~x176 & x832 ) | ( ~x176 & n6785 ) | ( x832 & n6785 ) ;
  assign n22584 = n22582 & ~n22583 ;
  assign n22585 = n22352 | n22584 ;
  assign n22586 = x177 | n14834 ;
  assign n22587 = n15141 & n22586 ;
  assign n22588 = x177 & n2032 ;
  assign n22589 = x757 | n17421 ;
  assign n22590 = ~n19618 & n22589 ;
  assign n22591 = x177 | n22590 ;
  assign n22592 = x177 | n17415 ;
  assign n22593 = ~x757 & n22592 ;
  assign n22594 = n22415 & n22593 ;
  assign n22595 = n22591 & ~n22594 ;
  assign n22596 = ~n2032 & n22595 ;
  assign n22597 = n22588 | n22596 ;
  assign n22598 = ~n15082 & n22597 ;
  assign n22599 = n15082 & n22586 ;
  assign n22600 = n22598 | n22599 ;
  assign n22601 = ~x785 & n22600 ;
  assign n22602 = ~n15088 & n22586 ;
  assign n22603 = x609 & n22598 ;
  assign n22604 = n22602 | n22603 ;
  assign n22605 = x1155 & n22604 ;
  assign n22606 = n15094 & n22586 ;
  assign n22607 = ~x609 & n22598 ;
  assign n22608 = n22606 | n22607 ;
  assign n22609 = ~x1155 & n22608 ;
  assign n22610 = n22605 | n22609 ;
  assign n22611 = x785 & n22610 ;
  assign n22612 = n22601 | n22611 ;
  assign n22613 = ~x781 & n22612 ;
  assign n22614 = ( x618 & x1154 ) | ( x618 & n22586 ) | ( x1154 & n22586 ) ;
  assign n22615 = ( ~x618 & x1154 ) | ( ~x618 & n22612 ) | ( x1154 & n22612 ) ;
  assign n22616 = n22614 & n22615 ;
  assign n22617 = ( x618 & x1154 ) | ( x618 & ~n22586 ) | ( x1154 & ~n22586 ) ;
  assign n22618 = ( x618 & ~x1154 ) | ( x618 & n22612 ) | ( ~x1154 & n22612 ) ;
  assign n22619 = ~n22617 & n22618 ;
  assign n22620 = n22616 | n22619 ;
  assign n22621 = x781 & n22620 ;
  assign n22622 = n22613 | n22621 ;
  assign n22623 = ~x789 & n22622 ;
  assign n22624 = ( x619 & x1159 ) | ( x619 & n22586 ) | ( x1159 & n22586 ) ;
  assign n22625 = ( ~x619 & x1159 ) | ( ~x619 & n22622 ) | ( x1159 & n22622 ) ;
  assign n22626 = n22624 & n22625 ;
  assign n22627 = ( x619 & x1159 ) | ( x619 & ~n22586 ) | ( x1159 & ~n22586 ) ;
  assign n22628 = ( x619 & ~x1159 ) | ( x619 & n22622 ) | ( ~x1159 & n22622 ) ;
  assign n22629 = ~n22627 & n22628 ;
  assign n22630 = n22626 | n22629 ;
  assign n22631 = x789 & n22630 ;
  assign n22632 = n22623 | n22631 ;
  assign n22633 = n16176 | n22632 ;
  assign n22634 = n16176 & ~n22586 ;
  assign n22635 = n22633 & ~n22634 ;
  assign n22636 = n15134 | n22635 ;
  assign n22637 = n15134 & ~n22586 ;
  assign n22638 = n22636 & ~n22637 ;
  assign n22639 = ~n15141 & n22638 ;
  assign n22640 = n22587 | n22639 ;
  assign n22641 = ( x644 & x715 ) | ( x644 & n22640 ) | ( x715 & n22640 ) ;
  assign n22642 = ( ~x644 & x715 ) | ( ~x644 & n22586 ) | ( x715 & n22586 ) ;
  assign n22643 = n22641 & n22642 ;
  assign n22644 = x1160 | n22643 ;
  assign n22645 = n15414 & n22586 ;
  assign n22646 = x177 | n15070 ;
  assign n22647 = n15375 & n22646 ;
  assign n22648 = x686 | n22647 ;
  assign n22649 = ( ~x38 & x177 ) | ( ~x38 & n16319 ) | ( x177 & n16319 ) ;
  assign n22650 = ( x38 & x177 ) | ( x38 & n16323 ) | ( x177 & n16323 ) ;
  assign n22651 = n22649 & ~n22650 ;
  assign n22652 = n22648 | n22651 ;
  assign n22653 = ~x177 & x686 ;
  assign n22654 = ~n15382 & n22653 ;
  assign n22655 = n2032 | n22654 ;
  assign n22656 = n22652 & ~n22655 ;
  assign n22657 = n22588 | n22656 ;
  assign n22658 = ~x778 & n22657 ;
  assign n22659 = ( x625 & x1153 ) | ( x625 & n22586 ) | ( x1153 & n22586 ) ;
  assign n22660 = ( ~x625 & x1153 ) | ( ~x625 & n22657 ) | ( x1153 & n22657 ) ;
  assign n22661 = n22659 & n22660 ;
  assign n22662 = ( x625 & x1153 ) | ( x625 & ~n22586 ) | ( x1153 & ~n22586 ) ;
  assign n22663 = ( x625 & ~x1153 ) | ( x625 & n22657 ) | ( ~x1153 & n22657 ) ;
  assign n22664 = ~n22662 & n22663 ;
  assign n22665 = n22661 | n22664 ;
  assign n22666 = x778 & n22665 ;
  assign n22667 = n22658 | n22666 ;
  assign n22668 = ~n15400 & n22667 ;
  assign n22669 = n15400 & n22586 ;
  assign n22670 = n22668 | n22669 ;
  assign n22671 = n15407 | n22670 ;
  assign n22672 = n15407 & ~n22586 ;
  assign n22673 = n22671 & ~n22672 ;
  assign n22674 = ~n15414 & n22673 ;
  assign n22675 = n22645 | n22674 ;
  assign n22676 = n15421 | n22675 ;
  assign n22677 = n15421 & ~n22586 ;
  assign n22678 = n22676 & ~n22677 ;
  assign n22679 = ~x792 & n22678 ;
  assign n22680 = ( x628 & x1156 ) | ( x628 & n22586 ) | ( x1156 & n22586 ) ;
  assign n22681 = ( ~x628 & x1156 ) | ( ~x628 & n22678 ) | ( x1156 & n22678 ) ;
  assign n22682 = n22680 & n22681 ;
  assign n22683 = ( x628 & x1156 ) | ( x628 & ~n22586 ) | ( x1156 & ~n22586 ) ;
  assign n22684 = ( x628 & ~x1156 ) | ( x628 & n22678 ) | ( ~x1156 & n22678 ) ;
  assign n22685 = ~n22683 & n22684 ;
  assign n22686 = n22682 | n22685 ;
  assign n22687 = x792 & n22686 ;
  assign n22688 = n22679 | n22687 ;
  assign n22689 = ~x787 & n22688 ;
  assign n22690 = ( x647 & x1157 ) | ( x647 & n22586 ) | ( x1157 & n22586 ) ;
  assign n22691 = ( ~x647 & x1157 ) | ( ~x647 & n22688 ) | ( x1157 & n22688 ) ;
  assign n22692 = n22690 & n22691 ;
  assign n22693 = ( x647 & x1157 ) | ( x647 & ~n22586 ) | ( x1157 & ~n22586 ) ;
  assign n22694 = ( x647 & ~x1157 ) | ( x647 & n22688 ) | ( ~x1157 & n22688 ) ;
  assign n22695 = ~n22693 & n22694 ;
  assign n22696 = n22692 | n22695 ;
  assign n22697 = x787 & n22696 ;
  assign n22698 = n22689 | n22697 ;
  assign n22699 = ( x644 & x715 ) | ( x644 & ~n22698 ) | ( x715 & ~n22698 ) ;
  assign n22700 = x630 | n22692 ;
  assign n22701 = ( x647 & x1157 ) | ( x647 & ~n22638 ) | ( x1157 & ~n22638 ) ;
  assign n22702 = x629 | n22682 ;
  assign n22703 = ( x628 & x1156 ) | ( x628 & ~n22635 ) | ( x1156 & ~n22635 ) ;
  assign n22704 = x648 | n22626 ;
  assign n22705 = ( x619 & x1159 ) | ( x619 & ~n22673 ) | ( x1159 & ~n22673 ) ;
  assign n22706 = x627 | n22616 ;
  assign n22707 = ( x618 & x1154 ) | ( x618 & ~n22670 ) | ( x1154 & ~n22670 ) ;
  assign n22708 = x660 | n22605 ;
  assign n22709 = ( x609 & x1155 ) | ( x609 & ~n22667 ) | ( x1155 & ~n22667 ) ;
  assign n22710 = x608 | n22661 ;
  assign n22711 = ( x625 & x1153 ) | ( x625 & ~n22597 ) | ( x1153 & ~n22597 ) ;
  assign n22712 = n16404 & n22646 ;
  assign n22713 = x757 & ~n22712 ;
  assign n22714 = ( ~x38 & x177 ) | ( ~x38 & n17577 ) | ( x177 & n17577 ) ;
  assign n22715 = ( x38 & x177 ) | ( x38 & n17568 ) | ( x177 & n17568 ) ;
  assign n22716 = n22714 & ~n22715 ;
  assign n22717 = n22713 & ~n22716 ;
  assign n22718 = ( x38 & x177 ) | ( x38 & n17550 ) | ( x177 & n17550 ) ;
  assign n22719 = ( ~x38 & x177 ) | ( ~x38 & n17556 ) | ( x177 & n17556 ) ;
  assign n22720 = n22718 & ~n22719 ;
  assign n22721 = x757 | n22720 ;
  assign n22722 = ~n17549 & n17552 ;
  assign n22723 = ( ~x38 & x177 ) | ( ~x38 & n22722 ) | ( x177 & n22722 ) ;
  assign n22724 = ( x38 & x177 ) | ( x38 & n17560 ) | ( x177 & n17560 ) ;
  assign n22725 = n22723 & ~n22724 ;
  assign n22726 = n22721 | n22725 ;
  assign n22727 = ~n22717 & n22726 ;
  assign n22728 = ( x686 & ~n2032 ) | ( x686 & n22727 ) | ( ~n2032 & n22727 ) ;
  assign n22729 = ( x686 & n2032 ) | ( x686 & ~n22595 ) | ( n2032 & ~n22595 ) ;
  assign n22730 = n22728 & ~n22729 ;
  assign n22731 = n22588 | n22730 ;
  assign n22732 = ( x625 & ~x1153 ) | ( x625 & n22731 ) | ( ~x1153 & n22731 ) ;
  assign n22733 = ~n22711 & n22732 ;
  assign n22734 = n22710 | n22733 ;
  assign n22735 = x608 & ~n22664 ;
  assign n22736 = ( x625 & x1153 ) | ( x625 & n22597 ) | ( x1153 & n22597 ) ;
  assign n22737 = ( ~x625 & x1153 ) | ( ~x625 & n22731 ) | ( x1153 & n22731 ) ;
  assign n22738 = n22736 & n22737 ;
  assign n22739 = n22735 & ~n22738 ;
  assign n22740 = n22734 & ~n22739 ;
  assign n22741 = x778 & ~n22740 ;
  assign n22742 = x778 | n22731 ;
  assign n22743 = ~n22741 & n22742 ;
  assign n22744 = ( x609 & ~x1155 ) | ( x609 & n22743 ) | ( ~x1155 & n22743 ) ;
  assign n22745 = ~n22709 & n22744 ;
  assign n22746 = n22708 | n22745 ;
  assign n22747 = x660 & ~n22609 ;
  assign n22748 = ( x609 & x1155 ) | ( x609 & n22667 ) | ( x1155 & n22667 ) ;
  assign n22749 = ( ~x609 & x1155 ) | ( ~x609 & n22743 ) | ( x1155 & n22743 ) ;
  assign n22750 = n22748 & n22749 ;
  assign n22751 = n22747 & ~n22750 ;
  assign n22752 = n22746 & ~n22751 ;
  assign n22753 = x785 & ~n22752 ;
  assign n22754 = x785 | n22743 ;
  assign n22755 = ~n22753 & n22754 ;
  assign n22756 = ( x618 & ~x1154 ) | ( x618 & n22755 ) | ( ~x1154 & n22755 ) ;
  assign n22757 = ~n22707 & n22756 ;
  assign n22758 = n22706 | n22757 ;
  assign n22759 = x627 & ~n22619 ;
  assign n22760 = ( x618 & x1154 ) | ( x618 & n22670 ) | ( x1154 & n22670 ) ;
  assign n22761 = ( ~x618 & x1154 ) | ( ~x618 & n22755 ) | ( x1154 & n22755 ) ;
  assign n22762 = n22760 & n22761 ;
  assign n22763 = n22759 & ~n22762 ;
  assign n22764 = n22758 & ~n22763 ;
  assign n22765 = x781 & ~n22764 ;
  assign n22766 = x781 | n22755 ;
  assign n22767 = ~n22765 & n22766 ;
  assign n22768 = ( x619 & ~x1159 ) | ( x619 & n22767 ) | ( ~x1159 & n22767 ) ;
  assign n22769 = ~n22705 & n22768 ;
  assign n22770 = n22704 | n22769 ;
  assign n22771 = x648 & ~n22629 ;
  assign n22772 = ( x619 & x1159 ) | ( x619 & n22673 ) | ( x1159 & n22673 ) ;
  assign n22773 = ( ~x619 & x1159 ) | ( ~x619 & n22767 ) | ( x1159 & n22767 ) ;
  assign n22774 = n22772 & n22773 ;
  assign n22775 = n22771 & ~n22774 ;
  assign n22776 = n22770 & ~n22775 ;
  assign n22777 = x789 & ~n22776 ;
  assign n22778 = x789 | n22767 ;
  assign n22779 = ~n22777 & n22778 ;
  assign n22780 = ~x788 & n22779 ;
  assign n22781 = ( x626 & x641 ) | ( x626 & ~n22632 ) | ( x641 & ~n22632 ) ;
  assign n22782 = ( x626 & ~x641 ) | ( x626 & n22586 ) | ( ~x641 & n22586 ) ;
  assign n22783 = n22781 & ~n22782 ;
  assign n22784 = x1158 | n22783 ;
  assign n22785 = ( x626 & x641 ) | ( x626 & n22675 ) | ( x641 & n22675 ) ;
  assign n22786 = ( ~x626 & x641 ) | ( ~x626 & n22779 ) | ( x641 & n22779 ) ;
  assign n22787 = n22785 | n22786 ;
  assign n22788 = ~n22784 & n22787 ;
  assign n22789 = ( x626 & x641 ) | ( x626 & n22632 ) | ( x641 & n22632 ) ;
  assign n22790 = ( ~x626 & x641 ) | ( ~x626 & n22586 ) | ( x641 & n22586 ) ;
  assign n22791 = n22789 | n22790 ;
  assign n22792 = x1158 & n22791 ;
  assign n22793 = ( x626 & x641 ) | ( x626 & ~n22675 ) | ( x641 & ~n22675 ) ;
  assign n22794 = ( x626 & ~x641 ) | ( x626 & n22779 ) | ( ~x641 & n22779 ) ;
  assign n22795 = n22793 & ~n22794 ;
  assign n22796 = n22792 & ~n22795 ;
  assign n22797 = n22788 | n22796 ;
  assign n22798 = x788 & n22797 ;
  assign n22799 = n22780 | n22798 ;
  assign n22800 = ( x628 & ~x1156 ) | ( x628 & n22799 ) | ( ~x1156 & n22799 ) ;
  assign n22801 = ~n22703 & n22800 ;
  assign n22802 = n22702 | n22801 ;
  assign n22803 = x629 & ~n22685 ;
  assign n22804 = ( x628 & x1156 ) | ( x628 & n22635 ) | ( x1156 & n22635 ) ;
  assign n22805 = ( ~x628 & x1156 ) | ( ~x628 & n22799 ) | ( x1156 & n22799 ) ;
  assign n22806 = n22804 & n22805 ;
  assign n22807 = n22803 & ~n22806 ;
  assign n22808 = n22802 & ~n22807 ;
  assign n22809 = x792 & ~n22808 ;
  assign n22810 = x792 | n22799 ;
  assign n22811 = ~n22809 & n22810 ;
  assign n22812 = ( x647 & ~x1157 ) | ( x647 & n22811 ) | ( ~x1157 & n22811 ) ;
  assign n22813 = ~n22701 & n22812 ;
  assign n22814 = n22700 | n22813 ;
  assign n22815 = x630 & ~n22695 ;
  assign n22816 = ( x647 & x1157 ) | ( x647 & n22638 ) | ( x1157 & n22638 ) ;
  assign n22817 = ( ~x647 & x1157 ) | ( ~x647 & n22811 ) | ( x1157 & n22811 ) ;
  assign n22818 = n22816 & n22817 ;
  assign n22819 = n22815 & ~n22818 ;
  assign n22820 = n22814 & ~n22819 ;
  assign n22821 = x787 & ~n22820 ;
  assign n22822 = x787 | n22811 ;
  assign n22823 = ~n22821 & n22822 ;
  assign n22824 = ( x644 & ~x715 ) | ( x644 & n22823 ) | ( ~x715 & n22823 ) ;
  assign n22825 = ~n22699 & n22824 ;
  assign n22826 = n22644 | n22825 ;
  assign n22827 = ( x644 & x715 ) | ( x644 & ~n22640 ) | ( x715 & ~n22640 ) ;
  assign n22828 = ( x644 & ~x715 ) | ( x644 & n22586 ) | ( ~x715 & n22586 ) ;
  assign n22829 = ~n22827 & n22828 ;
  assign n22830 = x1160 & ~n22829 ;
  assign n22831 = ( x644 & x715 ) | ( x644 & n22698 ) | ( x715 & n22698 ) ;
  assign n22832 = ( ~x644 & x715 ) | ( ~x644 & n22823 ) | ( x715 & n22823 ) ;
  assign n22833 = n22831 & n22832 ;
  assign n22834 = n22830 & ~n22833 ;
  assign n22835 = x790 & ~n22834 ;
  assign n22836 = n22826 & n22835 ;
  assign n22837 = ~x790 & n22823 ;
  assign n22838 = n6785 | n22837 ;
  assign n22839 = n22836 | n22838 ;
  assign n22840 = ~x177 & n6785 ;
  assign n22841 = x832 | n22840 ;
  assign n22842 = n22839 & ~n22841 ;
  assign n22843 = x177 | n1290 ;
  assign n22844 = ~x757 & n14840 ;
  assign n22845 = n22843 & ~n22844 ;
  assign n22846 = n16060 | n22845 ;
  assign n22847 = ~x785 & n22846 ;
  assign n22848 = n16065 | n22845 ;
  assign n22849 = x1155 & n22848 ;
  assign n22850 = n16068 | n22846 ;
  assign n22851 = ~x1155 & n22850 ;
  assign n22852 = n22849 | n22851 ;
  assign n22853 = x785 & n22852 ;
  assign n22854 = n22847 | n22853 ;
  assign n22855 = ~x781 & n22854 ;
  assign n22856 = n16075 | n22854 ;
  assign n22857 = x1154 & n22856 ;
  assign n22858 = n16078 | n22854 ;
  assign n22859 = ~x1154 & n22858 ;
  assign n22860 = n22857 | n22859 ;
  assign n22861 = x781 & n22860 ;
  assign n22862 = n22855 | n22861 ;
  assign n22863 = ~x789 & n22862 ;
  assign n22864 = ( x619 & x1159 ) | ( x619 & n22843 ) | ( x1159 & n22843 ) ;
  assign n22865 = ( ~x619 & x1159 ) | ( ~x619 & n22862 ) | ( x1159 & n22862 ) ;
  assign n22866 = n22864 & n22865 ;
  assign n22867 = ( x619 & x1159 ) | ( x619 & ~n22843 ) | ( x1159 & ~n22843 ) ;
  assign n22868 = ( x619 & ~x1159 ) | ( x619 & n22862 ) | ( ~x1159 & n22862 ) ;
  assign n22869 = ~n22867 & n22868 ;
  assign n22870 = n22866 | n22869 ;
  assign n22871 = x789 & n22870 ;
  assign n22872 = n22863 | n22871 ;
  assign n22873 = n16176 | n22872 ;
  assign n22874 = n16176 & ~n22843 ;
  assign n22875 = n22873 & ~n22874 ;
  assign n22876 = n15134 | n22875 ;
  assign n22877 = n15134 & ~n22843 ;
  assign n22878 = n22876 & ~n22877 ;
  assign n22879 = n18610 & n22878 ;
  assign n22880 = ( x647 & x1157 ) | ( x647 & ~n22843 ) | ( x1157 & ~n22843 ) ;
  assign n22881 = ~x686 & n15202 ;
  assign n22882 = n22843 & ~n22881 ;
  assign n22883 = ~x778 & n22882 ;
  assign n22884 = ~x625 & n22881 ;
  assign n22885 = n22882 | n22884 ;
  assign n22886 = x1153 & n22885 ;
  assign n22887 = ~x1153 & n22843 ;
  assign n22888 = ~n22884 & n22887 ;
  assign n22889 = n22886 | n22888 ;
  assign n22890 = x778 & n22889 ;
  assign n22891 = n22883 | n22890 ;
  assign n22892 = n16043 | n22891 ;
  assign n22893 = n16045 | n22892 ;
  assign n22894 = n16047 | n22893 ;
  assign n22895 = n16049 | n22894 ;
  assign n22896 = n16055 | n22895 ;
  assign n22897 = ( x647 & ~x1157 ) | ( x647 & n22896 ) | ( ~x1157 & n22896 ) ;
  assign n22898 = ~n22880 & n22897 ;
  assign n22899 = x630 & n22898 ;
  assign n22900 = x647 & n22896 ;
  assign n22901 = ~x647 & n22843 ;
  assign n22902 = n22900 | n22901 ;
  assign n22903 = n15138 & n22902 ;
  assign n22904 = n22899 | n22903 ;
  assign n22905 = n22879 | n22904 ;
  assign n22906 = x787 & n22905 ;
  assign n22907 = n16115 & ~n22894 ;
  assign n22908 = ( x626 & ~n15419 ) | ( x626 & n22843 ) | ( ~n15419 & n22843 ) ;
  assign n22909 = ( x626 & n15419 ) | ( x626 & ~n22872 ) | ( n15419 & ~n22872 ) ;
  assign n22910 = ~n22908 & n22909 ;
  assign n22911 = n22907 | n22910 ;
  assign n22912 = ( x626 & n15418 ) | ( x626 & ~n22843 ) | ( n15418 & ~n22843 ) ;
  assign n22913 = ( x626 & ~n15418 ) | ( x626 & n22872 ) | ( ~n15418 & n22872 ) ;
  assign n22914 = n22912 & ~n22913 ;
  assign n22915 = n22911 | n22914 ;
  assign n22916 = x788 & n22915 ;
  assign n22917 = x648 & ~n22869 ;
  assign n22918 = ( x619 & x1159 ) | ( x619 & n22893 ) | ( x1159 & n22893 ) ;
  assign n22919 = x627 | n22857 ;
  assign n22920 = ( x618 & x1154 ) | ( x618 & ~n22892 ) | ( x1154 & ~n22892 ) ;
  assign n22921 = x660 | n22849 ;
  assign n22922 = ( x609 & x1155 ) | ( x609 & ~n22891 ) | ( x1155 & ~n22891 ) ;
  assign n22923 = n14839 | n22882 ;
  assign n22924 = x625 & ~n22923 ;
  assign n22925 = n22845 & n22923 ;
  assign n22926 = n22924 | n22925 ;
  assign n22927 = n22887 & n22926 ;
  assign n22928 = x608 | n22886 ;
  assign n22929 = n22927 | n22928 ;
  assign n22930 = x1153 & n22845 ;
  assign n22931 = ~n22924 & n22930 ;
  assign n22932 = x608 & ~n22888 ;
  assign n22933 = ~n22931 & n22932 ;
  assign n22934 = n22929 & ~n22933 ;
  assign n22935 = x778 & ~n22934 ;
  assign n22936 = x778 | n22925 ;
  assign n22937 = ~n22935 & n22936 ;
  assign n22938 = ( x609 & ~x1155 ) | ( x609 & n22937 ) | ( ~x1155 & n22937 ) ;
  assign n22939 = ~n22922 & n22938 ;
  assign n22940 = n22921 | n22939 ;
  assign n22941 = x660 & ~n22851 ;
  assign n22942 = ( x609 & x1155 ) | ( x609 & n22891 ) | ( x1155 & n22891 ) ;
  assign n22943 = ( ~x609 & x1155 ) | ( ~x609 & n22937 ) | ( x1155 & n22937 ) ;
  assign n22944 = n22942 & n22943 ;
  assign n22945 = n22941 & ~n22944 ;
  assign n22946 = n22940 & ~n22945 ;
  assign n22947 = x785 & ~n22946 ;
  assign n22948 = x785 | n22937 ;
  assign n22949 = ~n22947 & n22948 ;
  assign n22950 = ( x618 & ~x1154 ) | ( x618 & n22949 ) | ( ~x1154 & n22949 ) ;
  assign n22951 = ~n22920 & n22950 ;
  assign n22952 = n22919 | n22951 ;
  assign n22953 = x627 & ~n22859 ;
  assign n22954 = ( x618 & x1154 ) | ( x618 & n22892 ) | ( x1154 & n22892 ) ;
  assign n22955 = ( ~x618 & x1154 ) | ( ~x618 & n22949 ) | ( x1154 & n22949 ) ;
  assign n22956 = n22954 & n22955 ;
  assign n22957 = n22953 & ~n22956 ;
  assign n22958 = n22952 & ~n22957 ;
  assign n22959 = x781 & ~n22958 ;
  assign n22960 = x781 | n22949 ;
  assign n22961 = ~n22959 & n22960 ;
  assign n22962 = ( ~x619 & x1159 ) | ( ~x619 & n22961 ) | ( x1159 & n22961 ) ;
  assign n22963 = n22918 & n22962 ;
  assign n22964 = n22917 & ~n22963 ;
  assign n22965 = x648 | n22866 ;
  assign n22966 = ( x619 & x1159 ) | ( x619 & ~n22893 ) | ( x1159 & ~n22893 ) ;
  assign n22967 = ( x619 & ~x1159 ) | ( x619 & n22961 ) | ( ~x1159 & n22961 ) ;
  assign n22968 = ~n22966 & n22967 ;
  assign n22969 = n22965 | n22968 ;
  assign n22970 = x789 & n22969 ;
  assign n22971 = ~n22964 & n22970 ;
  assign n22972 = ~x789 & n22961 ;
  assign n22973 = n16177 | n22972 ;
  assign n22974 = n22971 | n22973 ;
  assign n22975 = ~n22916 & n22974 ;
  assign n22976 = n18434 | n22975 ;
  assign n22977 = n16650 | n22895 ;
  assign n22978 = n16051 & ~n22875 ;
  assign n22979 = n22977 & ~n22978 ;
  assign n22980 = ( x629 & ~x792 ) | ( x629 & n22979 ) | ( ~x792 & n22979 ) ;
  assign n22981 = n16052 & ~n22875 ;
  assign n22982 = n16643 & ~n22895 ;
  assign n22983 = n22981 | n22982 ;
  assign n22984 = ( x629 & x792 ) | ( x629 & n22983 ) | ( x792 & n22983 ) ;
  assign n22985 = ~n22980 & n22984 ;
  assign n22986 = n18431 | n22985 ;
  assign n22987 = n22976 & ~n22986 ;
  assign n22988 = n22906 | n22987 ;
  assign n22989 = ( x790 & x832 ) | ( x790 & n22988 ) | ( x832 & n22988 ) ;
  assign n22990 = n15141 | n22878 ;
  assign n22991 = n15141 & ~n22843 ;
  assign n22992 = n22990 & ~n22991 ;
  assign n22993 = ( x644 & x715 ) | ( x644 & ~n22992 ) | ( x715 & ~n22992 ) ;
  assign n22994 = ( x644 & ~x715 ) | ( x644 & n22843 ) | ( ~x715 & n22843 ) ;
  assign n22995 = ~n22993 & n22994 ;
  assign n22996 = x1160 & ~n22995 ;
  assign n22997 = ~x787 & n22896 ;
  assign n22998 = x1157 & n22902 ;
  assign n22999 = n22898 | n22998 ;
  assign n23000 = x787 & n22999 ;
  assign n23001 = n22997 | n23000 ;
  assign n23002 = ( x644 & x715 ) | ( x644 & n23001 ) | ( x715 & n23001 ) ;
  assign n23003 = ( ~x644 & x715 ) | ( ~x644 & n22988 ) | ( x715 & n22988 ) ;
  assign n23004 = n23002 & n23003 ;
  assign n23005 = n22996 & ~n23004 ;
  assign n23006 = ( x644 & x715 ) | ( x644 & n22992 ) | ( x715 & n22992 ) ;
  assign n23007 = ( ~x644 & x715 ) | ( ~x644 & n22843 ) | ( x715 & n22843 ) ;
  assign n23008 = n23006 & n23007 ;
  assign n23009 = x1160 | n23008 ;
  assign n23010 = ( x644 & x715 ) | ( x644 & ~n23001 ) | ( x715 & ~n23001 ) ;
  assign n23011 = ( x644 & ~x715 ) | ( x644 & n22988 ) | ( ~x715 & n22988 ) ;
  assign n23012 = ~n23010 & n23011 ;
  assign n23013 = n23009 | n23012 ;
  assign n23014 = ~n23005 & n23013 ;
  assign n23015 = ( ~x790 & x832 ) | ( ~x790 & n23014 ) | ( x832 & n23014 ) ;
  assign n23016 = n22989 & n23015 ;
  assign n23017 = n22842 | n23016 ;
  assign n23018 = x178 | n1290 ;
  assign n23019 = ~x760 & n14840 ;
  assign n23020 = n23018 & ~n23019 ;
  assign n23021 = n16060 | n23020 ;
  assign n23022 = ~x785 & n23021 ;
  assign n23023 = ~n15094 & n23019 ;
  assign n23024 = n23021 | n23023 ;
  assign n23025 = x1155 & n23024 ;
  assign n23026 = ~x1155 & n23018 ;
  assign n23027 = ~n23023 & n23026 ;
  assign n23028 = n23025 | n23027 ;
  assign n23029 = x785 & n23028 ;
  assign n23030 = n23022 | n23029 ;
  assign n23031 = ~x781 & n23030 ;
  assign n23032 = n16075 | n23030 ;
  assign n23033 = x1154 & n23032 ;
  assign n23034 = n16078 | n23030 ;
  assign n23035 = ~x1154 & n23034 ;
  assign n23036 = n23033 | n23035 ;
  assign n23037 = x781 & n23036 ;
  assign n23038 = n23031 | n23037 ;
  assign n23039 = ~x789 & n23038 ;
  assign n23040 = n20948 | n23038 ;
  assign n23041 = x1159 & n23040 ;
  assign n23042 = n20951 | n23038 ;
  assign n23043 = ~x1159 & n23042 ;
  assign n23044 = n23041 | n23043 ;
  assign n23045 = x789 & n23044 ;
  assign n23046 = n23039 | n23045 ;
  assign n23047 = n16176 | n23046 ;
  assign n23048 = n16176 & ~n23018 ;
  assign n23049 = n23047 & ~n23048 ;
  assign n23050 = n15134 | n23049 ;
  assign n23051 = n15134 & ~n23018 ;
  assign n23052 = n23050 & ~n23051 ;
  assign n23053 = n18610 & n23052 ;
  assign n23054 = ( x647 & x1157 ) | ( x647 & ~n23018 ) | ( x1157 & ~n23018 ) ;
  assign n23055 = ~x688 & n15202 ;
  assign n23056 = n23018 & ~n23055 ;
  assign n23057 = x778 | n23056 ;
  assign n23058 = ~x625 & n23055 ;
  assign n23059 = n23056 | n23058 ;
  assign n23060 = x1153 & n23059 ;
  assign n23061 = ~x1153 & n23018 ;
  assign n23062 = ~n23058 & n23061 ;
  assign n23063 = x778 & ~n23062 ;
  assign n23064 = ~n23060 & n23063 ;
  assign n23065 = n23057 & ~n23064 ;
  assign n23066 = n16043 | n23065 ;
  assign n23067 = n16045 | n23066 ;
  assign n23068 = n16047 | n23067 ;
  assign n23069 = n16049 | n23068 ;
  assign n23070 = n16055 | n23069 ;
  assign n23071 = ( x647 & ~x1157 ) | ( x647 & n23070 ) | ( ~x1157 & n23070 ) ;
  assign n23072 = ~n23054 & n23071 ;
  assign n23073 = x630 & n23072 ;
  assign n23074 = x647 & n23070 ;
  assign n23075 = ~x647 & n23018 ;
  assign n23076 = n23074 | n23075 ;
  assign n23077 = n15138 & n23076 ;
  assign n23078 = n23073 | n23077 ;
  assign n23079 = n23053 | n23078 ;
  assign n23080 = x787 & n23079 ;
  assign n23081 = n16115 & ~n23068 ;
  assign n23082 = ( x626 & ~n15419 ) | ( x626 & n23018 ) | ( ~n15419 & n23018 ) ;
  assign n23083 = ( x626 & n15419 ) | ( x626 & ~n23046 ) | ( n15419 & ~n23046 ) ;
  assign n23084 = ~n23082 & n23083 ;
  assign n23085 = n23081 | n23084 ;
  assign n23086 = ( x626 & n15418 ) | ( x626 & ~n23018 ) | ( n15418 & ~n23018 ) ;
  assign n23087 = ( x626 & ~n15418 ) | ( x626 & n23046 ) | ( ~n15418 & n23046 ) ;
  assign n23088 = n23086 & ~n23087 ;
  assign n23089 = n23085 | n23088 ;
  assign n23090 = x788 & n23089 ;
  assign n23091 = x648 & ~n23043 ;
  assign n23092 = ( x619 & x1159 ) | ( x619 & n23067 ) | ( x1159 & n23067 ) ;
  assign n23093 = x627 | n23033 ;
  assign n23094 = ( x618 & x1154 ) | ( x618 & ~n23066 ) | ( x1154 & ~n23066 ) ;
  assign n23095 = x660 | n23025 ;
  assign n23096 = ( x609 & x1155 ) | ( x609 & ~n23065 ) | ( x1155 & ~n23065 ) ;
  assign n23097 = n14839 | n23056 ;
  assign n23098 = x625 & ~n23097 ;
  assign n23099 = n23020 & n23097 ;
  assign n23100 = n23098 | n23099 ;
  assign n23101 = n23061 & n23100 ;
  assign n23102 = x608 | n23060 ;
  assign n23103 = n23101 | n23102 ;
  assign n23104 = x1153 & n23020 ;
  assign n23105 = ~n23098 & n23104 ;
  assign n23106 = x608 & ~n23062 ;
  assign n23107 = ~n23105 & n23106 ;
  assign n23108 = n23103 & ~n23107 ;
  assign n23109 = x778 & ~n23108 ;
  assign n23110 = x778 | n23099 ;
  assign n23111 = ~n23109 & n23110 ;
  assign n23112 = ( x609 & ~x1155 ) | ( x609 & n23111 ) | ( ~x1155 & n23111 ) ;
  assign n23113 = ~n23096 & n23112 ;
  assign n23114 = n23095 | n23113 ;
  assign n23115 = x660 & ~n23027 ;
  assign n23116 = ( x609 & x1155 ) | ( x609 & n23065 ) | ( x1155 & n23065 ) ;
  assign n23117 = ( ~x609 & x1155 ) | ( ~x609 & n23111 ) | ( x1155 & n23111 ) ;
  assign n23118 = n23116 & n23117 ;
  assign n23119 = n23115 & ~n23118 ;
  assign n23120 = n23114 & ~n23119 ;
  assign n23121 = x785 & ~n23120 ;
  assign n23122 = x785 | n23111 ;
  assign n23123 = ~n23121 & n23122 ;
  assign n23124 = ( x618 & ~x1154 ) | ( x618 & n23123 ) | ( ~x1154 & n23123 ) ;
  assign n23125 = ~n23094 & n23124 ;
  assign n23126 = n23093 | n23125 ;
  assign n23127 = x627 & ~n23035 ;
  assign n23128 = ( x618 & x1154 ) | ( x618 & n23066 ) | ( x1154 & n23066 ) ;
  assign n23129 = ( ~x618 & x1154 ) | ( ~x618 & n23123 ) | ( x1154 & n23123 ) ;
  assign n23130 = n23128 & n23129 ;
  assign n23131 = n23127 & ~n23130 ;
  assign n23132 = n23126 & ~n23131 ;
  assign n23133 = x781 & ~n23132 ;
  assign n23134 = x781 | n23123 ;
  assign n23135 = ~n23133 & n23134 ;
  assign n23136 = ( ~x619 & x1159 ) | ( ~x619 & n23135 ) | ( x1159 & n23135 ) ;
  assign n23137 = n23092 & n23136 ;
  assign n23138 = n23091 & ~n23137 ;
  assign n23139 = x648 | n23041 ;
  assign n23140 = ( x619 & x1159 ) | ( x619 & ~n23067 ) | ( x1159 & ~n23067 ) ;
  assign n23141 = ( x619 & ~x1159 ) | ( x619 & n23135 ) | ( ~x1159 & n23135 ) ;
  assign n23142 = ~n23140 & n23141 ;
  assign n23143 = n23139 | n23142 ;
  assign n23144 = x789 & n23143 ;
  assign n23145 = ~n23138 & n23144 ;
  assign n23146 = ~x789 & n23135 ;
  assign n23147 = n16177 | n23146 ;
  assign n23148 = n23145 | n23147 ;
  assign n23149 = ~n23090 & n23148 ;
  assign n23150 = n18434 | n23149 ;
  assign n23151 = n16650 | n23069 ;
  assign n23152 = n16051 & ~n23049 ;
  assign n23153 = n23151 & ~n23152 ;
  assign n23154 = ( x629 & ~x792 ) | ( x629 & n23153 ) | ( ~x792 & n23153 ) ;
  assign n23155 = n16052 & ~n23049 ;
  assign n23156 = n16643 & ~n23069 ;
  assign n23157 = n23155 | n23156 ;
  assign n23158 = ( x629 & x792 ) | ( x629 & n23157 ) | ( x792 & n23157 ) ;
  assign n23159 = ~n23154 & n23158 ;
  assign n23160 = n18431 | n23159 ;
  assign n23161 = n23150 & ~n23160 ;
  assign n23162 = n23080 | n23161 ;
  assign n23163 = ( x790 & x832 ) | ( x790 & n23162 ) | ( x832 & n23162 ) ;
  assign n23164 = n15141 | n23052 ;
  assign n23165 = n15141 & ~n23018 ;
  assign n23166 = n23164 & ~n23165 ;
  assign n23167 = ( x644 & x715 ) | ( x644 & ~n23166 ) | ( x715 & ~n23166 ) ;
  assign n23168 = ( x644 & ~x715 ) | ( x644 & n23018 ) | ( ~x715 & n23018 ) ;
  assign n23169 = ~n23167 & n23168 ;
  assign n23170 = x1160 & ~n23169 ;
  assign n23171 = ~x787 & n23070 ;
  assign n23172 = x1157 & n23076 ;
  assign n23173 = n23072 | n23172 ;
  assign n23174 = x787 & n23173 ;
  assign n23175 = n23171 | n23174 ;
  assign n23176 = ( x644 & x715 ) | ( x644 & n23175 ) | ( x715 & n23175 ) ;
  assign n23177 = ( ~x644 & x715 ) | ( ~x644 & n23162 ) | ( x715 & n23162 ) ;
  assign n23178 = n23176 & n23177 ;
  assign n23179 = n23170 & ~n23178 ;
  assign n23180 = ( x644 & x715 ) | ( x644 & n23166 ) | ( x715 & n23166 ) ;
  assign n23181 = ( ~x644 & x715 ) | ( ~x644 & n23018 ) | ( x715 & n23018 ) ;
  assign n23182 = n23180 & n23181 ;
  assign n23183 = x1160 | n23182 ;
  assign n23184 = ( x644 & x715 ) | ( x644 & ~n23175 ) | ( x715 & ~n23175 ) ;
  assign n23185 = ( x644 & ~x715 ) | ( x644 & n23162 ) | ( ~x715 & n23162 ) ;
  assign n23186 = ~n23184 & n23185 ;
  assign n23187 = n23183 | n23186 ;
  assign n23188 = ~n23179 & n23187 ;
  assign n23189 = ( ~x790 & x832 ) | ( ~x790 & n23188 ) | ( x832 & n23188 ) ;
  assign n23190 = n23163 & n23189 ;
  assign n23191 = x178 | n14834 ;
  assign n23192 = n15414 & n23191 ;
  assign n23193 = x688 | n2032 ;
  assign n23194 = ~n23191 & n23193 ;
  assign n23195 = x178 & n16323 ;
  assign n23196 = x38 | n23195 ;
  assign n23197 = ~n2032 & n23196 ;
  assign n23198 = x178 | n16319 ;
  assign n23199 = ~n23197 & n23198 ;
  assign n23200 = x178 | n15070 ;
  assign n23201 = n15375 & n23200 ;
  assign n23202 = x688 | n23201 ;
  assign n23203 = n23199 | n23202 ;
  assign n23204 = ~n23194 & n23203 ;
  assign n23205 = ~x778 & n23204 ;
  assign n23206 = ( x625 & x1153 ) | ( x625 & n23191 ) | ( x1153 & n23191 ) ;
  assign n23207 = ( ~x625 & x1153 ) | ( ~x625 & n23204 ) | ( x1153 & n23204 ) ;
  assign n23208 = n23206 & n23207 ;
  assign n23209 = ( x625 & x1153 ) | ( x625 & ~n23191 ) | ( x1153 & ~n23191 ) ;
  assign n23210 = ( x625 & ~x1153 ) | ( x625 & n23204 ) | ( ~x1153 & n23204 ) ;
  assign n23211 = ~n23209 & n23210 ;
  assign n23212 = n23208 | n23211 ;
  assign n23213 = x778 & n23212 ;
  assign n23214 = n23205 | n23213 ;
  assign n23215 = ~n15400 & n23214 ;
  assign n23216 = n15400 & n23191 ;
  assign n23217 = n23215 | n23216 ;
  assign n23218 = n15407 | n23217 ;
  assign n23219 = n15407 & ~n23191 ;
  assign n23220 = n23218 & ~n23219 ;
  assign n23221 = ~n15414 & n23220 ;
  assign n23222 = n23192 | n23221 ;
  assign n23223 = n15421 | n23222 ;
  assign n23224 = n15421 & ~n23191 ;
  assign n23225 = n23223 & ~n23224 ;
  assign n23226 = ~x792 & n23225 ;
  assign n23227 = ( x628 & x1156 ) | ( x628 & n23191 ) | ( x1156 & n23191 ) ;
  assign n23228 = ( ~x628 & x1156 ) | ( ~x628 & n23225 ) | ( x1156 & n23225 ) ;
  assign n23229 = n23227 & n23228 ;
  assign n23230 = ( x628 & x1156 ) | ( x628 & ~n23191 ) | ( x1156 & ~n23191 ) ;
  assign n23231 = ( x628 & ~x1156 ) | ( x628 & n23225 ) | ( ~x1156 & n23225 ) ;
  assign n23232 = ~n23230 & n23231 ;
  assign n23233 = n23229 | n23232 ;
  assign n23234 = x792 & n23233 ;
  assign n23235 = n23226 | n23234 ;
  assign n23236 = x787 | n23235 ;
  assign n23237 = x647 & n23235 ;
  assign n23238 = ~x647 & n23191 ;
  assign n23239 = n23237 | n23238 ;
  assign n23240 = ( ~x787 & x1157 ) | ( ~x787 & n23239 ) | ( x1157 & n23239 ) ;
  assign n23241 = ~x647 & n23235 ;
  assign n23242 = x647 & n23191 ;
  assign n23243 = n23241 | n23242 ;
  assign n23244 = ( x787 & x1157 ) | ( x787 & ~n23243 ) | ( x1157 & ~n23243 ) ;
  assign n23245 = ~n23240 & n23244 ;
  assign n23246 = n23236 & ~n23245 ;
  assign n23247 = x644 | n23246 ;
  assign n23248 = x715 & n23247 ;
  assign n23249 = x178 & n2032 ;
  assign n23250 = ~x760 & n15072 ;
  assign n23251 = n23200 & ~n23250 ;
  assign n23252 = x38 & ~n23251 ;
  assign n23253 = ~x178 & x760 ;
  assign n23254 = ~n14936 & n23253 ;
  assign n23255 = ( ~x178 & x760 ) | ( ~x178 & n15063 ) | ( x760 & n15063 ) ;
  assign n23256 = ( x178 & x760 ) | ( x178 & ~n14933 ) | ( x760 & ~n14933 ) ;
  assign n23257 = n23255 | n23256 ;
  assign n23258 = ~n23254 & n23257 ;
  assign n23259 = x38 | n23258 ;
  assign n23260 = ~n23252 & n23259 ;
  assign n23261 = ~n2032 & n23260 ;
  assign n23262 = n23249 | n23261 ;
  assign n23263 = ~n15082 & n23262 ;
  assign n23264 = n15082 & n23191 ;
  assign n23265 = n23263 | n23264 ;
  assign n23266 = ~x785 & n23265 ;
  assign n23267 = ~n15088 & n23191 ;
  assign n23268 = x609 & n23263 ;
  assign n23269 = n23267 | n23268 ;
  assign n23270 = x1155 & n23269 ;
  assign n23271 = n15094 & n23191 ;
  assign n23272 = ~x609 & n23263 ;
  assign n23273 = n23271 | n23272 ;
  assign n23274 = ~x1155 & n23273 ;
  assign n23275 = n23270 | n23274 ;
  assign n23276 = x785 & n23275 ;
  assign n23277 = n23266 | n23276 ;
  assign n23278 = ~x781 & n23277 ;
  assign n23279 = ( x618 & x1154 ) | ( x618 & n23191 ) | ( x1154 & n23191 ) ;
  assign n23280 = ( ~x618 & x1154 ) | ( ~x618 & n23277 ) | ( x1154 & n23277 ) ;
  assign n23281 = n23279 & n23280 ;
  assign n23282 = ( x618 & x1154 ) | ( x618 & ~n23191 ) | ( x1154 & ~n23191 ) ;
  assign n23283 = ( x618 & ~x1154 ) | ( x618 & n23277 ) | ( ~x1154 & n23277 ) ;
  assign n23284 = ~n23282 & n23283 ;
  assign n23285 = n23281 | n23284 ;
  assign n23286 = x781 & n23285 ;
  assign n23287 = n23278 | n23286 ;
  assign n23288 = ~x789 & n23287 ;
  assign n23289 = ( x619 & x1159 ) | ( x619 & n23191 ) | ( x1159 & n23191 ) ;
  assign n23290 = ( ~x619 & x1159 ) | ( ~x619 & n23287 ) | ( x1159 & n23287 ) ;
  assign n23291 = n23289 & n23290 ;
  assign n23292 = ( x619 & x1159 ) | ( x619 & ~n23191 ) | ( x1159 & ~n23191 ) ;
  assign n23293 = ( x619 & ~x1159 ) | ( x619 & n23287 ) | ( ~x1159 & n23287 ) ;
  assign n23294 = ~n23292 & n23293 ;
  assign n23295 = n23291 | n23294 ;
  assign n23296 = x789 & n23295 ;
  assign n23297 = n23288 | n23296 ;
  assign n23298 = n16176 | n23297 ;
  assign n23299 = n16176 & ~n23191 ;
  assign n23300 = n23298 & ~n23299 ;
  assign n23301 = n15134 | n23300 ;
  assign n23302 = n15134 & ~n23191 ;
  assign n23303 = n23301 & ~n23302 ;
  assign n23304 = n15141 | n23303 ;
  assign n23305 = n15141 & ~n23191 ;
  assign n23306 = n23304 & ~n23305 ;
  assign n23307 = ( x644 & x715 ) | ( x644 & ~n23306 ) | ( x715 & ~n23306 ) ;
  assign n23308 = ( x644 & ~x715 ) | ( x644 & n23191 ) | ( ~x715 & n23191 ) ;
  assign n23309 = ~n23307 & n23308 ;
  assign n23310 = x1160 & ~n23309 ;
  assign n23311 = ~n23248 & n23310 ;
  assign n23312 = x644 & ~n23246 ;
  assign n23313 = x715 | n23312 ;
  assign n23314 = ( x644 & x715 ) | ( x644 & n23306 ) | ( x715 & n23306 ) ;
  assign n23315 = ( ~x644 & x715 ) | ( ~x644 & n23191 ) | ( x715 & n23191 ) ;
  assign n23316 = n23314 & n23315 ;
  assign n23317 = x1160 | n23316 ;
  assign n23318 = n23313 & ~n23317 ;
  assign n23319 = n23311 | n23318 ;
  assign n23320 = x790 & n23319 ;
  assign n23321 = n18621 & n23300 ;
  assign n23322 = ( x629 & n23232 ) | ( x629 & n23321 ) | ( n23232 & n23321 ) ;
  assign n23323 = ( ~x629 & n23229 ) | ( ~x629 & n23321 ) | ( n23229 & n23321 ) ;
  assign n23324 = n23322 | n23323 ;
  assign n23325 = x792 & n23324 ;
  assign n23326 = x648 & ~n23294 ;
  assign n23327 = ( x619 & x1159 ) | ( x619 & n23220 ) | ( x1159 & n23220 ) ;
  assign n23328 = x627 | n23281 ;
  assign n23329 = ( x618 & x1154 ) | ( x618 & ~n23217 ) | ( x1154 & ~n23217 ) ;
  assign n23330 = x660 | n23270 ;
  assign n23331 = ( x609 & x1155 ) | ( x609 & ~n23214 ) | ( x1155 & ~n23214 ) ;
  assign n23332 = x608 | n23208 ;
  assign n23333 = ( x625 & x1153 ) | ( x625 & ~n23262 ) | ( x1153 & ~n23262 ) ;
  assign n23334 = x688 & ~n23260 ;
  assign n23335 = ( x178 & ~x760 ) | ( x178 & n15797 ) | ( ~x760 & n15797 ) ;
  assign n23336 = ( x178 & x760 ) | ( x178 & n15872 ) | ( x760 & n15872 ) ;
  assign n23337 = n23335 & ~n23336 ;
  assign n23338 = x39 & ~n23337 ;
  assign n23339 = ( x178 & ~x760 ) | ( x178 & n15583 ) | ( ~x760 & n15583 ) ;
  assign n23340 = ( x178 & x760 ) | ( x178 & n15699 ) | ( x760 & n15699 ) ;
  assign n23341 = ~n23339 & n23340 ;
  assign n23342 = n23338 & ~n23341 ;
  assign n23343 = ( ~x178 & x760 ) | ( ~x178 & n15887 ) | ( x760 & n15887 ) ;
  assign n23344 = ( x178 & x760 ) | ( x178 & ~n15891 ) | ( x760 & ~n15891 ) ;
  assign n23345 = n23343 & n23344 ;
  assign n23346 = ( ~x178 & x760 ) | ( ~x178 & n15894 ) | ( x760 & n15894 ) ;
  assign n23347 = ( x178 & x760 ) | ( x178 & ~n15897 ) | ( x760 & ~n15897 ) ;
  assign n23348 = n23346 | n23347 ;
  assign n23349 = ~n23345 & n23348 ;
  assign n23350 = x39 | n23349 ;
  assign n23351 = ~x38 & n23350 ;
  assign n23352 = ~n23342 & n23351 ;
  assign n23353 = x760 | n15758 ;
  assign n23354 = n17573 & n23353 ;
  assign n23355 = x178 | n23354 ;
  assign n23356 = n15529 | n23019 ;
  assign n23357 = x178 & n23356 ;
  assign n23358 = ~n4810 & n23357 ;
  assign n23359 = x38 & ~n23358 ;
  assign n23360 = n23355 & n23359 ;
  assign n23361 = x688 | n23360 ;
  assign n23362 = n23352 | n23361 ;
  assign n23363 = ~n2032 & n23362 ;
  assign n23364 = ~n23334 & n23363 ;
  assign n23365 = n23249 | n23364 ;
  assign n23366 = ( x625 & ~x1153 ) | ( x625 & n23365 ) | ( ~x1153 & n23365 ) ;
  assign n23367 = ~n23333 & n23366 ;
  assign n23368 = n23332 | n23367 ;
  assign n23369 = x608 & ~n23211 ;
  assign n23370 = ( x625 & x1153 ) | ( x625 & n23262 ) | ( x1153 & n23262 ) ;
  assign n23371 = ( ~x625 & x1153 ) | ( ~x625 & n23365 ) | ( x1153 & n23365 ) ;
  assign n23372 = n23370 & n23371 ;
  assign n23373 = n23369 & ~n23372 ;
  assign n23374 = n23368 & ~n23373 ;
  assign n23375 = x778 & ~n23374 ;
  assign n23376 = x778 | n23365 ;
  assign n23377 = ~n23375 & n23376 ;
  assign n23378 = ( x609 & ~x1155 ) | ( x609 & n23377 ) | ( ~x1155 & n23377 ) ;
  assign n23379 = ~n23331 & n23378 ;
  assign n23380 = n23330 | n23379 ;
  assign n23381 = x660 & ~n23274 ;
  assign n23382 = ( x609 & x1155 ) | ( x609 & n23214 ) | ( x1155 & n23214 ) ;
  assign n23383 = ( ~x609 & x1155 ) | ( ~x609 & n23377 ) | ( x1155 & n23377 ) ;
  assign n23384 = n23382 & n23383 ;
  assign n23385 = n23381 & ~n23384 ;
  assign n23386 = n23380 & ~n23385 ;
  assign n23387 = x785 & ~n23386 ;
  assign n23388 = x785 | n23377 ;
  assign n23389 = ~n23387 & n23388 ;
  assign n23390 = ( x618 & ~x1154 ) | ( x618 & n23389 ) | ( ~x1154 & n23389 ) ;
  assign n23391 = ~n23329 & n23390 ;
  assign n23392 = n23328 | n23391 ;
  assign n23393 = x627 & ~n23284 ;
  assign n23394 = ( x618 & x1154 ) | ( x618 & n23217 ) | ( x1154 & n23217 ) ;
  assign n23395 = ( ~x618 & x1154 ) | ( ~x618 & n23389 ) | ( x1154 & n23389 ) ;
  assign n23396 = n23394 & n23395 ;
  assign n23397 = n23393 & ~n23396 ;
  assign n23398 = n23392 & ~n23397 ;
  assign n23399 = x781 & ~n23398 ;
  assign n23400 = x781 | n23389 ;
  assign n23401 = ~n23399 & n23400 ;
  assign n23402 = ( ~x619 & x1159 ) | ( ~x619 & n23401 ) | ( x1159 & n23401 ) ;
  assign n23403 = n23327 & n23402 ;
  assign n23404 = n23326 & ~n23403 ;
  assign n23405 = x648 | n23291 ;
  assign n23406 = ( x619 & x1159 ) | ( x619 & ~n23220 ) | ( x1159 & ~n23220 ) ;
  assign n23407 = ( x619 & ~x1159 ) | ( x619 & n23401 ) | ( ~x1159 & n23401 ) ;
  assign n23408 = ~n23406 & n23407 ;
  assign n23409 = n23405 | n23408 ;
  assign n23410 = x789 & n23409 ;
  assign n23411 = ~n23404 & n23410 ;
  assign n23412 = ~x789 & n23401 ;
  assign n23413 = n16177 | n23412 ;
  assign n23414 = n23411 | n23413 ;
  assign n23415 = n16115 & ~n23222 ;
  assign n23416 = ( x626 & ~n15419 ) | ( x626 & n23191 ) | ( ~n15419 & n23191 ) ;
  assign n23417 = ( x626 & n15419 ) | ( x626 & ~n23297 ) | ( n15419 & ~n23297 ) ;
  assign n23418 = ~n23416 & n23417 ;
  assign n23419 = n23415 | n23418 ;
  assign n23420 = ( x626 & n15418 ) | ( x626 & ~n23191 ) | ( n15418 & ~n23191 ) ;
  assign n23421 = ( x626 & ~n15418 ) | ( x626 & n23297 ) | ( ~n15418 & n23297 ) ;
  assign n23422 = n23420 & ~n23421 ;
  assign n23423 = n23419 | n23422 ;
  assign n23424 = x788 & n23423 ;
  assign n23425 = n18434 | n23424 ;
  assign n23426 = n23414 & ~n23425 ;
  assign n23427 = n23325 | n23426 ;
  assign n23428 = ~n18431 & n23427 ;
  assign n23429 = n18610 & n23303 ;
  assign n23430 = n15139 & n23243 ;
  assign n23431 = n15138 & n23239 ;
  assign n23432 = n23430 | n23431 ;
  assign n23433 = n23429 | n23432 ;
  assign n23434 = x787 & n23433 ;
  assign n23435 = n23428 | n23434 ;
  assign n23436 = ( x644 & ~x790 ) | ( x644 & n23310 ) | ( ~x790 & n23310 ) ;
  assign n23437 = ( x644 & x790 ) | ( x644 & n23317 ) | ( x790 & n23317 ) ;
  assign n23438 = ~n23436 & n23437 ;
  assign n23439 = n23435 | n23438 ;
  assign n23440 = ~n23320 & n23439 ;
  assign n23441 = ( ~x832 & n6785 ) | ( ~x832 & n23440 ) | ( n6785 & n23440 ) ;
  assign n23442 = ( ~x178 & x832 ) | ( ~x178 & n6785 ) | ( x832 & n6785 ) ;
  assign n23443 = n23441 & ~n23442 ;
  assign n23444 = n23190 | n23443 ;
  assign n23445 = x179 | n14834 ;
  assign n23446 = n15141 & n23445 ;
  assign n23447 = x179 & n2032 ;
  assign n23448 = ~x741 & n22415 ;
  assign n23449 = x179 & ~n23448 ;
  assign n23450 = x179 | x741 ;
  assign n23451 = n17415 | n23450 ;
  assign n23452 = n17421 & ~n23451 ;
  assign n23453 = n23449 | n23452 ;
  assign n23454 = n19643 | n23453 ;
  assign n23455 = ~n2032 & n23454 ;
  assign n23456 = n23447 | n23455 ;
  assign n23457 = ~n15082 & n23456 ;
  assign n23458 = n15082 & n23445 ;
  assign n23459 = n23457 | n23458 ;
  assign n23460 = ~x785 & n23459 ;
  assign n23461 = ~n15088 & n23445 ;
  assign n23462 = x609 & n23457 ;
  assign n23463 = n23461 | n23462 ;
  assign n23464 = x1155 & n23463 ;
  assign n23465 = n15094 & n23445 ;
  assign n23466 = ~x609 & n23457 ;
  assign n23467 = n23465 | n23466 ;
  assign n23468 = ~x1155 & n23467 ;
  assign n23469 = n23464 | n23468 ;
  assign n23470 = x785 & n23469 ;
  assign n23471 = n23460 | n23470 ;
  assign n23472 = ~x781 & n23471 ;
  assign n23473 = ( x618 & x1154 ) | ( x618 & n23445 ) | ( x1154 & n23445 ) ;
  assign n23474 = ( ~x618 & x1154 ) | ( ~x618 & n23471 ) | ( x1154 & n23471 ) ;
  assign n23475 = n23473 & n23474 ;
  assign n23476 = ( x618 & x1154 ) | ( x618 & ~n23445 ) | ( x1154 & ~n23445 ) ;
  assign n23477 = ( x618 & ~x1154 ) | ( x618 & n23471 ) | ( ~x1154 & n23471 ) ;
  assign n23478 = ~n23476 & n23477 ;
  assign n23479 = n23475 | n23478 ;
  assign n23480 = x781 & n23479 ;
  assign n23481 = n23472 | n23480 ;
  assign n23482 = ~x789 & n23481 ;
  assign n23483 = ( x619 & x1159 ) | ( x619 & n23445 ) | ( x1159 & n23445 ) ;
  assign n23484 = ( ~x619 & x1159 ) | ( ~x619 & n23481 ) | ( x1159 & n23481 ) ;
  assign n23485 = n23483 & n23484 ;
  assign n23486 = ( x619 & x1159 ) | ( x619 & ~n23445 ) | ( x1159 & ~n23445 ) ;
  assign n23487 = ( x619 & ~x1159 ) | ( x619 & n23481 ) | ( ~x1159 & n23481 ) ;
  assign n23488 = ~n23486 & n23487 ;
  assign n23489 = n23485 | n23488 ;
  assign n23490 = x789 & n23489 ;
  assign n23491 = n23482 | n23490 ;
  assign n23492 = n16176 | n23491 ;
  assign n23493 = n16176 & ~n23445 ;
  assign n23494 = n23492 & ~n23493 ;
  assign n23495 = n15134 | n23494 ;
  assign n23496 = n15134 & ~n23445 ;
  assign n23497 = n23495 & ~n23496 ;
  assign n23498 = ~n15141 & n23497 ;
  assign n23499 = n23446 | n23498 ;
  assign n23500 = ( x644 & x715 ) | ( x644 & n23499 ) | ( x715 & n23499 ) ;
  assign n23501 = ( ~x644 & x715 ) | ( ~x644 & n23445 ) | ( x715 & n23445 ) ;
  assign n23502 = n23500 & n23501 ;
  assign n23503 = x1160 | n23502 ;
  assign n23504 = n15414 & n23445 ;
  assign n23505 = x724 | n2032 ;
  assign n23506 = ~n23445 & n23505 ;
  assign n23507 = x179 | n16319 ;
  assign n23508 = x179 & n16323 ;
  assign n23509 = x38 | n23508 ;
  assign n23510 = ~n2032 & n23509 ;
  assign n23511 = n23507 & ~n23510 ;
  assign n23512 = x179 | n15070 ;
  assign n23513 = n15375 & n23512 ;
  assign n23514 = x724 | n23513 ;
  assign n23515 = n23511 | n23514 ;
  assign n23516 = ~n23506 & n23515 ;
  assign n23517 = ~x778 & n23516 ;
  assign n23518 = ( x625 & x1153 ) | ( x625 & n23445 ) | ( x1153 & n23445 ) ;
  assign n23519 = ( ~x625 & x1153 ) | ( ~x625 & n23516 ) | ( x1153 & n23516 ) ;
  assign n23520 = n23518 & n23519 ;
  assign n23521 = ( x625 & x1153 ) | ( x625 & ~n23445 ) | ( x1153 & ~n23445 ) ;
  assign n23522 = ( x625 & ~x1153 ) | ( x625 & n23516 ) | ( ~x1153 & n23516 ) ;
  assign n23523 = ~n23521 & n23522 ;
  assign n23524 = n23520 | n23523 ;
  assign n23525 = x778 & n23524 ;
  assign n23526 = n23517 | n23525 ;
  assign n23527 = ~n15400 & n23526 ;
  assign n23528 = n15400 & n23445 ;
  assign n23529 = n23527 | n23528 ;
  assign n23530 = n15407 | n23529 ;
  assign n23531 = n15407 & ~n23445 ;
  assign n23532 = n23530 & ~n23531 ;
  assign n23533 = ~n15414 & n23532 ;
  assign n23534 = n23504 | n23533 ;
  assign n23535 = n15421 | n23534 ;
  assign n23536 = n15421 & ~n23445 ;
  assign n23537 = n23535 & ~n23536 ;
  assign n23538 = ~x792 & n23537 ;
  assign n23539 = ( x628 & x1156 ) | ( x628 & n23445 ) | ( x1156 & n23445 ) ;
  assign n23540 = ( ~x628 & x1156 ) | ( ~x628 & n23537 ) | ( x1156 & n23537 ) ;
  assign n23541 = n23539 & n23540 ;
  assign n23542 = ( x628 & x1156 ) | ( x628 & ~n23445 ) | ( x1156 & ~n23445 ) ;
  assign n23543 = ( x628 & ~x1156 ) | ( x628 & n23537 ) | ( ~x1156 & n23537 ) ;
  assign n23544 = ~n23542 & n23543 ;
  assign n23545 = n23541 | n23544 ;
  assign n23546 = x792 & n23545 ;
  assign n23547 = n23538 | n23546 ;
  assign n23548 = ~x787 & n23547 ;
  assign n23549 = ( x647 & x1157 ) | ( x647 & n23445 ) | ( x1157 & n23445 ) ;
  assign n23550 = ( ~x647 & x1157 ) | ( ~x647 & n23547 ) | ( x1157 & n23547 ) ;
  assign n23551 = n23549 & n23550 ;
  assign n23552 = ( x647 & x1157 ) | ( x647 & ~n23445 ) | ( x1157 & ~n23445 ) ;
  assign n23553 = ( x647 & ~x1157 ) | ( x647 & n23547 ) | ( ~x1157 & n23547 ) ;
  assign n23554 = ~n23552 & n23553 ;
  assign n23555 = n23551 | n23554 ;
  assign n23556 = x787 & n23555 ;
  assign n23557 = n23548 | n23556 ;
  assign n23558 = ( x644 & x715 ) | ( x644 & ~n23557 ) | ( x715 & ~n23557 ) ;
  assign n23559 = x630 | n23551 ;
  assign n23560 = ( x647 & x1157 ) | ( x647 & ~n23497 ) | ( x1157 & ~n23497 ) ;
  assign n23561 = x629 | n23541 ;
  assign n23562 = ( x628 & x1156 ) | ( x628 & ~n23494 ) | ( x1156 & ~n23494 ) ;
  assign n23563 = x648 | n23485 ;
  assign n23564 = ( x619 & x1159 ) | ( x619 & ~n23532 ) | ( x1159 & ~n23532 ) ;
  assign n23565 = x627 | n23475 ;
  assign n23566 = ( x618 & x1154 ) | ( x618 & ~n23529 ) | ( x1154 & ~n23529 ) ;
  assign n23567 = x660 | n23464 ;
  assign n23568 = ( x609 & x1155 ) | ( x609 & ~n23526 ) | ( x1155 & ~n23526 ) ;
  assign n23569 = x608 | n23520 ;
  assign n23570 = ( x625 & x1153 ) | ( x625 & ~n23456 ) | ( x1153 & ~n23456 ) ;
  assign n23571 = n16404 & n23512 ;
  assign n23572 = ( x39 & x179 ) | ( x39 & n15699 ) | ( x179 & n15699 ) ;
  assign n23573 = ( ~x39 & x179 ) | ( ~x39 & n15583 ) | ( x179 & n15583 ) ;
  assign n23574 = n23572 & ~n23573 ;
  assign n23575 = ( ~x39 & x179 ) | ( ~x39 & n15891 ) | ( x179 & n15891 ) ;
  assign n23576 = ( x39 & x179 ) | ( x39 & n15887 ) | ( x179 & n15887 ) ;
  assign n23577 = n23575 & ~n23576 ;
  assign n23578 = n23574 | n23577 ;
  assign n23579 = ~x38 & n23578 ;
  assign n23580 = n23571 | n23579 ;
  assign n23581 = x741 & n23580 ;
  assign n23582 = ( x179 & ~x741 ) | ( x179 & n17554 ) | ( ~x741 & n17554 ) ;
  assign n23583 = ( x179 & x741 ) | ( x179 & n17562 ) | ( x741 & n17562 ) ;
  assign n23584 = n23582 & ~n23583 ;
  assign n23585 = x724 | n23584 ;
  assign n23586 = n23581 | n23585 ;
  assign n23587 = x724 & ~n23454 ;
  assign n23588 = n2032 | n23587 ;
  assign n23589 = n23586 & ~n23588 ;
  assign n23590 = n23447 | n23589 ;
  assign n23591 = ( x625 & ~x1153 ) | ( x625 & n23590 ) | ( ~x1153 & n23590 ) ;
  assign n23592 = ~n23570 & n23591 ;
  assign n23593 = n23569 | n23592 ;
  assign n23594 = x608 & ~n23523 ;
  assign n23595 = ( x625 & x1153 ) | ( x625 & n23456 ) | ( x1153 & n23456 ) ;
  assign n23596 = ( ~x625 & x1153 ) | ( ~x625 & n23590 ) | ( x1153 & n23590 ) ;
  assign n23597 = n23595 & n23596 ;
  assign n23598 = n23594 & ~n23597 ;
  assign n23599 = n23593 & ~n23598 ;
  assign n23600 = x778 & ~n23599 ;
  assign n23601 = x778 | n23590 ;
  assign n23602 = ~n23600 & n23601 ;
  assign n23603 = ( x609 & ~x1155 ) | ( x609 & n23602 ) | ( ~x1155 & n23602 ) ;
  assign n23604 = ~n23568 & n23603 ;
  assign n23605 = n23567 | n23604 ;
  assign n23606 = x660 & ~n23468 ;
  assign n23607 = ( x609 & x1155 ) | ( x609 & n23526 ) | ( x1155 & n23526 ) ;
  assign n23608 = ( ~x609 & x1155 ) | ( ~x609 & n23602 ) | ( x1155 & n23602 ) ;
  assign n23609 = n23607 & n23608 ;
  assign n23610 = n23606 & ~n23609 ;
  assign n23611 = n23605 & ~n23610 ;
  assign n23612 = x785 & ~n23611 ;
  assign n23613 = x785 | n23602 ;
  assign n23614 = ~n23612 & n23613 ;
  assign n23615 = ( x618 & ~x1154 ) | ( x618 & n23614 ) | ( ~x1154 & n23614 ) ;
  assign n23616 = ~n23566 & n23615 ;
  assign n23617 = n23565 | n23616 ;
  assign n23618 = x627 & ~n23478 ;
  assign n23619 = ( x618 & x1154 ) | ( x618 & n23529 ) | ( x1154 & n23529 ) ;
  assign n23620 = ( ~x618 & x1154 ) | ( ~x618 & n23614 ) | ( x1154 & n23614 ) ;
  assign n23621 = n23619 & n23620 ;
  assign n23622 = n23618 & ~n23621 ;
  assign n23623 = n23617 & ~n23622 ;
  assign n23624 = x781 & ~n23623 ;
  assign n23625 = x781 | n23614 ;
  assign n23626 = ~n23624 & n23625 ;
  assign n23627 = ( x619 & ~x1159 ) | ( x619 & n23626 ) | ( ~x1159 & n23626 ) ;
  assign n23628 = ~n23564 & n23627 ;
  assign n23629 = n23563 | n23628 ;
  assign n23630 = x648 & ~n23488 ;
  assign n23631 = ( x619 & x1159 ) | ( x619 & n23532 ) | ( x1159 & n23532 ) ;
  assign n23632 = ( ~x619 & x1159 ) | ( ~x619 & n23626 ) | ( x1159 & n23626 ) ;
  assign n23633 = n23631 & n23632 ;
  assign n23634 = n23630 & ~n23633 ;
  assign n23635 = n23629 & ~n23634 ;
  assign n23636 = x789 & ~n23635 ;
  assign n23637 = x789 | n23626 ;
  assign n23638 = ~n23636 & n23637 ;
  assign n23639 = ~x788 & n23638 ;
  assign n23640 = ( x626 & x641 ) | ( x626 & ~n23491 ) | ( x641 & ~n23491 ) ;
  assign n23641 = ( x626 & ~x641 ) | ( x626 & n23445 ) | ( ~x641 & n23445 ) ;
  assign n23642 = n23640 & ~n23641 ;
  assign n23643 = x1158 | n23642 ;
  assign n23644 = ( x626 & x641 ) | ( x626 & n23534 ) | ( x641 & n23534 ) ;
  assign n23645 = ( ~x626 & x641 ) | ( ~x626 & n23638 ) | ( x641 & n23638 ) ;
  assign n23646 = n23644 | n23645 ;
  assign n23647 = ~n23643 & n23646 ;
  assign n23648 = ( x626 & x641 ) | ( x626 & n23491 ) | ( x641 & n23491 ) ;
  assign n23649 = ( ~x626 & x641 ) | ( ~x626 & n23445 ) | ( x641 & n23445 ) ;
  assign n23650 = n23648 | n23649 ;
  assign n23651 = x1158 & n23650 ;
  assign n23652 = ( x626 & x641 ) | ( x626 & ~n23534 ) | ( x641 & ~n23534 ) ;
  assign n23653 = ( x626 & ~x641 ) | ( x626 & n23638 ) | ( ~x641 & n23638 ) ;
  assign n23654 = n23652 & ~n23653 ;
  assign n23655 = n23651 & ~n23654 ;
  assign n23656 = n23647 | n23655 ;
  assign n23657 = x788 & n23656 ;
  assign n23658 = n23639 | n23657 ;
  assign n23659 = ( x628 & ~x1156 ) | ( x628 & n23658 ) | ( ~x1156 & n23658 ) ;
  assign n23660 = ~n23562 & n23659 ;
  assign n23661 = n23561 | n23660 ;
  assign n23662 = x629 & ~n23544 ;
  assign n23663 = ( x628 & x1156 ) | ( x628 & n23494 ) | ( x1156 & n23494 ) ;
  assign n23664 = ( ~x628 & x1156 ) | ( ~x628 & n23658 ) | ( x1156 & n23658 ) ;
  assign n23665 = n23663 & n23664 ;
  assign n23666 = n23662 & ~n23665 ;
  assign n23667 = n23661 & ~n23666 ;
  assign n23668 = x792 & ~n23667 ;
  assign n23669 = x792 | n23658 ;
  assign n23670 = ~n23668 & n23669 ;
  assign n23671 = ( x647 & ~x1157 ) | ( x647 & n23670 ) | ( ~x1157 & n23670 ) ;
  assign n23672 = ~n23560 & n23671 ;
  assign n23673 = n23559 | n23672 ;
  assign n23674 = x630 & ~n23554 ;
  assign n23675 = ( x647 & x1157 ) | ( x647 & n23497 ) | ( x1157 & n23497 ) ;
  assign n23676 = ( ~x647 & x1157 ) | ( ~x647 & n23670 ) | ( x1157 & n23670 ) ;
  assign n23677 = n23675 & n23676 ;
  assign n23678 = n23674 & ~n23677 ;
  assign n23679 = n23673 & ~n23678 ;
  assign n23680 = x787 & ~n23679 ;
  assign n23681 = x787 | n23670 ;
  assign n23682 = ~n23680 & n23681 ;
  assign n23683 = ( x644 & ~x715 ) | ( x644 & n23682 ) | ( ~x715 & n23682 ) ;
  assign n23684 = ~n23558 & n23683 ;
  assign n23685 = n23503 | n23684 ;
  assign n23686 = ( x644 & x715 ) | ( x644 & ~n23499 ) | ( x715 & ~n23499 ) ;
  assign n23687 = ( x644 & ~x715 ) | ( x644 & n23445 ) | ( ~x715 & n23445 ) ;
  assign n23688 = ~n23686 & n23687 ;
  assign n23689 = x1160 & ~n23688 ;
  assign n23690 = ( x644 & x715 ) | ( x644 & n23557 ) | ( x715 & n23557 ) ;
  assign n23691 = ( ~x644 & x715 ) | ( ~x644 & n23682 ) | ( x715 & n23682 ) ;
  assign n23692 = n23690 & n23691 ;
  assign n23693 = n23689 & ~n23692 ;
  assign n23694 = x790 & ~n23693 ;
  assign n23695 = n23685 & n23694 ;
  assign n23696 = ~x790 & n23682 ;
  assign n23697 = n6785 | n23696 ;
  assign n23698 = n23695 | n23697 ;
  assign n23699 = ~x179 & n6785 ;
  assign n23700 = x832 | n23699 ;
  assign n23701 = n23698 & ~n23700 ;
  assign n23702 = x179 | n1290 ;
  assign n23703 = ~x741 & n14840 ;
  assign n23704 = n23702 & ~n23703 ;
  assign n23705 = n16060 | n23704 ;
  assign n23706 = ~x785 & n23705 ;
  assign n23707 = n16065 | n23704 ;
  assign n23708 = x1155 & n23707 ;
  assign n23709 = n16068 | n23705 ;
  assign n23710 = ~x1155 & n23709 ;
  assign n23711 = n23708 | n23710 ;
  assign n23712 = x785 & n23711 ;
  assign n23713 = n23706 | n23712 ;
  assign n23714 = ~x781 & n23713 ;
  assign n23715 = n16075 | n23713 ;
  assign n23716 = x1154 & n23715 ;
  assign n23717 = n16078 | n23713 ;
  assign n23718 = ~x1154 & n23717 ;
  assign n23719 = n23716 | n23718 ;
  assign n23720 = x781 & n23719 ;
  assign n23721 = n23714 | n23720 ;
  assign n23722 = ~x789 & n23721 ;
  assign n23723 = ( x619 & x1159 ) | ( x619 & n23702 ) | ( x1159 & n23702 ) ;
  assign n23724 = ( ~x619 & x1159 ) | ( ~x619 & n23721 ) | ( x1159 & n23721 ) ;
  assign n23725 = n23723 & n23724 ;
  assign n23726 = ( x619 & x1159 ) | ( x619 & ~n23702 ) | ( x1159 & ~n23702 ) ;
  assign n23727 = ( x619 & ~x1159 ) | ( x619 & n23721 ) | ( ~x1159 & n23721 ) ;
  assign n23728 = ~n23726 & n23727 ;
  assign n23729 = n23725 | n23728 ;
  assign n23730 = x789 & n23729 ;
  assign n23731 = n23722 | n23730 ;
  assign n23732 = n16176 | n23731 ;
  assign n23733 = n16176 & ~n23702 ;
  assign n23734 = n23732 & ~n23733 ;
  assign n23735 = n15134 | n23734 ;
  assign n23736 = n15134 & ~n23702 ;
  assign n23737 = n23735 & ~n23736 ;
  assign n23738 = n18610 & n23737 ;
  assign n23739 = ( x647 & x1157 ) | ( x647 & ~n23702 ) | ( x1157 & ~n23702 ) ;
  assign n23740 = ~x724 & n15202 ;
  assign n23741 = n23702 & ~n23740 ;
  assign n23742 = ~x778 & n23741 ;
  assign n23743 = ~x625 & n23740 ;
  assign n23744 = n23741 | n23743 ;
  assign n23745 = x1153 & n23744 ;
  assign n23746 = ~x1153 & n23702 ;
  assign n23747 = ~n23743 & n23746 ;
  assign n23748 = n23745 | n23747 ;
  assign n23749 = x778 & n23748 ;
  assign n23750 = n23742 | n23749 ;
  assign n23751 = n16043 | n23750 ;
  assign n23752 = n16045 | n23751 ;
  assign n23753 = n16047 | n23752 ;
  assign n23754 = n16049 | n23753 ;
  assign n23755 = n16055 | n23754 ;
  assign n23756 = ( x647 & ~x1157 ) | ( x647 & n23755 ) | ( ~x1157 & n23755 ) ;
  assign n23757 = ~n23739 & n23756 ;
  assign n23758 = x630 & n23757 ;
  assign n23759 = x647 & n23755 ;
  assign n23760 = ~x647 & n23702 ;
  assign n23761 = n23759 | n23760 ;
  assign n23762 = n15138 & n23761 ;
  assign n23763 = n23758 | n23762 ;
  assign n23764 = n23738 | n23763 ;
  assign n23765 = x787 & n23764 ;
  assign n23766 = n16115 & ~n23753 ;
  assign n23767 = ( x626 & ~n15419 ) | ( x626 & n23702 ) | ( ~n15419 & n23702 ) ;
  assign n23768 = ( x626 & n15419 ) | ( x626 & ~n23731 ) | ( n15419 & ~n23731 ) ;
  assign n23769 = ~n23767 & n23768 ;
  assign n23770 = n23766 | n23769 ;
  assign n23771 = ( x626 & n15418 ) | ( x626 & ~n23702 ) | ( n15418 & ~n23702 ) ;
  assign n23772 = ( x626 & ~n15418 ) | ( x626 & n23731 ) | ( ~n15418 & n23731 ) ;
  assign n23773 = n23771 & ~n23772 ;
  assign n23774 = n23770 | n23773 ;
  assign n23775 = x788 & n23774 ;
  assign n23776 = x648 & ~n23728 ;
  assign n23777 = ( x619 & x1159 ) | ( x619 & n23752 ) | ( x1159 & n23752 ) ;
  assign n23778 = x627 | n23716 ;
  assign n23779 = ( x618 & x1154 ) | ( x618 & ~n23751 ) | ( x1154 & ~n23751 ) ;
  assign n23780 = x660 | n23708 ;
  assign n23781 = ( x609 & x1155 ) | ( x609 & ~n23750 ) | ( x1155 & ~n23750 ) ;
  assign n23782 = n14839 | n23741 ;
  assign n23783 = x625 & ~n23782 ;
  assign n23784 = n23704 & n23782 ;
  assign n23785 = n23783 | n23784 ;
  assign n23786 = n23746 & n23785 ;
  assign n23787 = x608 | n23745 ;
  assign n23788 = n23786 | n23787 ;
  assign n23789 = x1153 & n23704 ;
  assign n23790 = ~n23783 & n23789 ;
  assign n23791 = x608 & ~n23747 ;
  assign n23792 = ~n23790 & n23791 ;
  assign n23793 = n23788 & ~n23792 ;
  assign n23794 = x778 & ~n23793 ;
  assign n23795 = x778 | n23784 ;
  assign n23796 = ~n23794 & n23795 ;
  assign n23797 = ( x609 & ~x1155 ) | ( x609 & n23796 ) | ( ~x1155 & n23796 ) ;
  assign n23798 = ~n23781 & n23797 ;
  assign n23799 = n23780 | n23798 ;
  assign n23800 = x660 & ~n23710 ;
  assign n23801 = ( x609 & x1155 ) | ( x609 & n23750 ) | ( x1155 & n23750 ) ;
  assign n23802 = ( ~x609 & x1155 ) | ( ~x609 & n23796 ) | ( x1155 & n23796 ) ;
  assign n23803 = n23801 & n23802 ;
  assign n23804 = n23800 & ~n23803 ;
  assign n23805 = n23799 & ~n23804 ;
  assign n23806 = x785 & ~n23805 ;
  assign n23807 = x785 | n23796 ;
  assign n23808 = ~n23806 & n23807 ;
  assign n23809 = ( x618 & ~x1154 ) | ( x618 & n23808 ) | ( ~x1154 & n23808 ) ;
  assign n23810 = ~n23779 & n23809 ;
  assign n23811 = n23778 | n23810 ;
  assign n23812 = x627 & ~n23718 ;
  assign n23813 = ( x618 & x1154 ) | ( x618 & n23751 ) | ( x1154 & n23751 ) ;
  assign n23814 = ( ~x618 & x1154 ) | ( ~x618 & n23808 ) | ( x1154 & n23808 ) ;
  assign n23815 = n23813 & n23814 ;
  assign n23816 = n23812 & ~n23815 ;
  assign n23817 = n23811 & ~n23816 ;
  assign n23818 = x781 & ~n23817 ;
  assign n23819 = x781 | n23808 ;
  assign n23820 = ~n23818 & n23819 ;
  assign n23821 = ( ~x619 & x1159 ) | ( ~x619 & n23820 ) | ( x1159 & n23820 ) ;
  assign n23822 = n23777 & n23821 ;
  assign n23823 = n23776 & ~n23822 ;
  assign n23824 = x648 | n23725 ;
  assign n23825 = ( x619 & x1159 ) | ( x619 & ~n23752 ) | ( x1159 & ~n23752 ) ;
  assign n23826 = ( x619 & ~x1159 ) | ( x619 & n23820 ) | ( ~x1159 & n23820 ) ;
  assign n23827 = ~n23825 & n23826 ;
  assign n23828 = n23824 | n23827 ;
  assign n23829 = x789 & n23828 ;
  assign n23830 = ~n23823 & n23829 ;
  assign n23831 = ~x789 & n23820 ;
  assign n23832 = n16177 | n23831 ;
  assign n23833 = n23830 | n23832 ;
  assign n23834 = ~n23775 & n23833 ;
  assign n23835 = n18434 | n23834 ;
  assign n23836 = n16650 | n23754 ;
  assign n23837 = n16051 & ~n23734 ;
  assign n23838 = n23836 & ~n23837 ;
  assign n23839 = ( x629 & ~x792 ) | ( x629 & n23838 ) | ( ~x792 & n23838 ) ;
  assign n23840 = n16052 & ~n23734 ;
  assign n23841 = n16643 & ~n23754 ;
  assign n23842 = n23840 | n23841 ;
  assign n23843 = ( x629 & x792 ) | ( x629 & n23842 ) | ( x792 & n23842 ) ;
  assign n23844 = ~n23839 & n23843 ;
  assign n23845 = n18431 | n23844 ;
  assign n23846 = n23835 & ~n23845 ;
  assign n23847 = n23765 | n23846 ;
  assign n23848 = ( x790 & x832 ) | ( x790 & n23847 ) | ( x832 & n23847 ) ;
  assign n23849 = n15141 | n23737 ;
  assign n23850 = n15141 & ~n23702 ;
  assign n23851 = n23849 & ~n23850 ;
  assign n23852 = ( x644 & x715 ) | ( x644 & ~n23851 ) | ( x715 & ~n23851 ) ;
  assign n23853 = ( x644 & ~x715 ) | ( x644 & n23702 ) | ( ~x715 & n23702 ) ;
  assign n23854 = ~n23852 & n23853 ;
  assign n23855 = x1160 & ~n23854 ;
  assign n23856 = ~x787 & n23755 ;
  assign n23857 = x1157 & n23761 ;
  assign n23858 = n23757 | n23857 ;
  assign n23859 = x787 & n23858 ;
  assign n23860 = n23856 | n23859 ;
  assign n23861 = ( x644 & x715 ) | ( x644 & n23860 ) | ( x715 & n23860 ) ;
  assign n23862 = ( ~x644 & x715 ) | ( ~x644 & n23847 ) | ( x715 & n23847 ) ;
  assign n23863 = n23861 & n23862 ;
  assign n23864 = n23855 & ~n23863 ;
  assign n23865 = ( x644 & x715 ) | ( x644 & n23851 ) | ( x715 & n23851 ) ;
  assign n23866 = ( ~x644 & x715 ) | ( ~x644 & n23702 ) | ( x715 & n23702 ) ;
  assign n23867 = n23865 & n23866 ;
  assign n23868 = x1160 | n23867 ;
  assign n23869 = ( x644 & x715 ) | ( x644 & ~n23860 ) | ( x715 & ~n23860 ) ;
  assign n23870 = ( x644 & ~x715 ) | ( x644 & n23847 ) | ( ~x715 & n23847 ) ;
  assign n23871 = ~n23869 & n23870 ;
  assign n23872 = n23868 | n23871 ;
  assign n23873 = ~n23864 & n23872 ;
  assign n23874 = ( ~x790 & x832 ) | ( ~x790 & n23873 ) | ( x832 & n23873 ) ;
  assign n23875 = n23848 & n23874 ;
  assign n23876 = n23701 | n23875 ;
  assign n23877 = x180 | n1290 ;
  assign n23878 = ~x753 & n14840 ;
  assign n23879 = n23877 & ~n23878 ;
  assign n23880 = n16060 | n23879 ;
  assign n23881 = ~x785 & n23880 ;
  assign n23882 = ~n15094 & n23878 ;
  assign n23883 = n23880 | n23882 ;
  assign n23884 = x1155 & n23883 ;
  assign n23885 = ~x1155 & n23877 ;
  assign n23886 = ~n23882 & n23885 ;
  assign n23887 = n23884 | n23886 ;
  assign n23888 = x785 & n23887 ;
  assign n23889 = n23881 | n23888 ;
  assign n23890 = ~x781 & n23889 ;
  assign n23891 = n16075 | n23889 ;
  assign n23892 = x1154 & n23891 ;
  assign n23893 = n16078 | n23889 ;
  assign n23894 = ~x1154 & n23893 ;
  assign n23895 = n23892 | n23894 ;
  assign n23896 = x781 & n23895 ;
  assign n23897 = n23890 | n23896 ;
  assign n23898 = ~x789 & n23897 ;
  assign n23899 = n20948 | n23897 ;
  assign n23900 = x1159 & n23899 ;
  assign n23901 = n20951 | n23897 ;
  assign n23902 = ~x1159 & n23901 ;
  assign n23903 = n23900 | n23902 ;
  assign n23904 = x789 & n23903 ;
  assign n23905 = n23898 | n23904 ;
  assign n23906 = n16176 | n23905 ;
  assign n23907 = n16176 & ~n23877 ;
  assign n23908 = n23906 & ~n23907 ;
  assign n23909 = n15134 | n23908 ;
  assign n23910 = n15134 & ~n23877 ;
  assign n23911 = n23909 & ~n23910 ;
  assign n23912 = n18610 & n23911 ;
  assign n23913 = ( x647 & x1157 ) | ( x647 & ~n23877 ) | ( x1157 & ~n23877 ) ;
  assign n23914 = ~x702 & n15202 ;
  assign n23915 = n23877 & ~n23914 ;
  assign n23916 = x778 | n23915 ;
  assign n23917 = ~x625 & n23914 ;
  assign n23918 = n23915 | n23917 ;
  assign n23919 = x1153 & n23918 ;
  assign n23920 = ~x1153 & n23877 ;
  assign n23921 = ~n23917 & n23920 ;
  assign n23922 = x778 & ~n23921 ;
  assign n23923 = ~n23919 & n23922 ;
  assign n23924 = n23916 & ~n23923 ;
  assign n23925 = n16043 | n23924 ;
  assign n23926 = n16045 | n23925 ;
  assign n23927 = n16047 | n23926 ;
  assign n23928 = n16049 | n23927 ;
  assign n23929 = n16055 | n23928 ;
  assign n23930 = ( x647 & ~x1157 ) | ( x647 & n23929 ) | ( ~x1157 & n23929 ) ;
  assign n23931 = ~n23913 & n23930 ;
  assign n23932 = x630 & n23931 ;
  assign n23933 = x647 & n23929 ;
  assign n23934 = ~x647 & n23877 ;
  assign n23935 = n23933 | n23934 ;
  assign n23936 = n15138 & n23935 ;
  assign n23937 = n23932 | n23936 ;
  assign n23938 = n23912 | n23937 ;
  assign n23939 = x787 & n23938 ;
  assign n23940 = n16115 & ~n23927 ;
  assign n23941 = ( x626 & ~n15419 ) | ( x626 & n23877 ) | ( ~n15419 & n23877 ) ;
  assign n23942 = ( x626 & n15419 ) | ( x626 & ~n23905 ) | ( n15419 & ~n23905 ) ;
  assign n23943 = ~n23941 & n23942 ;
  assign n23944 = n23940 | n23943 ;
  assign n23945 = ( x626 & n15418 ) | ( x626 & ~n23877 ) | ( n15418 & ~n23877 ) ;
  assign n23946 = ( x626 & ~n15418 ) | ( x626 & n23905 ) | ( ~n15418 & n23905 ) ;
  assign n23947 = n23945 & ~n23946 ;
  assign n23948 = n23944 | n23947 ;
  assign n23949 = x788 & n23948 ;
  assign n23950 = x648 & ~n23902 ;
  assign n23951 = ( x619 & x1159 ) | ( x619 & n23926 ) | ( x1159 & n23926 ) ;
  assign n23952 = x627 | n23892 ;
  assign n23953 = ( x618 & x1154 ) | ( x618 & ~n23925 ) | ( x1154 & ~n23925 ) ;
  assign n23954 = x660 | n23884 ;
  assign n23955 = ( x609 & x1155 ) | ( x609 & ~n23924 ) | ( x1155 & ~n23924 ) ;
  assign n23956 = n14839 | n23915 ;
  assign n23957 = x625 & ~n23956 ;
  assign n23958 = n23879 & n23956 ;
  assign n23959 = n23957 | n23958 ;
  assign n23960 = n23920 & n23959 ;
  assign n23961 = x608 | n23919 ;
  assign n23962 = n23960 | n23961 ;
  assign n23963 = x1153 & n23879 ;
  assign n23964 = ~n23957 & n23963 ;
  assign n23965 = x608 & ~n23921 ;
  assign n23966 = ~n23964 & n23965 ;
  assign n23967 = n23962 & ~n23966 ;
  assign n23968 = x778 & ~n23967 ;
  assign n23969 = x778 | n23958 ;
  assign n23970 = ~n23968 & n23969 ;
  assign n23971 = ( x609 & ~x1155 ) | ( x609 & n23970 ) | ( ~x1155 & n23970 ) ;
  assign n23972 = ~n23955 & n23971 ;
  assign n23973 = n23954 | n23972 ;
  assign n23974 = x660 & ~n23886 ;
  assign n23975 = ( x609 & x1155 ) | ( x609 & n23924 ) | ( x1155 & n23924 ) ;
  assign n23976 = ( ~x609 & x1155 ) | ( ~x609 & n23970 ) | ( x1155 & n23970 ) ;
  assign n23977 = n23975 & n23976 ;
  assign n23978 = n23974 & ~n23977 ;
  assign n23979 = n23973 & ~n23978 ;
  assign n23980 = x785 & ~n23979 ;
  assign n23981 = x785 | n23970 ;
  assign n23982 = ~n23980 & n23981 ;
  assign n23983 = ( x618 & ~x1154 ) | ( x618 & n23982 ) | ( ~x1154 & n23982 ) ;
  assign n23984 = ~n23953 & n23983 ;
  assign n23985 = n23952 | n23984 ;
  assign n23986 = x627 & ~n23894 ;
  assign n23987 = ( x618 & x1154 ) | ( x618 & n23925 ) | ( x1154 & n23925 ) ;
  assign n23988 = ( ~x618 & x1154 ) | ( ~x618 & n23982 ) | ( x1154 & n23982 ) ;
  assign n23989 = n23987 & n23988 ;
  assign n23990 = n23986 & ~n23989 ;
  assign n23991 = n23985 & ~n23990 ;
  assign n23992 = x781 & ~n23991 ;
  assign n23993 = x781 | n23982 ;
  assign n23994 = ~n23992 & n23993 ;
  assign n23995 = ( ~x619 & x1159 ) | ( ~x619 & n23994 ) | ( x1159 & n23994 ) ;
  assign n23996 = n23951 & n23995 ;
  assign n23997 = n23950 & ~n23996 ;
  assign n23998 = x648 | n23900 ;
  assign n23999 = ( x619 & x1159 ) | ( x619 & ~n23926 ) | ( x1159 & ~n23926 ) ;
  assign n24000 = ( x619 & ~x1159 ) | ( x619 & n23994 ) | ( ~x1159 & n23994 ) ;
  assign n24001 = ~n23999 & n24000 ;
  assign n24002 = n23998 | n24001 ;
  assign n24003 = x789 & n24002 ;
  assign n24004 = ~n23997 & n24003 ;
  assign n24005 = ~x789 & n23994 ;
  assign n24006 = n16177 | n24005 ;
  assign n24007 = n24004 | n24006 ;
  assign n24008 = ~n23949 & n24007 ;
  assign n24009 = n18434 | n24008 ;
  assign n24010 = n16650 | n23928 ;
  assign n24011 = n16051 & ~n23908 ;
  assign n24012 = n24010 & ~n24011 ;
  assign n24013 = ( x629 & ~x792 ) | ( x629 & n24012 ) | ( ~x792 & n24012 ) ;
  assign n24014 = n16052 & ~n23908 ;
  assign n24015 = n16643 & ~n23928 ;
  assign n24016 = n24014 | n24015 ;
  assign n24017 = ( x629 & x792 ) | ( x629 & n24016 ) | ( x792 & n24016 ) ;
  assign n24018 = ~n24013 & n24017 ;
  assign n24019 = n18431 | n24018 ;
  assign n24020 = n24009 & ~n24019 ;
  assign n24021 = n23939 | n24020 ;
  assign n24022 = ( x790 & x832 ) | ( x790 & n24021 ) | ( x832 & n24021 ) ;
  assign n24023 = n15141 | n23911 ;
  assign n24024 = n15141 & ~n23877 ;
  assign n24025 = n24023 & ~n24024 ;
  assign n24026 = ( x644 & x715 ) | ( x644 & ~n24025 ) | ( x715 & ~n24025 ) ;
  assign n24027 = ( x644 & ~x715 ) | ( x644 & n23877 ) | ( ~x715 & n23877 ) ;
  assign n24028 = ~n24026 & n24027 ;
  assign n24029 = x1160 & ~n24028 ;
  assign n24030 = ~x787 & n23929 ;
  assign n24031 = x1157 & n23935 ;
  assign n24032 = n23931 | n24031 ;
  assign n24033 = x787 & n24032 ;
  assign n24034 = n24030 | n24033 ;
  assign n24035 = ( x644 & x715 ) | ( x644 & n24034 ) | ( x715 & n24034 ) ;
  assign n24036 = ( ~x644 & x715 ) | ( ~x644 & n24021 ) | ( x715 & n24021 ) ;
  assign n24037 = n24035 & n24036 ;
  assign n24038 = n24029 & ~n24037 ;
  assign n24039 = ( x644 & x715 ) | ( x644 & n24025 ) | ( x715 & n24025 ) ;
  assign n24040 = ( ~x644 & x715 ) | ( ~x644 & n23877 ) | ( x715 & n23877 ) ;
  assign n24041 = n24039 & n24040 ;
  assign n24042 = x1160 | n24041 ;
  assign n24043 = ( x644 & x715 ) | ( x644 & ~n24034 ) | ( x715 & ~n24034 ) ;
  assign n24044 = ( x644 & ~x715 ) | ( x644 & n24021 ) | ( ~x715 & n24021 ) ;
  assign n24045 = ~n24043 & n24044 ;
  assign n24046 = n24042 | n24045 ;
  assign n24047 = ~n24038 & n24046 ;
  assign n24048 = ( ~x790 & x832 ) | ( ~x790 & n24047 ) | ( x832 & n24047 ) ;
  assign n24049 = n24022 & n24048 ;
  assign n24050 = x180 | n14834 ;
  assign n24051 = n15414 & n24050 ;
  assign n24052 = x702 | n2032 ;
  assign n24053 = ~n24050 & n24052 ;
  assign n24054 = x180 & n16323 ;
  assign n24055 = x38 | n24054 ;
  assign n24056 = ~n2032 & n24055 ;
  assign n24057 = x180 | n16319 ;
  assign n24058 = ~n24056 & n24057 ;
  assign n24059 = x180 | n15070 ;
  assign n24060 = n15375 & n24059 ;
  assign n24061 = x702 | n24060 ;
  assign n24062 = n24058 | n24061 ;
  assign n24063 = ~n24053 & n24062 ;
  assign n24064 = ~x778 & n24063 ;
  assign n24065 = ( x625 & x1153 ) | ( x625 & n24050 ) | ( x1153 & n24050 ) ;
  assign n24066 = ( ~x625 & x1153 ) | ( ~x625 & n24063 ) | ( x1153 & n24063 ) ;
  assign n24067 = n24065 & n24066 ;
  assign n24068 = ( x625 & x1153 ) | ( x625 & ~n24050 ) | ( x1153 & ~n24050 ) ;
  assign n24069 = ( x625 & ~x1153 ) | ( x625 & n24063 ) | ( ~x1153 & n24063 ) ;
  assign n24070 = ~n24068 & n24069 ;
  assign n24071 = n24067 | n24070 ;
  assign n24072 = x778 & n24071 ;
  assign n24073 = n24064 | n24072 ;
  assign n24074 = ~n15400 & n24073 ;
  assign n24075 = n15400 & n24050 ;
  assign n24076 = n24074 | n24075 ;
  assign n24077 = n15407 | n24076 ;
  assign n24078 = n15407 & ~n24050 ;
  assign n24079 = n24077 & ~n24078 ;
  assign n24080 = ~n15414 & n24079 ;
  assign n24081 = n24051 | n24080 ;
  assign n24082 = n15421 | n24081 ;
  assign n24083 = n15421 & ~n24050 ;
  assign n24084 = n24082 & ~n24083 ;
  assign n24085 = ~x792 & n24084 ;
  assign n24086 = ( x628 & x1156 ) | ( x628 & n24050 ) | ( x1156 & n24050 ) ;
  assign n24087 = ( ~x628 & x1156 ) | ( ~x628 & n24084 ) | ( x1156 & n24084 ) ;
  assign n24088 = n24086 & n24087 ;
  assign n24089 = ( x628 & x1156 ) | ( x628 & ~n24050 ) | ( x1156 & ~n24050 ) ;
  assign n24090 = ( x628 & ~x1156 ) | ( x628 & n24084 ) | ( ~x1156 & n24084 ) ;
  assign n24091 = ~n24089 & n24090 ;
  assign n24092 = n24088 | n24091 ;
  assign n24093 = x792 & n24092 ;
  assign n24094 = n24085 | n24093 ;
  assign n24095 = x787 | n24094 ;
  assign n24096 = x647 & n24094 ;
  assign n24097 = ~x647 & n24050 ;
  assign n24098 = n24096 | n24097 ;
  assign n24099 = ( ~x787 & x1157 ) | ( ~x787 & n24098 ) | ( x1157 & n24098 ) ;
  assign n24100 = ~x647 & n24094 ;
  assign n24101 = x647 & n24050 ;
  assign n24102 = n24100 | n24101 ;
  assign n24103 = ( x787 & x1157 ) | ( x787 & ~n24102 ) | ( x1157 & ~n24102 ) ;
  assign n24104 = ~n24099 & n24103 ;
  assign n24105 = n24095 & ~n24104 ;
  assign n24106 = x644 | n24105 ;
  assign n24107 = x715 & n24106 ;
  assign n24108 = x180 & n2032 ;
  assign n24109 = x753 & n14710 ;
  assign n24110 = x180 & ~n14907 ;
  assign n24111 = n24109 | n24110 ;
  assign n24112 = x39 & n24111 ;
  assign n24113 = x180 & ~x753 ;
  assign n24114 = x180 & ~n15896 ;
  assign n24115 = n19729 | n24114 ;
  assign n24116 = ~x39 & n24115 ;
  assign n24117 = ( ~x753 & n15063 ) | ( ~x753 & n24113 ) | ( n15063 & n24113 ) ;
  assign n24118 = ( ~n24113 & n24116 ) | ( ~n24113 & n24117 ) | ( n24116 & n24117 ) ;
  assign n24119 = ( x180 & ~n24113 ) | ( x180 & n24118 ) | ( ~n24113 & n24118 ) ;
  assign n24120 = n24112 | n24119 ;
  assign n24121 = ~x38 & n24120 ;
  assign n24122 = ~x753 & n15072 ;
  assign n24123 = x38 & n24059 ;
  assign n24124 = ~n24122 & n24123 ;
  assign n24125 = n24121 | n24124 ;
  assign n24126 = ~n2032 & n24125 ;
  assign n24127 = n24108 | n24126 ;
  assign n24128 = ~n15082 & n24127 ;
  assign n24129 = n15082 & n24050 ;
  assign n24130 = n24128 | n24129 ;
  assign n24131 = ~x785 & n24130 ;
  assign n24132 = ~n15088 & n24050 ;
  assign n24133 = x609 & n24128 ;
  assign n24134 = n24132 | n24133 ;
  assign n24135 = x1155 & n24134 ;
  assign n24136 = n15094 & n24050 ;
  assign n24137 = ~x609 & n24128 ;
  assign n24138 = n24136 | n24137 ;
  assign n24139 = ~x1155 & n24138 ;
  assign n24140 = n24135 | n24139 ;
  assign n24141 = x785 & n24140 ;
  assign n24142 = n24131 | n24141 ;
  assign n24143 = ~x781 & n24142 ;
  assign n24144 = ( x618 & x1154 ) | ( x618 & n24050 ) | ( x1154 & n24050 ) ;
  assign n24145 = ( ~x618 & x1154 ) | ( ~x618 & n24142 ) | ( x1154 & n24142 ) ;
  assign n24146 = n24144 & n24145 ;
  assign n24147 = ( x618 & x1154 ) | ( x618 & ~n24050 ) | ( x1154 & ~n24050 ) ;
  assign n24148 = ( x618 & ~x1154 ) | ( x618 & n24142 ) | ( ~x1154 & n24142 ) ;
  assign n24149 = ~n24147 & n24148 ;
  assign n24150 = n24146 | n24149 ;
  assign n24151 = x781 & n24150 ;
  assign n24152 = n24143 | n24151 ;
  assign n24153 = ~x789 & n24152 ;
  assign n24154 = ( x619 & x1159 ) | ( x619 & n24050 ) | ( x1159 & n24050 ) ;
  assign n24155 = ( ~x619 & x1159 ) | ( ~x619 & n24152 ) | ( x1159 & n24152 ) ;
  assign n24156 = n24154 & n24155 ;
  assign n24157 = ( x619 & x1159 ) | ( x619 & ~n24050 ) | ( x1159 & ~n24050 ) ;
  assign n24158 = ( x619 & ~x1159 ) | ( x619 & n24152 ) | ( ~x1159 & n24152 ) ;
  assign n24159 = ~n24157 & n24158 ;
  assign n24160 = n24156 | n24159 ;
  assign n24161 = x789 & n24160 ;
  assign n24162 = n24153 | n24161 ;
  assign n24163 = n16176 | n24162 ;
  assign n24164 = n16176 & ~n24050 ;
  assign n24165 = n24163 & ~n24164 ;
  assign n24166 = n15134 | n24165 ;
  assign n24167 = n15134 & ~n24050 ;
  assign n24168 = n24166 & ~n24167 ;
  assign n24169 = n15141 | n24168 ;
  assign n24170 = n15141 & ~n24050 ;
  assign n24171 = n24169 & ~n24170 ;
  assign n24172 = ( x644 & x715 ) | ( x644 & ~n24171 ) | ( x715 & ~n24171 ) ;
  assign n24173 = ( x644 & ~x715 ) | ( x644 & n24050 ) | ( ~x715 & n24050 ) ;
  assign n24174 = ~n24172 & n24173 ;
  assign n24175 = x1160 & ~n24174 ;
  assign n24176 = ~n24107 & n24175 ;
  assign n24177 = x644 & ~n24105 ;
  assign n24178 = x715 | n24177 ;
  assign n24179 = ( x644 & x715 ) | ( x644 & n24171 ) | ( x715 & n24171 ) ;
  assign n24180 = ( ~x644 & x715 ) | ( ~x644 & n24050 ) | ( x715 & n24050 ) ;
  assign n24181 = n24179 & n24180 ;
  assign n24182 = x1160 | n24181 ;
  assign n24183 = n24178 & ~n24182 ;
  assign n24184 = n24176 | n24183 ;
  assign n24185 = x790 & n24184 ;
  assign n24186 = n18621 & n24165 ;
  assign n24187 = ( x629 & n24091 ) | ( x629 & n24186 ) | ( n24091 & n24186 ) ;
  assign n24188 = ( ~x629 & n24088 ) | ( ~x629 & n24186 ) | ( n24088 & n24186 ) ;
  assign n24189 = n24187 | n24188 ;
  assign n24190 = x792 & n24189 ;
  assign n24191 = x648 & ~n24159 ;
  assign n24192 = ( x619 & x1159 ) | ( x619 & n24079 ) | ( x1159 & n24079 ) ;
  assign n24193 = x627 | n24146 ;
  assign n24194 = ( x618 & x1154 ) | ( x618 & ~n24076 ) | ( x1154 & ~n24076 ) ;
  assign n24195 = x660 | n24135 ;
  assign n24196 = ( x609 & x1155 ) | ( x609 & ~n24073 ) | ( x1155 & ~n24073 ) ;
  assign n24197 = x608 | n24067 ;
  assign n24198 = ( x625 & x1153 ) | ( x625 & ~n24127 ) | ( x1153 & ~n24127 ) ;
  assign n24199 = x702 & ~n24125 ;
  assign n24200 = ( x180 & ~x753 ) | ( x180 & n15797 ) | ( ~x753 & n15797 ) ;
  assign n24201 = ( x180 & x753 ) | ( x180 & n15872 ) | ( x753 & n15872 ) ;
  assign n24202 = n24200 & ~n24201 ;
  assign n24203 = x39 & ~n24202 ;
  assign n24204 = ( x180 & ~x753 ) | ( x180 & n15583 ) | ( ~x753 & n15583 ) ;
  assign n24205 = ( x180 & x753 ) | ( x180 & n15699 ) | ( x753 & n15699 ) ;
  assign n24206 = ~n24204 & n24205 ;
  assign n24207 = n24203 & ~n24206 ;
  assign n24208 = ( ~x180 & x753 ) | ( ~x180 & n15887 ) | ( x753 & n15887 ) ;
  assign n24209 = ( x180 & x753 ) | ( x180 & ~n15891 ) | ( x753 & ~n15891 ) ;
  assign n24210 = n24208 & n24209 ;
  assign n24211 = ( ~x180 & x753 ) | ( ~x180 & n15894 ) | ( x753 & n15894 ) ;
  assign n24212 = ( x180 & x753 ) | ( x180 & ~n15897 ) | ( x753 & ~n15897 ) ;
  assign n24213 = n24211 | n24212 ;
  assign n24214 = ~n24210 & n24213 ;
  assign n24215 = x39 | n24214 ;
  assign n24216 = ~x38 & n24215 ;
  assign n24217 = ~n24207 & n24216 ;
  assign n24218 = x753 | n15758 ;
  assign n24219 = n17573 & n24218 ;
  assign n24220 = x180 | n24219 ;
  assign n24221 = n15529 | n23878 ;
  assign n24222 = x180 & n24221 ;
  assign n24223 = ~n4810 & n24222 ;
  assign n24224 = x38 & ~n24223 ;
  assign n24225 = n24220 & n24224 ;
  assign n24226 = x702 | n24225 ;
  assign n24227 = n24217 | n24226 ;
  assign n24228 = ~n2032 & n24227 ;
  assign n24229 = ~n24199 & n24228 ;
  assign n24230 = n24108 | n24229 ;
  assign n24231 = ( x625 & ~x1153 ) | ( x625 & n24230 ) | ( ~x1153 & n24230 ) ;
  assign n24232 = ~n24198 & n24231 ;
  assign n24233 = n24197 | n24232 ;
  assign n24234 = x608 & ~n24070 ;
  assign n24235 = ( x625 & x1153 ) | ( x625 & n24127 ) | ( x1153 & n24127 ) ;
  assign n24236 = ( ~x625 & x1153 ) | ( ~x625 & n24230 ) | ( x1153 & n24230 ) ;
  assign n24237 = n24235 & n24236 ;
  assign n24238 = n24234 & ~n24237 ;
  assign n24239 = n24233 & ~n24238 ;
  assign n24240 = x778 & ~n24239 ;
  assign n24241 = x778 | n24230 ;
  assign n24242 = ~n24240 & n24241 ;
  assign n24243 = ( x609 & ~x1155 ) | ( x609 & n24242 ) | ( ~x1155 & n24242 ) ;
  assign n24244 = ~n24196 & n24243 ;
  assign n24245 = n24195 | n24244 ;
  assign n24246 = x660 & ~n24139 ;
  assign n24247 = ( x609 & x1155 ) | ( x609 & n24073 ) | ( x1155 & n24073 ) ;
  assign n24248 = ( ~x609 & x1155 ) | ( ~x609 & n24242 ) | ( x1155 & n24242 ) ;
  assign n24249 = n24247 & n24248 ;
  assign n24250 = n24246 & ~n24249 ;
  assign n24251 = n24245 & ~n24250 ;
  assign n24252 = x785 & ~n24251 ;
  assign n24253 = x785 | n24242 ;
  assign n24254 = ~n24252 & n24253 ;
  assign n24255 = ( x618 & ~x1154 ) | ( x618 & n24254 ) | ( ~x1154 & n24254 ) ;
  assign n24256 = ~n24194 & n24255 ;
  assign n24257 = n24193 | n24256 ;
  assign n24258 = x627 & ~n24149 ;
  assign n24259 = ( x618 & x1154 ) | ( x618 & n24076 ) | ( x1154 & n24076 ) ;
  assign n24260 = ( ~x618 & x1154 ) | ( ~x618 & n24254 ) | ( x1154 & n24254 ) ;
  assign n24261 = n24259 & n24260 ;
  assign n24262 = n24258 & ~n24261 ;
  assign n24263 = n24257 & ~n24262 ;
  assign n24264 = x781 & ~n24263 ;
  assign n24265 = x781 | n24254 ;
  assign n24266 = ~n24264 & n24265 ;
  assign n24267 = ( ~x619 & x1159 ) | ( ~x619 & n24266 ) | ( x1159 & n24266 ) ;
  assign n24268 = n24192 & n24267 ;
  assign n24269 = n24191 & ~n24268 ;
  assign n24270 = x648 | n24156 ;
  assign n24271 = ( x619 & x1159 ) | ( x619 & ~n24079 ) | ( x1159 & ~n24079 ) ;
  assign n24272 = ( x619 & ~x1159 ) | ( x619 & n24266 ) | ( ~x1159 & n24266 ) ;
  assign n24273 = ~n24271 & n24272 ;
  assign n24274 = n24270 | n24273 ;
  assign n24275 = x789 & n24274 ;
  assign n24276 = ~n24269 & n24275 ;
  assign n24277 = ~x789 & n24266 ;
  assign n24278 = n16177 | n24277 ;
  assign n24279 = n24276 | n24278 ;
  assign n24280 = n16115 & ~n24081 ;
  assign n24281 = ( x626 & ~n15419 ) | ( x626 & n24050 ) | ( ~n15419 & n24050 ) ;
  assign n24282 = ( x626 & n15419 ) | ( x626 & ~n24162 ) | ( n15419 & ~n24162 ) ;
  assign n24283 = ~n24281 & n24282 ;
  assign n24284 = n24280 | n24283 ;
  assign n24285 = ( x626 & n15418 ) | ( x626 & ~n24050 ) | ( n15418 & ~n24050 ) ;
  assign n24286 = ( x626 & ~n15418 ) | ( x626 & n24162 ) | ( ~n15418 & n24162 ) ;
  assign n24287 = n24285 & ~n24286 ;
  assign n24288 = n24284 | n24287 ;
  assign n24289 = x788 & n24288 ;
  assign n24290 = n18434 | n24289 ;
  assign n24291 = n24279 & ~n24290 ;
  assign n24292 = n24190 | n24291 ;
  assign n24293 = ~n18431 & n24292 ;
  assign n24294 = n18610 & n24168 ;
  assign n24295 = n15139 & n24102 ;
  assign n24296 = n15138 & n24098 ;
  assign n24297 = n24295 | n24296 ;
  assign n24298 = n24294 | n24297 ;
  assign n24299 = x787 & n24298 ;
  assign n24300 = n24293 | n24299 ;
  assign n24301 = ( x644 & ~x790 ) | ( x644 & n24175 ) | ( ~x790 & n24175 ) ;
  assign n24302 = ( x644 & x790 ) | ( x644 & n24182 ) | ( x790 & n24182 ) ;
  assign n24303 = ~n24301 & n24302 ;
  assign n24304 = n24300 | n24303 ;
  assign n24305 = ~n24185 & n24304 ;
  assign n24306 = ( ~x832 & n6785 ) | ( ~x832 & n24305 ) | ( n6785 & n24305 ) ;
  assign n24307 = ( ~x180 & x832 ) | ( ~x180 & n6785 ) | ( x832 & n6785 ) ;
  assign n24308 = n24306 & ~n24307 ;
  assign n24309 = n24049 | n24308 ;
  assign n24310 = x181 | n1290 ;
  assign n24311 = ~x754 & n14840 ;
  assign n24312 = n24310 & ~n24311 ;
  assign n24313 = n16060 | n24312 ;
  assign n24314 = ~x785 & n24313 ;
  assign n24315 = ~n15094 & n24311 ;
  assign n24316 = n24313 | n24315 ;
  assign n24317 = x1155 & n24316 ;
  assign n24318 = ~x1155 & n24310 ;
  assign n24319 = ~n24315 & n24318 ;
  assign n24320 = n24317 | n24319 ;
  assign n24321 = x785 & n24320 ;
  assign n24322 = n24314 | n24321 ;
  assign n24323 = ~x781 & n24322 ;
  assign n24324 = n16075 | n24322 ;
  assign n24325 = x1154 & n24324 ;
  assign n24326 = n16078 | n24322 ;
  assign n24327 = ~x1154 & n24326 ;
  assign n24328 = n24325 | n24327 ;
  assign n24329 = x781 & n24328 ;
  assign n24330 = n24323 | n24329 ;
  assign n24331 = ~x789 & n24330 ;
  assign n24332 = n20948 | n24330 ;
  assign n24333 = x1159 & n24332 ;
  assign n24334 = n20951 | n24330 ;
  assign n24335 = ~x1159 & n24334 ;
  assign n24336 = n24333 | n24335 ;
  assign n24337 = x789 & n24336 ;
  assign n24338 = n24331 | n24337 ;
  assign n24339 = n16176 | n24338 ;
  assign n24340 = n16176 & ~n24310 ;
  assign n24341 = n24339 & ~n24340 ;
  assign n24342 = n15134 | n24341 ;
  assign n24343 = n15134 & ~n24310 ;
  assign n24344 = n24342 & ~n24343 ;
  assign n24345 = n18610 & n24344 ;
  assign n24346 = ( x647 & x1157 ) | ( x647 & ~n24310 ) | ( x1157 & ~n24310 ) ;
  assign n24347 = ~x709 & n15202 ;
  assign n24348 = n24310 & ~n24347 ;
  assign n24349 = x778 | n24348 ;
  assign n24350 = ~x625 & n24347 ;
  assign n24351 = n24348 | n24350 ;
  assign n24352 = x1153 & n24351 ;
  assign n24353 = ~x1153 & n24310 ;
  assign n24354 = ~n24350 & n24353 ;
  assign n24355 = x778 & ~n24354 ;
  assign n24356 = ~n24352 & n24355 ;
  assign n24357 = n24349 & ~n24356 ;
  assign n24358 = n16043 | n24357 ;
  assign n24359 = n16045 | n24358 ;
  assign n24360 = n16047 | n24359 ;
  assign n24361 = n16049 | n24360 ;
  assign n24362 = n16055 | n24361 ;
  assign n24363 = ( x647 & ~x1157 ) | ( x647 & n24362 ) | ( ~x1157 & n24362 ) ;
  assign n24364 = ~n24346 & n24363 ;
  assign n24365 = x630 & n24364 ;
  assign n24366 = x647 & n24362 ;
  assign n24367 = ~x647 & n24310 ;
  assign n24368 = n24366 | n24367 ;
  assign n24369 = n15138 & n24368 ;
  assign n24370 = n24365 | n24369 ;
  assign n24371 = n24345 | n24370 ;
  assign n24372 = x787 & n24371 ;
  assign n24373 = n16115 & ~n24360 ;
  assign n24374 = ( x626 & ~n15419 ) | ( x626 & n24310 ) | ( ~n15419 & n24310 ) ;
  assign n24375 = ( x626 & n15419 ) | ( x626 & ~n24338 ) | ( n15419 & ~n24338 ) ;
  assign n24376 = ~n24374 & n24375 ;
  assign n24377 = n24373 | n24376 ;
  assign n24378 = ( x626 & n15418 ) | ( x626 & ~n24310 ) | ( n15418 & ~n24310 ) ;
  assign n24379 = ( x626 & ~n15418 ) | ( x626 & n24338 ) | ( ~n15418 & n24338 ) ;
  assign n24380 = n24378 & ~n24379 ;
  assign n24381 = n24377 | n24380 ;
  assign n24382 = x788 & n24381 ;
  assign n24383 = x648 & ~n24335 ;
  assign n24384 = ( x619 & x1159 ) | ( x619 & n24359 ) | ( x1159 & n24359 ) ;
  assign n24385 = x627 | n24325 ;
  assign n24386 = ( x618 & x1154 ) | ( x618 & ~n24358 ) | ( x1154 & ~n24358 ) ;
  assign n24387 = x660 | n24317 ;
  assign n24388 = ( x609 & x1155 ) | ( x609 & ~n24357 ) | ( x1155 & ~n24357 ) ;
  assign n24389 = n14839 | n24348 ;
  assign n24390 = x625 & ~n24389 ;
  assign n24391 = n24312 & n24389 ;
  assign n24392 = n24390 | n24391 ;
  assign n24393 = n24353 & n24392 ;
  assign n24394 = x608 | n24352 ;
  assign n24395 = n24393 | n24394 ;
  assign n24396 = x1153 & n24312 ;
  assign n24397 = ~n24390 & n24396 ;
  assign n24398 = x608 & ~n24354 ;
  assign n24399 = ~n24397 & n24398 ;
  assign n24400 = n24395 & ~n24399 ;
  assign n24401 = x778 & ~n24400 ;
  assign n24402 = x778 | n24391 ;
  assign n24403 = ~n24401 & n24402 ;
  assign n24404 = ( x609 & ~x1155 ) | ( x609 & n24403 ) | ( ~x1155 & n24403 ) ;
  assign n24405 = ~n24388 & n24404 ;
  assign n24406 = n24387 | n24405 ;
  assign n24407 = x660 & ~n24319 ;
  assign n24408 = ( x609 & x1155 ) | ( x609 & n24357 ) | ( x1155 & n24357 ) ;
  assign n24409 = ( ~x609 & x1155 ) | ( ~x609 & n24403 ) | ( x1155 & n24403 ) ;
  assign n24410 = n24408 & n24409 ;
  assign n24411 = n24407 & ~n24410 ;
  assign n24412 = n24406 & ~n24411 ;
  assign n24413 = x785 & ~n24412 ;
  assign n24414 = x785 | n24403 ;
  assign n24415 = ~n24413 & n24414 ;
  assign n24416 = ( x618 & ~x1154 ) | ( x618 & n24415 ) | ( ~x1154 & n24415 ) ;
  assign n24417 = ~n24386 & n24416 ;
  assign n24418 = n24385 | n24417 ;
  assign n24419 = x627 & ~n24327 ;
  assign n24420 = ( x618 & x1154 ) | ( x618 & n24358 ) | ( x1154 & n24358 ) ;
  assign n24421 = ( ~x618 & x1154 ) | ( ~x618 & n24415 ) | ( x1154 & n24415 ) ;
  assign n24422 = n24420 & n24421 ;
  assign n24423 = n24419 & ~n24422 ;
  assign n24424 = n24418 & ~n24423 ;
  assign n24425 = x781 & ~n24424 ;
  assign n24426 = x781 | n24415 ;
  assign n24427 = ~n24425 & n24426 ;
  assign n24428 = ( ~x619 & x1159 ) | ( ~x619 & n24427 ) | ( x1159 & n24427 ) ;
  assign n24429 = n24384 & n24428 ;
  assign n24430 = n24383 & ~n24429 ;
  assign n24431 = x648 | n24333 ;
  assign n24432 = ( x619 & x1159 ) | ( x619 & ~n24359 ) | ( x1159 & ~n24359 ) ;
  assign n24433 = ( x619 & ~x1159 ) | ( x619 & n24427 ) | ( ~x1159 & n24427 ) ;
  assign n24434 = ~n24432 & n24433 ;
  assign n24435 = n24431 | n24434 ;
  assign n24436 = x789 & n24435 ;
  assign n24437 = ~n24430 & n24436 ;
  assign n24438 = ~x789 & n24427 ;
  assign n24439 = n16177 | n24438 ;
  assign n24440 = n24437 | n24439 ;
  assign n24441 = ~n24382 & n24440 ;
  assign n24442 = n18434 | n24441 ;
  assign n24443 = n16650 | n24361 ;
  assign n24444 = n16051 & ~n24341 ;
  assign n24445 = n24443 & ~n24444 ;
  assign n24446 = ( x629 & ~x792 ) | ( x629 & n24445 ) | ( ~x792 & n24445 ) ;
  assign n24447 = n16052 & ~n24341 ;
  assign n24448 = n16643 & ~n24361 ;
  assign n24449 = n24447 | n24448 ;
  assign n24450 = ( x629 & x792 ) | ( x629 & n24449 ) | ( x792 & n24449 ) ;
  assign n24451 = ~n24446 & n24450 ;
  assign n24452 = n18431 | n24451 ;
  assign n24453 = n24442 & ~n24452 ;
  assign n24454 = n24372 | n24453 ;
  assign n24455 = ( x790 & x832 ) | ( x790 & n24454 ) | ( x832 & n24454 ) ;
  assign n24456 = n15141 | n24344 ;
  assign n24457 = n15141 & ~n24310 ;
  assign n24458 = n24456 & ~n24457 ;
  assign n24459 = ( x644 & x715 ) | ( x644 & ~n24458 ) | ( x715 & ~n24458 ) ;
  assign n24460 = ( x644 & ~x715 ) | ( x644 & n24310 ) | ( ~x715 & n24310 ) ;
  assign n24461 = ~n24459 & n24460 ;
  assign n24462 = x1160 & ~n24461 ;
  assign n24463 = ~x787 & n24362 ;
  assign n24464 = x1157 & n24368 ;
  assign n24465 = n24364 | n24464 ;
  assign n24466 = x787 & n24465 ;
  assign n24467 = n24463 | n24466 ;
  assign n24468 = ( x644 & x715 ) | ( x644 & n24467 ) | ( x715 & n24467 ) ;
  assign n24469 = ( ~x644 & x715 ) | ( ~x644 & n24454 ) | ( x715 & n24454 ) ;
  assign n24470 = n24468 & n24469 ;
  assign n24471 = n24462 & ~n24470 ;
  assign n24472 = ( x644 & x715 ) | ( x644 & n24458 ) | ( x715 & n24458 ) ;
  assign n24473 = ( ~x644 & x715 ) | ( ~x644 & n24310 ) | ( x715 & n24310 ) ;
  assign n24474 = n24472 & n24473 ;
  assign n24475 = x1160 | n24474 ;
  assign n24476 = ( x644 & x715 ) | ( x644 & ~n24467 ) | ( x715 & ~n24467 ) ;
  assign n24477 = ( x644 & ~x715 ) | ( x644 & n24454 ) | ( ~x715 & n24454 ) ;
  assign n24478 = ~n24476 & n24477 ;
  assign n24479 = n24475 | n24478 ;
  assign n24480 = ~n24471 & n24479 ;
  assign n24481 = ( ~x790 & x832 ) | ( ~x790 & n24480 ) | ( x832 & n24480 ) ;
  assign n24482 = n24455 & n24481 ;
  assign n24483 = x181 | n14834 ;
  assign n24484 = n15414 & n24483 ;
  assign n24485 = x709 | n2032 ;
  assign n24486 = ~n24483 & n24485 ;
  assign n24487 = x181 & n16323 ;
  assign n24488 = x38 | n24487 ;
  assign n24489 = ~n2032 & n24488 ;
  assign n24490 = x181 | n16319 ;
  assign n24491 = ~n24489 & n24490 ;
  assign n24492 = x181 | n15070 ;
  assign n24493 = n15375 & n24492 ;
  assign n24494 = x709 | n24493 ;
  assign n24495 = n24491 | n24494 ;
  assign n24496 = ~n24486 & n24495 ;
  assign n24497 = ~x778 & n24496 ;
  assign n24498 = ( x625 & x1153 ) | ( x625 & n24483 ) | ( x1153 & n24483 ) ;
  assign n24499 = ( ~x625 & x1153 ) | ( ~x625 & n24496 ) | ( x1153 & n24496 ) ;
  assign n24500 = n24498 & n24499 ;
  assign n24501 = ( x625 & x1153 ) | ( x625 & ~n24483 ) | ( x1153 & ~n24483 ) ;
  assign n24502 = ( x625 & ~x1153 ) | ( x625 & n24496 ) | ( ~x1153 & n24496 ) ;
  assign n24503 = ~n24501 & n24502 ;
  assign n24504 = n24500 | n24503 ;
  assign n24505 = x778 & n24504 ;
  assign n24506 = n24497 | n24505 ;
  assign n24507 = ~n15400 & n24506 ;
  assign n24508 = n15400 & n24483 ;
  assign n24509 = n24507 | n24508 ;
  assign n24510 = n15407 | n24509 ;
  assign n24511 = n15407 & ~n24483 ;
  assign n24512 = n24510 & ~n24511 ;
  assign n24513 = ~n15414 & n24512 ;
  assign n24514 = n24484 | n24513 ;
  assign n24515 = n15421 | n24514 ;
  assign n24516 = n15421 & ~n24483 ;
  assign n24517 = n24515 & ~n24516 ;
  assign n24518 = ~x792 & n24517 ;
  assign n24519 = ( x628 & x1156 ) | ( x628 & n24483 ) | ( x1156 & n24483 ) ;
  assign n24520 = ( ~x628 & x1156 ) | ( ~x628 & n24517 ) | ( x1156 & n24517 ) ;
  assign n24521 = n24519 & n24520 ;
  assign n24522 = ( x628 & x1156 ) | ( x628 & ~n24483 ) | ( x1156 & ~n24483 ) ;
  assign n24523 = ( x628 & ~x1156 ) | ( x628 & n24517 ) | ( ~x1156 & n24517 ) ;
  assign n24524 = ~n24522 & n24523 ;
  assign n24525 = n24521 | n24524 ;
  assign n24526 = x792 & n24525 ;
  assign n24527 = n24518 | n24526 ;
  assign n24528 = x787 | n24527 ;
  assign n24529 = x647 & n24527 ;
  assign n24530 = ~x647 & n24483 ;
  assign n24531 = n24529 | n24530 ;
  assign n24532 = ( ~x787 & x1157 ) | ( ~x787 & n24531 ) | ( x1157 & n24531 ) ;
  assign n24533 = ~x647 & n24527 ;
  assign n24534 = x647 & n24483 ;
  assign n24535 = n24533 | n24534 ;
  assign n24536 = ( x787 & x1157 ) | ( x787 & ~n24535 ) | ( x1157 & ~n24535 ) ;
  assign n24537 = ~n24532 & n24536 ;
  assign n24538 = n24528 & ~n24537 ;
  assign n24539 = x644 | n24538 ;
  assign n24540 = x715 & n24539 ;
  assign n24541 = x181 & n2032 ;
  assign n24542 = x754 & n14710 ;
  assign n24543 = x181 & ~n14907 ;
  assign n24544 = n24542 | n24543 ;
  assign n24545 = x39 & n24544 ;
  assign n24546 = x181 & ~x754 ;
  assign n24547 = x181 & ~n15896 ;
  assign n24548 = n19779 | n24547 ;
  assign n24549 = ~x39 & n24548 ;
  assign n24550 = ( ~x754 & n15063 ) | ( ~x754 & n24546 ) | ( n15063 & n24546 ) ;
  assign n24551 = ( ~n24546 & n24549 ) | ( ~n24546 & n24550 ) | ( n24549 & n24550 ) ;
  assign n24552 = ( x181 & ~n24546 ) | ( x181 & n24551 ) | ( ~n24546 & n24551 ) ;
  assign n24553 = n24545 | n24552 ;
  assign n24554 = ~x38 & n24553 ;
  assign n24555 = ~x754 & n15072 ;
  assign n24556 = x38 & n24492 ;
  assign n24557 = ~n24555 & n24556 ;
  assign n24558 = n24554 | n24557 ;
  assign n24559 = ~n2032 & n24558 ;
  assign n24560 = n24541 | n24559 ;
  assign n24561 = ~n15082 & n24560 ;
  assign n24562 = n15082 & n24483 ;
  assign n24563 = n24561 | n24562 ;
  assign n24564 = ~x785 & n24563 ;
  assign n24565 = ~n15088 & n24483 ;
  assign n24566 = x609 & n24561 ;
  assign n24567 = n24565 | n24566 ;
  assign n24568 = x1155 & n24567 ;
  assign n24569 = n15094 & n24483 ;
  assign n24570 = ~x609 & n24561 ;
  assign n24571 = n24569 | n24570 ;
  assign n24572 = ~x1155 & n24571 ;
  assign n24573 = n24568 | n24572 ;
  assign n24574 = x785 & n24573 ;
  assign n24575 = n24564 | n24574 ;
  assign n24576 = ~x781 & n24575 ;
  assign n24577 = ( x618 & x1154 ) | ( x618 & n24483 ) | ( x1154 & n24483 ) ;
  assign n24578 = ( ~x618 & x1154 ) | ( ~x618 & n24575 ) | ( x1154 & n24575 ) ;
  assign n24579 = n24577 & n24578 ;
  assign n24580 = ( x618 & x1154 ) | ( x618 & ~n24483 ) | ( x1154 & ~n24483 ) ;
  assign n24581 = ( x618 & ~x1154 ) | ( x618 & n24575 ) | ( ~x1154 & n24575 ) ;
  assign n24582 = ~n24580 & n24581 ;
  assign n24583 = n24579 | n24582 ;
  assign n24584 = x781 & n24583 ;
  assign n24585 = n24576 | n24584 ;
  assign n24586 = ~x789 & n24585 ;
  assign n24587 = ( x619 & x1159 ) | ( x619 & n24483 ) | ( x1159 & n24483 ) ;
  assign n24588 = ( ~x619 & x1159 ) | ( ~x619 & n24585 ) | ( x1159 & n24585 ) ;
  assign n24589 = n24587 & n24588 ;
  assign n24590 = ( x619 & x1159 ) | ( x619 & ~n24483 ) | ( x1159 & ~n24483 ) ;
  assign n24591 = ( x619 & ~x1159 ) | ( x619 & n24585 ) | ( ~x1159 & n24585 ) ;
  assign n24592 = ~n24590 & n24591 ;
  assign n24593 = n24589 | n24592 ;
  assign n24594 = x789 & n24593 ;
  assign n24595 = n24586 | n24594 ;
  assign n24596 = n16176 | n24595 ;
  assign n24597 = n16176 & ~n24483 ;
  assign n24598 = n24596 & ~n24597 ;
  assign n24599 = n15134 | n24598 ;
  assign n24600 = n15134 & ~n24483 ;
  assign n24601 = n24599 & ~n24600 ;
  assign n24602 = n15141 | n24601 ;
  assign n24603 = n15141 & ~n24483 ;
  assign n24604 = n24602 & ~n24603 ;
  assign n24605 = ( x644 & x715 ) | ( x644 & ~n24604 ) | ( x715 & ~n24604 ) ;
  assign n24606 = ( x644 & ~x715 ) | ( x644 & n24483 ) | ( ~x715 & n24483 ) ;
  assign n24607 = ~n24605 & n24606 ;
  assign n24608 = x1160 & ~n24607 ;
  assign n24609 = ~n24540 & n24608 ;
  assign n24610 = x644 & ~n24538 ;
  assign n24611 = x715 | n24610 ;
  assign n24612 = ( x644 & x715 ) | ( x644 & n24604 ) | ( x715 & n24604 ) ;
  assign n24613 = ( ~x644 & x715 ) | ( ~x644 & n24483 ) | ( x715 & n24483 ) ;
  assign n24614 = n24612 & n24613 ;
  assign n24615 = x1160 | n24614 ;
  assign n24616 = n24611 & ~n24615 ;
  assign n24617 = n24609 | n24616 ;
  assign n24618 = x790 & n24617 ;
  assign n24619 = n18621 & n24598 ;
  assign n24620 = ( x629 & n24524 ) | ( x629 & n24619 ) | ( n24524 & n24619 ) ;
  assign n24621 = ( ~x629 & n24521 ) | ( ~x629 & n24619 ) | ( n24521 & n24619 ) ;
  assign n24622 = n24620 | n24621 ;
  assign n24623 = x792 & n24622 ;
  assign n24624 = x648 & ~n24592 ;
  assign n24625 = ( x619 & x1159 ) | ( x619 & n24512 ) | ( x1159 & n24512 ) ;
  assign n24626 = x627 | n24579 ;
  assign n24627 = ( x618 & x1154 ) | ( x618 & ~n24509 ) | ( x1154 & ~n24509 ) ;
  assign n24628 = x660 | n24568 ;
  assign n24629 = ( x609 & x1155 ) | ( x609 & ~n24506 ) | ( x1155 & ~n24506 ) ;
  assign n24630 = x608 | n24500 ;
  assign n24631 = ( x625 & x1153 ) | ( x625 & ~n24560 ) | ( x1153 & ~n24560 ) ;
  assign n24632 = x709 & ~n24558 ;
  assign n24633 = ( x181 & ~x754 ) | ( x181 & n15797 ) | ( ~x754 & n15797 ) ;
  assign n24634 = ( x181 & x754 ) | ( x181 & n15872 ) | ( x754 & n15872 ) ;
  assign n24635 = n24633 & ~n24634 ;
  assign n24636 = x39 & ~n24635 ;
  assign n24637 = ( x181 & ~x754 ) | ( x181 & n15583 ) | ( ~x754 & n15583 ) ;
  assign n24638 = ( x181 & x754 ) | ( x181 & n15699 ) | ( x754 & n15699 ) ;
  assign n24639 = ~n24637 & n24638 ;
  assign n24640 = n24636 & ~n24639 ;
  assign n24641 = ( ~x181 & x754 ) | ( ~x181 & n15887 ) | ( x754 & n15887 ) ;
  assign n24642 = ( x181 & x754 ) | ( x181 & ~n15891 ) | ( x754 & ~n15891 ) ;
  assign n24643 = n24641 & n24642 ;
  assign n24644 = ( ~x181 & x754 ) | ( ~x181 & n15894 ) | ( x754 & n15894 ) ;
  assign n24645 = ( x181 & x754 ) | ( x181 & ~n15897 ) | ( x754 & ~n15897 ) ;
  assign n24646 = n24644 | n24645 ;
  assign n24647 = ~n24643 & n24646 ;
  assign n24648 = x39 | n24647 ;
  assign n24649 = ~x38 & n24648 ;
  assign n24650 = ~n24640 & n24649 ;
  assign n24651 = x754 | n15758 ;
  assign n24652 = n17573 & n24651 ;
  assign n24653 = x181 | n24652 ;
  assign n24654 = n15529 | n24311 ;
  assign n24655 = x181 & n24654 ;
  assign n24656 = ~n4810 & n24655 ;
  assign n24657 = x38 & ~n24656 ;
  assign n24658 = n24653 & n24657 ;
  assign n24659 = x709 | n24658 ;
  assign n24660 = n24650 | n24659 ;
  assign n24661 = ~n2032 & n24660 ;
  assign n24662 = ~n24632 & n24661 ;
  assign n24663 = n24541 | n24662 ;
  assign n24664 = ( x625 & ~x1153 ) | ( x625 & n24663 ) | ( ~x1153 & n24663 ) ;
  assign n24665 = ~n24631 & n24664 ;
  assign n24666 = n24630 | n24665 ;
  assign n24667 = x608 & ~n24503 ;
  assign n24668 = ( x625 & x1153 ) | ( x625 & n24560 ) | ( x1153 & n24560 ) ;
  assign n24669 = ( ~x625 & x1153 ) | ( ~x625 & n24663 ) | ( x1153 & n24663 ) ;
  assign n24670 = n24668 & n24669 ;
  assign n24671 = n24667 & ~n24670 ;
  assign n24672 = n24666 & ~n24671 ;
  assign n24673 = x778 & ~n24672 ;
  assign n24674 = x778 | n24663 ;
  assign n24675 = ~n24673 & n24674 ;
  assign n24676 = ( x609 & ~x1155 ) | ( x609 & n24675 ) | ( ~x1155 & n24675 ) ;
  assign n24677 = ~n24629 & n24676 ;
  assign n24678 = n24628 | n24677 ;
  assign n24679 = x660 & ~n24572 ;
  assign n24680 = ( x609 & x1155 ) | ( x609 & n24506 ) | ( x1155 & n24506 ) ;
  assign n24681 = ( ~x609 & x1155 ) | ( ~x609 & n24675 ) | ( x1155 & n24675 ) ;
  assign n24682 = n24680 & n24681 ;
  assign n24683 = n24679 & ~n24682 ;
  assign n24684 = n24678 & ~n24683 ;
  assign n24685 = x785 & ~n24684 ;
  assign n24686 = x785 | n24675 ;
  assign n24687 = ~n24685 & n24686 ;
  assign n24688 = ( x618 & ~x1154 ) | ( x618 & n24687 ) | ( ~x1154 & n24687 ) ;
  assign n24689 = ~n24627 & n24688 ;
  assign n24690 = n24626 | n24689 ;
  assign n24691 = x627 & ~n24582 ;
  assign n24692 = ( x618 & x1154 ) | ( x618 & n24509 ) | ( x1154 & n24509 ) ;
  assign n24693 = ( ~x618 & x1154 ) | ( ~x618 & n24687 ) | ( x1154 & n24687 ) ;
  assign n24694 = n24692 & n24693 ;
  assign n24695 = n24691 & ~n24694 ;
  assign n24696 = n24690 & ~n24695 ;
  assign n24697 = x781 & ~n24696 ;
  assign n24698 = x781 | n24687 ;
  assign n24699 = ~n24697 & n24698 ;
  assign n24700 = ( ~x619 & x1159 ) | ( ~x619 & n24699 ) | ( x1159 & n24699 ) ;
  assign n24701 = n24625 & n24700 ;
  assign n24702 = n24624 & ~n24701 ;
  assign n24703 = x648 | n24589 ;
  assign n24704 = ( x619 & x1159 ) | ( x619 & ~n24512 ) | ( x1159 & ~n24512 ) ;
  assign n24705 = ( x619 & ~x1159 ) | ( x619 & n24699 ) | ( ~x1159 & n24699 ) ;
  assign n24706 = ~n24704 & n24705 ;
  assign n24707 = n24703 | n24706 ;
  assign n24708 = x789 & n24707 ;
  assign n24709 = ~n24702 & n24708 ;
  assign n24710 = ~x789 & n24699 ;
  assign n24711 = n16177 | n24710 ;
  assign n24712 = n24709 | n24711 ;
  assign n24713 = n16115 & ~n24514 ;
  assign n24714 = ( x626 & ~n15419 ) | ( x626 & n24483 ) | ( ~n15419 & n24483 ) ;
  assign n24715 = ( x626 & n15419 ) | ( x626 & ~n24595 ) | ( n15419 & ~n24595 ) ;
  assign n24716 = ~n24714 & n24715 ;
  assign n24717 = n24713 | n24716 ;
  assign n24718 = ( x626 & n15418 ) | ( x626 & ~n24483 ) | ( n15418 & ~n24483 ) ;
  assign n24719 = ( x626 & ~n15418 ) | ( x626 & n24595 ) | ( ~n15418 & n24595 ) ;
  assign n24720 = n24718 & ~n24719 ;
  assign n24721 = n24717 | n24720 ;
  assign n24722 = x788 & n24721 ;
  assign n24723 = n18434 | n24722 ;
  assign n24724 = n24712 & ~n24723 ;
  assign n24725 = n24623 | n24724 ;
  assign n24726 = ~n18431 & n24725 ;
  assign n24727 = n18610 & n24601 ;
  assign n24728 = n15139 & n24535 ;
  assign n24729 = n15138 & n24531 ;
  assign n24730 = n24728 | n24729 ;
  assign n24731 = n24727 | n24730 ;
  assign n24732 = x787 & n24731 ;
  assign n24733 = n24726 | n24732 ;
  assign n24734 = ( x644 & ~x790 ) | ( x644 & n24608 ) | ( ~x790 & n24608 ) ;
  assign n24735 = ( x644 & x790 ) | ( x644 & n24615 ) | ( x790 & n24615 ) ;
  assign n24736 = ~n24734 & n24735 ;
  assign n24737 = n24733 | n24736 ;
  assign n24738 = ~n24618 & n24737 ;
  assign n24739 = ( ~x832 & n6785 ) | ( ~x832 & n24738 ) | ( n6785 & n24738 ) ;
  assign n24740 = ( ~x181 & x832 ) | ( ~x181 & n6785 ) | ( x832 & n6785 ) ;
  assign n24741 = n24739 & ~n24740 ;
  assign n24742 = n24482 | n24741 ;
  assign n24743 = x182 | n1290 ;
  assign n24744 = ~x756 & n14840 ;
  assign n24745 = n24743 & ~n24744 ;
  assign n24746 = n16060 | n24745 ;
  assign n24747 = ~x785 & n24746 ;
  assign n24748 = ~n15094 & n24744 ;
  assign n24749 = n24746 | n24748 ;
  assign n24750 = x1155 & n24749 ;
  assign n24751 = ~x1155 & n24743 ;
  assign n24752 = ~n24748 & n24751 ;
  assign n24753 = n24750 | n24752 ;
  assign n24754 = x785 & n24753 ;
  assign n24755 = n24747 | n24754 ;
  assign n24756 = ~x781 & n24755 ;
  assign n24757 = n16075 | n24755 ;
  assign n24758 = x1154 & n24757 ;
  assign n24759 = n16078 | n24755 ;
  assign n24760 = ~x1154 & n24759 ;
  assign n24761 = n24758 | n24760 ;
  assign n24762 = x781 & n24761 ;
  assign n24763 = n24756 | n24762 ;
  assign n24764 = ~x789 & n24763 ;
  assign n24765 = n20948 | n24763 ;
  assign n24766 = x1159 & n24765 ;
  assign n24767 = n20951 | n24763 ;
  assign n24768 = ~x1159 & n24767 ;
  assign n24769 = n24766 | n24768 ;
  assign n24770 = x789 & n24769 ;
  assign n24771 = n24764 | n24770 ;
  assign n24772 = n16176 | n24771 ;
  assign n24773 = n16176 & ~n24743 ;
  assign n24774 = n24772 & ~n24773 ;
  assign n24775 = n15134 | n24774 ;
  assign n24776 = n15134 & ~n24743 ;
  assign n24777 = n24775 & ~n24776 ;
  assign n24778 = n18610 & n24777 ;
  assign n24779 = ( x647 & x1157 ) | ( x647 & ~n24743 ) | ( x1157 & ~n24743 ) ;
  assign n24780 = ~x734 & n15202 ;
  assign n24781 = n24743 & ~n24780 ;
  assign n24782 = x778 | n24781 ;
  assign n24783 = ~x625 & n24780 ;
  assign n24784 = n24781 | n24783 ;
  assign n24785 = x1153 & n24784 ;
  assign n24786 = ~x1153 & n24743 ;
  assign n24787 = ~n24783 & n24786 ;
  assign n24788 = x778 & ~n24787 ;
  assign n24789 = ~n24785 & n24788 ;
  assign n24790 = n24782 & ~n24789 ;
  assign n24791 = n16043 | n24790 ;
  assign n24792 = n16045 | n24791 ;
  assign n24793 = n16047 | n24792 ;
  assign n24794 = n16049 | n24793 ;
  assign n24795 = n16055 | n24794 ;
  assign n24796 = ( x647 & ~x1157 ) | ( x647 & n24795 ) | ( ~x1157 & n24795 ) ;
  assign n24797 = ~n24779 & n24796 ;
  assign n24798 = x630 & n24797 ;
  assign n24799 = x647 & n24795 ;
  assign n24800 = ~x647 & n24743 ;
  assign n24801 = n24799 | n24800 ;
  assign n24802 = n15138 & n24801 ;
  assign n24803 = n24798 | n24802 ;
  assign n24804 = n24778 | n24803 ;
  assign n24805 = x787 & n24804 ;
  assign n24806 = n16115 & ~n24793 ;
  assign n24807 = ( x626 & ~n15419 ) | ( x626 & n24743 ) | ( ~n15419 & n24743 ) ;
  assign n24808 = ( x626 & n15419 ) | ( x626 & ~n24771 ) | ( n15419 & ~n24771 ) ;
  assign n24809 = ~n24807 & n24808 ;
  assign n24810 = n24806 | n24809 ;
  assign n24811 = ( x626 & n15418 ) | ( x626 & ~n24743 ) | ( n15418 & ~n24743 ) ;
  assign n24812 = ( x626 & ~n15418 ) | ( x626 & n24771 ) | ( ~n15418 & n24771 ) ;
  assign n24813 = n24811 & ~n24812 ;
  assign n24814 = n24810 | n24813 ;
  assign n24815 = x788 & n24814 ;
  assign n24816 = x648 & ~n24768 ;
  assign n24817 = ( x619 & x1159 ) | ( x619 & n24792 ) | ( x1159 & n24792 ) ;
  assign n24818 = x627 | n24758 ;
  assign n24819 = ( x618 & x1154 ) | ( x618 & ~n24791 ) | ( x1154 & ~n24791 ) ;
  assign n24820 = x660 | n24750 ;
  assign n24821 = ( x609 & x1155 ) | ( x609 & ~n24790 ) | ( x1155 & ~n24790 ) ;
  assign n24822 = n14839 | n24781 ;
  assign n24823 = x625 & ~n24822 ;
  assign n24824 = n24745 & n24822 ;
  assign n24825 = n24823 | n24824 ;
  assign n24826 = n24786 & n24825 ;
  assign n24827 = x608 | n24785 ;
  assign n24828 = n24826 | n24827 ;
  assign n24829 = x1153 & n24745 ;
  assign n24830 = ~n24823 & n24829 ;
  assign n24831 = x608 & ~n24787 ;
  assign n24832 = ~n24830 & n24831 ;
  assign n24833 = n24828 & ~n24832 ;
  assign n24834 = x778 & ~n24833 ;
  assign n24835 = x778 | n24824 ;
  assign n24836 = ~n24834 & n24835 ;
  assign n24837 = ( x609 & ~x1155 ) | ( x609 & n24836 ) | ( ~x1155 & n24836 ) ;
  assign n24838 = ~n24821 & n24837 ;
  assign n24839 = n24820 | n24838 ;
  assign n24840 = x660 & ~n24752 ;
  assign n24841 = ( x609 & x1155 ) | ( x609 & n24790 ) | ( x1155 & n24790 ) ;
  assign n24842 = ( ~x609 & x1155 ) | ( ~x609 & n24836 ) | ( x1155 & n24836 ) ;
  assign n24843 = n24841 & n24842 ;
  assign n24844 = n24840 & ~n24843 ;
  assign n24845 = n24839 & ~n24844 ;
  assign n24846 = x785 & ~n24845 ;
  assign n24847 = x785 | n24836 ;
  assign n24848 = ~n24846 & n24847 ;
  assign n24849 = ( x618 & ~x1154 ) | ( x618 & n24848 ) | ( ~x1154 & n24848 ) ;
  assign n24850 = ~n24819 & n24849 ;
  assign n24851 = n24818 | n24850 ;
  assign n24852 = x627 & ~n24760 ;
  assign n24853 = ( x618 & x1154 ) | ( x618 & n24791 ) | ( x1154 & n24791 ) ;
  assign n24854 = ( ~x618 & x1154 ) | ( ~x618 & n24848 ) | ( x1154 & n24848 ) ;
  assign n24855 = n24853 & n24854 ;
  assign n24856 = n24852 & ~n24855 ;
  assign n24857 = n24851 & ~n24856 ;
  assign n24858 = x781 & ~n24857 ;
  assign n24859 = x781 | n24848 ;
  assign n24860 = ~n24858 & n24859 ;
  assign n24861 = ( ~x619 & x1159 ) | ( ~x619 & n24860 ) | ( x1159 & n24860 ) ;
  assign n24862 = n24817 & n24861 ;
  assign n24863 = n24816 & ~n24862 ;
  assign n24864 = x648 | n24766 ;
  assign n24865 = ( x619 & x1159 ) | ( x619 & ~n24792 ) | ( x1159 & ~n24792 ) ;
  assign n24866 = ( x619 & ~x1159 ) | ( x619 & n24860 ) | ( ~x1159 & n24860 ) ;
  assign n24867 = ~n24865 & n24866 ;
  assign n24868 = n24864 | n24867 ;
  assign n24869 = x789 & n24868 ;
  assign n24870 = ~n24863 & n24869 ;
  assign n24871 = ~x789 & n24860 ;
  assign n24872 = n16177 | n24871 ;
  assign n24873 = n24870 | n24872 ;
  assign n24874 = ~n24815 & n24873 ;
  assign n24875 = n18434 | n24874 ;
  assign n24876 = n16650 | n24794 ;
  assign n24877 = n16051 & ~n24774 ;
  assign n24878 = n24876 & ~n24877 ;
  assign n24879 = ( x629 & ~x792 ) | ( x629 & n24878 ) | ( ~x792 & n24878 ) ;
  assign n24880 = n16052 & ~n24774 ;
  assign n24881 = n16643 & ~n24794 ;
  assign n24882 = n24880 | n24881 ;
  assign n24883 = ( x629 & x792 ) | ( x629 & n24882 ) | ( x792 & n24882 ) ;
  assign n24884 = ~n24879 & n24883 ;
  assign n24885 = n18431 | n24884 ;
  assign n24886 = n24875 & ~n24885 ;
  assign n24887 = n24805 | n24886 ;
  assign n24888 = ( x790 & x832 ) | ( x790 & n24887 ) | ( x832 & n24887 ) ;
  assign n24889 = n15141 | n24777 ;
  assign n24890 = n15141 & ~n24743 ;
  assign n24891 = n24889 & ~n24890 ;
  assign n24892 = ( x644 & x715 ) | ( x644 & ~n24891 ) | ( x715 & ~n24891 ) ;
  assign n24893 = ( x644 & ~x715 ) | ( x644 & n24743 ) | ( ~x715 & n24743 ) ;
  assign n24894 = ~n24892 & n24893 ;
  assign n24895 = x1160 & ~n24894 ;
  assign n24896 = ~x787 & n24795 ;
  assign n24897 = x1157 & n24801 ;
  assign n24898 = n24797 | n24897 ;
  assign n24899 = x787 & n24898 ;
  assign n24900 = n24896 | n24899 ;
  assign n24901 = ( x644 & x715 ) | ( x644 & n24900 ) | ( x715 & n24900 ) ;
  assign n24902 = ( ~x644 & x715 ) | ( ~x644 & n24887 ) | ( x715 & n24887 ) ;
  assign n24903 = n24901 & n24902 ;
  assign n24904 = n24895 & ~n24903 ;
  assign n24905 = ( x644 & x715 ) | ( x644 & n24891 ) | ( x715 & n24891 ) ;
  assign n24906 = ( ~x644 & x715 ) | ( ~x644 & n24743 ) | ( x715 & n24743 ) ;
  assign n24907 = n24905 & n24906 ;
  assign n24908 = x1160 | n24907 ;
  assign n24909 = ( x644 & x715 ) | ( x644 & ~n24900 ) | ( x715 & ~n24900 ) ;
  assign n24910 = ( x644 & ~x715 ) | ( x644 & n24887 ) | ( ~x715 & n24887 ) ;
  assign n24911 = ~n24909 & n24910 ;
  assign n24912 = n24908 | n24911 ;
  assign n24913 = ~n24904 & n24912 ;
  assign n24914 = ( ~x790 & x832 ) | ( ~x790 & n24913 ) | ( x832 & n24913 ) ;
  assign n24915 = n24888 & n24914 ;
  assign n24916 = x182 | n14834 ;
  assign n24917 = n15414 & n24916 ;
  assign n24918 = x734 | n2032 ;
  assign n24919 = ~n24916 & n24918 ;
  assign n24920 = x182 & n16323 ;
  assign n24921 = x38 | n24920 ;
  assign n24922 = ~n2032 & n24921 ;
  assign n24923 = x182 | n16319 ;
  assign n24924 = ~n24922 & n24923 ;
  assign n24925 = x182 | n15070 ;
  assign n24926 = n15375 & n24925 ;
  assign n24927 = x734 | n24926 ;
  assign n24928 = n24924 | n24927 ;
  assign n24929 = ~n24919 & n24928 ;
  assign n24930 = ~x778 & n24929 ;
  assign n24931 = ( x625 & x1153 ) | ( x625 & n24916 ) | ( x1153 & n24916 ) ;
  assign n24932 = ( ~x625 & x1153 ) | ( ~x625 & n24929 ) | ( x1153 & n24929 ) ;
  assign n24933 = n24931 & n24932 ;
  assign n24934 = ( x625 & x1153 ) | ( x625 & ~n24916 ) | ( x1153 & ~n24916 ) ;
  assign n24935 = ( x625 & ~x1153 ) | ( x625 & n24929 ) | ( ~x1153 & n24929 ) ;
  assign n24936 = ~n24934 & n24935 ;
  assign n24937 = n24933 | n24936 ;
  assign n24938 = x778 & n24937 ;
  assign n24939 = n24930 | n24938 ;
  assign n24940 = ~n15400 & n24939 ;
  assign n24941 = n15400 & n24916 ;
  assign n24942 = n24940 | n24941 ;
  assign n24943 = n15407 | n24942 ;
  assign n24944 = n15407 & ~n24916 ;
  assign n24945 = n24943 & ~n24944 ;
  assign n24946 = ~n15414 & n24945 ;
  assign n24947 = n24917 | n24946 ;
  assign n24948 = n15421 | n24947 ;
  assign n24949 = n15421 & ~n24916 ;
  assign n24950 = n24948 & ~n24949 ;
  assign n24951 = ~x792 & n24950 ;
  assign n24952 = ( x628 & x1156 ) | ( x628 & n24916 ) | ( x1156 & n24916 ) ;
  assign n24953 = ( ~x628 & x1156 ) | ( ~x628 & n24950 ) | ( x1156 & n24950 ) ;
  assign n24954 = n24952 & n24953 ;
  assign n24955 = ( x628 & x1156 ) | ( x628 & ~n24916 ) | ( x1156 & ~n24916 ) ;
  assign n24956 = ( x628 & ~x1156 ) | ( x628 & n24950 ) | ( ~x1156 & n24950 ) ;
  assign n24957 = ~n24955 & n24956 ;
  assign n24958 = n24954 | n24957 ;
  assign n24959 = x792 & n24958 ;
  assign n24960 = n24951 | n24959 ;
  assign n24961 = x787 | n24960 ;
  assign n24962 = x647 & n24960 ;
  assign n24963 = ~x647 & n24916 ;
  assign n24964 = n24962 | n24963 ;
  assign n24965 = ( ~x787 & x1157 ) | ( ~x787 & n24964 ) | ( x1157 & n24964 ) ;
  assign n24966 = ~x647 & n24960 ;
  assign n24967 = x647 & n24916 ;
  assign n24968 = n24966 | n24967 ;
  assign n24969 = ( x787 & x1157 ) | ( x787 & ~n24968 ) | ( x1157 & ~n24968 ) ;
  assign n24970 = ~n24965 & n24969 ;
  assign n24971 = n24961 & ~n24970 ;
  assign n24972 = x644 | n24971 ;
  assign n24973 = x715 & n24972 ;
  assign n24974 = x182 & n2032 ;
  assign n24975 = ~x756 & n15072 ;
  assign n24976 = n24925 & ~n24975 ;
  assign n24977 = x38 & ~n24976 ;
  assign n24978 = ~x182 & x756 ;
  assign n24979 = ~n14936 & n24978 ;
  assign n24980 = ( ~x182 & x756 ) | ( ~x182 & n15063 ) | ( x756 & n15063 ) ;
  assign n24981 = ( x182 & x756 ) | ( x182 & ~n14933 ) | ( x756 & ~n14933 ) ;
  assign n24982 = n24980 | n24981 ;
  assign n24983 = ~n24979 & n24982 ;
  assign n24984 = x38 | n24983 ;
  assign n24985 = ~n24977 & n24984 ;
  assign n24986 = ~n2032 & n24985 ;
  assign n24987 = n24974 | n24986 ;
  assign n24988 = ~n15082 & n24987 ;
  assign n24989 = n15082 & n24916 ;
  assign n24990 = n24988 | n24989 ;
  assign n24991 = ~x785 & n24990 ;
  assign n24992 = ~n15088 & n24916 ;
  assign n24993 = x609 & n24988 ;
  assign n24994 = n24992 | n24993 ;
  assign n24995 = x1155 & n24994 ;
  assign n24996 = n15094 & n24916 ;
  assign n24997 = ~x609 & n24988 ;
  assign n24998 = n24996 | n24997 ;
  assign n24999 = ~x1155 & n24998 ;
  assign n25000 = n24995 | n24999 ;
  assign n25001 = x785 & n25000 ;
  assign n25002 = n24991 | n25001 ;
  assign n25003 = ~x781 & n25002 ;
  assign n25004 = ( x618 & x1154 ) | ( x618 & n24916 ) | ( x1154 & n24916 ) ;
  assign n25005 = ( ~x618 & x1154 ) | ( ~x618 & n25002 ) | ( x1154 & n25002 ) ;
  assign n25006 = n25004 & n25005 ;
  assign n25007 = ( x618 & x1154 ) | ( x618 & ~n24916 ) | ( x1154 & ~n24916 ) ;
  assign n25008 = ( x618 & ~x1154 ) | ( x618 & n25002 ) | ( ~x1154 & n25002 ) ;
  assign n25009 = ~n25007 & n25008 ;
  assign n25010 = n25006 | n25009 ;
  assign n25011 = x781 & n25010 ;
  assign n25012 = n25003 | n25011 ;
  assign n25013 = ~x789 & n25012 ;
  assign n25014 = ( x619 & x1159 ) | ( x619 & n24916 ) | ( x1159 & n24916 ) ;
  assign n25015 = ( ~x619 & x1159 ) | ( ~x619 & n25012 ) | ( x1159 & n25012 ) ;
  assign n25016 = n25014 & n25015 ;
  assign n25017 = ( x619 & x1159 ) | ( x619 & ~n24916 ) | ( x1159 & ~n24916 ) ;
  assign n25018 = ( x619 & ~x1159 ) | ( x619 & n25012 ) | ( ~x1159 & n25012 ) ;
  assign n25019 = ~n25017 & n25018 ;
  assign n25020 = n25016 | n25019 ;
  assign n25021 = x789 & n25020 ;
  assign n25022 = n25013 | n25021 ;
  assign n25023 = n16176 | n25022 ;
  assign n25024 = n16176 & ~n24916 ;
  assign n25025 = n25023 & ~n25024 ;
  assign n25026 = n15134 | n25025 ;
  assign n25027 = n15134 & ~n24916 ;
  assign n25028 = n25026 & ~n25027 ;
  assign n25029 = n15141 | n25028 ;
  assign n25030 = n15141 & ~n24916 ;
  assign n25031 = n25029 & ~n25030 ;
  assign n25032 = ( x644 & x715 ) | ( x644 & ~n25031 ) | ( x715 & ~n25031 ) ;
  assign n25033 = ( x644 & ~x715 ) | ( x644 & n24916 ) | ( ~x715 & n24916 ) ;
  assign n25034 = ~n25032 & n25033 ;
  assign n25035 = x1160 & ~n25034 ;
  assign n25036 = ~n24973 & n25035 ;
  assign n25037 = x644 & ~n24971 ;
  assign n25038 = x715 | n25037 ;
  assign n25039 = ( x644 & x715 ) | ( x644 & n25031 ) | ( x715 & n25031 ) ;
  assign n25040 = ( ~x644 & x715 ) | ( ~x644 & n24916 ) | ( x715 & n24916 ) ;
  assign n25041 = n25039 & n25040 ;
  assign n25042 = x1160 | n25041 ;
  assign n25043 = n25038 & ~n25042 ;
  assign n25044 = n25036 | n25043 ;
  assign n25045 = x790 & n25044 ;
  assign n25046 = n18621 & n25025 ;
  assign n25047 = ( x629 & n24957 ) | ( x629 & n25046 ) | ( n24957 & n25046 ) ;
  assign n25048 = ( ~x629 & n24954 ) | ( ~x629 & n25046 ) | ( n24954 & n25046 ) ;
  assign n25049 = n25047 | n25048 ;
  assign n25050 = x792 & n25049 ;
  assign n25051 = x648 & ~n25019 ;
  assign n25052 = ( x619 & x1159 ) | ( x619 & n24945 ) | ( x1159 & n24945 ) ;
  assign n25053 = x627 | n25006 ;
  assign n25054 = ( x618 & x1154 ) | ( x618 & ~n24942 ) | ( x1154 & ~n24942 ) ;
  assign n25055 = x660 | n24995 ;
  assign n25056 = ( x609 & x1155 ) | ( x609 & ~n24939 ) | ( x1155 & ~n24939 ) ;
  assign n25057 = x608 | n24933 ;
  assign n25058 = ( x625 & x1153 ) | ( x625 & ~n24987 ) | ( x1153 & ~n24987 ) ;
  assign n25059 = x734 & ~n24985 ;
  assign n25060 = ( x182 & ~x756 ) | ( x182 & n15797 ) | ( ~x756 & n15797 ) ;
  assign n25061 = ( x182 & x756 ) | ( x182 & n15872 ) | ( x756 & n15872 ) ;
  assign n25062 = n25060 & ~n25061 ;
  assign n25063 = x39 & ~n25062 ;
  assign n25064 = ( x182 & ~x756 ) | ( x182 & n15583 ) | ( ~x756 & n15583 ) ;
  assign n25065 = ( x182 & x756 ) | ( x182 & n15699 ) | ( x756 & n15699 ) ;
  assign n25066 = ~n25064 & n25065 ;
  assign n25067 = n25063 & ~n25066 ;
  assign n25068 = ( ~x182 & x756 ) | ( ~x182 & n15887 ) | ( x756 & n15887 ) ;
  assign n25069 = ( x182 & x756 ) | ( x182 & ~n15891 ) | ( x756 & ~n15891 ) ;
  assign n25070 = n25068 & n25069 ;
  assign n25071 = ( ~x182 & x756 ) | ( ~x182 & n15894 ) | ( x756 & n15894 ) ;
  assign n25072 = ( x182 & x756 ) | ( x182 & ~n15897 ) | ( x756 & ~n15897 ) ;
  assign n25073 = n25071 | n25072 ;
  assign n25074 = ~n25070 & n25073 ;
  assign n25075 = x39 | n25074 ;
  assign n25076 = ~x38 & n25075 ;
  assign n25077 = ~n25067 & n25076 ;
  assign n25078 = x756 | n15758 ;
  assign n25079 = n17573 & n25078 ;
  assign n25080 = x182 | n25079 ;
  assign n25081 = n15529 | n24744 ;
  assign n25082 = x182 & n25081 ;
  assign n25083 = ~n4810 & n25082 ;
  assign n25084 = x38 & ~n25083 ;
  assign n25085 = n25080 & n25084 ;
  assign n25086 = x734 | n25085 ;
  assign n25087 = n25077 | n25086 ;
  assign n25088 = ~n2032 & n25087 ;
  assign n25089 = ~n25059 & n25088 ;
  assign n25090 = n24974 | n25089 ;
  assign n25091 = ( x625 & ~x1153 ) | ( x625 & n25090 ) | ( ~x1153 & n25090 ) ;
  assign n25092 = ~n25058 & n25091 ;
  assign n25093 = n25057 | n25092 ;
  assign n25094 = x608 & ~n24936 ;
  assign n25095 = ( x625 & x1153 ) | ( x625 & n24987 ) | ( x1153 & n24987 ) ;
  assign n25096 = ( ~x625 & x1153 ) | ( ~x625 & n25090 ) | ( x1153 & n25090 ) ;
  assign n25097 = n25095 & n25096 ;
  assign n25098 = n25094 & ~n25097 ;
  assign n25099 = n25093 & ~n25098 ;
  assign n25100 = x778 & ~n25099 ;
  assign n25101 = x778 | n25090 ;
  assign n25102 = ~n25100 & n25101 ;
  assign n25103 = ( x609 & ~x1155 ) | ( x609 & n25102 ) | ( ~x1155 & n25102 ) ;
  assign n25104 = ~n25056 & n25103 ;
  assign n25105 = n25055 | n25104 ;
  assign n25106 = x660 & ~n24999 ;
  assign n25107 = ( x609 & x1155 ) | ( x609 & n24939 ) | ( x1155 & n24939 ) ;
  assign n25108 = ( ~x609 & x1155 ) | ( ~x609 & n25102 ) | ( x1155 & n25102 ) ;
  assign n25109 = n25107 & n25108 ;
  assign n25110 = n25106 & ~n25109 ;
  assign n25111 = n25105 & ~n25110 ;
  assign n25112 = x785 & ~n25111 ;
  assign n25113 = x785 | n25102 ;
  assign n25114 = ~n25112 & n25113 ;
  assign n25115 = ( x618 & ~x1154 ) | ( x618 & n25114 ) | ( ~x1154 & n25114 ) ;
  assign n25116 = ~n25054 & n25115 ;
  assign n25117 = n25053 | n25116 ;
  assign n25118 = x627 & ~n25009 ;
  assign n25119 = ( x618 & x1154 ) | ( x618 & n24942 ) | ( x1154 & n24942 ) ;
  assign n25120 = ( ~x618 & x1154 ) | ( ~x618 & n25114 ) | ( x1154 & n25114 ) ;
  assign n25121 = n25119 & n25120 ;
  assign n25122 = n25118 & ~n25121 ;
  assign n25123 = n25117 & ~n25122 ;
  assign n25124 = x781 & ~n25123 ;
  assign n25125 = x781 | n25114 ;
  assign n25126 = ~n25124 & n25125 ;
  assign n25127 = ( ~x619 & x1159 ) | ( ~x619 & n25126 ) | ( x1159 & n25126 ) ;
  assign n25128 = n25052 & n25127 ;
  assign n25129 = n25051 & ~n25128 ;
  assign n25130 = x648 | n25016 ;
  assign n25131 = ( x619 & x1159 ) | ( x619 & ~n24945 ) | ( x1159 & ~n24945 ) ;
  assign n25132 = ( x619 & ~x1159 ) | ( x619 & n25126 ) | ( ~x1159 & n25126 ) ;
  assign n25133 = ~n25131 & n25132 ;
  assign n25134 = n25130 | n25133 ;
  assign n25135 = x789 & n25134 ;
  assign n25136 = ~n25129 & n25135 ;
  assign n25137 = ~x789 & n25126 ;
  assign n25138 = n16177 | n25137 ;
  assign n25139 = n25136 | n25138 ;
  assign n25140 = n16115 & ~n24947 ;
  assign n25141 = ( x626 & ~n15419 ) | ( x626 & n24916 ) | ( ~n15419 & n24916 ) ;
  assign n25142 = ( x626 & n15419 ) | ( x626 & ~n25022 ) | ( n15419 & ~n25022 ) ;
  assign n25143 = ~n25141 & n25142 ;
  assign n25144 = n25140 | n25143 ;
  assign n25145 = ( x626 & n15418 ) | ( x626 & ~n24916 ) | ( n15418 & ~n24916 ) ;
  assign n25146 = ( x626 & ~n15418 ) | ( x626 & n25022 ) | ( ~n15418 & n25022 ) ;
  assign n25147 = n25145 & ~n25146 ;
  assign n25148 = n25144 | n25147 ;
  assign n25149 = x788 & n25148 ;
  assign n25150 = n18434 | n25149 ;
  assign n25151 = n25139 & ~n25150 ;
  assign n25152 = n25050 | n25151 ;
  assign n25153 = ~n18431 & n25152 ;
  assign n25154 = n18610 & n25028 ;
  assign n25155 = n15139 & n24968 ;
  assign n25156 = n15138 & n24964 ;
  assign n25157 = n25155 | n25156 ;
  assign n25158 = n25154 | n25157 ;
  assign n25159 = x787 & n25158 ;
  assign n25160 = n25153 | n25159 ;
  assign n25161 = ( x644 & ~x790 ) | ( x644 & n25035 ) | ( ~x790 & n25035 ) ;
  assign n25162 = ( x644 & x790 ) | ( x644 & n25042 ) | ( x790 & n25042 ) ;
  assign n25163 = ~n25161 & n25162 ;
  assign n25164 = n25160 | n25163 ;
  assign n25165 = ~n25045 & n25164 ;
  assign n25166 = ( ~x832 & n6785 ) | ( ~x832 & n25165 ) | ( n6785 & n25165 ) ;
  assign n25167 = ( ~x182 & x832 ) | ( ~x182 & n6785 ) | ( x832 & n6785 ) ;
  assign n25168 = n25166 & ~n25167 ;
  assign n25169 = n24915 | n25168 ;
  assign n25170 = x183 | n1290 ;
  assign n25171 = ~x755 & n14840 ;
  assign n25172 = n25170 & ~n25171 ;
  assign n25173 = n16060 | n25172 ;
  assign n25174 = ~x785 & n25173 ;
  assign n25175 = ~n15094 & n25171 ;
  assign n25176 = n25173 | n25175 ;
  assign n25177 = x1155 & n25176 ;
  assign n25178 = ~x1155 & n25170 ;
  assign n25179 = ~n25175 & n25178 ;
  assign n25180 = n25177 | n25179 ;
  assign n25181 = x785 & n25180 ;
  assign n25182 = n25174 | n25181 ;
  assign n25183 = ~x781 & n25182 ;
  assign n25184 = n16075 | n25182 ;
  assign n25185 = x1154 & n25184 ;
  assign n25186 = n16078 | n25182 ;
  assign n25187 = ~x1154 & n25186 ;
  assign n25188 = n25185 | n25187 ;
  assign n25189 = x781 & n25188 ;
  assign n25190 = n25183 | n25189 ;
  assign n25191 = ~x789 & n25190 ;
  assign n25192 = n20948 | n25190 ;
  assign n25193 = x1159 & n25192 ;
  assign n25194 = n20951 | n25190 ;
  assign n25195 = ~x1159 & n25194 ;
  assign n25196 = n25193 | n25195 ;
  assign n25197 = x789 & n25196 ;
  assign n25198 = n25191 | n25197 ;
  assign n25199 = n16176 | n25198 ;
  assign n25200 = n16176 & ~n25170 ;
  assign n25201 = n25199 & ~n25200 ;
  assign n25202 = n15134 | n25201 ;
  assign n25203 = n15134 & ~n25170 ;
  assign n25204 = n25202 & ~n25203 ;
  assign n25205 = n18610 & n25204 ;
  assign n25206 = ( x647 & x1157 ) | ( x647 & ~n25170 ) | ( x1157 & ~n25170 ) ;
  assign n25207 = ~x725 & n15202 ;
  assign n25208 = n25170 & ~n25207 ;
  assign n25209 = x778 | n25208 ;
  assign n25210 = ~x625 & n25207 ;
  assign n25211 = n25208 | n25210 ;
  assign n25212 = x1153 & n25211 ;
  assign n25213 = ~x1153 & n25170 ;
  assign n25214 = ~n25210 & n25213 ;
  assign n25215 = x778 & ~n25214 ;
  assign n25216 = ~n25212 & n25215 ;
  assign n25217 = n25209 & ~n25216 ;
  assign n25218 = n16043 | n25217 ;
  assign n25219 = n16045 | n25218 ;
  assign n25220 = n16047 | n25219 ;
  assign n25221 = n16049 | n25220 ;
  assign n25222 = n16055 | n25221 ;
  assign n25223 = ( x647 & ~x1157 ) | ( x647 & n25222 ) | ( ~x1157 & n25222 ) ;
  assign n25224 = ~n25206 & n25223 ;
  assign n25225 = x630 & n25224 ;
  assign n25226 = x647 & n25222 ;
  assign n25227 = ~x647 & n25170 ;
  assign n25228 = n25226 | n25227 ;
  assign n25229 = n15138 & n25228 ;
  assign n25230 = n25225 | n25229 ;
  assign n25231 = n25205 | n25230 ;
  assign n25232 = x787 & n25231 ;
  assign n25233 = n16115 & ~n25220 ;
  assign n25234 = ( x626 & ~n15419 ) | ( x626 & n25170 ) | ( ~n15419 & n25170 ) ;
  assign n25235 = ( x626 & n15419 ) | ( x626 & ~n25198 ) | ( n15419 & ~n25198 ) ;
  assign n25236 = ~n25234 & n25235 ;
  assign n25237 = n25233 | n25236 ;
  assign n25238 = ( x626 & n15418 ) | ( x626 & ~n25170 ) | ( n15418 & ~n25170 ) ;
  assign n25239 = ( x626 & ~n15418 ) | ( x626 & n25198 ) | ( ~n15418 & n25198 ) ;
  assign n25240 = n25238 & ~n25239 ;
  assign n25241 = n25237 | n25240 ;
  assign n25242 = x788 & n25241 ;
  assign n25243 = x648 & ~n25195 ;
  assign n25244 = ( x619 & x1159 ) | ( x619 & n25219 ) | ( x1159 & n25219 ) ;
  assign n25245 = x627 | n25185 ;
  assign n25246 = ( x618 & x1154 ) | ( x618 & ~n25218 ) | ( x1154 & ~n25218 ) ;
  assign n25247 = x660 | n25177 ;
  assign n25248 = ( x609 & x1155 ) | ( x609 & ~n25217 ) | ( x1155 & ~n25217 ) ;
  assign n25249 = n14839 | n25208 ;
  assign n25250 = x625 & ~n25249 ;
  assign n25251 = n25172 & n25249 ;
  assign n25252 = n25250 | n25251 ;
  assign n25253 = n25213 & n25252 ;
  assign n25254 = x608 | n25212 ;
  assign n25255 = n25253 | n25254 ;
  assign n25256 = x1153 & n25172 ;
  assign n25257 = ~n25250 & n25256 ;
  assign n25258 = x608 & ~n25214 ;
  assign n25259 = ~n25257 & n25258 ;
  assign n25260 = n25255 & ~n25259 ;
  assign n25261 = x778 & ~n25260 ;
  assign n25262 = x778 | n25251 ;
  assign n25263 = ~n25261 & n25262 ;
  assign n25264 = ( x609 & ~x1155 ) | ( x609 & n25263 ) | ( ~x1155 & n25263 ) ;
  assign n25265 = ~n25248 & n25264 ;
  assign n25266 = n25247 | n25265 ;
  assign n25267 = x660 & ~n25179 ;
  assign n25268 = ( x609 & x1155 ) | ( x609 & n25217 ) | ( x1155 & n25217 ) ;
  assign n25269 = ( ~x609 & x1155 ) | ( ~x609 & n25263 ) | ( x1155 & n25263 ) ;
  assign n25270 = n25268 & n25269 ;
  assign n25271 = n25267 & ~n25270 ;
  assign n25272 = n25266 & ~n25271 ;
  assign n25273 = x785 & ~n25272 ;
  assign n25274 = x785 | n25263 ;
  assign n25275 = ~n25273 & n25274 ;
  assign n25276 = ( x618 & ~x1154 ) | ( x618 & n25275 ) | ( ~x1154 & n25275 ) ;
  assign n25277 = ~n25246 & n25276 ;
  assign n25278 = n25245 | n25277 ;
  assign n25279 = x627 & ~n25187 ;
  assign n25280 = ( x618 & x1154 ) | ( x618 & n25218 ) | ( x1154 & n25218 ) ;
  assign n25281 = ( ~x618 & x1154 ) | ( ~x618 & n25275 ) | ( x1154 & n25275 ) ;
  assign n25282 = n25280 & n25281 ;
  assign n25283 = n25279 & ~n25282 ;
  assign n25284 = n25278 & ~n25283 ;
  assign n25285 = x781 & ~n25284 ;
  assign n25286 = x781 | n25275 ;
  assign n25287 = ~n25285 & n25286 ;
  assign n25288 = ( ~x619 & x1159 ) | ( ~x619 & n25287 ) | ( x1159 & n25287 ) ;
  assign n25289 = n25244 & n25288 ;
  assign n25290 = n25243 & ~n25289 ;
  assign n25291 = x648 | n25193 ;
  assign n25292 = ( x619 & x1159 ) | ( x619 & ~n25219 ) | ( x1159 & ~n25219 ) ;
  assign n25293 = ( x619 & ~x1159 ) | ( x619 & n25287 ) | ( ~x1159 & n25287 ) ;
  assign n25294 = ~n25292 & n25293 ;
  assign n25295 = n25291 | n25294 ;
  assign n25296 = x789 & n25295 ;
  assign n25297 = ~n25290 & n25296 ;
  assign n25298 = ~x789 & n25287 ;
  assign n25299 = n16177 | n25298 ;
  assign n25300 = n25297 | n25299 ;
  assign n25301 = ~n25242 & n25300 ;
  assign n25302 = n18434 | n25301 ;
  assign n25303 = n16650 | n25221 ;
  assign n25304 = n16051 & ~n25201 ;
  assign n25305 = n25303 & ~n25304 ;
  assign n25306 = ( x629 & ~x792 ) | ( x629 & n25305 ) | ( ~x792 & n25305 ) ;
  assign n25307 = n16052 & ~n25201 ;
  assign n25308 = n16643 & ~n25221 ;
  assign n25309 = n25307 | n25308 ;
  assign n25310 = ( x629 & x792 ) | ( x629 & n25309 ) | ( x792 & n25309 ) ;
  assign n25311 = ~n25306 & n25310 ;
  assign n25312 = n18431 | n25311 ;
  assign n25313 = n25302 & ~n25312 ;
  assign n25314 = n25232 | n25313 ;
  assign n25315 = ( x790 & x832 ) | ( x790 & n25314 ) | ( x832 & n25314 ) ;
  assign n25316 = n15141 | n25204 ;
  assign n25317 = n15141 & ~n25170 ;
  assign n25318 = n25316 & ~n25317 ;
  assign n25319 = ( x644 & x715 ) | ( x644 & ~n25318 ) | ( x715 & ~n25318 ) ;
  assign n25320 = ( x644 & ~x715 ) | ( x644 & n25170 ) | ( ~x715 & n25170 ) ;
  assign n25321 = ~n25319 & n25320 ;
  assign n25322 = x1160 & ~n25321 ;
  assign n25323 = ~x787 & n25222 ;
  assign n25324 = x1157 & n25228 ;
  assign n25325 = n25224 | n25324 ;
  assign n25326 = x787 & n25325 ;
  assign n25327 = n25323 | n25326 ;
  assign n25328 = ( x644 & x715 ) | ( x644 & n25327 ) | ( x715 & n25327 ) ;
  assign n25329 = ( ~x644 & x715 ) | ( ~x644 & n25314 ) | ( x715 & n25314 ) ;
  assign n25330 = n25328 & n25329 ;
  assign n25331 = n25322 & ~n25330 ;
  assign n25332 = ( x644 & x715 ) | ( x644 & n25318 ) | ( x715 & n25318 ) ;
  assign n25333 = ( ~x644 & x715 ) | ( ~x644 & n25170 ) | ( x715 & n25170 ) ;
  assign n25334 = n25332 & n25333 ;
  assign n25335 = x1160 | n25334 ;
  assign n25336 = ( x644 & x715 ) | ( x644 & ~n25327 ) | ( x715 & ~n25327 ) ;
  assign n25337 = ( x644 & ~x715 ) | ( x644 & n25314 ) | ( ~x715 & n25314 ) ;
  assign n25338 = ~n25336 & n25337 ;
  assign n25339 = n25335 | n25338 ;
  assign n25340 = ~n25331 & n25339 ;
  assign n25341 = ( ~x790 & x832 ) | ( ~x790 & n25340 ) | ( x832 & n25340 ) ;
  assign n25342 = n25315 & n25341 ;
  assign n25343 = x183 | n14834 ;
  assign n25344 = n15414 & n25343 ;
  assign n25345 = x725 | n2032 ;
  assign n25346 = ~n25343 & n25345 ;
  assign n25347 = x183 & n16323 ;
  assign n25348 = x38 | n25347 ;
  assign n25349 = ~n2032 & n25348 ;
  assign n25350 = x183 | n16319 ;
  assign n25351 = ~n25349 & n25350 ;
  assign n25352 = x183 | n15070 ;
  assign n25353 = n15375 & n25352 ;
  assign n25354 = x725 | n25353 ;
  assign n25355 = n25351 | n25354 ;
  assign n25356 = ~n25346 & n25355 ;
  assign n25357 = ~x778 & n25356 ;
  assign n25358 = ( x625 & x1153 ) | ( x625 & n25343 ) | ( x1153 & n25343 ) ;
  assign n25359 = ( ~x625 & x1153 ) | ( ~x625 & n25356 ) | ( x1153 & n25356 ) ;
  assign n25360 = n25358 & n25359 ;
  assign n25361 = ( x625 & x1153 ) | ( x625 & ~n25343 ) | ( x1153 & ~n25343 ) ;
  assign n25362 = ( x625 & ~x1153 ) | ( x625 & n25356 ) | ( ~x1153 & n25356 ) ;
  assign n25363 = ~n25361 & n25362 ;
  assign n25364 = n25360 | n25363 ;
  assign n25365 = x778 & n25364 ;
  assign n25366 = n25357 | n25365 ;
  assign n25367 = ~n15400 & n25366 ;
  assign n25368 = n15400 & n25343 ;
  assign n25369 = n25367 | n25368 ;
  assign n25370 = n15407 | n25369 ;
  assign n25371 = n15407 & ~n25343 ;
  assign n25372 = n25370 & ~n25371 ;
  assign n25373 = ~n15414 & n25372 ;
  assign n25374 = n25344 | n25373 ;
  assign n25375 = n15421 | n25374 ;
  assign n25376 = n15421 & ~n25343 ;
  assign n25377 = n25375 & ~n25376 ;
  assign n25378 = ~x792 & n25377 ;
  assign n25379 = ( x628 & x1156 ) | ( x628 & n25343 ) | ( x1156 & n25343 ) ;
  assign n25380 = ( ~x628 & x1156 ) | ( ~x628 & n25377 ) | ( x1156 & n25377 ) ;
  assign n25381 = n25379 & n25380 ;
  assign n25382 = ( x628 & x1156 ) | ( x628 & ~n25343 ) | ( x1156 & ~n25343 ) ;
  assign n25383 = ( x628 & ~x1156 ) | ( x628 & n25377 ) | ( ~x1156 & n25377 ) ;
  assign n25384 = ~n25382 & n25383 ;
  assign n25385 = n25381 | n25384 ;
  assign n25386 = x792 & n25385 ;
  assign n25387 = n25378 | n25386 ;
  assign n25388 = x787 | n25387 ;
  assign n25389 = x647 & n25387 ;
  assign n25390 = ~x647 & n25343 ;
  assign n25391 = n25389 | n25390 ;
  assign n25392 = ( ~x787 & x1157 ) | ( ~x787 & n25391 ) | ( x1157 & n25391 ) ;
  assign n25393 = ~x647 & n25387 ;
  assign n25394 = x647 & n25343 ;
  assign n25395 = n25393 | n25394 ;
  assign n25396 = ( x787 & x1157 ) | ( x787 & ~n25395 ) | ( x1157 & ~n25395 ) ;
  assign n25397 = ~n25392 & n25396 ;
  assign n25398 = n25388 & ~n25397 ;
  assign n25399 = x644 | n25398 ;
  assign n25400 = x715 & n25399 ;
  assign n25401 = x183 & n2032 ;
  assign n25402 = ~x755 & n15072 ;
  assign n25403 = n25352 & ~n25402 ;
  assign n25404 = x38 & ~n25403 ;
  assign n25405 = ~x183 & x755 ;
  assign n25406 = ~n14936 & n25405 ;
  assign n25407 = ( ~x183 & x755 ) | ( ~x183 & n15063 ) | ( x755 & n15063 ) ;
  assign n25408 = ( x183 & x755 ) | ( x183 & ~n14933 ) | ( x755 & ~n14933 ) ;
  assign n25409 = n25407 | n25408 ;
  assign n25410 = ~n25406 & n25409 ;
  assign n25411 = x38 | n25410 ;
  assign n25412 = ~n25404 & n25411 ;
  assign n25413 = ~n2032 & n25412 ;
  assign n25414 = n25401 | n25413 ;
  assign n25415 = ~n15082 & n25414 ;
  assign n25416 = n15082 & n25343 ;
  assign n25417 = n25415 | n25416 ;
  assign n25418 = ~x785 & n25417 ;
  assign n25419 = ~n15088 & n25343 ;
  assign n25420 = x609 & n25415 ;
  assign n25421 = n25419 | n25420 ;
  assign n25422 = x1155 & n25421 ;
  assign n25423 = n15094 & n25343 ;
  assign n25424 = ~x609 & n25415 ;
  assign n25425 = n25423 | n25424 ;
  assign n25426 = ~x1155 & n25425 ;
  assign n25427 = n25422 | n25426 ;
  assign n25428 = x785 & n25427 ;
  assign n25429 = n25418 | n25428 ;
  assign n25430 = ~x781 & n25429 ;
  assign n25431 = ( x618 & x1154 ) | ( x618 & n25343 ) | ( x1154 & n25343 ) ;
  assign n25432 = ( ~x618 & x1154 ) | ( ~x618 & n25429 ) | ( x1154 & n25429 ) ;
  assign n25433 = n25431 & n25432 ;
  assign n25434 = ( x618 & x1154 ) | ( x618 & ~n25343 ) | ( x1154 & ~n25343 ) ;
  assign n25435 = ( x618 & ~x1154 ) | ( x618 & n25429 ) | ( ~x1154 & n25429 ) ;
  assign n25436 = ~n25434 & n25435 ;
  assign n25437 = n25433 | n25436 ;
  assign n25438 = x781 & n25437 ;
  assign n25439 = n25430 | n25438 ;
  assign n25440 = ~x789 & n25439 ;
  assign n25441 = ( x619 & x1159 ) | ( x619 & n25343 ) | ( x1159 & n25343 ) ;
  assign n25442 = ( ~x619 & x1159 ) | ( ~x619 & n25439 ) | ( x1159 & n25439 ) ;
  assign n25443 = n25441 & n25442 ;
  assign n25444 = ( x619 & x1159 ) | ( x619 & ~n25343 ) | ( x1159 & ~n25343 ) ;
  assign n25445 = ( x619 & ~x1159 ) | ( x619 & n25439 ) | ( ~x1159 & n25439 ) ;
  assign n25446 = ~n25444 & n25445 ;
  assign n25447 = n25443 | n25446 ;
  assign n25448 = x789 & n25447 ;
  assign n25449 = n25440 | n25448 ;
  assign n25450 = n16176 | n25449 ;
  assign n25451 = n16176 & ~n25343 ;
  assign n25452 = n25450 & ~n25451 ;
  assign n25453 = n15134 | n25452 ;
  assign n25454 = n15134 & ~n25343 ;
  assign n25455 = n25453 & ~n25454 ;
  assign n25456 = n15141 | n25455 ;
  assign n25457 = n15141 & ~n25343 ;
  assign n25458 = n25456 & ~n25457 ;
  assign n25459 = ( x644 & x715 ) | ( x644 & ~n25458 ) | ( x715 & ~n25458 ) ;
  assign n25460 = ( x644 & ~x715 ) | ( x644 & n25343 ) | ( ~x715 & n25343 ) ;
  assign n25461 = ~n25459 & n25460 ;
  assign n25462 = x1160 & ~n25461 ;
  assign n25463 = ~n25400 & n25462 ;
  assign n25464 = x644 & ~n25398 ;
  assign n25465 = x715 | n25464 ;
  assign n25466 = ( x644 & x715 ) | ( x644 & n25458 ) | ( x715 & n25458 ) ;
  assign n25467 = ( ~x644 & x715 ) | ( ~x644 & n25343 ) | ( x715 & n25343 ) ;
  assign n25468 = n25466 & n25467 ;
  assign n25469 = x1160 | n25468 ;
  assign n25470 = n25465 & ~n25469 ;
  assign n25471 = n25463 | n25470 ;
  assign n25472 = x790 & n25471 ;
  assign n25473 = n18621 & n25452 ;
  assign n25474 = ( x629 & n25384 ) | ( x629 & n25473 ) | ( n25384 & n25473 ) ;
  assign n25475 = ( ~x629 & n25381 ) | ( ~x629 & n25473 ) | ( n25381 & n25473 ) ;
  assign n25476 = n25474 | n25475 ;
  assign n25477 = x792 & n25476 ;
  assign n25478 = x648 & ~n25446 ;
  assign n25479 = ( x619 & x1159 ) | ( x619 & n25372 ) | ( x1159 & n25372 ) ;
  assign n25480 = x627 | n25433 ;
  assign n25481 = ( x618 & x1154 ) | ( x618 & ~n25369 ) | ( x1154 & ~n25369 ) ;
  assign n25482 = x660 | n25422 ;
  assign n25483 = ( x609 & x1155 ) | ( x609 & ~n25366 ) | ( x1155 & ~n25366 ) ;
  assign n25484 = x608 | n25360 ;
  assign n25485 = ( x625 & x1153 ) | ( x625 & ~n25414 ) | ( x1153 & ~n25414 ) ;
  assign n25486 = x725 & ~n25412 ;
  assign n25487 = ( x183 & ~x755 ) | ( x183 & n15797 ) | ( ~x755 & n15797 ) ;
  assign n25488 = ( x183 & x755 ) | ( x183 & n15872 ) | ( x755 & n15872 ) ;
  assign n25489 = n25487 & ~n25488 ;
  assign n25490 = x39 & ~n25489 ;
  assign n25491 = ( x183 & ~x755 ) | ( x183 & n15583 ) | ( ~x755 & n15583 ) ;
  assign n25492 = ( x183 & x755 ) | ( x183 & n15699 ) | ( x755 & n15699 ) ;
  assign n25493 = ~n25491 & n25492 ;
  assign n25494 = n25490 & ~n25493 ;
  assign n25495 = ( ~x183 & x755 ) | ( ~x183 & n15887 ) | ( x755 & n15887 ) ;
  assign n25496 = ( x183 & x755 ) | ( x183 & ~n15891 ) | ( x755 & ~n15891 ) ;
  assign n25497 = n25495 & n25496 ;
  assign n25498 = ( ~x183 & x755 ) | ( ~x183 & n15894 ) | ( x755 & n15894 ) ;
  assign n25499 = ( x183 & x755 ) | ( x183 & ~n15897 ) | ( x755 & ~n15897 ) ;
  assign n25500 = n25498 | n25499 ;
  assign n25501 = ~n25497 & n25500 ;
  assign n25502 = x39 | n25501 ;
  assign n25503 = ~x38 & n25502 ;
  assign n25504 = ~n25494 & n25503 ;
  assign n25505 = x755 | n15758 ;
  assign n25506 = n17573 & n25505 ;
  assign n25507 = x183 | n25506 ;
  assign n25508 = n15529 | n25171 ;
  assign n25509 = x183 & n25508 ;
  assign n25510 = ~n4810 & n25509 ;
  assign n25511 = x38 & ~n25510 ;
  assign n25512 = n25507 & n25511 ;
  assign n25513 = x725 | n25512 ;
  assign n25514 = n25504 | n25513 ;
  assign n25515 = ~n2032 & n25514 ;
  assign n25516 = ~n25486 & n25515 ;
  assign n25517 = n25401 | n25516 ;
  assign n25518 = ( x625 & ~x1153 ) | ( x625 & n25517 ) | ( ~x1153 & n25517 ) ;
  assign n25519 = ~n25485 & n25518 ;
  assign n25520 = n25484 | n25519 ;
  assign n25521 = x608 & ~n25363 ;
  assign n25522 = ( x625 & x1153 ) | ( x625 & n25414 ) | ( x1153 & n25414 ) ;
  assign n25523 = ( ~x625 & x1153 ) | ( ~x625 & n25517 ) | ( x1153 & n25517 ) ;
  assign n25524 = n25522 & n25523 ;
  assign n25525 = n25521 & ~n25524 ;
  assign n25526 = n25520 & ~n25525 ;
  assign n25527 = x778 & ~n25526 ;
  assign n25528 = x778 | n25517 ;
  assign n25529 = ~n25527 & n25528 ;
  assign n25530 = ( x609 & ~x1155 ) | ( x609 & n25529 ) | ( ~x1155 & n25529 ) ;
  assign n25531 = ~n25483 & n25530 ;
  assign n25532 = n25482 | n25531 ;
  assign n25533 = x660 & ~n25426 ;
  assign n25534 = ( x609 & x1155 ) | ( x609 & n25366 ) | ( x1155 & n25366 ) ;
  assign n25535 = ( ~x609 & x1155 ) | ( ~x609 & n25529 ) | ( x1155 & n25529 ) ;
  assign n25536 = n25534 & n25535 ;
  assign n25537 = n25533 & ~n25536 ;
  assign n25538 = n25532 & ~n25537 ;
  assign n25539 = x785 & ~n25538 ;
  assign n25540 = x785 | n25529 ;
  assign n25541 = ~n25539 & n25540 ;
  assign n25542 = ( x618 & ~x1154 ) | ( x618 & n25541 ) | ( ~x1154 & n25541 ) ;
  assign n25543 = ~n25481 & n25542 ;
  assign n25544 = n25480 | n25543 ;
  assign n25545 = x627 & ~n25436 ;
  assign n25546 = ( x618 & x1154 ) | ( x618 & n25369 ) | ( x1154 & n25369 ) ;
  assign n25547 = ( ~x618 & x1154 ) | ( ~x618 & n25541 ) | ( x1154 & n25541 ) ;
  assign n25548 = n25546 & n25547 ;
  assign n25549 = n25545 & ~n25548 ;
  assign n25550 = n25544 & ~n25549 ;
  assign n25551 = x781 & ~n25550 ;
  assign n25552 = x781 | n25541 ;
  assign n25553 = ~n25551 & n25552 ;
  assign n25554 = ( ~x619 & x1159 ) | ( ~x619 & n25553 ) | ( x1159 & n25553 ) ;
  assign n25555 = n25479 & n25554 ;
  assign n25556 = n25478 & ~n25555 ;
  assign n25557 = x648 | n25443 ;
  assign n25558 = ( x619 & x1159 ) | ( x619 & ~n25372 ) | ( x1159 & ~n25372 ) ;
  assign n25559 = ( x619 & ~x1159 ) | ( x619 & n25553 ) | ( ~x1159 & n25553 ) ;
  assign n25560 = ~n25558 & n25559 ;
  assign n25561 = n25557 | n25560 ;
  assign n25562 = x789 & n25561 ;
  assign n25563 = ~n25556 & n25562 ;
  assign n25564 = ~x789 & n25553 ;
  assign n25565 = n16177 | n25564 ;
  assign n25566 = n25563 | n25565 ;
  assign n25567 = n16115 & ~n25374 ;
  assign n25568 = ( x626 & ~n15419 ) | ( x626 & n25343 ) | ( ~n15419 & n25343 ) ;
  assign n25569 = ( x626 & n15419 ) | ( x626 & ~n25449 ) | ( n15419 & ~n25449 ) ;
  assign n25570 = ~n25568 & n25569 ;
  assign n25571 = n25567 | n25570 ;
  assign n25572 = ( x626 & n15418 ) | ( x626 & ~n25343 ) | ( n15418 & ~n25343 ) ;
  assign n25573 = ( x626 & ~n15418 ) | ( x626 & n25449 ) | ( ~n15418 & n25449 ) ;
  assign n25574 = n25572 & ~n25573 ;
  assign n25575 = n25571 | n25574 ;
  assign n25576 = x788 & n25575 ;
  assign n25577 = n18434 | n25576 ;
  assign n25578 = n25566 & ~n25577 ;
  assign n25579 = n25477 | n25578 ;
  assign n25580 = ~n18431 & n25579 ;
  assign n25581 = n18610 & n25455 ;
  assign n25582 = n15139 & n25395 ;
  assign n25583 = n15138 & n25391 ;
  assign n25584 = n25582 | n25583 ;
  assign n25585 = n25581 | n25584 ;
  assign n25586 = x787 & n25585 ;
  assign n25587 = n25580 | n25586 ;
  assign n25588 = ( x644 & ~x790 ) | ( x644 & n25462 ) | ( ~x790 & n25462 ) ;
  assign n25589 = ( x644 & x790 ) | ( x644 & n25469 ) | ( x790 & n25469 ) ;
  assign n25590 = ~n25588 & n25589 ;
  assign n25591 = n25587 | n25590 ;
  assign n25592 = ~n25472 & n25591 ;
  assign n25593 = ( ~x832 & n6785 ) | ( ~x832 & n25592 ) | ( n6785 & n25592 ) ;
  assign n25594 = ( ~x183 & x832 ) | ( ~x183 & n6785 ) | ( x832 & n6785 ) ;
  assign n25595 = n25593 & ~n25594 ;
  assign n25596 = n25342 | n25595 ;
  assign n25597 = x184 | n1290 ;
  assign n25598 = ~x777 & n14840 ;
  assign n25599 = n25597 & ~n25598 ;
  assign n25600 = n16060 | n25599 ;
  assign n25601 = ~x785 & n25600 ;
  assign n25602 = ~n15094 & n25598 ;
  assign n25603 = n25600 | n25602 ;
  assign n25604 = x1155 & n25603 ;
  assign n25605 = ~x1155 & n25597 ;
  assign n25606 = ~n25602 & n25605 ;
  assign n25607 = n25604 | n25606 ;
  assign n25608 = x785 & n25607 ;
  assign n25609 = n25601 | n25608 ;
  assign n25610 = ~x781 & n25609 ;
  assign n25611 = n16075 | n25609 ;
  assign n25612 = x1154 & n25611 ;
  assign n25613 = n16078 | n25609 ;
  assign n25614 = ~x1154 & n25613 ;
  assign n25615 = n25612 | n25614 ;
  assign n25616 = x781 & n25615 ;
  assign n25617 = n25610 | n25616 ;
  assign n25618 = ~x789 & n25617 ;
  assign n25619 = n20948 | n25617 ;
  assign n25620 = x1159 & n25619 ;
  assign n25621 = n20951 | n25617 ;
  assign n25622 = ~x1159 & n25621 ;
  assign n25623 = n25620 | n25622 ;
  assign n25624 = x789 & n25623 ;
  assign n25625 = n25618 | n25624 ;
  assign n25626 = n16176 | n25625 ;
  assign n25627 = n16176 & ~n25597 ;
  assign n25628 = n25626 & ~n25627 ;
  assign n25629 = n15134 | n25628 ;
  assign n25630 = n15134 & ~n25597 ;
  assign n25631 = n25629 & ~n25630 ;
  assign n25632 = n18610 & n25631 ;
  assign n25633 = ( x647 & x1157 ) | ( x647 & ~n25597 ) | ( x1157 & ~n25597 ) ;
  assign n25634 = ~x737 & n15202 ;
  assign n25635 = n25597 & ~n25634 ;
  assign n25636 = x778 | n25635 ;
  assign n25637 = ~x625 & n25634 ;
  assign n25638 = n25635 | n25637 ;
  assign n25639 = x1153 & n25638 ;
  assign n25640 = ~x1153 & n25597 ;
  assign n25641 = ~n25637 & n25640 ;
  assign n25642 = x778 & ~n25641 ;
  assign n25643 = ~n25639 & n25642 ;
  assign n25644 = n25636 & ~n25643 ;
  assign n25645 = n16043 | n25644 ;
  assign n25646 = n16045 | n25645 ;
  assign n25647 = n16047 | n25646 ;
  assign n25648 = n16049 | n25647 ;
  assign n25649 = n16055 | n25648 ;
  assign n25650 = ( x647 & ~x1157 ) | ( x647 & n25649 ) | ( ~x1157 & n25649 ) ;
  assign n25651 = ~n25633 & n25650 ;
  assign n25652 = x630 & n25651 ;
  assign n25653 = x647 & n25649 ;
  assign n25654 = ~x647 & n25597 ;
  assign n25655 = n25653 | n25654 ;
  assign n25656 = n15138 & n25655 ;
  assign n25657 = n25652 | n25656 ;
  assign n25658 = n25632 | n25657 ;
  assign n25659 = x787 & n25658 ;
  assign n25660 = n16115 & ~n25647 ;
  assign n25661 = ( x626 & ~n15419 ) | ( x626 & n25597 ) | ( ~n15419 & n25597 ) ;
  assign n25662 = ( x626 & n15419 ) | ( x626 & ~n25625 ) | ( n15419 & ~n25625 ) ;
  assign n25663 = ~n25661 & n25662 ;
  assign n25664 = n25660 | n25663 ;
  assign n25665 = ( x626 & n15418 ) | ( x626 & ~n25597 ) | ( n15418 & ~n25597 ) ;
  assign n25666 = ( x626 & ~n15418 ) | ( x626 & n25625 ) | ( ~n15418 & n25625 ) ;
  assign n25667 = n25665 & ~n25666 ;
  assign n25668 = n25664 | n25667 ;
  assign n25669 = x788 & n25668 ;
  assign n25670 = x648 & ~n25622 ;
  assign n25671 = ( x619 & x1159 ) | ( x619 & n25646 ) | ( x1159 & n25646 ) ;
  assign n25672 = x627 | n25612 ;
  assign n25673 = ( x618 & x1154 ) | ( x618 & ~n25645 ) | ( x1154 & ~n25645 ) ;
  assign n25674 = x660 | n25604 ;
  assign n25675 = ( x609 & x1155 ) | ( x609 & ~n25644 ) | ( x1155 & ~n25644 ) ;
  assign n25676 = n14839 | n25635 ;
  assign n25677 = x625 & ~n25676 ;
  assign n25678 = n25599 & n25676 ;
  assign n25679 = n25677 | n25678 ;
  assign n25680 = n25640 & n25679 ;
  assign n25681 = x608 | n25639 ;
  assign n25682 = n25680 | n25681 ;
  assign n25683 = x1153 & n25599 ;
  assign n25684 = ~n25677 & n25683 ;
  assign n25685 = x608 & ~n25641 ;
  assign n25686 = ~n25684 & n25685 ;
  assign n25687 = n25682 & ~n25686 ;
  assign n25688 = x778 & ~n25687 ;
  assign n25689 = x778 | n25678 ;
  assign n25690 = ~n25688 & n25689 ;
  assign n25691 = ( x609 & ~x1155 ) | ( x609 & n25690 ) | ( ~x1155 & n25690 ) ;
  assign n25692 = ~n25675 & n25691 ;
  assign n25693 = n25674 | n25692 ;
  assign n25694 = x660 & ~n25606 ;
  assign n25695 = ( x609 & x1155 ) | ( x609 & n25644 ) | ( x1155 & n25644 ) ;
  assign n25696 = ( ~x609 & x1155 ) | ( ~x609 & n25690 ) | ( x1155 & n25690 ) ;
  assign n25697 = n25695 & n25696 ;
  assign n25698 = n25694 & ~n25697 ;
  assign n25699 = n25693 & ~n25698 ;
  assign n25700 = x785 & ~n25699 ;
  assign n25701 = x785 | n25690 ;
  assign n25702 = ~n25700 & n25701 ;
  assign n25703 = ( x618 & ~x1154 ) | ( x618 & n25702 ) | ( ~x1154 & n25702 ) ;
  assign n25704 = ~n25673 & n25703 ;
  assign n25705 = n25672 | n25704 ;
  assign n25706 = x627 & ~n25614 ;
  assign n25707 = ( x618 & x1154 ) | ( x618 & n25645 ) | ( x1154 & n25645 ) ;
  assign n25708 = ( ~x618 & x1154 ) | ( ~x618 & n25702 ) | ( x1154 & n25702 ) ;
  assign n25709 = n25707 & n25708 ;
  assign n25710 = n25706 & ~n25709 ;
  assign n25711 = n25705 & ~n25710 ;
  assign n25712 = x781 & ~n25711 ;
  assign n25713 = x781 | n25702 ;
  assign n25714 = ~n25712 & n25713 ;
  assign n25715 = ( ~x619 & x1159 ) | ( ~x619 & n25714 ) | ( x1159 & n25714 ) ;
  assign n25716 = n25671 & n25715 ;
  assign n25717 = n25670 & ~n25716 ;
  assign n25718 = x648 | n25620 ;
  assign n25719 = ( x619 & x1159 ) | ( x619 & ~n25646 ) | ( x1159 & ~n25646 ) ;
  assign n25720 = ( x619 & ~x1159 ) | ( x619 & n25714 ) | ( ~x1159 & n25714 ) ;
  assign n25721 = ~n25719 & n25720 ;
  assign n25722 = n25718 | n25721 ;
  assign n25723 = x789 & n25722 ;
  assign n25724 = ~n25717 & n25723 ;
  assign n25725 = ~x789 & n25714 ;
  assign n25726 = n16177 | n25725 ;
  assign n25727 = n25724 | n25726 ;
  assign n25728 = ~n25669 & n25727 ;
  assign n25729 = n18434 | n25728 ;
  assign n25730 = n16650 | n25648 ;
  assign n25731 = n16051 & ~n25628 ;
  assign n25732 = n25730 & ~n25731 ;
  assign n25733 = ( x629 & ~x792 ) | ( x629 & n25732 ) | ( ~x792 & n25732 ) ;
  assign n25734 = n16052 & ~n25628 ;
  assign n25735 = n16643 & ~n25648 ;
  assign n25736 = n25734 | n25735 ;
  assign n25737 = ( x629 & x792 ) | ( x629 & n25736 ) | ( x792 & n25736 ) ;
  assign n25738 = ~n25733 & n25737 ;
  assign n25739 = n18431 | n25738 ;
  assign n25740 = n25729 & ~n25739 ;
  assign n25741 = n25659 | n25740 ;
  assign n25742 = ( x790 & x832 ) | ( x790 & n25741 ) | ( x832 & n25741 ) ;
  assign n25743 = n15141 | n25631 ;
  assign n25744 = n15141 & ~n25597 ;
  assign n25745 = n25743 & ~n25744 ;
  assign n25746 = ( x644 & x715 ) | ( x644 & ~n25745 ) | ( x715 & ~n25745 ) ;
  assign n25747 = ( x644 & ~x715 ) | ( x644 & n25597 ) | ( ~x715 & n25597 ) ;
  assign n25748 = ~n25746 & n25747 ;
  assign n25749 = x1160 & ~n25748 ;
  assign n25750 = ~x787 & n25649 ;
  assign n25751 = x1157 & n25655 ;
  assign n25752 = n25651 | n25751 ;
  assign n25753 = x787 & n25752 ;
  assign n25754 = n25750 | n25753 ;
  assign n25755 = ( x644 & x715 ) | ( x644 & n25754 ) | ( x715 & n25754 ) ;
  assign n25756 = ( ~x644 & x715 ) | ( ~x644 & n25741 ) | ( x715 & n25741 ) ;
  assign n25757 = n25755 & n25756 ;
  assign n25758 = n25749 & ~n25757 ;
  assign n25759 = ( x644 & x715 ) | ( x644 & n25745 ) | ( x715 & n25745 ) ;
  assign n25760 = ( ~x644 & x715 ) | ( ~x644 & n25597 ) | ( x715 & n25597 ) ;
  assign n25761 = n25759 & n25760 ;
  assign n25762 = x1160 | n25761 ;
  assign n25763 = ( x644 & x715 ) | ( x644 & ~n25754 ) | ( x715 & ~n25754 ) ;
  assign n25764 = ( x644 & ~x715 ) | ( x644 & n25741 ) | ( ~x715 & n25741 ) ;
  assign n25765 = ~n25763 & n25764 ;
  assign n25766 = n25762 | n25765 ;
  assign n25767 = ~n25758 & n25766 ;
  assign n25768 = ( ~x790 & x832 ) | ( ~x790 & n25767 ) | ( x832 & n25767 ) ;
  assign n25769 = n25742 & n25768 ;
  assign n25770 = x184 | n14834 ;
  assign n25771 = n15414 & n25770 ;
  assign n25772 = x737 | n2032 ;
  assign n25773 = ~n25770 & n25772 ;
  assign n25774 = x184 & n16323 ;
  assign n25775 = x38 | n25774 ;
  assign n25776 = ~n2032 & n25775 ;
  assign n25777 = x184 | n16319 ;
  assign n25778 = ~n25776 & n25777 ;
  assign n25779 = x184 | n15070 ;
  assign n25780 = n15375 & n25779 ;
  assign n25781 = x737 | n25780 ;
  assign n25782 = n25778 | n25781 ;
  assign n25783 = ~n25773 & n25782 ;
  assign n25784 = ~x778 & n25783 ;
  assign n25785 = ( x625 & x1153 ) | ( x625 & n25770 ) | ( x1153 & n25770 ) ;
  assign n25786 = ( ~x625 & x1153 ) | ( ~x625 & n25783 ) | ( x1153 & n25783 ) ;
  assign n25787 = n25785 & n25786 ;
  assign n25788 = ( x625 & x1153 ) | ( x625 & ~n25770 ) | ( x1153 & ~n25770 ) ;
  assign n25789 = ( x625 & ~x1153 ) | ( x625 & n25783 ) | ( ~x1153 & n25783 ) ;
  assign n25790 = ~n25788 & n25789 ;
  assign n25791 = n25787 | n25790 ;
  assign n25792 = x778 & n25791 ;
  assign n25793 = n25784 | n25792 ;
  assign n25794 = ~n15400 & n25793 ;
  assign n25795 = n15400 & n25770 ;
  assign n25796 = n25794 | n25795 ;
  assign n25797 = n15407 | n25796 ;
  assign n25798 = n15407 & ~n25770 ;
  assign n25799 = n25797 & ~n25798 ;
  assign n25800 = ~n15414 & n25799 ;
  assign n25801 = n25771 | n25800 ;
  assign n25802 = n15421 | n25801 ;
  assign n25803 = n15421 & ~n25770 ;
  assign n25804 = n25802 & ~n25803 ;
  assign n25805 = ~x792 & n25804 ;
  assign n25806 = ( x628 & x1156 ) | ( x628 & n25770 ) | ( x1156 & n25770 ) ;
  assign n25807 = ( ~x628 & x1156 ) | ( ~x628 & n25804 ) | ( x1156 & n25804 ) ;
  assign n25808 = n25806 & n25807 ;
  assign n25809 = ( x628 & x1156 ) | ( x628 & ~n25770 ) | ( x1156 & ~n25770 ) ;
  assign n25810 = ( x628 & ~x1156 ) | ( x628 & n25804 ) | ( ~x1156 & n25804 ) ;
  assign n25811 = ~n25809 & n25810 ;
  assign n25812 = n25808 | n25811 ;
  assign n25813 = x792 & n25812 ;
  assign n25814 = n25805 | n25813 ;
  assign n25815 = x787 | n25814 ;
  assign n25816 = x647 & n25814 ;
  assign n25817 = ~x647 & n25770 ;
  assign n25818 = n25816 | n25817 ;
  assign n25819 = ( ~x787 & x1157 ) | ( ~x787 & n25818 ) | ( x1157 & n25818 ) ;
  assign n25820 = ~x647 & n25814 ;
  assign n25821 = x647 & n25770 ;
  assign n25822 = n25820 | n25821 ;
  assign n25823 = ( x787 & x1157 ) | ( x787 & ~n25822 ) | ( x1157 & ~n25822 ) ;
  assign n25824 = ~n25819 & n25823 ;
  assign n25825 = n25815 & ~n25824 ;
  assign n25826 = x644 | n25825 ;
  assign n25827 = x715 & n25826 ;
  assign n25828 = x184 & n2032 ;
  assign n25829 = ~x777 & n15072 ;
  assign n25830 = n25779 & ~n25829 ;
  assign n25831 = x38 & ~n25830 ;
  assign n25832 = ~x184 & x777 ;
  assign n25833 = ~n14936 & n25832 ;
  assign n25834 = ( ~x184 & x777 ) | ( ~x184 & n15063 ) | ( x777 & n15063 ) ;
  assign n25835 = ( x184 & x777 ) | ( x184 & ~n14933 ) | ( x777 & ~n14933 ) ;
  assign n25836 = n25834 | n25835 ;
  assign n25837 = ~n25833 & n25836 ;
  assign n25838 = x38 | n25837 ;
  assign n25839 = ~n25831 & n25838 ;
  assign n25840 = ~n2032 & n25839 ;
  assign n25841 = n25828 | n25840 ;
  assign n25842 = ~n15082 & n25841 ;
  assign n25843 = n15082 & n25770 ;
  assign n25844 = n25842 | n25843 ;
  assign n25845 = ~x785 & n25844 ;
  assign n25846 = ~n15088 & n25770 ;
  assign n25847 = x609 & n25842 ;
  assign n25848 = n25846 | n25847 ;
  assign n25849 = x1155 & n25848 ;
  assign n25850 = n15094 & n25770 ;
  assign n25851 = ~x609 & n25842 ;
  assign n25852 = n25850 | n25851 ;
  assign n25853 = ~x1155 & n25852 ;
  assign n25854 = n25849 | n25853 ;
  assign n25855 = x785 & n25854 ;
  assign n25856 = n25845 | n25855 ;
  assign n25857 = ~x781 & n25856 ;
  assign n25858 = ( x618 & x1154 ) | ( x618 & n25770 ) | ( x1154 & n25770 ) ;
  assign n25859 = ( ~x618 & x1154 ) | ( ~x618 & n25856 ) | ( x1154 & n25856 ) ;
  assign n25860 = n25858 & n25859 ;
  assign n25861 = ( x618 & x1154 ) | ( x618 & ~n25770 ) | ( x1154 & ~n25770 ) ;
  assign n25862 = ( x618 & ~x1154 ) | ( x618 & n25856 ) | ( ~x1154 & n25856 ) ;
  assign n25863 = ~n25861 & n25862 ;
  assign n25864 = n25860 | n25863 ;
  assign n25865 = x781 & n25864 ;
  assign n25866 = n25857 | n25865 ;
  assign n25867 = ~x789 & n25866 ;
  assign n25868 = ( x619 & x1159 ) | ( x619 & n25770 ) | ( x1159 & n25770 ) ;
  assign n25869 = ( ~x619 & x1159 ) | ( ~x619 & n25866 ) | ( x1159 & n25866 ) ;
  assign n25870 = n25868 & n25869 ;
  assign n25871 = ( x619 & x1159 ) | ( x619 & ~n25770 ) | ( x1159 & ~n25770 ) ;
  assign n25872 = ( x619 & ~x1159 ) | ( x619 & n25866 ) | ( ~x1159 & n25866 ) ;
  assign n25873 = ~n25871 & n25872 ;
  assign n25874 = n25870 | n25873 ;
  assign n25875 = x789 & n25874 ;
  assign n25876 = n25867 | n25875 ;
  assign n25877 = n16176 | n25876 ;
  assign n25878 = n16176 & ~n25770 ;
  assign n25879 = n25877 & ~n25878 ;
  assign n25880 = n15134 | n25879 ;
  assign n25881 = n15134 & ~n25770 ;
  assign n25882 = n25880 & ~n25881 ;
  assign n25883 = n15141 | n25882 ;
  assign n25884 = n15141 & ~n25770 ;
  assign n25885 = n25883 & ~n25884 ;
  assign n25886 = ( x644 & x715 ) | ( x644 & ~n25885 ) | ( x715 & ~n25885 ) ;
  assign n25887 = ( x644 & ~x715 ) | ( x644 & n25770 ) | ( ~x715 & n25770 ) ;
  assign n25888 = ~n25886 & n25887 ;
  assign n25889 = x1160 & ~n25888 ;
  assign n25890 = ~n25827 & n25889 ;
  assign n25891 = x644 & ~n25825 ;
  assign n25892 = x715 | n25891 ;
  assign n25893 = ( x644 & x715 ) | ( x644 & n25885 ) | ( x715 & n25885 ) ;
  assign n25894 = ( ~x644 & x715 ) | ( ~x644 & n25770 ) | ( x715 & n25770 ) ;
  assign n25895 = n25893 & n25894 ;
  assign n25896 = x1160 | n25895 ;
  assign n25897 = n25892 & ~n25896 ;
  assign n25898 = n25890 | n25897 ;
  assign n25899 = x790 & n25898 ;
  assign n25900 = n18621 & n25879 ;
  assign n25901 = ( x629 & n25811 ) | ( x629 & n25900 ) | ( n25811 & n25900 ) ;
  assign n25902 = ( ~x629 & n25808 ) | ( ~x629 & n25900 ) | ( n25808 & n25900 ) ;
  assign n25903 = n25901 | n25902 ;
  assign n25904 = x792 & n25903 ;
  assign n25905 = x648 & ~n25873 ;
  assign n25906 = ( x619 & x1159 ) | ( x619 & n25799 ) | ( x1159 & n25799 ) ;
  assign n25907 = x627 | n25860 ;
  assign n25908 = ( x618 & x1154 ) | ( x618 & ~n25796 ) | ( x1154 & ~n25796 ) ;
  assign n25909 = x660 | n25849 ;
  assign n25910 = ( x609 & x1155 ) | ( x609 & ~n25793 ) | ( x1155 & ~n25793 ) ;
  assign n25911 = x608 | n25787 ;
  assign n25912 = ( x625 & x1153 ) | ( x625 & ~n25841 ) | ( x1153 & ~n25841 ) ;
  assign n25913 = x737 & ~n25839 ;
  assign n25914 = ( x184 & ~x777 ) | ( x184 & n15797 ) | ( ~x777 & n15797 ) ;
  assign n25915 = ( x184 & x777 ) | ( x184 & n15872 ) | ( x777 & n15872 ) ;
  assign n25916 = n25914 & ~n25915 ;
  assign n25917 = x39 & ~n25916 ;
  assign n25918 = ( x184 & ~x777 ) | ( x184 & n15583 ) | ( ~x777 & n15583 ) ;
  assign n25919 = ( x184 & x777 ) | ( x184 & n15699 ) | ( x777 & n15699 ) ;
  assign n25920 = ~n25918 & n25919 ;
  assign n25921 = n25917 & ~n25920 ;
  assign n25922 = ( ~x184 & x777 ) | ( ~x184 & n15887 ) | ( x777 & n15887 ) ;
  assign n25923 = ( x184 & x777 ) | ( x184 & ~n15891 ) | ( x777 & ~n15891 ) ;
  assign n25924 = n25922 & n25923 ;
  assign n25925 = ( ~x184 & x777 ) | ( ~x184 & n15894 ) | ( x777 & n15894 ) ;
  assign n25926 = ( x184 & x777 ) | ( x184 & ~n15897 ) | ( x777 & ~n15897 ) ;
  assign n25927 = n25925 | n25926 ;
  assign n25928 = ~n25924 & n25927 ;
  assign n25929 = x39 | n25928 ;
  assign n25930 = ~x38 & n25929 ;
  assign n25931 = ~n25921 & n25930 ;
  assign n25932 = x777 | n15758 ;
  assign n25933 = n17573 & n25932 ;
  assign n25934 = x184 | n25933 ;
  assign n25935 = n15529 | n25598 ;
  assign n25936 = x184 & n25935 ;
  assign n25937 = ~n4810 & n25936 ;
  assign n25938 = x38 & ~n25937 ;
  assign n25939 = n25934 & n25938 ;
  assign n25940 = x737 | n25939 ;
  assign n25941 = n25931 | n25940 ;
  assign n25942 = ~n2032 & n25941 ;
  assign n25943 = ~n25913 & n25942 ;
  assign n25944 = n25828 | n25943 ;
  assign n25945 = ( x625 & ~x1153 ) | ( x625 & n25944 ) | ( ~x1153 & n25944 ) ;
  assign n25946 = ~n25912 & n25945 ;
  assign n25947 = n25911 | n25946 ;
  assign n25948 = x608 & ~n25790 ;
  assign n25949 = ( x625 & x1153 ) | ( x625 & n25841 ) | ( x1153 & n25841 ) ;
  assign n25950 = ( ~x625 & x1153 ) | ( ~x625 & n25944 ) | ( x1153 & n25944 ) ;
  assign n25951 = n25949 & n25950 ;
  assign n25952 = n25948 & ~n25951 ;
  assign n25953 = n25947 & ~n25952 ;
  assign n25954 = x778 & ~n25953 ;
  assign n25955 = x778 | n25944 ;
  assign n25956 = ~n25954 & n25955 ;
  assign n25957 = ( x609 & ~x1155 ) | ( x609 & n25956 ) | ( ~x1155 & n25956 ) ;
  assign n25958 = ~n25910 & n25957 ;
  assign n25959 = n25909 | n25958 ;
  assign n25960 = x660 & ~n25853 ;
  assign n25961 = ( x609 & x1155 ) | ( x609 & n25793 ) | ( x1155 & n25793 ) ;
  assign n25962 = ( ~x609 & x1155 ) | ( ~x609 & n25956 ) | ( x1155 & n25956 ) ;
  assign n25963 = n25961 & n25962 ;
  assign n25964 = n25960 & ~n25963 ;
  assign n25965 = n25959 & ~n25964 ;
  assign n25966 = x785 & ~n25965 ;
  assign n25967 = x785 | n25956 ;
  assign n25968 = ~n25966 & n25967 ;
  assign n25969 = ( x618 & ~x1154 ) | ( x618 & n25968 ) | ( ~x1154 & n25968 ) ;
  assign n25970 = ~n25908 & n25969 ;
  assign n25971 = n25907 | n25970 ;
  assign n25972 = x627 & ~n25863 ;
  assign n25973 = ( x618 & x1154 ) | ( x618 & n25796 ) | ( x1154 & n25796 ) ;
  assign n25974 = ( ~x618 & x1154 ) | ( ~x618 & n25968 ) | ( x1154 & n25968 ) ;
  assign n25975 = n25973 & n25974 ;
  assign n25976 = n25972 & ~n25975 ;
  assign n25977 = n25971 & ~n25976 ;
  assign n25978 = x781 & ~n25977 ;
  assign n25979 = x781 | n25968 ;
  assign n25980 = ~n25978 & n25979 ;
  assign n25981 = ( ~x619 & x1159 ) | ( ~x619 & n25980 ) | ( x1159 & n25980 ) ;
  assign n25982 = n25906 & n25981 ;
  assign n25983 = n25905 & ~n25982 ;
  assign n25984 = x648 | n25870 ;
  assign n25985 = ( x619 & x1159 ) | ( x619 & ~n25799 ) | ( x1159 & ~n25799 ) ;
  assign n25986 = ( x619 & ~x1159 ) | ( x619 & n25980 ) | ( ~x1159 & n25980 ) ;
  assign n25987 = ~n25985 & n25986 ;
  assign n25988 = n25984 | n25987 ;
  assign n25989 = x789 & n25988 ;
  assign n25990 = ~n25983 & n25989 ;
  assign n25991 = ~x789 & n25980 ;
  assign n25992 = n16177 | n25991 ;
  assign n25993 = n25990 | n25992 ;
  assign n25994 = n16115 & ~n25801 ;
  assign n25995 = ( x626 & ~n15419 ) | ( x626 & n25770 ) | ( ~n15419 & n25770 ) ;
  assign n25996 = ( x626 & n15419 ) | ( x626 & ~n25876 ) | ( n15419 & ~n25876 ) ;
  assign n25997 = ~n25995 & n25996 ;
  assign n25998 = n25994 | n25997 ;
  assign n25999 = ( x626 & n15418 ) | ( x626 & ~n25770 ) | ( n15418 & ~n25770 ) ;
  assign n26000 = ( x626 & ~n15418 ) | ( x626 & n25876 ) | ( ~n15418 & n25876 ) ;
  assign n26001 = n25999 & ~n26000 ;
  assign n26002 = n25998 | n26001 ;
  assign n26003 = x788 & n26002 ;
  assign n26004 = n18434 | n26003 ;
  assign n26005 = n25993 & ~n26004 ;
  assign n26006 = n25904 | n26005 ;
  assign n26007 = ~n18431 & n26006 ;
  assign n26008 = n18610 & n25882 ;
  assign n26009 = n15139 & n25822 ;
  assign n26010 = n15138 & n25818 ;
  assign n26011 = n26009 | n26010 ;
  assign n26012 = n26008 | n26011 ;
  assign n26013 = x787 & n26012 ;
  assign n26014 = n26007 | n26013 ;
  assign n26015 = ( x644 & ~x790 ) | ( x644 & n25889 ) | ( ~x790 & n25889 ) ;
  assign n26016 = ( x644 & x790 ) | ( x644 & n25896 ) | ( x790 & n25896 ) ;
  assign n26017 = ~n26015 & n26016 ;
  assign n26018 = n26014 | n26017 ;
  assign n26019 = ~n25899 & n26018 ;
  assign n26020 = ( ~x832 & n6785 ) | ( ~x832 & n26019 ) | ( n6785 & n26019 ) ;
  assign n26021 = ( ~x184 & x832 ) | ( ~x184 & n6785 ) | ( x832 & n6785 ) ;
  assign n26022 = n26020 & ~n26021 ;
  assign n26023 = n25769 | n26022 ;
  assign n26024 = x185 | n1290 ;
  assign n26025 = ~x751 & n14840 ;
  assign n26026 = n26024 & ~n26025 ;
  assign n26027 = n16060 | n26026 ;
  assign n26028 = ~x785 & n26027 ;
  assign n26029 = ~n15094 & n26025 ;
  assign n26030 = n26027 | n26029 ;
  assign n26031 = x1155 & n26030 ;
  assign n26032 = ~x1155 & n26024 ;
  assign n26033 = ~n26029 & n26032 ;
  assign n26034 = n26031 | n26033 ;
  assign n26035 = x785 & n26034 ;
  assign n26036 = n26028 | n26035 ;
  assign n26037 = ~x781 & n26036 ;
  assign n26038 = n16075 | n26036 ;
  assign n26039 = x1154 & n26038 ;
  assign n26040 = n16078 | n26036 ;
  assign n26041 = ~x1154 & n26040 ;
  assign n26042 = n26039 | n26041 ;
  assign n26043 = x781 & n26042 ;
  assign n26044 = n26037 | n26043 ;
  assign n26045 = ~x789 & n26044 ;
  assign n26046 = n20948 | n26044 ;
  assign n26047 = x1159 & n26046 ;
  assign n26048 = n20951 | n26044 ;
  assign n26049 = ~x1159 & n26048 ;
  assign n26050 = n26047 | n26049 ;
  assign n26051 = x789 & n26050 ;
  assign n26052 = n26045 | n26051 ;
  assign n26053 = n16176 | n26052 ;
  assign n26054 = n16176 & ~n26024 ;
  assign n26055 = n26053 & ~n26054 ;
  assign n26056 = n15134 | n26055 ;
  assign n26057 = n15134 & ~n26024 ;
  assign n26058 = n26056 & ~n26057 ;
  assign n26059 = n18610 & n26058 ;
  assign n26060 = ( x647 & x1157 ) | ( x647 & ~n26024 ) | ( x1157 & ~n26024 ) ;
  assign n26061 = ~x701 & n15202 ;
  assign n26062 = n26024 & ~n26061 ;
  assign n26063 = x778 | n26062 ;
  assign n26064 = ~x625 & n26061 ;
  assign n26065 = n26062 | n26064 ;
  assign n26066 = x1153 & n26065 ;
  assign n26067 = ~x1153 & n26024 ;
  assign n26068 = ~n26064 & n26067 ;
  assign n26069 = x778 & ~n26068 ;
  assign n26070 = ~n26066 & n26069 ;
  assign n26071 = n26063 & ~n26070 ;
  assign n26072 = n16043 | n26071 ;
  assign n26073 = n16045 | n26072 ;
  assign n26074 = n16047 | n26073 ;
  assign n26075 = n16049 | n26074 ;
  assign n26076 = n16055 | n26075 ;
  assign n26077 = ( x647 & ~x1157 ) | ( x647 & n26076 ) | ( ~x1157 & n26076 ) ;
  assign n26078 = ~n26060 & n26077 ;
  assign n26079 = x630 & n26078 ;
  assign n26080 = x647 & n26076 ;
  assign n26081 = ~x647 & n26024 ;
  assign n26082 = n26080 | n26081 ;
  assign n26083 = n15138 & n26082 ;
  assign n26084 = n26079 | n26083 ;
  assign n26085 = n26059 | n26084 ;
  assign n26086 = x787 & n26085 ;
  assign n26087 = n16115 & ~n26074 ;
  assign n26088 = ( x626 & ~n15419 ) | ( x626 & n26024 ) | ( ~n15419 & n26024 ) ;
  assign n26089 = ( x626 & n15419 ) | ( x626 & ~n26052 ) | ( n15419 & ~n26052 ) ;
  assign n26090 = ~n26088 & n26089 ;
  assign n26091 = n26087 | n26090 ;
  assign n26092 = ( x626 & n15418 ) | ( x626 & ~n26024 ) | ( n15418 & ~n26024 ) ;
  assign n26093 = ( x626 & ~n15418 ) | ( x626 & n26052 ) | ( ~n15418 & n26052 ) ;
  assign n26094 = n26092 & ~n26093 ;
  assign n26095 = n26091 | n26094 ;
  assign n26096 = x788 & n26095 ;
  assign n26097 = x648 & ~n26049 ;
  assign n26098 = ( x619 & x1159 ) | ( x619 & n26073 ) | ( x1159 & n26073 ) ;
  assign n26099 = x627 | n26039 ;
  assign n26100 = ( x618 & x1154 ) | ( x618 & ~n26072 ) | ( x1154 & ~n26072 ) ;
  assign n26101 = x660 | n26031 ;
  assign n26102 = ( x609 & x1155 ) | ( x609 & ~n26071 ) | ( x1155 & ~n26071 ) ;
  assign n26103 = n14839 | n26062 ;
  assign n26104 = x625 & ~n26103 ;
  assign n26105 = n26026 & n26103 ;
  assign n26106 = n26104 | n26105 ;
  assign n26107 = n26067 & n26106 ;
  assign n26108 = x608 | n26066 ;
  assign n26109 = n26107 | n26108 ;
  assign n26110 = x1153 & n26026 ;
  assign n26111 = ~n26104 & n26110 ;
  assign n26112 = x608 & ~n26068 ;
  assign n26113 = ~n26111 & n26112 ;
  assign n26114 = n26109 & ~n26113 ;
  assign n26115 = x778 & ~n26114 ;
  assign n26116 = x778 | n26105 ;
  assign n26117 = ~n26115 & n26116 ;
  assign n26118 = ( x609 & ~x1155 ) | ( x609 & n26117 ) | ( ~x1155 & n26117 ) ;
  assign n26119 = ~n26102 & n26118 ;
  assign n26120 = n26101 | n26119 ;
  assign n26121 = x660 & ~n26033 ;
  assign n26122 = ( x609 & x1155 ) | ( x609 & n26071 ) | ( x1155 & n26071 ) ;
  assign n26123 = ( ~x609 & x1155 ) | ( ~x609 & n26117 ) | ( x1155 & n26117 ) ;
  assign n26124 = n26122 & n26123 ;
  assign n26125 = n26121 & ~n26124 ;
  assign n26126 = n26120 & ~n26125 ;
  assign n26127 = x785 & ~n26126 ;
  assign n26128 = x785 | n26117 ;
  assign n26129 = ~n26127 & n26128 ;
  assign n26130 = ( x618 & ~x1154 ) | ( x618 & n26129 ) | ( ~x1154 & n26129 ) ;
  assign n26131 = ~n26100 & n26130 ;
  assign n26132 = n26099 | n26131 ;
  assign n26133 = x627 & ~n26041 ;
  assign n26134 = ( x618 & x1154 ) | ( x618 & n26072 ) | ( x1154 & n26072 ) ;
  assign n26135 = ( ~x618 & x1154 ) | ( ~x618 & n26129 ) | ( x1154 & n26129 ) ;
  assign n26136 = n26134 & n26135 ;
  assign n26137 = n26133 & ~n26136 ;
  assign n26138 = n26132 & ~n26137 ;
  assign n26139 = x781 & ~n26138 ;
  assign n26140 = x781 | n26129 ;
  assign n26141 = ~n26139 & n26140 ;
  assign n26142 = ( ~x619 & x1159 ) | ( ~x619 & n26141 ) | ( x1159 & n26141 ) ;
  assign n26143 = n26098 & n26142 ;
  assign n26144 = n26097 & ~n26143 ;
  assign n26145 = x648 | n26047 ;
  assign n26146 = ( x619 & x1159 ) | ( x619 & ~n26073 ) | ( x1159 & ~n26073 ) ;
  assign n26147 = ( x619 & ~x1159 ) | ( x619 & n26141 ) | ( ~x1159 & n26141 ) ;
  assign n26148 = ~n26146 & n26147 ;
  assign n26149 = n26145 | n26148 ;
  assign n26150 = x789 & n26149 ;
  assign n26151 = ~n26144 & n26150 ;
  assign n26152 = ~x789 & n26141 ;
  assign n26153 = n16177 | n26152 ;
  assign n26154 = n26151 | n26153 ;
  assign n26155 = ~n26096 & n26154 ;
  assign n26156 = n18434 | n26155 ;
  assign n26157 = n16650 | n26075 ;
  assign n26158 = n16051 & ~n26055 ;
  assign n26159 = n26157 & ~n26158 ;
  assign n26160 = ( x629 & ~x792 ) | ( x629 & n26159 ) | ( ~x792 & n26159 ) ;
  assign n26161 = n16052 & ~n26055 ;
  assign n26162 = n16643 & ~n26075 ;
  assign n26163 = n26161 | n26162 ;
  assign n26164 = ( x629 & x792 ) | ( x629 & n26163 ) | ( x792 & n26163 ) ;
  assign n26165 = ~n26160 & n26164 ;
  assign n26166 = n18431 | n26165 ;
  assign n26167 = n26156 & ~n26166 ;
  assign n26168 = n26086 | n26167 ;
  assign n26169 = ( x790 & x832 ) | ( x790 & n26168 ) | ( x832 & n26168 ) ;
  assign n26170 = n15141 | n26058 ;
  assign n26171 = n15141 & ~n26024 ;
  assign n26172 = n26170 & ~n26171 ;
  assign n26173 = ( x644 & x715 ) | ( x644 & ~n26172 ) | ( x715 & ~n26172 ) ;
  assign n26174 = ( x644 & ~x715 ) | ( x644 & n26024 ) | ( ~x715 & n26024 ) ;
  assign n26175 = ~n26173 & n26174 ;
  assign n26176 = x1160 & ~n26175 ;
  assign n26177 = ~x787 & n26076 ;
  assign n26178 = x1157 & n26082 ;
  assign n26179 = n26078 | n26178 ;
  assign n26180 = x787 & n26179 ;
  assign n26181 = n26177 | n26180 ;
  assign n26182 = ( x644 & x715 ) | ( x644 & n26181 ) | ( x715 & n26181 ) ;
  assign n26183 = ( ~x644 & x715 ) | ( ~x644 & n26168 ) | ( x715 & n26168 ) ;
  assign n26184 = n26182 & n26183 ;
  assign n26185 = n26176 & ~n26184 ;
  assign n26186 = ( x644 & x715 ) | ( x644 & n26172 ) | ( x715 & n26172 ) ;
  assign n26187 = ( ~x644 & x715 ) | ( ~x644 & n26024 ) | ( x715 & n26024 ) ;
  assign n26188 = n26186 & n26187 ;
  assign n26189 = x1160 | n26188 ;
  assign n26190 = ( x644 & x715 ) | ( x644 & ~n26181 ) | ( x715 & ~n26181 ) ;
  assign n26191 = ( x644 & ~x715 ) | ( x644 & n26168 ) | ( ~x715 & n26168 ) ;
  assign n26192 = ~n26190 & n26191 ;
  assign n26193 = n26189 | n26192 ;
  assign n26194 = ~n26185 & n26193 ;
  assign n26195 = ( ~x790 & x832 ) | ( ~x790 & n26194 ) | ( x832 & n26194 ) ;
  assign n26196 = n26169 & n26195 ;
  assign n26197 = x185 | n14834 ;
  assign n26198 = n15414 & n26197 ;
  assign n26199 = x701 | n2032 ;
  assign n26200 = ~n26197 & n26199 ;
  assign n26201 = x185 & n16323 ;
  assign n26202 = x38 | n26201 ;
  assign n26203 = ~n2032 & n26202 ;
  assign n26204 = x185 | n16319 ;
  assign n26205 = ~n26203 & n26204 ;
  assign n26206 = x185 | n15070 ;
  assign n26207 = n15375 & n26206 ;
  assign n26208 = x701 | n26207 ;
  assign n26209 = n26205 | n26208 ;
  assign n26210 = ~n26200 & n26209 ;
  assign n26211 = ~x778 & n26210 ;
  assign n26212 = ( x625 & x1153 ) | ( x625 & n26197 ) | ( x1153 & n26197 ) ;
  assign n26213 = ( ~x625 & x1153 ) | ( ~x625 & n26210 ) | ( x1153 & n26210 ) ;
  assign n26214 = n26212 & n26213 ;
  assign n26215 = ( x625 & x1153 ) | ( x625 & ~n26197 ) | ( x1153 & ~n26197 ) ;
  assign n26216 = ( x625 & ~x1153 ) | ( x625 & n26210 ) | ( ~x1153 & n26210 ) ;
  assign n26217 = ~n26215 & n26216 ;
  assign n26218 = n26214 | n26217 ;
  assign n26219 = x778 & n26218 ;
  assign n26220 = n26211 | n26219 ;
  assign n26221 = ~n15400 & n26220 ;
  assign n26222 = n15400 & n26197 ;
  assign n26223 = n26221 | n26222 ;
  assign n26224 = n15407 | n26223 ;
  assign n26225 = n15407 & ~n26197 ;
  assign n26226 = n26224 & ~n26225 ;
  assign n26227 = ~n15414 & n26226 ;
  assign n26228 = n26198 | n26227 ;
  assign n26229 = n15421 | n26228 ;
  assign n26230 = n15421 & ~n26197 ;
  assign n26231 = n26229 & ~n26230 ;
  assign n26232 = ~x792 & n26231 ;
  assign n26233 = ( x628 & x1156 ) | ( x628 & n26197 ) | ( x1156 & n26197 ) ;
  assign n26234 = ( ~x628 & x1156 ) | ( ~x628 & n26231 ) | ( x1156 & n26231 ) ;
  assign n26235 = n26233 & n26234 ;
  assign n26236 = ( x628 & x1156 ) | ( x628 & ~n26197 ) | ( x1156 & ~n26197 ) ;
  assign n26237 = ( x628 & ~x1156 ) | ( x628 & n26231 ) | ( ~x1156 & n26231 ) ;
  assign n26238 = ~n26236 & n26237 ;
  assign n26239 = n26235 | n26238 ;
  assign n26240 = x792 & n26239 ;
  assign n26241 = n26232 | n26240 ;
  assign n26242 = x787 | n26241 ;
  assign n26243 = x647 & n26241 ;
  assign n26244 = ~x647 & n26197 ;
  assign n26245 = n26243 | n26244 ;
  assign n26246 = ( ~x787 & x1157 ) | ( ~x787 & n26245 ) | ( x1157 & n26245 ) ;
  assign n26247 = ~x647 & n26241 ;
  assign n26248 = x647 & n26197 ;
  assign n26249 = n26247 | n26248 ;
  assign n26250 = ( x787 & x1157 ) | ( x787 & ~n26249 ) | ( x1157 & ~n26249 ) ;
  assign n26251 = ~n26246 & n26250 ;
  assign n26252 = n26242 & ~n26251 ;
  assign n26253 = x644 | n26252 ;
  assign n26254 = x715 & n26253 ;
  assign n26255 = x185 & n2032 ;
  assign n26256 = x751 & n14710 ;
  assign n26257 = x185 & ~n14907 ;
  assign n26258 = n26256 | n26257 ;
  assign n26259 = x39 & n26258 ;
  assign n26260 = x185 & ~x751 ;
  assign n26261 = x185 & ~n15896 ;
  assign n26262 = n19258 | n26261 ;
  assign n26263 = ~x39 & n26262 ;
  assign n26264 = ( ~x751 & n15063 ) | ( ~x751 & n26260 ) | ( n15063 & n26260 ) ;
  assign n26265 = ( ~n26260 & n26263 ) | ( ~n26260 & n26264 ) | ( n26263 & n26264 ) ;
  assign n26266 = ( x185 & ~n26260 ) | ( x185 & n26265 ) | ( ~n26260 & n26265 ) ;
  assign n26267 = n26259 | n26266 ;
  assign n26268 = ~x38 & n26267 ;
  assign n26269 = ~x751 & n15072 ;
  assign n26270 = x38 & n26206 ;
  assign n26271 = ~n26269 & n26270 ;
  assign n26272 = n26268 | n26271 ;
  assign n26273 = ~n2032 & n26272 ;
  assign n26274 = n26255 | n26273 ;
  assign n26275 = ~n15082 & n26274 ;
  assign n26276 = n15082 & n26197 ;
  assign n26277 = n26275 | n26276 ;
  assign n26278 = ~x785 & n26277 ;
  assign n26279 = ~n15088 & n26197 ;
  assign n26280 = x609 & n26275 ;
  assign n26281 = n26279 | n26280 ;
  assign n26282 = x1155 & n26281 ;
  assign n26283 = n15094 & n26197 ;
  assign n26284 = ~x609 & n26275 ;
  assign n26285 = n26283 | n26284 ;
  assign n26286 = ~x1155 & n26285 ;
  assign n26287 = n26282 | n26286 ;
  assign n26288 = x785 & n26287 ;
  assign n26289 = n26278 | n26288 ;
  assign n26290 = ~x781 & n26289 ;
  assign n26291 = ( x618 & x1154 ) | ( x618 & n26197 ) | ( x1154 & n26197 ) ;
  assign n26292 = ( ~x618 & x1154 ) | ( ~x618 & n26289 ) | ( x1154 & n26289 ) ;
  assign n26293 = n26291 & n26292 ;
  assign n26294 = ( x618 & x1154 ) | ( x618 & ~n26197 ) | ( x1154 & ~n26197 ) ;
  assign n26295 = ( x618 & ~x1154 ) | ( x618 & n26289 ) | ( ~x1154 & n26289 ) ;
  assign n26296 = ~n26294 & n26295 ;
  assign n26297 = n26293 | n26296 ;
  assign n26298 = x781 & n26297 ;
  assign n26299 = n26290 | n26298 ;
  assign n26300 = ~x789 & n26299 ;
  assign n26301 = ( x619 & x1159 ) | ( x619 & n26197 ) | ( x1159 & n26197 ) ;
  assign n26302 = ( ~x619 & x1159 ) | ( ~x619 & n26299 ) | ( x1159 & n26299 ) ;
  assign n26303 = n26301 & n26302 ;
  assign n26304 = ( x619 & x1159 ) | ( x619 & ~n26197 ) | ( x1159 & ~n26197 ) ;
  assign n26305 = ( x619 & ~x1159 ) | ( x619 & n26299 ) | ( ~x1159 & n26299 ) ;
  assign n26306 = ~n26304 & n26305 ;
  assign n26307 = n26303 | n26306 ;
  assign n26308 = x789 & n26307 ;
  assign n26309 = n26300 | n26308 ;
  assign n26310 = n16176 | n26309 ;
  assign n26311 = n16176 & ~n26197 ;
  assign n26312 = n26310 & ~n26311 ;
  assign n26313 = n15134 | n26312 ;
  assign n26314 = n15134 & ~n26197 ;
  assign n26315 = n26313 & ~n26314 ;
  assign n26316 = n15141 | n26315 ;
  assign n26317 = n15141 & ~n26197 ;
  assign n26318 = n26316 & ~n26317 ;
  assign n26319 = ( x644 & x715 ) | ( x644 & ~n26318 ) | ( x715 & ~n26318 ) ;
  assign n26320 = ( x644 & ~x715 ) | ( x644 & n26197 ) | ( ~x715 & n26197 ) ;
  assign n26321 = ~n26319 & n26320 ;
  assign n26322 = x1160 & ~n26321 ;
  assign n26323 = ~n26254 & n26322 ;
  assign n26324 = x644 & ~n26252 ;
  assign n26325 = x715 | n26324 ;
  assign n26326 = ( x644 & x715 ) | ( x644 & n26318 ) | ( x715 & n26318 ) ;
  assign n26327 = ( ~x644 & x715 ) | ( ~x644 & n26197 ) | ( x715 & n26197 ) ;
  assign n26328 = n26326 & n26327 ;
  assign n26329 = x1160 | n26328 ;
  assign n26330 = n26325 & ~n26329 ;
  assign n26331 = n26323 | n26330 ;
  assign n26332 = x790 & n26331 ;
  assign n26333 = n18621 & n26312 ;
  assign n26334 = ( x629 & n26238 ) | ( x629 & n26333 ) | ( n26238 & n26333 ) ;
  assign n26335 = ( ~x629 & n26235 ) | ( ~x629 & n26333 ) | ( n26235 & n26333 ) ;
  assign n26336 = n26334 | n26335 ;
  assign n26337 = x792 & n26336 ;
  assign n26338 = x648 & ~n26306 ;
  assign n26339 = ( x619 & x1159 ) | ( x619 & n26226 ) | ( x1159 & n26226 ) ;
  assign n26340 = x627 | n26293 ;
  assign n26341 = ( x618 & x1154 ) | ( x618 & ~n26223 ) | ( x1154 & ~n26223 ) ;
  assign n26342 = x660 | n26282 ;
  assign n26343 = ( x609 & x1155 ) | ( x609 & ~n26220 ) | ( x1155 & ~n26220 ) ;
  assign n26344 = x608 | n26214 ;
  assign n26345 = ( x625 & x1153 ) | ( x625 & ~n26274 ) | ( x1153 & ~n26274 ) ;
  assign n26346 = x701 & ~n26272 ;
  assign n26347 = ( x185 & ~x751 ) | ( x185 & n15797 ) | ( ~x751 & n15797 ) ;
  assign n26348 = ( x185 & x751 ) | ( x185 & n15872 ) | ( x751 & n15872 ) ;
  assign n26349 = n26347 & ~n26348 ;
  assign n26350 = x39 & ~n26349 ;
  assign n26351 = ( x185 & ~x751 ) | ( x185 & n15583 ) | ( ~x751 & n15583 ) ;
  assign n26352 = ( x185 & x751 ) | ( x185 & n15699 ) | ( x751 & n15699 ) ;
  assign n26353 = ~n26351 & n26352 ;
  assign n26354 = n26350 & ~n26353 ;
  assign n26355 = ( ~x185 & x751 ) | ( ~x185 & n15887 ) | ( x751 & n15887 ) ;
  assign n26356 = ( x185 & x751 ) | ( x185 & ~n15891 ) | ( x751 & ~n15891 ) ;
  assign n26357 = n26355 & n26356 ;
  assign n26358 = ( ~x185 & x751 ) | ( ~x185 & n15894 ) | ( x751 & n15894 ) ;
  assign n26359 = ( x185 & x751 ) | ( x185 & ~n15897 ) | ( x751 & ~n15897 ) ;
  assign n26360 = n26358 | n26359 ;
  assign n26361 = ~n26357 & n26360 ;
  assign n26362 = x39 | n26361 ;
  assign n26363 = ~x38 & n26362 ;
  assign n26364 = ~n26354 & n26363 ;
  assign n26365 = x751 | n15758 ;
  assign n26366 = n17573 & n26365 ;
  assign n26367 = x185 | n26366 ;
  assign n26368 = n15529 | n26025 ;
  assign n26369 = x185 & n26368 ;
  assign n26370 = ~n4810 & n26369 ;
  assign n26371 = x38 & ~n26370 ;
  assign n26372 = n26367 & n26371 ;
  assign n26373 = x701 | n26372 ;
  assign n26374 = n26364 | n26373 ;
  assign n26375 = ~n2032 & n26374 ;
  assign n26376 = ~n26346 & n26375 ;
  assign n26377 = n26255 | n26376 ;
  assign n26378 = ( x625 & ~x1153 ) | ( x625 & n26377 ) | ( ~x1153 & n26377 ) ;
  assign n26379 = ~n26345 & n26378 ;
  assign n26380 = n26344 | n26379 ;
  assign n26381 = x608 & ~n26217 ;
  assign n26382 = ( x625 & x1153 ) | ( x625 & n26274 ) | ( x1153 & n26274 ) ;
  assign n26383 = ( ~x625 & x1153 ) | ( ~x625 & n26377 ) | ( x1153 & n26377 ) ;
  assign n26384 = n26382 & n26383 ;
  assign n26385 = n26381 & ~n26384 ;
  assign n26386 = n26380 & ~n26385 ;
  assign n26387 = x778 & ~n26386 ;
  assign n26388 = x778 | n26377 ;
  assign n26389 = ~n26387 & n26388 ;
  assign n26390 = ( x609 & ~x1155 ) | ( x609 & n26389 ) | ( ~x1155 & n26389 ) ;
  assign n26391 = ~n26343 & n26390 ;
  assign n26392 = n26342 | n26391 ;
  assign n26393 = x660 & ~n26286 ;
  assign n26394 = ( x609 & x1155 ) | ( x609 & n26220 ) | ( x1155 & n26220 ) ;
  assign n26395 = ( ~x609 & x1155 ) | ( ~x609 & n26389 ) | ( x1155 & n26389 ) ;
  assign n26396 = n26394 & n26395 ;
  assign n26397 = n26393 & ~n26396 ;
  assign n26398 = n26392 & ~n26397 ;
  assign n26399 = x785 & ~n26398 ;
  assign n26400 = x785 | n26389 ;
  assign n26401 = ~n26399 & n26400 ;
  assign n26402 = ( x618 & ~x1154 ) | ( x618 & n26401 ) | ( ~x1154 & n26401 ) ;
  assign n26403 = ~n26341 & n26402 ;
  assign n26404 = n26340 | n26403 ;
  assign n26405 = x627 & ~n26296 ;
  assign n26406 = ( x618 & x1154 ) | ( x618 & n26223 ) | ( x1154 & n26223 ) ;
  assign n26407 = ( ~x618 & x1154 ) | ( ~x618 & n26401 ) | ( x1154 & n26401 ) ;
  assign n26408 = n26406 & n26407 ;
  assign n26409 = n26405 & ~n26408 ;
  assign n26410 = n26404 & ~n26409 ;
  assign n26411 = x781 & ~n26410 ;
  assign n26412 = x781 | n26401 ;
  assign n26413 = ~n26411 & n26412 ;
  assign n26414 = ( ~x619 & x1159 ) | ( ~x619 & n26413 ) | ( x1159 & n26413 ) ;
  assign n26415 = n26339 & n26414 ;
  assign n26416 = n26338 & ~n26415 ;
  assign n26417 = x648 | n26303 ;
  assign n26418 = ( x619 & x1159 ) | ( x619 & ~n26226 ) | ( x1159 & ~n26226 ) ;
  assign n26419 = ( x619 & ~x1159 ) | ( x619 & n26413 ) | ( ~x1159 & n26413 ) ;
  assign n26420 = ~n26418 & n26419 ;
  assign n26421 = n26417 | n26420 ;
  assign n26422 = x789 & n26421 ;
  assign n26423 = ~n26416 & n26422 ;
  assign n26424 = ~x789 & n26413 ;
  assign n26425 = n16177 | n26424 ;
  assign n26426 = n26423 | n26425 ;
  assign n26427 = n16115 & ~n26228 ;
  assign n26428 = ( x626 & ~n15419 ) | ( x626 & n26197 ) | ( ~n15419 & n26197 ) ;
  assign n26429 = ( x626 & n15419 ) | ( x626 & ~n26309 ) | ( n15419 & ~n26309 ) ;
  assign n26430 = ~n26428 & n26429 ;
  assign n26431 = n26427 | n26430 ;
  assign n26432 = ( x626 & n15418 ) | ( x626 & ~n26197 ) | ( n15418 & ~n26197 ) ;
  assign n26433 = ( x626 & ~n15418 ) | ( x626 & n26309 ) | ( ~n15418 & n26309 ) ;
  assign n26434 = n26432 & ~n26433 ;
  assign n26435 = n26431 | n26434 ;
  assign n26436 = x788 & n26435 ;
  assign n26437 = n18434 | n26436 ;
  assign n26438 = n26426 & ~n26437 ;
  assign n26439 = n26337 | n26438 ;
  assign n26440 = ~n18431 & n26439 ;
  assign n26441 = n18610 & n26315 ;
  assign n26442 = n15139 & n26249 ;
  assign n26443 = n15138 & n26245 ;
  assign n26444 = n26442 | n26443 ;
  assign n26445 = n26441 | n26444 ;
  assign n26446 = x787 & n26445 ;
  assign n26447 = n26440 | n26446 ;
  assign n26448 = ( x644 & ~x790 ) | ( x644 & n26322 ) | ( ~x790 & n26322 ) ;
  assign n26449 = ( x644 & x790 ) | ( x644 & n26329 ) | ( x790 & n26329 ) ;
  assign n26450 = ~n26448 & n26449 ;
  assign n26451 = n26447 | n26450 ;
  assign n26452 = ~n26332 & n26451 ;
  assign n26453 = ( ~x832 & n6785 ) | ( ~x832 & n26452 ) | ( n6785 & n26452 ) ;
  assign n26454 = ( ~x185 & x832 ) | ( ~x185 & n6785 ) | ( x832 & n6785 ) ;
  assign n26455 = n26453 & ~n26454 ;
  assign n26456 = n26196 | n26455 ;
  assign n26457 = x186 | n14834 ;
  assign n26458 = n15141 & n26457 ;
  assign n26459 = x186 & n2032 ;
  assign n26460 = x186 | n15382 ;
  assign n26461 = x752 & n26460 ;
  assign n26462 = x186 & ~n17416 ;
  assign n26463 = x186 | x752 ;
  assign n26464 = n17421 & ~n26463 ;
  assign n26465 = n26462 | n26464 ;
  assign n26466 = ~n17415 & n26465 ;
  assign n26467 = n26461 | n26466 ;
  assign n26468 = ~n2032 & n26467 ;
  assign n26469 = n26459 | n26468 ;
  assign n26470 = ~n15082 & n26469 ;
  assign n26471 = n15082 & n26457 ;
  assign n26472 = n26470 | n26471 ;
  assign n26473 = ~x785 & n26472 ;
  assign n26474 = ~n15088 & n26457 ;
  assign n26475 = x609 & n26470 ;
  assign n26476 = n26474 | n26475 ;
  assign n26477 = x1155 & n26476 ;
  assign n26478 = n15094 & n26457 ;
  assign n26479 = ~x609 & n26470 ;
  assign n26480 = n26478 | n26479 ;
  assign n26481 = ~x1155 & n26480 ;
  assign n26482 = n26477 | n26481 ;
  assign n26483 = x785 & n26482 ;
  assign n26484 = n26473 | n26483 ;
  assign n26485 = ~x781 & n26484 ;
  assign n26486 = ( x618 & x1154 ) | ( x618 & n26457 ) | ( x1154 & n26457 ) ;
  assign n26487 = ( ~x618 & x1154 ) | ( ~x618 & n26484 ) | ( x1154 & n26484 ) ;
  assign n26488 = n26486 & n26487 ;
  assign n26489 = ( x618 & x1154 ) | ( x618 & ~n26457 ) | ( x1154 & ~n26457 ) ;
  assign n26490 = ( x618 & ~x1154 ) | ( x618 & n26484 ) | ( ~x1154 & n26484 ) ;
  assign n26491 = ~n26489 & n26490 ;
  assign n26492 = n26488 | n26491 ;
  assign n26493 = x781 & n26492 ;
  assign n26494 = n26485 | n26493 ;
  assign n26495 = ~x789 & n26494 ;
  assign n26496 = ( x619 & x1159 ) | ( x619 & n26457 ) | ( x1159 & n26457 ) ;
  assign n26497 = ( ~x619 & x1159 ) | ( ~x619 & n26494 ) | ( x1159 & n26494 ) ;
  assign n26498 = n26496 & n26497 ;
  assign n26499 = ( x619 & x1159 ) | ( x619 & ~n26457 ) | ( x1159 & ~n26457 ) ;
  assign n26500 = ( x619 & ~x1159 ) | ( x619 & n26494 ) | ( ~x1159 & n26494 ) ;
  assign n26501 = ~n26499 & n26500 ;
  assign n26502 = n26498 | n26501 ;
  assign n26503 = x789 & n26502 ;
  assign n26504 = n26495 | n26503 ;
  assign n26505 = n16176 | n26504 ;
  assign n26506 = n16176 & ~n26457 ;
  assign n26507 = n26505 & ~n26506 ;
  assign n26508 = n15134 | n26507 ;
  assign n26509 = n15134 & ~n26457 ;
  assign n26510 = n26508 & ~n26509 ;
  assign n26511 = ~n15141 & n26510 ;
  assign n26512 = n26458 | n26511 ;
  assign n26513 = ( x644 & x715 ) | ( x644 & n26512 ) | ( x715 & n26512 ) ;
  assign n26514 = ( ~x644 & x715 ) | ( ~x644 & n26457 ) | ( x715 & n26457 ) ;
  assign n26515 = n26513 & n26514 ;
  assign n26516 = x1160 | n26515 ;
  assign n26517 = n15414 & n26457 ;
  assign n26518 = x186 | n15070 ;
  assign n26519 = n15375 & n26518 ;
  assign n26520 = x703 & ~n26519 ;
  assign n26521 = ( ~x38 & x186 ) | ( ~x38 & n16319 ) | ( x186 & n16319 ) ;
  assign n26522 = ( x38 & x186 ) | ( x38 & n16323 ) | ( x186 & n16323 ) ;
  assign n26523 = n26521 & ~n26522 ;
  assign n26524 = n26520 & ~n26523 ;
  assign n26525 = x703 | n26460 ;
  assign n26526 = ~n2032 & n26525 ;
  assign n26527 = ~n26524 & n26526 ;
  assign n26528 = n26459 | n26527 ;
  assign n26529 = ~x778 & n26528 ;
  assign n26530 = ( x625 & x1153 ) | ( x625 & n26457 ) | ( x1153 & n26457 ) ;
  assign n26531 = ( ~x625 & x1153 ) | ( ~x625 & n26528 ) | ( x1153 & n26528 ) ;
  assign n26532 = n26530 & n26531 ;
  assign n26533 = ( x625 & x1153 ) | ( x625 & ~n26457 ) | ( x1153 & ~n26457 ) ;
  assign n26534 = ( x625 & ~x1153 ) | ( x625 & n26528 ) | ( ~x1153 & n26528 ) ;
  assign n26535 = ~n26533 & n26534 ;
  assign n26536 = n26532 | n26535 ;
  assign n26537 = x778 & n26536 ;
  assign n26538 = n26529 | n26537 ;
  assign n26539 = ~n15400 & n26538 ;
  assign n26540 = n15400 & n26457 ;
  assign n26541 = n26539 | n26540 ;
  assign n26542 = n15407 | n26541 ;
  assign n26543 = n15407 & ~n26457 ;
  assign n26544 = n26542 & ~n26543 ;
  assign n26545 = ~n15414 & n26544 ;
  assign n26546 = n26517 | n26545 ;
  assign n26547 = n15421 | n26546 ;
  assign n26548 = n15421 & ~n26457 ;
  assign n26549 = n26547 & ~n26548 ;
  assign n26550 = ~x792 & n26549 ;
  assign n26551 = ( x628 & x1156 ) | ( x628 & n26457 ) | ( x1156 & n26457 ) ;
  assign n26552 = ( ~x628 & x1156 ) | ( ~x628 & n26549 ) | ( x1156 & n26549 ) ;
  assign n26553 = n26551 & n26552 ;
  assign n26554 = ( x628 & x1156 ) | ( x628 & ~n26457 ) | ( x1156 & ~n26457 ) ;
  assign n26555 = ( x628 & ~x1156 ) | ( x628 & n26549 ) | ( ~x1156 & n26549 ) ;
  assign n26556 = ~n26554 & n26555 ;
  assign n26557 = n26553 | n26556 ;
  assign n26558 = x792 & n26557 ;
  assign n26559 = n26550 | n26558 ;
  assign n26560 = ~x787 & n26559 ;
  assign n26561 = ( x647 & x1157 ) | ( x647 & n26457 ) | ( x1157 & n26457 ) ;
  assign n26562 = ( ~x647 & x1157 ) | ( ~x647 & n26559 ) | ( x1157 & n26559 ) ;
  assign n26563 = n26561 & n26562 ;
  assign n26564 = ( x647 & x1157 ) | ( x647 & ~n26457 ) | ( x1157 & ~n26457 ) ;
  assign n26565 = ( x647 & ~x1157 ) | ( x647 & n26559 ) | ( ~x1157 & n26559 ) ;
  assign n26566 = ~n26564 & n26565 ;
  assign n26567 = n26563 | n26566 ;
  assign n26568 = x787 & n26567 ;
  assign n26569 = n26560 | n26568 ;
  assign n26570 = ( x644 & x715 ) | ( x644 & ~n26569 ) | ( x715 & ~n26569 ) ;
  assign n26571 = x630 | n26563 ;
  assign n26572 = ( x647 & x1157 ) | ( x647 & ~n26510 ) | ( x1157 & ~n26510 ) ;
  assign n26573 = x629 | n26553 ;
  assign n26574 = ( x628 & x1156 ) | ( x628 & ~n26507 ) | ( x1156 & ~n26507 ) ;
  assign n26575 = x648 | n26498 ;
  assign n26576 = ( x619 & x1159 ) | ( x619 & ~n26544 ) | ( x1159 & ~n26544 ) ;
  assign n26577 = x627 | n26488 ;
  assign n26578 = ( x618 & x1154 ) | ( x618 & ~n26541 ) | ( x1154 & ~n26541 ) ;
  assign n26579 = x660 | n26477 ;
  assign n26580 = ( x609 & x1155 ) | ( x609 & ~n26538 ) | ( x1155 & ~n26538 ) ;
  assign n26581 = x608 | n26532 ;
  assign n26582 = ( x625 & x1153 ) | ( x625 & ~n26469 ) | ( x1153 & ~n26469 ) ;
  assign n26583 = x703 | n26467 ;
  assign n26584 = ( x186 & ~x752 ) | ( x186 & n17554 ) | ( ~x752 & n17554 ) ;
  assign n26585 = ( x186 & x752 ) | ( x186 & n17562 ) | ( x752 & n17562 ) ;
  assign n26586 = n26584 & ~n26585 ;
  assign n26587 = x703 & ~n26586 ;
  assign n26588 = x752 & ~n17570 ;
  assign n26589 = ( x186 & n17569 ) | ( x186 & ~n26588 ) | ( n17569 & ~n26588 ) ;
  assign n26590 = ( x186 & n17579 ) | ( x186 & n26588 ) | ( n17579 & n26588 ) ;
  assign n26591 = ~n26589 & n26590 ;
  assign n26592 = n26587 & ~n26591 ;
  assign n26593 = n2032 | n26592 ;
  assign n26594 = n26583 & ~n26593 ;
  assign n26595 = n26459 | n26594 ;
  assign n26596 = ( x625 & ~x1153 ) | ( x625 & n26595 ) | ( ~x1153 & n26595 ) ;
  assign n26597 = ~n26582 & n26596 ;
  assign n26598 = n26581 | n26597 ;
  assign n26599 = x608 & ~n26535 ;
  assign n26600 = ( x625 & x1153 ) | ( x625 & n26469 ) | ( x1153 & n26469 ) ;
  assign n26601 = ( ~x625 & x1153 ) | ( ~x625 & n26595 ) | ( x1153 & n26595 ) ;
  assign n26602 = n26600 & n26601 ;
  assign n26603 = n26599 & ~n26602 ;
  assign n26604 = n26598 & ~n26603 ;
  assign n26605 = x778 & ~n26604 ;
  assign n26606 = x778 | n26595 ;
  assign n26607 = ~n26605 & n26606 ;
  assign n26608 = ( x609 & ~x1155 ) | ( x609 & n26607 ) | ( ~x1155 & n26607 ) ;
  assign n26609 = ~n26580 & n26608 ;
  assign n26610 = n26579 | n26609 ;
  assign n26611 = x660 & ~n26481 ;
  assign n26612 = ( x609 & x1155 ) | ( x609 & n26538 ) | ( x1155 & n26538 ) ;
  assign n26613 = ( ~x609 & x1155 ) | ( ~x609 & n26607 ) | ( x1155 & n26607 ) ;
  assign n26614 = n26612 & n26613 ;
  assign n26615 = n26611 & ~n26614 ;
  assign n26616 = n26610 & ~n26615 ;
  assign n26617 = x785 & ~n26616 ;
  assign n26618 = x785 | n26607 ;
  assign n26619 = ~n26617 & n26618 ;
  assign n26620 = ( x618 & ~x1154 ) | ( x618 & n26619 ) | ( ~x1154 & n26619 ) ;
  assign n26621 = ~n26578 & n26620 ;
  assign n26622 = n26577 | n26621 ;
  assign n26623 = x627 & ~n26491 ;
  assign n26624 = ( x618 & x1154 ) | ( x618 & n26541 ) | ( x1154 & n26541 ) ;
  assign n26625 = ( ~x618 & x1154 ) | ( ~x618 & n26619 ) | ( x1154 & n26619 ) ;
  assign n26626 = n26624 & n26625 ;
  assign n26627 = n26623 & ~n26626 ;
  assign n26628 = n26622 & ~n26627 ;
  assign n26629 = x781 & ~n26628 ;
  assign n26630 = x781 | n26619 ;
  assign n26631 = ~n26629 & n26630 ;
  assign n26632 = ( x619 & ~x1159 ) | ( x619 & n26631 ) | ( ~x1159 & n26631 ) ;
  assign n26633 = ~n26576 & n26632 ;
  assign n26634 = n26575 | n26633 ;
  assign n26635 = x648 & ~n26501 ;
  assign n26636 = ( x619 & x1159 ) | ( x619 & n26544 ) | ( x1159 & n26544 ) ;
  assign n26637 = ( ~x619 & x1159 ) | ( ~x619 & n26631 ) | ( x1159 & n26631 ) ;
  assign n26638 = n26636 & n26637 ;
  assign n26639 = n26635 & ~n26638 ;
  assign n26640 = n26634 & ~n26639 ;
  assign n26641 = x789 & ~n26640 ;
  assign n26642 = x789 | n26631 ;
  assign n26643 = ~n26641 & n26642 ;
  assign n26644 = ~x788 & n26643 ;
  assign n26645 = ( x626 & x641 ) | ( x626 & ~n26504 ) | ( x641 & ~n26504 ) ;
  assign n26646 = ( x626 & ~x641 ) | ( x626 & n26457 ) | ( ~x641 & n26457 ) ;
  assign n26647 = n26645 & ~n26646 ;
  assign n26648 = x1158 | n26647 ;
  assign n26649 = ( x626 & x641 ) | ( x626 & n26546 ) | ( x641 & n26546 ) ;
  assign n26650 = ( ~x626 & x641 ) | ( ~x626 & n26643 ) | ( x641 & n26643 ) ;
  assign n26651 = n26649 | n26650 ;
  assign n26652 = ~n26648 & n26651 ;
  assign n26653 = ( x626 & x641 ) | ( x626 & n26504 ) | ( x641 & n26504 ) ;
  assign n26654 = ( ~x626 & x641 ) | ( ~x626 & n26457 ) | ( x641 & n26457 ) ;
  assign n26655 = n26653 | n26654 ;
  assign n26656 = x1158 & n26655 ;
  assign n26657 = ( x626 & x641 ) | ( x626 & ~n26546 ) | ( x641 & ~n26546 ) ;
  assign n26658 = ( x626 & ~x641 ) | ( x626 & n26643 ) | ( ~x641 & n26643 ) ;
  assign n26659 = n26657 & ~n26658 ;
  assign n26660 = n26656 & ~n26659 ;
  assign n26661 = n26652 | n26660 ;
  assign n26662 = x788 & n26661 ;
  assign n26663 = n26644 | n26662 ;
  assign n26664 = ( x628 & ~x1156 ) | ( x628 & n26663 ) | ( ~x1156 & n26663 ) ;
  assign n26665 = ~n26574 & n26664 ;
  assign n26666 = n26573 | n26665 ;
  assign n26667 = x629 & ~n26556 ;
  assign n26668 = ( x628 & x1156 ) | ( x628 & n26507 ) | ( x1156 & n26507 ) ;
  assign n26669 = ( ~x628 & x1156 ) | ( ~x628 & n26663 ) | ( x1156 & n26663 ) ;
  assign n26670 = n26668 & n26669 ;
  assign n26671 = n26667 & ~n26670 ;
  assign n26672 = n26666 & ~n26671 ;
  assign n26673 = x792 & ~n26672 ;
  assign n26674 = x792 | n26663 ;
  assign n26675 = ~n26673 & n26674 ;
  assign n26676 = ( x647 & ~x1157 ) | ( x647 & n26675 ) | ( ~x1157 & n26675 ) ;
  assign n26677 = ~n26572 & n26676 ;
  assign n26678 = n26571 | n26677 ;
  assign n26679 = x630 & ~n26566 ;
  assign n26680 = ( x647 & x1157 ) | ( x647 & n26510 ) | ( x1157 & n26510 ) ;
  assign n26681 = ( ~x647 & x1157 ) | ( ~x647 & n26675 ) | ( x1157 & n26675 ) ;
  assign n26682 = n26680 & n26681 ;
  assign n26683 = n26679 & ~n26682 ;
  assign n26684 = n26678 & ~n26683 ;
  assign n26685 = x787 & ~n26684 ;
  assign n26686 = x787 | n26675 ;
  assign n26687 = ~n26685 & n26686 ;
  assign n26688 = ( x644 & ~x715 ) | ( x644 & n26687 ) | ( ~x715 & n26687 ) ;
  assign n26689 = ~n26570 & n26688 ;
  assign n26690 = n26516 | n26689 ;
  assign n26691 = ( x644 & x715 ) | ( x644 & ~n26512 ) | ( x715 & ~n26512 ) ;
  assign n26692 = ( x644 & ~x715 ) | ( x644 & n26457 ) | ( ~x715 & n26457 ) ;
  assign n26693 = ~n26691 & n26692 ;
  assign n26694 = x1160 & ~n26693 ;
  assign n26695 = ( x644 & x715 ) | ( x644 & n26569 ) | ( x715 & n26569 ) ;
  assign n26696 = ( ~x644 & x715 ) | ( ~x644 & n26687 ) | ( x715 & n26687 ) ;
  assign n26697 = n26695 & n26696 ;
  assign n26698 = n26694 & ~n26697 ;
  assign n26699 = x790 & ~n26698 ;
  assign n26700 = n26690 & n26699 ;
  assign n26701 = ~x790 & n26687 ;
  assign n26702 = n6785 | n26701 ;
  assign n26703 = n26700 | n26702 ;
  assign n26704 = ~x186 & n6785 ;
  assign n26705 = x832 | n26704 ;
  assign n26706 = n26703 & ~n26705 ;
  assign n26707 = x186 | n1290 ;
  assign n26708 = ~x752 & n14840 ;
  assign n26709 = n26707 & ~n26708 ;
  assign n26710 = n16060 | n26709 ;
  assign n26711 = ~x785 & n26710 ;
  assign n26712 = n16065 | n26709 ;
  assign n26713 = x1155 & n26712 ;
  assign n26714 = n16068 | n26710 ;
  assign n26715 = ~x1155 & n26714 ;
  assign n26716 = n26713 | n26715 ;
  assign n26717 = x785 & n26716 ;
  assign n26718 = n26711 | n26717 ;
  assign n26719 = ~x781 & n26718 ;
  assign n26720 = n16075 | n26718 ;
  assign n26721 = x1154 & n26720 ;
  assign n26722 = n16078 | n26718 ;
  assign n26723 = ~x1154 & n26722 ;
  assign n26724 = n26721 | n26723 ;
  assign n26725 = x781 & n26724 ;
  assign n26726 = n26719 | n26725 ;
  assign n26727 = ~x789 & n26726 ;
  assign n26728 = ( x619 & x1159 ) | ( x619 & n26707 ) | ( x1159 & n26707 ) ;
  assign n26729 = ( ~x619 & x1159 ) | ( ~x619 & n26726 ) | ( x1159 & n26726 ) ;
  assign n26730 = n26728 & n26729 ;
  assign n26731 = ( x619 & x1159 ) | ( x619 & ~n26707 ) | ( x1159 & ~n26707 ) ;
  assign n26732 = ( x619 & ~x1159 ) | ( x619 & n26726 ) | ( ~x1159 & n26726 ) ;
  assign n26733 = ~n26731 & n26732 ;
  assign n26734 = n26730 | n26733 ;
  assign n26735 = x789 & n26734 ;
  assign n26736 = n26727 | n26735 ;
  assign n26737 = n16176 | n26736 ;
  assign n26738 = n16176 & ~n26707 ;
  assign n26739 = n26737 & ~n26738 ;
  assign n26740 = n15134 | n26739 ;
  assign n26741 = n15134 & ~n26707 ;
  assign n26742 = n26740 & ~n26741 ;
  assign n26743 = n18610 & n26742 ;
  assign n26744 = ( x647 & x1157 ) | ( x647 & ~n26707 ) | ( x1157 & ~n26707 ) ;
  assign n26745 = x703 & n15202 ;
  assign n26746 = n26707 & ~n26745 ;
  assign n26747 = ~x778 & n26746 ;
  assign n26748 = ~x625 & n26745 ;
  assign n26749 = n26746 | n26748 ;
  assign n26750 = x1153 & n26749 ;
  assign n26751 = ~x1153 & n26707 ;
  assign n26752 = ~n26748 & n26751 ;
  assign n26753 = n26750 | n26752 ;
  assign n26754 = x778 & n26753 ;
  assign n26755 = n26747 | n26754 ;
  assign n26756 = n16043 | n26755 ;
  assign n26757 = n16045 | n26756 ;
  assign n26758 = n16047 | n26757 ;
  assign n26759 = n16049 | n26758 ;
  assign n26760 = n16055 | n26759 ;
  assign n26761 = ( x647 & ~x1157 ) | ( x647 & n26760 ) | ( ~x1157 & n26760 ) ;
  assign n26762 = ~n26744 & n26761 ;
  assign n26763 = x630 & n26762 ;
  assign n26764 = x647 & n26760 ;
  assign n26765 = ~x647 & n26707 ;
  assign n26766 = n26764 | n26765 ;
  assign n26767 = n15138 & n26766 ;
  assign n26768 = n26763 | n26767 ;
  assign n26769 = n26743 | n26768 ;
  assign n26770 = x787 & n26769 ;
  assign n26771 = n16115 & ~n26758 ;
  assign n26772 = ( x626 & ~n15419 ) | ( x626 & n26707 ) | ( ~n15419 & n26707 ) ;
  assign n26773 = ( x626 & n15419 ) | ( x626 & ~n26736 ) | ( n15419 & ~n26736 ) ;
  assign n26774 = ~n26772 & n26773 ;
  assign n26775 = n26771 | n26774 ;
  assign n26776 = ( x626 & n15418 ) | ( x626 & ~n26707 ) | ( n15418 & ~n26707 ) ;
  assign n26777 = ( x626 & ~n15418 ) | ( x626 & n26736 ) | ( ~n15418 & n26736 ) ;
  assign n26778 = n26776 & ~n26777 ;
  assign n26779 = n26775 | n26778 ;
  assign n26780 = x788 & n26779 ;
  assign n26781 = x648 & ~n26733 ;
  assign n26782 = ( x619 & x1159 ) | ( x619 & n26757 ) | ( x1159 & n26757 ) ;
  assign n26783 = x627 | n26721 ;
  assign n26784 = ( x618 & x1154 ) | ( x618 & ~n26756 ) | ( x1154 & ~n26756 ) ;
  assign n26785 = x660 | n26713 ;
  assign n26786 = ( x609 & x1155 ) | ( x609 & ~n26755 ) | ( x1155 & ~n26755 ) ;
  assign n26787 = n14839 | n26746 ;
  assign n26788 = x625 & ~n26787 ;
  assign n26789 = n26709 & n26787 ;
  assign n26790 = n26788 | n26789 ;
  assign n26791 = n26751 & n26790 ;
  assign n26792 = x608 | n26750 ;
  assign n26793 = n26791 | n26792 ;
  assign n26794 = x1153 & n26709 ;
  assign n26795 = ~n26788 & n26794 ;
  assign n26796 = x608 & ~n26752 ;
  assign n26797 = ~n26795 & n26796 ;
  assign n26798 = n26793 & ~n26797 ;
  assign n26799 = x778 & ~n26798 ;
  assign n26800 = x778 | n26789 ;
  assign n26801 = ~n26799 & n26800 ;
  assign n26802 = ( x609 & ~x1155 ) | ( x609 & n26801 ) | ( ~x1155 & n26801 ) ;
  assign n26803 = ~n26786 & n26802 ;
  assign n26804 = n26785 | n26803 ;
  assign n26805 = x660 & ~n26715 ;
  assign n26806 = ( x609 & x1155 ) | ( x609 & n26755 ) | ( x1155 & n26755 ) ;
  assign n26807 = ( ~x609 & x1155 ) | ( ~x609 & n26801 ) | ( x1155 & n26801 ) ;
  assign n26808 = n26806 & n26807 ;
  assign n26809 = n26805 & ~n26808 ;
  assign n26810 = n26804 & ~n26809 ;
  assign n26811 = x785 & ~n26810 ;
  assign n26812 = x785 | n26801 ;
  assign n26813 = ~n26811 & n26812 ;
  assign n26814 = ( x618 & ~x1154 ) | ( x618 & n26813 ) | ( ~x1154 & n26813 ) ;
  assign n26815 = ~n26784 & n26814 ;
  assign n26816 = n26783 | n26815 ;
  assign n26817 = x627 & ~n26723 ;
  assign n26818 = ( x618 & x1154 ) | ( x618 & n26756 ) | ( x1154 & n26756 ) ;
  assign n26819 = ( ~x618 & x1154 ) | ( ~x618 & n26813 ) | ( x1154 & n26813 ) ;
  assign n26820 = n26818 & n26819 ;
  assign n26821 = n26817 & ~n26820 ;
  assign n26822 = n26816 & ~n26821 ;
  assign n26823 = x781 & ~n26822 ;
  assign n26824 = x781 | n26813 ;
  assign n26825 = ~n26823 & n26824 ;
  assign n26826 = ( ~x619 & x1159 ) | ( ~x619 & n26825 ) | ( x1159 & n26825 ) ;
  assign n26827 = n26782 & n26826 ;
  assign n26828 = n26781 & ~n26827 ;
  assign n26829 = x648 | n26730 ;
  assign n26830 = ( x619 & x1159 ) | ( x619 & ~n26757 ) | ( x1159 & ~n26757 ) ;
  assign n26831 = ( x619 & ~x1159 ) | ( x619 & n26825 ) | ( ~x1159 & n26825 ) ;
  assign n26832 = ~n26830 & n26831 ;
  assign n26833 = n26829 | n26832 ;
  assign n26834 = x789 & n26833 ;
  assign n26835 = ~n26828 & n26834 ;
  assign n26836 = ~x789 & n26825 ;
  assign n26837 = n16177 | n26836 ;
  assign n26838 = n26835 | n26837 ;
  assign n26839 = ~n26780 & n26838 ;
  assign n26840 = n18434 | n26839 ;
  assign n26841 = n16650 | n26759 ;
  assign n26842 = n16051 & ~n26739 ;
  assign n26843 = n26841 & ~n26842 ;
  assign n26844 = ( x629 & ~x792 ) | ( x629 & n26843 ) | ( ~x792 & n26843 ) ;
  assign n26845 = n16052 & ~n26739 ;
  assign n26846 = n16643 & ~n26759 ;
  assign n26847 = n26845 | n26846 ;
  assign n26848 = ( x629 & x792 ) | ( x629 & n26847 ) | ( x792 & n26847 ) ;
  assign n26849 = ~n26844 & n26848 ;
  assign n26850 = n18431 | n26849 ;
  assign n26851 = n26840 & ~n26850 ;
  assign n26852 = n26770 | n26851 ;
  assign n26853 = ( x790 & x832 ) | ( x790 & n26852 ) | ( x832 & n26852 ) ;
  assign n26854 = n15141 | n26742 ;
  assign n26855 = n15141 & ~n26707 ;
  assign n26856 = n26854 & ~n26855 ;
  assign n26857 = ( x644 & x715 ) | ( x644 & ~n26856 ) | ( x715 & ~n26856 ) ;
  assign n26858 = ( x644 & ~x715 ) | ( x644 & n26707 ) | ( ~x715 & n26707 ) ;
  assign n26859 = ~n26857 & n26858 ;
  assign n26860 = x1160 & ~n26859 ;
  assign n26861 = ~x787 & n26760 ;
  assign n26862 = x1157 & n26766 ;
  assign n26863 = n26762 | n26862 ;
  assign n26864 = x787 & n26863 ;
  assign n26865 = n26861 | n26864 ;
  assign n26866 = ( x644 & x715 ) | ( x644 & n26865 ) | ( x715 & n26865 ) ;
  assign n26867 = ( ~x644 & x715 ) | ( ~x644 & n26852 ) | ( x715 & n26852 ) ;
  assign n26868 = n26866 & n26867 ;
  assign n26869 = n26860 & ~n26868 ;
  assign n26870 = ( x644 & x715 ) | ( x644 & n26856 ) | ( x715 & n26856 ) ;
  assign n26871 = ( ~x644 & x715 ) | ( ~x644 & n26707 ) | ( x715 & n26707 ) ;
  assign n26872 = n26870 & n26871 ;
  assign n26873 = x1160 | n26872 ;
  assign n26874 = ( x644 & x715 ) | ( x644 & ~n26865 ) | ( x715 & ~n26865 ) ;
  assign n26875 = ( x644 & ~x715 ) | ( x644 & n26852 ) | ( ~x715 & n26852 ) ;
  assign n26876 = ~n26874 & n26875 ;
  assign n26877 = n26873 | n26876 ;
  assign n26878 = ~n26869 & n26877 ;
  assign n26879 = ( ~x790 & x832 ) | ( ~x790 & n26878 ) | ( x832 & n26878 ) ;
  assign n26880 = n26853 & n26879 ;
  assign n26881 = n26706 | n26880 ;
  assign n26882 = x187 | n14834 ;
  assign n26883 = n15141 & n26882 ;
  assign n26884 = x187 & n2032 ;
  assign n26885 = x770 | n17421 ;
  assign n26886 = ~n19012 & n26885 ;
  assign n26887 = x187 | n26886 ;
  assign n26888 = x187 | n17415 ;
  assign n26889 = ~x770 & n26888 ;
  assign n26890 = n22415 & n26889 ;
  assign n26891 = n26887 & ~n26890 ;
  assign n26892 = ~n2032 & n26891 ;
  assign n26893 = n26884 | n26892 ;
  assign n26894 = ~n15082 & n26893 ;
  assign n26895 = n15082 & n26882 ;
  assign n26896 = n26894 | n26895 ;
  assign n26897 = ~x785 & n26896 ;
  assign n26898 = ~n15088 & n26882 ;
  assign n26899 = x609 & n26894 ;
  assign n26900 = n26898 | n26899 ;
  assign n26901 = x1155 & n26900 ;
  assign n26902 = n15094 & n26882 ;
  assign n26903 = ~x609 & n26894 ;
  assign n26904 = n26902 | n26903 ;
  assign n26905 = ~x1155 & n26904 ;
  assign n26906 = n26901 | n26905 ;
  assign n26907 = x785 & n26906 ;
  assign n26908 = n26897 | n26907 ;
  assign n26909 = ~x781 & n26908 ;
  assign n26910 = ( x618 & x1154 ) | ( x618 & n26882 ) | ( x1154 & n26882 ) ;
  assign n26911 = ( ~x618 & x1154 ) | ( ~x618 & n26908 ) | ( x1154 & n26908 ) ;
  assign n26912 = n26910 & n26911 ;
  assign n26913 = ( x618 & x1154 ) | ( x618 & ~n26882 ) | ( x1154 & ~n26882 ) ;
  assign n26914 = ( x618 & ~x1154 ) | ( x618 & n26908 ) | ( ~x1154 & n26908 ) ;
  assign n26915 = ~n26913 & n26914 ;
  assign n26916 = n26912 | n26915 ;
  assign n26917 = x781 & n26916 ;
  assign n26918 = n26909 | n26917 ;
  assign n26919 = ~x789 & n26918 ;
  assign n26920 = ( x619 & x1159 ) | ( x619 & n26882 ) | ( x1159 & n26882 ) ;
  assign n26921 = ( ~x619 & x1159 ) | ( ~x619 & n26918 ) | ( x1159 & n26918 ) ;
  assign n26922 = n26920 & n26921 ;
  assign n26923 = ( x619 & x1159 ) | ( x619 & ~n26882 ) | ( x1159 & ~n26882 ) ;
  assign n26924 = ( x619 & ~x1159 ) | ( x619 & n26918 ) | ( ~x1159 & n26918 ) ;
  assign n26925 = ~n26923 & n26924 ;
  assign n26926 = n26922 | n26925 ;
  assign n26927 = x789 & n26926 ;
  assign n26928 = n26919 | n26927 ;
  assign n26929 = n16176 | n26928 ;
  assign n26930 = n16176 & ~n26882 ;
  assign n26931 = n26929 & ~n26930 ;
  assign n26932 = n15134 | n26931 ;
  assign n26933 = n15134 & ~n26882 ;
  assign n26934 = n26932 & ~n26933 ;
  assign n26935 = ~n15141 & n26934 ;
  assign n26936 = n26883 | n26935 ;
  assign n26937 = ( x644 & x715 ) | ( x644 & n26936 ) | ( x715 & n26936 ) ;
  assign n26938 = ( ~x644 & x715 ) | ( ~x644 & n26882 ) | ( x715 & n26882 ) ;
  assign n26939 = n26937 & n26938 ;
  assign n26940 = x1160 | n26939 ;
  assign n26941 = n15414 & n26882 ;
  assign n26942 = x187 | n15070 ;
  assign n26943 = n15375 & n26942 ;
  assign n26944 = x726 & ~n26943 ;
  assign n26945 = ( ~x38 & x187 ) | ( ~x38 & n16319 ) | ( x187 & n16319 ) ;
  assign n26946 = ( x38 & x187 ) | ( x38 & n16323 ) | ( x187 & n16323 ) ;
  assign n26947 = n26945 & ~n26946 ;
  assign n26948 = n26944 & ~n26947 ;
  assign n26949 = x187 | x726 ;
  assign n26950 = n15382 | n26949 ;
  assign n26951 = ~n2032 & n26950 ;
  assign n26952 = ~n26948 & n26951 ;
  assign n26953 = n26884 | n26952 ;
  assign n26954 = ~x778 & n26953 ;
  assign n26955 = ( x625 & x1153 ) | ( x625 & n26882 ) | ( x1153 & n26882 ) ;
  assign n26956 = ( ~x625 & x1153 ) | ( ~x625 & n26953 ) | ( x1153 & n26953 ) ;
  assign n26957 = n26955 & n26956 ;
  assign n26958 = ( x625 & x1153 ) | ( x625 & ~n26882 ) | ( x1153 & ~n26882 ) ;
  assign n26959 = ( x625 & ~x1153 ) | ( x625 & n26953 ) | ( ~x1153 & n26953 ) ;
  assign n26960 = ~n26958 & n26959 ;
  assign n26961 = n26957 | n26960 ;
  assign n26962 = x778 & n26961 ;
  assign n26963 = n26954 | n26962 ;
  assign n26964 = ~n15400 & n26963 ;
  assign n26965 = n15400 & n26882 ;
  assign n26966 = n26964 | n26965 ;
  assign n26967 = n15407 | n26966 ;
  assign n26968 = n15407 & ~n26882 ;
  assign n26969 = n26967 & ~n26968 ;
  assign n26970 = ~n15414 & n26969 ;
  assign n26971 = n26941 | n26970 ;
  assign n26972 = n15421 | n26971 ;
  assign n26973 = n15421 & ~n26882 ;
  assign n26974 = n26972 & ~n26973 ;
  assign n26975 = ~x792 & n26974 ;
  assign n26976 = ( x628 & x1156 ) | ( x628 & n26882 ) | ( x1156 & n26882 ) ;
  assign n26977 = ( ~x628 & x1156 ) | ( ~x628 & n26974 ) | ( x1156 & n26974 ) ;
  assign n26978 = n26976 & n26977 ;
  assign n26979 = ( x628 & x1156 ) | ( x628 & ~n26882 ) | ( x1156 & ~n26882 ) ;
  assign n26980 = ( x628 & ~x1156 ) | ( x628 & n26974 ) | ( ~x1156 & n26974 ) ;
  assign n26981 = ~n26979 & n26980 ;
  assign n26982 = n26978 | n26981 ;
  assign n26983 = x792 & n26982 ;
  assign n26984 = n26975 | n26983 ;
  assign n26985 = ~x787 & n26984 ;
  assign n26986 = ( x647 & x1157 ) | ( x647 & n26882 ) | ( x1157 & n26882 ) ;
  assign n26987 = ( ~x647 & x1157 ) | ( ~x647 & n26984 ) | ( x1157 & n26984 ) ;
  assign n26988 = n26986 & n26987 ;
  assign n26989 = ( x647 & x1157 ) | ( x647 & ~n26882 ) | ( x1157 & ~n26882 ) ;
  assign n26990 = ( x647 & ~x1157 ) | ( x647 & n26984 ) | ( ~x1157 & n26984 ) ;
  assign n26991 = ~n26989 & n26990 ;
  assign n26992 = n26988 | n26991 ;
  assign n26993 = x787 & n26992 ;
  assign n26994 = n26985 | n26993 ;
  assign n26995 = ( x644 & x715 ) | ( x644 & ~n26994 ) | ( x715 & ~n26994 ) ;
  assign n26996 = x630 | n26988 ;
  assign n26997 = ( x647 & x1157 ) | ( x647 & ~n26934 ) | ( x1157 & ~n26934 ) ;
  assign n26998 = x629 | n26978 ;
  assign n26999 = ( x628 & x1156 ) | ( x628 & ~n26931 ) | ( x1156 & ~n26931 ) ;
  assign n27000 = x648 | n26922 ;
  assign n27001 = ( x619 & x1159 ) | ( x619 & ~n26969 ) | ( x1159 & ~n26969 ) ;
  assign n27002 = x627 | n26912 ;
  assign n27003 = ( x618 & x1154 ) | ( x618 & ~n26966 ) | ( x1154 & ~n26966 ) ;
  assign n27004 = x660 | n26901 ;
  assign n27005 = ( x609 & x1155 ) | ( x609 & ~n26963 ) | ( x1155 & ~n26963 ) ;
  assign n27006 = x608 | n26957 ;
  assign n27007 = ( x625 & x1153 ) | ( x625 & ~n26893 ) | ( x1153 & ~n26893 ) ;
  assign n27008 = x726 | n26891 ;
  assign n27009 = ( x187 & ~x770 ) | ( x187 & n17554 ) | ( ~x770 & n17554 ) ;
  assign n27010 = ( x187 & x770 ) | ( x187 & n17562 ) | ( x770 & n17562 ) ;
  assign n27011 = n27009 & ~n27010 ;
  assign n27012 = x726 & ~n27011 ;
  assign n27013 = x770 & ~n17570 ;
  assign n27014 = ( x187 & n17569 ) | ( x187 & ~n27013 ) | ( n17569 & ~n27013 ) ;
  assign n27015 = ( x187 & n17579 ) | ( x187 & n27013 ) | ( n17579 & n27013 ) ;
  assign n27016 = ~n27014 & n27015 ;
  assign n27017 = n27012 & ~n27016 ;
  assign n27018 = n2032 | n27017 ;
  assign n27019 = n27008 & ~n27018 ;
  assign n27020 = n26884 | n27019 ;
  assign n27021 = ( x625 & ~x1153 ) | ( x625 & n27020 ) | ( ~x1153 & n27020 ) ;
  assign n27022 = ~n27007 & n27021 ;
  assign n27023 = n27006 | n27022 ;
  assign n27024 = x608 & ~n26960 ;
  assign n27025 = ( x625 & x1153 ) | ( x625 & n26893 ) | ( x1153 & n26893 ) ;
  assign n27026 = ( ~x625 & x1153 ) | ( ~x625 & n27020 ) | ( x1153 & n27020 ) ;
  assign n27027 = n27025 & n27026 ;
  assign n27028 = n27024 & ~n27027 ;
  assign n27029 = n27023 & ~n27028 ;
  assign n27030 = x778 & ~n27029 ;
  assign n27031 = x778 | n27020 ;
  assign n27032 = ~n27030 & n27031 ;
  assign n27033 = ( x609 & ~x1155 ) | ( x609 & n27032 ) | ( ~x1155 & n27032 ) ;
  assign n27034 = ~n27005 & n27033 ;
  assign n27035 = n27004 | n27034 ;
  assign n27036 = x660 & ~n26905 ;
  assign n27037 = ( x609 & x1155 ) | ( x609 & n26963 ) | ( x1155 & n26963 ) ;
  assign n27038 = ( ~x609 & x1155 ) | ( ~x609 & n27032 ) | ( x1155 & n27032 ) ;
  assign n27039 = n27037 & n27038 ;
  assign n27040 = n27036 & ~n27039 ;
  assign n27041 = n27035 & ~n27040 ;
  assign n27042 = x785 & ~n27041 ;
  assign n27043 = x785 | n27032 ;
  assign n27044 = ~n27042 & n27043 ;
  assign n27045 = ( x618 & ~x1154 ) | ( x618 & n27044 ) | ( ~x1154 & n27044 ) ;
  assign n27046 = ~n27003 & n27045 ;
  assign n27047 = n27002 | n27046 ;
  assign n27048 = x627 & ~n26915 ;
  assign n27049 = ( x618 & x1154 ) | ( x618 & n26966 ) | ( x1154 & n26966 ) ;
  assign n27050 = ( ~x618 & x1154 ) | ( ~x618 & n27044 ) | ( x1154 & n27044 ) ;
  assign n27051 = n27049 & n27050 ;
  assign n27052 = n27048 & ~n27051 ;
  assign n27053 = n27047 & ~n27052 ;
  assign n27054 = x781 & ~n27053 ;
  assign n27055 = x781 | n27044 ;
  assign n27056 = ~n27054 & n27055 ;
  assign n27057 = ( x619 & ~x1159 ) | ( x619 & n27056 ) | ( ~x1159 & n27056 ) ;
  assign n27058 = ~n27001 & n27057 ;
  assign n27059 = n27000 | n27058 ;
  assign n27060 = x648 & ~n26925 ;
  assign n27061 = ( x619 & x1159 ) | ( x619 & n26969 ) | ( x1159 & n26969 ) ;
  assign n27062 = ( ~x619 & x1159 ) | ( ~x619 & n27056 ) | ( x1159 & n27056 ) ;
  assign n27063 = n27061 & n27062 ;
  assign n27064 = n27060 & ~n27063 ;
  assign n27065 = n27059 & ~n27064 ;
  assign n27066 = x789 & ~n27065 ;
  assign n27067 = x789 | n27056 ;
  assign n27068 = ~n27066 & n27067 ;
  assign n27069 = ~x788 & n27068 ;
  assign n27070 = ( x626 & x641 ) | ( x626 & ~n26928 ) | ( x641 & ~n26928 ) ;
  assign n27071 = ( x626 & ~x641 ) | ( x626 & n26882 ) | ( ~x641 & n26882 ) ;
  assign n27072 = n27070 & ~n27071 ;
  assign n27073 = x1158 | n27072 ;
  assign n27074 = ( x626 & x641 ) | ( x626 & n26971 ) | ( x641 & n26971 ) ;
  assign n27075 = ( ~x626 & x641 ) | ( ~x626 & n27068 ) | ( x641 & n27068 ) ;
  assign n27076 = n27074 | n27075 ;
  assign n27077 = ~n27073 & n27076 ;
  assign n27078 = ( x626 & x641 ) | ( x626 & n26928 ) | ( x641 & n26928 ) ;
  assign n27079 = ( ~x626 & x641 ) | ( ~x626 & n26882 ) | ( x641 & n26882 ) ;
  assign n27080 = n27078 | n27079 ;
  assign n27081 = x1158 & n27080 ;
  assign n27082 = ( x626 & x641 ) | ( x626 & ~n26971 ) | ( x641 & ~n26971 ) ;
  assign n27083 = ( x626 & ~x641 ) | ( x626 & n27068 ) | ( ~x641 & n27068 ) ;
  assign n27084 = n27082 & ~n27083 ;
  assign n27085 = n27081 & ~n27084 ;
  assign n27086 = n27077 | n27085 ;
  assign n27087 = x788 & n27086 ;
  assign n27088 = n27069 | n27087 ;
  assign n27089 = ( x628 & ~x1156 ) | ( x628 & n27088 ) | ( ~x1156 & n27088 ) ;
  assign n27090 = ~n26999 & n27089 ;
  assign n27091 = n26998 | n27090 ;
  assign n27092 = x629 & ~n26981 ;
  assign n27093 = ( x628 & x1156 ) | ( x628 & n26931 ) | ( x1156 & n26931 ) ;
  assign n27094 = ( ~x628 & x1156 ) | ( ~x628 & n27088 ) | ( x1156 & n27088 ) ;
  assign n27095 = n27093 & n27094 ;
  assign n27096 = n27092 & ~n27095 ;
  assign n27097 = n27091 & ~n27096 ;
  assign n27098 = x792 & ~n27097 ;
  assign n27099 = x792 | n27088 ;
  assign n27100 = ~n27098 & n27099 ;
  assign n27101 = ( x647 & ~x1157 ) | ( x647 & n27100 ) | ( ~x1157 & n27100 ) ;
  assign n27102 = ~n26997 & n27101 ;
  assign n27103 = n26996 | n27102 ;
  assign n27104 = x630 & ~n26991 ;
  assign n27105 = ( x647 & x1157 ) | ( x647 & n26934 ) | ( x1157 & n26934 ) ;
  assign n27106 = ( ~x647 & x1157 ) | ( ~x647 & n27100 ) | ( x1157 & n27100 ) ;
  assign n27107 = n27105 & n27106 ;
  assign n27108 = n27104 & ~n27107 ;
  assign n27109 = n27103 & ~n27108 ;
  assign n27110 = x787 & ~n27109 ;
  assign n27111 = x787 | n27100 ;
  assign n27112 = ~n27110 & n27111 ;
  assign n27113 = ( x644 & ~x715 ) | ( x644 & n27112 ) | ( ~x715 & n27112 ) ;
  assign n27114 = ~n26995 & n27113 ;
  assign n27115 = n26940 | n27114 ;
  assign n27116 = ( x644 & x715 ) | ( x644 & ~n26936 ) | ( x715 & ~n26936 ) ;
  assign n27117 = ( x644 & ~x715 ) | ( x644 & n26882 ) | ( ~x715 & n26882 ) ;
  assign n27118 = ~n27116 & n27117 ;
  assign n27119 = x1160 & ~n27118 ;
  assign n27120 = ( x644 & x715 ) | ( x644 & n26994 ) | ( x715 & n26994 ) ;
  assign n27121 = ( ~x644 & x715 ) | ( ~x644 & n27112 ) | ( x715 & n27112 ) ;
  assign n27122 = n27120 & n27121 ;
  assign n27123 = n27119 & ~n27122 ;
  assign n27124 = x790 & ~n27123 ;
  assign n27125 = n27115 & n27124 ;
  assign n27126 = ~x790 & n27112 ;
  assign n27127 = n6785 | n27126 ;
  assign n27128 = n27125 | n27127 ;
  assign n27129 = ~x187 & n6785 ;
  assign n27130 = x832 | n27129 ;
  assign n27131 = n27128 & ~n27130 ;
  assign n27132 = x187 | n1290 ;
  assign n27133 = ~x770 & n14840 ;
  assign n27134 = n27132 & ~n27133 ;
  assign n27135 = n16060 | n27134 ;
  assign n27136 = ~x785 & n27135 ;
  assign n27137 = n16065 | n27134 ;
  assign n27138 = x1155 & n27137 ;
  assign n27139 = n16068 | n27135 ;
  assign n27140 = ~x1155 & n27139 ;
  assign n27141 = n27138 | n27140 ;
  assign n27142 = x785 & n27141 ;
  assign n27143 = n27136 | n27142 ;
  assign n27144 = ~x781 & n27143 ;
  assign n27145 = n16075 | n27143 ;
  assign n27146 = x1154 & n27145 ;
  assign n27147 = n16078 | n27143 ;
  assign n27148 = ~x1154 & n27147 ;
  assign n27149 = n27146 | n27148 ;
  assign n27150 = x781 & n27149 ;
  assign n27151 = n27144 | n27150 ;
  assign n27152 = ~x789 & n27151 ;
  assign n27153 = ( x619 & x1159 ) | ( x619 & n27132 ) | ( x1159 & n27132 ) ;
  assign n27154 = ( ~x619 & x1159 ) | ( ~x619 & n27151 ) | ( x1159 & n27151 ) ;
  assign n27155 = n27153 & n27154 ;
  assign n27156 = ( x619 & x1159 ) | ( x619 & ~n27132 ) | ( x1159 & ~n27132 ) ;
  assign n27157 = ( x619 & ~x1159 ) | ( x619 & n27151 ) | ( ~x1159 & n27151 ) ;
  assign n27158 = ~n27156 & n27157 ;
  assign n27159 = n27155 | n27158 ;
  assign n27160 = x789 & n27159 ;
  assign n27161 = n27152 | n27160 ;
  assign n27162 = n16176 | n27161 ;
  assign n27163 = n16176 & ~n27132 ;
  assign n27164 = n27162 & ~n27163 ;
  assign n27165 = n15134 | n27164 ;
  assign n27166 = n15134 & ~n27132 ;
  assign n27167 = n27165 & ~n27166 ;
  assign n27168 = n18610 & n27167 ;
  assign n27169 = ( x647 & x1157 ) | ( x647 & ~n27132 ) | ( x1157 & ~n27132 ) ;
  assign n27170 = x726 & n15202 ;
  assign n27171 = n27132 & ~n27170 ;
  assign n27172 = ~x778 & n27171 ;
  assign n27173 = ~x625 & n27170 ;
  assign n27174 = n27171 | n27173 ;
  assign n27175 = x1153 & n27174 ;
  assign n27176 = ~x1153 & n27132 ;
  assign n27177 = ~n27173 & n27176 ;
  assign n27178 = n27175 | n27177 ;
  assign n27179 = x778 & n27178 ;
  assign n27180 = n27172 | n27179 ;
  assign n27181 = n16043 | n27180 ;
  assign n27182 = n16045 | n27181 ;
  assign n27183 = n16047 | n27182 ;
  assign n27184 = n16049 | n27183 ;
  assign n27185 = n16055 | n27184 ;
  assign n27186 = ( x647 & ~x1157 ) | ( x647 & n27185 ) | ( ~x1157 & n27185 ) ;
  assign n27187 = ~n27169 & n27186 ;
  assign n27188 = x630 & n27187 ;
  assign n27189 = x647 & n27185 ;
  assign n27190 = ~x647 & n27132 ;
  assign n27191 = n27189 | n27190 ;
  assign n27192 = n15138 & n27191 ;
  assign n27193 = n27188 | n27192 ;
  assign n27194 = n27168 | n27193 ;
  assign n27195 = x787 & n27194 ;
  assign n27196 = n16115 & ~n27183 ;
  assign n27197 = ( x626 & ~n15419 ) | ( x626 & n27132 ) | ( ~n15419 & n27132 ) ;
  assign n27198 = ( x626 & n15419 ) | ( x626 & ~n27161 ) | ( n15419 & ~n27161 ) ;
  assign n27199 = ~n27197 & n27198 ;
  assign n27200 = n27196 | n27199 ;
  assign n27201 = ( x626 & n15418 ) | ( x626 & ~n27132 ) | ( n15418 & ~n27132 ) ;
  assign n27202 = ( x626 & ~n15418 ) | ( x626 & n27161 ) | ( ~n15418 & n27161 ) ;
  assign n27203 = n27201 & ~n27202 ;
  assign n27204 = n27200 | n27203 ;
  assign n27205 = x788 & n27204 ;
  assign n27206 = x648 & ~n27158 ;
  assign n27207 = ( x619 & x1159 ) | ( x619 & n27182 ) | ( x1159 & n27182 ) ;
  assign n27208 = x627 | n27146 ;
  assign n27209 = ( x618 & x1154 ) | ( x618 & ~n27181 ) | ( x1154 & ~n27181 ) ;
  assign n27210 = x660 | n27138 ;
  assign n27211 = ( x609 & x1155 ) | ( x609 & ~n27180 ) | ( x1155 & ~n27180 ) ;
  assign n27212 = n14839 | n27171 ;
  assign n27213 = x625 & ~n27212 ;
  assign n27214 = n27134 & n27212 ;
  assign n27215 = n27213 | n27214 ;
  assign n27216 = n27176 & n27215 ;
  assign n27217 = x608 | n27175 ;
  assign n27218 = n27216 | n27217 ;
  assign n27219 = x1153 & n27134 ;
  assign n27220 = ~n27213 & n27219 ;
  assign n27221 = x608 & ~n27177 ;
  assign n27222 = ~n27220 & n27221 ;
  assign n27223 = n27218 & ~n27222 ;
  assign n27224 = x778 & ~n27223 ;
  assign n27225 = x778 | n27214 ;
  assign n27226 = ~n27224 & n27225 ;
  assign n27227 = ( x609 & ~x1155 ) | ( x609 & n27226 ) | ( ~x1155 & n27226 ) ;
  assign n27228 = ~n27211 & n27227 ;
  assign n27229 = n27210 | n27228 ;
  assign n27230 = x660 & ~n27140 ;
  assign n27231 = ( x609 & x1155 ) | ( x609 & n27180 ) | ( x1155 & n27180 ) ;
  assign n27232 = ( ~x609 & x1155 ) | ( ~x609 & n27226 ) | ( x1155 & n27226 ) ;
  assign n27233 = n27231 & n27232 ;
  assign n27234 = n27230 & ~n27233 ;
  assign n27235 = n27229 & ~n27234 ;
  assign n27236 = x785 & ~n27235 ;
  assign n27237 = x785 | n27226 ;
  assign n27238 = ~n27236 & n27237 ;
  assign n27239 = ( x618 & ~x1154 ) | ( x618 & n27238 ) | ( ~x1154 & n27238 ) ;
  assign n27240 = ~n27209 & n27239 ;
  assign n27241 = n27208 | n27240 ;
  assign n27242 = x627 & ~n27148 ;
  assign n27243 = ( x618 & x1154 ) | ( x618 & n27181 ) | ( x1154 & n27181 ) ;
  assign n27244 = ( ~x618 & x1154 ) | ( ~x618 & n27238 ) | ( x1154 & n27238 ) ;
  assign n27245 = n27243 & n27244 ;
  assign n27246 = n27242 & ~n27245 ;
  assign n27247 = n27241 & ~n27246 ;
  assign n27248 = x781 & ~n27247 ;
  assign n27249 = x781 | n27238 ;
  assign n27250 = ~n27248 & n27249 ;
  assign n27251 = ( ~x619 & x1159 ) | ( ~x619 & n27250 ) | ( x1159 & n27250 ) ;
  assign n27252 = n27207 & n27251 ;
  assign n27253 = n27206 & ~n27252 ;
  assign n27254 = x648 | n27155 ;
  assign n27255 = ( x619 & x1159 ) | ( x619 & ~n27182 ) | ( x1159 & ~n27182 ) ;
  assign n27256 = ( x619 & ~x1159 ) | ( x619 & n27250 ) | ( ~x1159 & n27250 ) ;
  assign n27257 = ~n27255 & n27256 ;
  assign n27258 = n27254 | n27257 ;
  assign n27259 = x789 & n27258 ;
  assign n27260 = ~n27253 & n27259 ;
  assign n27261 = ~x789 & n27250 ;
  assign n27262 = n16177 | n27261 ;
  assign n27263 = n27260 | n27262 ;
  assign n27264 = ~n27205 & n27263 ;
  assign n27265 = n18434 | n27264 ;
  assign n27266 = n16650 | n27184 ;
  assign n27267 = n16051 & ~n27164 ;
  assign n27268 = n27266 & ~n27267 ;
  assign n27269 = ( x629 & ~x792 ) | ( x629 & n27268 ) | ( ~x792 & n27268 ) ;
  assign n27270 = n16052 & ~n27164 ;
  assign n27271 = n16643 & ~n27184 ;
  assign n27272 = n27270 | n27271 ;
  assign n27273 = ( x629 & x792 ) | ( x629 & n27272 ) | ( x792 & n27272 ) ;
  assign n27274 = ~n27269 & n27273 ;
  assign n27275 = n18431 | n27274 ;
  assign n27276 = n27265 & ~n27275 ;
  assign n27277 = n27195 | n27276 ;
  assign n27278 = ( x790 & x832 ) | ( x790 & n27277 ) | ( x832 & n27277 ) ;
  assign n27279 = n15141 | n27167 ;
  assign n27280 = n15141 & ~n27132 ;
  assign n27281 = n27279 & ~n27280 ;
  assign n27282 = ( x644 & x715 ) | ( x644 & ~n27281 ) | ( x715 & ~n27281 ) ;
  assign n27283 = ( x644 & ~x715 ) | ( x644 & n27132 ) | ( ~x715 & n27132 ) ;
  assign n27284 = ~n27282 & n27283 ;
  assign n27285 = x1160 & ~n27284 ;
  assign n27286 = ~x787 & n27185 ;
  assign n27287 = x1157 & n27191 ;
  assign n27288 = n27187 | n27287 ;
  assign n27289 = x787 & n27288 ;
  assign n27290 = n27286 | n27289 ;
  assign n27291 = ( x644 & x715 ) | ( x644 & n27290 ) | ( x715 & n27290 ) ;
  assign n27292 = ( ~x644 & x715 ) | ( ~x644 & n27277 ) | ( x715 & n27277 ) ;
  assign n27293 = n27291 & n27292 ;
  assign n27294 = n27285 & ~n27293 ;
  assign n27295 = ( x644 & x715 ) | ( x644 & n27281 ) | ( x715 & n27281 ) ;
  assign n27296 = ( ~x644 & x715 ) | ( ~x644 & n27132 ) | ( x715 & n27132 ) ;
  assign n27297 = n27295 & n27296 ;
  assign n27298 = x1160 | n27297 ;
  assign n27299 = ( x644 & x715 ) | ( x644 & ~n27290 ) | ( x715 & ~n27290 ) ;
  assign n27300 = ( x644 & ~x715 ) | ( x644 & n27277 ) | ( ~x715 & n27277 ) ;
  assign n27301 = ~n27299 & n27300 ;
  assign n27302 = n27298 | n27301 ;
  assign n27303 = ~n27294 & n27302 ;
  assign n27304 = ( ~x790 & x832 ) | ( ~x790 & n27303 ) | ( x832 & n27303 ) ;
  assign n27305 = n27278 & n27304 ;
  assign n27306 = n27131 | n27305 ;
  assign n27307 = x188 | n14834 ;
  assign n27308 = n15141 & n27307 ;
  assign n27309 = x188 & n2032 ;
  assign n27310 = x768 | n17421 ;
  assign n27311 = ~n20256 & n27310 ;
  assign n27312 = x188 | n27311 ;
  assign n27313 = x188 | n17415 ;
  assign n27314 = ~x768 & n27313 ;
  assign n27315 = n22415 & n27314 ;
  assign n27316 = n27312 & ~n27315 ;
  assign n27317 = ~n2032 & n27316 ;
  assign n27318 = n27309 | n27317 ;
  assign n27319 = ~n15082 & n27318 ;
  assign n27320 = n15082 & n27307 ;
  assign n27321 = n27319 | n27320 ;
  assign n27322 = ~x785 & n27321 ;
  assign n27323 = ~n15088 & n27307 ;
  assign n27324 = x609 & n27319 ;
  assign n27325 = n27323 | n27324 ;
  assign n27326 = x1155 & n27325 ;
  assign n27327 = n15094 & n27307 ;
  assign n27328 = ~x609 & n27319 ;
  assign n27329 = n27327 | n27328 ;
  assign n27330 = ~x1155 & n27329 ;
  assign n27331 = n27326 | n27330 ;
  assign n27332 = x785 & n27331 ;
  assign n27333 = n27322 | n27332 ;
  assign n27334 = ~x781 & n27333 ;
  assign n27335 = ( x618 & x1154 ) | ( x618 & n27307 ) | ( x1154 & n27307 ) ;
  assign n27336 = ( ~x618 & x1154 ) | ( ~x618 & n27333 ) | ( x1154 & n27333 ) ;
  assign n27337 = n27335 & n27336 ;
  assign n27338 = ( x618 & x1154 ) | ( x618 & ~n27307 ) | ( x1154 & ~n27307 ) ;
  assign n27339 = ( x618 & ~x1154 ) | ( x618 & n27333 ) | ( ~x1154 & n27333 ) ;
  assign n27340 = ~n27338 & n27339 ;
  assign n27341 = n27337 | n27340 ;
  assign n27342 = x781 & n27341 ;
  assign n27343 = n27334 | n27342 ;
  assign n27344 = ~x789 & n27343 ;
  assign n27345 = ( x619 & x1159 ) | ( x619 & n27307 ) | ( x1159 & n27307 ) ;
  assign n27346 = ( ~x619 & x1159 ) | ( ~x619 & n27343 ) | ( x1159 & n27343 ) ;
  assign n27347 = n27345 & n27346 ;
  assign n27348 = ( x619 & x1159 ) | ( x619 & ~n27307 ) | ( x1159 & ~n27307 ) ;
  assign n27349 = ( x619 & ~x1159 ) | ( x619 & n27343 ) | ( ~x1159 & n27343 ) ;
  assign n27350 = ~n27348 & n27349 ;
  assign n27351 = n27347 | n27350 ;
  assign n27352 = x789 & n27351 ;
  assign n27353 = n27344 | n27352 ;
  assign n27354 = n16176 | n27353 ;
  assign n27355 = n16176 & ~n27307 ;
  assign n27356 = n27354 & ~n27355 ;
  assign n27357 = n15134 | n27356 ;
  assign n27358 = n15134 & ~n27307 ;
  assign n27359 = n27357 & ~n27358 ;
  assign n27360 = ~n15141 & n27359 ;
  assign n27361 = n27308 | n27360 ;
  assign n27362 = ( x644 & x715 ) | ( x644 & n27361 ) | ( x715 & n27361 ) ;
  assign n27363 = ( ~x644 & x715 ) | ( ~x644 & n27307 ) | ( x715 & n27307 ) ;
  assign n27364 = n27362 & n27363 ;
  assign n27365 = x1160 | n27364 ;
  assign n27366 = n15414 & n27307 ;
  assign n27367 = x188 | n15070 ;
  assign n27368 = n15375 & n27367 ;
  assign n27369 = x705 & ~n27368 ;
  assign n27370 = ( ~x38 & x188 ) | ( ~x38 & n16319 ) | ( x188 & n16319 ) ;
  assign n27371 = ( x38 & x188 ) | ( x38 & n16323 ) | ( x188 & n16323 ) ;
  assign n27372 = n27370 & ~n27371 ;
  assign n27373 = n27369 & ~n27372 ;
  assign n27374 = x188 | x705 ;
  assign n27375 = n15382 | n27374 ;
  assign n27376 = ~n2032 & n27375 ;
  assign n27377 = ~n27373 & n27376 ;
  assign n27378 = n27309 | n27377 ;
  assign n27379 = ~x778 & n27378 ;
  assign n27380 = ( x625 & x1153 ) | ( x625 & n27307 ) | ( x1153 & n27307 ) ;
  assign n27381 = ( ~x625 & x1153 ) | ( ~x625 & n27378 ) | ( x1153 & n27378 ) ;
  assign n27382 = n27380 & n27381 ;
  assign n27383 = ( x625 & x1153 ) | ( x625 & ~n27307 ) | ( x1153 & ~n27307 ) ;
  assign n27384 = ( x625 & ~x1153 ) | ( x625 & n27378 ) | ( ~x1153 & n27378 ) ;
  assign n27385 = ~n27383 & n27384 ;
  assign n27386 = n27382 | n27385 ;
  assign n27387 = x778 & n27386 ;
  assign n27388 = n27379 | n27387 ;
  assign n27389 = ~n15400 & n27388 ;
  assign n27390 = n15400 & n27307 ;
  assign n27391 = n27389 | n27390 ;
  assign n27392 = n15407 | n27391 ;
  assign n27393 = n15407 & ~n27307 ;
  assign n27394 = n27392 & ~n27393 ;
  assign n27395 = ~n15414 & n27394 ;
  assign n27396 = n27366 | n27395 ;
  assign n27397 = n15421 | n27396 ;
  assign n27398 = n15421 & ~n27307 ;
  assign n27399 = n27397 & ~n27398 ;
  assign n27400 = ~x792 & n27399 ;
  assign n27401 = ( x628 & x1156 ) | ( x628 & n27307 ) | ( x1156 & n27307 ) ;
  assign n27402 = ( ~x628 & x1156 ) | ( ~x628 & n27399 ) | ( x1156 & n27399 ) ;
  assign n27403 = n27401 & n27402 ;
  assign n27404 = ( x628 & x1156 ) | ( x628 & ~n27307 ) | ( x1156 & ~n27307 ) ;
  assign n27405 = ( x628 & ~x1156 ) | ( x628 & n27399 ) | ( ~x1156 & n27399 ) ;
  assign n27406 = ~n27404 & n27405 ;
  assign n27407 = n27403 | n27406 ;
  assign n27408 = x792 & n27407 ;
  assign n27409 = n27400 | n27408 ;
  assign n27410 = ~x787 & n27409 ;
  assign n27411 = ( x647 & x1157 ) | ( x647 & n27307 ) | ( x1157 & n27307 ) ;
  assign n27412 = ( ~x647 & x1157 ) | ( ~x647 & n27409 ) | ( x1157 & n27409 ) ;
  assign n27413 = n27411 & n27412 ;
  assign n27414 = ( x647 & x1157 ) | ( x647 & ~n27307 ) | ( x1157 & ~n27307 ) ;
  assign n27415 = ( x647 & ~x1157 ) | ( x647 & n27409 ) | ( ~x1157 & n27409 ) ;
  assign n27416 = ~n27414 & n27415 ;
  assign n27417 = n27413 | n27416 ;
  assign n27418 = x787 & n27417 ;
  assign n27419 = n27410 | n27418 ;
  assign n27420 = ( x644 & x715 ) | ( x644 & ~n27419 ) | ( x715 & ~n27419 ) ;
  assign n27421 = x630 | n27413 ;
  assign n27422 = ( x647 & x1157 ) | ( x647 & ~n27359 ) | ( x1157 & ~n27359 ) ;
  assign n27423 = x629 | n27403 ;
  assign n27424 = ( x628 & x1156 ) | ( x628 & ~n27356 ) | ( x1156 & ~n27356 ) ;
  assign n27425 = x648 | n27347 ;
  assign n27426 = ( x619 & x1159 ) | ( x619 & ~n27394 ) | ( x1159 & ~n27394 ) ;
  assign n27427 = x627 | n27337 ;
  assign n27428 = ( x618 & x1154 ) | ( x618 & ~n27391 ) | ( x1154 & ~n27391 ) ;
  assign n27429 = x660 | n27326 ;
  assign n27430 = ( x609 & x1155 ) | ( x609 & ~n27388 ) | ( x1155 & ~n27388 ) ;
  assign n27431 = x608 | n27382 ;
  assign n27432 = ( x625 & x1153 ) | ( x625 & ~n27318 ) | ( x1153 & ~n27318 ) ;
  assign n27433 = x705 | n27316 ;
  assign n27434 = ( x188 & ~x768 ) | ( x188 & n17554 ) | ( ~x768 & n17554 ) ;
  assign n27435 = ( x188 & x768 ) | ( x188 & n17562 ) | ( x768 & n17562 ) ;
  assign n27436 = n27434 & ~n27435 ;
  assign n27437 = x705 & ~n27436 ;
  assign n27438 = x768 & ~n17570 ;
  assign n27439 = ( x188 & n17569 ) | ( x188 & ~n27438 ) | ( n17569 & ~n27438 ) ;
  assign n27440 = ( x188 & n17579 ) | ( x188 & n27438 ) | ( n17579 & n27438 ) ;
  assign n27441 = ~n27439 & n27440 ;
  assign n27442 = n27437 & ~n27441 ;
  assign n27443 = n2032 | n27442 ;
  assign n27444 = n27433 & ~n27443 ;
  assign n27445 = n27309 | n27444 ;
  assign n27446 = ( x625 & ~x1153 ) | ( x625 & n27445 ) | ( ~x1153 & n27445 ) ;
  assign n27447 = ~n27432 & n27446 ;
  assign n27448 = n27431 | n27447 ;
  assign n27449 = x608 & ~n27385 ;
  assign n27450 = ( x625 & x1153 ) | ( x625 & n27318 ) | ( x1153 & n27318 ) ;
  assign n27451 = ( ~x625 & x1153 ) | ( ~x625 & n27445 ) | ( x1153 & n27445 ) ;
  assign n27452 = n27450 & n27451 ;
  assign n27453 = n27449 & ~n27452 ;
  assign n27454 = n27448 & ~n27453 ;
  assign n27455 = x778 & ~n27454 ;
  assign n27456 = x778 | n27445 ;
  assign n27457 = ~n27455 & n27456 ;
  assign n27458 = ( x609 & ~x1155 ) | ( x609 & n27457 ) | ( ~x1155 & n27457 ) ;
  assign n27459 = ~n27430 & n27458 ;
  assign n27460 = n27429 | n27459 ;
  assign n27461 = x660 & ~n27330 ;
  assign n27462 = ( x609 & x1155 ) | ( x609 & n27388 ) | ( x1155 & n27388 ) ;
  assign n27463 = ( ~x609 & x1155 ) | ( ~x609 & n27457 ) | ( x1155 & n27457 ) ;
  assign n27464 = n27462 & n27463 ;
  assign n27465 = n27461 & ~n27464 ;
  assign n27466 = n27460 & ~n27465 ;
  assign n27467 = x785 & ~n27466 ;
  assign n27468 = x785 | n27457 ;
  assign n27469 = ~n27467 & n27468 ;
  assign n27470 = ( x618 & ~x1154 ) | ( x618 & n27469 ) | ( ~x1154 & n27469 ) ;
  assign n27471 = ~n27428 & n27470 ;
  assign n27472 = n27427 | n27471 ;
  assign n27473 = x627 & ~n27340 ;
  assign n27474 = ( x618 & x1154 ) | ( x618 & n27391 ) | ( x1154 & n27391 ) ;
  assign n27475 = ( ~x618 & x1154 ) | ( ~x618 & n27469 ) | ( x1154 & n27469 ) ;
  assign n27476 = n27474 & n27475 ;
  assign n27477 = n27473 & ~n27476 ;
  assign n27478 = n27472 & ~n27477 ;
  assign n27479 = x781 & ~n27478 ;
  assign n27480 = x781 | n27469 ;
  assign n27481 = ~n27479 & n27480 ;
  assign n27482 = ( x619 & ~x1159 ) | ( x619 & n27481 ) | ( ~x1159 & n27481 ) ;
  assign n27483 = ~n27426 & n27482 ;
  assign n27484 = n27425 | n27483 ;
  assign n27485 = x648 & ~n27350 ;
  assign n27486 = ( x619 & x1159 ) | ( x619 & n27394 ) | ( x1159 & n27394 ) ;
  assign n27487 = ( ~x619 & x1159 ) | ( ~x619 & n27481 ) | ( x1159 & n27481 ) ;
  assign n27488 = n27486 & n27487 ;
  assign n27489 = n27485 & ~n27488 ;
  assign n27490 = n27484 & ~n27489 ;
  assign n27491 = x789 & ~n27490 ;
  assign n27492 = x789 | n27481 ;
  assign n27493 = ~n27491 & n27492 ;
  assign n27494 = ~x788 & n27493 ;
  assign n27495 = ( x626 & x641 ) | ( x626 & ~n27353 ) | ( x641 & ~n27353 ) ;
  assign n27496 = ( x626 & ~x641 ) | ( x626 & n27307 ) | ( ~x641 & n27307 ) ;
  assign n27497 = n27495 & ~n27496 ;
  assign n27498 = x1158 | n27497 ;
  assign n27499 = ( x626 & x641 ) | ( x626 & n27396 ) | ( x641 & n27396 ) ;
  assign n27500 = ( ~x626 & x641 ) | ( ~x626 & n27493 ) | ( x641 & n27493 ) ;
  assign n27501 = n27499 | n27500 ;
  assign n27502 = ~n27498 & n27501 ;
  assign n27503 = ( x626 & x641 ) | ( x626 & n27353 ) | ( x641 & n27353 ) ;
  assign n27504 = ( ~x626 & x641 ) | ( ~x626 & n27307 ) | ( x641 & n27307 ) ;
  assign n27505 = n27503 | n27504 ;
  assign n27506 = x1158 & n27505 ;
  assign n27507 = ( x626 & x641 ) | ( x626 & ~n27396 ) | ( x641 & ~n27396 ) ;
  assign n27508 = ( x626 & ~x641 ) | ( x626 & n27493 ) | ( ~x641 & n27493 ) ;
  assign n27509 = n27507 & ~n27508 ;
  assign n27510 = n27506 & ~n27509 ;
  assign n27511 = n27502 | n27510 ;
  assign n27512 = x788 & n27511 ;
  assign n27513 = n27494 | n27512 ;
  assign n27514 = ( x628 & ~x1156 ) | ( x628 & n27513 ) | ( ~x1156 & n27513 ) ;
  assign n27515 = ~n27424 & n27514 ;
  assign n27516 = n27423 | n27515 ;
  assign n27517 = x629 & ~n27406 ;
  assign n27518 = ( x628 & x1156 ) | ( x628 & n27356 ) | ( x1156 & n27356 ) ;
  assign n27519 = ( ~x628 & x1156 ) | ( ~x628 & n27513 ) | ( x1156 & n27513 ) ;
  assign n27520 = n27518 & n27519 ;
  assign n27521 = n27517 & ~n27520 ;
  assign n27522 = n27516 & ~n27521 ;
  assign n27523 = x792 & ~n27522 ;
  assign n27524 = x792 | n27513 ;
  assign n27525 = ~n27523 & n27524 ;
  assign n27526 = ( x647 & ~x1157 ) | ( x647 & n27525 ) | ( ~x1157 & n27525 ) ;
  assign n27527 = ~n27422 & n27526 ;
  assign n27528 = n27421 | n27527 ;
  assign n27529 = x630 & ~n27416 ;
  assign n27530 = ( x647 & x1157 ) | ( x647 & n27359 ) | ( x1157 & n27359 ) ;
  assign n27531 = ( ~x647 & x1157 ) | ( ~x647 & n27525 ) | ( x1157 & n27525 ) ;
  assign n27532 = n27530 & n27531 ;
  assign n27533 = n27529 & ~n27532 ;
  assign n27534 = n27528 & ~n27533 ;
  assign n27535 = x787 & ~n27534 ;
  assign n27536 = x787 | n27525 ;
  assign n27537 = ~n27535 & n27536 ;
  assign n27538 = ( x644 & ~x715 ) | ( x644 & n27537 ) | ( ~x715 & n27537 ) ;
  assign n27539 = ~n27420 & n27538 ;
  assign n27540 = n27365 | n27539 ;
  assign n27541 = ( x644 & x715 ) | ( x644 & ~n27361 ) | ( x715 & ~n27361 ) ;
  assign n27542 = ( x644 & ~x715 ) | ( x644 & n27307 ) | ( ~x715 & n27307 ) ;
  assign n27543 = ~n27541 & n27542 ;
  assign n27544 = x1160 & ~n27543 ;
  assign n27545 = ( x644 & x715 ) | ( x644 & n27419 ) | ( x715 & n27419 ) ;
  assign n27546 = ( ~x644 & x715 ) | ( ~x644 & n27537 ) | ( x715 & n27537 ) ;
  assign n27547 = n27545 & n27546 ;
  assign n27548 = n27544 & ~n27547 ;
  assign n27549 = x790 & ~n27548 ;
  assign n27550 = n27540 & n27549 ;
  assign n27551 = ~x790 & n27537 ;
  assign n27552 = n6785 | n27551 ;
  assign n27553 = n27550 | n27552 ;
  assign n27554 = ~x188 & n6785 ;
  assign n27555 = x832 | n27554 ;
  assign n27556 = n27553 & ~n27555 ;
  assign n27557 = x188 | n1290 ;
  assign n27558 = ~x768 & n14840 ;
  assign n27559 = n27557 & ~n27558 ;
  assign n27560 = n16060 | n27559 ;
  assign n27561 = ~x785 & n27560 ;
  assign n27562 = n16065 | n27559 ;
  assign n27563 = x1155 & n27562 ;
  assign n27564 = n16068 | n27560 ;
  assign n27565 = ~x1155 & n27564 ;
  assign n27566 = n27563 | n27565 ;
  assign n27567 = x785 & n27566 ;
  assign n27568 = n27561 | n27567 ;
  assign n27569 = ~x781 & n27568 ;
  assign n27570 = n16075 | n27568 ;
  assign n27571 = x1154 & n27570 ;
  assign n27572 = n16078 | n27568 ;
  assign n27573 = ~x1154 & n27572 ;
  assign n27574 = n27571 | n27573 ;
  assign n27575 = x781 & n27574 ;
  assign n27576 = n27569 | n27575 ;
  assign n27577 = ~x789 & n27576 ;
  assign n27578 = ( x619 & x1159 ) | ( x619 & n27557 ) | ( x1159 & n27557 ) ;
  assign n27579 = ( ~x619 & x1159 ) | ( ~x619 & n27576 ) | ( x1159 & n27576 ) ;
  assign n27580 = n27578 & n27579 ;
  assign n27581 = ( x619 & x1159 ) | ( x619 & ~n27557 ) | ( x1159 & ~n27557 ) ;
  assign n27582 = ( x619 & ~x1159 ) | ( x619 & n27576 ) | ( ~x1159 & n27576 ) ;
  assign n27583 = ~n27581 & n27582 ;
  assign n27584 = n27580 | n27583 ;
  assign n27585 = x789 & n27584 ;
  assign n27586 = n27577 | n27585 ;
  assign n27587 = n16176 | n27586 ;
  assign n27588 = n16176 & ~n27557 ;
  assign n27589 = n27587 & ~n27588 ;
  assign n27590 = n15134 | n27589 ;
  assign n27591 = n15134 & ~n27557 ;
  assign n27592 = n27590 & ~n27591 ;
  assign n27593 = n18610 & n27592 ;
  assign n27594 = ( x647 & x1157 ) | ( x647 & ~n27557 ) | ( x1157 & ~n27557 ) ;
  assign n27595 = x705 & n15202 ;
  assign n27596 = n27557 & ~n27595 ;
  assign n27597 = ~x778 & n27596 ;
  assign n27598 = ~x625 & n27595 ;
  assign n27599 = n27596 | n27598 ;
  assign n27600 = x1153 & n27599 ;
  assign n27601 = ~x1153 & n27557 ;
  assign n27602 = ~n27598 & n27601 ;
  assign n27603 = n27600 | n27602 ;
  assign n27604 = x778 & n27603 ;
  assign n27605 = n27597 | n27604 ;
  assign n27606 = n16043 | n27605 ;
  assign n27607 = n16045 | n27606 ;
  assign n27608 = n16047 | n27607 ;
  assign n27609 = n16049 | n27608 ;
  assign n27610 = n16055 | n27609 ;
  assign n27611 = ( x647 & ~x1157 ) | ( x647 & n27610 ) | ( ~x1157 & n27610 ) ;
  assign n27612 = ~n27594 & n27611 ;
  assign n27613 = x630 & n27612 ;
  assign n27614 = x647 & n27610 ;
  assign n27615 = ~x647 & n27557 ;
  assign n27616 = n27614 | n27615 ;
  assign n27617 = n15138 & n27616 ;
  assign n27618 = n27613 | n27617 ;
  assign n27619 = n27593 | n27618 ;
  assign n27620 = x787 & n27619 ;
  assign n27621 = n16115 & ~n27608 ;
  assign n27622 = ( x626 & ~n15419 ) | ( x626 & n27557 ) | ( ~n15419 & n27557 ) ;
  assign n27623 = ( x626 & n15419 ) | ( x626 & ~n27586 ) | ( n15419 & ~n27586 ) ;
  assign n27624 = ~n27622 & n27623 ;
  assign n27625 = n27621 | n27624 ;
  assign n27626 = ( x626 & n15418 ) | ( x626 & ~n27557 ) | ( n15418 & ~n27557 ) ;
  assign n27627 = ( x626 & ~n15418 ) | ( x626 & n27586 ) | ( ~n15418 & n27586 ) ;
  assign n27628 = n27626 & ~n27627 ;
  assign n27629 = n27625 | n27628 ;
  assign n27630 = x788 & n27629 ;
  assign n27631 = x648 & ~n27583 ;
  assign n27632 = ( x619 & x1159 ) | ( x619 & n27607 ) | ( x1159 & n27607 ) ;
  assign n27633 = x627 | n27571 ;
  assign n27634 = ( x618 & x1154 ) | ( x618 & ~n27606 ) | ( x1154 & ~n27606 ) ;
  assign n27635 = x660 | n27563 ;
  assign n27636 = ( x609 & x1155 ) | ( x609 & ~n27605 ) | ( x1155 & ~n27605 ) ;
  assign n27637 = n14839 | n27596 ;
  assign n27638 = x625 & ~n27637 ;
  assign n27639 = n27559 & n27637 ;
  assign n27640 = n27638 | n27639 ;
  assign n27641 = n27601 & n27640 ;
  assign n27642 = x608 | n27600 ;
  assign n27643 = n27641 | n27642 ;
  assign n27644 = x1153 & n27559 ;
  assign n27645 = ~n27638 & n27644 ;
  assign n27646 = x608 & ~n27602 ;
  assign n27647 = ~n27645 & n27646 ;
  assign n27648 = n27643 & ~n27647 ;
  assign n27649 = x778 & ~n27648 ;
  assign n27650 = x778 | n27639 ;
  assign n27651 = ~n27649 & n27650 ;
  assign n27652 = ( x609 & ~x1155 ) | ( x609 & n27651 ) | ( ~x1155 & n27651 ) ;
  assign n27653 = ~n27636 & n27652 ;
  assign n27654 = n27635 | n27653 ;
  assign n27655 = x660 & ~n27565 ;
  assign n27656 = ( x609 & x1155 ) | ( x609 & n27605 ) | ( x1155 & n27605 ) ;
  assign n27657 = ( ~x609 & x1155 ) | ( ~x609 & n27651 ) | ( x1155 & n27651 ) ;
  assign n27658 = n27656 & n27657 ;
  assign n27659 = n27655 & ~n27658 ;
  assign n27660 = n27654 & ~n27659 ;
  assign n27661 = x785 & ~n27660 ;
  assign n27662 = x785 | n27651 ;
  assign n27663 = ~n27661 & n27662 ;
  assign n27664 = ( x618 & ~x1154 ) | ( x618 & n27663 ) | ( ~x1154 & n27663 ) ;
  assign n27665 = ~n27634 & n27664 ;
  assign n27666 = n27633 | n27665 ;
  assign n27667 = x627 & ~n27573 ;
  assign n27668 = ( x618 & x1154 ) | ( x618 & n27606 ) | ( x1154 & n27606 ) ;
  assign n27669 = ( ~x618 & x1154 ) | ( ~x618 & n27663 ) | ( x1154 & n27663 ) ;
  assign n27670 = n27668 & n27669 ;
  assign n27671 = n27667 & ~n27670 ;
  assign n27672 = n27666 & ~n27671 ;
  assign n27673 = x781 & ~n27672 ;
  assign n27674 = x781 | n27663 ;
  assign n27675 = ~n27673 & n27674 ;
  assign n27676 = ( ~x619 & x1159 ) | ( ~x619 & n27675 ) | ( x1159 & n27675 ) ;
  assign n27677 = n27632 & n27676 ;
  assign n27678 = n27631 & ~n27677 ;
  assign n27679 = x648 | n27580 ;
  assign n27680 = ( x619 & x1159 ) | ( x619 & ~n27607 ) | ( x1159 & ~n27607 ) ;
  assign n27681 = ( x619 & ~x1159 ) | ( x619 & n27675 ) | ( ~x1159 & n27675 ) ;
  assign n27682 = ~n27680 & n27681 ;
  assign n27683 = n27679 | n27682 ;
  assign n27684 = x789 & n27683 ;
  assign n27685 = ~n27678 & n27684 ;
  assign n27686 = ~x789 & n27675 ;
  assign n27687 = n16177 | n27686 ;
  assign n27688 = n27685 | n27687 ;
  assign n27689 = ~n27630 & n27688 ;
  assign n27690 = n18434 | n27689 ;
  assign n27691 = n16650 | n27609 ;
  assign n27692 = n16051 & ~n27589 ;
  assign n27693 = n27691 & ~n27692 ;
  assign n27694 = ( x629 & ~x792 ) | ( x629 & n27693 ) | ( ~x792 & n27693 ) ;
  assign n27695 = n16052 & ~n27589 ;
  assign n27696 = n16643 & ~n27609 ;
  assign n27697 = n27695 | n27696 ;
  assign n27698 = ( x629 & x792 ) | ( x629 & n27697 ) | ( x792 & n27697 ) ;
  assign n27699 = ~n27694 & n27698 ;
  assign n27700 = n18431 | n27699 ;
  assign n27701 = n27690 & ~n27700 ;
  assign n27702 = n27620 | n27701 ;
  assign n27703 = ( x790 & x832 ) | ( x790 & n27702 ) | ( x832 & n27702 ) ;
  assign n27704 = n15141 | n27592 ;
  assign n27705 = n15141 & ~n27557 ;
  assign n27706 = n27704 & ~n27705 ;
  assign n27707 = ( x644 & x715 ) | ( x644 & ~n27706 ) | ( x715 & ~n27706 ) ;
  assign n27708 = ( x644 & ~x715 ) | ( x644 & n27557 ) | ( ~x715 & n27557 ) ;
  assign n27709 = ~n27707 & n27708 ;
  assign n27710 = x1160 & ~n27709 ;
  assign n27711 = ~x787 & n27610 ;
  assign n27712 = x1157 & n27616 ;
  assign n27713 = n27612 | n27712 ;
  assign n27714 = x787 & n27713 ;
  assign n27715 = n27711 | n27714 ;
  assign n27716 = ( x644 & x715 ) | ( x644 & n27715 ) | ( x715 & n27715 ) ;
  assign n27717 = ( ~x644 & x715 ) | ( ~x644 & n27702 ) | ( x715 & n27702 ) ;
  assign n27718 = n27716 & n27717 ;
  assign n27719 = n27710 & ~n27718 ;
  assign n27720 = ( x644 & x715 ) | ( x644 & n27706 ) | ( x715 & n27706 ) ;
  assign n27721 = ( ~x644 & x715 ) | ( ~x644 & n27557 ) | ( x715 & n27557 ) ;
  assign n27722 = n27720 & n27721 ;
  assign n27723 = x1160 | n27722 ;
  assign n27724 = ( x644 & x715 ) | ( x644 & ~n27715 ) | ( x715 & ~n27715 ) ;
  assign n27725 = ( x644 & ~x715 ) | ( x644 & n27702 ) | ( ~x715 & n27702 ) ;
  assign n27726 = ~n27724 & n27725 ;
  assign n27727 = n27723 | n27726 ;
  assign n27728 = ~n27719 & n27727 ;
  assign n27729 = ( ~x790 & x832 ) | ( ~x790 & n27728 ) | ( x832 & n27728 ) ;
  assign n27730 = n27703 & n27729 ;
  assign n27731 = n27556 | n27730 ;
  assign n27732 = x189 & ~n14834 ;
  assign n27733 = n15141 & ~n27732 ;
  assign n27734 = n15082 & ~n27732 ;
  assign n27735 = x189 & n2032 ;
  assign n27736 = x772 & ~n15061 ;
  assign n27737 = n20169 & ~n27736 ;
  assign n27738 = x39 & ~n27737 ;
  assign n27739 = ( x39 & x772 ) | ( x39 & n14956 ) | ( x772 & n14956 ) ;
  assign n27740 = ( x39 & ~x772 ) | ( x39 & n14822 ) | ( ~x772 & n14822 ) ;
  assign n27741 = n27739 | n27740 ;
  assign n27742 = ~n27738 & n27741 ;
  assign n27743 = x189 & ~n27742 ;
  assign n27744 = ~x189 & x772 ;
  assign n27745 = n14933 & n27744 ;
  assign n27746 = n27743 | n27745 ;
  assign n27747 = ~x38 & n27746 ;
  assign n27748 = x772 & n14839 ;
  assign n27749 = n15070 & ~n27748 ;
  assign n27750 = x189 | n15070 ;
  assign n27751 = x38 & n27750 ;
  assign n27752 = ~n27749 & n27751 ;
  assign n27753 = n27747 | n27752 ;
  assign n27754 = ~n2032 & n27753 ;
  assign n27755 = n27735 | n27754 ;
  assign n27756 = n15082 | n27755 ;
  assign n27757 = ~n27734 & n27756 ;
  assign n27758 = ~x785 & n27757 ;
  assign n27759 = ( x609 & x1155 ) | ( x609 & n27732 ) | ( x1155 & n27732 ) ;
  assign n27760 = ( ~x609 & x1155 ) | ( ~x609 & n27757 ) | ( x1155 & n27757 ) ;
  assign n27761 = n27759 & n27760 ;
  assign n27762 = ( x609 & x1155 ) | ( x609 & ~n27732 ) | ( x1155 & ~n27732 ) ;
  assign n27763 = ( x609 & ~x1155 ) | ( x609 & n27757 ) | ( ~x1155 & n27757 ) ;
  assign n27764 = ~n27762 & n27763 ;
  assign n27765 = n27761 | n27764 ;
  assign n27766 = x785 & n27765 ;
  assign n27767 = n27758 | n27766 ;
  assign n27768 = ~x781 & n27767 ;
  assign n27769 = ( x618 & x1154 ) | ( x618 & n27732 ) | ( x1154 & n27732 ) ;
  assign n27770 = ( ~x618 & x1154 ) | ( ~x618 & n27767 ) | ( x1154 & n27767 ) ;
  assign n27771 = n27769 & n27770 ;
  assign n27772 = ( x618 & x1154 ) | ( x618 & ~n27732 ) | ( x1154 & ~n27732 ) ;
  assign n27773 = ( x618 & ~x1154 ) | ( x618 & n27767 ) | ( ~x1154 & n27767 ) ;
  assign n27774 = ~n27772 & n27773 ;
  assign n27775 = n27771 | n27774 ;
  assign n27776 = x781 & n27775 ;
  assign n27777 = n27768 | n27776 ;
  assign n27778 = ~x789 & n27777 ;
  assign n27779 = ( x619 & x1159 ) | ( x619 & n27732 ) | ( x1159 & n27732 ) ;
  assign n27780 = ( ~x619 & x1159 ) | ( ~x619 & n27777 ) | ( x1159 & n27777 ) ;
  assign n27781 = n27779 & n27780 ;
  assign n27782 = ( x619 & x1159 ) | ( x619 & ~n27732 ) | ( x1159 & ~n27732 ) ;
  assign n27783 = ( x619 & ~x1159 ) | ( x619 & n27777 ) | ( ~x1159 & n27777 ) ;
  assign n27784 = ~n27782 & n27783 ;
  assign n27785 = n27781 | n27784 ;
  assign n27786 = x789 & n27785 ;
  assign n27787 = n27778 | n27786 ;
  assign n27788 = ~n16176 & n27787 ;
  assign n27789 = n16176 & n27732 ;
  assign n27790 = n27788 | n27789 ;
  assign n27791 = ~n15134 & n27790 ;
  assign n27792 = n15134 & n27732 ;
  assign n27793 = n27791 | n27792 ;
  assign n27794 = n15141 | n27793 ;
  assign n27795 = ~n27733 & n27794 ;
  assign n27796 = ( x644 & x715 ) | ( x644 & n27795 ) | ( x715 & n27795 ) ;
  assign n27797 = ( ~x644 & x715 ) | ( ~x644 & n27732 ) | ( x715 & n27732 ) ;
  assign n27798 = n27796 & n27797 ;
  assign n27799 = x1160 | n27798 ;
  assign n27800 = n15414 & ~n27732 ;
  assign n27801 = n15400 & ~n27732 ;
  assign n27802 = x727 & ~n2032 ;
  assign n27803 = n27732 | n27802 ;
  assign n27804 = n17892 & n27750 ;
  assign n27805 = n27802 & ~n27804 ;
  assign n27806 = ( ~x38 & x189 ) | ( ~x38 & n16323 ) | ( x189 & n16323 ) ;
  assign n27807 = ( x38 & x189 ) | ( x38 & n16319 ) | ( x189 & n16319 ) ;
  assign n27808 = n27806 & ~n27807 ;
  assign n27809 = n27805 & ~n27808 ;
  assign n27810 = n27803 & ~n27809 ;
  assign n27811 = ~x778 & n27810 ;
  assign n27812 = ( x625 & x1153 ) | ( x625 & n27732 ) | ( x1153 & n27732 ) ;
  assign n27813 = ( ~x625 & x1153 ) | ( ~x625 & n27810 ) | ( x1153 & n27810 ) ;
  assign n27814 = n27812 & n27813 ;
  assign n27815 = ( x625 & x1153 ) | ( x625 & ~n27732 ) | ( x1153 & ~n27732 ) ;
  assign n27816 = ( x625 & ~x1153 ) | ( x625 & n27810 ) | ( ~x1153 & n27810 ) ;
  assign n27817 = ~n27815 & n27816 ;
  assign n27818 = n27814 | n27817 ;
  assign n27819 = x778 & n27818 ;
  assign n27820 = n27811 | n27819 ;
  assign n27821 = n15400 | n27820 ;
  assign n27822 = ~n27801 & n27821 ;
  assign n27823 = ~n15407 & n27822 ;
  assign n27824 = n15407 & n27732 ;
  assign n27825 = n27823 | n27824 ;
  assign n27826 = n15414 | n27825 ;
  assign n27827 = ~n27800 & n27826 ;
  assign n27828 = ~n15421 & n27827 ;
  assign n27829 = n15421 & n27732 ;
  assign n27830 = n27828 | n27829 ;
  assign n27831 = ~x792 & n27830 ;
  assign n27832 = ( x628 & x1156 ) | ( x628 & n27732 ) | ( x1156 & n27732 ) ;
  assign n27833 = ( ~x628 & x1156 ) | ( ~x628 & n27830 ) | ( x1156 & n27830 ) ;
  assign n27834 = n27832 & n27833 ;
  assign n27835 = ( x628 & x1156 ) | ( x628 & ~n27732 ) | ( x1156 & ~n27732 ) ;
  assign n27836 = ( x628 & ~x1156 ) | ( x628 & n27830 ) | ( ~x1156 & n27830 ) ;
  assign n27837 = ~n27835 & n27836 ;
  assign n27838 = n27834 | n27837 ;
  assign n27839 = x792 & n27838 ;
  assign n27840 = n27831 | n27839 ;
  assign n27841 = ~x787 & n27840 ;
  assign n27842 = ( x647 & x1157 ) | ( x647 & n27732 ) | ( x1157 & n27732 ) ;
  assign n27843 = ( ~x647 & x1157 ) | ( ~x647 & n27840 ) | ( x1157 & n27840 ) ;
  assign n27844 = n27842 & n27843 ;
  assign n27845 = ( x647 & x1157 ) | ( x647 & ~n27732 ) | ( x1157 & ~n27732 ) ;
  assign n27846 = ( x647 & ~x1157 ) | ( x647 & n27840 ) | ( ~x1157 & n27840 ) ;
  assign n27847 = ~n27845 & n27846 ;
  assign n27848 = n27844 | n27847 ;
  assign n27849 = x787 & n27848 ;
  assign n27850 = n27841 | n27849 ;
  assign n27851 = ( x644 & x715 ) | ( x644 & ~n27850 ) | ( x715 & ~n27850 ) ;
  assign n27852 = x630 | n27844 ;
  assign n27853 = ( x647 & x1157 ) | ( x647 & ~n27793 ) | ( x1157 & ~n27793 ) ;
  assign n27854 = x629 | n27834 ;
  assign n27855 = ( x628 & x1156 ) | ( x628 & ~n27790 ) | ( x1156 & ~n27790 ) ;
  assign n27856 = x648 | n27781 ;
  assign n27857 = ( x619 & x1159 ) | ( x619 & ~n27825 ) | ( x1159 & ~n27825 ) ;
  assign n27858 = x627 | n27771 ;
  assign n27859 = ( x618 & x1154 ) | ( x618 & ~n27822 ) | ( x1154 & ~n27822 ) ;
  assign n27860 = x660 | n27761 ;
  assign n27861 = ( x609 & x1155 ) | ( x609 & ~n27820 ) | ( x1155 & ~n27820 ) ;
  assign n27862 = x608 | n27814 ;
  assign n27863 = ( x625 & x1153 ) | ( x625 & ~n27755 ) | ( x1153 & ~n27755 ) ;
  assign n27864 = x727 | n27753 ;
  assign n27865 = ( x189 & ~x772 ) | ( x189 & n15797 ) | ( ~x772 & n15797 ) ;
  assign n27866 = ( x189 & x772 ) | ( x189 & n15872 ) | ( x772 & n15872 ) ;
  assign n27867 = ~n27865 & n27866 ;
  assign n27868 = x39 & ~n27867 ;
  assign n27869 = ( x189 & ~x772 ) | ( x189 & n15583 ) | ( ~x772 & n15583 ) ;
  assign n27870 = ( x189 & x772 ) | ( x189 & n15699 ) | ( x772 & n15699 ) ;
  assign n27871 = n27869 & ~n27870 ;
  assign n27872 = n27868 & ~n27871 ;
  assign n27873 = ( x189 & ~x772 ) | ( x189 & n15887 ) | ( ~x772 & n15887 ) ;
  assign n27874 = ( x189 & x772 ) | ( x189 & n15891 ) | ( x772 & n15891 ) ;
  assign n27875 = n27873 & ~n27874 ;
  assign n27876 = ( x189 & ~x772 ) | ( x189 & n15894 ) | ( ~x772 & n15894 ) ;
  assign n27877 = ( x189 & x772 ) | ( x189 & n15897 ) | ( x772 & n15897 ) ;
  assign n27878 = ~n27876 & n27877 ;
  assign n27879 = n27875 | n27878 ;
  assign n27880 = ( ~x38 & n9138 ) | ( ~x38 & n27879 ) | ( n9138 & n27879 ) ;
  assign n27881 = ~n27872 & n27880 ;
  assign n27882 = x727 & ~n17570 ;
  assign n27883 = ~n27752 & n27882 ;
  assign n27884 = ~n27881 & n27883 ;
  assign n27885 = n2032 | n27884 ;
  assign n27886 = n27864 & ~n27885 ;
  assign n27887 = n27735 | n27886 ;
  assign n27888 = ( x625 & ~x1153 ) | ( x625 & n27887 ) | ( ~x1153 & n27887 ) ;
  assign n27889 = ~n27863 & n27888 ;
  assign n27890 = n27862 | n27889 ;
  assign n27891 = x608 & ~n27817 ;
  assign n27892 = ( x625 & x1153 ) | ( x625 & n27755 ) | ( x1153 & n27755 ) ;
  assign n27893 = ( ~x625 & x1153 ) | ( ~x625 & n27887 ) | ( x1153 & n27887 ) ;
  assign n27894 = n27892 & n27893 ;
  assign n27895 = n27891 & ~n27894 ;
  assign n27896 = n27890 & ~n27895 ;
  assign n27897 = x778 & ~n27896 ;
  assign n27898 = x778 | n27887 ;
  assign n27899 = ~n27897 & n27898 ;
  assign n27900 = ( x609 & ~x1155 ) | ( x609 & n27899 ) | ( ~x1155 & n27899 ) ;
  assign n27901 = ~n27861 & n27900 ;
  assign n27902 = n27860 | n27901 ;
  assign n27903 = x660 & ~n27764 ;
  assign n27904 = ( x609 & x1155 ) | ( x609 & n27820 ) | ( x1155 & n27820 ) ;
  assign n27905 = ( ~x609 & x1155 ) | ( ~x609 & n27899 ) | ( x1155 & n27899 ) ;
  assign n27906 = n27904 & n27905 ;
  assign n27907 = n27903 & ~n27906 ;
  assign n27908 = n27902 & ~n27907 ;
  assign n27909 = x785 & ~n27908 ;
  assign n27910 = x785 | n27899 ;
  assign n27911 = ~n27909 & n27910 ;
  assign n27912 = ( x618 & ~x1154 ) | ( x618 & n27911 ) | ( ~x1154 & n27911 ) ;
  assign n27913 = ~n27859 & n27912 ;
  assign n27914 = n27858 | n27913 ;
  assign n27915 = x627 & ~n27774 ;
  assign n27916 = ( x618 & x1154 ) | ( x618 & n27822 ) | ( x1154 & n27822 ) ;
  assign n27917 = ( ~x618 & x1154 ) | ( ~x618 & n27911 ) | ( x1154 & n27911 ) ;
  assign n27918 = n27916 & n27917 ;
  assign n27919 = n27915 & ~n27918 ;
  assign n27920 = n27914 & ~n27919 ;
  assign n27921 = x781 & ~n27920 ;
  assign n27922 = x781 | n27911 ;
  assign n27923 = ~n27921 & n27922 ;
  assign n27924 = ( x619 & ~x1159 ) | ( x619 & n27923 ) | ( ~x1159 & n27923 ) ;
  assign n27925 = ~n27857 & n27924 ;
  assign n27926 = n27856 | n27925 ;
  assign n27927 = x648 & ~n27784 ;
  assign n27928 = ( x619 & x1159 ) | ( x619 & n27825 ) | ( x1159 & n27825 ) ;
  assign n27929 = ( ~x619 & x1159 ) | ( ~x619 & n27923 ) | ( x1159 & n27923 ) ;
  assign n27930 = n27928 & n27929 ;
  assign n27931 = n27927 & ~n27930 ;
  assign n27932 = n27926 & ~n27931 ;
  assign n27933 = x789 & ~n27932 ;
  assign n27934 = x789 | n27923 ;
  assign n27935 = ~n27933 & n27934 ;
  assign n27936 = ~x788 & n27935 ;
  assign n27937 = ( x626 & x641 ) | ( x626 & ~n27787 ) | ( x641 & ~n27787 ) ;
  assign n27938 = ( x626 & ~x641 ) | ( x626 & n27732 ) | ( ~x641 & n27732 ) ;
  assign n27939 = n27937 & ~n27938 ;
  assign n27940 = x1158 | n27939 ;
  assign n27941 = ( x626 & x641 ) | ( x626 & n27827 ) | ( x641 & n27827 ) ;
  assign n27942 = ( ~x626 & x641 ) | ( ~x626 & n27935 ) | ( x641 & n27935 ) ;
  assign n27943 = n27941 | n27942 ;
  assign n27944 = ~n27940 & n27943 ;
  assign n27945 = ( x626 & x641 ) | ( x626 & n27787 ) | ( x641 & n27787 ) ;
  assign n27946 = ( ~x626 & x641 ) | ( ~x626 & n27732 ) | ( x641 & n27732 ) ;
  assign n27947 = n27945 | n27946 ;
  assign n27948 = x1158 & n27947 ;
  assign n27949 = ( x626 & x641 ) | ( x626 & ~n27827 ) | ( x641 & ~n27827 ) ;
  assign n27950 = ( x626 & ~x641 ) | ( x626 & n27935 ) | ( ~x641 & n27935 ) ;
  assign n27951 = n27949 & ~n27950 ;
  assign n27952 = n27948 & ~n27951 ;
  assign n27953 = n27944 | n27952 ;
  assign n27954 = x788 & n27953 ;
  assign n27955 = n27936 | n27954 ;
  assign n27956 = ( x628 & ~x1156 ) | ( x628 & n27955 ) | ( ~x1156 & n27955 ) ;
  assign n27957 = ~n27855 & n27956 ;
  assign n27958 = n27854 | n27957 ;
  assign n27959 = x629 & ~n27837 ;
  assign n27960 = ( x628 & x1156 ) | ( x628 & n27790 ) | ( x1156 & n27790 ) ;
  assign n27961 = ( ~x628 & x1156 ) | ( ~x628 & n27955 ) | ( x1156 & n27955 ) ;
  assign n27962 = n27960 & n27961 ;
  assign n27963 = n27959 & ~n27962 ;
  assign n27964 = n27958 & ~n27963 ;
  assign n27965 = x792 & ~n27964 ;
  assign n27966 = x792 | n27955 ;
  assign n27967 = ~n27965 & n27966 ;
  assign n27968 = ( x647 & ~x1157 ) | ( x647 & n27967 ) | ( ~x1157 & n27967 ) ;
  assign n27969 = ~n27853 & n27968 ;
  assign n27970 = n27852 | n27969 ;
  assign n27971 = x630 & ~n27847 ;
  assign n27972 = ( x647 & x1157 ) | ( x647 & n27793 ) | ( x1157 & n27793 ) ;
  assign n27973 = ( ~x647 & x1157 ) | ( ~x647 & n27967 ) | ( x1157 & n27967 ) ;
  assign n27974 = n27972 & n27973 ;
  assign n27975 = n27971 & ~n27974 ;
  assign n27976 = n27970 & ~n27975 ;
  assign n27977 = x787 & ~n27976 ;
  assign n27978 = x787 | n27967 ;
  assign n27979 = ~n27977 & n27978 ;
  assign n27980 = ( x644 & ~x715 ) | ( x644 & n27979 ) | ( ~x715 & n27979 ) ;
  assign n27981 = ~n27851 & n27980 ;
  assign n27982 = n27799 | n27981 ;
  assign n27983 = ( x644 & x715 ) | ( x644 & ~n27795 ) | ( x715 & ~n27795 ) ;
  assign n27984 = ( x644 & ~x715 ) | ( x644 & n27732 ) | ( ~x715 & n27732 ) ;
  assign n27985 = ~n27983 & n27984 ;
  assign n27986 = x1160 & ~n27985 ;
  assign n27987 = ( x644 & x715 ) | ( x644 & n27850 ) | ( x715 & n27850 ) ;
  assign n27988 = ( ~x644 & x715 ) | ( ~x644 & n27979 ) | ( x715 & n27979 ) ;
  assign n27989 = n27987 & n27988 ;
  assign n27990 = n27986 & ~n27989 ;
  assign n27991 = x790 & ~n27990 ;
  assign n27992 = n27982 & n27991 ;
  assign n27993 = ~x790 & n27979 ;
  assign n27994 = n4832 | n27993 ;
  assign n27995 = n27992 | n27994 ;
  assign n27996 = ~x189 & n4832 ;
  assign n27997 = x57 | n27996 ;
  assign n27998 = n27995 & ~n27997 ;
  assign n27999 = x57 & x189 ;
  assign n28000 = x832 | n27999 ;
  assign n28001 = n27998 | n28000 ;
  assign n28002 = x189 & ~n1290 ;
  assign n28003 = x727 & n15202 ;
  assign n28004 = n28002 | n28003 ;
  assign n28005 = x778 | n28004 ;
  assign n28006 = x625 & n28003 ;
  assign n28007 = x1153 & ~n28002 ;
  assign n28008 = ~n28006 & n28007 ;
  assign n28009 = n28004 & ~n28006 ;
  assign n28010 = x1153 | n28009 ;
  assign n28011 = ~n28008 & n28010 ;
  assign n28012 = x778 & ~n28011 ;
  assign n28013 = n28005 & ~n28012 ;
  assign n28014 = ~n17214 & n28013 ;
  assign n28015 = n21632 & ~n28014 ;
  assign n28016 = x772 & n14840 ;
  assign n28017 = ~n18257 & n28016 ;
  assign n28018 = ~n18249 & n28017 ;
  assign n28019 = ~n18302 & n28018 ;
  assign n28020 = n15412 & ~n28019 ;
  assign n28021 = n18383 & n28018 ;
  assign n28022 = n15411 & ~n28021 ;
  assign n28023 = n28020 | n28022 ;
  assign n28024 = n28015 | n28023 ;
  assign n28025 = x789 & ~n28002 ;
  assign n28026 = n28024 & n28025 ;
  assign n28027 = n16177 | n28026 ;
  assign n28028 = ~n15400 & n28013 ;
  assign n28029 = n28002 | n28028 ;
  assign n28030 = ( x618 & x1154 ) | ( x618 & ~n28029 ) | ( x1154 & ~n28029 ) ;
  assign n28031 = ( x609 & x1155 ) | ( x609 & n28013 ) | ( x1155 & n28013 ) ;
  assign n28032 = n28002 | n28016 ;
  assign n28033 = x727 & n15529 ;
  assign n28034 = n28032 | n28033 ;
  assign n28035 = x625 & n28033 ;
  assign n28036 = n28034 & ~n28035 ;
  assign n28037 = x1153 | n28036 ;
  assign n28038 = x608 | n28008 ;
  assign n28039 = n28037 & ~n28038 ;
  assign n28040 = x1153 & ~n28032 ;
  assign n28041 = ~n28035 & n28040 ;
  assign n28042 = x608 & n28010 ;
  assign n28043 = ~n28041 & n28042 ;
  assign n28044 = n28039 | n28043 ;
  assign n28045 = x778 & n28044 ;
  assign n28046 = ~x778 & n28034 ;
  assign n28047 = n28045 | n28046 ;
  assign n28048 = ( ~x609 & x1155 ) | ( ~x609 & n28047 ) | ( x1155 & n28047 ) ;
  assign n28049 = n28031 | n28048 ;
  assign n28050 = n15088 & n28016 ;
  assign n28051 = n28002 | n28050 ;
  assign n28052 = ( x660 & n15397 ) | ( x660 & ~n28051 ) | ( n15397 & ~n28051 ) ;
  assign n28053 = n28049 & ~n28052 ;
  assign n28054 = ( x609 & x1155 ) | ( x609 & ~n28013 ) | ( x1155 & ~n28013 ) ;
  assign n28055 = ( x609 & ~x1155 ) | ( x609 & n28047 ) | ( ~x1155 & n28047 ) ;
  assign n28056 = n28054 & ~n28055 ;
  assign n28057 = ~n15094 & n28016 ;
  assign n28058 = n28002 | n28057 ;
  assign n28059 = ( x660 & n15398 ) | ( x660 & n28058 ) | ( n15398 & n28058 ) ;
  assign n28060 = ~n28056 & n28059 ;
  assign n28061 = n28053 | n28060 ;
  assign n28062 = x785 & n28061 ;
  assign n28063 = ~x785 & n28047 ;
  assign n28064 = n28062 | n28063 ;
  assign n28065 = ( x618 & ~x1154 ) | ( x618 & n28064 ) | ( ~x1154 & n28064 ) ;
  assign n28066 = n28030 & ~n28065 ;
  assign n28067 = ~n18366 & n28017 ;
  assign n28068 = n28002 | n28067 ;
  assign n28069 = ( x627 & n15405 ) | ( x627 & n28068 ) | ( n15405 & n28068 ) ;
  assign n28070 = ~n28066 & n28069 ;
  assign n28071 = ( x618 & x1154 ) | ( x618 & n28029 ) | ( x1154 & n28029 ) ;
  assign n28072 = ( ~x618 & x1154 ) | ( ~x618 & n28064 ) | ( x1154 & n28064 ) ;
  assign n28073 = n28071 | n28072 ;
  assign n28074 = n18315 & n28017 ;
  assign n28075 = n28002 | n28074 ;
  assign n28076 = ( x627 & n15404 ) | ( x627 & ~n28075 ) | ( n15404 & ~n28075 ) ;
  assign n28077 = n28073 & ~n28076 ;
  assign n28078 = n28070 | n28077 ;
  assign n28079 = ( x781 & n21647 ) | ( x781 & n28078 ) | ( n21647 & n28078 ) ;
  assign n28080 = ( ~x781 & n21647 ) | ( ~x781 & n28064 ) | ( n21647 & n28064 ) ;
  assign n28081 = n28079 | n28080 ;
  assign n28082 = ~n28027 & n28081 ;
  assign n28083 = ~n15414 & n28014 ;
  assign n28084 = n28002 | n28083 ;
  assign n28085 = n16110 & n28084 ;
  assign n28086 = ~n18255 & n28017 ;
  assign n28087 = x626 & n28086 ;
  assign n28088 = n28002 | n28087 ;
  assign n28089 = x1158 & n28088 ;
  assign n28090 = x641 | n28089 ;
  assign n28091 = n28085 | n28090 ;
  assign n28092 = n16109 & n28084 ;
  assign n28093 = ~x626 & n28086 ;
  assign n28094 = n28002 | n28093 ;
  assign n28095 = ~x1158 & n28094 ;
  assign n28096 = x641 & ~n28095 ;
  assign n28097 = ~n28092 & n28096 ;
  assign n28098 = x788 & ~n28097 ;
  assign n28099 = n28091 & n28098 ;
  assign n28100 = n18434 | n28099 ;
  assign n28101 = n28082 | n28100 ;
  assign n28102 = ~n17215 & n28013 ;
  assign n28103 = x629 & ~n28102 ;
  assign n28104 = ~n16176 & n28086 ;
  assign n28105 = ( x628 & n18420 ) | ( x628 & ~n28104 ) | ( n18420 & ~n28104 ) ;
  assign n28106 = n28103 | n28105 ;
  assign n28107 = ~x1156 & n28106 ;
  assign n28108 = x628 & n28102 ;
  assign n28109 = x628 | n28104 ;
  assign n28110 = x629 & n28109 ;
  assign n28111 = x1156 & ~n28110 ;
  assign n28112 = ~n28108 & n28111 ;
  assign n28113 = n28107 | n28112 ;
  assign n28114 = x792 & ~n28002 ;
  assign n28115 = n28113 & n28114 ;
  assign n28116 = n28101 & ~n28115 ;
  assign n28117 = n18431 | n28116 ;
  assign n28118 = ~n15134 & n28104 ;
  assign n28119 = ~x630 & n28118 ;
  assign n28120 = ~n17220 & n28102 ;
  assign n28121 = x630 & ~n28120 ;
  assign n28122 = ( x647 & ~n28119 ) | ( x647 & n28121 ) | ( ~n28119 & n28121 ) ;
  assign n28123 = ~x1157 & n28122 ;
  assign n28124 = x630 | n28120 ;
  assign n28125 = x647 & n28124 ;
  assign n28126 = x630 & n28118 ;
  assign n28127 = x1157 & ~n28126 ;
  assign n28128 = ~n28125 & n28127 ;
  assign n28129 = n28123 | n28128 ;
  assign n28130 = x787 & ~n28002 ;
  assign n28131 = n28129 & n28130 ;
  assign n28132 = n28117 & ~n28131 ;
  assign n28133 = ( x790 & x832 ) | ( x790 & ~n28132 ) | ( x832 & ~n28132 ) ;
  assign n28134 = n16176 | n18264 ;
  assign n28135 = n28086 & ~n28134 ;
  assign n28136 = x644 & n28135 ;
  assign n28137 = x715 | n28002 ;
  assign n28138 = n28136 | n28137 ;
  assign n28139 = x1160 & n28138 ;
  assign n28140 = ~n17389 & n28120 ;
  assign n28141 = n28002 | n28140 ;
  assign n28142 = ( x644 & x715 ) | ( x644 & ~n28141 ) | ( x715 & ~n28141 ) ;
  assign n28143 = ( x644 & ~x715 ) | ( x644 & n28132 ) | ( ~x715 & n28132 ) ;
  assign n28144 = n28142 & ~n28143 ;
  assign n28145 = n28139 & ~n28144 ;
  assign n28146 = ~x644 & n28135 ;
  assign n28147 = x715 & ~n28002 ;
  assign n28148 = ~n28146 & n28147 ;
  assign n28149 = x1160 | n28148 ;
  assign n28150 = ( x644 & x715 ) | ( x644 & n28141 ) | ( x715 & n28141 ) ;
  assign n28151 = ( ~x644 & x715 ) | ( ~x644 & n28132 ) | ( x715 & n28132 ) ;
  assign n28152 = n28150 | n28151 ;
  assign n28153 = ~n28149 & n28152 ;
  assign n28154 = n28145 | n28153 ;
  assign n28155 = ( x790 & ~x832 ) | ( x790 & n28154 ) | ( ~x832 & n28154 ) ;
  assign n28156 = n28133 & ~n28155 ;
  assign n28157 = n28001 & ~n28156 ;
  assign n28158 = x190 | n1290 ;
  assign n28159 = x763 & n14840 ;
  assign n28160 = n28158 & ~n28159 ;
  assign n28161 = n16060 | n28160 ;
  assign n28162 = ~x785 & n28161 ;
  assign n28163 = ~n15094 & n28159 ;
  assign n28164 = n28161 | n28163 ;
  assign n28165 = x1155 & n28164 ;
  assign n28166 = ~x1155 & n28158 ;
  assign n28167 = ~n28163 & n28166 ;
  assign n28168 = n28165 | n28167 ;
  assign n28169 = x785 & n28168 ;
  assign n28170 = n28162 | n28169 ;
  assign n28171 = ~x781 & n28170 ;
  assign n28172 = n16075 | n28170 ;
  assign n28173 = x1154 & n28172 ;
  assign n28174 = n16078 | n28170 ;
  assign n28175 = ~x1154 & n28174 ;
  assign n28176 = n28173 | n28175 ;
  assign n28177 = x781 & n28176 ;
  assign n28178 = n28171 | n28177 ;
  assign n28179 = ~x789 & n28178 ;
  assign n28180 = n20948 | n28178 ;
  assign n28181 = x1159 & n28180 ;
  assign n28182 = n20951 | n28178 ;
  assign n28183 = ~x1159 & n28182 ;
  assign n28184 = n28181 | n28183 ;
  assign n28185 = x789 & n28184 ;
  assign n28186 = n28179 | n28185 ;
  assign n28187 = n16176 | n28186 ;
  assign n28188 = n16176 & ~n28158 ;
  assign n28189 = n28187 & ~n28188 ;
  assign n28190 = n15134 | n28189 ;
  assign n28191 = n15134 & ~n28158 ;
  assign n28192 = n28190 & ~n28191 ;
  assign n28193 = n18610 & n28192 ;
  assign n28194 = ( x647 & x1157 ) | ( x647 & ~n28158 ) | ( x1157 & ~n28158 ) ;
  assign n28195 = x699 & n15202 ;
  assign n28196 = n28158 & ~n28195 ;
  assign n28197 = x778 | n28196 ;
  assign n28198 = ~x625 & n28195 ;
  assign n28199 = n28196 | n28198 ;
  assign n28200 = x1153 & n28199 ;
  assign n28201 = ~x1153 & n28158 ;
  assign n28202 = ~n28198 & n28201 ;
  assign n28203 = x778 & ~n28202 ;
  assign n28204 = ~n28200 & n28203 ;
  assign n28205 = n28197 & ~n28204 ;
  assign n28206 = n16043 | n28205 ;
  assign n28207 = n16045 | n28206 ;
  assign n28208 = n16047 | n28207 ;
  assign n28209 = n16049 | n28208 ;
  assign n28210 = n16055 | n28209 ;
  assign n28211 = ( x647 & ~x1157 ) | ( x647 & n28210 ) | ( ~x1157 & n28210 ) ;
  assign n28212 = ~n28194 & n28211 ;
  assign n28213 = x630 & n28212 ;
  assign n28214 = x647 & n28210 ;
  assign n28215 = ~x647 & n28158 ;
  assign n28216 = n28214 | n28215 ;
  assign n28217 = n15138 & n28216 ;
  assign n28218 = n28213 | n28217 ;
  assign n28219 = n28193 | n28218 ;
  assign n28220 = x787 & n28219 ;
  assign n28221 = n16115 & ~n28208 ;
  assign n28222 = ( x626 & ~n15419 ) | ( x626 & n28158 ) | ( ~n15419 & n28158 ) ;
  assign n28223 = ( x626 & n15419 ) | ( x626 & ~n28186 ) | ( n15419 & ~n28186 ) ;
  assign n28224 = ~n28222 & n28223 ;
  assign n28225 = n28221 | n28224 ;
  assign n28226 = ( x626 & n15418 ) | ( x626 & ~n28158 ) | ( n15418 & ~n28158 ) ;
  assign n28227 = ( x626 & ~n15418 ) | ( x626 & n28186 ) | ( ~n15418 & n28186 ) ;
  assign n28228 = n28226 & ~n28227 ;
  assign n28229 = n28225 | n28228 ;
  assign n28230 = x788 & n28229 ;
  assign n28231 = x648 & ~n28183 ;
  assign n28232 = ( x619 & x1159 ) | ( x619 & n28207 ) | ( x1159 & n28207 ) ;
  assign n28233 = x627 | n28173 ;
  assign n28234 = ( x618 & x1154 ) | ( x618 & ~n28206 ) | ( x1154 & ~n28206 ) ;
  assign n28235 = x660 | n28165 ;
  assign n28236 = ( x609 & x1155 ) | ( x609 & ~n28205 ) | ( x1155 & ~n28205 ) ;
  assign n28237 = n14839 | n28196 ;
  assign n28238 = x625 & ~n28237 ;
  assign n28239 = n28160 & n28237 ;
  assign n28240 = n28238 | n28239 ;
  assign n28241 = n28201 & n28240 ;
  assign n28242 = x608 | n28200 ;
  assign n28243 = n28241 | n28242 ;
  assign n28244 = x1153 & n28160 ;
  assign n28245 = ~n28238 & n28244 ;
  assign n28246 = x608 & ~n28202 ;
  assign n28247 = ~n28245 & n28246 ;
  assign n28248 = n28243 & ~n28247 ;
  assign n28249 = x778 & ~n28248 ;
  assign n28250 = x778 | n28239 ;
  assign n28251 = ~n28249 & n28250 ;
  assign n28252 = ( x609 & ~x1155 ) | ( x609 & n28251 ) | ( ~x1155 & n28251 ) ;
  assign n28253 = ~n28236 & n28252 ;
  assign n28254 = n28235 | n28253 ;
  assign n28255 = x660 & ~n28167 ;
  assign n28256 = ( x609 & x1155 ) | ( x609 & n28205 ) | ( x1155 & n28205 ) ;
  assign n28257 = ( ~x609 & x1155 ) | ( ~x609 & n28251 ) | ( x1155 & n28251 ) ;
  assign n28258 = n28256 & n28257 ;
  assign n28259 = n28255 & ~n28258 ;
  assign n28260 = n28254 & ~n28259 ;
  assign n28261 = x785 & ~n28260 ;
  assign n28262 = x785 | n28251 ;
  assign n28263 = ~n28261 & n28262 ;
  assign n28264 = ( x618 & ~x1154 ) | ( x618 & n28263 ) | ( ~x1154 & n28263 ) ;
  assign n28265 = ~n28234 & n28264 ;
  assign n28266 = n28233 | n28265 ;
  assign n28267 = x627 & ~n28175 ;
  assign n28268 = ( x618 & x1154 ) | ( x618 & n28206 ) | ( x1154 & n28206 ) ;
  assign n28269 = ( ~x618 & x1154 ) | ( ~x618 & n28263 ) | ( x1154 & n28263 ) ;
  assign n28270 = n28268 & n28269 ;
  assign n28271 = n28267 & ~n28270 ;
  assign n28272 = n28266 & ~n28271 ;
  assign n28273 = x781 & ~n28272 ;
  assign n28274 = x781 | n28263 ;
  assign n28275 = ~n28273 & n28274 ;
  assign n28276 = ( ~x619 & x1159 ) | ( ~x619 & n28275 ) | ( x1159 & n28275 ) ;
  assign n28277 = n28232 & n28276 ;
  assign n28278 = n28231 & ~n28277 ;
  assign n28279 = x648 | n28181 ;
  assign n28280 = ( x619 & x1159 ) | ( x619 & ~n28207 ) | ( x1159 & ~n28207 ) ;
  assign n28281 = ( x619 & ~x1159 ) | ( x619 & n28275 ) | ( ~x1159 & n28275 ) ;
  assign n28282 = ~n28280 & n28281 ;
  assign n28283 = n28279 | n28282 ;
  assign n28284 = x789 & n28283 ;
  assign n28285 = ~n28278 & n28284 ;
  assign n28286 = ~x789 & n28275 ;
  assign n28287 = n16177 | n28286 ;
  assign n28288 = n28285 | n28287 ;
  assign n28289 = ~n28230 & n28288 ;
  assign n28290 = n18434 | n28289 ;
  assign n28291 = n16650 | n28209 ;
  assign n28292 = n16051 & ~n28189 ;
  assign n28293 = n28291 & ~n28292 ;
  assign n28294 = ( x629 & ~x792 ) | ( x629 & n28293 ) | ( ~x792 & n28293 ) ;
  assign n28295 = n16052 & ~n28189 ;
  assign n28296 = n16643 & ~n28209 ;
  assign n28297 = n28295 | n28296 ;
  assign n28298 = ( x629 & x792 ) | ( x629 & n28297 ) | ( x792 & n28297 ) ;
  assign n28299 = ~n28294 & n28298 ;
  assign n28300 = n18431 | n28299 ;
  assign n28301 = n28290 & ~n28300 ;
  assign n28302 = n28220 | n28301 ;
  assign n28303 = ( x790 & x832 ) | ( x790 & n28302 ) | ( x832 & n28302 ) ;
  assign n28304 = n15141 | n28192 ;
  assign n28305 = n15141 & ~n28158 ;
  assign n28306 = n28304 & ~n28305 ;
  assign n28307 = ( x644 & x715 ) | ( x644 & ~n28306 ) | ( x715 & ~n28306 ) ;
  assign n28308 = ( x644 & ~x715 ) | ( x644 & n28158 ) | ( ~x715 & n28158 ) ;
  assign n28309 = ~n28307 & n28308 ;
  assign n28310 = x1160 & ~n28309 ;
  assign n28311 = ~x787 & n28210 ;
  assign n28312 = x1157 & n28216 ;
  assign n28313 = n28212 | n28312 ;
  assign n28314 = x787 & n28313 ;
  assign n28315 = n28311 | n28314 ;
  assign n28316 = ( x644 & x715 ) | ( x644 & n28315 ) | ( x715 & n28315 ) ;
  assign n28317 = ( ~x644 & x715 ) | ( ~x644 & n28302 ) | ( x715 & n28302 ) ;
  assign n28318 = n28316 & n28317 ;
  assign n28319 = n28310 & ~n28318 ;
  assign n28320 = ( x644 & x715 ) | ( x644 & n28306 ) | ( x715 & n28306 ) ;
  assign n28321 = ( ~x644 & x715 ) | ( ~x644 & n28158 ) | ( x715 & n28158 ) ;
  assign n28322 = n28320 & n28321 ;
  assign n28323 = x1160 | n28322 ;
  assign n28324 = ( x644 & x715 ) | ( x644 & ~n28315 ) | ( x715 & ~n28315 ) ;
  assign n28325 = ( x644 & ~x715 ) | ( x644 & n28302 ) | ( ~x715 & n28302 ) ;
  assign n28326 = ~n28324 & n28325 ;
  assign n28327 = n28323 | n28326 ;
  assign n28328 = ~n28319 & n28327 ;
  assign n28329 = ( ~x790 & x832 ) | ( ~x790 & n28328 ) | ( x832 & n28328 ) ;
  assign n28330 = n28303 & n28329 ;
  assign n28331 = x190 | n14834 ;
  assign n28332 = n15414 & n28331 ;
  assign n28333 = x190 & n2032 ;
  assign n28334 = x190 | n15070 ;
  assign n28335 = n15375 & n28334 ;
  assign n28336 = x699 & ~n28335 ;
  assign n28337 = ( ~x38 & x190 ) | ( ~x38 & n16319 ) | ( x190 & n16319 ) ;
  assign n28338 = ( x38 & x190 ) | ( x38 & n16323 ) | ( x190 & n16323 ) ;
  assign n28339 = n28337 & ~n28338 ;
  assign n28340 = n28336 & ~n28339 ;
  assign n28341 = x190 | x699 ;
  assign n28342 = n15382 | n28341 ;
  assign n28343 = ~n2032 & n28342 ;
  assign n28344 = ~n28340 & n28343 ;
  assign n28345 = n28333 | n28344 ;
  assign n28346 = ~x778 & n28345 ;
  assign n28347 = ( x625 & x1153 ) | ( x625 & n28331 ) | ( x1153 & n28331 ) ;
  assign n28348 = ( ~x625 & x1153 ) | ( ~x625 & n28345 ) | ( x1153 & n28345 ) ;
  assign n28349 = n28347 & n28348 ;
  assign n28350 = ( x625 & x1153 ) | ( x625 & ~n28331 ) | ( x1153 & ~n28331 ) ;
  assign n28351 = ( x625 & ~x1153 ) | ( x625 & n28345 ) | ( ~x1153 & n28345 ) ;
  assign n28352 = ~n28350 & n28351 ;
  assign n28353 = n28349 | n28352 ;
  assign n28354 = x778 & n28353 ;
  assign n28355 = n28346 | n28354 ;
  assign n28356 = ~n15400 & n28355 ;
  assign n28357 = n15400 & n28331 ;
  assign n28358 = n28356 | n28357 ;
  assign n28359 = n15407 | n28358 ;
  assign n28360 = n15407 & ~n28331 ;
  assign n28361 = n28359 & ~n28360 ;
  assign n28362 = ~n15414 & n28361 ;
  assign n28363 = n28332 | n28362 ;
  assign n28364 = n15421 | n28363 ;
  assign n28365 = n15421 & ~n28331 ;
  assign n28366 = n28364 & ~n28365 ;
  assign n28367 = x792 | n28366 ;
  assign n28368 = x628 & ~n28366 ;
  assign n28369 = x628 | n28331 ;
  assign n28370 = ~n28368 & n28369 ;
  assign n28371 = ( ~x792 & x1156 ) | ( ~x792 & n28370 ) | ( x1156 & n28370 ) ;
  assign n28372 = x628 | n28366 ;
  assign n28373 = x628 & ~n28331 ;
  assign n28374 = n28372 & ~n28373 ;
  assign n28375 = ( x792 & x1156 ) | ( x792 & ~n28374 ) | ( x1156 & ~n28374 ) ;
  assign n28376 = ~n28371 & n28375 ;
  assign n28377 = n28367 & ~n28376 ;
  assign n28378 = x787 | n28377 ;
  assign n28379 = x647 & ~n28377 ;
  assign n28380 = x647 | n28331 ;
  assign n28381 = ~n28379 & n28380 ;
  assign n28382 = ( ~x787 & x1157 ) | ( ~x787 & n28381 ) | ( x1157 & n28381 ) ;
  assign n28383 = x647 | n28377 ;
  assign n28384 = x647 & ~n28331 ;
  assign n28385 = n28383 & ~n28384 ;
  assign n28386 = ( x787 & x1157 ) | ( x787 & ~n28385 ) | ( x1157 & ~n28385 ) ;
  assign n28387 = ~n28382 & n28386 ;
  assign n28388 = n28378 & ~n28387 ;
  assign n28389 = x644 | n28388 ;
  assign n28390 = x715 & n28389 ;
  assign n28391 = ~x763 & n14710 ;
  assign n28392 = x190 & ~n14907 ;
  assign n28393 = n28391 | n28392 ;
  assign n28394 = x39 & n28393 ;
  assign n28395 = ~x190 & x763 ;
  assign n28396 = n15063 & n28395 ;
  assign n28397 = x763 & n14932 ;
  assign n28398 = x190 & ~n28397 ;
  assign n28399 = n20280 | n28398 ;
  assign n28400 = n28396 | n28399 ;
  assign n28401 = n28394 | n28400 ;
  assign n28402 = ~x38 & n28401 ;
  assign n28403 = x763 & n15072 ;
  assign n28404 = x38 & n28334 ;
  assign n28405 = ~n28403 & n28404 ;
  assign n28406 = n28402 | n28405 ;
  assign n28407 = ~n2032 & n28406 ;
  assign n28408 = n28333 | n28407 ;
  assign n28409 = ~n15082 & n28408 ;
  assign n28410 = n15082 & n28331 ;
  assign n28411 = n28409 | n28410 ;
  assign n28412 = ~x785 & n28411 ;
  assign n28413 = ~n15088 & n28331 ;
  assign n28414 = x609 & n28409 ;
  assign n28415 = n28413 | n28414 ;
  assign n28416 = x1155 & n28415 ;
  assign n28417 = n15094 & n28331 ;
  assign n28418 = ~x609 & n28409 ;
  assign n28419 = n28417 | n28418 ;
  assign n28420 = ~x1155 & n28419 ;
  assign n28421 = n28416 | n28420 ;
  assign n28422 = x785 & n28421 ;
  assign n28423 = n28412 | n28422 ;
  assign n28424 = ~x781 & n28423 ;
  assign n28425 = ( x618 & x1154 ) | ( x618 & n28331 ) | ( x1154 & n28331 ) ;
  assign n28426 = ( ~x618 & x1154 ) | ( ~x618 & n28423 ) | ( x1154 & n28423 ) ;
  assign n28427 = n28425 & n28426 ;
  assign n28428 = ( x618 & x1154 ) | ( x618 & ~n28331 ) | ( x1154 & ~n28331 ) ;
  assign n28429 = ( x618 & ~x1154 ) | ( x618 & n28423 ) | ( ~x1154 & n28423 ) ;
  assign n28430 = ~n28428 & n28429 ;
  assign n28431 = n28427 | n28430 ;
  assign n28432 = x781 & n28431 ;
  assign n28433 = n28424 | n28432 ;
  assign n28434 = ~x789 & n28433 ;
  assign n28435 = ( x619 & x1159 ) | ( x619 & n28331 ) | ( x1159 & n28331 ) ;
  assign n28436 = ( ~x619 & x1159 ) | ( ~x619 & n28433 ) | ( x1159 & n28433 ) ;
  assign n28437 = n28435 & n28436 ;
  assign n28438 = ( x619 & x1159 ) | ( x619 & ~n28331 ) | ( x1159 & ~n28331 ) ;
  assign n28439 = ( x619 & ~x1159 ) | ( x619 & n28433 ) | ( ~x1159 & n28433 ) ;
  assign n28440 = ~n28438 & n28439 ;
  assign n28441 = n28437 | n28440 ;
  assign n28442 = x789 & n28441 ;
  assign n28443 = n28434 | n28442 ;
  assign n28444 = n16176 | n28443 ;
  assign n28445 = n16176 & ~n28331 ;
  assign n28446 = n28444 & ~n28445 ;
  assign n28447 = n15134 | n28446 ;
  assign n28448 = n15134 & ~n28331 ;
  assign n28449 = n28447 & ~n28448 ;
  assign n28450 = n15141 | n28449 ;
  assign n28451 = n15141 & ~n28331 ;
  assign n28452 = n28450 & ~n28451 ;
  assign n28453 = ( x644 & x715 ) | ( x644 & ~n28452 ) | ( x715 & ~n28452 ) ;
  assign n28454 = ( x644 & ~x715 ) | ( x644 & n28331 ) | ( ~x715 & n28331 ) ;
  assign n28455 = ~n28453 & n28454 ;
  assign n28456 = x1160 & ~n28455 ;
  assign n28457 = ~n28390 & n28456 ;
  assign n28458 = x644 & ~n28388 ;
  assign n28459 = x715 | n28458 ;
  assign n28460 = ( x644 & x715 ) | ( x644 & n28452 ) | ( x715 & n28452 ) ;
  assign n28461 = ( ~x644 & x715 ) | ( ~x644 & n28331 ) | ( x715 & n28331 ) ;
  assign n28462 = n28460 & n28461 ;
  assign n28463 = x1160 | n28462 ;
  assign n28464 = n28459 & ~n28463 ;
  assign n28465 = n28457 | n28464 ;
  assign n28466 = x790 & n28465 ;
  assign n28467 = n18621 & n28446 ;
  assign n28468 = n15132 & n28374 ;
  assign n28469 = n15131 & n28370 ;
  assign n28470 = n28468 | n28469 ;
  assign n28471 = n28467 | n28470 ;
  assign n28472 = x792 & n28471 ;
  assign n28473 = x648 & ~n28440 ;
  assign n28474 = ( x619 & x1159 ) | ( x619 & n28361 ) | ( x1159 & n28361 ) ;
  assign n28475 = x627 | n28427 ;
  assign n28476 = ( x618 & x1154 ) | ( x618 & ~n28358 ) | ( x1154 & ~n28358 ) ;
  assign n28477 = x660 | n28416 ;
  assign n28478 = ( x609 & x1155 ) | ( x609 & ~n28355 ) | ( x1155 & ~n28355 ) ;
  assign n28479 = x608 | n28349 ;
  assign n28480 = ( x625 & x1153 ) | ( x625 & ~n28408 ) | ( x1153 & ~n28408 ) ;
  assign n28481 = x699 | n28406 ;
  assign n28482 = ( x190 & ~x763 ) | ( x190 & n15872 ) | ( ~x763 & n15872 ) ;
  assign n28483 = ( x190 & x763 ) | ( x190 & n15797 ) | ( x763 & n15797 ) ;
  assign n28484 = ~n28482 & n28483 ;
  assign n28485 = x39 & ~n28484 ;
  assign n28486 = ( x190 & ~x763 ) | ( x190 & n15699 ) | ( ~x763 & n15699 ) ;
  assign n28487 = ( x190 & x763 ) | ( x190 & n15583 ) | ( x763 & n15583 ) ;
  assign n28488 = n28486 & ~n28487 ;
  assign n28489 = n28485 & ~n28488 ;
  assign n28490 = ( x190 & ~x763 ) | ( x190 & n15891 ) | ( ~x763 & n15891 ) ;
  assign n28491 = ( x190 & x763 ) | ( x190 & n15887 ) | ( x763 & n15887 ) ;
  assign n28492 = n28490 & ~n28491 ;
  assign n28493 = ( x190 & ~x763 ) | ( x190 & n15897 ) | ( ~x763 & n15897 ) ;
  assign n28494 = ( x190 & x763 ) | ( x190 & n15894 ) | ( x763 & n15894 ) ;
  assign n28495 = ~n28493 & n28494 ;
  assign n28496 = n28492 | n28495 ;
  assign n28497 = ( ~x38 & n9138 ) | ( ~x38 & n28496 ) | ( n9138 & n28496 ) ;
  assign n28498 = ~n28489 & n28497 ;
  assign n28499 = ~x763 & n22085 ;
  assign n28500 = n15758 | n28499 ;
  assign n28501 = ~x39 & n28500 ;
  assign n28502 = x190 | n28501 ;
  assign n28503 = n15529 | n28159 ;
  assign n28504 = x190 & n28503 ;
  assign n28505 = ~n4810 & n28504 ;
  assign n28506 = x38 & ~n28505 ;
  assign n28507 = n28502 & n28506 ;
  assign n28508 = x699 & ~n28507 ;
  assign n28509 = ~n28498 & n28508 ;
  assign n28510 = n2032 | n28509 ;
  assign n28511 = n28481 & ~n28510 ;
  assign n28512 = n28333 | n28511 ;
  assign n28513 = ( x625 & ~x1153 ) | ( x625 & n28512 ) | ( ~x1153 & n28512 ) ;
  assign n28514 = ~n28480 & n28513 ;
  assign n28515 = n28479 | n28514 ;
  assign n28516 = x608 & ~n28352 ;
  assign n28517 = ( x625 & x1153 ) | ( x625 & n28408 ) | ( x1153 & n28408 ) ;
  assign n28518 = ( ~x625 & x1153 ) | ( ~x625 & n28512 ) | ( x1153 & n28512 ) ;
  assign n28519 = n28517 & n28518 ;
  assign n28520 = n28516 & ~n28519 ;
  assign n28521 = n28515 & ~n28520 ;
  assign n28522 = x778 & ~n28521 ;
  assign n28523 = x778 | n28512 ;
  assign n28524 = ~n28522 & n28523 ;
  assign n28525 = ( x609 & ~x1155 ) | ( x609 & n28524 ) | ( ~x1155 & n28524 ) ;
  assign n28526 = ~n28478 & n28525 ;
  assign n28527 = n28477 | n28526 ;
  assign n28528 = x660 & ~n28420 ;
  assign n28529 = ( x609 & x1155 ) | ( x609 & n28355 ) | ( x1155 & n28355 ) ;
  assign n28530 = ( ~x609 & x1155 ) | ( ~x609 & n28524 ) | ( x1155 & n28524 ) ;
  assign n28531 = n28529 & n28530 ;
  assign n28532 = n28528 & ~n28531 ;
  assign n28533 = n28527 & ~n28532 ;
  assign n28534 = x785 & ~n28533 ;
  assign n28535 = x785 | n28524 ;
  assign n28536 = ~n28534 & n28535 ;
  assign n28537 = ( x618 & ~x1154 ) | ( x618 & n28536 ) | ( ~x1154 & n28536 ) ;
  assign n28538 = ~n28476 & n28537 ;
  assign n28539 = n28475 | n28538 ;
  assign n28540 = x627 & ~n28430 ;
  assign n28541 = ( x618 & x1154 ) | ( x618 & n28358 ) | ( x1154 & n28358 ) ;
  assign n28542 = ( ~x618 & x1154 ) | ( ~x618 & n28536 ) | ( x1154 & n28536 ) ;
  assign n28543 = n28541 & n28542 ;
  assign n28544 = n28540 & ~n28543 ;
  assign n28545 = n28539 & ~n28544 ;
  assign n28546 = x781 & ~n28545 ;
  assign n28547 = x781 | n28536 ;
  assign n28548 = ~n28546 & n28547 ;
  assign n28549 = ( ~x619 & x1159 ) | ( ~x619 & n28548 ) | ( x1159 & n28548 ) ;
  assign n28550 = n28474 & n28549 ;
  assign n28551 = n28473 & ~n28550 ;
  assign n28552 = x648 | n28437 ;
  assign n28553 = ( x619 & x1159 ) | ( x619 & ~n28361 ) | ( x1159 & ~n28361 ) ;
  assign n28554 = ( x619 & ~x1159 ) | ( x619 & n28548 ) | ( ~x1159 & n28548 ) ;
  assign n28555 = ~n28553 & n28554 ;
  assign n28556 = n28552 | n28555 ;
  assign n28557 = x789 & n28556 ;
  assign n28558 = ~n28551 & n28557 ;
  assign n28559 = ~x789 & n28548 ;
  assign n28560 = n16177 | n28559 ;
  assign n28561 = n28558 | n28560 ;
  assign n28562 = n16115 & ~n28363 ;
  assign n28563 = ( x626 & ~n15419 ) | ( x626 & n28331 ) | ( ~n15419 & n28331 ) ;
  assign n28564 = ( x626 & n15419 ) | ( x626 & ~n28443 ) | ( n15419 & ~n28443 ) ;
  assign n28565 = ~n28563 & n28564 ;
  assign n28566 = n28562 | n28565 ;
  assign n28567 = ( x626 & n15418 ) | ( x626 & ~n28331 ) | ( n15418 & ~n28331 ) ;
  assign n28568 = ( x626 & ~n15418 ) | ( x626 & n28443 ) | ( ~n15418 & n28443 ) ;
  assign n28569 = n28567 & ~n28568 ;
  assign n28570 = n28566 | n28569 ;
  assign n28571 = x788 & n28570 ;
  assign n28572 = n18434 | n28571 ;
  assign n28573 = n28561 & ~n28572 ;
  assign n28574 = n28472 | n28573 ;
  assign n28575 = ~n18431 & n28574 ;
  assign n28576 = n15138 & n28381 ;
  assign n28577 = n15139 & n28385 ;
  assign n28578 = n18610 & n28449 ;
  assign n28579 = n28577 | n28578 ;
  assign n28580 = n28576 | n28579 ;
  assign n28581 = x787 & n28580 ;
  assign n28582 = n28575 | n28581 ;
  assign n28583 = ( x644 & ~x790 ) | ( x644 & n28456 ) | ( ~x790 & n28456 ) ;
  assign n28584 = ( x644 & x790 ) | ( x644 & n28463 ) | ( x790 & n28463 ) ;
  assign n28585 = ~n28583 & n28584 ;
  assign n28586 = n28582 | n28585 ;
  assign n28587 = ~n28466 & n28586 ;
  assign n28588 = ( ~x832 & n6785 ) | ( ~x832 & n28587 ) | ( n6785 & n28587 ) ;
  assign n28589 = ( ~x190 & x832 ) | ( ~x190 & n6785 ) | ( x832 & n6785 ) ;
  assign n28590 = n28588 & ~n28589 ;
  assign n28591 = n28330 | n28590 ;
  assign n28592 = x191 | n1290 ;
  assign n28593 = x746 & n14840 ;
  assign n28594 = n28592 & ~n28593 ;
  assign n28595 = n16060 | n28594 ;
  assign n28596 = ~x785 & n28595 ;
  assign n28597 = ~n15094 & n28593 ;
  assign n28598 = n28595 | n28597 ;
  assign n28599 = x1155 & n28598 ;
  assign n28600 = ~x1155 & n28592 ;
  assign n28601 = ~n28597 & n28600 ;
  assign n28602 = n28599 | n28601 ;
  assign n28603 = x785 & n28602 ;
  assign n28604 = n28596 | n28603 ;
  assign n28605 = ~x781 & n28604 ;
  assign n28606 = n16075 | n28604 ;
  assign n28607 = x1154 & n28606 ;
  assign n28608 = n16078 | n28604 ;
  assign n28609 = ~x1154 & n28608 ;
  assign n28610 = n28607 | n28609 ;
  assign n28611 = x781 & n28610 ;
  assign n28612 = n28605 | n28611 ;
  assign n28613 = ~x789 & n28612 ;
  assign n28614 = n20948 | n28612 ;
  assign n28615 = x1159 & n28614 ;
  assign n28616 = n20951 | n28612 ;
  assign n28617 = ~x1159 & n28616 ;
  assign n28618 = n28615 | n28617 ;
  assign n28619 = x789 & n28618 ;
  assign n28620 = n28613 | n28619 ;
  assign n28621 = n16176 | n28620 ;
  assign n28622 = n16176 & ~n28592 ;
  assign n28623 = n28621 & ~n28622 ;
  assign n28624 = n15134 | n28623 ;
  assign n28625 = n15134 & ~n28592 ;
  assign n28626 = n28624 & ~n28625 ;
  assign n28627 = n18610 & n28626 ;
  assign n28628 = ( x647 & x1157 ) | ( x647 & ~n28592 ) | ( x1157 & ~n28592 ) ;
  assign n28629 = x729 & n15202 ;
  assign n28630 = n28592 & ~n28629 ;
  assign n28631 = x778 | n28630 ;
  assign n28632 = ~x625 & n28629 ;
  assign n28633 = n28630 | n28632 ;
  assign n28634 = x1153 & n28633 ;
  assign n28635 = ~x1153 & n28592 ;
  assign n28636 = ~n28632 & n28635 ;
  assign n28637 = x778 & ~n28636 ;
  assign n28638 = ~n28634 & n28637 ;
  assign n28639 = n28631 & ~n28638 ;
  assign n28640 = n16043 | n28639 ;
  assign n28641 = n16045 | n28640 ;
  assign n28642 = n16047 | n28641 ;
  assign n28643 = n16049 | n28642 ;
  assign n28644 = n16055 | n28643 ;
  assign n28645 = ( x647 & ~x1157 ) | ( x647 & n28644 ) | ( ~x1157 & n28644 ) ;
  assign n28646 = ~n28628 & n28645 ;
  assign n28647 = x630 & n28646 ;
  assign n28648 = x647 & n28644 ;
  assign n28649 = ~x647 & n28592 ;
  assign n28650 = n28648 | n28649 ;
  assign n28651 = n15138 & n28650 ;
  assign n28652 = n28647 | n28651 ;
  assign n28653 = n28627 | n28652 ;
  assign n28654 = x787 & n28653 ;
  assign n28655 = n16115 & ~n28642 ;
  assign n28656 = ( x626 & ~n15419 ) | ( x626 & n28592 ) | ( ~n15419 & n28592 ) ;
  assign n28657 = ( x626 & n15419 ) | ( x626 & ~n28620 ) | ( n15419 & ~n28620 ) ;
  assign n28658 = ~n28656 & n28657 ;
  assign n28659 = n28655 | n28658 ;
  assign n28660 = ( x626 & n15418 ) | ( x626 & ~n28592 ) | ( n15418 & ~n28592 ) ;
  assign n28661 = ( x626 & ~n15418 ) | ( x626 & n28620 ) | ( ~n15418 & n28620 ) ;
  assign n28662 = n28660 & ~n28661 ;
  assign n28663 = n28659 | n28662 ;
  assign n28664 = x788 & n28663 ;
  assign n28665 = x648 & ~n28617 ;
  assign n28666 = ( x619 & x1159 ) | ( x619 & n28641 ) | ( x1159 & n28641 ) ;
  assign n28667 = x627 | n28607 ;
  assign n28668 = ( x618 & x1154 ) | ( x618 & ~n28640 ) | ( x1154 & ~n28640 ) ;
  assign n28669 = x660 | n28599 ;
  assign n28670 = ( x609 & x1155 ) | ( x609 & ~n28639 ) | ( x1155 & ~n28639 ) ;
  assign n28671 = n14839 | n28630 ;
  assign n28672 = x625 & ~n28671 ;
  assign n28673 = n28594 & n28671 ;
  assign n28674 = n28672 | n28673 ;
  assign n28675 = n28635 & n28674 ;
  assign n28676 = x608 | n28634 ;
  assign n28677 = n28675 | n28676 ;
  assign n28678 = x1153 & n28594 ;
  assign n28679 = ~n28672 & n28678 ;
  assign n28680 = x608 & ~n28636 ;
  assign n28681 = ~n28679 & n28680 ;
  assign n28682 = n28677 & ~n28681 ;
  assign n28683 = x778 & ~n28682 ;
  assign n28684 = x778 | n28673 ;
  assign n28685 = ~n28683 & n28684 ;
  assign n28686 = ( x609 & ~x1155 ) | ( x609 & n28685 ) | ( ~x1155 & n28685 ) ;
  assign n28687 = ~n28670 & n28686 ;
  assign n28688 = n28669 | n28687 ;
  assign n28689 = x660 & ~n28601 ;
  assign n28690 = ( x609 & x1155 ) | ( x609 & n28639 ) | ( x1155 & n28639 ) ;
  assign n28691 = ( ~x609 & x1155 ) | ( ~x609 & n28685 ) | ( x1155 & n28685 ) ;
  assign n28692 = n28690 & n28691 ;
  assign n28693 = n28689 & ~n28692 ;
  assign n28694 = n28688 & ~n28693 ;
  assign n28695 = x785 & ~n28694 ;
  assign n28696 = x785 | n28685 ;
  assign n28697 = ~n28695 & n28696 ;
  assign n28698 = ( x618 & ~x1154 ) | ( x618 & n28697 ) | ( ~x1154 & n28697 ) ;
  assign n28699 = ~n28668 & n28698 ;
  assign n28700 = n28667 | n28699 ;
  assign n28701 = x627 & ~n28609 ;
  assign n28702 = ( x618 & x1154 ) | ( x618 & n28640 ) | ( x1154 & n28640 ) ;
  assign n28703 = ( ~x618 & x1154 ) | ( ~x618 & n28697 ) | ( x1154 & n28697 ) ;
  assign n28704 = n28702 & n28703 ;
  assign n28705 = n28701 & ~n28704 ;
  assign n28706 = n28700 & ~n28705 ;
  assign n28707 = x781 & ~n28706 ;
  assign n28708 = x781 | n28697 ;
  assign n28709 = ~n28707 & n28708 ;
  assign n28710 = ( ~x619 & x1159 ) | ( ~x619 & n28709 ) | ( x1159 & n28709 ) ;
  assign n28711 = n28666 & n28710 ;
  assign n28712 = n28665 & ~n28711 ;
  assign n28713 = x648 | n28615 ;
  assign n28714 = ( x619 & x1159 ) | ( x619 & ~n28641 ) | ( x1159 & ~n28641 ) ;
  assign n28715 = ( x619 & ~x1159 ) | ( x619 & n28709 ) | ( ~x1159 & n28709 ) ;
  assign n28716 = ~n28714 & n28715 ;
  assign n28717 = n28713 | n28716 ;
  assign n28718 = x789 & n28717 ;
  assign n28719 = ~n28712 & n28718 ;
  assign n28720 = ~x789 & n28709 ;
  assign n28721 = n16177 | n28720 ;
  assign n28722 = n28719 | n28721 ;
  assign n28723 = ~n28664 & n28722 ;
  assign n28724 = n18434 | n28723 ;
  assign n28725 = n16650 | n28643 ;
  assign n28726 = n16051 & ~n28623 ;
  assign n28727 = n28725 & ~n28726 ;
  assign n28728 = ( x629 & ~x792 ) | ( x629 & n28727 ) | ( ~x792 & n28727 ) ;
  assign n28729 = n16052 & ~n28623 ;
  assign n28730 = n16643 & ~n28643 ;
  assign n28731 = n28729 | n28730 ;
  assign n28732 = ( x629 & x792 ) | ( x629 & n28731 ) | ( x792 & n28731 ) ;
  assign n28733 = ~n28728 & n28732 ;
  assign n28734 = n18431 | n28733 ;
  assign n28735 = n28724 & ~n28734 ;
  assign n28736 = n28654 | n28735 ;
  assign n28737 = ( x790 & x832 ) | ( x790 & n28736 ) | ( x832 & n28736 ) ;
  assign n28738 = n15141 | n28626 ;
  assign n28739 = n15141 & ~n28592 ;
  assign n28740 = n28738 & ~n28739 ;
  assign n28741 = ( x644 & x715 ) | ( x644 & ~n28740 ) | ( x715 & ~n28740 ) ;
  assign n28742 = ( x644 & ~x715 ) | ( x644 & n28592 ) | ( ~x715 & n28592 ) ;
  assign n28743 = ~n28741 & n28742 ;
  assign n28744 = x1160 & ~n28743 ;
  assign n28745 = ~x787 & n28644 ;
  assign n28746 = x1157 & n28650 ;
  assign n28747 = n28646 | n28746 ;
  assign n28748 = x787 & n28747 ;
  assign n28749 = n28745 | n28748 ;
  assign n28750 = ( x644 & x715 ) | ( x644 & n28749 ) | ( x715 & n28749 ) ;
  assign n28751 = ( ~x644 & x715 ) | ( ~x644 & n28736 ) | ( x715 & n28736 ) ;
  assign n28752 = n28750 & n28751 ;
  assign n28753 = n28744 & ~n28752 ;
  assign n28754 = ( x644 & x715 ) | ( x644 & n28740 ) | ( x715 & n28740 ) ;
  assign n28755 = ( ~x644 & x715 ) | ( ~x644 & n28592 ) | ( x715 & n28592 ) ;
  assign n28756 = n28754 & n28755 ;
  assign n28757 = x1160 | n28756 ;
  assign n28758 = ( x644 & x715 ) | ( x644 & ~n28749 ) | ( x715 & ~n28749 ) ;
  assign n28759 = ( x644 & ~x715 ) | ( x644 & n28736 ) | ( ~x715 & n28736 ) ;
  assign n28760 = ~n28758 & n28759 ;
  assign n28761 = n28757 | n28760 ;
  assign n28762 = ~n28753 & n28761 ;
  assign n28763 = ( ~x790 & x832 ) | ( ~x790 & n28762 ) | ( x832 & n28762 ) ;
  assign n28764 = n28737 & n28763 ;
  assign n28765 = x191 | n14834 ;
  assign n28766 = n15414 & n28765 ;
  assign n28767 = x191 & n2032 ;
  assign n28768 = x191 | n15070 ;
  assign n28769 = n15375 & n28768 ;
  assign n28770 = x729 & ~n28769 ;
  assign n28771 = ( ~x38 & x191 ) | ( ~x38 & n16319 ) | ( x191 & n16319 ) ;
  assign n28772 = ( x38 & x191 ) | ( x38 & n16323 ) | ( x191 & n16323 ) ;
  assign n28773 = n28771 & ~n28772 ;
  assign n28774 = n28770 & ~n28773 ;
  assign n28775 = x191 | x729 ;
  assign n28776 = n15382 | n28775 ;
  assign n28777 = ~n2032 & n28776 ;
  assign n28778 = ~n28774 & n28777 ;
  assign n28779 = n28767 | n28778 ;
  assign n28780 = ~x778 & n28779 ;
  assign n28781 = ( x625 & x1153 ) | ( x625 & n28765 ) | ( x1153 & n28765 ) ;
  assign n28782 = ( ~x625 & x1153 ) | ( ~x625 & n28779 ) | ( x1153 & n28779 ) ;
  assign n28783 = n28781 & n28782 ;
  assign n28784 = ( x625 & x1153 ) | ( x625 & ~n28765 ) | ( x1153 & ~n28765 ) ;
  assign n28785 = ( x625 & ~x1153 ) | ( x625 & n28779 ) | ( ~x1153 & n28779 ) ;
  assign n28786 = ~n28784 & n28785 ;
  assign n28787 = n28783 | n28786 ;
  assign n28788 = x778 & n28787 ;
  assign n28789 = n28780 | n28788 ;
  assign n28790 = ~n15400 & n28789 ;
  assign n28791 = n15400 & n28765 ;
  assign n28792 = n28790 | n28791 ;
  assign n28793 = n15407 | n28792 ;
  assign n28794 = n15407 & ~n28765 ;
  assign n28795 = n28793 & ~n28794 ;
  assign n28796 = ~n15414 & n28795 ;
  assign n28797 = n28766 | n28796 ;
  assign n28798 = n15421 | n28797 ;
  assign n28799 = n15421 & ~n28765 ;
  assign n28800 = n28798 & ~n28799 ;
  assign n28801 = x792 | n28800 ;
  assign n28802 = x628 & ~n28800 ;
  assign n28803 = x628 | n28765 ;
  assign n28804 = ~n28802 & n28803 ;
  assign n28805 = ( ~x792 & x1156 ) | ( ~x792 & n28804 ) | ( x1156 & n28804 ) ;
  assign n28806 = x628 | n28800 ;
  assign n28807 = x628 & ~n28765 ;
  assign n28808 = n28806 & ~n28807 ;
  assign n28809 = ( x792 & x1156 ) | ( x792 & ~n28808 ) | ( x1156 & ~n28808 ) ;
  assign n28810 = ~n28805 & n28809 ;
  assign n28811 = n28801 & ~n28810 ;
  assign n28812 = x787 | n28811 ;
  assign n28813 = x647 & ~n28811 ;
  assign n28814 = x647 | n28765 ;
  assign n28815 = ~n28813 & n28814 ;
  assign n28816 = ( ~x787 & x1157 ) | ( ~x787 & n28815 ) | ( x1157 & n28815 ) ;
  assign n28817 = x647 | n28811 ;
  assign n28818 = x647 & ~n28765 ;
  assign n28819 = n28817 & ~n28818 ;
  assign n28820 = ( x787 & x1157 ) | ( x787 & ~n28819 ) | ( x1157 & ~n28819 ) ;
  assign n28821 = ~n28816 & n28820 ;
  assign n28822 = n28812 & ~n28821 ;
  assign n28823 = x644 | n28822 ;
  assign n28824 = x715 & n28823 ;
  assign n28825 = ~x746 & n14710 ;
  assign n28826 = x191 & ~n14907 ;
  assign n28827 = n28825 | n28826 ;
  assign n28828 = x39 & n28827 ;
  assign n28829 = ~x191 & x746 ;
  assign n28830 = n15063 & n28829 ;
  assign n28831 = x746 & n14932 ;
  assign n28832 = x191 & ~n28831 ;
  assign n28833 = n20361 | n28832 ;
  assign n28834 = n28830 | n28833 ;
  assign n28835 = n28828 | n28834 ;
  assign n28836 = ~x38 & n28835 ;
  assign n28837 = x746 & n15072 ;
  assign n28838 = x38 & n28768 ;
  assign n28839 = ~n28837 & n28838 ;
  assign n28840 = n28836 | n28839 ;
  assign n28841 = ~n2032 & n28840 ;
  assign n28842 = n28767 | n28841 ;
  assign n28843 = ~n15082 & n28842 ;
  assign n28844 = n15082 & n28765 ;
  assign n28845 = n28843 | n28844 ;
  assign n28846 = ~x785 & n28845 ;
  assign n28847 = ~n15088 & n28765 ;
  assign n28848 = x609 & n28843 ;
  assign n28849 = n28847 | n28848 ;
  assign n28850 = x1155 & n28849 ;
  assign n28851 = n15094 & n28765 ;
  assign n28852 = ~x609 & n28843 ;
  assign n28853 = n28851 | n28852 ;
  assign n28854 = ~x1155 & n28853 ;
  assign n28855 = n28850 | n28854 ;
  assign n28856 = x785 & n28855 ;
  assign n28857 = n28846 | n28856 ;
  assign n28858 = ~x781 & n28857 ;
  assign n28859 = ( x618 & x1154 ) | ( x618 & n28765 ) | ( x1154 & n28765 ) ;
  assign n28860 = ( ~x618 & x1154 ) | ( ~x618 & n28857 ) | ( x1154 & n28857 ) ;
  assign n28861 = n28859 & n28860 ;
  assign n28862 = ( x618 & x1154 ) | ( x618 & ~n28765 ) | ( x1154 & ~n28765 ) ;
  assign n28863 = ( x618 & ~x1154 ) | ( x618 & n28857 ) | ( ~x1154 & n28857 ) ;
  assign n28864 = ~n28862 & n28863 ;
  assign n28865 = n28861 | n28864 ;
  assign n28866 = x781 & n28865 ;
  assign n28867 = n28858 | n28866 ;
  assign n28868 = ~x789 & n28867 ;
  assign n28869 = ( x619 & x1159 ) | ( x619 & n28765 ) | ( x1159 & n28765 ) ;
  assign n28870 = ( ~x619 & x1159 ) | ( ~x619 & n28867 ) | ( x1159 & n28867 ) ;
  assign n28871 = n28869 & n28870 ;
  assign n28872 = ( x619 & x1159 ) | ( x619 & ~n28765 ) | ( x1159 & ~n28765 ) ;
  assign n28873 = ( x619 & ~x1159 ) | ( x619 & n28867 ) | ( ~x1159 & n28867 ) ;
  assign n28874 = ~n28872 & n28873 ;
  assign n28875 = n28871 | n28874 ;
  assign n28876 = x789 & n28875 ;
  assign n28877 = n28868 | n28876 ;
  assign n28878 = n16176 | n28877 ;
  assign n28879 = n16176 & ~n28765 ;
  assign n28880 = n28878 & ~n28879 ;
  assign n28881 = n15134 | n28880 ;
  assign n28882 = n15134 & ~n28765 ;
  assign n28883 = n28881 & ~n28882 ;
  assign n28884 = n15141 | n28883 ;
  assign n28885 = n15141 & ~n28765 ;
  assign n28886 = n28884 & ~n28885 ;
  assign n28887 = ( x644 & x715 ) | ( x644 & ~n28886 ) | ( x715 & ~n28886 ) ;
  assign n28888 = ( x644 & ~x715 ) | ( x644 & n28765 ) | ( ~x715 & n28765 ) ;
  assign n28889 = ~n28887 & n28888 ;
  assign n28890 = x1160 & ~n28889 ;
  assign n28891 = ~n28824 & n28890 ;
  assign n28892 = x644 & ~n28822 ;
  assign n28893 = x715 | n28892 ;
  assign n28894 = ( x644 & x715 ) | ( x644 & n28886 ) | ( x715 & n28886 ) ;
  assign n28895 = ( ~x644 & x715 ) | ( ~x644 & n28765 ) | ( x715 & n28765 ) ;
  assign n28896 = n28894 & n28895 ;
  assign n28897 = x1160 | n28896 ;
  assign n28898 = n28893 & ~n28897 ;
  assign n28899 = n28891 | n28898 ;
  assign n28900 = x790 & n28899 ;
  assign n28901 = n18621 & n28880 ;
  assign n28902 = n15132 & n28808 ;
  assign n28903 = n15131 & n28804 ;
  assign n28904 = n28902 | n28903 ;
  assign n28905 = n28901 | n28904 ;
  assign n28906 = x792 & n28905 ;
  assign n28907 = x648 & ~n28874 ;
  assign n28908 = ( x619 & x1159 ) | ( x619 & n28795 ) | ( x1159 & n28795 ) ;
  assign n28909 = x627 | n28861 ;
  assign n28910 = ( x618 & x1154 ) | ( x618 & ~n28792 ) | ( x1154 & ~n28792 ) ;
  assign n28911 = x660 | n28850 ;
  assign n28912 = ( x609 & x1155 ) | ( x609 & ~n28789 ) | ( x1155 & ~n28789 ) ;
  assign n28913 = x608 | n28783 ;
  assign n28914 = ( x625 & x1153 ) | ( x625 & ~n28842 ) | ( x1153 & ~n28842 ) ;
  assign n28915 = x729 | n28840 ;
  assign n28916 = ( x191 & ~x746 ) | ( x191 & n15872 ) | ( ~x746 & n15872 ) ;
  assign n28917 = ( x191 & x746 ) | ( x191 & n15797 ) | ( x746 & n15797 ) ;
  assign n28918 = ~n28916 & n28917 ;
  assign n28919 = x39 & ~n28918 ;
  assign n28920 = ( x191 & ~x746 ) | ( x191 & n15699 ) | ( ~x746 & n15699 ) ;
  assign n28921 = ( x191 & x746 ) | ( x191 & n15583 ) | ( x746 & n15583 ) ;
  assign n28922 = n28920 & ~n28921 ;
  assign n28923 = n28919 & ~n28922 ;
  assign n28924 = ( x191 & ~x746 ) | ( x191 & n15891 ) | ( ~x746 & n15891 ) ;
  assign n28925 = ( x191 & x746 ) | ( x191 & n15887 ) | ( x746 & n15887 ) ;
  assign n28926 = n28924 & ~n28925 ;
  assign n28927 = ( x191 & ~x746 ) | ( x191 & n15897 ) | ( ~x746 & n15897 ) ;
  assign n28928 = ( x191 & x746 ) | ( x191 & n15894 ) | ( x746 & n15894 ) ;
  assign n28929 = ~n28927 & n28928 ;
  assign n28930 = n28926 | n28929 ;
  assign n28931 = ( ~x38 & n9138 ) | ( ~x38 & n28930 ) | ( n9138 & n28930 ) ;
  assign n28932 = ~n28923 & n28931 ;
  assign n28933 = ~x746 & n22085 ;
  assign n28934 = n15758 | n28933 ;
  assign n28935 = ~x39 & n28934 ;
  assign n28936 = x191 | n28935 ;
  assign n28937 = n15529 | n28593 ;
  assign n28938 = x191 & n28937 ;
  assign n28939 = ~n4810 & n28938 ;
  assign n28940 = x38 & ~n28939 ;
  assign n28941 = n28936 & n28940 ;
  assign n28942 = x729 & ~n28941 ;
  assign n28943 = ~n28932 & n28942 ;
  assign n28944 = n2032 | n28943 ;
  assign n28945 = n28915 & ~n28944 ;
  assign n28946 = n28767 | n28945 ;
  assign n28947 = ( x625 & ~x1153 ) | ( x625 & n28946 ) | ( ~x1153 & n28946 ) ;
  assign n28948 = ~n28914 & n28947 ;
  assign n28949 = n28913 | n28948 ;
  assign n28950 = x608 & ~n28786 ;
  assign n28951 = ( x625 & x1153 ) | ( x625 & n28842 ) | ( x1153 & n28842 ) ;
  assign n28952 = ( ~x625 & x1153 ) | ( ~x625 & n28946 ) | ( x1153 & n28946 ) ;
  assign n28953 = n28951 & n28952 ;
  assign n28954 = n28950 & ~n28953 ;
  assign n28955 = n28949 & ~n28954 ;
  assign n28956 = x778 & ~n28955 ;
  assign n28957 = x778 | n28946 ;
  assign n28958 = ~n28956 & n28957 ;
  assign n28959 = ( x609 & ~x1155 ) | ( x609 & n28958 ) | ( ~x1155 & n28958 ) ;
  assign n28960 = ~n28912 & n28959 ;
  assign n28961 = n28911 | n28960 ;
  assign n28962 = x660 & ~n28854 ;
  assign n28963 = ( x609 & x1155 ) | ( x609 & n28789 ) | ( x1155 & n28789 ) ;
  assign n28964 = ( ~x609 & x1155 ) | ( ~x609 & n28958 ) | ( x1155 & n28958 ) ;
  assign n28965 = n28963 & n28964 ;
  assign n28966 = n28962 & ~n28965 ;
  assign n28967 = n28961 & ~n28966 ;
  assign n28968 = x785 & ~n28967 ;
  assign n28969 = x785 | n28958 ;
  assign n28970 = ~n28968 & n28969 ;
  assign n28971 = ( x618 & ~x1154 ) | ( x618 & n28970 ) | ( ~x1154 & n28970 ) ;
  assign n28972 = ~n28910 & n28971 ;
  assign n28973 = n28909 | n28972 ;
  assign n28974 = x627 & ~n28864 ;
  assign n28975 = ( x618 & x1154 ) | ( x618 & n28792 ) | ( x1154 & n28792 ) ;
  assign n28976 = ( ~x618 & x1154 ) | ( ~x618 & n28970 ) | ( x1154 & n28970 ) ;
  assign n28977 = n28975 & n28976 ;
  assign n28978 = n28974 & ~n28977 ;
  assign n28979 = n28973 & ~n28978 ;
  assign n28980 = x781 & ~n28979 ;
  assign n28981 = x781 | n28970 ;
  assign n28982 = ~n28980 & n28981 ;
  assign n28983 = ( ~x619 & x1159 ) | ( ~x619 & n28982 ) | ( x1159 & n28982 ) ;
  assign n28984 = n28908 & n28983 ;
  assign n28985 = n28907 & ~n28984 ;
  assign n28986 = x648 | n28871 ;
  assign n28987 = ( x619 & x1159 ) | ( x619 & ~n28795 ) | ( x1159 & ~n28795 ) ;
  assign n28988 = ( x619 & ~x1159 ) | ( x619 & n28982 ) | ( ~x1159 & n28982 ) ;
  assign n28989 = ~n28987 & n28988 ;
  assign n28990 = n28986 | n28989 ;
  assign n28991 = x789 & n28990 ;
  assign n28992 = ~n28985 & n28991 ;
  assign n28993 = ~x789 & n28982 ;
  assign n28994 = n16177 | n28993 ;
  assign n28995 = n28992 | n28994 ;
  assign n28996 = n16115 & ~n28797 ;
  assign n28997 = ( x626 & ~n15419 ) | ( x626 & n28765 ) | ( ~n15419 & n28765 ) ;
  assign n28998 = ( x626 & n15419 ) | ( x626 & ~n28877 ) | ( n15419 & ~n28877 ) ;
  assign n28999 = ~n28997 & n28998 ;
  assign n29000 = n28996 | n28999 ;
  assign n29001 = ( x626 & n15418 ) | ( x626 & ~n28765 ) | ( n15418 & ~n28765 ) ;
  assign n29002 = ( x626 & ~n15418 ) | ( x626 & n28877 ) | ( ~n15418 & n28877 ) ;
  assign n29003 = n29001 & ~n29002 ;
  assign n29004 = n29000 | n29003 ;
  assign n29005 = x788 & n29004 ;
  assign n29006 = n18434 | n29005 ;
  assign n29007 = n28995 & ~n29006 ;
  assign n29008 = n28906 | n29007 ;
  assign n29009 = ~n18431 & n29008 ;
  assign n29010 = n15138 & n28815 ;
  assign n29011 = n15139 & n28819 ;
  assign n29012 = n18610 & n28883 ;
  assign n29013 = n29011 | n29012 ;
  assign n29014 = n29010 | n29013 ;
  assign n29015 = x787 & n29014 ;
  assign n29016 = n29009 | n29015 ;
  assign n29017 = ( x644 & ~x790 ) | ( x644 & n28890 ) | ( ~x790 & n28890 ) ;
  assign n29018 = ( x644 & x790 ) | ( x644 & n28897 ) | ( x790 & n28897 ) ;
  assign n29019 = ~n29017 & n29018 ;
  assign n29020 = n29016 | n29019 ;
  assign n29021 = ~n28900 & n29020 ;
  assign n29022 = ( ~x832 & n6785 ) | ( ~x832 & n29021 ) | ( n6785 & n29021 ) ;
  assign n29023 = ( ~x191 & x832 ) | ( ~x191 & n6785 ) | ( x832 & n6785 ) ;
  assign n29024 = n29022 & ~n29023 ;
  assign n29025 = n28764 | n29024 ;
  assign n29026 = x192 | n1290 ;
  assign n29027 = x764 & n14840 ;
  assign n29028 = n29026 & ~n29027 ;
  assign n29029 = n16060 | n29028 ;
  assign n29030 = ~x785 & n29029 ;
  assign n29031 = ~n15094 & n29027 ;
  assign n29032 = n29029 | n29031 ;
  assign n29033 = x1155 & n29032 ;
  assign n29034 = ~x1155 & n29026 ;
  assign n29035 = ~n29031 & n29034 ;
  assign n29036 = n29033 | n29035 ;
  assign n29037 = x785 & n29036 ;
  assign n29038 = n29030 | n29037 ;
  assign n29039 = ~x781 & n29038 ;
  assign n29040 = n16075 | n29038 ;
  assign n29041 = x1154 & n29040 ;
  assign n29042 = n16078 | n29038 ;
  assign n29043 = ~x1154 & n29042 ;
  assign n29044 = n29041 | n29043 ;
  assign n29045 = x781 & n29044 ;
  assign n29046 = n29039 | n29045 ;
  assign n29047 = ~x789 & n29046 ;
  assign n29048 = n20948 | n29046 ;
  assign n29049 = x1159 & n29048 ;
  assign n29050 = n20951 | n29046 ;
  assign n29051 = ~x1159 & n29050 ;
  assign n29052 = n29049 | n29051 ;
  assign n29053 = x789 & n29052 ;
  assign n29054 = n29047 | n29053 ;
  assign n29055 = n16176 | n29054 ;
  assign n29056 = n16176 & ~n29026 ;
  assign n29057 = n29055 & ~n29056 ;
  assign n29058 = n15134 | n29057 ;
  assign n29059 = n15134 & ~n29026 ;
  assign n29060 = n29058 & ~n29059 ;
  assign n29061 = n18610 & n29060 ;
  assign n29062 = ( x647 & x1157 ) | ( x647 & ~n29026 ) | ( x1157 & ~n29026 ) ;
  assign n29063 = x691 & n15202 ;
  assign n29064 = n29026 & ~n29063 ;
  assign n29065 = x778 | n29064 ;
  assign n29066 = ~x625 & n29063 ;
  assign n29067 = n29064 | n29066 ;
  assign n29068 = x1153 & n29067 ;
  assign n29069 = ~x1153 & n29026 ;
  assign n29070 = ~n29066 & n29069 ;
  assign n29071 = x778 & ~n29070 ;
  assign n29072 = ~n29068 & n29071 ;
  assign n29073 = n29065 & ~n29072 ;
  assign n29074 = n16043 | n29073 ;
  assign n29075 = n16045 | n29074 ;
  assign n29076 = n16047 | n29075 ;
  assign n29077 = n16049 | n29076 ;
  assign n29078 = n16055 | n29077 ;
  assign n29079 = ( x647 & ~x1157 ) | ( x647 & n29078 ) | ( ~x1157 & n29078 ) ;
  assign n29080 = ~n29062 & n29079 ;
  assign n29081 = x630 & n29080 ;
  assign n29082 = x647 & n29078 ;
  assign n29083 = ~x647 & n29026 ;
  assign n29084 = n29082 | n29083 ;
  assign n29085 = n15138 & n29084 ;
  assign n29086 = n29081 | n29085 ;
  assign n29087 = n29061 | n29086 ;
  assign n29088 = x787 & n29087 ;
  assign n29089 = n16115 & ~n29076 ;
  assign n29090 = ( x626 & ~n15419 ) | ( x626 & n29026 ) | ( ~n15419 & n29026 ) ;
  assign n29091 = ( x626 & n15419 ) | ( x626 & ~n29054 ) | ( n15419 & ~n29054 ) ;
  assign n29092 = ~n29090 & n29091 ;
  assign n29093 = n29089 | n29092 ;
  assign n29094 = ( x626 & n15418 ) | ( x626 & ~n29026 ) | ( n15418 & ~n29026 ) ;
  assign n29095 = ( x626 & ~n15418 ) | ( x626 & n29054 ) | ( ~n15418 & n29054 ) ;
  assign n29096 = n29094 & ~n29095 ;
  assign n29097 = n29093 | n29096 ;
  assign n29098 = x788 & n29097 ;
  assign n29099 = x648 & ~n29051 ;
  assign n29100 = ( x619 & x1159 ) | ( x619 & n29075 ) | ( x1159 & n29075 ) ;
  assign n29101 = x627 | n29041 ;
  assign n29102 = ( x618 & x1154 ) | ( x618 & ~n29074 ) | ( x1154 & ~n29074 ) ;
  assign n29103 = x660 | n29033 ;
  assign n29104 = ( x609 & x1155 ) | ( x609 & ~n29073 ) | ( x1155 & ~n29073 ) ;
  assign n29105 = n14839 | n29064 ;
  assign n29106 = x625 & ~n29105 ;
  assign n29107 = n29028 & n29105 ;
  assign n29108 = n29106 | n29107 ;
  assign n29109 = n29069 & n29108 ;
  assign n29110 = x608 | n29068 ;
  assign n29111 = n29109 | n29110 ;
  assign n29112 = x1153 & n29028 ;
  assign n29113 = ~n29106 & n29112 ;
  assign n29114 = x608 & ~n29070 ;
  assign n29115 = ~n29113 & n29114 ;
  assign n29116 = n29111 & ~n29115 ;
  assign n29117 = x778 & ~n29116 ;
  assign n29118 = x778 | n29107 ;
  assign n29119 = ~n29117 & n29118 ;
  assign n29120 = ( x609 & ~x1155 ) | ( x609 & n29119 ) | ( ~x1155 & n29119 ) ;
  assign n29121 = ~n29104 & n29120 ;
  assign n29122 = n29103 | n29121 ;
  assign n29123 = x660 & ~n29035 ;
  assign n29124 = ( x609 & x1155 ) | ( x609 & n29073 ) | ( x1155 & n29073 ) ;
  assign n29125 = ( ~x609 & x1155 ) | ( ~x609 & n29119 ) | ( x1155 & n29119 ) ;
  assign n29126 = n29124 & n29125 ;
  assign n29127 = n29123 & ~n29126 ;
  assign n29128 = n29122 & ~n29127 ;
  assign n29129 = x785 & ~n29128 ;
  assign n29130 = x785 | n29119 ;
  assign n29131 = ~n29129 & n29130 ;
  assign n29132 = ( x618 & ~x1154 ) | ( x618 & n29131 ) | ( ~x1154 & n29131 ) ;
  assign n29133 = ~n29102 & n29132 ;
  assign n29134 = n29101 | n29133 ;
  assign n29135 = x627 & ~n29043 ;
  assign n29136 = ( x618 & x1154 ) | ( x618 & n29074 ) | ( x1154 & n29074 ) ;
  assign n29137 = ( ~x618 & x1154 ) | ( ~x618 & n29131 ) | ( x1154 & n29131 ) ;
  assign n29138 = n29136 & n29137 ;
  assign n29139 = n29135 & ~n29138 ;
  assign n29140 = n29134 & ~n29139 ;
  assign n29141 = x781 & ~n29140 ;
  assign n29142 = x781 | n29131 ;
  assign n29143 = ~n29141 & n29142 ;
  assign n29144 = ( ~x619 & x1159 ) | ( ~x619 & n29143 ) | ( x1159 & n29143 ) ;
  assign n29145 = n29100 & n29144 ;
  assign n29146 = n29099 & ~n29145 ;
  assign n29147 = x648 | n29049 ;
  assign n29148 = ( x619 & x1159 ) | ( x619 & ~n29075 ) | ( x1159 & ~n29075 ) ;
  assign n29149 = ( x619 & ~x1159 ) | ( x619 & n29143 ) | ( ~x1159 & n29143 ) ;
  assign n29150 = ~n29148 & n29149 ;
  assign n29151 = n29147 | n29150 ;
  assign n29152 = x789 & n29151 ;
  assign n29153 = ~n29146 & n29152 ;
  assign n29154 = ~x789 & n29143 ;
  assign n29155 = n16177 | n29154 ;
  assign n29156 = n29153 | n29155 ;
  assign n29157 = ~n29098 & n29156 ;
  assign n29158 = n18434 | n29157 ;
  assign n29159 = n16650 | n29077 ;
  assign n29160 = n16051 & ~n29057 ;
  assign n29161 = n29159 & ~n29160 ;
  assign n29162 = ( x629 & ~x792 ) | ( x629 & n29161 ) | ( ~x792 & n29161 ) ;
  assign n29163 = n16052 & ~n29057 ;
  assign n29164 = n16643 & ~n29077 ;
  assign n29165 = n29163 | n29164 ;
  assign n29166 = ( x629 & x792 ) | ( x629 & n29165 ) | ( x792 & n29165 ) ;
  assign n29167 = ~n29162 & n29166 ;
  assign n29168 = n18431 | n29167 ;
  assign n29169 = n29158 & ~n29168 ;
  assign n29170 = n29088 | n29169 ;
  assign n29171 = ( x790 & x832 ) | ( x790 & n29170 ) | ( x832 & n29170 ) ;
  assign n29172 = n15141 | n29060 ;
  assign n29173 = n15141 & ~n29026 ;
  assign n29174 = n29172 & ~n29173 ;
  assign n29175 = ( x644 & x715 ) | ( x644 & ~n29174 ) | ( x715 & ~n29174 ) ;
  assign n29176 = ( x644 & ~x715 ) | ( x644 & n29026 ) | ( ~x715 & n29026 ) ;
  assign n29177 = ~n29175 & n29176 ;
  assign n29178 = x1160 & ~n29177 ;
  assign n29179 = ~x787 & n29078 ;
  assign n29180 = x1157 & n29084 ;
  assign n29181 = n29080 | n29180 ;
  assign n29182 = x787 & n29181 ;
  assign n29183 = n29179 | n29182 ;
  assign n29184 = ( x644 & x715 ) | ( x644 & n29183 ) | ( x715 & n29183 ) ;
  assign n29185 = ( ~x644 & x715 ) | ( ~x644 & n29170 ) | ( x715 & n29170 ) ;
  assign n29186 = n29184 & n29185 ;
  assign n29187 = n29178 & ~n29186 ;
  assign n29188 = ( x644 & x715 ) | ( x644 & n29174 ) | ( x715 & n29174 ) ;
  assign n29189 = ( ~x644 & x715 ) | ( ~x644 & n29026 ) | ( x715 & n29026 ) ;
  assign n29190 = n29188 & n29189 ;
  assign n29191 = x1160 | n29190 ;
  assign n29192 = ( x644 & x715 ) | ( x644 & ~n29183 ) | ( x715 & ~n29183 ) ;
  assign n29193 = ( x644 & ~x715 ) | ( x644 & n29170 ) | ( ~x715 & n29170 ) ;
  assign n29194 = ~n29192 & n29193 ;
  assign n29195 = n29191 | n29194 ;
  assign n29196 = ~n29187 & n29195 ;
  assign n29197 = ( ~x790 & x832 ) | ( ~x790 & n29196 ) | ( x832 & n29196 ) ;
  assign n29198 = n29171 & n29197 ;
  assign n29199 = x192 | n14834 ;
  assign n29200 = n15414 & n29199 ;
  assign n29201 = x192 & n2032 ;
  assign n29202 = x192 | n15070 ;
  assign n29203 = n15375 & n29202 ;
  assign n29204 = x691 & ~n29203 ;
  assign n29205 = ( ~x38 & x192 ) | ( ~x38 & n16319 ) | ( x192 & n16319 ) ;
  assign n29206 = ( x38 & x192 ) | ( x38 & n16323 ) | ( x192 & n16323 ) ;
  assign n29207 = n29205 & ~n29206 ;
  assign n29208 = n29204 & ~n29207 ;
  assign n29209 = x192 | x691 ;
  assign n29210 = n15382 | n29209 ;
  assign n29211 = ~n2032 & n29210 ;
  assign n29212 = ~n29208 & n29211 ;
  assign n29213 = n29201 | n29212 ;
  assign n29214 = ~x778 & n29213 ;
  assign n29215 = ( x625 & x1153 ) | ( x625 & n29199 ) | ( x1153 & n29199 ) ;
  assign n29216 = ( ~x625 & x1153 ) | ( ~x625 & n29213 ) | ( x1153 & n29213 ) ;
  assign n29217 = n29215 & n29216 ;
  assign n29218 = ( x625 & x1153 ) | ( x625 & ~n29199 ) | ( x1153 & ~n29199 ) ;
  assign n29219 = ( x625 & ~x1153 ) | ( x625 & n29213 ) | ( ~x1153 & n29213 ) ;
  assign n29220 = ~n29218 & n29219 ;
  assign n29221 = n29217 | n29220 ;
  assign n29222 = x778 & n29221 ;
  assign n29223 = n29214 | n29222 ;
  assign n29224 = ~n15400 & n29223 ;
  assign n29225 = n15400 & n29199 ;
  assign n29226 = n29224 | n29225 ;
  assign n29227 = n15407 | n29226 ;
  assign n29228 = n15407 & ~n29199 ;
  assign n29229 = n29227 & ~n29228 ;
  assign n29230 = ~n15414 & n29229 ;
  assign n29231 = n29200 | n29230 ;
  assign n29232 = n15421 | n29231 ;
  assign n29233 = n15421 & ~n29199 ;
  assign n29234 = n29232 & ~n29233 ;
  assign n29235 = x792 | n29234 ;
  assign n29236 = x628 & ~n29234 ;
  assign n29237 = x628 | n29199 ;
  assign n29238 = ~n29236 & n29237 ;
  assign n29239 = ( ~x792 & x1156 ) | ( ~x792 & n29238 ) | ( x1156 & n29238 ) ;
  assign n29240 = x628 | n29234 ;
  assign n29241 = x628 & ~n29199 ;
  assign n29242 = n29240 & ~n29241 ;
  assign n29243 = ( x792 & x1156 ) | ( x792 & ~n29242 ) | ( x1156 & ~n29242 ) ;
  assign n29244 = ~n29239 & n29243 ;
  assign n29245 = n29235 & ~n29244 ;
  assign n29246 = x787 | n29245 ;
  assign n29247 = x647 & ~n29245 ;
  assign n29248 = x647 | n29199 ;
  assign n29249 = ~n29247 & n29248 ;
  assign n29250 = ( ~x787 & x1157 ) | ( ~x787 & n29249 ) | ( x1157 & n29249 ) ;
  assign n29251 = x647 | n29245 ;
  assign n29252 = x647 & ~n29199 ;
  assign n29253 = n29251 & ~n29252 ;
  assign n29254 = ( x787 & x1157 ) | ( x787 & ~n29253 ) | ( x1157 & ~n29253 ) ;
  assign n29255 = ~n29250 & n29254 ;
  assign n29256 = n29246 & ~n29255 ;
  assign n29257 = x644 | n29256 ;
  assign n29258 = x715 & n29257 ;
  assign n29259 = ~x764 & n14710 ;
  assign n29260 = x192 & ~n14907 ;
  assign n29261 = n29259 | n29260 ;
  assign n29262 = x39 & n29261 ;
  assign n29263 = ~x192 & x764 ;
  assign n29264 = n15063 & n29263 ;
  assign n29265 = x764 & n14932 ;
  assign n29266 = x192 & ~n29265 ;
  assign n29267 = n20522 | n29266 ;
  assign n29268 = n29264 | n29267 ;
  assign n29269 = n29262 | n29268 ;
  assign n29270 = ~x38 & n29269 ;
  assign n29271 = x764 & n15072 ;
  assign n29272 = x38 & n29202 ;
  assign n29273 = ~n29271 & n29272 ;
  assign n29274 = n29270 | n29273 ;
  assign n29275 = ~n2032 & n29274 ;
  assign n29276 = n29201 | n29275 ;
  assign n29277 = ~n15082 & n29276 ;
  assign n29278 = n15082 & n29199 ;
  assign n29279 = n29277 | n29278 ;
  assign n29280 = ~x785 & n29279 ;
  assign n29281 = ~n15088 & n29199 ;
  assign n29282 = x609 & n29277 ;
  assign n29283 = n29281 | n29282 ;
  assign n29284 = x1155 & n29283 ;
  assign n29285 = n15094 & n29199 ;
  assign n29286 = ~x609 & n29277 ;
  assign n29287 = n29285 | n29286 ;
  assign n29288 = ~x1155 & n29287 ;
  assign n29289 = n29284 | n29288 ;
  assign n29290 = x785 & n29289 ;
  assign n29291 = n29280 | n29290 ;
  assign n29292 = ~x781 & n29291 ;
  assign n29293 = ( x618 & x1154 ) | ( x618 & n29199 ) | ( x1154 & n29199 ) ;
  assign n29294 = ( ~x618 & x1154 ) | ( ~x618 & n29291 ) | ( x1154 & n29291 ) ;
  assign n29295 = n29293 & n29294 ;
  assign n29296 = ( x618 & x1154 ) | ( x618 & ~n29199 ) | ( x1154 & ~n29199 ) ;
  assign n29297 = ( x618 & ~x1154 ) | ( x618 & n29291 ) | ( ~x1154 & n29291 ) ;
  assign n29298 = ~n29296 & n29297 ;
  assign n29299 = n29295 | n29298 ;
  assign n29300 = x781 & n29299 ;
  assign n29301 = n29292 | n29300 ;
  assign n29302 = ~x789 & n29301 ;
  assign n29303 = ( x619 & x1159 ) | ( x619 & n29199 ) | ( x1159 & n29199 ) ;
  assign n29304 = ( ~x619 & x1159 ) | ( ~x619 & n29301 ) | ( x1159 & n29301 ) ;
  assign n29305 = n29303 & n29304 ;
  assign n29306 = ( x619 & x1159 ) | ( x619 & ~n29199 ) | ( x1159 & ~n29199 ) ;
  assign n29307 = ( x619 & ~x1159 ) | ( x619 & n29301 ) | ( ~x1159 & n29301 ) ;
  assign n29308 = ~n29306 & n29307 ;
  assign n29309 = n29305 | n29308 ;
  assign n29310 = x789 & n29309 ;
  assign n29311 = n29302 | n29310 ;
  assign n29312 = n16176 | n29311 ;
  assign n29313 = n16176 & ~n29199 ;
  assign n29314 = n29312 & ~n29313 ;
  assign n29315 = n15134 | n29314 ;
  assign n29316 = n15134 & ~n29199 ;
  assign n29317 = n29315 & ~n29316 ;
  assign n29318 = n15141 | n29317 ;
  assign n29319 = n15141 & ~n29199 ;
  assign n29320 = n29318 & ~n29319 ;
  assign n29321 = ( x644 & x715 ) | ( x644 & ~n29320 ) | ( x715 & ~n29320 ) ;
  assign n29322 = ( x644 & ~x715 ) | ( x644 & n29199 ) | ( ~x715 & n29199 ) ;
  assign n29323 = ~n29321 & n29322 ;
  assign n29324 = x1160 & ~n29323 ;
  assign n29325 = ~n29258 & n29324 ;
  assign n29326 = x644 & ~n29256 ;
  assign n29327 = x715 | n29326 ;
  assign n29328 = ( x644 & x715 ) | ( x644 & n29320 ) | ( x715 & n29320 ) ;
  assign n29329 = ( ~x644 & x715 ) | ( ~x644 & n29199 ) | ( x715 & n29199 ) ;
  assign n29330 = n29328 & n29329 ;
  assign n29331 = x1160 | n29330 ;
  assign n29332 = n29327 & ~n29331 ;
  assign n29333 = n29325 | n29332 ;
  assign n29334 = x790 & n29333 ;
  assign n29335 = n18621 & n29314 ;
  assign n29336 = n15132 & n29242 ;
  assign n29337 = n15131 & n29238 ;
  assign n29338 = n29336 | n29337 ;
  assign n29339 = n29335 | n29338 ;
  assign n29340 = x792 & n29339 ;
  assign n29341 = x648 & ~n29308 ;
  assign n29342 = ( x619 & x1159 ) | ( x619 & n29229 ) | ( x1159 & n29229 ) ;
  assign n29343 = x627 | n29295 ;
  assign n29344 = ( x618 & x1154 ) | ( x618 & ~n29226 ) | ( x1154 & ~n29226 ) ;
  assign n29345 = x660 | n29284 ;
  assign n29346 = ( x609 & x1155 ) | ( x609 & ~n29223 ) | ( x1155 & ~n29223 ) ;
  assign n29347 = x608 | n29217 ;
  assign n29348 = ( x625 & x1153 ) | ( x625 & ~n29276 ) | ( x1153 & ~n29276 ) ;
  assign n29349 = x691 | n29274 ;
  assign n29350 = ( x192 & ~x764 ) | ( x192 & n15872 ) | ( ~x764 & n15872 ) ;
  assign n29351 = ( x192 & x764 ) | ( x192 & n15797 ) | ( x764 & n15797 ) ;
  assign n29352 = ~n29350 & n29351 ;
  assign n29353 = x39 & ~n29352 ;
  assign n29354 = ( x192 & ~x764 ) | ( x192 & n15699 ) | ( ~x764 & n15699 ) ;
  assign n29355 = ( x192 & x764 ) | ( x192 & n15583 ) | ( x764 & n15583 ) ;
  assign n29356 = n29354 & ~n29355 ;
  assign n29357 = n29353 & ~n29356 ;
  assign n29358 = ( x192 & ~x764 ) | ( x192 & n15891 ) | ( ~x764 & n15891 ) ;
  assign n29359 = ( x192 & x764 ) | ( x192 & n15887 ) | ( x764 & n15887 ) ;
  assign n29360 = n29358 & ~n29359 ;
  assign n29361 = ( x192 & ~x764 ) | ( x192 & n15897 ) | ( ~x764 & n15897 ) ;
  assign n29362 = ( x192 & x764 ) | ( x192 & n15894 ) | ( x764 & n15894 ) ;
  assign n29363 = ~n29361 & n29362 ;
  assign n29364 = n29360 | n29363 ;
  assign n29365 = ( ~x38 & n9138 ) | ( ~x38 & n29364 ) | ( n9138 & n29364 ) ;
  assign n29366 = ~n29357 & n29365 ;
  assign n29367 = ~x764 & n22085 ;
  assign n29368 = n15758 | n29367 ;
  assign n29369 = ~x39 & n29368 ;
  assign n29370 = x192 | n29369 ;
  assign n29371 = n15529 | n29027 ;
  assign n29372 = x192 & n29371 ;
  assign n29373 = ~n4810 & n29372 ;
  assign n29374 = x38 & ~n29373 ;
  assign n29375 = n29370 & n29374 ;
  assign n29376 = x691 & ~n29375 ;
  assign n29377 = ~n29366 & n29376 ;
  assign n29378 = n2032 | n29377 ;
  assign n29379 = n29349 & ~n29378 ;
  assign n29380 = n29201 | n29379 ;
  assign n29381 = ( x625 & ~x1153 ) | ( x625 & n29380 ) | ( ~x1153 & n29380 ) ;
  assign n29382 = ~n29348 & n29381 ;
  assign n29383 = n29347 | n29382 ;
  assign n29384 = x608 & ~n29220 ;
  assign n29385 = ( x625 & x1153 ) | ( x625 & n29276 ) | ( x1153 & n29276 ) ;
  assign n29386 = ( ~x625 & x1153 ) | ( ~x625 & n29380 ) | ( x1153 & n29380 ) ;
  assign n29387 = n29385 & n29386 ;
  assign n29388 = n29384 & ~n29387 ;
  assign n29389 = n29383 & ~n29388 ;
  assign n29390 = x778 & ~n29389 ;
  assign n29391 = x778 | n29380 ;
  assign n29392 = ~n29390 & n29391 ;
  assign n29393 = ( x609 & ~x1155 ) | ( x609 & n29392 ) | ( ~x1155 & n29392 ) ;
  assign n29394 = ~n29346 & n29393 ;
  assign n29395 = n29345 | n29394 ;
  assign n29396 = x660 & ~n29288 ;
  assign n29397 = ( x609 & x1155 ) | ( x609 & n29223 ) | ( x1155 & n29223 ) ;
  assign n29398 = ( ~x609 & x1155 ) | ( ~x609 & n29392 ) | ( x1155 & n29392 ) ;
  assign n29399 = n29397 & n29398 ;
  assign n29400 = n29396 & ~n29399 ;
  assign n29401 = n29395 & ~n29400 ;
  assign n29402 = x785 & ~n29401 ;
  assign n29403 = x785 | n29392 ;
  assign n29404 = ~n29402 & n29403 ;
  assign n29405 = ( x618 & ~x1154 ) | ( x618 & n29404 ) | ( ~x1154 & n29404 ) ;
  assign n29406 = ~n29344 & n29405 ;
  assign n29407 = n29343 | n29406 ;
  assign n29408 = x627 & ~n29298 ;
  assign n29409 = ( x618 & x1154 ) | ( x618 & n29226 ) | ( x1154 & n29226 ) ;
  assign n29410 = ( ~x618 & x1154 ) | ( ~x618 & n29404 ) | ( x1154 & n29404 ) ;
  assign n29411 = n29409 & n29410 ;
  assign n29412 = n29408 & ~n29411 ;
  assign n29413 = n29407 & ~n29412 ;
  assign n29414 = x781 & ~n29413 ;
  assign n29415 = x781 | n29404 ;
  assign n29416 = ~n29414 & n29415 ;
  assign n29417 = ( ~x619 & x1159 ) | ( ~x619 & n29416 ) | ( x1159 & n29416 ) ;
  assign n29418 = n29342 & n29417 ;
  assign n29419 = n29341 & ~n29418 ;
  assign n29420 = x648 | n29305 ;
  assign n29421 = ( x619 & x1159 ) | ( x619 & ~n29229 ) | ( x1159 & ~n29229 ) ;
  assign n29422 = ( x619 & ~x1159 ) | ( x619 & n29416 ) | ( ~x1159 & n29416 ) ;
  assign n29423 = ~n29421 & n29422 ;
  assign n29424 = n29420 | n29423 ;
  assign n29425 = x789 & n29424 ;
  assign n29426 = ~n29419 & n29425 ;
  assign n29427 = ~x789 & n29416 ;
  assign n29428 = n16177 | n29427 ;
  assign n29429 = n29426 | n29428 ;
  assign n29430 = n16115 & ~n29231 ;
  assign n29431 = ( x626 & ~n15419 ) | ( x626 & n29199 ) | ( ~n15419 & n29199 ) ;
  assign n29432 = ( x626 & n15419 ) | ( x626 & ~n29311 ) | ( n15419 & ~n29311 ) ;
  assign n29433 = ~n29431 & n29432 ;
  assign n29434 = n29430 | n29433 ;
  assign n29435 = ( x626 & n15418 ) | ( x626 & ~n29199 ) | ( n15418 & ~n29199 ) ;
  assign n29436 = ( x626 & ~n15418 ) | ( x626 & n29311 ) | ( ~n15418 & n29311 ) ;
  assign n29437 = n29435 & ~n29436 ;
  assign n29438 = n29434 | n29437 ;
  assign n29439 = x788 & n29438 ;
  assign n29440 = n18434 | n29439 ;
  assign n29441 = n29429 & ~n29440 ;
  assign n29442 = n29340 | n29441 ;
  assign n29443 = ~n18431 & n29442 ;
  assign n29444 = n15138 & n29249 ;
  assign n29445 = n15139 & n29253 ;
  assign n29446 = n18610 & n29317 ;
  assign n29447 = n29445 | n29446 ;
  assign n29448 = n29444 | n29447 ;
  assign n29449 = x787 & n29448 ;
  assign n29450 = n29443 | n29449 ;
  assign n29451 = ( x644 & ~x790 ) | ( x644 & n29324 ) | ( ~x790 & n29324 ) ;
  assign n29452 = ( x644 & x790 ) | ( x644 & n29331 ) | ( x790 & n29331 ) ;
  assign n29453 = ~n29451 & n29452 ;
  assign n29454 = n29450 | n29453 ;
  assign n29455 = ~n29334 & n29454 ;
  assign n29456 = ( ~x832 & n6785 ) | ( ~x832 & n29455 ) | ( n6785 & n29455 ) ;
  assign n29457 = ( ~x192 & x832 ) | ( ~x192 & n6785 ) | ( x832 & n6785 ) ;
  assign n29458 = n29456 & ~n29457 ;
  assign n29459 = n29198 | n29458 ;
  assign n29460 = x193 | n1290 ;
  assign n29461 = x739 & n14840 ;
  assign n29462 = n29460 & ~n29461 ;
  assign n29463 = n16060 | n29462 ;
  assign n29464 = ~x785 & n29463 ;
  assign n29465 = ~n15094 & n29461 ;
  assign n29466 = n29463 | n29465 ;
  assign n29467 = x1155 & n29466 ;
  assign n29468 = ~x1155 & n29460 ;
  assign n29469 = ~n29465 & n29468 ;
  assign n29470 = n29467 | n29469 ;
  assign n29471 = x785 & n29470 ;
  assign n29472 = n29464 | n29471 ;
  assign n29473 = ~x781 & n29472 ;
  assign n29474 = n16075 | n29472 ;
  assign n29475 = x1154 & n29474 ;
  assign n29476 = n16078 | n29472 ;
  assign n29477 = ~x1154 & n29476 ;
  assign n29478 = n29475 | n29477 ;
  assign n29479 = x781 & n29478 ;
  assign n29480 = n29473 | n29479 ;
  assign n29481 = ~x789 & n29480 ;
  assign n29482 = n20948 | n29480 ;
  assign n29483 = x1159 & n29482 ;
  assign n29484 = n20951 | n29480 ;
  assign n29485 = ~x1159 & n29484 ;
  assign n29486 = n29483 | n29485 ;
  assign n29487 = x789 & n29486 ;
  assign n29488 = n29481 | n29487 ;
  assign n29489 = n16176 | n29488 ;
  assign n29490 = n16176 & ~n29460 ;
  assign n29491 = n29489 & ~n29490 ;
  assign n29492 = n15134 | n29491 ;
  assign n29493 = n15134 & ~n29460 ;
  assign n29494 = n29492 & ~n29493 ;
  assign n29495 = n18610 & n29494 ;
  assign n29496 = ( x647 & x1157 ) | ( x647 & ~n29460 ) | ( x1157 & ~n29460 ) ;
  assign n29497 = x690 & n15202 ;
  assign n29498 = n29460 & ~n29497 ;
  assign n29499 = x778 | n29498 ;
  assign n29500 = ~x625 & n29497 ;
  assign n29501 = n29498 | n29500 ;
  assign n29502 = x1153 & n29501 ;
  assign n29503 = ~x1153 & n29460 ;
  assign n29504 = ~n29500 & n29503 ;
  assign n29505 = x778 & ~n29504 ;
  assign n29506 = ~n29502 & n29505 ;
  assign n29507 = n29499 & ~n29506 ;
  assign n29508 = n16043 | n29507 ;
  assign n29509 = n16045 | n29508 ;
  assign n29510 = n16047 | n29509 ;
  assign n29511 = n16049 | n29510 ;
  assign n29512 = n16055 | n29511 ;
  assign n29513 = ( x647 & ~x1157 ) | ( x647 & n29512 ) | ( ~x1157 & n29512 ) ;
  assign n29514 = ~n29496 & n29513 ;
  assign n29515 = x630 & n29514 ;
  assign n29516 = x647 & n29512 ;
  assign n29517 = ~x647 & n29460 ;
  assign n29518 = n29516 | n29517 ;
  assign n29519 = n15138 & n29518 ;
  assign n29520 = n29515 | n29519 ;
  assign n29521 = n29495 | n29520 ;
  assign n29522 = x787 & n29521 ;
  assign n29523 = n16115 & ~n29510 ;
  assign n29524 = ( x626 & ~n15419 ) | ( x626 & n29460 ) | ( ~n15419 & n29460 ) ;
  assign n29525 = ( x626 & n15419 ) | ( x626 & ~n29488 ) | ( n15419 & ~n29488 ) ;
  assign n29526 = ~n29524 & n29525 ;
  assign n29527 = n29523 | n29526 ;
  assign n29528 = ( x626 & n15418 ) | ( x626 & ~n29460 ) | ( n15418 & ~n29460 ) ;
  assign n29529 = ( x626 & ~n15418 ) | ( x626 & n29488 ) | ( ~n15418 & n29488 ) ;
  assign n29530 = n29528 & ~n29529 ;
  assign n29531 = n29527 | n29530 ;
  assign n29532 = x788 & n29531 ;
  assign n29533 = x648 & ~n29485 ;
  assign n29534 = ( x619 & x1159 ) | ( x619 & n29509 ) | ( x1159 & n29509 ) ;
  assign n29535 = x627 | n29475 ;
  assign n29536 = ( x618 & x1154 ) | ( x618 & ~n29508 ) | ( x1154 & ~n29508 ) ;
  assign n29537 = x660 | n29467 ;
  assign n29538 = ( x609 & x1155 ) | ( x609 & ~n29507 ) | ( x1155 & ~n29507 ) ;
  assign n29539 = n14839 | n29498 ;
  assign n29540 = x625 & ~n29539 ;
  assign n29541 = n29462 & n29539 ;
  assign n29542 = n29540 | n29541 ;
  assign n29543 = n29503 & n29542 ;
  assign n29544 = x608 | n29502 ;
  assign n29545 = n29543 | n29544 ;
  assign n29546 = x1153 & n29462 ;
  assign n29547 = ~n29540 & n29546 ;
  assign n29548 = x608 & ~n29504 ;
  assign n29549 = ~n29547 & n29548 ;
  assign n29550 = n29545 & ~n29549 ;
  assign n29551 = x778 & ~n29550 ;
  assign n29552 = x778 | n29541 ;
  assign n29553 = ~n29551 & n29552 ;
  assign n29554 = ( x609 & ~x1155 ) | ( x609 & n29553 ) | ( ~x1155 & n29553 ) ;
  assign n29555 = ~n29538 & n29554 ;
  assign n29556 = n29537 | n29555 ;
  assign n29557 = x660 & ~n29469 ;
  assign n29558 = ( x609 & x1155 ) | ( x609 & n29507 ) | ( x1155 & n29507 ) ;
  assign n29559 = ( ~x609 & x1155 ) | ( ~x609 & n29553 ) | ( x1155 & n29553 ) ;
  assign n29560 = n29558 & n29559 ;
  assign n29561 = n29557 & ~n29560 ;
  assign n29562 = n29556 & ~n29561 ;
  assign n29563 = x785 & ~n29562 ;
  assign n29564 = x785 | n29553 ;
  assign n29565 = ~n29563 & n29564 ;
  assign n29566 = ( x618 & ~x1154 ) | ( x618 & n29565 ) | ( ~x1154 & n29565 ) ;
  assign n29567 = ~n29536 & n29566 ;
  assign n29568 = n29535 | n29567 ;
  assign n29569 = x627 & ~n29477 ;
  assign n29570 = ( x618 & x1154 ) | ( x618 & n29508 ) | ( x1154 & n29508 ) ;
  assign n29571 = ( ~x618 & x1154 ) | ( ~x618 & n29565 ) | ( x1154 & n29565 ) ;
  assign n29572 = n29570 & n29571 ;
  assign n29573 = n29569 & ~n29572 ;
  assign n29574 = n29568 & ~n29573 ;
  assign n29575 = x781 & ~n29574 ;
  assign n29576 = x781 | n29565 ;
  assign n29577 = ~n29575 & n29576 ;
  assign n29578 = ( ~x619 & x1159 ) | ( ~x619 & n29577 ) | ( x1159 & n29577 ) ;
  assign n29579 = n29534 & n29578 ;
  assign n29580 = n29533 & ~n29579 ;
  assign n29581 = x648 | n29483 ;
  assign n29582 = ( x619 & x1159 ) | ( x619 & ~n29509 ) | ( x1159 & ~n29509 ) ;
  assign n29583 = ( x619 & ~x1159 ) | ( x619 & n29577 ) | ( ~x1159 & n29577 ) ;
  assign n29584 = ~n29582 & n29583 ;
  assign n29585 = n29581 | n29584 ;
  assign n29586 = x789 & n29585 ;
  assign n29587 = ~n29580 & n29586 ;
  assign n29588 = ~x789 & n29577 ;
  assign n29589 = n16177 | n29588 ;
  assign n29590 = n29587 | n29589 ;
  assign n29591 = ~n29532 & n29590 ;
  assign n29592 = n18434 | n29591 ;
  assign n29593 = n16650 | n29511 ;
  assign n29594 = n16051 & ~n29491 ;
  assign n29595 = n29593 & ~n29594 ;
  assign n29596 = ( x629 & ~x792 ) | ( x629 & n29595 ) | ( ~x792 & n29595 ) ;
  assign n29597 = n16052 & ~n29491 ;
  assign n29598 = n16643 & ~n29511 ;
  assign n29599 = n29597 | n29598 ;
  assign n29600 = ( x629 & x792 ) | ( x629 & n29599 ) | ( x792 & n29599 ) ;
  assign n29601 = ~n29596 & n29600 ;
  assign n29602 = n18431 | n29601 ;
  assign n29603 = n29592 & ~n29602 ;
  assign n29604 = n29522 | n29603 ;
  assign n29605 = ( x790 & x832 ) | ( x790 & n29604 ) | ( x832 & n29604 ) ;
  assign n29606 = n15141 | n29494 ;
  assign n29607 = n15141 & ~n29460 ;
  assign n29608 = n29606 & ~n29607 ;
  assign n29609 = ( x644 & x715 ) | ( x644 & ~n29608 ) | ( x715 & ~n29608 ) ;
  assign n29610 = ( x644 & ~x715 ) | ( x644 & n29460 ) | ( ~x715 & n29460 ) ;
  assign n29611 = ~n29609 & n29610 ;
  assign n29612 = x1160 & ~n29611 ;
  assign n29613 = ~x787 & n29512 ;
  assign n29614 = x1157 & n29518 ;
  assign n29615 = n29514 | n29614 ;
  assign n29616 = x787 & n29615 ;
  assign n29617 = n29613 | n29616 ;
  assign n29618 = ( x644 & x715 ) | ( x644 & n29617 ) | ( x715 & n29617 ) ;
  assign n29619 = ( ~x644 & x715 ) | ( ~x644 & n29604 ) | ( x715 & n29604 ) ;
  assign n29620 = n29618 & n29619 ;
  assign n29621 = n29612 & ~n29620 ;
  assign n29622 = ( x644 & x715 ) | ( x644 & n29608 ) | ( x715 & n29608 ) ;
  assign n29623 = ( ~x644 & x715 ) | ( ~x644 & n29460 ) | ( x715 & n29460 ) ;
  assign n29624 = n29622 & n29623 ;
  assign n29625 = x1160 | n29624 ;
  assign n29626 = ( x644 & x715 ) | ( x644 & ~n29617 ) | ( x715 & ~n29617 ) ;
  assign n29627 = ( x644 & ~x715 ) | ( x644 & n29604 ) | ( ~x715 & n29604 ) ;
  assign n29628 = ~n29626 & n29627 ;
  assign n29629 = n29625 | n29628 ;
  assign n29630 = ~n29621 & n29629 ;
  assign n29631 = ( ~x790 & x832 ) | ( ~x790 & n29630 ) | ( x832 & n29630 ) ;
  assign n29632 = n29605 & n29631 ;
  assign n29633 = x193 | n14834 ;
  assign n29634 = n15414 & n29633 ;
  assign n29635 = x690 & ~n2032 ;
  assign n29636 = n29633 | n29635 ;
  assign n29637 = x193 & n16323 ;
  assign n29638 = x38 | n29637 ;
  assign n29639 = ~n2032 & n29638 ;
  assign n29640 = x193 | n16319 ;
  assign n29641 = ~n29639 & n29640 ;
  assign n29642 = x193 | n15070 ;
  assign n29643 = n15375 & n29642 ;
  assign n29644 = x690 & ~n29643 ;
  assign n29645 = ~n29641 & n29644 ;
  assign n29646 = n29636 & ~n29645 ;
  assign n29647 = ~x778 & n29646 ;
  assign n29648 = ( x625 & x1153 ) | ( x625 & n29633 ) | ( x1153 & n29633 ) ;
  assign n29649 = ( ~x625 & x1153 ) | ( ~x625 & n29646 ) | ( x1153 & n29646 ) ;
  assign n29650 = n29648 & n29649 ;
  assign n29651 = ( x625 & x1153 ) | ( x625 & ~n29633 ) | ( x1153 & ~n29633 ) ;
  assign n29652 = ( x625 & ~x1153 ) | ( x625 & n29646 ) | ( ~x1153 & n29646 ) ;
  assign n29653 = ~n29651 & n29652 ;
  assign n29654 = n29650 | n29653 ;
  assign n29655 = x778 & n29654 ;
  assign n29656 = n29647 | n29655 ;
  assign n29657 = ~n15400 & n29656 ;
  assign n29658 = n15400 & n29633 ;
  assign n29659 = n29657 | n29658 ;
  assign n29660 = n15407 | n29659 ;
  assign n29661 = n15407 & ~n29633 ;
  assign n29662 = n29660 & ~n29661 ;
  assign n29663 = ~n15414 & n29662 ;
  assign n29664 = n29634 | n29663 ;
  assign n29665 = n15421 | n29664 ;
  assign n29666 = n15421 & ~n29633 ;
  assign n29667 = n29665 & ~n29666 ;
  assign n29668 = ~x792 & n29667 ;
  assign n29669 = ( x628 & x1156 ) | ( x628 & n29633 ) | ( x1156 & n29633 ) ;
  assign n29670 = ( ~x628 & x1156 ) | ( ~x628 & n29667 ) | ( x1156 & n29667 ) ;
  assign n29671 = n29669 & n29670 ;
  assign n29672 = ( x628 & x1156 ) | ( x628 & ~n29633 ) | ( x1156 & ~n29633 ) ;
  assign n29673 = ( x628 & ~x1156 ) | ( x628 & n29667 ) | ( ~x1156 & n29667 ) ;
  assign n29674 = ~n29672 & n29673 ;
  assign n29675 = n29671 | n29674 ;
  assign n29676 = x792 & n29675 ;
  assign n29677 = n29668 | n29676 ;
  assign n29678 = x787 | n29677 ;
  assign n29679 = x647 & n29677 ;
  assign n29680 = ~x647 & n29633 ;
  assign n29681 = n29679 | n29680 ;
  assign n29682 = ( ~x787 & x1157 ) | ( ~x787 & n29681 ) | ( x1157 & n29681 ) ;
  assign n29683 = ~x647 & n29677 ;
  assign n29684 = x647 & n29633 ;
  assign n29685 = n29683 | n29684 ;
  assign n29686 = ( x787 & x1157 ) | ( x787 & ~n29685 ) | ( x1157 & ~n29685 ) ;
  assign n29687 = ~n29682 & n29686 ;
  assign n29688 = n29678 & ~n29687 ;
  assign n29689 = x644 | n29688 ;
  assign n29690 = x715 & n29689 ;
  assign n29691 = x193 & n2032 ;
  assign n29692 = x739 & n15072 ;
  assign n29693 = n29642 & ~n29692 ;
  assign n29694 = x38 & ~n29693 ;
  assign n29695 = x193 | x739 ;
  assign n29696 = n14936 | n29695 ;
  assign n29697 = ( ~x193 & x739 ) | ( ~x193 & n14933 ) | ( x739 & n14933 ) ;
  assign n29698 = ( x193 & x739 ) | ( x193 & ~n15063 ) | ( x739 & ~n15063 ) ;
  assign n29699 = n29697 & n29698 ;
  assign n29700 = n29696 & ~n29699 ;
  assign n29701 = x38 | n29700 ;
  assign n29702 = ~n29694 & n29701 ;
  assign n29703 = ~n2032 & n29702 ;
  assign n29704 = n29691 | n29703 ;
  assign n29705 = ~n15082 & n29704 ;
  assign n29706 = n15082 & n29633 ;
  assign n29707 = n29705 | n29706 ;
  assign n29708 = ~x785 & n29707 ;
  assign n29709 = ~n15088 & n29633 ;
  assign n29710 = x609 & n29705 ;
  assign n29711 = n29709 | n29710 ;
  assign n29712 = x1155 & n29711 ;
  assign n29713 = n15094 & n29633 ;
  assign n29714 = ~x609 & n29705 ;
  assign n29715 = n29713 | n29714 ;
  assign n29716 = ~x1155 & n29715 ;
  assign n29717 = n29712 | n29716 ;
  assign n29718 = x785 & n29717 ;
  assign n29719 = n29708 | n29718 ;
  assign n29720 = ~x781 & n29719 ;
  assign n29721 = ( x618 & x1154 ) | ( x618 & n29633 ) | ( x1154 & n29633 ) ;
  assign n29722 = ( ~x618 & x1154 ) | ( ~x618 & n29719 ) | ( x1154 & n29719 ) ;
  assign n29723 = n29721 & n29722 ;
  assign n29724 = ( x618 & x1154 ) | ( x618 & ~n29633 ) | ( x1154 & ~n29633 ) ;
  assign n29725 = ( x618 & ~x1154 ) | ( x618 & n29719 ) | ( ~x1154 & n29719 ) ;
  assign n29726 = ~n29724 & n29725 ;
  assign n29727 = n29723 | n29726 ;
  assign n29728 = x781 & n29727 ;
  assign n29729 = n29720 | n29728 ;
  assign n29730 = ~x789 & n29729 ;
  assign n29731 = ( x619 & x1159 ) | ( x619 & n29633 ) | ( x1159 & n29633 ) ;
  assign n29732 = ( ~x619 & x1159 ) | ( ~x619 & n29729 ) | ( x1159 & n29729 ) ;
  assign n29733 = n29731 & n29732 ;
  assign n29734 = ( x619 & x1159 ) | ( x619 & ~n29633 ) | ( x1159 & ~n29633 ) ;
  assign n29735 = ( x619 & ~x1159 ) | ( x619 & n29729 ) | ( ~x1159 & n29729 ) ;
  assign n29736 = ~n29734 & n29735 ;
  assign n29737 = n29733 | n29736 ;
  assign n29738 = x789 & n29737 ;
  assign n29739 = n29730 | n29738 ;
  assign n29740 = n16176 | n29739 ;
  assign n29741 = n16176 & ~n29633 ;
  assign n29742 = n29740 & ~n29741 ;
  assign n29743 = n15134 | n29742 ;
  assign n29744 = n15134 & ~n29633 ;
  assign n29745 = n29743 & ~n29744 ;
  assign n29746 = n15141 | n29745 ;
  assign n29747 = n15141 & ~n29633 ;
  assign n29748 = n29746 & ~n29747 ;
  assign n29749 = ( x644 & x715 ) | ( x644 & ~n29748 ) | ( x715 & ~n29748 ) ;
  assign n29750 = ( x644 & ~x715 ) | ( x644 & n29633 ) | ( ~x715 & n29633 ) ;
  assign n29751 = ~n29749 & n29750 ;
  assign n29752 = x1160 & ~n29751 ;
  assign n29753 = ~n29690 & n29752 ;
  assign n29754 = x644 & ~n29688 ;
  assign n29755 = x715 | n29754 ;
  assign n29756 = ( x644 & x715 ) | ( x644 & n29748 ) | ( x715 & n29748 ) ;
  assign n29757 = ( ~x644 & x715 ) | ( ~x644 & n29633 ) | ( x715 & n29633 ) ;
  assign n29758 = n29756 & n29757 ;
  assign n29759 = x1160 | n29758 ;
  assign n29760 = n29755 & ~n29759 ;
  assign n29761 = n29753 | n29760 ;
  assign n29762 = x790 & n29761 ;
  assign n29763 = n18621 & n29742 ;
  assign n29764 = ( x629 & n29674 ) | ( x629 & n29763 ) | ( n29674 & n29763 ) ;
  assign n29765 = ( ~x629 & n29671 ) | ( ~x629 & n29763 ) | ( n29671 & n29763 ) ;
  assign n29766 = n29764 | n29765 ;
  assign n29767 = x792 & n29766 ;
  assign n29768 = x648 & ~n29736 ;
  assign n29769 = ( x619 & x1159 ) | ( x619 & n29662 ) | ( x1159 & n29662 ) ;
  assign n29770 = x627 | n29723 ;
  assign n29771 = ( x618 & x1154 ) | ( x618 & ~n29659 ) | ( x1154 & ~n29659 ) ;
  assign n29772 = x660 | n29712 ;
  assign n29773 = ( x609 & x1155 ) | ( x609 & ~n29656 ) | ( x1155 & ~n29656 ) ;
  assign n29774 = x608 | n29650 ;
  assign n29775 = ( x625 & x1153 ) | ( x625 & ~n29704 ) | ( x1153 & ~n29704 ) ;
  assign n29776 = x690 | n29702 ;
  assign n29777 = ( x193 & ~x739 ) | ( x193 & n15872 ) | ( ~x739 & n15872 ) ;
  assign n29778 = ( x193 & x739 ) | ( x193 & n15797 ) | ( x739 & n15797 ) ;
  assign n29779 = ~n29777 & n29778 ;
  assign n29780 = x39 & ~n29779 ;
  assign n29781 = ( x193 & ~x739 ) | ( x193 & n15699 ) | ( ~x739 & n15699 ) ;
  assign n29782 = ( x193 & x739 ) | ( x193 & n15583 ) | ( x739 & n15583 ) ;
  assign n29783 = n29781 & ~n29782 ;
  assign n29784 = n29780 & ~n29783 ;
  assign n29785 = ( ~x193 & x739 ) | ( ~x193 & n15897 ) | ( x739 & n15897 ) ;
  assign n29786 = ( x193 & x739 ) | ( x193 & ~n15894 ) | ( x739 & ~n15894 ) ;
  assign n29787 = n29785 & n29786 ;
  assign n29788 = ( ~x193 & x739 ) | ( ~x193 & n15891 ) | ( x739 & n15891 ) ;
  assign n29789 = ( x193 & x739 ) | ( x193 & ~n15887 ) | ( x739 & ~n15887 ) ;
  assign n29790 = n29788 | n29789 ;
  assign n29791 = ~n29787 & n29790 ;
  assign n29792 = x39 | n29791 ;
  assign n29793 = ~x38 & n29792 ;
  assign n29794 = ~n29784 & n29793 ;
  assign n29795 = ~x739 & n22085 ;
  assign n29796 = n15758 | n29795 ;
  assign n29797 = ~x39 & n29796 ;
  assign n29798 = x193 | n29797 ;
  assign n29799 = n15529 | n29461 ;
  assign n29800 = x193 & n29799 ;
  assign n29801 = ~n4810 & n29800 ;
  assign n29802 = x38 & ~n29801 ;
  assign n29803 = n29798 & n29802 ;
  assign n29804 = x690 & ~n29803 ;
  assign n29805 = ~n29794 & n29804 ;
  assign n29806 = n2032 | n29805 ;
  assign n29807 = n29776 & ~n29806 ;
  assign n29808 = n29691 | n29807 ;
  assign n29809 = ( x625 & ~x1153 ) | ( x625 & n29808 ) | ( ~x1153 & n29808 ) ;
  assign n29810 = ~n29775 & n29809 ;
  assign n29811 = n29774 | n29810 ;
  assign n29812 = x608 & ~n29653 ;
  assign n29813 = ( x625 & x1153 ) | ( x625 & n29704 ) | ( x1153 & n29704 ) ;
  assign n29814 = ( ~x625 & x1153 ) | ( ~x625 & n29808 ) | ( x1153 & n29808 ) ;
  assign n29815 = n29813 & n29814 ;
  assign n29816 = n29812 & ~n29815 ;
  assign n29817 = n29811 & ~n29816 ;
  assign n29818 = x778 & ~n29817 ;
  assign n29819 = x778 | n29808 ;
  assign n29820 = ~n29818 & n29819 ;
  assign n29821 = ( x609 & ~x1155 ) | ( x609 & n29820 ) | ( ~x1155 & n29820 ) ;
  assign n29822 = ~n29773 & n29821 ;
  assign n29823 = n29772 | n29822 ;
  assign n29824 = x660 & ~n29716 ;
  assign n29825 = ( x609 & x1155 ) | ( x609 & n29656 ) | ( x1155 & n29656 ) ;
  assign n29826 = ( ~x609 & x1155 ) | ( ~x609 & n29820 ) | ( x1155 & n29820 ) ;
  assign n29827 = n29825 & n29826 ;
  assign n29828 = n29824 & ~n29827 ;
  assign n29829 = n29823 & ~n29828 ;
  assign n29830 = x785 & ~n29829 ;
  assign n29831 = x785 | n29820 ;
  assign n29832 = ~n29830 & n29831 ;
  assign n29833 = ( x618 & ~x1154 ) | ( x618 & n29832 ) | ( ~x1154 & n29832 ) ;
  assign n29834 = ~n29771 & n29833 ;
  assign n29835 = n29770 | n29834 ;
  assign n29836 = x627 & ~n29726 ;
  assign n29837 = ( x618 & x1154 ) | ( x618 & n29659 ) | ( x1154 & n29659 ) ;
  assign n29838 = ( ~x618 & x1154 ) | ( ~x618 & n29832 ) | ( x1154 & n29832 ) ;
  assign n29839 = n29837 & n29838 ;
  assign n29840 = n29836 & ~n29839 ;
  assign n29841 = n29835 & ~n29840 ;
  assign n29842 = x781 & ~n29841 ;
  assign n29843 = x781 | n29832 ;
  assign n29844 = ~n29842 & n29843 ;
  assign n29845 = ( ~x619 & x1159 ) | ( ~x619 & n29844 ) | ( x1159 & n29844 ) ;
  assign n29846 = n29769 & n29845 ;
  assign n29847 = n29768 & ~n29846 ;
  assign n29848 = x648 | n29733 ;
  assign n29849 = ( x619 & x1159 ) | ( x619 & ~n29662 ) | ( x1159 & ~n29662 ) ;
  assign n29850 = ( x619 & ~x1159 ) | ( x619 & n29844 ) | ( ~x1159 & n29844 ) ;
  assign n29851 = ~n29849 & n29850 ;
  assign n29852 = n29848 | n29851 ;
  assign n29853 = x789 & n29852 ;
  assign n29854 = ~n29847 & n29853 ;
  assign n29855 = ~x789 & n29844 ;
  assign n29856 = n16177 | n29855 ;
  assign n29857 = n29854 | n29856 ;
  assign n29858 = n16115 & ~n29664 ;
  assign n29859 = ( x626 & ~n15419 ) | ( x626 & n29633 ) | ( ~n15419 & n29633 ) ;
  assign n29860 = ( x626 & n15419 ) | ( x626 & ~n29739 ) | ( n15419 & ~n29739 ) ;
  assign n29861 = ~n29859 & n29860 ;
  assign n29862 = n29858 | n29861 ;
  assign n29863 = ( x626 & n15418 ) | ( x626 & ~n29633 ) | ( n15418 & ~n29633 ) ;
  assign n29864 = ( x626 & ~n15418 ) | ( x626 & n29739 ) | ( ~n15418 & n29739 ) ;
  assign n29865 = n29863 & ~n29864 ;
  assign n29866 = n29862 | n29865 ;
  assign n29867 = x788 & n29866 ;
  assign n29868 = n18434 | n29867 ;
  assign n29869 = n29857 & ~n29868 ;
  assign n29870 = n29767 | n29869 ;
  assign n29871 = ~n18431 & n29870 ;
  assign n29872 = n18610 & n29745 ;
  assign n29873 = n15139 & n29685 ;
  assign n29874 = n15138 & n29681 ;
  assign n29875 = n29873 | n29874 ;
  assign n29876 = n29872 | n29875 ;
  assign n29877 = x787 & n29876 ;
  assign n29878 = n29871 | n29877 ;
  assign n29879 = ( x644 & ~x790 ) | ( x644 & n29752 ) | ( ~x790 & n29752 ) ;
  assign n29880 = ( x644 & x790 ) | ( x644 & n29759 ) | ( x790 & n29759 ) ;
  assign n29881 = ~n29879 & n29880 ;
  assign n29882 = n29878 | n29881 ;
  assign n29883 = ~n29762 & n29882 ;
  assign n29884 = ( ~x832 & n6785 ) | ( ~x832 & n29883 ) | ( n6785 & n29883 ) ;
  assign n29885 = ( ~x193 & x832 ) | ( ~x193 & n6785 ) | ( x832 & n6785 ) ;
  assign n29886 = n29884 & ~n29885 ;
  assign n29887 = n29632 | n29886 ;
  assign n29888 = x194 | n14834 ;
  assign n29889 = n15141 & n29888 ;
  assign n29890 = x194 & n2032 ;
  assign n29891 = x194 | n15382 ;
  assign n29892 = ~x748 & n29891 ;
  assign n29893 = ( x194 & ~x748 ) | ( x194 & n22415 ) | ( ~x748 & n22415 ) ;
  assign n29894 = ( x194 & x748 ) | ( x194 & n17421 ) | ( x748 & n17421 ) ;
  assign n29895 = ~n29893 & n29894 ;
  assign n29896 = n29892 | n29895 ;
  assign n29897 = ~n2032 & n29896 ;
  assign n29898 = n29890 | n29897 ;
  assign n29899 = ~n15082 & n29898 ;
  assign n29900 = n15082 & n29888 ;
  assign n29901 = n29899 | n29900 ;
  assign n29902 = ~x785 & n29901 ;
  assign n29903 = ~n15088 & n29888 ;
  assign n29904 = x609 & n29899 ;
  assign n29905 = n29903 | n29904 ;
  assign n29906 = x1155 & n29905 ;
  assign n29907 = n15094 & n29888 ;
  assign n29908 = ~x609 & n29899 ;
  assign n29909 = n29907 | n29908 ;
  assign n29910 = ~x1155 & n29909 ;
  assign n29911 = n29906 | n29910 ;
  assign n29912 = x785 & n29911 ;
  assign n29913 = n29902 | n29912 ;
  assign n29914 = ~x781 & n29913 ;
  assign n29915 = ( x618 & x1154 ) | ( x618 & n29888 ) | ( x1154 & n29888 ) ;
  assign n29916 = ( ~x618 & x1154 ) | ( ~x618 & n29913 ) | ( x1154 & n29913 ) ;
  assign n29917 = n29915 & n29916 ;
  assign n29918 = ( x618 & x1154 ) | ( x618 & ~n29888 ) | ( x1154 & ~n29888 ) ;
  assign n29919 = ( x618 & ~x1154 ) | ( x618 & n29913 ) | ( ~x1154 & n29913 ) ;
  assign n29920 = ~n29918 & n29919 ;
  assign n29921 = n29917 | n29920 ;
  assign n29922 = x781 & n29921 ;
  assign n29923 = n29914 | n29922 ;
  assign n29924 = ~x789 & n29923 ;
  assign n29925 = ( x619 & x1159 ) | ( x619 & n29888 ) | ( x1159 & n29888 ) ;
  assign n29926 = ( ~x619 & x1159 ) | ( ~x619 & n29923 ) | ( x1159 & n29923 ) ;
  assign n29927 = n29925 & n29926 ;
  assign n29928 = ( x619 & x1159 ) | ( x619 & ~n29888 ) | ( x1159 & ~n29888 ) ;
  assign n29929 = ( x619 & ~x1159 ) | ( x619 & n29923 ) | ( ~x1159 & n29923 ) ;
  assign n29930 = ~n29928 & n29929 ;
  assign n29931 = n29927 | n29930 ;
  assign n29932 = x789 & n29931 ;
  assign n29933 = n29924 | n29932 ;
  assign n29934 = n16176 | n29933 ;
  assign n29935 = n16176 & ~n29888 ;
  assign n29936 = n29934 & ~n29935 ;
  assign n29937 = n15134 | n29936 ;
  assign n29938 = n15134 & ~n29888 ;
  assign n29939 = n29937 & ~n29938 ;
  assign n29940 = ~n15141 & n29939 ;
  assign n29941 = n29889 | n29940 ;
  assign n29942 = ( x644 & x715 ) | ( x644 & n29941 ) | ( x715 & n29941 ) ;
  assign n29943 = ( ~x644 & x715 ) | ( ~x644 & n29888 ) | ( x715 & n29888 ) ;
  assign n29944 = n29942 & n29943 ;
  assign n29945 = x1160 | n29944 ;
  assign n29946 = n15414 & n29888 ;
  assign n29947 = x194 & ~n22357 ;
  assign n29948 = ( x730 & ~n2032 ) | ( x730 & n29891 ) | ( ~n2032 & n29891 ) ;
  assign n29949 = ~x194 & n22362 ;
  assign n29950 = ( x730 & n2032 ) | ( x730 & ~n29949 ) | ( n2032 & ~n29949 ) ;
  assign n29951 = n29948 & ~n29950 ;
  assign n29952 = n29947 | n29951 ;
  assign n29953 = ~x778 & n29952 ;
  assign n29954 = ( x625 & x1153 ) | ( x625 & n29888 ) | ( x1153 & n29888 ) ;
  assign n29955 = ( ~x625 & x1153 ) | ( ~x625 & n29952 ) | ( x1153 & n29952 ) ;
  assign n29956 = n29954 & n29955 ;
  assign n29957 = ( x625 & x1153 ) | ( x625 & ~n29888 ) | ( x1153 & ~n29888 ) ;
  assign n29958 = ( x625 & ~x1153 ) | ( x625 & n29952 ) | ( ~x1153 & n29952 ) ;
  assign n29959 = ~n29957 & n29958 ;
  assign n29960 = n29956 | n29959 ;
  assign n29961 = x778 & n29960 ;
  assign n29962 = n29953 | n29961 ;
  assign n29963 = ~n15400 & n29962 ;
  assign n29964 = n15400 & n29888 ;
  assign n29965 = n29963 | n29964 ;
  assign n29966 = n15407 | n29965 ;
  assign n29967 = n15407 & ~n29888 ;
  assign n29968 = n29966 & ~n29967 ;
  assign n29969 = ~n15414 & n29968 ;
  assign n29970 = n29946 | n29969 ;
  assign n29971 = n15421 | n29970 ;
  assign n29972 = n15421 & ~n29888 ;
  assign n29973 = n29971 & ~n29972 ;
  assign n29974 = ~x792 & n29973 ;
  assign n29975 = ( x628 & x1156 ) | ( x628 & n29888 ) | ( x1156 & n29888 ) ;
  assign n29976 = ( ~x628 & x1156 ) | ( ~x628 & n29973 ) | ( x1156 & n29973 ) ;
  assign n29977 = n29975 & n29976 ;
  assign n29978 = ( x628 & x1156 ) | ( x628 & ~n29888 ) | ( x1156 & ~n29888 ) ;
  assign n29979 = ( x628 & ~x1156 ) | ( x628 & n29973 ) | ( ~x1156 & n29973 ) ;
  assign n29980 = ~n29978 & n29979 ;
  assign n29981 = n29977 | n29980 ;
  assign n29982 = x792 & n29981 ;
  assign n29983 = n29974 | n29982 ;
  assign n29984 = ~x787 & n29983 ;
  assign n29985 = ( x647 & x1157 ) | ( x647 & n29888 ) | ( x1157 & n29888 ) ;
  assign n29986 = ( ~x647 & x1157 ) | ( ~x647 & n29983 ) | ( x1157 & n29983 ) ;
  assign n29987 = n29985 & n29986 ;
  assign n29988 = ( x647 & x1157 ) | ( x647 & ~n29888 ) | ( x1157 & ~n29888 ) ;
  assign n29989 = ( x647 & ~x1157 ) | ( x647 & n29983 ) | ( ~x1157 & n29983 ) ;
  assign n29990 = ~n29988 & n29989 ;
  assign n29991 = n29987 | n29990 ;
  assign n29992 = x787 & n29991 ;
  assign n29993 = n29984 | n29992 ;
  assign n29994 = ( x644 & x715 ) | ( x644 & ~n29993 ) | ( x715 & ~n29993 ) ;
  assign n29995 = x630 | n29987 ;
  assign n29996 = ( x647 & x1157 ) | ( x647 & ~n29939 ) | ( x1157 & ~n29939 ) ;
  assign n29997 = x629 | n29977 ;
  assign n29998 = ( x628 & x1156 ) | ( x628 & ~n29936 ) | ( x1156 & ~n29936 ) ;
  assign n29999 = x648 | n29927 ;
  assign n30000 = ( x619 & x1159 ) | ( x619 & ~n29968 ) | ( x1159 & ~n29968 ) ;
  assign n30001 = x627 | n29917 ;
  assign n30002 = ( x618 & x1154 ) | ( x618 & ~n29965 ) | ( x1154 & ~n29965 ) ;
  assign n30003 = x660 | n29906 ;
  assign n30004 = ( x609 & x1155 ) | ( x609 & ~n29962 ) | ( x1155 & ~n29962 ) ;
  assign n30005 = x608 | n29956 ;
  assign n30006 = ( x625 & x1153 ) | ( x625 & ~n29898 ) | ( x1153 & ~n29898 ) ;
  assign n30007 = ( x194 & ~x748 ) | ( x194 & n17562 ) | ( ~x748 & n17562 ) ;
  assign n30008 = ( x194 & x748 ) | ( x194 & n17554 ) | ( x748 & n17554 ) ;
  assign n30009 = ~n30007 & n30008 ;
  assign n30010 = x730 & ~n30009 ;
  assign n30011 = ( x194 & ~x748 ) | ( x194 & n17579 ) | ( ~x748 & n17579 ) ;
  assign n30012 = ( x194 & x748 ) | ( x194 & n22514 ) | ( x748 & n22514 ) ;
  assign n30013 = n30011 & ~n30012 ;
  assign n30014 = n30010 & ~n30013 ;
  assign n30015 = x730 | n29896 ;
  assign n30016 = ~n2032 & n30015 ;
  assign n30017 = ~n30014 & n30016 ;
  assign n30018 = n29890 | n30017 ;
  assign n30019 = ( x625 & ~x1153 ) | ( x625 & n30018 ) | ( ~x1153 & n30018 ) ;
  assign n30020 = ~n30006 & n30019 ;
  assign n30021 = n30005 | n30020 ;
  assign n30022 = x608 & ~n29959 ;
  assign n30023 = ( x625 & x1153 ) | ( x625 & n29898 ) | ( x1153 & n29898 ) ;
  assign n30024 = ( ~x625 & x1153 ) | ( ~x625 & n30018 ) | ( x1153 & n30018 ) ;
  assign n30025 = n30023 & n30024 ;
  assign n30026 = n30022 & ~n30025 ;
  assign n30027 = n30021 & ~n30026 ;
  assign n30028 = x778 & ~n30027 ;
  assign n30029 = x778 | n30018 ;
  assign n30030 = ~n30028 & n30029 ;
  assign n30031 = ( x609 & ~x1155 ) | ( x609 & n30030 ) | ( ~x1155 & n30030 ) ;
  assign n30032 = ~n30004 & n30031 ;
  assign n30033 = n30003 | n30032 ;
  assign n30034 = x660 & ~n29910 ;
  assign n30035 = ( x609 & x1155 ) | ( x609 & n29962 ) | ( x1155 & n29962 ) ;
  assign n30036 = ( ~x609 & x1155 ) | ( ~x609 & n30030 ) | ( x1155 & n30030 ) ;
  assign n30037 = n30035 & n30036 ;
  assign n30038 = n30034 & ~n30037 ;
  assign n30039 = n30033 & ~n30038 ;
  assign n30040 = x785 & ~n30039 ;
  assign n30041 = x785 | n30030 ;
  assign n30042 = ~n30040 & n30041 ;
  assign n30043 = ( x618 & ~x1154 ) | ( x618 & n30042 ) | ( ~x1154 & n30042 ) ;
  assign n30044 = ~n30002 & n30043 ;
  assign n30045 = n30001 | n30044 ;
  assign n30046 = x627 & ~n29920 ;
  assign n30047 = ( x618 & x1154 ) | ( x618 & n29965 ) | ( x1154 & n29965 ) ;
  assign n30048 = ( ~x618 & x1154 ) | ( ~x618 & n30042 ) | ( x1154 & n30042 ) ;
  assign n30049 = n30047 & n30048 ;
  assign n30050 = n30046 & ~n30049 ;
  assign n30051 = n30045 & ~n30050 ;
  assign n30052 = x781 & ~n30051 ;
  assign n30053 = x781 | n30042 ;
  assign n30054 = ~n30052 & n30053 ;
  assign n30055 = ( x619 & ~x1159 ) | ( x619 & n30054 ) | ( ~x1159 & n30054 ) ;
  assign n30056 = ~n30000 & n30055 ;
  assign n30057 = n29999 | n30056 ;
  assign n30058 = x648 & ~n29930 ;
  assign n30059 = ( x619 & x1159 ) | ( x619 & n29968 ) | ( x1159 & n29968 ) ;
  assign n30060 = ( ~x619 & x1159 ) | ( ~x619 & n30054 ) | ( x1159 & n30054 ) ;
  assign n30061 = n30059 & n30060 ;
  assign n30062 = n30058 & ~n30061 ;
  assign n30063 = n30057 & ~n30062 ;
  assign n30064 = x789 & ~n30063 ;
  assign n30065 = x789 | n30054 ;
  assign n30066 = ~n30064 & n30065 ;
  assign n30067 = ~x788 & n30066 ;
  assign n30068 = ( x626 & x641 ) | ( x626 & ~n29933 ) | ( x641 & ~n29933 ) ;
  assign n30069 = ( x626 & ~x641 ) | ( x626 & n29888 ) | ( ~x641 & n29888 ) ;
  assign n30070 = n30068 & ~n30069 ;
  assign n30071 = x1158 | n30070 ;
  assign n30072 = ( x626 & x641 ) | ( x626 & n29970 ) | ( x641 & n29970 ) ;
  assign n30073 = ( ~x626 & x641 ) | ( ~x626 & n30066 ) | ( x641 & n30066 ) ;
  assign n30074 = n30072 | n30073 ;
  assign n30075 = ~n30071 & n30074 ;
  assign n30076 = ( x626 & x641 ) | ( x626 & n29933 ) | ( x641 & n29933 ) ;
  assign n30077 = ( ~x626 & x641 ) | ( ~x626 & n29888 ) | ( x641 & n29888 ) ;
  assign n30078 = n30076 | n30077 ;
  assign n30079 = x1158 & n30078 ;
  assign n30080 = ( x626 & x641 ) | ( x626 & ~n29970 ) | ( x641 & ~n29970 ) ;
  assign n30081 = ( x626 & ~x641 ) | ( x626 & n30066 ) | ( ~x641 & n30066 ) ;
  assign n30082 = n30080 & ~n30081 ;
  assign n30083 = n30079 & ~n30082 ;
  assign n30084 = n30075 | n30083 ;
  assign n30085 = x788 & n30084 ;
  assign n30086 = n30067 | n30085 ;
  assign n30087 = ( x628 & ~x1156 ) | ( x628 & n30086 ) | ( ~x1156 & n30086 ) ;
  assign n30088 = ~n29998 & n30087 ;
  assign n30089 = n29997 | n30088 ;
  assign n30090 = x629 & ~n29980 ;
  assign n30091 = ( x628 & x1156 ) | ( x628 & n29936 ) | ( x1156 & n29936 ) ;
  assign n30092 = ( ~x628 & x1156 ) | ( ~x628 & n30086 ) | ( x1156 & n30086 ) ;
  assign n30093 = n30091 & n30092 ;
  assign n30094 = n30090 & ~n30093 ;
  assign n30095 = n30089 & ~n30094 ;
  assign n30096 = x792 & ~n30095 ;
  assign n30097 = x792 | n30086 ;
  assign n30098 = ~n30096 & n30097 ;
  assign n30099 = ( x647 & ~x1157 ) | ( x647 & n30098 ) | ( ~x1157 & n30098 ) ;
  assign n30100 = ~n29996 & n30099 ;
  assign n30101 = n29995 | n30100 ;
  assign n30102 = x630 & ~n29990 ;
  assign n30103 = ( x647 & x1157 ) | ( x647 & n29939 ) | ( x1157 & n29939 ) ;
  assign n30104 = ( ~x647 & x1157 ) | ( ~x647 & n30098 ) | ( x1157 & n30098 ) ;
  assign n30105 = n30103 & n30104 ;
  assign n30106 = n30102 & ~n30105 ;
  assign n30107 = n30101 & ~n30106 ;
  assign n30108 = x787 & ~n30107 ;
  assign n30109 = x787 | n30098 ;
  assign n30110 = ~n30108 & n30109 ;
  assign n30111 = ( x644 & ~x715 ) | ( x644 & n30110 ) | ( ~x715 & n30110 ) ;
  assign n30112 = ~n29994 & n30111 ;
  assign n30113 = n29945 | n30112 ;
  assign n30114 = ( x644 & x715 ) | ( x644 & ~n29941 ) | ( x715 & ~n29941 ) ;
  assign n30115 = ( x644 & ~x715 ) | ( x644 & n29888 ) | ( ~x715 & n29888 ) ;
  assign n30116 = ~n30114 & n30115 ;
  assign n30117 = x1160 & ~n30116 ;
  assign n30118 = ( x644 & x715 ) | ( x644 & n29993 ) | ( x715 & n29993 ) ;
  assign n30119 = ( ~x644 & x715 ) | ( ~x644 & n30110 ) | ( x715 & n30110 ) ;
  assign n30120 = n30118 & n30119 ;
  assign n30121 = n30117 & ~n30120 ;
  assign n30122 = x790 & ~n30121 ;
  assign n30123 = n30113 & n30122 ;
  assign n30124 = ~x790 & n30110 ;
  assign n30125 = n6785 | n30124 ;
  assign n30126 = n30123 | n30125 ;
  assign n30127 = ~x194 & n6785 ;
  assign n30128 = x832 | n30127 ;
  assign n30129 = n30126 & ~n30128 ;
  assign n30130 = x194 | n1290 ;
  assign n30131 = x748 & n14840 ;
  assign n30132 = n30130 & ~n30131 ;
  assign n30133 = n16060 | n30132 ;
  assign n30134 = ~x785 & n30133 ;
  assign n30135 = n16065 | n30132 ;
  assign n30136 = x1155 & n30135 ;
  assign n30137 = n16068 | n30133 ;
  assign n30138 = ~x1155 & n30137 ;
  assign n30139 = n30136 | n30138 ;
  assign n30140 = x785 & n30139 ;
  assign n30141 = n30134 | n30140 ;
  assign n30142 = ~x781 & n30141 ;
  assign n30143 = n16075 | n30141 ;
  assign n30144 = x1154 & n30143 ;
  assign n30145 = n16078 | n30141 ;
  assign n30146 = ~x1154 & n30145 ;
  assign n30147 = n30144 | n30146 ;
  assign n30148 = x781 & n30147 ;
  assign n30149 = n30142 | n30148 ;
  assign n30150 = ~x789 & n30149 ;
  assign n30151 = ( x619 & x1159 ) | ( x619 & n30130 ) | ( x1159 & n30130 ) ;
  assign n30152 = ( ~x619 & x1159 ) | ( ~x619 & n30149 ) | ( x1159 & n30149 ) ;
  assign n30153 = n30151 & n30152 ;
  assign n30154 = ( x619 & x1159 ) | ( x619 & ~n30130 ) | ( x1159 & ~n30130 ) ;
  assign n30155 = ( x619 & ~x1159 ) | ( x619 & n30149 ) | ( ~x1159 & n30149 ) ;
  assign n30156 = ~n30154 & n30155 ;
  assign n30157 = n30153 | n30156 ;
  assign n30158 = x789 & n30157 ;
  assign n30159 = n30150 | n30158 ;
  assign n30160 = n16176 | n30159 ;
  assign n30161 = n16176 & ~n30130 ;
  assign n30162 = n30160 & ~n30161 ;
  assign n30163 = n15134 | n30162 ;
  assign n30164 = n15134 & ~n30130 ;
  assign n30165 = n30163 & ~n30164 ;
  assign n30166 = n18610 & n30165 ;
  assign n30167 = ( x647 & x1157 ) | ( x647 & ~n30130 ) | ( x1157 & ~n30130 ) ;
  assign n30168 = x730 & n15202 ;
  assign n30169 = n30130 & ~n30168 ;
  assign n30170 = ~x778 & n30169 ;
  assign n30171 = ~x625 & n30168 ;
  assign n30172 = n30169 | n30171 ;
  assign n30173 = x1153 & n30172 ;
  assign n30174 = ~x1153 & n30130 ;
  assign n30175 = ~n30171 & n30174 ;
  assign n30176 = n30173 | n30175 ;
  assign n30177 = x778 & n30176 ;
  assign n30178 = n30170 | n30177 ;
  assign n30179 = n16043 | n30178 ;
  assign n30180 = n16045 | n30179 ;
  assign n30181 = n16047 | n30180 ;
  assign n30182 = n16049 | n30181 ;
  assign n30183 = n16055 | n30182 ;
  assign n30184 = ( x647 & ~x1157 ) | ( x647 & n30183 ) | ( ~x1157 & n30183 ) ;
  assign n30185 = ~n30167 & n30184 ;
  assign n30186 = x630 & n30185 ;
  assign n30187 = x647 & n30183 ;
  assign n30188 = ~x647 & n30130 ;
  assign n30189 = n30187 | n30188 ;
  assign n30190 = n15138 & n30189 ;
  assign n30191 = n30186 | n30190 ;
  assign n30192 = n30166 | n30191 ;
  assign n30193 = x787 & n30192 ;
  assign n30194 = n16115 & ~n30181 ;
  assign n30195 = ( x626 & ~n15419 ) | ( x626 & n30130 ) | ( ~n15419 & n30130 ) ;
  assign n30196 = ( x626 & n15419 ) | ( x626 & ~n30159 ) | ( n15419 & ~n30159 ) ;
  assign n30197 = ~n30195 & n30196 ;
  assign n30198 = n30194 | n30197 ;
  assign n30199 = ( x626 & n15418 ) | ( x626 & ~n30130 ) | ( n15418 & ~n30130 ) ;
  assign n30200 = ( x626 & ~n15418 ) | ( x626 & n30159 ) | ( ~n15418 & n30159 ) ;
  assign n30201 = n30199 & ~n30200 ;
  assign n30202 = n30198 | n30201 ;
  assign n30203 = x788 & n30202 ;
  assign n30204 = x648 & ~n30156 ;
  assign n30205 = ( x619 & x1159 ) | ( x619 & n30180 ) | ( x1159 & n30180 ) ;
  assign n30206 = x627 | n30144 ;
  assign n30207 = ( x618 & x1154 ) | ( x618 & ~n30179 ) | ( x1154 & ~n30179 ) ;
  assign n30208 = x660 | n30136 ;
  assign n30209 = ( x609 & x1155 ) | ( x609 & ~n30178 ) | ( x1155 & ~n30178 ) ;
  assign n30210 = n14839 | n30169 ;
  assign n30211 = x625 & ~n30210 ;
  assign n30212 = n30132 & n30210 ;
  assign n30213 = n30211 | n30212 ;
  assign n30214 = n30174 & n30213 ;
  assign n30215 = x608 | n30173 ;
  assign n30216 = n30214 | n30215 ;
  assign n30217 = x1153 & n30132 ;
  assign n30218 = ~n30211 & n30217 ;
  assign n30219 = x608 & ~n30175 ;
  assign n30220 = ~n30218 & n30219 ;
  assign n30221 = n30216 & ~n30220 ;
  assign n30222 = x778 & ~n30221 ;
  assign n30223 = x778 | n30212 ;
  assign n30224 = ~n30222 & n30223 ;
  assign n30225 = ( x609 & ~x1155 ) | ( x609 & n30224 ) | ( ~x1155 & n30224 ) ;
  assign n30226 = ~n30209 & n30225 ;
  assign n30227 = n30208 | n30226 ;
  assign n30228 = x660 & ~n30138 ;
  assign n30229 = ( x609 & x1155 ) | ( x609 & n30178 ) | ( x1155 & n30178 ) ;
  assign n30230 = ( ~x609 & x1155 ) | ( ~x609 & n30224 ) | ( x1155 & n30224 ) ;
  assign n30231 = n30229 & n30230 ;
  assign n30232 = n30228 & ~n30231 ;
  assign n30233 = n30227 & ~n30232 ;
  assign n30234 = x785 & ~n30233 ;
  assign n30235 = x785 | n30224 ;
  assign n30236 = ~n30234 & n30235 ;
  assign n30237 = ( x618 & ~x1154 ) | ( x618 & n30236 ) | ( ~x1154 & n30236 ) ;
  assign n30238 = ~n30207 & n30237 ;
  assign n30239 = n30206 | n30238 ;
  assign n30240 = x627 & ~n30146 ;
  assign n30241 = ( x618 & x1154 ) | ( x618 & n30179 ) | ( x1154 & n30179 ) ;
  assign n30242 = ( ~x618 & x1154 ) | ( ~x618 & n30236 ) | ( x1154 & n30236 ) ;
  assign n30243 = n30241 & n30242 ;
  assign n30244 = n30240 & ~n30243 ;
  assign n30245 = n30239 & ~n30244 ;
  assign n30246 = x781 & ~n30245 ;
  assign n30247 = x781 | n30236 ;
  assign n30248 = ~n30246 & n30247 ;
  assign n30249 = ( ~x619 & x1159 ) | ( ~x619 & n30248 ) | ( x1159 & n30248 ) ;
  assign n30250 = n30205 & n30249 ;
  assign n30251 = n30204 & ~n30250 ;
  assign n30252 = x648 | n30153 ;
  assign n30253 = ( x619 & x1159 ) | ( x619 & ~n30180 ) | ( x1159 & ~n30180 ) ;
  assign n30254 = ( x619 & ~x1159 ) | ( x619 & n30248 ) | ( ~x1159 & n30248 ) ;
  assign n30255 = ~n30253 & n30254 ;
  assign n30256 = n30252 | n30255 ;
  assign n30257 = x789 & n30256 ;
  assign n30258 = ~n30251 & n30257 ;
  assign n30259 = ~x789 & n30248 ;
  assign n30260 = n16177 | n30259 ;
  assign n30261 = n30258 | n30260 ;
  assign n30262 = ~n30203 & n30261 ;
  assign n30263 = n18434 | n30262 ;
  assign n30264 = n16650 | n30182 ;
  assign n30265 = n16051 & ~n30162 ;
  assign n30266 = n30264 & ~n30265 ;
  assign n30267 = ( x629 & ~x792 ) | ( x629 & n30266 ) | ( ~x792 & n30266 ) ;
  assign n30268 = n16052 & ~n30162 ;
  assign n30269 = n16643 & ~n30182 ;
  assign n30270 = n30268 | n30269 ;
  assign n30271 = ( x629 & x792 ) | ( x629 & n30270 ) | ( x792 & n30270 ) ;
  assign n30272 = ~n30267 & n30271 ;
  assign n30273 = n18431 | n30272 ;
  assign n30274 = n30263 & ~n30273 ;
  assign n30275 = n30193 | n30274 ;
  assign n30276 = ( x790 & x832 ) | ( x790 & n30275 ) | ( x832 & n30275 ) ;
  assign n30277 = n15141 | n30165 ;
  assign n30278 = n15141 & ~n30130 ;
  assign n30279 = n30277 & ~n30278 ;
  assign n30280 = ( x644 & x715 ) | ( x644 & ~n30279 ) | ( x715 & ~n30279 ) ;
  assign n30281 = ( x644 & ~x715 ) | ( x644 & n30130 ) | ( ~x715 & n30130 ) ;
  assign n30282 = ~n30280 & n30281 ;
  assign n30283 = x1160 & ~n30282 ;
  assign n30284 = ~x787 & n30183 ;
  assign n30285 = x1157 & n30189 ;
  assign n30286 = n30185 | n30285 ;
  assign n30287 = x787 & n30286 ;
  assign n30288 = n30284 | n30287 ;
  assign n30289 = ( x644 & x715 ) | ( x644 & n30288 ) | ( x715 & n30288 ) ;
  assign n30290 = ( ~x644 & x715 ) | ( ~x644 & n30275 ) | ( x715 & n30275 ) ;
  assign n30291 = n30289 & n30290 ;
  assign n30292 = n30283 & ~n30291 ;
  assign n30293 = ( x644 & x715 ) | ( x644 & n30279 ) | ( x715 & n30279 ) ;
  assign n30294 = ( ~x644 & x715 ) | ( ~x644 & n30130 ) | ( x715 & n30130 ) ;
  assign n30295 = n30293 & n30294 ;
  assign n30296 = x1160 | n30295 ;
  assign n30297 = ( x644 & x715 ) | ( x644 & ~n30288 ) | ( x715 & ~n30288 ) ;
  assign n30298 = ( x644 & ~x715 ) | ( x644 & n30275 ) | ( ~x715 & n30275 ) ;
  assign n30299 = ~n30297 & n30298 ;
  assign n30300 = n30296 | n30299 ;
  assign n30301 = ~n30292 & n30300 ;
  assign n30302 = ( ~x790 & x832 ) | ( ~x790 & n30301 ) | ( x832 & n30301 ) ;
  assign n30303 = n30276 & n30302 ;
  assign n30304 = n30129 | n30303 ;
  assign n30305 = n7614 & ~n14012 ;
  assign n30306 = x171 & n11725 ;
  assign n30307 = n30305 | n30306 ;
  assign n30308 = x299 & n30307 ;
  assign n30309 = ( x192 & x232 ) | ( x192 & ~n14331 ) | ( x232 & ~n14331 ) ;
  assign n30310 = ( x192 & ~x232 ) | ( x192 & n14335 ) | ( ~x232 & n14335 ) ;
  assign n30311 = n30309 & ~n30310 ;
  assign n30312 = ~n30308 & n30311 ;
  assign n30313 = n14341 & ~n30312 ;
  assign n30314 = x171 | n7301 ;
  assign n30315 = n14352 & n30314 ;
  assign n30316 = n7296 & ~n30315 ;
  assign n30317 = n7298 & ~n30316 ;
  assign n30318 = ( x192 & n14358 ) | ( x192 & n30317 ) | ( n14358 & n30317 ) ;
  assign n30319 = ( ~x192 & n14345 ) | ( ~x192 & n30317 ) | ( n14345 & n30317 ) ;
  assign n30320 = n30318 | n30319 ;
  assign n30321 = x232 & n30320 ;
  assign n30322 = n14351 | n30321 ;
  assign n30323 = x39 & n30322 ;
  assign n30324 = n1975 | n30323 ;
  assign n30325 = n30313 | n30324 ;
  assign n30326 = ~x87 & n30325 ;
  assign n30327 = n14326 | n30326 ;
  assign n30328 = ~x92 & n30327 ;
  assign n30329 = n14325 | n30328 ;
  assign n30330 = ~x55 & n30329 ;
  assign n30331 = n14373 | n30330 ;
  assign n30332 = ~n2058 & n30331 ;
  assign n30333 = x138 | n14378 ;
  assign n30334 = x196 | n30333 ;
  assign n30335 = x195 & n30334 ;
  assign n30336 = ~n8073 & n30335 ;
  assign n30337 = ~n30332 & n30336 ;
  assign n30338 = ~n14045 & n14380 ;
  assign n30339 = n8366 | n30335 ;
  assign n30340 = ( x39 & n30338 ) | ( x39 & ~n30339 ) | ( n30338 & ~n30339 ) ;
  assign n30341 = ~n4714 & n14043 ;
  assign n30342 = n9616 | n30341 ;
  assign n30343 = n9613 | n14021 ;
  assign n30344 = n14018 & ~n14385 ;
  assign n30345 = n30343 & ~n30344 ;
  assign n30346 = ~n30342 & n30345 ;
  assign n30347 = x232 & ~n30346 ;
  assign n30348 = n14383 & ~n30347 ;
  assign n30349 = ( x39 & n30339 ) | ( x39 & ~n30348 ) | ( n30339 & ~n30348 ) ;
  assign n30350 = n30340 & ~n30349 ;
  assign n30351 = n30337 | n30350 ;
  assign n30352 = x170 | n7301 ;
  assign n30353 = n14352 & n30352 ;
  assign n30354 = n7296 & ~n30353 ;
  assign n30355 = n7298 & ~n30354 ;
  assign n30356 = n14345 | n30355 ;
  assign n30357 = x232 & n30356 ;
  assign n30358 = n14351 | n30357 ;
  assign n30359 = x232 & n14358 ;
  assign n30360 = n30358 | n30359 ;
  assign n30361 = x39 & n30360 ;
  assign n30362 = ~x38 & x194 ;
  assign n30363 = ~n30361 & n30362 ;
  assign n30364 = x39 & n30358 ;
  assign n30365 = x38 | x194 ;
  assign n30366 = n30364 | n30365 ;
  assign n30367 = ~n30363 & n30366 ;
  assign n30368 = n14341 | n30367 ;
  assign n30369 = ~n14335 & n30363 ;
  assign n30370 = n14331 | n30366 ;
  assign n30371 = ~n30369 & n30370 ;
  assign n30372 = n7614 & ~n14117 ;
  assign n30373 = x170 & n11725 ;
  assign n30374 = n30372 | n30373 ;
  assign n30375 = x299 & n30374 ;
  assign n30376 = x232 & ~n30375 ;
  assign n30377 = ~n30371 & n30376 ;
  assign n30378 = n30368 & ~n30377 ;
  assign n30379 = n1924 | n30378 ;
  assign n30380 = ( ~x87 & n14326 ) | ( ~x87 & n30379 ) | ( n14326 & n30379 ) ;
  assign n30381 = ~x92 & n30380 ;
  assign n30382 = n14325 | n30381 ;
  assign n30383 = ~x55 & n30382 ;
  assign n30384 = n14373 | n30383 ;
  assign n30385 = ~n2058 & n30384 ;
  assign n30386 = n8073 | n30385 ;
  assign n30387 = ( x196 & ~n30333 ) | ( x196 & n30386 ) | ( ~n30333 & n30386 ) ;
  assign n30388 = ~x170 & n7759 ;
  assign n30389 = n14384 | n30388 ;
  assign n30390 = n11170 & n30389 ;
  assign n30391 = n11172 & n14384 ;
  assign n30392 = x232 & ~n30391 ;
  assign n30393 = ~n30390 & n30392 ;
  assign n30394 = n14383 & ~n30393 ;
  assign n30395 = ( x38 & x39 ) | ( x38 & ~n30394 ) | ( x39 & ~n30394 ) ;
  assign n30396 = ~n14172 & n14380 ;
  assign n30397 = ( ~x38 & x39 ) | ( ~x38 & n30396 ) | ( x39 & n30396 ) ;
  assign n30398 = ~n30395 & n30397 ;
  assign n30399 = ( x194 & n8359 ) | ( x194 & ~n30398 ) | ( n8359 & ~n30398 ) ;
  assign n30400 = x299 & ~n30394 ;
  assign n30401 = n9614 & ~n30400 ;
  assign n30402 = ( x38 & x39 ) | ( x38 & ~n30401 ) | ( x39 & ~n30401 ) ;
  assign n30403 = ~n14118 & n14380 ;
  assign n30404 = ( ~x38 & x39 ) | ( ~x38 & n30403 ) | ( x39 & n30403 ) ;
  assign n30405 = ~n30402 & n30404 ;
  assign n30406 = ( x194 & ~n8359 ) | ( x194 & n30405 ) | ( ~n8359 & n30405 ) ;
  assign n30407 = ~n30399 & n30406 ;
  assign n30408 = ( x196 & n30333 ) | ( x196 & n30407 ) | ( n30333 & n30407 ) ;
  assign n30409 = ~n30387 & n30408 ;
  assign n30410 = x195 & ~x196 ;
  assign n30411 = ( ~n30333 & n30407 ) | ( ~n30333 & n30410 ) | ( n30407 & n30410 ) ;
  assign n30412 = ( n30333 & n30386 ) | ( n30333 & n30410 ) | ( n30386 & n30410 ) ;
  assign n30413 = n30411 & ~n30412 ;
  assign n30414 = n30409 | n30413 ;
  assign n30415 = ~x767 & x947 ;
  assign n30416 = ~x698 & n18913 ;
  assign n30417 = n30415 | n30416 ;
  assign n30418 = ( ~x832 & n1290 ) | ( ~x832 & n30417 ) | ( n1290 & n30417 ) ;
  assign n30419 = ( x197 & x832 ) | ( x197 & n1290 ) | ( x832 & n1290 ) ;
  assign n30420 = ~n30418 & n30419 ;
  assign n30421 = x197 & ~n14827 ;
  assign n30422 = n15070 & ~n30415 ;
  assign n30423 = x38 & ~n30422 ;
  assign n30424 = ~n30421 & n30423 ;
  assign n30425 = x197 | n18988 ;
  assign n30426 = ~n19019 & n30425 ;
  assign n30427 = x767 | n30426 ;
  assign n30428 = ( x197 & ~x299 ) | ( x197 & n19161 ) | ( ~x299 & n19161 ) ;
  assign n30429 = ( x197 & x299 ) | ( x197 & n19001 ) | ( x299 & n19001 ) ;
  assign n30430 = ~n30428 & n30429 ;
  assign n30431 = n30427 | n30430 ;
  assign n30432 = ~x197 & x767 ;
  assign n30433 = ~n14710 & n30432 ;
  assign n30434 = x39 & ~n30433 ;
  assign n30435 = n30431 & n30434 ;
  assign n30436 = ( x39 & n14822 ) | ( x39 & n30415 ) | ( n14822 & n30415 ) ;
  assign n30437 = ( ~x39 & x197 ) | ( ~x39 & n14822 ) | ( x197 & n14822 ) ;
  assign n30438 = ~n30436 & n30437 ;
  assign n30439 = x38 | n30438 ;
  assign n30440 = n30435 | n30439 ;
  assign n30441 = ~n30424 & n30440 ;
  assign n30442 = x698 & ~n30441 ;
  assign n30443 = ~n19072 & n30438 ;
  assign n30444 = ~n19069 & n30425 ;
  assign n30445 = x767 & ~n30444 ;
  assign n30446 = ( x197 & ~x299 ) | ( x197 & n19066 ) | ( ~x299 & n19066 ) ;
  assign n30447 = ( x197 & x299 ) | ( x197 & n19050 ) | ( x299 & n19050 ) ;
  assign n30448 = ~n30446 & n30447 ;
  assign n30449 = n30445 & ~n30448 ;
  assign n30450 = x39 & ~n30449 ;
  assign n30451 = ( ~x197 & x767 ) | ( ~x197 & n19099 ) | ( x767 & n19099 ) ;
  assign n30452 = ( x197 & x767 ) | ( x197 & ~n19114 ) | ( x767 & ~n19114 ) ;
  assign n30453 = n30451 | n30452 ;
  assign n30454 = n30450 & n30453 ;
  assign n30455 = n30443 | n30454 ;
  assign n30456 = ~x38 & n30455 ;
  assign n30457 = x767 & x947 ;
  assign n30458 = x39 | n30457 ;
  assign n30459 = n19236 & ~n30458 ;
  assign n30460 = x197 | n15070 ;
  assign n30461 = x38 & n30460 ;
  assign n30462 = ~n30459 & n30461 ;
  assign n30463 = x698 | n30462 ;
  assign n30464 = n30456 | n30463 ;
  assign n30465 = ~n30442 & n30464 ;
  assign n30466 = ( ~x832 & n8359 ) | ( ~x832 & n30465 ) | ( n8359 & n30465 ) ;
  assign n30467 = ( ~x197 & x832 ) | ( ~x197 & n8359 ) | ( x832 & n8359 ) ;
  assign n30468 = n30466 & ~n30467 ;
  assign n30469 = n30420 | n30468 ;
  assign n30470 = n1925 | n14822 ;
  assign n30471 = ~n14828 & n30470 ;
  assign n30472 = x198 & ~n30471 ;
  assign n30473 = x198 & ~n16705 ;
  assign n30474 = n1823 | n30473 ;
  assign n30475 = ~x223 & n30474 ;
  assign n30476 = x198 & ~n14997 ;
  assign n30477 = ( ~n1823 & n4764 ) | ( ~n1823 & n30476 ) | ( n4764 & n30476 ) ;
  assign n30478 = n4712 | n30473 ;
  assign n30479 = x198 & ~n14641 ;
  assign n30480 = n4712 & ~n30479 ;
  assign n30481 = n30478 & ~n30480 ;
  assign n30482 = ( n1823 & n4764 ) | ( n1823 & ~n30481 ) | ( n4764 & ~n30481 ) ;
  assign n30483 = ~n30477 & n30482 ;
  assign n30484 = n30475 & ~n30483 ;
  assign n30485 = ( n14475 & n14484 ) | ( n14475 & n14490 ) | ( n14484 & n14490 ) ;
  assign n30486 = x198 & ~n30485 ;
  assign n30487 = n30478 & n30486 ;
  assign n30488 = ~n4708 & n14521 ;
  assign n30489 = n4708 & n14475 ;
  assign n30490 = x198 & ~n30489 ;
  assign n30491 = ~n30488 & n30490 ;
  assign n30492 = n4764 & n30491 ;
  assign n30493 = n30487 | n30492 ;
  assign n30494 = x223 & n30493 ;
  assign n30495 = x299 | n30494 ;
  assign n30496 = n30484 | n30495 ;
  assign n30497 = n2203 | n30473 ;
  assign n30498 = ~x215 & n30497 ;
  assign n30499 = ( ~n2203 & n4721 ) | ( ~n2203 & n30476 ) | ( n4721 & n30476 ) ;
  assign n30500 = ( n2203 & n4721 ) | ( n2203 & ~n30481 ) | ( n4721 & ~n30481 ) ;
  assign n30501 = ~n30499 & n30500 ;
  assign n30502 = n30498 & ~n30501 ;
  assign n30503 = n4721 & n30491 ;
  assign n30504 = n30487 | n30503 ;
  assign n30505 = x215 & n30504 ;
  assign n30506 = x299 & ~n30505 ;
  assign n30507 = ~n30502 & n30506 ;
  assign n30508 = ~n2032 & n9138 ;
  assign n30509 = ~n30507 & n30508 ;
  assign n30510 = n30496 & n30509 ;
  assign n30511 = n30472 | n30510 ;
  assign n30512 = n15134 & n30511 ;
  assign n30513 = x198 & n2032 ;
  assign n30514 = x198 & ~n14814 ;
  assign n30515 = x603 & x633 ;
  assign n30516 = n30514 | n30515 ;
  assign n30517 = ~n14941 & n14943 ;
  assign n30518 = x198 & ~n30517 ;
  assign n30519 = ~n14914 & n14918 ;
  assign n30520 = ~x198 & n30519 ;
  assign n30521 = n30518 | n30520 ;
  assign n30522 = n30515 & ~n30521 ;
  assign n30523 = n30516 & ~n30522 ;
  assign n30524 = ( x39 & x299 ) | ( x39 & n30523 ) | ( x299 & n30523 ) ;
  assign n30525 = n14783 & ~n14925 ;
  assign n30526 = n14951 | n30525 ;
  assign n30527 = x633 & n30526 ;
  assign n30528 = n14819 | n30527 ;
  assign n30529 = ~n14950 & n30528 ;
  assign n30530 = ( x39 & ~x299 ) | ( x39 & n30529 ) | ( ~x299 & n30529 ) ;
  assign n30531 = n30524 | n30530 ;
  assign n30532 = x633 & n16705 ;
  assign n30533 = ~n14838 & n30532 ;
  assign n30534 = n30473 | n30533 ;
  assign n30535 = x603 & n30534 ;
  assign n30536 = ~x603 & n30473 ;
  assign n30537 = n30535 | n30536 ;
  assign n30538 = n2203 | n30537 ;
  assign n30539 = ~x215 & n30538 ;
  assign n30540 = n14599 | n14604 ;
  assign n30541 = x198 & ~n30540 ;
  assign n30542 = x633 & n15019 ;
  assign n30543 = n30541 | n30542 ;
  assign n30544 = n4713 | n30543 ;
  assign n30545 = n4713 & ~n30534 ;
  assign n30546 = x603 & n14855 ;
  assign n30547 = ~n30545 & n30546 ;
  assign n30548 = n30544 & n30547 ;
  assign n30549 = x603 & n30543 ;
  assign n30550 = ~n14855 & n30549 ;
  assign n30551 = x198 & ~n15009 ;
  assign n30552 = n30550 | n30551 ;
  assign n30553 = n30548 | n30552 ;
  assign n30554 = n4711 | n30553 ;
  assign n30555 = n4711 & ~n30541 ;
  assign n30556 = ~n30549 & n30555 ;
  assign n30557 = n30554 & ~n30556 ;
  assign n30558 = ( ~n2203 & n4721 ) | ( ~n2203 & n30557 ) | ( n4721 & n30557 ) ;
  assign n30559 = n4707 & n30535 ;
  assign n30560 = n30536 | n30559 ;
  assign n30561 = ( x642 & n4707 ) | ( x642 & ~n30535 ) | ( n4707 & ~n30535 ) ;
  assign n30562 = ~n4713 & n30534 ;
  assign n30563 = n4713 & n30543 ;
  assign n30564 = n30562 | n30563 ;
  assign n30565 = x603 & n30564 ;
  assign n30566 = ( x642 & ~n4707 ) | ( x642 & n30565 ) | ( ~n4707 & n30565 ) ;
  assign n30567 = ~n30561 & n30566 ;
  assign n30568 = n30560 | n30567 ;
  assign n30569 = n4711 | n30568 ;
  assign n30570 = ~x603 & n30479 ;
  assign n30571 = n4711 & ~n30570 ;
  assign n30572 = ~n30565 & n30571 ;
  assign n30573 = n30569 & ~n30572 ;
  assign n30574 = ( n2203 & n4721 ) | ( n2203 & ~n30573 ) | ( n4721 & ~n30573 ) ;
  assign n30575 = ~n30558 & n30574 ;
  assign n30576 = n30539 & ~n30575 ;
  assign n30577 = n14876 & ~n14879 ;
  assign n30578 = x633 & n30577 ;
  assign n30579 = n30491 | n30578 ;
  assign n30580 = ~n4711 & n30579 ;
  assign n30581 = n14475 & n30533 ;
  assign n30582 = x198 & ~n14475 ;
  assign n30583 = n30581 | n30582 ;
  assign n30584 = n14965 & n30583 ;
  assign n30585 = n30580 | n30584 ;
  assign n30586 = ( x215 & ~n4721 ) | ( x215 & n30585 ) | ( ~n4721 & n30585 ) ;
  assign n30587 = n30486 | n30581 ;
  assign n30588 = n30562 | n30587 ;
  assign n30589 = x603 & n30588 ;
  assign n30590 = ( ~n14855 & n30536 ) | ( ~n14855 & n30589 ) | ( n30536 & n30589 ) ;
  assign n30591 = ( n14855 & n30535 ) | ( n14855 & n30536 ) | ( n30535 & n30536 ) ;
  assign n30592 = n30590 | n30591 ;
  assign n30593 = ~n4711 & n30592 ;
  assign n30594 = n30486 | n30589 ;
  assign n30595 = n4711 & n30594 ;
  assign n30596 = n30593 | n30595 ;
  assign n30597 = ( x215 & n4721 ) | ( x215 & n30596 ) | ( n4721 & n30596 ) ;
  assign n30598 = n30586 & n30597 ;
  assign n30599 = n30576 | n30598 ;
  assign n30600 = ( ~x39 & x299 ) | ( ~x39 & n30599 ) | ( x299 & n30599 ) ;
  assign n30601 = n1823 | n30537 ;
  assign n30602 = ~x223 & n30601 ;
  assign n30603 = ( ~n1823 & n4764 ) | ( ~n1823 & n30557 ) | ( n4764 & n30557 ) ;
  assign n30604 = ( n1823 & n4764 ) | ( n1823 & ~n30573 ) | ( n4764 & ~n30573 ) ;
  assign n30605 = ~n30603 & n30604 ;
  assign n30606 = n30602 & ~n30605 ;
  assign n30607 = ( x223 & ~n4764 ) | ( x223 & n30585 ) | ( ~n4764 & n30585 ) ;
  assign n30608 = ( x223 & n4764 ) | ( x223 & n30596 ) | ( n4764 & n30596 ) ;
  assign n30609 = n30607 & n30608 ;
  assign n30610 = n30606 | n30609 ;
  assign n30611 = ( x39 & x299 ) | ( x39 & ~n30610 ) | ( x299 & ~n30610 ) ;
  assign n30612 = ~n30600 & n30611 ;
  assign n30613 = n30531 & ~n30612 ;
  assign n30614 = x38 | n30613 ;
  assign n30615 = x39 & x198 ;
  assign n30616 = x38 & ~n30615 ;
  assign n30617 = x198 & ~n15756 ;
  assign n30618 = x633 & n14839 ;
  assign n30619 = n15756 & n30618 ;
  assign n30620 = n30617 | n30619 ;
  assign n30621 = ~x39 & n30620 ;
  assign n30622 = n30616 & ~n30621 ;
  assign n30623 = n2032 | n30622 ;
  assign n30624 = n30614 & ~n30623 ;
  assign n30625 = n30513 | n30624 ;
  assign n30626 = ~n15082 & n30625 ;
  assign n30627 = n15082 & n30511 ;
  assign n30628 = n30626 | n30627 ;
  assign n30629 = ~x785 & n30628 ;
  assign n30630 = ~n15088 & n30511 ;
  assign n30631 = x609 & n30626 ;
  assign n30632 = n30630 | n30631 ;
  assign n30633 = x1155 & n30632 ;
  assign n30634 = n15094 & n30511 ;
  assign n30635 = ~x609 & n30626 ;
  assign n30636 = n30634 | n30635 ;
  assign n30637 = ~x1155 & n30636 ;
  assign n30638 = n30633 | n30637 ;
  assign n30639 = x785 & n30638 ;
  assign n30640 = n30629 | n30639 ;
  assign n30641 = ~x781 & n30640 ;
  assign n30642 = ( x618 & x1154 ) | ( x618 & n30511 ) | ( x1154 & n30511 ) ;
  assign n30643 = ( ~x618 & x1154 ) | ( ~x618 & n30640 ) | ( x1154 & n30640 ) ;
  assign n30644 = n30642 & n30643 ;
  assign n30645 = ( x618 & x1154 ) | ( x618 & ~n30511 ) | ( x1154 & ~n30511 ) ;
  assign n30646 = ( x618 & ~x1154 ) | ( x618 & n30640 ) | ( ~x1154 & n30640 ) ;
  assign n30647 = ~n30645 & n30646 ;
  assign n30648 = n30644 | n30647 ;
  assign n30649 = x781 & n30648 ;
  assign n30650 = n30641 | n30649 ;
  assign n30651 = ~x789 & n30650 ;
  assign n30652 = ( x619 & x1159 ) | ( x619 & n30511 ) | ( x1159 & n30511 ) ;
  assign n30653 = ( ~x619 & x1159 ) | ( ~x619 & n30650 ) | ( x1159 & n30650 ) ;
  assign n30654 = n30652 & n30653 ;
  assign n30655 = ( x619 & x1159 ) | ( x619 & ~n30511 ) | ( x1159 & ~n30511 ) ;
  assign n30656 = ( x619 & ~x1159 ) | ( x619 & n30650 ) | ( ~x1159 & n30650 ) ;
  assign n30657 = ~n30655 & n30656 ;
  assign n30658 = n30654 | n30657 ;
  assign n30659 = x789 & n30658 ;
  assign n30660 = n30651 | n30659 ;
  assign n30661 = n16176 | n30660 ;
  assign n30662 = n16176 & ~n30511 ;
  assign n30663 = n30661 & ~n30662 ;
  assign n30664 = ~n15134 & n30663 ;
  assign n30665 = n30512 | n30664 ;
  assign n30666 = n18610 & n30665 ;
  assign n30667 = ( x647 & x1157 ) | ( x647 & ~n30511 ) | ( x1157 & ~n30511 ) ;
  assign n30668 = n17213 & ~n30511 ;
  assign n30669 = n15407 & n30511 ;
  assign n30670 = n15151 | n30473 ;
  assign n30671 = x634 & x680 ;
  assign n30672 = ( n30473 & n30670 ) | ( n30473 & n30671 ) | ( n30670 & n30671 ) ;
  assign n30673 = n1823 | n30672 ;
  assign n30674 = ~x223 & n30673 ;
  assign n30675 = x198 & ~n15285 ;
  assign n30676 = x634 & n15156 ;
  assign n30677 = n30541 | n30676 ;
  assign n30678 = n4711 & n30677 ;
  assign n30679 = n30675 | n30678 ;
  assign n30680 = x634 & n30670 ;
  assign n30681 = n30473 | n30680 ;
  assign n30682 = n4713 & ~n30681 ;
  assign n30683 = n4713 | n30677 ;
  assign n30684 = ~n30682 & n30683 ;
  assign n30685 = ( n4708 & n15160 ) | ( n4708 & n30684 ) | ( n15160 & n30684 ) ;
  assign n30686 = ( ~n4708 & n15160 ) | ( ~n4708 & n30677 ) | ( n15160 & n30677 ) ;
  assign n30687 = n30685 & n30686 ;
  assign n30688 = n30679 | n30687 ;
  assign n30689 = ( ~n1823 & n4764 ) | ( ~n1823 & n30688 ) | ( n4764 & n30688 ) ;
  assign n30690 = n4708 | n30681 ;
  assign n30691 = n15160 & n30690 ;
  assign n30692 = ~n4713 & n30681 ;
  assign n30693 = n4713 & n30677 ;
  assign n30694 = n30692 | n30693 ;
  assign n30695 = n4708 & ~n30694 ;
  assign n30696 = n30691 & ~n30695 ;
  assign n30697 = n4711 & n30694 ;
  assign n30698 = ( x680 & n4708 ) | ( x680 & ~n30479 ) | ( n4708 & ~n30479 ) ;
  assign n30699 = ( ~x680 & n4708 ) | ( ~x680 & n30473 ) | ( n4708 & n30473 ) ;
  assign n30700 = ~n30698 & n30699 ;
  assign n30701 = n30697 | n30700 ;
  assign n30702 = n30696 | n30701 ;
  assign n30703 = ( n1823 & n4764 ) | ( n1823 & ~n30702 ) | ( n4764 & ~n30702 ) ;
  assign n30704 = ~n30689 & n30703 ;
  assign n30705 = n30674 & ~n30704 ;
  assign n30706 = ~x680 & n30491 ;
  assign n30707 = x634 & n14475 ;
  assign n30708 = n15151 & n30707 ;
  assign n30709 = n30582 | n30708 ;
  assign n30710 = n4711 & n30709 ;
  assign n30711 = n30706 | n30710 ;
  assign n30712 = n4713 | n30709 ;
  assign n30713 = ~n30682 & n30712 ;
  assign n30714 = ( n4708 & n15160 ) | ( n4708 & n30713 ) | ( n15160 & n30713 ) ;
  assign n30715 = ( ~n4708 & n15160 ) | ( ~n4708 & n30709 ) | ( n15160 & n30709 ) ;
  assign n30716 = n30714 & n30715 ;
  assign n30717 = n30711 | n30716 ;
  assign n30718 = ( x223 & ~n4764 ) | ( x223 & n30717 ) | ( ~n4764 & n30717 ) ;
  assign n30719 = n4713 & n30709 ;
  assign n30720 = n30692 | n30719 ;
  assign n30721 = n4708 & ~n30720 ;
  assign n30722 = n30691 & ~n30721 ;
  assign n30723 = n30486 & n30706 ;
  assign n30724 = n4711 & n30720 ;
  assign n30725 = n30723 | n30724 ;
  assign n30726 = n30722 | n30725 ;
  assign n30727 = ( x223 & n4764 ) | ( x223 & n30726 ) | ( n4764 & n30726 ) ;
  assign n30728 = n30718 & n30727 ;
  assign n30729 = x299 | n30728 ;
  assign n30730 = n30705 | n30729 ;
  assign n30731 = n2203 | n30672 ;
  assign n30732 = ~x215 & n30731 ;
  assign n30733 = ( ~n2203 & n4721 ) | ( ~n2203 & n30688 ) | ( n4721 & n30688 ) ;
  assign n30734 = ( n2203 & n4721 ) | ( n2203 & ~n30702 ) | ( n4721 & ~n30702 ) ;
  assign n30735 = ~n30733 & n30734 ;
  assign n30736 = n30732 & ~n30735 ;
  assign n30737 = ( x215 & ~n4721 ) | ( x215 & n30717 ) | ( ~n4721 & n30717 ) ;
  assign n30738 = ( x215 & n4721 ) | ( x215 & n30726 ) | ( n4721 & n30726 ) ;
  assign n30739 = n30737 & n30738 ;
  assign n30740 = x299 & ~n30739 ;
  assign n30741 = ~n30736 & n30740 ;
  assign n30742 = n30730 & ~n30741 ;
  assign n30743 = x39 & ~n30742 ;
  assign n30744 = x198 & n15330 ;
  assign n30745 = n15350 & n30671 ;
  assign n30746 = ~n30744 & n30745 ;
  assign n30747 = n14819 | n30746 ;
  assign n30748 = ~x299 & n30747 ;
  assign n30749 = x39 | n30748 ;
  assign n30750 = ( x299 & n30514 ) | ( x299 & n30671 ) | ( n30514 & n30671 ) ;
  assign n30751 = ~x198 & n15366 ;
  assign n30752 = ~n15338 & n15340 ;
  assign n30753 = x198 & ~n30752 ;
  assign n30754 = n30751 | n30753 ;
  assign n30755 = ( x299 & ~n30671 ) | ( x299 & n30754 ) | ( ~n30671 & n30754 ) ;
  assign n30756 = n30750 & n30755 ;
  assign n30757 = n30749 | n30756 ;
  assign n30758 = ~n30743 & n30757 ;
  assign n30759 = x38 | n30758 ;
  assign n30760 = x634 & n15171 ;
  assign n30761 = n15756 & n30760 ;
  assign n30762 = n30617 | n30761 ;
  assign n30763 = ~x39 & n30762 ;
  assign n30764 = n30616 & ~n30763 ;
  assign n30765 = n2032 | n30764 ;
  assign n30766 = n30759 & ~n30765 ;
  assign n30767 = n30513 | n30766 ;
  assign n30768 = ~x778 & n30767 ;
  assign n30769 = ( x625 & x1153 ) | ( x625 & n30511 ) | ( x1153 & n30511 ) ;
  assign n30770 = ( ~x625 & x1153 ) | ( ~x625 & n30767 ) | ( x1153 & n30767 ) ;
  assign n30771 = n30769 & n30770 ;
  assign n30772 = ( x625 & x1153 ) | ( x625 & ~n30511 ) | ( x1153 & ~n30511 ) ;
  assign n30773 = ( x625 & ~x1153 ) | ( x625 & n30767 ) | ( ~x1153 & n30767 ) ;
  assign n30774 = ~n30772 & n30773 ;
  assign n30775 = n30771 | n30774 ;
  assign n30776 = x778 & n30775 ;
  assign n30777 = n30768 | n30776 ;
  assign n30778 = n15400 | n30777 ;
  assign n30779 = n15400 & ~n30511 ;
  assign n30780 = n30778 & ~n30779 ;
  assign n30781 = ~n15407 & n30780 ;
  assign n30782 = n30669 | n30781 ;
  assign n30783 = n15414 | n30782 ;
  assign n30784 = n15421 | n30783 ;
  assign n30785 = ~n30668 & n30784 ;
  assign n30786 = ~x792 & n30785 ;
  assign n30787 = x628 & ~n30785 ;
  assign n30788 = x628 | n30511 ;
  assign n30789 = ~n30787 & n30788 ;
  assign n30790 = x1156 & n30789 ;
  assign n30791 = ( x628 & x1156 ) | ( x628 & ~n30511 ) | ( x1156 & ~n30511 ) ;
  assign n30792 = ( x628 & ~x1156 ) | ( x628 & n30785 ) | ( ~x1156 & n30785 ) ;
  assign n30793 = ~n30791 & n30792 ;
  assign n30794 = n30790 | n30793 ;
  assign n30795 = x792 & n30794 ;
  assign n30796 = n30786 | n30795 ;
  assign n30797 = ( x647 & ~x1157 ) | ( x647 & n30796 ) | ( ~x1157 & n30796 ) ;
  assign n30798 = ~n30667 & n30797 ;
  assign n30799 = x630 & n30798 ;
  assign n30800 = x647 & n30796 ;
  assign n30801 = ~x647 & n30511 ;
  assign n30802 = n30800 | n30801 ;
  assign n30803 = n15138 & n30802 ;
  assign n30804 = n30799 | n30803 ;
  assign n30805 = n30666 | n30804 ;
  assign n30806 = x787 & n30805 ;
  assign n30807 = n18621 & n30663 ;
  assign n30808 = x629 & n30793 ;
  assign n30809 = n15131 & n30789 ;
  assign n30810 = n30808 | n30809 ;
  assign n30811 = n30807 | n30810 ;
  assign n30812 = x792 & n30811 ;
  assign n30813 = n15414 & ~n30511 ;
  assign n30814 = n30783 & ~n30813 ;
  assign n30815 = n16115 & ~n30814 ;
  assign n30816 = ( x626 & ~n15419 ) | ( x626 & n30511 ) | ( ~n15419 & n30511 ) ;
  assign n30817 = ( x626 & n15419 ) | ( x626 & ~n30660 ) | ( n15419 & ~n30660 ) ;
  assign n30818 = ~n30816 & n30817 ;
  assign n30819 = n30815 | n30818 ;
  assign n30820 = ( x626 & n15418 ) | ( x626 & ~n30511 ) | ( n15418 & ~n30511 ) ;
  assign n30821 = ( x626 & ~n15418 ) | ( x626 & n30660 ) | ( ~n15418 & n30660 ) ;
  assign n30822 = n30820 & ~n30821 ;
  assign n30823 = n30819 | n30822 ;
  assign n30824 = x788 & n30823 ;
  assign n30825 = x648 & ~n30657 ;
  assign n30826 = ( x619 & x1159 ) | ( x619 & n30782 ) | ( x1159 & n30782 ) ;
  assign n30827 = x627 | n30644 ;
  assign n30828 = ( x618 & x1154 ) | ( x618 & ~n30780 ) | ( x1154 & ~n30780 ) ;
  assign n30829 = x660 | n30633 ;
  assign n30830 = ( x609 & x1155 ) | ( x609 & ~n30777 ) | ( x1155 & ~n30777 ) ;
  assign n30831 = x608 | n30771 ;
  assign n30832 = ( x625 & x1153 ) | ( x625 & ~n30625 ) | ( x1153 & ~n30625 ) ;
  assign n30833 = ~x634 & n14819 ;
  assign n30834 = x634 & n15331 ;
  assign n30835 = ~n14913 & n30834 ;
  assign n30836 = n30833 | n30835 ;
  assign n30837 = ~x633 & n30836 ;
  assign n30838 = x198 & ~x633 ;
  assign n30839 = x634 & ~x665 ;
  assign n30840 = ~n30838 & n30839 ;
  assign n30841 = ( x603 & n15877 ) | ( x603 & ~n30840 ) | ( n15877 & ~n30840 ) ;
  assign n30842 = ~n30527 & n30841 ;
  assign n30843 = ~n30837 & n30842 ;
  assign n30844 = x603 | n30747 ;
  assign n30845 = x680 & n30844 ;
  assign n30846 = ~n30843 & n30845 ;
  assign n30847 = ~x680 & n30529 ;
  assign n30848 = x299 | n30847 ;
  assign n30849 = n30846 | n30848 ;
  assign n30850 = ~x603 & n30754 ;
  assign n30851 = x198 & ~x665 ;
  assign n30852 = x633 & ~n30851 ;
  assign n30853 = ~n30751 & n30852 ;
  assign n30854 = ~n30521 & n30853 ;
  assign n30855 = ~n30519 & n30753 ;
  assign n30856 = ~n15332 & n30517 ;
  assign n30857 = n30855 | n30856 ;
  assign n30858 = ( x603 & n30515 ) | ( x603 & n30857 ) | ( n30515 & n30857 ) ;
  assign n30859 = ~n30854 & n30858 ;
  assign n30860 = n30850 | n30859 ;
  assign n30861 = ( ~x299 & n30671 ) | ( ~x299 & n30860 ) | ( n30671 & n30860 ) ;
  assign n30862 = ( x299 & ~n30523 ) | ( x299 & n30671 ) | ( ~n30523 & n30671 ) ;
  assign n30863 = ~n30861 & n30862 ;
  assign n30864 = n30849 & ~n30863 ;
  assign n30865 = x39 | n30864 ;
  assign n30866 = ~x603 & n30684 ;
  assign n30867 = ~n14481 & n14971 ;
  assign n30868 = n30839 & n30867 ;
  assign n30869 = n30534 | n30868 ;
  assign n30870 = x603 & n30869 ;
  assign n30871 = n14855 & n30870 ;
  assign n30872 = n30547 | n30871 ;
  assign n30873 = n4708 | n30872 ;
  assign n30874 = ( n14595 & n15505 ) | ( n14595 & n15507 ) | ( n15505 & n15507 ) ;
  assign n30875 = x634 & n30874 ;
  assign n30876 = n30543 | n30875 ;
  assign n30877 = n4713 & n30872 ;
  assign n30878 = n30876 | n30877 ;
  assign n30879 = n30873 & n30878 ;
  assign n30880 = n30866 | n30879 ;
  assign n30881 = n15160 & n30880 ;
  assign n30882 = ~x680 & n30553 ;
  assign n30883 = ~n14839 & n30677 ;
  assign n30884 = n30549 | n30883 ;
  assign n30885 = n4711 & n30884 ;
  assign n30886 = n30882 | n30885 ;
  assign n30887 = n30881 | n30886 ;
  assign n30888 = ( ~n2203 & n4721 ) | ( ~n2203 & n30887 ) | ( n4721 & n30887 ) ;
  assign n30889 = x680 | n30568 ;
  assign n30890 = ~n4713 & n30869 ;
  assign n30891 = n4713 & n30876 ;
  assign n30892 = n30890 | n30891 ;
  assign n30893 = x603 & n30892 ;
  assign n30894 = ~x603 & n30694 ;
  assign n30895 = n14553 | n30894 ;
  assign n30896 = n30893 | n30895 ;
  assign n30897 = ~x603 & n30681 ;
  assign n30898 = ( x642 & n30870 ) | ( x642 & n30897 ) | ( n30870 & n30897 ) ;
  assign n30899 = ( ~x642 & n30893 ) | ( ~x642 & n30897 ) | ( n30893 & n30897 ) ;
  assign n30900 = n30898 | n30899 ;
  assign n30901 = ( n4707 & n14553 ) | ( n4707 & ~n30900 ) | ( n14553 & ~n30900 ) ;
  assign n30902 = n30870 | n30897 ;
  assign n30903 = ( n4707 & ~n14553 ) | ( n4707 & n30902 ) | ( ~n14553 & n30902 ) ;
  assign n30904 = n30901 & ~n30903 ;
  assign n30905 = n30896 & ~n30904 ;
  assign n30906 = x680 & ~n30905 ;
  assign n30907 = n30889 & ~n30906 ;
  assign n30908 = ( n2203 & n4721 ) | ( n2203 & ~n30907 ) | ( n4721 & ~n30907 ) ;
  assign n30909 = ~n30888 & n30908 ;
  assign n30910 = n15477 & n30680 ;
  assign n30911 = n30537 | n30910 ;
  assign n30912 = ( ~x215 & n14841 ) | ( ~x215 & n30911 ) | ( n14841 & n30911 ) ;
  assign n30913 = ~n30909 & n30912 ;
  assign n30914 = ~x603 & n30713 ;
  assign n30915 = n30877 | n30914 ;
  assign n30916 = x621 & n14465 ;
  assign n30917 = ~n15332 & n30916 ;
  assign n30918 = n14838 & n30851 ;
  assign n30919 = n30582 | n30918 ;
  assign n30920 = n30917 | n30919 ;
  assign n30921 = ( x634 & n30581 ) | ( x634 & n30920 ) | ( n30581 & n30920 ) ;
  assign n30922 = ( ~x634 & n30581 ) | ( ~x634 & n30582 ) | ( n30581 & n30582 ) ;
  assign n30923 = n30921 | n30922 ;
  assign n30924 = x603 & n30923 ;
  assign n30925 = ~n14855 & n30924 ;
  assign n30926 = n30872 & n30923 ;
  assign n30927 = n30925 | n30926 ;
  assign n30928 = n30915 | n30927 ;
  assign n30929 = n15160 & n30928 ;
  assign n30930 = ~x680 & n30579 ;
  assign n30931 = ~x603 & n30709 ;
  assign n30932 = n30924 | n30931 ;
  assign n30933 = n4711 & n30932 ;
  assign n30934 = n30930 | n30933 ;
  assign n30935 = n30929 | n30934 ;
  assign n30936 = ( x215 & ~n4721 ) | ( x215 & n30935 ) | ( ~n4721 & n30935 ) ;
  assign n30937 = n4713 & n30923 ;
  assign n30938 = n30890 | n30937 ;
  assign n30939 = x603 & n30938 ;
  assign n30940 = n14855 | n30897 ;
  assign n30941 = n30939 | n30940 ;
  assign n30942 = n14855 & ~n30902 ;
  assign n30943 = n15160 & ~n30942 ;
  assign n30944 = n30941 & n30943 ;
  assign n30945 = ~x680 & n30592 ;
  assign n30946 = ~x603 & n30720 ;
  assign n30947 = n30939 | n30946 ;
  assign n30948 = n4711 & n30947 ;
  assign n30949 = n30945 | n30948 ;
  assign n30950 = n30944 | n30949 ;
  assign n30951 = ( x215 & n4721 ) | ( x215 & n30950 ) | ( n4721 & n30950 ) ;
  assign n30952 = n30936 & n30951 ;
  assign n30953 = n30913 | n30952 ;
  assign n30954 = ( ~x39 & x299 ) | ( ~x39 & n30953 ) | ( x299 & n30953 ) ;
  assign n30955 = n1823 | n30911 ;
  assign n30956 = ~x223 & n30955 ;
  assign n30957 = ( ~n1823 & n4764 ) | ( ~n1823 & n30887 ) | ( n4764 & n30887 ) ;
  assign n30958 = ( n1823 & n4764 ) | ( n1823 & ~n30907 ) | ( n4764 & ~n30907 ) ;
  assign n30959 = ~n30957 & n30958 ;
  assign n30960 = n30956 & ~n30959 ;
  assign n30961 = ( x223 & ~n4764 ) | ( x223 & n30935 ) | ( ~n4764 & n30935 ) ;
  assign n30962 = ( x223 & n4764 ) | ( x223 & n30950 ) | ( n4764 & n30950 ) ;
  assign n30963 = n30961 & n30962 ;
  assign n30964 = n30960 | n30963 ;
  assign n30965 = ( x39 & x299 ) | ( x39 & ~n30964 ) | ( x299 & ~n30964 ) ;
  assign n30966 = ~n30954 & n30965 ;
  assign n30967 = n30865 & ~n30966 ;
  assign n30968 = x38 | n30967 ;
  assign n30969 = x634 & n15913 ;
  assign n30970 = n30620 | n30969 ;
  assign n30971 = ~x39 & n30970 ;
  assign n30972 = n30616 & ~n30971 ;
  assign n30973 = n2032 | n30972 ;
  assign n30974 = n30968 & ~n30973 ;
  assign n30975 = n30513 | n30974 ;
  assign n30976 = ( x625 & ~x1153 ) | ( x625 & n30975 ) | ( ~x1153 & n30975 ) ;
  assign n30977 = ~n30832 & n30976 ;
  assign n30978 = n30831 | n30977 ;
  assign n30979 = x608 & ~n30774 ;
  assign n30980 = ( x625 & x1153 ) | ( x625 & n30625 ) | ( x1153 & n30625 ) ;
  assign n30981 = ( ~x625 & x1153 ) | ( ~x625 & n30975 ) | ( x1153 & n30975 ) ;
  assign n30982 = n30980 & n30981 ;
  assign n30983 = n30979 & ~n30982 ;
  assign n30984 = n30978 & ~n30983 ;
  assign n30985 = x778 & ~n30984 ;
  assign n30986 = x778 | n30975 ;
  assign n30987 = ~n30985 & n30986 ;
  assign n30988 = ( x609 & ~x1155 ) | ( x609 & n30987 ) | ( ~x1155 & n30987 ) ;
  assign n30989 = ~n30830 & n30988 ;
  assign n30990 = n30829 | n30989 ;
  assign n30991 = x660 & ~n30637 ;
  assign n30992 = ( x609 & x1155 ) | ( x609 & n30777 ) | ( x1155 & n30777 ) ;
  assign n30993 = ( ~x609 & x1155 ) | ( ~x609 & n30987 ) | ( x1155 & n30987 ) ;
  assign n30994 = n30992 & n30993 ;
  assign n30995 = n30991 & ~n30994 ;
  assign n30996 = n30990 & ~n30995 ;
  assign n30997 = x785 & ~n30996 ;
  assign n30998 = x785 | n30987 ;
  assign n30999 = ~n30997 & n30998 ;
  assign n31000 = ( x618 & ~x1154 ) | ( x618 & n30999 ) | ( ~x1154 & n30999 ) ;
  assign n31001 = ~n30828 & n31000 ;
  assign n31002 = n30827 | n31001 ;
  assign n31003 = x627 & ~n30647 ;
  assign n31004 = ( x618 & x1154 ) | ( x618 & n30780 ) | ( x1154 & n30780 ) ;
  assign n31005 = ( ~x618 & x1154 ) | ( ~x618 & n30999 ) | ( x1154 & n30999 ) ;
  assign n31006 = n31004 & n31005 ;
  assign n31007 = n31003 & ~n31006 ;
  assign n31008 = n31002 & ~n31007 ;
  assign n31009 = x781 & ~n31008 ;
  assign n31010 = x781 | n30999 ;
  assign n31011 = ~n31009 & n31010 ;
  assign n31012 = ( ~x619 & x1159 ) | ( ~x619 & n31011 ) | ( x1159 & n31011 ) ;
  assign n31013 = n30826 & n31012 ;
  assign n31014 = n30825 & ~n31013 ;
  assign n31015 = x648 | n30654 ;
  assign n31016 = ( x619 & x1159 ) | ( x619 & ~n30782 ) | ( x1159 & ~n30782 ) ;
  assign n31017 = ( x619 & ~x1159 ) | ( x619 & n31011 ) | ( ~x1159 & n31011 ) ;
  assign n31018 = ~n31016 & n31017 ;
  assign n31019 = n31015 | n31018 ;
  assign n31020 = x789 & n31019 ;
  assign n31021 = ~n31014 & n31020 ;
  assign n31022 = ~x789 & n31011 ;
  assign n31023 = n16177 | n31022 ;
  assign n31024 = n31021 | n31023 ;
  assign n31025 = ~n30824 & n31024 ;
  assign n31026 = n30812 | n31025 ;
  assign n31027 = ( n18431 & n22573 ) | ( n18431 & ~n30811 ) | ( n22573 & ~n30811 ) ;
  assign n31028 = n31026 & ~n31027 ;
  assign n31029 = n30806 | n31028 ;
  assign n31030 = ~x790 & n31029 ;
  assign n31031 = n15141 | n30665 ;
  assign n31032 = n15141 & ~n30511 ;
  assign n31033 = n31031 & ~n31032 ;
  assign n31034 = ( x644 & x715 ) | ( x644 & n31033 ) | ( x715 & n31033 ) ;
  assign n31035 = ( ~x644 & x715 ) | ( ~x644 & n30511 ) | ( x715 & n30511 ) ;
  assign n31036 = n31034 & n31035 ;
  assign n31037 = x1160 | n31036 ;
  assign n31038 = ~x787 & n30796 ;
  assign n31039 = x1157 & n30802 ;
  assign n31040 = n30798 | n31039 ;
  assign n31041 = x787 & n31040 ;
  assign n31042 = n31038 | n31041 ;
  assign n31043 = ( x644 & x715 ) | ( x644 & ~n31042 ) | ( x715 & ~n31042 ) ;
  assign n31044 = ( x644 & ~x715 ) | ( x644 & n31029 ) | ( ~x715 & n31029 ) ;
  assign n31045 = ~n31043 & n31044 ;
  assign n31046 = n31037 | n31045 ;
  assign n31047 = ( x644 & x715 ) | ( x644 & ~n31033 ) | ( x715 & ~n31033 ) ;
  assign n31048 = ( x644 & ~x715 ) | ( x644 & n30511 ) | ( ~x715 & n30511 ) ;
  assign n31049 = ~n31047 & n31048 ;
  assign n31050 = x1160 & ~n31049 ;
  assign n31051 = ( x644 & x715 ) | ( x644 & n31042 ) | ( x715 & n31042 ) ;
  assign n31052 = ( ~x644 & x715 ) | ( ~x644 & n31029 ) | ( x715 & n31029 ) ;
  assign n31053 = n31051 & n31052 ;
  assign n31054 = n31050 & ~n31053 ;
  assign n31055 = x790 & ~n31054 ;
  assign n31056 = n31046 & n31055 ;
  assign n31057 = n31030 | n31056 ;
  assign n31058 = ~n6785 & n31057 ;
  assign n31059 = x198 & n6785 ;
  assign n31060 = n31058 | n31059 ;
  assign n31061 = x199 & ~n14834 ;
  assign n31062 = ( x647 & x1157 ) | ( x647 & n31061 ) | ( x1157 & n31061 ) ;
  assign n31063 = n15414 & ~n31061 ;
  assign n31064 = n15400 & ~n31061 ;
  assign n31065 = x637 | n31061 ;
  assign n31066 = x199 | n15070 ;
  assign n31067 = n17892 & n31066 ;
  assign n31068 = ( x39 & ~x199 ) | ( x39 & n15369 ) | ( ~x199 & n15369 ) ;
  assign n31069 = ( x39 & x199 ) | ( x39 & ~n15345 ) | ( x199 & ~n15345 ) ;
  assign n31070 = n31068 | n31069 ;
  assign n31071 = ~x38 & n31070 ;
  assign n31072 = ( x39 & x199 ) | ( x39 & ~n15221 ) | ( x199 & ~n15221 ) ;
  assign n31073 = ( x39 & ~x199 ) | ( x39 & n15324 ) | ( ~x199 & n15324 ) ;
  assign n31074 = n31072 & n31073 ;
  assign n31075 = n31071 & ~n31074 ;
  assign n31076 = n31067 | n31075 ;
  assign n31077 = ~n2032 & n31076 ;
  assign n31078 = x199 & n2032 ;
  assign n31079 = x637 & ~n31078 ;
  assign n31080 = ~n31077 & n31079 ;
  assign n31081 = n31065 & ~n31080 ;
  assign n31082 = ~x778 & n31081 ;
  assign n31083 = ( x625 & x1153 ) | ( x625 & n31061 ) | ( x1153 & n31061 ) ;
  assign n31084 = ( ~x625 & x1153 ) | ( ~x625 & n31081 ) | ( x1153 & n31081 ) ;
  assign n31085 = n31083 & n31084 ;
  assign n31086 = ( x625 & x1153 ) | ( x625 & ~n31061 ) | ( x1153 & ~n31061 ) ;
  assign n31087 = ( x625 & ~x1153 ) | ( x625 & n31081 ) | ( ~x1153 & n31081 ) ;
  assign n31088 = ~n31086 & n31087 ;
  assign n31089 = n31085 | n31088 ;
  assign n31090 = x778 & n31089 ;
  assign n31091 = n31082 | n31090 ;
  assign n31092 = n15400 | n31091 ;
  assign n31093 = ~n31064 & n31092 ;
  assign n31094 = ~n15407 & n31093 ;
  assign n31095 = n15407 & n31061 ;
  assign n31096 = n31094 | n31095 ;
  assign n31097 = n15414 | n31096 ;
  assign n31098 = ~n31063 & n31097 ;
  assign n31099 = ~n15421 & n31098 ;
  assign n31100 = n15421 & n31061 ;
  assign n31101 = n31099 | n31100 ;
  assign n31102 = ~x792 & n31101 ;
  assign n31103 = ( x628 & x1156 ) | ( x628 & n31061 ) | ( x1156 & n31061 ) ;
  assign n31104 = ( ~x628 & x1156 ) | ( ~x628 & n31101 ) | ( x1156 & n31101 ) ;
  assign n31105 = n31103 & n31104 ;
  assign n31106 = ( x628 & x1156 ) | ( x628 & ~n31061 ) | ( x1156 & ~n31061 ) ;
  assign n31107 = ( x628 & ~x1156 ) | ( x628 & n31101 ) | ( ~x1156 & n31101 ) ;
  assign n31108 = ~n31106 & n31107 ;
  assign n31109 = n31105 | n31108 ;
  assign n31110 = x792 & n31109 ;
  assign n31111 = n31102 | n31110 ;
  assign n31112 = ( ~x647 & x1157 ) | ( ~x647 & n31111 ) | ( x1157 & n31111 ) ;
  assign n31113 = n31062 & n31112 ;
  assign n31114 = x630 | n31113 ;
  assign n31115 = x617 | n31061 ;
  assign n31116 = x199 | n17414 ;
  assign n31117 = n17420 & n31116 ;
  assign n31118 = ( ~x38 & x199 ) | ( ~x38 & n14933 ) | ( x199 & n14933 ) ;
  assign n31119 = ( x38 & x199 ) | ( x38 & n15063 ) | ( x199 & n15063 ) ;
  assign n31120 = n31118 & ~n31119 ;
  assign n31121 = n31117 | n31120 ;
  assign n31122 = ~n2032 & n31121 ;
  assign n31123 = x617 & ~n31078 ;
  assign n31124 = ~n31122 & n31123 ;
  assign n31125 = n31115 & ~n31124 ;
  assign n31126 = n15082 | n31125 ;
  assign n31127 = n15082 & ~n31061 ;
  assign n31128 = n31126 & ~n31127 ;
  assign n31129 = ~x785 & n31128 ;
  assign n31130 = ( x609 & x1155 ) | ( x609 & n31061 ) | ( x1155 & n31061 ) ;
  assign n31131 = ( ~x609 & x1155 ) | ( ~x609 & n31128 ) | ( x1155 & n31128 ) ;
  assign n31132 = n31130 & n31131 ;
  assign n31133 = ( x609 & x1155 ) | ( x609 & ~n31061 ) | ( x1155 & ~n31061 ) ;
  assign n31134 = ( x609 & ~x1155 ) | ( x609 & n31128 ) | ( ~x1155 & n31128 ) ;
  assign n31135 = ~n31133 & n31134 ;
  assign n31136 = n31132 | n31135 ;
  assign n31137 = x785 & n31136 ;
  assign n31138 = n31129 | n31137 ;
  assign n31139 = ~x781 & n31138 ;
  assign n31140 = ( x618 & x1154 ) | ( x618 & n31061 ) | ( x1154 & n31061 ) ;
  assign n31141 = ( ~x618 & x1154 ) | ( ~x618 & n31138 ) | ( x1154 & n31138 ) ;
  assign n31142 = n31140 & n31141 ;
  assign n31143 = ( x618 & x1154 ) | ( x618 & ~n31061 ) | ( x1154 & ~n31061 ) ;
  assign n31144 = ( x618 & ~x1154 ) | ( x618 & n31138 ) | ( ~x1154 & n31138 ) ;
  assign n31145 = ~n31143 & n31144 ;
  assign n31146 = n31142 | n31145 ;
  assign n31147 = x781 & n31146 ;
  assign n31148 = n31139 | n31147 ;
  assign n31149 = ~x789 & n31148 ;
  assign n31150 = ( x619 & x1159 ) | ( x619 & n31061 ) | ( x1159 & n31061 ) ;
  assign n31151 = ( ~x619 & x1159 ) | ( ~x619 & n31148 ) | ( x1159 & n31148 ) ;
  assign n31152 = n31150 & n31151 ;
  assign n31153 = ( x619 & x1159 ) | ( x619 & ~n31061 ) | ( x1159 & ~n31061 ) ;
  assign n31154 = ( x619 & ~x1159 ) | ( x619 & n31148 ) | ( ~x1159 & n31148 ) ;
  assign n31155 = ~n31153 & n31154 ;
  assign n31156 = n31152 | n31155 ;
  assign n31157 = x789 & n31156 ;
  assign n31158 = n31149 | n31157 ;
  assign n31159 = ~n16176 & n31158 ;
  assign n31160 = n16176 & n31061 ;
  assign n31161 = n31159 | n31160 ;
  assign n31162 = ~n15134 & n31161 ;
  assign n31163 = n15134 & n31061 ;
  assign n31164 = n31162 | n31163 ;
  assign n31165 = ( x647 & x1157 ) | ( x647 & ~n31164 ) | ( x1157 & ~n31164 ) ;
  assign n31166 = x629 | n31105 ;
  assign n31167 = ( x628 & x1156 ) | ( x628 & ~n31161 ) | ( x1156 & ~n31161 ) ;
  assign n31168 = x648 | n31152 ;
  assign n31169 = ( x619 & x1159 ) | ( x619 & ~n31096 ) | ( x1159 & ~n31096 ) ;
  assign n31170 = x627 | n31142 ;
  assign n31171 = ( x618 & x1154 ) | ( x618 & ~n31093 ) | ( x1154 & ~n31093 ) ;
  assign n31172 = x660 | n31132 ;
  assign n31173 = ( x609 & x1155 ) | ( x609 & ~n31091 ) | ( x1155 & ~n31091 ) ;
  assign n31174 = x608 | n31085 ;
  assign n31175 = ( x625 & x1153 ) | ( x625 & ~n31125 ) | ( x1153 & ~n31125 ) ;
  assign n31176 = ~x637 & n31125 ;
  assign n31177 = ( x199 & ~x617 ) | ( x199 & n17554 ) | ( ~x617 & n17554 ) ;
  assign n31178 = ~n2032 & n17562 ;
  assign n31179 = ( x199 & x617 ) | ( x199 & n31178 ) | ( x617 & n31178 ) ;
  assign n31180 = ~n31177 & n31179 ;
  assign n31181 = n31078 | n31180 ;
  assign n31182 = ~n2032 & n22514 ;
  assign n31183 = x617 | n17574 ;
  assign n31184 = ( x199 & n31182 ) | ( x199 & ~n31183 ) | ( n31182 & ~n31183 ) ;
  assign n31185 = ( x199 & n17578 ) | ( x199 & n31183 ) | ( n17578 & n31183 ) ;
  assign n31186 = n31184 & ~n31185 ;
  assign n31187 = n31181 | n31186 ;
  assign n31188 = x637 & n31187 ;
  assign n31189 = n31176 | n31188 ;
  assign n31190 = ( x625 & ~x1153 ) | ( x625 & n31189 ) | ( ~x1153 & n31189 ) ;
  assign n31191 = ~n31175 & n31190 ;
  assign n31192 = n31174 | n31191 ;
  assign n31193 = x608 & ~n31088 ;
  assign n31194 = ( x625 & x1153 ) | ( x625 & n31125 ) | ( x1153 & n31125 ) ;
  assign n31195 = ( ~x625 & x1153 ) | ( ~x625 & n31189 ) | ( x1153 & n31189 ) ;
  assign n31196 = n31194 & n31195 ;
  assign n31197 = n31193 & ~n31196 ;
  assign n31198 = n31192 & ~n31197 ;
  assign n31199 = x778 & ~n31198 ;
  assign n31200 = x778 | n31189 ;
  assign n31201 = ~n31199 & n31200 ;
  assign n31202 = ( x609 & ~x1155 ) | ( x609 & n31201 ) | ( ~x1155 & n31201 ) ;
  assign n31203 = ~n31173 & n31202 ;
  assign n31204 = n31172 | n31203 ;
  assign n31205 = x660 & ~n31135 ;
  assign n31206 = ( x609 & x1155 ) | ( x609 & n31091 ) | ( x1155 & n31091 ) ;
  assign n31207 = ( ~x609 & x1155 ) | ( ~x609 & n31201 ) | ( x1155 & n31201 ) ;
  assign n31208 = n31206 & n31207 ;
  assign n31209 = n31205 & ~n31208 ;
  assign n31210 = n31204 & ~n31209 ;
  assign n31211 = x785 & ~n31210 ;
  assign n31212 = x785 | n31201 ;
  assign n31213 = ~n31211 & n31212 ;
  assign n31214 = ( x618 & ~x1154 ) | ( x618 & n31213 ) | ( ~x1154 & n31213 ) ;
  assign n31215 = ~n31171 & n31214 ;
  assign n31216 = n31170 | n31215 ;
  assign n31217 = x627 & ~n31145 ;
  assign n31218 = ( x618 & x1154 ) | ( x618 & n31093 ) | ( x1154 & n31093 ) ;
  assign n31219 = ( ~x618 & x1154 ) | ( ~x618 & n31213 ) | ( x1154 & n31213 ) ;
  assign n31220 = n31218 & n31219 ;
  assign n31221 = n31217 & ~n31220 ;
  assign n31222 = n31216 & ~n31221 ;
  assign n31223 = x781 & ~n31222 ;
  assign n31224 = x781 | n31213 ;
  assign n31225 = ~n31223 & n31224 ;
  assign n31226 = ( x619 & ~x1159 ) | ( x619 & n31225 ) | ( ~x1159 & n31225 ) ;
  assign n31227 = ~n31169 & n31226 ;
  assign n31228 = n31168 | n31227 ;
  assign n31229 = x648 & ~n31155 ;
  assign n31230 = ( x619 & x1159 ) | ( x619 & n31096 ) | ( x1159 & n31096 ) ;
  assign n31231 = ( ~x619 & x1159 ) | ( ~x619 & n31225 ) | ( x1159 & n31225 ) ;
  assign n31232 = n31230 & n31231 ;
  assign n31233 = n31229 & ~n31232 ;
  assign n31234 = n31228 & ~n31233 ;
  assign n31235 = x789 & ~n31234 ;
  assign n31236 = x789 | n31225 ;
  assign n31237 = ~n31235 & n31236 ;
  assign n31238 = ~x788 & n31237 ;
  assign n31239 = ( x626 & x641 ) | ( x626 & ~n31158 ) | ( x641 & ~n31158 ) ;
  assign n31240 = ( x626 & ~x641 ) | ( x626 & n31061 ) | ( ~x641 & n31061 ) ;
  assign n31241 = n31239 & ~n31240 ;
  assign n31242 = x1158 | n31241 ;
  assign n31243 = ( x626 & x641 ) | ( x626 & n31098 ) | ( x641 & n31098 ) ;
  assign n31244 = ( ~x626 & x641 ) | ( ~x626 & n31237 ) | ( x641 & n31237 ) ;
  assign n31245 = n31243 | n31244 ;
  assign n31246 = ~n31242 & n31245 ;
  assign n31247 = ( x626 & x641 ) | ( x626 & n31158 ) | ( x641 & n31158 ) ;
  assign n31248 = ( ~x626 & x641 ) | ( ~x626 & n31061 ) | ( x641 & n31061 ) ;
  assign n31249 = n31247 | n31248 ;
  assign n31250 = x1158 & n31249 ;
  assign n31251 = ( x626 & x641 ) | ( x626 & ~n31098 ) | ( x641 & ~n31098 ) ;
  assign n31252 = ( x626 & ~x641 ) | ( x626 & n31237 ) | ( ~x641 & n31237 ) ;
  assign n31253 = n31251 & ~n31252 ;
  assign n31254 = n31250 & ~n31253 ;
  assign n31255 = n31246 | n31254 ;
  assign n31256 = x788 & n31255 ;
  assign n31257 = n31238 | n31256 ;
  assign n31258 = ( x628 & ~x1156 ) | ( x628 & n31257 ) | ( ~x1156 & n31257 ) ;
  assign n31259 = ~n31167 & n31258 ;
  assign n31260 = n31166 | n31259 ;
  assign n31261 = x629 & ~n31108 ;
  assign n31262 = ( x628 & x1156 ) | ( x628 & n31161 ) | ( x1156 & n31161 ) ;
  assign n31263 = ( ~x628 & x1156 ) | ( ~x628 & n31257 ) | ( x1156 & n31257 ) ;
  assign n31264 = n31262 & n31263 ;
  assign n31265 = n31261 & ~n31264 ;
  assign n31266 = n31260 & ~n31265 ;
  assign n31267 = x792 & ~n31266 ;
  assign n31268 = x792 | n31257 ;
  assign n31269 = ~n31267 & n31268 ;
  assign n31270 = ( x647 & ~x1157 ) | ( x647 & n31269 ) | ( ~x1157 & n31269 ) ;
  assign n31271 = ~n31165 & n31270 ;
  assign n31272 = n31114 | n31271 ;
  assign n31273 = ( x647 & x1157 ) | ( x647 & ~n31061 ) | ( x1157 & ~n31061 ) ;
  assign n31274 = ( x647 & ~x1157 ) | ( x647 & n31111 ) | ( ~x1157 & n31111 ) ;
  assign n31275 = ~n31273 & n31274 ;
  assign n31276 = x630 & ~n31275 ;
  assign n31277 = ( x647 & x1157 ) | ( x647 & n31164 ) | ( x1157 & n31164 ) ;
  assign n31278 = ( ~x647 & x1157 ) | ( ~x647 & n31269 ) | ( x1157 & n31269 ) ;
  assign n31279 = n31277 & n31278 ;
  assign n31280 = n31276 & ~n31279 ;
  assign n31281 = n31272 & ~n31280 ;
  assign n31282 = x787 & ~n31281 ;
  assign n31283 = x787 | n31269 ;
  assign n31284 = ~n31282 & n31283 ;
  assign n31285 = ~x790 & n31284 ;
  assign n31286 = n15141 & ~n31061 ;
  assign n31287 = n15141 | n31164 ;
  assign n31288 = ~n31286 & n31287 ;
  assign n31289 = ( x644 & x715 ) | ( x644 & n31288 ) | ( x715 & n31288 ) ;
  assign n31290 = ( ~x644 & x715 ) | ( ~x644 & n31061 ) | ( x715 & n31061 ) ;
  assign n31291 = n31289 & n31290 ;
  assign n31292 = x1160 | n31291 ;
  assign n31293 = ~x787 & n31111 ;
  assign n31294 = n31113 | n31275 ;
  assign n31295 = x787 & n31294 ;
  assign n31296 = n31293 | n31295 ;
  assign n31297 = ( x644 & x715 ) | ( x644 & ~n31296 ) | ( x715 & ~n31296 ) ;
  assign n31298 = ( x644 & ~x715 ) | ( x644 & n31284 ) | ( ~x715 & n31284 ) ;
  assign n31299 = ~n31297 & n31298 ;
  assign n31300 = n31292 | n31299 ;
  assign n31301 = ( x644 & x715 ) | ( x644 & ~n31288 ) | ( x715 & ~n31288 ) ;
  assign n31302 = ( x644 & ~x715 ) | ( x644 & n31061 ) | ( ~x715 & n31061 ) ;
  assign n31303 = ~n31301 & n31302 ;
  assign n31304 = x1160 & ~n31303 ;
  assign n31305 = ( x644 & x715 ) | ( x644 & n31296 ) | ( x715 & n31296 ) ;
  assign n31306 = ( ~x644 & x715 ) | ( ~x644 & n31284 ) | ( x715 & n31284 ) ;
  assign n31307 = n31305 & n31306 ;
  assign n31308 = n31304 & ~n31307 ;
  assign n31309 = x790 & ~n31308 ;
  assign n31310 = n31300 & n31309 ;
  assign n31311 = n31285 | n31310 ;
  assign n31312 = ~n6785 & n31311 ;
  assign n31313 = x199 & n6785 ;
  assign n31314 = n31312 | n31313 ;
  assign n31315 = ~x200 & n6785 ;
  assign n31316 = x200 & ~n14834 ;
  assign n31317 = x606 | n31316 ;
  assign n31318 = x200 | n17414 ;
  assign n31319 = n17420 & n31318 ;
  assign n31320 = ( ~x38 & x200 ) | ( ~x38 & n14933 ) | ( x200 & n14933 ) ;
  assign n31321 = ( x38 & x200 ) | ( x38 & n15063 ) | ( x200 & n15063 ) ;
  assign n31322 = n31320 & ~n31321 ;
  assign n31323 = n31319 | n31322 ;
  assign n31324 = ~n2032 & n31323 ;
  assign n31325 = x200 & n2032 ;
  assign n31326 = x606 & ~n31325 ;
  assign n31327 = ~n31324 & n31326 ;
  assign n31328 = n31317 & ~n31327 ;
  assign n31329 = n15082 | n31328 ;
  assign n31330 = n15082 & ~n31316 ;
  assign n31331 = n31329 & ~n31330 ;
  assign n31332 = ~x785 & n31331 ;
  assign n31333 = ( x609 & x1155 ) | ( x609 & n31316 ) | ( x1155 & n31316 ) ;
  assign n31334 = ( ~x609 & x1155 ) | ( ~x609 & n31331 ) | ( x1155 & n31331 ) ;
  assign n31335 = n31333 & n31334 ;
  assign n31336 = ( x609 & x1155 ) | ( x609 & ~n31316 ) | ( x1155 & ~n31316 ) ;
  assign n31337 = ( x609 & ~x1155 ) | ( x609 & n31331 ) | ( ~x1155 & n31331 ) ;
  assign n31338 = ~n31336 & n31337 ;
  assign n31339 = n31335 | n31338 ;
  assign n31340 = x785 & n31339 ;
  assign n31341 = n31332 | n31340 ;
  assign n31342 = ~x781 & n31341 ;
  assign n31343 = ( x618 & x1154 ) | ( x618 & n31316 ) | ( x1154 & n31316 ) ;
  assign n31344 = ( ~x618 & x1154 ) | ( ~x618 & n31341 ) | ( x1154 & n31341 ) ;
  assign n31345 = n31343 & n31344 ;
  assign n31346 = ( x618 & x1154 ) | ( x618 & ~n31316 ) | ( x1154 & ~n31316 ) ;
  assign n31347 = ( x618 & ~x1154 ) | ( x618 & n31341 ) | ( ~x1154 & n31341 ) ;
  assign n31348 = ~n31346 & n31347 ;
  assign n31349 = n31345 | n31348 ;
  assign n31350 = x781 & n31349 ;
  assign n31351 = n31342 | n31350 ;
  assign n31352 = ~x789 & n31351 ;
  assign n31353 = ( x619 & x1159 ) | ( x619 & n31316 ) | ( x1159 & n31316 ) ;
  assign n31354 = ( ~x619 & x1159 ) | ( ~x619 & n31351 ) | ( x1159 & n31351 ) ;
  assign n31355 = n31353 & n31354 ;
  assign n31356 = ( x619 & x1159 ) | ( x619 & ~n31316 ) | ( x1159 & ~n31316 ) ;
  assign n31357 = ( x619 & ~x1159 ) | ( x619 & n31351 ) | ( ~x1159 & n31351 ) ;
  assign n31358 = ~n31356 & n31357 ;
  assign n31359 = n31355 | n31358 ;
  assign n31360 = x789 & n31359 ;
  assign n31361 = n31352 | n31360 ;
  assign n31362 = ~n16176 & n31361 ;
  assign n31363 = n16176 & n31316 ;
  assign n31364 = n31362 | n31363 ;
  assign n31365 = ~n15134 & n31364 ;
  assign n31366 = n15134 & n31316 ;
  assign n31367 = n31365 | n31366 ;
  assign n31368 = ~n15141 & n31367 ;
  assign n31369 = n15141 & n31316 ;
  assign n31370 = n31368 | n31369 ;
  assign n31371 = ( x644 & x715 ) | ( x644 & n31370 ) | ( x715 & n31370 ) ;
  assign n31372 = ( ~x644 & x715 ) | ( ~x644 & n31316 ) | ( x715 & n31316 ) ;
  assign n31373 = n31371 & n31372 ;
  assign n31374 = x1160 | n31373 ;
  assign n31375 = n15414 & ~n31316 ;
  assign n31376 = n15400 & ~n31316 ;
  assign n31377 = x643 | n31316 ;
  assign n31378 = x200 | n15070 ;
  assign n31379 = n17892 & n31378 ;
  assign n31380 = ( x200 & ~x299 ) | ( x200 & n15199 ) | ( ~x299 & n15199 ) ;
  assign n31381 = ( x200 & x299 ) | ( x200 & n15303 ) | ( x299 & n15303 ) ;
  assign n31382 = n31380 & ~n31381 ;
  assign n31383 = ( x200 & ~x299 ) | ( x200 & n15322 ) | ( ~x299 & n15322 ) ;
  assign n31384 = ( x200 & x299 ) | ( x200 & n15219 ) | ( x299 & n15219 ) ;
  assign n31385 = ~n31383 & n31384 ;
  assign n31386 = n31382 | n31385 ;
  assign n31387 = x39 & n31386 ;
  assign n31388 = ( ~x39 & x200 ) | ( ~x39 & n15369 ) | ( x200 & n15369 ) ;
  assign n31389 = ( x39 & x200 ) | ( x39 & n15345 ) | ( x200 & n15345 ) ;
  assign n31390 = n31388 & ~n31389 ;
  assign n31391 = n31387 | n31390 ;
  assign n31392 = ~x38 & n31391 ;
  assign n31393 = n31379 | n31392 ;
  assign n31394 = ~n2032 & n31393 ;
  assign n31395 = x643 & ~n31325 ;
  assign n31396 = ~n31394 & n31395 ;
  assign n31397 = n31377 & ~n31396 ;
  assign n31398 = ~x778 & n31397 ;
  assign n31399 = ( x625 & x1153 ) | ( x625 & n31316 ) | ( x1153 & n31316 ) ;
  assign n31400 = ( ~x625 & x1153 ) | ( ~x625 & n31397 ) | ( x1153 & n31397 ) ;
  assign n31401 = n31399 & n31400 ;
  assign n31402 = ( x625 & x1153 ) | ( x625 & ~n31316 ) | ( x1153 & ~n31316 ) ;
  assign n31403 = ( x625 & ~x1153 ) | ( x625 & n31397 ) | ( ~x1153 & n31397 ) ;
  assign n31404 = ~n31402 & n31403 ;
  assign n31405 = n31401 | n31404 ;
  assign n31406 = x778 & n31405 ;
  assign n31407 = n31398 | n31406 ;
  assign n31408 = n15400 | n31407 ;
  assign n31409 = ~n31376 & n31408 ;
  assign n31410 = ~n15407 & n31409 ;
  assign n31411 = n15407 & n31316 ;
  assign n31412 = n31410 | n31411 ;
  assign n31413 = n15414 | n31412 ;
  assign n31414 = ~n31375 & n31413 ;
  assign n31415 = ~n15421 & n31414 ;
  assign n31416 = n15421 & n31316 ;
  assign n31417 = n31415 | n31416 ;
  assign n31418 = ~x792 & n31417 ;
  assign n31419 = ( x628 & x1156 ) | ( x628 & n31316 ) | ( x1156 & n31316 ) ;
  assign n31420 = ( ~x628 & x1156 ) | ( ~x628 & n31417 ) | ( x1156 & n31417 ) ;
  assign n31421 = n31419 & n31420 ;
  assign n31422 = ( x628 & x1156 ) | ( x628 & ~n31316 ) | ( x1156 & ~n31316 ) ;
  assign n31423 = ( x628 & ~x1156 ) | ( x628 & n31417 ) | ( ~x1156 & n31417 ) ;
  assign n31424 = ~n31422 & n31423 ;
  assign n31425 = n31421 | n31424 ;
  assign n31426 = x792 & n31425 ;
  assign n31427 = n31418 | n31426 ;
  assign n31428 = ~x787 & n31427 ;
  assign n31429 = x647 & n31427 ;
  assign n31430 = ~x647 & n31316 ;
  assign n31431 = n31429 | n31430 ;
  assign n31432 = x1157 & n31431 ;
  assign n31433 = ( x647 & x1157 ) | ( x647 & ~n31316 ) | ( x1157 & ~n31316 ) ;
  assign n31434 = ( x647 & ~x1157 ) | ( x647 & n31427 ) | ( ~x1157 & n31427 ) ;
  assign n31435 = ~n31433 & n31434 ;
  assign n31436 = n31432 | n31435 ;
  assign n31437 = x787 & n31436 ;
  assign n31438 = n31428 | n31437 ;
  assign n31439 = ( x644 & x715 ) | ( x644 & ~n31438 ) | ( x715 & ~n31438 ) ;
  assign n31440 = n18621 & n31364 ;
  assign n31441 = ( x629 & n31424 ) | ( x629 & n31440 ) | ( n31424 & n31440 ) ;
  assign n31442 = ( ~x629 & n31421 ) | ( ~x629 & n31440 ) | ( n31421 & n31440 ) ;
  assign n31443 = n31441 | n31442 ;
  assign n31444 = x792 & n31443 ;
  assign n31445 = x648 & ~n31358 ;
  assign n31446 = ( x619 & x1159 ) | ( x619 & n31412 ) | ( x1159 & n31412 ) ;
  assign n31447 = x627 | n31345 ;
  assign n31448 = ( x618 & x1154 ) | ( x618 & ~n31409 ) | ( x1154 & ~n31409 ) ;
  assign n31449 = x660 | n31335 ;
  assign n31450 = ( x609 & x1155 ) | ( x609 & ~n31407 ) | ( x1155 & ~n31407 ) ;
  assign n31451 = x608 | n31401 ;
  assign n31452 = ( x625 & x1153 ) | ( x625 & ~n31328 ) | ( x1153 & ~n31328 ) ;
  assign n31453 = ~x643 & n31328 ;
  assign n31454 = n15375 | n15477 ;
  assign n31455 = n31379 & n31454 ;
  assign n31456 = ( ~x38 & x200 ) | ( ~x38 & n17568 ) | ( x200 & n17568 ) ;
  assign n31457 = ( x38 & x200 ) | ( x38 & n17577 ) | ( x200 & n17577 ) ;
  assign n31458 = n31456 & ~n31457 ;
  assign n31459 = n31455 | n31458 ;
  assign n31460 = x606 | n2032 ;
  assign n31461 = n31459 & ~n31460 ;
  assign n31462 = n17557 | n17558 ;
  assign n31463 = ~x200 & n31462 ;
  assign n31464 = x38 & x200 ;
  assign n31465 = n17550 & n31464 ;
  assign n31466 = x606 & ~n2032 ;
  assign n31467 = ~n31465 & n31466 ;
  assign n31468 = ~n31463 & n31467 ;
  assign n31469 = ( x38 & ~x200 ) | ( x38 & n17559 ) | ( ~x200 & n17559 ) ;
  assign n31470 = ( x38 & x200 ) | ( x38 & ~n22722 ) | ( x200 & ~n22722 ) ;
  assign n31471 = n31469 | n31470 ;
  assign n31472 = n31468 & n31471 ;
  assign n31473 = n31325 | n31472 ;
  assign n31474 = n31461 | n31473 ;
  assign n31475 = x643 & n31474 ;
  assign n31476 = n31453 | n31475 ;
  assign n31477 = ( x625 & ~x1153 ) | ( x625 & n31476 ) | ( ~x1153 & n31476 ) ;
  assign n31478 = ~n31452 & n31477 ;
  assign n31479 = n31451 | n31478 ;
  assign n31480 = x608 & ~n31404 ;
  assign n31481 = ( x625 & x1153 ) | ( x625 & n31328 ) | ( x1153 & n31328 ) ;
  assign n31482 = ( ~x625 & x1153 ) | ( ~x625 & n31476 ) | ( x1153 & n31476 ) ;
  assign n31483 = n31481 & n31482 ;
  assign n31484 = n31480 & ~n31483 ;
  assign n31485 = n31479 & ~n31484 ;
  assign n31486 = x778 & ~n31485 ;
  assign n31487 = x778 | n31476 ;
  assign n31488 = ~n31486 & n31487 ;
  assign n31489 = ( x609 & ~x1155 ) | ( x609 & n31488 ) | ( ~x1155 & n31488 ) ;
  assign n31490 = ~n31450 & n31489 ;
  assign n31491 = n31449 | n31490 ;
  assign n31492 = x660 & ~n31338 ;
  assign n31493 = ( x609 & x1155 ) | ( x609 & n31407 ) | ( x1155 & n31407 ) ;
  assign n31494 = ( ~x609 & x1155 ) | ( ~x609 & n31488 ) | ( x1155 & n31488 ) ;
  assign n31495 = n31493 & n31494 ;
  assign n31496 = n31492 & ~n31495 ;
  assign n31497 = n31491 & ~n31496 ;
  assign n31498 = x785 & ~n31497 ;
  assign n31499 = x785 | n31488 ;
  assign n31500 = ~n31498 & n31499 ;
  assign n31501 = ( x618 & ~x1154 ) | ( x618 & n31500 ) | ( ~x1154 & n31500 ) ;
  assign n31502 = ~n31448 & n31501 ;
  assign n31503 = n31447 | n31502 ;
  assign n31504 = x627 & ~n31348 ;
  assign n31505 = ( x618 & x1154 ) | ( x618 & n31409 ) | ( x1154 & n31409 ) ;
  assign n31506 = ( ~x618 & x1154 ) | ( ~x618 & n31500 ) | ( x1154 & n31500 ) ;
  assign n31507 = n31505 & n31506 ;
  assign n31508 = n31504 & ~n31507 ;
  assign n31509 = n31503 & ~n31508 ;
  assign n31510 = x781 & ~n31509 ;
  assign n31511 = x781 | n31500 ;
  assign n31512 = ~n31510 & n31511 ;
  assign n31513 = ( ~x619 & x1159 ) | ( ~x619 & n31512 ) | ( x1159 & n31512 ) ;
  assign n31514 = n31446 & n31513 ;
  assign n31515 = n31445 & ~n31514 ;
  assign n31516 = x648 | n31355 ;
  assign n31517 = ( x619 & x1159 ) | ( x619 & ~n31412 ) | ( x1159 & ~n31412 ) ;
  assign n31518 = ( x619 & ~x1159 ) | ( x619 & n31512 ) | ( ~x1159 & n31512 ) ;
  assign n31519 = ~n31517 & n31518 ;
  assign n31520 = n31516 | n31519 ;
  assign n31521 = x789 & n31520 ;
  assign n31522 = ~n31515 & n31521 ;
  assign n31523 = ~x789 & n31512 ;
  assign n31524 = n16177 | n31523 ;
  assign n31525 = n31522 | n31524 ;
  assign n31526 = n16115 & ~n31414 ;
  assign n31527 = ( x626 & ~n15419 ) | ( x626 & n31316 ) | ( ~n15419 & n31316 ) ;
  assign n31528 = ( x626 & n15419 ) | ( x626 & ~n31361 ) | ( n15419 & ~n31361 ) ;
  assign n31529 = ~n31527 & n31528 ;
  assign n31530 = n31526 | n31529 ;
  assign n31531 = ( x626 & n15418 ) | ( x626 & ~n31316 ) | ( n15418 & ~n31316 ) ;
  assign n31532 = ( x626 & ~n15418 ) | ( x626 & n31361 ) | ( ~n15418 & n31361 ) ;
  assign n31533 = n31531 & ~n31532 ;
  assign n31534 = n31530 | n31533 ;
  assign n31535 = x788 & n31534 ;
  assign n31536 = n18434 | n31535 ;
  assign n31537 = n31525 & ~n31536 ;
  assign n31538 = n31444 | n31537 ;
  assign n31539 = ~n18431 & n31538 ;
  assign n31540 = n15138 & n31431 ;
  assign n31541 = x630 & n31435 ;
  assign n31542 = n18610 & n31367 ;
  assign n31543 = n31541 | n31542 ;
  assign n31544 = n31540 | n31543 ;
  assign n31545 = x787 & n31544 ;
  assign n31546 = n31539 | n31545 ;
  assign n31547 = ( x644 & ~x715 ) | ( x644 & n31546 ) | ( ~x715 & n31546 ) ;
  assign n31548 = ~n31439 & n31547 ;
  assign n31549 = n31374 | n31548 ;
  assign n31550 = ( x644 & x715 ) | ( x644 & ~n31370 ) | ( x715 & ~n31370 ) ;
  assign n31551 = ( x644 & ~x715 ) | ( x644 & n31316 ) | ( ~x715 & n31316 ) ;
  assign n31552 = ~n31550 & n31551 ;
  assign n31553 = x1160 & ~n31552 ;
  assign n31554 = ( x644 & x715 ) | ( x644 & n31438 ) | ( x715 & n31438 ) ;
  assign n31555 = ( ~x644 & x715 ) | ( ~x644 & n31546 ) | ( x715 & n31546 ) ;
  assign n31556 = n31554 & n31555 ;
  assign n31557 = n31553 & ~n31556 ;
  assign n31558 = n31549 & ~n31557 ;
  assign n31559 = ( x790 & n6785 ) | ( x790 & n31558 ) | ( n6785 & n31558 ) ;
  assign n31560 = ( ~x790 & n6785 ) | ( ~x790 & n31546 ) | ( n6785 & n31546 ) ;
  assign n31561 = n31559 | n31560 ;
  assign n31562 = ~n31315 & n31561 ;
  assign n31563 = x233 & x237 ;
  assign n31564 = x96 & x210 ;
  assign n31565 = n14313 & ~n31564 ;
  assign n31566 = ~n5094 & n14313 ;
  assign n31567 = x96 & x198 ;
  assign n31568 = n5107 & n31567 ;
  assign n31569 = n14313 | n31568 ;
  assign n31570 = ~n31566 & n31569 ;
  assign n31571 = ~n31565 & n31570 ;
  assign n31572 = n31563 & n31571 ;
  assign n31573 = x201 & ~n31572 ;
  assign n31574 = x332 | n4708 ;
  assign n31575 = ~x947 & n31574 ;
  assign n31576 = x332 & n31564 ;
  assign n31577 = x32 & n11142 ;
  assign n31578 = x32 | x70 ;
  assign n31579 = ~n31577 & n31578 ;
  assign n31580 = ~x210 & n31579 ;
  assign n31581 = x32 | x96 ;
  assign n31582 = x70 & ~n31581 ;
  assign n31583 = x332 | n31582 ;
  assign n31584 = n31580 | n31583 ;
  assign n31585 = ~n31576 & n31584 ;
  assign n31586 = n4713 & n31585 ;
  assign n31587 = n4708 & ~n31586 ;
  assign n31588 = n31575 & ~n31587 ;
  assign n31589 = ( x947 & ~n4708 ) | ( x947 & n31585 ) | ( ~n4708 & n31585 ) ;
  assign n31590 = x332 & x468 ;
  assign n31591 = ~x468 & n31584 ;
  assign n31592 = n31590 | n31591 ;
  assign n31593 = ( x947 & n4708 ) | ( x947 & n31592 ) | ( n4708 & n31592 ) ;
  assign n31594 = n31589 & n31593 ;
  assign n31595 = n31588 | n31594 ;
  assign n31596 = x57 & n31595 ;
  assign n31597 = ~n1526 & n1592 ;
  assign n31598 = x95 | n1212 ;
  assign n31599 = n31597 & ~n31598 ;
  assign n31600 = x70 | n31599 ;
  assign n31601 = ~n31581 & n31600 ;
  assign n31602 = ( x210 & x332 ) | ( x210 & n31601 ) | ( x332 & n31601 ) ;
  assign n31603 = x95 | n1682 ;
  assign n31604 = n31577 | n31603 ;
  assign n31605 = n31597 & ~n31604 ;
  assign n31606 = n31579 | n31605 ;
  assign n31607 = ( ~x210 & x332 ) | ( ~x210 & n31606 ) | ( x332 & n31606 ) ;
  assign n31608 = n31602 | n31607 ;
  assign n31609 = ~n31576 & n31608 ;
  assign n31610 = n4713 & n31609 ;
  assign n31611 = n4708 & ~n31610 ;
  assign n31612 = n31575 & ~n31611 ;
  assign n31613 = x299 & ~n31612 ;
  assign n31614 = ( x947 & ~n4708 ) | ( x947 & n31609 ) | ( ~n4708 & n31609 ) ;
  assign n31615 = ~x468 & n31608 ;
  assign n31616 = n31590 | n31615 ;
  assign n31617 = ( x947 & n4708 ) | ( x947 & n31616 ) | ( n4708 & n31616 ) ;
  assign n31618 = n31614 & n31617 ;
  assign n31619 = n31613 & ~n31618 ;
  assign n31620 = ( x198 & x332 ) | ( x198 & n31601 ) | ( x332 & n31601 ) ;
  assign n31621 = ( ~x198 & x332 ) | ( ~x198 & n31606 ) | ( x332 & n31606 ) ;
  assign n31622 = n31620 | n31621 ;
  assign n31623 = ~x468 & n31622 ;
  assign n31624 = n4708 | n31590 ;
  assign n31625 = n31623 | n31624 ;
  assign n31626 = x332 & n31567 ;
  assign n31627 = n31622 & ~n31626 ;
  assign n31628 = n4708 & ~n31627 ;
  assign n31629 = x587 & ~n31628 ;
  assign n31630 = n31625 & n31629 ;
  assign n31631 = ~x587 & n31574 ;
  assign n31632 = n5150 & n31627 ;
  assign n31633 = ( ~n4708 & n31631 ) | ( ~n4708 & n31632 ) | ( n31631 & n31632 ) ;
  assign n31634 = x299 | n31633 ;
  assign n31635 = n31630 | n31634 ;
  assign n31636 = ~n31619 & n31635 ;
  assign n31637 = n5844 | n31636 ;
  assign n31638 = x95 | n1642 ;
  assign n31639 = ~x70 & n31638 ;
  assign n31640 = n31581 | n31639 ;
  assign n31641 = ( x210 & x332 ) | ( x210 & ~n31640 ) | ( x332 & ~n31640 ) ;
  assign n31642 = n1257 | n31604 ;
  assign n31643 = n1273 | n31642 ;
  assign n31644 = ~n31579 & n31643 ;
  assign n31645 = ( x210 & ~x332 ) | ( x210 & n31644 ) | ( ~x332 & n31644 ) ;
  assign n31646 = ~n31641 & n31645 ;
  assign n31647 = n31576 | n31646 ;
  assign n31648 = n4713 & ~n31647 ;
  assign n31649 = n4708 & ~n31648 ;
  assign n31650 = n31575 & ~n31649 ;
  assign n31651 = ( ~x947 & n4708 ) | ( ~x947 & n31647 ) | ( n4708 & n31647 ) ;
  assign n31652 = x468 | n31646 ;
  assign n31653 = ~n31590 & n31652 ;
  assign n31654 = ( x947 & n4708 ) | ( x947 & ~n31653 ) | ( n4708 & ~n31653 ) ;
  assign n31655 = ~n31651 & n31654 ;
  assign n31656 = n31650 | n31655 ;
  assign n31657 = ( x299 & ~n13580 ) | ( x299 & n31656 ) | ( ~n13580 & n31656 ) ;
  assign n31658 = ( x198 & x332 ) | ( x198 & ~n31640 ) | ( x332 & ~n31640 ) ;
  assign n31659 = ( x198 & ~x332 ) | ( x198 & n31644 ) | ( ~x332 & n31644 ) ;
  assign n31660 = ~n31658 & n31659 ;
  assign n31661 = x468 | n31660 ;
  assign n31662 = ~n31624 & n31661 ;
  assign n31663 = n31626 | n31660 ;
  assign n31664 = n4708 & n31663 ;
  assign n31665 = x587 & ~n31664 ;
  assign n31666 = ~n31662 & n31665 ;
  assign n31667 = n5150 & ~n31663 ;
  assign n31668 = ( ~n4708 & n31631 ) | ( ~n4708 & n31667 ) | ( n31631 & n31667 ) ;
  assign n31669 = n31666 | n31668 ;
  assign n31670 = ( x299 & n13580 ) | ( x299 & ~n31669 ) | ( n13580 & ~n31669 ) ;
  assign n31671 = ~n31657 & n31670 ;
  assign n31672 = n31637 & ~n31671 ;
  assign n31673 = x74 | n31672 ;
  assign n31674 = x299 & n31595 ;
  assign n31675 = x74 | n2005 ;
  assign n31676 = ~x198 & n31579 ;
  assign n31677 = n31583 | n31676 ;
  assign n31678 = n5107 & n31677 ;
  assign n31679 = n31574 | n31678 ;
  assign n31680 = ~n31626 & n31677 ;
  assign n31681 = n4708 & ~n31680 ;
  assign n31682 = ~x299 & n5106 ;
  assign n31683 = ~n31681 & n31682 ;
  assign n31684 = n31679 & n31683 ;
  assign n31685 = n31675 & ~n31684 ;
  assign n31686 = ~n31674 & n31685 ;
  assign n31687 = x55 | n31686 ;
  assign n31688 = n31673 & ~n31687 ;
  assign n31689 = n2033 & ~n31595 ;
  assign n31690 = n2033 | n31656 ;
  assign n31691 = ~n31689 & n31690 ;
  assign n31692 = x55 & n31691 ;
  assign n31693 = n2058 | n31692 ;
  assign n31694 = n31688 | n31693 ;
  assign n31695 = n2058 & ~n31595 ;
  assign n31696 = x59 | n31695 ;
  assign n31697 = n31694 & ~n31696 ;
  assign n31698 = ( x59 & ~n5086 ) | ( x59 & n31595 ) | ( ~n5086 & n31595 ) ;
  assign n31699 = ( x59 & n5086 ) | ( x59 & n31691 ) | ( n5086 & n31691 ) ;
  assign n31700 = n31698 & n31699 ;
  assign n31701 = n31697 | n31700 ;
  assign n31702 = ~x57 & n31701 ;
  assign n31703 = n31596 | n31702 ;
  assign n31704 = ( x201 & n31563 ) | ( x201 & ~n31703 ) | ( n31563 & ~n31703 ) ;
  assign n31705 = x57 & x332 ;
  assign n31706 = x332 & n2058 ;
  assign n31707 = x59 | n31706 ;
  assign n31708 = x74 & x332 ;
  assign n31709 = x55 | n31708 ;
  assign n31710 = n1592 & ~n9243 ;
  assign n31711 = ~x299 & x587 ;
  assign n31712 = n19097 | n31711 ;
  assign n31713 = ( x468 & n31710 ) | ( x468 & n31712 ) | ( n31710 & n31712 ) ;
  assign n31714 = ( ~x468 & n4708 ) | ( ~x468 & n31710 ) | ( n4708 & n31710 ) ;
  assign n31715 = n31713 & n31714 ;
  assign n31716 = x332 | n31715 ;
  assign n31717 = ~n5844 & n31716 ;
  assign n31718 = ~n1868 & n5135 ;
  assign n31719 = x332 | n31718 ;
  assign n31720 = n13580 & n31719 ;
  assign n31721 = x332 & n2005 ;
  assign n31722 = n31720 | n31721 ;
  assign n31723 = n31717 | n31722 ;
  assign n31724 = ~x74 & n31723 ;
  assign n31725 = n31709 | n31724 ;
  assign n31726 = ~n2033 & n5094 ;
  assign n31727 = ~n1868 & n31726 ;
  assign n31728 = x332 | n31727 ;
  assign n31729 = x55 & ~n31728 ;
  assign n31730 = n2058 | n31729 ;
  assign n31731 = n31725 & ~n31730 ;
  assign n31732 = n31707 | n31731 ;
  assign n31733 = ~n5086 & n31728 ;
  assign n31734 = x332 & n5086 ;
  assign n31735 = x59 & ~n31734 ;
  assign n31736 = ~n31733 & n31735 ;
  assign n31737 = x57 | n31736 ;
  assign n31738 = n31732 & ~n31737 ;
  assign n31739 = n31705 | n31738 ;
  assign n31740 = ( ~x201 & n31563 ) | ( ~x201 & n31739 ) | ( n31563 & n31739 ) ;
  assign n31741 = ~n31704 & n31740 ;
  assign n31742 = n31573 | n31741 ;
  assign n31743 = ~x233 & x237 ;
  assign n31744 = n31571 & n31743 ;
  assign n31745 = x202 & ~n31744 ;
  assign n31746 = ( x202 & ~n31703 ) | ( x202 & n31743 ) | ( ~n31703 & n31743 ) ;
  assign n31747 = ( ~x202 & n31739 ) | ( ~x202 & n31743 ) | ( n31739 & n31743 ) ;
  assign n31748 = ~n31746 & n31747 ;
  assign n31749 = n31745 | n31748 ;
  assign n31750 = x233 | x237 ;
  assign n31751 = n31571 & ~n31750 ;
  assign n31752 = x203 & ~n31751 ;
  assign n31753 = ( x203 & ~n31739 ) | ( x203 & n31750 ) | ( ~n31739 & n31750 ) ;
  assign n31754 = ( ~x203 & n31703 ) | ( ~x203 & n31750 ) | ( n31703 & n31750 ) ;
  assign n31755 = ~n31753 & n31754 ;
  assign n31756 = n31752 | n31755 ;
  assign n31757 = ~n4837 & n14313 ;
  assign n31758 = n31565 | n31757 ;
  assign n31759 = n4845 | n14313 ;
  assign n31760 = ( n14313 & n31567 ) | ( n14313 & n31759 ) | ( n31567 & n31759 ) ;
  assign n31761 = ~n31758 & n31760 ;
  assign n31762 = n31563 & n31761 ;
  assign n31763 = x204 & ~n31762 ;
  assign n31764 = x332 | n4711 ;
  assign n31765 = ~x907 & n31764 ;
  assign n31766 = n4711 & ~n31586 ;
  assign n31767 = n31765 & ~n31766 ;
  assign n31768 = ( x907 & ~n4711 ) | ( x907 & n31585 ) | ( ~n4711 & n31585 ) ;
  assign n31769 = ( x907 & n4711 ) | ( x907 & n31592 ) | ( n4711 & n31592 ) ;
  assign n31770 = n31768 & n31769 ;
  assign n31771 = n31767 | n31770 ;
  assign n31772 = x57 & n31771 ;
  assign n31773 = x332 & n14553 ;
  assign n31774 = x680 & ~n31773 ;
  assign n31775 = ~n31648 & n31774 ;
  assign n31776 = n31765 & ~n31775 ;
  assign n31777 = ( ~x907 & n4711 ) | ( ~x907 & n31647 ) | ( n4711 & n31647 ) ;
  assign n31778 = ( x907 & n4711 ) | ( x907 & ~n31653 ) | ( n4711 & ~n31653 ) ;
  assign n31779 = ~n31777 & n31778 ;
  assign n31780 = n31776 | n31779 ;
  assign n31781 = x299 & ~n31780 ;
  assign n31782 = n4711 & n31567 ;
  assign n31783 = x332 & ~n31782 ;
  assign n31784 = x299 | n31783 ;
  assign n31785 = n4845 & ~n31663 ;
  assign n31786 = n31784 | n31785 ;
  assign n31787 = ~n31781 & n31786 ;
  assign n31788 = n13580 & ~n31787 ;
  assign n31789 = n4845 & n31627 ;
  assign n31790 = n31784 | n31789 ;
  assign n31791 = n4711 & ~n31610 ;
  assign n31792 = n31765 & ~n31791 ;
  assign n31793 = x299 & ~n31792 ;
  assign n31794 = ( x907 & ~n4711 ) | ( x907 & n31609 ) | ( ~n4711 & n31609 ) ;
  assign n31795 = ( x907 & n4711 ) | ( x907 & n31616 ) | ( n4711 & n31616 ) ;
  assign n31796 = n31794 & n31795 ;
  assign n31797 = n31793 & ~n31796 ;
  assign n31798 = n31790 & ~n31797 ;
  assign n31799 = n5844 | n31798 ;
  assign n31800 = ~n31788 & n31799 ;
  assign n31801 = x74 | n31800 ;
  assign n31802 = ~x468 & x602 ;
  assign n31803 = x468 & n4711 ;
  assign n31804 = n31802 | n31803 ;
  assign n31805 = n31680 & n31804 ;
  assign n31806 = n31783 | n31805 ;
  assign n31807 = ( x299 & n31675 ) | ( x299 & ~n31806 ) | ( n31675 & ~n31806 ) ;
  assign n31808 = ( x299 & ~n31675 ) | ( x299 & n31771 ) | ( ~n31675 & n31771 ) ;
  assign n31809 = n31807 & ~n31808 ;
  assign n31810 = x55 | n31809 ;
  assign n31811 = n31801 & ~n31810 ;
  assign n31812 = n2033 & ~n31771 ;
  assign n31813 = n2033 | n31780 ;
  assign n31814 = ~n31812 & n31813 ;
  assign n31815 = x55 & n31814 ;
  assign n31816 = n2058 | n31815 ;
  assign n31817 = n31811 | n31816 ;
  assign n31818 = n2058 & ~n31771 ;
  assign n31819 = x59 | n31818 ;
  assign n31820 = n31817 & ~n31819 ;
  assign n31821 = ( x59 & ~n5086 ) | ( x59 & n31771 ) | ( ~n5086 & n31771 ) ;
  assign n31822 = ( x59 & n5086 ) | ( x59 & n31814 ) | ( n5086 & n31814 ) ;
  assign n31823 = n31821 & n31822 ;
  assign n31824 = n31820 | n31823 ;
  assign n31825 = ~x57 & n31824 ;
  assign n31826 = n31772 | n31825 ;
  assign n31827 = ( x204 & n31563 ) | ( x204 & ~n31826 ) | ( n31563 & ~n31826 ) ;
  assign n31828 = ~x299 & n31804 ;
  assign n31829 = n5013 | n31828 ;
  assign n31830 = ~n1868 & n31829 ;
  assign n31831 = x332 | n31830 ;
  assign n31832 = n13580 & n31831 ;
  assign n31833 = ( x299 & x468 ) | ( x299 & ~x907 ) | ( x468 & ~x907 ) ;
  assign n31834 = ( x299 & ~x468 ) | ( x299 & x602 ) | ( ~x468 & x602 ) ;
  assign n31835 = ~n31833 & n31834 ;
  assign n31836 = n31803 | n31835 ;
  assign n31837 = n31710 & n31836 ;
  assign n31838 = x332 | n31837 ;
  assign n31839 = ~n5844 & n31838 ;
  assign n31840 = n31832 | n31839 ;
  assign n31841 = ~x74 & n31840 ;
  assign n31842 = n31709 | n31721 ;
  assign n31843 = n31841 | n31842 ;
  assign n31844 = ~n2033 & n4837 ;
  assign n31845 = ~n1868 & n31844 ;
  assign n31846 = x332 | n31845 ;
  assign n31847 = x55 & ~n31846 ;
  assign n31848 = n2058 | n31847 ;
  assign n31849 = n31843 & ~n31848 ;
  assign n31850 = n31707 | n31849 ;
  assign n31851 = ~n5086 & n31846 ;
  assign n31852 = n31735 & ~n31851 ;
  assign n31853 = x57 | n31852 ;
  assign n31854 = n31850 & ~n31853 ;
  assign n31855 = n31705 | n31854 ;
  assign n31856 = ( ~x204 & n31563 ) | ( ~x204 & n31855 ) | ( n31563 & n31855 ) ;
  assign n31857 = ~n31827 & n31856 ;
  assign n31858 = n31763 | n31857 ;
  assign n31859 = n31743 & n31761 ;
  assign n31860 = x205 & ~n31859 ;
  assign n31861 = ( x205 & n31743 ) | ( x205 & ~n31826 ) | ( n31743 & ~n31826 ) ;
  assign n31862 = ( ~x205 & n31743 ) | ( ~x205 & n31855 ) | ( n31743 & n31855 ) ;
  assign n31863 = ~n31861 & n31862 ;
  assign n31864 = n31860 | n31863 ;
  assign n31865 = x233 & ~x237 ;
  assign n31866 = n31761 & n31865 ;
  assign n31867 = x206 & ~n31866 ;
  assign n31868 = ( x206 & ~n31826 ) | ( x206 & n31865 ) | ( ~n31826 & n31865 ) ;
  assign n31869 = ( ~x206 & n31855 ) | ( ~x206 & n31865 ) | ( n31855 & n31865 ) ;
  assign n31870 = ~n31868 & n31869 ;
  assign n31871 = n31867 | n31870 ;
  assign n31872 = ~x207 & n6785 ;
  assign n31873 = x207 | n14834 ;
  assign n31874 = n15141 & n31873 ;
  assign n31875 = x623 | n31873 ;
  assign n31876 = ~n2032 & n22415 ;
  assign n31877 = ~n15082 & n31876 ;
  assign n31878 = ~n18257 & n31877 ;
  assign n31879 = ~n18249 & n31878 ;
  assign n31880 = ~n18253 & n31879 ;
  assign n31881 = ~n16176 & n31880 ;
  assign n31882 = ~n15134 & n31881 ;
  assign n31883 = ( ~x207 & x623 ) | ( ~x207 & n31882 ) | ( x623 & n31882 ) ;
  assign n31884 = ~n14834 & n15082 ;
  assign n31885 = ~n2032 & n17421 ;
  assign n31886 = n15082 | n31885 ;
  assign n31887 = ~n31884 & n31886 ;
  assign n31888 = x785 | n31887 ;
  assign n31889 = ~n14834 & n15094 ;
  assign n31890 = x609 | n31886 ;
  assign n31891 = ~n31889 & n31890 ;
  assign n31892 = x1155 | n31891 ;
  assign n31893 = n14834 | n15088 ;
  assign n31894 = x609 & ~n31886 ;
  assign n31895 = n31893 & ~n31894 ;
  assign n31896 = x1155 & ~n31895 ;
  assign n31897 = n31892 & ~n31896 ;
  assign n31898 = x785 & ~n31897 ;
  assign n31899 = n31888 & ~n31898 ;
  assign n31900 = x781 | n31899 ;
  assign n31901 = ( x618 & x1154 ) | ( x618 & n14834 ) | ( x1154 & n14834 ) ;
  assign n31902 = ( ~x618 & x1154 ) | ( ~x618 & n31899 ) | ( x1154 & n31899 ) ;
  assign n31903 = n31901 | n31902 ;
  assign n31904 = ( x618 & x1154 ) | ( x618 & ~n14834 ) | ( x1154 & ~n14834 ) ;
  assign n31905 = ( x618 & ~x1154 ) | ( x618 & n31899 ) | ( ~x1154 & n31899 ) ;
  assign n31906 = n31904 & ~n31905 ;
  assign n31907 = n31903 & ~n31906 ;
  assign n31908 = x781 & ~n31907 ;
  assign n31909 = n31900 & ~n31908 ;
  assign n31910 = x789 | n31909 ;
  assign n31911 = ( x619 & x1159 ) | ( x619 & n14834 ) | ( x1159 & n14834 ) ;
  assign n31912 = ( ~x619 & x1159 ) | ( ~x619 & n31909 ) | ( x1159 & n31909 ) ;
  assign n31913 = n31911 | n31912 ;
  assign n31914 = ( x619 & x1159 ) | ( x619 & ~n14834 ) | ( x1159 & ~n14834 ) ;
  assign n31915 = ( x619 & ~x1159 ) | ( x619 & n31909 ) | ( ~x1159 & n31909 ) ;
  assign n31916 = n31914 & ~n31915 ;
  assign n31917 = n31913 & ~n31916 ;
  assign n31918 = x789 & ~n31917 ;
  assign n31919 = n31910 & ~n31918 ;
  assign n31920 = ~n16176 & n31919 ;
  assign n31921 = n14834 & n16176 ;
  assign n31922 = n31920 | n31921 ;
  assign n31923 = ~n15134 & n31922 ;
  assign n31924 = n14834 & n15134 ;
  assign n31925 = n31923 | n31924 ;
  assign n31926 = ( x207 & x623 ) | ( x207 & ~n31925 ) | ( x623 & ~n31925 ) ;
  assign n31927 = n31883 & n31926 ;
  assign n31928 = n31875 & ~n31927 ;
  assign n31929 = ~n15141 & n31928 ;
  assign n31930 = n31874 | n31929 ;
  assign n31931 = ( x644 & x715 ) | ( x644 & ~n31930 ) | ( x715 & ~n31930 ) ;
  assign n31932 = ( x644 & ~x715 ) | ( x644 & n31873 ) | ( ~x715 & n31873 ) ;
  assign n31933 = ~n31931 & n31932 ;
  assign n31934 = x1160 & ~n31933 ;
  assign n31935 = ~x710 & n31873 ;
  assign n31936 = ~n17210 & n22357 ;
  assign n31937 = ~n17215 & n31936 ;
  assign n31938 = ~n17220 & n31937 ;
  assign n31939 = ( x207 & ~x710 ) | ( x207 & n31938 ) | ( ~x710 & n31938 ) ;
  assign n31940 = ~n14834 & n15414 ;
  assign n31941 = ~n2032 & n22362 ;
  assign n31942 = x778 | n31941 ;
  assign n31943 = x625 | n14834 ;
  assign n31944 = x625 & ~n31941 ;
  assign n31945 = n31943 & ~n31944 ;
  assign n31946 = x1153 & ~n31945 ;
  assign n31947 = x625 & ~n14834 ;
  assign n31948 = x625 | n31941 ;
  assign n31949 = ~n31947 & n31948 ;
  assign n31950 = x1153 | n31949 ;
  assign n31951 = ~n31946 & n31950 ;
  assign n31952 = x778 & ~n31951 ;
  assign n31953 = n31942 & ~n31952 ;
  assign n31954 = n15400 | n31953 ;
  assign n31955 = ~n14834 & n15400 ;
  assign n31956 = n31954 & ~n31955 ;
  assign n31957 = ~n15407 & n31956 ;
  assign n31958 = n14834 & n15407 ;
  assign n31959 = n31957 | n31958 ;
  assign n31960 = n15414 | n31959 ;
  assign n31961 = ~n31940 & n31960 ;
  assign n31962 = ~n15421 & n31961 ;
  assign n31963 = n14834 & n15421 ;
  assign n31964 = n31962 | n31963 ;
  assign n31965 = ~n17220 & n31964 ;
  assign n31966 = n14834 & n16054 ;
  assign n31967 = n31965 | n31966 ;
  assign n31968 = ( x207 & x710 ) | ( x207 & n31967 ) | ( x710 & n31967 ) ;
  assign n31969 = ~n31939 & n31968 ;
  assign n31970 = n31935 | n31969 ;
  assign n31971 = ~x787 & n31970 ;
  assign n31972 = ( x647 & x1157 ) | ( x647 & ~n31873 ) | ( x1157 & ~n31873 ) ;
  assign n31973 = ( x647 & ~x1157 ) | ( x647 & n31970 ) | ( ~x1157 & n31970 ) ;
  assign n31974 = ~n31972 & n31973 ;
  assign n31975 = ( x647 & x1157 ) | ( x647 & n31873 ) | ( x1157 & n31873 ) ;
  assign n31976 = ( ~x647 & x1157 ) | ( ~x647 & n31970 ) | ( x1157 & n31970 ) ;
  assign n31977 = n31975 & n31976 ;
  assign n31978 = n31974 | n31977 ;
  assign n31979 = x787 & n31978 ;
  assign n31980 = n31971 | n31979 ;
  assign n31981 = ( x644 & x715 ) | ( x644 & n31980 ) | ( x715 & n31980 ) ;
  assign n31982 = n18610 & n31928 ;
  assign n31983 = ( x630 & n31974 ) | ( x630 & n31982 ) | ( n31974 & n31982 ) ;
  assign n31984 = ( ~x630 & n31977 ) | ( ~x630 & n31982 ) | ( n31977 & n31982 ) ;
  assign n31985 = n31983 | n31984 ;
  assign n31986 = x787 & n31985 ;
  assign n31987 = x1156 | n31937 ;
  assign n31988 = n18617 & n31987 ;
  assign n31989 = x1156 & ~n31937 ;
  assign n31990 = n18619 & ~n31989 ;
  assign n31991 = ( x1156 & n31881 ) | ( x1156 & n31990 ) | ( n31881 & n31990 ) ;
  assign n31992 = x1156 & ~n31990 ;
  assign n31993 = ( n31988 & n31991 ) | ( n31988 & ~n31992 ) | ( n31991 & ~n31992 ) ;
  assign n31994 = x792 & n31993 ;
  assign n31995 = ~n17214 & n31936 ;
  assign n31996 = ~n15414 & n31995 ;
  assign n31997 = x626 & ~n31996 ;
  assign n31998 = x641 | n31997 ;
  assign n31999 = ~x619 & x648 ;
  assign n32000 = ( x1159 & n31879 ) | ( x1159 & n31999 ) | ( n31879 & n31999 ) ;
  assign n32001 = ( ~x1159 & n31995 ) | ( ~x1159 & n31999 ) | ( n31995 & n31999 ) ;
  assign n32002 = n32000 & n32001 ;
  assign n32003 = x789 & ~n32002 ;
  assign n32004 = x619 & ~x648 ;
  assign n32005 = ( ~x1159 & n31879 ) | ( ~x1159 & n32004 ) | ( n31879 & n32004 ) ;
  assign n32006 = ( x1159 & n31995 ) | ( x1159 & n32004 ) | ( n31995 & n32004 ) ;
  assign n32007 = n32005 & n32006 ;
  assign n32008 = n32003 & ~n32007 ;
  assign n32009 = x789 & ~n32008 ;
  assign n32010 = ~n15400 & n31936 ;
  assign n32011 = x618 & ~n32010 ;
  assign n32012 = x1154 | n32011 ;
  assign n32013 = n18246 & n31878 ;
  assign n32014 = x627 | n32013 ;
  assign n32015 = n32012 & ~n32014 ;
  assign n32016 = x778 | n31178 ;
  assign n32017 = ~x625 & n22357 ;
  assign n32018 = x1153 | n32017 ;
  assign n32019 = x608 & n32018 ;
  assign n32020 = ( x625 & x1153 ) | ( x625 & ~n31876 ) | ( x1153 & ~n31876 ) ;
  assign n32021 = ( x625 & ~x1153 ) | ( x625 & n31178 ) | ( ~x1153 & n31178 ) ;
  assign n32022 = n32020 & ~n32021 ;
  assign n32023 = n32019 & ~n32022 ;
  assign n32024 = x625 & n22357 ;
  assign n32025 = x1153 & ~n32024 ;
  assign n32026 = x608 | n32025 ;
  assign n32027 = ( x625 & x1153 ) | ( x625 & n31876 ) | ( x1153 & n31876 ) ;
  assign n32028 = ( ~x625 & x1153 ) | ( ~x625 & n31178 ) | ( x1153 & n31178 ) ;
  assign n32029 = n32027 | n32028 ;
  assign n32030 = ~n32026 & n32029 ;
  assign n32031 = x778 & ~n32030 ;
  assign n32032 = ~n32023 & n32031 ;
  assign n32033 = n32016 & ~n32032 ;
  assign n32034 = x785 | n32033 ;
  assign n32035 = x609 | n32033 ;
  assign n32036 = x609 & ~n31936 ;
  assign n32037 = x1155 | n32036 ;
  assign n32038 = n32035 & ~n32037 ;
  assign n32039 = n18136 & n31877 ;
  assign n32040 = x660 | n32039 ;
  assign n32041 = n32038 | n32040 ;
  assign n32042 = x609 & ~n32033 ;
  assign n32043 = x609 | n31936 ;
  assign n32044 = x1155 & n32043 ;
  assign n32045 = ~n32042 & n32044 ;
  assign n32046 = ~n18085 & n31877 ;
  assign n32047 = x660 & ~n32046 ;
  assign n32048 = ~n32045 & n32047 ;
  assign n32049 = n32041 & ~n32048 ;
  assign n32050 = x785 & ~n32049 ;
  assign n32051 = n32034 & ~n32050 ;
  assign n32052 = x618 & ~n32051 ;
  assign n32053 = x618 | n32010 ;
  assign n32054 = x1154 & n32053 ;
  assign n32055 = ~n32052 & n32054 ;
  assign n32056 = ~n18247 & n31878 ;
  assign n32057 = x627 & ~n32056 ;
  assign n32058 = ~n32055 & n32057 ;
  assign n32059 = n32015 | n32058 ;
  assign n32060 = x781 & n32059 ;
  assign n32061 = x618 | x627 ;
  assign n32062 = x781 & n32061 ;
  assign n32063 = n32051 | n32062 ;
  assign n32064 = n15413 | n21632 ;
  assign n32065 = n32008 & n32064 ;
  assign n32066 = n32063 & ~n32065 ;
  assign n32067 = ~n32060 & n32066 ;
  assign n32068 = n32009 | n32067 ;
  assign n32069 = x626 | n32068 ;
  assign n32070 = ~n31998 & n32069 ;
  assign n32071 = n16112 & n31880 ;
  assign n32072 = x1158 | n32071 ;
  assign n32073 = n32070 | n32072 ;
  assign n32074 = x626 | n31996 ;
  assign n32075 = x641 & n32074 ;
  assign n32076 = x626 & ~n32068 ;
  assign n32077 = n32075 & ~n32076 ;
  assign n32078 = n16113 & n31880 ;
  assign n32079 = x1158 & ~n32078 ;
  assign n32080 = ~n32077 & n32079 ;
  assign n32081 = n32073 & ~n32080 ;
  assign n32082 = ( x788 & n18434 ) | ( x788 & ~n32081 ) | ( n18434 & ~n32081 ) ;
  assign n32083 = ( x788 & ~n18434 ) | ( x788 & n32068 ) | ( ~n18434 & n32068 ) ;
  assign n32084 = ~n32082 & n32083 ;
  assign n32085 = n31994 | n32084 ;
  assign n32086 = ( x207 & ~x623 ) | ( x207 & n32085 ) | ( ~x623 & n32085 ) ;
  assign n32087 = x619 | n31959 ;
  assign n32088 = x618 & ~n31956 ;
  assign n32089 = x609 & ~n31953 ;
  assign n32090 = ~n2032 & n17554 ;
  assign n32091 = x778 | n32090 ;
  assign n32092 = x608 | n31946 ;
  assign n32093 = ( x625 & x1153 ) | ( x625 & n31885 ) | ( x1153 & n31885 ) ;
  assign n32094 = ( ~x625 & x1153 ) | ( ~x625 & n32090 ) | ( x1153 & n32090 ) ;
  assign n32095 = n32093 | n32094 ;
  assign n32096 = ~n32092 & n32095 ;
  assign n32097 = x608 & n31950 ;
  assign n32098 = ( x625 & x1153 ) | ( x625 & ~n31885 ) | ( x1153 & ~n31885 ) ;
  assign n32099 = ( x625 & ~x1153 ) | ( x625 & n32090 ) | ( ~x1153 & n32090 ) ;
  assign n32100 = n32098 & ~n32099 ;
  assign n32101 = n32097 & ~n32100 ;
  assign n32102 = x778 & ~n32101 ;
  assign n32103 = ~n32096 & n32102 ;
  assign n32104 = n32091 & ~n32103 ;
  assign n32105 = x609 | n32104 ;
  assign n32106 = ~n32089 & n32105 ;
  assign n32107 = x1155 | n32106 ;
  assign n32108 = x660 | n31896 ;
  assign n32109 = n32107 & ~n32108 ;
  assign n32110 = x609 | n31953 ;
  assign n32111 = x609 & ~n32104 ;
  assign n32112 = n32110 & ~n32111 ;
  assign n32113 = x1155 & ~n32112 ;
  assign n32114 = x660 & n31892 ;
  assign n32115 = ~n32113 & n32114 ;
  assign n32116 = n32109 | n32115 ;
  assign n32117 = x785 & n32116 ;
  assign n32118 = ~x785 & n32104 ;
  assign n32119 = n32117 | n32118 ;
  assign n32120 = x618 | n32119 ;
  assign n32121 = ~n32088 & n32120 ;
  assign n32122 = x1154 | n32121 ;
  assign n32123 = x627 | n31906 ;
  assign n32124 = n32122 & ~n32123 ;
  assign n32125 = x618 | n31956 ;
  assign n32126 = x618 & ~n32119 ;
  assign n32127 = n32125 & ~n32126 ;
  assign n32128 = x1154 & ~n32127 ;
  assign n32129 = x627 & n31903 ;
  assign n32130 = ~n32128 & n32129 ;
  assign n32131 = n32124 | n32130 ;
  assign n32132 = x781 & n32131 ;
  assign n32133 = ~x781 & n32119 ;
  assign n32134 = n32132 | n32133 ;
  assign n32135 = x619 & ~n32134 ;
  assign n32136 = n32087 & ~n32135 ;
  assign n32137 = x1159 & ~n32136 ;
  assign n32138 = x648 & n31913 ;
  assign n32139 = ~n32137 & n32138 ;
  assign n32140 = x619 & ~n31959 ;
  assign n32141 = x619 | n32134 ;
  assign n32142 = ~n32140 & n32141 ;
  assign n32143 = x1159 | n32142 ;
  assign n32144 = x648 | n31916 ;
  assign n32145 = n32143 & ~n32144 ;
  assign n32146 = x789 & ~n32145 ;
  assign n32147 = ~n32139 & n32146 ;
  assign n32148 = x789 | n32134 ;
  assign n32149 = ~n16177 & n32148 ;
  assign n32150 = ~n32147 & n32149 ;
  assign n32151 = n15420 & n16114 ;
  assign n32152 = n31919 & n32151 ;
  assign n32153 = x641 | n14834 ;
  assign n32154 = n16109 & n32153 ;
  assign n32155 = x641 & ~n14834 ;
  assign n32156 = n16110 & ~n32155 ;
  assign n32157 = ( x641 & n31961 ) | ( x641 & n32156 ) | ( n31961 & n32156 ) ;
  assign n32158 = x641 & ~n32156 ;
  assign n32159 = ( n32154 & n32157 ) | ( n32154 & ~n32158 ) | ( n32157 & ~n32158 ) ;
  assign n32160 = n32152 | n32159 ;
  assign n32161 = x788 & n32160 ;
  assign n32162 = n18434 | n32161 ;
  assign n32163 = n32150 | n32162 ;
  assign n32164 = x628 | n14834 ;
  assign n32165 = x628 & ~n31964 ;
  assign n32166 = n32164 & ~n32165 ;
  assign n32167 = x629 | n32166 ;
  assign n32168 = x1156 & ~n32167 ;
  assign n32169 = x628 & ~n14834 ;
  assign n32170 = x628 | n31964 ;
  assign n32171 = ~n32169 & n32170 ;
  assign n32172 = n15132 & ~n32171 ;
  assign n32173 = n18621 & ~n31922 ;
  assign n32174 = n32172 | n32173 ;
  assign n32175 = n32168 | n32174 ;
  assign n32176 = x792 & n32175 ;
  assign n32177 = n32163 & ~n32176 ;
  assign n32178 = ( x207 & x623 ) | ( x207 & n32177 ) | ( x623 & n32177 ) ;
  assign n32179 = ~n32086 & n32178 ;
  assign n32180 = x710 & ~n32179 ;
  assign n32181 = ( ~x1156 & n32169 ) | ( ~x1156 & n32172 ) | ( n32169 & n32172 ) ;
  assign n32182 = n32164 & n32167 ;
  assign n32183 = ( x1156 & n32172 ) | ( x1156 & ~n32182 ) | ( n32172 & ~n32182 ) ;
  assign n32184 = n32181 | n32183 ;
  assign n32185 = x792 & n32184 ;
  assign n32186 = x1158 | n32155 ;
  assign n32187 = ( x626 & x641 ) | ( x626 & n31961 ) | ( x641 & n31961 ) ;
  assign n32188 = ( x648 & x1159 ) | ( x648 & ~n14834 ) | ( x1159 & ~n14834 ) ;
  assign n32189 = ( x627 & x1154 ) | ( x627 & ~n14834 ) | ( x1154 & ~n14834 ) ;
  assign n32190 = ( x660 & x1155 ) | ( x660 & ~n14834 ) | ( x1155 & ~n14834 ) ;
  assign n32191 = ~n2032 & n17579 ;
  assign n32192 = x778 | n32191 ;
  assign n32193 = x625 & ~n32191 ;
  assign n32194 = n31943 & ~n32193 ;
  assign n32195 = x1153 & ~n32194 ;
  assign n32196 = n32097 & ~n32195 ;
  assign n32197 = x625 | n32191 ;
  assign n32198 = ~n31947 & n32197 ;
  assign n32199 = x1153 | n32198 ;
  assign n32200 = ~n32092 & n32199 ;
  assign n32201 = x778 & ~n32200 ;
  assign n32202 = ~n32196 & n32201 ;
  assign n32203 = n32192 & ~n32202 ;
  assign n32204 = x609 | n32203 ;
  assign n32205 = ~n32089 & n32204 ;
  assign n32206 = ( ~x660 & x1155 ) | ( ~x660 & n32205 ) | ( x1155 & n32205 ) ;
  assign n32207 = ~n32190 & n32206 ;
  assign n32208 = x609 & ~n32203 ;
  assign n32209 = n32110 & ~n32208 ;
  assign n32210 = ( x660 & ~x1155 ) | ( x660 & n32209 ) | ( ~x1155 & n32209 ) ;
  assign n32211 = ( x660 & x1155 ) | ( x660 & n14834 ) | ( x1155 & n14834 ) ;
  assign n32212 = n32210 & n32211 ;
  assign n32213 = n32207 | n32212 ;
  assign n32214 = x785 & n32213 ;
  assign n32215 = ~x785 & n32203 ;
  assign n32216 = n32214 | n32215 ;
  assign n32217 = x618 | n32216 ;
  assign n32218 = ~n32088 & n32217 ;
  assign n32219 = ( ~x627 & x1154 ) | ( ~x627 & n32218 ) | ( x1154 & n32218 ) ;
  assign n32220 = ~n32189 & n32219 ;
  assign n32221 = x618 & ~n32216 ;
  assign n32222 = n32125 & ~n32221 ;
  assign n32223 = ( x627 & ~x1154 ) | ( x627 & n32222 ) | ( ~x1154 & n32222 ) ;
  assign n32224 = ( x627 & x1154 ) | ( x627 & n14834 ) | ( x1154 & n14834 ) ;
  assign n32225 = n32223 & n32224 ;
  assign n32226 = n32220 | n32225 ;
  assign n32227 = x781 & n32226 ;
  assign n32228 = ~x781 & n32216 ;
  assign n32229 = n32227 | n32228 ;
  assign n32230 = x619 | n32229 ;
  assign n32231 = ~n32140 & n32230 ;
  assign n32232 = ( ~x648 & x1159 ) | ( ~x648 & n32231 ) | ( x1159 & n32231 ) ;
  assign n32233 = ~n32188 & n32232 ;
  assign n32234 = x619 & ~n32229 ;
  assign n32235 = n32087 & ~n32234 ;
  assign n32236 = ( x648 & ~x1159 ) | ( x648 & n32235 ) | ( ~x1159 & n32235 ) ;
  assign n32237 = ( x648 & x1159 ) | ( x648 & n14834 ) | ( x1159 & n14834 ) ;
  assign n32238 = n32236 & n32237 ;
  assign n32239 = n32233 | n32238 ;
  assign n32240 = x789 & n32239 ;
  assign n32241 = ~x789 & n32229 ;
  assign n32242 = n32240 | n32241 ;
  assign n32243 = ( ~x626 & x641 ) | ( ~x626 & n32242 ) | ( x641 & n32242 ) ;
  assign n32244 = n32187 | n32243 ;
  assign n32245 = ~n32186 & n32244 ;
  assign n32246 = x1158 & n32153 ;
  assign n32247 = ( x626 & x641 ) | ( x626 & ~n31961 ) | ( x641 & ~n31961 ) ;
  assign n32248 = ( x626 & ~x641 ) | ( x626 & n32242 ) | ( ~x641 & n32242 ) ;
  assign n32249 = n32247 & ~n32248 ;
  assign n32250 = n32246 & ~n32249 ;
  assign n32251 = n32245 | n32250 ;
  assign n32252 = ( x788 & n18434 ) | ( x788 & n32251 ) | ( n18434 & n32251 ) ;
  assign n32253 = ( ~x788 & n18434 ) | ( ~x788 & n32242 ) | ( n18434 & n32242 ) ;
  assign n32254 = n32252 | n32253 ;
  assign n32255 = ~n32185 & n32254 ;
  assign n32256 = ( x207 & ~x623 ) | ( x207 & n32255 ) | ( ~x623 & n32255 ) ;
  assign n32257 = n15397 | n32036 ;
  assign n32258 = x778 | n31182 ;
  assign n32259 = x625 & n31182 ;
  assign n32260 = x1153 & ~n32259 ;
  assign n32261 = n32019 & ~n32260 ;
  assign n32262 = ~x625 & n31182 ;
  assign n32263 = x1153 | n32262 ;
  assign n32264 = ~n32026 & n32263 ;
  assign n32265 = x778 & ~n32264 ;
  assign n32266 = ~n32261 & n32265 ;
  assign n32267 = n32258 & ~n32266 ;
  assign n32268 = n15398 & n32043 ;
  assign n32269 = ( ~x609 & n32267 ) | ( ~x609 & n32268 ) | ( n32267 & n32268 ) ;
  assign n32270 = x609 | n32268 ;
  assign n32271 = ( ~n32257 & n32269 ) | ( ~n32257 & n32270 ) | ( n32269 & n32270 ) ;
  assign n32272 = x785 & n32271 ;
  assign n32273 = ~x785 & n32267 ;
  assign n32274 = n32272 | n32273 ;
  assign n32275 = x618 & ~n32274 ;
  assign n32276 = n15405 & n32053 ;
  assign n32277 = ~n32275 & n32276 ;
  assign n32278 = x618 | n32274 ;
  assign n32279 = n15404 | n32011 ;
  assign n32280 = n32278 & ~n32279 ;
  assign n32281 = x781 & ~n32280 ;
  assign n32282 = ~n32277 & n32281 ;
  assign n32283 = x781 | n32274 ;
  assign n32284 = ~n21647 & n32283 ;
  assign n32285 = ~n32282 & n32284 ;
  assign n32286 = ~n15413 & n18253 ;
  assign n32287 = n31995 & n32286 ;
  assign n32288 = n32285 | n32287 ;
  assign n32289 = x626 & ~n32288 ;
  assign n32290 = x1158 & n32075 ;
  assign n32291 = ~n32289 & n32290 ;
  assign n32292 = x626 | n32288 ;
  assign n32293 = x1158 | n31998 ;
  assign n32294 = n32292 & ~n32293 ;
  assign n32295 = x788 & ~n32294 ;
  assign n32296 = ~n32291 & n32295 ;
  assign n32297 = x788 | n32288 ;
  assign n32298 = ~n18434 & n32297 ;
  assign n32299 = ~n32296 & n32298 ;
  assign n32300 = n15134 & ~n16053 ;
  assign n32301 = n31937 & n32300 ;
  assign n32302 = n32299 | n32301 ;
  assign n32303 = ( x207 & x623 ) | ( x207 & n32302 ) | ( x623 & n32302 ) ;
  assign n32304 = n32256 & ~n32303 ;
  assign n32305 = n32180 & ~n32304 ;
  assign n32306 = x710 | n31928 ;
  assign n32307 = ~n18431 & n32306 ;
  assign n32308 = ~n32305 & n32307 ;
  assign n32309 = n31986 | n32308 ;
  assign n32310 = ( ~x644 & x715 ) | ( ~x644 & n32309 ) | ( x715 & n32309 ) ;
  assign n32311 = n31981 & n32310 ;
  assign n32312 = n31934 & ~n32311 ;
  assign n32313 = ( x644 & x715 ) | ( x644 & n31930 ) | ( x715 & n31930 ) ;
  assign n32314 = ( ~x644 & x715 ) | ( ~x644 & n31873 ) | ( x715 & n31873 ) ;
  assign n32315 = n32313 & n32314 ;
  assign n32316 = x1160 | n32315 ;
  assign n32317 = ( x644 & x715 ) | ( x644 & ~n31980 ) | ( x715 & ~n31980 ) ;
  assign n32318 = ( x644 & ~x715 ) | ( x644 & n32309 ) | ( ~x715 & n32309 ) ;
  assign n32319 = ~n32317 & n32318 ;
  assign n32320 = n32316 | n32319 ;
  assign n32321 = ~n32312 & n32320 ;
  assign n32322 = ( x790 & n6785 ) | ( x790 & n32321 ) | ( n6785 & n32321 ) ;
  assign n32323 = ( ~x790 & n6785 ) | ( ~x790 & n32309 ) | ( n6785 & n32309 ) ;
  assign n32324 = n32322 | n32323 ;
  assign n32325 = ~n31872 & n32324 ;
  assign n32326 = ~x208 & n6785 ;
  assign n32327 = x208 | n14834 ;
  assign n32328 = n15141 & n32327 ;
  assign n32329 = x607 | n32327 ;
  assign n32330 = ( ~x208 & x607 ) | ( ~x208 & n31882 ) | ( x607 & n31882 ) ;
  assign n32331 = ( x208 & x607 ) | ( x208 & ~n31925 ) | ( x607 & ~n31925 ) ;
  assign n32332 = n32330 & n32331 ;
  assign n32333 = n32329 & ~n32332 ;
  assign n32334 = ~n15141 & n32333 ;
  assign n32335 = n32328 | n32334 ;
  assign n32336 = ( x644 & x715 ) | ( x644 & ~n32335 ) | ( x715 & ~n32335 ) ;
  assign n32337 = ( x644 & ~x715 ) | ( x644 & n32327 ) | ( ~x715 & n32327 ) ;
  assign n32338 = ~n32336 & n32337 ;
  assign n32339 = x1160 & ~n32338 ;
  assign n32340 = ~x638 & n32327 ;
  assign n32341 = ( x208 & ~x638 ) | ( x208 & n31938 ) | ( ~x638 & n31938 ) ;
  assign n32342 = ( x208 & x638 ) | ( x208 & n31967 ) | ( x638 & n31967 ) ;
  assign n32343 = ~n32341 & n32342 ;
  assign n32344 = n32340 | n32343 ;
  assign n32345 = ~x787 & n32344 ;
  assign n32346 = ( x647 & x1157 ) | ( x647 & ~n32327 ) | ( x1157 & ~n32327 ) ;
  assign n32347 = ( x647 & ~x1157 ) | ( x647 & n32344 ) | ( ~x1157 & n32344 ) ;
  assign n32348 = ~n32346 & n32347 ;
  assign n32349 = ( x647 & x1157 ) | ( x647 & n32327 ) | ( x1157 & n32327 ) ;
  assign n32350 = ( ~x647 & x1157 ) | ( ~x647 & n32344 ) | ( x1157 & n32344 ) ;
  assign n32351 = n32349 & n32350 ;
  assign n32352 = n32348 | n32351 ;
  assign n32353 = x787 & n32352 ;
  assign n32354 = n32345 | n32353 ;
  assign n32355 = ( x644 & x715 ) | ( x644 & n32354 ) | ( x715 & n32354 ) ;
  assign n32356 = n18610 & n32333 ;
  assign n32357 = ( x630 & n32348 ) | ( x630 & n32356 ) | ( n32348 & n32356 ) ;
  assign n32358 = ( ~x630 & n32351 ) | ( ~x630 & n32356 ) | ( n32351 & n32356 ) ;
  assign n32359 = n32357 | n32358 ;
  assign n32360 = x787 & n32359 ;
  assign n32361 = ( x208 & ~x607 ) | ( x208 & n32085 ) | ( ~x607 & n32085 ) ;
  assign n32362 = ( x208 & x607 ) | ( x208 & n32177 ) | ( x607 & n32177 ) ;
  assign n32363 = ~n32361 & n32362 ;
  assign n32364 = x638 & ~n32363 ;
  assign n32365 = ( x208 & ~x607 ) | ( x208 & n32255 ) | ( ~x607 & n32255 ) ;
  assign n32366 = ( x208 & x607 ) | ( x208 & n32302 ) | ( x607 & n32302 ) ;
  assign n32367 = n32365 & ~n32366 ;
  assign n32368 = n32364 & ~n32367 ;
  assign n32369 = x638 | n32333 ;
  assign n32370 = ~n18431 & n32369 ;
  assign n32371 = ~n32368 & n32370 ;
  assign n32372 = n32360 | n32371 ;
  assign n32373 = ( ~x644 & x715 ) | ( ~x644 & n32372 ) | ( x715 & n32372 ) ;
  assign n32374 = n32355 & n32373 ;
  assign n32375 = n32339 & ~n32374 ;
  assign n32376 = ( x644 & x715 ) | ( x644 & n32335 ) | ( x715 & n32335 ) ;
  assign n32377 = ( ~x644 & x715 ) | ( ~x644 & n32327 ) | ( x715 & n32327 ) ;
  assign n32378 = n32376 & n32377 ;
  assign n32379 = x1160 | n32378 ;
  assign n32380 = ( x644 & x715 ) | ( x644 & ~n32354 ) | ( x715 & ~n32354 ) ;
  assign n32381 = ( x644 & ~x715 ) | ( x644 & n32372 ) | ( ~x715 & n32372 ) ;
  assign n32382 = ~n32380 & n32381 ;
  assign n32383 = n32379 | n32382 ;
  assign n32384 = ~n32375 & n32383 ;
  assign n32385 = ( x790 & n6785 ) | ( x790 & n32384 ) | ( n6785 & n32384 ) ;
  assign n32386 = ( ~x790 & n6785 ) | ( ~x790 & n32372 ) | ( n6785 & n32372 ) ;
  assign n32387 = n32385 | n32386 ;
  assign n32388 = ~n32326 & n32387 ;
  assign n32389 = n18431 | n32177 ;
  assign n32390 = x647 | n14834 ;
  assign n32391 = x647 & ~n31967 ;
  assign n32392 = n32390 & ~n32391 ;
  assign n32393 = x630 | n32392 ;
  assign n32394 = x1157 & ~n32393 ;
  assign n32395 = x647 & ~n14834 ;
  assign n32396 = x647 | n31967 ;
  assign n32397 = ~n32395 & n32396 ;
  assign n32398 = n15139 & ~n32397 ;
  assign n32399 = n18610 & ~n31925 ;
  assign n32400 = n32398 | n32399 ;
  assign n32401 = n32394 | n32400 ;
  assign n32402 = x787 & n32401 ;
  assign n32403 = n32389 & ~n32402 ;
  assign n32404 = ( x790 & ~n6785 ) | ( x790 & n32403 ) | ( ~n6785 & n32403 ) ;
  assign n32405 = n17389 | n31967 ;
  assign n32406 = ~n14834 & n17389 ;
  assign n32407 = n32405 & ~n32406 ;
  assign n32408 = x644 & ~n32407 ;
  assign n32409 = x715 | n32408 ;
  assign n32410 = x644 | n32403 ;
  assign n32411 = ~n32409 & n32410 ;
  assign n32412 = ~n14834 & n15141 ;
  assign n32413 = n15141 | n31925 ;
  assign n32414 = ~n32412 & n32413 ;
  assign n32415 = x644 | n32414 ;
  assign n32416 = x644 & ~n14834 ;
  assign n32417 = n32415 & ~n32416 ;
  assign n32418 = x715 & n32417 ;
  assign n32419 = x1160 | n32418 ;
  assign n32420 = n32411 | n32419 ;
  assign n32421 = x644 | n32407 ;
  assign n32422 = x715 & n32421 ;
  assign n32423 = x644 & ~n32403 ;
  assign n32424 = n32422 & ~n32423 ;
  assign n32425 = x644 & ~n32414 ;
  assign n32426 = x644 | n14834 ;
  assign n32427 = ~n32425 & n32426 ;
  assign n32428 = ~x715 & n32427 ;
  assign n32429 = x1160 & ~n32428 ;
  assign n32430 = ~n32424 & n32429 ;
  assign n32431 = n32420 & ~n32430 ;
  assign n32432 = ( x790 & n6785 ) | ( x790 & ~n32431 ) | ( n6785 & ~n32431 ) ;
  assign n32433 = n32404 & ~n32432 ;
  assign n32434 = x639 & n32433 ;
  assign n32435 = x790 | n32414 ;
  assign n32436 = ~n6785 & n32435 ;
  assign n32437 = ( ~x790 & x1160 ) | ( ~x790 & n32427 ) | ( x1160 & n32427 ) ;
  assign n32438 = ( x790 & x1160 ) | ( x790 & ~n32417 ) | ( x1160 & ~n32417 ) ;
  assign n32439 = ~n32437 & n32438 ;
  assign n32440 = n32436 & ~n32439 ;
  assign n32441 = x622 & x639 ;
  assign n32442 = ( x622 & ~n32440 ) | ( x622 & n32441 ) | ( ~n32440 & n32441 ) ;
  assign n32443 = ~n32434 & n32442 ;
  assign n32444 = n18431 | n32255 ;
  assign n32445 = ( ~x1157 & n32395 ) | ( ~x1157 & n32398 ) | ( n32395 & n32398 ) ;
  assign n32446 = n32390 & n32393 ;
  assign n32447 = ( x1157 & n32398 ) | ( x1157 & ~n32446 ) | ( n32398 & ~n32446 ) ;
  assign n32448 = n32445 | n32447 ;
  assign n32449 = x787 & n32448 ;
  assign n32450 = n32444 & ~n32449 ;
  assign n32451 = ( x790 & ~n6785 ) | ( x790 & n32450 ) | ( ~n6785 & n32450 ) ;
  assign n32452 = x644 | n32450 ;
  assign n32453 = ~n32409 & n32452 ;
  assign n32454 = x715 & n14834 ;
  assign n32455 = x1160 | n32454 ;
  assign n32456 = n32453 | n32455 ;
  assign n32457 = x644 & ~n32450 ;
  assign n32458 = n32422 & ~n32457 ;
  assign n32459 = ~x715 & n14834 ;
  assign n32460 = x1160 & ~n32459 ;
  assign n32461 = ~n32458 & n32460 ;
  assign n32462 = n32456 & ~n32461 ;
  assign n32463 = ( x790 & n6785 ) | ( x790 & ~n32462 ) | ( n6785 & ~n32462 ) ;
  assign n32464 = n32451 & ~n32463 ;
  assign n32465 = ( x622 & x639 ) | ( x622 & n32464 ) | ( x639 & n32464 ) ;
  assign n32466 = ~n8359 & n15382 ;
  assign n32467 = ( x622 & ~x639 ) | ( x622 & n32466 ) | ( ~x639 & n32466 ) ;
  assign n32468 = n32465 | n32467 ;
  assign n32469 = ~n32443 & n32468 ;
  assign n32470 = x209 | n32469 ;
  assign n32471 = x647 & n31938 ;
  assign n32472 = x1157 & ~n32471 ;
  assign n32473 = x630 | n32472 ;
  assign n32474 = ( x647 & x1157 ) | ( x647 & n31882 ) | ( x1157 & n31882 ) ;
  assign n32475 = ( ~x647 & x1157 ) | ( ~x647 & n32085 ) | ( x1157 & n32085 ) ;
  assign n32476 = n32474 | n32475 ;
  assign n32477 = ~n32473 & n32476 ;
  assign n32478 = ~x647 & n31938 ;
  assign n32479 = x1157 | n32478 ;
  assign n32480 = x630 & n32479 ;
  assign n32481 = ( x647 & x1157 ) | ( x647 & ~n31882 ) | ( x1157 & ~n31882 ) ;
  assign n32482 = ( x647 & ~x1157 ) | ( x647 & n32085 ) | ( ~x1157 & n32085 ) ;
  assign n32483 = n32481 & ~n32482 ;
  assign n32484 = n32480 & ~n32483 ;
  assign n32485 = n32477 | n32484 ;
  assign n32486 = x787 & n32485 ;
  assign n32487 = ~x787 & n32085 ;
  assign n32488 = n32486 | n32487 ;
  assign n32489 = ( x790 & ~n6785 ) | ( x790 & n32488 ) | ( ~n6785 & n32488 ) ;
  assign n32490 = ~n17389 & n31938 ;
  assign n32491 = x644 & ~n32490 ;
  assign n32492 = x715 | n32491 ;
  assign n32493 = x644 | n32488 ;
  assign n32494 = ~n32492 & n32493 ;
  assign n32495 = ~n18264 & n31881 ;
  assign n32496 = n21195 & n32495 ;
  assign n32497 = x1160 | n32496 ;
  assign n32498 = n32494 | n32497 ;
  assign n32499 = x644 | n32490 ;
  assign n32500 = x715 & n32499 ;
  assign n32501 = x644 & ~n32488 ;
  assign n32502 = n32500 & ~n32501 ;
  assign n32503 = n21513 & n32495 ;
  assign n32504 = x1160 & ~n32503 ;
  assign n32505 = ~n32502 & n32504 ;
  assign n32506 = n32498 & ~n32505 ;
  assign n32507 = ( x790 & n6785 ) | ( x790 & ~n32506 ) | ( n6785 & ~n32506 ) ;
  assign n32508 = n32489 & ~n32507 ;
  assign n32509 = n32441 & ~n32508 ;
  assign n32510 = ~n18431 & n32302 ;
  assign n32511 = n15141 & ~n17388 ;
  assign n32512 = n31938 & n32511 ;
  assign n32513 = n32510 | n32512 ;
  assign n32514 = x644 | n32513 ;
  assign n32515 = x1160 | n32492 ;
  assign n32516 = n32514 & ~n32515 ;
  assign n32517 = x644 & ~n32513 ;
  assign n32518 = x1160 & n32500 ;
  assign n32519 = ~n32517 & n32518 ;
  assign n32520 = x790 & ~n32519 ;
  assign n32521 = ~n32516 & n32520 ;
  assign n32522 = x790 | n32513 ;
  assign n32523 = ~n6785 & n32522 ;
  assign n32524 = ~n32521 & n32523 ;
  assign n32525 = x622 | n32524 ;
  assign n32526 = ~x644 & x1160 ;
  assign n32527 = ( x790 & ~x1160 ) | ( x790 & n32526 ) | ( ~x1160 & n32526 ) ;
  assign n32528 = ( x644 & n32526 ) | ( x644 & n32527 ) | ( n32526 & n32527 ) ;
  assign n32529 = n6785 | n32528 ;
  assign n32530 = n32495 & ~n32529 ;
  assign n32531 = x622 & n32530 ;
  assign n32532 = x639 | n32531 ;
  assign n32533 = x209 & n32532 ;
  assign n32534 = n32525 & n32533 ;
  assign n32535 = ~n32509 & n32534 ;
  assign n32536 = n32470 & ~n32535 ;
  assign n32537 = x210 & ~n16705 ;
  assign n32538 = ~n4712 & n32537 ;
  assign n32539 = x210 & n4712 ;
  assign n32540 = ~n30485 & n32539 ;
  assign n32541 = n32538 | n32540 ;
  assign n32542 = x907 | n32541 ;
  assign n32543 = x634 & n16705 ;
  assign n32544 = n32537 | n32543 ;
  assign n32545 = ~n4714 & n32544 ;
  assign n32546 = x907 & ~n32545 ;
  assign n32547 = x210 & ~n14475 ;
  assign n32548 = n30707 | n32547 ;
  assign n32549 = n4714 & n32548 ;
  assign n32550 = n32546 & ~n32549 ;
  assign n32551 = x947 | n32550 ;
  assign n32552 = n32542 & ~n32551 ;
  assign n32553 = n30532 | n32537 ;
  assign n32554 = n4712 | n32553 ;
  assign n32555 = x947 & n32554 ;
  assign n32556 = n4712 & ~n32553 ;
  assign n32557 = n4714 | n32556 ;
  assign n32558 = x633 & n14475 ;
  assign n32559 = n32547 | n32558 ;
  assign n32560 = n4713 & n32559 ;
  assign n32561 = n32557 & ~n32560 ;
  assign n32562 = n32555 & ~n32561 ;
  assign n32563 = n4764 | n32562 ;
  assign n32564 = n32552 | n32563 ;
  assign n32565 = n4751 & ~n32544 ;
  assign n32566 = x907 & ~n32565 ;
  assign n32567 = n4751 | n32548 ;
  assign n32568 = n32566 & n32567 ;
  assign n32569 = n4751 & ~n14481 ;
  assign n32570 = n1290 & n32569 ;
  assign n32571 = n32547 & ~n32570 ;
  assign n32572 = n32568 | n32571 ;
  assign n32573 = ~x947 & n32572 ;
  assign n32574 = n4751 & ~n32553 ;
  assign n32575 = x947 & ~n32574 ;
  assign n32576 = n4751 | n32559 ;
  assign n32577 = n32575 & n32576 ;
  assign n32578 = n32573 | n32577 ;
  assign n32579 = ( x223 & n15044 ) | ( x223 & n32578 ) | ( n15044 & n32578 ) ;
  assign n32580 = n32564 & n32579 ;
  assign n32581 = x299 | n32580 ;
  assign n32582 = ~n14641 & n32539 ;
  assign n32583 = n32538 | n32582 ;
  assign n32584 = x907 | n32583 ;
  assign n32585 = x210 & ~n30540 ;
  assign n32586 = x634 & n30540 ;
  assign n32587 = n32585 | n32586 ;
  assign n32588 = n4714 & n32587 ;
  assign n32589 = n32546 & ~n32588 ;
  assign n32590 = x947 | n32589 ;
  assign n32591 = n32584 & ~n32590 ;
  assign n32592 = x633 & n30540 ;
  assign n32593 = n32585 | n32592 ;
  assign n32594 = n4713 & n32593 ;
  assign n32595 = n32557 & ~n32594 ;
  assign n32596 = n32555 & ~n32595 ;
  assign n32597 = n4764 | n32596 ;
  assign n32598 = n32591 | n32597 ;
  assign n32599 = n4751 | n32587 ;
  assign n32600 = n32566 & n32599 ;
  assign n32601 = x210 & ~n14997 ;
  assign n32602 = ~x907 & n32601 ;
  assign n32603 = n32600 | n32602 ;
  assign n32604 = ~x947 & n32603 ;
  assign n32605 = n4751 | n32593 ;
  assign n32606 = n32575 & n32605 ;
  assign n32607 = n4764 & ~n32606 ;
  assign n32608 = ~n32604 & n32607 ;
  assign n32609 = n32598 & ~n32608 ;
  assign n32610 = ( x223 & n1823 ) | ( x223 & ~n32609 ) | ( n1823 & ~n32609 ) ;
  assign n32611 = x634 & n18913 ;
  assign n32612 = x633 & x947 ;
  assign n32613 = n32611 | n32612 ;
  assign n32614 = n16705 & n32613 ;
  assign n32615 = n32537 | n32614 ;
  assign n32616 = ( ~x223 & n1823 ) | ( ~x223 & n32615 ) | ( n1823 & n32615 ) ;
  assign n32617 = ~n32610 & n32616 ;
  assign n32618 = n32581 | n32617 ;
  assign n32619 = ( x907 & n14450 ) | ( x907 & ~n32601 ) | ( n14450 & ~n32601 ) ;
  assign n32620 = ( ~x907 & n14450 ) | ( ~x907 & n32583 ) | ( n14450 & n32583 ) ;
  assign n32621 = ~n32619 & n32620 ;
  assign n32622 = n32600 | n32621 ;
  assign n32623 = ~x947 & n32622 ;
  assign n32624 = n2203 & ~n32606 ;
  assign n32625 = ~n32623 & n32624 ;
  assign n32626 = ( ~x215 & n14841 ) | ( ~x215 & n32615 ) | ( n14841 & n32615 ) ;
  assign n32627 = ~n32625 & n32626 ;
  assign n32628 = ( x907 & n14450 ) | ( x907 & ~n32571 ) | ( n14450 & ~n32571 ) ;
  assign n32629 = ( ~x907 & n14450 ) | ( ~x907 & n32541 ) | ( n14450 & n32541 ) ;
  assign n32630 = ~n32628 & n32629 ;
  assign n32631 = n32568 | n32630 ;
  assign n32632 = ~x947 & n32631 ;
  assign n32633 = n32577 | n32632 ;
  assign n32634 = x215 & n32633 ;
  assign n32635 = x299 & ~n32634 ;
  assign n32636 = ~n32627 & n32635 ;
  assign n32637 = x39 & ~n32636 ;
  assign n32638 = n32618 & n32637 ;
  assign n32639 = n14784 & n32613 ;
  assign n32640 = x299 & ~n32639 ;
  assign n32641 = ~n14813 & n32640 ;
  assign n32642 = ( x299 & n14820 ) | ( x299 & n32613 ) | ( n14820 & n32613 ) ;
  assign n32643 = ( x210 & x299 ) | ( x210 & ~n14820 ) | ( x299 & ~n14820 ) ;
  assign n32644 = n32642 | n32643 ;
  assign n32645 = ~n32641 & n32644 ;
  assign n32646 = ( x38 & ~n9138 ) | ( x38 & n32645 ) | ( ~n9138 & n32645 ) ;
  assign n32647 = n32638 | n32646 ;
  assign n32648 = ( ~x38 & n15070 ) | ( ~x38 & n32613 ) | ( n15070 & n32613 ) ;
  assign n32649 = ( x38 & ~x210 ) | ( x38 & n15070 ) | ( ~x210 & n15070 ) ;
  assign n32650 = ~n32648 & n32649 ;
  assign n32651 = n32647 & ~n32650 ;
  assign n32652 = n8359 | n32651 ;
  assign n32653 = ~x210 & n8359 ;
  assign n32654 = n32652 & ~n32653 ;
  assign n32655 = ~n2032 & n19010 ;
  assign n32656 = ( x606 & x643 ) | ( x606 & n32655 ) | ( x643 & n32655 ) ;
  assign n32657 = ( ~x606 & x643 ) | ( ~x606 & n14834 ) | ( x643 & n14834 ) ;
  assign n32658 = n32656 | n32657 ;
  assign n32659 = ~n6785 & n32658 ;
  assign n32660 = ~n2032 & n19623 ;
  assign n32661 = ( x606 & x643 ) | ( x606 & ~n32660 ) | ( x643 & ~n32660 ) ;
  assign n32662 = ~n2032 & n19627 ;
  assign n32663 = ( x606 & ~x643 ) | ( x606 & n32662 ) | ( ~x643 & n32662 ) ;
  assign n32664 = n32661 & ~n32663 ;
  assign n32665 = n32659 & ~n32664 ;
  assign n32666 = x211 & ~n32665 ;
  assign n32667 = ~n2032 & n19034 ;
  assign n32668 = x606 & ~x643 ;
  assign n32669 = n32667 & n32668 ;
  assign n32670 = ~n2032 & n19609 ;
  assign n32671 = ( x606 & x643 ) | ( x606 & n32670 ) | ( x643 & n32670 ) ;
  assign n32672 = ~n2032 & n19612 ;
  assign n32673 = ( ~x606 & x643 ) | ( ~x606 & n32672 ) | ( x643 & n32672 ) ;
  assign n32674 = n32671 & n32673 ;
  assign n32675 = n32669 | n32674 ;
  assign n32676 = x211 | n6785 ;
  assign n32677 = n32675 & ~n32676 ;
  assign n32678 = n32666 | n32677 ;
  assign n32679 = ( x607 & x638 ) | ( x607 & n32655 ) | ( x638 & n32655 ) ;
  assign n32680 = ( ~x607 & x638 ) | ( ~x607 & n14834 ) | ( x638 & n14834 ) ;
  assign n32681 = n32679 | n32680 ;
  assign n32682 = ~n6785 & n32681 ;
  assign n32683 = ( x607 & x638 ) | ( x607 & ~n32660 ) | ( x638 & ~n32660 ) ;
  assign n32684 = ( x607 & ~x638 ) | ( x607 & n32662 ) | ( ~x638 & n32662 ) ;
  assign n32685 = n32683 & ~n32684 ;
  assign n32686 = n32682 & ~n32685 ;
  assign n32687 = x212 | n32686 ;
  assign n32688 = x607 & ~x638 ;
  assign n32689 = n32667 & n32688 ;
  assign n32690 = ( x607 & x638 ) | ( x607 & n32670 ) | ( x638 & n32670 ) ;
  assign n32691 = ( ~x607 & x638 ) | ( ~x607 & n32672 ) | ( x638 & n32672 ) ;
  assign n32692 = n32690 & n32691 ;
  assign n32693 = n32689 | n32692 ;
  assign n32694 = x212 & ~n6785 ;
  assign n32695 = n32693 & n32694 ;
  assign n32696 = n32687 & ~n32695 ;
  assign n32697 = x213 & ~n6785 ;
  assign n32698 = x622 & ~x639 ;
  assign n32699 = n32667 & n32698 ;
  assign n32700 = ( x622 & x639 ) | ( x622 & n32670 ) | ( x639 & n32670 ) ;
  assign n32701 = ( ~x622 & x639 ) | ( ~x622 & n32672 ) | ( x639 & n32672 ) ;
  assign n32702 = n32700 & n32701 ;
  assign n32703 = n32699 | n32702 ;
  assign n32704 = n32697 & n32703 ;
  assign n32705 = x639 & n32662 ;
  assign n32706 = ( x622 & n32441 ) | ( x622 & ~n32655 ) | ( n32441 & ~n32655 ) ;
  assign n32707 = ~n32705 & n32706 ;
  assign n32708 = ( x622 & x639 ) | ( x622 & n32660 ) | ( x639 & n32660 ) ;
  assign n32709 = ( x622 & ~x639 ) | ( x622 & n14834 ) | ( ~x639 & n14834 ) ;
  assign n32710 = n32708 | n32709 ;
  assign n32711 = ~n6785 & n32710 ;
  assign n32712 = ~n32707 & n32711 ;
  assign n32713 = x213 | n32712 ;
  assign n32714 = ~n32704 & n32713 ;
  assign n32715 = ( x623 & x710 ) | ( x623 & n32655 ) | ( x710 & n32655 ) ;
  assign n32716 = ( ~x623 & x710 ) | ( ~x623 & n14834 ) | ( x710 & n14834 ) ;
  assign n32717 = n32715 | n32716 ;
  assign n32718 = ~n6785 & n32717 ;
  assign n32719 = ( x623 & x710 ) | ( x623 & ~n32660 ) | ( x710 & ~n32660 ) ;
  assign n32720 = ( x623 & ~x710 ) | ( x623 & n32662 ) | ( ~x710 & n32662 ) ;
  assign n32721 = n32719 & ~n32720 ;
  assign n32722 = n32718 & ~n32721 ;
  assign n32723 = x214 | n32722 ;
  assign n32724 = x623 & ~x710 ;
  assign n32725 = n32667 & n32724 ;
  assign n32726 = ( x623 & x710 ) | ( x623 & n32670 ) | ( x710 & n32670 ) ;
  assign n32727 = ( ~x623 & x710 ) | ( ~x623 & n32672 ) | ( x710 & n32672 ) ;
  assign n32728 = n32726 & n32727 ;
  assign n32729 = n32725 | n32728 ;
  assign n32730 = x214 & ~n6785 ;
  assign n32731 = n32729 & n32730 ;
  assign n32732 = n32723 & ~n32731 ;
  assign n32733 = x215 & n8359 ;
  assign n32734 = x947 | n19310 ;
  assign n32735 = x681 & x907 ;
  assign n32736 = ~x947 & n32735 ;
  assign n32737 = ( n14515 & n14519 ) | ( n14515 & n14521 ) | ( n14519 & n14521 ) ;
  assign n32738 = n4711 | n32737 ;
  assign n32739 = ~n4710 & n14507 ;
  assign n32740 = x642 | n32739 ;
  assign n32741 = n32738 & ~n32740 ;
  assign n32742 = x947 & ~n32741 ;
  assign n32743 = n32736 | n32742 ;
  assign n32744 = n32734 & ~n32743 ;
  assign n32745 = x299 & ~n32744 ;
  assign n32746 = n19384 & ~n32735 ;
  assign n32747 = ~x642 & n14997 ;
  assign n32748 = ( x947 & ~n4764 ) | ( x947 & n32747 ) | ( ~n4764 & n32747 ) ;
  assign n32749 = ~x642 & n14641 ;
  assign n32750 = n4711 & ~n32749 ;
  assign n32751 = ( ~n14624 & n14647 ) | ( ~n14624 & n14650 ) | ( n14647 & n14650 ) ;
  assign n32752 = ~n14855 & n32751 ;
  assign n32753 = n4707 & n16705 ;
  assign n32754 = ~x642 & n32753 ;
  assign n32755 = n4711 | n32754 ;
  assign n32756 = n32752 | n32755 ;
  assign n32757 = ~n32750 & n32756 ;
  assign n32758 = ( x947 & n4764 ) | ( x947 & n32757 ) | ( n4764 & n32757 ) ;
  assign n32759 = n32748 & n32758 ;
  assign n32760 = n1823 & ~n32759 ;
  assign n32761 = ~n32746 & n32760 ;
  assign n32762 = n1823 | n16705 ;
  assign n32763 = x642 & x947 ;
  assign n32764 = n32736 | n32763 ;
  assign n32765 = ~n1823 & n32764 ;
  assign n32766 = x223 | n32765 ;
  assign n32767 = n32762 & ~n32766 ;
  assign n32768 = ~n32761 & n32767 ;
  assign n32769 = ( x947 & ~n4764 ) | ( x947 & n32741 ) | ( ~n4764 & n32741 ) ;
  assign n32770 = n4711 | n14504 ;
  assign n32771 = n4711 & ~n30485 ;
  assign n32772 = x642 | n32771 ;
  assign n32773 = n32770 & ~n32772 ;
  assign n32774 = ( x947 & n4764 ) | ( x947 & n32773 ) | ( n4764 & n32773 ) ;
  assign n32775 = n32769 & n32774 ;
  assign n32776 = n19090 | n32775 ;
  assign n32777 = x223 & ~n32736 ;
  assign n32778 = n32776 & n32777 ;
  assign n32779 = x299 | n32778 ;
  assign n32780 = n32768 | n32779 ;
  assign n32781 = ~n32745 & n32780 ;
  assign n32782 = x215 & ~n32781 ;
  assign n32783 = n14678 & n32736 ;
  assign n32784 = x642 & n14553 ;
  assign n32785 = n16705 & n32784 ;
  assign n32786 = ( x680 & ~n14481 ) | ( x680 & n14544 ) | ( ~n14481 & n14544 ) ;
  assign n32787 = x642 & ~n14553 ;
  assign n32788 = n32786 & n32787 ;
  assign n32789 = ( x680 & n14533 ) | ( x680 & n14624 ) | ( n14533 & n14624 ) ;
  assign n32790 = n32788 & ~n32789 ;
  assign n32791 = n32785 | n32790 ;
  assign n32792 = x947 & n32791 ;
  assign n32793 = n4764 | n32792 ;
  assign n32794 = n32783 | n32793 ;
  assign n32795 = n4711 | n15503 ;
  assign n32796 = ~n14848 & n32795 ;
  assign n32797 = n32787 & n32796 ;
  assign n32798 = n15503 & n32784 ;
  assign n32799 = x947 & ~n32798 ;
  assign n32800 = ~n32797 & n32799 ;
  assign n32801 = n14614 & n32736 ;
  assign n32802 = ( x947 & ~n32800 ) | ( x947 & n32801 ) | ( ~n32800 & n32801 ) ;
  assign n32803 = n4764 & ~n32802 ;
  assign n32804 = n1823 & ~n32803 ;
  assign n32805 = n32794 & n32804 ;
  assign n32806 = n16705 & n32765 ;
  assign n32807 = x223 | n32806 ;
  assign n32808 = n32805 | n32807 ;
  assign n32809 = x947 & ~n14521 ;
  assign n32810 = ( x947 & n32737 ) | ( x947 & ~n32809 ) | ( n32737 & ~n32809 ) ;
  assign n32811 = n4764 & ~n32810 ;
  assign n32812 = ~n14534 & n32788 ;
  assign n32813 = x947 & ~n32785 ;
  assign n32814 = ~n32812 & n32813 ;
  assign n32815 = n32811 | n32814 ;
  assign n32816 = n4764 | n14504 ;
  assign n32817 = n32736 & n32816 ;
  assign n32818 = ( x947 & ~n32815 ) | ( x947 & n32817 ) | ( ~n32815 & n32817 ) ;
  assign n32819 = x223 & ~n32818 ;
  assign n32820 = n32808 & ~n32819 ;
  assign n32821 = x299 | n32820 ;
  assign n32822 = n2203 & n32802 ;
  assign n32823 = n18991 & n32764 ;
  assign n32824 = x299 & ~n32823 ;
  assign n32825 = ~n32822 & n32824 ;
  assign n32826 = x215 | n32825 ;
  assign n32827 = n32821 & ~n32826 ;
  assign n32828 = n32782 | n32827 ;
  assign n32829 = x39 & n32828 ;
  assign n32830 = ( x299 & n14820 ) | ( x299 & n32764 ) | ( n14820 & n32764 ) ;
  assign n32831 = ( x215 & x299 ) | ( x215 & ~n14820 ) | ( x299 & ~n14820 ) ;
  assign n32832 = n32830 | n32831 ;
  assign n32833 = ( ~x299 & n14814 ) | ( ~x299 & n32764 ) | ( n14814 & n32764 ) ;
  assign n32834 = ( ~x215 & x299 ) | ( ~x215 & n14814 ) | ( x299 & n14814 ) ;
  assign n32835 = ~n32833 & n32834 ;
  assign n32836 = n32832 & ~n32835 ;
  assign n32837 = ( x38 & ~n9138 ) | ( x38 & n32836 ) | ( ~n9138 & n32836 ) ;
  assign n32838 = n32829 | n32837 ;
  assign n32839 = ( ~x38 & n15070 ) | ( ~x38 & n32764 ) | ( n15070 & n32764 ) ;
  assign n32840 = ( x38 & ~x215 ) | ( x38 & n15070 ) | ( ~x215 & n15070 ) ;
  assign n32841 = ~n32839 & n32840 ;
  assign n32842 = n8359 | n32841 ;
  assign n32843 = n32838 & ~n32842 ;
  assign n32844 = n32733 | n32843 ;
  assign n32845 = x947 | n18994 ;
  assign n32846 = x662 & x907 ;
  assign n32847 = ~x947 & n32846 ;
  assign n32848 = ~x614 & n14997 ;
  assign n32849 = x947 & ~n32848 ;
  assign n32850 = n32847 | n32849 ;
  assign n32851 = n32845 & ~n32850 ;
  assign n32852 = x216 & ~n32851 ;
  assign n32853 = x614 & x947 ;
  assign n32854 = n32796 & n32853 ;
  assign n32855 = n14614 & n32847 ;
  assign n32856 = n32854 | n32855 ;
  assign n32857 = n4322 & n32856 ;
  assign n32858 = n32847 | n32853 ;
  assign n32859 = n18991 & n32858 ;
  assign n32860 = n32857 | n32859 ;
  assign n32861 = n32852 | n32860 ;
  assign n32862 = ~x215 & n32861 ;
  assign n32863 = n14495 | n30489 ;
  assign n32864 = n30488 | n32863 ;
  assign n32865 = ~n14653 & n32864 ;
  assign n32866 = ~x614 & n14475 ;
  assign n32867 = n4711 & n32866 ;
  assign n32868 = n32865 | n32867 ;
  assign n32869 = x947 & ~n32868 ;
  assign n32870 = x216 & ~n32847 ;
  assign n32871 = ~n32869 & n32870 ;
  assign n32872 = n32734 & n32871 ;
  assign n32873 = ~n14534 & n14632 ;
  assign n32874 = x947 & ~n14627 ;
  assign n32875 = ~n32873 & n32874 ;
  assign n32876 = ( x947 & ~n14521 ) | ( x947 & n32875 ) | ( ~n14521 & n32875 ) ;
  assign n32877 = n32737 & n32846 ;
  assign n32878 = ( x947 & ~n32875 ) | ( x947 & n32877 ) | ( ~n32875 & n32877 ) ;
  assign n32879 = ~n32876 & n32878 ;
  assign n32880 = x216 | n32879 ;
  assign n32881 = x215 & n32880 ;
  assign n32882 = ~n32872 & n32881 ;
  assign n32883 = x299 & ~n32882 ;
  assign n32884 = ~n32862 & n32883 ;
  assign n32885 = x947 & n14665 ;
  assign n32886 = ~x947 & n16712 ;
  assign n32887 = ~n32846 & n32886 ;
  assign n32888 = n32885 | n32887 ;
  assign n32889 = ~n4764 & n32888 ;
  assign n32890 = n4764 & ~n32850 ;
  assign n32891 = n18925 & n32890 ;
  assign n32892 = n1823 & ~n32891 ;
  assign n32893 = ~n32889 & n32892 ;
  assign n32894 = ~n1823 & n32858 ;
  assign n32895 = x223 | n32894 ;
  assign n32896 = n32762 & ~n32895 ;
  assign n32897 = ~n32893 & n32896 ;
  assign n32898 = ( x947 & ~n4764 ) | ( x947 & n32868 ) | ( ~n4764 & n32868 ) ;
  assign n32899 = ~x616 & n14492 ;
  assign n32900 = ~n14481 & n14554 ;
  assign n32901 = n4711 | n32900 ;
  assign n32902 = n32899 | n32901 ;
  assign n32903 = x614 | n32771 ;
  assign n32904 = n32902 & ~n32903 ;
  assign n32905 = ( x947 & n4764 ) | ( x947 & n32904 ) | ( n4764 & n32904 ) ;
  assign n32906 = n32898 & n32905 ;
  assign n32907 = n19090 | n32906 ;
  assign n32908 = x223 & ~n32847 ;
  assign n32909 = n32907 & n32908 ;
  assign n32910 = x216 & ~n32909 ;
  assign n32911 = ~n32897 & n32910 ;
  assign n32912 = n14678 & n32847 ;
  assign n32913 = x947 & n14639 ;
  assign n32914 = n4764 | n32913 ;
  assign n32915 = n32912 | n32914 ;
  assign n32916 = ( n1823 & n15052 ) | ( n1823 & n32856 ) | ( n15052 & n32856 ) ;
  assign n32917 = n32915 & n32916 ;
  assign n32918 = n16705 & n32894 ;
  assign n32919 = x223 | n32918 ;
  assign n32920 = n32917 | n32919 ;
  assign n32921 = n32816 & n32846 ;
  assign n32922 = x947 | n32921 ;
  assign n32923 = n32811 | n32875 ;
  assign n32924 = n32922 & ~n32923 ;
  assign n32925 = x223 & ~n32924 ;
  assign n32926 = x216 | n32925 ;
  assign n32927 = n32920 & ~n32926 ;
  assign n32928 = n32911 | n32927 ;
  assign n32929 = ( x39 & n4757 ) | ( x39 & n32928 ) | ( n4757 & n32928 ) ;
  assign n32930 = ~n32884 & n32929 ;
  assign n32931 = ( x299 & n14820 ) | ( x299 & n32858 ) | ( n14820 & n32858 ) ;
  assign n32932 = ( x216 & x299 ) | ( x216 & ~n14820 ) | ( x299 & ~n14820 ) ;
  assign n32933 = n32931 | n32932 ;
  assign n32934 = ( ~x299 & n14814 ) | ( ~x299 & n32858 ) | ( n14814 & n32858 ) ;
  assign n32935 = ( ~x216 & x299 ) | ( ~x216 & n14814 ) | ( x299 & n14814 ) ;
  assign n32936 = ~n32934 & n32935 ;
  assign n32937 = n32933 & ~n32936 ;
  assign n32938 = ( x38 & ~n9138 ) | ( x38 & n32937 ) | ( ~n9138 & n32937 ) ;
  assign n32939 = n32930 | n32938 ;
  assign n32940 = ( ~x38 & n15070 ) | ( ~x38 & n32858 ) | ( n15070 & n32858 ) ;
  assign n32941 = ( x38 & ~x216 ) | ( x38 & n15070 ) | ( ~x216 & n15070 ) ;
  assign n32942 = ~n32940 & n32941 ;
  assign n32943 = n32939 & ~n32942 ;
  assign n32944 = n8359 | n32943 ;
  assign n32945 = ~x216 & n8359 ;
  assign n32946 = n32944 & ~n32945 ;
  assign n32947 = ~x695 & n32524 ;
  assign n32948 = x217 & ~n32947 ;
  assign n32949 = x612 | n32948 ;
  assign n32950 = ( x217 & x695 ) | ( x217 & ~n32466 ) | ( x695 & ~n32466 ) ;
  assign n32951 = ( ~x217 & x695 ) | ( ~x217 & n32464 ) | ( x695 & n32464 ) ;
  assign n32952 = ~n32950 & n32951 ;
  assign n32953 = n32949 | n32952 ;
  assign n32954 = ( ~x217 & x695 ) | ( ~x217 & n32530 ) | ( x695 & n32530 ) ;
  assign n32955 = ( x217 & x695 ) | ( x217 & ~n32508 ) | ( x695 & ~n32508 ) ;
  assign n32956 = ~n32954 & n32955 ;
  assign n32957 = x612 & ~n32956 ;
  assign n32958 = ( x217 & x695 ) | ( x217 & ~n32440 ) | ( x695 & ~n32440 ) ;
  assign n32959 = ( ~x217 & x695 ) | ( ~x217 & n32433 ) | ( x695 & n32433 ) ;
  assign n32960 = ~n32958 & n32959 ;
  assign n32961 = n32957 & ~n32960 ;
  assign n32962 = n32953 & ~n32961 ;
  assign n32963 = ~n31750 & n31761 ;
  assign n32964 = x218 & ~n32963 ;
  assign n32965 = ( x218 & n31750 ) | ( x218 & ~n31855 ) | ( n31750 & ~n31855 ) ;
  assign n32966 = ( ~x218 & n31750 ) | ( ~x218 & n31826 ) | ( n31750 & n31826 ) ;
  assign n32967 = ~n32965 & n32966 ;
  assign n32968 = n32964 | n32967 ;
  assign n32969 = x219 | n6785 ;
  assign n32970 = x617 & ~x637 ;
  assign n32971 = n32667 & n32970 ;
  assign n32972 = ( x617 & x637 ) | ( x617 & n32670 ) | ( x637 & n32670 ) ;
  assign n32973 = ( ~x617 & x637 ) | ( ~x617 & n32672 ) | ( x637 & n32672 ) ;
  assign n32974 = n32972 & n32973 ;
  assign n32975 = n32971 | n32974 ;
  assign n32976 = ~n32969 & n32975 ;
  assign n32977 = x219 & n6785 ;
  assign n32978 = ( x617 & x637 ) | ( x617 & ~n32660 ) | ( x637 & ~n32660 ) ;
  assign n32979 = ( x617 & ~x637 ) | ( x617 & n32662 ) | ( ~x637 & n32662 ) ;
  assign n32980 = n32978 & ~n32979 ;
  assign n32981 = ( x617 & x637 ) | ( x617 & n32655 ) | ( x637 & n32655 ) ;
  assign n32982 = ( ~x617 & x637 ) | ( ~x617 & n14834 ) | ( x637 & n14834 ) ;
  assign n32983 = n32981 | n32982 ;
  assign n32984 = ~n32980 & n32983 ;
  assign n32985 = ( x219 & n32977 ) | ( x219 & ~n32984 ) | ( n32977 & ~n32984 ) ;
  assign n32986 = n32976 | n32985 ;
  assign n32987 = n31571 & n31865 ;
  assign n32988 = x220 & ~n32987 ;
  assign n32989 = ( x220 & ~n31703 ) | ( x220 & n31865 ) | ( ~n31703 & n31865 ) ;
  assign n32990 = ( ~x220 & n31739 ) | ( ~x220 & n31865 ) | ( n31739 & n31865 ) ;
  assign n32991 = ~n32989 & n32990 ;
  assign n32992 = n32988 | n32991 ;
  assign n32993 = x661 & x907 ;
  assign n32994 = n18994 & ~n32993 ;
  assign n32995 = x947 | n32994 ;
  assign n32996 = ~n14481 & n14674 ;
  assign n32997 = ( n14652 & n14671 ) | ( n14652 & n32996 ) | ( n14671 & n32996 ) ;
  assign n32998 = n4713 & n32997 ;
  assign n32999 = n14609 | n32998 ;
  assign n33000 = n14563 & n32999 ;
  assign n33001 = n32747 | n32797 ;
  assign n33002 = ~n14536 & n33001 ;
  assign n33003 = x947 & ~n33002 ;
  assign n33004 = ~n33000 & n33003 ;
  assign n33005 = x221 & ~n33004 ;
  assign n33006 = n32995 & n33005 ;
  assign n33007 = x616 & x947 ;
  assign n33008 = n32796 & n33007 ;
  assign n33009 = ~x947 & n32993 ;
  assign n33010 = n14614 & n33009 ;
  assign n33011 = n33008 | n33010 ;
  assign n33012 = ( x216 & x221 ) | ( x216 & n33011 ) | ( x221 & n33011 ) ;
  assign n33013 = n33007 | n33009 ;
  assign n33014 = n16705 & n33013 ;
  assign n33015 = ( ~x216 & x221 ) | ( ~x216 & n33014 ) | ( x221 & n33014 ) ;
  assign n33016 = n33012 | n33015 ;
  assign n33017 = ~x215 & n33016 ;
  assign n33018 = ~n33006 & n33017 ;
  assign n33019 = n14515 & n14521 ;
  assign n33020 = n4711 | n33019 ;
  assign n33021 = x616 | n32739 ;
  assign n33022 = n33020 & ~n33021 ;
  assign n33023 = x947 & ~n33022 ;
  assign n33024 = x221 & ~n33009 ;
  assign n33025 = ~n33023 & n33024 ;
  assign n33026 = n32734 & n33025 ;
  assign n33027 = ( ~n14552 & n14557 ) | ( ~n14552 & n14559 ) | ( n14557 & n14559 ) ;
  assign n33028 = x947 & n33027 ;
  assign n33029 = n33009 | n33028 ;
  assign n33030 = n32810 & n33029 ;
  assign n33031 = x221 | n33030 ;
  assign n33032 = x215 & n33031 ;
  assign n33033 = ~n33026 & n33032 ;
  assign n33034 = x299 & ~n33033 ;
  assign n33035 = ~n33018 & n33034 ;
  assign n33036 = n14563 & n32997 ;
  assign n33037 = ( ~n14624 & n14633 ) | ( ~n14624 & n14637 ) | ( n14633 & n14637 ) ;
  assign n33038 = n14665 | n33037 ;
  assign n33039 = ~n14536 & n33038 ;
  assign n33040 = n33036 | n33039 ;
  assign n33041 = x947 & n33040 ;
  assign n33042 = n4764 | n32886 ;
  assign n33043 = n33041 | n33042 ;
  assign n33044 = n18925 & ~n33004 ;
  assign n33045 = n4764 & ~n33044 ;
  assign n33046 = n33009 | n33045 ;
  assign n33047 = n33043 & ~n33046 ;
  assign n33048 = n1823 & ~n33047 ;
  assign n33049 = ( x223 & ~n15629 ) | ( x223 & n33014 ) | ( ~n15629 & n33014 ) ;
  assign n33050 = n32762 & ~n33049 ;
  assign n33051 = ~n33048 & n33050 ;
  assign n33052 = x947 | n14528 ;
  assign n33053 = ~n33023 & n33052 ;
  assign n33054 = n4764 & ~n33053 ;
  assign n33055 = x223 & ~n33009 ;
  assign n33056 = n14543 | n14568 ;
  assign n33057 = ( x947 & n4764 ) | ( x947 & n33056 ) | ( n4764 & n33056 ) ;
  assign n33058 = ( ~x947 & n4764 ) | ( ~x947 & n16719 ) | ( n4764 & n16719 ) ;
  assign n33059 = n33057 | n33058 ;
  assign n33060 = n33055 & n33059 ;
  assign n33061 = ~n33054 & n33060 ;
  assign n33062 = x221 & ~n33061 ;
  assign n33063 = ~n33051 & n33062 ;
  assign n33064 = n14678 & n33009 ;
  assign n33065 = n14549 & ~n32789 ;
  assign n33066 = n14556 | n33065 ;
  assign n33067 = x947 & n33066 ;
  assign n33068 = n4764 | n33067 ;
  assign n33069 = n33064 | n33068 ;
  assign n33070 = ( n1823 & n15052 ) | ( n1823 & n33011 ) | ( n15052 & n33011 ) ;
  assign n33071 = n33069 & n33070 ;
  assign n33072 = n33049 | n33071 ;
  assign n33073 = n32816 | n33028 ;
  assign n33074 = ~n32811 & n33029 ;
  assign n33075 = n33073 & n33074 ;
  assign n33076 = x223 & ~n33075 ;
  assign n33077 = x221 | n33076 ;
  assign n33078 = n33072 & ~n33077 ;
  assign n33079 = n33063 | n33078 ;
  assign n33080 = ( x39 & n4757 ) | ( x39 & n33079 ) | ( n4757 & n33079 ) ;
  assign n33081 = ~n33035 & n33080 ;
  assign n33082 = ( x299 & n14820 ) | ( x299 & n33013 ) | ( n14820 & n33013 ) ;
  assign n33083 = ( x221 & x299 ) | ( x221 & ~n14820 ) | ( x299 & ~n14820 ) ;
  assign n33084 = n33082 | n33083 ;
  assign n33085 = ( ~x299 & n14814 ) | ( ~x299 & n33013 ) | ( n14814 & n33013 ) ;
  assign n33086 = ( ~x221 & x299 ) | ( ~x221 & n14814 ) | ( x299 & n14814 ) ;
  assign n33087 = ~n33085 & n33086 ;
  assign n33088 = n33084 & ~n33087 ;
  assign n33089 = ( x38 & ~n9138 ) | ( x38 & n33088 ) | ( ~n9138 & n33088 ) ;
  assign n33090 = n33081 | n33089 ;
  assign n33091 = ( ~x38 & n15070 ) | ( ~x38 & n33013 ) | ( n15070 & n33013 ) ;
  assign n33092 = ( x38 & ~x221 ) | ( x38 & n15070 ) | ( ~x221 & n15070 ) ;
  assign n33093 = ~n33091 & n33092 ;
  assign n33094 = n33090 & ~n33093 ;
  assign n33095 = n8359 | n33094 ;
  assign n33096 = ~x221 & n8359 ;
  assign n33097 = n33095 & ~n33096 ;
  assign n33098 = ~x222 & n6785 ;
  assign n33099 = x223 | n19382 ;
  assign n33100 = ~n14707 & n33099 ;
  assign n33101 = x299 | n33100 ;
  assign n33102 = x39 & n33101 ;
  assign n33103 = ~n14692 & n33102 ;
  assign n33104 = x38 | n14823 ;
  assign n33105 = n33103 | n33104 ;
  assign n33106 = ~n14828 & n33105 ;
  assign n33107 = x222 & ~n33106 ;
  assign n33108 = n15141 & ~n33107 ;
  assign n33109 = n16176 & ~n33107 ;
  assign n33110 = x222 & n2032 ;
  assign n33111 = n14839 & n32900 ;
  assign n33112 = x224 | n33111 ;
  assign n33113 = ~x222 & n33112 ;
  assign n33114 = x616 & n14839 ;
  assign n33115 = n15503 & n33114 ;
  assign n33116 = n4710 & ~n33115 ;
  assign n33117 = ~n4709 & n33115 ;
  assign n33118 = x616 & n4709 ;
  assign n33119 = n15815 & n33118 ;
  assign n33120 = n4710 | n33119 ;
  assign n33121 = n33117 | n33120 ;
  assign n33122 = ~n33116 & n33121 ;
  assign n33123 = ( ~x224 & n4764 ) | ( ~x224 & n33122 ) | ( n4764 & n33122 ) ;
  assign n33124 = ~n4711 & n14874 ;
  assign n33125 = n14869 | n33124 ;
  assign n33126 = x616 & n33125 ;
  assign n33127 = ( x224 & n4764 ) | ( x224 & ~n33126 ) | ( n4764 & ~n33126 ) ;
  assign n33128 = ~n33123 & n33127 ;
  assign n33129 = n33113 & ~n33128 ;
  assign n33130 = x223 | n33129 ;
  assign n33131 = x616 & ~n15010 ;
  assign n33132 = x616 | n32999 ;
  assign n33133 = ~n33131 & n33132 ;
  assign n33134 = n4710 & ~n33133 ;
  assign n33135 = n15019 & ~n33114 ;
  assign n33136 = n15011 | n33135 ;
  assign n33137 = ( n4709 & n4710 ) | ( n4709 & n33136 ) | ( n4710 & n33136 ) ;
  assign n33138 = ( ~n4709 & n4710 ) | ( ~n4709 & n33133 ) | ( n4710 & n33133 ) ;
  assign n33139 = n33137 | n33138 ;
  assign n33140 = ~n33134 & n33139 ;
  assign n33141 = ( ~x222 & n4764 ) | ( ~x222 & n33140 ) | ( n4764 & n33140 ) ;
  assign n33142 = ( n14652 & n14672 ) | ( n14652 & n14676 ) | ( n14672 & n14676 ) ;
  assign n33143 = ~n14481 & n14959 ;
  assign n33144 = x616 & ~n33143 ;
  assign n33145 = n33142 & ~n33144 ;
  assign n33146 = n4710 & ~n33145 ;
  assign n33147 = ~n4709 & n33145 ;
  assign n33148 = n4709 & ~n33114 ;
  assign n33149 = n14641 & n33148 ;
  assign n33150 = n4710 | n33149 ;
  assign n33151 = n33147 | n33150 ;
  assign n33152 = ~n33146 & n33151 ;
  assign n33153 = ( x222 & n4764 ) | ( x222 & ~n33152 ) | ( n4764 & ~n33152 ) ;
  assign n33154 = ~n33141 & n33153 ;
  assign n33155 = n33130 | n33154 ;
  assign n33156 = n14884 | n33124 ;
  assign n33157 = x616 & n33156 ;
  assign n33158 = ~x222 & n33157 ;
  assign n33159 = ~n14900 & n33158 ;
  assign n33160 = x223 & ~n33159 ;
  assign n33161 = x616 & ~n14959 ;
  assign n33162 = n32737 & ~n33161 ;
  assign n33163 = n4710 & ~n33162 ;
  assign n33164 = n4709 | n32737 ;
  assign n33165 = ~n33161 & n33164 ;
  assign n33166 = ( n4710 & ~n32739 ) | ( n4710 & n33165 ) | ( ~n32739 & n33165 ) ;
  assign n33167 = ~n33163 & n33166 ;
  assign n33168 = ( ~x222 & n4764 ) | ( ~x222 & n33167 ) | ( n4764 & n33167 ) ;
  assign n33169 = ( n14492 & ~n14538 ) | ( n14492 & n14540 ) | ( ~n14538 & n14540 ) ;
  assign n33170 = ~n33144 & n33169 ;
  assign n33171 = n4710 & ~n33170 ;
  assign n33172 = ~n4709 & n33170 ;
  assign n33173 = n30485 & n33148 ;
  assign n33174 = n4710 | n33173 ;
  assign n33175 = n33172 | n33174 ;
  assign n33176 = ~n33171 & n33175 ;
  assign n33177 = ( x222 & n4764 ) | ( x222 & ~n33176 ) | ( n4764 & ~n33176 ) ;
  assign n33178 = ~n33168 & n33177 ;
  assign n33179 = n33160 & ~n33178 ;
  assign n33180 = n33155 & ~n33179 ;
  assign n33181 = x299 | n33180 ;
  assign n33182 = ( x222 & n4721 ) | ( x222 & ~n33122 ) | ( n4721 & ~n33122 ) ;
  assign n33183 = ( ~x222 & n4721 ) | ( ~x222 & n33126 ) | ( n4721 & n33126 ) ;
  assign n33184 = ~n33182 & n33183 ;
  assign n33185 = n2203 & ~n33184 ;
  assign n33186 = ( ~x222 & n4721 ) | ( ~x222 & n33140 ) | ( n4721 & n33140 ) ;
  assign n33187 = ( x222 & n4721 ) | ( x222 & ~n33152 ) | ( n4721 & ~n33152 ) ;
  assign n33188 = ~n33186 & n33187 ;
  assign n33189 = n33185 & ~n33188 ;
  assign n33190 = x222 & ~n16705 ;
  assign n33191 = n2203 | n33190 ;
  assign n33192 = n33111 | n33191 ;
  assign n33193 = ~x215 & n33192 ;
  assign n33194 = ~n33189 & n33193 ;
  assign n33195 = ~n14873 & n33158 ;
  assign n33196 = ( ~x222 & n4721 ) | ( ~x222 & n33167 ) | ( n4721 & n33167 ) ;
  assign n33197 = ( x222 & n4721 ) | ( x222 & ~n33176 ) | ( n4721 & ~n33176 ) ;
  assign n33198 = ~n33196 & n33197 ;
  assign n33199 = n33195 | n33198 ;
  assign n33200 = x215 & n33199 ;
  assign n33201 = x299 & ~n33200 ;
  assign n33202 = ~n33194 & n33201 ;
  assign n33203 = x39 & ~n33202 ;
  assign n33204 = n33181 & n33203 ;
  assign n33205 = ~x39 & x616 ;
  assign n33206 = ( x39 & n15896 ) | ( x39 & ~n33205 ) | ( n15896 & ~n33205 ) ;
  assign n33207 = ( x222 & n15896 ) | ( x222 & ~n33206 ) | ( n15896 & ~n33206 ) ;
  assign n33208 = ( x222 & n14956 ) | ( x222 & n33206 ) | ( n14956 & n33206 ) ;
  assign n33209 = n33207 & ~n33208 ;
  assign n33210 = x38 | n33209 ;
  assign n33211 = n33204 | n33210 ;
  assign n33212 = x222 & ~n15070 ;
  assign n33213 = x38 & ~n33212 ;
  assign n33214 = x616 & n15072 ;
  assign n33215 = n33213 & ~n33214 ;
  assign n33216 = n2032 | n33215 ;
  assign n33217 = n33211 & ~n33216 ;
  assign n33218 = n33110 | n33217 ;
  assign n33219 = ~n15082 & n33218 ;
  assign n33220 = n15082 & n33107 ;
  assign n33221 = n33219 | n33220 ;
  assign n33222 = ~x785 & n33221 ;
  assign n33223 = ( x609 & x1155 ) | ( x609 & n33107 ) | ( x1155 & n33107 ) ;
  assign n33224 = ( ~x609 & x1155 ) | ( ~x609 & n33221 ) | ( x1155 & n33221 ) ;
  assign n33225 = n33223 & n33224 ;
  assign n33226 = ( x609 & x1155 ) | ( x609 & ~n33107 ) | ( x1155 & ~n33107 ) ;
  assign n33227 = ( x609 & ~x1155 ) | ( x609 & n33221 ) | ( ~x1155 & n33221 ) ;
  assign n33228 = ~n33226 & n33227 ;
  assign n33229 = n33225 | n33228 ;
  assign n33230 = x785 & n33229 ;
  assign n33231 = n33222 | n33230 ;
  assign n33232 = ~x781 & n33231 ;
  assign n33233 = ( x618 & x1154 ) | ( x618 & n33107 ) | ( x1154 & n33107 ) ;
  assign n33234 = ( ~x618 & x1154 ) | ( ~x618 & n33231 ) | ( x1154 & n33231 ) ;
  assign n33235 = n33233 & n33234 ;
  assign n33236 = ( x618 & x1154 ) | ( x618 & ~n33107 ) | ( x1154 & ~n33107 ) ;
  assign n33237 = ( x618 & ~x1154 ) | ( x618 & n33231 ) | ( ~x1154 & n33231 ) ;
  assign n33238 = ~n33236 & n33237 ;
  assign n33239 = n33235 | n33238 ;
  assign n33240 = x781 & n33239 ;
  assign n33241 = n33232 | n33240 ;
  assign n33242 = ~x789 & n33241 ;
  assign n33243 = ( x619 & x1159 ) | ( x619 & n33107 ) | ( x1159 & n33107 ) ;
  assign n33244 = ( ~x619 & x1159 ) | ( ~x619 & n33241 ) | ( x1159 & n33241 ) ;
  assign n33245 = n33243 & n33244 ;
  assign n33246 = ( x619 & x1159 ) | ( x619 & ~n33107 ) | ( x1159 & ~n33107 ) ;
  assign n33247 = ( x619 & ~x1159 ) | ( x619 & n33241 ) | ( ~x1159 & n33241 ) ;
  assign n33248 = ~n33246 & n33247 ;
  assign n33249 = n33245 | n33248 ;
  assign n33250 = x789 & n33249 ;
  assign n33251 = n33242 | n33250 ;
  assign n33252 = n16176 | n33251 ;
  assign n33253 = ~n33109 & n33252 ;
  assign n33254 = ~n15134 & n33253 ;
  assign n33255 = n15134 & n33107 ;
  assign n33256 = n33254 | n33255 ;
  assign n33257 = n15141 | n33256 ;
  assign n33258 = ~n33108 & n33257 ;
  assign n33259 = ( x644 & x715 ) | ( x644 & ~n33258 ) | ( x715 & ~n33258 ) ;
  assign n33260 = ( x644 & ~x715 ) | ( x644 & n33107 ) | ( ~x715 & n33107 ) ;
  assign n33261 = ~n33259 & n33260 ;
  assign n33262 = x1160 & ~n33261 ;
  assign n33263 = n17213 & ~n33107 ;
  assign n33264 = x661 & x680 ;
  assign n33265 = ~n15331 & n15333 ;
  assign n33266 = x222 & n33265 ;
  assign n33267 = x299 | n33266 ;
  assign n33268 = ( n15356 & ~n33264 ) | ( n15356 & n33267 ) | ( ~n33264 & n33267 ) ;
  assign n33269 = ( x222 & n15356 ) | ( x222 & ~n33267 ) | ( n15356 & ~n33267 ) ;
  assign n33270 = ~n33268 & n33269 ;
  assign n33271 = x39 | n33270 ;
  assign n33272 = x222 & n30752 ;
  assign n33273 = x299 & ~n33272 ;
  assign n33274 = ( ~n15366 & n33264 ) | ( ~n15366 & n33273 ) | ( n33264 & n33273 ) ;
  assign n33275 = ( x222 & n15366 ) | ( x222 & n33273 ) | ( n15366 & n33273 ) ;
  assign n33276 = n33274 & n33275 ;
  assign n33277 = n33271 | n33276 ;
  assign n33278 = ~n14481 & n15202 ;
  assign n33279 = x661 & n33278 ;
  assign n33280 = x224 | n33279 ;
  assign n33281 = ~x222 & n33280 ;
  assign n33282 = x661 & n15175 ;
  assign n33283 = ( ~x224 & n4764 ) | ( ~x224 & n33282 ) | ( n4764 & n33282 ) ;
  assign n33284 = ( n15158 & n15164 ) | ( n15158 & n15166 ) | ( n15164 & n15166 ) ;
  assign n33285 = n33264 & n33284 ;
  assign n33286 = ( x224 & n4764 ) | ( x224 & ~n33285 ) | ( n4764 & ~n33285 ) ;
  assign n33287 = ~n33283 & n33286 ;
  assign n33288 = n33281 & ~n33287 ;
  assign n33289 = x223 | n33288 ;
  assign n33290 = x661 | n16709 ;
  assign n33291 = n15259 | n15293 ;
  assign n33292 = x680 & ~n33291 ;
  assign n33293 = n15285 & ~n33292 ;
  assign n33294 = x661 & ~n33293 ;
  assign n33295 = n33290 & ~n33294 ;
  assign n33296 = ( ~x222 & n4764 ) | ( ~x222 & n33295 ) | ( n4764 & n33295 ) ;
  assign n33297 = ( n14678 & n15242 ) | ( n14678 & ~n15245 ) | ( n15242 & ~n15245 ) ;
  assign n33298 = n4709 | n14678 ;
  assign n33299 = ~x662 & n32789 ;
  assign n33300 = n33298 & ~n33299 ;
  assign n33301 = n4710 | n33300 ;
  assign n33302 = ( ~x661 & n33297 ) | ( ~x661 & n33301 ) | ( n33297 & n33301 ) ;
  assign n33303 = ( x661 & ~n14679 ) | ( x661 & n33301 ) | ( ~n14679 & n33301 ) ;
  assign n33304 = n33302 & n33303 ;
  assign n33305 = ( x222 & n4764 ) | ( x222 & ~n33304 ) | ( n4764 & ~n33304 ) ;
  assign n33306 = ~n33296 & n33305 ;
  assign n33307 = n33289 | n33306 ;
  assign n33308 = ~n14900 & n15188 ;
  assign n33309 = ~x222 & x661 ;
  assign n33310 = n33308 & n33309 ;
  assign n33311 = x223 & ~n33310 ;
  assign n33312 = ( n14505 & n14510 ) | ( n14505 & n14511 ) | ( n14510 & n14511 ) ;
  assign n33313 = n4710 | n33312 ;
  assign n33314 = ( ~x661 & n15264 ) | ( ~x661 & n33313 ) | ( n15264 & n33313 ) ;
  assign n33315 = ( x661 & ~n14523 ) | ( x661 & n33313 ) | ( ~n14523 & n33313 ) ;
  assign n33316 = n33314 & n33315 ;
  assign n33317 = ( ~x222 & n4764 ) | ( ~x222 & n33316 ) | ( n4764 & n33316 ) ;
  assign n33318 = x661 | n16719 ;
  assign n33319 = ~n15271 & n15275 ;
  assign n33320 = x661 & ~n33319 ;
  assign n33321 = n33318 & ~n33320 ;
  assign n33322 = ( x222 & n4764 ) | ( x222 & ~n33321 ) | ( n4764 & ~n33321 ) ;
  assign n33323 = ~n33317 & n33322 ;
  assign n33324 = n33311 & ~n33323 ;
  assign n33325 = n33307 & ~n33324 ;
  assign n33326 = x299 | n33325 ;
  assign n33327 = ( x222 & n4721 ) | ( x222 & ~n33282 ) | ( n4721 & ~n33282 ) ;
  assign n33328 = ( ~x222 & n4721 ) | ( ~x222 & n33285 ) | ( n4721 & n33285 ) ;
  assign n33329 = ~n33327 & n33328 ;
  assign n33330 = n2203 & ~n33329 ;
  assign n33331 = ( ~x222 & n4721 ) | ( ~x222 & n33295 ) | ( n4721 & n33295 ) ;
  assign n33332 = ( x222 & n4721 ) | ( x222 & ~n33304 ) | ( n4721 & ~n33304 ) ;
  assign n33333 = ~n33331 & n33332 ;
  assign n33334 = n33330 & ~n33333 ;
  assign n33335 = n33191 | n33279 ;
  assign n33336 = ~x215 & n33335 ;
  assign n33337 = ~n33334 & n33336 ;
  assign n33338 = ~n14873 & n15188 ;
  assign n33339 = n33309 & n33338 ;
  assign n33340 = ( ~x222 & n4721 ) | ( ~x222 & n33316 ) | ( n4721 & n33316 ) ;
  assign n33341 = ( x222 & n4721 ) | ( x222 & ~n33321 ) | ( n4721 & ~n33321 ) ;
  assign n33342 = ~n33340 & n33341 ;
  assign n33343 = n33339 | n33342 ;
  assign n33344 = x215 & n33343 ;
  assign n33345 = x299 & ~n33344 ;
  assign n33346 = ~n33337 & n33345 ;
  assign n33347 = n33326 & ~n33346 ;
  assign n33348 = x39 & ~n33347 ;
  assign n33349 = n33277 & ~n33348 ;
  assign n33350 = x38 | n33349 ;
  assign n33351 = x661 & n15374 ;
  assign n33352 = n33213 & ~n33351 ;
  assign n33353 = n2032 | n33352 ;
  assign n33354 = n33350 & ~n33353 ;
  assign n33355 = n33110 | n33354 ;
  assign n33356 = ~x778 & n33355 ;
  assign n33357 = ( x625 & x1153 ) | ( x625 & n33107 ) | ( x1153 & n33107 ) ;
  assign n33358 = ( ~x625 & x1153 ) | ( ~x625 & n33355 ) | ( x1153 & n33355 ) ;
  assign n33359 = n33357 & n33358 ;
  assign n33360 = ( x625 & x1153 ) | ( x625 & ~n33107 ) | ( x1153 & ~n33107 ) ;
  assign n33361 = ( x625 & ~x1153 ) | ( x625 & n33355 ) | ( ~x1153 & n33355 ) ;
  assign n33362 = ~n33360 & n33361 ;
  assign n33363 = n33359 | n33362 ;
  assign n33364 = x778 & n33363 ;
  assign n33365 = n33356 | n33364 ;
  assign n33366 = ~n15400 & n33365 ;
  assign n33367 = n15400 & n33107 ;
  assign n33368 = n33366 | n33367 ;
  assign n33369 = ~n15407 & n33368 ;
  assign n33370 = n15407 & n33107 ;
  assign n33371 = n33369 | n33370 ;
  assign n33372 = n15414 | n33371 ;
  assign n33373 = n15421 | n33372 ;
  assign n33374 = ~n33263 & n33373 ;
  assign n33375 = n17220 | n33374 ;
  assign n33376 = n16054 & ~n33107 ;
  assign n33377 = n33375 & ~n33376 ;
  assign n33378 = ~x787 & n33377 ;
  assign n33379 = ( x647 & x1157 ) | ( x647 & n33107 ) | ( x1157 & n33107 ) ;
  assign n33380 = ( ~x647 & x1157 ) | ( ~x647 & n33377 ) | ( x1157 & n33377 ) ;
  assign n33381 = n33379 & n33380 ;
  assign n33382 = ( x647 & x1157 ) | ( x647 & ~n33107 ) | ( x1157 & ~n33107 ) ;
  assign n33383 = ( x647 & ~x1157 ) | ( x647 & n33377 ) | ( ~x1157 & n33377 ) ;
  assign n33384 = ~n33382 & n33383 ;
  assign n33385 = n33381 | n33384 ;
  assign n33386 = x787 & n33385 ;
  assign n33387 = n33378 | n33386 ;
  assign n33388 = ( x644 & x715 ) | ( x644 & n33387 ) | ( x715 & n33387 ) ;
  assign n33389 = n18621 & n33253 ;
  assign n33390 = x628 | n33107 ;
  assign n33391 = n15131 & n33390 ;
  assign n33392 = x628 & ~n33107 ;
  assign n33393 = n15132 & ~n33392 ;
  assign n33394 = ( x628 & n33374 ) | ( x628 & n33393 ) | ( n33374 & n33393 ) ;
  assign n33395 = x628 & ~n33393 ;
  assign n33396 = ( n33391 & n33394 ) | ( n33391 & ~n33395 ) | ( n33394 & ~n33395 ) ;
  assign n33397 = n33389 | n33396 ;
  assign n33398 = x792 & n33397 ;
  assign n33399 = x648 & ~n33248 ;
  assign n33400 = ( x619 & x1159 ) | ( x619 & n33371 ) | ( x1159 & n33371 ) ;
  assign n33401 = x627 | n33235 ;
  assign n33402 = ( x618 & x1154 ) | ( x618 & ~n33368 ) | ( x1154 & ~n33368 ) ;
  assign n33403 = x660 | n33225 ;
  assign n33404 = ( x609 & x1155 ) | ( x609 & ~n33365 ) | ( x1155 & ~n33365 ) ;
  assign n33405 = x608 | n33359 ;
  assign n33406 = ( x625 & x1153 ) | ( x625 & ~n33218 ) | ( x1153 & ~n33218 ) ;
  assign n33407 = ~x680 & n33133 ;
  assign n33408 = ( n14595 & n15234 ) | ( n14595 & n15238 ) | ( n15234 & n15238 ) ;
  assign n33409 = ~n4713 & n33408 ;
  assign n33410 = n15642 | n33409 ;
  assign n33411 = n15821 | n33410 ;
  assign n33412 = n14495 & ~n33411 ;
  assign n33413 = n15705 & n33410 ;
  assign n33414 = x616 & ~n33413 ;
  assign n33415 = x680 & ~n33414 ;
  assign n33416 = ~n33412 & n33415 ;
  assign n33417 = ( x603 & n15535 ) | ( x603 & ~n30540 ) | ( n15535 & ~n30540 ) ;
  assign n33418 = ( x603 & ~n15535 ) | ( x603 & n33410 ) | ( ~n15535 & n33410 ) ;
  assign n33419 = ~n33417 & n33418 ;
  assign n33420 = ( ~x642 & n4707 ) | ( ~x642 & n33419 ) | ( n4707 & n33419 ) ;
  assign n33421 = ( x642 & n4707 ) | ( x642 & n33411 ) | ( n4707 & n33411 ) ;
  assign n33422 = n33420 | n33421 ;
  assign n33423 = n33416 & n33422 ;
  assign n33424 = x661 & ~n33423 ;
  assign n33425 = ~n33407 & n33424 ;
  assign n33426 = ~x661 & x681 ;
  assign n33427 = ~n33133 & n33426 ;
  assign n33428 = n33139 & ~n33427 ;
  assign n33429 = ~n33425 & n33428 ;
  assign n33430 = ( x222 & ~n4721 ) | ( x222 & n33429 ) | ( ~n4721 & n33429 ) ;
  assign n33431 = ( n15603 & n15612 ) | ( n15603 & ~n15622 ) | ( n15612 & ~n15622 ) ;
  assign n33432 = ~n14481 & n15713 ;
  assign n33433 = x616 & ~n33432 ;
  assign n33434 = x680 & ~n33433 ;
  assign n33435 = n33431 & n33434 ;
  assign n33436 = ( x661 & ~n33145 ) | ( x661 & n33264 ) | ( ~n33145 & n33264 ) ;
  assign n33437 = ~n33435 & n33436 ;
  assign n33438 = ~n33145 & n33426 ;
  assign n33439 = n33151 & ~n33438 ;
  assign n33440 = ~n33437 & n33439 ;
  assign n33441 = ( x222 & n4721 ) | ( x222 & n33440 ) | ( n4721 & n33440 ) ;
  assign n33442 = n33430 & n33441 ;
  assign n33443 = n15504 | n15821 ;
  assign n33444 = x616 & ~n33443 ;
  assign n33445 = x680 & ~n33444 ;
  assign n33446 = n15520 & n33445 ;
  assign n33447 = ( x661 & ~n33115 ) | ( x661 & n33264 ) | ( ~n33115 & n33264 ) ;
  assign n33448 = ~n33446 & n33447 ;
  assign n33449 = ~n33115 & n33426 ;
  assign n33450 = n33121 & ~n33449 ;
  assign n33451 = ~n33448 & n33450 ;
  assign n33452 = ( x222 & n4721 ) | ( x222 & n33451 ) | ( n4721 & n33451 ) ;
  assign n33453 = ~n14481 & n15802 ;
  assign n33454 = x616 & ~n33453 ;
  assign n33455 = ( n15549 & ~n15553 ) | ( n15549 & n15555 ) | ( ~n15553 & n15555 ) ;
  assign n33456 = x680 & n33455 ;
  assign n33457 = ~n33454 & n33456 ;
  assign n33458 = ( x661 & ~n33111 ) | ( x661 & n33264 ) | ( ~n33111 & n33264 ) ;
  assign n33459 = ~n33457 & n33458 ;
  assign n33460 = n15799 & n33118 ;
  assign n33461 = ~n4709 & n33111 ;
  assign n33462 = n4710 | n33461 ;
  assign n33463 = n33460 | n33462 ;
  assign n33464 = ~n33111 & n33426 ;
  assign n33465 = n33463 & ~n33464 ;
  assign n33466 = ~n33459 & n33465 ;
  assign n33467 = ( x222 & ~n4721 ) | ( x222 & n33466 ) | ( ~n4721 & n33466 ) ;
  assign n33468 = n33452 | n33467 ;
  assign n33469 = ~n33442 & n33468 ;
  assign n33470 = n2203 & ~n33469 ;
  assign n33471 = n33114 | n33264 ;
  assign n33472 = ~n14481 & n15490 ;
  assign n33473 = x616 | n33472 ;
  assign n33474 = ~n33454 & n33473 ;
  assign n33475 = n33471 & n33474 ;
  assign n33476 = n33191 | n33475 ;
  assign n33477 = ~x215 & n33476 ;
  assign n33478 = ~n33470 & n33477 ;
  assign n33479 = n15472 & ~n15473 ;
  assign n33480 = n14876 | n15848 ;
  assign n33481 = x616 & ~n33480 ;
  assign n33482 = x680 & ~n33481 ;
  assign n33483 = n33479 & n33482 ;
  assign n33484 = x616 & n14876 ;
  assign n33485 = ( x661 & n33264 ) | ( x661 & ~n33484 ) | ( n33264 & ~n33484 ) ;
  assign n33486 = ~n33483 & n33485 ;
  assign n33487 = x661 | n33484 ;
  assign n33488 = n14475 & n33111 ;
  assign n33489 = n4711 & ~n33488 ;
  assign n33490 = n33487 & ~n33489 ;
  assign n33491 = ~n33486 & n33490 ;
  assign n33492 = ( x222 & n4721 ) | ( x222 & n33491 ) | ( n4721 & n33491 ) ;
  assign n33493 = n14988 & ~n15149 ;
  assign n33494 = n33264 & n33493 ;
  assign n33495 = n33157 | n33494 ;
  assign n33496 = ( x222 & ~n4721 ) | ( x222 & n33495 ) | ( ~n4721 & n33495 ) ;
  assign n33497 = n33492 | n33496 ;
  assign n33498 = x215 & n33497 ;
  assign n33499 = ~x680 & n33162 ;
  assign n33500 = n15643 & n15705 ;
  assign n33501 = x616 & ~n33500 ;
  assign n33502 = x680 & ~n33501 ;
  assign n33503 = n15646 & n33502 ;
  assign n33504 = x661 & ~n33503 ;
  assign n33505 = ~n33499 & n33504 ;
  assign n33506 = ~n33162 & n33426 ;
  assign n33507 = n33166 & ~n33506 ;
  assign n33508 = ~n33505 & n33507 ;
  assign n33509 = ( x222 & ~n4721 ) | ( x222 & n33508 ) | ( ~n4721 & n33508 ) ;
  assign n33510 = ( ~n15622 & n15667 ) | ( ~n15622 & n15673 ) | ( n15667 & n15673 ) ;
  assign n33511 = n33434 & n33510 ;
  assign n33512 = ( x661 & ~n33170 ) | ( x661 & n33264 ) | ( ~n33170 & n33264 ) ;
  assign n33513 = ~n33511 & n33512 ;
  assign n33514 = ~n33170 & n33426 ;
  assign n33515 = n33175 & ~n33514 ;
  assign n33516 = ~n33513 & n33515 ;
  assign n33517 = ( x222 & n4721 ) | ( x222 & n33516 ) | ( n4721 & n33516 ) ;
  assign n33518 = n33509 & n33517 ;
  assign n33519 = n33498 & ~n33518 ;
  assign n33520 = x299 & ~n33519 ;
  assign n33521 = ~n33478 & n33520 ;
  assign n33522 = ( ~x222 & n33111 ) | ( ~x222 & n33264 ) | ( n33111 & n33264 ) ;
  assign n33523 = ( x222 & n33264 ) | ( x222 & ~n33474 ) | ( n33264 & ~n33474 ) ;
  assign n33524 = n33522 & ~n33523 ;
  assign n33525 = n1817 | n33524 ;
  assign n33526 = ( ~x224 & n4764 ) | ( ~x224 & n33451 ) | ( n4764 & n33451 ) ;
  assign n33527 = ( x224 & n4764 ) | ( x224 & ~n33466 ) | ( n4764 & ~n33466 ) ;
  assign n33528 = ~n33526 & n33527 ;
  assign n33529 = n33525 & ~n33528 ;
  assign n33530 = ( ~x222 & n4764 ) | ( ~x222 & n33429 ) | ( n4764 & n33429 ) ;
  assign n33531 = ( x222 & n4764 ) | ( x222 & ~n33440 ) | ( n4764 & ~n33440 ) ;
  assign n33532 = ~n33530 & n33531 ;
  assign n33533 = n33529 | n33532 ;
  assign n33534 = ~x223 & n33533 ;
  assign n33535 = ( x222 & n4764 ) | ( x222 & n33491 ) | ( n4764 & n33491 ) ;
  assign n33536 = ( x222 & ~n4764 ) | ( x222 & n33495 ) | ( ~n4764 & n33495 ) ;
  assign n33537 = n33535 | n33536 ;
  assign n33538 = x223 & n33537 ;
  assign n33539 = ( x222 & ~n4764 ) | ( x222 & n33508 ) | ( ~n4764 & n33508 ) ;
  assign n33540 = ( x222 & n4764 ) | ( x222 & n33516 ) | ( n4764 & n33516 ) ;
  assign n33541 = n33539 & n33540 ;
  assign n33542 = n33538 & ~n33541 ;
  assign n33543 = n33534 | n33542 ;
  assign n33544 = ( x39 & n4757 ) | ( x39 & n33543 ) | ( n4757 & n33543 ) ;
  assign n33545 = ~n33521 & n33544 ;
  assign n33546 = ~x616 & n14920 ;
  assign n33547 = x603 | n30752 ;
  assign n33548 = n14945 | n15463 ;
  assign n33549 = n33547 & ~n33548 ;
  assign n33550 = n33546 | n33549 ;
  assign n33551 = x661 & n16998 ;
  assign n33552 = ( n15885 & n33550 ) | ( n15885 & ~n33551 ) | ( n33550 & ~n33551 ) ;
  assign n33553 = x222 & n33552 ;
  assign n33554 = x616 & n14920 ;
  assign n33555 = x222 | n33554 ;
  assign n33556 = n33551 | n33555 ;
  assign n33557 = ~n33553 & n33556 ;
  assign n33558 = ( x39 & x299 ) | ( x39 & ~n33557 ) | ( x299 & ~n33557 ) ;
  assign n33559 = x661 & n16990 ;
  assign n33560 = x616 & n16781 ;
  assign n33561 = x222 | n33560 ;
  assign n33562 = n33559 | n33561 ;
  assign n33563 = n15881 & ~n33264 ;
  assign n33564 = ~x616 & n16781 ;
  assign n33565 = x603 | n33265 ;
  assign n33566 = n15463 | n15878 ;
  assign n33567 = n33565 & ~n33566 ;
  assign n33568 = n33564 | n33567 ;
  assign n33569 = n33563 | n33568 ;
  assign n33570 = x222 & n33569 ;
  assign n33571 = n33562 & ~n33570 ;
  assign n33572 = ( ~x39 & x299 ) | ( ~x39 & n33571 ) | ( x299 & n33571 ) ;
  assign n33573 = ~n33558 & n33572 ;
  assign n33574 = x38 | n33573 ;
  assign n33575 = n33545 | n33574 ;
  assign n33576 = n15705 & n15756 ;
  assign n33577 = x222 | x616 ;
  assign n33578 = n33205 & n33264 ;
  assign n33579 = n33577 & ~n33578 ;
  assign n33580 = n33576 & ~n33579 ;
  assign n33581 = x616 | n15477 ;
  assign n33582 = n33471 & n33581 ;
  assign n33583 = n15070 & n33582 ;
  assign n33584 = n33212 | n33583 ;
  assign n33585 = ~n33580 & n33584 ;
  assign n33586 = x38 & ~n33585 ;
  assign n33587 = n2032 | n33586 ;
  assign n33588 = n33575 & ~n33587 ;
  assign n33589 = n33110 | n33588 ;
  assign n33590 = ( x625 & ~x1153 ) | ( x625 & n33589 ) | ( ~x1153 & n33589 ) ;
  assign n33591 = ~n33406 & n33590 ;
  assign n33592 = n33405 | n33591 ;
  assign n33593 = x608 & ~n33362 ;
  assign n33594 = ( x625 & x1153 ) | ( x625 & n33218 ) | ( x1153 & n33218 ) ;
  assign n33595 = ( ~x625 & x1153 ) | ( ~x625 & n33589 ) | ( x1153 & n33589 ) ;
  assign n33596 = n33594 & n33595 ;
  assign n33597 = n33593 & ~n33596 ;
  assign n33598 = n33592 & ~n33597 ;
  assign n33599 = x778 & ~n33598 ;
  assign n33600 = x778 | n33589 ;
  assign n33601 = ~n33599 & n33600 ;
  assign n33602 = ( x609 & ~x1155 ) | ( x609 & n33601 ) | ( ~x1155 & n33601 ) ;
  assign n33603 = ~n33404 & n33602 ;
  assign n33604 = n33403 | n33603 ;
  assign n33605 = x660 & ~n33228 ;
  assign n33606 = ( x609 & x1155 ) | ( x609 & n33365 ) | ( x1155 & n33365 ) ;
  assign n33607 = ( ~x609 & x1155 ) | ( ~x609 & n33601 ) | ( x1155 & n33601 ) ;
  assign n33608 = n33606 & n33607 ;
  assign n33609 = n33605 & ~n33608 ;
  assign n33610 = n33604 & ~n33609 ;
  assign n33611 = x785 & ~n33610 ;
  assign n33612 = x785 | n33601 ;
  assign n33613 = ~n33611 & n33612 ;
  assign n33614 = ( x618 & ~x1154 ) | ( x618 & n33613 ) | ( ~x1154 & n33613 ) ;
  assign n33615 = ~n33402 & n33614 ;
  assign n33616 = n33401 | n33615 ;
  assign n33617 = x627 & ~n33238 ;
  assign n33618 = ( x618 & x1154 ) | ( x618 & n33368 ) | ( x1154 & n33368 ) ;
  assign n33619 = ( ~x618 & x1154 ) | ( ~x618 & n33613 ) | ( x1154 & n33613 ) ;
  assign n33620 = n33618 & n33619 ;
  assign n33621 = n33617 & ~n33620 ;
  assign n33622 = n33616 & ~n33621 ;
  assign n33623 = x781 & ~n33622 ;
  assign n33624 = x781 | n33613 ;
  assign n33625 = ~n33623 & n33624 ;
  assign n33626 = ( ~x619 & x1159 ) | ( ~x619 & n33625 ) | ( x1159 & n33625 ) ;
  assign n33627 = n33400 & n33626 ;
  assign n33628 = n33399 & ~n33627 ;
  assign n33629 = x648 | n33245 ;
  assign n33630 = ( x619 & x1159 ) | ( x619 & ~n33371 ) | ( x1159 & ~n33371 ) ;
  assign n33631 = ( x619 & ~x1159 ) | ( x619 & n33625 ) | ( ~x1159 & n33625 ) ;
  assign n33632 = ~n33630 & n33631 ;
  assign n33633 = n33629 | n33632 ;
  assign n33634 = x789 & n33633 ;
  assign n33635 = ~n33628 & n33634 ;
  assign n33636 = ~x789 & n33625 ;
  assign n33637 = n15414 & ~n33107 ;
  assign n33638 = n16115 & ~n33637 ;
  assign n33639 = n33372 & n33638 ;
  assign n33640 = ( ~x626 & n15419 ) | ( ~x626 & n33107 ) | ( n15419 & n33107 ) ;
  assign n33641 = ( x626 & n15419 ) | ( x626 & n33251 ) | ( n15419 & n33251 ) ;
  assign n33642 = n33640 & n33641 ;
  assign n33643 = n33639 | n33642 ;
  assign n33644 = ( x626 & n15418 ) | ( x626 & n33107 ) | ( n15418 & n33107 ) ;
  assign n33645 = ( ~x626 & n15418 ) | ( ~x626 & n33251 ) | ( n15418 & n33251 ) ;
  assign n33646 = n33644 & n33645 ;
  assign n33647 = n33643 | n33646 ;
  assign n33648 = x788 & n33647 ;
  assign n33649 = n33636 | n33648 ;
  assign n33650 = n33635 | n33649 ;
  assign n33651 = n16177 & ~n33647 ;
  assign n33652 = n18434 | n33651 ;
  assign n33653 = n33650 & ~n33652 ;
  assign n33654 = n33398 | n33653 ;
  assign n33655 = ~n18431 & n33654 ;
  assign n33656 = n18610 & n33256 ;
  assign n33657 = ( x630 & n33384 ) | ( x630 & n33656 ) | ( n33384 & n33656 ) ;
  assign n33658 = ( ~x630 & n33381 ) | ( ~x630 & n33656 ) | ( n33381 & n33656 ) ;
  assign n33659 = n33657 | n33658 ;
  assign n33660 = x787 & n33659 ;
  assign n33661 = n33655 | n33660 ;
  assign n33662 = ( ~x644 & x715 ) | ( ~x644 & n33661 ) | ( x715 & n33661 ) ;
  assign n33663 = n33388 & n33662 ;
  assign n33664 = n33262 & ~n33663 ;
  assign n33665 = ( x644 & x715 ) | ( x644 & n33258 ) | ( x715 & n33258 ) ;
  assign n33666 = ( ~x644 & x715 ) | ( ~x644 & n33107 ) | ( x715 & n33107 ) ;
  assign n33667 = n33665 & n33666 ;
  assign n33668 = x1160 | n33667 ;
  assign n33669 = ( x644 & x715 ) | ( x644 & ~n33387 ) | ( x715 & ~n33387 ) ;
  assign n33670 = ( x644 & ~x715 ) | ( x644 & n33661 ) | ( ~x715 & n33661 ) ;
  assign n33671 = ~n33669 & n33670 ;
  assign n33672 = n33668 | n33671 ;
  assign n33673 = ~n33664 & n33672 ;
  assign n33674 = ( x790 & n6785 ) | ( x790 & n33673 ) | ( n6785 & n33673 ) ;
  assign n33675 = ( ~x790 & n6785 ) | ( ~x790 & n33661 ) | ( n6785 & n33661 ) ;
  assign n33676 = n33674 | n33675 ;
  assign n33677 = ~n33098 & n33676 ;
  assign n33678 = ~x223 & n6785 ;
  assign n33679 = x299 | n19089 ;
  assign n33680 = x39 & n33679 ;
  assign n33681 = ~n14692 & n33680 ;
  assign n33682 = n12808 | n14823 ;
  assign n33683 = n33681 | n33682 ;
  assign n33684 = ~n14828 & n33683 ;
  assign n33685 = x223 & ~n33684 ;
  assign n33686 = n15141 & ~n33685 ;
  assign n33687 = n16176 & ~n33685 ;
  assign n33688 = n15082 & ~n33685 ;
  assign n33689 = x223 & n2032 ;
  assign n33690 = x642 & n14839 ;
  assign n33691 = n32753 & ~n33690 ;
  assign n33692 = x642 & ~n33143 ;
  assign n33693 = n4707 | n33692 ;
  assign n33694 = n14652 & ~n33693 ;
  assign n33695 = n33691 | n33694 ;
  assign n33696 = x681 & ~n33695 ;
  assign n33697 = n14641 & ~n15027 ;
  assign n33698 = n32749 | n33697 ;
  assign n33699 = ( x681 & n14580 ) | ( x681 & n33698 ) | ( n14580 & n33698 ) ;
  assign n33700 = ( x681 & ~n14580 ) | ( x681 & n33695 ) | ( ~n14580 & n33695 ) ;
  assign n33701 = n33699 | n33700 ;
  assign n33702 = ~n4721 & n33701 ;
  assign n33703 = ~n33696 & n33702 ;
  assign n33704 = x642 & ~n15010 ;
  assign n33705 = x642 | n14614 ;
  assign n33706 = ~n33704 & n33705 ;
  assign n33707 = x681 & ~n33706 ;
  assign n33708 = ~n14580 & n33706 ;
  assign n33709 = n14606 & ~n33690 ;
  assign n33710 = x681 | n33709 ;
  assign n33711 = n33708 | n33710 ;
  assign n33712 = n4721 & n33711 ;
  assign n33713 = ~n33707 & n33712 ;
  assign n33714 = x223 & ~n33713 ;
  assign n33715 = ~n33703 & n33714 ;
  assign n33716 = n15503 & n33690 ;
  assign n33717 = x681 & ~n33716 ;
  assign n33718 = ~n14580 & n33716 ;
  assign n33719 = x642 & n14580 ;
  assign n33720 = n15815 & n33719 ;
  assign n33721 = x681 | n33720 ;
  assign n33722 = n33718 | n33721 ;
  assign n33723 = ~n33717 & n33722 ;
  assign n33724 = x947 & ~n33723 ;
  assign n33725 = x223 | n33724 ;
  assign n33726 = ( x947 & n18919 ) | ( x947 & n33723 ) | ( n18919 & n33723 ) ;
  assign n33727 = x642 & n14874 ;
  assign n33728 = ~n14580 & n33727 ;
  assign n33729 = x681 | n33728 ;
  assign n33730 = n15799 & n33719 ;
  assign n33731 = n33729 | n33730 ;
  assign n33732 = x681 & ~n33727 ;
  assign n33733 = n33731 & ~n33732 ;
  assign n33734 = ( x947 & ~n18919 ) | ( x947 & n33733 ) | ( ~n18919 & n33733 ) ;
  assign n33735 = n33726 | n33734 ;
  assign n33736 = ~n33725 & n33735 ;
  assign n33737 = n2203 & ~n33736 ;
  assign n33738 = ~n33715 & n33737 ;
  assign n33739 = x223 & ~n16705 ;
  assign n33740 = n2203 | n33739 ;
  assign n33741 = n33727 | n33740 ;
  assign n33742 = ~x215 & n33741 ;
  assign n33743 = ~n33738 & n33742 ;
  assign n33744 = n14884 & n33719 ;
  assign n33745 = n33729 | n33744 ;
  assign n33746 = x642 & ~n14959 ;
  assign n33747 = n14580 & ~n33746 ;
  assign n33748 = n14475 & n33747 ;
  assign n33749 = x681 | n33748 ;
  assign n33750 = n14521 | n33749 ;
  assign n33751 = n33745 & n33750 ;
  assign n33752 = x642 & n14876 ;
  assign n33753 = x681 & ~n33752 ;
  assign n33754 = n33751 & ~n33753 ;
  assign n33755 = n18919 & n33754 ;
  assign n33756 = ~n4721 & n33745 ;
  assign n33757 = n33727 & n33756 ;
  assign n33758 = x947 | n33757 ;
  assign n33759 = n33755 | n33758 ;
  assign n33760 = x947 & ~n33754 ;
  assign n33761 = x223 | n33760 ;
  assign n33762 = n33759 & ~n33761 ;
  assign n33763 = x642 | n32737 ;
  assign n33764 = x642 & ~n14961 ;
  assign n33765 = n33763 & ~n33764 ;
  assign n33766 = ~n14580 & n33765 ;
  assign n33767 = n33749 | n33766 ;
  assign n33768 = x681 & ~n33765 ;
  assign n33769 = n33767 & ~n33768 ;
  assign n33770 = ( ~x223 & n4721 ) | ( ~x223 & n33769 ) | ( n4721 & n33769 ) ;
  assign n33771 = n33170 & ~n33692 ;
  assign n33772 = n33691 | n33771 ;
  assign n33773 = x681 & ~n33772 ;
  assign n33774 = ~n14580 & n33772 ;
  assign n33775 = n15756 & ~n33690 ;
  assign n33776 = n14580 & n33775 ;
  assign n33777 = n30485 & n33776 ;
  assign n33778 = x681 | n33777 ;
  assign n33779 = n33774 | n33778 ;
  assign n33780 = ~n33773 & n33779 ;
  assign n33781 = ( x223 & n4721 ) | ( x223 & ~n33780 ) | ( n4721 & ~n33780 ) ;
  assign n33782 = ~n33770 & n33781 ;
  assign n33783 = n33762 | n33782 ;
  assign n33784 = x215 & n33783 ;
  assign n33785 = x299 & ~n33784 ;
  assign n33786 = ~n33743 & n33785 ;
  assign n33787 = n4764 & n33723 ;
  assign n33788 = ( n1823 & n14897 ) | ( n1823 & ~n33733 ) | ( n14897 & ~n33733 ) ;
  assign n33789 = ~n33787 & n33788 ;
  assign n33790 = n1823 | n33727 ;
  assign n33791 = ~x223 & n33790 ;
  assign n33792 = ~n33789 & n33791 ;
  assign n33793 = ~n4764 & n33780 ;
  assign n33794 = ( x223 & n15044 ) | ( x223 & ~n33769 ) | ( n15044 & ~n33769 ) ;
  assign n33795 = ~n33793 & n33794 ;
  assign n33796 = n33792 | n33795 ;
  assign n33797 = ( x39 & n4757 ) | ( x39 & n33796 ) | ( n4757 & n33796 ) ;
  assign n33798 = ~n33786 & n33797 ;
  assign n33799 = ~x223 & x642 ;
  assign n33800 = n16781 & n33799 ;
  assign n33801 = x299 | n33800 ;
  assign n33802 = ~x642 & n16781 ;
  assign n33803 = x223 & ~n33802 ;
  assign n33804 = ~n16779 & n33803 ;
  assign n33805 = n33801 | n33804 ;
  assign n33806 = n14920 & n33799 ;
  assign n33807 = x299 & ~n33806 ;
  assign n33808 = n4706 & n30519 ;
  assign n33809 = x223 & ~n14946 ;
  assign n33810 = ~n33808 & n33809 ;
  assign n33811 = n33807 & ~n33810 ;
  assign n33812 = n33805 & ~n33811 ;
  assign n33813 = ( x38 & ~n9138 ) | ( x38 & n33812 ) | ( ~n9138 & n33812 ) ;
  assign n33814 = n33798 | n33813 ;
  assign n33815 = x39 & x223 ;
  assign n33816 = x38 & ~n33815 ;
  assign n33817 = x223 | n15756 ;
  assign n33818 = ~x39 & n33817 ;
  assign n33819 = ~n33775 & n33818 ;
  assign n33820 = n33816 & ~n33819 ;
  assign n33821 = n2032 | n33820 ;
  assign n33822 = n33814 & ~n33821 ;
  assign n33823 = n33689 | n33822 ;
  assign n33824 = n15082 | n33823 ;
  assign n33825 = ~n33688 & n33824 ;
  assign n33826 = ~x785 & n33825 ;
  assign n33827 = ( x609 & x1155 ) | ( x609 & n33685 ) | ( x1155 & n33685 ) ;
  assign n33828 = ( ~x609 & x1155 ) | ( ~x609 & n33825 ) | ( x1155 & n33825 ) ;
  assign n33829 = n33827 & n33828 ;
  assign n33830 = ( x609 & x1155 ) | ( x609 & ~n33685 ) | ( x1155 & ~n33685 ) ;
  assign n33831 = ( x609 & ~x1155 ) | ( x609 & n33825 ) | ( ~x1155 & n33825 ) ;
  assign n33832 = ~n33830 & n33831 ;
  assign n33833 = n33829 | n33832 ;
  assign n33834 = x785 & n33833 ;
  assign n33835 = n33826 | n33834 ;
  assign n33836 = ~x781 & n33835 ;
  assign n33837 = ( x618 & x1154 ) | ( x618 & n33685 ) | ( x1154 & n33685 ) ;
  assign n33838 = ( ~x618 & x1154 ) | ( ~x618 & n33835 ) | ( x1154 & n33835 ) ;
  assign n33839 = n33837 & n33838 ;
  assign n33840 = ( x618 & x1154 ) | ( x618 & ~n33685 ) | ( x1154 & ~n33685 ) ;
  assign n33841 = ( x618 & ~x1154 ) | ( x618 & n33835 ) | ( ~x1154 & n33835 ) ;
  assign n33842 = ~n33840 & n33841 ;
  assign n33843 = n33839 | n33842 ;
  assign n33844 = x781 & n33843 ;
  assign n33845 = n33836 | n33844 ;
  assign n33846 = ~x789 & n33845 ;
  assign n33847 = ( x619 & x1159 ) | ( x619 & n33685 ) | ( x1159 & n33685 ) ;
  assign n33848 = ( ~x619 & x1159 ) | ( ~x619 & n33845 ) | ( x1159 & n33845 ) ;
  assign n33849 = n33847 & n33848 ;
  assign n33850 = ( x619 & x1159 ) | ( x619 & ~n33685 ) | ( x1159 & ~n33685 ) ;
  assign n33851 = ( x619 & ~x1159 ) | ( x619 & n33845 ) | ( ~x1159 & n33845 ) ;
  assign n33852 = ~n33850 & n33851 ;
  assign n33853 = n33849 | n33852 ;
  assign n33854 = x789 & n33853 ;
  assign n33855 = n33846 | n33854 ;
  assign n33856 = n16176 | n33855 ;
  assign n33857 = ~n33687 & n33856 ;
  assign n33858 = ~n15134 & n33857 ;
  assign n33859 = n15134 & n33685 ;
  assign n33860 = n33858 | n33859 ;
  assign n33861 = n15141 | n33860 ;
  assign n33862 = ~n33686 & n33861 ;
  assign n33863 = ( x644 & x715 ) | ( x644 & ~n33862 ) | ( x715 & ~n33862 ) ;
  assign n33864 = ( x644 & ~x715 ) | ( x644 & n33685 ) | ( ~x715 & n33685 ) ;
  assign n33865 = ~n33863 & n33864 ;
  assign n33866 = x1160 & ~n33865 ;
  assign n33867 = n17213 & ~n33685 ;
  assign n33868 = n15400 & ~n33685 ;
  assign n33869 = x680 & x681 ;
  assign n33870 = x223 & n33265 ;
  assign n33871 = x299 | n33870 ;
  assign n33872 = ( n15356 & ~n33869 ) | ( n15356 & n33871 ) | ( ~n33869 & n33871 ) ;
  assign n33873 = ( x223 & n15356 ) | ( x223 & ~n33871 ) | ( n15356 & ~n33871 ) ;
  assign n33874 = ~n33872 & n33873 ;
  assign n33875 = x39 | n33874 ;
  assign n33876 = x223 & n30752 ;
  assign n33877 = x299 & ~n33876 ;
  assign n33878 = ( ~n15366 & n33869 ) | ( ~n15366 & n33877 ) | ( n33869 & n33877 ) ;
  assign n33879 = ( x223 & n15366 ) | ( x223 & n33877 ) | ( n15366 & n33877 ) ;
  assign n33880 = n33878 & n33879 ;
  assign n33881 = n33875 | n33880 ;
  assign n33882 = x681 & n33278 ;
  assign n33883 = n33740 | n33882 ;
  assign n33884 = x681 & ~n33297 ;
  assign n33885 = ~n4721 & n14666 ;
  assign n33886 = ~n33884 & n33885 ;
  assign n33887 = x681 & ~n33293 ;
  assign n33888 = n4721 & n14617 ;
  assign n33889 = ~n33887 & n33888 ;
  assign n33890 = x223 & ~n33889 ;
  assign n33891 = ~n33886 & n33890 ;
  assign n33892 = x681 & n15175 ;
  assign n33893 = ( x223 & n4721 ) | ( x223 & ~n33892 ) | ( n4721 & ~n33892 ) ;
  assign n33894 = n33284 & n33869 ;
  assign n33895 = ( ~x223 & n4721 ) | ( ~x223 & n33894 ) | ( n4721 & n33894 ) ;
  assign n33896 = ~n33893 & n33895 ;
  assign n33897 = n2203 & ~n33896 ;
  assign n33898 = ~n33891 & n33897 ;
  assign n33899 = n33883 & ~n33898 ;
  assign n33900 = x215 | n33899 ;
  assign n33901 = ~x223 & x681 ;
  assign n33902 = n33338 & n33901 ;
  assign n33903 = x215 & ~n33902 ;
  assign n33904 = n14514 | n14526 ;
  assign n33905 = x681 & ~n15264 ;
  assign n33906 = n33904 & ~n33905 ;
  assign n33907 = ( ~x223 & n4721 ) | ( ~x223 & n33906 ) | ( n4721 & n33906 ) ;
  assign n33908 = x681 & ~n33319 ;
  assign n33909 = n14570 & ~n33908 ;
  assign n33910 = ( x223 & n4721 ) | ( x223 & ~n33909 ) | ( n4721 & ~n33909 ) ;
  assign n33911 = ~n33907 & n33910 ;
  assign n33912 = n33903 & ~n33911 ;
  assign n33913 = x299 & ~n33912 ;
  assign n33914 = n33900 & n33913 ;
  assign n33915 = n1823 | n33882 ;
  assign n33916 = n4764 & n33892 ;
  assign n33917 = ( n1823 & n14897 ) | ( n1823 & ~n33894 ) | ( n14897 & ~n33894 ) ;
  assign n33918 = ~n33916 & n33917 ;
  assign n33919 = n33915 & ~n33918 ;
  assign n33920 = x223 | n33919 ;
  assign n33921 = ( x223 & ~n4764 ) | ( x223 & n33906 ) | ( ~n4764 & n33906 ) ;
  assign n33922 = ( x223 & n4764 ) | ( x223 & n33909 ) | ( n4764 & n33909 ) ;
  assign n33923 = n33921 & n33922 ;
  assign n33924 = n33920 & ~n33923 ;
  assign n33925 = ( x39 & n4757 ) | ( x39 & ~n33924 ) | ( n4757 & ~n33924 ) ;
  assign n33926 = ~n33914 & n33925 ;
  assign n33927 = n33881 & ~n33926 ;
  assign n33928 = x38 | n33927 ;
  assign n33929 = x223 & ~n15070 ;
  assign n33930 = x681 & n15374 ;
  assign n33931 = x38 & ~n33930 ;
  assign n33932 = ~n33929 & n33931 ;
  assign n33933 = n2032 | n33932 ;
  assign n33934 = n33928 & ~n33933 ;
  assign n33935 = n33689 | n33934 ;
  assign n33936 = ~x778 & n33935 ;
  assign n33937 = ( x625 & x1153 ) | ( x625 & n33685 ) | ( x1153 & n33685 ) ;
  assign n33938 = ( ~x625 & x1153 ) | ( ~x625 & n33935 ) | ( x1153 & n33935 ) ;
  assign n33939 = n33937 & n33938 ;
  assign n33940 = ( x625 & x1153 ) | ( x625 & ~n33685 ) | ( x1153 & ~n33685 ) ;
  assign n33941 = ( x625 & ~x1153 ) | ( x625 & n33935 ) | ( ~x1153 & n33935 ) ;
  assign n33942 = ~n33940 & n33941 ;
  assign n33943 = n33939 | n33942 ;
  assign n33944 = x778 & n33943 ;
  assign n33945 = n33936 | n33944 ;
  assign n33946 = n15400 | n33945 ;
  assign n33947 = ~n33868 & n33946 ;
  assign n33948 = ~n15407 & n33947 ;
  assign n33949 = n15407 & n33685 ;
  assign n33950 = n33948 | n33949 ;
  assign n33951 = n15414 | n33950 ;
  assign n33952 = n15421 | n33951 ;
  assign n33953 = ~n33867 & n33952 ;
  assign n33954 = n17220 | n33953 ;
  assign n33955 = n16054 & ~n33685 ;
  assign n33956 = n33954 & ~n33955 ;
  assign n33957 = ~x787 & n33956 ;
  assign n33958 = ( x647 & x1157 ) | ( x647 & n33685 ) | ( x1157 & n33685 ) ;
  assign n33959 = ( ~x647 & x1157 ) | ( ~x647 & n33956 ) | ( x1157 & n33956 ) ;
  assign n33960 = n33958 & n33959 ;
  assign n33961 = ( x647 & x1157 ) | ( x647 & ~n33685 ) | ( x1157 & ~n33685 ) ;
  assign n33962 = ( x647 & ~x1157 ) | ( x647 & n33956 ) | ( ~x1157 & n33956 ) ;
  assign n33963 = ~n33961 & n33962 ;
  assign n33964 = n33960 | n33963 ;
  assign n33965 = x787 & n33964 ;
  assign n33966 = n33957 | n33965 ;
  assign n33967 = ( x644 & x715 ) | ( x644 & n33966 ) | ( x715 & n33966 ) ;
  assign n33968 = n18610 & n33860 ;
  assign n33969 = ( x630 & n33963 ) | ( x630 & n33968 ) | ( n33963 & n33968 ) ;
  assign n33970 = ( ~x630 & n33960 ) | ( ~x630 & n33968 ) | ( n33960 & n33968 ) ;
  assign n33971 = n33969 | n33970 ;
  assign n33972 = x787 & n33971 ;
  assign n33973 = n18621 & n33857 ;
  assign n33974 = x628 | n33685 ;
  assign n33975 = n15131 & n33974 ;
  assign n33976 = x628 & ~n33685 ;
  assign n33977 = n15132 & ~n33976 ;
  assign n33978 = ( x628 & n33953 ) | ( x628 & n33977 ) | ( n33953 & n33977 ) ;
  assign n33979 = x628 & ~n33977 ;
  assign n33980 = ( n33975 & n33978 ) | ( n33975 & ~n33979 ) | ( n33978 & ~n33979 ) ;
  assign n33981 = n33973 | n33980 ;
  assign n33982 = x792 & n33981 ;
  assign n33983 = n15414 & ~n33685 ;
  assign n33984 = n33951 & ~n33983 ;
  assign n33985 = n16115 & ~n33984 ;
  assign n33986 = ( x626 & n15418 ) | ( x626 & ~n33685 ) | ( n15418 & ~n33685 ) ;
  assign n33987 = ( x626 & ~n15418 ) | ( x626 & n33855 ) | ( ~n15418 & n33855 ) ;
  assign n33988 = n33986 & ~n33987 ;
  assign n33989 = n33985 | n33988 ;
  assign n33990 = ( x626 & ~n15419 ) | ( x626 & n33685 ) | ( ~n15419 & n33685 ) ;
  assign n33991 = ( x626 & n15419 ) | ( x626 & ~n33855 ) | ( n15419 & ~n33855 ) ;
  assign n33992 = ~n33990 & n33991 ;
  assign n33993 = n33989 | n33992 ;
  assign n33994 = x788 & n33993 ;
  assign n33995 = x648 & ~n33852 ;
  assign n33996 = ( x619 & x1159 ) | ( x619 & n33950 ) | ( x1159 & n33950 ) ;
  assign n33997 = x627 | n33839 ;
  assign n33998 = ( x618 & x1154 ) | ( x618 & ~n33947 ) | ( x1154 & ~n33947 ) ;
  assign n33999 = x660 | n33829 ;
  assign n34000 = ( x609 & x1155 ) | ( x609 & ~n33945 ) | ( x1155 & ~n33945 ) ;
  assign n34001 = ( x625 & x1153 ) | ( x625 & ~n33823 ) | ( x1153 & ~n33823 ) ;
  assign n34002 = n33696 | n33869 ;
  assign n34003 = ~x642 & n15585 ;
  assign n34004 = x642 & n15705 ;
  assign n34005 = n34003 | n34004 ;
  assign n34006 = n15756 & n34005 ;
  assign n34007 = ~n14479 & n34006 ;
  assign n34008 = n4707 & ~n34007 ;
  assign n34009 = x680 & ~n34008 ;
  assign n34010 = x642 & ~n33432 ;
  assign n34011 = x642 | n15603 ;
  assign n34012 = ~n34010 & n34011 ;
  assign n34013 = n4707 | n34012 ;
  assign n34014 = n34009 & n34013 ;
  assign n34015 = n34002 & ~n34014 ;
  assign n34016 = n33702 & ~n34015 ;
  assign n34017 = n33707 | n33869 ;
  assign n34018 = ~x642 & n4707 ;
  assign n34019 = ~n33411 & n34018 ;
  assign n34020 = n14855 | n33419 ;
  assign n34021 = x642 & ~n33413 ;
  assign n34022 = x680 & ~n34021 ;
  assign n34023 = n34020 & n34022 ;
  assign n34024 = ~n34019 & n34023 ;
  assign n34025 = n34017 & ~n34024 ;
  assign n34026 = n33712 & ~n34025 ;
  assign n34027 = x223 & ~n34026 ;
  assign n34028 = ~n34016 & n34027 ;
  assign n34029 = n2203 & ~n34028 ;
  assign n34030 = n33717 | n33869 ;
  assign n34031 = ~n15502 & n34018 ;
  assign n34032 = x642 & ~n33443 ;
  assign n34033 = x680 & ~n34032 ;
  assign n34034 = n15513 & n34033 ;
  assign n34035 = ~n34031 & n34034 ;
  assign n34036 = n34030 & ~n34035 ;
  assign n34037 = n33722 & ~n34036 ;
  assign n34038 = ( x223 & n4721 ) | ( x223 & ~n34037 ) | ( n4721 & ~n34037 ) ;
  assign n34039 = x680 | n33727 ;
  assign n34040 = n15585 & ~n34010 ;
  assign n34041 = n32753 & ~n34040 ;
  assign n34042 = x680 & ~n34041 ;
  assign n34043 = x642 & ~n33453 ;
  assign n34044 = n4707 | n34043 ;
  assign n34045 = x642 | n15549 ;
  assign n34046 = ~n34044 & n34045 ;
  assign n34047 = n34042 & ~n34046 ;
  assign n34048 = n34039 & ~n34047 ;
  assign n34049 = x681 & ~n34048 ;
  assign n34050 = n33731 & ~n34049 ;
  assign n34051 = ( ~x223 & n4721 ) | ( ~x223 & n34050 ) | ( n4721 & n34050 ) ;
  assign n34052 = ~n34038 & n34051 ;
  assign n34053 = n34029 & ~n34052 ;
  assign n34054 = n33690 & ~n33869 ;
  assign n34055 = n33869 & ~n34003 ;
  assign n34056 = ~n33576 & n34055 ;
  assign n34057 = n34054 | n34056 ;
  assign n34058 = n16705 & n34057 ;
  assign n34059 = ~x223 & n34058 ;
  assign n34060 = ( ~x223 & n33869 ) | ( ~x223 & n34006 ) | ( n33869 & n34006 ) ;
  assign n34061 = ( x223 & ~n33775 ) | ( x223 & n33869 ) | ( ~n33775 & n33869 ) ;
  assign n34062 = ~n34060 & n34061 ;
  assign n34063 = n33740 | n34062 ;
  assign n34064 = n34059 | n34063 ;
  assign n34065 = ~x215 & n34064 ;
  assign n34066 = ~n34053 & n34065 ;
  assign n34067 = n33753 | n33869 ;
  assign n34068 = n15487 & n15848 ;
  assign n34069 = n14855 | n34068 ;
  assign n34070 = x642 & ~n33480 ;
  assign n34071 = ~n15467 & n34018 ;
  assign n34072 = x680 & ~n34071 ;
  assign n34073 = ~n34070 & n34072 ;
  assign n34074 = n34069 & n34073 ;
  assign n34075 = n34067 & ~n34074 ;
  assign n34076 = n4721 & n33751 ;
  assign n34077 = ~n34075 & n34076 ;
  assign n34078 = n15470 & ~n34044 ;
  assign n34079 = n34042 & ~n34078 ;
  assign n34080 = n34039 & ~n34079 ;
  assign n34081 = x681 & ~n34080 ;
  assign n34082 = n33756 & ~n34081 ;
  assign n34083 = x223 | n34082 ;
  assign n34084 = n34077 | n34083 ;
  assign n34085 = x215 & n34084 ;
  assign n34086 = ~x680 & n33765 ;
  assign n34087 = n14876 | n15643 ;
  assign n34088 = n4707 & ~n34087 ;
  assign n34089 = x642 & ~n33500 ;
  assign n34090 = x680 & n15641 ;
  assign n34091 = ~n34089 & n34090 ;
  assign n34092 = ~n34088 & n34091 ;
  assign n34093 = x681 & ~n34092 ;
  assign n34094 = ~n34086 & n34093 ;
  assign n34095 = n33767 & ~n34094 ;
  assign n34096 = ( x223 & ~n4721 ) | ( x223 & n34095 ) | ( ~n4721 & n34095 ) ;
  assign n34097 = n33773 | n33869 ;
  assign n34098 = x614 | n15667 ;
  assign n34099 = ~n34010 & n34098 ;
  assign n34100 = x616 | n34099 ;
  assign n34101 = n34009 & n34100 ;
  assign n34102 = n34097 & ~n34101 ;
  assign n34103 = n33779 & ~n34102 ;
  assign n34104 = ( x223 & n4721 ) | ( x223 & n34103 ) | ( n4721 & n34103 ) ;
  assign n34105 = n34096 & n34104 ;
  assign n34106 = n34085 & ~n34105 ;
  assign n34107 = x299 & ~n34106 ;
  assign n34108 = ~n34066 & n34107 ;
  assign n34109 = ~n4764 & n34050 ;
  assign n34110 = ( n1823 & n15052 ) | ( n1823 & ~n34037 ) | ( n15052 & ~n34037 ) ;
  assign n34111 = ~n34109 & n34110 ;
  assign n34112 = n1823 | n34058 ;
  assign n34113 = ~x223 & n34112 ;
  assign n34114 = ~n34111 & n34113 ;
  assign n34115 = ~n4764 & n34103 ;
  assign n34116 = ( x223 & n15044 ) | ( x223 & ~n34095 ) | ( n15044 & ~n34095 ) ;
  assign n34117 = ~n34115 & n34116 ;
  assign n34118 = n34114 | n34117 ;
  assign n34119 = ( x39 & n4757 ) | ( x39 & n34118 ) | ( n4757 & n34118 ) ;
  assign n34120 = ~n34108 & n34119 ;
  assign n34121 = n15885 & ~n33869 ;
  assign n34122 = x223 & ~n33808 ;
  assign n34123 = ~n33549 & n34122 ;
  assign n34124 = ~n34121 & n34123 ;
  assign n34125 = n16998 & n33901 ;
  assign n34126 = n33807 & ~n34125 ;
  assign n34127 = ~n34124 & n34126 ;
  assign n34128 = n15881 & ~n33869 ;
  assign n34129 = ~n33567 & n33803 ;
  assign n34130 = ~n34128 & n34129 ;
  assign n34131 = n16990 & n33901 ;
  assign n34132 = n33801 | n34131 ;
  assign n34133 = n34130 | n34132 ;
  assign n34134 = ~n34127 & n34133 ;
  assign n34135 = ( x38 & ~n9138 ) | ( x38 & n34134 ) | ( ~n9138 & n34134 ) ;
  assign n34136 = n34120 | n34135 ;
  assign n34137 = n34057 | n34062 ;
  assign n34138 = n33818 & n34137 ;
  assign n34139 = n33816 & ~n34138 ;
  assign n34140 = n2032 | n34139 ;
  assign n34141 = n34136 & ~n34140 ;
  assign n34142 = n33689 | n34141 ;
  assign n34143 = ( x625 & ~x1153 ) | ( x625 & n34142 ) | ( ~x1153 & n34142 ) ;
  assign n34144 = ~n34001 & n34143 ;
  assign n34145 = x608 | n34144 ;
  assign n34146 = n33939 | n34145 ;
  assign n34147 = ( x625 & x1153 ) | ( x625 & n33823 ) | ( x1153 & n33823 ) ;
  assign n34148 = ( ~x625 & x1153 ) | ( ~x625 & n34142 ) | ( x1153 & n34142 ) ;
  assign n34149 = n34147 & n34148 ;
  assign n34150 = x608 & ~n34149 ;
  assign n34151 = ~n33942 & n34150 ;
  assign n34152 = n34146 & ~n34151 ;
  assign n34153 = x778 & ~n34152 ;
  assign n34154 = x778 | n34142 ;
  assign n34155 = ~n34153 & n34154 ;
  assign n34156 = ( x609 & ~x1155 ) | ( x609 & n34155 ) | ( ~x1155 & n34155 ) ;
  assign n34157 = ~n34000 & n34156 ;
  assign n34158 = n33999 | n34157 ;
  assign n34159 = x660 & ~n33832 ;
  assign n34160 = ( x609 & x1155 ) | ( x609 & n33945 ) | ( x1155 & n33945 ) ;
  assign n34161 = ( ~x609 & x1155 ) | ( ~x609 & n34155 ) | ( x1155 & n34155 ) ;
  assign n34162 = n34160 & n34161 ;
  assign n34163 = n34159 & ~n34162 ;
  assign n34164 = n34158 & ~n34163 ;
  assign n34165 = x785 & ~n34164 ;
  assign n34166 = x785 | n34155 ;
  assign n34167 = ~n34165 & n34166 ;
  assign n34168 = ( x618 & ~x1154 ) | ( x618 & n34167 ) | ( ~x1154 & n34167 ) ;
  assign n34169 = ~n33998 & n34168 ;
  assign n34170 = n33997 | n34169 ;
  assign n34171 = x627 & ~n33842 ;
  assign n34172 = ( x618 & x1154 ) | ( x618 & n33947 ) | ( x1154 & n33947 ) ;
  assign n34173 = ( ~x618 & x1154 ) | ( ~x618 & n34167 ) | ( x1154 & n34167 ) ;
  assign n34174 = n34172 & n34173 ;
  assign n34175 = n34171 & ~n34174 ;
  assign n34176 = n34170 & ~n34175 ;
  assign n34177 = x781 & ~n34176 ;
  assign n34178 = x781 | n34167 ;
  assign n34179 = ~n34177 & n34178 ;
  assign n34180 = ( ~x619 & x1159 ) | ( ~x619 & n34179 ) | ( x1159 & n34179 ) ;
  assign n34181 = n33996 & n34180 ;
  assign n34182 = n33995 & ~n34181 ;
  assign n34183 = x648 | n33849 ;
  assign n34184 = ( x619 & x1159 ) | ( x619 & ~n33950 ) | ( x1159 & ~n33950 ) ;
  assign n34185 = ( x619 & ~x1159 ) | ( x619 & n34179 ) | ( ~x1159 & n34179 ) ;
  assign n34186 = ~n34184 & n34185 ;
  assign n34187 = n34183 | n34186 ;
  assign n34188 = x789 & n34187 ;
  assign n34189 = ~n34182 & n34188 ;
  assign n34190 = ~x789 & n34179 ;
  assign n34191 = n16177 | n34190 ;
  assign n34192 = n34189 | n34191 ;
  assign n34193 = ~n33994 & n34192 ;
  assign n34194 = n33982 | n34193 ;
  assign n34195 = ( n18431 & n22573 ) | ( n18431 & ~n33981 ) | ( n22573 & ~n33981 ) ;
  assign n34196 = n34194 & ~n34195 ;
  assign n34197 = n33972 | n34196 ;
  assign n34198 = ( ~x644 & x715 ) | ( ~x644 & n34197 ) | ( x715 & n34197 ) ;
  assign n34199 = n33967 & n34198 ;
  assign n34200 = n33866 & ~n34199 ;
  assign n34201 = ( x644 & x715 ) | ( x644 & n33862 ) | ( x715 & n33862 ) ;
  assign n34202 = ( ~x644 & x715 ) | ( ~x644 & n33685 ) | ( x715 & n33685 ) ;
  assign n34203 = n34201 & n34202 ;
  assign n34204 = x1160 | n34203 ;
  assign n34205 = ( x644 & x715 ) | ( x644 & ~n33966 ) | ( x715 & ~n33966 ) ;
  assign n34206 = ( x644 & ~x715 ) | ( x644 & n34197 ) | ( ~x715 & n34197 ) ;
  assign n34207 = ~n34205 & n34206 ;
  assign n34208 = n34204 | n34207 ;
  assign n34209 = ~n34200 & n34208 ;
  assign n34210 = ( x790 & n6785 ) | ( x790 & n34209 ) | ( n6785 & n34209 ) ;
  assign n34211 = ( ~x790 & n6785 ) | ( ~x790 & n34197 ) | ( n6785 & n34197 ) ;
  assign n34212 = n34210 | n34211 ;
  assign n34213 = ~n33678 & n34212 ;
  assign n34214 = ~x224 & n6785 ;
  assign n34215 = x224 & ~n33106 ;
  assign n34216 = n15141 & ~n34215 ;
  assign n34217 = n16176 & ~n34215 ;
  assign n34218 = x224 & n2032 ;
  assign n34219 = x614 & n33156 ;
  assign n34220 = ~x224 & n34219 ;
  assign n34221 = ~n14900 & n34220 ;
  assign n34222 = x223 & ~n34221 ;
  assign n34223 = x614 & ~n14961 ;
  assign n34224 = n32864 & ~n34223 ;
  assign n34225 = x680 | n34224 ;
  assign n34226 = x680 & ~n14964 ;
  assign n34227 = ~n32866 & n34226 ;
  assign n34228 = n34225 & ~n34227 ;
  assign n34229 = n14553 | n34228 ;
  assign n34230 = n14553 & ~n34224 ;
  assign n34231 = n34229 & ~n34230 ;
  assign n34232 = ( ~x224 & n4764 ) | ( ~x224 & n34231 ) | ( n4764 & n34231 ) ;
  assign n34233 = x614 & n14839 ;
  assign n34234 = n16705 & ~n34233 ;
  assign n34235 = n4708 | n34234 ;
  assign n34236 = n33169 & n34235 ;
  assign n34237 = n14553 & ~n34236 ;
  assign n34238 = x680 | n34236 ;
  assign n34239 = x680 & n34233 ;
  assign n34240 = n14534 | n34239 ;
  assign n34241 = n34238 & ~n34240 ;
  assign n34242 = n14553 | n34241 ;
  assign n34243 = ~n34237 & n34242 ;
  assign n34244 = ( x224 & n4764 ) | ( x224 & ~n34243 ) | ( n4764 & ~n34243 ) ;
  assign n34245 = ~n34232 & n34244 ;
  assign n34246 = n34222 & ~n34245 ;
  assign n34247 = ~n14481 & n14891 ;
  assign n34248 = x614 & n34247 ;
  assign n34249 = x223 | n34248 ;
  assign n34250 = x614 & n33125 ;
  assign n34251 = ( n4346 & n4764 ) | ( n4346 & n34250 ) | ( n4764 & n34250 ) ;
  assign n34252 = x614 & n15815 ;
  assign n34253 = x680 & ~n34252 ;
  assign n34254 = n15503 & n34233 ;
  assign n34255 = x680 | n34254 ;
  assign n34256 = ~n34253 & n34255 ;
  assign n34257 = n14553 | n34256 ;
  assign n34258 = n14553 & ~n34254 ;
  assign n34259 = n34257 & ~n34258 ;
  assign n34260 = ( n4346 & ~n4764 ) | ( n4346 & n34259 ) | ( ~n4764 & n34259 ) ;
  assign n34261 = n34251 & n34260 ;
  assign n34262 = n34249 | n34261 ;
  assign n34263 = n14486 & n14652 ;
  assign n34264 = n4713 & n34263 ;
  assign n34265 = n4707 | n14609 ;
  assign n34266 = n34264 | n34265 ;
  assign n34267 = x614 & ~n15010 ;
  assign n34268 = ~x614 & x616 ;
  assign n34269 = ~n15503 & n34268 ;
  assign n34270 = n34267 | n34269 ;
  assign n34271 = n34266 & ~n34270 ;
  assign n34272 = n14553 & ~n34271 ;
  assign n34273 = x680 | n34271 ;
  assign n34274 = ~n30540 & n34253 ;
  assign n34275 = n34239 | n34274 ;
  assign n34276 = n34273 & ~n34275 ;
  assign n34277 = n14553 | n34276 ;
  assign n34278 = ~n34272 & n34277 ;
  assign n34279 = ( ~x224 & n4764 ) | ( ~x224 & n34278 ) | ( n4764 & n34278 ) ;
  assign n34280 = n33142 & n34235 ;
  assign n34281 = n14553 & ~n34280 ;
  assign n34282 = x680 | n34280 ;
  assign n34283 = n32789 | n34239 ;
  assign n34284 = n34282 & ~n34283 ;
  assign n34285 = n14553 | n34284 ;
  assign n34286 = ~n34281 & n34285 ;
  assign n34287 = ( x224 & n4764 ) | ( x224 & ~n34286 ) | ( n4764 & ~n34286 ) ;
  assign n34288 = ~n34279 & n34287 ;
  assign n34289 = n34262 | n34288 ;
  assign n34290 = ~n34246 & n34289 ;
  assign n34291 = x299 | n34290 ;
  assign n34292 = ( x224 & n4721 ) | ( x224 & ~n34259 ) | ( n4721 & ~n34259 ) ;
  assign n34293 = ( ~x224 & n4721 ) | ( ~x224 & n34250 ) | ( n4721 & n34250 ) ;
  assign n34294 = ~n34292 & n34293 ;
  assign n34295 = n2203 & ~n34294 ;
  assign n34296 = ( ~x224 & n4721 ) | ( ~x224 & n34278 ) | ( n4721 & n34278 ) ;
  assign n34297 = ( x224 & n4721 ) | ( x224 & ~n34286 ) | ( n4721 & ~n34286 ) ;
  assign n34298 = ~n34296 & n34297 ;
  assign n34299 = n34295 & ~n34298 ;
  assign n34300 = x224 & ~n16705 ;
  assign n34301 = n2203 | n34300 ;
  assign n34302 = ~n14481 & n14625 ;
  assign n34303 = n14839 & n34302 ;
  assign n34304 = n34301 | n34303 ;
  assign n34305 = ~x215 & n34304 ;
  assign n34306 = ~n34299 & n34305 ;
  assign n34307 = ~n14873 & n34220 ;
  assign n34308 = ( ~x224 & n4721 ) | ( ~x224 & n34231 ) | ( n4721 & n34231 ) ;
  assign n34309 = ( x224 & n4721 ) | ( x224 & ~n34243 ) | ( n4721 & ~n34243 ) ;
  assign n34310 = ~n34308 & n34309 ;
  assign n34311 = n34307 | n34310 ;
  assign n34312 = x215 & n34311 ;
  assign n34313 = x299 & ~n34312 ;
  assign n34314 = ~n34306 & n34313 ;
  assign n34315 = x39 & ~n34314 ;
  assign n34316 = n34291 & n34315 ;
  assign n34317 = x614 & n14920 ;
  assign n34318 = x224 & n30517 ;
  assign n34319 = n34317 & ~n34318 ;
  assign n34320 = x224 & ~n14814 ;
  assign n34321 = n34319 | n34320 ;
  assign n34322 = x299 & ~n34321 ;
  assign n34323 = ~x614 & n16781 ;
  assign n34324 = x224 & ~n34323 ;
  assign n34325 = ~n16779 & n34324 ;
  assign n34326 = x614 & n16781 ;
  assign n34327 = ~x224 & n34326 ;
  assign n34328 = x299 | n34327 ;
  assign n34329 = n34325 | n34328 ;
  assign n34330 = ~n34322 & n34329 ;
  assign n34331 = ( x38 & ~n9138 ) | ( x38 & n34330 ) | ( ~n9138 & n34330 ) ;
  assign n34332 = n34316 | n34331 ;
  assign n34333 = x224 & ~n15070 ;
  assign n34334 = x38 & ~n34333 ;
  assign n34335 = x614 & n15072 ;
  assign n34336 = n34334 & ~n34335 ;
  assign n34337 = n2032 | n34336 ;
  assign n34338 = n34332 & ~n34337 ;
  assign n34339 = n34218 | n34338 ;
  assign n34340 = ~n15082 & n34339 ;
  assign n34341 = n15082 & n34215 ;
  assign n34342 = n34340 | n34341 ;
  assign n34343 = ~x785 & n34342 ;
  assign n34344 = ( x609 & x1155 ) | ( x609 & n34215 ) | ( x1155 & n34215 ) ;
  assign n34345 = ( ~x609 & x1155 ) | ( ~x609 & n34342 ) | ( x1155 & n34342 ) ;
  assign n34346 = n34344 & n34345 ;
  assign n34347 = ( x609 & x1155 ) | ( x609 & ~n34215 ) | ( x1155 & ~n34215 ) ;
  assign n34348 = ( x609 & ~x1155 ) | ( x609 & n34342 ) | ( ~x1155 & n34342 ) ;
  assign n34349 = ~n34347 & n34348 ;
  assign n34350 = n34346 | n34349 ;
  assign n34351 = x785 & n34350 ;
  assign n34352 = n34343 | n34351 ;
  assign n34353 = ~x781 & n34352 ;
  assign n34354 = ( x618 & x1154 ) | ( x618 & n34215 ) | ( x1154 & n34215 ) ;
  assign n34355 = ( ~x618 & x1154 ) | ( ~x618 & n34352 ) | ( x1154 & n34352 ) ;
  assign n34356 = n34354 & n34355 ;
  assign n34357 = ( x618 & x1154 ) | ( x618 & ~n34215 ) | ( x1154 & ~n34215 ) ;
  assign n34358 = ( x618 & ~x1154 ) | ( x618 & n34352 ) | ( ~x1154 & n34352 ) ;
  assign n34359 = ~n34357 & n34358 ;
  assign n34360 = n34356 | n34359 ;
  assign n34361 = x781 & n34360 ;
  assign n34362 = n34353 | n34361 ;
  assign n34363 = ~x789 & n34362 ;
  assign n34364 = ( x619 & x1159 ) | ( x619 & n34215 ) | ( x1159 & n34215 ) ;
  assign n34365 = ( ~x619 & x1159 ) | ( ~x619 & n34362 ) | ( x1159 & n34362 ) ;
  assign n34366 = n34364 & n34365 ;
  assign n34367 = ( x619 & x1159 ) | ( x619 & ~n34215 ) | ( x1159 & ~n34215 ) ;
  assign n34368 = ( x619 & ~x1159 ) | ( x619 & n34362 ) | ( ~x1159 & n34362 ) ;
  assign n34369 = ~n34367 & n34368 ;
  assign n34370 = n34366 | n34369 ;
  assign n34371 = x789 & n34370 ;
  assign n34372 = n34363 | n34371 ;
  assign n34373 = n16176 | n34372 ;
  assign n34374 = ~n34217 & n34373 ;
  assign n34375 = ~n15134 & n34374 ;
  assign n34376 = n15134 & n34215 ;
  assign n34377 = n34375 | n34376 ;
  assign n34378 = n15141 | n34377 ;
  assign n34379 = ~n34216 & n34378 ;
  assign n34380 = ( x644 & x715 ) | ( x644 & ~n34379 ) | ( x715 & ~n34379 ) ;
  assign n34381 = ( x644 & ~x715 ) | ( x644 & n34215 ) | ( ~x715 & n34215 ) ;
  assign n34382 = ~n34380 & n34381 ;
  assign n34383 = x1160 & ~n34382 ;
  assign n34384 = n17213 & ~n34215 ;
  assign n34385 = x224 & n33265 ;
  assign n34386 = x299 | n34385 ;
  assign n34387 = ( ~n15159 & n15356 ) | ( ~n15159 & n34386 ) | ( n15356 & n34386 ) ;
  assign n34388 = ( x224 & n15356 ) | ( x224 & ~n34386 ) | ( n15356 & ~n34386 ) ;
  assign n34389 = ~n34387 & n34388 ;
  assign n34390 = x39 | n34389 ;
  assign n34391 = x224 & n30752 ;
  assign n34392 = x299 & ~n34391 ;
  assign n34393 = ( n15159 & ~n15366 ) | ( n15159 & n34392 ) | ( ~n15366 & n34392 ) ;
  assign n34394 = ( x224 & n15366 ) | ( x224 & n34392 ) | ( n15366 & n34392 ) ;
  assign n34395 = n34393 & n34394 ;
  assign n34396 = n34390 | n34395 ;
  assign n34397 = n15151 & n15159 ;
  assign n34398 = n34301 | n34397 ;
  assign n34399 = x662 & n15175 ;
  assign n34400 = ( x224 & n4721 ) | ( x224 & ~n34399 ) | ( n4721 & ~n34399 ) ;
  assign n34401 = n15159 & n33284 ;
  assign n34402 = ( ~x224 & n4721 ) | ( ~x224 & n34401 ) | ( n4721 & n34401 ) ;
  assign n34403 = ~n34400 & n34402 ;
  assign n34404 = n2203 & ~n34403 ;
  assign n34405 = n4709 | n33293 ;
  assign n34406 = n16709 & n34405 ;
  assign n34407 = ( ~x224 & n4721 ) | ( ~x224 & n34406 ) | ( n4721 & n34406 ) ;
  assign n34408 = x662 & ~n33297 ;
  assign n34409 = x662 | n16712 ;
  assign n34410 = ~n34408 & n34409 ;
  assign n34411 = ( x224 & n4721 ) | ( x224 & ~n34410 ) | ( n4721 & ~n34410 ) ;
  assign n34412 = ~n34407 & n34411 ;
  assign n34413 = n34404 & ~n34412 ;
  assign n34414 = n34398 & ~n34413 ;
  assign n34415 = x215 | n34414 ;
  assign n34416 = ~x224 & x662 ;
  assign n34417 = n33338 & n34416 ;
  assign n34418 = x215 & ~n34417 ;
  assign n34419 = x662 | n14528 ;
  assign n34420 = x662 & ~n15264 ;
  assign n34421 = n34419 & ~n34420 ;
  assign n34422 = ( ~x224 & n4721 ) | ( ~x224 & n34421 ) | ( n4721 & n34421 ) ;
  assign n34423 = x662 | n16719 ;
  assign n34424 = x662 & ~n33319 ;
  assign n34425 = n34423 & ~n34424 ;
  assign n34426 = ( x224 & n4721 ) | ( x224 & ~n34425 ) | ( n4721 & ~n34425 ) ;
  assign n34427 = ~n34422 & n34426 ;
  assign n34428 = n34418 & ~n34427 ;
  assign n34429 = x299 & ~n34428 ;
  assign n34430 = n34415 & n34429 ;
  assign n34431 = x662 & n15173 ;
  assign n34432 = x223 | n34431 ;
  assign n34433 = ( n4346 & ~n4764 ) | ( n4346 & n34399 ) | ( ~n4764 & n34399 ) ;
  assign n34434 = ( n4346 & n4764 ) | ( n4346 & n34401 ) | ( n4764 & n34401 ) ;
  assign n34435 = n34433 & n34434 ;
  assign n34436 = n34432 | n34435 ;
  assign n34437 = ( ~x224 & n4764 ) | ( ~x224 & n34406 ) | ( n4764 & n34406 ) ;
  assign n34438 = ( x224 & n4764 ) | ( x224 & ~n34410 ) | ( n4764 & ~n34410 ) ;
  assign n34439 = ~n34437 & n34438 ;
  assign n34440 = n34436 | n34439 ;
  assign n34441 = n33308 & n34416 ;
  assign n34442 = x223 & ~n34441 ;
  assign n34443 = ( ~x224 & n4764 ) | ( ~x224 & n34421 ) | ( n4764 & n34421 ) ;
  assign n34444 = ( x224 & n4764 ) | ( x224 & ~n34425 ) | ( n4764 & ~n34425 ) ;
  assign n34445 = ~n34443 & n34444 ;
  assign n34446 = n34442 & ~n34445 ;
  assign n34447 = n34440 & ~n34446 ;
  assign n34448 = ( x39 & n4757 ) | ( x39 & ~n34447 ) | ( n4757 & ~n34447 ) ;
  assign n34449 = ~n34430 & n34448 ;
  assign n34450 = n34396 & ~n34449 ;
  assign n34451 = x38 | n34450 ;
  assign n34452 = x662 & n15374 ;
  assign n34453 = n34334 & ~n34452 ;
  assign n34454 = n2032 | n34453 ;
  assign n34455 = n34451 & ~n34454 ;
  assign n34456 = n34218 | n34455 ;
  assign n34457 = ~x778 & n34456 ;
  assign n34458 = ( x625 & x1153 ) | ( x625 & n34215 ) | ( x1153 & n34215 ) ;
  assign n34459 = ( ~x625 & x1153 ) | ( ~x625 & n34456 ) | ( x1153 & n34456 ) ;
  assign n34460 = n34458 & n34459 ;
  assign n34461 = ( x625 & x1153 ) | ( x625 & ~n34215 ) | ( x1153 & ~n34215 ) ;
  assign n34462 = ( x625 & ~x1153 ) | ( x625 & n34456 ) | ( ~x1153 & n34456 ) ;
  assign n34463 = ~n34461 & n34462 ;
  assign n34464 = n34460 | n34463 ;
  assign n34465 = x778 & n34464 ;
  assign n34466 = n34457 | n34465 ;
  assign n34467 = ~n15400 & n34466 ;
  assign n34468 = n15400 & n34215 ;
  assign n34469 = n34467 | n34468 ;
  assign n34470 = ~n15407 & n34469 ;
  assign n34471 = n15407 & n34215 ;
  assign n34472 = n34470 | n34471 ;
  assign n34473 = n15414 | n34472 ;
  assign n34474 = n15421 | n34473 ;
  assign n34475 = ~n34384 & n34474 ;
  assign n34476 = n17220 | n34475 ;
  assign n34477 = n16054 & ~n34215 ;
  assign n34478 = n34476 & ~n34477 ;
  assign n34479 = ~x787 & n34478 ;
  assign n34480 = ( x647 & x1157 ) | ( x647 & n34215 ) | ( x1157 & n34215 ) ;
  assign n34481 = ( ~x647 & x1157 ) | ( ~x647 & n34478 ) | ( x1157 & n34478 ) ;
  assign n34482 = n34480 & n34481 ;
  assign n34483 = ( x647 & x1157 ) | ( x647 & ~n34215 ) | ( x1157 & ~n34215 ) ;
  assign n34484 = ( x647 & ~x1157 ) | ( x647 & n34478 ) | ( ~x1157 & n34478 ) ;
  assign n34485 = ~n34483 & n34484 ;
  assign n34486 = n34482 | n34485 ;
  assign n34487 = x787 & n34486 ;
  assign n34488 = n34479 | n34487 ;
  assign n34489 = ( x644 & x715 ) | ( x644 & n34488 ) | ( x715 & n34488 ) ;
  assign n34490 = n18621 & n34374 ;
  assign n34491 = x628 | n34215 ;
  assign n34492 = n15131 & n34491 ;
  assign n34493 = x628 & ~n34215 ;
  assign n34494 = n15132 & ~n34493 ;
  assign n34495 = ( x628 & n34475 ) | ( x628 & n34494 ) | ( n34475 & n34494 ) ;
  assign n34496 = x628 & ~n34494 ;
  assign n34497 = ( n34492 & n34495 ) | ( n34492 & ~n34496 ) | ( n34495 & ~n34496 ) ;
  assign n34498 = n34490 | n34497 ;
  assign n34499 = x792 & n34498 ;
  assign n34500 = x648 & ~n34369 ;
  assign n34501 = ( x619 & x1159 ) | ( x619 & n34472 ) | ( x1159 & n34472 ) ;
  assign n34502 = x627 | n34356 ;
  assign n34503 = ( x618 & x1154 ) | ( x618 & ~n34469 ) | ( x1154 & ~n34469 ) ;
  assign n34504 = x660 | n34346 ;
  assign n34505 = ( x609 & x1155 ) | ( x609 & ~n34466 ) | ( x1155 & ~n34466 ) ;
  assign n34506 = x608 | n34460 ;
  assign n34507 = ( x625 & x1153 ) | ( x625 & ~n34339 ) | ( x1153 & ~n34339 ) ;
  assign n34508 = ~n33472 & n34268 ;
  assign n34509 = n33454 | n34508 ;
  assign n34510 = x680 & n34509 ;
  assign n34511 = n33456 | n34303 ;
  assign n34512 = ~n34510 & n34511 ;
  assign n34513 = x662 & ~n34512 ;
  assign n34514 = x662 | n34250 ;
  assign n34515 = ~n34513 & n34514 ;
  assign n34516 = ( x224 & ~n4721 ) | ( x224 & n34515 ) | ( ~n4721 & n34515 ) ;
  assign n34517 = x614 | n22085 ;
  assign n34518 = x614 & ~n33576 ;
  assign n34519 = n34517 & ~n34518 ;
  assign n34520 = ~n14479 & n34519 ;
  assign n34521 = x616 & ~n34520 ;
  assign n34522 = x614 & ~n33432 ;
  assign n34523 = ( n15603 & n15610 ) | ( n15603 & ~n15620 ) | ( n15610 & ~n15620 ) ;
  assign n34524 = ~n34522 & n34523 ;
  assign n34525 = x616 | n34524 ;
  assign n34526 = ~n34521 & n34525 ;
  assign n34527 = x680 & ~n34526 ;
  assign n34528 = n34282 & ~n34527 ;
  assign n34529 = x662 & ~n34528 ;
  assign n34530 = ~x662 & n4710 ;
  assign n34531 = ~n34280 & n34530 ;
  assign n34532 = n34285 & ~n34531 ;
  assign n34533 = ~n34529 & n34532 ;
  assign n34534 = ( x224 & n4721 ) | ( x224 & n34533 ) | ( n4721 & n34533 ) ;
  assign n34535 = n34516 & ~n34534 ;
  assign n34536 = n2203 & ~n34535 ;
  assign n34537 = x614 & ~n33413 ;
  assign n34538 = ~n33411 & n34268 ;
  assign n34539 = n34537 | n34538 ;
  assign n34540 = n33422 & ~n34539 ;
  assign n34541 = x680 & ~n34540 ;
  assign n34542 = n34273 & ~n34541 ;
  assign n34543 = x662 & ~n34542 ;
  assign n34544 = ~n34271 & n34530 ;
  assign n34545 = n34277 & ~n34544 ;
  assign n34546 = ~n34543 & n34545 ;
  assign n34547 = ( x224 & ~n4721 ) | ( x224 & n34546 ) | ( ~n4721 & n34546 ) ;
  assign n34548 = n15520 & ~n15524 ;
  assign n34549 = ( x614 & x680 ) | ( x614 & ~n34548 ) | ( x680 & ~n34548 ) ;
  assign n34550 = ( x614 & ~x680 ) | ( x614 & n33443 ) | ( ~x680 & n33443 ) ;
  assign n34551 = n34549 & ~n34550 ;
  assign n34552 = n34255 & ~n34551 ;
  assign n34553 = x662 & ~n34552 ;
  assign n34554 = ~n34254 & n34530 ;
  assign n34555 = n34257 & ~n34554 ;
  assign n34556 = ~n34553 & n34555 ;
  assign n34557 = ( x224 & n4721 ) | ( x224 & n34556 ) | ( n4721 & n34556 ) ;
  assign n34558 = ~n34547 & n34557 ;
  assign n34559 = n34536 & ~n34558 ;
  assign n34560 = n15159 & n33472 ;
  assign n34561 = n34303 | n34560 ;
  assign n34562 = ~x224 & n34561 ;
  assign n34563 = n15159 & n34519 ;
  assign n34564 = n15159 | n34233 ;
  assign n34565 = n15756 & ~n34564 ;
  assign n34566 = x224 & ~n34565 ;
  assign n34567 = ~n34563 & n34566 ;
  assign n34568 = n34301 | n34567 ;
  assign n34569 = n34562 | n34568 ;
  assign n34570 = ~x215 & n34569 ;
  assign n34571 = ~n34559 & n34570 ;
  assign n34572 = n14521 & n34219 ;
  assign n34573 = x662 | n34572 ;
  assign n34574 = ( ~x614 & x680 ) | ( ~x614 & n33480 ) | ( x680 & n33480 ) ;
  assign n34575 = ( x614 & x680 ) | ( x614 & ~n15476 ) | ( x680 & ~n15476 ) ;
  assign n34576 = n34574 & n34575 ;
  assign n34577 = n15472 & n34576 ;
  assign n34578 = x614 & n14876 ;
  assign n34579 = ( x662 & n15159 ) | ( x662 & ~n34578 ) | ( n15159 & ~n34578 ) ;
  assign n34580 = ~n34577 & n34579 ;
  assign n34581 = n34573 & ~n34580 ;
  assign n34582 = ( x224 & n4721 ) | ( x224 & n34581 ) | ( n4721 & n34581 ) ;
  assign n34583 = ( x616 & n14988 ) | ( x616 & ~n15489 ) | ( n14988 & ~n15489 ) ;
  assign n34584 = x680 & n34583 ;
  assign n34585 = n34303 | n34584 ;
  assign n34586 = ~n34510 & n34585 ;
  assign n34587 = x662 & ~n34586 ;
  assign n34588 = x662 | n34219 ;
  assign n34589 = ~n34587 & n34588 ;
  assign n34590 = ( x224 & ~n4721 ) | ( x224 & n34589 ) | ( ~n4721 & n34589 ) ;
  assign n34591 = n34582 | n34590 ;
  assign n34592 = x215 & n34591 ;
  assign n34593 = x614 & ~n33500 ;
  assign n34594 = n15646 & ~n34593 ;
  assign n34595 = x680 & ~n34594 ;
  assign n34596 = n34225 & ~n34595 ;
  assign n34597 = x662 & ~n34596 ;
  assign n34598 = ~n34224 & n34530 ;
  assign n34599 = n34229 & ~n34598 ;
  assign n34600 = ~n34597 & n34599 ;
  assign n34601 = ( x224 & ~n4721 ) | ( x224 & n34600 ) | ( ~n4721 & n34600 ) ;
  assign n34602 = ( x614 & ~n15620 ) | ( x614 & n15667 ) | ( ~n15620 & n15667 ) ;
  assign n34603 = ~n34522 & n34602 ;
  assign n34604 = x616 | n34603 ;
  assign n34605 = ~n34521 & n34604 ;
  assign n34606 = x680 & ~n34605 ;
  assign n34607 = n34238 & ~n34606 ;
  assign n34608 = x662 & ~n34607 ;
  assign n34609 = ~n34236 & n34530 ;
  assign n34610 = n34242 & ~n34609 ;
  assign n34611 = ~n34608 & n34610 ;
  assign n34612 = ( x224 & n4721 ) | ( x224 & n34611 ) | ( n4721 & n34611 ) ;
  assign n34613 = n34601 & n34612 ;
  assign n34614 = n34592 & ~n34613 ;
  assign n34615 = x299 & ~n34614 ;
  assign n34616 = ~n34571 & n34615 ;
  assign n34617 = ~x222 & n34562 ;
  assign n34618 = x223 | n34617 ;
  assign n34619 = ( n4346 & n4764 ) | ( n4346 & n34515 ) | ( n4764 & n34515 ) ;
  assign n34620 = ( n4346 & ~n4764 ) | ( n4346 & n34556 ) | ( ~n4764 & n34556 ) ;
  assign n34621 = n34619 & n34620 ;
  assign n34622 = n34618 | n34621 ;
  assign n34623 = ( ~x224 & n4764 ) | ( ~x224 & n34546 ) | ( n4764 & n34546 ) ;
  assign n34624 = ( x224 & n4764 ) | ( x224 & ~n34533 ) | ( n4764 & ~n34533 ) ;
  assign n34625 = ~n34623 & n34624 ;
  assign n34626 = n34622 | n34625 ;
  assign n34627 = ( x224 & ~n4764 ) | ( x224 & n34600 ) | ( ~n4764 & n34600 ) ;
  assign n34628 = ( x224 & n4764 ) | ( x224 & n34581 ) | ( n4764 & n34581 ) ;
  assign n34629 = ~n34627 & n34628 ;
  assign n34630 = x223 & ~n34629 ;
  assign n34631 = ( x224 & ~n4764 ) | ( x224 & n34589 ) | ( ~n4764 & n34589 ) ;
  assign n34632 = ( x224 & n4764 ) | ( x224 & n34611 ) | ( n4764 & n34611 ) ;
  assign n34633 = n34631 & ~n34632 ;
  assign n34634 = n34630 & ~n34633 ;
  assign n34635 = n34626 & ~n34634 ;
  assign n34636 = x299 | n34635 ;
  assign n34637 = x39 & n34636 ;
  assign n34638 = ~n34616 & n34637 ;
  assign n34639 = n15159 & n15881 ;
  assign n34640 = n34326 | n34639 ;
  assign n34641 = ~x224 & n34640 ;
  assign n34642 = ~n15159 & n15881 ;
  assign n34643 = ~n33567 & n34324 ;
  assign n34644 = ~n34642 & n34643 ;
  assign n34645 = n34641 | n34644 ;
  assign n34646 = ~x299 & n34645 ;
  assign n34647 = ~x614 & n14920 ;
  assign n34648 = n33549 | n34647 ;
  assign n34649 = x224 & n34648 ;
  assign n34650 = x224 | n15885 ;
  assign n34651 = n34317 | n34650 ;
  assign n34652 = ~n34649 & n34651 ;
  assign n34653 = ( x299 & ~n15159 ) | ( x299 & n34652 ) | ( ~n15159 & n34652 ) ;
  assign n34654 = ( x299 & n15159 ) | ( x299 & n34321 ) | ( n15159 & n34321 ) ;
  assign n34655 = n34653 & n34654 ;
  assign n34656 = n34646 | n34655 ;
  assign n34657 = ~x39 & n34656 ;
  assign n34658 = x38 | n34657 ;
  assign n34659 = n34638 | n34658 ;
  assign n34660 = x662 & n15477 ;
  assign n34661 = n15070 & n34660 ;
  assign n34662 = n34336 & ~n34661 ;
  assign n34663 = n2032 | n34662 ;
  assign n34664 = n34659 & ~n34663 ;
  assign n34665 = n34218 | n34664 ;
  assign n34666 = ( x625 & ~x1153 ) | ( x625 & n34665 ) | ( ~x1153 & n34665 ) ;
  assign n34667 = ~n34507 & n34666 ;
  assign n34668 = n34506 | n34667 ;
  assign n34669 = x608 & ~n34463 ;
  assign n34670 = ( x625 & x1153 ) | ( x625 & n34339 ) | ( x1153 & n34339 ) ;
  assign n34671 = ( ~x625 & x1153 ) | ( ~x625 & n34665 ) | ( x1153 & n34665 ) ;
  assign n34672 = n34670 & n34671 ;
  assign n34673 = n34669 & ~n34672 ;
  assign n34674 = n34668 & ~n34673 ;
  assign n34675 = x778 & ~n34674 ;
  assign n34676 = x778 | n34665 ;
  assign n34677 = ~n34675 & n34676 ;
  assign n34678 = ( x609 & ~x1155 ) | ( x609 & n34677 ) | ( ~x1155 & n34677 ) ;
  assign n34679 = ~n34505 & n34678 ;
  assign n34680 = n34504 | n34679 ;
  assign n34681 = x660 & ~n34349 ;
  assign n34682 = ( x609 & x1155 ) | ( x609 & n34466 ) | ( x1155 & n34466 ) ;
  assign n34683 = ( ~x609 & x1155 ) | ( ~x609 & n34677 ) | ( x1155 & n34677 ) ;
  assign n34684 = n34682 & n34683 ;
  assign n34685 = n34681 & ~n34684 ;
  assign n34686 = n34680 & ~n34685 ;
  assign n34687 = x785 & ~n34686 ;
  assign n34688 = x785 | n34677 ;
  assign n34689 = ~n34687 & n34688 ;
  assign n34690 = ( x618 & ~x1154 ) | ( x618 & n34689 ) | ( ~x1154 & n34689 ) ;
  assign n34691 = ~n34503 & n34690 ;
  assign n34692 = n34502 | n34691 ;
  assign n34693 = x627 & ~n34359 ;
  assign n34694 = ( x618 & x1154 ) | ( x618 & n34469 ) | ( x1154 & n34469 ) ;
  assign n34695 = ( ~x618 & x1154 ) | ( ~x618 & n34689 ) | ( x1154 & n34689 ) ;
  assign n34696 = n34694 & n34695 ;
  assign n34697 = n34693 & ~n34696 ;
  assign n34698 = n34692 & ~n34697 ;
  assign n34699 = x781 & ~n34698 ;
  assign n34700 = x781 | n34689 ;
  assign n34701 = ~n34699 & n34700 ;
  assign n34702 = ( ~x619 & x1159 ) | ( ~x619 & n34701 ) | ( x1159 & n34701 ) ;
  assign n34703 = n34501 & n34702 ;
  assign n34704 = n34500 & ~n34703 ;
  assign n34705 = x648 | n34366 ;
  assign n34706 = ( x619 & x1159 ) | ( x619 & ~n34472 ) | ( x1159 & ~n34472 ) ;
  assign n34707 = ( x619 & ~x1159 ) | ( x619 & n34701 ) | ( ~x1159 & n34701 ) ;
  assign n34708 = ~n34706 & n34707 ;
  assign n34709 = n34705 | n34708 ;
  assign n34710 = x789 & n34709 ;
  assign n34711 = ~n34704 & n34710 ;
  assign n34712 = ~x789 & n34701 ;
  assign n34713 = n16177 | n34712 ;
  assign n34714 = n34711 | n34713 ;
  assign n34715 = n15414 & ~n34215 ;
  assign n34716 = n34473 & ~n34715 ;
  assign n34717 = n16115 & ~n34716 ;
  assign n34718 = ( x626 & n15418 ) | ( x626 & ~n34215 ) | ( n15418 & ~n34215 ) ;
  assign n34719 = ( x626 & ~n15418 ) | ( x626 & n34372 ) | ( ~n15418 & n34372 ) ;
  assign n34720 = n34718 & ~n34719 ;
  assign n34721 = n34717 | n34720 ;
  assign n34722 = ( x626 & ~n15419 ) | ( x626 & n34215 ) | ( ~n15419 & n34215 ) ;
  assign n34723 = ( x626 & n15419 ) | ( x626 & ~n34372 ) | ( n15419 & ~n34372 ) ;
  assign n34724 = ~n34722 & n34723 ;
  assign n34725 = n34721 | n34724 ;
  assign n34726 = x788 & n34725 ;
  assign n34727 = n18434 | n34726 ;
  assign n34728 = n34714 & ~n34727 ;
  assign n34729 = n34499 | n34728 ;
  assign n34730 = ~n18431 & n34729 ;
  assign n34731 = n18610 & n34377 ;
  assign n34732 = ( x630 & n34485 ) | ( x630 & n34731 ) | ( n34485 & n34731 ) ;
  assign n34733 = ( ~x630 & n34482 ) | ( ~x630 & n34731 ) | ( n34482 & n34731 ) ;
  assign n34734 = n34732 | n34733 ;
  assign n34735 = x787 & n34734 ;
  assign n34736 = n34730 | n34735 ;
  assign n34737 = ( ~x644 & x715 ) | ( ~x644 & n34736 ) | ( x715 & n34736 ) ;
  assign n34738 = n34489 & n34737 ;
  assign n34739 = n34383 & ~n34738 ;
  assign n34740 = ( x644 & x715 ) | ( x644 & n34379 ) | ( x715 & n34379 ) ;
  assign n34741 = ( ~x644 & x715 ) | ( ~x644 & n34215 ) | ( x715 & n34215 ) ;
  assign n34742 = n34740 & n34741 ;
  assign n34743 = x1160 | n34742 ;
  assign n34744 = ( x644 & x715 ) | ( x644 & ~n34488 ) | ( x715 & ~n34488 ) ;
  assign n34745 = ( x644 & ~x715 ) | ( x644 & n34736 ) | ( ~x715 & n34736 ) ;
  assign n34746 = ~n34744 & n34745 ;
  assign n34747 = n34743 | n34746 ;
  assign n34748 = ~n34739 & n34747 ;
  assign n34749 = ( x790 & n6785 ) | ( x790 & n34748 ) | ( n6785 & n34748 ) ;
  assign n34750 = ( ~x790 & n6785 ) | ( ~x790 & n34736 ) | ( n6785 & n34736 ) ;
  assign n34751 = n34749 | n34750 ;
  assign n34752 = ~n34214 & n34751 ;
  assign n34753 = n1880 & ~n1976 ;
  assign n34754 = ~n2192 & n34753 ;
  assign n34755 = ~x62 & n34754 ;
  assign n34756 = n2057 & ~n34755 ;
  assign n34757 = n13509 | n34756 ;
  assign n34758 = ( x62 & n2057 ) | ( x62 & n34754 ) | ( n2057 & n34754 ) ;
  assign n34759 = n4694 | n4784 ;
  assign n34760 = ~x137 & n34759 ;
  assign n34761 = n4811 & ~n34760 ;
  assign n34762 = ~n1496 & n1746 ;
  assign n34763 = x137 & ~n34762 ;
  assign n34764 = n1711 & ~n34763 ;
  assign n34765 = x332 | n34764 ;
  assign n34766 = ~n1212 & n9552 ;
  assign n34767 = n1684 | n34766 ;
  assign n34768 = x137 | n1706 ;
  assign n34769 = n34767 & ~n34768 ;
  assign n34770 = x332 & ~n34769 ;
  assign n34771 = n1539 | n9552 ;
  assign n34772 = n1740 | n34771 ;
  assign n34773 = ~n1302 & n34772 ;
  assign n34774 = n1300 | n34773 ;
  assign n34775 = ~n1706 & n34774 ;
  assign n34776 = ( x95 & n1674 ) | ( x95 & n34775 ) | ( n1674 & n34775 ) ;
  assign n34777 = n34770 & ~n34776 ;
  assign n34778 = n34765 & ~n34777 ;
  assign n34779 = x210 & ~n34778 ;
  assign n34780 = x299 & ~n34779 ;
  assign n34781 = ~n1610 & n34774 ;
  assign n34782 = x95 | n34781 ;
  assign n34783 = ~n1496 & n34782 ;
  assign n34784 = x137 & ~n34783 ;
  assign n34785 = ~n1635 & n34767 ;
  assign n34786 = x137 | n34785 ;
  assign n34787 = ~n34784 & n34786 ;
  assign n34788 = x332 & ~n34787 ;
  assign n34789 = ~n1496 & n1753 ;
  assign n34790 = x137 & ~n34789 ;
  assign n34791 = n1686 & ~n34790 ;
  assign n34792 = x332 | n34791 ;
  assign n34793 = ~n34788 & n34792 ;
  assign n34794 = ( x210 & n1615 ) | ( x210 & n34793 ) | ( n1615 & n34793 ) ;
  assign n34795 = x1093 & ~n34785 ;
  assign n34796 = ~n1635 & n1693 ;
  assign n34797 = n1212 | n5910 ;
  assign n34798 = n1597 & ~n34797 ;
  assign n34799 = x32 | n34798 ;
  assign n34800 = n34796 & n34799 ;
  assign n34801 = x1093 | n34800 ;
  assign n34802 = ~n1693 & n34785 ;
  assign n34803 = n9551 & ~n34797 ;
  assign n34804 = n34796 & n34803 ;
  assign n34805 = n34802 | n34804 ;
  assign n34806 = n34801 | n34805 ;
  assign n34807 = ~n34795 & n34806 ;
  assign n34808 = n9680 | n34807 ;
  assign n34809 = n1685 & ~n1693 ;
  assign n34810 = n34801 | n34809 ;
  assign n34811 = n1632 & ~n34797 ;
  assign n34812 = x32 | n34811 ;
  assign n34813 = n34796 & n34812 ;
  assign n34814 = x1093 & ~n34809 ;
  assign n34815 = ~n34813 & n34814 ;
  assign n34816 = n34810 & ~n34815 ;
  assign n34817 = n9648 & ~n34816 ;
  assign n34818 = ~n34805 & n34817 ;
  assign n34819 = n34808 & ~n34818 ;
  assign n34820 = ~n34784 & n34819 ;
  assign n34821 = x332 & ~n34820 ;
  assign n34822 = x1093 & ~n1685 ;
  assign n34823 = n34810 & ~n34822 ;
  assign n34824 = n9680 | n34823 ;
  assign n34825 = ~n34817 & n34824 ;
  assign n34826 = ~n34790 & n34825 ;
  assign n34827 = x332 | n34826 ;
  assign n34828 = ~n34821 & n34827 ;
  assign n34829 = ( x210 & ~n1615 ) | ( x210 & n34828 ) | ( ~n1615 & n34828 ) ;
  assign n34830 = n34794 | n34829 ;
  assign n34831 = n34780 & n34830 ;
  assign n34832 = x198 & ~n34778 ;
  assign n34833 = x299 | n34832 ;
  assign n34834 = ( x198 & n4781 ) | ( x198 & n34793 ) | ( n4781 & n34793 ) ;
  assign n34835 = ( x198 & ~n4781 ) | ( x198 & n34828 ) | ( ~n4781 & n34828 ) ;
  assign n34836 = n34834 | n34835 ;
  assign n34837 = ~n34833 & n34836 ;
  assign n34838 = n34831 | n34837 ;
  assign n34839 = ~x39 & n34838 ;
  assign n34840 = ( x38 & n1880 ) | ( x38 & n1925 ) | ( n1880 & n1925 ) ;
  assign n34841 = n34839 | n34840 ;
  assign n34842 = x38 & ~x137 ;
  assign n34843 = n4662 | n34842 ;
  assign n34844 = n34841 & ~n34843 ;
  assign n34845 = n34761 | n34844 ;
  assign n34846 = ~x87 & n34845 ;
  assign n34847 = ( x75 & n1998 ) | ( x75 & n34753 ) | ( n1998 & n34753 ) ;
  assign n34848 = n34846 | n34847 ;
  assign n34849 = n5762 | n34760 ;
  assign n34850 = x75 & n34849 ;
  assign n34851 = x92 | n34850 ;
  assign n34852 = n34848 & ~n34851 ;
  assign n34853 = ~n1998 & n34753 ;
  assign n34854 = ( x54 & n4817 ) | ( x54 & n34853 ) | ( n4817 & n34853 ) ;
  assign n34855 = n34852 | n34854 ;
  assign n34856 = ~n2042 & n34753 ;
  assign n34857 = x54 & ~n34856 ;
  assign n34858 = x74 | n34857 ;
  assign n34859 = n34855 & ~n34858 ;
  assign n34860 = ~n4654 & n34753 ;
  assign n34861 = ( x55 & n5073 ) | ( x55 & n34860 ) | ( n5073 & n34860 ) ;
  assign n34862 = n34859 | n34861 ;
  assign n34863 = ~n5760 & n34862 ;
  assign n34864 = x56 & ~n2044 ;
  assign n34865 = n34753 & n34864 ;
  assign n34866 = n34863 | n34865 ;
  assign n34867 = ( ~x62 & n2057 ) | ( ~x62 & n34866 ) | ( n2057 & n34866 ) ;
  assign n34868 = n34758 | n34867 ;
  assign n34869 = ~n34757 & n34868 ;
  assign n34870 = x228 & x231 ;
  assign n34871 = n5845 & ~n34870 ;
  assign n34872 = x74 & ~n34871 ;
  assign n34873 = x55 | n34872 ;
  assign n34874 = ( x54 & x74 ) | ( x54 & ~n34870 ) | ( x74 & ~n34870 ) ;
  assign n34875 = n1274 | n1460 ;
  assign n34876 = ~n1294 & n34875 ;
  assign n34877 = ( x51 & ~n1465 ) | ( x51 & n34876 ) | ( ~n1465 & n34876 ) ;
  assign n34878 = n1539 | n34877 ;
  assign n34879 = ~n1302 & n34878 ;
  assign n34880 = n1300 | n34879 ;
  assign n34881 = ~n4701 & n34880 ;
  assign n34882 = x95 | n34881 ;
  assign n34883 = ~n1497 & n34882 ;
  assign n34884 = x39 | n34883 ;
  assign n34885 = x38 | n2120 ;
  assign n34886 = n34884 & ~n34885 ;
  assign n34887 = ~x228 & n34886 ;
  assign n34888 = n34870 | n34887 ;
  assign n34889 = ( x87 & ~x100 ) | ( x87 & n34888 ) | ( ~x100 & n34888 ) ;
  assign n34890 = n11995 & ~n34870 ;
  assign n34891 = ( x87 & x100 ) | ( x87 & ~n34890 ) | ( x100 & ~n34890 ) ;
  assign n34892 = n34889 | n34891 ;
  assign n34893 = n5811 & ~n34870 ;
  assign n34894 = ( x75 & n1998 ) | ( x75 & n34893 ) | ( n1998 & n34893 ) ;
  assign n34895 = n34892 & ~n34894 ;
  assign n34896 = n12000 & ~n34870 ;
  assign n34897 = x75 & ~n34896 ;
  assign n34898 = x92 | n34897 ;
  assign n34899 = n34895 | n34898 ;
  assign n34900 = x92 & ~n34870 ;
  assign n34901 = n5836 & n34900 ;
  assign n34902 = n34899 & ~n34901 ;
  assign n34903 = ( x54 & ~x74 ) | ( x54 & n34902 ) | ( ~x74 & n34902 ) ;
  assign n34904 = ~n34874 & n34903 ;
  assign n34905 = n34873 | n34904 ;
  assign n34906 = x55 & ~n34870 ;
  assign n34907 = x56 | n34906 ;
  assign n34908 = n34905 & ~n34907 ;
  assign n34909 = n5851 & ~n34870 ;
  assign n34910 = x56 & ~n34909 ;
  assign n34911 = x62 | n34910 ;
  assign n34912 = n34908 | n34911 ;
  assign n34913 = x62 & ~n34870 ;
  assign n34914 = n5812 & n34913 ;
  assign n34915 = n34912 & ~n34914 ;
  assign n34916 = n2057 | n34915 ;
  assign n34917 = n2057 & ~n34870 ;
  assign n34918 = n34916 & ~n34917 ;
  assign n34919 = n1259 | n4884 ;
  assign n34920 = ~n1312 & n9190 ;
  assign n34921 = n9188 & n34920 ;
  assign n34922 = x91 | n4678 ;
  assign n34923 = ~n1692 & n9180 ;
  assign n34924 = n34922 | n34923 ;
  assign n34925 = n34921 | n34924 ;
  assign n34926 = ~n34919 & n34925 ;
  assign n34927 = x72 | n34926 ;
  assign n34928 = ~n4905 & n34927 ;
  assign n34929 = n4742 & ~n34928 ;
  assign n34930 = n11122 & n11156 ;
  assign n34931 = ~n4905 & n34930 ;
  assign n34932 = n4987 | n34931 ;
  assign n34933 = x1093 & n34932 ;
  assign n34934 = n9180 & ~n34919 ;
  assign n34935 = ~n5950 & n34934 ;
  assign n34936 = ~n34919 & n34922 ;
  assign n34937 = x72 | n34936 ;
  assign n34938 = n7134 | n34937 ;
  assign n34939 = n34935 | n34938 ;
  assign n34940 = ~n4905 & n34939 ;
  assign n34941 = n34933 | n34940 ;
  assign n34942 = n34934 | n34937 ;
  assign n34943 = ~n4905 & n34942 ;
  assign n34944 = n8243 & ~n34943 ;
  assign n34945 = n34941 & ~n34944 ;
  assign n34946 = ~n34929 & n34945 ;
  assign n34947 = x39 | n34946 ;
  assign n34948 = ~n9607 & n34947 ;
  assign n34949 = n9555 | n9560 ;
  assign n34950 = x39 & n34949 ;
  assign n34951 = n4996 & n34950 ;
  assign n34952 = n1690 | n7135 ;
  assign n34953 = x32 | n4658 ;
  assign n34954 = n34952 & ~n34953 ;
  assign n34955 = ~n1599 & n34954 ;
  assign n34956 = n9622 & n34955 ;
  assign n34957 = n34951 | n34956 ;
  assign n34958 = ~n8366 & n34957 ;
  assign n34959 = n8693 | n34958 ;
  assign n34960 = n4661 | n8359 ;
  assign n34961 = ( n14786 & n14794 ) | ( n14786 & n14796 ) | ( n14794 & n14796 ) ;
  assign n34962 = x824 & ~n34961 ;
  assign n34963 = x829 & x1091 ;
  assign n34964 = ( x32 & ~n14736 ) | ( x32 & n14800 ) | ( ~n14736 & n14800 ) ;
  assign n34965 = n14796 & n34964 ;
  assign n34966 = n34963 & n34965 ;
  assign n34967 = x824 | n34966 ;
  assign n34968 = n34963 & ~n34967 ;
  assign n34969 = n34962 | n34968 ;
  assign n34970 = n1692 & ~n4992 ;
  assign n34971 = n34969 & n34970 ;
  assign n34972 = n4694 | n4992 ;
  assign n34973 = ~n14736 & n14744 ;
  assign n34974 = ~n4992 & n34967 ;
  assign n34975 = ~n34962 & n34974 ;
  assign n34976 = n34973 | n34975 ;
  assign n34977 = n34972 & n34976 ;
  assign n34978 = ~n34971 & n34977 ;
  assign n34979 = ~n5950 & n34973 ;
  assign n34980 = n14775 | n34979 ;
  assign n34981 = ~n34972 & n34980 ;
  assign n34982 = x1093 & ~n34981 ;
  assign n34983 = ~n34978 & n34982 ;
  assign n34984 = ~n4799 & n34973 ;
  assign n34985 = n4695 | n14711 ;
  assign n34986 = n14729 & ~n34985 ;
  assign n34987 = x40 | n34986 ;
  assign n34988 = ~n8462 & n34987 ;
  assign n34989 = x252 & ~n34988 ;
  assign n34990 = n4799 & n14743 ;
  assign n34991 = ~n34989 & n34990 ;
  assign n34992 = x1093 | n34991 ;
  assign n34993 = n34984 | n34992 ;
  assign n34994 = ~x39 & n34993 ;
  assign n34995 = ~n34983 & n34994 ;
  assign n34996 = n4798 & n5949 ;
  assign n34997 = ( x1091 & n14584 ) | ( x1091 & ~n34996 ) | ( n14584 & ~n34996 ) ;
  assign n34998 = ( x1091 & n14478 ) | ( x1091 & n34996 ) | ( n14478 & n34996 ) ;
  assign n34999 = n34997 & n34998 ;
  assign n35000 = ( x1091 & n4983 ) | ( x1091 & ~n14584 ) | ( n4983 & ~n14584 ) ;
  assign n35001 = ( ~x1091 & n4983 ) | ( ~x1091 & n14478 ) | ( n4983 & n14478 ) ;
  assign n35002 = ~n35000 & n35001 ;
  assign n35003 = n34999 | n35002 ;
  assign n35004 = ~x120 & n35003 ;
  assign n35005 = n14480 | n35004 ;
  assign n35006 = n4751 | n35005 ;
  assign n35007 = ~n32569 & n35006 ;
  assign n35008 = ( ~n1823 & n4764 ) | ( ~n1823 & n35007 ) | ( n4764 & n35007 ) ;
  assign n35009 = n4714 | n14481 ;
  assign n35010 = n4714 & ~n35005 ;
  assign n35011 = n35009 & ~n35010 ;
  assign n35012 = ( n1823 & n4764 ) | ( n1823 & ~n35011 ) | ( n4764 & ~n35011 ) ;
  assign n35013 = ~n35008 & n35012 ;
  assign n35014 = ( ~x223 & n14481 ) | ( ~x223 & n15629 ) | ( n14481 & n15629 ) ;
  assign n35015 = ~n35013 & n35014 ;
  assign n35016 = x120 & n4745 ;
  assign n35017 = n14481 | n35016 ;
  assign n35018 = ~n32569 & n35017 ;
  assign n35019 = ( x223 & ~n4764 ) | ( x223 & n35018 ) | ( ~n4764 & n35018 ) ;
  assign n35020 = n35009 & n35017 ;
  assign n35021 = ( x223 & n4764 ) | ( x223 & n35020 ) | ( n4764 & n35020 ) ;
  assign n35022 = n35019 & n35021 ;
  assign n35023 = x299 | n35022 ;
  assign n35024 = n35015 | n35023 ;
  assign n35025 = n2203 | n14481 ;
  assign n35026 = ~x215 & n35025 ;
  assign n35027 = ( ~n2203 & n4721 ) | ( ~n2203 & n35007 ) | ( n4721 & n35007 ) ;
  assign n35028 = ( n2203 & n4721 ) | ( n2203 & ~n35011 ) | ( n4721 & ~n35011 ) ;
  assign n35029 = ~n35027 & n35028 ;
  assign n35030 = n35026 & ~n35029 ;
  assign n35031 = ( x215 & ~n4721 ) | ( x215 & n35018 ) | ( ~n4721 & n35018 ) ;
  assign n35032 = ( x215 & n4721 ) | ( x215 & n35020 ) | ( n4721 & n35020 ) ;
  assign n35033 = n35031 & n35032 ;
  assign n35034 = x299 & ~n35033 ;
  assign n35035 = ~n35030 & n35034 ;
  assign n35036 = n35024 & ~n35035 ;
  assign n35037 = x39 & ~n35036 ;
  assign n35038 = x38 | n35037 ;
  assign n35039 = n34995 | n35038 ;
  assign n35040 = ~n34960 & n35039 ;
  assign n35041 = x81 | n1427 ;
  assign n35042 = ~n4869 & n35041 ;
  assign n35043 = n1243 | n35042 ;
  assign n35044 = ~n1439 & n35043 ;
  assign n35045 = n1350 | n35044 ;
  assign n35046 = ~n1443 & n35045 ;
  assign n35047 = n1582 | n35046 ;
  assign n35048 = ~n1584 & n35047 ;
  assign n35049 = x86 | n35048 ;
  assign n35050 = ~n1347 & n35049 ;
  assign n35051 = n1345 | n35050 ;
  assign n35052 = ~n1337 & n35051 ;
  assign n35053 = x108 | n35052 ;
  assign n35054 = ~n1334 & n35053 ;
  assign n35055 = n1731 | n35054 ;
  assign n35056 = ~n1454 & n35055 ;
  assign n35057 = ( ~n1324 & n1325 ) | ( ~n1324 & n35056 ) | ( n1325 & n35056 ) ;
  assign n35058 = n1315 | n35057 ;
  assign n35059 = ~n1310 & n35058 ;
  assign n35060 = n1278 | n35059 ;
  assign n35061 = ~n13522 & n35060 ;
  assign n35062 = x70 | n35061 ;
  assign n35063 = ~n1280 & n35062 ;
  assign n35064 = x51 | n35063 ;
  assign n35065 = ~n1465 & n35064 ;
  assign n35066 = n1539 | n35065 ;
  assign n35067 = ~n1302 & n35066 ;
  assign n35068 = ~x1082 & n1299 ;
  assign n35069 = x32 | n35068 ;
  assign n35070 = n35067 | n35069 ;
  assign n35071 = ~n2129 & n35070 ;
  assign n35072 = x95 | n35071 ;
  assign n35073 = ~n1496 & n35072 ;
  assign n35074 = x39 | n35073 ;
  assign n35075 = n5771 | n5773 ;
  assign n35076 = n1692 & n4744 ;
  assign n35077 = n4978 & n35076 ;
  assign n35078 = n35075 & n35077 ;
  assign n35079 = n4729 & n9505 ;
  assign n35080 = ~n35078 & n35079 ;
  assign n35081 = n2120 | n35080 ;
  assign n35082 = n35074 & ~n35081 ;
  assign n35083 = x38 | n35082 ;
  assign n35084 = ~n4662 & n35083 ;
  assign n35085 = n4812 | n35084 ;
  assign n35086 = ~n4815 & n35085 ;
  assign n35087 = n2004 | n35086 ;
  assign n35088 = ~n5767 & n35087 ;
  assign n35089 = x54 | n35088 ;
  assign n35090 = ~n5801 & n35089 ;
  assign n35091 = n5073 | n35090 ;
  assign n35092 = ~n13596 & n35091 ;
  assign n35093 = x56 | n35092 ;
  assign n35094 = ~n4653 & n35093 ;
  assign n35095 = x62 | n35094 ;
  assign n35096 = ~n4826 & n35095 ;
  assign n35097 = n2057 | n35096 ;
  assign n35098 = ~n4649 & n35097 ;
  assign n35099 = x230 | x233 ;
  assign n35100 = x212 | x214 ;
  assign n35101 = ~x211 & n35100 ;
  assign n35102 = x219 & ~n35101 ;
  assign n35103 = n6785 & ~n35102 ;
  assign n35104 = x1142 & n8654 ;
  assign n35105 = x211 & x1143 ;
  assign n35106 = ~x211 & x1144 ;
  assign n35107 = n35105 | n35106 ;
  assign n35108 = ~x212 & x214 ;
  assign n35109 = x212 & ~x214 ;
  assign n35110 = n35108 | n35109 ;
  assign n35111 = n35107 & n35110 ;
  assign n35112 = ~x211 & x1143 ;
  assign n35113 = n8894 & n35112 ;
  assign n35114 = n35111 | n35113 ;
  assign n35115 = ~x219 & n35114 ;
  assign n35116 = n35104 | n35115 ;
  assign n35117 = n35103 & n35116 ;
  assign n35118 = x299 & n35107 ;
  assign n35119 = x199 & x1142 ;
  assign n35120 = x200 | n35119 ;
  assign n35121 = ~x199 & x1143 ;
  assign n35122 = n35120 | n35121 ;
  assign n35123 = x207 & ~x299 ;
  assign n35124 = ~x199 & x1142 ;
  assign n35125 = x200 & ~n35124 ;
  assign n35126 = n35123 & ~n35125 ;
  assign n35127 = n35122 & n35126 ;
  assign n35128 = ~x199 & x1144 ;
  assign n35129 = n35120 | n35128 ;
  assign n35130 = x200 & ~n35121 ;
  assign n35131 = n35129 & ~n35130 ;
  assign n35132 = x207 | x299 ;
  assign n35133 = n35131 | n35132 ;
  assign n35134 = ( ~x207 & n35127 ) | ( ~x207 & n35133 ) | ( n35127 & n35133 ) ;
  assign n35135 = x208 & n35134 ;
  assign n35136 = x207 & ~x208 ;
  assign n35137 = n35131 & n35136 ;
  assign n35138 = n35135 | n35137 ;
  assign n35139 = ~x299 & n35138 ;
  assign n35140 = n35118 | n35139 ;
  assign n35141 = x214 | n35139 ;
  assign n35142 = ~x212 & n35141 ;
  assign n35143 = n35140 & n35142 ;
  assign n35144 = n35118 | n35141 ;
  assign n35145 = x211 & x1142 ;
  assign n35146 = n35112 | n35145 ;
  assign n35147 = x299 & n35146 ;
  assign n35148 = n35139 | n35147 ;
  assign n35149 = ( x212 & n35109 ) | ( x212 & n35148 ) | ( n35109 & n35148 ) ;
  assign n35150 = n35144 & n35149 ;
  assign n35151 = x219 | n35150 ;
  assign n35152 = n35143 | n35151 ;
  assign n35153 = x299 | n35138 ;
  assign n35154 = x299 & ~x1142 ;
  assign n35155 = n35101 & ~n35154 ;
  assign n35156 = n35153 & n35155 ;
  assign n35157 = ~n35101 & n35139 ;
  assign n35158 = x219 & ~n35157 ;
  assign n35159 = ~n35156 & n35158 ;
  assign n35160 = n6785 | n35159 ;
  assign n35161 = n35152 & ~n35160 ;
  assign n35162 = n35117 | n35161 ;
  assign n35163 = x213 & ~n35162 ;
  assign n35164 = ~x211 & x1156 ;
  assign n35165 = x211 & x1155 ;
  assign n35166 = n35164 | n35165 ;
  assign n35167 = ~x214 & n35166 ;
  assign n35168 = ~x211 & x1155 ;
  assign n35169 = x211 & x1154 ;
  assign n35170 = n35168 | n35169 ;
  assign n35171 = x214 & n35170 ;
  assign n35172 = n35167 | n35171 ;
  assign n35173 = x212 & n35172 ;
  assign n35174 = ~x211 & x1157 ;
  assign n35175 = x211 & x1156 ;
  assign n35176 = n35174 | n35175 ;
  assign n35177 = x214 & n35176 ;
  assign n35178 = ~x212 & n35177 ;
  assign n35179 = n35173 | n35178 ;
  assign n35180 = ( x219 & n6785 ) | ( x219 & n35179 ) | ( n6785 & n35179 ) ;
  assign n35181 = ~x211 & x1154 ;
  assign n35182 = x214 | n35181 ;
  assign n35183 = ~x211 & x1153 ;
  assign n35184 = n8894 & ~n35183 ;
  assign n35185 = n35182 & ~n35184 ;
  assign n35186 = ( x212 & n35100 ) | ( x212 & n35168 ) | ( n35100 & n35168 ) ;
  assign n35187 = n35185 & n35186 ;
  assign n35188 = ( ~x219 & n6785 ) | ( ~x219 & n35187 ) | ( n6785 & n35187 ) ;
  assign n35189 = n35180 & n35188 ;
  assign n35190 = x213 | n35189 ;
  assign n35191 = ~x219 & x299 ;
  assign n35192 = n35179 & n35191 ;
  assign n35193 = x299 & x1155 ;
  assign n35194 = n35108 & n35193 ;
  assign n35195 = x299 & x1153 ;
  assign n35196 = ( x212 & ~x214 ) | ( x212 & n35195 ) | ( ~x214 & n35195 ) ;
  assign n35197 = x299 & x1154 ;
  assign n35198 = ( x212 & x214 ) | ( x212 & n35197 ) | ( x214 & n35197 ) ;
  assign n35199 = n35196 & n35198 ;
  assign n35200 = n35194 | n35199 ;
  assign n35201 = ~x211 & x219 ;
  assign n35202 = n35200 & n35201 ;
  assign n35203 = n35192 | n35202 ;
  assign n35204 = n35139 | n35203 ;
  assign n35205 = ~n6785 & n35204 ;
  assign n35206 = n35190 | n35205 ;
  assign n35207 = x209 & n35206 ;
  assign n35208 = ~n35163 & n35207 ;
  assign n35209 = ~x200 & x1155 ;
  assign n35210 = x199 & n35209 ;
  assign n35211 = ~x299 & n35210 ;
  assign n35212 = x1156 | n35211 ;
  assign n35213 = x200 | x1155 ;
  assign n35214 = x199 & x200 ;
  assign n35215 = n8980 & ~n35214 ;
  assign n35216 = ~x299 & n35215 ;
  assign n35217 = n35213 & n35216 ;
  assign n35218 = n35212 & n35217 ;
  assign n35219 = x207 & n35218 ;
  assign n35220 = x208 | n35219 ;
  assign n35221 = x299 | n35214 ;
  assign n35222 = x1153 & n35221 ;
  assign n35223 = x1154 & ~n35222 ;
  assign n35224 = ~n9520 & n35209 ;
  assign n35225 = ~x1153 & n9520 ;
  assign n35226 = x1154 & n35215 ;
  assign n35227 = ~n35225 & n35226 ;
  assign n35228 = n35224 | n35227 ;
  assign n35229 = n35223 & n35228 ;
  assign n35230 = x200 | x299 ;
  assign n35231 = x199 & ~x1153 ;
  assign n35232 = n35230 | n35231 ;
  assign n35233 = x199 | x1155 ;
  assign n35234 = ~x1154 & n35233 ;
  assign n35235 = ~n35232 & n35234 ;
  assign n35236 = n35229 | n35235 ;
  assign n35237 = x207 & ~n35236 ;
  assign n35238 = x200 & ~x299 ;
  assign n35239 = ~x199 & x1155 ;
  assign n35240 = n35238 & n35239 ;
  assign n35241 = x1154 | n35240 ;
  assign n35242 = x200 & ~n35239 ;
  assign n35243 = n8981 & ~n35242 ;
  assign n35244 = n35241 & n35243 ;
  assign n35245 = x200 & ~x1155 ;
  assign n35246 = n9520 | n35245 ;
  assign n35247 = x1156 & ~n35246 ;
  assign n35248 = n35244 | n35247 ;
  assign n35249 = x207 | n35248 ;
  assign n35250 = ~n35237 & n35249 ;
  assign n35251 = x208 & ~n35250 ;
  assign n35252 = n35220 & ~n35251 ;
  assign n35253 = x1157 | n35252 ;
  assign n35254 = x199 & ~x1155 ;
  assign n35255 = x1156 & ~n35254 ;
  assign n35256 = ~n35221 & n35255 ;
  assign n35257 = x1156 | n35254 ;
  assign n35258 = n35230 | n35257 ;
  assign n35259 = ~n35256 & n35258 ;
  assign n35260 = x207 & ~n35259 ;
  assign n35261 = x208 | n35260 ;
  assign n35262 = ~n35251 & n35261 ;
  assign n35263 = x1157 & ~n35262 ;
  assign n35264 = n35253 & ~n35263 ;
  assign n35265 = x211 & ~n35264 ;
  assign n35266 = x214 | n35264 ;
  assign n35267 = ~x212 & n35266 ;
  assign n35268 = ~x211 & x214 ;
  assign n35269 = n9515 & ~n35213 ;
  assign n35270 = x1153 & n35269 ;
  assign n35271 = x1153 & ~n35238 ;
  assign n35272 = x1153 | n8981 ;
  assign n35273 = ~n35271 & n35272 ;
  assign n35274 = x1155 & ~n35273 ;
  assign n35275 = n35270 | n35274 ;
  assign n35276 = ~x1154 & n35275 ;
  assign n35277 = x1155 & ~n9515 ;
  assign n35278 = n35216 & ~n35231 ;
  assign n35279 = n35277 | n35278 ;
  assign n35280 = x1154 & n35279 ;
  assign n35281 = n35276 | n35280 ;
  assign n35282 = x207 & ~n35281 ;
  assign n35283 = x207 | n35193 ;
  assign n35284 = n35248 | n35283 ;
  assign n35285 = x208 & n35284 ;
  assign n35286 = ~n35282 & n35285 ;
  assign n35287 = x1155 & ~n35238 ;
  assign n35288 = n9520 & ~n35287 ;
  assign n35289 = x1156 & ~n35288 ;
  assign n35290 = x199 & ~x200 ;
  assign n35291 = x299 | n35290 ;
  assign n35292 = ~x1155 & n35291 ;
  assign n35293 = x1156 | n35238 ;
  assign n35294 = n35292 | n35293 ;
  assign n35295 = ~n35289 & n35294 ;
  assign n35296 = x207 & n35295 ;
  assign n35297 = ~x208 & n35283 ;
  assign n35298 = x1157 & n35297 ;
  assign n35299 = ~n35296 & n35298 ;
  assign n35300 = x299 | n35212 ;
  assign n35301 = x299 | n35215 ;
  assign n35302 = ~x1155 & n9520 ;
  assign n35303 = n35301 & ~n35302 ;
  assign n35304 = n35300 & n35303 ;
  assign n35305 = n35297 & n35304 ;
  assign n35306 = n35299 | n35305 ;
  assign n35307 = n35286 | n35306 ;
  assign n35308 = n35268 & ~n35307 ;
  assign n35309 = n35267 & ~n35308 ;
  assign n35310 = x1155 | n8981 ;
  assign n35311 = ~n35287 & n35310 ;
  assign n35312 = x1156 | n35311 ;
  assign n35313 = n9515 & ~n35209 ;
  assign n35314 = x1156 & ~n35313 ;
  assign n35315 = n35312 & ~n35314 ;
  assign n35316 = x207 & n35315 ;
  assign n35317 = ~x208 & n35132 ;
  assign n35318 = ~n35316 & n35317 ;
  assign n35319 = x1157 & ~n35318 ;
  assign n35320 = x299 | n9578 ;
  assign n35321 = x1156 & ~n35210 ;
  assign n35322 = ~n35320 & n35321 ;
  assign n35323 = n35212 & ~n35322 ;
  assign n35324 = n35123 & n35323 ;
  assign n35325 = ( ~x208 & x299 ) | ( ~x208 & n35324 ) | ( x299 & n35324 ) ;
  assign n35326 = x1157 | n35325 ;
  assign n35327 = x299 & ~x1153 ;
  assign n35328 = n35326 & ~n35327 ;
  assign n35329 = ~n35319 & n35328 ;
  assign n35330 = x1153 & n35291 ;
  assign n35331 = n35228 | n35330 ;
  assign n35332 = x207 & n35331 ;
  assign n35333 = ~n35277 & n35310 ;
  assign n35334 = x1156 & ~n35333 ;
  assign n35335 = x1155 & n35301 ;
  assign n35336 = n35292 | n35335 ;
  assign n35337 = x1154 & n35336 ;
  assign n35338 = n35334 | n35337 ;
  assign n35339 = x299 & ~x1155 ;
  assign n35340 = x1155 & n35320 ;
  assign n35341 = n35339 | n35340 ;
  assign n35342 = n35338 | n35341 ;
  assign n35343 = x207 | n35327 ;
  assign n35344 = n35342 & ~n35343 ;
  assign n35345 = n35332 | n35344 ;
  assign n35346 = x208 & n35345 ;
  assign n35347 = n35268 & ~n35346 ;
  assign n35348 = ~n35329 & n35347 ;
  assign n35349 = n35248 | n35337 ;
  assign n35350 = ~x207 & n35349 ;
  assign n35351 = x299 | n35279 ;
  assign n35352 = x1154 & n35351 ;
  assign n35353 = n35235 | n35352 ;
  assign n35354 = x207 & n35353 ;
  assign n35355 = n35350 | n35354 ;
  assign n35356 = x208 & n35355 ;
  assign n35357 = x299 & ~x1154 ;
  assign n35358 = x1157 & ~n35357 ;
  assign n35359 = n35318 & n35358 ;
  assign n35360 = n35197 | n35219 ;
  assign n35361 = ~x208 & n35360 ;
  assign n35362 = ~x1157 & n35361 ;
  assign n35363 = n35359 | n35362 ;
  assign n35364 = n35356 | n35363 ;
  assign n35365 = x211 | x214 ;
  assign n35366 = x212 & n35365 ;
  assign n35367 = ( x212 & n35364 ) | ( x212 & n35366 ) | ( n35364 & n35366 ) ;
  assign n35368 = ~n35348 & n35367 ;
  assign n35369 = n35309 | n35368 ;
  assign n35370 = ~n35265 & n35369 ;
  assign n35371 = x219 & ~n35370 ;
  assign n35372 = x207 | n35342 ;
  assign n35373 = n35123 & ~n35331 ;
  assign n35374 = x208 & ~n35373 ;
  assign n35375 = n35372 & n35374 ;
  assign n35376 = n35319 & ~n35375 ;
  assign n35377 = x211 | n35376 ;
  assign n35378 = n35253 & ~n35377 ;
  assign n35379 = x207 & n35236 ;
  assign n35380 = n35244 | n35334 ;
  assign n35381 = ~x207 & n35380 ;
  assign n35382 = x299 & x1156 ;
  assign n35383 = x207 & n35382 ;
  assign n35384 = n35381 | n35383 ;
  assign n35385 = n35379 | n35384 ;
  assign n35386 = x208 & n35385 ;
  assign n35387 = n35212 & n35325 ;
  assign n35388 = ~x208 & x1157 ;
  assign n35389 = n35260 | n35382 ;
  assign n35390 = n35388 & n35389 ;
  assign n35391 = n35387 | n35390 ;
  assign n35392 = n35386 | n35391 ;
  assign n35393 = x211 & n35392 ;
  assign n35394 = x214 & ~n35393 ;
  assign n35395 = ~n35378 & n35394 ;
  assign n35396 = n35267 & ~n35395 ;
  assign n35397 = n8652 & n35364 ;
  assign n35398 = ~n8652 & n35365 ;
  assign n35399 = n35307 & n35398 ;
  assign n35400 = ~n35365 & n35392 ;
  assign n35401 = n35399 | n35400 ;
  assign n35402 = n35397 | n35401 ;
  assign n35403 = x212 & n35402 ;
  assign n35404 = x219 | n35403 ;
  assign n35405 = n35396 | n35404 ;
  assign n35406 = ~n6785 & n35405 ;
  assign n35407 = ~n35371 & n35406 ;
  assign n35408 = n35190 | n35407 ;
  assign n35409 = ~x211 & n8894 ;
  assign n35410 = x299 & ~x1143 ;
  assign n35411 = n35335 & ~n35410 ;
  assign n35412 = x299 & x1143 ;
  assign n35413 = ~x1155 & n35412 ;
  assign n35414 = x1154 & ~n35269 ;
  assign n35415 = ~n35413 & n35414 ;
  assign n35416 = ~n35411 & n35415 ;
  assign n35417 = n35241 | n35412 ;
  assign n35418 = ~x1156 & n35417 ;
  assign n35419 = ~n35416 & n35418 ;
  assign n35420 = n35333 | n35410 ;
  assign n35421 = ~x1154 & n35420 ;
  assign n35422 = x299 | n35242 ;
  assign n35423 = x1154 & n35422 ;
  assign n35424 = ~n35412 & n35423 ;
  assign n35425 = x1156 & ~n35424 ;
  assign n35426 = ~n35421 & n35425 ;
  assign n35427 = n35419 | n35426 ;
  assign n35428 = x207 | n35427 ;
  assign n35429 = n35237 & ~n35412 ;
  assign n35430 = x208 & ~n35429 ;
  assign n35431 = n35428 & n35430 ;
  assign n35432 = ~x1157 & n35325 ;
  assign n35433 = ~n35410 & n35432 ;
  assign n35434 = ~n35256 & n35311 ;
  assign n35435 = x207 & ~n35410 ;
  assign n35436 = ~n35434 & n35435 ;
  assign n35437 = n35412 | n35436 ;
  assign n35438 = n35388 & n35437 ;
  assign n35439 = n35433 | n35438 ;
  assign n35440 = n35431 | n35439 ;
  assign n35441 = n35409 & ~n35440 ;
  assign n35442 = ~n8894 & n35100 ;
  assign n35443 = ( x211 & n35440 ) | ( x211 & ~n35442 ) | ( n35440 & ~n35442 ) ;
  assign n35444 = x299 & ~x1144 ;
  assign n35445 = n35335 & ~n35444 ;
  assign n35446 = x299 & x1144 ;
  assign n35447 = ~x1155 & n35446 ;
  assign n35448 = n35414 & ~n35447 ;
  assign n35449 = ~n35445 & n35448 ;
  assign n35450 = n35241 | n35446 ;
  assign n35451 = ~x1156 & n35450 ;
  assign n35452 = ~n35449 & n35451 ;
  assign n35453 = n35333 | n35444 ;
  assign n35454 = ~x1154 & n35453 ;
  assign n35455 = n35423 & ~n35446 ;
  assign n35456 = x1156 & ~n35455 ;
  assign n35457 = ~n35454 & n35456 ;
  assign n35458 = n35452 | n35457 ;
  assign n35459 = x207 | n35458 ;
  assign n35460 = n35237 & ~n35446 ;
  assign n35461 = x208 & ~n35460 ;
  assign n35462 = n35459 & n35461 ;
  assign n35463 = n35432 & ~n35444 ;
  assign n35464 = x207 & ~n35444 ;
  assign n35465 = ~n35434 & n35464 ;
  assign n35466 = n35446 | n35465 ;
  assign n35467 = n35388 & n35466 ;
  assign n35468 = n35463 | n35467 ;
  assign n35469 = n35462 | n35468 ;
  assign n35470 = ( x211 & n35442 ) | ( x211 & ~n35469 ) | ( n35442 & ~n35469 ) ;
  assign n35471 = ~n35443 & n35470 ;
  assign n35472 = n35441 | n35471 ;
  assign n35473 = ~x219 & n35472 ;
  assign n35474 = ~x219 & n35100 ;
  assign n35475 = n35101 | n35474 ;
  assign n35476 = n35264 | n35475 ;
  assign n35477 = ~x299 & n35281 ;
  assign n35478 = x299 & x1142 ;
  assign n35479 = x207 & ~n35478 ;
  assign n35480 = ~n35477 & n35479 ;
  assign n35481 = ~n35154 & n35338 ;
  assign n35482 = n35240 | n35478 ;
  assign n35483 = x1154 | x1156 ;
  assign n35484 = n35482 & ~n35483 ;
  assign n35485 = x207 | n35484 ;
  assign n35486 = n35481 | n35485 ;
  assign n35487 = x208 & n35486 ;
  assign n35488 = ~n35480 & n35487 ;
  assign n35489 = ~n35154 & n35326 ;
  assign n35490 = ~n35319 & n35489 ;
  assign n35491 = n8654 & n35475 ;
  assign n35492 = ~n35490 & n35491 ;
  assign n35493 = ~n35488 & n35492 ;
  assign n35494 = n6785 | n35493 ;
  assign n35495 = n35476 & ~n35494 ;
  assign n35496 = ~n35473 & n35495 ;
  assign n35497 = x213 & ~n35117 ;
  assign n35498 = ~n35496 & n35497 ;
  assign n35499 = x209 | n35498 ;
  assign n35500 = n35408 & ~n35499 ;
  assign n35501 = n35208 | n35500 ;
  assign n35502 = x230 & n35501 ;
  assign n35503 = n35099 & ~n35502 ;
  assign n35504 = x1153 & n35365 ;
  assign n35505 = n35182 & ~n35268 ;
  assign n35506 = n35504 | n35505 ;
  assign n35507 = x212 & n35506 ;
  assign n35508 = x211 & x1153 ;
  assign n35509 = n35181 | n35508 ;
  assign n35510 = n35108 & n35509 ;
  assign n35511 = x219 | n35510 ;
  assign n35512 = n35507 | n35511 ;
  assign n35513 = n35103 & n35512 ;
  assign n35514 = x1152 & ~n35513 ;
  assign n35515 = n8790 | n35248 ;
  assign n35516 = x207 | x208 ;
  assign n35517 = ~n8790 & n35516 ;
  assign n35518 = x1154 | n35224 ;
  assign n35519 = x199 | n35213 ;
  assign n35520 = ~n35221 & n35519 ;
  assign n35521 = n35518 & n35520 ;
  assign n35522 = x207 & n35521 ;
  assign n35523 = n35517 | n35522 ;
  assign n35524 = n35515 & n35523 ;
  assign n35525 = x214 | n35524 ;
  assign n35526 = ~x212 & n35525 ;
  assign n35527 = ~x207 & n35197 ;
  assign n35528 = x207 & n35349 ;
  assign n35529 = n35527 | n35528 ;
  assign n35530 = ~x208 & n35529 ;
  assign n35531 = x1155 | n8980 ;
  assign n35532 = ~n35214 & n35531 ;
  assign n35533 = x299 | n35532 ;
  assign n35534 = n35518 & n35533 ;
  assign n35535 = x207 & n35534 ;
  assign n35536 = n35350 | n35535 ;
  assign n35537 = x208 & n35536 ;
  assign n35538 = n35530 | n35537 ;
  assign n35539 = ~x211 & n35538 ;
  assign n35540 = x207 & ~n35341 ;
  assign n35541 = ~n35338 & n35540 ;
  assign n35542 = n35317 & ~n35541 ;
  assign n35543 = n35123 & ~n35534 ;
  assign n35544 = x208 & ~n35543 ;
  assign n35545 = n35372 & n35544 ;
  assign n35546 = n35542 | n35545 ;
  assign n35547 = ~n35327 & n35546 ;
  assign n35548 = x211 & n35547 ;
  assign n35549 = n35539 | n35548 ;
  assign n35550 = x214 & ~n35549 ;
  assign n35551 = n35526 & ~n35550 ;
  assign n35552 = x219 | n35551 ;
  assign n35553 = ~x214 & n35549 ;
  assign n35554 = x211 | n35547 ;
  assign n35555 = x214 & n35554 ;
  assign n35556 = n35546 & n35555 ;
  assign n35557 = n35553 | n35556 ;
  assign n35558 = x212 & n35557 ;
  assign n35559 = n35552 | n35558 ;
  assign n35560 = ~n35101 & n35524 ;
  assign n35561 = x219 & ~n35560 ;
  assign n35562 = n35101 & n35546 ;
  assign n35563 = n35561 & ~n35562 ;
  assign n35564 = n6785 | n35563 ;
  assign n35565 = n35559 & ~n35564 ;
  assign n35566 = n35514 & ~n35565 ;
  assign n35567 = x211 & ~n35524 ;
  assign n35568 = n35555 & ~n35567 ;
  assign n35569 = n35553 | n35568 ;
  assign n35570 = x212 & n35569 ;
  assign n35571 = n35552 | n35570 ;
  assign n35572 = x219 & ~n35524 ;
  assign n35573 = n6785 | n35572 ;
  assign n35574 = n35571 & ~n35573 ;
  assign n35575 = n8894 | n35509 ;
  assign n35576 = n35474 & n35575 ;
  assign n35577 = ~n35184 & n35576 ;
  assign n35578 = x1152 | n6785 ;
  assign n35579 = ( x1152 & n35577 ) | ( x1152 & n35578 ) | ( n35577 & n35578 ) ;
  assign n35580 = n35574 | n35579 ;
  assign n35581 = ~x213 & n35580 ;
  assign n35582 = ~n35566 & n35581 ;
  assign n35583 = x207 & n35380 ;
  assign n35584 = n35382 | n35583 ;
  assign n35585 = ~x208 & n35584 ;
  assign n35586 = n35384 | n35522 ;
  assign n35587 = x208 & n35586 ;
  assign n35588 = n35585 | n35587 ;
  assign n35589 = ~x211 & n35588 ;
  assign n35590 = n35193 | n35248 ;
  assign n35591 = n35297 & n35590 ;
  assign n35592 = x207 & ~n35193 ;
  assign n35593 = ( n35285 & n35521 ) | ( n35285 & ~n35592 ) | ( n35521 & ~n35592 ) ;
  assign n35594 = n35285 & n35593 ;
  assign n35595 = n35591 | n35594 ;
  assign n35596 = x211 & n35595 ;
  assign n35597 = n35589 | n35596 ;
  assign n35598 = x214 | n35597 ;
  assign n35599 = ( x211 & x214 ) | ( x211 & ~n35595 ) | ( x214 & ~n35595 ) ;
  assign n35600 = ( x211 & ~x214 ) | ( x211 & n35538 ) | ( ~x214 & n35538 ) ;
  assign n35601 = n35599 & ~n35600 ;
  assign n35602 = x212 & ~n35601 ;
  assign n35603 = n35598 & n35602 ;
  assign n35604 = x214 & ~n35597 ;
  assign n35605 = n35526 & ~n35604 ;
  assign n35606 = x219 | n35605 ;
  assign n35607 = n35603 | n35606 ;
  assign n35608 = n35100 & n35539 ;
  assign n35609 = n35561 & ~n35608 ;
  assign n35610 = n32697 & ~n35609 ;
  assign n35611 = n35607 & n35610 ;
  assign n35612 = x209 & ~n35611 ;
  assign n35613 = ~n35582 & n35612 ;
  assign n35614 = x299 | n8980 ;
  assign n35615 = ~x1153 & n35614 ;
  assign n35616 = n35223 & ~n35615 ;
  assign n35617 = x199 | x1153 ;
  assign n35618 = n35216 & n35617 ;
  assign n35619 = n35616 | n35618 ;
  assign n35620 = ( n8790 & n35516 ) | ( n8790 & n35619 ) | ( n35516 & n35619 ) ;
  assign n35621 = x1153 | n8980 ;
  assign n35622 = ~n35221 & n35621 ;
  assign n35623 = ( ~n8790 & n35516 ) | ( ~n8790 & n35622 ) | ( n35516 & n35622 ) ;
  assign n35624 = n35620 & n35623 ;
  assign n35625 = ~n35101 & n35624 ;
  assign n35626 = x200 | x1153 ;
  assign n35627 = ~x199 & n35626 ;
  assign n35628 = x299 | n35627 ;
  assign n35629 = n35290 | n35628 ;
  assign n35630 = x207 & n35629 ;
  assign n35631 = ~n35357 & n35630 ;
  assign n35632 = x1154 & ~n8981 ;
  assign n35633 = n35616 | n35632 ;
  assign n35634 = n35618 | n35633 ;
  assign n35635 = ~x207 & n35634 ;
  assign n35636 = n35631 | n35635 ;
  assign n35637 = x208 & n35636 ;
  assign n35638 = x207 & n35619 ;
  assign n35639 = x208 | n35197 ;
  assign n35640 = n35638 | n35639 ;
  assign n35641 = ( ~x208 & n35637 ) | ( ~x208 & n35640 ) | ( n35637 & n35640 ) ;
  assign n35642 = ~x211 & n35641 ;
  assign n35643 = n35100 & n35642 ;
  assign n35644 = n35625 | n35643 ;
  assign n35645 = x219 & n35644 ;
  assign n35646 = ~x199 & x1153 ;
  assign n35647 = x200 & n35646 ;
  assign n35648 = ~x299 & n35647 ;
  assign n35649 = x1154 | n35648 ;
  assign n35650 = x1154 & n35238 ;
  assign n35651 = ~n35646 & n35650 ;
  assign n35652 = n35649 & ~n35651 ;
  assign n35653 = n35291 | n35652 ;
  assign n35654 = x207 | n35653 ;
  assign n35655 = x207 & ~n35629 ;
  assign n35656 = x208 & ~n35655 ;
  assign n35657 = n35654 & n35656 ;
  assign n35658 = n35297 & n35653 ;
  assign n35659 = n35657 | n35658 ;
  assign n35660 = x199 | x1154 ;
  assign n35661 = x200 | n35660 ;
  assign n35662 = n35132 | n35661 ;
  assign n35663 = ~n35339 & n35662 ;
  assign n35664 = n35659 & n35663 ;
  assign n35665 = x211 & n35664 ;
  assign n35666 = n35382 | n35619 ;
  assign n35667 = ~x207 & n35666 ;
  assign n35668 = x299 & ~x1156 ;
  assign n35669 = n35630 & ~n35668 ;
  assign n35670 = x208 & ~n35669 ;
  assign n35671 = ~n35667 & n35670 ;
  assign n35672 = x208 | n35382 ;
  assign n35673 = n35638 | n35672 ;
  assign n35674 = ~x211 & n35673 ;
  assign n35675 = ~n35671 & n35674 ;
  assign n35676 = n35110 & ~n35675 ;
  assign n35677 = ~n35665 & n35676 ;
  assign n35678 = x214 | n35624 ;
  assign n35679 = x212 | n35678 ;
  assign n35680 = ~x219 & n35679 ;
  assign n35681 = ~n35677 & n35680 ;
  assign n35682 = ( x211 & n8894 ) | ( x211 & ~n35664 ) | ( n8894 & ~n35664 ) ;
  assign n35683 = ( x211 & ~n8894 ) | ( x211 & n35641 ) | ( ~n8894 & n35641 ) ;
  assign n35684 = n35682 & ~n35683 ;
  assign n35685 = n35681 & ~n35684 ;
  assign n35686 = n35645 | n35685 ;
  assign n35687 = ( x1152 & n6785 ) | ( x1152 & ~n35686 ) | ( n6785 & ~n35686 ) ;
  assign n35688 = x299 | n35647 ;
  assign n35689 = ~x1154 & n35688 ;
  assign n35690 = ~n35339 & n35689 ;
  assign n35691 = x1153 & ~n9515 ;
  assign n35692 = n35272 & ~n35691 ;
  assign n35693 = x1154 & ~n35692 ;
  assign n35694 = ~n35302 & n35693 ;
  assign n35695 = n35690 | n35694 ;
  assign n35696 = x299 | x1153 ;
  assign n35697 = ~n8981 & n35696 ;
  assign n35698 = ~n35339 & n35697 ;
  assign n35699 = x207 & ~n35698 ;
  assign n35700 = x208 & ~n35699 ;
  assign n35701 = ( x207 & n35695 ) | ( x207 & n35700 ) | ( n35695 & n35700 ) ;
  assign n35702 = x207 & ~n35700 ;
  assign n35703 = ( n35297 & n35701 ) | ( n35297 & ~n35702 ) | ( n35701 & ~n35702 ) ;
  assign n35704 = x211 & ~n35703 ;
  assign n35705 = x200 & ~x1153 ;
  assign n35706 = n9520 | n35705 ;
  assign n35707 = x1154 & n35706 ;
  assign n35708 = n35649 & ~n35707 ;
  assign n35709 = n35517 & n35708 ;
  assign n35710 = x208 & n35123 ;
  assign n35711 = x1153 & ~n8981 ;
  assign n35712 = n35710 & n35711 ;
  assign n35713 = n35709 | n35712 ;
  assign n35714 = x211 | n35382 ;
  assign n35715 = n35713 | n35714 ;
  assign n35716 = n35110 & n35715 ;
  assign n35717 = ~n35704 & n35716 ;
  assign n35718 = ( x211 & n8894 ) | ( x211 & n35703 ) | ( n8894 & n35703 ) ;
  assign n35719 = n35648 | n35693 ;
  assign n35720 = x207 & n35719 ;
  assign n35721 = n35527 | n35720 ;
  assign n35722 = ~x208 & n35721 ;
  assign n35723 = ( x207 & x208 ) | ( x207 & n35719 ) | ( x208 & n35719 ) ;
  assign n35724 = ~n35357 & n35697 ;
  assign n35725 = ( ~x207 & x208 ) | ( ~x207 & n35724 ) | ( x208 & n35724 ) ;
  assign n35726 = n35723 & n35725 ;
  assign n35727 = n35722 | n35726 ;
  assign n35728 = ( ~x211 & n8894 ) | ( ~x211 & n35727 ) | ( n8894 & n35727 ) ;
  assign n35729 = n35718 & n35728 ;
  assign n35730 = n35717 | n35729 ;
  assign n35731 = ~x219 & n35730 ;
  assign n35732 = ~n35100 & n35713 ;
  assign n35733 = x211 | n35727 ;
  assign n35734 = x219 & n35100 ;
  assign n35735 = x211 & ~n35713 ;
  assign n35736 = n35734 & ~n35735 ;
  assign n35737 = n35733 & n35736 ;
  assign n35738 = n35732 | n35737 ;
  assign n35739 = n35731 | n35738 ;
  assign n35740 = ( x1152 & ~n6785 ) | ( x1152 & n35739 ) | ( ~n6785 & n35739 ) ;
  assign n35741 = ~n35687 & n35740 ;
  assign n35742 = ( x209 & x213 ) | ( x209 & n35741 ) | ( x213 & n35741 ) ;
  assign n35743 = n35317 & n35653 ;
  assign n35744 = n35657 | n35743 ;
  assign n35745 = x211 | n35744 ;
  assign n35746 = x211 & ~n35624 ;
  assign n35747 = n35745 & ~n35746 ;
  assign n35748 = n35100 & n35747 ;
  assign n35749 = x219 & ~n35624 ;
  assign n35750 = n35734 | n35749 ;
  assign n35751 = ~n35748 & n35750 ;
  assign n35752 = n6785 | n35751 ;
  assign n35753 = ~x212 & n35678 ;
  assign n35754 = ~x207 & n35195 ;
  assign n35755 = ~x1153 & n35230 ;
  assign n35756 = n35301 & ~n35755 ;
  assign n35757 = x1154 & ~n9515 ;
  assign n35758 = ~n35755 & n35757 ;
  assign n35759 = n35756 | n35758 ;
  assign n35760 = x207 & n35759 ;
  assign n35761 = n35754 | n35760 ;
  assign n35762 = ~x208 & n35761 ;
  assign n35763 = ~x207 & n35759 ;
  assign n35764 = ~x299 & n35214 ;
  assign n35765 = x207 & ~n35764 ;
  assign n35766 = n35272 & n35765 ;
  assign n35767 = n35763 | n35766 ;
  assign n35768 = x208 & n35767 ;
  assign n35769 = n35762 | n35768 ;
  assign n35770 = x211 & n35769 ;
  assign n35771 = n35642 | n35770 ;
  assign n35772 = x214 & ~n35771 ;
  assign n35773 = n35753 & ~n35772 ;
  assign n35774 = x214 | n35771 ;
  assign n35775 = x211 & n35744 ;
  assign n35776 = ~x211 & n35769 ;
  assign n35777 = n35775 | n35776 ;
  assign n35778 = ( x212 & n35109 ) | ( x212 & n35777 ) | ( n35109 & n35777 ) ;
  assign n35779 = n35774 & n35778 ;
  assign n35780 = x219 | n35779 ;
  assign n35781 = n35773 | n35780 ;
  assign n35782 = ~n35752 & n35781 ;
  assign n35783 = n35514 & ~n35782 ;
  assign n35784 = x1153 & ~x1154 ;
  assign n35785 = n35320 & n35784 ;
  assign n35786 = n35758 | n35785 ;
  assign n35787 = x207 & n35786 ;
  assign n35788 = n35754 | n35787 ;
  assign n35789 = ~x208 & n35788 ;
  assign n35790 = ~x207 & n35786 ;
  assign n35791 = x207 & ~n8981 ;
  assign n35792 = x1153 & n35791 ;
  assign n35793 = n35790 | n35792 ;
  assign n35794 = x208 & n35793 ;
  assign n35795 = n35789 | n35794 ;
  assign n35796 = n35409 & ~n35795 ;
  assign n35797 = x211 & ~n35795 ;
  assign n35798 = n35733 & ~n35797 ;
  assign n35799 = n35442 & ~n35798 ;
  assign n35800 = n35796 | n35799 ;
  assign n35801 = ~x219 & n35800 ;
  assign n35802 = x219 & ~n35713 ;
  assign n35803 = n6785 | n35802 ;
  assign n35804 = n35268 | n35442 ;
  assign n35805 = n35713 | n35804 ;
  assign n35806 = ~n35803 & n35805 ;
  assign n35807 = ~n35801 & n35806 ;
  assign n35808 = n35579 | n35807 ;
  assign n35809 = ~n35783 & n35808 ;
  assign n35810 = ( x209 & ~x213 ) | ( x209 & n35809 ) | ( ~x213 & n35809 ) ;
  assign n35811 = n35742 | n35810 ;
  assign n35812 = ~n35613 & n35811 ;
  assign n35813 = x214 & n35166 ;
  assign n35814 = ~x212 & n35813 ;
  assign n35815 = x219 | n35814 ;
  assign n35816 = n35173 | n35815 ;
  assign n35817 = x219 & ~n35181 ;
  assign n35818 = x213 & ~n35817 ;
  assign n35819 = n35103 & n35818 ;
  assign n35820 = n35816 & n35819 ;
  assign n35821 = n35812 | n35820 ;
  assign n35822 = x230 & n35821 ;
  assign n35823 = ~x230 & x234 ;
  assign n35824 = n35822 | n35823 ;
  assign n35825 = ~x1156 & n35240 ;
  assign n35826 = n8790 & ~n35247 ;
  assign n35827 = ~n35825 & n35826 ;
  assign n35828 = x207 | n35218 ;
  assign n35829 = ~n35827 & n35828 ;
  assign n35830 = n35220 & n35829 ;
  assign n35831 = x1157 | n35830 ;
  assign n35832 = ~x207 & n35259 ;
  assign n35833 = n35827 | n35832 ;
  assign n35834 = n35261 & ~n35833 ;
  assign n35835 = x1157 & ~n35834 ;
  assign n35836 = n35831 & ~n35835 ;
  assign n35837 = n35100 | n35836 ;
  assign n35838 = n35334 | n35825 ;
  assign n35839 = x207 & n35838 ;
  assign n35840 = ~x207 & n35323 ;
  assign n35841 = x208 & ~n35840 ;
  assign n35842 = ~n35839 & n35841 ;
  assign n35843 = ( x208 & n35387 ) | ( x208 & ~n35842 ) | ( n35387 & ~n35842 ) ;
  assign n35844 = ~x1157 & n35843 ;
  assign n35845 = x208 & x1157 ;
  assign n35846 = n35258 & ~n35314 ;
  assign n35847 = x207 | n35846 ;
  assign n35848 = ~n35839 & n35847 ;
  assign n35849 = n35845 & ~n35848 ;
  assign n35850 = n35390 | n35849 ;
  assign n35851 = n35844 | n35850 ;
  assign n35852 = x211 & n35851 ;
  assign n35853 = ~x207 & n35315 ;
  assign n35854 = x208 & ~n35853 ;
  assign n35855 = ~n35334 & n35540 ;
  assign n35856 = n35854 & ~n35855 ;
  assign n35857 = n35318 | n35856 ;
  assign n35858 = x1157 & ~n35857 ;
  assign n35859 = ~x211 & n35831 ;
  assign n35860 = ~n35858 & n35859 ;
  assign n35861 = n35442 & ~n35860 ;
  assign n35862 = ~n35852 & n35861 ;
  assign n35863 = n35837 & ~n35862 ;
  assign n35864 = n35247 | n35340 ;
  assign n35865 = x207 & n35864 ;
  assign n35866 = ~x207 & n35304 ;
  assign n35867 = n35865 | n35866 ;
  assign n35868 = x208 & n35867 ;
  assign n35869 = n35305 | n35868 ;
  assign n35870 = ~x1157 & n35869 ;
  assign n35871 = x207 | n35295 ;
  assign n35872 = ~n35865 & n35871 ;
  assign n35873 = n35845 & ~n35872 ;
  assign n35874 = n35299 | n35873 ;
  assign n35875 = n35870 | n35874 ;
  assign n35876 = ( x211 & ~n8894 ) | ( x211 & n35875 ) | ( ~n8894 & n35875 ) ;
  assign n35877 = ( x211 & n8894 ) | ( x211 & ~n35851 ) | ( n8894 & ~n35851 ) ;
  assign n35878 = ~n35876 & n35877 ;
  assign n35879 = n35863 & ~n35878 ;
  assign n35880 = x219 | n35879 ;
  assign n35881 = x211 | n35875 ;
  assign n35882 = x211 & ~n35836 ;
  assign n35883 = n35110 & ~n35882 ;
  assign n35884 = n35881 & n35883 ;
  assign n35885 = ~n35110 & n35836 ;
  assign n35886 = x219 & ~n35885 ;
  assign n35887 = ~n35884 & n35886 ;
  assign n35888 = x209 & ~n35887 ;
  assign n35889 = n35880 & n35888 ;
  assign n35890 = n8790 & ~n35708 ;
  assign n35891 = ( x207 & x208 ) | ( x207 & n35236 ) | ( x208 & n35236 ) ;
  assign n35892 = ~n35890 & n35891 ;
  assign n35893 = n35382 | n35892 ;
  assign n35894 = x211 & ~n35893 ;
  assign n35895 = n35317 & ~n35373 ;
  assign n35896 = n35689 | n35693 ;
  assign n35897 = x207 & ~n35896 ;
  assign n35898 = n35132 | n35331 ;
  assign n35899 = x208 & n35898 ;
  assign n35900 = ~n35897 & n35899 ;
  assign n35901 = n35895 | n35900 ;
  assign n35902 = ( x211 & x1157 ) | ( x211 & n35901 ) | ( x1157 & n35901 ) ;
  assign n35903 = ( x211 & ~x1157 ) | ( x211 & n35892 ) | ( ~x1157 & n35892 ) ;
  assign n35904 = n35902 | n35903 ;
  assign n35905 = ~n35894 & n35904 ;
  assign n35906 = n35442 & ~n35905 ;
  assign n35907 = n35100 | n35892 ;
  assign n35908 = n35281 & n35297 ;
  assign n35909 = x207 | n35281 ;
  assign n35910 = x207 & ~n35695 ;
  assign n35911 = x208 & ~n35910 ;
  assign n35912 = n35909 & n35911 ;
  assign n35913 = n35908 | n35912 ;
  assign n35914 = ( x211 & ~n8894 ) | ( x211 & n35913 ) | ( ~n8894 & n35913 ) ;
  assign n35915 = ( x211 & n8894 ) | ( x211 & ~n35893 ) | ( n8894 & ~n35893 ) ;
  assign n35916 = ~n35914 & n35915 ;
  assign n35917 = n35907 & ~n35916 ;
  assign n35918 = ~n35906 & n35917 ;
  assign n35919 = x219 | n35918 ;
  assign n35920 = x211 | n35913 ;
  assign n35921 = x211 & ~n35892 ;
  assign n35922 = n35110 & ~n35921 ;
  assign n35923 = n35920 & n35922 ;
  assign n35924 = ~n35110 & n35892 ;
  assign n35925 = x219 & ~n35924 ;
  assign n35926 = ~n35923 & n35925 ;
  assign n35927 = x209 | n35926 ;
  assign n35928 = n35919 & ~n35927 ;
  assign n35929 = n35889 | n35928 ;
  assign n35930 = ~n6785 & n35929 ;
  assign n35931 = ~x214 & n35176 ;
  assign n35932 = n35813 | n35931 ;
  assign n35933 = x212 & n35932 ;
  assign n35934 = x219 | n35933 ;
  assign n35935 = n35178 | n35934 ;
  assign n35936 = x219 & ~n35168 ;
  assign n35937 = x219 & ~n35442 ;
  assign n35938 = n35936 | n35937 ;
  assign n35939 = n35935 & ~n35938 ;
  assign n35940 = ( x213 & n32697 ) | ( x213 & ~n35939 ) | ( n32697 & ~n35939 ) ;
  assign n35941 = ~n35930 & n35940 ;
  assign n35942 = n8894 & n35509 ;
  assign n35943 = n35170 & n35442 ;
  assign n35944 = x219 | n35943 ;
  assign n35945 = n35942 | n35944 ;
  assign n35946 = x219 & ~n35183 ;
  assign n35947 = n6785 & ~n35946 ;
  assign n35948 = ~n35937 & n35947 ;
  assign n35949 = n35945 & n35948 ;
  assign n35950 = x213 | n35949 ;
  assign n35951 = n35332 | n35754 ;
  assign n35952 = ~x208 & n35951 ;
  assign n35953 = ~x207 & n35331 ;
  assign n35954 = n35787 | n35953 ;
  assign n35955 = x208 & n35954 ;
  assign n35956 = n35952 | n35955 ;
  assign n35957 = x211 | n35956 ;
  assign n35958 = n35922 & n35957 ;
  assign n35959 = n35925 & ~n35958 ;
  assign n35960 = n35354 | n35527 ;
  assign n35961 = ~x208 & n35960 ;
  assign n35962 = ~x207 & n35353 ;
  assign n35963 = n35720 | n35962 ;
  assign n35964 = x208 & n35963 ;
  assign n35965 = n35961 | n35964 ;
  assign n35966 = x211 & ~n35965 ;
  assign n35967 = n35920 & ~n35966 ;
  assign n35968 = n35110 & ~n35967 ;
  assign n35969 = ( x211 & ~n8894 ) | ( x211 & n35956 ) | ( ~n8894 & n35956 ) ;
  assign n35970 = ( x211 & n8894 ) | ( x211 & ~n35965 ) | ( n8894 & ~n35965 ) ;
  assign n35971 = ~n35969 & n35970 ;
  assign n35972 = n35907 & ~n35971 ;
  assign n35973 = ~n35968 & n35972 ;
  assign n35974 = x219 | n35973 ;
  assign n35975 = ~n35959 & n35974 ;
  assign n35976 = ( x209 & ~n6785 ) | ( x209 & n35975 ) | ( ~n6785 & n35975 ) ;
  assign n35977 = ( x1157 & n35844 ) | ( x1157 & n35857 ) | ( n35844 & n35857 ) ;
  assign n35978 = ( x299 & ~x1157 ) | ( x299 & n35844 ) | ( ~x1157 & n35844 ) ;
  assign n35979 = n35977 | n35978 ;
  assign n35980 = ~n35327 & n35979 ;
  assign n35981 = x211 | n35980 ;
  assign n35982 = n35883 & n35981 ;
  assign n35983 = n35886 & ~n35982 ;
  assign n35984 = n35241 & n35341 ;
  assign n35985 = n35247 | n35984 ;
  assign n35986 = x207 & n35985 ;
  assign n35987 = x1154 & ~n35322 ;
  assign n35988 = n35217 | n35987 ;
  assign n35989 = ~x207 & n35300 ;
  assign n35990 = n35988 & n35989 ;
  assign n35991 = n35986 | n35990 ;
  assign n35992 = x208 & n35991 ;
  assign n35993 = n35361 | n35992 ;
  assign n35994 = ~x1157 & n35993 ;
  assign n35995 = n35358 & n35857 ;
  assign n35996 = n35994 | n35995 ;
  assign n35997 = x211 & ~n35996 ;
  assign n35998 = n35881 & ~n35997 ;
  assign n35999 = n35442 & ~n35998 ;
  assign n36000 = n35837 & ~n35999 ;
  assign n36001 = ( x211 & n8894 ) | ( x211 & ~n35996 ) | ( n8894 & ~n35996 ) ;
  assign n36002 = ( x211 & ~n8894 ) | ( x211 & n35980 ) | ( ~n8894 & n35980 ) ;
  assign n36003 = n36001 & ~n36002 ;
  assign n36004 = n36000 & ~n36003 ;
  assign n36005 = x219 | n36004 ;
  assign n36006 = ~n35983 & n36005 ;
  assign n36007 = ( x209 & n6785 ) | ( x209 & ~n36006 ) | ( n6785 & ~n36006 ) ;
  assign n36008 = n35976 & ~n36007 ;
  assign n36009 = n35950 | n36008 ;
  assign n36010 = ~n35941 & n36009 ;
  assign n36011 = x230 & ~n36010 ;
  assign n36012 = x230 | x235 ;
  assign n36013 = ~n36011 & n36012 ;
  assign n36014 = ~x100 & n34886 ;
  assign n36015 = n4812 | n36014 ;
  assign n36016 = ~n4816 & n36015 ;
  assign n36017 = ( x75 & ~n5763 ) | ( x75 & n36016 ) | ( ~n5763 & n36016 ) ;
  assign n36018 = x92 | n36017 ;
  assign n36019 = ~n11665 & n36018 ;
  assign n36020 = x74 | n36019 ;
  assign n36021 = ~n4657 & n36020 ;
  assign n36022 = x56 | n36021 ;
  assign n36023 = ~n4653 & n36022 ;
  assign n36024 = x62 | n36023 ;
  assign n36025 = ~n4828 & n36024 ;
  assign n36026 = ~x211 & x1145 ;
  assign n36027 = x211 & x1144 ;
  assign n36028 = n36026 | n36027 ;
  assign n36029 = ( n8894 & n35100 ) | ( n8894 & n36028 ) | ( n35100 & n36028 ) ;
  assign n36030 = ( ~n8894 & n35100 ) | ( ~n8894 & n35107 ) | ( n35100 & n35107 ) ;
  assign n36031 = n36029 & n36030 ;
  assign n36032 = x219 | n36031 ;
  assign n36033 = x219 & ~n35112 ;
  assign n36034 = n35103 & ~n36033 ;
  assign n36035 = n36032 & n36034 ;
  assign n36036 = n35191 & n36031 ;
  assign n36037 = x199 & x1143 ;
  assign n36038 = x200 | n36037 ;
  assign n36039 = n35128 | n36038 ;
  assign n36040 = ~n35130 & n35710 ;
  assign n36041 = n36039 & n36040 ;
  assign n36042 = ~x199 & x1145 ;
  assign n36043 = n36038 | n36042 ;
  assign n36044 = x200 & ~n35128 ;
  assign n36045 = n35517 & ~n36044 ;
  assign n36046 = n36043 & n36045 ;
  assign n36047 = n36041 | n36046 ;
  assign n36048 = ~x299 & n36047 ;
  assign n36049 = x299 & n35734 ;
  assign n36050 = n35112 & n36049 ;
  assign n36051 = n36048 | n36050 ;
  assign n36052 = n36036 | n36051 ;
  assign n36053 = ~n6785 & n36052 ;
  assign n36054 = n36035 | n36053 ;
  assign n36055 = x213 & ~n36054 ;
  assign n36056 = x211 & x1157 ;
  assign n36057 = ~x211 & x1158 ;
  assign n36058 = n36056 | n36057 ;
  assign n36059 = n35108 & n36058 ;
  assign n36060 = n35934 | n36059 ;
  assign n36061 = ~x219 & n6785 ;
  assign n36062 = n35108 & n35164 ;
  assign n36063 = n6785 & n36062 ;
  assign n36064 = n36061 | n36063 ;
  assign n36065 = x214 & n35181 ;
  assign n36066 = x1155 & ~n35365 ;
  assign n36067 = n36065 | n36066 ;
  assign n36068 = x212 & n36067 ;
  assign n36069 = n6785 & n36068 ;
  assign n36070 = n36064 | n36069 ;
  assign n36071 = n36060 & n36070 ;
  assign n36072 = x213 | n36071 ;
  assign n36073 = n35191 & n36060 ;
  assign n36074 = n35108 & n35382 ;
  assign n36075 = ( x212 & ~x214 ) | ( x212 & n35197 ) | ( ~x214 & n35197 ) ;
  assign n36076 = ( x212 & x214 ) | ( x212 & n35193 ) | ( x214 & n35193 ) ;
  assign n36077 = n36075 & n36076 ;
  assign n36078 = n36074 | n36077 ;
  assign n36079 = n35201 & n36078 ;
  assign n36080 = n36048 | n36079 ;
  assign n36081 = n36073 | n36080 ;
  assign n36082 = ~n6785 & n36081 ;
  assign n36083 = n36072 | n36082 ;
  assign n36084 = x209 & n36083 ;
  assign n36085 = ~n36055 & n36084 ;
  assign n36086 = n35136 & ~n35230 ;
  assign n36087 = x1158 & ~n35614 ;
  assign n36088 = x199 | x1158 ;
  assign n36089 = x1156 & n36088 ;
  assign n36090 = n36087 | n36089 ;
  assign n36091 = n36086 & n36090 ;
  assign n36092 = x207 & ~n35248 ;
  assign n36093 = x208 & n35828 ;
  assign n36094 = ~n36092 & n36093 ;
  assign n36095 = n36091 | n36094 ;
  assign n36096 = ~x1157 & n36095 ;
  assign n36097 = ~n35541 & n35854 ;
  assign n36098 = x1156 & n35290 ;
  assign n36099 = x200 | x1158 ;
  assign n36100 = ~x199 & n36099 ;
  assign n36101 = n36098 | n36100 ;
  assign n36102 = n35123 & n36101 ;
  assign n36103 = ( ~x208 & x299 ) | ( ~x208 & n36102 ) | ( x299 & n36102 ) ;
  assign n36104 = n36097 | n36103 ;
  assign n36105 = x1157 & n36104 ;
  assign n36106 = n36096 | n36105 ;
  assign n36107 = x211 & ~n36106 ;
  assign n36108 = x207 | n35315 ;
  assign n36109 = x299 & ~x1158 ;
  assign n36110 = n36108 | n36109 ;
  assign n36111 = ( x207 & ~x1158 ) | ( x207 & n35342 ) | ( ~x1158 & n35342 ) ;
  assign n36112 = ( x207 & x1158 ) | ( x207 & n35248 ) | ( x1158 & n35248 ) ;
  assign n36113 = n36111 & n36112 ;
  assign n36114 = n36110 & ~n36113 ;
  assign n36115 = n35845 & ~n36114 ;
  assign n36116 = x299 | n35323 ;
  assign n36117 = x207 | n36109 ;
  assign n36118 = n36116 & ~n36117 ;
  assign n36119 = x208 & ~n36118 ;
  assign n36120 = ~n36113 & n36119 ;
  assign n36121 = x299 | n35791 ;
  assign n36122 = x1158 & n36121 ;
  assign n36123 = n35123 & n36098 ;
  assign n36124 = x208 | n36123 ;
  assign n36125 = n36122 | n36124 ;
  assign n36126 = ~x1157 & n36125 ;
  assign n36127 = ~n36120 & n36126 ;
  assign n36128 = n35216 & n35293 ;
  assign n36129 = x1157 & ~n36087 ;
  assign n36130 = ~n36128 & n36129 ;
  assign n36131 = x207 & ~n36130 ;
  assign n36132 = n36122 | n36131 ;
  assign n36133 = n35388 & n36132 ;
  assign n36134 = x211 | n36133 ;
  assign n36135 = n36127 | n36134 ;
  assign n36136 = n36115 | n36135 ;
  assign n36137 = ~n36107 & n36136 ;
  assign n36138 = x214 & ~n36137 ;
  assign n36139 = ~x208 & n36102 ;
  assign n36140 = x208 & ~n35832 ;
  assign n36141 = ~n36092 & n36140 ;
  assign n36142 = n36139 | n36141 ;
  assign n36143 = x1157 & n36142 ;
  assign n36144 = n36096 | n36143 ;
  assign n36145 = ( ~x212 & n35108 ) | ( ~x212 & n36144 ) | ( n35108 & n36144 ) ;
  assign n36146 = ~n36138 & n36145 ;
  assign n36147 = ~n35365 & n36106 ;
  assign n36148 = ~n35583 & n35841 ;
  assign n36149 = ~x200 & x207 ;
  assign n36150 = n36090 & n36149 ;
  assign n36151 = n35672 | n36150 ;
  assign n36152 = ~x1157 & n36151 ;
  assign n36153 = ~n36148 & n36152 ;
  assign n36154 = ~n35583 & n35847 ;
  assign n36155 = n35845 & ~n36154 ;
  assign n36156 = n35382 | n36102 ;
  assign n36157 = n35388 & n36156 ;
  assign n36158 = n36155 | n36157 ;
  assign n36159 = n36153 | n36158 ;
  assign n36160 = n35398 & n36159 ;
  assign n36161 = x207 & n35590 ;
  assign n36162 = n35866 | n36161 ;
  assign n36163 = ( x208 & n36091 ) | ( x208 & n36162 ) | ( n36091 & n36162 ) ;
  assign n36164 = ( ~x208 & n35193 ) | ( ~x208 & n36091 ) | ( n35193 & n36091 ) ;
  assign n36165 = n36163 | n36164 ;
  assign n36166 = ~x1157 & n36165 ;
  assign n36167 = n35871 & ~n36161 ;
  assign n36168 = n35845 & ~n36167 ;
  assign n36169 = x1156 & ~n35764 ;
  assign n36170 = x1158 | n35216 ;
  assign n36171 = n36169 & n36170 ;
  assign n36172 = n36100 | n36171 ;
  assign n36173 = n35123 & n36172 ;
  assign n36174 = n35193 | n36173 ;
  assign n36175 = n35388 & n36174 ;
  assign n36176 = n36168 | n36175 ;
  assign n36177 = n36166 | n36176 ;
  assign n36178 = n8652 & n36177 ;
  assign n36179 = n36160 | n36178 ;
  assign n36180 = n36147 | n36179 ;
  assign n36181 = x212 & n36180 ;
  assign n36182 = x219 | n36181 ;
  assign n36183 = n36146 | n36182 ;
  assign n36184 = n35101 | n36144 ;
  assign n36185 = n35108 & ~n36159 ;
  assign n36186 = ~x214 & n36177 ;
  assign n36187 = x208 & ~n35528 ;
  assign n36188 = x1157 | n36091 ;
  assign n36189 = n35990 | n36188 ;
  assign n36190 = n35358 & ~n36108 ;
  assign n36191 = ( ~x1157 & n36189 ) | ( ~x1157 & n36190 ) | ( n36189 & n36190 ) ;
  assign n36192 = n36187 & ~n36191 ;
  assign n36193 = n36173 & n36188 ;
  assign n36194 = n35639 | n36193 ;
  assign n36195 = ~n36192 & n36194 ;
  assign n36196 = ( x212 & n35109 ) | ( x212 & ~n36195 ) | ( n35109 & ~n36195 ) ;
  assign n36197 = ~n36186 & n36196 ;
  assign n36198 = n36185 | n36197 ;
  assign n36199 = ~x211 & n36198 ;
  assign n36200 = n36184 & ~n36199 ;
  assign n36201 = x219 & ~n36200 ;
  assign n36202 = n6785 | n36201 ;
  assign n36203 = n36183 & ~n36202 ;
  assign n36204 = n36072 | n36203 ;
  assign n36205 = x299 & ~x1145 ;
  assign n36206 = n35333 | n36205 ;
  assign n36207 = ~x1154 & n36206 ;
  assign n36208 = x299 & x1145 ;
  assign n36209 = n35423 & ~n36208 ;
  assign n36210 = x1156 & ~n36209 ;
  assign n36211 = ~n36207 & n36210 ;
  assign n36212 = n35241 | n36208 ;
  assign n36213 = ~x1156 & n36212 ;
  assign n36214 = n35337 & ~n36205 ;
  assign n36215 = ( ~x1154 & n36213 ) | ( ~x1154 & n36214 ) | ( n36213 & n36214 ) ;
  assign n36216 = n36211 | n36215 ;
  assign n36217 = x207 & n36216 ;
  assign n36218 = ~x200 & x1157 ;
  assign n36219 = ~x199 & n36218 ;
  assign n36220 = n36116 | n36219 ;
  assign n36221 = x207 | n36205 ;
  assign n36222 = n36220 & ~n36221 ;
  assign n36223 = x208 & ~n36222 ;
  assign n36224 = ~n36217 & n36223 ;
  assign n36225 = ~x299 & n36098 ;
  assign n36226 = x1157 | n36087 ;
  assign n36227 = n36225 | n36226 ;
  assign n36228 = n36131 & n36227 ;
  assign n36229 = x208 | n36208 ;
  assign n36230 = n36228 | n36229 ;
  assign n36231 = ~n36224 & n36230 ;
  assign n36232 = x211 | n36231 ;
  assign n36233 = x1157 | n36150 ;
  assign n36234 = ~x208 & n36233 ;
  assign n36235 = n36173 & n36234 ;
  assign n36236 = x208 | n36235 ;
  assign n36237 = n35446 | n36236 ;
  assign n36238 = x207 & n35458 ;
  assign n36239 = x207 | n35444 ;
  assign n36240 = n36220 & ~n36239 ;
  assign n36241 = x208 & ~n36240 ;
  assign n36242 = ~n36238 & n36241 ;
  assign n36243 = n36237 & ~n36242 ;
  assign n36244 = x211 & ~n36243 ;
  assign n36245 = n36232 & ~n36244 ;
  assign n36246 = x214 | n36245 ;
  assign n36247 = ( x211 & x214 ) | ( x211 & ~n36243 ) | ( x214 & ~n36243 ) ;
  assign n36248 = n35412 | n36236 ;
  assign n36249 = x207 & n35427 ;
  assign n36250 = x207 | n35410 ;
  assign n36251 = n36220 & ~n36250 ;
  assign n36252 = x208 & ~n36251 ;
  assign n36253 = ~n36249 & n36252 ;
  assign n36254 = n36248 & ~n36253 ;
  assign n36255 = ( x211 & ~x214 ) | ( x211 & n36254 ) | ( ~x214 & n36254 ) ;
  assign n36256 = n36247 & ~n36255 ;
  assign n36257 = x212 & ~n36256 ;
  assign n36258 = n36246 & n36257 ;
  assign n36259 = x214 & ~n36245 ;
  assign n36260 = n36145 & ~n36259 ;
  assign n36261 = x219 | n36260 ;
  assign n36262 = n36258 | n36261 ;
  assign n36263 = n35101 & ~n36254 ;
  assign n36264 = n36184 & ~n36263 ;
  assign n36265 = x219 & ~n36264 ;
  assign n36266 = n6785 | n36265 ;
  assign n36267 = n36262 & ~n36266 ;
  assign n36268 = x213 & ~n36035 ;
  assign n36269 = ~n36267 & n36268 ;
  assign n36270 = x209 | n36269 ;
  assign n36271 = n36204 & ~n36270 ;
  assign n36272 = n36085 | n36271 ;
  assign n36273 = x230 & n36272 ;
  assign n36274 = x230 | x237 ;
  assign n36275 = ~n36273 & n36274 ;
  assign n36276 = x211 | x1153 ;
  assign n36277 = x219 & ~n36276 ;
  assign n36278 = n35103 & ~n36277 ;
  assign n36279 = n35945 & n36278 ;
  assign n36280 = n35216 & n35784 ;
  assign n36281 = n35633 | n36280 ;
  assign n36282 = x207 & n36281 ;
  assign n36283 = n35962 | n36282 ;
  assign n36284 = x208 & n36283 ;
  assign n36285 = n35961 | n36284 ;
  assign n36286 = n35398 & n36285 ;
  assign n36287 = n35221 & n35699 ;
  assign n36288 = ~x1154 & n35696 ;
  assign n36289 = n35301 & n36288 ;
  assign n36290 = x207 & ~n36289 ;
  assign n36291 = ~n35633 & n36290 ;
  assign n36292 = x208 & ~n36291 ;
  assign n36293 = ~n36287 & n36292 ;
  assign n36294 = n35909 & n36293 ;
  assign n36295 = n35908 | n36294 ;
  assign n36296 = ~n35365 & n36295 ;
  assign n36297 = x1153 & n35301 ;
  assign n36298 = n35616 | n36297 ;
  assign n36299 = x207 & n36298 ;
  assign n36300 = n35953 | n36299 ;
  assign n36301 = x208 & n36300 ;
  assign n36302 = n35952 | n36301 ;
  assign n36303 = n8652 & n36302 ;
  assign n36304 = x212 & ~n36303 ;
  assign n36305 = ~n36296 & n36304 ;
  assign n36306 = ~n36286 & n36305 ;
  assign n36307 = ( x211 & n35108 ) | ( x211 & ~n36295 ) | ( n35108 & ~n36295 ) ;
  assign n36308 = ( x211 & ~n35108 ) | ( x211 & n36285 ) | ( ~n35108 & n36285 ) ;
  assign n36309 = n36307 & ~n36308 ;
  assign n36310 = n36306 | n36309 ;
  assign n36311 = ~x219 & n36310 ;
  assign n36312 = n8790 & ~n36280 ;
  assign n36313 = ~n35616 & n36312 ;
  assign n36314 = n35891 & ~n36313 ;
  assign n36315 = x211 & n36314 ;
  assign n36316 = ~x211 & n36302 ;
  assign n36317 = n36315 | n36316 ;
  assign n36318 = n35734 & ~n36317 ;
  assign n36319 = x214 | n36314 ;
  assign n36320 = x212 | n36319 ;
  assign n36321 = ~n6785 & n36320 ;
  assign n36322 = ~n36318 & n36321 ;
  assign n36323 = ~n36311 & n36322 ;
  assign n36324 = ( x209 & n36279 ) | ( x209 & n36323 ) | ( n36279 & n36323 ) ;
  assign n36325 = n8790 | n35230 ;
  assign n36326 = n35516 & ~n36325 ;
  assign n36327 = n35215 & n35710 ;
  assign n36328 = n36326 | n36327 ;
  assign n36329 = n35621 & n36328 ;
  assign n36330 = x214 | n36329 ;
  assign n36331 = ~x212 & n36330 ;
  assign n36332 = ~n35230 & n35617 ;
  assign n36333 = ~x1153 & n35291 ;
  assign n36334 = n35271 | n36333 ;
  assign n36335 = x1155 & n36334 ;
  assign n36336 = n36332 | n36335 ;
  assign n36337 = n35123 & ~n35215 ;
  assign n36338 = x208 & ~n36337 ;
  assign n36339 = n35297 | n36338 ;
  assign n36340 = n36336 & n36339 ;
  assign n36341 = n36327 | n36340 ;
  assign n36342 = ~x299 & n36341 ;
  assign n36343 = x299 & n35170 ;
  assign n36344 = x214 & ~n36343 ;
  assign n36345 = ~n36342 & n36344 ;
  assign n36346 = n36331 & ~n36345 ;
  assign n36347 = n35365 | n36341 ;
  assign n36348 = x299 | n36149 ;
  assign n36349 = ~x208 & n36348 ;
  assign n36350 = x200 & ~n35132 ;
  assign n36351 = n36338 & ~n36350 ;
  assign n36352 = n36349 | n36351 ;
  assign n36353 = n35272 & n36352 ;
  assign n36354 = n8652 & ~n36353 ;
  assign n36355 = ~n35197 & n35398 ;
  assign n36356 = ~n36329 & n36355 ;
  assign n36357 = x212 & ~n36356 ;
  assign n36358 = ~n36354 & n36357 ;
  assign n36359 = n36347 & n36358 ;
  assign n36360 = x219 | n36359 ;
  assign n36361 = n36346 | n36360 ;
  assign n36362 = x1151 & ~n6785 ;
  assign n36363 = ~x211 & n36352 ;
  assign n36364 = x211 & n36328 ;
  assign n36365 = n36363 | n36364 ;
  assign n36366 = n35272 & n36365 ;
  assign n36367 = n35100 | n36329 ;
  assign n36368 = n36366 & n36367 ;
  assign n36369 = x219 & ~n36368 ;
  assign n36370 = n36362 & ~n36369 ;
  assign n36371 = n36361 & n36370 ;
  assign n36372 = n35517 & ~n35614 ;
  assign n36373 = x1153 & n36372 ;
  assign n36374 = n35110 & ~n36343 ;
  assign n36375 = ~n36373 & n36374 ;
  assign n36376 = ~n8980 & n35517 ;
  assign n36377 = x299 | n36376 ;
  assign n36378 = n35508 & n36377 ;
  assign n36379 = n8894 & ~n36378 ;
  assign n36380 = x211 | n35197 ;
  assign n36381 = n36373 | n36380 ;
  assign n36382 = ( x211 & n36379 ) | ( x211 & ~n36381 ) | ( n36379 & ~n36381 ) ;
  assign n36383 = n36375 | n36382 ;
  assign n36384 = ~x219 & n36383 ;
  assign n36385 = x1151 | n6785 ;
  assign n36386 = ~n11103 & n36377 ;
  assign n36387 = x214 | n36372 ;
  assign n36388 = x212 | n36387 ;
  assign n36389 = n36386 & n36388 ;
  assign n36390 = x1153 & n36389 ;
  assign n36391 = n35474 | n36390 ;
  assign n36392 = ~n36385 & n36391 ;
  assign n36393 = ~n36384 & n36392 ;
  assign n36394 = x1152 | n36393 ;
  assign n36395 = n36371 | n36394 ;
  assign n36396 = n9579 | n35691 ;
  assign n36397 = x207 & n36396 ;
  assign n36398 = n35754 | n36397 ;
  assign n36399 = ~x208 & n36398 ;
  assign n36400 = x200 & x207 ;
  assign n36401 = x199 | n36400 ;
  assign n36402 = ~x299 & n36401 ;
  assign n36403 = x208 & ~n36402 ;
  assign n36404 = x207 | n8980 ;
  assign n36405 = ~x299 & n36404 ;
  assign n36406 = x1153 | n36405 ;
  assign n36407 = n36403 & n36406 ;
  assign n36408 = n36399 | n36407 ;
  assign n36409 = x211 & n36408 ;
  assign n36410 = ~x207 & n35628 ;
  assign n36411 = n35791 | n36410 ;
  assign n36412 = x208 & n36411 ;
  assign n36413 = n35317 & n35628 ;
  assign n36414 = n36412 | n36413 ;
  assign n36415 = x211 | n35357 ;
  assign n36416 = n36414 & ~n36415 ;
  assign n36417 = n36409 | n36416 ;
  assign n36418 = n8894 & n36417 ;
  assign n36419 = x299 & ~n35170 ;
  assign n36420 = n35110 & n36414 ;
  assign n36421 = ~n36419 & n36420 ;
  assign n36422 = n36418 | n36421 ;
  assign n36423 = ~x219 & n36422 ;
  assign n36424 = n8790 | n35626 ;
  assign n36425 = n35517 | n36149 ;
  assign n36426 = ~n9520 & n36425 ;
  assign n36427 = n36424 & n36426 ;
  assign n36428 = ~x211 & n35195 ;
  assign n36429 = n35100 & n36428 ;
  assign n36430 = n36427 | n36429 ;
  assign n36431 = ~n35474 & n36430 ;
  assign n36432 = n36423 | n36431 ;
  assign n36433 = ~n36385 & n36432 ;
  assign n36434 = n35629 | n35765 ;
  assign n36435 = x208 & n36434 ;
  assign n36436 = n35317 & ~n35655 ;
  assign n36437 = n36435 | n36436 ;
  assign n36438 = ~x211 & n36437 ;
  assign n36439 = ~n35339 & n36438 ;
  assign n36440 = x211 & n36437 ;
  assign n36441 = ~n35357 & n36440 ;
  assign n36442 = n36439 | n36441 ;
  assign n36443 = n35110 & n36442 ;
  assign n36444 = n35123 & n35215 ;
  assign n36445 = x208 & ~n35221 ;
  assign n36446 = n36404 & n36445 ;
  assign n36447 = n36444 | n36446 ;
  assign n36448 = n36378 | n36447 ;
  assign n36449 = n36416 | n36448 ;
  assign n36450 = n8894 & n36449 ;
  assign n36451 = x214 | n36447 ;
  assign n36452 = n36373 | n36451 ;
  assign n36453 = ~x212 & n36452 ;
  assign n36454 = ~x214 & n36453 ;
  assign n36455 = x219 | n36454 ;
  assign n36456 = n36450 | n36455 ;
  assign n36457 = n36443 | n36456 ;
  assign n36458 = x219 & ~n36447 ;
  assign n36459 = ~n36390 & n36458 ;
  assign n36460 = n36362 & ~n36459 ;
  assign n36461 = n36457 & n36460 ;
  assign n36462 = x1152 & ~n36461 ;
  assign n36463 = ~n36433 & n36462 ;
  assign n36464 = n36395 & ~n36463 ;
  assign n36465 = ( ~x209 & n36279 ) | ( ~x209 & n36464 ) | ( n36279 & n36464 ) ;
  assign n36466 = n36324 | n36465 ;
  assign n36467 = x213 & n36466 ;
  assign n36468 = ~n8653 & n35474 ;
  assign n36469 = n6785 & n36468 ;
  assign n36470 = ~n8894 & n36276 ;
  assign n36471 = n35409 | n36470 ;
  assign n36472 = n36469 & n36471 ;
  assign n36473 = n8654 & n35103 ;
  assign n36474 = x1151 & ~n36473 ;
  assign n36475 = ~n36472 & n36474 ;
  assign n36476 = n35898 & n36292 ;
  assign n36477 = n35895 | n36476 ;
  assign n36478 = ~x211 & n36477 ;
  assign n36479 = n36315 | n36478 ;
  assign n36480 = n35100 & ~n36479 ;
  assign n36481 = n36320 & ~n36480 ;
  assign n36482 = x219 & ~n36481 ;
  assign n36483 = n6785 | n36482 ;
  assign n36484 = x211 & n36477 ;
  assign n36485 = n36316 | n36484 ;
  assign n36486 = x214 & ~n36485 ;
  assign n36487 = ~x212 & n36319 ;
  assign n36488 = ~n36486 & n36487 ;
  assign n36489 = x219 | n36488 ;
  assign n36490 = ~x214 & n36485 ;
  assign n36491 = x214 & n36477 ;
  assign n36492 = n36490 | n36491 ;
  assign n36493 = x212 & n36492 ;
  assign n36494 = n36489 | n36493 ;
  assign n36495 = ~n36483 & n36494 ;
  assign n36496 = n36475 & ~n36495 ;
  assign n36497 = x1151 | n36472 ;
  assign n36498 = x214 & n36479 ;
  assign n36499 = n36490 | n36498 ;
  assign n36500 = x212 & n36499 ;
  assign n36501 = n36489 | n36500 ;
  assign n36502 = x219 & ~n36314 ;
  assign n36503 = n6785 | n36502 ;
  assign n36504 = n36501 & ~n36503 ;
  assign n36505 = n36497 | n36504 ;
  assign n36506 = x1152 & n36505 ;
  assign n36507 = ~n36496 & n36506 ;
  assign n36508 = ~x211 & n35442 ;
  assign n36509 = x1153 & n36508 ;
  assign n36510 = n8654 | n36509 ;
  assign n36511 = n35103 & n36510 ;
  assign n36512 = x1151 & ~n36511 ;
  assign n36513 = ~x211 & n36314 ;
  assign n36514 = n36484 | n36513 ;
  assign n36515 = ( ~x212 & x214 ) | ( ~x212 & n36514 ) | ( x214 & n36514 ) ;
  assign n36516 = ( x212 & x214 ) | ( x212 & ~n36317 ) | ( x214 & ~n36317 ) ;
  assign n36517 = ~n36515 & n36516 ;
  assign n36518 = x214 & ~n36317 ;
  assign n36519 = n36487 & ~n36518 ;
  assign n36520 = ( x212 & ~n36517 ) | ( x212 & n36519 ) | ( ~n36517 & n36519 ) ;
  assign n36521 = x219 | n36520 ;
  assign n36522 = ~n36483 & n36521 ;
  assign n36523 = n36512 & ~n36522 ;
  assign n36524 = n36061 & n36509 ;
  assign n36525 = x1151 | n36524 ;
  assign n36526 = ~x219 & n35442 ;
  assign n36527 = ( ~n6785 & n36314 ) | ( ~n6785 & n36526 ) | ( n36314 & n36526 ) ;
  assign n36528 = ( n6785 & ~n36317 ) | ( n6785 & n36526 ) | ( ~n36317 & n36526 ) ;
  assign n36529 = n36527 & ~n36528 ;
  assign n36530 = n36525 | n36529 ;
  assign n36531 = ~x1152 & n36530 ;
  assign n36532 = ~n36523 & n36531 ;
  assign n36533 = x209 & ~n36532 ;
  assign n36534 = ~n36507 & n36533 ;
  assign n36535 = ~x214 & n36366 ;
  assign n36536 = n11103 | n36373 ;
  assign n36537 = n36329 | n36536 ;
  assign n36538 = x214 & n36537 ;
  assign n36539 = x212 & ~n36538 ;
  assign n36540 = ~n36535 & n36539 ;
  assign n36541 = x212 | n36368 ;
  assign n36542 = ~n36540 & n36541 ;
  assign n36543 = x219 | n36542 ;
  assign n36544 = ~x211 & x299 ;
  assign n36545 = n36373 | n36544 ;
  assign n36546 = n36329 | n36545 ;
  assign n36547 = n36367 & n36546 ;
  assign n36548 = x219 & ~n36547 ;
  assign n36549 = n6785 | n36548 ;
  assign n36550 = n36543 & ~n36549 ;
  assign n36551 = n36512 & ~n36550 ;
  assign n36552 = ~n36387 & n36390 ;
  assign n36553 = x212 & n36387 ;
  assign n36554 = n36536 & n36553 ;
  assign n36555 = x219 | n36554 ;
  assign n36556 = n35108 & n36428 ;
  assign n36557 = n36372 | n36556 ;
  assign n36558 = n36555 | n36557 ;
  assign n36559 = n36552 | n36558 ;
  assign n36560 = x219 & ~n36372 ;
  assign n36561 = n6785 | n36560 ;
  assign n36562 = n36390 & ~n36561 ;
  assign n36563 = n36559 & n36562 ;
  assign n36564 = n36525 | n36563 ;
  assign n36565 = ~x1152 & n36564 ;
  assign n36566 = ~n36551 & n36565 ;
  assign n36567 = n36373 | n36447 ;
  assign n36568 = n36438 | n36567 ;
  assign n36569 = x214 & ~n36568 ;
  assign n36570 = n36452 & ~n36569 ;
  assign n36571 = x212 | n36570 ;
  assign n36572 = n36568 & n36571 ;
  assign n36573 = x219 & ~n36572 ;
  assign n36574 = n6785 | n36573 ;
  assign n36575 = x1153 & n36377 ;
  assign n36576 = n36440 | n36575 ;
  assign n36577 = n36451 | n36576 ;
  assign n36578 = x214 & ~n36437 ;
  assign n36579 = x212 & ~n36578 ;
  assign n36580 = n36577 & n36579 ;
  assign n36581 = x214 & ~n36447 ;
  assign n36582 = ~n36576 & n36581 ;
  assign n36583 = n36453 & ~n36582 ;
  assign n36584 = x219 | n36583 ;
  assign n36585 = n36580 | n36584 ;
  assign n36586 = ~n36574 & n36585 ;
  assign n36587 = n36475 & ~n36586 ;
  assign n36588 = x219 & ~n36427 ;
  assign n36589 = n6785 | n36588 ;
  assign n36590 = x211 | n36408 ;
  assign n36591 = n36420 & n36590 ;
  assign n36592 = ~n35442 & n36427 ;
  assign n36593 = x299 & n35409 ;
  assign n36594 = x219 | n36593 ;
  assign n36595 = n36592 | n36594 ;
  assign n36596 = n36591 | n36595 ;
  assign n36597 = ~n36589 & n36596 ;
  assign n36598 = n36497 | n36597 ;
  assign n36599 = x1152 & n36598 ;
  assign n36600 = ~n36587 & n36599 ;
  assign n36601 = n36566 | n36600 ;
  assign n36602 = x209 | n36601 ;
  assign n36603 = ~x213 & n36602 ;
  assign n36604 = ~n36534 & n36603 ;
  assign n36605 = n36467 | n36604 ;
  assign n36606 = x230 & n36605 ;
  assign n36607 = ~x230 & x238 ;
  assign n36608 = n36606 | n36607 ;
  assign n36609 = n35136 & n35248 ;
  assign n36610 = ( x212 & ~n35108 ) | ( x212 & n36609 ) | ( ~n35108 & n36609 ) ;
  assign n36611 = x219 | n36610 ;
  assign n36612 = x299 & x1158 ;
  assign n36613 = ~n35136 & n36612 ;
  assign n36614 = ~x208 & n36113 ;
  assign n36615 = n36613 | n36614 ;
  assign n36616 = ~x211 & n36615 ;
  assign n36617 = x208 & x299 ;
  assign n36618 = x1157 & ~n36617 ;
  assign n36619 = ~n35542 & n36618 ;
  assign n36620 = x1157 | n36609 ;
  assign n36621 = x211 & n36620 ;
  assign n36622 = ~n36619 & n36621 ;
  assign n36623 = n36616 | n36622 ;
  assign n36624 = x214 & n36623 ;
  assign n36625 = n36611 | n36624 ;
  assign n36626 = x219 & ~n36610 ;
  assign n36627 = x211 & ~n36609 ;
  assign n36628 = x214 & ~n36627 ;
  assign n36629 = n35585 | n35714 ;
  assign n36630 = n36628 & n36629 ;
  assign n36631 = n36626 & ~n36630 ;
  assign n36632 = x212 & ~n36609 ;
  assign n36633 = n6785 | n36632 ;
  assign n36634 = x209 | n36633 ;
  assign n36635 = n36631 | n36634 ;
  assign n36636 = n36625 & ~n36635 ;
  assign n36637 = n36139 & n36188 ;
  assign n36638 = ( x212 & ~n35108 ) | ( x212 & n36637 ) | ( ~n35108 & n36637 ) ;
  assign n36639 = x219 | n36638 ;
  assign n36640 = x208 & ~n36612 ;
  assign n36641 = n35388 | n36640 ;
  assign n36642 = n36125 & ~n36641 ;
  assign n36643 = n36134 | n36642 ;
  assign n36644 = ~n36103 & n36618 ;
  assign n36645 = n36188 & ~n36644 ;
  assign n36646 = x211 & ~n36645 ;
  assign n36647 = x214 & ~n36646 ;
  assign n36648 = n36643 & n36647 ;
  assign n36649 = n36639 | n36648 ;
  assign n36650 = x219 & ~n36638 ;
  assign n36651 = x211 & ~n36637 ;
  assign n36652 = n35714 | n36637 ;
  assign n36653 = x214 & n36652 ;
  assign n36654 = ~n36651 & n36653 ;
  assign n36655 = n36650 & ~n36654 ;
  assign n36656 = x212 & ~n36637 ;
  assign n36657 = n6785 | n36656 ;
  assign n36658 = x209 & ~n36657 ;
  assign n36659 = ~n36655 & n36658 ;
  assign n36660 = n36649 & n36659 ;
  assign n36661 = x219 | n36059 ;
  assign n36662 = n36064 & n36661 ;
  assign n36663 = x213 & ~n36662 ;
  assign n36664 = ~n36660 & n36663 ;
  assign n36665 = ~n36636 & n36664 ;
  assign n36666 = n36235 | n36380 ;
  assign n36667 = x214 & ~n36651 ;
  assign n36668 = n36666 & n36667 ;
  assign n36669 = n36650 & ~n36668 ;
  assign n36670 = x211 & ~n35193 ;
  assign n36671 = ~n36235 & n36670 ;
  assign n36672 = n36653 & ~n36671 ;
  assign n36673 = n36639 | n36672 ;
  assign n36674 = ~n36657 & n36673 ;
  assign n36675 = ~n36669 & n36674 ;
  assign n36676 = n6785 & ~n35817 ;
  assign n36677 = n35108 & n35815 ;
  assign n36678 = n36676 & n36677 ;
  assign n36679 = x213 | n36678 ;
  assign n36680 = ( x209 & n36675 ) | ( x209 & n36679 ) | ( n36675 & n36679 ) ;
  assign n36681 = n35197 | n35530 ;
  assign n36682 = n36628 & n36681 ;
  assign n36683 = n36626 & ~n36682 ;
  assign n36684 = ~n35591 & n36670 ;
  assign n36685 = x214 & ~n36684 ;
  assign n36686 = n36629 & n36685 ;
  assign n36687 = n36611 | n36686 ;
  assign n36688 = ~n36633 & n36687 ;
  assign n36689 = ~n36683 & n36688 ;
  assign n36690 = ( ~x209 & n36679 ) | ( ~x209 & n36689 ) | ( n36679 & n36689 ) ;
  assign n36691 = n36680 | n36690 ;
  assign n36692 = ~n36665 & n36691 ;
  assign n36693 = x230 & ~n36692 ;
  assign n36694 = x230 | x239 ;
  assign n36695 = ~n36693 & n36694 ;
  assign n36696 = ~n6785 & n36426 ;
  assign n36697 = n36561 & ~n36696 ;
  assign n36698 = x214 | n36426 ;
  assign n36699 = ~x212 & n36698 ;
  assign n36700 = ~n9520 & n35136 ;
  assign n36701 = x299 | n36700 ;
  assign n36702 = n36403 | n36701 ;
  assign n36703 = x214 & ~n36702 ;
  assign n36704 = n36699 & ~n36703 ;
  assign n36705 = x219 | n36704 ;
  assign n36706 = ~x211 & n36702 ;
  assign n36707 = x211 & n36426 ;
  assign n36708 = x214 & ~n36707 ;
  assign n36709 = ~n36706 & n36708 ;
  assign n36710 = x212 & ~n36709 ;
  assign n36711 = n36702 & n36710 ;
  assign n36712 = n36705 | n36711 ;
  assign n36713 = ~n36697 & n36712 ;
  assign n36714 = n36469 | n36713 ;
  assign n36715 = ( x1147 & x1149 ) | ( x1147 & n36714 ) | ( x1149 & n36714 ) ;
  assign n36716 = ~x211 & n6785 ;
  assign n36717 = n36061 | n36716 ;
  assign n36718 = n35100 & n36717 ;
  assign n36719 = x299 & n35100 ;
  assign n36720 = n6785 | n35102 ;
  assign n36721 = n36719 & ~n36720 ;
  assign n36722 = ~n35221 & n35516 ;
  assign n36723 = ~n6785 & n36722 ;
  assign n36724 = n36721 | n36723 ;
  assign n36725 = n36718 | n36724 ;
  assign n36726 = ( ~x1147 & x1149 ) | ( ~x1147 & n36725 ) | ( x1149 & n36725 ) ;
  assign n36727 = n36715 & n36726 ;
  assign n36728 = x211 & n35108 ;
  assign n36729 = x219 | n36728 ;
  assign n36730 = n35366 | n36729 ;
  assign n36731 = n36721 & n36730 ;
  assign n36732 = ~n6785 & n36447 ;
  assign n36733 = n35103 & n36730 ;
  assign n36734 = n36732 | n36733 ;
  assign n36735 = n36731 | n36734 ;
  assign n36736 = ( x1147 & x1149 ) | ( x1147 & ~n36735 ) | ( x1149 & ~n36735 ) ;
  assign n36737 = x212 & n35398 ;
  assign n36738 = n36728 | n36737 ;
  assign n36739 = n36061 & n36738 ;
  assign n36740 = n35517 | n35791 ;
  assign n36741 = n8790 | n35320 ;
  assign n36742 = n36740 & n36741 ;
  assign n36743 = n36405 & n36742 ;
  assign n36744 = x299 & n8652 ;
  assign n36745 = n36743 | n36744 ;
  assign n36746 = ~x212 & n36745 ;
  assign n36747 = x219 | n36746 ;
  assign n36748 = x299 | n36742 ;
  assign n36749 = x214 & n36748 ;
  assign n36750 = n11103 | n36743 ;
  assign n36751 = n36749 | n36750 ;
  assign n36752 = x212 & n36751 ;
  assign n36753 = ( x212 & ~n35108 ) | ( x212 & n36743 ) | ( ~n35108 & n36743 ) ;
  assign n36754 = ~x211 & n36748 ;
  assign n36755 = n36743 | n36754 ;
  assign n36756 = x214 & n36755 ;
  assign n36757 = x212 & ~n36756 ;
  assign n36758 = ( x214 & ~n36748 ) | ( x214 & n36757 ) | ( ~n36748 & n36757 ) ;
  assign n36759 = x214 & ~n36757 ;
  assign n36760 = ( n36753 & ~n36758 ) | ( n36753 & n36759 ) | ( ~n36758 & n36759 ) ;
  assign n36761 = n36752 & n36760 ;
  assign n36762 = n36747 | n36761 ;
  assign n36763 = x219 & ~n36743 ;
  assign n36764 = n6785 | n36763 ;
  assign n36765 = n36762 & ~n36764 ;
  assign n36766 = n36739 | n36765 ;
  assign n36767 = ( x1147 & ~x1149 ) | ( x1147 & n36766 ) | ( ~x1149 & n36766 ) ;
  assign n36768 = ~n36736 & n36767 ;
  assign n36769 = n36727 | n36768 ;
  assign n36770 = x1148 & n36769 ;
  assign n36771 = x212 | n36744 ;
  assign n36772 = n36447 | n36771 ;
  assign n36773 = n36447 | n36544 ;
  assign n36774 = n36451 & n36773 ;
  assign n36775 = ( x212 & n8894 ) | ( x212 & ~n11103 ) | ( n8894 & ~n11103 ) ;
  assign n36776 = ~n36774 & n36775 ;
  assign n36777 = n36772 & ~n36776 ;
  assign n36778 = x219 | n36777 ;
  assign n36779 = n35291 | n36400 ;
  assign n36780 = x208 & n36779 ;
  assign n36781 = x199 | n36780 ;
  assign n36782 = n36447 & n36781 ;
  assign n36783 = x299 | n36782 ;
  assign n36784 = x219 | n36783 ;
  assign n36785 = n36778 & n36784 ;
  assign n36786 = x211 | n36785 ;
  assign n36787 = ~n11103 & n36581 ;
  assign n36788 = ( x212 & n8894 ) | ( x212 & n36773 ) | ( n8894 & n36773 ) ;
  assign n36789 = ~n36787 & n36788 ;
  assign n36790 = ~x212 & n36774 ;
  assign n36791 = x219 | n36790 ;
  assign n36792 = n36789 | n36791 ;
  assign n36793 = x219 & ~n36544 ;
  assign n36794 = n36720 | n36793 ;
  assign n36795 = ~n36732 & n36794 ;
  assign n36796 = n36792 & ~n36795 ;
  assign n36797 = n36783 & n36796 ;
  assign n36798 = n36786 & n36797 ;
  assign n36799 = n36473 | n36798 ;
  assign n36800 = x1147 & ~x1149 ;
  assign n36801 = n36799 & n36800 ;
  assign n36802 = ~n14313 & n36376 ;
  assign n36803 = ~x219 & n14313 ;
  assign n36804 = n36508 & n36803 ;
  assign n36805 = n36802 | n36804 ;
  assign n36806 = ( x1147 & x1149 ) | ( x1147 & n36805 ) | ( x1149 & n36805 ) ;
  assign n36807 = n8654 | n36508 ;
  assign n36808 = n35103 & n36807 ;
  assign n36809 = ~x211 & n36328 ;
  assign n36810 = x211 & n36352 ;
  assign n36811 = x214 & ~n36810 ;
  assign n36812 = ~n36809 & n36811 ;
  assign n36813 = n8894 & ~n36812 ;
  assign n36814 = x214 | n36328 ;
  assign n36815 = ~x212 & n36814 ;
  assign n36816 = x214 & ~n36365 ;
  assign n36817 = n36815 & ~n36816 ;
  assign n36818 = x219 | n36817 ;
  assign n36819 = x212 & ~n36812 ;
  assign n36820 = n36365 & n36819 ;
  assign n36821 = n36818 | n36820 ;
  assign n36822 = n36813 | n36821 ;
  assign n36823 = x212 & n36365 ;
  assign n36824 = x219 & ~n36823 ;
  assign n36825 = ~n36817 & n36824 ;
  assign n36826 = n6785 | n36825 ;
  assign n36827 = n36822 & ~n36826 ;
  assign n36828 = n36808 | n36827 ;
  assign n36829 = ( ~x1147 & x1149 ) | ( ~x1147 & n36828 ) | ( x1149 & n36828 ) ;
  assign n36830 = n36806 & n36829 ;
  assign n36831 = n36801 | n36830 ;
  assign n36832 = ~x1148 & n36831 ;
  assign n36833 = n36770 | n36832 ;
  assign n36834 = x213 & n36833 ;
  assign n36835 = ~x211 & x1146 ;
  assign n36836 = x211 & x1145 ;
  assign n36837 = n36835 | n36836 ;
  assign n36838 = x214 & n36837 ;
  assign n36839 = x211 & x1146 ;
  assign n36840 = ~x214 & n36839 ;
  assign n36841 = n36838 | n36840 ;
  assign n36842 = x212 & n36841 ;
  assign n36843 = n35108 & n36839 ;
  assign n36844 = n36842 | n36843 ;
  assign n36845 = n35734 | n36844 ;
  assign n36846 = n6785 & n36026 ;
  assign n36847 = n36061 | n36846 ;
  assign n36848 = n36845 & n36847 ;
  assign n36849 = ~n8897 & n35474 ;
  assign n36850 = n6785 & n36849 ;
  assign n36851 = x1147 & ~n36850 ;
  assign n36852 = ~n36848 & n36851 ;
  assign n36853 = ~x211 & n36208 ;
  assign n36854 = x219 & ~n36853 ;
  assign n36855 = n36720 | n36854 ;
  assign n36856 = x219 & ~n36328 ;
  assign n36857 = n6785 | n36856 ;
  assign n36858 = n36855 & n36857 ;
  assign n36859 = x299 & x1146 ;
  assign n36860 = ~x299 & n36351 ;
  assign n36861 = n36086 | n36860 ;
  assign n36862 = n36859 | n36861 ;
  assign n36863 = x211 & n36862 ;
  assign n36864 = n36363 | n36863 ;
  assign n36865 = x214 | n36864 ;
  assign n36866 = x299 & n36837 ;
  assign n36867 = x214 & ~n36866 ;
  assign n36868 = ~n36861 & n36867 ;
  assign n36869 = x212 & ~n36868 ;
  assign n36870 = n36865 & n36869 ;
  assign n36871 = x214 & ~n36864 ;
  assign n36872 = n36815 & ~n36871 ;
  assign n36873 = x219 | n36872 ;
  assign n36874 = n36870 | n36873 ;
  assign n36875 = ~n36858 & n36874 ;
  assign n36876 = n36852 & ~n36875 ;
  assign n36877 = x1147 | n36848 ;
  assign n36878 = x219 & ~n36855 ;
  assign n36879 = x299 & n36844 ;
  assign n36880 = ~n32969 & n36879 ;
  assign n36881 = n36878 | n36880 ;
  assign n36882 = n36877 | n36881 ;
  assign n36883 = n36802 | n36882 ;
  assign n36884 = ~x1148 & n36883 ;
  assign n36885 = ~n36876 & n36884 ;
  assign n36886 = n35100 & n36706 ;
  assign n36887 = ~n35101 & n36426 ;
  assign n36888 = x219 & ~n36887 ;
  assign n36889 = ~n36886 & n36888 ;
  assign n36890 = n6785 | n36889 ;
  assign n36891 = n9520 | n36890 ;
  assign n36892 = n36855 & n36891 ;
  assign n36893 = x212 & n36702 ;
  assign n36894 = n36426 | n36841 ;
  assign n36895 = n36893 & n36894 ;
  assign n36896 = x211 & n36859 ;
  assign n36897 = n36426 | n36896 ;
  assign n36898 = n36699 & n36897 ;
  assign n36899 = x219 | n36898 ;
  assign n36900 = n36895 | n36899 ;
  assign n36901 = ~n36892 & n36900 ;
  assign n36902 = n36877 | n36901 ;
  assign n36903 = x219 & ~n36722 ;
  assign n36904 = n6785 | n36903 ;
  assign n36905 = x299 & n35366 ;
  assign n36906 = ( x212 & x299 ) | ( x212 & n36722 ) | ( x299 & n36722 ) ;
  assign n36907 = ~n36905 & n36906 ;
  assign n36908 = x211 & ~n36722 ;
  assign n36909 = x214 & x299 ;
  assign n36910 = n36722 | n36909 ;
  assign n36911 = ~x212 & n36910 ;
  assign n36912 = ~n36908 & n36911 ;
  assign n36913 = x219 | n36912 ;
  assign n36914 = n36907 | n36913 ;
  assign n36915 = ~n36904 & n36914 ;
  assign n36916 = n36852 & ~n36881 ;
  assign n36917 = ~n36915 & n36916 ;
  assign n36918 = x1148 & ~n36917 ;
  assign n36919 = n36902 & n36918 ;
  assign n36920 = n36885 | n36919 ;
  assign n36921 = ( x213 & x1149 ) | ( x213 & ~n36920 ) | ( x1149 & ~n36920 ) ;
  assign n36922 = ~n6785 & n36743 ;
  assign n36923 = n36882 | n36922 ;
  assign n36924 = ~n36732 & n36855 ;
  assign n36925 = n36544 | n36896 ;
  assign n36926 = n36447 | n36925 ;
  assign n36927 = n35442 & n36926 ;
  assign n36928 = ~n35100 & n36447 ;
  assign n36929 = x219 | n36928 ;
  assign n36930 = n36447 | n36866 ;
  assign n36931 = n8894 & n36930 ;
  assign n36932 = n36929 | n36931 ;
  assign n36933 = n36927 | n36932 ;
  assign n36934 = ~n36924 & n36933 ;
  assign n36935 = n36852 & ~n36934 ;
  assign n36936 = x1148 & ~n36935 ;
  assign n36937 = n36923 & n36936 ;
  assign n36938 = ~x1146 & n11103 ;
  assign n36939 = n35442 & ~n36938 ;
  assign n36940 = n36931 | n36939 ;
  assign n36941 = ~x219 & n36783 ;
  assign n36942 = n36940 & n36941 ;
  assign n36943 = n36026 & n36049 ;
  assign n36944 = ~n35474 & n36782 ;
  assign n36945 = n36943 | n36944 ;
  assign n36946 = n36942 | n36945 ;
  assign n36947 = ~n6785 & n36946 ;
  assign n36948 = n36852 & ~n36947 ;
  assign n36949 = ~x1148 & n36882 ;
  assign n36950 = ~n36948 & n36949 ;
  assign n36951 = n36937 | n36950 ;
  assign n36952 = ( ~x213 & x1149 ) | ( ~x213 & n36951 ) | ( x1149 & n36951 ) ;
  assign n36953 = ~n36921 & n36952 ;
  assign n36954 = x209 & ~n36953 ;
  assign n36955 = ~n36834 & n36954 ;
  assign n36956 = ~x199 & x1146 ;
  assign n36957 = x200 & ~n36956 ;
  assign n36958 = x299 | n36957 ;
  assign n36959 = x199 & x1145 ;
  assign n36960 = n35290 & ~n36959 ;
  assign n36961 = n36958 | n36960 ;
  assign n36962 = x207 | n36961 ;
  assign n36963 = x200 | n36959 ;
  assign n36964 = n36956 | n36963 ;
  assign n36965 = x200 & ~n36042 ;
  assign n36966 = n35123 & ~n36965 ;
  assign n36967 = n36964 & n36966 ;
  assign n36968 = n36859 | n36967 ;
  assign n36969 = n36962 & ~n36968 ;
  assign n36970 = x208 & ~n36969 ;
  assign n36971 = n35136 & ~n36961 ;
  assign n36972 = n36970 | n36971 ;
  assign n36973 = x299 | n36972 ;
  assign n36974 = x211 & n36973 ;
  assign n36975 = n36962 | n36963 ;
  assign n36976 = n36970 & n36975 ;
  assign n36977 = ~n36958 & n36963 ;
  assign n36978 = n35136 & n36977 ;
  assign n36979 = n36976 | n36978 ;
  assign n36980 = x299 | n36979 ;
  assign n36981 = x214 & n36980 ;
  assign n36982 = n36974 | n36981 ;
  assign n36983 = x212 & n36982 ;
  assign n36984 = n8652 & n36973 ;
  assign n36985 = n35517 | n36967 ;
  assign n36986 = ~n8790 & n36961 ;
  assign n36987 = n36985 & ~n36986 ;
  assign n36988 = x219 | n36987 ;
  assign n36989 = n36984 | n36988 ;
  assign n36990 = n36983 | n36989 ;
  assign n36991 = n8790 | n36977 ;
  assign n36992 = n36985 & n36991 ;
  assign n36993 = ~n35100 & n36992 ;
  assign n36994 = n36990 | n36993 ;
  assign n36995 = ( x219 & n6785 ) | ( x219 & ~n36992 ) | ( n6785 & ~n36992 ) ;
  assign n36996 = ~x211 & n36973 ;
  assign n36997 = n36987 | n36996 ;
  assign n36998 = x214 & ~n36997 ;
  assign n36999 = n36980 & ~n36998 ;
  assign n37000 = x212 & ~n36999 ;
  assign n37001 = ( x212 & ~n35108 ) | ( x212 & n36992 ) | ( ~n35108 & n36992 ) ;
  assign n37002 = n36981 | n37001 ;
  assign n37003 = ~n37000 & n37002 ;
  assign n37004 = ( x219 & ~n6785 ) | ( x219 & n37003 ) | ( ~n6785 & n37003 ) ;
  assign n37005 = ~n36995 & n37004 ;
  assign n37006 = n36994 & n37005 ;
  assign n37007 = x1147 | n36739 ;
  assign n37008 = n37006 | n37007 ;
  assign n37009 = ~n35101 & n36987 ;
  assign n37010 = x219 & ~n37009 ;
  assign n37011 = n35100 & n36996 ;
  assign n37012 = n37010 & ~n37011 ;
  assign n37013 = n6785 | n37012 ;
  assign n37014 = n36990 & ~n37013 ;
  assign n37015 = x1147 & ~n36733 ;
  assign n37016 = ~n37014 & n37015 ;
  assign n37017 = x1149 | n37016 ;
  assign n37018 = n37008 & ~n37017 ;
  assign n37019 = x1147 | n36469 ;
  assign n37020 = n37005 | n37019 ;
  assign n37021 = n36719 | n36988 ;
  assign n37022 = ~n37013 & n37021 ;
  assign n37023 = x1147 & ~n36718 ;
  assign n37024 = ~n37022 & n37023 ;
  assign n37025 = x1149 & ~n37024 ;
  assign n37026 = n37020 & n37025 ;
  assign n37027 = x1148 & ~n37026 ;
  assign n37028 = ~n37018 & n37027 ;
  assign n37029 = x213 & ~n37028 ;
  assign n37030 = x214 | n36987 ;
  assign n37031 = n36996 | n37030 ;
  assign n37032 = n36974 | n36987 ;
  assign n37033 = ( x212 & n35109 ) | ( x212 & n37032 ) | ( n35109 & n37032 ) ;
  assign n37034 = n37031 & n37033 ;
  assign n37035 = ~x212 & n37030 ;
  assign n37036 = n36997 & n37035 ;
  assign n37037 = x219 | n37036 ;
  assign n37038 = n37034 | n37037 ;
  assign n37039 = ~n37013 & n37038 ;
  assign n37040 = n36808 | n37039 ;
  assign n37041 = x1147 & n37040 ;
  assign n37042 = x1147 | n6785 ;
  assign n37043 = n36992 & ~n37042 ;
  assign n37044 = ~x1147 & n36849 ;
  assign n37045 = n37043 | n37044 ;
  assign n37046 = ~n14313 & n36849 ;
  assign n37047 = ~n36979 & n37046 ;
  assign n37048 = n37045 & ~n37047 ;
  assign n37049 = n37041 | n37048 ;
  assign n37050 = ( x1148 & x1149 ) | ( x1148 & n37049 ) | ( x1149 & n37049 ) ;
  assign n37051 = n37014 & n37038 ;
  assign n37052 = n36473 | n37051 ;
  assign n37053 = x1147 & n37052 ;
  assign n37054 = n37043 | n37053 ;
  assign n37055 = ( x1148 & ~x1149 ) | ( x1148 & n37054 ) | ( ~x1149 & n37054 ) ;
  assign n37056 = n37050 | n37055 ;
  assign n37057 = n37029 & n37056 ;
  assign n37058 = n36896 | n36992 ;
  assign n37059 = x214 | n36992 ;
  assign n37060 = ~x212 & n37059 ;
  assign n37061 = n37058 & n37060 ;
  assign n37062 = x219 | n37061 ;
  assign n37063 = ~x299 & n36979 ;
  assign n37064 = n36867 & ~n37063 ;
  assign n37065 = ( x212 & n8894 ) | ( x212 & n37058 ) | ( n8894 & n37058 ) ;
  assign n37066 = ~n37064 & n37065 ;
  assign n37067 = n37062 | n37066 ;
  assign n37068 = x219 & ~n36993 ;
  assign n37069 = x211 | n36208 ;
  assign n37070 = n37063 | n37069 ;
  assign n37071 = ( n35100 & n35101 ) | ( n35100 & n36992 ) | ( n35101 & n36992 ) ;
  assign n37072 = n37070 & n37071 ;
  assign n37073 = n37068 & ~n37072 ;
  assign n37074 = n6785 | n37073 ;
  assign n37075 = n37067 & ~n37074 ;
  assign n37076 = n36877 | n37075 ;
  assign n37077 = ~n36205 & n36974 ;
  assign n37078 = n36867 & ~n36972 ;
  assign n37079 = n36984 | n37078 ;
  assign n37080 = ~n37077 & n37079 ;
  assign n37081 = n36925 | n36972 ;
  assign n37082 = ( x212 & n8894 ) | ( x212 & n37081 ) | ( n8894 & n37081 ) ;
  assign n37083 = ~n37080 & n37082 ;
  assign n37084 = n37036 | n37062 ;
  assign n37085 = n37083 | n37084 ;
  assign n37086 = ~n36205 & n36996 ;
  assign n37087 = n35100 & n37086 ;
  assign n37088 = n37010 & ~n37087 ;
  assign n37089 = n6785 | n37088 ;
  assign n37090 = n37085 & ~n37089 ;
  assign n37091 = n36852 & ~n37090 ;
  assign n37092 = n37076 & ~n37091 ;
  assign n37093 = ~x213 & n37092 ;
  assign n37094 = x209 | n37093 ;
  assign n37095 = n37057 | n37094 ;
  assign n37096 = ~n36955 & n37095 ;
  assign n37097 = x230 & ~n37096 ;
  assign n37098 = x230 | x240 ;
  assign n37099 = ~n37097 & n37098 ;
  assign n37100 = x213 & n36601 ;
  assign n37101 = x209 & ~n37100 ;
  assign n37102 = ~n35398 & n36437 ;
  assign n37103 = x212 & ~n36567 ;
  assign n37104 = ~n37102 & n37103 ;
  assign n37105 = n36571 & ~n37104 ;
  assign n37106 = x219 | n37105 ;
  assign n37107 = x1152 & n37106 ;
  assign n37108 = ~n36574 & n37107 ;
  assign n37109 = x1151 & ~n36808 ;
  assign n37110 = ~x214 & n36546 ;
  assign n37111 = n36539 & ~n37110 ;
  assign n37112 = x212 | n36547 ;
  assign n37113 = ~n37111 & n37112 ;
  assign n37114 = x219 | n37113 ;
  assign n37115 = x1152 | n36549 ;
  assign n37116 = n37114 & ~n37115 ;
  assign n37117 = n37109 & ~n37116 ;
  assign n37118 = ~n37108 & n37117 ;
  assign n37119 = n36427 | n36555 ;
  assign n37120 = x219 & ~n36373 ;
  assign n37121 = n6785 | n37120 ;
  assign n37122 = n36794 & n37121 ;
  assign n37123 = n36589 & n37122 ;
  assign n37124 = x1152 & ~n37123 ;
  assign n37125 = n37119 & n37124 ;
  assign n37126 = x1151 | n36473 ;
  assign n37127 = n36373 | n36555 ;
  assign n37128 = ~n37122 & n37127 ;
  assign n37129 = ~x1152 & n37128 ;
  assign n37130 = n37126 | n37129 ;
  assign n37131 = n37125 | n37130 ;
  assign n37132 = ~x1150 & n37131 ;
  assign n37133 = ~n37118 & n37132 ;
  assign n37134 = n36453 & ~n36578 ;
  assign n37135 = x219 | n37134 ;
  assign n37136 = x212 & n36437 ;
  assign n37137 = n37135 | n37136 ;
  assign n37138 = x1152 & n37137 ;
  assign n37139 = ~n36574 & n37138 ;
  assign n37140 = x1151 & ~n36718 ;
  assign n37141 = x299 | n36353 ;
  assign n37142 = n36367 & n37141 ;
  assign n37143 = x219 | n37142 ;
  assign n37144 = ~n37115 & n37143 ;
  assign n37145 = n37140 & ~n37144 ;
  assign n37146 = ~n37139 & n37145 ;
  assign n37147 = x1151 | n36733 ;
  assign n37148 = ~x212 & n36377 ;
  assign n37149 = n36387 & n37148 ;
  assign n37150 = ~n36544 & n37149 ;
  assign n37151 = x219 | n37150 ;
  assign n37152 = x214 & ~n36386 ;
  assign n37153 = x211 | n36387 ;
  assign n37154 = x212 & n36377 ;
  assign n37155 = n37153 & n37154 ;
  assign n37156 = ~n37152 & n37155 ;
  assign n37157 = n37151 | n37156 ;
  assign n37158 = x299 | n37127 ;
  assign n37159 = n37157 & n37158 ;
  assign n37160 = ~n37121 & n37159 ;
  assign n37161 = x1152 | n37160 ;
  assign n37162 = n37128 | n37161 ;
  assign n37163 = n8894 & ~n36414 ;
  assign n37164 = n36388 & n36536 ;
  assign n37165 = n8894 | n36427 ;
  assign n37166 = n37164 | n37165 ;
  assign n37167 = ~n37163 & n37166 ;
  assign n37168 = x219 | n37167 ;
  assign n37169 = n37124 & n37168 ;
  assign n37170 = ( ~x1152 & n37162 ) | ( ~x1152 & n37169 ) | ( n37162 & n37169 ) ;
  assign n37171 = n37147 | n37170 ;
  assign n37172 = x1150 & n37171 ;
  assign n37173 = ~n37146 & n37172 ;
  assign n37174 = n37133 | n37173 ;
  assign n37175 = ( x213 & x1149 ) | ( x213 & ~n37174 ) | ( x1149 & ~n37174 ) ;
  assign n37176 = n6785 & ~n36849 ;
  assign n37177 = x1151 & ~n37176 ;
  assign n37178 = n36437 & n36849 ;
  assign n37179 = n36567 | n37178 ;
  assign n37180 = x1152 & n37179 ;
  assign n37181 = n6785 | n37180 ;
  assign n37182 = n37177 & n37181 ;
  assign n37183 = n36373 & ~n36385 ;
  assign n37184 = n35191 & n36508 ;
  assign n37185 = n36329 | n37184 ;
  assign n37186 = n37177 & n37185 ;
  assign n37187 = n37183 | n37186 ;
  assign n37188 = ~x1152 & n37187 ;
  assign n37189 = x1152 & ~n36385 ;
  assign n37190 = n36427 & n37189 ;
  assign n37191 = n37188 | n37190 ;
  assign n37192 = n37182 | n37191 ;
  assign n37193 = ~x1150 & n37192 ;
  assign n37194 = x1151 & ~n36469 ;
  assign n37195 = ~n36732 & n37121 ;
  assign n37196 = ( x212 & n8894 ) | ( x212 & n36437 ) | ( n8894 & n36437 ) ;
  assign n37197 = ~n36569 & n37196 ;
  assign n37198 = n37135 | n37197 ;
  assign n37199 = x1152 & n37198 ;
  assign n37200 = ( x212 & n8894 ) | ( x212 & n36352 ) | ( n8894 & n36352 ) ;
  assign n37201 = ~n36816 & n37200 ;
  assign n37202 = n36331 | n37201 ;
  assign n37203 = n37141 & n37202 ;
  assign n37204 = x219 | n37203 ;
  assign n37205 = x1152 | n36856 ;
  assign n37206 = n37204 & ~n37205 ;
  assign n37207 = n37199 | n37206 ;
  assign n37208 = ~n37195 & n37207 ;
  assign n37209 = n37194 & ~n37208 ;
  assign n37210 = x1151 | n36739 ;
  assign n37211 = n36427 | n37159 ;
  assign n37212 = ~n36589 & n37211 ;
  assign n37213 = x1152 & ~n37212 ;
  assign n37214 = n37161 & ~n37213 ;
  assign n37215 = n37210 | n37214 ;
  assign n37216 = x1150 & n37215 ;
  assign n37217 = ~n37209 & n37216 ;
  assign n37218 = n37193 | n37217 ;
  assign n37219 = ( ~x213 & x1149 ) | ( ~x213 & n37218 ) | ( x1149 & n37218 ) ;
  assign n37220 = ~n37175 & n37219 ;
  assign n37221 = n37101 & ~n37220 ;
  assign n37222 = n36815 | n36819 ;
  assign n37223 = ~n35327 & n36363 ;
  assign n37224 = n36364 | n37223 ;
  assign n37225 = n36813 | n37224 ;
  assign n37226 = n37222 & n37225 ;
  assign n37227 = x219 | n37226 ;
  assign n37228 = ~n36826 & n37227 ;
  assign n37229 = n36512 & ~n37228 ;
  assign n37230 = x299 & ~n36276 ;
  assign n37231 = n36782 | n37184 ;
  assign n37232 = ~n6785 & n37231 ;
  assign n37233 = ~n37230 & n37232 ;
  assign n37234 = n36525 | n37233 ;
  assign n37235 = ~x1152 & n37234 ;
  assign n37236 = ~n37229 & n37235 ;
  assign n37237 = ~n36812 & n36814 ;
  assign n37238 = x219 | n36905 ;
  assign n37239 = n36368 | n37238 ;
  assign n37240 = n37237 | n37239 ;
  assign n37241 = ~n36826 & n37240 ;
  assign n37242 = n36475 & ~n37241 ;
  assign n37243 = n36719 | n36782 ;
  assign n37244 = n35216 | n36471 ;
  assign n37245 = n37243 & n37244 ;
  assign n37246 = x219 | n37245 ;
  assign n37247 = x219 & ~n36782 ;
  assign n37248 = n6785 | n37247 ;
  assign n37249 = n37246 & ~n37248 ;
  assign n37250 = n36497 | n37249 ;
  assign n37251 = x1152 & n37250 ;
  assign n37252 = ~n37242 & n37251 ;
  assign n37253 = x1150 | n37252 ;
  assign n37254 = n37236 | n37253 ;
  assign n37255 = x1149 & ~x1150 ;
  assign n37256 = x219 | n36722 ;
  assign n37257 = n36905 | n37256 ;
  assign n37258 = x1153 | n37257 ;
  assign n37259 = x299 & n8653 ;
  assign n37260 = x219 | n37259 ;
  assign n37261 = ~n36794 & n37260 ;
  assign n37262 = n36915 | n37261 ;
  assign n37263 = n37258 & n37262 ;
  assign n37264 = x211 | n37257 ;
  assign n37265 = n36724 & n37264 ;
  assign n37266 = n36475 & ~n37265 ;
  assign n37267 = ~n37263 & n37266 ;
  assign n37268 = n6785 | n36458 ;
  assign n37269 = x299 | n36447 ;
  assign n37270 = n35110 & ~n37230 ;
  assign n37271 = n37269 & n37270 ;
  assign n37272 = n8894 & n36773 ;
  assign n37273 = n36929 | n37272 ;
  assign n37274 = n37271 | n37273 ;
  assign n37275 = ~n37268 & n37274 ;
  assign n37276 = n36497 | n37275 ;
  assign n37277 = x1152 & n37276 ;
  assign n37278 = ~n37267 & n37277 ;
  assign n37279 = n36512 & ~n37263 ;
  assign n37280 = x1153 & n37184 ;
  assign n37281 = n36525 | n37280 ;
  assign n37282 = ~x1152 & n37281 ;
  assign n37283 = x1151 | n36732 ;
  assign n37284 = ~x1152 & n37283 ;
  assign n37285 = n37282 | n37284 ;
  assign n37286 = ~n37279 & n37285 ;
  assign n37287 = n37278 | n37286 ;
  assign n37288 = ( x1149 & n37255 ) | ( x1149 & n37287 ) | ( n37255 & n37287 ) ;
  assign n37289 = n37254 & n37288 ;
  assign n37290 = n36748 & ~n37230 ;
  assign n37291 = ( x214 & n36757 ) | ( x214 & ~n37290 ) | ( n36757 & ~n37290 ) ;
  assign n37292 = ( n36753 & n36759 ) | ( n36753 & ~n37291 ) | ( n36759 & ~n37291 ) ;
  assign n37293 = x219 | n37292 ;
  assign n37294 = ~n36764 & n37293 ;
  assign n37295 = n36497 | n37294 ;
  assign n37296 = x211 & n36702 ;
  assign n37297 = ~n9515 & n35317 ;
  assign n37298 = n36403 | n37297 ;
  assign n37299 = x211 | n35327 ;
  assign n37300 = n37298 & ~n37299 ;
  assign n37301 = n37296 | n37300 ;
  assign n37302 = x214 | n37301 ;
  assign n37303 = n36893 & n37302 ;
  assign n37304 = x214 & ~n37301 ;
  assign n37305 = n36699 & ~n37304 ;
  assign n37306 = x219 | n37305 ;
  assign n37307 = n37303 | n37306 ;
  assign n37308 = ~n36890 & n37307 ;
  assign n37309 = n36475 & ~n37308 ;
  assign n37310 = x1152 & ~n37309 ;
  assign n37311 = n37295 & n37310 ;
  assign n37312 = n36426 | n37296 ;
  assign n37313 = x214 & ~n37312 ;
  assign n37314 = n36698 | n36706 ;
  assign n37315 = x212 & n37314 ;
  assign n37316 = ~n37313 & n37315 ;
  assign n37317 = n37301 & n37316 ;
  assign n37318 = n36707 | n37300 ;
  assign n37319 = n36699 & n37318 ;
  assign n37320 = x219 | n37319 ;
  assign n37321 = n37317 | n37320 ;
  assign n37322 = ~n36890 & n37321 ;
  assign n37323 = n36512 & ~n37322 ;
  assign n37324 = ~n36526 & n36743 ;
  assign n37325 = ~n35327 & n36748 ;
  assign n37326 = x211 | n37325 ;
  assign n37327 = n36526 & n36755 ;
  assign n37328 = n37326 & n37327 ;
  assign n37329 = n37324 | n37328 ;
  assign n37330 = ~n6785 & n37329 ;
  assign n37331 = n36525 | n37330 ;
  assign n37332 = ~x1152 & n37331 ;
  assign n37333 = ~n37323 & n37332 ;
  assign n37334 = x1150 & ~n37333 ;
  assign n37335 = ~n37311 & n37334 ;
  assign n37336 = ~x1149 & x1150 ;
  assign n37337 = x219 & ~n36389 ;
  assign n37338 = n6785 | n37337 ;
  assign n37339 = n37151 | n37155 ;
  assign n37340 = ~n37338 & n37339 ;
  assign n37341 = n36559 & ~n37338 ;
  assign n37342 = n36475 & ~n37341 ;
  assign n37343 = ~n37340 & n37342 ;
  assign n37344 = x299 & n36468 ;
  assign n37345 = n36471 & n37344 ;
  assign n37346 = n36497 | n37345 ;
  assign n37347 = x1152 & n37346 ;
  assign n37348 = ~n37343 & n37347 ;
  assign n37349 = n36512 & ~n37341 ;
  assign n37350 = n37282 & ~n37349 ;
  assign n37351 = n37348 | n37350 ;
  assign n37352 = ( ~x1149 & n37336 ) | ( ~x1149 & n37351 ) | ( n37336 & n37351 ) ;
  assign n37353 = ~n37335 & n37352 ;
  assign n37354 = n37289 | n37353 ;
  assign n37355 = ( x209 & x213 ) | ( x209 & n37354 ) | ( x213 & n37354 ) ;
  assign n37356 = n36765 | n37210 ;
  assign n37357 = ~n36713 & n37194 ;
  assign n37358 = x1150 & ~n37357 ;
  assign n37359 = n37356 & n37358 ;
  assign n37360 = ~x1150 & x1151 ;
  assign n37361 = n36805 & n37360 ;
  assign n37362 = x1149 | n37361 ;
  assign n37363 = n37359 | n37362 ;
  assign n37364 = ~n36827 & n37109 ;
  assign n37365 = n36798 | n37126 ;
  assign n37366 = ~x1150 & n37365 ;
  assign n37367 = ~n37364 & n37366 ;
  assign n37368 = x1151 | n36735 ;
  assign n37369 = ~n36724 & n37140 ;
  assign n37370 = n37368 & ~n37369 ;
  assign n37371 = ( x1149 & n37255 ) | ( x1149 & ~n37370 ) | ( n37255 & ~n37370 ) ;
  assign n37372 = ~n37367 & n37371 ;
  assign n37373 = n37363 & ~n37372 ;
  assign n37374 = ( x209 & ~x213 ) | ( x209 & n37373 ) | ( ~x213 & n37373 ) ;
  assign n37375 = n37355 | n37374 ;
  assign n37376 = ~n37221 & n37375 ;
  assign n37377 = x230 & ~n37376 ;
  assign n37378 = x230 | x241 ;
  assign n37379 = ~n37377 & n37378 ;
  assign n37380 = x230 | x242 ;
  assign n37381 = x219 & ~n35106 ;
  assign n37382 = n35103 & ~n37381 ;
  assign n37383 = x214 & n36028 ;
  assign n37384 = ~x214 & n36837 ;
  assign n37385 = n37383 | n37384 ;
  assign n37386 = ( x212 & x219 ) | ( x212 & n37385 ) | ( x219 & n37385 ) ;
  assign n37387 = ( ~x212 & x219 ) | ( ~x212 & n36838 ) | ( x219 & n36838 ) ;
  assign n37388 = n37386 | n37387 ;
  assign n37389 = n37382 & n37388 ;
  assign n37390 = x199 & x1144 ;
  assign n37391 = x200 | n37390 ;
  assign n37392 = n36956 | n37391 ;
  assign n37393 = x299 | n36965 ;
  assign n37394 = n37392 & ~n37393 ;
  assign n37395 = n35136 & n37394 ;
  assign n37396 = n36859 | n37395 ;
  assign n37397 = ( x207 & x208 ) | ( x207 & n37394 ) | ( x208 & n37394 ) ;
  assign n37398 = x299 | n36044 ;
  assign n37399 = n36042 | n37391 ;
  assign n37400 = ~n37398 & n37399 ;
  assign n37401 = ( ~x207 & x208 ) | ( ~x207 & n37400 ) | ( x208 & n37400 ) ;
  assign n37402 = n37397 & n37401 ;
  assign n37403 = n37396 | n37402 ;
  assign n37404 = ~x211 & n37403 ;
  assign n37405 = n36208 | n37395 ;
  assign n37406 = n37402 | n37405 ;
  assign n37407 = x211 & n37406 ;
  assign n37408 = n37404 | n37407 ;
  assign n37409 = x214 | n37408 ;
  assign n37410 = ( x211 & x214 ) | ( x211 & ~n37406 ) | ( x214 & ~n37406 ) ;
  assign n37411 = n35446 | n37395 ;
  assign n37412 = n37402 | n37411 ;
  assign n37413 = ( x211 & ~x214 ) | ( x211 & n37412 ) | ( ~x214 & n37412 ) ;
  assign n37414 = n37410 & ~n37413 ;
  assign n37415 = x212 & ~n37414 ;
  assign n37416 = n37409 & n37415 ;
  assign n37417 = n35517 & n37394 ;
  assign n37418 = n37402 | n37417 ;
  assign n37419 = x214 | n37418 ;
  assign n37420 = ~x212 & n37419 ;
  assign n37421 = x214 & ~n37408 ;
  assign n37422 = n37420 & ~n37421 ;
  assign n37423 = x219 | n37422 ;
  assign n37424 = n37416 | n37423 ;
  assign n37425 = ~n35101 & n37418 ;
  assign n37426 = x219 & ~n37425 ;
  assign n37427 = n35101 & n37412 ;
  assign n37428 = n37426 & ~n37427 ;
  assign n37429 = n6785 | n37428 ;
  assign n37430 = n37424 & ~n37429 ;
  assign n37431 = n37389 | n37430 ;
  assign n37432 = x213 & ~n37431 ;
  assign n37433 = x211 & ~n37417 ;
  assign n37434 = n35101 & ~n35478 ;
  assign n37435 = ~n37395 & n37434 ;
  assign n37436 = n37433 | n37435 ;
  assign n37437 = x219 & n37436 ;
  assign n37438 = n35100 | n37417 ;
  assign n37439 = n8894 & ~n35147 ;
  assign n37440 = ~n35118 & n35442 ;
  assign n37441 = n37439 | n37440 ;
  assign n37442 = x219 | n37395 ;
  assign n37443 = n37441 & ~n37442 ;
  assign n37444 = n37438 & ~n37443 ;
  assign n37445 = ~n37437 & n37444 ;
  assign n37446 = n37402 | n37445 ;
  assign n37447 = ~n6785 & n37446 ;
  assign n37448 = x213 | n35117 ;
  assign n37449 = n37447 | n37448 ;
  assign n37450 = ~n37432 & n37449 ;
  assign n37451 = x209 & ~n37450 ;
  assign n37452 = n35106 & n35734 ;
  assign n37453 = ( ~x219 & n37388 ) | ( ~x219 & n37452 ) | ( n37388 & n37452 ) ;
  assign n37454 = x299 & ~n37453 ;
  assign n37455 = n6785 | n37454 ;
  assign n37456 = n35153 & ~n37455 ;
  assign n37457 = n37389 | n37456 ;
  assign n37458 = ( x209 & x213 ) | ( x209 & n37457 ) | ( x213 & n37457 ) ;
  assign n37459 = ( x209 & ~x213 ) | ( x209 & n35162 ) | ( ~x213 & n35162 ) ;
  assign n37460 = n37458 | n37459 ;
  assign n37461 = ~n37451 & n37460 ;
  assign n37462 = x230 & ~n37461 ;
  assign n37463 = n37380 & ~n37462 ;
  assign n37464 = x243 & ~x1091 ;
  assign n37465 = x83 | x85 ;
  assign n37466 = x314 & n37465 ;
  assign n37467 = x802 & n37466 ;
  assign n37468 = x276 & n37467 ;
  assign n37469 = x1091 | n37468 ;
  assign n37470 = x271 & n37469 ;
  assign n37471 = x1091 | n37470 ;
  assign n37472 = x273 & n37471 ;
  assign n37473 = x1091 | n37472 ;
  assign n37474 = ~x200 & n37473 ;
  assign n37475 = x199 & n37473 ;
  assign n37476 = x81 | n37465 ;
  assign n37477 = x314 & n37476 ;
  assign n37478 = x802 & n37477 ;
  assign n37479 = x276 & n37478 ;
  assign n37480 = ~x1091 & n37479 ;
  assign n37481 = x271 & n37480 ;
  assign n37482 = x273 & n37481 ;
  assign n37483 = n37472 | n37482 ;
  assign n37484 = x1091 | n37483 ;
  assign n37485 = ~x199 & n37484 ;
  assign n37486 = n37475 | n37485 ;
  assign n37487 = n37480 & n37486 ;
  assign n37488 = x299 | n37487 ;
  assign n37489 = n37475 | n37488 ;
  assign n37490 = n37474 | n37489 ;
  assign n37491 = x299 & ~n37482 ;
  assign n37492 = n37490 & ~n37491 ;
  assign n37493 = n37464 | n37492 ;
  assign n37494 = x200 | n37480 ;
  assign n37495 = n37486 & n37494 ;
  assign n37496 = x299 | n37495 ;
  assign n37497 = n37475 | n37496 ;
  assign n37498 = ~x1091 & n37468 ;
  assign n37499 = x271 & n37498 ;
  assign n37500 = x273 & n37499 ;
  assign n37501 = x299 & ~n37500 ;
  assign n37502 = n37474 | n37488 ;
  assign n37503 = n37485 | n37502 ;
  assign n37504 = ~n37501 & n37503 ;
  assign n37505 = n37497 & n37504 ;
  assign n37506 = x299 & ~n37473 ;
  assign n37507 = n37502 & ~n37506 ;
  assign n37508 = x243 & ~n37507 ;
  assign n37509 = ~n37505 & n37508 ;
  assign n37510 = x1155 & ~n37509 ;
  assign n37511 = ~n37482 & n37506 ;
  assign n37512 = n37503 & ~n37511 ;
  assign n37513 = x1155 & n37512 ;
  assign n37514 = n37510 | n37513 ;
  assign n37515 = ~n37491 & n37496 ;
  assign n37516 = ~x243 & n37515 ;
  assign n37517 = n37490 & n37516 ;
  assign n37518 = n37514 & ~n37517 ;
  assign n37519 = n37485 | n37496 ;
  assign n37520 = n37490 & n37519 ;
  assign n37521 = ~n37511 & n37520 ;
  assign n37522 = x243 | n37521 ;
  assign n37523 = ~n37491 & n37497 ;
  assign n37524 = x243 & n37503 ;
  assign n37525 = n37523 & n37524 ;
  assign n37526 = n37522 & ~n37525 ;
  assign n37527 = x1155 | n37526 ;
  assign n37528 = ~n37518 & n37527 ;
  assign n37529 = n37493 & n37528 ;
  assign n37530 = x1156 & ~n37529 ;
  assign n37531 = ~n37506 & n37519 ;
  assign n37532 = x243 | n37531 ;
  assign n37533 = ~x1155 & n37532 ;
  assign n37534 = n37488 & ~n37491 ;
  assign n37535 = ~x1155 & n37534 ;
  assign n37536 = n37533 | n37535 ;
  assign n37537 = ~n37491 & n37502 ;
  assign n37538 = x243 & n37537 ;
  assign n37539 = n37489 & n37538 ;
  assign n37540 = n37536 & ~n37539 ;
  assign n37541 = x1156 | n37540 ;
  assign n37542 = n37496 & ~n37511 ;
  assign n37543 = x243 | n37542 ;
  assign n37544 = x1155 & n37543 ;
  assign n37545 = ~n37538 & n37544 ;
  assign n37546 = n37541 | n37545 ;
  assign n37547 = x1157 & n37546 ;
  assign n37548 = ~n37530 & n37547 ;
  assign n37549 = x243 & n37534 ;
  assign n37550 = x243 | x1091 ;
  assign n37551 = n37488 & ~n37501 ;
  assign n37552 = n37550 | n37551 ;
  assign n37553 = ~x1155 & n37552 ;
  assign n37554 = n37535 | n37553 ;
  assign n37555 = ~n37549 & n37554 ;
  assign n37556 = x1156 | n37555 ;
  assign n37557 = x1155 & ~n37464 ;
  assign n37558 = n37475 & n37557 ;
  assign n37559 = n37545 | n37558 ;
  assign n37560 = n37556 | n37559 ;
  assign n37561 = n37485 | n37488 ;
  assign n37562 = ~n37511 & n37561 ;
  assign n37563 = x243 & ~n37562 ;
  assign n37564 = n37489 & ~n37491 ;
  assign n37565 = ~x243 & n37564 ;
  assign n37566 = n37563 | n37565 ;
  assign n37567 = ~x1155 & n37537 ;
  assign n37568 = ~n37480 & n37567 ;
  assign n37569 = x1156 & ~n37568 ;
  assign n37570 = ~n37566 & n37569 ;
  assign n37571 = n37560 & ~n37570 ;
  assign n37572 = ( x211 & n36056 ) | ( x211 & ~n37571 ) | ( n36056 & ~n37571 ) ;
  assign n37573 = ~n37548 & n37572 ;
  assign n37574 = x1156 & ~n37528 ;
  assign n37575 = n37502 & ~n37511 ;
  assign n37576 = x243 & ~n37575 ;
  assign n37577 = n37516 | n37576 ;
  assign n37578 = n37541 | n37577 ;
  assign n37579 = x1157 & n37578 ;
  assign n37580 = ~n37574 & n37579 ;
  assign n37581 = n37566 | n37577 ;
  assign n37582 = x1155 & n37581 ;
  assign n37583 = n37556 | n37582 ;
  assign n37584 = ~x1155 & n37575 ;
  assign n37585 = ~n37515 & n37584 ;
  assign n37586 = n37570 & ~n37585 ;
  assign n37587 = n37583 & ~n37586 ;
  assign n37588 = ( x211 & ~n35174 ) | ( x211 & n37587 ) | ( ~n35174 & n37587 ) ;
  assign n37589 = n37580 | n37588 ;
  assign n37590 = ~x219 & n37589 ;
  assign n37591 = ~n37573 & n37590 ;
  assign n37592 = x253 & x254 ;
  assign n37593 = x267 & n37592 ;
  assign n37594 = ~x263 & n37593 ;
  assign n37595 = n37490 & ~n37506 ;
  assign n37596 = ~x243 & n37595 ;
  assign n37597 = n37496 & ~n37501 ;
  assign n37598 = n37596 & n37597 ;
  assign n37599 = n37510 & ~n37598 ;
  assign n37600 = x243 & ~n37505 ;
  assign n37601 = n37596 | n37600 ;
  assign n37602 = n37493 & n37532 ;
  assign n37603 = n37601 & n37602 ;
  assign n37604 = x1155 | n37603 ;
  assign n37605 = ~n37599 & n37604 ;
  assign n37606 = x1156 & ~n37605 ;
  assign n37607 = ~x243 & x1155 ;
  assign n37608 = n37597 & n37607 ;
  assign n37609 = x1156 | n37608 ;
  assign n37610 = n37508 | n37609 ;
  assign n37611 = ~n37501 & n37519 ;
  assign n37612 = ( x243 & ~x1155 ) | ( x243 & n37611 ) | ( ~x1155 & n37611 ) ;
  assign n37613 = ( x243 & x1155 ) | ( x243 & n37489 ) | ( x1155 & n37489 ) ;
  assign n37614 = n37612 & ~n37613 ;
  assign n37615 = n37610 | n37614 ;
  assign n37616 = n35174 & n37615 ;
  assign n37617 = ~n37606 & n37616 ;
  assign n37618 = ~n37501 & n37561 ;
  assign n37619 = x1155 & n37618 ;
  assign n37620 = n37496 & n37618 ;
  assign n37621 = n37619 | n37620 ;
  assign n37622 = x243 & n37621 ;
  assign n37623 = n37489 & ~n37506 ;
  assign n37624 = x243 | n37623 ;
  assign n37625 = n37568 | n37624 ;
  assign n37626 = ~n37622 & n37625 ;
  assign n37627 = x1156 & ~n37626 ;
  assign n37628 = ~n37501 & n37502 ;
  assign n37629 = x243 & n37628 ;
  assign n37630 = n37561 & n37629 ;
  assign n37631 = n37497 & ~n37506 ;
  assign n37632 = x243 | n37631 ;
  assign n37633 = x1155 & n37632 ;
  assign n37634 = ~n37630 & n37633 ;
  assign n37635 = x243 & n37551 ;
  assign n37636 = n37553 & ~n37635 ;
  assign n37637 = x1156 | n37636 ;
  assign n37638 = n37634 | n37637 ;
  assign n37639 = ~x1157 & n37638 ;
  assign n37640 = ~n37627 & n37639 ;
  assign n37641 = n37489 & n37628 ;
  assign n37642 = x243 & n37641 ;
  assign n37643 = n37532 & ~n37642 ;
  assign n37644 = n37544 & ~n37629 ;
  assign n37645 = ( ~x1155 & n37643 ) | ( ~x1155 & n37644 ) | ( n37643 & n37644 ) ;
  assign n37646 = ( x1156 & n36056 ) | ( x1156 & n37645 ) | ( n36056 & n37645 ) ;
  assign n37647 = x243 & n37504 ;
  assign n37648 = n37544 & ~n37647 ;
  assign n37649 = n37533 | n37648 ;
  assign n37650 = n37601 & n37649 ;
  assign n37651 = ( ~x1156 & n36056 ) | ( ~x1156 & n37650 ) | ( n36056 & n37650 ) ;
  assign n37652 = n37646 & n37651 ;
  assign n37653 = n37640 | n37652 ;
  assign n37654 = n37617 | n37653 ;
  assign n37655 = x219 & n37654 ;
  assign n37656 = n37594 & ~n37655 ;
  assign n37657 = ~n37591 & n37656 ;
  assign n37658 = ~x299 & x1091 ;
  assign n37659 = n35532 & n37658 ;
  assign n37660 = n37550 & ~n37659 ;
  assign n37661 = x1156 & ~n37660 ;
  assign n37662 = x1091 & n35614 ;
  assign n37663 = n36169 & n37662 ;
  assign n37664 = n37661 | n37663 ;
  assign n37665 = ~x299 & n35290 ;
  assign n37666 = x1091 & ~n37665 ;
  assign n37667 = n37464 | n37666 ;
  assign n37668 = ~x1155 & n37550 ;
  assign n37669 = n37464 | n37668 ;
  assign n37670 = n35230 | n37669 ;
  assign n37671 = n37667 & n37670 ;
  assign n37672 = x1156 | n37671 ;
  assign n37673 = ~n37664 & n37672 ;
  assign n37674 = x1157 & ~n37673 ;
  assign n37675 = x199 & x1091 ;
  assign n37676 = ~x299 & n37675 ;
  assign n37677 = n37557 & ~n37676 ;
  assign n37678 = x1156 & ~n37677 ;
  assign n37679 = x1155 | n37464 ;
  assign n37680 = ~n9578 & n37658 ;
  assign n37681 = n37679 | n37680 ;
  assign n37682 = n37678 & n37681 ;
  assign n37683 = n37662 | n37669 ;
  assign n37684 = ~x1156 & n37683 ;
  assign n37685 = x1157 | n37684 ;
  assign n37686 = n37682 | n37685 ;
  assign n37687 = ~n37674 & n37686 ;
  assign n37688 = x211 & ~n37687 ;
  assign n37689 = n37660 & n37678 ;
  assign n37690 = x1155 | n37667 ;
  assign n37691 = x200 & x1091 ;
  assign n37692 = ~x299 & n37691 ;
  assign n37693 = n37557 & ~n37692 ;
  assign n37694 = x1156 | n37693 ;
  assign n37695 = n37690 & ~n37694 ;
  assign n37696 = n37689 | n37695 ;
  assign n37697 = ( x211 & x1157 ) | ( x211 & n37696 ) | ( x1157 & n37696 ) ;
  assign n37698 = x1091 & ~n9579 ;
  assign n37699 = n37679 | n37698 ;
  assign n37700 = ~n37677 & n37699 ;
  assign n37701 = x200 & ~x1156 ;
  assign n37702 = n37658 & n37701 ;
  assign n37703 = n37700 | n37702 ;
  assign n37704 = ( x211 & ~x1157 ) | ( x211 & n37703 ) | ( ~x1157 & n37703 ) ;
  assign n37705 = n37697 | n37704 ;
  assign n37706 = ~n37688 & n37705 ;
  assign n37707 = x219 | n37706 ;
  assign n37708 = n36056 & ~n37661 ;
  assign n37709 = n37672 & n37708 ;
  assign n37710 = x219 & ~n37709 ;
  assign n37711 = x299 & x1091 ;
  assign n37712 = n37703 | n37711 ;
  assign n37713 = ~x1157 & n37712 ;
  assign n37714 = x1091 & ~n35291 ;
  assign n37715 = n37679 | n37714 ;
  assign n37716 = ~n37693 & n37715 ;
  assign n37717 = x1156 | n37716 ;
  assign n37718 = n35174 & n37717 ;
  assign n37719 = ~n37664 & n37718 ;
  assign n37720 = n37713 | n37719 ;
  assign n37721 = n37710 & ~n37720 ;
  assign n37722 = n37707 & ~n37721 ;
  assign n37723 = n37594 | n37722 ;
  assign n37724 = ~n6785 & n37723 ;
  assign n37725 = ~n37657 & n37724 ;
  assign n37726 = x272 & x283 ;
  assign n37727 = x275 & n37726 ;
  assign n37728 = x268 & n37727 ;
  assign n37729 = n35174 & ~n37464 ;
  assign n37730 = ~n37498 & n37729 ;
  assign n37731 = ( x243 & n37473 ) | ( x243 & ~n37730 ) | ( n37473 & ~n37730 ) ;
  assign n37732 = ( x243 & n37500 ) | ( x243 & n37730 ) | ( n37500 & n37730 ) ;
  assign n37733 = n37731 & ~n37732 ;
  assign n37734 = x219 & ~n37733 ;
  assign n37735 = n37464 & ~n37483 ;
  assign n37736 = ~x243 & n37482 ;
  assign n37737 = n35168 | n35175 ;
  assign n37738 = x1091 & ~n37737 ;
  assign n37739 = x219 | n37738 ;
  assign n37740 = n37736 | n37739 ;
  assign n37741 = n37735 | n37740 ;
  assign n37742 = ~n37734 & n37741 ;
  assign n37743 = ( n6785 & ~n37594 ) | ( n6785 & n37742 ) | ( ~n37594 & n37742 ) ;
  assign n37744 = ~x219 & n37737 ;
  assign n37745 = x1157 & n35201 ;
  assign n37746 = n37744 | n37745 ;
  assign n37747 = x1091 & n37746 ;
  assign n37748 = n37550 & ~n37747 ;
  assign n37749 = ( n6785 & n37594 ) | ( n6785 & n37748 ) | ( n37594 & n37748 ) ;
  assign n37750 = n37743 & n37749 ;
  assign n37751 = n37728 & ~n37750 ;
  assign n37752 = ~n37725 & n37751 ;
  assign n37753 = ( n6785 & n37728 ) | ( n6785 & n37748 ) | ( n37728 & n37748 ) ;
  assign n37754 = ( ~n6785 & n37722 ) | ( ~n6785 & n37728 ) | ( n37722 & n37728 ) ;
  assign n37755 = n37753 | n37754 ;
  assign n37756 = ~x230 & n37755 ;
  assign n37757 = ~n37752 & n37756 ;
  assign n37758 = ( ~x230 & n14313 ) | ( ~x230 & n37746 ) | ( n14313 & n37746 ) ;
  assign n37759 = x199 & ~n36218 ;
  assign n37760 = n35531 & ~n37701 ;
  assign n37761 = ~n37759 & n37760 ;
  assign n37762 = ( x230 & n14313 ) | ( x230 & ~n37761 ) | ( n14313 & ~n37761 ) ;
  assign n37763 = ~n37758 & n37762 ;
  assign n37764 = n37757 | n37763 ;
  assign n37765 = x230 | x244 ;
  assign n37766 = x213 & ~n37092 ;
  assign n37767 = ~n35444 & n36974 ;
  assign n37768 = n37086 | n37767 ;
  assign n37769 = x214 | n37768 ;
  assign n37770 = ~n35107 & n36909 ;
  assign n37771 = x212 & ~n37770 ;
  assign n37772 = n37769 & n37771 ;
  assign n37773 = n36980 & n37772 ;
  assign n37774 = n36981 & n37768 ;
  assign n37775 = ( ~x214 & n37060 ) | ( ~x214 & n37774 ) | ( n37060 & n37774 ) ;
  assign n37776 = x219 | n37775 ;
  assign n37777 = n37773 | n37776 ;
  assign n37778 = x211 | n35412 ;
  assign n37779 = n37063 | n37778 ;
  assign n37780 = n37071 & n37779 ;
  assign n37781 = n37068 & ~n37780 ;
  assign n37782 = n37042 | n37781 ;
  assign n37783 = n37777 & ~n37782 ;
  assign n37784 = n36973 & n37772 ;
  assign n37785 = x214 & ~n37768 ;
  assign n37786 = n37035 & ~n37785 ;
  assign n37787 = x219 | n37786 ;
  assign n37788 = n37784 | n37787 ;
  assign n37789 = x299 & n36033 ;
  assign n37790 = x1147 & ~n37789 ;
  assign n37791 = ~n37013 & n37790 ;
  assign n37792 = n37788 & n37791 ;
  assign n37793 = x213 | n36035 ;
  assign n37794 = n37792 | n37793 ;
  assign n37795 = n37783 | n37794 ;
  assign n37796 = ~n37766 & n37795 ;
  assign n37797 = x209 & ~n37796 ;
  assign n37798 = n36877 | n36880 ;
  assign n37799 = ~n36852 & n37798 ;
  assign n37800 = n36877 | n36879 ;
  assign n37801 = ( n8894 & n35474 ) | ( n8894 & n36925 ) | ( n35474 & n36925 ) ;
  assign n37802 = ( ~n8894 & n35474 ) | ( ~n8894 & n36866 ) | ( n35474 & n36866 ) ;
  assign n37803 = n37801 & n37802 ;
  assign n37804 = n37800 & n37803 ;
  assign n37805 = n36048 | n36943 ;
  assign n37806 = n37804 | n37805 ;
  assign n37807 = ~n6785 & n37806 ;
  assign n37808 = n37799 | n37807 ;
  assign n37809 = ( x209 & x213 ) | ( x209 & n37808 ) | ( x213 & n37808 ) ;
  assign n37810 = ( x209 & ~x213 ) | ( x209 & n36054 ) | ( ~x213 & n36054 ) ;
  assign n37811 = n37809 | n37810 ;
  assign n37812 = ~n37797 & n37811 ;
  assign n37813 = x230 & ~n37812 ;
  assign n37814 = n37765 & ~n37813 ;
  assign n37815 = x1146 & n36473 ;
  assign n37816 = x1147 | n37815 ;
  assign n37817 = n36469 & n36807 ;
  assign n37818 = n37816 | n37817 ;
  assign n37819 = x199 & x1146 ;
  assign n37820 = n35290 & ~n37819 ;
  assign n37821 = n36958 | n37820 ;
  assign n37822 = x208 & ~n37821 ;
  assign n37823 = x207 | n37822 ;
  assign n37824 = n36325 | n37820 ;
  assign n37825 = n37823 & ~n37824 ;
  assign n37826 = ~x208 & n36859 ;
  assign n37827 = x200 | n37819 ;
  assign n37828 = ~n36958 & n37827 ;
  assign n37829 = x207 & n37828 ;
  assign n37830 = x1146 & n35291 ;
  assign n37831 = n37829 | n37830 ;
  assign n37832 = x208 & n37831 ;
  assign n37833 = n37826 | n37832 ;
  assign n37834 = n37825 | n37833 ;
  assign n37835 = ~x299 & n37834 ;
  assign n37836 = x214 | n37835 ;
  assign n37837 = ~x212 & n37836 ;
  assign n37838 = ( n8790 & n36326 ) | ( n8790 & n37828 ) | ( n36326 & n37828 ) ;
  assign n37839 = x211 & ~n37838 ;
  assign n37840 = x299 | n37828 ;
  assign n37841 = n37834 & n37840 ;
  assign n37842 = x299 | n37841 ;
  assign n37843 = x211 | n37842 ;
  assign n37844 = ~n37839 & n37843 ;
  assign n37845 = n37835 | n37844 ;
  assign n37846 = n37837 & n37845 ;
  assign n37847 = x219 | n37846 ;
  assign n37848 = x214 & ~n36896 ;
  assign n37849 = ~n37835 & n37848 ;
  assign n37850 = ( x212 & n8894 ) | ( x212 & n37845 ) | ( n8894 & n37845 ) ;
  assign n37851 = ~n37849 & n37850 ;
  assign n37852 = n37847 | n37851 ;
  assign n37853 = ~n35101 & n37835 ;
  assign n37854 = x219 & ~n37853 ;
  assign n37855 = n35101 & n37834 ;
  assign n37856 = n37854 & ~n37855 ;
  assign n37857 = n6785 | n37856 ;
  assign n37858 = n37852 & ~n37857 ;
  assign n37859 = n37818 | n37858 ;
  assign n37860 = x1147 & ~n36469 ;
  assign n37861 = ~n37815 & n37860 ;
  assign n37862 = n35221 | n37820 ;
  assign n37863 = ~n8790 & n37862 ;
  assign n37864 = x207 & ~n37821 ;
  assign n37865 = n35517 | n37864 ;
  assign n37866 = ~n37863 & n37865 ;
  assign n37867 = x214 | n37866 ;
  assign n37868 = ~x212 & n37867 ;
  assign n37869 = ~n35221 & n37827 ;
  assign n37870 = ~x207 & n37869 ;
  assign n37871 = n36859 | n37870 ;
  assign n37872 = n37864 | n37871 ;
  assign n37873 = x208 & n37872 ;
  assign n37874 = ~x299 & n37873 ;
  assign n37875 = n35136 & ~n37862 ;
  assign n37876 = n37822 | n37875 ;
  assign n37877 = n37874 | n37876 ;
  assign n37878 = x299 | n37877 ;
  assign n37879 = n37868 & n37878 ;
  assign n37880 = x219 | n37879 ;
  assign n37881 = x212 & n37878 ;
  assign n37882 = n36859 | n37877 ;
  assign n37883 = n8652 & ~n37882 ;
  assign n37884 = n37881 & ~n37883 ;
  assign n37885 = n37880 | n37884 ;
  assign n37886 = ~n35101 & n37866 ;
  assign n37887 = x219 & ~n37886 ;
  assign n37888 = n35101 & n37882 ;
  assign n37889 = n37887 & ~n37888 ;
  assign n37890 = n6785 | n37889 ;
  assign n37891 = n37885 & ~n37890 ;
  assign n37892 = n37861 & ~n37891 ;
  assign n37893 = x1148 & ~n37892 ;
  assign n37894 = n37859 & n37893 ;
  assign n37895 = n37015 | n37861 ;
  assign n37896 = n8790 | n37869 ;
  assign n37897 = n37865 & n37896 ;
  assign n37898 = ~x214 & n37897 ;
  assign n37899 = x212 | n37898 ;
  assign n37900 = n11103 | n37897 ;
  assign n37901 = n35136 & n37869 ;
  assign n37902 = n37826 | n37901 ;
  assign n37903 = n37873 | n37902 ;
  assign n37904 = x299 | n37903 ;
  assign n37905 = x214 & n37904 ;
  assign n37906 = ~x211 & n37878 ;
  assign n37907 = n37866 | n37906 ;
  assign n37908 = n37905 & n37907 ;
  assign n37909 = x212 & ~n37908 ;
  assign n37910 = ( x214 & ~n37900 ) | ( x214 & n37909 ) | ( ~n37900 & n37909 ) ;
  assign n37911 = x214 & ~n37909 ;
  assign n37912 = ( n37899 & ~n37910 ) | ( n37899 & n37911 ) | ( ~n37910 & n37911 ) ;
  assign n37913 = x219 | n37912 ;
  assign n37914 = x1146 | n35398 ;
  assign n37915 = n36905 & n37914 ;
  assign n37916 = n37913 | n37915 ;
  assign n37917 = n35100 & n37897 ;
  assign n37918 = n35101 | n37917 ;
  assign n37919 = n37903 & n37918 ;
  assign n37920 = x219 & ~n37897 ;
  assign n37921 = ( x219 & n35100 ) | ( x219 & n37920 ) | ( n35100 & n37920 ) ;
  assign n37922 = ~n37919 & n37921 ;
  assign n37923 = n6785 | n37922 ;
  assign n37924 = n37916 & ~n37923 ;
  assign n37925 = n37895 & ~n37924 ;
  assign n37926 = n37259 | n37835 ;
  assign n37927 = n37831 & n37926 ;
  assign n37928 = x219 | n37927 ;
  assign n37929 = x219 & ~n37838 ;
  assign n37930 = n35734 | n37929 ;
  assign n37931 = n35100 & ~n37839 ;
  assign n37932 = n37841 & n37931 ;
  assign n37933 = n37930 & ~n37932 ;
  assign n37934 = n6785 | n37933 ;
  assign n37935 = n37928 & ~n37934 ;
  assign n37936 = n37816 | n37935 ;
  assign n37937 = ~x1148 & n37936 ;
  assign n37938 = ~n37925 & n37937 ;
  assign n37939 = n37894 | n37938 ;
  assign n37940 = x213 & n37939 ;
  assign n37941 = ~n35444 & n37842 ;
  assign n37942 = x211 | n37941 ;
  assign n37943 = n37931 & n37942 ;
  assign n37944 = n37930 & ~n37943 ;
  assign n37945 = n37042 | n37944 ;
  assign n37946 = x299 & n37385 ;
  assign n37947 = n37835 | n37946 ;
  assign n37948 = x212 & n37947 ;
  assign n37949 = n37840 & n37948 ;
  assign n37950 = x219 | n37949 ;
  assign n37951 = n36866 | n37835 ;
  assign n37952 = x214 & n37842 ;
  assign n37953 = n37951 & n37952 ;
  assign n37954 = ~x214 & n37838 ;
  assign n37955 = x212 | n37954 ;
  assign n37956 = n37953 | n37955 ;
  assign n37957 = ( ~x212 & n37950 ) | ( ~x212 & n37956 ) | ( n37950 & n37956 ) ;
  assign n37958 = ~n37945 & n37957 ;
  assign n37959 = n35446 | n37877 ;
  assign n37960 = n37904 & n37959 ;
  assign n37961 = x211 | n37960 ;
  assign n37962 = n37918 & n37961 ;
  assign n37963 = n37921 & ~n37962 ;
  assign n37964 = x1147 & ~n6785 ;
  assign n37965 = n37877 | n37946 ;
  assign n37966 = x212 & n37965 ;
  assign n37967 = n37904 & n37966 ;
  assign n37968 = x219 | n37967 ;
  assign n37969 = n36866 | n37877 ;
  assign n37970 = n37905 & n37969 ;
  assign n37971 = n37899 | n37970 ;
  assign n37972 = ( ~x212 & n37968 ) | ( ~x212 & n37971 ) | ( n37968 & n37971 ) ;
  assign n37973 = n37964 & n37972 ;
  assign n37974 = ~n37963 & n37973 ;
  assign n37975 = x1148 | n37389 ;
  assign n37976 = n37974 | n37975 ;
  assign n37977 = n37958 | n37976 ;
  assign n37978 = n37837 & n37951 ;
  assign n37979 = x219 | n37948 ;
  assign n37980 = n37978 | n37979 ;
  assign n37981 = x299 | n37834 ;
  assign n37982 = n35101 & n37981 ;
  assign n37983 = ~n35444 & n37982 ;
  assign n37984 = n37854 & ~n37983 ;
  assign n37985 = n37042 | n37984 ;
  assign n37986 = n37980 & ~n37985 ;
  assign n37987 = x214 & ~n37969 ;
  assign n37988 = n37868 & ~n37987 ;
  assign n37989 = x219 | n37966 ;
  assign n37990 = n37988 | n37989 ;
  assign n37991 = n35101 & n37959 ;
  assign n37992 = n37887 & ~n37991 ;
  assign n37993 = n37964 & ~n37992 ;
  assign n37994 = n37990 & n37993 ;
  assign n37995 = x1148 & ~n37389 ;
  assign n37996 = ~n37994 & n37995 ;
  assign n37997 = ~n37986 & n37996 ;
  assign n37998 = x213 | n37997 ;
  assign n37999 = n37977 & ~n37998 ;
  assign n38000 = x209 & ~n37999 ;
  assign n38001 = ~n37940 & n38000 ;
  assign n38002 = n35100 & n37404 ;
  assign n38003 = n37426 & ~n38002 ;
  assign n38004 = n6785 | n38003 ;
  assign n38005 = x299 | n37406 ;
  assign n38006 = ~x211 & n38005 ;
  assign n38007 = x211 & n37403 ;
  assign n38008 = n38006 | n38007 ;
  assign n38009 = x214 & n38008 ;
  assign n38010 = ~x214 & n38005 ;
  assign n38011 = n38009 | n38010 ;
  assign n38012 = x212 & n38011 ;
  assign n38013 = n37420 & n38005 ;
  assign n38014 = x219 | n38013 ;
  assign n38015 = n38012 | n38014 ;
  assign n38016 = ~n38004 & n38015 ;
  assign n38017 = n37861 & ~n38016 ;
  assign n38018 = ~x299 & n37408 ;
  assign n38019 = n37848 & ~n38018 ;
  assign n38020 = x212 & ~n38019 ;
  assign n38021 = n37418 | n38006 ;
  assign n38022 = x214 | n38021 ;
  assign n38023 = n38020 & n38022 ;
  assign n38024 = n37420 & n38021 ;
  assign n38025 = x219 | n38024 ;
  assign n38026 = n38023 | n38025 ;
  assign n38027 = ~n38004 & n38026 ;
  assign n38028 = n37818 | n38027 ;
  assign n38029 = x1148 & n38028 ;
  assign n38030 = ~n38017 & n38029 ;
  assign n38031 = n37419 & n38020 ;
  assign n38032 = ~x212 & n37418 ;
  assign n38033 = x219 | n38032 ;
  assign n38034 = n38031 | n38033 ;
  assign n38035 = ~n38004 & n38034 ;
  assign n38036 = n37816 | n38035 ;
  assign n38037 = n11103 | n37418 ;
  assign n38038 = ~x214 & n38037 ;
  assign n38039 = n38009 | n38038 ;
  assign n38040 = x212 & n38039 ;
  assign n38041 = n37420 & n38037 ;
  assign n38042 = x219 | n38041 ;
  assign n38043 = n38040 | n38042 ;
  assign n38044 = ~n38004 & n38043 ;
  assign n38045 = n37895 & ~n38044 ;
  assign n38046 = x1148 | n38045 ;
  assign n38047 = n38036 & ~n38046 ;
  assign n38048 = n38030 | n38047 ;
  assign n38049 = ( x209 & x213 ) | ( x209 & n38048 ) | ( x213 & n38048 ) ;
  assign n38050 = ( x209 & ~x213 ) | ( x209 & n37431 ) | ( ~x213 & n37431 ) ;
  assign n38051 = n38049 | n38050 ;
  assign n38052 = ~n38001 & n38051 ;
  assign n38053 = x230 & ~n38052 ;
  assign n38054 = x230 | x245 ;
  assign n38055 = ~n38053 & n38054 ;
  assign n38056 = n11103 | n37838 ;
  assign n38057 = ( x212 & n35109 ) | ( x212 & ~n37844 ) | ( n35109 & ~n37844 ) ;
  assign n38058 = ( x214 & ~n38056 ) | ( x214 & n38057 ) | ( ~n38056 & n38057 ) ;
  assign n38059 = x214 & ~n38057 ;
  assign n38060 = ( n37955 & ~n38058 ) | ( n37955 & n38059 ) | ( ~n38058 & n38059 ) ;
  assign n38061 = x219 | n38060 ;
  assign n38062 = n37042 | n37929 ;
  assign n38063 = n38061 & ~n38062 ;
  assign n38064 = ~n37920 & n37964 ;
  assign n38065 = n37913 & n38064 ;
  assign n38066 = x1150 | n36739 ;
  assign n38067 = n38065 | n38066 ;
  assign n38068 = n38063 | n38067 ;
  assign n38069 = x1150 & ~n36469 ;
  assign n38070 = ( x214 & ~n37904 ) | ( x214 & n37909 ) | ( ~n37904 & n37909 ) ;
  assign n38071 = ( n37899 & n37911 ) | ( n37899 & ~n38070 ) | ( n37911 & ~n38070 ) ;
  assign n38072 = x219 | n38071 ;
  assign n38073 = ~n37920 & n38072 ;
  assign n38074 = ( x1147 & n6785 ) | ( x1147 & ~n38073 ) | ( n6785 & ~n38073 ) ;
  assign n38075 = ( x214 & ~n37842 ) | ( x214 & n38057 ) | ( ~n37842 & n38057 ) ;
  assign n38076 = ( n37955 & n38059 ) | ( n37955 & ~n38075 ) | ( n38059 & ~n38075 ) ;
  assign n38077 = x219 | n38076 ;
  assign n38078 = ~n37929 & n38077 ;
  assign n38079 = ( x1147 & ~n6785 ) | ( x1147 & n38078 ) | ( ~n6785 & n38078 ) ;
  assign n38080 = ~n38074 & n38079 ;
  assign n38081 = n38069 & ~n38080 ;
  assign n38082 = n38068 & ~n38081 ;
  assign n38083 = x1149 & ~n38082 ;
  assign n38084 = x1150 & n36849 ;
  assign n38085 = ~x1147 & n37841 ;
  assign n38086 = n14313 | n38085 ;
  assign n38087 = n38084 & n38086 ;
  assign n38088 = n37838 & ~n38084 ;
  assign n38089 = ( x1147 & ~n6785 ) | ( x1147 & n38088 ) | ( ~n6785 & n38088 ) ;
  assign n38090 = ( x1147 & n6785 ) | ( x1147 & ~n37897 ) | ( n6785 & ~n37897 ) ;
  assign n38091 = n38089 & ~n38090 ;
  assign n38092 = x1149 | n38091 ;
  assign n38093 = n38087 | n38092 ;
  assign n38094 = ~n38083 & n38093 ;
  assign n38095 = x1148 | n38094 ;
  assign n38096 = n37854 & ~n37982 ;
  assign n38097 = n37042 | n38096 ;
  assign n38098 = n37835 | n38056 ;
  assign n38099 = x214 & ~n38098 ;
  assign n38100 = n37850 & ~n38099 ;
  assign n38101 = n37847 | n38100 ;
  assign n38102 = ~n38097 & n38101 ;
  assign n38103 = n35100 & n37906 ;
  assign n38104 = n37887 & ~n38103 ;
  assign n38105 = n37964 & ~n38104 ;
  assign n38106 = x214 | n37907 ;
  assign n38107 = n11103 | n37877 ;
  assign n38108 = ( x212 & n35109 ) | ( x212 & n38107 ) | ( n35109 & n38107 ) ;
  assign n38109 = n38106 & n38108 ;
  assign n38110 = n37868 & n37907 ;
  assign n38111 = x219 | n38110 ;
  assign n38112 = n38109 | n38111 ;
  assign n38113 = n38105 & n38112 ;
  assign n38114 = x1150 & ~n36808 ;
  assign n38115 = ~n38113 & n38114 ;
  assign n38116 = ~n38102 & n38115 ;
  assign n38117 = x219 | n37926 ;
  assign n38118 = ~n38097 & n38117 ;
  assign n38119 = n37867 & n38108 ;
  assign n38120 = ~x212 & n37866 ;
  assign n38121 = x219 | n38120 ;
  assign n38122 = n38119 | n38121 ;
  assign n38123 = n38105 & n38122 ;
  assign n38124 = x1150 | n36473 ;
  assign n38125 = n38123 | n38124 ;
  assign n38126 = n38118 | n38125 ;
  assign n38127 = ~x1149 & n38126 ;
  assign n38128 = ~n38116 & n38127 ;
  assign n38129 = n37880 | n37881 ;
  assign n38130 = ~n38104 & n38129 ;
  assign n38131 = ~n4832 & n38130 ;
  assign n38132 = n4832 & n35475 ;
  assign n38133 = ~x57 & x1147 ;
  assign n38134 = ~n38132 & n38133 ;
  assign n38135 = ~n38131 & n38134 ;
  assign n38136 = x57 & ~n35475 ;
  assign n38137 = n4832 | n35474 ;
  assign n38138 = n37853 & ~n38137 ;
  assign n38139 = n35475 & n37981 ;
  assign n38140 = x57 | x1147 ;
  assign n38141 = n38132 | n38140 ;
  assign n38142 = n38139 | n38141 ;
  assign n38143 = n38138 | n38142 ;
  assign n38144 = ~n38136 & n38143 ;
  assign n38145 = ~n38135 & n38144 ;
  assign n38146 = x1150 & ~n38145 ;
  assign n38147 = n37952 | n38098 ;
  assign n38148 = x212 & n38147 ;
  assign n38149 = n37837 & ~n38099 ;
  assign n38150 = x219 | n38149 ;
  assign n38151 = n38148 | n38150 ;
  assign n38152 = ~n38097 & n38151 ;
  assign n38153 = n37264 & n37964 ;
  assign n38154 = n38130 & n38153 ;
  assign n38155 = x1150 | n36733 ;
  assign n38156 = n38154 | n38155 ;
  assign n38157 = n38152 | n38156 ;
  assign n38158 = x1149 & n38157 ;
  assign n38159 = ~n38146 & n38158 ;
  assign n38160 = x1148 & ~n38159 ;
  assign n38161 = ~n38128 & n38160 ;
  assign n38162 = x213 & ~n38161 ;
  assign n38163 = n38095 & n38162 ;
  assign n38164 = ~x213 & n37939 ;
  assign n38165 = x209 | n38164 ;
  assign n38166 = n38163 | n38165 ;
  assign n38167 = x1150 & ~n36828 ;
  assign n38168 = ( ~x1149 & n36799 ) | ( ~x1149 & n37336 ) | ( n36799 & n37336 ) ;
  assign n38169 = ~n38167 & n38168 ;
  assign n38170 = ( x1149 & ~x1150 ) | ( x1149 & n36725 ) | ( ~x1150 & n36725 ) ;
  assign n38171 = ( x1149 & x1150 ) | ( x1149 & n36735 ) | ( x1150 & n36735 ) ;
  assign n38172 = n38170 & n38171 ;
  assign n38173 = n38169 | n38172 ;
  assign n38174 = x1148 & n38173 ;
  assign n38175 = x1150 | n36766 ;
  assign n38176 = ( x1149 & n36714 ) | ( x1149 & n37255 ) | ( n36714 & n37255 ) ;
  assign n38177 = n38175 & n38176 ;
  assign n38178 = n36805 & n37336 ;
  assign n38179 = n38177 | n38178 ;
  assign n38180 = ~x1148 & n38179 ;
  assign n38181 = n38174 | n38180 ;
  assign n38182 = ( ~x209 & x213 ) | ( ~x209 & n38181 ) | ( x213 & n38181 ) ;
  assign n38183 = n37818 & ~n37861 ;
  assign n38184 = x219 & ~n36859 ;
  assign n38185 = n36720 | n38184 ;
  assign n38186 = n36732 & n36781 ;
  assign n38187 = n38185 & ~n38186 ;
  assign n38188 = n36783 & ~n36938 ;
  assign n38189 = n35110 | n38188 ;
  assign n38190 = n37243 & n38189 ;
  assign n38191 = x219 | n38190 ;
  assign n38192 = ~n38187 & n38191 ;
  assign n38193 = n38183 | n38192 ;
  assign n38194 = n36784 & n36792 ;
  assign n38195 = n37818 | n38194 ;
  assign n38196 = ~x1150 & n38195 ;
  assign n38197 = n38193 & n38196 ;
  assign n38198 = n36857 & n38185 ;
  assign n38199 = ~n36871 & n37200 ;
  assign n38200 = ~x212 & n36328 ;
  assign n38201 = x219 | n38200 ;
  assign n38202 = n37149 | n38201 ;
  assign n38203 = n38199 | n38202 ;
  assign n38204 = ~n38198 & n38203 ;
  assign n38205 = n37861 & ~n38204 ;
  assign n38206 = x214 & ~n36809 ;
  assign n38207 = ~n36863 & n38206 ;
  assign n38208 = ( x212 & n8894 ) | ( x212 & n36365 ) | ( n8894 & n36365 ) ;
  assign n38209 = ~n38207 & n38208 ;
  assign n38210 = n36818 | n38209 ;
  assign n38211 = ~n38198 & n38210 ;
  assign n38212 = n37818 | n38211 ;
  assign n38213 = x1150 & n38212 ;
  assign n38214 = ~n38205 & n38213 ;
  assign n38215 = n38197 | n38214 ;
  assign n38216 = x1148 & n38215 ;
  assign n38217 = x1150 & n36802 ;
  assign n38218 = x219 | n36839 ;
  assign n38219 = n37260 & n38218 ;
  assign n38220 = ~n38185 & n38219 ;
  assign n38221 = n37895 & n38185 ;
  assign n38222 = ( n37816 & n38220 ) | ( n37816 & ~n38221 ) | ( n38220 & ~n38221 ) ;
  assign n38223 = n38217 | n38222 ;
  assign n38224 = x1150 & n36372 ;
  assign n38225 = x299 & n36728 ;
  assign n38226 = x219 | n38225 ;
  assign n38227 = n37915 | n38226 ;
  assign n38228 = n38224 | n38227 ;
  assign n38229 = n37895 & ~n38228 ;
  assign n38230 = x1148 | n38229 ;
  assign n38231 = n38223 & ~n38230 ;
  assign n38232 = n38216 | n38231 ;
  assign n38233 = ~x1149 & n38232 ;
  assign n38234 = n36839 & n36909 ;
  assign n38235 = n36743 | n38234 ;
  assign n38236 = n36762 | n38235 ;
  assign n38237 = ~x1146 & n36763 ;
  assign n38238 = ~n36720 & n36748 ;
  assign n38239 = n36764 & ~n38238 ;
  assign n38240 = n38237 | n38239 ;
  assign n38241 = n38236 & ~n38240 ;
  assign n38242 = n37895 & ~n38241 ;
  assign n38243 = n36745 & ~n37148 ;
  assign n38244 = x219 | n38243 ;
  assign n38245 = ~n38239 & n38244 ;
  assign n38246 = x1146 | n36743 ;
  assign n38247 = n38245 & n38246 ;
  assign n38248 = n37816 | n38247 ;
  assign n38249 = ~x1150 & n38248 ;
  assign n38250 = ~n38242 & n38249 ;
  assign n38251 = x214 | n37312 ;
  assign n38252 = n36710 & n38251 ;
  assign n38253 = x219 | n38252 ;
  assign n38254 = n36698 & n37312 ;
  assign n38255 = ~x212 & n38254 ;
  assign n38256 = n38253 | n38255 ;
  assign n38257 = ~x299 & n36403 ;
  assign n38258 = n36700 | n36859 ;
  assign n38259 = n38257 | n38258 ;
  assign n38260 = n38256 | n38259 ;
  assign n38261 = n36891 & n38185 ;
  assign n38262 = n38253 | n38254 ;
  assign n38263 = ~n38261 & n38262 ;
  assign n38264 = n38260 & n38263 ;
  assign n38265 = n36696 | n38264 ;
  assign n38266 = n36699 & ~n36709 ;
  assign n38267 = x219 | n38266 ;
  assign n38268 = n37316 | n38267 ;
  assign n38269 = ~n36890 & n38268 ;
  assign n38270 = n38265 & n38269 ;
  assign n38271 = n37816 | n38270 ;
  assign n38272 = n37895 & ~n38264 ;
  assign n38273 = x1150 & ~n38272 ;
  assign n38274 = n38271 & n38273 ;
  assign n38275 = x1148 | n38274 ;
  assign n38276 = n38250 | n38275 ;
  assign n38277 = ~n36732 & n38185 ;
  assign n38278 = n36773 & n36789 ;
  assign n38279 = n36777 | n38278 ;
  assign n38280 = n37818 & n38279 ;
  assign n38281 = ~n36447 & n37848 ;
  assign n38282 = n36788 & ~n38281 ;
  assign n38283 = n36791 | n38282 ;
  assign n38284 = n38280 | n38283 ;
  assign n38285 = ~n38277 & n38284 ;
  assign n38286 = n38183 | n38285 ;
  assign n38287 = ~x1150 & n38286 ;
  assign n38288 = n36915 | n38220 ;
  assign n38289 = n37818 | n38288 ;
  assign n38290 = x214 & n36908 ;
  assign n38291 = n36906 & ~n38290 ;
  assign n38292 = x219 | n36911 ;
  assign n38293 = n38291 | n38292 ;
  assign n38294 = ~n36904 & n38293 ;
  assign n38295 = x1146 & n36721 ;
  assign n38296 = n37861 & ~n38295 ;
  assign n38297 = ~n38294 & n38296 ;
  assign n38298 = x1150 & ~n38297 ;
  assign n38299 = n38289 & n38298 ;
  assign n38300 = x1148 & ~n38299 ;
  assign n38301 = ~n38287 & n38300 ;
  assign n38302 = x1149 & ~n38301 ;
  assign n38303 = n38276 & n38302 ;
  assign n38304 = n38233 | n38303 ;
  assign n38305 = ( x209 & x213 ) | ( x209 & ~n38304 ) | ( x213 & ~n38304 ) ;
  assign n38306 = ~n38182 & n38305 ;
  assign n38307 = n38166 & ~n38306 ;
  assign n38308 = x230 & ~n38307 ;
  assign n38309 = x230 | x246 ;
  assign n38310 = ~n38308 & n38309 ;
  assign n38311 = ( ~x209 & x213 ) | ( ~x209 & n37373 ) | ( x213 & n37373 ) ;
  assign n38312 = ~x1147 & n37356 ;
  assign n38313 = x1151 & ~n36739 ;
  assign n38314 = ~n36697 & n38256 ;
  assign n38315 = n38313 & ~n38314 ;
  assign n38316 = n38312 & ~n38315 ;
  assign n38317 = n36747 | n36752 ;
  assign n38318 = ~n38239 & n38317 ;
  assign n38319 = n36733 | n38318 ;
  assign n38320 = x1151 | n38319 ;
  assign n38321 = x1151 & ~n36733 ;
  assign n38322 = ~n36890 & n38262 ;
  assign n38323 = n38321 & ~n38322 ;
  assign n38324 = x1147 & ~n38323 ;
  assign n38325 = n38320 & n38324 ;
  assign n38326 = x1149 | n38325 ;
  assign n38327 = n38316 | n38326 ;
  assign n38328 = x1151 | n36469 ;
  assign n38329 = n36791 | n38278 ;
  assign n38330 = ~n37268 & n38329 ;
  assign n38331 = n36778 & ~n37268 ;
  assign n38332 = n38330 | n38331 ;
  assign n38333 = n38328 | n38332 ;
  assign n38334 = n37194 & ~n38294 ;
  assign n38335 = x1147 | n38334 ;
  assign n38336 = n38333 & ~n38335 ;
  assign n38337 = x1147 & ~n37369 ;
  assign n38338 = n36718 | n36721 ;
  assign n38339 = n37283 | n38338 ;
  assign n38340 = n38337 & n38339 ;
  assign n38341 = x1149 & ~n38340 ;
  assign n38342 = ~n38336 & n38341 ;
  assign n38343 = x1150 & ~n38342 ;
  assign n38344 = n38327 & n38343 ;
  assign n38345 = x212 & n36352 ;
  assign n38346 = n38202 | n38345 ;
  assign n38347 = ~n36826 & n38346 ;
  assign n38348 = n37140 & ~n38347 ;
  assign n38349 = x1147 & ~n38348 ;
  assign n38350 = n35110 | n36774 ;
  assign n38351 = n36783 & ~n37248 ;
  assign n38352 = n38350 & n38351 ;
  assign n38353 = x1151 | n36718 ;
  assign n38354 = n38352 | n38353 ;
  assign n38355 = n36797 | n38354 ;
  assign n38356 = n38349 & n38355 ;
  assign n38357 = n37201 | n38202 ;
  assign n38358 = ~n36857 & n38357 ;
  assign n38359 = n36469 | n38358 ;
  assign n38360 = x1151 & ~n38359 ;
  assign n38361 = n38328 | n38352 ;
  assign n38362 = ~x1147 & n38361 ;
  assign n38363 = ~n38360 & n38362 ;
  assign n38364 = x1149 & ~n38363 ;
  assign n38365 = ~n38356 & n38364 ;
  assign n38366 = ~n37340 & n38321 ;
  assign n38367 = n36731 | n37147 ;
  assign n38368 = x1147 & n38367 ;
  assign n38369 = ~n38366 & n38368 ;
  assign n38370 = n36738 & n36803 ;
  assign n38371 = x1151 | n38370 ;
  assign n38372 = ~x1147 & n38371 ;
  assign n38373 = ~n36561 & n37157 ;
  assign n38374 = n38313 & ~n38373 ;
  assign n38375 = n38372 & ~n38374 ;
  assign n38376 = x1149 | n38375 ;
  assign n38377 = n38369 | n38376 ;
  assign n38378 = ~x1150 & n38377 ;
  assign n38379 = ~n38365 & n38378 ;
  assign n38380 = n38344 | n38379 ;
  assign n38381 = x1148 & n38380 ;
  assign n38382 = x1147 & ~n37364 ;
  assign n38383 = x1151 | n36808 ;
  assign n38384 = n36797 | n38383 ;
  assign n38385 = n38382 & n38384 ;
  assign n38386 = n36821 & ~n36857 ;
  assign n38387 = n36850 | n38386 ;
  assign n38388 = x1151 & ~n38387 ;
  assign n38389 = x1151 | n36850 ;
  assign n38390 = n37232 | n38389 ;
  assign n38391 = ~x1147 & n38390 ;
  assign n38392 = ~n38388 & n38391 ;
  assign n38393 = x1150 | n38392 ;
  assign n38394 = n38385 | n38393 ;
  assign n38395 = n38330 | n38389 ;
  assign n38396 = x1151 & ~n36850 ;
  assign n38397 = ~n36915 & n38396 ;
  assign n38398 = x1147 | n38397 ;
  assign n38399 = n38395 & ~n38398 ;
  assign n38400 = n37109 & ~n37262 ;
  assign n38401 = x1147 & ~n38400 ;
  assign n38402 = n36796 | n36808 ;
  assign n38403 = x1151 | n38402 ;
  assign n38404 = n38401 & n38403 ;
  assign n38405 = x1150 & ~n38404 ;
  assign n38406 = ~n38399 & n38405 ;
  assign n38407 = n38394 & ~n38406 ;
  assign n38408 = ( x1148 & x1149 ) | ( x1148 & ~n38407 ) | ( x1149 & ~n38407 ) ;
  assign n38409 = n38268 & n38322 ;
  assign n38410 = n36474 & ~n38409 ;
  assign n38411 = n36473 | n38245 ;
  assign n38412 = x1151 | n38411 ;
  assign n38413 = x1147 & n38412 ;
  assign n38414 = ~n38410 & n38413 ;
  assign n38415 = x1151 | n36922 ;
  assign n38416 = ~x1147 & n38415 ;
  assign n38417 = x1151 & ~n36696 ;
  assign n38418 = n38416 & ~n38417 ;
  assign n38419 = x1150 & ~n38418 ;
  assign n38420 = ~n38414 & n38419 ;
  assign n38421 = n36372 | n37260 ;
  assign n38422 = ~n37338 & n38421 ;
  assign n38423 = n36474 & ~n38422 ;
  assign n38424 = n37126 | n37261 ;
  assign n38425 = x1147 & n38424 ;
  assign n38426 = ~n38423 & n38425 ;
  assign n38427 = ~x1147 & x1151 ;
  assign n38428 = n36802 & n38427 ;
  assign n38429 = x1150 | n38428 ;
  assign n38430 = n38426 | n38429 ;
  assign n38431 = ~n38420 & n38430 ;
  assign n38432 = ( ~x1148 & x1149 ) | ( ~x1148 & n38431 ) | ( x1149 & n38431 ) ;
  assign n38433 = ~n38408 & n38432 ;
  assign n38434 = n38381 | n38433 ;
  assign n38435 = ( x209 & x213 ) | ( x209 & ~n38434 ) | ( x213 & ~n38434 ) ;
  assign n38436 = ~n38311 & n38435 ;
  assign n38437 = n37126 | n38409 ;
  assign n38438 = n36808 | n38269 ;
  assign n38439 = x1151 & ~n38438 ;
  assign n38440 = x1147 | n38439 ;
  assign n38441 = n38437 & ~n38440 ;
  assign n38442 = n36723 | n38424 ;
  assign n38443 = n38401 & n38442 ;
  assign n38444 = x1150 | n38443 ;
  assign n38445 = n38441 | n38444 ;
  assign n38446 = n37147 | n38322 ;
  assign n38447 = n36705 | n36893 ;
  assign n38448 = ~n36890 & n38447 ;
  assign n38449 = n37140 & ~n38448 ;
  assign n38450 = x1147 | n38449 ;
  assign n38451 = n38446 & ~n38450 ;
  assign n38452 = n36733 | n37265 ;
  assign n38453 = x1151 | n38452 ;
  assign n38454 = n38337 & n38453 ;
  assign n38455 = x1150 & ~n38454 ;
  assign n38456 = ~n38451 & n38455 ;
  assign n38457 = n38445 & ~n38456 ;
  assign n38458 = ( x1148 & ~x1149 ) | ( x1148 & n38457 ) | ( ~x1149 & n38457 ) ;
  assign n38459 = ~n38330 & n38396 ;
  assign n38460 = x1147 & n37283 ;
  assign n38461 = ~n38459 & n38460 ;
  assign n38462 = n6785 | n37324 ;
  assign n38463 = n37327 | n38462 ;
  assign n38464 = ~n37176 & n38463 ;
  assign n38465 = n38416 & n38464 ;
  assign n38466 = x1150 | n38465 ;
  assign n38467 = n38461 | n38466 ;
  assign n38468 = n36760 & ~n36764 ;
  assign n38469 = n37194 & ~n38468 ;
  assign n38470 = n38312 & ~n38469 ;
  assign n38471 = n37194 & ~n38332 ;
  assign n38472 = n37210 | n38331 ;
  assign n38473 = x1147 & n38472 ;
  assign n38474 = ~n38471 & n38473 ;
  assign n38475 = x1150 & ~n38474 ;
  assign n38476 = ~n38470 & n38475 ;
  assign n38477 = n38467 & ~n38476 ;
  assign n38478 = ( x1148 & x1149 ) | ( x1148 & n38477 ) | ( x1149 & n38477 ) ;
  assign n38479 = n38458 & n38478 ;
  assign n38480 = x219 | n37155 ;
  assign n38481 = n37237 | n38480 ;
  assign n38482 = ~n36826 & n38481 ;
  assign n38483 = n36822 & n38482 ;
  assign n38484 = n37126 | n38483 ;
  assign n38485 = n38382 & n38484 ;
  assign n38486 = n36389 & ~n36561 ;
  assign n38487 = ~n8894 & n38486 ;
  assign n38488 = n38422 | n38487 ;
  assign n38489 = n37109 & ~n38488 ;
  assign n38490 = n37126 | n38422 ;
  assign n38491 = ~x1147 & n38490 ;
  assign n38492 = ~n38489 & n38491 ;
  assign n38493 = x1150 | n38492 ;
  assign n38494 = n38485 | n38493 ;
  assign n38495 = n36733 | n38482 ;
  assign n38496 = x1151 | n38495 ;
  assign n38497 = n38349 & n38496 ;
  assign n38498 = n37147 | n37340 ;
  assign n38499 = n37140 & ~n38486 ;
  assign n38500 = ~n37340 & n38499 ;
  assign n38501 = x1147 | n38500 ;
  assign n38502 = n38498 & ~n38501 ;
  assign n38503 = x1150 & ~n38502 ;
  assign n38504 = ~n38497 & n38503 ;
  assign n38505 = n38494 & ~n38504 ;
  assign n38506 = ( x1148 & x1149 ) | ( x1148 & ~n38505 ) | ( x1149 & ~n38505 ) ;
  assign n38507 = n36785 & ~n37248 ;
  assign n38508 = n36739 | n38507 ;
  assign n38509 = x1151 | n38508 ;
  assign n38510 = n37194 & ~n38352 ;
  assign n38511 = x1147 & ~n38510 ;
  assign n38512 = n38509 & n38511 ;
  assign n38513 = n14313 & n36468 ;
  assign n38514 = x1151 & ~n38513 ;
  assign n38515 = n38372 & ~n38514 ;
  assign n38516 = x1150 & ~n38515 ;
  assign n38517 = ~n38512 & n38516 ;
  assign n38518 = n36850 | n37232 ;
  assign n38519 = x1151 | n38186 ;
  assign n38520 = x1147 & n38519 ;
  assign n38521 = n38518 & n38520 ;
  assign n38522 = n36804 & n38427 ;
  assign n38523 = x1150 | n38522 ;
  assign n38524 = n38521 | n38523 ;
  assign n38525 = ~n38517 & n38524 ;
  assign n38526 = ( ~x1148 & x1149 ) | ( ~x1148 & n38525 ) | ( x1149 & n38525 ) ;
  assign n38527 = ~n38506 & n38526 ;
  assign n38528 = n38479 | n38527 ;
  assign n38529 = ( x209 & x213 ) | ( x209 & n38528 ) | ( x213 & n38528 ) ;
  assign n38530 = ( x209 & ~x213 ) | ( x209 & n36833 ) | ( ~x213 & n36833 ) ;
  assign n38531 = n38529 | n38530 ;
  assign n38532 = ~n38436 & n38531 ;
  assign n38533 = x230 & ~n38532 ;
  assign n38534 = x230 | x247 ;
  assign n38535 = ~n38533 & n38534 ;
  assign n38536 = x1151 & ~n38495 ;
  assign n38537 = ~x1152 & n38484 ;
  assign n38538 = ~n38536 & n38537 ;
  assign n38539 = n36827 | n38383 ;
  assign n38540 = x1152 & n38539 ;
  assign n38541 = ~n38348 & n38540 ;
  assign n38542 = x1150 & ~n38541 ;
  assign n38543 = ~n38538 & n38542 ;
  assign n38544 = x1151 & ~n38508 ;
  assign n38545 = ~x1152 & n38519 ;
  assign n38546 = ~n38544 & n38545 ;
  assign n38547 = x1152 & n38390 ;
  assign n38548 = ~n38510 & n38547 ;
  assign n38549 = n38546 | n38548 ;
  assign n38550 = ( ~x1149 & n37336 ) | ( ~x1149 & n38549 ) | ( n37336 & n38549 ) ;
  assign n38551 = ~n38543 & n38550 ;
  assign n38552 = x1152 & n38395 ;
  assign n38553 = ~n38471 & n38552 ;
  assign n38554 = n38313 & ~n38331 ;
  assign n38555 = n37284 & ~n38554 ;
  assign n38556 = x1150 | n38555 ;
  assign n38557 = n38553 | n38556 ;
  assign n38558 = x1152 & ~n37369 ;
  assign n38559 = n37262 | n38383 ;
  assign n38560 = n38558 & n38559 ;
  assign n38561 = x1151 & ~n38452 ;
  assign n38562 = ~x1152 & n38442 ;
  assign n38563 = ~n38561 & n38562 ;
  assign n38564 = n38560 | n38563 ;
  assign n38565 = ( x1149 & n37255 ) | ( x1149 & n38564 ) | ( n37255 & n38564 ) ;
  assign n38566 = n38557 & n38565 ;
  assign n38567 = x1148 & ~n38566 ;
  assign n38568 = ~n38551 & n38567 ;
  assign n38569 = ~n36765 & n38313 ;
  assign n38570 = x1152 | n38569 ;
  assign n38571 = n38415 & ~n38570 ;
  assign n38572 = x1151 | n38464 ;
  assign n38573 = x1152 & n38572 ;
  assign n38574 = ~n38469 & n38573 ;
  assign n38575 = x1150 | n38574 ;
  assign n38576 = n38571 | n38575 ;
  assign n38577 = x1152 | n38323 ;
  assign n38578 = n38437 & ~n38577 ;
  assign n38579 = x1151 | n38438 ;
  assign n38580 = x1152 & ~n38449 ;
  assign n38581 = n38579 & n38580 ;
  assign n38582 = n38578 | n38581 ;
  assign n38583 = ( x1149 & n37255 ) | ( x1149 & n38582 ) | ( n37255 & n38582 ) ;
  assign n38584 = n38576 & n38583 ;
  assign n38585 = n38383 | n38488 ;
  assign n38586 = x1152 & ~n38500 ;
  assign n38587 = n38585 & n38586 ;
  assign n38588 = ~x1152 & n38490 ;
  assign n38589 = ~n38366 & n38588 ;
  assign n38590 = x1150 & ~n38589 ;
  assign n38591 = ~n38587 & n38590 ;
  assign n38592 = x1151 | n36804 ;
  assign n38593 = x1152 & ~n38514 ;
  assign n38594 = n38592 & n38593 ;
  assign n38595 = x1151 & ~x1152 ;
  assign n38596 = n38370 & n38595 ;
  assign n38597 = n38594 | n38596 ;
  assign n38598 = ( ~x1149 & n37336 ) | ( ~x1149 & n38597 ) | ( n37336 & n38597 ) ;
  assign n38599 = ~n38591 & n38598 ;
  assign n38600 = x1148 | n38599 ;
  assign n38601 = n38584 | n38600 ;
  assign n38602 = x213 & n38601 ;
  assign n38603 = ~n38568 & n38602 ;
  assign n38604 = ~x213 & n38181 ;
  assign n38605 = x209 | n38604 ;
  assign n38606 = n38603 | n38605 ;
  assign n38607 = n36766 & n38595 ;
  assign n38608 = n36802 | n38592 ;
  assign n38609 = x1152 & n38608 ;
  assign n38610 = ~n37357 & n38609 ;
  assign n38611 = x1150 | n38610 ;
  assign n38612 = n38607 | n38611 ;
  assign n38613 = n38539 & n38558 ;
  assign n38614 = x1151 & ~n36735 ;
  assign n38615 = x1152 | n38614 ;
  assign n38616 = n37365 & ~n38615 ;
  assign n38617 = x1150 & ~n38616 ;
  assign n38618 = ~n38613 & n38617 ;
  assign n38619 = n38612 & ~n38618 ;
  assign n38620 = ( ~x209 & x213 ) | ( ~x209 & n38619 ) | ( x213 & n38619 ) ;
  assign n38621 = n38347 | n38353 ;
  assign n38622 = n38558 & n38621 ;
  assign n38623 = x1151 & ~n36732 ;
  assign n38624 = ~n38338 & n38623 ;
  assign n38625 = x1152 | n38624 ;
  assign n38626 = n38355 & ~n38625 ;
  assign n38627 = x1150 & ~n38626 ;
  assign n38628 = ~n38622 & n38627 ;
  assign n38629 = x1151 & ~n38319 ;
  assign n38630 = ~x1152 & n38367 ;
  assign n38631 = ~n38629 & n38630 ;
  assign n38632 = x1152 & n38498 ;
  assign n38633 = ~n38323 & n38632 ;
  assign n38634 = x1150 | n38633 ;
  assign n38635 = n38631 | n38634 ;
  assign n38636 = x1148 & n38635 ;
  assign n38637 = ~n38628 & n38636 ;
  assign n38638 = n38371 & ~n38570 ;
  assign n38639 = n37210 | n38373 ;
  assign n38640 = x1152 & n38639 ;
  assign n38641 = ~n38315 & n38640 ;
  assign n38642 = x1150 | n38641 ;
  assign n38643 = n38638 | n38642 ;
  assign n38644 = ~x1152 & n38361 ;
  assign n38645 = ~n38471 & n38644 ;
  assign n38646 = x1151 | n38359 ;
  assign n38647 = x1152 & ~n38334 ;
  assign n38648 = n38646 & n38647 ;
  assign n38649 = x1150 & ~n38648 ;
  assign n38650 = ~n38645 & n38649 ;
  assign n38651 = x1148 | n38650 ;
  assign n38652 = n38643 & ~n38651 ;
  assign n38653 = n38637 | n38652 ;
  assign n38654 = x1149 & n38653 ;
  assign n38655 = ~n38400 & n38540 ;
  assign n38656 = x1151 & ~n38402 ;
  assign n38657 = ~x1152 & n38384 ;
  assign n38658 = ~n38656 & n38657 ;
  assign n38659 = n38655 | n38658 ;
  assign n38660 = x1150 & n38659 ;
  assign n38661 = ~n38410 & n38490 ;
  assign n38662 = ( x1150 & x1152 ) | ( x1150 & ~n38661 ) | ( x1152 & ~n38661 ) ;
  assign n38663 = x1151 & ~n38411 ;
  assign n38664 = n38424 & ~n38663 ;
  assign n38665 = ( ~x1150 & x1152 ) | ( ~x1150 & n38664 ) | ( x1152 & n38664 ) ;
  assign n38666 = ~n38662 & n38665 ;
  assign n38667 = x1148 & ~n38666 ;
  assign n38668 = ~n38660 & n38667 ;
  assign n38669 = x1151 | n38387 ;
  assign n38670 = x1152 & ~n38397 ;
  assign n38671 = n38669 & n38670 ;
  assign n38672 = ~x1152 & n38390 ;
  assign n38673 = ~n38459 & n38672 ;
  assign n38674 = x1150 & ~n38673 ;
  assign n38675 = ~n38671 & n38674 ;
  assign n38676 = x1151 | n36802 ;
  assign n38677 = x1152 & ~n38417 ;
  assign n38678 = n38676 & n38677 ;
  assign n38679 = n36922 & n38595 ;
  assign n38680 = x1150 | n38679 ;
  assign n38681 = n38678 | n38680 ;
  assign n38682 = ~n38675 & n38681 ;
  assign n38683 = x1148 | n38682 ;
  assign n38684 = ~x1149 & n38683 ;
  assign n38685 = ~n38668 & n38684 ;
  assign n38686 = n38654 | n38685 ;
  assign n38687 = ( x209 & x213 ) | ( x209 & ~n38686 ) | ( x213 & ~n38686 ) ;
  assign n38688 = ~n38620 & n38687 ;
  assign n38689 = n38606 & ~n38688 ;
  assign n38690 = x230 & ~n38689 ;
  assign n38691 = x230 | x248 ;
  assign n38692 = ~n38690 & n38691 ;
  assign n38693 = x213 & n35809 ;
  assign n38694 = x209 & ~n38693 ;
  assign n38695 = x207 & ~n35327 ;
  assign n38696 = ~n35711 & n38695 ;
  assign n38697 = x208 & ~n38696 ;
  assign n38698 = ( x207 & n35896 ) | ( x207 & n38697 ) | ( n35896 & n38697 ) ;
  assign n38699 = x207 & ~n38697 ;
  assign n38700 = ( n35317 & n38698 ) | ( n35317 & ~n38699 ) | ( n38698 & ~n38699 ) ;
  assign n38701 = x211 | n38700 ;
  assign n38702 = ~n35735 & n38701 ;
  assign n38703 = n35100 & n38702 ;
  assign n38704 = x219 & ~n35732 ;
  assign n38705 = ~n38703 & n38704 ;
  assign n38706 = n6785 | n38705 ;
  assign n38707 = ~n8652 & n35713 ;
  assign n38708 = x211 & n38700 ;
  assign n38709 = x214 & n38708 ;
  assign n38710 = n38707 | n38709 ;
  assign n38711 = ~x212 & n38710 ;
  assign n38712 = x219 | n38711 ;
  assign n38713 = x214 & ~n38700 ;
  assign n38714 = ~x211 & n35713 ;
  assign n38715 = n38708 | n38714 ;
  assign n38716 = ( x212 & n8894 ) | ( x212 & n38715 ) | ( n8894 & n38715 ) ;
  assign n38717 = ~n38713 & n38716 ;
  assign n38718 = n38712 | n38717 ;
  assign n38719 = ~n38706 & n38718 ;
  assign n38720 = n38321 & ~n38719 ;
  assign n38721 = ( x212 & x219 ) | ( x212 & n38710 ) | ( x219 & n38710 ) ;
  assign n38722 = ( ~x212 & x219 ) | ( ~x212 & n35713 ) | ( x219 & n35713 ) ;
  assign n38723 = n38721 | n38722 ;
  assign n38724 = ~n38706 & n38723 ;
  assign n38725 = n37126 | n38724 ;
  assign n38726 = ~x1152 & n38725 ;
  assign n38727 = ~n38720 & n38726 ;
  assign n38728 = ~x211 & n35624 ;
  assign n38729 = n35775 | n38728 ;
  assign n38730 = ( ~x212 & x214 ) | ( ~x212 & n38729 ) | ( x214 & n38729 ) ;
  assign n38731 = ( x212 & x214 ) | ( x212 & ~n35747 ) | ( x214 & ~n35747 ) ;
  assign n38732 = ~n38730 & n38731 ;
  assign n38733 = x214 & ~n35747 ;
  assign n38734 = n35753 & ~n38733 ;
  assign n38735 = ( x212 & ~n38732 ) | ( x212 & n38734 ) | ( ~n38732 & n38734 ) ;
  assign n38736 = x219 | n38735 ;
  assign n38737 = ~n35752 & n38736 ;
  assign n38738 = n38383 | n38737 ;
  assign n38739 = x214 & ~n35744 ;
  assign n38740 = n35753 & ~n38739 ;
  assign n38741 = x219 | n38740 ;
  assign n38742 = x212 & n35744 ;
  assign n38743 = n38741 | n38742 ;
  assign n38744 = ~n35752 & n38743 ;
  assign n38745 = n37140 & ~n38744 ;
  assign n38746 = x1152 & ~n38745 ;
  assign n38747 = n38738 & n38746 ;
  assign n38748 = n38727 | n38747 ;
  assign n38749 = ( x213 & x1150 ) | ( x213 & ~n38748 ) | ( x1150 & ~n38748 ) ;
  assign n38750 = x214 & ~n38702 ;
  assign n38751 = n38716 & ~n38750 ;
  assign n38752 = n38712 | n38751 ;
  assign n38753 = ~n35803 & n38752 ;
  assign n38754 = n38313 & ~n38753 ;
  assign n38755 = ~n35578 & n35713 ;
  assign n38756 = n38595 | n38755 ;
  assign n38757 = ~n38754 & n38756 ;
  assign n38758 = ( x212 & n8894 ) | ( x212 & n35744 ) | ( n8894 & n35744 ) ;
  assign n38759 = ~n38733 & n38758 ;
  assign n38760 = n38741 | n38759 ;
  assign n38761 = n6785 | n35749 ;
  assign n38762 = n38760 & ~n38761 ;
  assign n38763 = n37194 & ~n38762 ;
  assign n38764 = ( ~n6785 & n35624 ) | ( ~n6785 & n36526 ) | ( n35624 & n36526 ) ;
  assign n38765 = ( n6785 & ~n35747 ) | ( n6785 & n36526 ) | ( ~n35747 & n36526 ) ;
  assign n38766 = n38764 & ~n38765 ;
  assign n38767 = n38389 | n38766 ;
  assign n38768 = x1152 & n38767 ;
  assign n38769 = ~n38763 & n38768 ;
  assign n38770 = n38757 | n38769 ;
  assign n38771 = ( ~x213 & x1150 ) | ( ~x213 & n38770 ) | ( x1150 & n38770 ) ;
  assign n38772 = ~n38749 & n38771 ;
  assign n38773 = n38694 & ~n38772 ;
  assign n38774 = x299 & ~n35509 ;
  assign n38775 = n36783 & ~n38774 ;
  assign n38776 = ~x214 & n38775 ;
  assign n38777 = n36544 | n36782 ;
  assign n38778 = ~n37230 & n38777 ;
  assign n38779 = ( x212 & n35109 ) | ( x212 & ~n38778 ) | ( n35109 & ~n38778 ) ;
  assign n38780 = ~n38776 & n38779 ;
  assign n38781 = ~x212 & n36451 ;
  assign n38782 = n38775 & n38781 ;
  assign n38783 = ( x212 & ~n38780 ) | ( x212 & n38782 ) | ( ~n38780 & n38782 ) ;
  assign n38784 = x219 | n38783 ;
  assign n38785 = n4832 | n37247 ;
  assign n38786 = n38784 & ~n38785 ;
  assign n38787 = n4832 & n35577 ;
  assign n38788 = x57 | x1151 ;
  assign n38789 = n38787 | n38788 ;
  assign n38790 = n38786 | n38789 ;
  assign n38791 = x57 & ~n35577 ;
  assign n38792 = n37269 & ~n38774 ;
  assign n38793 = x214 & ~n38792 ;
  assign n38794 = n38781 & ~n38793 ;
  assign n38795 = x214 | n38792 ;
  assign n38796 = ~n36428 & n36581 ;
  assign n38797 = x212 & ~n38796 ;
  assign n38798 = n38795 & n38797 ;
  assign n38799 = x219 | n38798 ;
  assign n38800 = n38794 | n38799 ;
  assign n38801 = n4832 | n36458 ;
  assign n38802 = n38800 & ~n38801 ;
  assign n38803 = ~x57 & x1151 ;
  assign n38804 = ~n38787 & n38803 ;
  assign n38805 = ~n38802 & n38804 ;
  assign n38806 = n38791 | n38805 ;
  assign n38807 = n38790 & ~n38806 ;
  assign n38808 = x1152 | n38807 ;
  assign n38809 = n36811 & ~n37223 ;
  assign n38810 = n36352 & ~n38774 ;
  assign n38811 = x214 | n38810 ;
  assign n38812 = x212 & n38811 ;
  assign n38813 = ~n38809 & n38812 ;
  assign n38814 = n37149 & ~n38774 ;
  assign n38815 = n38201 | n38814 ;
  assign n38816 = n38813 | n38815 ;
  assign n38817 = ~x1151 & n38816 ;
  assign n38818 = ~n36826 & n38817 ;
  assign n38819 = x299 & n35509 ;
  assign n38820 = ~n8894 & n38819 ;
  assign n38821 = n35507 | n38820 ;
  assign n38822 = n36719 & n38821 ;
  assign n38823 = n37256 | n38822 ;
  assign n38824 = n36794 & n36904 ;
  assign n38825 = x1151 & ~n38824 ;
  assign n38826 = n38823 & n38825 ;
  assign n38827 = n35514 & ~n38826 ;
  assign n38828 = ~n38818 & n38827 ;
  assign n38829 = x1150 & ~n38828 ;
  assign n38830 = n38808 & n38829 ;
  assign n38831 = x211 & n37325 ;
  assign n38832 = ~n35357 & n36754 ;
  assign n38833 = n35442 & ~n38832 ;
  assign n38834 = ~n38831 & n38833 ;
  assign n38835 = n8894 & ~n37326 ;
  assign n38836 = n35804 | n36743 ;
  assign n38837 = ~n38835 & n38836 ;
  assign n38838 = ~n38834 & n38837 ;
  assign n38839 = x219 | n38838 ;
  assign n38840 = x1151 & ~n36764 ;
  assign n38841 = n38839 & n38840 ;
  assign n38842 = n36428 | n38820 ;
  assign n38843 = n35576 & ~n36385 ;
  assign n38844 = n38842 & n38843 ;
  assign n38845 = n35579 | n38844 ;
  assign n38846 = n38841 | n38845 ;
  assign n38847 = n36698 | n38819 ;
  assign n38848 = x212 & n38847 ;
  assign n38849 = ~n37304 & n38848 ;
  assign n38850 = ~x212 & n36426 ;
  assign n38851 = x219 | n38850 ;
  assign n38852 = n38814 | n38851 ;
  assign n38853 = n38849 | n38852 ;
  assign n38854 = n36362 & ~n36889 ;
  assign n38855 = n38853 & n38854 ;
  assign n38856 = ~x1151 & n38422 ;
  assign n38857 = n35514 & ~n38844 ;
  assign n38858 = ~n38856 & n38857 ;
  assign n38859 = ~n38855 & n38858 ;
  assign n38860 = x1150 | n38859 ;
  assign n38861 = n38846 & ~n38860 ;
  assign n38862 = n38830 | n38861 ;
  assign n38863 = ( x209 & x213 ) | ( x209 & n38862 ) | ( x213 & n38862 ) ;
  assign n38864 = ( x209 & ~x213 ) | ( x209 & n38619 ) | ( ~x213 & n38619 ) ;
  assign n38865 = n38863 | n38864 ;
  assign n38866 = ~n38773 & n38865 ;
  assign n38867 = x230 & ~n38866 ;
  assign n38868 = x230 | x249 ;
  assign n38869 = ~n38867 & n38868 ;
  assign n38870 = ~n2041 & n9644 ;
  assign n38871 = n4811 | n38870 ;
  assign n38872 = ~x75 & n38871 ;
  assign n38873 = ~n5768 & n7196 ;
  assign n38874 = n38872 | n38873 ;
  assign n38875 = x87 | x250 ;
  assign n38876 = n7113 | n38875 ;
  assign n38877 = n38874 & ~n38876 ;
  assign n38878 = x897 & ~n8980 ;
  assign n38879 = ~x476 & n9578 ;
  assign n38880 = n38878 | n38879 ;
  assign n38881 = ( x199 & x200 ) | ( x199 & x1039 ) | ( x200 & x1039 ) ;
  assign n38882 = ( x199 & ~x200 ) | ( x199 & x1053 ) | ( ~x200 & x1053 ) ;
  assign n38883 = n38881 | n38882 ;
  assign n38884 = n38880 & n38883 ;
  assign n38885 = x251 & ~n38880 ;
  assign n38886 = n38884 | n38885 ;
  assign n38887 = x979 | x984 ;
  assign n38888 = x1001 & ~n38887 ;
  assign n38889 = n4724 & n38888 ;
  assign n38890 = n4798 & n38889 ;
  assign n38891 = ~n4981 & n38890 ;
  assign n38892 = x252 | n38891 ;
  assign n38893 = x1092 & ~x1093 ;
  assign n38894 = n38892 & n38893 ;
  assign n38895 = n4997 | n38894 ;
  assign n38896 = n4996 & n38894 ;
  assign n38897 = n38895 & ~n38896 ;
  assign n38898 = ~n4751 & n38897 ;
  assign n38899 = n4751 & n9683 ;
  assign n38900 = n38898 | n38899 ;
  assign n38901 = ( ~x299 & n4721 ) | ( ~x299 & n38900 ) | ( n4721 & n38900 ) ;
  assign n38902 = ~n4714 & n9683 ;
  assign n38903 = n4714 & n38897 ;
  assign n38904 = n38902 | n38903 ;
  assign n38905 = ( x299 & n4721 ) | ( x299 & ~n38904 ) | ( n4721 & ~n38904 ) ;
  assign n38906 = ~n38901 & n38905 ;
  assign n38907 = n9139 & ~n38906 ;
  assign n38908 = ( x299 & n4764 ) | ( x299 & n38900 ) | ( n4764 & n38900 ) ;
  assign n38909 = ( x299 & ~n4764 ) | ( x299 & n38904 ) | ( ~n4764 & n38904 ) ;
  assign n38910 = n38908 | n38909 ;
  assign n38911 = n38907 & n38910 ;
  assign n38912 = ~n9139 & n9683 ;
  assign n38913 = n7103 & ~n38912 ;
  assign n38914 = ~n38911 & n38913 ;
  assign n38915 = n9138 & n38889 ;
  assign n38916 = ~n19157 & n38915 ;
  assign n38917 = n4744 & n38916 ;
  assign n38918 = n35075 & n38917 ;
  assign n38919 = ~n4981 & n38918 ;
  assign n38920 = x252 | n38919 ;
  assign n38921 = ~x57 & x1092 ;
  assign n38922 = n38920 & n38921 ;
  assign n38923 = x57 & n9682 ;
  assign n38924 = n7103 | n38923 ;
  assign n38925 = n38922 | n38924 ;
  assign n38926 = ~n38914 & n38925 ;
  assign n38927 = n11103 | n35191 ;
  assign n38928 = n35291 & ~n38927 ;
  assign n38929 = ~n6785 & n38928 ;
  assign n38930 = x219 & n36716 ;
  assign n38931 = n38929 | n38930 ;
  assign n38932 = x1153 & n38931 ;
  assign n38933 = x1151 | n38932 ;
  assign n38934 = ~n8895 & n35273 ;
  assign n38935 = x211 & n35232 ;
  assign n38936 = n38934 | n38935 ;
  assign n38937 = n35225 | n35238 ;
  assign n38938 = n35201 & n38937 ;
  assign n38939 = n6785 | n38938 ;
  assign n38940 = n38936 | n38939 ;
  assign n38941 = ~n9580 & n35947 ;
  assign n38942 = x1151 & ~n38941 ;
  assign n38943 = n38940 & n38942 ;
  assign n38944 = n38933 & ~n38943 ;
  assign n38945 = x1152 | n38944 ;
  assign n38946 = n35201 & n36297 ;
  assign n38947 = x1151 | n9581 ;
  assign n38948 = n35278 | n38947 ;
  assign n38949 = n38946 | n38948 ;
  assign n38950 = n35230 & ~n36544 ;
  assign n38951 = x1153 & ~n38950 ;
  assign n38952 = n9520 & ~n35191 ;
  assign n38953 = x1151 & n38952 ;
  assign n38954 = ~n38951 & n38953 ;
  assign n38955 = n6785 | n38954 ;
  assign n38956 = n38949 & ~n38955 ;
  assign n38957 = ( x1151 & n8895 ) | ( x1151 & n35947 ) | ( n8895 & n35947 ) ;
  assign n38958 = n35947 & n38957 ;
  assign n38959 = x1152 & ~n38958 ;
  assign n38960 = ~n38956 & n38959 ;
  assign n38961 = n38945 & ~n38960 ;
  assign n38962 = x230 & ~n38961 ;
  assign n38963 = n37497 & ~n37511 ;
  assign n38964 = ~x211 & n37491 ;
  assign n38965 = n38963 & ~n38964 ;
  assign n38966 = n37490 & n37531 ;
  assign n38967 = n38965 & n38966 ;
  assign n38968 = x1153 & ~n38967 ;
  assign n38969 = x1153 | n37623 ;
  assign n38970 = x219 & n38969 ;
  assign n38971 = ~n38968 & n38970 ;
  assign n38972 = n37492 & n37542 ;
  assign n38973 = x1153 & ~n38972 ;
  assign n38974 = x1153 | n37564 ;
  assign n38975 = ~x219 & n38974 ;
  assign n38976 = ~n38973 & n38975 ;
  assign n38977 = x253 & ~n38976 ;
  assign n38978 = ~n38971 & n38977 ;
  assign n38979 = n37502 & n37623 ;
  assign n38980 = ~x211 & n38979 ;
  assign n38981 = n37504 | n38980 ;
  assign n38982 = x1153 & n38981 ;
  assign n38983 = n37618 | n38982 ;
  assign n38984 = x219 & ~n38983 ;
  assign n38985 = x1153 & n37512 ;
  assign n38986 = ~x1153 & n37562 ;
  assign n38987 = x219 | n38986 ;
  assign n38988 = n38985 | n38987 ;
  assign n38989 = ~x253 & n38988 ;
  assign n38990 = ~n38984 & n38989 ;
  assign n38991 = n38978 | n38990 ;
  assign n38992 = ~n6785 & n38991 ;
  assign n38993 = ~x219 & n37484 ;
  assign n38994 = x211 | n37482 ;
  assign n38995 = n38993 & n38994 ;
  assign n38996 = x219 | n38995 ;
  assign n38997 = n6785 & ~n38996 ;
  assign n38998 = n37473 & n38997 ;
  assign n38999 = x1151 & ~n38998 ;
  assign n39000 = x219 & x1091 ;
  assign n39001 = ~n35183 & n39000 ;
  assign n39002 = n37500 | n39001 ;
  assign n39003 = n38993 | n39002 ;
  assign n39004 = ( x253 & ~n6785 ) | ( x253 & n39003 ) | ( ~n6785 & n39003 ) ;
  assign n39005 = ~x211 & n37473 ;
  assign n39006 = x211 & n37500 ;
  assign n39007 = x219 & ~n39006 ;
  assign n39008 = ~n39005 & n39007 ;
  assign n39009 = x219 | n37482 ;
  assign n39010 = ~n39001 & n39009 ;
  assign n39011 = ~n39008 & n39010 ;
  assign n39012 = ( x253 & n6785 ) | ( x253 & n39011 ) | ( n6785 & n39011 ) ;
  assign n39013 = ~n39004 & n39012 ;
  assign n39014 = n38999 & ~n39013 ;
  assign n39015 = ~n38992 & n39014 ;
  assign n39016 = n37492 | n38980 ;
  assign n39017 = n38993 & n39016 ;
  assign n39018 = ~n37511 & n37519 ;
  assign n39019 = x1153 | n39018 ;
  assign n39020 = ~n37520 & n39019 ;
  assign n39021 = n39017 & ~n39020 ;
  assign n39022 = x219 & n37595 ;
  assign n39023 = ~n37611 & n38968 ;
  assign n39024 = n39022 & ~n39023 ;
  assign n39025 = n39021 | n39024 ;
  assign n39026 = ( x253 & n6785 ) | ( x253 & n39025 ) | ( n6785 & n39025 ) ;
  assign n39027 = ( x219 & ~n37497 ) | ( x219 & n38984 ) | ( ~n37497 & n38984 ) ;
  assign n39028 = n37503 & n38965 ;
  assign n39029 = n39019 & n39028 ;
  assign n39030 = ( x219 & ~n38984 ) | ( x219 & n39029 ) | ( ~n38984 & n39029 ) ;
  assign n39031 = ~n39027 & n39030 ;
  assign n39032 = ( x253 & ~n6785 ) | ( x253 & n39031 ) | ( ~n6785 & n39031 ) ;
  assign n39033 = ~n39026 & n39032 ;
  assign n39034 = x1151 | n39033 ;
  assign n39035 = ~n39015 & n39034 ;
  assign n39036 = n39005 | n39009 ;
  assign n39037 = n38993 & n39036 ;
  assign n39038 = x219 & n37473 ;
  assign n39039 = n6785 & ~n39038 ;
  assign n39040 = ~n39037 & n39039 ;
  assign n39041 = n37473 & n39040 ;
  assign n39042 = n39013 | n39041 ;
  assign n39043 = n39035 | n39042 ;
  assign n39044 = x1152 & n39043 ;
  assign n39045 = x1153 & ~n37542 ;
  assign n39046 = n38965 & n38993 ;
  assign n39047 = ~n39045 & n39046 ;
  assign n39048 = n37597 | n38967 ;
  assign n39049 = x1153 & ~n39048 ;
  assign n39050 = x1153 | n37631 ;
  assign n39051 = x219 & n39050 ;
  assign n39052 = ~n39049 & n39051 ;
  assign n39053 = n39047 | n39052 ;
  assign n39054 = ( x253 & n6785 ) | ( x253 & n39053 ) | ( n6785 & n39053 ) ;
  assign n39055 = x219 & n38983 ;
  assign n39056 = n38988 & n39017 ;
  assign n39057 = n39055 | n39056 ;
  assign n39058 = n37502 & n39057 ;
  assign n39059 = ( x253 & ~n6785 ) | ( x253 & n39058 ) | ( ~n6785 & n39058 ) ;
  assign n39060 = ~n39054 & n39059 ;
  assign n39061 = n39014 & ~n39060 ;
  assign n39062 = n37489 & n39055 ;
  assign n39063 = x1153 | n37534 ;
  assign n39064 = n37502 & n39063 ;
  assign n39065 = ~x219 & n37564 ;
  assign n39066 = n39064 & n39065 ;
  assign n39067 = x253 | n39066 ;
  assign n39068 = n39062 | n39067 ;
  assign n39069 = n37611 | n38967 ;
  assign n39070 = x1091 | n37618 ;
  assign n39071 = ~x1153 & n39070 ;
  assign n39072 = ~x219 & n39018 ;
  assign n39073 = n39071 | n39072 ;
  assign n39074 = n39069 | n39073 ;
  assign n39075 = x253 & n39074 ;
  assign n39076 = n6785 | n39075 ;
  assign n39077 = n39068 & ~n39076 ;
  assign n39078 = x1151 | n39013 ;
  assign n39079 = n39077 | n39078 ;
  assign n39080 = ~x1152 & n39079 ;
  assign n39081 = ~n39061 & n39080 ;
  assign n39082 = n39044 | n39081 ;
  assign n39083 = n37728 & n39082 ;
  assign n39084 = x253 | x1091 ;
  assign n39085 = n6785 & n39084 ;
  assign n39086 = x211 & x1091 ;
  assign n39087 = x1091 & ~x1153 ;
  assign n39088 = x219 & n39087 ;
  assign n39089 = n39086 | n39088 ;
  assign n39090 = n39085 & ~n39089 ;
  assign n39091 = x1151 & ~n39090 ;
  assign n39092 = n11106 & ~n38951 ;
  assign n39093 = x1091 & ~n39092 ;
  assign n39094 = ( x253 & ~n6785 ) | ( x253 & n39093 ) | ( ~n6785 & n39093 ) ;
  assign n39095 = x1091 & n38936 ;
  assign n39096 = x1153 | n37662 ;
  assign n39097 = x1153 & ~n37692 ;
  assign n39098 = n35201 & ~n39097 ;
  assign n39099 = n39096 & n39098 ;
  assign n39100 = n39095 | n39099 ;
  assign n39101 = ( x253 & n6785 ) | ( x253 & n39100 ) | ( n6785 & n39100 ) ;
  assign n39102 = n39094 & ~n39101 ;
  assign n39103 = n39091 & ~n39102 ;
  assign n39104 = ~n39001 & n39085 ;
  assign n39105 = x219 & n39104 ;
  assign n39106 = x1091 & x1153 ;
  assign n39107 = n38929 & n39106 ;
  assign n39108 = x253 & ~x1091 ;
  assign n39109 = x1151 | n39108 ;
  assign n39110 = n39107 | n39109 ;
  assign n39111 = n39105 | n39110 ;
  assign n39112 = ~n39103 & n39111 ;
  assign n39113 = x1152 | n39112 ;
  assign n39114 = x1153 | n37698 ;
  assign n39115 = ~n35215 & n37658 ;
  assign n39116 = x1153 & ~n39115 ;
  assign n39117 = n35201 & ~n39116 ;
  assign n39118 = n39114 & n39117 ;
  assign n39119 = n9580 & n37658 ;
  assign n39120 = ~n35278 & n39119 ;
  assign n39121 = x253 & ~n39120 ;
  assign n39122 = ~n39118 & n39121 ;
  assign n39123 = x1091 & n35278 ;
  assign n39124 = x211 & ~n37711 ;
  assign n39125 = ~n39123 & n39124 ;
  assign n39126 = x1091 & n36297 ;
  assign n39127 = x1091 & n35238 ;
  assign n39128 = ~n35617 & n39127 ;
  assign n39129 = n35201 & ~n39128 ;
  assign n39130 = ~n39126 & n39129 ;
  assign n39131 = x253 | n39130 ;
  assign n39132 = n39125 | n39131 ;
  assign n39133 = ~n39122 & n39132 ;
  assign n39134 = n9580 | n35201 ;
  assign n39135 = n39108 | n39134 ;
  assign n39136 = n39123 | n39135 ;
  assign n39137 = ~n36385 & n39136 ;
  assign n39138 = ~n39133 & n39137 ;
  assign n39139 = n38950 & ~n39108 ;
  assign n39140 = n39087 | n39139 ;
  assign n39141 = n38952 & n39140 ;
  assign n39142 = ~n6785 & n39084 ;
  assign n39143 = ~n39141 & n39142 ;
  assign n39144 = n39104 | n39143 ;
  assign n39145 = x1151 & n39144 ;
  assign n39146 = ~x211 & x1091 ;
  assign n39147 = ~x219 & n39146 ;
  assign n39148 = n39104 & ~n39147 ;
  assign n39149 = x1152 & ~n39148 ;
  assign n39150 = ~n39145 & n39149 ;
  assign n39151 = ~n39138 & n39150 ;
  assign n39152 = n37728 | n39151 ;
  assign n39153 = n39113 & ~n39152 ;
  assign n39154 = x230 | n39153 ;
  assign n39155 = n39083 | n39154 ;
  assign n39156 = ~n38962 & n39155 ;
  assign n39157 = x1154 & n35756 ;
  assign n39158 = n35785 | n39157 ;
  assign n39159 = n9580 & n39158 ;
  assign n39160 = x299 & n35201 ;
  assign n39161 = ~n9580 & n35618 ;
  assign n39162 = n39160 | n39161 ;
  assign n39163 = n35649 & n39162 ;
  assign n39164 = n39159 | n39163 ;
  assign n39165 = ~n6785 & n39164 ;
  assign n39166 = x219 | n35508 ;
  assign n39167 = ~n35817 & n39166 ;
  assign n39168 = ( x1152 & n35578 ) | ( x1152 & n39167 ) | ( n35578 & n39167 ) ;
  assign n39169 = n39165 | n39168 ;
  assign n39170 = n35222 | n35755 ;
  assign n39171 = n35169 & n39170 ;
  assign n39172 = ~x1154 & n35706 ;
  assign n39173 = n35651 | n39172 ;
  assign n39174 = n39171 | n39173 ;
  assign n39175 = x219 & n39174 ;
  assign n39176 = ~x200 & x1154 ;
  assign n39177 = n9515 & ~n39176 ;
  assign n39178 = n35755 & ~n36544 ;
  assign n39179 = n39177 | n39178 ;
  assign n39180 = ~x219 & n39179 ;
  assign n39181 = n6785 | n39180 ;
  assign n39182 = n39175 | n39181 ;
  assign n39183 = n9580 & ~n35508 ;
  assign n39184 = n36676 & ~n39183 ;
  assign n39185 = x1152 & ~n39184 ;
  assign n39186 = n39182 & n39185 ;
  assign n39187 = n39169 & ~n39186 ;
  assign n39188 = x230 & ~n39187 ;
  assign n39189 = x211 | n35272 ;
  assign n39190 = x1153 & ~n37676 ;
  assign n39191 = x1154 | n39190 ;
  assign n39192 = n39096 & ~n39191 ;
  assign n39193 = n39189 & n39192 ;
  assign n39194 = x1091 & n35169 ;
  assign n39195 = n35230 & n39194 ;
  assign n39196 = ~n35691 & n39195 ;
  assign n39197 = n39193 | n39196 ;
  assign n39198 = ~x219 & n39197 ;
  assign n39199 = x1154 & n39146 ;
  assign n39200 = n39000 | n39199 ;
  assign n39201 = n39174 & n39200 ;
  assign n39202 = n39198 | n39201 ;
  assign n39203 = x254 & n39202 ;
  assign n39204 = x254 | x1091 ;
  assign n39205 = x1154 & ~n38950 ;
  assign n39206 = x219 & n35706 ;
  assign n39207 = ~n39205 & n39206 ;
  assign n39208 = n39180 | n39207 ;
  assign n39209 = ( x254 & n39204 ) | ( x254 & ~n39208 ) | ( n39204 & ~n39208 ) ;
  assign n39210 = ~n39203 & n39209 ;
  assign n39211 = x253 | n39210 ;
  assign n39212 = ~n6785 & n39211 ;
  assign n39213 = x1154 & n37496 ;
  assign n39214 = n38965 & n39213 ;
  assign n39215 = ~n38973 & n39214 ;
  assign n39216 = x254 & ~n39215 ;
  assign n39217 = ~n38974 & n39029 ;
  assign n39218 = ( ~x1154 & n37564 ) | ( ~x1154 & n39217 ) | ( n37564 & n39217 ) ;
  assign n39219 = n39216 & ~n39218 ;
  assign n39220 = n37503 & n37631 ;
  assign n39221 = x1154 & n39220 ;
  assign n39222 = n37562 | n39221 ;
  assign n39223 = x211 & n37491 ;
  assign n39224 = n37502 & ~n39223 ;
  assign n39225 = x1153 | n39224 ;
  assign n39226 = ~x254 & n39225 ;
  assign n39227 = n39222 & n39226 ;
  assign n39228 = n39219 | n39227 ;
  assign n39229 = ( x219 & x253 ) | ( x219 & ~n39228 ) | ( x253 & ~n39228 ) ;
  assign n39230 = x1154 & ~n38968 ;
  assign n39231 = n39048 & n39230 ;
  assign n39232 = x254 & x1154 ;
  assign n39233 = x1153 & ~n37623 ;
  assign n39234 = n39050 & ~n39233 ;
  assign n39235 = ( x254 & n39232 ) | ( x254 & ~n39234 ) | ( n39232 & ~n39234 ) ;
  assign n39236 = ~n39231 & n39235 ;
  assign n39237 = x1153 | n37551 ;
  assign n39238 = n37620 & n39237 ;
  assign n39239 = x1154 | n39238 ;
  assign n39240 = n37502 & n37618 ;
  assign n39241 = n39239 | n39240 ;
  assign n39242 = n38969 & n39220 ;
  assign n39243 = n35181 & ~n39242 ;
  assign n39244 = ~n37474 & n39243 ;
  assign n39245 = x1153 & n37504 ;
  assign n39246 = n35169 & ~n37628 ;
  assign n39247 = ~n39245 & n39246 ;
  assign n39248 = x254 | n39247 ;
  assign n39249 = n39244 | n39248 ;
  assign n39250 = n39241 & ~n39249 ;
  assign n39251 = n39236 | n39250 ;
  assign n39252 = ( x219 & ~x253 ) | ( x219 & n39251 ) | ( ~x253 & n39251 ) ;
  assign n39253 = n39229 & ~n39252 ;
  assign n39254 = n39212 & ~n39253 ;
  assign n39255 = n39036 | n39106 ;
  assign n39256 = x1091 & n35817 ;
  assign n39257 = x254 | n39256 ;
  assign n39258 = n39008 | n39257 ;
  assign n39259 = n39255 & ~n39258 ;
  assign n39260 = x211 | n37498 ;
  assign n39261 = n39038 & n39260 ;
  assign n39262 = ~x219 & n37482 ;
  assign n39263 = n39261 | n39262 ;
  assign n39264 = n9580 & n39087 ;
  assign n39265 = x254 & ~n39264 ;
  assign n39266 = ~n39256 & n39265 ;
  assign n39267 = ~n39263 & n39266 ;
  assign n39268 = x253 & ~n39267 ;
  assign n39269 = ~n39259 & n39268 ;
  assign n39270 = x1091 & ~n39167 ;
  assign n39271 = n6785 & n39204 ;
  assign n39272 = ~n39270 & n39271 ;
  assign n39273 = n6785 & n39147 ;
  assign n39274 = n39272 | n39273 ;
  assign n39275 = x253 & n6785 ;
  assign n39276 = n39274 | n39275 ;
  assign n39277 = ~n39269 & n39276 ;
  assign n39278 = x1152 & ~n39277 ;
  assign n39279 = ~n39254 & n39278 ;
  assign n39280 = n39272 | n39275 ;
  assign n39281 = n38996 & n39259 ;
  assign n39282 = ~n39037 & n39267 ;
  assign n39283 = x253 & ~n39282 ;
  assign n39284 = ~n39281 & n39283 ;
  assign n39285 = n39280 & ~n39284 ;
  assign n39286 = x1152 | n39285 ;
  assign n39287 = n37665 & n39087 ;
  assign n39288 = n39126 | n39287 ;
  assign n39289 = x211 & n39191 ;
  assign n39290 = n39288 & n39289 ;
  assign n39291 = x1091 & n35618 ;
  assign n39292 = x1154 & ~n39291 ;
  assign n39293 = n9579 & n39106 ;
  assign n39294 = x1154 | n39293 ;
  assign n39295 = ~x211 & n39294 ;
  assign n39296 = ~n39292 & n39295 ;
  assign n39297 = n39290 | n39296 ;
  assign n39298 = ~x219 & n39297 ;
  assign n39299 = x211 & n39292 ;
  assign n39300 = x1091 & n36333 ;
  assign n39301 = n35181 & ~n39300 ;
  assign n39302 = ~n39126 & n39301 ;
  assign n39303 = x219 & n39294 ;
  assign n39304 = ~n39302 & n39303 ;
  assign n39305 = ~n39299 & n39304 ;
  assign n39306 = n39298 | n39305 ;
  assign n39307 = ~x254 & n39306 ;
  assign n39308 = x1153 | n37666 ;
  assign n39309 = ~n39116 & n39308 ;
  assign n39310 = x1091 & ~x1154 ;
  assign n39311 = ~n35320 & n39310 ;
  assign n39312 = n39309 | n39311 ;
  assign n39313 = n9580 & n39312 ;
  assign n39314 = x254 & ~n39313 ;
  assign n39315 = x1091 & ~n35216 ;
  assign n39316 = n39309 | n39315 ;
  assign n39317 = ~n39134 & n39316 ;
  assign n39318 = n37714 & n39117 ;
  assign n39319 = x1154 & ~n39318 ;
  assign n39320 = ~n39317 & n39319 ;
  assign n39321 = x1091 & ~n9580 ;
  assign n39322 = ~n35649 & n39321 ;
  assign n39323 = ( x1154 & ~n39320 ) | ( x1154 & n39322 ) | ( ~n39320 & n39322 ) ;
  assign n39324 = n39314 & ~n39323 ;
  assign n39325 = n39307 | n39324 ;
  assign n39326 = ( x253 & ~n6785 ) | ( x253 & n39325 ) | ( ~n6785 & n39325 ) ;
  assign n39327 = x1154 | n37641 ;
  assign n39328 = ~x1154 & n39327 ;
  assign n39329 = ~x1153 & n37531 ;
  assign n39330 = n38966 | n39329 ;
  assign n39331 = n39328 | n39330 ;
  assign n39332 = n35181 & ~n37611 ;
  assign n39333 = x219 & ~n39332 ;
  assign n39334 = n39331 & n39333 ;
  assign n39335 = n39016 | n39329 ;
  assign n39336 = x1154 & ~n37519 ;
  assign n39337 = x219 | n39336 ;
  assign n39338 = n39335 & ~n39337 ;
  assign n39339 = n39334 | n39338 ;
  assign n39340 = x254 & n39339 ;
  assign n39341 = n37505 & n38969 ;
  assign n39342 = n35169 & ~n39341 ;
  assign n39343 = x219 & ~n39243 ;
  assign n39344 = n39239 & n39343 ;
  assign n39345 = ~n39342 & n39344 ;
  assign n39346 = n37496 & n37562 ;
  assign n39347 = n39063 & n39346 ;
  assign n39348 = x1154 & ~n37497 ;
  assign n39349 = n37491 | n39348 ;
  assign n39350 = ~x211 & n39349 ;
  assign n39351 = x219 | n39350 ;
  assign n39352 = n37502 & n37564 ;
  assign n39353 = ~n39347 & n39352 ;
  assign n39354 = x1154 & n39353 ;
  assign n39355 = ( n39347 & ~n39351 ) | ( n39347 & n39354 ) | ( ~n39351 & n39354 ) ;
  assign n39356 = x254 | n39355 ;
  assign n39357 = n39345 | n39356 ;
  assign n39358 = ~n39340 & n39357 ;
  assign n39359 = ( x253 & n6785 ) | ( x253 & ~n39358 ) | ( n6785 & ~n39358 ) ;
  assign n39360 = n39326 & ~n39359 ;
  assign n39361 = n39286 | n39360 ;
  assign n39362 = n37728 & n39361 ;
  assign n39363 = ~n39279 & n39362 ;
  assign n39364 = ~n6785 & n39325 ;
  assign n39365 = x1152 | n39272 ;
  assign n39366 = n39364 | n39365 ;
  assign n39367 = ~n6785 & n39210 ;
  assign n39368 = x1152 & ~n39274 ;
  assign n39369 = ~n39367 & n39368 ;
  assign n39370 = n37728 | n39369 ;
  assign n39371 = n39366 & ~n39370 ;
  assign n39372 = x230 | n39371 ;
  assign n39373 = n39363 | n39372 ;
  assign n39374 = ~n39188 & n39373 ;
  assign n39375 = ~x200 & x1049 ;
  assign n39376 = x200 & x1036 ;
  assign n39377 = n39375 | n39376 ;
  assign n39378 = n38880 & ~n39377 ;
  assign n39379 = x255 | n38880 ;
  assign n39380 = ~n39378 & n39379 ;
  assign n39381 = ~x200 & x1048 ;
  assign n39382 = x200 & x1070 ;
  assign n39383 = n39381 | n39382 ;
  assign n39384 = n38880 & ~n39383 ;
  assign n39385 = x256 | n38880 ;
  assign n39386 = ~n39384 & n39385 ;
  assign n39387 = ~x200 & x1084 ;
  assign n39388 = x200 & x1065 ;
  assign n39389 = n39387 | n39388 ;
  assign n39390 = n38880 & ~n39389 ;
  assign n39391 = x257 | n38880 ;
  assign n39392 = ~n39390 & n39391 ;
  assign n39393 = ~x200 & x1072 ;
  assign n39394 = x200 & x1062 ;
  assign n39395 = n39393 | n39394 ;
  assign n39396 = n38880 & ~n39395 ;
  assign n39397 = x258 | n38880 ;
  assign n39398 = ~n39396 & n39397 ;
  assign n39399 = ~x200 & x1059 ;
  assign n39400 = x200 & x1069 ;
  assign n39401 = n39399 | n39400 ;
  assign n39402 = n38880 & ~n39401 ;
  assign n39403 = x259 | n38880 ;
  assign n39404 = ~n39402 & n39403 ;
  assign n39405 = ( x199 & x200 ) | ( x199 & x1067 ) | ( x200 & x1067 ) ;
  assign n39406 = ( x199 & ~x200 ) | ( x199 & x1044 ) | ( ~x200 & x1044 ) ;
  assign n39407 = n39405 | n39406 ;
  assign n39408 = n38880 & n39407 ;
  assign n39409 = x260 & ~n38880 ;
  assign n39410 = n39408 | n39409 ;
  assign n39411 = ( x199 & x200 ) | ( x199 & x1040 ) | ( x200 & x1040 ) ;
  assign n39412 = ( x199 & ~x200 ) | ( x199 & x1037 ) | ( ~x200 & x1037 ) ;
  assign n39413 = n39411 | n39412 ;
  assign n39414 = n38880 & n39413 ;
  assign n39415 = x261 & ~n38880 ;
  assign n39416 = n39414 | n39415 ;
  assign n39417 = x1093 & x1142 ;
  assign n39418 = x262 | x1093 ;
  assign n39419 = ~n39417 & n39418 ;
  assign n39420 = x228 | n39419 ;
  assign n39421 = ( x123 & ~x228 ) | ( x123 & x262 ) | ( ~x228 & x262 ) ;
  assign n39422 = ( x123 & x228 ) | ( x123 & x1142 ) | ( x228 & x1142 ) ;
  assign n39423 = ~n39421 & n39422 ;
  assign n39424 = n39420 & ~n39423 ;
  assign n39425 = x228 | x1093 ;
  assign n39426 = x123 & x228 ;
  assign n39427 = n39425 & ~n39426 ;
  assign n39428 = x262 | n39427 ;
  assign n39429 = ~n37344 & n39428 ;
  assign n39430 = x199 & n39427 ;
  assign n39431 = n35123 & ~n39430 ;
  assign n39432 = n39429 & ~n39431 ;
  assign n39433 = n39424 | n39432 ;
  assign n39434 = x207 | n39428 ;
  assign n39435 = ~x208 & n39434 ;
  assign n39436 = n37344 | n39435 ;
  assign n39437 = n39433 & n39436 ;
  assign n39438 = x299 & ~n39429 ;
  assign n39439 = n36401 & n39427 ;
  assign n39440 = n39424 | n39439 ;
  assign n39441 = ( x208 & n36617 ) | ( x208 & n39440 ) | ( n36617 & n39440 ) ;
  assign n39442 = ~n39438 & n39441 ;
  assign n39443 = n6785 | n39442 ;
  assign n39444 = n39437 | n39443 ;
  assign n39445 = ~n36468 & n39427 ;
  assign n39446 = n6785 & ~n39424 ;
  assign n39447 = ~n39445 & n39446 ;
  assign n39448 = n39444 & ~n39447 ;
  assign n39449 = x1154 & ~n37513 ;
  assign n39450 = ~n37567 & n39449 ;
  assign n39451 = x1156 & n39352 ;
  assign n39452 = x1154 | n37535 ;
  assign n39453 = x1155 & n39346 ;
  assign n39454 = n39452 | n39453 ;
  assign n39455 = ~n37584 & n39449 ;
  assign n39456 = x1156 | n39336 ;
  assign n39457 = n39455 | n39456 ;
  assign n39458 = ( x1156 & n39454 ) | ( x1156 & ~n39457 ) | ( n39454 & ~n39457 ) ;
  assign n39459 = n39451 | n39458 ;
  assign n39460 = ~n39450 & n39459 ;
  assign n39461 = x211 & ~n39460 ;
  assign n39462 = n37515 & n37561 ;
  assign n39463 = x1155 & n39462 ;
  assign n39464 = n39452 | n39463 ;
  assign n39465 = ~n39457 & n39464 ;
  assign n39466 = ( x1156 & n39451 ) | ( x1156 & n39464 ) | ( n39451 & n39464 ) ;
  assign n39467 = ~n39455 & n39466 ;
  assign n39468 = x211 | n39467 ;
  assign n39469 = n39465 | n39468 ;
  assign n39470 = ~x219 & n39469 ;
  assign n39471 = ~n39461 & n39470 ;
  assign n39472 = n37507 | n37619 ;
  assign n39473 = n37505 | n39348 ;
  assign n39474 = n39472 & n39473 ;
  assign n39475 = n37561 & n39474 ;
  assign n39476 = x1156 | n39475 ;
  assign n39477 = n35175 & ~n39474 ;
  assign n39478 = x219 & ~n35164 ;
  assign n39479 = x1155 | n38979 ;
  assign n39480 = x1155 & ~n39220 ;
  assign n39481 = x1154 | n39480 ;
  assign n39482 = n39479 & ~n39481 ;
  assign n39483 = x1154 & n39472 ;
  assign n39484 = n39482 | n39483 ;
  assign n39485 = ( x219 & n39478 ) | ( x219 & n39484 ) | ( n39478 & n39484 ) ;
  assign n39486 = ~n39477 & n39485 ;
  assign n39487 = n39476 & n39486 ;
  assign n39488 = x263 & ~n39487 ;
  assign n39489 = ~n39471 & n39488 ;
  assign n39490 = x1155 | n39070 ;
  assign n39491 = n37562 | n39490 ;
  assign n39492 = x1155 & ~n37492 ;
  assign n39493 = x1154 | n39492 ;
  assign n39494 = n39491 & ~n39493 ;
  assign n39495 = x1156 | n39494 ;
  assign n39496 = x1155 & ~n37564 ;
  assign n39497 = x1154 & ~n39496 ;
  assign n39498 = n38963 & n39497 ;
  assign n39499 = n39495 | n39498 ;
  assign n39500 = ~x1155 & n37531 ;
  assign n39501 = ~n37491 & n37520 ;
  assign n39502 = n39500 | n39501 ;
  assign n39503 = ~x1154 & n39502 ;
  assign n39504 = x1156 & ~n39503 ;
  assign n39505 = n37542 & n39497 ;
  assign n39506 = n39504 & ~n39505 ;
  assign n39507 = x211 & ~n39506 ;
  assign n39508 = n39499 & n39507 ;
  assign n39509 = x1155 & ~n37595 ;
  assign n39510 = x1154 | n39509 ;
  assign n39511 = n37531 & ~n39510 ;
  assign n39512 = n37523 & n39497 ;
  assign n39513 = n37494 & n39512 ;
  assign n39514 = n39511 | n39513 ;
  assign n39515 = n39504 & ~n39514 ;
  assign n39516 = n39490 & ~n39510 ;
  assign n39517 = n39512 | n39516 ;
  assign n39518 = n39495 | n39517 ;
  assign n39519 = ~x211 & n39518 ;
  assign n39520 = ~n39515 & n39519 ;
  assign n39521 = x219 | n39520 ;
  assign n39522 = n39508 | n39521 ;
  assign n39523 = x1155 & ~n37490 ;
  assign n39524 = x1154 & n37631 ;
  assign n39525 = ~n39523 & n39524 ;
  assign n39526 = n39516 | n39525 ;
  assign n39527 = ~x1156 & n39526 ;
  assign n39528 = n37496 & n39525 ;
  assign n39529 = n39511 | n39528 ;
  assign n39530 = n35175 & n39529 ;
  assign n39531 = ~x1154 & n37618 ;
  assign n39532 = n37597 | n39531 ;
  assign n39533 = ~n39523 & n39532 ;
  assign n39534 = ( x219 & n39478 ) | ( x219 & ~n39533 ) | ( n39478 & ~n39533 ) ;
  assign n39535 = ~n39530 & n39534 ;
  assign n39536 = ~n39527 & n39535 ;
  assign n39537 = x263 | n39536 ;
  assign n39538 = n39522 & ~n39537 ;
  assign n39539 = n37593 & ~n39538 ;
  assign n39540 = ~n39489 & n39539 ;
  assign n39541 = x1155 & ~n35764 ;
  assign n39542 = n37692 & ~n39541 ;
  assign n39543 = ~x1154 & n39315 ;
  assign n39544 = n39542 | n39543 ;
  assign n39545 = n37711 | n39544 ;
  assign n39546 = n35175 & n39545 ;
  assign n39547 = ~x1154 & n35336 ;
  assign n39548 = x1091 & n35164 ;
  assign n39549 = ~n35239 & n35650 ;
  assign n39550 = ( ~x1154 & n39548 ) | ( ~x1154 & n39549 ) | ( n39548 & n39549 ) ;
  assign n39551 = ~n39547 & n39550 ;
  assign n39552 = n37662 | n39310 ;
  assign n39553 = x1156 | n35240 ;
  assign n39554 = n39552 & ~n39553 ;
  assign n39555 = x219 & ~n39554 ;
  assign n39556 = ~n39551 & n39555 ;
  assign n39557 = ~n39546 & n39556 ;
  assign n39558 = ~x211 & n39544 ;
  assign n39559 = ~n35230 & n35660 ;
  assign n39560 = n39086 & ~n39559 ;
  assign n39561 = ~n35340 & n39560 ;
  assign n39562 = n39558 | n39561 ;
  assign n39563 = ( x219 & x1156 ) | ( x219 & n39562 ) | ( x1156 & n39562 ) ;
  assign n39564 = ~n35340 & n39552 ;
  assign n39565 = x211 & n39564 ;
  assign n39566 = n35240 | n35632 ;
  assign n39567 = n39146 & ~n39566 ;
  assign n39568 = n39565 | n39567 ;
  assign n39569 = ( x219 & ~x1156 ) | ( x219 & n39568 ) | ( ~x1156 & n39568 ) ;
  assign n39570 = n39563 | n39569 ;
  assign n39571 = ~n39557 & n39570 ;
  assign n39572 = x263 | n39571 ;
  assign n39573 = n35310 & n39547 ;
  assign n39574 = n35230 & ~n35277 ;
  assign n39575 = x1154 & ~n39574 ;
  assign n39576 = x1156 & ~n39575 ;
  assign n39577 = ~n39573 & n39576 ;
  assign n39578 = ( x211 & n35175 ) | ( x211 & ~n39564 ) | ( n35175 & ~n39564 ) ;
  assign n39579 = ~n39577 & n39578 ;
  assign n39580 = ~n35245 & n36128 ;
  assign n39581 = n35632 | n39580 ;
  assign n39582 = ~x211 & n39581 ;
  assign n39583 = x219 | n39582 ;
  assign n39584 = n39579 | n39583 ;
  assign n39585 = x1154 & ~n35242 ;
  assign n39586 = x1156 & ~n39585 ;
  assign n39587 = x299 | n39586 ;
  assign n39588 = n39566 & ~n39587 ;
  assign n39589 = x219 & ~n39588 ;
  assign n39590 = x1156 & n36544 ;
  assign n39591 = ~x1154 & n35243 ;
  assign n39592 = n39587 & ~n39591 ;
  assign n39593 = ( x1156 & n39590 ) | ( x1156 & ~n39592 ) | ( n39590 & ~n39592 ) ;
  assign n39594 = n39589 & ~n39593 ;
  assign n39595 = x263 & x1091 ;
  assign n39596 = ~n39594 & n39595 ;
  assign n39597 = n39584 & n39596 ;
  assign n39598 = n39572 & ~n39597 ;
  assign n39599 = n37593 | n39598 ;
  assign n39600 = ~n6785 & n39599 ;
  assign n39601 = ~n39540 & n39600 ;
  assign n39602 = x211 & ~n37473 ;
  assign n39603 = n35165 | n39199 ;
  assign n39604 = ~n39602 & n39603 ;
  assign n39605 = n39009 | n39604 ;
  assign n39606 = x263 & ~n39008 ;
  assign n39607 = n39605 & n39606 ;
  assign n39608 = x263 | n39261 ;
  assign n39609 = x211 | n39310 ;
  assign n39610 = ~n35165 & n39609 ;
  assign n39611 = ~n39602 & n39610 ;
  assign n39612 = n39009 | n39611 ;
  assign n39613 = ( ~x219 & n39608 ) | ( ~x219 & n39612 ) | ( n39608 & n39612 ) ;
  assign n39614 = ~n39607 & n39613 ;
  assign n39615 = x1091 & n39478 ;
  assign n39616 = n37593 & ~n39615 ;
  assign n39617 = ~n39614 & n39616 ;
  assign n39618 = x219 | n35165 ;
  assign n39619 = n35181 | n39618 ;
  assign n39620 = ~n39478 & n39619 ;
  assign n39621 = x1091 & ~n39620 ;
  assign n39622 = x263 & ~x1091 ;
  assign n39623 = n39621 | n39622 ;
  assign n39624 = n6785 & n39623 ;
  assign n39625 = ( n6785 & n37593 ) | ( n6785 & n39624 ) | ( n37593 & n39624 ) ;
  assign n39626 = ~n39617 & n39625 ;
  assign n39627 = n37728 & ~n39626 ;
  assign n39628 = ~n39601 & n39627 ;
  assign n39629 = ( n6785 & n37728 ) | ( n6785 & n39623 ) | ( n37728 & n39623 ) ;
  assign n39630 = ( ~n6785 & n37728 ) | ( ~n6785 & n39598 ) | ( n37728 & n39598 ) ;
  assign n39631 = n39629 | n39630 ;
  assign n39632 = ~x230 & n39631 ;
  assign n39633 = ~n39628 & n39632 ;
  assign n39634 = n35241 & ~n35246 ;
  assign n39635 = x1156 | n39634 ;
  assign n39636 = ~n35422 & n35661 ;
  assign n39637 = n39635 & n39636 ;
  assign n39638 = x219 & ~n39590 ;
  assign n39639 = ~n39637 & n39638 ;
  assign n39640 = n6785 | n39639 ;
  assign n39641 = n36670 & ~n39637 ;
  assign n39642 = ( x211 & n39583 ) | ( x211 & ~n39641 ) | ( n39583 & ~n39641 ) ;
  assign n39643 = ~n39640 & n39642 ;
  assign n39644 = n6785 & n39620 ;
  assign n39645 = x230 & ~n39644 ;
  assign n39646 = ~n39643 & n39645 ;
  assign n39647 = n39633 | n39646 ;
  assign n39648 = ( ~x796 & x1091 ) | ( ~x796 & n37466 ) | ( x1091 & n37466 ) ;
  assign n39649 = ( x264 & x1091 ) | ( x264 & ~n37466 ) | ( x1091 & ~n37466 ) ;
  assign n39650 = n39648 | n39649 ;
  assign n39651 = x1091 & x1143 ;
  assign n39652 = ( x199 & n35214 ) | ( x199 & ~n39651 ) | ( n35214 & ~n39651 ) ;
  assign n39653 = n39650 & n39652 ;
  assign n39654 = n14313 | n39653 ;
  assign n39655 = x1091 & x1142 ;
  assign n39656 = ( ~x796 & x1091 ) | ( ~x796 & n37477 ) | ( x1091 & n37477 ) ;
  assign n39657 = ( x264 & x1091 ) | ( x264 & ~n37477 ) | ( x1091 & ~n37477 ) ;
  assign n39658 = n39656 | n39657 ;
  assign n39659 = ~n39655 & n39658 ;
  assign n39660 = ( x199 & x200 ) | ( x199 & ~n39659 ) | ( x200 & ~n39659 ) ;
  assign n39661 = x1091 & x1141 ;
  assign n39662 = n39658 & ~n39661 ;
  assign n39663 = ( ~x199 & x200 ) | ( ~x199 & n39662 ) | ( x200 & n39662 ) ;
  assign n39664 = ~n39660 & n39663 ;
  assign n39665 = n39654 | n39664 ;
  assign n39666 = x219 & ~n39146 ;
  assign n39667 = n36033 | n39666 ;
  assign n39668 = n39650 & n39667 ;
  assign n39669 = n14313 & ~n39668 ;
  assign n39670 = ( x211 & x219 ) | ( x211 & ~n39659 ) | ( x219 & ~n39659 ) ;
  assign n39671 = ( x211 & ~x219 ) | ( x211 & n39662 ) | ( ~x219 & n39662 ) ;
  assign n39672 = ~n39670 & n39671 ;
  assign n39673 = n39669 & ~n39672 ;
  assign n39674 = n39665 & ~n39673 ;
  assign n39675 = x230 | n39674 ;
  assign n39676 = ~x211 & x1141 ;
  assign n39677 = x219 | n35145 ;
  assign n39678 = n39676 | n39677 ;
  assign n39679 = ~n36033 & n39678 ;
  assign n39680 = ( x230 & ~n14313 ) | ( x230 & n39679 ) | ( ~n14313 & n39679 ) ;
  assign n39681 = ~x199 & x1141 ;
  assign n39682 = n36038 | n39681 ;
  assign n39683 = ~n35125 & n39682 ;
  assign n39684 = ( x230 & n14313 ) | ( x230 & n39683 ) | ( n14313 & n39683 ) ;
  assign n39685 = n39680 & n39684 ;
  assign n39686 = n39675 & ~n39685 ;
  assign n39687 = x1091 & x1144 ;
  assign n39688 = ~x200 & n39687 ;
  assign n39689 = x199 & ~n39688 ;
  assign n39690 = ( ~x819 & x1091 ) | ( ~x819 & n37466 ) | ( x1091 & n37466 ) ;
  assign n39691 = ( x265 & x1091 ) | ( x265 & ~n37466 ) | ( x1091 & ~n37466 ) ;
  assign n39692 = n39690 | n39691 ;
  assign n39693 = n39689 & n39692 ;
  assign n39694 = n14313 | n39693 ;
  assign n39695 = ( ~x819 & x1091 ) | ( ~x819 & n37477 ) | ( x1091 & n37477 ) ;
  assign n39696 = ( x265 & x1091 ) | ( x265 & ~n37477 ) | ( x1091 & ~n37477 ) ;
  assign n39697 = n39695 | n39696 ;
  assign n39698 = ~n39651 & n39697 ;
  assign n39699 = ( x199 & x200 ) | ( x199 & ~n39698 ) | ( x200 & ~n39698 ) ;
  assign n39700 = ~n39655 & n39697 ;
  assign n39701 = ( ~x199 & x200 ) | ( ~x199 & n39700 ) | ( x200 & n39700 ) ;
  assign n39702 = ~n39699 & n39701 ;
  assign n39703 = n39694 | n39702 ;
  assign n39704 = n37381 | n39666 ;
  assign n39705 = n39692 & n39704 ;
  assign n39706 = n14313 & ~n39705 ;
  assign n39707 = ( x211 & x219 ) | ( x211 & ~n39698 ) | ( x219 & ~n39698 ) ;
  assign n39708 = ( x211 & ~x219 ) | ( x211 & n39700 ) | ( ~x219 & n39700 ) ;
  assign n39709 = ~n39707 & n39708 ;
  assign n39710 = n39706 & ~n39709 ;
  assign n39711 = n39703 & ~n39710 ;
  assign n39712 = x230 | n39711 ;
  assign n39713 = ~x211 & x1142 ;
  assign n39714 = x219 | n35105 ;
  assign n39715 = n39713 | n39714 ;
  assign n39716 = ~n37381 & n39715 ;
  assign n39717 = ( x230 & ~n14313 ) | ( x230 & n39716 ) | ( ~n14313 & n39716 ) ;
  assign n39718 = n35124 | n37391 ;
  assign n39719 = ~n35130 & n39718 ;
  assign n39720 = ( x230 & n14313 ) | ( x230 & n39719 ) | ( n14313 & n39719 ) ;
  assign n39721 = n39717 & n39720 ;
  assign n39722 = n39712 & ~n39721 ;
  assign n39723 = ( ~x948 & x1091 ) | ( ~x948 & n37477 ) | ( x1091 & n37477 ) ;
  assign n39724 = ( x266 & ~x1091 ) | ( x266 & n37477 ) | ( ~x1091 & n37477 ) ;
  assign n39725 = ~n39723 & n39724 ;
  assign n39726 = x199 | n39725 ;
  assign n39727 = x1091 & x1136 ;
  assign n39728 = ( ~x948 & x1091 ) | ( ~x948 & n37466 ) | ( x1091 & n37466 ) ;
  assign n39729 = ( x266 & ~x1091 ) | ( x266 & n37466 ) | ( ~x1091 & n37466 ) ;
  assign n39730 = ~n39728 & n39729 ;
  assign n39731 = x199 & ~n39730 ;
  assign n39732 = ~n39727 & n39731 ;
  assign n39733 = n39726 & ~n39732 ;
  assign n39734 = ~x200 & n39733 ;
  assign n39735 = x1091 & x1135 ;
  assign n39736 = n39726 | n39735 ;
  assign n39737 = x200 & ~n39731 ;
  assign n39738 = n39736 & n39737 ;
  assign n39739 = n39734 | n39738 ;
  assign n39740 = ~n14313 & n39739 ;
  assign n39741 = ~x211 & x1136 ;
  assign n39742 = x219 & ~n39741 ;
  assign n39743 = n39666 | n39742 ;
  assign n39744 = ~n39730 & n39743 ;
  assign n39745 = n14313 & ~n39744 ;
  assign n39746 = x219 | n39725 ;
  assign n39747 = x1135 & n39086 ;
  assign n39748 = n39746 | n39747 ;
  assign n39749 = n39745 & n39748 ;
  assign n39750 = x230 | n39749 ;
  assign n39751 = n39740 | n39750 ;
  assign n39752 = x211 & ~x1135 ;
  assign n39753 = n39742 | n39752 ;
  assign n39754 = n8895 & ~n39753 ;
  assign n39755 = ( ~x230 & n6785 ) | ( ~x230 & n39754 ) | ( n6785 & n39754 ) ;
  assign n39756 = x299 & n39754 ;
  assign n39757 = x199 & x1136 ;
  assign n39758 = x200 | n39757 ;
  assign n39759 = ~x199 & x1135 ;
  assign n39760 = x200 & ~n39759 ;
  assign n39761 = x299 | n39760 ;
  assign n39762 = n39758 & ~n39761 ;
  assign n39763 = n39756 | n39762 ;
  assign n39764 = ( x230 & n6785 ) | ( x230 & ~n39763 ) | ( n6785 & ~n39763 ) ;
  assign n39765 = ~n39755 & n39764 ;
  assign n39766 = n39751 & ~n39765 ;
  assign n39767 = x1134 | n39766 ;
  assign n39768 = ~x199 & x1091 ;
  assign n39769 = n39733 | n39768 ;
  assign n39770 = ~x200 & n39769 ;
  assign n39771 = n39738 | n39770 ;
  assign n39772 = ~n14313 & n39771 ;
  assign n39773 = x1091 & ~n39752 ;
  assign n39774 = n39746 | n39773 ;
  assign n39775 = n39745 & n39774 ;
  assign n39776 = x230 | n39775 ;
  assign n39777 = n39772 | n39776 ;
  assign n39778 = ( x230 & ~n14313 ) | ( x230 & n39753 ) | ( ~n14313 & n39753 ) ;
  assign n39779 = n35290 & ~n39757 ;
  assign n39780 = n39760 | n39779 ;
  assign n39781 = ( x230 & n14313 ) | ( x230 & n39780 ) | ( n14313 & n39780 ) ;
  assign n39782 = n39778 & n39781 ;
  assign n39783 = n39777 & ~n39782 ;
  assign n39784 = x1134 & ~n39783 ;
  assign n39785 = n39767 & ~n39784 ;
  assign n39786 = x267 & ~n39263 ;
  assign n39787 = ~x267 & n37484 ;
  assign n39788 = ~n39008 & n39787 ;
  assign n39789 = n37592 & ~n39788 ;
  assign n39790 = ~n39786 & n39789 ;
  assign n39791 = x219 | n35169 ;
  assign n39792 = n35183 | n39791 ;
  assign n39793 = ~n35936 & n39792 ;
  assign n39794 = x1091 & ~n39793 ;
  assign n39795 = x267 | x1091 ;
  assign n39796 = n37592 | n39795 ;
  assign n39797 = ~n39794 & n39796 ;
  assign n39798 = ~n39790 & n39797 ;
  assign n39799 = n6785 & ~n39798 ;
  assign n39800 = n37728 & ~n39799 ;
  assign n39801 = x1091 & n39541 ;
  assign n39802 = n39096 & n39801 ;
  assign n39803 = x1154 & ~n39802 ;
  assign n39804 = ~x299 & n35627 ;
  assign n39805 = x1091 & ~n39804 ;
  assign n39806 = n39803 & n39805 ;
  assign n39807 = x1153 & ~n35614 ;
  assign n39808 = n39310 & ~n39807 ;
  assign n39809 = ~n36335 & n39808 ;
  assign n39810 = x219 & ~n39809 ;
  assign n39811 = ~n39806 & n39810 ;
  assign n39812 = x1155 & ~n39097 ;
  assign n39813 = n39315 & n39812 ;
  assign n39814 = x1155 | n39190 ;
  assign n39815 = n39114 & ~n39814 ;
  assign n39816 = n39813 | n39815 ;
  assign n39817 = ( x219 & x1154 ) | ( x219 & n39816 ) | ( x1154 & n39816 ) ;
  assign n39818 = n39308 & n39812 ;
  assign n39819 = x1155 | n35711 ;
  assign n39820 = x1091 & ~n39819 ;
  assign n39821 = n39818 | n39820 ;
  assign n39822 = ( x219 & ~x1154 ) | ( x219 & n39821 ) | ( ~x1154 & n39821 ) ;
  assign n39823 = n39817 | n39822 ;
  assign n39824 = ~n39811 & n39823 ;
  assign n39825 = x211 | n39824 ;
  assign n39826 = ~x1155 & n35628 ;
  assign n39827 = n35335 | n39826 ;
  assign n39828 = ~n11104 & n39827 ;
  assign n39829 = x1155 & n35622 ;
  assign n39830 = x1154 & ~n39829 ;
  assign n39831 = x1091 & n39830 ;
  assign n39832 = ~n39828 & n39831 ;
  assign n39833 = n35292 | n37666 ;
  assign n39834 = n39808 & n39833 ;
  assign n39835 = x211 & ~n39834 ;
  assign n39836 = ~n39832 & n39835 ;
  assign n39837 = n39825 & ~n39836 ;
  assign n39838 = x267 & ~n39837 ;
  assign n39839 = x1091 & ~x1155 ;
  assign n39840 = n39804 & n39839 ;
  assign n39841 = n39803 & ~n39840 ;
  assign n39842 = n39541 & n39830 ;
  assign n39843 = n39841 | n39842 ;
  assign n39844 = x211 & n39843 ;
  assign n39845 = x219 & ~n39844 ;
  assign n39846 = ~n35292 & n39310 ;
  assign n39847 = n36334 & n39846 ;
  assign n39848 = x211 | n39847 ;
  assign n39849 = ( x1154 & ~n39841 ) | ( x1154 & n39848 ) | ( ~n39841 & n39848 ) ;
  assign n39850 = n39845 & n39849 ;
  assign n39851 = n35628 & n39839 ;
  assign n39852 = n39802 | n39851 ;
  assign n39853 = ( x219 & n39791 ) | ( x219 & ~n39852 ) | ( n39791 & ~n39852 ) ;
  assign n39854 = ~x1154 & n35238 ;
  assign n39855 = n35313 | n39854 ;
  assign n39856 = n35272 & ~n39855 ;
  assign n39857 = n39146 & n39856 ;
  assign n39858 = ( x211 & ~n39853 ) | ( x211 & n39857 ) | ( ~n39853 & n39857 ) ;
  assign n39859 = n39850 | n39858 ;
  assign n39860 = ~n35230 & n39106 ;
  assign n39861 = n39287 | n39860 ;
  assign n39862 = n39819 & n39861 ;
  assign n39863 = x211 & ~x1154 ;
  assign n39864 = ~n39862 & n39863 ;
  assign n39865 = x267 | n39864 ;
  assign n39866 = n39859 & ~n39865 ;
  assign n39867 = n39838 | n39866 ;
  assign n39868 = ( n6785 & ~n37592 ) | ( n6785 & n39867 ) | ( ~n37592 & n39867 ) ;
  assign n39869 = n39237 & n39240 ;
  assign n39870 = n39327 | n39869 ;
  assign n39871 = x1154 & x1155 ;
  assign n39872 = ~n37505 & n39871 ;
  assign n39873 = ~n39245 & n39872 ;
  assign n39874 = n39870 & ~n39873 ;
  assign n39875 = x211 & ~n39874 ;
  assign n39876 = x1153 & n37507 ;
  assign n39877 = n35168 & ~n38979 ;
  assign n39878 = ~n39876 & n39877 ;
  assign n39879 = ~n39221 & n39878 ;
  assign n39880 = n37618 & n39213 ;
  assign n39881 = x1155 | n39880 ;
  assign n39882 = n39869 | n39881 ;
  assign n39883 = ~x267 & n39882 ;
  assign n39884 = ~n39879 & n39883 ;
  assign n39885 = ~n39875 & n39884 ;
  assign n39886 = n38963 | n38986 ;
  assign n39887 = n37595 & n39886 ;
  assign n39888 = x1154 & ~n39887 ;
  assign n39889 = x1154 | n37631 ;
  assign n39890 = n39071 | n39889 ;
  assign n39891 = ~x1155 & n39890 ;
  assign n39892 = ~n39888 & n39891 ;
  assign n39893 = x1155 & ~n39045 ;
  assign n39894 = n37490 | n39531 ;
  assign n39895 = n39893 & n39894 ;
  assign n39896 = n39069 & n39895 ;
  assign n39897 = x267 & ~n39896 ;
  assign n39898 = ~n39892 & n39897 ;
  assign n39899 = n39885 | n39898 ;
  assign n39900 = x219 & n39899 ;
  assign n39901 = n37492 & ~n39887 ;
  assign n39902 = n39480 & ~n39901 ;
  assign n39903 = x1154 & ~n39902 ;
  assign n39904 = ~x1154 & n38974 ;
  assign n39905 = x1155 & ~n39904 ;
  assign n39906 = n37537 & ~n39905 ;
  assign n39907 = n39903 | n39906 ;
  assign n39908 = n39346 | n39869 ;
  assign n39909 = ( x211 & n35165 ) | ( x211 & n39908 ) | ( n35165 & n39908 ) ;
  assign n39910 = n39907 & n39909 ;
  assign n39911 = x1153 & ~n37562 ;
  assign n39912 = x1155 | n39911 ;
  assign n39913 = x1153 | n39462 ;
  assign n39914 = ~n39912 & n39913 ;
  assign n39915 = n39352 | n39876 ;
  assign n39916 = x1155 & n39915 ;
  assign n39917 = x1154 & ~n39463 ;
  assign n39918 = ~n39916 & n39917 ;
  assign n39919 = ~n39914 & n39918 ;
  assign n39920 = n39064 & ~n39912 ;
  assign n39921 = n39916 | n39920 ;
  assign n39922 = ( ~x211 & n35181 ) | ( ~x211 & n39921 ) | ( n35181 & n39921 ) ;
  assign n39923 = ~n39919 & n39922 ;
  assign n39924 = x267 | n39923 ;
  assign n39925 = n39910 | n39924 ;
  assign n39926 = n39501 & n39893 ;
  assign n39927 = ~x1153 & n37575 ;
  assign n39928 = n37564 | n39927 ;
  assign n39929 = n37492 & n39928 ;
  assign n39930 = ( x1154 & n39871 ) | ( x1154 & ~n39929 ) | ( n39871 & ~n39929 ) ;
  assign n39931 = ~n39926 & n39930 ;
  assign n39932 = x1154 | n38986 ;
  assign n39933 = n37523 | n39932 ;
  assign n39934 = ~x1155 & n39933 ;
  assign n39935 = n37542 | n39932 ;
  assign n39936 = n39934 | n39935 ;
  assign n39937 = ~n39931 & n39936 ;
  assign n39938 = x211 & ~n39937 ;
  assign n39939 = x1154 & ~n39928 ;
  assign n39940 = n39934 & ~n39939 ;
  assign n39941 = n37515 | n39329 ;
  assign n39942 = x1154 & ~n37490 ;
  assign n39943 = x1155 & ~n39942 ;
  assign n39944 = n39941 & n39943 ;
  assign n39945 = x211 | n39944 ;
  assign n39946 = n39940 | n39945 ;
  assign n39947 = x267 & n39946 ;
  assign n39948 = ~n39938 & n39947 ;
  assign n39949 = x219 | n39948 ;
  assign n39950 = n39925 & ~n39949 ;
  assign n39951 = n39900 | n39950 ;
  assign n39952 = ( n6785 & n37592 ) | ( n6785 & n39951 ) | ( n37592 & n39951 ) ;
  assign n39953 = n39868 | n39952 ;
  assign n39954 = n39800 & n39953 ;
  assign n39955 = ~n39794 & n39795 ;
  assign n39956 = ( n6785 & n37728 ) | ( n6785 & ~n39955 ) | ( n37728 & ~n39955 ) ;
  assign n39957 = ( n6785 & ~n37728 ) | ( n6785 & n39867 ) | ( ~n37728 & n39867 ) ;
  assign n39958 = ~n39956 & n39957 ;
  assign n39959 = x230 | n39958 ;
  assign n39960 = n39954 | n39959 ;
  assign n39961 = x219 & ~n35622 ;
  assign n39962 = ~x1155 & n39807 ;
  assign n39963 = x1154 | n39962 ;
  assign n39964 = n35628 & n39963 ;
  assign n39965 = x1155 & n36332 ;
  assign n39966 = n39964 | n39965 ;
  assign n39967 = ~n39961 & n39966 ;
  assign n39968 = x211 & ~n39967 ;
  assign n39969 = ~x199 & x1154 ;
  assign n39970 = x200 & ~n39969 ;
  assign n39971 = ~n35302 & n35621 ;
  assign n39972 = ~n39970 & n39971 ;
  assign n39973 = n35193 | n39972 ;
  assign n39974 = x219 & n39973 ;
  assign n39975 = ( x211 & ~n35201 ) | ( x211 & n39856 ) | ( ~n35201 & n39856 ) ;
  assign n39976 = n39974 | n39975 ;
  assign n39977 = ~n6785 & n39976 ;
  assign n39978 = ~n39968 & n39977 ;
  assign n39979 = n6785 & n39793 ;
  assign n39980 = x230 & ~n39979 ;
  assign n39981 = ~n39978 & n39980 ;
  assign n39982 = n39960 & ~n39981 ;
  assign n39983 = x199 | n14313 ;
  assign n39984 = ~n36803 & n39983 ;
  assign n39985 = ~x211 & n14313 ;
  assign n39986 = n6785 | n35230 ;
  assign n39987 = ~n39985 & n39986 ;
  assign n39988 = x1152 & ~n39987 ;
  assign n39989 = n39984 & ~n39988 ;
  assign n39990 = ~x1151 & n39987 ;
  assign n39991 = x1150 & ~n39990 ;
  assign n39992 = ~n39989 & n39991 ;
  assign n39993 = x230 & ~n39992 ;
  assign n39994 = ~n6785 & n9582 ;
  assign n39995 = n6785 & n9580 ;
  assign n39996 = n39994 | n39995 ;
  assign n39997 = x1151 & n39996 ;
  assign n39998 = ( ~x1150 & n37360 ) | ( ~x1150 & n38931 ) | ( n37360 & n38931 ) ;
  assign n39999 = ( x1152 & n39997 ) | ( x1152 & n39998 ) | ( n39997 & n39998 ) ;
  assign n40000 = n14313 & ~n39134 ;
  assign n40001 = n6785 | n35301 ;
  assign n40002 = ~n40000 & n40001 ;
  assign n40003 = x1151 & ~n40002 ;
  assign n40004 = ( x1152 & ~n39998 ) | ( x1152 & n40003 ) | ( ~n39998 & n40003 ) ;
  assign n40005 = n39999 & ~n40004 ;
  assign n40006 = n39993 & ~n40005 ;
  assign n40007 = ~n38995 & n39039 ;
  assign n40008 = n37503 & n39046 ;
  assign n40009 = x219 & n38981 ;
  assign n40010 = n37497 & n40009 ;
  assign n40011 = n40008 | n40010 ;
  assign n40012 = n6785 | n38967 ;
  assign n40013 = n40011 | n40012 ;
  assign n40014 = ~n40007 & n40013 ;
  assign n40015 = x1151 | n40014 ;
  assign n40016 = n6785 | n39065 ;
  assign n40017 = x219 & n37623 ;
  assign n40018 = n40016 | n40017 ;
  assign n40019 = n39039 & ~n39262 ;
  assign n40020 = n40018 & ~n40019 ;
  assign n40021 = x1151 & ~n40020 ;
  assign n40022 = n40015 & ~n40021 ;
  assign n40023 = x268 & ~n40022 ;
  assign n40024 = n37473 & ~n40020 ;
  assign n40025 = n37551 | n40016 ;
  assign n40026 = n32977 & ~n37500 ;
  assign n40027 = n39009 & ~n40026 ;
  assign n40028 = n40025 & n40027 ;
  assign n40029 = n40024 | n40028 ;
  assign n40030 = ( x268 & x1151 ) | ( x268 & ~n40029 ) | ( x1151 & ~n40029 ) ;
  assign n40031 = n6785 & ~n39008 ;
  assign n40032 = n39036 & n40031 ;
  assign n40033 = n6785 & ~n39261 ;
  assign n40034 = ~n38993 & n40033 ;
  assign n40035 = n40032 & ~n40034 ;
  assign n40036 = x219 & ~n37501 ;
  assign n40037 = n39017 | n40036 ;
  assign n40038 = n37502 & n40037 ;
  assign n40039 = ~n6785 & n37561 ;
  assign n40040 = n40038 & n40039 ;
  assign n40041 = n40035 | n40040 ;
  assign n40042 = ( ~x268 & x1151 ) | ( ~x268 & n40041 ) | ( x1151 & n40041 ) ;
  assign n40043 = ~n40030 & n40042 ;
  assign n40044 = n40023 | n40043 ;
  assign n40045 = ~x1152 & n40044 ;
  assign n40046 = ~n38995 & n40033 ;
  assign n40047 = n37597 | n39072 ;
  assign n40048 = n40011 & n40047 ;
  assign n40049 = n6785 | n40048 ;
  assign n40050 = ~n37500 & n39048 ;
  assign n40051 = n40049 | n40050 ;
  assign n40052 = ~n40046 & n40051 ;
  assign n40053 = x1151 | n40052 ;
  assign n40054 = n37469 & ~n40012 ;
  assign n40055 = ~n39262 & n40033 ;
  assign n40056 = n40018 & ~n40055 ;
  assign n40057 = ~n40054 & n40056 ;
  assign n40058 = x1151 & ~n40057 ;
  assign n40059 = x268 & ~n40058 ;
  assign n40060 = n40053 & n40059 ;
  assign n40061 = ~x219 & n37512 ;
  assign n40062 = n40009 | n40061 ;
  assign n40063 = ~n6785 & n40062 ;
  assign n40064 = n38996 & n40031 ;
  assign n40065 = n40035 | n40064 ;
  assign n40066 = n40063 | n40065 ;
  assign n40067 = ( x268 & x1151 ) | ( x268 & n40066 ) | ( x1151 & n40066 ) ;
  assign n40068 = n38980 | n40038 ;
  assign n40069 = ~n6785 & n40068 ;
  assign n40070 = n40032 | n40069 ;
  assign n40071 = ( x268 & ~x1151 ) | ( x268 & n40070 ) | ( ~x1151 & n40070 ) ;
  assign n40072 = n40067 | n40071 ;
  assign n40073 = x1152 & n40072 ;
  assign n40074 = ~n40060 & n40073 ;
  assign n40075 = n40045 | n40074 ;
  assign n40076 = x1150 & n40075 ;
  assign n40077 = n39009 & n40031 ;
  assign n40078 = x219 | n37537 ;
  assign n40079 = n37489 & n40078 ;
  assign n40080 = n40063 & n40079 ;
  assign n40081 = n40077 | n40080 ;
  assign n40082 = ( x1151 & x1152 ) | ( x1151 & ~n40081 ) | ( x1152 & ~n40081 ) ;
  assign n40083 = ~n6785 & n40011 ;
  assign n40084 = n40064 | n40083 ;
  assign n40085 = ( x1151 & ~x1152 ) | ( x1151 & n40084 ) | ( ~x1152 & n40084 ) ;
  assign n40086 = n40082 & ~n40085 ;
  assign n40087 = n38997 | n40026 ;
  assign n40088 = n40049 & ~n40087 ;
  assign n40089 = ( x1151 & x1152 ) | ( x1151 & n40088 ) | ( x1152 & n40088 ) ;
  assign n40090 = ( ~x1151 & x1152 ) | ( ~x1151 & n40028 ) | ( x1152 & n40028 ) ;
  assign n40091 = n40089 | n40090 ;
  assign n40092 = ~n40086 & n40091 ;
  assign n40093 = x268 | n40092 ;
  assign n40094 = n6785 | n39022 ;
  assign n40095 = n39017 | n40094 ;
  assign n40096 = ~n39040 & n40095 ;
  assign n40097 = ( x1151 & x1152 ) | ( x1151 & n40096 ) | ( x1152 & n40096 ) ;
  assign n40098 = n37473 | n40020 ;
  assign n40099 = ( ~x1151 & x1152 ) | ( ~x1151 & n40098 ) | ( x1152 & n40098 ) ;
  assign n40100 = n40097 | n40099 ;
  assign n40101 = x268 & n40100 ;
  assign n40102 = x219 & n39069 ;
  assign n40103 = n6785 | n39072 ;
  assign n40104 = n40102 | n40103 ;
  assign n40105 = ~n40034 & n40104 ;
  assign n40106 = ( x1151 & x1152 ) | ( x1151 & ~n40105 ) | ( x1152 & ~n40105 ) ;
  assign n40107 = ~n39037 & n40033 ;
  assign n40108 = n39017 | n40102 ;
  assign n40109 = n37520 & n40108 ;
  assign n40110 = n6785 | n40109 ;
  assign n40111 = ~n40107 & n40110 ;
  assign n40112 = ( x1151 & ~x1152 ) | ( x1151 & n40111 ) | ( ~x1152 & n40111 ) ;
  assign n40113 = n40106 & ~n40112 ;
  assign n40114 = n40101 & ~n40113 ;
  assign n40115 = x1150 | n40114 ;
  assign n40116 = n40093 & ~n40115 ;
  assign n40117 = n40076 | n40116 ;
  assign n40118 = ( x230 & n37727 ) | ( x230 & n40117 ) | ( n37727 & n40117 ) ;
  assign n40119 = x1152 & n39992 ;
  assign n40120 = x268 & n40119 ;
  assign n40121 = ( n39992 & n40005 ) | ( n39992 & ~n40120 ) | ( n40005 & ~n40120 ) ;
  assign n40122 = x1091 & n40121 ;
  assign n40123 = x1091 & ~n40119 ;
  assign n40124 = x268 & ~n40123 ;
  assign n40125 = n40122 | n40124 ;
  assign n40126 = ( x230 & ~n37727 ) | ( x230 & n40125 ) | ( ~n37727 & n40125 ) ;
  assign n40127 = n40118 | n40126 ;
  assign n40128 = ~n40006 & n40127 ;
  assign n40129 = ~x199 & x1137 ;
  assign n40130 = x200 & ~n40129 ;
  assign n40131 = ~x199 & x1136 ;
  assign n40132 = x199 & x1138 ;
  assign n40133 = x200 | n40132 ;
  assign n40134 = n40131 | n40133 ;
  assign n40135 = ~n40130 & n40134 ;
  assign n40136 = n14313 | n40135 ;
  assign n40137 = x211 & x1137 ;
  assign n40138 = n39741 | n40137 ;
  assign n40139 = ( x219 & n14313 ) | ( x219 & ~n40138 ) | ( n14313 & ~n40138 ) ;
  assign n40140 = ~x211 & x1138 ;
  assign n40141 = ( x219 & ~n14313 ) | ( x219 & n40140 ) | ( ~n14313 & n40140 ) ;
  assign n40142 = n40139 & ~n40141 ;
  assign n40143 = n40136 & ~n40142 ;
  assign n40144 = x230 & ~n40143 ;
  assign n40145 = ~x200 & n39727 ;
  assign n40146 = x1137 & n37691 ;
  assign n40147 = n40145 | n40146 ;
  assign n40148 = n39983 | n40147 ;
  assign n40149 = x1091 & n40138 ;
  assign n40150 = n36803 & ~n40149 ;
  assign n40151 = n40148 & ~n40150 ;
  assign n40152 = ( ~x817 & x1091 ) | ( ~x817 & n37477 ) | ( x1091 & n37477 ) ;
  assign n40153 = ( x269 & x1091 ) | ( x269 & ~n37477 ) | ( x1091 & ~n37477 ) ;
  assign n40154 = n40152 | n40153 ;
  assign n40155 = ~n40151 & n40154 ;
  assign n40156 = x1138 & n39146 ;
  assign n40157 = x219 & n14313 ;
  assign n40158 = ~n40156 & n40157 ;
  assign n40159 = ~x200 & x1091 ;
  assign n40160 = x1138 & n40159 ;
  assign n40161 = x199 & ~n40160 ;
  assign n40162 = ~n14313 & n40161 ;
  assign n40163 = n40158 | n40162 ;
  assign n40164 = ( ~x817 & x1091 ) | ( ~x817 & n37466 ) | ( x1091 & n37466 ) ;
  assign n40165 = ( x269 & x1091 ) | ( x269 & ~n37466 ) | ( x1091 & ~n37466 ) ;
  assign n40166 = n40164 | n40165 ;
  assign n40167 = n40163 & n40166 ;
  assign n40168 = n40155 | n40167 ;
  assign n40169 = ~x230 & n40168 ;
  assign n40170 = n40144 | n40169 ;
  assign n40171 = ~x211 & x1139 ;
  assign n40172 = x211 & x1140 ;
  assign n40173 = n40171 | n40172 ;
  assign n40174 = x1091 & n40173 ;
  assign n40175 = n36803 & ~n40174 ;
  assign n40176 = x1091 & x1140 ;
  assign n40177 = x200 & n40176 ;
  assign n40178 = x1139 & n40159 ;
  assign n40179 = n40177 | n40178 ;
  assign n40180 = n39983 | n40179 ;
  assign n40181 = ~n40175 & n40180 ;
  assign n40182 = ( ~x805 & x1091 ) | ( ~x805 & n37477 ) | ( x1091 & n37477 ) ;
  assign n40183 = ( x270 & x1091 ) | ( x270 & ~n37477 ) | ( x1091 & ~n37477 ) ;
  assign n40184 = n40182 | n40183 ;
  assign n40185 = ~n40181 & n40184 ;
  assign n40186 = n39146 & n39676 ;
  assign n40187 = n40157 & ~n40186 ;
  assign n40188 = ( x199 & n35214 ) | ( x199 & ~n39661 ) | ( n35214 & ~n39661 ) ;
  assign n40189 = ~n14313 & n40188 ;
  assign n40190 = n40187 | n40189 ;
  assign n40191 = ( ~x805 & x1091 ) | ( ~x805 & n37466 ) | ( x1091 & n37466 ) ;
  assign n40192 = ( x270 & x1091 ) | ( x270 & ~n37466 ) | ( x1091 & ~n37466 ) ;
  assign n40193 = n40191 | n40192 ;
  assign n40194 = n40190 & n40193 ;
  assign n40195 = x230 | n40194 ;
  assign n40196 = n40185 | n40195 ;
  assign n40197 = ~x199 & x1140 ;
  assign n40198 = x200 & ~n40197 ;
  assign n40199 = ~x199 & x1139 ;
  assign n40200 = x199 & x1141 ;
  assign n40201 = x200 | n40200 ;
  assign n40202 = n40199 | n40201 ;
  assign n40203 = ~n40198 & n40202 ;
  assign n40204 = n14313 | n40203 ;
  assign n40205 = ( x219 & n14313 ) | ( x219 & ~n40173 ) | ( n14313 & ~n40173 ) ;
  assign n40206 = ( x219 & ~n14313 ) | ( x219 & n39676 ) | ( ~n14313 & n39676 ) ;
  assign n40207 = n40205 & ~n40206 ;
  assign n40208 = x230 & ~n40207 ;
  assign n40209 = n40204 & n40208 ;
  assign n40210 = n40196 & ~n40209 ;
  assign n40211 = x271 | n37498 ;
  assign n40212 = ~n37470 & n40211 ;
  assign n40213 = x219 & ~n40212 ;
  assign n40214 = x1091 | n37479 ;
  assign n40215 = x271 & n40214 ;
  assign n40216 = x271 | n37480 ;
  assign n40217 = ~n40215 & n40216 ;
  assign n40218 = x1091 & x1146 ;
  assign n40219 = n40217 | n40218 ;
  assign n40220 = ~x211 & n40218 ;
  assign n40221 = n40219 & ~n40220 ;
  assign n40222 = x1091 & n36026 ;
  assign n40223 = x219 | n40222 ;
  assign n40224 = n40221 | n40223 ;
  assign n40225 = ~n40213 & n40224 ;
  assign n40226 = ~x211 & x1147 ;
  assign n40227 = n39000 & n40226 ;
  assign n40228 = n14313 & ~n40227 ;
  assign n40229 = ~n40225 & n40228 ;
  assign n40230 = x199 & ~n40212 ;
  assign n40231 = x199 | n40219 ;
  assign n40232 = ~n40230 & n40231 ;
  assign n40233 = x200 & ~n40232 ;
  assign n40234 = x1091 & x1145 ;
  assign n40235 = x199 | n40234 ;
  assign n40236 = n40217 | n40235 ;
  assign n40237 = ~n40230 & n40236 ;
  assign n40238 = x1147 & n37675 ;
  assign n40239 = x200 | n40238 ;
  assign n40240 = n40237 | n40239 ;
  assign n40241 = ~n40233 & n40240 ;
  assign n40242 = n14313 | n40241 ;
  assign n40243 = ~n40229 & n40242 ;
  assign n40244 = x230 | n40243 ;
  assign n40245 = x219 & ~n40226 ;
  assign n40246 = n36026 | n38218 ;
  assign n40247 = ~n40245 & n40246 ;
  assign n40248 = ( ~x230 & n6785 ) | ( ~x230 & n40247 ) | ( n6785 & n40247 ) ;
  assign n40249 = x200 | n36042 ;
  assign n40250 = ~n36958 & n40249 ;
  assign n40251 = x1147 & n38928 ;
  assign n40252 = n36853 | n36896 ;
  assign n40253 = ~x219 & n40252 ;
  assign n40254 = n40251 | n40253 ;
  assign n40255 = n40250 | n40254 ;
  assign n40256 = ( x230 & n6785 ) | ( x230 & ~n40255 ) | ( n6785 & ~n40255 ) ;
  assign n40257 = ~n40248 & n40256 ;
  assign n40258 = n40244 & ~n40257 ;
  assign n40259 = x1150 & n40066 ;
  assign n40260 = ~x1150 & n40029 ;
  assign n40261 = x1149 & ~n40260 ;
  assign n40262 = ~n40259 & n40261 ;
  assign n40263 = x1150 & n40070 ;
  assign n40264 = ~x1150 & n40041 ;
  assign n40265 = x1149 | n40264 ;
  assign n40266 = n40263 | n40265 ;
  assign n40267 = ~n40262 & n40266 ;
  assign n40268 = x1148 & ~n40267 ;
  assign n40269 = x1150 | n40088 ;
  assign n40270 = x1150 & ~n40084 ;
  assign n40271 = x1149 & ~n40270 ;
  assign n40272 = n40269 & n40271 ;
  assign n40273 = x1150 & ~n40081 ;
  assign n40274 = x1150 | n40028 ;
  assign n40275 = ~x1149 & n40274 ;
  assign n40276 = ~n40273 & n40275 ;
  assign n40277 = x1148 | n40276 ;
  assign n40278 = n40272 | n40277 ;
  assign n40279 = ~n40268 & n40278 ;
  assign n40280 = x283 & ~n40279 ;
  assign n40281 = n6785 | n35221 ;
  assign n40282 = ~n36803 & n40281 ;
  assign n40283 = ~n39985 & n40282 ;
  assign n40284 = x1150 & ~n40283 ;
  assign n40285 = x1149 & ~n40284 ;
  assign n40286 = n39984 & n40285 ;
  assign n40287 = n6785 & ~n8895 ;
  assign n40288 = n11107 & ~n40287 ;
  assign n40289 = ~x1150 & n40288 ;
  assign n40290 = n39987 | n40289 ;
  assign n40291 = ~x1149 & n40290 ;
  assign n40292 = x1148 & ~n40291 ;
  assign n40293 = ~n40286 & n40292 ;
  assign n40294 = x1091 & n40293 ;
  assign n40295 = x1150 & n38931 ;
  assign n40296 = x1149 | n40295 ;
  assign n40297 = ~x1148 & n40296 ;
  assign n40298 = x1150 & n40002 ;
  assign n40299 = ~x1150 & n39996 ;
  assign n40300 = x1149 & ~n40299 ;
  assign n40301 = ~n40298 & n40300 ;
  assign n40302 = x1091 & ~n40301 ;
  assign n40303 = n40297 & n40302 ;
  assign n40304 = x283 | n40303 ;
  assign n40305 = n40294 | n40304 ;
  assign n40306 = ~x272 & n40305 ;
  assign n40307 = ~n40280 & n40306 ;
  assign n40308 = x1150 & n40052 ;
  assign n40309 = ( x1149 & ~n37336 ) | ( x1149 & n40014 ) | ( ~n37336 & n40014 ) ;
  assign n40310 = n40308 | n40309 ;
  assign n40311 = ( ~x1149 & x1150 ) | ( ~x1149 & n40057 ) | ( x1150 & n40057 ) ;
  assign n40312 = ( x1149 & x1150 ) | ( x1149 & ~n40020 ) | ( x1150 & ~n40020 ) ;
  assign n40313 = ~n40311 & n40312 ;
  assign n40314 = n40310 & ~n40313 ;
  assign n40315 = ( x283 & ~x1148 ) | ( x283 & n40314 ) | ( ~x1148 & n40314 ) ;
  assign n40316 = x1150 & n40105 ;
  assign n40317 = ~x1150 & n40098 ;
  assign n40318 = x1149 | n40317 ;
  assign n40319 = n40316 | n40318 ;
  assign n40320 = x1150 & n40111 ;
  assign n40321 = ~x1150 & n40096 ;
  assign n40322 = x1149 & ~n40321 ;
  assign n40323 = ~n40320 & n40322 ;
  assign n40324 = n40319 & ~n40323 ;
  assign n40325 = ( x283 & x1148 ) | ( x283 & n40324 ) | ( x1148 & n40324 ) ;
  assign n40326 = n40315 & n40325 ;
  assign n40327 = x1091 & ~n40296 ;
  assign n40328 = x1148 | n40327 ;
  assign n40329 = x1091 & ~n40002 ;
  assign n40330 = ( x1149 & ~x1150 ) | ( x1149 & n40329 ) | ( ~x1150 & n40329 ) ;
  assign n40331 = n14313 & n39321 ;
  assign n40332 = ~n6785 & n37680 ;
  assign n40333 = n40331 | n40332 ;
  assign n40334 = ( x1149 & x1150 ) | ( x1149 & n40333 ) | ( x1150 & n40333 ) ;
  assign n40335 = n40330 & n40334 ;
  assign n40336 = n40328 | n40335 ;
  assign n40337 = n37255 | n39987 ;
  assign n40338 = n39984 & n40337 ;
  assign n40339 = n40291 | n40338 ;
  assign n40340 = x1091 & n40339 ;
  assign n40341 = x1148 & ~n40340 ;
  assign n40342 = n40336 & ~n40341 ;
  assign n40343 = ( x272 & n37726 ) | ( x272 & ~n40342 ) | ( n37726 & ~n40342 ) ;
  assign n40344 = ~n40326 & n40343 ;
  assign n40345 = x230 | n40344 ;
  assign n40346 = n40307 | n40345 ;
  assign n40347 = x1149 & ~n40002 ;
  assign n40348 = n40285 | n40347 ;
  assign n40349 = ~n40299 & n40348 ;
  assign n40350 = n40297 & ~n40349 ;
  assign n40351 = x230 & ~n40293 ;
  assign n40352 = ~n40350 & n40351 ;
  assign n40353 = n40346 & ~n40352 ;
  assign n40354 = x273 | n37499 ;
  assign n40355 = ~n37472 & n40354 ;
  assign n40356 = x219 & ~n40355 ;
  assign n40357 = x273 | n37481 ;
  assign n40358 = ~n37483 & n40357 ;
  assign n40359 = x219 | n40220 ;
  assign n40360 = n40358 | n40359 ;
  assign n40361 = ~n40356 & n40360 ;
  assign n40362 = x299 & n40361 ;
  assign n40363 = ~x200 & n40218 ;
  assign n40364 = x199 | n40363 ;
  assign n40365 = n40358 | n40364 ;
  assign n40366 = x199 & ~n40355 ;
  assign n40367 = x299 | n40366 ;
  assign n40368 = n40365 & ~n40367 ;
  assign n40369 = n40362 | n40368 ;
  assign n40370 = n9581 | n37620 ;
  assign n40371 = x1091 & n40370 ;
  assign n40372 = n40369 | n40371 ;
  assign n40373 = ~n6785 & n40372 ;
  assign n40374 = x1091 & n39040 ;
  assign n40375 = n40373 | n40374 ;
  assign n40376 = x1147 & n40375 ;
  assign n40377 = n6785 & n40361 ;
  assign n40378 = ~n37042 & n40369 ;
  assign n40379 = x1148 | n40378 ;
  assign n40380 = x1091 & n35201 ;
  assign n40381 = n40361 | n40380 ;
  assign n40382 = x299 & n40381 ;
  assign n40383 = n37676 & ~n40233 ;
  assign n40384 = n40368 | n40383 ;
  assign n40385 = n40382 | n40384 ;
  assign n40386 = ~n6785 & n40385 ;
  assign n40387 = n36716 & n39000 ;
  assign n40388 = x1148 & ~n40387 ;
  assign n40389 = ~n40386 & n40388 ;
  assign n40390 = n40379 & ~n40389 ;
  assign n40391 = n40377 | n40390 ;
  assign n40392 = n40376 | n40391 ;
  assign n40393 = ~x230 & n40392 ;
  assign n40394 = x1146 | n8895 ;
  assign n40395 = x1147 & n36803 ;
  assign n40396 = n39985 | n40395 ;
  assign n40397 = n40394 & n40396 ;
  assign n40398 = x1146 | n8980 ;
  assign n40399 = ~x199 & x1147 ;
  assign n40400 = x200 & ~n40399 ;
  assign n40401 = n40398 & ~n40400 ;
  assign n40402 = ~n14313 & n40401 ;
  assign n40403 = x1148 & ~n40402 ;
  assign n40404 = ~n40397 & n40403 ;
  assign n40405 = x211 | n36859 ;
  assign n40406 = n36803 & n40405 ;
  assign n40407 = ~n39983 & n40398 ;
  assign n40408 = n40406 | n40407 ;
  assign n40409 = x1147 & n40408 ;
  assign n40410 = x1146 & ~n37964 ;
  assign n40411 = ~n40288 & n40410 ;
  assign n40412 = x1148 | n40411 ;
  assign n40413 = n40409 | n40412 ;
  assign n40414 = x230 & n40413 ;
  assign n40415 = ~n40404 & n40414 ;
  assign n40416 = n40393 | n40415 ;
  assign n40417 = x219 & ~n40222 ;
  assign n40418 = ( ~x659 & x1091 ) | ( ~x659 & n37466 ) | ( x1091 & n37466 ) ;
  assign n40419 = ( x274 & x1091 ) | ( x274 & ~n37466 ) | ( x1091 & ~n37466 ) ;
  assign n40420 = n40418 | n40419 ;
  assign n40421 = n40417 & n40420 ;
  assign n40422 = n14313 & ~n40421 ;
  assign n40423 = ( ~x659 & x1091 ) | ( ~x659 & n37477 ) | ( x1091 & n37477 ) ;
  assign n40424 = ( x274 & x1091 ) | ( x274 & ~n37477 ) | ( x1091 & ~n37477 ) ;
  assign n40425 = n40423 | n40424 ;
  assign n40426 = ~n39687 & n40425 ;
  assign n40427 = ( x211 & x219 ) | ( x211 & ~n40426 ) | ( x219 & ~n40426 ) ;
  assign n40428 = ~n39651 & n40425 ;
  assign n40429 = ( x211 & ~x219 ) | ( x211 & n40428 ) | ( ~x219 & n40428 ) ;
  assign n40430 = ~n40427 & n40429 ;
  assign n40431 = n40422 & ~n40430 ;
  assign n40432 = ( x199 & n35214 ) | ( x199 & ~n40234 ) | ( n35214 & ~n40234 ) ;
  assign n40433 = n40420 & n40432 ;
  assign n40434 = n14313 | n40433 ;
  assign n40435 = ( x199 & x200 ) | ( x199 & ~n40426 ) | ( x200 & ~n40426 ) ;
  assign n40436 = ( ~x199 & x200 ) | ( ~x199 & n40428 ) | ( x200 & n40428 ) ;
  assign n40437 = ~n40435 & n40436 ;
  assign n40438 = n40434 | n40437 ;
  assign n40439 = ~x230 & n40438 ;
  assign n40440 = ~n40431 & n40439 ;
  assign n40441 = x219 | n35112 ;
  assign n40442 = n36027 | n40441 ;
  assign n40443 = n36847 & n40442 ;
  assign n40444 = n35191 | n36853 ;
  assign n40445 = n40442 & n40444 ;
  assign n40446 = n35121 | n36963 ;
  assign n40447 = ~n37398 & n40446 ;
  assign n40448 = n40445 | n40447 ;
  assign n40449 = ~n6785 & n40448 ;
  assign n40450 = x230 & ~n40449 ;
  assign n40451 = ~n40443 & n40450 ;
  assign n40452 = n40440 | n40451 ;
  assign n40453 = x1151 & ~n40052 ;
  assign n40454 = ~x1150 & n40015 ;
  assign n40455 = ~n40453 & n40454 ;
  assign n40456 = x1151 | n40020 ;
  assign n40457 = x1150 & n40456 ;
  assign n40458 = ~n40058 & n40457 ;
  assign n40459 = x275 & ~n40458 ;
  assign n40460 = ~n40455 & n40459 ;
  assign n40461 = ~x1150 & n40070 ;
  assign n40462 = x1151 & ~n40259 ;
  assign n40463 = ~n40461 & n40462 ;
  assign n40464 = x1150 & n40029 ;
  assign n40465 = x1151 | n40464 ;
  assign n40466 = n40264 | n40465 ;
  assign n40467 = ~x275 & n40466 ;
  assign n40468 = ~n40463 & n40467 ;
  assign n40469 = x1149 & ~n40468 ;
  assign n40470 = ~n40460 & n40469 ;
  assign n40471 = x1150 | n40081 ;
  assign n40472 = x1151 & ~n40270 ;
  assign n40473 = n40471 & n40472 ;
  assign n40474 = x1150 & ~n40088 ;
  assign n40475 = ~x1151 & n40274 ;
  assign n40476 = ~n40474 & n40475 ;
  assign n40477 = n40473 | n40476 ;
  assign n40478 = ~x275 & n40477 ;
  assign n40479 = ~x1150 & n40105 ;
  assign n40480 = n40320 | n40479 ;
  assign n40481 = ( ~x275 & x1151 ) | ( ~x275 & n40480 ) | ( x1151 & n40480 ) ;
  assign n40482 = x1150 & n40096 ;
  assign n40483 = n40317 | n40482 ;
  assign n40484 = ( x275 & x1151 ) | ( x275 & ~n40483 ) | ( x1151 & ~n40483 ) ;
  assign n40485 = ~n40481 & n40484 ;
  assign n40486 = x1149 | n40485 ;
  assign n40487 = n40478 | n40486 ;
  assign n40488 = n37726 & n40487 ;
  assign n40489 = ~n40470 & n40488 ;
  assign n40490 = x1151 | n39996 ;
  assign n40491 = x1150 & n40490 ;
  assign n40492 = ~n40003 & n40491 ;
  assign n40493 = n37360 & n38931 ;
  assign n40494 = x1149 | n40493 ;
  assign n40495 = n40492 | n40494 ;
  assign n40496 = x1151 & ~n39987 ;
  assign n40497 = x1149 & n39984 ;
  assign n40498 = ~n40496 & n40497 ;
  assign n40499 = n37255 & n39987 ;
  assign n40500 = n40498 | n40499 ;
  assign n40501 = n40495 & ~n40500 ;
  assign n40502 = x1091 & n40501 ;
  assign n40503 = ( x275 & ~n37726 ) | ( x275 & n40502 ) | ( ~n37726 & n40502 ) ;
  assign n40504 = ~x1149 & n40003 ;
  assign n40505 = n40498 | n40504 ;
  assign n40506 = x1150 & n40505 ;
  assign n40507 = ~x1151 & n40288 ;
  assign n40508 = x1149 & ~n39987 ;
  assign n40509 = ~n40507 & n40508 ;
  assign n40510 = ~x1149 & x1151 ;
  assign n40511 = n38931 & n40510 ;
  assign n40512 = x1150 | n40511 ;
  assign n40513 = n40509 | n40512 ;
  assign n40514 = ~n40506 & n40513 ;
  assign n40515 = x1091 & ~n40514 ;
  assign n40516 = ~x1151 & n37336 ;
  assign n40517 = n40333 & n40516 ;
  assign n40518 = n40515 | n40517 ;
  assign n40519 = ( x275 & n37726 ) | ( x275 & n40518 ) | ( n37726 & n40518 ) ;
  assign n40520 = n40503 & ~n40519 ;
  assign n40521 = n40489 | n40520 ;
  assign n40522 = ~x230 & n40521 ;
  assign n40523 = x230 & n40501 ;
  assign n40524 = n40522 | n40523 ;
  assign n40525 = x276 | n37478 ;
  assign n40526 = ~n40214 & n40525 ;
  assign n40527 = n35106 | n36836 ;
  assign n40528 = x1091 & n40527 ;
  assign n40529 = n36803 & ~n40528 ;
  assign n40530 = x1145 & n37691 ;
  assign n40531 = n39688 | n40530 ;
  assign n40532 = n39983 | n40531 ;
  assign n40533 = ~n40529 & n40532 ;
  assign n40534 = n40526 | n40533 ;
  assign n40535 = ~x230 & n40534 ;
  assign n40536 = n40157 & ~n40220 ;
  assign n40537 = x199 & ~n40363 ;
  assign n40538 = ~n14313 & n40537 ;
  assign n40539 = n40536 | n40538 ;
  assign n40540 = ( x276 & ~x1091 ) | ( x276 & n37467 ) | ( ~x1091 & n37467 ) ;
  assign n40541 = ( n37468 & n40539 ) | ( n37468 & ~n40540 ) | ( n40539 & ~n40540 ) ;
  assign n40542 = n40535 & ~n40541 ;
  assign n40543 = ~x219 & n40527 ;
  assign n40544 = x1146 & n35201 ;
  assign n40545 = n40543 | n40544 ;
  assign n40546 = ( x230 & ~n14313 ) | ( x230 & n40545 ) | ( ~n14313 & n40545 ) ;
  assign n40547 = n35128 | n37827 ;
  assign n40548 = ~n36965 & n40547 ;
  assign n40549 = ( x230 & n14313 ) | ( x230 & n40548 ) | ( n14313 & n40548 ) ;
  assign n40550 = n40546 & n40549 ;
  assign n40551 = n40542 | n40550 ;
  assign n40552 = ( ~x820 & x1091 ) | ( ~x820 & n37466 ) | ( x1091 & n37466 ) ;
  assign n40553 = ( x277 & x1091 ) | ( x277 & ~n37466 ) | ( x1091 & ~n37466 ) ;
  assign n40554 = n40552 | n40553 ;
  assign n40555 = ( x199 & n35214 ) | ( x199 & ~n39655 ) | ( n35214 & ~n39655 ) ;
  assign n40556 = n40554 & n40555 ;
  assign n40557 = n14313 | n40556 ;
  assign n40558 = ( ~x820 & x1091 ) | ( ~x820 & n37477 ) | ( x1091 & n37477 ) ;
  assign n40559 = ( x277 & x1091 ) | ( x277 & ~n37477 ) | ( x1091 & ~n37477 ) ;
  assign n40560 = n40558 | n40559 ;
  assign n40561 = ~n39661 & n40560 ;
  assign n40562 = ( x199 & x200 ) | ( x199 & ~n40561 ) | ( x200 & ~n40561 ) ;
  assign n40563 = ~n40176 & n40560 ;
  assign n40564 = ( ~x199 & x200 ) | ( ~x199 & n40563 ) | ( x200 & n40563 ) ;
  assign n40565 = ~n40562 & n40564 ;
  assign n40566 = n40557 | n40565 ;
  assign n40567 = x219 & ~n39713 ;
  assign n40568 = n39666 | n40567 ;
  assign n40569 = n40554 & n40568 ;
  assign n40570 = n14313 & ~n40569 ;
  assign n40571 = ( x211 & x219 ) | ( x211 & ~n40561 ) | ( x219 & ~n40561 ) ;
  assign n40572 = ( x211 & ~x219 ) | ( x211 & n40563 ) | ( ~x219 & n40563 ) ;
  assign n40573 = ~n40571 & n40572 ;
  assign n40574 = n40570 & ~n40573 ;
  assign n40575 = n40566 & ~n40574 ;
  assign n40576 = x230 | n40575 ;
  assign n40577 = ~x211 & x1140 ;
  assign n40578 = x211 & x1141 ;
  assign n40579 = x219 | n40578 ;
  assign n40580 = n40577 | n40579 ;
  assign n40581 = ~n40567 & n40580 ;
  assign n40582 = ( x230 & ~n14313 ) | ( x230 & n40581 ) | ( ~n14313 & n40581 ) ;
  assign n40583 = n35120 | n40197 ;
  assign n40584 = x200 & ~n39681 ;
  assign n40585 = n40583 & ~n40584 ;
  assign n40586 = ( x230 & n14313 ) | ( x230 & n40585 ) | ( n14313 & n40585 ) ;
  assign n40587 = n40582 & n40586 ;
  assign n40588 = n40576 & ~n40587 ;
  assign n40589 = ( ~x976 & x1091 ) | ( ~x976 & n37466 ) | ( x1091 & n37466 ) ;
  assign n40590 = ( x278 & ~x1091 ) | ( x278 & n37466 ) | ( ~x1091 & n37466 ) ;
  assign n40591 = ~n40589 & n40590 ;
  assign n40592 = x199 & ~n40591 ;
  assign n40593 = x1091 & ~x1132 ;
  assign n40594 = ( x976 & x1091 ) | ( x976 & n37477 ) | ( x1091 & n37477 ) ;
  assign n40595 = ( x278 & x1091 ) | ( x278 & ~n37477 ) | ( x1091 & ~n37477 ) ;
  assign n40596 = n40594 | n40595 ;
  assign n40597 = ~n40593 & n40596 ;
  assign n40598 = x199 | n40597 ;
  assign n40599 = ~n40592 & n40598 ;
  assign n40600 = x200 | n40599 ;
  assign n40601 = x1091 & ~x1133 ;
  assign n40602 = n40596 & ~n40601 ;
  assign n40603 = x199 | n40602 ;
  assign n40604 = ~n40592 & n40603 ;
  assign n40605 = x200 & ~n40604 ;
  assign n40606 = x299 | n40605 ;
  assign n40607 = n40600 & ~n40606 ;
  assign n40608 = x219 & ~n40591 ;
  assign n40609 = x211 & ~x1133 ;
  assign n40610 = x211 | x1132 ;
  assign n40611 = ~n40609 & n40610 ;
  assign n40612 = x1091 & ~n40611 ;
  assign n40613 = n40596 & ~n40612 ;
  assign n40614 = x219 | n40613 ;
  assign n40615 = ~n40608 & n40614 ;
  assign n40616 = x299 & n40615 ;
  assign n40617 = n40607 | n40616 ;
  assign n40618 = ~n6785 & n40617 ;
  assign n40619 = n6785 & n40615 ;
  assign n40620 = x230 | n40619 ;
  assign n40621 = n40618 | n40620 ;
  assign n40622 = ~x199 & x1132 ;
  assign n40623 = x200 | n40622 ;
  assign n40624 = ~x199 & x1133 ;
  assign n40625 = x200 & ~n40624 ;
  assign n40626 = x299 | n40625 ;
  assign n40627 = n40623 & ~n40626 ;
  assign n40628 = n35191 & n40611 ;
  assign n40629 = n40627 | n40628 ;
  assign n40630 = ~n6785 & n40629 ;
  assign n40631 = n36061 & n40611 ;
  assign n40632 = x230 & ~n40631 ;
  assign n40633 = ~n40630 & n40632 ;
  assign n40634 = n40621 & ~n40633 ;
  assign n40635 = x1134 | n40634 ;
  assign n40636 = x219 | n40611 ;
  assign n40637 = n36717 & n40636 ;
  assign n40638 = n8980 | n40622 ;
  assign n40639 = ~n40626 & n40638 ;
  assign n40640 = n39160 | n40628 ;
  assign n40641 = n40639 | n40640 ;
  assign n40642 = ~n6785 & n40641 ;
  assign n40643 = x230 & ~n40642 ;
  assign n40644 = ~n40637 & n40643 ;
  assign n40645 = n37675 | n40600 ;
  assign n40646 = ~n40606 & n40645 ;
  assign n40647 = n11104 & n39146 ;
  assign n40648 = n40616 | n40647 ;
  assign n40649 = n40646 | n40648 ;
  assign n40650 = ~n6785 & n40649 ;
  assign n40651 = n40387 | n40620 ;
  assign n40652 = n40650 | n40651 ;
  assign n40653 = ~n40644 & n40652 ;
  assign n40654 = x1134 & ~n40653 ;
  assign n40655 = n40635 & ~n40654 ;
  assign n40656 = x1135 & n40159 ;
  assign n40657 = ( ~x958 & x1091 ) | ( ~x958 & n37466 ) | ( x1091 & n37466 ) ;
  assign n40658 = ( x279 & ~x1091 ) | ( x279 & n37466 ) | ( ~x1091 & n37466 ) ;
  assign n40659 = ~n40657 & n40658 ;
  assign n40660 = n40656 | n40659 ;
  assign n40661 = x199 & n40660 ;
  assign n40662 = ( x958 & x1091 ) | ( x958 & n37477 ) | ( x1091 & n37477 ) ;
  assign n40663 = ( x279 & x1091 ) | ( x279 & ~n37477 ) | ( x1091 & ~n37477 ) ;
  assign n40664 = n40662 | n40663 ;
  assign n40665 = ( x199 & ~n9578 ) | ( x199 & n40601 ) | ( ~n9578 & n40601 ) ;
  assign n40666 = n40664 & ~n40665 ;
  assign n40667 = n40661 | n40666 ;
  assign n40668 = ~n14313 & n40667 ;
  assign n40669 = ~n37691 & n40668 ;
  assign n40670 = n39086 | n40601 ;
  assign n40671 = n40664 & ~n40670 ;
  assign n40672 = x219 | n40671 ;
  assign n40673 = x1135 & n39146 ;
  assign n40674 = x219 & ~n40673 ;
  assign n40675 = ~n40659 & n40674 ;
  assign n40676 = n14313 & ~n40675 ;
  assign n40677 = n40672 & n40676 ;
  assign n40678 = x230 | n40677 ;
  assign n40679 = n40669 | n40678 ;
  assign n40680 = x1135 & n35201 ;
  assign n40681 = x211 | x1133 ;
  assign n40682 = ~x219 & n40681 ;
  assign n40683 = ~x211 & n40682 ;
  assign n40684 = n40680 | n40683 ;
  assign n40685 = ( ~x230 & n6785 ) | ( ~x230 & n40684 ) | ( n6785 & n40684 ) ;
  assign n40686 = x199 & x1135 ;
  assign n40687 = n40624 | n40686 ;
  assign n40688 = ~n35230 & n40687 ;
  assign n40689 = x299 & n40684 ;
  assign n40690 = n40688 | n40689 ;
  assign n40691 = ( x230 & n6785 ) | ( x230 & ~n40690 ) | ( n6785 & ~n40690 ) ;
  assign n40692 = ~n40685 & n40691 ;
  assign n40693 = n40679 & ~n40692 ;
  assign n40694 = x1134 | n40693 ;
  assign n40695 = x1091 & n40681 ;
  assign n40696 = n36803 & n40695 ;
  assign n40697 = n40668 | n40696 ;
  assign n40698 = n40678 | n40697 ;
  assign n40699 = n40680 | n40682 ;
  assign n40700 = ( ~x230 & n14313 ) | ( ~x230 & n40699 ) | ( n14313 & n40699 ) ;
  assign n40701 = x1133 | n8980 ;
  assign n40702 = ~x200 & x1135 ;
  assign n40703 = x199 & ~n40702 ;
  assign n40704 = n40701 & ~n40703 ;
  assign n40705 = ( x230 & n14313 ) | ( x230 & ~n40704 ) | ( n14313 & ~n40704 ) ;
  assign n40706 = ~n40700 & n40705 ;
  assign n40707 = n40698 & ~n40706 ;
  assign n40708 = x1134 & ~n40707 ;
  assign n40709 = n40694 & ~n40708 ;
  assign n40710 = ~x211 & x1135 ;
  assign n40711 = x211 & x1136 ;
  assign n40712 = n40710 | n40711 ;
  assign n40713 = x1091 & ~n40712 ;
  assign n40714 = ( x914 & x1091 ) | ( x914 & n37477 ) | ( x1091 & n37477 ) ;
  assign n40715 = ( x280 & ~x1091 ) | ( x280 & n37477 ) | ( ~x1091 & n37477 ) ;
  assign n40716 = ~n40714 & n40715 ;
  assign n40717 = n40713 | n40716 ;
  assign n40718 = ~x219 & n40717 ;
  assign n40719 = ~x211 & x1137 ;
  assign n40720 = x219 & ~n40719 ;
  assign n40721 = n39666 | n40720 ;
  assign n40722 = ( ~x914 & x1091 ) | ( ~x914 & n37466 ) | ( x1091 & n37466 ) ;
  assign n40723 = ( x280 & x1091 ) | ( x280 & ~n37466 ) | ( x1091 & ~n37466 ) ;
  assign n40724 = n40722 | n40723 ;
  assign n40725 = n40721 & n40724 ;
  assign n40726 = n40718 | n40725 ;
  assign n40727 = n14313 & n40726 ;
  assign n40728 = x200 & x1136 ;
  assign n40729 = x1091 & ~n40702 ;
  assign n40730 = ~n40728 & n40729 ;
  assign n40731 = x199 | n40730 ;
  assign n40732 = n40716 | n40731 ;
  assign n40733 = x1137 & n40159 ;
  assign n40734 = n40724 & ~n40733 ;
  assign n40735 = x199 & ~n40734 ;
  assign n40736 = n14313 | n40735 ;
  assign n40737 = n40732 & ~n40736 ;
  assign n40738 = n40727 | n40737 ;
  assign n40739 = ~x230 & n40738 ;
  assign n40740 = x219 | n40712 ;
  assign n40741 = ~n40720 & n40740 ;
  assign n40742 = ( ~x230 & n14313 ) | ( ~x230 & n40741 ) | ( n14313 & n40741 ) ;
  assign n40743 = x200 & ~n40131 ;
  assign n40744 = x199 & x1137 ;
  assign n40745 = x200 | n39759 ;
  assign n40746 = n40744 | n40745 ;
  assign n40747 = ~n40743 & n40746 ;
  assign n40748 = ( x230 & n14313 ) | ( x230 & ~n40747 ) | ( n14313 & ~n40747 ) ;
  assign n40749 = ~n40742 & n40748 ;
  assign n40750 = n40739 | n40749 ;
  assign n40751 = ~x199 & x1138 ;
  assign n40752 = x200 & ~n40751 ;
  assign n40753 = x199 & x1139 ;
  assign n40754 = x200 | n40129 ;
  assign n40755 = n40753 | n40754 ;
  assign n40756 = ~n40752 & n40755 ;
  assign n40757 = n14313 | n40756 ;
  assign n40758 = x211 & x1138 ;
  assign n40759 = n40719 | n40758 ;
  assign n40760 = ( x219 & n14313 ) | ( x219 & ~n40759 ) | ( n14313 & ~n40759 ) ;
  assign n40761 = ( x219 & ~n14313 ) | ( x219 & n40171 ) | ( ~n14313 & n40171 ) ;
  assign n40762 = n40760 & ~n40761 ;
  assign n40763 = n40757 & ~n40762 ;
  assign n40764 = x230 & ~n40763 ;
  assign n40765 = x1091 & n40759 ;
  assign n40766 = n36803 & ~n40765 ;
  assign n40767 = x1138 & n37691 ;
  assign n40768 = n40733 | n40767 ;
  assign n40769 = n39983 | n40768 ;
  assign n40770 = ~n40766 & n40769 ;
  assign n40771 = ( ~x830 & x1091 ) | ( ~x830 & n37477 ) | ( x1091 & n37477 ) ;
  assign n40772 = ( x281 & x1091 ) | ( x281 & ~n37477 ) | ( x1091 & ~n37477 ) ;
  assign n40773 = n40771 | n40772 ;
  assign n40774 = ~n40770 & n40773 ;
  assign n40775 = x1139 & n39146 ;
  assign n40776 = n40157 & ~n40775 ;
  assign n40777 = x199 & ~n40178 ;
  assign n40778 = ~n14313 & n40777 ;
  assign n40779 = n40776 | n40778 ;
  assign n40780 = ( ~x830 & x1091 ) | ( ~x830 & n37466 ) | ( x1091 & n37466 ) ;
  assign n40781 = ( x281 & x1091 ) | ( x281 & ~n37466 ) | ( x1091 & ~n37466 ) ;
  assign n40782 = n40780 | n40781 ;
  assign n40783 = n40779 & n40782 ;
  assign n40784 = n40774 | n40783 ;
  assign n40785 = ~x230 & n40784 ;
  assign n40786 = n40764 | n40785 ;
  assign n40787 = x200 & ~n40199 ;
  assign n40788 = x199 & x1140 ;
  assign n40789 = x200 | n40751 ;
  assign n40790 = n40788 | n40789 ;
  assign n40791 = ~n40787 & n40790 ;
  assign n40792 = n14313 | n40791 ;
  assign n40793 = x211 & x1139 ;
  assign n40794 = n40140 | n40793 ;
  assign n40795 = ( x219 & n14313 ) | ( x219 & ~n40794 ) | ( n14313 & ~n40794 ) ;
  assign n40796 = ( x219 & ~n14313 ) | ( x219 & n40577 ) | ( ~n14313 & n40577 ) ;
  assign n40797 = n40795 & ~n40796 ;
  assign n40798 = n40792 & ~n40797 ;
  assign n40799 = x230 & ~n40798 ;
  assign n40800 = x1091 & n40794 ;
  assign n40801 = n36803 & ~n40800 ;
  assign n40802 = x1139 & n37691 ;
  assign n40803 = n40160 | n40802 ;
  assign n40804 = n39983 | n40803 ;
  assign n40805 = ~n40801 & n40804 ;
  assign n40806 = ( ~x836 & x1091 ) | ( ~x836 & n37477 ) | ( x1091 & n37477 ) ;
  assign n40807 = ( x282 & x1091 ) | ( x282 & ~n37477 ) | ( x1091 & ~n37477 ) ;
  assign n40808 = n40806 | n40807 ;
  assign n40809 = ~n40805 & n40808 ;
  assign n40810 = x1140 & n39146 ;
  assign n40811 = n40157 & ~n40810 ;
  assign n40812 = ( x199 & n35214 ) | ( x199 & ~n40176 ) | ( n35214 & ~n40176 ) ;
  assign n40813 = ~n14313 & n40812 ;
  assign n40814 = n40811 | n40813 ;
  assign n40815 = ( ~x836 & x1091 ) | ( ~x836 & n37466 ) | ( x1091 & n37466 ) ;
  assign n40816 = ( x282 & x1091 ) | ( x282 & ~n37466 ) | ( x1091 & ~n37466 ) ;
  assign n40817 = n40815 | n40816 ;
  assign n40818 = n40814 & n40817 ;
  assign n40819 = n40809 | n40818 ;
  assign n40820 = ~x230 & n40819 ;
  assign n40821 = n40799 | n40820 ;
  assign n40822 = x1147 & ~n39984 ;
  assign n40823 = x1149 | n39996 ;
  assign n40824 = n40822 | n40823 ;
  assign n40825 = x1147 & ~n40288 ;
  assign n40826 = n40347 & ~n40825 ;
  assign n40827 = x1148 & ~n40826 ;
  assign n40828 = n40824 & n40827 ;
  assign n40829 = x1149 & n38931 ;
  assign n40830 = n40825 | n40829 ;
  assign n40831 = ~x1148 & n40830 ;
  assign n40832 = x230 & ~n40831 ;
  assign n40833 = ~n40828 & n40832 ;
  assign n40834 = ( x1147 & x1149 ) | ( x1147 & n40084 ) | ( x1149 & n40084 ) ;
  assign n40835 = ( ~x1147 & x1149 ) | ( ~x1147 & n40066 ) | ( x1149 & n40066 ) ;
  assign n40836 = n40834 & n40835 ;
  assign n40837 = x1148 & ~n40836 ;
  assign n40838 = ( x1147 & x1149 ) | ( x1147 & ~n40029 ) | ( x1149 & ~n40029 ) ;
  assign n40839 = ( x1147 & ~x1149 ) | ( x1147 & n40088 ) | ( ~x1149 & n40088 ) ;
  assign n40840 = ~n40838 & n40839 ;
  assign n40841 = n40837 & ~n40840 ;
  assign n40842 = ( x1147 & x1149 ) | ( x1147 & ~n40041 ) | ( x1149 & ~n40041 ) ;
  assign n40843 = ( x1147 & ~x1149 ) | ( x1147 & n40028 ) | ( ~x1149 & n40028 ) ;
  assign n40844 = ~n40842 & n40843 ;
  assign n40845 = x1148 | n40844 ;
  assign n40846 = ( x1147 & x1149 ) | ( x1147 & n40081 ) | ( x1149 & n40081 ) ;
  assign n40847 = ( ~x1147 & x1149 ) | ( ~x1147 & n40070 ) | ( x1149 & n40070 ) ;
  assign n40848 = n40846 & n40847 ;
  assign n40849 = n40845 | n40848 ;
  assign n40850 = ~x283 & n40849 ;
  assign n40851 = ~n40841 & n40850 ;
  assign n40852 = ( x1147 & x1148 ) | ( x1147 & ~n40111 ) | ( x1148 & ~n40111 ) ;
  assign n40853 = ( x1147 & ~x1148 ) | ( x1147 & n40057 ) | ( ~x1148 & n40057 ) ;
  assign n40854 = n40852 & ~n40853 ;
  assign n40855 = x1149 & ~n40854 ;
  assign n40856 = ( x1147 & x1148 ) | ( x1147 & n40052 ) | ( x1148 & n40052 ) ;
  assign n40857 = ( ~x1147 & x1148 ) | ( ~x1147 & n40105 ) | ( x1148 & n40105 ) ;
  assign n40858 = n40856 | n40857 ;
  assign n40859 = n40855 & n40858 ;
  assign n40860 = ( x1147 & x1148 ) | ( x1147 & ~n40096 ) | ( x1148 & ~n40096 ) ;
  assign n40861 = ( x1147 & ~x1148 ) | ( x1147 & n40020 ) | ( ~x1148 & n40020 ) ;
  assign n40862 = n40860 & ~n40861 ;
  assign n40863 = x1149 | n40862 ;
  assign n40864 = ( x1147 & x1148 ) | ( x1147 & n40014 ) | ( x1148 & n40014 ) ;
  assign n40865 = ( ~x1147 & x1148 ) | ( ~x1147 & n40098 ) | ( x1148 & n40098 ) ;
  assign n40866 = n40864 | n40865 ;
  assign n40867 = ~n40863 & n40866 ;
  assign n40868 = x283 & ~n40867 ;
  assign n40869 = ~n40859 & n40868 ;
  assign n40870 = x230 | n40869 ;
  assign n40871 = n40851 | n40870 ;
  assign n40872 = ~n40833 & n40871 ;
  assign n40873 = x284 | n39427 ;
  assign n40874 = x1143 & n39427 ;
  assign n40875 = n36805 & n40874 ;
  assign n40876 = n40873 & ~n40875 ;
  assign n40877 = ~n2033 & n8593 ;
  assign n40878 = ~n6412 & n40877 ;
  assign n40879 = x286 & n40878 ;
  assign n40880 = x288 & x289 ;
  assign n40881 = n40879 & n40880 ;
  assign n40882 = ~n6785 & n40881 ;
  assign n40883 = ~x286 & n6412 ;
  assign n40884 = ~x288 & n40883 ;
  assign n40885 = ~x289 & n40884 ;
  assign n40886 = x285 & ~n40885 ;
  assign n40887 = ~n40882 & n40886 ;
  assign n40888 = x285 & ~n40881 ;
  assign n40889 = n40877 & ~n40881 ;
  assign n40890 = ( x285 & n6785 ) | ( x285 & ~n40889 ) | ( n6785 & ~n40889 ) ;
  assign n40891 = ( n40881 & n40888 ) | ( n40881 & ~n40890 ) | ( n40888 & ~n40890 ) ;
  assign n40892 = n40887 | n40891 ;
  assign n40893 = ~x793 & n40892 ;
  assign n40894 = x286 | n40878 ;
  assign n40895 = x288 & ~n40879 ;
  assign n40896 = n40894 & n40895 ;
  assign n40897 = ~x288 & n6152 ;
  assign n40898 = n6412 & ~n40877 ;
  assign n40899 = x286 & ~n40898 ;
  assign n40900 = ~n40877 & n40883 ;
  assign n40901 = n40899 | n40900 ;
  assign n40902 = n40897 & n40901 ;
  assign n40903 = n6785 | n40902 ;
  assign n40904 = n40896 | n40903 ;
  assign n40905 = n6412 & n40897 ;
  assign n40906 = ~x286 & n40905 ;
  assign n40907 = ( ~x286 & n6785 ) | ( ~x286 & n40905 ) | ( n6785 & n40905 ) ;
  assign n40908 = ( x793 & ~n40906 ) | ( x793 & n40907 ) | ( ~n40906 & n40907 ) ;
  assign n40909 = n40904 & ~n40908 ;
  assign n40910 = ~x287 & x457 ;
  assign n40911 = x332 | n40910 ;
  assign n40912 = ~n6785 & n40877 ;
  assign n40913 = x288 & ~n6412 ;
  assign n40914 = n40905 | n40913 ;
  assign n40915 = ~n40912 & n40914 ;
  assign n40916 = ( x793 & n40914 ) | ( x793 & ~n40915 ) | ( n40914 & ~n40915 ) ;
  assign n40917 = ( n40912 & n40915 ) | ( n40912 & ~n40916 ) | ( n40915 & ~n40916 ) ;
  assign n40918 = x285 & ~x289 ;
  assign n40919 = ( ~n6785 & n40884 ) | ( ~n6785 & n40918 ) | ( n40884 & n40918 ) ;
  assign n40920 = ( ~x289 & n6785 ) | ( ~x289 & n40884 ) | ( n6785 & n40884 ) ;
  assign n40921 = ~n40919 & n40920 ;
  assign n40922 = x793 | n40921 ;
  assign n40923 = ~x289 & n40895 ;
  assign n40924 = ( x288 & n40900 ) | ( x288 & n40918 ) | ( n40900 & n40918 ) ;
  assign n40925 = ( x288 & x289 ) | ( x288 & ~n40900 ) | ( x289 & ~n40900 ) ;
  assign n40926 = n40924 | n40925 ;
  assign n40927 = ~n40923 & n40926 ;
  assign n40928 = ( n6785 & ~n40882 ) | ( n6785 & n40927 ) | ( ~n40882 & n40927 ) ;
  assign n40929 = ~n40922 & n40928 ;
  assign n40930 = ~x290 & x476 ;
  assign n40931 = x476 | x1048 ;
  assign n40932 = ~n40930 & n40931 ;
  assign n40933 = ~x291 & x476 ;
  assign n40934 = x476 | x1049 ;
  assign n40935 = ~n40933 & n40934 ;
  assign n40936 = ~x292 & x476 ;
  assign n40937 = x476 | x1084 ;
  assign n40938 = ~n40936 & n40937 ;
  assign n40939 = ~x293 & x476 ;
  assign n40940 = x476 | x1059 ;
  assign n40941 = ~n40939 & n40940 ;
  assign n40942 = ~x294 & x476 ;
  assign n40943 = x476 | x1072 ;
  assign n40944 = ~n40942 & n40943 ;
  assign n40945 = ~x295 & x476 ;
  assign n40946 = x476 | x1053 ;
  assign n40947 = ~n40945 & n40946 ;
  assign n40948 = ~x296 & x476 ;
  assign n40949 = x476 | x1037 ;
  assign n40950 = ~n40948 & n40949 ;
  assign n40951 = ~x297 & x476 ;
  assign n40952 = x476 | x1044 ;
  assign n40953 = ~n40951 & n40952 ;
  assign n40954 = ~x478 & x1044 ;
  assign n40955 = x298 & x478 ;
  assign n40956 = n40954 | n40955 ;
  assign n40957 = x54 & ~n1868 ;
  assign n40958 = x54 | n11191 ;
  assign n40959 = n11432 & ~n40958 ;
  assign n40960 = n40957 | n40959 ;
  assign n40961 = n2008 | n7112 ;
  assign n40962 = n40960 & ~n40961 ;
  assign n40963 = x39 | n40962 ;
  assign n40964 = ~n9407 & n40963 ;
  assign n40965 = x57 & ~x59 ;
  assign n40966 = ~n8309 & n40965 ;
  assign n40967 = ~x312 & n40966 ;
  assign n40968 = x300 & ~n40967 ;
  assign n40969 = ~x300 & n40967 ;
  assign n40970 = x55 | n40969 ;
  assign n40971 = n40968 | n40970 ;
  assign n40972 = x301 | n40970 ;
  assign n40973 = ~x55 & x301 ;
  assign n40974 = n40969 & n40973 ;
  assign n40975 = n40972 & ~n40974 ;
  assign n40976 = n4353 | n6785 ;
  assign n40977 = ~n4364 & n14313 ;
  assign n40978 = n40976 & ~n40977 ;
  assign n40979 = ~x1148 & n40978 ;
  assign n40980 = x222 | x223 ;
  assign n40981 = x937 & n40980 ;
  assign n40982 = x273 & n1817 ;
  assign n40983 = n40981 | n40982 ;
  assign n40984 = n40976 | n40983 ;
  assign n40985 = ~n2204 & n14313 ;
  assign n40986 = n40984 & ~n40985 ;
  assign n40987 = x237 & ~n40986 ;
  assign n40988 = n1823 & ~n40984 ;
  assign n40989 = ~x215 & n2085 ;
  assign n40990 = ~x273 & n40989 ;
  assign n40991 = x833 & n6433 ;
  assign n40992 = ~x937 & n40991 ;
  assign n40993 = n40990 | n40992 ;
  assign n40994 = n14313 & n40993 ;
  assign n40995 = n40988 | n40994 ;
  assign n40996 = n40987 | n40995 ;
  assign n40997 = n40979 | n40996 ;
  assign n40998 = ~x478 & x1049 ;
  assign n40999 = x303 & x478 ;
  assign n41000 = n40998 | n40999 ;
  assign n41001 = ~x478 & x1048 ;
  assign n41002 = x304 & x478 ;
  assign n41003 = n41001 | n41002 ;
  assign n41004 = ~x478 & x1084 ;
  assign n41005 = x305 & x478 ;
  assign n41006 = n41004 | n41005 ;
  assign n41007 = ~x478 & x1059 ;
  assign n41008 = x306 & x478 ;
  assign n41009 = n41007 | n41008 ;
  assign n41010 = ~x478 & x1053 ;
  assign n41011 = x307 & x478 ;
  assign n41012 = n41010 | n41011 ;
  assign n41013 = ~x478 & x1037 ;
  assign n41014 = x308 & x478 ;
  assign n41015 = n41013 | n41014 ;
  assign n41016 = ~x478 & x1072 ;
  assign n41017 = x309 & x478 ;
  assign n41018 = n41016 | n41017 ;
  assign n41019 = x1147 & n40978 ;
  assign n41020 = n2203 & n40977 ;
  assign n41021 = x934 & n1908 ;
  assign n41022 = x271 & n2085 ;
  assign n41023 = n41021 | n41022 ;
  assign n41024 = n41020 & n41023 ;
  assign n41025 = x222 & ~x934 ;
  assign n41026 = ~x271 & n1817 ;
  assign n41027 = n41025 | n41026 ;
  assign n41028 = n40976 | n41027 ;
  assign n41029 = ~n40985 & n41028 ;
  assign n41030 = ~n41024 & n41029 ;
  assign n41031 = ~n41019 & n41030 ;
  assign n41032 = x233 | n41031 ;
  assign n41033 = n40977 & ~n41023 ;
  assign n41034 = ~n40976 & n41027 ;
  assign n41035 = n1873 | n14313 ;
  assign n41036 = x1147 & n41035 ;
  assign n41037 = ~n41034 & n41036 ;
  assign n41038 = ~n41033 & n41037 ;
  assign n41039 = n1823 & ~n40976 ;
  assign n41040 = n41020 | n41039 ;
  assign n41041 = ~x1147 & n41040 ;
  assign n41042 = ~n41030 & n41041 ;
  assign n41043 = n41038 | n41042 ;
  assign n41044 = x233 & n41043 ;
  assign n41045 = n41032 & ~n41044 ;
  assign n41046 = x55 | x311 ;
  assign n41047 = ~n40974 & n41046 ;
  assign n41048 = ~x311 & n40974 ;
  assign n41049 = n41047 | n41048 ;
  assign n41050 = x312 & ~n40966 ;
  assign n41051 = n40967 | n41050 ;
  assign n41052 = ~x55 & n41051 ;
  assign n41053 = n8582 | n11466 ;
  assign n41054 = n4800 & ~n11472 ;
  assign n41055 = n8332 | n41054 ;
  assign n41056 = n41053 & ~n41055 ;
  assign n41057 = x954 | n41056 ;
  assign n41058 = x313 & x954 ;
  assign n41059 = n41057 & ~n41058 ;
  assign n41060 = n5075 | n7112 ;
  assign n41061 = ~n12404 & n41060 ;
  assign n41062 = ( x39 & n1975 ) | ( x39 & n13214 ) | ( n1975 & n13214 ) ;
  assign n41063 = ( ~x39 & n1975 ) | ( ~x39 & n12461 ) | ( n1975 & n12461 ) ;
  assign n41064 = n41062 | n41063 ;
  assign n41065 = ~n13485 & n41064 ;
  assign n41066 = n2042 | n8329 ;
  assign n41067 = n41065 | n41066 ;
  assign n41068 = ~n41061 & n41067 ;
  assign n41069 = n12396 | n12397 ;
  assign n41070 = n41068 | n41069 ;
  assign n41071 = ~x340 & n40877 ;
  assign n41072 = ~n6785 & n41071 ;
  assign n41073 = x315 & ~n41072 ;
  assign n41074 = x1080 & n41072 ;
  assign n41075 = n41073 | n41074 ;
  assign n41076 = x316 & ~n41072 ;
  assign n41077 = x1047 & n41072 ;
  assign n41078 = n41076 | n41077 ;
  assign n41079 = ~x330 & n40912 ;
  assign n41080 = x317 & ~n41079 ;
  assign n41081 = x1078 & n41079 ;
  assign n41082 = n41080 | n41081 ;
  assign n41083 = ~x341 & n40877 ;
  assign n41084 = ~n6785 & n41083 ;
  assign n41085 = x318 & ~n41084 ;
  assign n41086 = x1074 & n41084 ;
  assign n41087 = n41085 | n41086 ;
  assign n41088 = x319 & ~n41084 ;
  assign n41089 = x1072 & n41084 ;
  assign n41090 = n41088 | n41089 ;
  assign n41091 = x320 & ~n41072 ;
  assign n41092 = x1048 & n41072 ;
  assign n41093 = n41091 | n41092 ;
  assign n41094 = x321 & ~n41072 ;
  assign n41095 = x1058 & n41072 ;
  assign n41096 = n41094 | n41095 ;
  assign n41097 = x322 & ~n41072 ;
  assign n41098 = x1051 & n41072 ;
  assign n41099 = n41097 | n41098 ;
  assign n41100 = x323 & ~n41072 ;
  assign n41101 = x1065 & n41072 ;
  assign n41102 = n41100 | n41101 ;
  assign n41103 = x324 & ~n41084 ;
  assign n41104 = x1086 & n41084 ;
  assign n41105 = n41103 | n41104 ;
  assign n41106 = x325 & ~n41084 ;
  assign n41107 = x1063 & n41084 ;
  assign n41108 = n41106 | n41107 ;
  assign n41109 = x326 & ~n41084 ;
  assign n41110 = x1057 & n41084 ;
  assign n41111 = n41109 | n41110 ;
  assign n41112 = x327 & ~n41072 ;
  assign n41113 = x1040 & n41072 ;
  assign n41114 = n41112 | n41113 ;
  assign n41115 = x328 & ~n41084 ;
  assign n41116 = x1058 & n41084 ;
  assign n41117 = n41115 | n41116 ;
  assign n41118 = x329 & ~n41084 ;
  assign n41119 = x1043 & n41084 ;
  assign n41120 = n41118 | n41119 ;
  assign n41121 = x1092 & ~n1690 ;
  assign n41122 = n6785 & n41121 ;
  assign n41123 = ~x330 & n41122 ;
  assign n41124 = ~n6785 & n41121 ;
  assign n41125 = x330 | n40877 ;
  assign n41126 = ~n41071 & n41125 ;
  assign n41127 = n41124 & ~n41126 ;
  assign n41128 = n41123 | n41127 ;
  assign n41129 = ~x331 & n41122 ;
  assign n41130 = x331 | n40877 ;
  assign n41131 = ~n41083 & n41130 ;
  assign n41132 = n41124 & ~n41131 ;
  assign n41133 = n41129 | n41132 ;
  assign n41134 = n9158 & ~n11209 ;
  assign n41135 = x332 & ~n7777 ;
  assign n41136 = n9158 | n11145 ;
  assign n41137 = ~n5900 & n41136 ;
  assign n41138 = ( x70 & n41135 ) | ( x70 & n41137 ) | ( n41135 & n41137 ) ;
  assign n41139 = n41134 | n41138 ;
  assign n41140 = ~x39 & n41139 ;
  assign n41141 = ( x38 & n1925 ) | ( x38 & n8609 ) | ( n1925 & n8609 ) ;
  assign n41142 = n41140 | n41141 ;
  assign n41143 = ~n34960 & n41142 ;
  assign n41144 = x333 & ~n41084 ;
  assign n41145 = x1040 & n41084 ;
  assign n41146 = n41144 | n41145 ;
  assign n41147 = x334 & ~n41084 ;
  assign n41148 = x1065 & n41084 ;
  assign n41149 = n41147 | n41148 ;
  assign n41150 = x335 & ~n41084 ;
  assign n41151 = x1069 & n41084 ;
  assign n41152 = n41150 | n41151 ;
  assign n41153 = x336 & ~n41079 ;
  assign n41154 = x1070 & n41079 ;
  assign n41155 = n41153 | n41154 ;
  assign n41156 = x337 & ~n41079 ;
  assign n41157 = x1044 & n41079 ;
  assign n41158 = n41156 | n41157 ;
  assign n41159 = x338 & ~n41079 ;
  assign n41160 = x1072 & n41079 ;
  assign n41161 = n41159 | n41160 ;
  assign n41162 = x339 & ~n41079 ;
  assign n41163 = x1086 & n41079 ;
  assign n41164 = n41162 | n41163 ;
  assign n41165 = x340 & n41122 ;
  assign n41166 = ~x331 & n40877 ;
  assign n41167 = x340 | n40877 ;
  assign n41168 = n41124 & n41167 ;
  assign n41169 = ~n41166 & n41168 ;
  assign n41170 = n41165 | n41169 ;
  assign n41171 = x341 | n40912 ;
  assign n41172 = ~n41079 & n41171 ;
  assign n41173 = n41121 & ~n41172 ;
  assign n41174 = x342 & ~n41072 ;
  assign n41175 = x1049 & n41072 ;
  assign n41176 = n41174 | n41175 ;
  assign n41177 = x343 & ~n41072 ;
  assign n41178 = x1062 & n41072 ;
  assign n41179 = n41177 | n41178 ;
  assign n41180 = x344 & ~n41072 ;
  assign n41181 = x1069 & n41072 ;
  assign n41182 = n41180 | n41181 ;
  assign n41183 = x345 & ~n41072 ;
  assign n41184 = x1039 & n41072 ;
  assign n41185 = n41183 | n41184 ;
  assign n41186 = x346 & ~n41072 ;
  assign n41187 = x1067 & n41072 ;
  assign n41188 = n41186 | n41187 ;
  assign n41189 = x347 & ~n41072 ;
  assign n41190 = x1055 & n41072 ;
  assign n41191 = n41189 | n41190 ;
  assign n41192 = x348 & ~n41072 ;
  assign n41193 = x1087 & n41072 ;
  assign n41194 = n41192 | n41193 ;
  assign n41195 = x349 & ~n41072 ;
  assign n41196 = x1043 & n41072 ;
  assign n41197 = n41195 | n41196 ;
  assign n41198 = x350 & ~n41072 ;
  assign n41199 = x1035 & n41072 ;
  assign n41200 = n41198 | n41199 ;
  assign n41201 = x351 & ~n41072 ;
  assign n41202 = x1079 & n41072 ;
  assign n41203 = n41201 | n41202 ;
  assign n41204 = x352 & ~n41072 ;
  assign n41205 = x1078 & n41072 ;
  assign n41206 = n41204 | n41205 ;
  assign n41207 = x353 & ~n41072 ;
  assign n41208 = x1063 & n41072 ;
  assign n41209 = n41207 | n41208 ;
  assign n41210 = x354 & ~n41072 ;
  assign n41211 = x1045 & n41072 ;
  assign n41212 = n41210 | n41211 ;
  assign n41213 = x355 & ~n41072 ;
  assign n41214 = x1084 & n41072 ;
  assign n41215 = n41213 | n41214 ;
  assign n41216 = x356 & ~n41072 ;
  assign n41217 = x1081 & n41072 ;
  assign n41218 = n41216 | n41217 ;
  assign n41219 = x357 & ~n41072 ;
  assign n41220 = x1076 & n41072 ;
  assign n41221 = n41219 | n41220 ;
  assign n41222 = x358 & ~n41072 ;
  assign n41223 = x1071 & n41072 ;
  assign n41224 = n41222 | n41223 ;
  assign n41225 = x359 & ~n41072 ;
  assign n41226 = x1068 & n41072 ;
  assign n41227 = n41225 | n41226 ;
  assign n41228 = x360 & ~n41072 ;
  assign n41229 = x1042 & n41072 ;
  assign n41230 = n41228 | n41229 ;
  assign n41231 = x361 & ~n41072 ;
  assign n41232 = x1059 & n41072 ;
  assign n41233 = n41231 | n41232 ;
  assign n41234 = x362 & ~n41072 ;
  assign n41235 = x1070 & n41072 ;
  assign n41236 = n41234 | n41235 ;
  assign n41237 = x363 & ~n41079 ;
  assign n41238 = x1049 & n41079 ;
  assign n41239 = n41237 | n41238 ;
  assign n41240 = x364 & ~n41079 ;
  assign n41241 = x1062 & n41079 ;
  assign n41242 = n41240 | n41241 ;
  assign n41243 = x365 & ~n41079 ;
  assign n41244 = x1065 & n41079 ;
  assign n41245 = n41243 | n41244 ;
  assign n41246 = x366 & ~n41079 ;
  assign n41247 = x1069 & n41079 ;
  assign n41248 = n41246 | n41247 ;
  assign n41249 = x367 & ~n41079 ;
  assign n41250 = x1039 & n41079 ;
  assign n41251 = n41249 | n41250 ;
  assign n41252 = x368 & ~n41079 ;
  assign n41253 = x1067 & n41079 ;
  assign n41254 = n41252 | n41253 ;
  assign n41255 = x369 & ~n41079 ;
  assign n41256 = x1080 & n41079 ;
  assign n41257 = n41255 | n41256 ;
  assign n41258 = x370 & ~n41079 ;
  assign n41259 = x1055 & n41079 ;
  assign n41260 = n41258 | n41259 ;
  assign n41261 = x371 & ~n41079 ;
  assign n41262 = x1051 & n41079 ;
  assign n41263 = n41261 | n41262 ;
  assign n41264 = x372 & ~n41079 ;
  assign n41265 = x1048 & n41079 ;
  assign n41266 = n41264 | n41265 ;
  assign n41267 = x373 & ~n41079 ;
  assign n41268 = x1087 & n41079 ;
  assign n41269 = n41267 | n41268 ;
  assign n41270 = x374 & ~n41079 ;
  assign n41271 = x1035 & n41079 ;
  assign n41272 = n41270 | n41271 ;
  assign n41273 = x375 & ~n41079 ;
  assign n41274 = x1047 & n41079 ;
  assign n41275 = n41273 | n41274 ;
  assign n41276 = x376 & ~n41079 ;
  assign n41277 = x1079 & n41079 ;
  assign n41278 = n41276 | n41277 ;
  assign n41279 = x377 & ~n41079 ;
  assign n41280 = x1074 & n41079 ;
  assign n41281 = n41279 | n41280 ;
  assign n41282 = x378 & ~n41079 ;
  assign n41283 = x1063 & n41079 ;
  assign n41284 = n41282 | n41283 ;
  assign n41285 = x379 & ~n41079 ;
  assign n41286 = x1045 & n41079 ;
  assign n41287 = n41285 | n41286 ;
  assign n41288 = x380 & ~n41079 ;
  assign n41289 = x1084 & n41079 ;
  assign n41290 = n41288 | n41289 ;
  assign n41291 = x381 & ~n41079 ;
  assign n41292 = x1081 & n41079 ;
  assign n41293 = n41291 | n41292 ;
  assign n41294 = x382 & ~n41079 ;
  assign n41295 = x1076 & n41079 ;
  assign n41296 = n41294 | n41295 ;
  assign n41297 = x383 & ~n41079 ;
  assign n41298 = x1071 & n41079 ;
  assign n41299 = n41297 | n41298 ;
  assign n41300 = x384 & ~n41079 ;
  assign n41301 = x1068 & n41079 ;
  assign n41302 = n41300 | n41301 ;
  assign n41303 = x385 & ~n41079 ;
  assign n41304 = x1042 & n41079 ;
  assign n41305 = n41303 | n41304 ;
  assign n41306 = x386 & ~n41079 ;
  assign n41307 = x1059 & n41079 ;
  assign n41308 = n41306 | n41307 ;
  assign n41309 = x387 & ~n41079 ;
  assign n41310 = x1053 & n41079 ;
  assign n41311 = n41309 | n41310 ;
  assign n41312 = x388 & ~n41079 ;
  assign n41313 = x1037 & n41079 ;
  assign n41314 = n41312 | n41313 ;
  assign n41315 = x389 & ~n41079 ;
  assign n41316 = x1036 & n41079 ;
  assign n41317 = n41315 | n41316 ;
  assign n41318 = x390 & ~n41084 ;
  assign n41319 = x1049 & n41084 ;
  assign n41320 = n41318 | n41319 ;
  assign n41321 = x391 & ~n41084 ;
  assign n41322 = x1062 & n41084 ;
  assign n41323 = n41321 | n41322 ;
  assign n41324 = x392 & ~n41084 ;
  assign n41325 = x1039 & n41084 ;
  assign n41326 = n41324 | n41325 ;
  assign n41327 = x393 & ~n41084 ;
  assign n41328 = x1067 & n41084 ;
  assign n41329 = n41327 | n41328 ;
  assign n41330 = x394 & ~n41084 ;
  assign n41331 = x1080 & n41084 ;
  assign n41332 = n41330 | n41331 ;
  assign n41333 = x395 & ~n41084 ;
  assign n41334 = x1055 & n41084 ;
  assign n41335 = n41333 | n41334 ;
  assign n41336 = x396 & ~n41084 ;
  assign n41337 = x1051 & n41084 ;
  assign n41338 = n41336 | n41337 ;
  assign n41339 = x397 & ~n41084 ;
  assign n41340 = x1048 & n41084 ;
  assign n41341 = n41339 | n41340 ;
  assign n41342 = x398 & ~n41084 ;
  assign n41343 = x1087 & n41084 ;
  assign n41344 = n41342 | n41343 ;
  assign n41345 = x399 & ~n41084 ;
  assign n41346 = x1047 & n41084 ;
  assign n41347 = n41345 | n41346 ;
  assign n41348 = x400 & ~n41084 ;
  assign n41349 = x1035 & n41084 ;
  assign n41350 = n41348 | n41349 ;
  assign n41351 = x401 & ~n41084 ;
  assign n41352 = x1079 & n41084 ;
  assign n41353 = n41351 | n41352 ;
  assign n41354 = x402 & ~n41084 ;
  assign n41355 = x1078 & n41084 ;
  assign n41356 = n41354 | n41355 ;
  assign n41357 = x403 & ~n41084 ;
  assign n41358 = x1045 & n41084 ;
  assign n41359 = n41357 | n41358 ;
  assign n41360 = x404 & ~n41084 ;
  assign n41361 = x1084 & n41084 ;
  assign n41362 = n41360 | n41361 ;
  assign n41363 = x405 & ~n41084 ;
  assign n41364 = x1081 & n41084 ;
  assign n41365 = n41363 | n41364 ;
  assign n41366 = x406 & ~n41084 ;
  assign n41367 = x1076 & n41084 ;
  assign n41368 = n41366 | n41367 ;
  assign n41369 = x407 & ~n41084 ;
  assign n41370 = x1071 & n41084 ;
  assign n41371 = n41369 | n41370 ;
  assign n41372 = x408 & ~n41084 ;
  assign n41373 = x1068 & n41084 ;
  assign n41374 = n41372 | n41373 ;
  assign n41375 = x409 & ~n41084 ;
  assign n41376 = x1042 & n41084 ;
  assign n41377 = n41375 | n41376 ;
  assign n41378 = x410 & ~n41084 ;
  assign n41379 = x1059 & n41084 ;
  assign n41380 = n41378 | n41379 ;
  assign n41381 = x411 & ~n41084 ;
  assign n41382 = x1053 & n41084 ;
  assign n41383 = n41381 | n41382 ;
  assign n41384 = x412 & ~n41084 ;
  assign n41385 = x1037 & n41084 ;
  assign n41386 = n41384 | n41385 ;
  assign n41387 = x413 & ~n41084 ;
  assign n41388 = x1036 & n41084 ;
  assign n41389 = n41387 | n41388 ;
  assign n41390 = ~n6785 & n41166 ;
  assign n41391 = x414 & ~n41390 ;
  assign n41392 = x1049 & n41390 ;
  assign n41393 = n41391 | n41392 ;
  assign n41394 = x415 & ~n41390 ;
  assign n41395 = x1062 & n41390 ;
  assign n41396 = n41394 | n41395 ;
  assign n41397 = x416 & ~n41390 ;
  assign n41398 = x1069 & n41390 ;
  assign n41399 = n41397 | n41398 ;
  assign n41400 = x417 & ~n41390 ;
  assign n41401 = x1039 & n41390 ;
  assign n41402 = n41400 | n41401 ;
  assign n41403 = x418 & ~n41390 ;
  assign n41404 = x1067 & n41390 ;
  assign n41405 = n41403 | n41404 ;
  assign n41406 = x419 & ~n41390 ;
  assign n41407 = x1080 & n41390 ;
  assign n41408 = n41406 | n41407 ;
  assign n41409 = x420 & ~n41390 ;
  assign n41410 = x1055 & n41390 ;
  assign n41411 = n41409 | n41410 ;
  assign n41412 = x421 & ~n41390 ;
  assign n41413 = x1051 & n41390 ;
  assign n41414 = n41412 | n41413 ;
  assign n41415 = x422 & ~n41390 ;
  assign n41416 = x1048 & n41390 ;
  assign n41417 = n41415 | n41416 ;
  assign n41418 = x423 & ~n41390 ;
  assign n41419 = x1087 & n41390 ;
  assign n41420 = n41418 | n41419 ;
  assign n41421 = x424 & ~n41390 ;
  assign n41422 = x1047 & n41390 ;
  assign n41423 = n41421 | n41422 ;
  assign n41424 = x425 & ~n41390 ;
  assign n41425 = x1035 & n41390 ;
  assign n41426 = n41424 | n41425 ;
  assign n41427 = x426 & ~n41390 ;
  assign n41428 = x1079 & n41390 ;
  assign n41429 = n41427 | n41428 ;
  assign n41430 = x427 & ~n41390 ;
  assign n41431 = x1078 & n41390 ;
  assign n41432 = n41430 | n41431 ;
  assign n41433 = x428 & ~n41390 ;
  assign n41434 = x1045 & n41390 ;
  assign n41435 = n41433 | n41434 ;
  assign n41436 = x429 & ~n41390 ;
  assign n41437 = x1084 & n41390 ;
  assign n41438 = n41436 | n41437 ;
  assign n41439 = x430 & ~n41390 ;
  assign n41440 = x1076 & n41390 ;
  assign n41441 = n41439 | n41440 ;
  assign n41442 = x431 & ~n41390 ;
  assign n41443 = x1071 & n41390 ;
  assign n41444 = n41442 | n41443 ;
  assign n41445 = x432 & ~n41390 ;
  assign n41446 = x1068 & n41390 ;
  assign n41447 = n41445 | n41446 ;
  assign n41448 = x433 & ~n41390 ;
  assign n41449 = x1042 & n41390 ;
  assign n41450 = n41448 | n41449 ;
  assign n41451 = x434 & ~n41390 ;
  assign n41452 = x1059 & n41390 ;
  assign n41453 = n41451 | n41452 ;
  assign n41454 = x435 & ~n41390 ;
  assign n41455 = x1053 & n41390 ;
  assign n41456 = n41454 | n41455 ;
  assign n41457 = x436 & ~n41390 ;
  assign n41458 = x1037 & n41390 ;
  assign n41459 = n41457 | n41458 ;
  assign n41460 = x437 & ~n41390 ;
  assign n41461 = x1070 & n41390 ;
  assign n41462 = n41460 | n41461 ;
  assign n41463 = x438 & ~n41390 ;
  assign n41464 = x1036 & n41390 ;
  assign n41465 = n41463 | n41464 ;
  assign n41466 = x439 & ~n41079 ;
  assign n41467 = x1057 & n41079 ;
  assign n41468 = n41466 | n41467 ;
  assign n41469 = x440 & ~n41079 ;
  assign n41470 = x1043 & n41079 ;
  assign n41471 = n41469 | n41470 ;
  assign n41472 = x441 & ~n41072 ;
  assign n41473 = x1044 & n41072 ;
  assign n41474 = n41472 | n41473 ;
  assign n41475 = x442 & ~n41079 ;
  assign n41476 = x1058 & n41079 ;
  assign n41477 = n41475 | n41476 ;
  assign n41478 = x443 & ~n41390 ;
  assign n41479 = x1044 & n41390 ;
  assign n41480 = n41478 | n41479 ;
  assign n41481 = x444 & ~n41390 ;
  assign n41482 = x1072 & n41390 ;
  assign n41483 = n41481 | n41482 ;
  assign n41484 = x445 & ~n41390 ;
  assign n41485 = x1081 & n41390 ;
  assign n41486 = n41484 | n41485 ;
  assign n41487 = x446 & ~n41390 ;
  assign n41488 = x1086 & n41390 ;
  assign n41489 = n41487 | n41488 ;
  assign n41490 = x447 & ~n41079 ;
  assign n41491 = x1040 & n41079 ;
  assign n41492 = n41490 | n41491 ;
  assign n41493 = x448 & ~n41390 ;
  assign n41494 = x1074 & n41390 ;
  assign n41495 = n41493 | n41494 ;
  assign n41496 = x449 & ~n41390 ;
  assign n41497 = x1057 & n41390 ;
  assign n41498 = n41496 | n41497 ;
  assign n41499 = x450 & ~n41072 ;
  assign n41500 = x1036 & n41072 ;
  assign n41501 = n41499 | n41500 ;
  assign n41502 = x451 & ~n41390 ;
  assign n41503 = x1063 & n41390 ;
  assign n41504 = n41502 | n41503 ;
  assign n41505 = x452 & ~n41072 ;
  assign n41506 = x1053 & n41072 ;
  assign n41507 = n41505 | n41506 ;
  assign n41508 = x453 & ~n41390 ;
  assign n41509 = x1040 & n41390 ;
  assign n41510 = n41508 | n41509 ;
  assign n41511 = x454 & ~n41390 ;
  assign n41512 = x1043 & n41390 ;
  assign n41513 = n41511 | n41512 ;
  assign n41514 = x455 & ~n41072 ;
  assign n41515 = x1037 & n41072 ;
  assign n41516 = n41514 | n41515 ;
  assign n41517 = x456 & ~n41084 ;
  assign n41518 = x1044 & n41084 ;
  assign n41519 = n41517 | n41518 ;
  assign n41520 = x594 & x600 ;
  assign n41521 = x597 & n41520 ;
  assign n41522 = x601 & n41521 ;
  assign n41523 = x804 | x810 ;
  assign n41524 = x595 | n41523 ;
  assign n41525 = ~x599 & x810 ;
  assign n41526 = x596 & ~n41525 ;
  assign n41527 = x804 & ~n41526 ;
  assign n41528 = x595 & x815 ;
  assign n41529 = ~n41527 & n41528 ;
  assign n41530 = n41524 & ~n41529 ;
  assign n41531 = n41522 & ~n41530 ;
  assign n41532 = ~x601 & n41523 ;
  assign n41533 = x600 & ~x810 ;
  assign n41534 = x804 & ~n41533 ;
  assign n41535 = x815 | n41534 ;
  assign n41536 = n41532 | n41535 ;
  assign n41537 = ~n41531 & n41536 ;
  assign n41538 = x605 & ~n41537 ;
  assign n41539 = x990 & n41520 ;
  assign n41540 = ~x815 & n41534 ;
  assign n41541 = n41539 & n41540 ;
  assign n41542 = n41538 | n41541 ;
  assign n41543 = x821 & n41542 ;
  assign n41544 = x458 & ~n41072 ;
  assign n41545 = x1072 & n41072 ;
  assign n41546 = n41544 | n41545 ;
  assign n41547 = x459 & ~n41390 ;
  assign n41548 = x1058 & n41390 ;
  assign n41549 = n41547 | n41548 ;
  assign n41550 = x460 & ~n41072 ;
  assign n41551 = x1086 & n41072 ;
  assign n41552 = n41550 | n41551 ;
  assign n41553 = x461 & ~n41072 ;
  assign n41554 = x1057 & n41072 ;
  assign n41555 = n41553 | n41554 ;
  assign n41556 = x462 & ~n41072 ;
  assign n41557 = x1074 & n41072 ;
  assign n41558 = n41556 | n41557 ;
  assign n41559 = x463 & ~n41084 ;
  assign n41560 = x1070 & n41084 ;
  assign n41561 = n41559 | n41560 ;
  assign n41562 = x464 & ~n41390 ;
  assign n41563 = x1065 & n41390 ;
  assign n41564 = n41562 | n41563 ;
  assign n41565 = n9531 | n9534 ;
  assign n41566 = ~x243 & n41565 ;
  assign n41567 = x299 | n40980 ;
  assign n41568 = ~n9558 & n41567 ;
  assign n41569 = ~x243 & x1157 ;
  assign n41570 = n41568 | n41569 ;
  assign n41571 = n41566 | n41570 ;
  assign n41572 = n2214 & ~n9559 ;
  assign n41573 = x926 & n41569 ;
  assign n41574 = ~n41572 & n41573 ;
  assign n41575 = n41571 & ~n41574 ;
  assign n41576 = ~n4344 & n4353 ;
  assign n41577 = ( x1157 & n41566 ) | ( x1157 & n41576 ) | ( n41566 & n41576 ) ;
  assign n41578 = ( x926 & n41566 ) | ( x926 & ~n41576 ) | ( n41566 & ~n41576 ) ;
  assign n41579 = n41577 | n41578 ;
  assign n41580 = n41575 & n41579 ;
  assign n41581 = n6785 | n41580 ;
  assign n41582 = ~x243 & n40989 ;
  assign n41583 = n6785 & ~n41582 ;
  assign n41584 = x926 & n40991 ;
  assign n41585 = x1157 & n4364 ;
  assign n41586 = n41584 | n41585 ;
  assign n41587 = n41583 & ~n41586 ;
  assign n41588 = n41581 & ~n41587 ;
  assign n41589 = n6785 & ~n40989 ;
  assign n41590 = n6785 | n41565 ;
  assign n41591 = ~n41589 & n41590 ;
  assign n41592 = x943 | n41591 ;
  assign n41593 = x943 & ~n41040 ;
  assign n41594 = n41592 & ~n41593 ;
  assign n41595 = x1151 | n41594 ;
  assign n41596 = ~n40985 & n41035 ;
  assign n41597 = x943 & x1151 ;
  assign n41598 = ~n41596 & n41597 ;
  assign n41599 = n40978 | n41592 ;
  assign n41600 = n6785 | n41568 ;
  assign n41601 = ~n1908 & n6785 ;
  assign n41602 = n41600 & ~n41601 ;
  assign n41603 = x275 | n41602 ;
  assign n41604 = n41599 & n41603 ;
  assign n41605 = ~n41598 & n41604 ;
  assign n41606 = n41595 & n41605 ;
  assign n41607 = x40 & ~x287 ;
  assign n41608 = n38888 & n41607 ;
  assign n41609 = ~n35076 & n41608 ;
  assign n41610 = n8331 & ~n41609 ;
  assign n41611 = x102 | n11404 ;
  assign n41612 = n7130 | n8328 ;
  assign n41613 = n14716 | n41612 ;
  assign n41614 = n41611 & ~n41613 ;
  assign n41615 = ~n14726 & n41614 ;
  assign n41616 = n41608 & ~n41615 ;
  assign n41617 = ~n41608 & n41615 ;
  assign n41618 = n41616 | n41617 ;
  assign n41619 = ~n4799 & n41618 ;
  assign n41620 = n4799 & n41615 ;
  assign n41621 = n41619 | n41620 ;
  assign n41622 = ~x1093 & n41621 ;
  assign n41623 = x1091 | n41622 ;
  assign n41624 = ( x1093 & ~n5950 ) | ( x1093 & n41615 ) | ( ~n5950 & n41615 ) ;
  assign n41625 = ( x1093 & n5950 ) | ( x1093 & n41618 ) | ( n5950 & n41618 ) ;
  assign n41626 = n41624 & n41625 ;
  assign n41627 = n41623 | n41626 ;
  assign n41628 = ( ~x1091 & n5997 ) | ( ~x1091 & n41618 ) | ( n5997 & n41618 ) ;
  assign n41629 = ( x1091 & n5997 ) | ( x1091 & ~n41621 ) | ( n5997 & ~n41621 ) ;
  assign n41630 = ~n41628 & n41629 ;
  assign n41631 = n41627 & ~n41630 ;
  assign n41632 = n1984 | n41060 ;
  assign n41633 = n41631 | n41632 ;
  assign n41634 = ~n41610 & n41633 ;
  assign n41635 = ~n8366 & n9477 ;
  assign n41636 = n1919 & ~n8359 ;
  assign n41637 = ~n7192 & n41636 ;
  assign n41638 = x468 & ~n41637 ;
  assign n41639 = n41635 | n41638 ;
  assign n41640 = ~x263 & n41565 ;
  assign n41641 = ~x263 & x1156 ;
  assign n41642 = n41568 | n41641 ;
  assign n41643 = n41640 | n41642 ;
  assign n41644 = x942 & n41641 ;
  assign n41645 = ~n41572 & n41644 ;
  assign n41646 = n41643 & ~n41645 ;
  assign n41647 = ( x1156 & n41576 ) | ( x1156 & n41640 ) | ( n41576 & n41640 ) ;
  assign n41648 = ( x942 & ~n41576 ) | ( x942 & n41640 ) | ( ~n41576 & n41640 ) ;
  assign n41649 = n41647 | n41648 ;
  assign n41650 = n41646 & n41649 ;
  assign n41651 = n6785 | n41650 ;
  assign n41652 = ~x263 & n40989 ;
  assign n41653 = n6785 & ~n41652 ;
  assign n41654 = x1156 & n4364 ;
  assign n41655 = x942 & n40991 ;
  assign n41656 = n41654 | n41655 ;
  assign n41657 = n41653 & ~n41656 ;
  assign n41658 = n41651 & ~n41657 ;
  assign n41659 = x267 & n41565 ;
  assign n41660 = x267 & x1155 ;
  assign n41661 = n41568 | n41660 ;
  assign n41662 = n41659 | n41661 ;
  assign n41663 = x925 & n41660 ;
  assign n41664 = ~n41572 & n41663 ;
  assign n41665 = n41662 & ~n41664 ;
  assign n41666 = ( x1155 & n41576 ) | ( x1155 & n41659 ) | ( n41576 & n41659 ) ;
  assign n41667 = ( x925 & ~n41576 ) | ( x925 & n41659 ) | ( ~n41576 & n41659 ) ;
  assign n41668 = n41666 | n41667 ;
  assign n41669 = n41665 & n41668 ;
  assign n41670 = n6785 | n41669 ;
  assign n41671 = x267 & n40989 ;
  assign n41672 = n6785 & ~n41671 ;
  assign n41673 = x1155 & n4364 ;
  assign n41674 = x925 & n40991 ;
  assign n41675 = n41673 | n41674 ;
  assign n41676 = n41672 & ~n41675 ;
  assign n41677 = n41670 & ~n41676 ;
  assign n41678 = x253 & n41565 ;
  assign n41679 = x253 & x1153 ;
  assign n41680 = n41568 | n41679 ;
  assign n41681 = n41678 | n41680 ;
  assign n41682 = x941 & n41679 ;
  assign n41683 = ~n41572 & n41682 ;
  assign n41684 = n41681 & ~n41683 ;
  assign n41685 = ( x1153 & n41576 ) | ( x1153 & n41678 ) | ( n41576 & n41678 ) ;
  assign n41686 = ( x941 & ~n41576 ) | ( x941 & n41678 ) | ( ~n41576 & n41678 ) ;
  assign n41687 = n41685 | n41686 ;
  assign n41688 = n41684 & n41687 ;
  assign n41689 = n6785 | n41688 ;
  assign n41690 = x253 & n40989 ;
  assign n41691 = n6785 & ~n41690 ;
  assign n41692 = x1153 & n4364 ;
  assign n41693 = x941 & n40991 ;
  assign n41694 = n41692 | n41693 ;
  assign n41695 = n41691 & ~n41694 ;
  assign n41696 = n41689 & ~n41695 ;
  assign n41697 = x254 & n41565 ;
  assign n41698 = n39232 | n41568 ;
  assign n41699 = n41697 | n41698 ;
  assign n41700 = x923 & n39232 ;
  assign n41701 = ~n41572 & n41700 ;
  assign n41702 = n41699 & ~n41701 ;
  assign n41703 = ( x1154 & n41576 ) | ( x1154 & n41697 ) | ( n41576 & n41697 ) ;
  assign n41704 = ( x923 & ~n41576 ) | ( x923 & n41697 ) | ( ~n41576 & n41697 ) ;
  assign n41705 = n41703 | n41704 ;
  assign n41706 = n41702 & n41705 ;
  assign n41707 = n6785 | n41706 ;
  assign n41708 = x254 & n40989 ;
  assign n41709 = n6785 & ~n41708 ;
  assign n41710 = x1154 & n4364 ;
  assign n41711 = x923 & n40991 ;
  assign n41712 = n41710 | n41711 ;
  assign n41713 = n41709 & ~n41712 ;
  assign n41714 = n41707 & ~n41713 ;
  assign n41715 = x922 | n41591 ;
  assign n41716 = x922 & ~n41040 ;
  assign n41717 = n41715 & ~n41716 ;
  assign n41718 = x1152 | n41717 ;
  assign n41719 = x922 & x1152 ;
  assign n41720 = ~n41596 & n41719 ;
  assign n41721 = n40978 | n41715 ;
  assign n41722 = x268 | n41602 ;
  assign n41723 = n41721 & n41722 ;
  assign n41724 = ~n41720 & n41723 ;
  assign n41725 = n41718 & n41724 ;
  assign n41726 = x931 | n41591 ;
  assign n41727 = x931 & ~n41040 ;
  assign n41728 = n41726 & ~n41727 ;
  assign n41729 = x1150 | n41728 ;
  assign n41730 = x931 & x1150 ;
  assign n41731 = ~n41596 & n41730 ;
  assign n41732 = n40978 | n41726 ;
  assign n41733 = x272 | n41602 ;
  assign n41734 = n41732 & n41733 ;
  assign n41735 = ~n41731 & n41734 ;
  assign n41736 = n41729 & n41735 ;
  assign n41737 = x936 | n41591 ;
  assign n41738 = x936 & ~n41040 ;
  assign n41739 = n41737 & ~n41738 ;
  assign n41740 = x1149 | n41739 ;
  assign n41741 = x936 & x1149 ;
  assign n41742 = ~n41596 & n41741 ;
  assign n41743 = n40978 | n41737 ;
  assign n41744 = x283 | n41602 ;
  assign n41745 = n41743 & n41744 ;
  assign n41746 = ~n41742 & n41745 ;
  assign n41747 = n41740 & n41746 ;
  assign n41748 = x71 & n39995 ;
  assign n41749 = x71 & n9582 ;
  assign n41750 = n9582 | n11091 ;
  assign n41751 = ~n8317 & n9582 ;
  assign n41752 = ~n8313 & n41751 ;
  assign n41753 = n41750 & ~n41752 ;
  assign n41754 = n2033 | n8328 ;
  assign n41755 = n41753 | n41754 ;
  assign n41756 = n11095 & ~n41755 ;
  assign n41757 = n41749 | n41756 ;
  assign n41758 = ~n6785 & n41757 ;
  assign n41759 = n41748 | n41758 ;
  assign n41760 = x71 & ~n40288 ;
  assign n41761 = x481 & ~n31572 ;
  assign n41762 = x248 & n31572 ;
  assign n41763 = n41761 | n41762 ;
  assign n41764 = x482 & ~n31751 ;
  assign n41765 = x249 & n31751 ;
  assign n41766 = n41764 | n41765 ;
  assign n41767 = x483 & ~n31866 ;
  assign n41768 = x242 & n31866 ;
  assign n41769 = n41767 | n41768 ;
  assign n41770 = x484 & ~n31866 ;
  assign n41771 = x249 & n31866 ;
  assign n41772 = n41770 | n41771 ;
  assign n41773 = x485 & ~n32963 ;
  assign n41774 = x234 & n32963 ;
  assign n41775 = n41773 | n41774 ;
  assign n41776 = x486 & ~n32963 ;
  assign n41777 = x244 & n32963 ;
  assign n41778 = n41776 | n41777 ;
  assign n41779 = x487 & ~n31572 ;
  assign n41780 = x246 & n31572 ;
  assign n41781 = n41779 | n41780 ;
  assign n41782 = x488 & ~n31572 ;
  assign n41783 = ~x239 & n31572 ;
  assign n41784 = n41782 | n41783 ;
  assign n41785 = x489 & ~n32963 ;
  assign n41786 = x242 & n32963 ;
  assign n41787 = n41785 | n41786 ;
  assign n41788 = x490 & ~n31866 ;
  assign n41789 = x241 & n31866 ;
  assign n41790 = n41788 | n41789 ;
  assign n41791 = x491 & ~n31866 ;
  assign n41792 = x238 & n31866 ;
  assign n41793 = n41791 | n41792 ;
  assign n41794 = x492 & ~n31866 ;
  assign n41795 = x240 & n31866 ;
  assign n41796 = n41794 | n41795 ;
  assign n41797 = x493 & ~n31866 ;
  assign n41798 = x244 & n31866 ;
  assign n41799 = n41797 | n41798 ;
  assign n41800 = x494 & ~n31866 ;
  assign n41801 = ~x239 & n31866 ;
  assign n41802 = n41800 | n41801 ;
  assign n41803 = x495 & ~n31866 ;
  assign n41804 = x235 & n31866 ;
  assign n41805 = n41803 | n41804 ;
  assign n41806 = x496 & ~n31859 ;
  assign n41807 = x249 & n31859 ;
  assign n41808 = n41806 | n41807 ;
  assign n41809 = x497 & ~n31859 ;
  assign n41810 = ~x239 & n31859 ;
  assign n41811 = n41809 | n41810 ;
  assign n41812 = x498 & ~n31751 ;
  assign n41813 = x238 & n31751 ;
  assign n41814 = n41812 | n41813 ;
  assign n41815 = x499 & ~n31859 ;
  assign n41816 = x246 & n31859 ;
  assign n41817 = n41815 | n41816 ;
  assign n41818 = x500 & ~n31859 ;
  assign n41819 = x241 & n31859 ;
  assign n41820 = n41818 | n41819 ;
  assign n41821 = x501 & ~n31859 ;
  assign n41822 = x248 & n31859 ;
  assign n41823 = n41821 | n41822 ;
  assign n41824 = x502 & ~n31859 ;
  assign n41825 = x247 & n31859 ;
  assign n41826 = n41824 | n41825 ;
  assign n41827 = x503 & ~n31859 ;
  assign n41828 = x245 & n31859 ;
  assign n41829 = n41827 | n41828 ;
  assign n41830 = x504 & ~n31762 ;
  assign n41831 = x242 & n31762 ;
  assign n41832 = n41830 | n41831 ;
  assign n41833 = ~n31757 & n31759 ;
  assign n41834 = ~x234 & n41833 ;
  assign n41835 = n31859 & n41834 ;
  assign n41836 = x505 & ~n41835 ;
  assign n41837 = x234 & n31761 ;
  assign n41838 = ~x505 & n31743 ;
  assign n41839 = n41837 & n41838 ;
  assign n41840 = n41836 | n41839 ;
  assign n41841 = x506 & ~n31762 ;
  assign n41842 = x241 & n31762 ;
  assign n41843 = n41841 | n41842 ;
  assign n41844 = x507 & ~n31762 ;
  assign n41845 = x238 & n31762 ;
  assign n41846 = n41844 | n41845 ;
  assign n41847 = x508 & ~n31762 ;
  assign n41848 = x247 & n31762 ;
  assign n41849 = n41847 | n41848 ;
  assign n41850 = x509 & ~n31762 ;
  assign n41851 = x245 & n31762 ;
  assign n41852 = n41850 | n41851 ;
  assign n41853 = x510 & ~n31572 ;
  assign n41854 = x242 & n31572 ;
  assign n41855 = n41853 | n41854 ;
  assign n41856 = n5134 | n6785 ;
  assign n41857 = ~n31566 & n41856 ;
  assign n41858 = ~x234 & n41857 ;
  assign n41859 = n31572 & ~n41858 ;
  assign n41860 = x511 & ~n31572 ;
  assign n41861 = n41859 | n41860 ;
  assign n41862 = x512 & ~n31572 ;
  assign n41863 = x235 & n31572 ;
  assign n41864 = n41862 | n41863 ;
  assign n41865 = x513 & ~n31572 ;
  assign n41866 = x244 & n31572 ;
  assign n41867 = n41865 | n41866 ;
  assign n41868 = x514 & ~n31572 ;
  assign n41869 = x245 & n31572 ;
  assign n41870 = n41868 | n41869 ;
  assign n41871 = x515 & ~n31572 ;
  assign n41872 = x240 & n31572 ;
  assign n41873 = n41871 | n41872 ;
  assign n41874 = x516 & ~n31572 ;
  assign n41875 = x247 & n31572 ;
  assign n41876 = n41874 | n41875 ;
  assign n41877 = x517 & ~n31572 ;
  assign n41878 = x238 & n31572 ;
  assign n41879 = n41877 | n41878 ;
  assign n41880 = n31744 & n41858 ;
  assign n41881 = x518 & ~n41880 ;
  assign n41882 = x234 & n31571 ;
  assign n41883 = ~x518 & n31743 ;
  assign n41884 = n41882 & n41883 ;
  assign n41885 = n41881 | n41884 ;
  assign n41886 = x519 & ~n31744 ;
  assign n41887 = ~x239 & n31744 ;
  assign n41888 = n41886 | n41887 ;
  assign n41889 = x520 & ~n31744 ;
  assign n41890 = x246 & n31744 ;
  assign n41891 = n41889 | n41890 ;
  assign n41892 = x521 & ~n31744 ;
  assign n41893 = x248 & n31744 ;
  assign n41894 = n41892 | n41893 ;
  assign n41895 = x522 & ~n31744 ;
  assign n41896 = x238 & n31744 ;
  assign n41897 = n41895 | n41896 ;
  assign n41898 = n32987 & n41858 ;
  assign n41899 = x523 & ~n41898 ;
  assign n41900 = ~x523 & n31865 ;
  assign n41901 = n41882 & n41900 ;
  assign n41902 = n41899 | n41901 ;
  assign n41903 = x524 & ~n32987 ;
  assign n41904 = ~x239 & n32987 ;
  assign n41905 = n41903 | n41904 ;
  assign n41906 = x525 & ~n32987 ;
  assign n41907 = x245 & n32987 ;
  assign n41908 = n41906 | n41907 ;
  assign n41909 = x526 & ~n32987 ;
  assign n41910 = x246 & n32987 ;
  assign n41911 = n41909 | n41910 ;
  assign n41912 = x527 & ~n32987 ;
  assign n41913 = x247 & n32987 ;
  assign n41914 = n41912 | n41913 ;
  assign n41915 = x528 & ~n32987 ;
  assign n41916 = x249 & n32987 ;
  assign n41917 = n41915 | n41916 ;
  assign n41918 = x529 & ~n32987 ;
  assign n41919 = x238 & n32987 ;
  assign n41920 = n41918 | n41919 ;
  assign n41921 = x530 & ~n32987 ;
  assign n41922 = x240 & n32987 ;
  assign n41923 = n41921 | n41922 ;
  assign n41924 = x531 & ~n31751 ;
  assign n41925 = x235 & n31751 ;
  assign n41926 = n41924 | n41925 ;
  assign n41927 = x532 & ~n31751 ;
  assign n41928 = x247 & n31751 ;
  assign n41929 = n41927 | n41928 ;
  assign n41930 = x533 & ~n31762 ;
  assign n41931 = x235 & n31762 ;
  assign n41932 = n41930 | n41931 ;
  assign n41933 = x534 & ~n31762 ;
  assign n41934 = ~x239 & n31762 ;
  assign n41935 = n41933 | n41934 ;
  assign n41936 = x535 & ~n31762 ;
  assign n41937 = x240 & n31762 ;
  assign n41938 = n41936 | n41937 ;
  assign n41939 = x536 & ~n31762 ;
  assign n41940 = x246 & n31762 ;
  assign n41941 = n41939 | n41940 ;
  assign n41942 = x537 & ~n31762 ;
  assign n41943 = x248 & n31762 ;
  assign n41944 = n41942 | n41943 ;
  assign n41945 = x538 & ~n31762 ;
  assign n41946 = x249 & n31762 ;
  assign n41947 = n41945 | n41946 ;
  assign n41948 = x539 & ~n31859 ;
  assign n41949 = x242 & n31859 ;
  assign n41950 = n41948 | n41949 ;
  assign n41951 = x540 & ~n31859 ;
  assign n41952 = x235 & n31859 ;
  assign n41953 = n41951 | n41952 ;
  assign n41954 = x541 & ~n31859 ;
  assign n41955 = x244 & n31859 ;
  assign n41956 = n41954 | n41955 ;
  assign n41957 = x542 & ~n31859 ;
  assign n41958 = x240 & n31859 ;
  assign n41959 = n41957 | n41958 ;
  assign n41960 = x543 & ~n31859 ;
  assign n41961 = x238 & n31859 ;
  assign n41962 = n41960 | n41961 ;
  assign n41963 = n31866 & n41834 ;
  assign n41964 = x544 & ~n41963 ;
  assign n41965 = ~x544 & n31865 ;
  assign n41966 = n41837 & n41965 ;
  assign n41967 = n41964 | n41966 ;
  assign n41968 = x545 & ~n31866 ;
  assign n41969 = x245 & n31866 ;
  assign n41970 = n41968 | n41969 ;
  assign n41971 = x546 & ~n31866 ;
  assign n41972 = x246 & n31866 ;
  assign n41973 = n41971 | n41972 ;
  assign n41974 = x547 & ~n31866 ;
  assign n41975 = x247 & n31866 ;
  assign n41976 = n41974 | n41975 ;
  assign n41977 = x548 & ~n31866 ;
  assign n41978 = x248 & n31866 ;
  assign n41979 = n41977 | n41978 ;
  assign n41980 = x549 & ~n32963 ;
  assign n41981 = x235 & n32963 ;
  assign n41982 = n41980 | n41981 ;
  assign n41983 = x550 & ~n32963 ;
  assign n41984 = ~x239 & n32963 ;
  assign n41985 = n41983 | n41984 ;
  assign n41986 = x551 & ~n32963 ;
  assign n41987 = x240 & n32963 ;
  assign n41988 = n41986 | n41987 ;
  assign n41989 = x552 & ~n32963 ;
  assign n41990 = x247 & n32963 ;
  assign n41991 = n41989 | n41990 ;
  assign n41992 = x553 & ~n32963 ;
  assign n41993 = x241 & n32963 ;
  assign n41994 = n41992 | n41993 ;
  assign n41995 = x554 & ~n32963 ;
  assign n41996 = x248 & n32963 ;
  assign n41997 = n41995 | n41996 ;
  assign n41998 = x555 & ~n32963 ;
  assign n41999 = x249 & n32963 ;
  assign n42000 = n41998 | n41999 ;
  assign n42001 = x556 & ~n31751 ;
  assign n42002 = x242 & n31751 ;
  assign n42003 = n42001 | n42002 ;
  assign n42004 = n31762 & n41834 ;
  assign n42005 = x557 & ~n42004 ;
  assign n42006 = ~x557 & n31563 ;
  assign n42007 = n41837 & n42006 ;
  assign n42008 = n42005 | n42007 ;
  assign n42009 = x558 & ~n31762 ;
  assign n42010 = x244 & n31762 ;
  assign n42011 = n42009 | n42010 ;
  assign n42012 = x559 & ~n31572 ;
  assign n42013 = x241 & n31572 ;
  assign n42014 = n42012 | n42013 ;
  assign n42015 = x560 & ~n31751 ;
  assign n42016 = x240 & n31751 ;
  assign n42017 = n42015 | n42016 ;
  assign n42018 = x561 & ~n31744 ;
  assign n42019 = x247 & n31744 ;
  assign n42020 = n42018 | n42019 ;
  assign n42021 = x562 & ~n31751 ;
  assign n42022 = x241 & n31751 ;
  assign n42023 = n42021 | n42022 ;
  assign n42024 = x563 & ~n32963 ;
  assign n42025 = x246 & n32963 ;
  assign n42026 = n42024 | n42025 ;
  assign n42027 = x564 & ~n31751 ;
  assign n42028 = x246 & n31751 ;
  assign n42029 = n42027 | n42028 ;
  assign n42030 = x565 & ~n31751 ;
  assign n42031 = x248 & n31751 ;
  assign n42032 = n42030 | n42031 ;
  assign n42033 = x566 & ~n31751 ;
  assign n42034 = x244 & n31751 ;
  assign n42035 = n42033 | n42034 ;
  assign n42036 = ~x567 & x1092 ;
  assign n42037 = ~x1093 & n42036 ;
  assign n42038 = x680 & n15313 ;
  assign n42039 = ~n17210 & n42038 ;
  assign n42040 = n42037 | n42039 ;
  assign n42041 = ~n17215 & n42040 ;
  assign n42042 = ~n17220 & n42041 ;
  assign n42043 = x647 & n42042 ;
  assign n42044 = x1157 & ~n42037 ;
  assign n42045 = ~n42043 & n42044 ;
  assign n42046 = x630 | n42045 ;
  assign n42047 = x603 & ~n15082 ;
  assign n42048 = n14959 & ~n18257 ;
  assign n42049 = ~n18249 & n42048 ;
  assign n42050 = n42047 & n42049 ;
  assign n42051 = x789 | n42037 ;
  assign n42052 = n42050 | n42051 ;
  assign n42053 = x619 & n42050 ;
  assign n42054 = n42037 | n42053 ;
  assign n42055 = ( ~x789 & x1159 ) | ( ~x789 & n42054 ) | ( x1159 & n42054 ) ;
  assign n42056 = ~x619 & n42050 ;
  assign n42057 = n42037 | n42056 ;
  assign n42058 = ( x789 & x1159 ) | ( x789 & ~n42057 ) | ( x1159 & ~n42057 ) ;
  assign n42059 = ~n42055 & n42058 ;
  assign n42060 = n42052 & ~n42059 ;
  assign n42061 = ~n16176 & n42060 ;
  assign n42062 = n16176 & n42037 ;
  assign n42063 = n42061 | n42062 ;
  assign n42064 = ~n15134 & n42063 ;
  assign n42065 = n15134 & n42037 ;
  assign n42066 = n42064 | n42065 ;
  assign n42067 = ( x647 & x1157 ) | ( x647 & n42066 ) | ( x1157 & n42066 ) ;
  assign n42068 = ~n17214 & n42040 ;
  assign n42069 = n15413 & n42059 ;
  assign n42070 = n42068 & ~n42069 ;
  assign n42071 = n42060 | n42070 ;
  assign n42072 = ~n16177 & n42071 ;
  assign n42073 = n32151 & n42060 ;
  assign n42074 = ~n15414 & n42068 ;
  assign n42075 = x641 & n42074 ;
  assign n42076 = n42037 | n42075 ;
  assign n42077 = n16109 & n42076 ;
  assign n42078 = ~x641 & n42074 ;
  assign n42079 = n42037 | n42078 ;
  assign n42080 = n16110 & n42079 ;
  assign n42081 = n42077 | n42080 ;
  assign n42082 = n42073 | n42081 ;
  assign n42083 = x788 & n42082 ;
  assign n42084 = n42072 | n42083 ;
  assign n42085 = ~n18434 & n42084 ;
  assign n42086 = n16051 & n42063 ;
  assign n42087 = ~x628 & n42041 ;
  assign n42088 = n42037 | n42087 ;
  assign n42089 = ~x1156 & n42088 ;
  assign n42090 = x629 & ~n42089 ;
  assign n42091 = ~n42086 & n42090 ;
  assign n42092 = n16052 & n42063 ;
  assign n42093 = x628 & n42041 ;
  assign n42094 = n42037 | n42093 ;
  assign n42095 = x1156 & n42094 ;
  assign n42096 = x629 | n42095 ;
  assign n42097 = n42092 | n42096 ;
  assign n42098 = x792 & n42097 ;
  assign n42099 = ~n42091 & n42098 ;
  assign n42100 = n42085 | n42099 ;
  assign n42101 = ( ~x647 & x1157 ) | ( ~x647 & n42100 ) | ( x1157 & n42100 ) ;
  assign n42102 = n42067 | n42101 ;
  assign n42103 = ~n42046 & n42102 ;
  assign n42104 = ~x647 & n42042 ;
  assign n42105 = x1157 | n42037 ;
  assign n42106 = n42104 | n42105 ;
  assign n42107 = x630 & n42106 ;
  assign n42108 = ( x647 & x1157 ) | ( x647 & ~n42066 ) | ( x1157 & ~n42066 ) ;
  assign n42109 = ( x647 & ~x1157 ) | ( x647 & n42100 ) | ( ~x1157 & n42100 ) ;
  assign n42110 = n42108 & ~n42109 ;
  assign n42111 = n42107 & ~n42110 ;
  assign n42112 = n42103 | n42111 ;
  assign n42113 = x787 & n42112 ;
  assign n42114 = ~x787 & n42100 ;
  assign n42115 = n42113 | n42114 ;
  assign n42116 = ~x790 & n42115 ;
  assign n42117 = ~n15141 & n42064 ;
  assign n42118 = ~x644 & n42117 ;
  assign n42119 = x715 & ~n42037 ;
  assign n42120 = ~n42118 & n42119 ;
  assign n42121 = ~n17389 & n42042 ;
  assign n42122 = n42037 | n42121 ;
  assign n42123 = ( x644 & x715 ) | ( x644 & n42122 ) | ( x715 & n42122 ) ;
  assign n42124 = ( ~x644 & x715 ) | ( ~x644 & n42115 ) | ( x715 & n42115 ) ;
  assign n42125 = n42123 | n42124 ;
  assign n42126 = ~n42120 & n42125 ;
  assign n42127 = x1160 | n42126 ;
  assign n42128 = x644 & n42117 ;
  assign n42129 = n42037 | n42128 ;
  assign n42130 = ~x715 & n42129 ;
  assign n42131 = x1160 & ~n42130 ;
  assign n42132 = n42123 & n42124 ;
  assign n42133 = n42131 & ~n42132 ;
  assign n42134 = x790 & ~n42133 ;
  assign n42135 = n42127 & n42134 ;
  assign n42136 = n42116 | n42135 ;
  assign n42137 = x230 & n42136 ;
  assign n42138 = ~x230 & n42036 ;
  assign n42139 = n42137 | n42138 ;
  assign n42140 = x568 & ~n31751 ;
  assign n42141 = x245 & n31751 ;
  assign n42142 = n42140 | n42141 ;
  assign n42143 = x569 & ~n31751 ;
  assign n42144 = ~x239 & n31751 ;
  assign n42145 = n42143 | n42144 ;
  assign n42146 = n31751 & n41858 ;
  assign n42147 = x570 & ~n42146 ;
  assign n42148 = x570 | n31750 ;
  assign n42149 = n41882 & ~n42148 ;
  assign n42150 = n42147 | n42149 ;
  assign n42151 = x571 & ~n32987 ;
  assign n42152 = x241 & n32987 ;
  assign n42153 = n42151 | n42152 ;
  assign n42154 = x572 & ~n32987 ;
  assign n42155 = x244 & n32987 ;
  assign n42156 = n42154 | n42155 ;
  assign n42157 = x573 & ~n32987 ;
  assign n42158 = x242 & n32987 ;
  assign n42159 = n42157 | n42158 ;
  assign n42160 = x574 & ~n31744 ;
  assign n42161 = x241 & n31744 ;
  assign n42162 = n42160 | n42161 ;
  assign n42163 = x575 & ~n32987 ;
  assign n42164 = x235 & n32987 ;
  assign n42165 = n42163 | n42164 ;
  assign n42166 = x576 & ~n32987 ;
  assign n42167 = x248 & n32987 ;
  assign n42168 = n42166 | n42167 ;
  assign n42169 = x577 & ~n32963 ;
  assign n42170 = x238 & n32963 ;
  assign n42171 = n42169 | n42170 ;
  assign n42172 = x578 & ~n31744 ;
  assign n42173 = x249 & n31744 ;
  assign n42174 = n42172 | n42173 ;
  assign n42175 = x579 & ~n31572 ;
  assign n42176 = x249 & n31572 ;
  assign n42177 = n42175 | n42176 ;
  assign n42178 = x580 & ~n32963 ;
  assign n42179 = x245 & n32963 ;
  assign n42180 = n42178 | n42179 ;
  assign n42181 = x581 & ~n31744 ;
  assign n42182 = x235 & n31744 ;
  assign n42183 = n42181 | n42182 ;
  assign n42184 = x582 & ~n31744 ;
  assign n42185 = x240 & n31744 ;
  assign n42186 = n42184 | n42185 ;
  assign n42187 = x584 & ~n31744 ;
  assign n42188 = x245 & n31744 ;
  assign n42189 = n42187 | n42188 ;
  assign n42190 = x585 & ~n31744 ;
  assign n42191 = x244 & n31744 ;
  assign n42192 = n42190 | n42191 ;
  assign n42193 = x586 & ~n31744 ;
  assign n42194 = x242 & n31744 ;
  assign n42195 = n42193 | n42194 ;
  assign n42196 = ~x230 & x587 ;
  assign n42197 = x230 & n14839 ;
  assign n42198 = ~n18257 & n42197 ;
  assign n42199 = ~n32528 & n42198 ;
  assign n42200 = ~n18255 & n42199 ;
  assign n42201 = ~n28134 & n42200 ;
  assign n42202 = n42196 | n42201 ;
  assign n42203 = ~x123 & n10310 ;
  assign n42204 = ( x588 & n41121 ) | ( x588 & n42203 ) | ( n41121 & n42203 ) ;
  assign n42205 = ( x591 & n41121 ) | ( x591 & ~n42203 ) | ( n41121 & ~n42203 ) ;
  assign n42206 = n42204 & n42205 ;
  assign n42207 = ~x201 & n41857 ;
  assign n42208 = ~x204 & n41833 ;
  assign n42209 = x233 & ~n42208 ;
  assign n42210 = ~n42207 & n42209 ;
  assign n42211 = ~x202 & n41857 ;
  assign n42212 = ~x205 & n41833 ;
  assign n42213 = x233 | n42212 ;
  assign n42214 = n42211 | n42213 ;
  assign n42215 = ~n42210 & n42214 ;
  assign n42216 = x237 & ~n42215 ;
  assign n42217 = ~x220 & n41857 ;
  assign n42218 = ~x206 & n41833 ;
  assign n42219 = x233 & ~n42218 ;
  assign n42220 = ~n42217 & n42219 ;
  assign n42221 = ~x203 & n41857 ;
  assign n42222 = ~x218 & n41833 ;
  assign n42223 = x233 | n42222 ;
  assign n42224 = n42221 | n42223 ;
  assign n42225 = ~n42220 & n42224 ;
  assign n42226 = x237 | n42225 ;
  assign n42227 = ~n42216 & n42226 ;
  assign n42228 = ( x588 & ~n41121 ) | ( x588 & n42203 ) | ( ~n41121 & n42203 ) ;
  assign n42229 = ( ~x590 & n41121 ) | ( ~x590 & n42203 ) | ( n41121 & n42203 ) ;
  assign n42230 = ~n42228 & n42229 ;
  assign n42231 = ( x591 & n41121 ) | ( x591 & n42203 ) | ( n41121 & n42203 ) ;
  assign n42232 = ( x592 & n41121 ) | ( x592 & ~n42203 ) | ( n41121 & ~n42203 ) ;
  assign n42233 = n42231 & n42232 ;
  assign n42234 = ( x592 & n41121 ) | ( x592 & n42203 ) | ( n41121 & n42203 ) ;
  assign n42235 = ( x590 & n41121 ) | ( x590 & ~n42203 ) | ( n41121 & ~n42203 ) ;
  assign n42236 = n42234 & n42235 ;
  assign n42237 = x247 | x561 ;
  assign n42238 = x245 | x503 ;
  assign n42239 = x244 | x541 ;
  assign n42240 = x240 | x542 ;
  assign n42241 = x241 | x500 ;
  assign n42242 = x241 & x500 ;
  assign n42243 = n42241 & ~n42242 ;
  assign n42244 = x234 & n41833 ;
  assign n42245 = x246 & x499 ;
  assign n42246 = ~x249 & x496 ;
  assign n42247 = ( ~x248 & x501 ) | ( ~x248 & n42246 ) | ( x501 & n42246 ) ;
  assign n42248 = x249 & ~x496 ;
  assign n42249 = ( x248 & ~x501 ) | ( x248 & n42248 ) | ( ~x501 & n42248 ) ;
  assign n42250 = n42247 | n42249 ;
  assign n42251 = ( x499 & ~n42245 ) | ( x499 & n42250 ) | ( ~n42245 & n42250 ) ;
  assign n42252 = ( x246 & ~n42245 ) | ( x246 & n42251 ) | ( ~n42245 & n42251 ) ;
  assign n42253 = ( x505 & ~n42244 ) | ( x505 & n42252 ) | ( ~n42244 & n42252 ) ;
  assign n42254 = ( x505 & n41834 ) | ( x505 & ~n42252 ) | ( n41834 & ~n42252 ) ;
  assign n42255 = ~n42253 & n42254 ;
  assign n42256 = ~n42243 & n42255 ;
  assign n42257 = ( x542 & ~n42240 ) | ( x542 & n42256 ) | ( ~n42240 & n42256 ) ;
  assign n42258 = ( x240 & ~n42240 ) | ( x240 & n42257 ) | ( ~n42240 & n42257 ) ;
  assign n42259 = x497 & n42258 ;
  assign n42260 = x239 | n42259 ;
  assign n42261 = ~x497 & n42258 ;
  assign n42262 = x239 & ~n42261 ;
  assign n42263 = n42260 & ~n42262 ;
  assign n42264 = x539 & n42263 ;
  assign n42265 = x242 & ~n42264 ;
  assign n42266 = ~x539 & n42263 ;
  assign n42267 = x242 | n42266 ;
  assign n42268 = ~n42265 & n42267 ;
  assign n42269 = x540 & n42268 ;
  assign n42270 = x235 & ~n42269 ;
  assign n42271 = ~x540 & n42268 ;
  assign n42272 = x235 | n42271 ;
  assign n42273 = ~n42270 & n42272 ;
  assign n42274 = ( x541 & ~n42239 ) | ( x541 & n42273 ) | ( ~n42239 & n42273 ) ;
  assign n42275 = ( x244 & ~n42239 ) | ( x244 & n42274 ) | ( ~n42239 & n42274 ) ;
  assign n42276 = ( x503 & ~n42238 ) | ( x503 & n42275 ) | ( ~n42238 & n42275 ) ;
  assign n42277 = ( x245 & ~n42238 ) | ( x245 & n42276 ) | ( ~n42238 & n42276 ) ;
  assign n42278 = ~x502 & n42277 ;
  assign n42279 = x247 | n42278 ;
  assign n42280 = n42237 & n42279 ;
  assign n42281 = x235 | x581 ;
  assign n42282 = x242 | x586 ;
  assign n42283 = x239 & ~x519 ;
  assign n42284 = x234 & n41857 ;
  assign n42285 = ~x249 & x578 ;
  assign n42286 = ( ~x248 & x521 ) | ( ~x248 & n42285 ) | ( x521 & n42285 ) ;
  assign n42287 = x249 & ~x578 ;
  assign n42288 = ( x248 & ~x521 ) | ( x248 & n42287 ) | ( ~x521 & n42287 ) ;
  assign n42289 = n42286 | n42288 ;
  assign n42290 = ~x246 & x520 ;
  assign n42291 = ( ~x241 & x574 ) | ( ~x241 & n42290 ) | ( x574 & n42290 ) ;
  assign n42292 = x246 & ~x520 ;
  assign n42293 = ( x241 & ~x574 ) | ( x241 & n42292 ) | ( ~x574 & n42292 ) ;
  assign n42294 = n42291 | n42293 ;
  assign n42295 = n42289 | n42294 ;
  assign n42296 = ( x518 & ~n42284 ) | ( x518 & n42295 ) | ( ~n42284 & n42295 ) ;
  assign n42297 = ( x518 & n41858 ) | ( x518 & ~n42295 ) | ( n41858 & ~n42295 ) ;
  assign n42298 = ~n42296 & n42297 ;
  assign n42299 = x582 & n42298 ;
  assign n42300 = x240 & ~n42299 ;
  assign n42301 = ~x582 & n42298 ;
  assign n42302 = x240 | n42301 ;
  assign n42303 = ~n42300 & n42302 ;
  assign n42304 = ( x519 & n42283 ) | ( x519 & n42303 ) | ( n42283 & n42303 ) ;
  assign n42305 = ( ~x239 & n42283 ) | ( ~x239 & n42304 ) | ( n42283 & n42304 ) ;
  assign n42306 = ( x586 & ~n42282 ) | ( x586 & n42305 ) | ( ~n42282 & n42305 ) ;
  assign n42307 = ( x242 & ~n42282 ) | ( x242 & n42306 ) | ( ~n42282 & n42306 ) ;
  assign n42308 = ( x581 & ~n42281 ) | ( x581 & n42307 ) | ( ~n42281 & n42307 ) ;
  assign n42309 = ( x235 & ~n42281 ) | ( x235 & n42308 ) | ( ~n42281 & n42308 ) ;
  assign n42310 = x585 & n42309 ;
  assign n42311 = x244 & ~n42310 ;
  assign n42312 = ~x585 & n42309 ;
  assign n42313 = x244 | n42312 ;
  assign n42314 = ~n42311 & n42313 ;
  assign n42315 = x584 & n42314 ;
  assign n42316 = x245 & ~n42315 ;
  assign n42317 = ~x584 & n42314 ;
  assign n42318 = x245 | n42317 ;
  assign n42319 = ~n42316 & n42318 ;
  assign n42320 = ( x502 & x561 ) | ( x502 & ~n42319 ) | ( x561 & ~n42319 ) ;
  assign n42321 = ( x245 & x584 ) | ( x245 & n42275 ) | ( x584 & n42275 ) ;
  assign n42322 = ( x244 & x585 ) | ( x244 & n42273 ) | ( x585 & n42273 ) ;
  assign n42323 = ( x235 & x540 ) | ( x235 & n42307 ) | ( x540 & n42307 ) ;
  assign n42324 = ( x242 & x539 ) | ( x242 & n42305 ) | ( x539 & n42305 ) ;
  assign n42325 = ( ~x239 & x497 ) | ( ~x239 & n42303 ) | ( x497 & n42303 ) ;
  assign n42326 = ( x240 & x582 ) | ( x240 & n42256 ) | ( x582 & n42256 ) ;
  assign n42327 = ( x241 & ~x500 ) | ( x241 & n42255 ) | ( ~x500 & n42255 ) ;
  assign n42328 = x241 & ~x500 ;
  assign n42329 = ( n42298 & n42327 ) | ( n42298 & ~n42328 ) | ( n42327 & ~n42328 ) ;
  assign n42330 = ( x240 & ~x582 ) | ( x240 & n42329 ) | ( ~x582 & n42329 ) ;
  assign n42331 = n42326 | n42330 ;
  assign n42332 = ~n42300 & n42331 ;
  assign n42333 = x542 | n42332 ;
  assign n42334 = ( ~x240 & x582 ) | ( ~x240 & n42329 ) | ( x582 & n42329 ) ;
  assign n42335 = ( x240 & x582 ) | ( x240 & ~n42256 ) | ( x582 & ~n42256 ) ;
  assign n42336 = ~n42334 & n42335 ;
  assign n42337 = n42302 & ~n42336 ;
  assign n42338 = x542 & ~n42337 ;
  assign n42339 = n42333 & ~n42338 ;
  assign n42340 = ( x239 & x497 ) | ( x239 & ~n42339 ) | ( x497 & ~n42339 ) ;
  assign n42341 = ~n42325 & n42340 ;
  assign n42342 = n42260 & ~n42341 ;
  assign n42343 = x519 | n42342 ;
  assign n42344 = ( x239 & x497 ) | ( x239 & n42339 ) | ( x497 & n42339 ) ;
  assign n42345 = ( x239 & ~x497 ) | ( x239 & n42303 ) | ( ~x497 & n42303 ) ;
  assign n42346 = n42344 | n42345 ;
  assign n42347 = ~n42262 & n42346 ;
  assign n42348 = x519 & ~n42347 ;
  assign n42349 = n42343 & ~n42348 ;
  assign n42350 = ( x242 & ~x539 ) | ( x242 & n42349 ) | ( ~x539 & n42349 ) ;
  assign n42351 = n42324 | n42350 ;
  assign n42352 = ~n42265 & n42351 ;
  assign n42353 = x586 | n42352 ;
  assign n42354 = ( ~x242 & x539 ) | ( ~x242 & n42349 ) | ( x539 & n42349 ) ;
  assign n42355 = ( x242 & x539 ) | ( x242 & ~n42305 ) | ( x539 & ~n42305 ) ;
  assign n42356 = ~n42354 & n42355 ;
  assign n42357 = n42267 & ~n42356 ;
  assign n42358 = x586 & ~n42357 ;
  assign n42359 = n42353 & ~n42358 ;
  assign n42360 = ( x235 & ~x540 ) | ( x235 & n42359 ) | ( ~x540 & n42359 ) ;
  assign n42361 = n42323 | n42360 ;
  assign n42362 = ~n42270 & n42361 ;
  assign n42363 = x581 | n42362 ;
  assign n42364 = ( ~x235 & x540 ) | ( ~x235 & n42359 ) | ( x540 & n42359 ) ;
  assign n42365 = ( x235 & x540 ) | ( x235 & ~n42307 ) | ( x540 & ~n42307 ) ;
  assign n42366 = ~n42364 & n42365 ;
  assign n42367 = n42272 & ~n42366 ;
  assign n42368 = x581 & ~n42367 ;
  assign n42369 = n42363 & ~n42368 ;
  assign n42370 = ( x244 & ~x585 ) | ( x244 & n42369 ) | ( ~x585 & n42369 ) ;
  assign n42371 = n42322 | n42370 ;
  assign n42372 = ~n42311 & n42371 ;
  assign n42373 = x541 | n42372 ;
  assign n42374 = ( ~x244 & x585 ) | ( ~x244 & n42369 ) | ( x585 & n42369 ) ;
  assign n42375 = ( x244 & x585 ) | ( x244 & ~n42273 ) | ( x585 & ~n42273 ) ;
  assign n42376 = ~n42374 & n42375 ;
  assign n42377 = n42313 & ~n42376 ;
  assign n42378 = x541 & ~n42377 ;
  assign n42379 = n42373 & ~n42378 ;
  assign n42380 = ( x245 & ~x584 ) | ( x245 & n42379 ) | ( ~x584 & n42379 ) ;
  assign n42381 = n42321 | n42380 ;
  assign n42382 = ~n42316 & n42381 ;
  assign n42383 = x503 | n42382 ;
  assign n42384 = ( ~x245 & x584 ) | ( ~x245 & n42379 ) | ( x584 & n42379 ) ;
  assign n42385 = ( x245 & x584 ) | ( x245 & ~n42275 ) | ( x584 & ~n42275 ) ;
  assign n42386 = ~n42384 & n42385 ;
  assign n42387 = n42318 & ~n42386 ;
  assign n42388 = x503 & ~n42387 ;
  assign n42389 = n42383 & ~n42388 ;
  assign n42390 = ( x502 & ~x561 ) | ( x502 & n42389 ) | ( ~x561 & n42389 ) ;
  assign n42391 = ~n42320 & n42390 ;
  assign n42392 = n42280 | n42391 ;
  assign n42393 = x247 & x561 ;
  assign n42394 = x502 & n42277 ;
  assign n42395 = x247 & ~n42394 ;
  assign n42396 = n42393 | n42395 ;
  assign n42397 = ( x502 & x561 ) | ( x502 & n42319 ) | ( x561 & n42319 ) ;
  assign n42398 = ( ~x502 & x561 ) | ( ~x502 & n42389 ) | ( x561 & n42389 ) ;
  assign n42399 = n42397 & n42398 ;
  assign n42400 = n42396 & ~n42399 ;
  assign n42401 = n42392 & ~n42400 ;
  assign n42402 = ~x238 & n42401 ;
  assign n42403 = x522 | n42402 ;
  assign n42404 = n42279 & ~n42395 ;
  assign n42405 = ( x238 & x522 ) | ( x238 & ~n42404 ) | ( x522 & ~n42404 ) ;
  assign n42406 = n42237 & ~n42393 ;
  assign n42407 = n42319 & ~n42406 ;
  assign n42408 = ( x238 & ~x522 ) | ( x238 & n42407 ) | ( ~x522 & n42407 ) ;
  assign n42409 = n42405 & ~n42408 ;
  assign n42410 = x543 | n42409 ;
  assign n42411 = n42403 & ~n42410 ;
  assign n42412 = x238 & n42401 ;
  assign n42413 = x522 & ~n42412 ;
  assign n42414 = ( x238 & x522 ) | ( x238 & n42404 ) | ( x522 & n42404 ) ;
  assign n42415 = ( ~x238 & x522 ) | ( ~x238 & n42407 ) | ( x522 & n42407 ) ;
  assign n42416 = n42414 | n42415 ;
  assign n42417 = x543 & n42416 ;
  assign n42418 = ~n42413 & n42417 ;
  assign n42419 = n42411 | n42418 ;
  assign n42420 = ( x233 & x237 ) | ( x233 & ~n42419 ) | ( x237 & ~n42419 ) ;
  assign n42421 = x240 | x535 ;
  assign n42422 = x241 | x506 ;
  assign n42423 = x557 & ~n42244 ;
  assign n42424 = ( x246 & ~x536 ) | ( x246 & n42423 ) | ( ~x536 & n42423 ) ;
  assign n42425 = x557 | n41834 ;
  assign n42426 = ( x246 & ~x536 ) | ( x246 & n42425 ) | ( ~x536 & n42425 ) ;
  assign n42427 = ~n42424 & n42426 ;
  assign n42428 = ~x538 & n42427 ;
  assign n42429 = x249 | n42428 ;
  assign n42430 = x538 & n42427 ;
  assign n42431 = x249 & ~n42430 ;
  assign n42432 = n42429 & ~n42431 ;
  assign n42433 = ~x537 & n42432 ;
  assign n42434 = x248 | n42433 ;
  assign n42435 = x537 & n42432 ;
  assign n42436 = x248 & ~n42435 ;
  assign n42437 = n42434 & ~n42436 ;
  assign n42438 = ( x506 & ~n42422 ) | ( x506 & n42437 ) | ( ~n42422 & n42437 ) ;
  assign n42439 = ( x241 & ~n42422 ) | ( x241 & n42438 ) | ( ~n42422 & n42438 ) ;
  assign n42440 = ( x535 & ~n42421 ) | ( x535 & n42439 ) | ( ~n42421 & n42439 ) ;
  assign n42441 = ( x240 & ~n42421 ) | ( x240 & n42440 ) | ( ~n42421 & n42440 ) ;
  assign n42442 = x534 & n42441 ;
  assign n42443 = x239 | n42442 ;
  assign n42444 = ~x534 & n42441 ;
  assign n42445 = x239 & ~n42444 ;
  assign n42446 = n42443 & ~n42445 ;
  assign n42447 = x504 & n42446 ;
  assign n42448 = x242 & ~n42447 ;
  assign n42449 = ~x504 & n42446 ;
  assign n42450 = x242 | n42449 ;
  assign n42451 = ~n42448 & n42450 ;
  assign n42452 = x533 & n42451 ;
  assign n42453 = x235 & ~n42452 ;
  assign n42454 = ~x533 & n42451 ;
  assign n42455 = x235 | n42454 ;
  assign n42456 = ~n42453 & n42455 ;
  assign n42457 = x558 & n42456 ;
  assign n42458 = x244 & ~n42457 ;
  assign n42459 = ~x558 & n42456 ;
  assign n42460 = x244 | n42459 ;
  assign n42461 = ~n42458 & n42460 ;
  assign n42462 = x509 & n42461 ;
  assign n42463 = x245 & ~n42462 ;
  assign n42464 = ~x509 & n42461 ;
  assign n42465 = x245 | n42464 ;
  assign n42466 = ~n42463 & n42465 ;
  assign n42467 = x508 & n42466 ;
  assign n42468 = x247 & ~n42467 ;
  assign n42469 = x245 | x514 ;
  assign n42470 = x244 | x513 ;
  assign n42471 = x235 | x512 ;
  assign n42472 = x242 | x510 ;
  assign n42473 = x239 & ~x488 ;
  assign n42474 = x248 | x481 ;
  assign n42475 = x249 | x579 ;
  assign n42476 = x511 & ~n42284 ;
  assign n42477 = ( x246 & ~x487 ) | ( x246 & n42476 ) | ( ~x487 & n42476 ) ;
  assign n42478 = x511 | n41858 ;
  assign n42479 = ( x246 & ~x487 ) | ( x246 & n42478 ) | ( ~x487 & n42478 ) ;
  assign n42480 = ~n42477 & n42479 ;
  assign n42481 = ( x579 & ~n42475 ) | ( x579 & n42480 ) | ( ~n42475 & n42480 ) ;
  assign n42482 = ( x249 & ~n42475 ) | ( x249 & n42481 ) | ( ~n42475 & n42481 ) ;
  assign n42483 = ( x481 & ~n42474 ) | ( x481 & n42482 ) | ( ~n42474 & n42482 ) ;
  assign n42484 = ( x248 & ~n42474 ) | ( x248 & n42483 ) | ( ~n42474 & n42483 ) ;
  assign n42485 = x559 & n42484 ;
  assign n42486 = x241 & ~n42485 ;
  assign n42487 = ~x559 & n42484 ;
  assign n42488 = x241 | n42487 ;
  assign n42489 = ~n42486 & n42488 ;
  assign n42490 = x515 & n42489 ;
  assign n42491 = x240 & ~n42490 ;
  assign n42492 = ~x515 & n42489 ;
  assign n42493 = x240 | n42492 ;
  assign n42494 = ~n42491 & n42493 ;
  assign n42495 = ( x488 & n42473 ) | ( x488 & n42494 ) | ( n42473 & n42494 ) ;
  assign n42496 = ( ~x239 & n42473 ) | ( ~x239 & n42495 ) | ( n42473 & n42495 ) ;
  assign n42497 = ( x510 & ~n42472 ) | ( x510 & n42496 ) | ( ~n42472 & n42496 ) ;
  assign n42498 = ( x242 & ~n42472 ) | ( x242 & n42497 ) | ( ~n42472 & n42497 ) ;
  assign n42499 = ( x512 & ~n42471 ) | ( x512 & n42498 ) | ( ~n42471 & n42498 ) ;
  assign n42500 = ( x235 & ~n42471 ) | ( x235 & n42499 ) | ( ~n42471 & n42499 ) ;
  assign n42501 = ( x513 & ~n42470 ) | ( x513 & n42500 ) | ( ~n42470 & n42500 ) ;
  assign n42502 = ( x244 & ~n42470 ) | ( x244 & n42501 ) | ( ~n42470 & n42501 ) ;
  assign n42503 = ( x514 & ~n42469 ) | ( x514 & n42502 ) | ( ~n42469 & n42502 ) ;
  assign n42504 = ( x245 & ~n42469 ) | ( x245 & n42503 ) | ( ~n42469 & n42503 ) ;
  assign n42505 = ( x247 & x508 ) | ( x247 & n42504 ) | ( x508 & n42504 ) ;
  assign n42506 = ( x245 & x509 ) | ( x245 & n42502 ) | ( x509 & n42502 ) ;
  assign n42507 = ( x244 & x558 ) | ( x244 & n42500 ) | ( x558 & n42500 ) ;
  assign n42508 = ( x235 & x533 ) | ( x235 & n42498 ) | ( x533 & n42498 ) ;
  assign n42509 = ( x242 & x504 ) | ( x242 & n42496 ) | ( x504 & n42496 ) ;
  assign n42510 = ( ~x239 & x534 ) | ( ~x239 & n42494 ) | ( x534 & n42494 ) ;
  assign n42511 = ( x240 & x515 ) | ( x240 & n42439 ) | ( x515 & n42439 ) ;
  assign n42512 = ( x241 & x559 ) | ( x241 & n42437 ) | ( x559 & n42437 ) ;
  assign n42513 = ( x248 & x537 ) | ( x248 & n42482 ) | ( x537 & n42482 ) ;
  assign n42514 = n42429 & n42480 ;
  assign n42515 = ( x579 & n42432 ) | ( x579 & n42514 ) | ( n42432 & n42514 ) ;
  assign n42516 = ( ~x579 & n42432 ) | ( ~x579 & n42482 ) | ( n42432 & n42482 ) ;
  assign n42517 = n42515 | n42516 ;
  assign n42518 = ( x248 & ~x537 ) | ( x248 & n42517 ) | ( ~x537 & n42517 ) ;
  assign n42519 = n42513 | n42518 ;
  assign n42520 = ~n42436 & n42519 ;
  assign n42521 = x481 | n42520 ;
  assign n42522 = ( ~x248 & x537 ) | ( ~x248 & n42517 ) | ( x537 & n42517 ) ;
  assign n42523 = ( x248 & x537 ) | ( x248 & ~n42482 ) | ( x537 & ~n42482 ) ;
  assign n42524 = ~n42522 & n42523 ;
  assign n42525 = n42434 & ~n42524 ;
  assign n42526 = x481 & ~n42525 ;
  assign n42527 = n42521 & ~n42526 ;
  assign n42528 = ( x241 & ~x559 ) | ( x241 & n42527 ) | ( ~x559 & n42527 ) ;
  assign n42529 = n42512 | n42528 ;
  assign n42530 = ~n42486 & n42529 ;
  assign n42531 = x506 | n42530 ;
  assign n42532 = ( ~x241 & x559 ) | ( ~x241 & n42527 ) | ( x559 & n42527 ) ;
  assign n42533 = ( x241 & x559 ) | ( x241 & ~n42437 ) | ( x559 & ~n42437 ) ;
  assign n42534 = ~n42532 & n42533 ;
  assign n42535 = n42488 & ~n42534 ;
  assign n42536 = x506 & ~n42535 ;
  assign n42537 = n42531 & ~n42536 ;
  assign n42538 = ( x240 & ~x515 ) | ( x240 & n42537 ) | ( ~x515 & n42537 ) ;
  assign n42539 = n42511 | n42538 ;
  assign n42540 = ~n42491 & n42539 ;
  assign n42541 = x535 | n42540 ;
  assign n42542 = ( ~x240 & x515 ) | ( ~x240 & n42537 ) | ( x515 & n42537 ) ;
  assign n42543 = ( x240 & x515 ) | ( x240 & ~n42439 ) | ( x515 & ~n42439 ) ;
  assign n42544 = ~n42542 & n42543 ;
  assign n42545 = n42493 & ~n42544 ;
  assign n42546 = x535 & ~n42545 ;
  assign n42547 = n42541 & ~n42546 ;
  assign n42548 = ( x239 & x534 ) | ( x239 & ~n42547 ) | ( x534 & ~n42547 ) ;
  assign n42549 = ~n42510 & n42548 ;
  assign n42550 = n42443 & ~n42549 ;
  assign n42551 = x488 | n42550 ;
  assign n42552 = ( x239 & x534 ) | ( x239 & n42547 ) | ( x534 & n42547 ) ;
  assign n42553 = ( x239 & ~x534 ) | ( x239 & n42494 ) | ( ~x534 & n42494 ) ;
  assign n42554 = n42552 | n42553 ;
  assign n42555 = ~n42445 & n42554 ;
  assign n42556 = x488 & ~n42555 ;
  assign n42557 = n42551 & ~n42556 ;
  assign n42558 = ( x242 & ~x504 ) | ( x242 & n42557 ) | ( ~x504 & n42557 ) ;
  assign n42559 = n42509 | n42558 ;
  assign n42560 = ~n42448 & n42559 ;
  assign n42561 = x510 | n42560 ;
  assign n42562 = ( ~x242 & x504 ) | ( ~x242 & n42557 ) | ( x504 & n42557 ) ;
  assign n42563 = ( x242 & x504 ) | ( x242 & ~n42496 ) | ( x504 & ~n42496 ) ;
  assign n42564 = ~n42562 & n42563 ;
  assign n42565 = n42450 & ~n42564 ;
  assign n42566 = x510 & ~n42565 ;
  assign n42567 = n42561 & ~n42566 ;
  assign n42568 = ( x235 & ~x533 ) | ( x235 & n42567 ) | ( ~x533 & n42567 ) ;
  assign n42569 = n42508 | n42568 ;
  assign n42570 = ~n42453 & n42569 ;
  assign n42571 = x512 | n42570 ;
  assign n42572 = ( ~x235 & x533 ) | ( ~x235 & n42567 ) | ( x533 & n42567 ) ;
  assign n42573 = ( x235 & x533 ) | ( x235 & ~n42498 ) | ( x533 & ~n42498 ) ;
  assign n42574 = ~n42572 & n42573 ;
  assign n42575 = n42455 & ~n42574 ;
  assign n42576 = x512 & ~n42575 ;
  assign n42577 = n42571 & ~n42576 ;
  assign n42578 = ( x244 & ~x558 ) | ( x244 & n42577 ) | ( ~x558 & n42577 ) ;
  assign n42579 = n42507 | n42578 ;
  assign n42580 = ~n42458 & n42579 ;
  assign n42581 = x513 | n42580 ;
  assign n42582 = ( ~x244 & x558 ) | ( ~x244 & n42577 ) | ( x558 & n42577 ) ;
  assign n42583 = ( x244 & x558 ) | ( x244 & ~n42500 ) | ( x558 & ~n42500 ) ;
  assign n42584 = ~n42582 & n42583 ;
  assign n42585 = n42460 & ~n42584 ;
  assign n42586 = x513 & ~n42585 ;
  assign n42587 = n42581 & ~n42586 ;
  assign n42588 = ( x245 & ~x509 ) | ( x245 & n42587 ) | ( ~x509 & n42587 ) ;
  assign n42589 = n42506 | n42588 ;
  assign n42590 = ~n42463 & n42589 ;
  assign n42591 = x514 | n42590 ;
  assign n42592 = ( ~x245 & x509 ) | ( ~x245 & n42587 ) | ( x509 & n42587 ) ;
  assign n42593 = ( x245 & x509 ) | ( x245 & ~n42502 ) | ( x509 & ~n42502 ) ;
  assign n42594 = ~n42592 & n42593 ;
  assign n42595 = n42465 & ~n42594 ;
  assign n42596 = x514 & ~n42595 ;
  assign n42597 = n42591 & ~n42596 ;
  assign n42598 = ( x247 & ~x508 ) | ( x247 & n42597 ) | ( ~x508 & n42597 ) ;
  assign n42599 = n42505 | n42598 ;
  assign n42600 = ~n42468 & n42599 ;
  assign n42601 = x516 | n42600 ;
  assign n42602 = ~x508 & n42466 ;
  assign n42603 = x247 | n42602 ;
  assign n42604 = ( ~x247 & x508 ) | ( ~x247 & n42597 ) | ( x508 & n42597 ) ;
  assign n42605 = ( x247 & x508 ) | ( x247 & ~n42504 ) | ( x508 & ~n42504 ) ;
  assign n42606 = ~n42604 & n42605 ;
  assign n42607 = n42603 & ~n42606 ;
  assign n42608 = x516 & ~n42607 ;
  assign n42609 = n42601 & ~n42608 ;
  assign n42610 = ~x238 & n42609 ;
  assign n42611 = x517 | n42610 ;
  assign n42612 = ~n42468 & n42603 ;
  assign n42613 = ( x238 & x517 ) | ( x238 & ~n42612 ) | ( x517 & ~n42612 ) ;
  assign n42614 = x247 | x516 ;
  assign n42615 = ( x516 & n42504 ) | ( x516 & ~n42614 ) | ( n42504 & ~n42614 ) ;
  assign n42616 = ( x247 & ~n42614 ) | ( x247 & n42615 ) | ( ~n42614 & n42615 ) ;
  assign n42617 = ( x238 & ~x517 ) | ( x238 & n42616 ) | ( ~x517 & n42616 ) ;
  assign n42618 = n42613 & ~n42617 ;
  assign n42619 = x507 | n42618 ;
  assign n42620 = n42611 & ~n42619 ;
  assign n42621 = x238 & n42609 ;
  assign n42622 = x517 & ~n42621 ;
  assign n42623 = ( x238 & x517 ) | ( x238 & n42612 ) | ( x517 & n42612 ) ;
  assign n42624 = ( ~x238 & x517 ) | ( ~x238 & n42616 ) | ( x517 & n42616 ) ;
  assign n42625 = n42623 | n42624 ;
  assign n42626 = x507 & n42625 ;
  assign n42627 = ~n42622 & n42626 ;
  assign n42628 = n42620 | n42627 ;
  assign n42629 = ( x233 & ~x237 ) | ( x233 & n42628 ) | ( ~x237 & n42628 ) ;
  assign n42630 = n42420 & ~n42629 ;
  assign n42631 = x244 | x493 ;
  assign n42632 = x240 | x492 ;
  assign n42633 = x240 & x492 ;
  assign n42634 = n42632 & ~n42633 ;
  assign n42635 = x241 | x490 ;
  assign n42636 = x544 & ~n42244 ;
  assign n42637 = x544 | n41834 ;
  assign n42638 = ( ~x246 & x546 ) | ( ~x246 & n42637 ) | ( x546 & n42637 ) ;
  assign n42639 = ~x249 & x484 ;
  assign n42640 = ( ~x248 & x548 ) | ( ~x248 & n42639 ) | ( x548 & n42639 ) ;
  assign n42641 = x249 & ~x484 ;
  assign n42642 = ( x248 & ~x548 ) | ( x248 & n42641 ) | ( ~x548 & n42641 ) ;
  assign n42643 = n42640 | n42642 ;
  assign n42644 = ( ~x246 & x546 ) | ( ~x246 & n42643 ) | ( x546 & n42643 ) ;
  assign n42645 = n42638 & ~n42644 ;
  assign n42646 = ~n42636 & n42645 ;
  assign n42647 = ( x490 & ~n42635 ) | ( x490 & n42646 ) | ( ~n42635 & n42646 ) ;
  assign n42648 = ( x241 & ~n42635 ) | ( x241 & n42647 ) | ( ~n42635 & n42647 ) ;
  assign n42649 = ~n42634 & n42648 ;
  assign n42650 = x494 & n42649 ;
  assign n42651 = x239 | n42650 ;
  assign n42652 = ~x494 & n42649 ;
  assign n42653 = x239 & ~n42652 ;
  assign n42654 = n42651 & ~n42653 ;
  assign n42655 = x483 & n42654 ;
  assign n42656 = x242 & ~n42655 ;
  assign n42657 = ~x483 & n42654 ;
  assign n42658 = x242 | n42657 ;
  assign n42659 = ~n42656 & n42658 ;
  assign n42660 = x495 & n42659 ;
  assign n42661 = x235 & ~n42660 ;
  assign n42662 = ~x495 & n42659 ;
  assign n42663 = x235 | n42662 ;
  assign n42664 = ~n42661 & n42663 ;
  assign n42665 = ( x493 & ~n42631 ) | ( x493 & n42664 ) | ( ~n42631 & n42664 ) ;
  assign n42666 = ( x244 & ~n42631 ) | ( x244 & n42665 ) | ( ~n42631 & n42665 ) ;
  assign n42667 = x545 & n42666 ;
  assign n42668 = x245 & ~n42667 ;
  assign n42669 = ~x545 & n42666 ;
  assign n42670 = x245 | n42669 ;
  assign n42671 = ~n42668 & n42670 ;
  assign n42672 = x547 & n42671 ;
  assign n42673 = x247 & ~n42672 ;
  assign n42674 = x245 | x525 ;
  assign n42675 = x235 | x575 ;
  assign n42676 = x242 | x573 ;
  assign n42677 = x239 & ~x524 ;
  assign n42678 = x246 & x526 ;
  assign n42679 = ~x249 & x528 ;
  assign n42680 = ( ~x248 & x576 ) | ( ~x248 & n42679 ) | ( x576 & n42679 ) ;
  assign n42681 = x249 & ~x528 ;
  assign n42682 = ( x248 & ~x576 ) | ( x248 & n42681 ) | ( ~x576 & n42681 ) ;
  assign n42683 = n42680 | n42682 ;
  assign n42684 = ( x526 & ~n42678 ) | ( x526 & n42683 ) | ( ~n42678 & n42683 ) ;
  assign n42685 = ( x246 & ~n42678 ) | ( x246 & n42684 ) | ( ~n42678 & n42684 ) ;
  assign n42686 = ( x523 & ~n42284 ) | ( x523 & n42685 ) | ( ~n42284 & n42685 ) ;
  assign n42687 = ( x523 & n41858 ) | ( x523 & ~n42685 ) | ( n41858 & ~n42685 ) ;
  assign n42688 = ~n42686 & n42687 ;
  assign n42689 = x571 & n42688 ;
  assign n42690 = x241 & ~n42689 ;
  assign n42691 = ~x571 & n42688 ;
  assign n42692 = x241 | n42691 ;
  assign n42693 = ~n42690 & n42692 ;
  assign n42694 = ~x530 & n42693 ;
  assign n42695 = x240 | n42694 ;
  assign n42696 = x530 & n42693 ;
  assign n42697 = x240 & ~n42696 ;
  assign n42698 = n42695 & ~n42697 ;
  assign n42699 = ( x524 & n42677 ) | ( x524 & n42698 ) | ( n42677 & n42698 ) ;
  assign n42700 = ( ~x239 & n42677 ) | ( ~x239 & n42699 ) | ( n42677 & n42699 ) ;
  assign n42701 = ( x573 & ~n42676 ) | ( x573 & n42700 ) | ( ~n42676 & n42700 ) ;
  assign n42702 = ( x242 & ~n42676 ) | ( x242 & n42701 ) | ( ~n42676 & n42701 ) ;
  assign n42703 = ( x575 & ~n42675 ) | ( x575 & n42702 ) | ( ~n42675 & n42702 ) ;
  assign n42704 = ( x235 & ~n42675 ) | ( x235 & n42703 ) | ( ~n42675 & n42703 ) ;
  assign n42705 = x572 & n42704 ;
  assign n42706 = x244 & ~n42705 ;
  assign n42707 = ~x572 & n42704 ;
  assign n42708 = x244 | n42707 ;
  assign n42709 = ~n42706 & n42708 ;
  assign n42710 = ( x525 & ~n42674 ) | ( x525 & n42709 ) | ( ~n42674 & n42709 ) ;
  assign n42711 = ( x245 & ~n42674 ) | ( x245 & n42710 ) | ( ~n42674 & n42710 ) ;
  assign n42712 = ( x247 & x547 ) | ( x247 & n42711 ) | ( x547 & n42711 ) ;
  assign n42713 = ( x245 & x545 ) | ( x245 & n42709 ) | ( x545 & n42709 ) ;
  assign n42714 = ( x244 & x572 ) | ( x244 & n42664 ) | ( x572 & n42664 ) ;
  assign n42715 = ( x235 & x495 ) | ( x235 & n42702 ) | ( x495 & n42702 ) ;
  assign n42716 = ( x242 & x483 ) | ( x242 & n42700 ) | ( x483 & n42700 ) ;
  assign n42717 = ( ~x239 & x494 ) | ( ~x239 & n42698 ) | ( x494 & n42698 ) ;
  assign n42718 = n42632 & n42695 ;
  assign n42719 = ( x492 & x530 ) | ( x492 & ~n42648 ) | ( x530 & ~n42648 ) ;
  assign n42720 = x241 | n42646 ;
  assign n42721 = n42691 | n42720 ;
  assign n42722 = ~n42690 & n42721 ;
  assign n42723 = x490 | n42722 ;
  assign n42724 = x241 & ~n42646 ;
  assign n42725 = ~n42689 & n42724 ;
  assign n42726 = n42692 & ~n42725 ;
  assign n42727 = x490 & ~n42726 ;
  assign n42728 = n42723 & ~n42727 ;
  assign n42729 = ( ~x492 & x530 ) | ( ~x492 & n42728 ) | ( x530 & n42728 ) ;
  assign n42730 = ~n42719 & n42729 ;
  assign n42731 = n42718 | n42730 ;
  assign n42732 = n42633 | n42697 ;
  assign n42733 = ( x492 & ~x530 ) | ( x492 & n42728 ) | ( ~x530 & n42728 ) ;
  assign n42734 = ( x492 & x530 ) | ( x492 & n42648 ) | ( x530 & n42648 ) ;
  assign n42735 = n42733 & n42734 ;
  assign n42736 = n42732 & ~n42735 ;
  assign n42737 = n42731 & ~n42736 ;
  assign n42738 = ( x239 & x494 ) | ( x239 & ~n42737 ) | ( x494 & ~n42737 ) ;
  assign n42739 = ~n42717 & n42738 ;
  assign n42740 = n42651 & ~n42739 ;
  assign n42741 = x524 | n42740 ;
  assign n42742 = ( x239 & x494 ) | ( x239 & n42737 ) | ( x494 & n42737 ) ;
  assign n42743 = ( x239 & ~x494 ) | ( x239 & n42698 ) | ( ~x494 & n42698 ) ;
  assign n42744 = n42742 | n42743 ;
  assign n42745 = ~n42653 & n42744 ;
  assign n42746 = x524 & ~n42745 ;
  assign n42747 = n42741 & ~n42746 ;
  assign n42748 = ( x242 & ~x483 ) | ( x242 & n42747 ) | ( ~x483 & n42747 ) ;
  assign n42749 = n42716 | n42748 ;
  assign n42750 = ~n42656 & n42749 ;
  assign n42751 = x573 | n42750 ;
  assign n42752 = ( ~x242 & x483 ) | ( ~x242 & n42747 ) | ( x483 & n42747 ) ;
  assign n42753 = ( x242 & x483 ) | ( x242 & ~n42700 ) | ( x483 & ~n42700 ) ;
  assign n42754 = ~n42752 & n42753 ;
  assign n42755 = n42658 & ~n42754 ;
  assign n42756 = x573 & ~n42755 ;
  assign n42757 = n42751 & ~n42756 ;
  assign n42758 = ( x235 & ~x495 ) | ( x235 & n42757 ) | ( ~x495 & n42757 ) ;
  assign n42759 = n42715 | n42758 ;
  assign n42760 = ~n42661 & n42759 ;
  assign n42761 = x575 | n42760 ;
  assign n42762 = ( ~x235 & x495 ) | ( ~x235 & n42757 ) | ( x495 & n42757 ) ;
  assign n42763 = ( x235 & x495 ) | ( x235 & ~n42702 ) | ( x495 & ~n42702 ) ;
  assign n42764 = ~n42762 & n42763 ;
  assign n42765 = n42663 & ~n42764 ;
  assign n42766 = x575 & ~n42765 ;
  assign n42767 = n42761 & ~n42766 ;
  assign n42768 = ( x244 & ~x572 ) | ( x244 & n42767 ) | ( ~x572 & n42767 ) ;
  assign n42769 = n42714 | n42768 ;
  assign n42770 = ~n42706 & n42769 ;
  assign n42771 = x493 | n42770 ;
  assign n42772 = ( ~x244 & x572 ) | ( ~x244 & n42767 ) | ( x572 & n42767 ) ;
  assign n42773 = ( x244 & x572 ) | ( x244 & ~n42664 ) | ( x572 & ~n42664 ) ;
  assign n42774 = ~n42772 & n42773 ;
  assign n42775 = n42708 & ~n42774 ;
  assign n42776 = x493 & ~n42775 ;
  assign n42777 = n42771 & ~n42776 ;
  assign n42778 = ( x245 & ~x545 ) | ( x245 & n42777 ) | ( ~x545 & n42777 ) ;
  assign n42779 = n42713 | n42778 ;
  assign n42780 = ~n42668 & n42779 ;
  assign n42781 = x525 | n42780 ;
  assign n42782 = ( ~x245 & x545 ) | ( ~x245 & n42777 ) | ( x545 & n42777 ) ;
  assign n42783 = ( x245 & x545 ) | ( x245 & ~n42709 ) | ( x545 & ~n42709 ) ;
  assign n42784 = ~n42782 & n42783 ;
  assign n42785 = n42670 & ~n42784 ;
  assign n42786 = x525 & ~n42785 ;
  assign n42787 = n42781 & ~n42786 ;
  assign n42788 = ( x247 & ~x547 ) | ( x247 & n42787 ) | ( ~x547 & n42787 ) ;
  assign n42789 = n42712 | n42788 ;
  assign n42790 = ~n42673 & n42789 ;
  assign n42791 = x527 | n42790 ;
  assign n42792 = ~x547 & n42671 ;
  assign n42793 = x247 | n42792 ;
  assign n42794 = ( ~x247 & x547 ) | ( ~x247 & n42787 ) | ( x547 & n42787 ) ;
  assign n42795 = ( x247 & x547 ) | ( x247 & ~n42711 ) | ( x547 & ~n42711 ) ;
  assign n42796 = ~n42794 & n42795 ;
  assign n42797 = n42793 & ~n42796 ;
  assign n42798 = x527 & ~n42797 ;
  assign n42799 = n42791 & ~n42798 ;
  assign n42800 = ~x238 & n42799 ;
  assign n42801 = x529 | n42800 ;
  assign n42802 = ~n42673 & n42793 ;
  assign n42803 = ( x238 & x529 ) | ( x238 & ~n42802 ) | ( x529 & ~n42802 ) ;
  assign n42804 = x247 | x527 ;
  assign n42805 = ( x527 & n42711 ) | ( x527 & ~n42804 ) | ( n42711 & ~n42804 ) ;
  assign n42806 = ( x247 & ~n42804 ) | ( x247 & n42805 ) | ( ~n42804 & n42805 ) ;
  assign n42807 = ( x238 & ~x529 ) | ( x238 & n42806 ) | ( ~x529 & n42806 ) ;
  assign n42808 = n42803 & ~n42807 ;
  assign n42809 = x491 | n42808 ;
  assign n42810 = n42801 & ~n42809 ;
  assign n42811 = x238 & n42799 ;
  assign n42812 = x529 & ~n42811 ;
  assign n42813 = ( x238 & x529 ) | ( x238 & n42802 ) | ( x529 & n42802 ) ;
  assign n42814 = ( ~x238 & x529 ) | ( ~x238 & n42806 ) | ( x529 & n42806 ) ;
  assign n42815 = n42813 | n42814 ;
  assign n42816 = x491 & n42815 ;
  assign n42817 = ~n42812 & n42816 ;
  assign n42818 = n42810 | n42817 ;
  assign n42819 = ( x233 & x237 ) | ( x233 & n42818 ) | ( x237 & n42818 ) ;
  assign n42820 = x245 | x580 ;
  assign n42821 = ~x248 & x554 ;
  assign n42822 = ( ~x246 & x563 ) | ( ~x246 & n42821 ) | ( x563 & n42821 ) ;
  assign n42823 = x248 & ~x554 ;
  assign n42824 = ( x246 & ~x563 ) | ( x246 & n42823 ) | ( ~x563 & n42823 ) ;
  assign n42825 = n42822 | n42824 ;
  assign n42826 = ( ~x240 & x551 ) | ( ~x240 & n42825 ) | ( x551 & n42825 ) ;
  assign n42827 = ~x249 & x555 ;
  assign n42828 = ( ~x241 & x553 ) | ( ~x241 & n42827 ) | ( x553 & n42827 ) ;
  assign n42829 = x249 & ~x555 ;
  assign n42830 = ( x241 & ~x553 ) | ( x241 & n42829 ) | ( ~x553 & n42829 ) ;
  assign n42831 = n42828 | n42830 ;
  assign n42832 = ( x240 & ~x551 ) | ( x240 & n42831 ) | ( ~x551 & n42831 ) ;
  assign n42833 = n42826 | n42832 ;
  assign n42834 = ( x485 & ~n42244 ) | ( x485 & n42833 ) | ( ~n42244 & n42833 ) ;
  assign n42835 = ( x485 & n41834 ) | ( x485 & ~n42833 ) | ( n41834 & ~n42833 ) ;
  assign n42836 = ~n42834 & n42835 ;
  assign n42837 = x550 & n42836 ;
  assign n42838 = x239 | n42837 ;
  assign n42839 = ~x550 & n42836 ;
  assign n42840 = x239 & ~n42839 ;
  assign n42841 = n42838 & ~n42840 ;
  assign n42842 = ~x489 & n42841 ;
  assign n42843 = x242 | n42842 ;
  assign n42844 = x489 & n42841 ;
  assign n42845 = x242 & ~n42844 ;
  assign n42846 = n42843 & ~n42845 ;
  assign n42847 = x549 & n42846 ;
  assign n42848 = x235 & ~n42847 ;
  assign n42849 = ~x549 & n42846 ;
  assign n42850 = x235 | n42849 ;
  assign n42851 = ~n42848 & n42850 ;
  assign n42852 = x486 & n42851 ;
  assign n42853 = x244 & ~n42852 ;
  assign n42854 = ~x486 & n42851 ;
  assign n42855 = x244 | n42854 ;
  assign n42856 = ~n42853 & n42855 ;
  assign n42857 = ( x580 & ~n42820 ) | ( x580 & n42856 ) | ( ~n42820 & n42856 ) ;
  assign n42858 = ( x245 & ~n42820 ) | ( x245 & n42857 ) | ( ~n42820 & n42857 ) ;
  assign n42859 = x552 & n42858 ;
  assign n42860 = x247 & ~n42859 ;
  assign n42861 = x244 | x566 ;
  assign n42862 = x235 | x531 ;
  assign n42863 = x242 | x556 ;
  assign n42864 = x242 & x556 ;
  assign n42865 = n42863 & ~n42864 ;
  assign n42866 = x239 & ~x569 ;
  assign n42867 = ~x246 & x564 ;
  assign n42868 = ( x249 & ~x482 ) | ( x249 & n42867 ) | ( ~x482 & n42867 ) ;
  assign n42869 = x241 & x562 ;
  assign n42870 = x241 | x562 ;
  assign n42871 = ~n42869 & n42870 ;
  assign n42872 = ( ~x249 & x482 ) | ( ~x249 & n42871 ) | ( x482 & n42871 ) ;
  assign n42873 = n42868 | n42872 ;
  assign n42874 = ( x570 & ~n42284 ) | ( x570 & n42873 ) | ( ~n42284 & n42873 ) ;
  assign n42875 = ( x570 & n41858 ) | ( x570 & ~n42873 ) | ( n41858 & ~n42873 ) ;
  assign n42876 = ~n42874 & n42875 ;
  assign n42877 = x246 & ~x564 ;
  assign n42878 = x248 & ~x565 ;
  assign n42879 = ~x248 & x565 ;
  assign n42880 = n42878 | n42879 ;
  assign n42881 = n42877 | n42880 ;
  assign n42882 = x560 & ~n42881 ;
  assign n42883 = ( ~x240 & n42876 ) | ( ~x240 & n42882 ) | ( n42876 & n42882 ) ;
  assign n42884 = ( ~x240 & x560 ) | ( ~x240 & n42877 ) | ( x560 & n42877 ) ;
  assign n42885 = ( x240 & ~x560 ) | ( x240 & n42880 ) | ( ~x560 & n42880 ) ;
  assign n42886 = n42884 | n42885 ;
  assign n42887 = ( x240 & n42876 ) | ( x240 & ~n42886 ) | ( n42876 & ~n42886 ) ;
  assign n42888 = n42883 & n42887 ;
  assign n42889 = ( x569 & n42866 ) | ( x569 & n42888 ) | ( n42866 & n42888 ) ;
  assign n42890 = ( ~x239 & n42866 ) | ( ~x239 & n42889 ) | ( n42866 & n42889 ) ;
  assign n42891 = ~n42865 & n42890 ;
  assign n42892 = ( x531 & ~n42862 ) | ( x531 & n42891 ) | ( ~n42862 & n42891 ) ;
  assign n42893 = ( x235 & ~n42862 ) | ( x235 & n42892 ) | ( ~n42862 & n42892 ) ;
  assign n42894 = ( x566 & ~n42861 ) | ( x566 & n42893 ) | ( ~n42861 & n42893 ) ;
  assign n42895 = ( x244 & ~n42861 ) | ( x244 & n42894 ) | ( ~n42861 & n42894 ) ;
  assign n42896 = x568 & n42895 ;
  assign n42897 = x245 & ~n42896 ;
  assign n42898 = ~x568 & n42895 ;
  assign n42899 = x245 | n42898 ;
  assign n42900 = ~n42897 & n42899 ;
  assign n42901 = ( x247 & x552 ) | ( x247 & n42900 ) | ( x552 & n42900 ) ;
  assign n42902 = ( x245 & x568 ) | ( x245 & n42856 ) | ( x568 & n42856 ) ;
  assign n42903 = ( x244 & x486 ) | ( x244 & n42893 ) | ( x486 & n42893 ) ;
  assign n42904 = ( x235 & x549 ) | ( x235 & n42891 ) | ( x549 & n42891 ) ;
  assign n42905 = n42843 & n42863 ;
  assign n42906 = ( x489 & x556 ) | ( x489 & ~n42890 ) | ( x556 & ~n42890 ) ;
  assign n42907 = x569 & ~n42840 ;
  assign n42908 = n42888 & n42907 ;
  assign n42909 = n42876 & ~n42886 ;
  assign n42910 = n42866 & n42909 ;
  assign n42911 = n42841 | n42910 ;
  assign n42912 = n42908 | n42911 ;
  assign n42913 = ( x489 & ~x556 ) | ( x489 & n42912 ) | ( ~x556 & n42912 ) ;
  assign n42914 = ~n42906 & n42913 ;
  assign n42915 = n42905 | n42914 ;
  assign n42916 = n42845 | n42864 ;
  assign n42917 = ( x489 & x556 ) | ( x489 & n42890 ) | ( x556 & n42890 ) ;
  assign n42918 = ( ~x489 & x556 ) | ( ~x489 & n42912 ) | ( x556 & n42912 ) ;
  assign n42919 = n42917 & n42918 ;
  assign n42920 = n42916 & ~n42919 ;
  assign n42921 = n42915 & ~n42920 ;
  assign n42922 = ( x235 & ~x549 ) | ( x235 & n42921 ) | ( ~x549 & n42921 ) ;
  assign n42923 = n42904 | n42922 ;
  assign n42924 = ~n42848 & n42923 ;
  assign n42925 = x531 | n42924 ;
  assign n42926 = ( ~x235 & x549 ) | ( ~x235 & n42921 ) | ( x549 & n42921 ) ;
  assign n42927 = ( x235 & x549 ) | ( x235 & ~n42891 ) | ( x549 & ~n42891 ) ;
  assign n42928 = ~n42926 & n42927 ;
  assign n42929 = n42850 & ~n42928 ;
  assign n42930 = x531 & ~n42929 ;
  assign n42931 = n42925 & ~n42930 ;
  assign n42932 = ( x244 & ~x486 ) | ( x244 & n42931 ) | ( ~x486 & n42931 ) ;
  assign n42933 = n42903 | n42932 ;
  assign n42934 = ~n42853 & n42933 ;
  assign n42935 = x566 | n42934 ;
  assign n42936 = ( ~x244 & x486 ) | ( ~x244 & n42931 ) | ( x486 & n42931 ) ;
  assign n42937 = ( x244 & x486 ) | ( x244 & ~n42893 ) | ( x486 & ~n42893 ) ;
  assign n42938 = ~n42936 & n42937 ;
  assign n42939 = n42855 & ~n42938 ;
  assign n42940 = x566 & ~n42939 ;
  assign n42941 = n42935 & ~n42940 ;
  assign n42942 = ( x245 & ~x568 ) | ( x245 & n42941 ) | ( ~x568 & n42941 ) ;
  assign n42943 = n42902 | n42942 ;
  assign n42944 = ~n42897 & n42943 ;
  assign n42945 = x580 | n42944 ;
  assign n42946 = ( ~x245 & x568 ) | ( ~x245 & n42941 ) | ( x568 & n42941 ) ;
  assign n42947 = ( x245 & x568 ) | ( x245 & ~n42856 ) | ( x568 & ~n42856 ) ;
  assign n42948 = ~n42946 & n42947 ;
  assign n42949 = n42899 & ~n42948 ;
  assign n42950 = x580 & ~n42949 ;
  assign n42951 = n42945 & ~n42950 ;
  assign n42952 = ( x247 & ~x552 ) | ( x247 & n42951 ) | ( ~x552 & n42951 ) ;
  assign n42953 = n42901 | n42952 ;
  assign n42954 = ~n42860 & n42953 ;
  assign n42955 = x532 | n42954 ;
  assign n42956 = ~x552 & n42858 ;
  assign n42957 = x247 | n42956 ;
  assign n42958 = ( ~x247 & x552 ) | ( ~x247 & n42951 ) | ( x552 & n42951 ) ;
  assign n42959 = ( x247 & x552 ) | ( x247 & ~n42900 ) | ( x552 & ~n42900 ) ;
  assign n42960 = ~n42958 & n42959 ;
  assign n42961 = n42957 & ~n42960 ;
  assign n42962 = x532 & ~n42961 ;
  assign n42963 = n42955 & ~n42962 ;
  assign n42964 = ~x238 & n42963 ;
  assign n42965 = x577 | n42964 ;
  assign n42966 = x247 | x532 ;
  assign n42967 = ( x532 & n42900 ) | ( x532 & ~n42966 ) | ( n42900 & ~n42966 ) ;
  assign n42968 = ( x247 & ~n42966 ) | ( x247 & n42967 ) | ( ~n42966 & n42967 ) ;
  assign n42969 = ( x238 & x577 ) | ( x238 & ~n42968 ) | ( x577 & ~n42968 ) ;
  assign n42970 = ~n42860 & n42957 ;
  assign n42971 = ( x238 & ~x577 ) | ( x238 & n42970 ) | ( ~x577 & n42970 ) ;
  assign n42972 = n42969 & ~n42971 ;
  assign n42973 = x498 | n42972 ;
  assign n42974 = n42965 & ~n42973 ;
  assign n42975 = x238 & n42963 ;
  assign n42976 = x577 & ~n42975 ;
  assign n42977 = ( x238 & x577 ) | ( x238 & n42968 ) | ( x577 & n42968 ) ;
  assign n42978 = ( ~x238 & x577 ) | ( ~x238 & n42970 ) | ( x577 & n42970 ) ;
  assign n42979 = n42977 | n42978 ;
  assign n42980 = x498 & n42979 ;
  assign n42981 = ~n42976 & n42980 ;
  assign n42982 = n42974 | n42981 ;
  assign n42983 = ( ~x233 & x237 ) | ( ~x233 & n42982 ) | ( x237 & n42982 ) ;
  assign n42984 = n42819 | n42983 ;
  assign n42985 = ~n42630 & n42984 ;
  assign n42986 = ~x806 & n41539 ;
  assign n42987 = x332 | x806 ;
  assign n42988 = x990 & ~n42987 ;
  assign n42989 = x600 & n42988 ;
  assign n42990 = ~x332 & x594 ;
  assign n42991 = n42989 | n42990 ;
  assign n42992 = ~n42986 & n42991 ;
  assign n42993 = x605 & ~x806 ;
  assign n42994 = n41522 & n42993 ;
  assign n42995 = x595 & ~n42994 ;
  assign n42996 = ( x332 & x595 ) | ( x332 & ~n42995 ) | ( x595 & ~n42995 ) ;
  assign n42997 = ( n42994 & n42995 ) | ( n42994 & ~n42996 ) | ( n42995 & ~n42996 ) ;
  assign n42998 = ~x332 & x596 ;
  assign n42999 = x595 & n41521 ;
  assign n43000 = n42988 & n42999 ;
  assign n43001 = n42998 | n43000 ;
  assign n43002 = x596 & n43000 ;
  assign n43003 = n43001 & ~n43002 ;
  assign n43004 = x597 & ~n42986 ;
  assign n43005 = ( x332 & x597 ) | ( x332 & ~n43004 ) | ( x597 & ~n43004 ) ;
  assign n43006 = ( n42986 & n43004 ) | ( n42986 & ~n43005 ) | ( n43004 & ~n43005 ) ;
  assign n43007 = x882 | n6785 ;
  assign n43008 = x947 & ~n43007 ;
  assign n43009 = x598 & ~n43008 ;
  assign n43010 = x740 & x780 ;
  assign n43011 = n4708 & n43010 ;
  assign n43012 = n43009 | n43011 ;
  assign n43013 = ~x332 & x599 ;
  assign n43014 = n43002 | n43013 ;
  assign n43015 = x599 & n43002 ;
  assign n43016 = n43014 & ~n43015 ;
  assign n43017 = ~x332 & x600 ;
  assign n43018 = n42988 | n43017 ;
  assign n43019 = ~n42989 & n43018 ;
  assign n43020 = ( ~x332 & x806 ) | ( ~x332 & x989 ) | ( x806 & x989 ) ;
  assign n43021 = ( x332 & ~x601 ) | ( x332 & x806 ) | ( ~x601 & x806 ) ;
  assign n43022 = n43020 & ~n43021 ;
  assign n43023 = ~x230 & x602 ;
  assign n43024 = x230 & n15171 ;
  assign n43025 = ~n16054 & n43024 ;
  assign n43026 = x715 | x1160 ;
  assign n43027 = n17210 | n17389 ;
  assign n43028 = ( x715 & ~x790 ) | ( x715 & x1160 ) | ( ~x790 & x1160 ) ;
  assign n43029 = ( n43026 & n43027 ) | ( n43026 & ~n43028 ) | ( n43027 & ~n43028 ) ;
  assign n43030 = n43025 & ~n43029 ;
  assign n43031 = ~n17215 & n43030 ;
  assign n43032 = n43023 | n43031 ;
  assign n43033 = ~x980 & x1038 ;
  assign n43034 = x1060 & n43033 ;
  assign n43035 = x952 & ~x1061 ;
  assign n43036 = n43034 & n43035 ;
  assign n43037 = x832 & n43036 ;
  assign n43038 = x603 | n43037 ;
  assign n43039 = x832 & ~x1100 ;
  assign n43040 = n43036 & n43039 ;
  assign n43041 = x966 | n43040 ;
  assign n43042 = n43038 & ~n43041 ;
  assign n43043 = x871 & x966 ;
  assign n43044 = x872 & x966 ;
  assign n43045 = n43043 | n43044 ;
  assign n43046 = n43042 | n43045 ;
  assign n43047 = x823 & ~n14553 ;
  assign n43048 = ~x779 & n43047 ;
  assign n43049 = ~x299 & x983 ;
  assign n43050 = x907 & n43049 ;
  assign n43051 = x604 & ~n43050 ;
  assign n43052 = ~n43047 & n43051 ;
  assign n43053 = n43048 | n43052 ;
  assign n43054 = ~x605 & n42987 ;
  assign n43055 = x332 | n42993 ;
  assign n43056 = n43054 | n43055 ;
  assign n43057 = ~x837 & x966 ;
  assign n43058 = ( x966 & x1104 ) | ( x966 & n43037 ) | ( x1104 & n43037 ) ;
  assign n43059 = ( x606 & x966 ) | ( x606 & ~n43037 ) | ( x966 & ~n43037 ) ;
  assign n43060 = n43058 | n43059 ;
  assign n43061 = ~n43057 & n43060 ;
  assign n43062 = ( x966 & ~x1107 ) | ( x966 & n43037 ) | ( ~x1107 & n43037 ) ;
  assign n43063 = ( x607 & ~x966 ) | ( x607 & n43037 ) | ( ~x966 & n43037 ) ;
  assign n43064 = ~n43062 & n43063 ;
  assign n43065 = ( x966 & ~x1116 ) | ( x966 & n43037 ) | ( ~x1116 & n43037 ) ;
  assign n43066 = ( x608 & ~x966 ) | ( x608 & n43037 ) | ( ~x966 & n43037 ) ;
  assign n43067 = ~n43065 & n43066 ;
  assign n43068 = ( x966 & ~x1118 ) | ( x966 & n43037 ) | ( ~x1118 & n43037 ) ;
  assign n43069 = ( x609 & ~x966 ) | ( x609 & n43037 ) | ( ~x966 & n43037 ) ;
  assign n43070 = ~n43068 & n43069 ;
  assign n43071 = ( x966 & ~x1113 ) | ( x966 & n43037 ) | ( ~x1113 & n43037 ) ;
  assign n43072 = ( x610 & ~x966 ) | ( x610 & n43037 ) | ( ~x966 & n43037 ) ;
  assign n43073 = ~n43071 & n43072 ;
  assign n43074 = ( x966 & ~x1114 ) | ( x966 & n43037 ) | ( ~x1114 & n43037 ) ;
  assign n43075 = ( x611 & ~x966 ) | ( x611 & n43037 ) | ( ~x966 & n43037 ) ;
  assign n43076 = ~n43074 & n43075 ;
  assign n43077 = ( x966 & ~x1111 ) | ( x966 & n43037 ) | ( ~x1111 & n43037 ) ;
  assign n43078 = ( x612 & ~x966 ) | ( x612 & n43037 ) | ( ~x966 & n43037 ) ;
  assign n43079 = ~n43077 & n43078 ;
  assign n43080 = ( x966 & ~x1115 ) | ( x966 & n43037 ) | ( ~x1115 & n43037 ) ;
  assign n43081 = ( x613 & ~x966 ) | ( x613 & n43037 ) | ( ~x966 & n43037 ) ;
  assign n43082 = ~n43080 & n43081 ;
  assign n43083 = ( x966 & ~x1102 ) | ( x966 & n43037 ) | ( ~x1102 & n43037 ) ;
  assign n43084 = ( x614 & ~x966 ) | ( x614 & n43037 ) | ( ~x966 & n43037 ) ;
  assign n43085 = ~n43083 & n43084 ;
  assign n43086 = n43043 | n43085 ;
  assign n43087 = x907 & ~n43007 ;
  assign n43088 = x615 | n43087 ;
  assign n43089 = x779 & x797 ;
  assign n43090 = n4711 & n43089 ;
  assign n43091 = n43088 & ~n43090 ;
  assign n43092 = ( x966 & ~x1101 ) | ( x966 & n43037 ) | ( ~x1101 & n43037 ) ;
  assign n43093 = ( x616 & ~x966 ) | ( x616 & n43037 ) | ( ~x966 & n43037 ) ;
  assign n43094 = ~n43092 & n43093 ;
  assign n43095 = n43044 | n43094 ;
  assign n43096 = ~x850 & x966 ;
  assign n43097 = ( x966 & x1105 ) | ( x966 & n43037 ) | ( x1105 & n43037 ) ;
  assign n43098 = ( x617 & x966 ) | ( x617 & ~n43037 ) | ( x966 & ~n43037 ) ;
  assign n43099 = n43097 | n43098 ;
  assign n43100 = ~n43096 & n43099 ;
  assign n43101 = ( x966 & ~x1117 ) | ( x966 & n43037 ) | ( ~x1117 & n43037 ) ;
  assign n43102 = ( x618 & ~x966 ) | ( x618 & n43037 ) | ( ~x966 & n43037 ) ;
  assign n43103 = ~n43101 & n43102 ;
  assign n43104 = ( x966 & ~x1122 ) | ( x966 & n43037 ) | ( ~x1122 & n43037 ) ;
  assign n43105 = ( x619 & ~x966 ) | ( x619 & n43037 ) | ( ~x966 & n43037 ) ;
  assign n43106 = ~n43104 & n43105 ;
  assign n43107 = ( x966 & ~x1112 ) | ( x966 & n43037 ) | ( ~x1112 & n43037 ) ;
  assign n43108 = ( x620 & ~x966 ) | ( x620 & n43037 ) | ( ~x966 & n43037 ) ;
  assign n43109 = ~n43107 & n43108 ;
  assign n43110 = ( x966 & ~x1108 ) | ( x966 & n43037 ) | ( ~x1108 & n43037 ) ;
  assign n43111 = ( x621 & ~x966 ) | ( x621 & n43037 ) | ( ~x966 & n43037 ) ;
  assign n43112 = ~n43110 & n43111 ;
  assign n43113 = ( x966 & ~x1109 ) | ( x966 & n43037 ) | ( ~x1109 & n43037 ) ;
  assign n43114 = ( x622 & ~x966 ) | ( x622 & n43037 ) | ( ~x966 & n43037 ) ;
  assign n43115 = ~n43113 & n43114 ;
  assign n43116 = ( x966 & ~x1106 ) | ( x966 & n43037 ) | ( ~x1106 & n43037 ) ;
  assign n43117 = ( x623 & ~x966 ) | ( x623 & n43037 ) | ( ~x966 & n43037 ) ;
  assign n43118 = ~n43116 & n43117 ;
  assign n43119 = x831 & ~n14855 ;
  assign n43120 = ~x780 & n43119 ;
  assign n43121 = x947 & n43049 ;
  assign n43122 = x624 & ~n43121 ;
  assign n43123 = ~n43119 & n43122 ;
  assign n43124 = n43120 | n43123 ;
  assign n43125 = x832 & ~x973 ;
  assign n43126 = ~x1054 & x1066 ;
  assign n43127 = x1088 & n43126 ;
  assign n43128 = n43125 & n43127 ;
  assign n43129 = ~x953 & n43128 ;
  assign n43130 = ( x962 & ~x1116 ) | ( x962 & n43129 ) | ( ~x1116 & n43129 ) ;
  assign n43131 = ( x625 & ~x962 ) | ( x625 & n43129 ) | ( ~x962 & n43129 ) ;
  assign n43132 = ~n43130 & n43131 ;
  assign n43133 = ( x966 & ~x1121 ) | ( x966 & n43037 ) | ( ~x1121 & n43037 ) ;
  assign n43134 = ( x626 & ~x966 ) | ( x626 & n43037 ) | ( ~x966 & n43037 ) ;
  assign n43135 = ~n43133 & n43134 ;
  assign n43136 = ( x962 & ~x1117 ) | ( x962 & n43129 ) | ( ~x1117 & n43129 ) ;
  assign n43137 = ( x627 & ~x962 ) | ( x627 & n43129 ) | ( ~x962 & n43129 ) ;
  assign n43138 = ~n43136 & n43137 ;
  assign n43139 = ( x962 & ~x1119 ) | ( x962 & n43129 ) | ( ~x1119 & n43129 ) ;
  assign n43140 = ( x628 & ~x962 ) | ( x628 & n43129 ) | ( ~x962 & n43129 ) ;
  assign n43141 = ~n43139 & n43140 ;
  assign n43142 = ( x966 & ~x1119 ) | ( x966 & n43037 ) | ( ~x1119 & n43037 ) ;
  assign n43143 = ( x629 & ~x966 ) | ( x629 & n43037 ) | ( ~x966 & n43037 ) ;
  assign n43144 = ~n43142 & n43143 ;
  assign n43145 = ( x966 & ~x1120 ) | ( x966 & n43037 ) | ( ~x1120 & n43037 ) ;
  assign n43146 = ( x630 & ~x966 ) | ( x630 & n43037 ) | ( ~x966 & n43037 ) ;
  assign n43147 = ~n43145 & n43146 ;
  assign n43148 = ( x962 & ~x1113 ) | ( x962 & n43129 ) | ( ~x1113 & n43129 ) ;
  assign n43149 = ( x631 & x962 ) | ( x631 & ~n43129 ) | ( x962 & ~n43129 ) ;
  assign n43150 = n43148 | n43149 ;
  assign n43151 = ( x962 & ~x1115 ) | ( x962 & n43129 ) | ( ~x1115 & n43129 ) ;
  assign n43152 = ( x632 & x962 ) | ( x632 & ~n43129 ) | ( x962 & ~n43129 ) ;
  assign n43153 = n43151 | n43152 ;
  assign n43154 = ( x966 & ~x1110 ) | ( x966 & n43037 ) | ( ~x1110 & n43037 ) ;
  assign n43155 = ( x633 & ~x966 ) | ( x633 & n43037 ) | ( ~x966 & n43037 ) ;
  assign n43156 = ~n43154 & n43155 ;
  assign n43157 = ( x962 & ~x1110 ) | ( x962 & n43129 ) | ( ~x1110 & n43129 ) ;
  assign n43158 = ( x634 & ~x962 ) | ( x634 & n43129 ) | ( ~x962 & n43129 ) ;
  assign n43159 = ~n43157 & n43158 ;
  assign n43160 = ( x962 & ~x1112 ) | ( x962 & n43129 ) | ( ~x1112 & n43129 ) ;
  assign n43161 = ( x635 & x962 ) | ( x635 & ~n43129 ) | ( x962 & ~n43129 ) ;
  assign n43162 = n43160 | n43161 ;
  assign n43163 = ( x966 & ~x1127 ) | ( x966 & n43037 ) | ( ~x1127 & n43037 ) ;
  assign n43164 = ( x636 & ~x966 ) | ( x636 & n43037 ) | ( ~x966 & n43037 ) ;
  assign n43165 = ~n43163 & n43164 ;
  assign n43166 = ( x962 & ~x1105 ) | ( x962 & n43129 ) | ( ~x1105 & n43129 ) ;
  assign n43167 = ( x637 & ~x962 ) | ( x637 & n43129 ) | ( ~x962 & n43129 ) ;
  assign n43168 = ~n43166 & n43167 ;
  assign n43169 = ( x962 & ~x1107 ) | ( x962 & n43129 ) | ( ~x1107 & n43129 ) ;
  assign n43170 = ( x638 & ~x962 ) | ( x638 & n43129 ) | ( ~x962 & n43129 ) ;
  assign n43171 = ~n43169 & n43170 ;
  assign n43172 = ( x962 & ~x1109 ) | ( x962 & n43129 ) | ( ~x1109 & n43129 ) ;
  assign n43173 = ( x639 & ~x962 ) | ( x639 & n43129 ) | ( ~x962 & n43129 ) ;
  assign n43174 = ~n43172 & n43173 ;
  assign n43175 = ( x966 & ~x1128 ) | ( x966 & n43037 ) | ( ~x1128 & n43037 ) ;
  assign n43176 = ( x640 & ~x966 ) | ( x640 & n43037 ) | ( ~x966 & n43037 ) ;
  assign n43177 = ~n43175 & n43176 ;
  assign n43178 = ( x962 & ~x1121 ) | ( x962 & n43129 ) | ( ~x1121 & n43129 ) ;
  assign n43179 = ( x641 & ~x962 ) | ( x641 & n43129 ) | ( ~x962 & n43129 ) ;
  assign n43180 = ~n43178 & n43179 ;
  assign n43181 = ( x966 & ~x1103 ) | ( x966 & n43037 ) | ( ~x1103 & n43037 ) ;
  assign n43182 = ( x642 & ~x966 ) | ( x642 & n43037 ) | ( ~x966 & n43037 ) ;
  assign n43183 = ~n43181 & n43182 ;
  assign n43184 = ( x962 & ~x1104 ) | ( x962 & n43129 ) | ( ~x1104 & n43129 ) ;
  assign n43185 = ( x643 & ~x962 ) | ( x643 & n43129 ) | ( ~x962 & n43129 ) ;
  assign n43186 = ~n43184 & n43185 ;
  assign n43187 = ( x966 & ~x1123 ) | ( x966 & n43037 ) | ( ~x1123 & n43037 ) ;
  assign n43188 = ( x644 & ~x966 ) | ( x644 & n43037 ) | ( ~x966 & n43037 ) ;
  assign n43189 = ~n43187 & n43188 ;
  assign n43190 = ( x966 & ~x1125 ) | ( x966 & n43037 ) | ( ~x1125 & n43037 ) ;
  assign n43191 = ( x645 & ~x966 ) | ( x645 & n43037 ) | ( ~x966 & n43037 ) ;
  assign n43192 = ~n43190 & n43191 ;
  assign n43193 = ( x962 & ~x1114 ) | ( x962 & n43129 ) | ( ~x1114 & n43129 ) ;
  assign n43194 = ( x646 & x962 ) | ( x646 & ~n43129 ) | ( x962 & ~n43129 ) ;
  assign n43195 = n43193 | n43194 ;
  assign n43196 = ( x962 & ~x1120 ) | ( x962 & n43129 ) | ( ~x1120 & n43129 ) ;
  assign n43197 = ( x647 & ~x962 ) | ( x647 & n43129 ) | ( ~x962 & n43129 ) ;
  assign n43198 = ~n43196 & n43197 ;
  assign n43199 = ( x962 & ~x1122 ) | ( x962 & n43129 ) | ( ~x1122 & n43129 ) ;
  assign n43200 = ( x648 & ~x962 ) | ( x648 & n43129 ) | ( ~x962 & n43129 ) ;
  assign n43201 = ~n43199 & n43200 ;
  assign n43202 = ( x962 & ~x1126 ) | ( x962 & n43129 ) | ( ~x1126 & n43129 ) ;
  assign n43203 = ( x649 & x962 ) | ( x649 & ~n43129 ) | ( x962 & ~n43129 ) ;
  assign n43204 = n43202 | n43203 ;
  assign n43205 = ( x962 & ~x1127 ) | ( x962 & n43129 ) | ( ~x1127 & n43129 ) ;
  assign n43206 = ( x650 & x962 ) | ( x650 & ~n43129 ) | ( x962 & ~n43129 ) ;
  assign n43207 = n43205 | n43206 ;
  assign n43208 = ( x966 & ~x1130 ) | ( x966 & n43037 ) | ( ~x1130 & n43037 ) ;
  assign n43209 = ( x651 & ~x966 ) | ( x651 & n43037 ) | ( ~x966 & n43037 ) ;
  assign n43210 = ~n43208 & n43209 ;
  assign n43211 = ( x966 & ~x1131 ) | ( x966 & n43037 ) | ( ~x1131 & n43037 ) ;
  assign n43212 = ( x652 & ~x966 ) | ( x652 & n43037 ) | ( ~x966 & n43037 ) ;
  assign n43213 = ~n43211 & n43212 ;
  assign n43214 = ( x966 & ~x1129 ) | ( x966 & n43037 ) | ( ~x1129 & n43037 ) ;
  assign n43215 = ( x653 & ~x966 ) | ( x653 & n43037 ) | ( ~x966 & n43037 ) ;
  assign n43216 = ~n43214 & n43215 ;
  assign n43217 = ( x962 & ~x1130 ) | ( x962 & n43129 ) | ( ~x1130 & n43129 ) ;
  assign n43218 = ( x654 & x962 ) | ( x654 & ~n43129 ) | ( x962 & ~n43129 ) ;
  assign n43219 = n43217 | n43218 ;
  assign n43220 = ( x962 & ~x1124 ) | ( x962 & n43129 ) | ( ~x1124 & n43129 ) ;
  assign n43221 = ( x655 & x962 ) | ( x655 & ~n43129 ) | ( x962 & ~n43129 ) ;
  assign n43222 = n43220 | n43221 ;
  assign n43223 = ( x966 & ~x1126 ) | ( x966 & n43037 ) | ( ~x1126 & n43037 ) ;
  assign n43224 = ( x656 & ~x966 ) | ( x656 & n43037 ) | ( ~x966 & n43037 ) ;
  assign n43225 = ~n43223 & n43224 ;
  assign n43226 = ( x962 & ~x1131 ) | ( x962 & n43129 ) | ( ~x1131 & n43129 ) ;
  assign n43227 = ( x657 & x962 ) | ( x657 & ~n43129 ) | ( x962 & ~n43129 ) ;
  assign n43228 = n43226 | n43227 ;
  assign n43229 = ( x966 & ~x1124 ) | ( x966 & n43037 ) | ( ~x1124 & n43037 ) ;
  assign n43230 = ( x658 & ~x966 ) | ( x658 & n43037 ) | ( ~x966 & n43037 ) ;
  assign n43231 = ~n43229 & n43230 ;
  assign n43232 = x266 & x992 ;
  assign n43233 = ~x280 & n43232 ;
  assign n43234 = ~x269 & n43233 ;
  assign n43235 = ~x281 & n43234 ;
  assign n43236 = x270 | x277 ;
  assign n43237 = x282 | n43236 ;
  assign n43238 = n43235 & ~n43237 ;
  assign n43239 = ~x264 & n43238 ;
  assign n43240 = ~x265 & n43239 ;
  assign n43241 = ~x274 & n43240 ;
  assign n43242 = x274 & ~n43240 ;
  assign n43243 = n43241 | n43242 ;
  assign n43244 = ( x962 & ~x1118 ) | ( x962 & n43129 ) | ( ~x1118 & n43129 ) ;
  assign n43245 = ( x660 & ~x962 ) | ( x660 & n43129 ) | ( ~x962 & n43129 ) ;
  assign n43246 = ~n43244 & n43245 ;
  assign n43247 = ( x962 & ~x1101 ) | ( x962 & n43129 ) | ( ~x1101 & n43129 ) ;
  assign n43248 = ( x661 & ~x962 ) | ( x661 & n43129 ) | ( ~x962 & n43129 ) ;
  assign n43249 = ~n43247 & n43248 ;
  assign n43250 = ( x962 & ~x1102 ) | ( x962 & n43129 ) | ( ~x1102 & n43129 ) ;
  assign n43251 = ( x662 & ~x962 ) | ( x662 & n43129 ) | ( ~x962 & n43129 ) ;
  assign n43252 = ~n43250 & n43251 ;
  assign n43253 = ~x591 & x592 ;
  assign n43254 = x365 & n43253 ;
  assign n43255 = x334 & x591 ;
  assign n43256 = ~x592 & n43255 ;
  assign n43257 = n43254 | n43256 ;
  assign n43258 = ~x590 & n43257 ;
  assign n43259 = x591 | x592 ;
  assign n43260 = x590 & ~n43259 ;
  assign n43261 = x323 & n43260 ;
  assign n43262 = x588 | n43261 ;
  assign n43263 = n43258 | n43262 ;
  assign n43264 = x223 | x224 ;
  assign n43265 = x592 | n6278 ;
  assign n43266 = x464 & ~n43265 ;
  assign n43267 = x588 & ~n43266 ;
  assign n43268 = n43264 | n43267 ;
  assign n43269 = n43263 & ~n43268 ;
  assign n43270 = ( x199 & x257 ) | ( x199 & n43264 ) | ( x257 & n43264 ) ;
  assign n43271 = ( ~x199 & x1065 ) | ( ~x199 & n43264 ) | ( x1065 & n43264 ) ;
  assign n43272 = n43270 & n43271 ;
  assign n43273 = n43269 | n43272 ;
  assign n43274 = ~n7103 & n43273 ;
  assign n43275 = x1137 | x1138 ;
  assign n43276 = x1134 | n43275 ;
  assign n43277 = ( x634 & x1135 ) | ( x634 & ~x1136 ) | ( x1135 & ~x1136 ) ;
  assign n43278 = ( x784 & x1135 ) | ( x784 & x1136 ) | ( x1135 & x1136 ) ;
  assign n43279 = n43277 & n43278 ;
  assign n43280 = ( ~x633 & x1135 ) | ( ~x633 & x1136 ) | ( x1135 & x1136 ) ;
  assign n43281 = ( x815 & ~x1135 ) | ( x815 & x1136 ) | ( ~x1135 & x1136 ) ;
  assign n43282 = ~n43280 & n43281 ;
  assign n43283 = n43279 | n43282 ;
  assign n43284 = ~n43276 & n43283 ;
  assign n43285 = x1135 & ~n43275 ;
  assign n43286 = x1136 & ~n43285 ;
  assign n43287 = ~x766 & n43286 ;
  assign n43288 = x1135 & ~x1136 ;
  assign n43289 = x1134 & ~n43275 ;
  assign n43290 = ~n43288 & n43289 ;
  assign n43291 = x855 | x1136 ;
  assign n43292 = ~x700 & x1135 ;
  assign n43293 = n43291 & ~n43292 ;
  assign n43294 = n43290 & n43293 ;
  assign n43295 = ~n43287 & n43294 ;
  assign n43296 = n43284 | n43295 ;
  assign n43297 = n7103 & n43296 ;
  assign n43298 = n43274 | n43297 ;
  assign n43299 = x355 & n43260 ;
  assign n43300 = x404 & n10558 ;
  assign n43301 = ~x590 & x592 ;
  assign n43302 = x588 | n43301 ;
  assign n43303 = n43300 | n43302 ;
  assign n43304 = x380 & n43253 ;
  assign n43305 = ( ~x592 & n43303 ) | ( ~x592 & n43304 ) | ( n43303 & n43304 ) ;
  assign n43306 = n43299 | n43305 ;
  assign n43307 = x429 & ~n43265 ;
  assign n43308 = x588 & ~n43307 ;
  assign n43309 = n43264 | n43308 ;
  assign n43310 = n43306 & ~n43309 ;
  assign n43311 = ( x199 & x292 ) | ( x199 & n43264 ) | ( x292 & n43264 ) ;
  assign n43312 = ( ~x199 & x1084 ) | ( ~x199 & n43264 ) | ( x1084 & n43264 ) ;
  assign n43313 = n43311 & n43312 ;
  assign n43314 = n43310 | n43313 ;
  assign n43315 = ~n7103 & n43314 ;
  assign n43316 = ( ~x614 & x1135 ) | ( ~x614 & x1136 ) | ( x1135 & x1136 ) ;
  assign n43317 = ( x662 & x1135 ) | ( x662 & ~x1136 ) | ( x1135 & ~x1136 ) ;
  assign n43318 = n43316 & ~n43317 ;
  assign n43319 = ( x785 & x1135 ) | ( x785 & x1136 ) | ( x1135 & x1136 ) ;
  assign n43320 = ( x811 & ~x1135 ) | ( x811 & x1136 ) | ( ~x1135 & x1136 ) ;
  assign n43321 = n43319 | n43320 ;
  assign n43322 = ~n43318 & n43321 ;
  assign n43323 = x1134 | n43322 ;
  assign n43324 = x1135 | x1136 ;
  assign n43325 = x872 & ~n43324 ;
  assign n43326 = x1134 & ~n43325 ;
  assign n43327 = ( x772 & x1135 ) | ( x772 & x1136 ) | ( x1135 & x1136 ) ;
  assign n43328 = ( x727 & ~x1135 ) | ( x727 & x1136 ) | ( ~x1135 & x1136 ) ;
  assign n43329 = n43327 & n43328 ;
  assign n43330 = n43326 & ~n43329 ;
  assign n43331 = n7103 & ~n43275 ;
  assign n43332 = ~n43330 & n43331 ;
  assign n43333 = n43323 & n43332 ;
  assign n43334 = n43315 | n43333 ;
  assign n43335 = ( x962 & ~x1108 ) | ( x962 & n43129 ) | ( ~x1108 & n43129 ) ;
  assign n43336 = ( x665 & ~x962 ) | ( x665 & n43129 ) | ( ~x962 & n43129 ) ;
  assign n43337 = ~n43335 & n43336 ;
  assign n43338 = ( x607 & x1135 ) | ( x607 & x1136 ) | ( x1135 & x1136 ) ;
  assign n43339 = ( x638 & ~x1135 ) | ( x638 & x1136 ) | ( ~x1135 & x1136 ) ;
  assign n43340 = n43338 & n43339 ;
  assign n43341 = ( ~x790 & x1135 ) | ( ~x790 & x1136 ) | ( x1135 & x1136 ) ;
  assign n43342 = ( x799 & ~x1135 ) | ( x799 & x1136 ) | ( ~x1135 & x1136 ) ;
  assign n43343 = n43341 | n43342 ;
  assign n43344 = ~n43340 & n43343 ;
  assign n43345 = n43276 | n43344 ;
  assign n43346 = ~x764 & n43286 ;
  assign n43347 = ~x691 & x1135 ;
  assign n43348 = x873 | x1136 ;
  assign n43349 = ~n43347 & n43348 ;
  assign n43350 = n43290 & n43349 ;
  assign n43351 = ~n43346 & n43350 ;
  assign n43352 = n43345 & ~n43351 ;
  assign n43353 = n7103 & ~n43352 ;
  assign n43354 = x441 & n43260 ;
  assign n43355 = x456 & n10558 ;
  assign n43356 = n43302 | n43355 ;
  assign n43357 = x337 & n43253 ;
  assign n43358 = ( ~x592 & n43356 ) | ( ~x592 & n43357 ) | ( n43356 & n43357 ) ;
  assign n43359 = n43354 | n43358 ;
  assign n43360 = x443 & ~n43265 ;
  assign n43361 = x588 & ~n43360 ;
  assign n43362 = n43264 | n43361 ;
  assign n43363 = n43359 & ~n43362 ;
  assign n43364 = ( x199 & x297 ) | ( x199 & n43264 ) | ( x297 & n43264 ) ;
  assign n43365 = ( ~x199 & x1044 ) | ( ~x199 & n43264 ) | ( x1044 & n43264 ) ;
  assign n43366 = n43364 & n43365 ;
  assign n43367 = n43363 | n43366 ;
  assign n43368 = ~n7103 & n43367 ;
  assign n43369 = n43353 | n43368 ;
  assign n43370 = x458 & n43260 ;
  assign n43371 = x319 & n10558 ;
  assign n43372 = n43302 | n43371 ;
  assign n43373 = x338 & n43253 ;
  assign n43374 = ( ~x592 & n43372 ) | ( ~x592 & n43373 ) | ( n43372 & n43373 ) ;
  assign n43375 = n43370 | n43374 ;
  assign n43376 = x444 & ~n43265 ;
  assign n43377 = x588 & ~n43376 ;
  assign n43378 = n43264 | n43377 ;
  assign n43379 = n43375 & ~n43378 ;
  assign n43380 = ( x199 & x294 ) | ( x199 & n43264 ) | ( x294 & n43264 ) ;
  assign n43381 = ( ~x199 & x1072 ) | ( ~x199 & n43264 ) | ( x1072 & n43264 ) ;
  assign n43382 = n43380 & n43381 ;
  assign n43383 = n43379 | n43382 ;
  assign n43384 = ~n7103 & n43383 ;
  assign n43385 = ( x681 & ~x1135 ) | ( x681 & x1136 ) | ( ~x1135 & x1136 ) ;
  assign n43386 = ( ~x792 & x1135 ) | ( ~x792 & x1136 ) | ( x1135 & x1136 ) ;
  assign n43387 = ~n43385 & n43386 ;
  assign n43388 = ( x642 & x1135 ) | ( x642 & x1136 ) | ( x1135 & x1136 ) ;
  assign n43389 = ( x809 & ~x1135 ) | ( x809 & x1136 ) | ( ~x1135 & x1136 ) ;
  assign n43390 = ~n43388 & n43389 ;
  assign n43391 = n43387 | n43390 ;
  assign n43392 = ~x1134 & n43391 ;
  assign n43393 = x871 & ~n43324 ;
  assign n43394 = x1134 & ~n43393 ;
  assign n43395 = ( x763 & x1135 ) | ( x763 & x1136 ) | ( x1135 & x1136 ) ;
  assign n43396 = ( x699 & ~x1135 ) | ( x699 & x1136 ) | ( ~x1135 & x1136 ) ;
  assign n43397 = n43395 & n43396 ;
  assign n43398 = n43394 & ~n43397 ;
  assign n43399 = n43331 & ~n43398 ;
  assign n43400 = ~n43392 & n43399 ;
  assign n43401 = n43384 | n43400 ;
  assign n43402 = ( x603 & x1135 ) | ( x603 & x1136 ) | ( x1135 & x1136 ) ;
  assign n43403 = ( x680 & ~x1135 ) | ( x680 & x1136 ) | ( ~x1135 & x1136 ) ;
  assign n43404 = n43402 & n43403 ;
  assign n43405 = ( ~x778 & x1135 ) | ( ~x778 & x1136 ) | ( x1135 & x1136 ) ;
  assign n43406 = ( x981 & x1135 ) | ( x981 & ~x1136 ) | ( x1135 & ~x1136 ) ;
  assign n43407 = ~n43405 & n43406 ;
  assign n43408 = n43404 | n43407 ;
  assign n43409 = ~n43276 & n43408 ;
  assign n43410 = ~x759 & n43286 ;
  assign n43411 = ~x696 & x1135 ;
  assign n43412 = x837 | x1136 ;
  assign n43413 = ~n43411 & n43412 ;
  assign n43414 = n43290 & n43413 ;
  assign n43415 = ~n43410 & n43414 ;
  assign n43416 = n43409 | n43415 ;
  assign n43417 = n7103 & n43416 ;
  assign n43418 = x342 & n43260 ;
  assign n43419 = x390 & n10558 ;
  assign n43420 = n43302 | n43419 ;
  assign n43421 = x363 & n43253 ;
  assign n43422 = ( ~x592 & n43420 ) | ( ~x592 & n43421 ) | ( n43420 & n43421 ) ;
  assign n43423 = n43418 | n43422 ;
  assign n43424 = x414 & ~n43265 ;
  assign n43425 = x588 & ~n43424 ;
  assign n43426 = n43264 | n43425 ;
  assign n43427 = n43423 & ~n43426 ;
  assign n43428 = ( x199 & x291 ) | ( x199 & n43264 ) | ( x291 & n43264 ) ;
  assign n43429 = ( ~x199 & x1049 ) | ( ~x199 & n43264 ) | ( x1049 & n43264 ) ;
  assign n43430 = n43428 & n43429 ;
  assign n43431 = n43427 | n43430 ;
  assign n43432 = ~n7103 & n43431 ;
  assign n43433 = n43417 | n43432 ;
  assign n43434 = ( x962 & ~x1125 ) | ( x962 & n43129 ) | ( ~x1125 & n43129 ) ;
  assign n43435 = ( x669 & x962 ) | ( x669 & ~n43129 ) | ( x962 & ~n43129 ) ;
  assign n43436 = n43434 | n43435 ;
  assign n43437 = x364 & n43253 ;
  assign n43438 = x391 & x591 ;
  assign n43439 = ~x592 & n43438 ;
  assign n43440 = n43437 | n43439 ;
  assign n43441 = ~x590 & n43440 ;
  assign n43442 = x343 & n43260 ;
  assign n43443 = x588 | n43442 ;
  assign n43444 = n43441 | n43443 ;
  assign n43445 = x415 & ~n43265 ;
  assign n43446 = x588 & ~n43445 ;
  assign n43447 = n43264 | n43446 ;
  assign n43448 = n43444 & ~n43447 ;
  assign n43449 = ( x199 & x258 ) | ( x199 & n43264 ) | ( x258 & n43264 ) ;
  assign n43450 = ( ~x199 & x1062 ) | ( ~x199 & n43264 ) | ( x1062 & n43264 ) ;
  assign n43451 = n43449 & n43450 ;
  assign n43452 = n43448 | n43451 ;
  assign n43453 = ~n7103 & n43452 ;
  assign n43454 = x745 & n43286 ;
  assign n43455 = x723 & x1135 ;
  assign n43456 = x852 | x1136 ;
  assign n43457 = ~n43455 & n43456 ;
  assign n43458 = n43290 & n43457 ;
  assign n43459 = ~n43454 & n43458 ;
  assign n43460 = x1136 & ~n43275 ;
  assign n43461 = ( x695 & x1134 ) | ( x695 & x1135 ) | ( x1134 & x1135 ) ;
  assign n43462 = ( x612 & ~x1134 ) | ( x612 & x1135 ) | ( ~x1134 & x1135 ) ;
  assign n43463 = ~n43461 & n43462 ;
  assign n43464 = n43460 & n43463 ;
  assign n43465 = n43459 | n43464 ;
  assign n43466 = n7103 & n43465 ;
  assign n43467 = n43453 | n43466 ;
  assign n43468 = x447 & n43253 ;
  assign n43469 = x333 & x591 ;
  assign n43470 = ~x592 & n43469 ;
  assign n43471 = n43468 | n43470 ;
  assign n43472 = ~x590 & n43471 ;
  assign n43473 = x327 & n43260 ;
  assign n43474 = x588 | n43473 ;
  assign n43475 = n43472 | n43474 ;
  assign n43476 = x453 & ~n43265 ;
  assign n43477 = x588 & ~n43476 ;
  assign n43478 = n43264 | n43477 ;
  assign n43479 = n43475 & ~n43478 ;
  assign n43480 = ( x199 & x261 ) | ( x199 & n43264 ) | ( x261 & n43264 ) ;
  assign n43481 = ( ~x199 & x1040 ) | ( ~x199 & n43264 ) | ( x1040 & n43264 ) ;
  assign n43482 = n43480 & n43481 ;
  assign n43483 = n43479 | n43482 ;
  assign n43484 = ~n7103 & n43483 ;
  assign n43485 = x741 & n43286 ;
  assign n43486 = x724 & x1135 ;
  assign n43487 = x865 | x1136 ;
  assign n43488 = ~n43486 & n43487 ;
  assign n43489 = n43290 & n43488 ;
  assign n43490 = ~n43485 & n43489 ;
  assign n43491 = ( x646 & x1134 ) | ( x646 & x1135 ) | ( x1134 & x1135 ) ;
  assign n43492 = ( x611 & ~x1134 ) | ( x611 & x1135 ) | ( ~x1134 & x1135 ) ;
  assign n43493 = ~n43491 & n43492 ;
  assign n43494 = n43460 & n43493 ;
  assign n43495 = n43490 | n43494 ;
  assign n43496 = n7103 & n43495 ;
  assign n43497 = n43484 | n43496 ;
  assign n43498 = ( x616 & x1135 ) | ( x616 & x1136 ) | ( x1135 & x1136 ) ;
  assign n43499 = ( x661 & ~x1135 ) | ( x661 & x1136 ) | ( ~x1135 & x1136 ) ;
  assign n43500 = n43498 & n43499 ;
  assign n43501 = ( ~x781 & x1135 ) | ( ~x781 & x1136 ) | ( x1135 & x1136 ) ;
  assign n43502 = ( x808 & x1135 ) | ( x808 & ~x1136 ) | ( x1135 & ~x1136 ) ;
  assign n43503 = ~n43501 & n43502 ;
  assign n43504 = n43500 | n43503 ;
  assign n43505 = ~n43276 & n43504 ;
  assign n43506 = ~x758 & n43286 ;
  assign n43507 = ~x736 & x1135 ;
  assign n43508 = x850 | x1136 ;
  assign n43509 = ~n43507 & n43508 ;
  assign n43510 = n43290 & n43509 ;
  assign n43511 = ~n43506 & n43510 ;
  assign n43512 = n43505 | n43511 ;
  assign n43513 = n7103 & n43512 ;
  assign n43514 = x320 & n43260 ;
  assign n43515 = x397 & n10558 ;
  assign n43516 = n43302 | n43515 ;
  assign n43517 = x372 & n43253 ;
  assign n43518 = ( ~x592 & n43516 ) | ( ~x592 & n43517 ) | ( n43516 & n43517 ) ;
  assign n43519 = n43514 | n43518 ;
  assign n43520 = x422 & ~n43265 ;
  assign n43521 = x588 & ~n43520 ;
  assign n43522 = n43264 | n43521 ;
  assign n43523 = n43519 & ~n43522 ;
  assign n43524 = ( x199 & x290 ) | ( x199 & n43264 ) | ( x290 & n43264 ) ;
  assign n43525 = ( ~x199 & x1048 ) | ( ~x199 & n43264 ) | ( x1048 & n43264 ) ;
  assign n43526 = n43524 & n43525 ;
  assign n43527 = n43523 | n43526 ;
  assign n43528 = ~n7103 & n43527 ;
  assign n43529 = n43513 | n43528 ;
  assign n43530 = ( x617 & x1135 ) | ( x617 & x1136 ) | ( x1135 & x1136 ) ;
  assign n43531 = ( x637 & ~x1135 ) | ( x637 & x1136 ) | ( ~x1135 & x1136 ) ;
  assign n43532 = n43530 & n43531 ;
  assign n43533 = ( ~x788 & x1135 ) | ( ~x788 & x1136 ) | ( x1135 & x1136 ) ;
  assign n43534 = ( x814 & ~x1135 ) | ( x814 & x1136 ) | ( ~x1135 & x1136 ) ;
  assign n43535 = n43533 | n43534 ;
  assign n43536 = ~n43532 & n43535 ;
  assign n43537 = n43276 | n43536 ;
  assign n43538 = ~x749 & n43286 ;
  assign n43539 = ~x706 & x1135 ;
  assign n43540 = x866 | x1136 ;
  assign n43541 = ~n43539 & n43540 ;
  assign n43542 = n43290 & n43541 ;
  assign n43543 = ~n43538 & n43542 ;
  assign n43544 = n43537 & ~n43543 ;
  assign n43545 = n7103 & ~n43544 ;
  assign n43546 = x452 & n43260 ;
  assign n43547 = x411 & n10558 ;
  assign n43548 = n43302 | n43547 ;
  assign n43549 = x387 & n43253 ;
  assign n43550 = ( ~x592 & n43548 ) | ( ~x592 & n43549 ) | ( n43548 & n43549 ) ;
  assign n43551 = n43546 | n43550 ;
  assign n43552 = x435 & ~n43265 ;
  assign n43553 = x588 & ~n43552 ;
  assign n43554 = n43264 | n43553 ;
  assign n43555 = n43551 & ~n43554 ;
  assign n43556 = ( x199 & x295 ) | ( x199 & n43264 ) | ( x295 & n43264 ) ;
  assign n43557 = ( ~x199 & x1053 ) | ( ~x199 & n43264 ) | ( x1053 & n43264 ) ;
  assign n43558 = n43556 & n43557 ;
  assign n43559 = n43555 | n43558 ;
  assign n43560 = ~n7103 & n43559 ;
  assign n43561 = n43545 | n43560 ;
  assign n43562 = x336 & n43253 ;
  assign n43563 = x463 & x591 ;
  assign n43564 = ~x592 & n43563 ;
  assign n43565 = n43562 | n43564 ;
  assign n43566 = ~x590 & n43565 ;
  assign n43567 = x362 & n43260 ;
  assign n43568 = x588 | n43567 ;
  assign n43569 = n43566 | n43568 ;
  assign n43570 = x437 & ~n43265 ;
  assign n43571 = x588 & ~n43570 ;
  assign n43572 = n43264 | n43571 ;
  assign n43573 = n43569 & ~n43572 ;
  assign n43574 = ( x199 & x256 ) | ( x199 & n43264 ) | ( x256 & n43264 ) ;
  assign n43575 = ( ~x199 & x1070 ) | ( ~x199 & n43264 ) | ( x1070 & n43264 ) ;
  assign n43576 = n43574 & n43575 ;
  assign n43577 = n43573 | n43576 ;
  assign n43578 = ~n7103 & n43577 ;
  assign n43579 = ( ~x622 & x1135 ) | ( ~x622 & x1136 ) | ( x1135 & x1136 ) ;
  assign n43580 = ( x639 & x1135 ) | ( x639 & ~x1136 ) | ( x1135 & ~x1136 ) ;
  assign n43581 = n43579 & ~n43580 ;
  assign n43582 = ( x783 & x1135 ) | ( x783 & x1136 ) | ( x1135 & x1136 ) ;
  assign n43583 = ( x804 & ~x1135 ) | ( x804 & x1136 ) | ( ~x1135 & x1136 ) ;
  assign n43584 = n43582 | n43583 ;
  assign n43585 = ~n43581 & n43584 ;
  assign n43586 = x1134 | n43585 ;
  assign n43587 = x859 & ~n43324 ;
  assign n43588 = x1134 & ~n43587 ;
  assign n43589 = ( x743 & x1135 ) | ( x743 & x1136 ) | ( x1135 & x1136 ) ;
  assign n43590 = ( x735 & ~x1135 ) | ( x735 & x1136 ) | ( ~x1135 & x1136 ) ;
  assign n43591 = n43589 & n43590 ;
  assign n43592 = n43588 & ~n43591 ;
  assign n43593 = n43331 & ~n43592 ;
  assign n43594 = n43586 & n43593 ;
  assign n43595 = n43578 | n43594 ;
  assign n43596 = x876 & ~n43324 ;
  assign n43597 = ( x748 & x1135 ) | ( x748 & x1136 ) | ( x1135 & x1136 ) ;
  assign n43598 = ( x730 & ~x1135 ) | ( x730 & x1136 ) | ( ~x1135 & x1136 ) ;
  assign n43599 = n43597 & n43598 ;
  assign n43600 = n43596 | n43599 ;
  assign n43601 = n43289 & n43600 ;
  assign n43602 = ~x623 & n43286 ;
  assign n43603 = n43276 | n43602 ;
  assign n43604 = x789 & n43288 ;
  assign n43605 = x803 | x1135 ;
  assign n43606 = ~n43604 & n43605 ;
  assign n43607 = x1135 & x1136 ;
  assign n43608 = ~x710 & n43607 ;
  assign n43609 = ( ~x1136 & n43606 ) | ( ~x1136 & n43608 ) | ( n43606 & n43608 ) ;
  assign n43610 = n43603 | n43609 ;
  assign n43611 = ~n43601 & n43610 ;
  assign n43612 = n7103 & ~n43611 ;
  assign n43613 = x455 & n43260 ;
  assign n43614 = x412 & n10558 ;
  assign n43615 = n43302 | n43614 ;
  assign n43616 = x388 & n43253 ;
  assign n43617 = ( ~x592 & n43615 ) | ( ~x592 & n43616 ) | ( n43615 & n43616 ) ;
  assign n43618 = n43613 | n43617 ;
  assign n43619 = x436 & ~n43265 ;
  assign n43620 = x588 & ~n43619 ;
  assign n43621 = n43264 | n43620 ;
  assign n43622 = n43618 & ~n43621 ;
  assign n43623 = ( x199 & x296 ) | ( x199 & n43264 ) | ( x296 & n43264 ) ;
  assign n43624 = ( ~x199 & x1037 ) | ( ~x199 & n43264 ) | ( x1037 & n43264 ) ;
  assign n43625 = n43623 & n43624 ;
  assign n43626 = n43622 | n43625 ;
  assign n43627 = ~n7103 & n43626 ;
  assign n43628 = n43612 | n43627 ;
  assign n43629 = ( x606 & x1135 ) | ( x606 & x1136 ) | ( x1135 & x1136 ) ;
  assign n43630 = ( x643 & ~x1135 ) | ( x643 & x1136 ) | ( ~x1135 & x1136 ) ;
  assign n43631 = n43629 & n43630 ;
  assign n43632 = ( ~x787 & x1135 ) | ( ~x787 & x1136 ) | ( x1135 & x1136 ) ;
  assign n43633 = ( x812 & ~x1135 ) | ( x812 & x1136 ) | ( ~x1135 & x1136 ) ;
  assign n43634 = n43632 | n43633 ;
  assign n43635 = ~n43631 & n43634 ;
  assign n43636 = n43276 | n43635 ;
  assign n43637 = ~x746 & n43286 ;
  assign n43638 = ~x729 & x1135 ;
  assign n43639 = x881 | x1136 ;
  assign n43640 = ~n43638 & n43639 ;
  assign n43641 = n43290 & n43640 ;
  assign n43642 = ~n43637 & n43641 ;
  assign n43643 = n43636 & ~n43642 ;
  assign n43644 = n7103 & ~n43643 ;
  assign n43645 = x361 & n43260 ;
  assign n43646 = x410 & n10558 ;
  assign n43647 = n43302 | n43646 ;
  assign n43648 = x386 & n43253 ;
  assign n43649 = ( ~x592 & n43647 ) | ( ~x592 & n43648 ) | ( n43647 & n43648 ) ;
  assign n43650 = n43645 | n43649 ;
  assign n43651 = x434 & ~n43265 ;
  assign n43652 = x588 & ~n43651 ;
  assign n43653 = n43264 | n43652 ;
  assign n43654 = n43650 & ~n43653 ;
  assign n43655 = ( x199 & x293 ) | ( x199 & n43264 ) | ( x293 & n43264 ) ;
  assign n43656 = ( ~x199 & x1059 ) | ( ~x199 & n43264 ) | ( x1059 & n43264 ) ;
  assign n43657 = n43655 & n43656 ;
  assign n43658 = n43654 | n43657 ;
  assign n43659 = ~n7103 & n43658 ;
  assign n43660 = n43644 | n43659 ;
  assign n43661 = x366 & n43253 ;
  assign n43662 = x335 & x591 ;
  assign n43663 = ~x592 & n43662 ;
  assign n43664 = n43661 | n43663 ;
  assign n43665 = ~x590 & n43664 ;
  assign n43666 = x344 & n43260 ;
  assign n43667 = x588 | n43666 ;
  assign n43668 = n43665 | n43667 ;
  assign n43669 = x416 & ~n43265 ;
  assign n43670 = x588 & ~n43669 ;
  assign n43671 = n43264 | n43670 ;
  assign n43672 = n43668 & ~n43671 ;
  assign n43673 = ( x199 & x259 ) | ( x199 & n43264 ) | ( x259 & n43264 ) ;
  assign n43674 = ( ~x199 & x1069 ) | ( ~x199 & n43264 ) | ( x1069 & n43264 ) ;
  assign n43675 = n43673 & n43674 ;
  assign n43676 = n43672 | n43675 ;
  assign n43677 = ~n7103 & n43676 ;
  assign n43678 = x742 & n43286 ;
  assign n43679 = x704 & x1135 ;
  assign n43680 = x870 | x1136 ;
  assign n43681 = ~n43679 & n43680 ;
  assign n43682 = n43290 & n43681 ;
  assign n43683 = ~n43678 & n43682 ;
  assign n43684 = ( x635 & x1134 ) | ( x635 & x1135 ) | ( x1134 & x1135 ) ;
  assign n43685 = ( x620 & ~x1134 ) | ( x620 & x1135 ) | ( ~x1134 & x1135 ) ;
  assign n43686 = ~n43684 & n43685 ;
  assign n43687 = n43460 & n43686 ;
  assign n43688 = n43683 | n43687 ;
  assign n43689 = n7103 & n43688 ;
  assign n43690 = n43677 | n43689 ;
  assign n43691 = x368 & n43253 ;
  assign n43692 = x393 & x591 ;
  assign n43693 = ~x592 & n43692 ;
  assign n43694 = n43691 | n43693 ;
  assign n43695 = ~x590 & n43694 ;
  assign n43696 = x346 & n43260 ;
  assign n43697 = x588 | n43696 ;
  assign n43698 = n43695 | n43697 ;
  assign n43699 = x418 & ~n43265 ;
  assign n43700 = x588 & ~n43699 ;
  assign n43701 = n43264 | n43700 ;
  assign n43702 = n43698 & ~n43701 ;
  assign n43703 = ( x199 & x260 ) | ( x199 & n43264 ) | ( x260 & n43264 ) ;
  assign n43704 = ( ~x199 & x1067 ) | ( ~x199 & n43264 ) | ( x1067 & n43264 ) ;
  assign n43705 = n43703 & n43704 ;
  assign n43706 = n43702 | n43705 ;
  assign n43707 = ~n7103 & n43706 ;
  assign n43708 = x760 & n43286 ;
  assign n43709 = x688 & x1135 ;
  assign n43710 = x856 | x1136 ;
  assign n43711 = ~n43709 & n43710 ;
  assign n43712 = n43290 & n43711 ;
  assign n43713 = ~n43708 & n43712 ;
  assign n43714 = ( x632 & x1134 ) | ( x632 & x1135 ) | ( x1134 & x1135 ) ;
  assign n43715 = ( x613 & ~x1134 ) | ( x613 & x1135 ) | ( ~x1134 & x1135 ) ;
  assign n43716 = ~n43714 & n43715 ;
  assign n43717 = n43460 & n43716 ;
  assign n43718 = n43713 | n43717 ;
  assign n43719 = n7103 & n43718 ;
  assign n43720 = n43707 | n43719 ;
  assign n43721 = x389 & n43253 ;
  assign n43722 = x413 & x591 ;
  assign n43723 = ~x592 & n43722 ;
  assign n43724 = n43721 | n43723 ;
  assign n43725 = ~x590 & n43724 ;
  assign n43726 = x450 & n43260 ;
  assign n43727 = x588 | n43726 ;
  assign n43728 = n43725 | n43727 ;
  assign n43729 = x438 & ~n43265 ;
  assign n43730 = x588 & ~n43729 ;
  assign n43731 = n43264 | n43730 ;
  assign n43732 = n43728 & ~n43731 ;
  assign n43733 = ( x199 & x255 ) | ( x199 & n43264 ) | ( x255 & n43264 ) ;
  assign n43734 = ( ~x199 & x1036 ) | ( ~x199 & n43264 ) | ( x1036 & n43264 ) ;
  assign n43735 = n43733 & n43734 ;
  assign n43736 = n43732 | n43735 ;
  assign n43737 = ~n7103 & n43736 ;
  assign n43738 = ( x665 & x1135 ) | ( x665 & ~x1136 ) | ( x1135 & ~x1136 ) ;
  assign n43739 = ( x791 & x1135 ) | ( x791 & x1136 ) | ( x1135 & x1136 ) ;
  assign n43740 = n43738 & n43739 ;
  assign n43741 = ( ~x621 & x1135 ) | ( ~x621 & x1136 ) | ( x1135 & x1136 ) ;
  assign n43742 = ( x810 & ~x1135 ) | ( x810 & x1136 ) | ( ~x1135 & x1136 ) ;
  assign n43743 = ~n43741 & n43742 ;
  assign n43744 = n43740 | n43743 ;
  assign n43745 = ~n43276 & n43744 ;
  assign n43746 = ~x739 & n43286 ;
  assign n43747 = x874 | x1136 ;
  assign n43748 = ~x690 & x1135 ;
  assign n43749 = n43747 & ~n43748 ;
  assign n43750 = n43290 & n43749 ;
  assign n43751 = ~n43746 & n43750 ;
  assign n43752 = n43745 | n43751 ;
  assign n43753 = n7103 & n43752 ;
  assign n43754 = n43737 | n43753 ;
  assign n43755 = ( x962 & ~x1100 ) | ( x962 & n43129 ) | ( ~x1100 & n43129 ) ;
  assign n43756 = ( x680 & ~x962 ) | ( x680 & n43129 ) | ( ~x962 & n43129 ) ;
  assign n43757 = ~n43755 & n43756 ;
  assign n43758 = ( x962 & ~x1103 ) | ( x962 & n43129 ) | ( ~x1103 & n43129 ) ;
  assign n43759 = ( x681 & ~x962 ) | ( x681 & n43129 ) | ( ~x962 & n43129 ) ;
  assign n43760 = ~n43758 & n43759 ;
  assign n43761 = x367 & n43253 ;
  assign n43762 = x392 & x591 ;
  assign n43763 = ~x592 & n43762 ;
  assign n43764 = n43761 | n43763 ;
  assign n43765 = ~x590 & n43764 ;
  assign n43766 = x345 & n43260 ;
  assign n43767 = x588 | n43766 ;
  assign n43768 = n43765 | n43767 ;
  assign n43769 = x417 & ~n43265 ;
  assign n43770 = x588 & ~n43769 ;
  assign n43771 = n43264 | n43770 ;
  assign n43772 = n43768 & ~n43771 ;
  assign n43773 = ( x199 & x251 ) | ( x199 & n43264 ) | ( x251 & n43264 ) ;
  assign n43774 = ( ~x199 & x1039 ) | ( ~x199 & n43264 ) | ( x1039 & n43264 ) ;
  assign n43775 = n43773 & n43774 ;
  assign n43776 = n43772 | n43775 ;
  assign n43777 = ~n7103 & n43776 ;
  assign n43778 = x757 & n43286 ;
  assign n43779 = x686 & x1135 ;
  assign n43780 = x848 | x1136 ;
  assign n43781 = ~n43779 & n43780 ;
  assign n43782 = n43290 & n43781 ;
  assign n43783 = ~n43778 & n43782 ;
  assign n43784 = ( x631 & x1134 ) | ( x631 & x1135 ) | ( x1134 & x1135 ) ;
  assign n43785 = ( x610 & ~x1134 ) | ( x610 & x1135 ) | ( ~x1134 & x1135 ) ;
  assign n43786 = ~n43784 & n43785 ;
  assign n43787 = n43460 & n43786 ;
  assign n43788 = n43783 | n43787 ;
  assign n43789 = n7103 & n43788 ;
  assign n43790 = n43777 | n43789 ;
  assign n43791 = x953 & n43128 ;
  assign n43792 = ( x962 & ~x1130 ) | ( x962 & n43791 ) | ( ~x1130 & n43791 ) ;
  assign n43793 = ( x684 & x962 ) | ( x684 & ~n43791 ) | ( x962 & ~n43791 ) ;
  assign n43794 = n43792 | n43793 ;
  assign n43795 = x590 & ~x592 ;
  assign n43796 = x357 & n43795 ;
  assign n43797 = x382 & n43301 ;
  assign n43798 = n43796 | n43797 ;
  assign n43799 = ~x591 & n43798 ;
  assign n43800 = x406 & ~x592 ;
  assign n43801 = n10558 & n43800 ;
  assign n43802 = n43799 | n43801 ;
  assign n43803 = ~x588 & n43802 ;
  assign n43804 = x588 & ~x590 ;
  assign n43805 = x430 & ~n43259 ;
  assign n43806 = n43804 & n43805 ;
  assign n43807 = n43803 | n43806 ;
  assign n43808 = ~n43264 & n43807 ;
  assign n43809 = x199 & ~x1076 ;
  assign n43810 = n43264 & ~n43809 ;
  assign n43811 = n39407 & n43810 ;
  assign n43812 = n43808 | n43811 ;
  assign n43813 = ~n7103 & n43812 ;
  assign n43814 = x860 & ~n43324 ;
  assign n43815 = ( ~x744 & x1135 ) | ( ~x744 & x1136 ) | ( x1135 & x1136 ) ;
  assign n43816 = ( x728 & x1135 ) | ( x728 & ~x1136 ) | ( x1135 & ~x1136 ) ;
  assign n43817 = n43815 & ~n43816 ;
  assign n43818 = n43814 | n43817 ;
  assign n43819 = n43289 & n43818 ;
  assign n43820 = x1136 & n43275 ;
  assign n43821 = x1134 | n43820 ;
  assign n43822 = x813 & ~n43275 ;
  assign n43823 = ~n43324 & n43822 ;
  assign n43824 = ( x652 & x1135 ) | ( x652 & x1136 ) | ( x1135 & x1136 ) ;
  assign n43825 = ( x657 & x1135 ) | ( x657 & ~x1136 ) | ( x1135 & ~x1136 ) ;
  assign n43826 = n43824 & ~n43825 ;
  assign n43827 = n43823 | n43826 ;
  assign n43828 = ~n43821 & n43827 ;
  assign n43829 = n43819 | n43828 ;
  assign n43830 = n7103 & n43829 ;
  assign n43831 = n43813 | n43830 ;
  assign n43832 = ( x962 & ~x1113 ) | ( x962 & n43791 ) | ( ~x1113 & n43791 ) ;
  assign n43833 = ( x686 & x962 ) | ( x686 & ~n43791 ) | ( x962 & ~n43791 ) ;
  assign n43834 = n43832 | n43833 ;
  assign n43835 = ( x962 & ~x1127 ) | ( x962 & n43791 ) | ( ~x1127 & n43791 ) ;
  assign n43836 = ( x687 & ~x962 ) | ( x687 & n43791 ) | ( ~x962 & n43791 ) ;
  assign n43837 = ~n43835 & n43836 ;
  assign n43838 = ( x962 & ~x1115 ) | ( x962 & n43791 ) | ( ~x1115 & n43791 ) ;
  assign n43839 = ( x688 & x962 ) | ( x688 & ~n43791 ) | ( x962 & ~n43791 ) ;
  assign n43840 = n43838 | n43839 ;
  assign n43841 = x351 & n43795 ;
  assign n43842 = x376 & n43301 ;
  assign n43843 = n43841 | n43842 ;
  assign n43844 = ~x591 & n43843 ;
  assign n43845 = x401 & ~x592 ;
  assign n43846 = n10558 & n43845 ;
  assign n43847 = n43844 | n43846 ;
  assign n43848 = ~x588 & n43847 ;
  assign n43849 = x426 & ~n43259 ;
  assign n43850 = n43804 & n43849 ;
  assign n43851 = n43848 | n43850 ;
  assign n43852 = ~n43264 & n43851 ;
  assign n43853 = ( x199 & n39377 ) | ( x199 & n43264 ) | ( n39377 & n43264 ) ;
  assign n43854 = ( ~x199 & x1079 ) | ( ~x199 & n43264 ) | ( x1079 & n43264 ) ;
  assign n43855 = n43853 & n43854 ;
  assign n43856 = n43852 | n43855 ;
  assign n43857 = ~n7103 & n43856 ;
  assign n43858 = x798 & ~n43324 ;
  assign n43859 = ( x658 & x1135 ) | ( x658 & x1136 ) | ( x1135 & x1136 ) ;
  assign n43860 = ( x655 & x1135 ) | ( x655 & ~x1136 ) | ( x1135 & ~x1136 ) ;
  assign n43861 = n43859 & ~n43860 ;
  assign n43862 = n43858 | n43861 ;
  assign n43863 = ~n43276 & n43862 ;
  assign n43864 = x752 & n43286 ;
  assign n43865 = ~x703 & x1135 ;
  assign n43866 = x843 | x1136 ;
  assign n43867 = ~n43865 & n43866 ;
  assign n43868 = n43290 & n43867 ;
  assign n43869 = ~n43864 & n43868 ;
  assign n43870 = n43863 | n43869 ;
  assign n43871 = n7103 & n43870 ;
  assign n43872 = n43857 | n43871 ;
  assign n43873 = ( x962 & ~x1108 ) | ( x962 & n43791 ) | ( ~x1108 & n43791 ) ;
  assign n43874 = ( x690 & ~x962 ) | ( x690 & n43791 ) | ( ~x962 & n43791 ) ;
  assign n43875 = ~n43873 & n43874 ;
  assign n43876 = ( x962 & ~x1107 ) | ( x962 & n43791 ) | ( ~x1107 & n43791 ) ;
  assign n43877 = ( x691 & ~x962 ) | ( x691 & n43791 ) | ( ~x962 & n43791 ) ;
  assign n43878 = ~n43876 & n43877 ;
  assign n43879 = x352 & n43795 ;
  assign n43880 = x317 & n43301 ;
  assign n43881 = n43879 | n43880 ;
  assign n43882 = ~x591 & n43881 ;
  assign n43883 = x402 & ~x592 ;
  assign n43884 = n10558 & n43883 ;
  assign n43885 = n43882 | n43884 ;
  assign n43886 = ~x588 & n43885 ;
  assign n43887 = x427 & ~n43259 ;
  assign n43888 = n43804 & n43887 ;
  assign n43889 = n43886 | n43888 ;
  assign n43890 = ~n43264 & n43889 ;
  assign n43891 = ( x199 & n39389 ) | ( x199 & n43264 ) | ( n39389 & n43264 ) ;
  assign n43892 = ( ~x199 & x1078 ) | ( ~x199 & n43264 ) | ( x1078 & n43264 ) ;
  assign n43893 = n43891 & n43892 ;
  assign n43894 = n43890 | n43893 ;
  assign n43895 = ~n7103 & n43894 ;
  assign n43896 = x801 & ~n43324 ;
  assign n43897 = x1134 | n43896 ;
  assign n43898 = ( x656 & x1135 ) | ( x656 & x1136 ) | ( x1135 & x1136 ) ;
  assign n43899 = ( x649 & x1135 ) | ( x649 & ~x1136 ) | ( x1135 & ~x1136 ) ;
  assign n43900 = n43898 & ~n43899 ;
  assign n43901 = n43897 | n43900 ;
  assign n43902 = x844 & ~n43324 ;
  assign n43903 = x1134 & ~n43902 ;
  assign n43904 = ( ~x770 & x1135 ) | ( ~x770 & x1136 ) | ( x1135 & x1136 ) ;
  assign n43905 = ( x726 & ~x1135 ) | ( x726 & x1136 ) | ( ~x1135 & x1136 ) ;
  assign n43906 = n43904 & n43905 ;
  assign n43907 = n43903 & ~n43906 ;
  assign n43908 = n43331 & ~n43907 ;
  assign n43909 = n43901 & n43908 ;
  assign n43910 = n43895 | n43909 ;
  assign n43911 = ( x962 & ~x1129 ) | ( x962 & n43129 ) | ( ~x1129 & n43129 ) ;
  assign n43912 = ( x693 & x962 ) | ( x693 & ~n43129 ) | ( x962 & ~n43129 ) ;
  assign n43913 = n43911 | n43912 ;
  assign n43914 = ( x962 & ~x1128 ) | ( x962 & n43791 ) | ( ~x1128 & n43791 ) ;
  assign n43915 = ( x694 & x962 ) | ( x694 & ~n43791 ) | ( x962 & ~n43791 ) ;
  assign n43916 = n43914 | n43915 ;
  assign n43917 = ( x962 & ~x1111 ) | ( x962 & n43129 ) | ( ~x1111 & n43129 ) ;
  assign n43918 = ( x695 & x962 ) | ( x695 & ~n43129 ) | ( x962 & ~n43129 ) ;
  assign n43919 = n43917 | n43918 ;
  assign n43920 = ( x962 & ~x1100 ) | ( x962 & n43791 ) | ( ~x1100 & n43791 ) ;
  assign n43921 = ( x696 & ~x962 ) | ( x696 & n43791 ) | ( ~x962 & n43791 ) ;
  assign n43922 = ~n43920 & n43921 ;
  assign n43923 = ( x962 & ~x1129 ) | ( x962 & n43791 ) | ( ~x1129 & n43791 ) ;
  assign n43924 = ( x697 & x962 ) | ( x697 & ~n43791 ) | ( x962 & ~n43791 ) ;
  assign n43925 = n43923 | n43924 ;
  assign n43926 = ( x962 & ~x1116 ) | ( x962 & n43791 ) | ( ~x1116 & n43791 ) ;
  assign n43927 = ( x698 & x962 ) | ( x698 & ~n43791 ) | ( x962 & ~n43791 ) ;
  assign n43928 = n43926 | n43927 ;
  assign n43929 = ( x962 & ~x1103 ) | ( x962 & n43791 ) | ( ~x1103 & n43791 ) ;
  assign n43930 = ( x699 & ~x962 ) | ( x699 & n43791 ) | ( ~x962 & n43791 ) ;
  assign n43931 = ~n43929 & n43930 ;
  assign n43932 = ( x962 & ~x1110 ) | ( x962 & n43791 ) | ( ~x1110 & n43791 ) ;
  assign n43933 = ( x700 & ~x962 ) | ( x700 & n43791 ) | ( ~x962 & n43791 ) ;
  assign n43934 = ~n43932 & n43933 ;
  assign n43935 = ( x962 & ~x1123 ) | ( x962 & n43791 ) | ( ~x1123 & n43791 ) ;
  assign n43936 = ( x701 & x962 ) | ( x701 & ~n43791 ) | ( x962 & ~n43791 ) ;
  assign n43937 = n43935 | n43936 ;
  assign n43938 = ( x962 & ~x1117 ) | ( x962 & n43791 ) | ( ~x1117 & n43791 ) ;
  assign n43939 = ( x702 & x962 ) | ( x702 & ~n43791 ) | ( x962 & ~n43791 ) ;
  assign n43940 = n43938 | n43939 ;
  assign n43941 = ( x962 & ~x1124 ) | ( x962 & n43791 ) | ( ~x1124 & n43791 ) ;
  assign n43942 = ( x703 & ~x962 ) | ( x703 & n43791 ) | ( ~x962 & n43791 ) ;
  assign n43943 = ~n43941 & n43942 ;
  assign n43944 = ( x962 & ~x1112 ) | ( x962 & n43791 ) | ( ~x1112 & n43791 ) ;
  assign n43945 = ( x704 & x962 ) | ( x704 & ~n43791 ) | ( x962 & ~n43791 ) ;
  assign n43946 = n43944 | n43945 ;
  assign n43947 = ( x962 & ~x1125 ) | ( x962 & n43791 ) | ( ~x1125 & n43791 ) ;
  assign n43948 = ( x705 & ~x962 ) | ( x705 & n43791 ) | ( ~x962 & n43791 ) ;
  assign n43949 = ~n43947 & n43948 ;
  assign n43950 = ( x962 & ~x1105 ) | ( x962 & n43791 ) | ( ~x1105 & n43791 ) ;
  assign n43951 = ( x706 & ~x962 ) | ( x706 & n43791 ) | ( ~x962 & n43791 ) ;
  assign n43952 = ~n43950 & n43951 ;
  assign n43953 = x370 & n43253 ;
  assign n43954 = x395 & x591 ;
  assign n43955 = ~x592 & n43954 ;
  assign n43956 = n43953 | n43955 ;
  assign n43957 = ~x590 & n43956 ;
  assign n43958 = x347 & n43260 ;
  assign n43959 = n43957 | n43958 ;
  assign n43960 = x588 | n43264 ;
  assign n43961 = n43959 & ~n43960 ;
  assign n43962 = x199 & ~x1055 ;
  assign n43963 = n43264 & ~n43962 ;
  assign n43964 = ( x199 & x200 ) | ( x199 & x1048 ) | ( x200 & x1048 ) ;
  assign n43965 = ( x199 & ~x200 ) | ( x199 & x304 ) | ( ~x200 & x304 ) ;
  assign n43966 = n43964 | n43965 ;
  assign n43967 = n43963 & n43966 ;
  assign n43968 = n43264 | n43265 ;
  assign n43969 = x420 & x588 ;
  assign n43970 = ~n43968 & n43969 ;
  assign n43971 = n43967 | n43970 ;
  assign n43972 = n43961 | n43971 ;
  assign n43973 = ~n7103 & n43972 ;
  assign n43974 = ( ~x627 & x1134 ) | ( ~x627 & x1135 ) | ( x1134 & x1135 ) ;
  assign n43975 = ( x618 & ~x1134 ) | ( x618 & x1135 ) | ( ~x1134 & x1135 ) ;
  assign n43976 = ~n43974 & n43975 ;
  assign n43977 = n43460 & n43976 ;
  assign n43978 = x753 & n43286 ;
  assign n43979 = x702 & x1135 ;
  assign n43980 = x847 | x1136 ;
  assign n43981 = ~n43979 & n43980 ;
  assign n43982 = n43290 & n43981 ;
  assign n43983 = ~n43978 & n43982 ;
  assign n43984 = n43977 | n43983 ;
  assign n43985 = n7103 & n43984 ;
  assign n43986 = n43973 | n43985 ;
  assign n43987 = n43253 & ~n43264 ;
  assign n43988 = x442 & n43987 ;
  assign n43989 = x592 | n43264 ;
  assign n43990 = x328 & x591 ;
  assign n43991 = ~n43989 & n43990 ;
  assign n43992 = n43988 | n43991 ;
  assign n43993 = ~x590 & n43992 ;
  assign n43994 = x321 & ~n43264 ;
  assign n43995 = n43260 & n43994 ;
  assign n43996 = n43993 | n43995 ;
  assign n43997 = ~x588 & n43996 ;
  assign n43998 = x199 & ~x1058 ;
  assign n43999 = n43264 & ~n43998 ;
  assign n44000 = ( x199 & x200 ) | ( x199 & x1084 ) | ( x200 & x1084 ) ;
  assign n44001 = ( x199 & ~x200 ) | ( x199 & x305 ) | ( ~x200 & x305 ) ;
  assign n44002 = n44000 | n44001 ;
  assign n44003 = n43999 & n44002 ;
  assign n44004 = n43259 | n43264 ;
  assign n44005 = x459 & n43804 ;
  assign n44006 = ~n44004 & n44005 ;
  assign n44007 = n7103 | n44006 ;
  assign n44008 = n44003 | n44007 ;
  assign n44009 = n43997 | n44008 ;
  assign n44010 = x754 & n43286 ;
  assign n44011 = n43275 | n43288 ;
  assign n44012 = x857 | x1136 ;
  assign n44013 = x709 & x1135 ;
  assign n44014 = x1134 & ~n44013 ;
  assign n44015 = n44012 & n44014 ;
  assign n44016 = ~n44011 & n44015 ;
  assign n44017 = ~n44010 & n44016 ;
  assign n44018 = ( ~x660 & x1134 ) | ( ~x660 & x1135 ) | ( x1134 & x1135 ) ;
  assign n44019 = ( x609 & ~x1134 ) | ( x609 & x1135 ) | ( ~x1134 & x1135 ) ;
  assign n44020 = ~n44018 & n44019 ;
  assign n44021 = n43460 & n44020 ;
  assign n44022 = n7103 & ~n44021 ;
  assign n44023 = ~n44017 & n44022 ;
  assign n44024 = n44009 & ~n44023 ;
  assign n44025 = ( x962 & ~x1118 ) | ( x962 & n43791 ) | ( ~x1118 & n43791 ) ;
  assign n44026 = ( x709 & x962 ) | ( x709 & ~n43791 ) | ( x962 & ~n43791 ) ;
  assign n44027 = n44025 | n44026 ;
  assign n44028 = ( x962 & ~x1106 ) | ( x962 & n43129 ) | ( ~x1106 & n43129 ) ;
  assign n44029 = ( x710 & ~x962 ) | ( x710 & n43129 ) | ( ~x962 & n43129 ) ;
  assign n44030 = ~n44028 & n44029 ;
  assign n44031 = x373 & n43253 ;
  assign n44032 = x398 & x591 ;
  assign n44033 = ~x592 & n44032 ;
  assign n44034 = n44031 | n44033 ;
  assign n44035 = ~x590 & n44034 ;
  assign n44036 = x348 & n43260 ;
  assign n44037 = n44035 | n44036 ;
  assign n44038 = ~n43960 & n44037 ;
  assign n44039 = x199 & ~x1087 ;
  assign n44040 = n43264 & ~n44039 ;
  assign n44041 = ( x199 & x200 ) | ( x199 & x1059 ) | ( x200 & x1059 ) ;
  assign n44042 = ( x199 & ~x200 ) | ( x199 & x306 ) | ( ~x200 & x306 ) ;
  assign n44043 = n44041 | n44042 ;
  assign n44044 = n44040 & n44043 ;
  assign n44045 = x423 & x588 ;
  assign n44046 = ~n43968 & n44045 ;
  assign n44047 = n44044 | n44046 ;
  assign n44048 = n44038 | n44047 ;
  assign n44049 = ~n7103 & n44048 ;
  assign n44050 = ( ~x647 & x1134 ) | ( ~x647 & x1135 ) | ( x1134 & x1135 ) ;
  assign n44051 = ( x630 & ~x1134 ) | ( x630 & x1135 ) | ( ~x1134 & x1135 ) ;
  assign n44052 = ~n44050 & n44051 ;
  assign n44053 = n43460 & n44052 ;
  assign n44054 = x755 & n43286 ;
  assign n44055 = x725 & x1135 ;
  assign n44056 = x858 | x1136 ;
  assign n44057 = ~n44055 & n44056 ;
  assign n44058 = n43290 & n44057 ;
  assign n44059 = ~n44054 & n44058 ;
  assign n44060 = n44053 | n44059 ;
  assign n44061 = n7103 & n44060 ;
  assign n44062 = n44049 | n44061 ;
  assign n44063 = x751 & n43286 ;
  assign n44064 = x842 | x1136 ;
  assign n44065 = x701 & x1135 ;
  assign n44066 = x1134 & ~n44065 ;
  assign n44067 = n44064 & n44066 ;
  assign n44068 = ~n44011 & n44067 ;
  assign n44069 = ~n44063 & n44068 ;
  assign n44070 = ( ~x715 & x1134 ) | ( ~x715 & x1135 ) | ( x1134 & x1135 ) ;
  assign n44071 = ( x644 & ~x1134 ) | ( x644 & x1135 ) | ( ~x1134 & x1135 ) ;
  assign n44072 = ~n44070 & n44071 ;
  assign n44073 = n43460 & n44072 ;
  assign n44074 = n44069 | n44073 ;
  assign n44075 = n7103 & n44074 ;
  assign n44076 = x374 & n43253 ;
  assign n44077 = x400 & x591 ;
  assign n44078 = ~x592 & n44077 ;
  assign n44079 = n44076 | n44078 ;
  assign n44080 = ~x590 & n44079 ;
  assign n44081 = x350 & n43260 ;
  assign n44082 = n44080 | n44081 ;
  assign n44083 = ~x588 & n44082 ;
  assign n44084 = x425 & ~n43259 ;
  assign n44085 = n43804 & n44084 ;
  assign n44086 = n43264 | n44085 ;
  assign n44087 = n44083 | n44086 ;
  assign n44088 = x1044 & n9578 ;
  assign n44089 = x298 & ~n8980 ;
  assign n44090 = x199 & x1035 ;
  assign n44091 = n43264 & ~n44090 ;
  assign n44092 = ~n44089 & n44091 ;
  assign n44093 = ~n44088 & n44092 ;
  assign n44094 = n7103 | n44093 ;
  assign n44095 = n44087 & ~n44094 ;
  assign n44096 = n44075 | n44095 ;
  assign n44097 = x371 & n43253 ;
  assign n44098 = x396 & x591 ;
  assign n44099 = ~x592 & n44098 ;
  assign n44100 = n44097 | n44099 ;
  assign n44101 = ~x590 & n44100 ;
  assign n44102 = x322 & n43260 ;
  assign n44103 = n44101 | n44102 ;
  assign n44104 = ~n43960 & n44103 ;
  assign n44105 = x199 & ~x1051 ;
  assign n44106 = n43264 & ~n44105 ;
  assign n44107 = ( x199 & x200 ) | ( x199 & x1072 ) | ( x200 & x1072 ) ;
  assign n44108 = ( x199 & ~x200 ) | ( x199 & x309 ) | ( ~x200 & x309 ) ;
  assign n44109 = n44107 | n44108 ;
  assign n44110 = n44106 & n44109 ;
  assign n44111 = x421 & x588 ;
  assign n44112 = ~n43968 & n44111 ;
  assign n44113 = n44110 | n44112 ;
  assign n44114 = n44104 | n44113 ;
  assign n44115 = ~n7103 & n44114 ;
  assign n44116 = ( ~x628 & x1134 ) | ( ~x628 & x1135 ) | ( x1134 & x1135 ) ;
  assign n44117 = ( x629 & ~x1134 ) | ( x629 & x1135 ) | ( ~x1134 & x1135 ) ;
  assign n44118 = ~n44116 & n44117 ;
  assign n44119 = n43460 & n44118 ;
  assign n44120 = x756 & n43286 ;
  assign n44121 = x734 & x1135 ;
  assign n44122 = x854 | x1136 ;
  assign n44123 = ~n44121 & n44122 ;
  assign n44124 = n43290 & n44123 ;
  assign n44125 = ~n44120 & n44124 ;
  assign n44126 = n44119 | n44125 ;
  assign n44127 = n7103 & n44126 ;
  assign n44128 = n44115 | n44127 ;
  assign n44129 = x461 & n43795 ;
  assign n44130 = x439 & n43301 ;
  assign n44131 = n44129 | n44130 ;
  assign n44132 = ~x591 & n44131 ;
  assign n44133 = x326 & ~x592 ;
  assign n44134 = n10558 & n44133 ;
  assign n44135 = n44132 | n44134 ;
  assign n44136 = ~x588 & n44135 ;
  assign n44137 = x449 & ~n43259 ;
  assign n44138 = n43804 & n44137 ;
  assign n44139 = n44136 | n44138 ;
  assign n44140 = ~n43264 & n44139 ;
  assign n44141 = x199 & ~x1057 ;
  assign n44142 = n43264 & ~n44141 ;
  assign n44143 = n38883 & n44142 ;
  assign n44144 = n44140 | n44143 ;
  assign n44145 = ~n7103 & n44144 ;
  assign n44146 = x867 & ~n43324 ;
  assign n44147 = ( ~x762 & x1135 ) | ( ~x762 & x1136 ) | ( x1135 & x1136 ) ;
  assign n44148 = ( x697 & x1135 ) | ( x697 & ~x1136 ) | ( x1135 & ~x1136 ) ;
  assign n44149 = n44147 & ~n44148 ;
  assign n44150 = n44146 | n44149 ;
  assign n44151 = n43289 & n44150 ;
  assign n44152 = x816 & ~n43275 ;
  assign n44153 = ~n43324 & n44152 ;
  assign n44154 = ( x653 & x1135 ) | ( x653 & x1136 ) | ( x1135 & x1136 ) ;
  assign n44155 = ( x693 & x1135 ) | ( x693 & ~x1136 ) | ( x1135 & ~x1136 ) ;
  assign n44156 = n44154 & ~n44155 ;
  assign n44157 = n44153 | n44156 ;
  assign n44158 = ~n43821 & n44157 ;
  assign n44159 = n44151 | n44158 ;
  assign n44160 = n7103 & n44159 ;
  assign n44161 = n44145 | n44160 ;
  assign n44162 = ( x962 & ~x1123 ) | ( x962 & n43129 ) | ( ~x1123 & n43129 ) ;
  assign n44163 = ( x715 & ~x962 ) | ( x715 & n43129 ) | ( ~x962 & n43129 ) ;
  assign n44164 = ~n44162 & n44163 ;
  assign n44165 = x440 & n43987 ;
  assign n44166 = x329 & x591 ;
  assign n44167 = ~n43989 & n44166 ;
  assign n44168 = n44165 | n44167 ;
  assign n44169 = ~x590 & n44168 ;
  assign n44170 = x349 & ~n43264 ;
  assign n44171 = n43260 & n44170 ;
  assign n44172 = n44169 | n44171 ;
  assign n44173 = ~x588 & n44172 ;
  assign n44174 = x199 & ~x1043 ;
  assign n44175 = n43264 & ~n44174 ;
  assign n44176 = ( x199 & x200 ) | ( x199 & x1053 ) | ( x200 & x1053 ) ;
  assign n44177 = ( x199 & ~x200 ) | ( x199 & x307 ) | ( ~x200 & x307 ) ;
  assign n44178 = n44176 | n44177 ;
  assign n44179 = n44175 & n44178 ;
  assign n44180 = x454 & n43804 ;
  assign n44181 = ~n44004 & n44180 ;
  assign n44182 = n7103 | n44181 ;
  assign n44183 = n44179 | n44182 ;
  assign n44184 = n44173 | n44183 ;
  assign n44185 = x761 & n43286 ;
  assign n44186 = x845 | x1136 ;
  assign n44187 = x738 & x1135 ;
  assign n44188 = x1134 & ~n44187 ;
  assign n44189 = n44186 & n44188 ;
  assign n44190 = ~n44011 & n44189 ;
  assign n44191 = ~n44185 & n44190 ;
  assign n44192 = ( ~x641 & x1134 ) | ( ~x641 & x1135 ) | ( x1134 & x1135 ) ;
  assign n44193 = ( x626 & ~x1134 ) | ( x626 & x1135 ) | ( ~x1134 & x1135 ) ;
  assign n44194 = ~n44192 & n44193 ;
  assign n44195 = n43460 & n44194 ;
  assign n44196 = n7103 & ~n44195 ;
  assign n44197 = ~n44191 & n44196 ;
  assign n44198 = n44184 & ~n44197 ;
  assign n44199 = x318 & x591 ;
  assign n44200 = ~x592 & n44199 ;
  assign n44201 = ~x591 & n6192 ;
  assign n44202 = n44200 | n44201 ;
  assign n44203 = ~x590 & n44202 ;
  assign n44204 = x462 & n43260 ;
  assign n44205 = n44203 | n44204 ;
  assign n44206 = ~n43960 & n44205 ;
  assign n44207 = x448 & x588 ;
  assign n44208 = ~n43968 & n44207 ;
  assign n44209 = ( x199 & n39383 ) | ( x199 & n43264 ) | ( n39383 & n43264 ) ;
  assign n44210 = ( ~x199 & x1074 ) | ( ~x199 & n43264 ) | ( x1074 & n43264 ) ;
  assign n44211 = n44209 & n44210 ;
  assign n44212 = n44208 | n44211 ;
  assign n44213 = n44206 | n44212 ;
  assign n44214 = ~n7103 & n44213 ;
  assign n44215 = x768 & n43286 ;
  assign n44216 = x839 | x1136 ;
  assign n44217 = ~x705 & x1135 ;
  assign n44218 = x1134 & ~n44217 ;
  assign n44219 = n44216 & n44218 ;
  assign n44220 = ~n44011 & n44219 ;
  assign n44221 = ~n44215 & n44220 ;
  assign n44222 = x800 & ~n43324 ;
  assign n44223 = ( x645 & x1135 ) | ( x645 & x1136 ) | ( x1135 & x1136 ) ;
  assign n44224 = ( x669 & x1135 ) | ( x669 & ~x1136 ) | ( x1135 & ~x1136 ) ;
  assign n44225 = n44223 & ~n44224 ;
  assign n44226 = n44222 | n44225 ;
  assign n44227 = ~n43276 & n44226 ;
  assign n44228 = n44221 | n44227 ;
  assign n44229 = n7103 & n44228 ;
  assign n44230 = n44214 | n44229 ;
  assign n44231 = x369 & n43987 ;
  assign n44232 = x394 & x591 ;
  assign n44233 = ~n43989 & n44232 ;
  assign n44234 = n44231 | n44233 ;
  assign n44235 = ~x590 & n44234 ;
  assign n44236 = x315 & ~n43264 ;
  assign n44237 = n43260 & n44236 ;
  assign n44238 = n44235 | n44237 ;
  assign n44239 = ~x588 & n44238 ;
  assign n44240 = x199 & ~x1080 ;
  assign n44241 = n43264 & ~n44240 ;
  assign n44242 = ( x199 & x200 ) | ( x199 & x1049 ) | ( x200 & x1049 ) ;
  assign n44243 = ( x199 & ~x200 ) | ( x199 & x303 ) | ( ~x200 & x303 ) ;
  assign n44244 = n44242 | n44243 ;
  assign n44245 = n44241 & n44244 ;
  assign n44246 = x419 & n43804 ;
  assign n44247 = ~n44004 & n44246 ;
  assign n44248 = n7103 | n44247 ;
  assign n44249 = n44245 | n44248 ;
  assign n44250 = n44239 | n44249 ;
  assign n44251 = x767 & n43286 ;
  assign n44252 = x853 | x1136 ;
  assign n44253 = x698 & x1135 ;
  assign n44254 = x1134 & ~n44253 ;
  assign n44255 = n44252 & n44254 ;
  assign n44256 = ~n44011 & n44255 ;
  assign n44257 = ~n44251 & n44256 ;
  assign n44258 = ( ~x625 & x1134 ) | ( ~x625 & x1135 ) | ( x1134 & x1135 ) ;
  assign n44259 = ( x608 & ~x1134 ) | ( x608 & x1135 ) | ( ~x1134 & x1135 ) ;
  assign n44260 = ~n44258 & n44259 ;
  assign n44261 = n43460 & n44260 ;
  assign n44262 = n7103 & ~n44261 ;
  assign n44263 = ~n44257 & n44262 ;
  assign n44264 = n44250 & ~n44263 ;
  assign n44265 = x378 & n43253 ;
  assign n44266 = x325 & x591 ;
  assign n44267 = ~x592 & n44266 ;
  assign n44268 = n44265 | n44267 ;
  assign n44269 = ~x590 & n44268 ;
  assign n44270 = x353 & n43260 ;
  assign n44271 = n44269 | n44270 ;
  assign n44272 = ~n43960 & n44271 ;
  assign n44273 = x451 & x588 ;
  assign n44274 = ~n43968 & n44273 ;
  assign n44275 = ( x199 & n39395 ) | ( x199 & n43264 ) | ( n39395 & n43264 ) ;
  assign n44276 = ( ~x199 & x1063 ) | ( ~x199 & n43264 ) | ( x1063 & n43264 ) ;
  assign n44277 = n44275 & n44276 ;
  assign n44278 = n44274 | n44277 ;
  assign n44279 = n44272 | n44278 ;
  assign n44280 = ~n7103 & n44279 ;
  assign n44281 = x774 & n43286 ;
  assign n44282 = x868 | x1136 ;
  assign n44283 = ~x687 & x1135 ;
  assign n44284 = x1134 & ~n44283 ;
  assign n44285 = n44282 & n44284 ;
  assign n44286 = ~n44011 & n44285 ;
  assign n44287 = ~n44281 & n44286 ;
  assign n44288 = x807 & ~n43324 ;
  assign n44289 = ( x636 & x1135 ) | ( x636 & x1136 ) | ( x1135 & x1136 ) ;
  assign n44290 = ( x650 & x1135 ) | ( x650 & ~x1136 ) | ( x1135 & ~x1136 ) ;
  assign n44291 = n44289 & ~n44290 ;
  assign n44292 = n44288 | n44291 ;
  assign n44293 = ~n43276 & n44292 ;
  assign n44294 = n44287 | n44293 ;
  assign n44295 = n7103 & n44294 ;
  assign n44296 = n44280 | n44295 ;
  assign n44297 = x356 & n43795 ;
  assign n44298 = x381 & n43301 ;
  assign n44299 = n44297 | n44298 ;
  assign n44300 = ~x591 & n44299 ;
  assign n44301 = x405 & ~x592 ;
  assign n44302 = n10558 & n44301 ;
  assign n44303 = n44300 | n44302 ;
  assign n44304 = ~x588 & n44303 ;
  assign n44305 = x445 & ~n43259 ;
  assign n44306 = n43804 & n44305 ;
  assign n44307 = n44304 | n44306 ;
  assign n44308 = ~n43264 & n44307 ;
  assign n44309 = x199 & ~x1081 ;
  assign n44310 = n43264 & ~n44309 ;
  assign n44311 = n39413 & n44310 ;
  assign n44312 = n44308 | n44311 ;
  assign n44313 = ~n7103 & n44312 ;
  assign n44314 = x880 & ~n43324 ;
  assign n44315 = ( ~x750 & x1135 ) | ( ~x750 & x1136 ) | ( x1135 & x1136 ) ;
  assign n44316 = ( x684 & x1135 ) | ( x684 & ~x1136 ) | ( x1135 & ~x1136 ) ;
  assign n44317 = n44315 & ~n44316 ;
  assign n44318 = n44314 | n44317 ;
  assign n44319 = n43289 & n44318 ;
  assign n44320 = x794 & ~n43275 ;
  assign n44321 = ~n43324 & n44320 ;
  assign n44322 = ( x651 & x1135 ) | ( x651 & x1136 ) | ( x1135 & x1136 ) ;
  assign n44323 = ( x654 & x1135 ) | ( x654 & ~x1136 ) | ( x1135 & ~x1136 ) ;
  assign n44324 = n44322 & ~n44323 ;
  assign n44325 = n44321 | n44324 ;
  assign n44326 = ~n43821 & n44325 ;
  assign n44327 = n44319 | n44326 ;
  assign n44328 = n7103 & n44327 ;
  assign n44329 = n44313 | n44328 ;
  assign n44330 = x721 & x813 ;
  assign n44331 = x773 | x801 ;
  assign n44332 = x773 & x801 ;
  assign n44333 = n44331 & ~n44332 ;
  assign n44334 = x771 | x800 ;
  assign n44335 = x771 & x800 ;
  assign n44336 = n44334 & ~n44335 ;
  assign n44337 = x769 | x794 ;
  assign n44338 = x769 & x794 ;
  assign n44339 = n44337 & ~n44338 ;
  assign n44340 = x765 | x798 ;
  assign n44341 = x765 & x798 ;
  assign n44342 = n44340 & ~n44341 ;
  assign n44343 = x807 & ~n44342 ;
  assign n44344 = x747 & n44343 ;
  assign n44345 = x747 | x807 ;
  assign n44346 = n44342 | n44345 ;
  assign n44347 = ~n44344 & n44346 ;
  assign n44348 = n44339 | n44347 ;
  assign n44349 = n44336 | n44348 ;
  assign n44350 = n44333 | n44349 ;
  assign n44351 = n44330 & ~n44350 ;
  assign n44352 = ~n44336 & n44343 ;
  assign n44353 = x721 | x813 ;
  assign n44354 = x794 & x801 ;
  assign n44355 = ~n44353 & n44354 ;
  assign n44356 = n44352 & n44355 ;
  assign n44357 = n44351 | n44356 ;
  assign n44358 = x816 & n44357 ;
  assign n44359 = x747 & x773 ;
  assign n44360 = x769 & n44359 ;
  assign n44361 = ~x721 & n44360 ;
  assign n44362 = ( x775 & ~n44360 ) | ( x775 & n44361 ) | ( ~n44360 & n44361 ) ;
  assign n44363 = ( x721 & n44361 ) | ( x721 & n44362 ) | ( n44361 & n44362 ) ;
  assign n44364 = ~n44358 & n44363 ;
  assign n44365 = x795 & ~n44364 ;
  assign n44366 = ~x945 & x988 ;
  assign n44367 = x731 & n44366 ;
  assign n44368 = x721 & ~x775 ;
  assign n44369 = n44363 | n44368 ;
  assign n44370 = n44367 & n44369 ;
  assign n44371 = ~n44365 & n44370 ;
  assign n44372 = x775 | x816 ;
  assign n44373 = x775 & x816 ;
  assign n44374 = n44372 & ~n44373 ;
  assign n44375 = n44351 & ~n44374 ;
  assign n44376 = n44368 & ~n44375 ;
  assign n44377 = x731 | x795 ;
  assign n44378 = x731 & x795 ;
  assign n44379 = n44377 & ~n44378 ;
  assign n44380 = n44375 & ~n44379 ;
  assign n44381 = x721 & ~n44367 ;
  assign n44382 = ( n44376 & ~n44380 ) | ( n44376 & n44381 ) | ( ~n44380 & n44381 ) ;
  assign n44383 = n44371 | n44382 ;
  assign n44384 = x379 & n43253 ;
  assign n44385 = x403 & x591 ;
  assign n44386 = ~x592 & n44385 ;
  assign n44387 = n44384 | n44386 ;
  assign n44388 = ~x590 & n44387 ;
  assign n44389 = x354 & n43260 ;
  assign n44390 = n44388 | n44389 ;
  assign n44391 = ~n43960 & n44390 ;
  assign n44392 = x428 & x588 ;
  assign n44393 = ~n43968 & n44392 ;
  assign n44394 = ( x199 & n39401 ) | ( x199 & n43264 ) | ( n39401 & n43264 ) ;
  assign n44395 = ( ~x199 & x1045 ) | ( ~x199 & n43264 ) | ( x1045 & n43264 ) ;
  assign n44396 = n44394 & n44395 ;
  assign n44397 = n44393 | n44396 ;
  assign n44398 = n44391 | n44397 ;
  assign n44399 = ~n7103 & n44398 ;
  assign n44400 = ( ~x851 & x1134 ) | ( ~x851 & x1136 ) | ( x1134 & x1136 ) ;
  assign n44401 = ( x795 & x1134 ) | ( x795 & ~x1136 ) | ( x1134 & ~x1136 ) ;
  assign n44402 = ~n44400 & n44401 ;
  assign n44403 = ( x640 & x1134 ) | ( x640 & x1136 ) | ( x1134 & x1136 ) ;
  assign n44404 = ( x776 & x1134 ) | ( x776 & ~x1136 ) | ( x1134 & ~x1136 ) ;
  assign n44405 = n44403 & ~n44404 ;
  assign n44406 = n44402 | n44405 ;
  assign n44407 = ~x1135 & n44406 ;
  assign n44408 = ( x694 & x1134 ) | ( x694 & ~n43607 ) | ( x1134 & ~n43607 ) ;
  assign n44409 = ( ~x732 & x1134 ) | ( ~x732 & n43607 ) | ( x1134 & n43607 ) ;
  assign n44410 = ~n44408 & n44409 ;
  assign n44411 = n44407 | n44410 ;
  assign n44412 = n43331 & n44411 ;
  assign n44413 = n44399 | n44412 ;
  assign n44414 = ( x962 & ~x1111 ) | ( x962 & n43791 ) | ( ~x1111 & n43791 ) ;
  assign n44415 = ( x723 & x962 ) | ( x723 & ~n43791 ) | ( x962 & ~n43791 ) ;
  assign n44416 = n44414 | n44415 ;
  assign n44417 = ( x962 & ~x1114 ) | ( x962 & n43791 ) | ( ~x1114 & n43791 ) ;
  assign n44418 = ( x724 & x962 ) | ( x724 & ~n43791 ) | ( x962 & ~n43791 ) ;
  assign n44419 = n44417 | n44418 ;
  assign n44420 = ( x962 & ~x1120 ) | ( x962 & n43791 ) | ( ~x1120 & n43791 ) ;
  assign n44421 = ( x725 & x962 ) | ( x725 & ~n43791 ) | ( x962 & ~n43791 ) ;
  assign n44422 = n44420 | n44421 ;
  assign n44423 = ( x962 & ~x1126 ) | ( x962 & n43791 ) | ( ~x1126 & n43791 ) ;
  assign n44424 = ( x726 & ~x962 ) | ( x726 & n43791 ) | ( ~x962 & n43791 ) ;
  assign n44425 = ~n44423 & n44424 ;
  assign n44426 = ( x962 & ~x1102 ) | ( x962 & n43791 ) | ( ~x1102 & n43791 ) ;
  assign n44427 = ( x727 & ~x962 ) | ( x727 & n43791 ) | ( ~x962 & n43791 ) ;
  assign n44428 = ~n44426 & n44427 ;
  assign n44429 = ( x962 & ~x1131 ) | ( x962 & n43791 ) | ( ~x1131 & n43791 ) ;
  assign n44430 = ( x728 & x962 ) | ( x728 & ~n43791 ) | ( x962 & ~n43791 ) ;
  assign n44431 = n44429 | n44430 ;
  assign n44432 = ( x962 & ~x1104 ) | ( x962 & n43791 ) | ( ~x1104 & n43791 ) ;
  assign n44433 = ( x729 & ~x962 ) | ( x729 & n43791 ) | ( ~x962 & n43791 ) ;
  assign n44434 = ~n44432 & n44433 ;
  assign n44435 = ( x962 & ~x1106 ) | ( x962 & n43791 ) | ( ~x1106 & n43791 ) ;
  assign n44436 = ( x730 & ~x962 ) | ( x730 & n43791 ) | ( ~x962 & n43791 ) ;
  assign n44437 = ~n44435 & n44436 ;
  assign n44438 = ~n44330 & n44353 ;
  assign n44439 = n44350 | n44438 ;
  assign n44440 = x795 & ~n44374 ;
  assign n44441 = ~n44439 & n44440 ;
  assign n44442 = n44359 | n44441 ;
  assign n44443 = n44367 & n44442 ;
  assign n44444 = x731 & ~n44441 ;
  assign n44445 = n44374 | n44438 ;
  assign n44446 = ~x795 & x801 ;
  assign n44447 = ~n44339 & n44446 ;
  assign n44448 = ~n44445 & n44447 ;
  assign n44449 = n44352 & n44448 ;
  assign n44450 = n44359 & ~n44449 ;
  assign n44451 = x731 | n44450 ;
  assign n44452 = ( n44366 & n44444 ) | ( n44366 & n44451 ) | ( n44444 & n44451 ) ;
  assign n44453 = ~n44443 & n44452 ;
  assign n44454 = ( x962 & ~x1128 ) | ( x962 & n43129 ) | ( ~x1128 & n43129 ) ;
  assign n44455 = ( x732 & x962 ) | ( x732 & ~n43129 ) | ( x962 & ~n43129 ) ;
  assign n44456 = n44454 | n44455 ;
  assign n44457 = x375 & n43987 ;
  assign n44458 = x399 & x591 ;
  assign n44459 = ~n43989 & n44458 ;
  assign n44460 = n44457 | n44459 ;
  assign n44461 = ~x590 & n44460 ;
  assign n44462 = x316 & ~n43264 ;
  assign n44463 = n43260 & n44462 ;
  assign n44464 = n44461 | n44463 ;
  assign n44465 = ~x588 & n44464 ;
  assign n44466 = x199 & ~x1047 ;
  assign n44467 = n43264 & ~n44466 ;
  assign n44468 = ( x199 & x200 ) | ( x199 & x1037 ) | ( x200 & x1037 ) ;
  assign n44469 = ( x199 & ~x200 ) | ( x199 & x308 ) | ( ~x200 & x308 ) ;
  assign n44470 = n44468 | n44469 ;
  assign n44471 = n44467 & n44470 ;
  assign n44472 = x424 & n43804 ;
  assign n44473 = ~n44004 & n44472 ;
  assign n44474 = n7103 | n44473 ;
  assign n44475 = n44471 | n44474 ;
  assign n44476 = n44465 | n44475 ;
  assign n44477 = x777 & n43286 ;
  assign n44478 = x838 | x1136 ;
  assign n44479 = x737 & x1135 ;
  assign n44480 = x1134 & ~n44479 ;
  assign n44481 = n44478 & n44480 ;
  assign n44482 = ~n44011 & n44481 ;
  assign n44483 = ~n44477 & n44482 ;
  assign n44484 = ( ~x648 & x1134 ) | ( ~x648 & x1135 ) | ( x1134 & x1135 ) ;
  assign n44485 = ( x619 & ~x1134 ) | ( x619 & x1135 ) | ( ~x1134 & x1135 ) ;
  assign n44486 = ~n44484 & n44485 ;
  assign n44487 = n43460 & n44486 ;
  assign n44488 = n7103 & ~n44487 ;
  assign n44489 = ~n44483 & n44488 ;
  assign n44490 = n44476 & ~n44489 ;
  assign n44491 = ( x962 & ~x1119 ) | ( x962 & n43791 ) | ( ~x1119 & n43791 ) ;
  assign n44492 = ( x734 & x962 ) | ( x734 & ~n43791 ) | ( x962 & ~n43791 ) ;
  assign n44493 = n44491 | n44492 ;
  assign n44494 = ( x962 & ~x1109 ) | ( x962 & n43791 ) | ( ~x1109 & n43791 ) ;
  assign n44495 = ( x735 & ~x962 ) | ( x735 & n43791 ) | ( ~x962 & n43791 ) ;
  assign n44496 = ~n44494 & n44495 ;
  assign n44497 = ( x962 & ~x1101 ) | ( x962 & n43791 ) | ( ~x1101 & n43791 ) ;
  assign n44498 = ( x736 & ~x962 ) | ( x736 & n43791 ) | ( ~x962 & n43791 ) ;
  assign n44499 = ~n44497 & n44498 ;
  assign n44500 = ( x962 & ~x1122 ) | ( x962 & n43791 ) | ( ~x1122 & n43791 ) ;
  assign n44501 = ( x737 & x962 ) | ( x737 & ~n43791 ) | ( x962 & ~n43791 ) ;
  assign n44502 = n44500 | n44501 ;
  assign n44503 = ( x962 & ~x1121 ) | ( x962 & n43791 ) | ( ~x1121 & n43791 ) ;
  assign n44504 = ( x738 & x962 ) | ( x738 & ~n43791 ) | ( x962 & ~n43791 ) ;
  assign n44505 = n44503 | n44504 ;
  assign n44506 = x952 | x1061 ;
  assign n44507 = n43034 & ~n44506 ;
  assign n44508 = x832 & n44507 ;
  assign n44509 = ( x966 & x1108 ) | ( x966 & n44508 ) | ( x1108 & n44508 ) ;
  assign n44510 = ( x739 & x966 ) | ( x739 & ~n44508 ) | ( x966 & ~n44508 ) ;
  assign n44511 = n44509 | n44510 ;
  assign n44512 = ( x966 & x1114 ) | ( x966 & n44508 ) | ( x1114 & n44508 ) ;
  assign n44513 = ( x741 & ~x966 ) | ( x741 & n44508 ) | ( ~x966 & n44508 ) ;
  assign n44514 = ~n44512 & n44513 ;
  assign n44515 = ( x966 & x1112 ) | ( x966 & n44508 ) | ( x1112 & n44508 ) ;
  assign n44516 = ( x742 & ~x966 ) | ( x742 & n44508 ) | ( ~x966 & n44508 ) ;
  assign n44517 = ~n44515 & n44516 ;
  assign n44518 = ( x966 & x1109 ) | ( x966 & n44508 ) | ( x1109 & n44508 ) ;
  assign n44519 = ( x743 & x966 ) | ( x743 & ~n44508 ) | ( x966 & ~n44508 ) ;
  assign n44520 = n44518 | n44519 ;
  assign n44521 = ( x966 & x1131 ) | ( x966 & n44508 ) | ( x1131 & n44508 ) ;
  assign n44522 = ( x744 & ~x966 ) | ( x744 & n44508 ) | ( ~x966 & n44508 ) ;
  assign n44523 = ~n44521 & n44522 ;
  assign n44524 = ( x966 & x1111 ) | ( x966 & n44508 ) | ( x1111 & n44508 ) ;
  assign n44525 = ( x745 & ~x966 ) | ( x745 & n44508 ) | ( ~x966 & n44508 ) ;
  assign n44526 = ~n44524 & n44525 ;
  assign n44527 = ( x966 & x1104 ) | ( x966 & n44508 ) | ( x1104 & n44508 ) ;
  assign n44528 = ( x746 & x966 ) | ( x746 & ~n44508 ) | ( x966 & ~n44508 ) ;
  assign n44529 = n44527 | n44528 ;
  assign n44530 = x773 & n44366 ;
  assign n44531 = x747 | n44530 ;
  assign n44532 = x801 & ~n44346 ;
  assign n44533 = n44333 | n44530 ;
  assign n44534 = n44343 & ~n44533 ;
  assign n44535 = n44532 | n44534 ;
  assign n44536 = n44379 | n44445 ;
  assign n44537 = n44336 | n44339 ;
  assign n44538 = n44536 | n44537 ;
  assign n44539 = n44535 & ~n44538 ;
  assign n44540 = ( x747 & n44530 ) | ( x747 & n44539 ) | ( n44530 & n44539 ) ;
  assign n44541 = n44531 & ~n44540 ;
  assign n44542 = ( x966 & x1106 ) | ( x966 & n44508 ) | ( x1106 & n44508 ) ;
  assign n44543 = ( x748 & x966 ) | ( x748 & ~n44508 ) | ( x966 & ~n44508 ) ;
  assign n44544 = n44542 | n44543 ;
  assign n44545 = ( x966 & x1105 ) | ( x966 & n44508 ) | ( x1105 & n44508 ) ;
  assign n44546 = ( x749 & x966 ) | ( x749 & ~n44508 ) | ( x966 & ~n44508 ) ;
  assign n44547 = n44545 | n44546 ;
  assign n44548 = ( x966 & x1130 ) | ( x966 & n44508 ) | ( x1130 & n44508 ) ;
  assign n44549 = ( x750 & ~x966 ) | ( x750 & n44508 ) | ( ~x966 & n44508 ) ;
  assign n44550 = ~n44548 & n44549 ;
  assign n44551 = ( x966 & x1123 ) | ( x966 & n44508 ) | ( x1123 & n44508 ) ;
  assign n44552 = ( x751 & ~x966 ) | ( x751 & n44508 ) | ( ~x966 & n44508 ) ;
  assign n44553 = ~n44551 & n44552 ;
  assign n44554 = ( x966 & x1124 ) | ( x966 & n44508 ) | ( x1124 & n44508 ) ;
  assign n44555 = ( x752 & ~x966 ) | ( x752 & n44508 ) | ( ~x966 & n44508 ) ;
  assign n44556 = ~n44554 & n44555 ;
  assign n44557 = ( x966 & x1117 ) | ( x966 & n44508 ) | ( x1117 & n44508 ) ;
  assign n44558 = ( x753 & ~x966 ) | ( x753 & n44508 ) | ( ~x966 & n44508 ) ;
  assign n44559 = ~n44557 & n44558 ;
  assign n44560 = ( x966 & x1118 ) | ( x966 & n44508 ) | ( x1118 & n44508 ) ;
  assign n44561 = ( x754 & ~x966 ) | ( x754 & n44508 ) | ( ~x966 & n44508 ) ;
  assign n44562 = ~n44560 & n44561 ;
  assign n44563 = ( x966 & x1120 ) | ( x966 & n44508 ) | ( x1120 & n44508 ) ;
  assign n44564 = ( x755 & ~x966 ) | ( x755 & n44508 ) | ( ~x966 & n44508 ) ;
  assign n44565 = ~n44563 & n44564 ;
  assign n44566 = ( x966 & x1119 ) | ( x966 & n44508 ) | ( x1119 & n44508 ) ;
  assign n44567 = ( x756 & ~x966 ) | ( x756 & n44508 ) | ( ~x966 & n44508 ) ;
  assign n44568 = ~n44566 & n44567 ;
  assign n44569 = ( x966 & x1113 ) | ( x966 & n44508 ) | ( x1113 & n44508 ) ;
  assign n44570 = ( x757 & ~x966 ) | ( x757 & n44508 ) | ( ~x966 & n44508 ) ;
  assign n44571 = ~n44569 & n44570 ;
  assign n44572 = ( x966 & x1101 ) | ( x966 & n44508 ) | ( x1101 & n44508 ) ;
  assign n44573 = ( x758 & x966 ) | ( x758 & ~n44508 ) | ( x966 & ~n44508 ) ;
  assign n44574 = n44572 | n44573 ;
  assign n44575 = x759 | n44508 ;
  assign n44576 = n43039 & n44507 ;
  assign n44577 = n44575 & ~n44576 ;
  assign n44578 = x966 | n44577 ;
  assign n44579 = ( x966 & x1115 ) | ( x966 & n44508 ) | ( x1115 & n44508 ) ;
  assign n44580 = ( x760 & ~x966 ) | ( x760 & n44508 ) | ( ~x966 & n44508 ) ;
  assign n44581 = ~n44579 & n44580 ;
  assign n44582 = ( x966 & x1121 ) | ( x966 & n44508 ) | ( x1121 & n44508 ) ;
  assign n44583 = ( x761 & ~x966 ) | ( x761 & n44508 ) | ( ~x966 & n44508 ) ;
  assign n44584 = ~n44582 & n44583 ;
  assign n44585 = ( x966 & x1129 ) | ( x966 & n44508 ) | ( x1129 & n44508 ) ;
  assign n44586 = ( x762 & ~x966 ) | ( x762 & n44508 ) | ( ~x966 & n44508 ) ;
  assign n44587 = ~n44585 & n44586 ;
  assign n44588 = ( x966 & x1103 ) | ( x966 & n44508 ) | ( x1103 & n44508 ) ;
  assign n44589 = ( x763 & x966 ) | ( x763 & ~n44508 ) | ( x966 & ~n44508 ) ;
  assign n44590 = n44588 | n44589 ;
  assign n44591 = ( x966 & x1107 ) | ( x966 & n44508 ) | ( x1107 & n44508 ) ;
  assign n44592 = ( x764 & x966 ) | ( x764 & ~n44508 ) | ( x966 & ~n44508 ) ;
  assign n44593 = n44591 | n44592 ;
  assign n44594 = n44350 | n44536 ;
  assign n44595 = x765 & n44594 ;
  assign n44596 = x945 & ~n44595 ;
  assign n44597 = ~n44351 & n44353 ;
  assign n44598 = x765 | n44335 ;
  assign n44599 = n44338 | n44598 ;
  assign n44600 = n44344 | n44599 ;
  assign n44601 = ~n44331 & n44600 ;
  assign n44602 = n44332 | n44601 ;
  assign n44603 = ~n44349 & n44602 ;
  assign n44604 = x721 | n44603 ;
  assign n44605 = ~n44372 & n44604 ;
  assign n44606 = ~n44597 & n44605 ;
  assign n44607 = n44373 & ~n44439 ;
  assign n44608 = x765 | n44607 ;
  assign n44609 = n44606 | n44608 ;
  assign n44610 = ~x795 & n44609 ;
  assign n44611 = x731 | n44610 ;
  assign n44612 = x795 | n44611 ;
  assign n44613 = ~n44444 & n44611 ;
  assign n44614 = ( x765 & n44612 ) | ( x765 & n44613 ) | ( n44612 & n44613 ) ;
  assign n44615 = ~x945 & n44614 ;
  assign n44616 = n44596 | n44615 ;
  assign n44617 = ( x966 & x1110 ) | ( x966 & n44508 ) | ( x1110 & n44508 ) ;
  assign n44618 = ( x766 & x966 ) | ( x766 & ~n44508 ) | ( x966 & ~n44508 ) ;
  assign n44619 = n44617 | n44618 ;
  assign n44620 = ( x966 & x1116 ) | ( x966 & n44508 ) | ( x1116 & n44508 ) ;
  assign n44621 = ( x767 & ~x966 ) | ( x767 & n44508 ) | ( ~x966 & n44508 ) ;
  assign n44622 = ~n44620 & n44621 ;
  assign n44623 = ( x966 & x1125 ) | ( x966 & n44508 ) | ( x1125 & n44508 ) ;
  assign n44624 = ( x768 & ~x966 ) | ( x768 & n44508 ) | ( ~x966 & n44508 ) ;
  assign n44625 = ~n44623 & n44624 ;
  assign n44626 = x794 & ~n44333 ;
  assign n44627 = ~n44336 & n44626 ;
  assign n44628 = ~n44445 & n44627 ;
  assign n44629 = ~n44347 & n44628 ;
  assign n44630 = ~n44379 & n44629 ;
  assign n44631 = x769 & ~n44367 ;
  assign n44632 = ~n44630 & n44631 ;
  assign n44633 = x775 & n44359 ;
  assign n44634 = ( x769 & ~n44367 ) | ( x769 & n44633 ) | ( ~n44367 & n44633 ) ;
  assign n44635 = ~x775 & n44629 ;
  assign n44636 = n44607 | n44635 ;
  assign n44637 = x795 & n44636 ;
  assign n44638 = ( x769 & n44633 ) | ( x769 & ~n44637 ) | ( n44633 & ~n44637 ) ;
  assign n44639 = ~n44634 & n44638 ;
  assign n44640 = n44632 | n44639 ;
  assign n44641 = ( x966 & x1126 ) | ( x966 & n44508 ) | ( x1126 & n44508 ) ;
  assign n44642 = ( x770 & ~x966 ) | ( x770 & n44508 ) | ( ~x966 & n44508 ) ;
  assign n44643 = ~n44641 & n44642 ;
  assign n44644 = n44373 | n44605 ;
  assign n44645 = ~n44377 & n44644 ;
  assign n44646 = ~n44374 & n44378 ;
  assign n44647 = n44645 | n44646 ;
  assign n44648 = ~n44439 & n44647 ;
  assign n44649 = ~x945 & x987 ;
  assign n44650 = ~n44648 & n44649 ;
  assign n44651 = x771 & x945 ;
  assign n44652 = n44594 & n44651 ;
  assign n44653 = n44650 | n44652 ;
  assign n44654 = ( x966 & x1102 ) | ( x966 & n44508 ) | ( x1102 & n44508 ) ;
  assign n44655 = ( x772 & x966 ) | ( x772 & ~n44508 ) | ( x966 & ~n44508 ) ;
  assign n44656 = n44654 | n44655 ;
  assign n44657 = x801 | n44349 ;
  assign n44658 = n44648 & ~n44657 ;
  assign n44659 = n44366 & ~n44658 ;
  assign n44660 = x801 & n44536 ;
  assign n44661 = n44350 | n44660 ;
  assign n44662 = x773 & n44661 ;
  assign n44663 = n44659 | n44662 ;
  assign n44664 = ~n44530 & n44663 ;
  assign n44665 = ( x966 & x1127 ) | ( x966 & n44508 ) | ( x1127 & n44508 ) ;
  assign n44666 = ( x774 & ~x966 ) | ( x774 & n44508 ) | ( ~x966 & n44508 ) ;
  assign n44667 = ~n44665 & n44666 ;
  assign n44668 = x765 & x771 ;
  assign n44669 = n44359 & n44668 ;
  assign n44670 = n44441 | n44669 ;
  assign n44671 = x731 & ~x945 ;
  assign n44672 = x775 & n44671 ;
  assign n44673 = n44670 & n44672 ;
  assign n44674 = n44594 | n44671 ;
  assign n44675 = x795 & x800 ;
  assign n44676 = x801 & ~x816 ;
  assign n44677 = n44675 & n44676 ;
  assign n44678 = ~n44438 & n44677 ;
  assign n44679 = ~n44348 & n44678 ;
  assign n44680 = n44669 & ~n44679 ;
  assign n44681 = n44671 & n44680 ;
  assign n44682 = ( x775 & n44674 ) | ( x775 & n44681 ) | ( n44674 & n44681 ) ;
  assign n44683 = ~n44673 & n44682 ;
  assign n44684 = ( x966 & x1128 ) | ( x966 & n44508 ) | ( x1128 & n44508 ) ;
  assign n44685 = ( x776 & ~x966 ) | ( x776 & n44508 ) | ( ~x966 & n44508 ) ;
  assign n44686 = ~n44684 & n44685 ;
  assign n44687 = ( x966 & x1122 ) | ( x966 & n44508 ) | ( x1122 & n44508 ) ;
  assign n44688 = ( x777 & ~x966 ) | ( x777 & n44508 ) | ( ~x966 & n44508 ) ;
  assign n44689 = ~n44687 & n44688 ;
  assign n44690 = x832 & x956 ;
  assign n44691 = x1046 | x1083 ;
  assign n44692 = x1085 & ~n44691 ;
  assign n44693 = n44690 & n44692 ;
  assign n44694 = ~x968 & n44693 ;
  assign n44695 = x778 & ~n44694 ;
  assign n44696 = x1100 & n44694 ;
  assign n44697 = n44695 | n44696 ;
  assign n44698 = x779 & ~n43087 ;
  assign n44699 = x780 & ~n43008 ;
  assign n44700 = x781 & ~n44694 ;
  assign n44701 = x1101 & n44694 ;
  assign n44702 = n44700 | n44701 ;
  assign n44703 = n38887 & ~n43049 ;
  assign n44704 = n43007 & n44703 ;
  assign n44705 = x783 & ~n44694 ;
  assign n44706 = x1109 & n44694 ;
  assign n44707 = n44705 | n44706 ;
  assign n44708 = x784 & ~n44694 ;
  assign n44709 = x1110 & n44694 ;
  assign n44710 = n44708 | n44709 ;
  assign n44711 = x785 & ~n44694 ;
  assign n44712 = x1102 & n44694 ;
  assign n44713 = n44711 | n44712 ;
  assign n44714 = x24 & ~x954 ;
  assign n44715 = x786 & x954 ;
  assign n44716 = n44714 | n44715 ;
  assign n44717 = x787 & ~n44694 ;
  assign n44718 = x1104 & n44694 ;
  assign n44719 = n44717 | n44718 ;
  assign n44720 = x788 & ~n44694 ;
  assign n44721 = x1105 & n44694 ;
  assign n44722 = n44720 | n44721 ;
  assign n44723 = x789 & ~n44694 ;
  assign n44724 = x1106 & n44694 ;
  assign n44725 = n44723 | n44724 ;
  assign n44726 = x790 & ~n44694 ;
  assign n44727 = x1107 & n44694 ;
  assign n44728 = n44726 | n44727 ;
  assign n44729 = x791 & ~n44694 ;
  assign n44730 = x1108 & n44694 ;
  assign n44731 = n44729 | n44730 ;
  assign n44732 = x792 & ~n44694 ;
  assign n44733 = x1103 & n44694 ;
  assign n44734 = n44732 | n44733 ;
  assign n44735 = x968 & n44693 ;
  assign n44736 = x794 & ~n44735 ;
  assign n44737 = x1130 & n44735 ;
  assign n44738 = n44736 | n44737 ;
  assign n44739 = x795 & ~n44735 ;
  assign n44740 = x1128 & n44735 ;
  assign n44741 = n44739 | n44740 ;
  assign n44742 = x266 & ~x269 ;
  assign n44743 = x278 & x279 ;
  assign n44744 = ~x280 & n44743 ;
  assign n44745 = n44742 & n44744 ;
  assign n44746 = ~x281 & n44745 ;
  assign n44747 = ~n43237 & n44746 ;
  assign n44748 = x264 & ~n44747 ;
  assign n44749 = ~x264 & n44747 ;
  assign n44750 = n44748 | n44749 ;
  assign n44751 = x798 & ~n44735 ;
  assign n44752 = x1124 & n44735 ;
  assign n44753 = n44751 | n44752 ;
  assign n44754 = x799 & ~n44735 ;
  assign n44755 = ~x1107 & n44735 ;
  assign n44756 = n44754 | n44755 ;
  assign n44757 = x800 & ~n44735 ;
  assign n44758 = x1125 & n44735 ;
  assign n44759 = n44757 | n44758 ;
  assign n44760 = x801 & ~n44735 ;
  assign n44761 = x1126 & n44735 ;
  assign n44762 = n44760 | n44761 ;
  assign n44763 = x803 & ~n44735 ;
  assign n44764 = ~x1106 & n44735 ;
  assign n44765 = n44763 | n44764 ;
  assign n44766 = x804 & ~n44735 ;
  assign n44767 = x1109 & n44735 ;
  assign n44768 = n44766 | n44767 ;
  assign n44769 = ~x282 & n43235 ;
  assign n44770 = ~x270 & n44769 ;
  assign n44771 = x270 & ~n44769 ;
  assign n44772 = n44770 | n44771 ;
  assign n44773 = x807 & ~n44735 ;
  assign n44774 = x1127 & n44735 ;
  assign n44775 = n44773 | n44774 ;
  assign n44776 = x808 & ~n44735 ;
  assign n44777 = x1101 & n44735 ;
  assign n44778 = n44776 | n44777 ;
  assign n44779 = x809 & ~n44735 ;
  assign n44780 = ~x1103 & n44735 ;
  assign n44781 = n44779 | n44780 ;
  assign n44782 = x810 & ~n44735 ;
  assign n44783 = x1108 & n44735 ;
  assign n44784 = n44782 | n44783 ;
  assign n44785 = x811 & ~n44735 ;
  assign n44786 = x1102 & n44735 ;
  assign n44787 = n44785 | n44786 ;
  assign n44788 = x812 & ~n44735 ;
  assign n44789 = ~x1104 & n44735 ;
  assign n44790 = n44788 | n44789 ;
  assign n44791 = x813 & ~n44735 ;
  assign n44792 = x1131 & n44735 ;
  assign n44793 = n44791 | n44792 ;
  assign n44794 = x814 & ~n44735 ;
  assign n44795 = ~x1105 & n44735 ;
  assign n44796 = n44794 | n44795 ;
  assign n44797 = x815 & ~n44735 ;
  assign n44798 = x1110 & n44735 ;
  assign n44799 = n44797 | n44798 ;
  assign n44800 = x816 & ~n44735 ;
  assign n44801 = x1129 & n44735 ;
  assign n44802 = n44800 | n44801 ;
  assign n44803 = x269 & ~n43233 ;
  assign n44804 = n43234 | n44803 ;
  assign n44805 = ~n7103 & n12151 ;
  assign n44806 = n12011 | n44805 ;
  assign n44807 = x265 & ~n43239 ;
  assign n44808 = n43240 | n44807 ;
  assign n44809 = x277 & ~n44770 ;
  assign n44810 = n43238 | n44809 ;
  assign n44811 = x811 | x893 ;
  assign n44812 = x982 | n8243 ;
  assign n44813 = n5995 & ~n7103 ;
  assign n44814 = n44812 & ~n44813 ;
  assign n44815 = n1692 & ~n44814 ;
  assign n44816 = x123 & ~n1873 ;
  assign n44817 = x1131 & ~n44816 ;
  assign n44818 = x1127 & ~n44816 ;
  assign n44819 = n44817 | n44818 ;
  assign n44820 = ~x825 & n44816 ;
  assign n44821 = n44819 | n44820 ;
  assign n44822 = x1131 & n44818 ;
  assign n44823 = n44821 & ~n44822 ;
  assign n44824 = x1125 | x1126 ;
  assign n44825 = x1125 & x1126 ;
  assign n44826 = n44824 & ~n44825 ;
  assign n44827 = ( x1128 & ~x1129 ) | ( x1128 & n44826 ) | ( ~x1129 & n44826 ) ;
  assign n44828 = ( ~x1128 & x1129 ) | ( ~x1128 & n44827 ) | ( x1129 & n44827 ) ;
  assign n44829 = ( ~n44826 & n44827 ) | ( ~n44826 & n44828 ) | ( n44827 & n44828 ) ;
  assign n44830 = ( x1124 & ~x1130 ) | ( x1124 & n44829 ) | ( ~x1130 & n44829 ) ;
  assign n44831 = ( ~x1124 & x1130 ) | ( ~x1124 & n44830 ) | ( x1130 & n44830 ) ;
  assign n44832 = ( ~n44829 & n44830 ) | ( ~n44829 & n44831 ) | ( n44830 & n44831 ) ;
  assign n44833 = n44823 | n44832 ;
  assign n44834 = x825 & n44816 ;
  assign n44835 = n44819 | n44834 ;
  assign n44836 = ~n44822 & n44832 ;
  assign n44837 = n44835 & n44836 ;
  assign n44838 = n44833 & ~n44837 ;
  assign n44839 = x1123 & ~n44816 ;
  assign n44840 = x1122 & ~n44816 ;
  assign n44841 = n44839 | n44840 ;
  assign n44842 = ~x826 & n44816 ;
  assign n44843 = n44841 | n44842 ;
  assign n44844 = x1123 & n44840 ;
  assign n44845 = n44843 & ~n44844 ;
  assign n44846 = x1116 | x1117 ;
  assign n44847 = x1116 & x1117 ;
  assign n44848 = n44846 & ~n44847 ;
  assign n44849 = ( x1120 & ~x1121 ) | ( x1120 & n44848 ) | ( ~x1121 & n44848 ) ;
  assign n44850 = ( ~x1120 & x1121 ) | ( ~x1120 & n44849 ) | ( x1121 & n44849 ) ;
  assign n44851 = ( ~n44848 & n44849 ) | ( ~n44848 & n44850 ) | ( n44849 & n44850 ) ;
  assign n44852 = ( x1118 & ~x1119 ) | ( x1118 & n44851 ) | ( ~x1119 & n44851 ) ;
  assign n44853 = ( ~x1118 & x1119 ) | ( ~x1118 & n44852 ) | ( x1119 & n44852 ) ;
  assign n44854 = ( ~n44851 & n44852 ) | ( ~n44851 & n44853 ) | ( n44852 & n44853 ) ;
  assign n44855 = n44845 | n44854 ;
  assign n44856 = x826 & n44816 ;
  assign n44857 = n44841 | n44856 ;
  assign n44858 = ~n44844 & n44854 ;
  assign n44859 = n44857 & n44858 ;
  assign n44860 = n44855 & ~n44859 ;
  assign n44861 = x1100 & ~n44816 ;
  assign n44862 = x1107 & ~n44816 ;
  assign n44863 = n44861 | n44862 ;
  assign n44864 = ~x827 & n44816 ;
  assign n44865 = n44863 | n44864 ;
  assign n44866 = x1100 & n44862 ;
  assign n44867 = n44865 & ~n44866 ;
  assign n44868 = x1104 | x1106 ;
  assign n44869 = x1104 & x1106 ;
  assign n44870 = n44868 & ~n44869 ;
  assign n44871 = ( x1101 & ~x1102 ) | ( x1101 & n44870 ) | ( ~x1102 & n44870 ) ;
  assign n44872 = ( ~x1101 & x1102 ) | ( ~x1101 & n44871 ) | ( x1102 & n44871 ) ;
  assign n44873 = ( ~n44870 & n44871 ) | ( ~n44870 & n44872 ) | ( n44871 & n44872 ) ;
  assign n44874 = ( x1103 & ~x1105 ) | ( x1103 & n44873 ) | ( ~x1105 & n44873 ) ;
  assign n44875 = ( ~x1103 & x1105 ) | ( ~x1103 & n44874 ) | ( x1105 & n44874 ) ;
  assign n44876 = ( ~n44873 & n44874 ) | ( ~n44873 & n44875 ) | ( n44874 & n44875 ) ;
  assign n44877 = n44867 | n44876 ;
  assign n44878 = x827 & n44816 ;
  assign n44879 = n44863 | n44878 ;
  assign n44880 = ~n44866 & n44876 ;
  assign n44881 = n44879 & n44880 ;
  assign n44882 = n44877 & ~n44881 ;
  assign n44883 = x1115 & ~n44816 ;
  assign n44884 = x1114 & ~n44816 ;
  assign n44885 = n44883 | n44884 ;
  assign n44886 = ~x828 & n44816 ;
  assign n44887 = n44885 | n44886 ;
  assign n44888 = x1115 & n44884 ;
  assign n44889 = n44887 & ~n44888 ;
  assign n44890 = x1108 | x1109 ;
  assign n44891 = x1108 & x1109 ;
  assign n44892 = n44890 & ~n44891 ;
  assign n44893 = ( x1112 & ~x1113 ) | ( x1112 & n44892 ) | ( ~x1113 & n44892 ) ;
  assign n44894 = ( ~x1112 & x1113 ) | ( ~x1112 & n44893 ) | ( x1113 & n44893 ) ;
  assign n44895 = ( ~n44892 & n44893 ) | ( ~n44892 & n44894 ) | ( n44893 & n44894 ) ;
  assign n44896 = ( x1110 & ~x1111 ) | ( x1110 & n44895 ) | ( ~x1111 & n44895 ) ;
  assign n44897 = ( ~x1110 & x1111 ) | ( ~x1110 & n44896 ) | ( x1111 & n44896 ) ;
  assign n44898 = ( ~n44895 & n44896 ) | ( ~n44895 & n44897 ) | ( n44896 & n44897 ) ;
  assign n44899 = n44889 | n44898 ;
  assign n44900 = x828 & n44816 ;
  assign n44901 = n44885 | n44900 ;
  assign n44902 = ~n44888 & n44898 ;
  assign n44903 = n44901 & n44902 ;
  assign n44904 = n44899 & ~n44903 ;
  assign n44905 = n1690 & ~n7103 ;
  assign n44906 = x951 & ~n44905 ;
  assign n44907 = x1092 & ~n44906 ;
  assign n44908 = x281 & ~n44745 ;
  assign n44909 = n44746 | n44908 ;
  assign n44910 = ~x832 & x1091 ;
  assign n44911 = x1162 & n44910 ;
  assign n44912 = n7107 & n44911 ;
  assign n44913 = x833 & ~n1290 ;
  assign n44914 = n14745 | n44913 ;
  assign n44915 = x946 & n1290 ;
  assign n44916 = x282 & ~n43235 ;
  assign n44917 = n44769 | n44916 ;
  assign n44918 = ~x955 & x1049 ;
  assign n44919 = x837 & x955 ;
  assign n44920 = n44918 | n44919 ;
  assign n44921 = ~x955 & x1047 ;
  assign n44922 = x838 & x955 ;
  assign n44923 = n44921 | n44922 ;
  assign n44924 = ~x955 & x1074 ;
  assign n44925 = x839 & x955 ;
  assign n44926 = n44924 | n44925 ;
  assign n44927 = x840 & ~n1290 ;
  assign n44928 = x1196 & n1290 ;
  assign n44929 = n44927 | n44928 ;
  assign n44930 = x33 | n7209 ;
  assign n44931 = ~x955 & x1035 ;
  assign n44932 = x842 & x955 ;
  assign n44933 = n44931 | n44932 ;
  assign n44934 = ~x955 & x1079 ;
  assign n44935 = x843 & x955 ;
  assign n44936 = n44934 | n44935 ;
  assign n44937 = ~x955 & x1078 ;
  assign n44938 = x844 & x955 ;
  assign n44939 = n44937 | n44938 ;
  assign n44940 = ~x955 & x1043 ;
  assign n44941 = x845 & x955 ;
  assign n44942 = n44940 | n44941 ;
  assign n44943 = x846 & ~n39427 ;
  assign n44944 = x1134 & n39427 ;
  assign n44945 = n44943 | n44944 ;
  assign n44946 = ~x955 & x1055 ;
  assign n44947 = x847 & x955 ;
  assign n44948 = n44946 | n44947 ;
  assign n44949 = ~x955 & x1039 ;
  assign n44950 = x848 & x955 ;
  assign n44951 = n44949 | n44950 ;
  assign n44952 = x849 & ~n1290 ;
  assign n44953 = x1198 & n1290 ;
  assign n44954 = n44952 | n44953 ;
  assign n44955 = ~x955 & x1048 ;
  assign n44956 = x850 & x955 ;
  assign n44957 = n44955 | n44956 ;
  assign n44958 = ~x955 & x1045 ;
  assign n44959 = x851 & x955 ;
  assign n44960 = n44958 | n44959 ;
  assign n44961 = ~x955 & x1062 ;
  assign n44962 = x852 & x955 ;
  assign n44963 = n44961 | n44962 ;
  assign n44964 = ~x955 & x1080 ;
  assign n44965 = x853 & x955 ;
  assign n44966 = n44964 | n44965 ;
  assign n44967 = ~x955 & x1051 ;
  assign n44968 = x854 & x955 ;
  assign n44969 = n44967 | n44968 ;
  assign n44970 = ~x955 & x1065 ;
  assign n44971 = x855 & x955 ;
  assign n44972 = n44970 | n44971 ;
  assign n44973 = ~x955 & x1067 ;
  assign n44974 = x856 & x955 ;
  assign n44975 = n44973 | n44974 ;
  assign n44976 = ~x955 & x1058 ;
  assign n44977 = x857 & x955 ;
  assign n44978 = n44976 | n44977 ;
  assign n44979 = ~x955 & x1087 ;
  assign n44980 = x858 & x955 ;
  assign n44981 = n44979 | n44980 ;
  assign n44982 = ~x955 & x1070 ;
  assign n44983 = x859 & x955 ;
  assign n44984 = n44982 | n44983 ;
  assign n44985 = ~x955 & x1076 ;
  assign n44986 = x860 & x955 ;
  assign n44987 = n44985 | n44986 ;
  assign n44988 = x1093 & x1141 ;
  assign n44989 = x861 & ~x1093 ;
  assign n44990 = n44988 | n44989 ;
  assign n44991 = ~x228 & n44990 ;
  assign n44992 = ( x123 & x228 ) | ( x123 & x1141 ) | ( x228 & x1141 ) ;
  assign n44993 = ( ~x123 & x228 ) | ( ~x123 & x861 ) | ( x228 & x861 ) ;
  assign n44994 = n44992 & n44993 ;
  assign n44995 = n44991 | n44994 ;
  assign n44996 = x862 & ~n39427 ;
  assign n44997 = x1139 & n39427 ;
  assign n44998 = n44996 | n44997 ;
  assign n44999 = x863 & ~n1290 ;
  assign n45000 = x1199 & n1290 ;
  assign n45001 = n44999 | n45000 ;
  assign n45002 = x864 & ~n1290 ;
  assign n45003 = x1197 & n1290 ;
  assign n45004 = n45002 | n45003 ;
  assign n45005 = ~x955 & x1040 ;
  assign n45006 = x865 & x955 ;
  assign n45007 = n45005 | n45006 ;
  assign n45008 = ~x955 & x1053 ;
  assign n45009 = x866 & x955 ;
  assign n45010 = n45008 | n45009 ;
  assign n45011 = ~x955 & x1057 ;
  assign n45012 = x867 & x955 ;
  assign n45013 = n45011 | n45012 ;
  assign n45014 = ~x955 & x1063 ;
  assign n45015 = x868 & x955 ;
  assign n45016 = n45014 | n45015 ;
  assign n45017 = x1093 & x1140 ;
  assign n45018 = x869 & ~x1093 ;
  assign n45019 = n45017 | n45018 ;
  assign n45020 = ~x228 & n45019 ;
  assign n45021 = ( x123 & x228 ) | ( x123 & x1140 ) | ( x228 & x1140 ) ;
  assign n45022 = ( ~x123 & x228 ) | ( ~x123 & x869 ) | ( x228 & x869 ) ;
  assign n45023 = n45021 & n45022 ;
  assign n45024 = n45020 | n45023 ;
  assign n45025 = ~x955 & x1069 ;
  assign n45026 = x870 & x955 ;
  assign n45027 = n45025 | n45026 ;
  assign n45028 = ~x955 & x1072 ;
  assign n45029 = x871 & x955 ;
  assign n45030 = n45028 | n45029 ;
  assign n45031 = ~x955 & x1084 ;
  assign n45032 = x872 & x955 ;
  assign n45033 = n45031 | n45032 ;
  assign n45034 = ~x955 & x1044 ;
  assign n45035 = x873 & x955 ;
  assign n45036 = n45034 | n45035 ;
  assign n45037 = ~x955 & x1036 ;
  assign n45038 = x874 & x955 ;
  assign n45039 = n45037 | n45038 ;
  assign n45040 = x1093 & ~x1136 ;
  assign n45041 = x875 | x1093 ;
  assign n45042 = ~n45040 & n45041 ;
  assign n45043 = x228 | n45042 ;
  assign n45044 = ( x123 & x228 ) | ( x123 & ~x1136 ) | ( x228 & ~x1136 ) ;
  assign n45045 = ( x123 & ~x228 ) | ( x123 & x875 ) | ( ~x228 & x875 ) ;
  assign n45046 = n45044 & ~n45045 ;
  assign n45047 = n45043 & ~n45046 ;
  assign n45048 = ~x955 & x1037 ;
  assign n45049 = x876 & x955 ;
  assign n45050 = n45048 | n45049 ;
  assign n45051 = x1093 & x1138 ;
  assign n45052 = x877 & ~x1093 ;
  assign n45053 = n45051 | n45052 ;
  assign n45054 = ~x228 & n45053 ;
  assign n45055 = ( x123 & x228 ) | ( x123 & x1138 ) | ( x228 & x1138 ) ;
  assign n45056 = ( ~x123 & x228 ) | ( ~x123 & x877 ) | ( x228 & x877 ) ;
  assign n45057 = n45055 & n45056 ;
  assign n45058 = n45054 | n45057 ;
  assign n45059 = x1093 & x1137 ;
  assign n45060 = x878 & ~x1093 ;
  assign n45061 = n45059 | n45060 ;
  assign n45062 = ~x228 & n45061 ;
  assign n45063 = ( x123 & x228 ) | ( x123 & x1137 ) | ( x228 & x1137 ) ;
  assign n45064 = ( ~x123 & x228 ) | ( ~x123 & x878 ) | ( x228 & x878 ) ;
  assign n45065 = n45063 & n45064 ;
  assign n45066 = n45062 | n45065 ;
  assign n45067 = x1093 & x1135 ;
  assign n45068 = x879 & ~x1093 ;
  assign n45069 = n45067 | n45068 ;
  assign n45070 = ~x228 & n45069 ;
  assign n45071 = ( x123 & x228 ) | ( x123 & x1135 ) | ( x228 & x1135 ) ;
  assign n45072 = ( ~x123 & x228 ) | ( ~x123 & x879 ) | ( x228 & x879 ) ;
  assign n45073 = n45071 & n45072 ;
  assign n45074 = n45070 | n45073 ;
  assign n45075 = ~x955 & x1081 ;
  assign n45076 = x880 & x955 ;
  assign n45077 = n45075 | n45076 ;
  assign n45078 = ~x955 & x1059 ;
  assign n45079 = x881 & x955 ;
  assign n45080 = n45078 | n45079 ;
  assign n45081 = ~x883 & n44816 ;
  assign n45082 = n44862 | n45081 ;
  assign n45083 = x1124 & ~n44816 ;
  assign n45084 = ~x884 & n44816 ;
  assign n45085 = n45083 | n45084 ;
  assign n45086 = x1125 & ~n44816 ;
  assign n45087 = ~x885 & n44816 ;
  assign n45088 = n45086 | n45087 ;
  assign n45089 = x1109 & ~n44816 ;
  assign n45090 = ~x886 & n44816 ;
  assign n45091 = n45089 | n45090 ;
  assign n45092 = ~x887 & n44816 ;
  assign n45093 = n44861 | n45092 ;
  assign n45094 = x1120 & ~n44816 ;
  assign n45095 = ~x888 & n44816 ;
  assign n45096 = n45094 | n45095 ;
  assign n45097 = x1103 & ~n44816 ;
  assign n45098 = ~x889 & n44816 ;
  assign n45099 = n45097 | n45098 ;
  assign n45100 = x1126 & ~n44816 ;
  assign n45101 = ~x890 & n44816 ;
  assign n45102 = n45100 | n45101 ;
  assign n45103 = x1116 & ~n44816 ;
  assign n45104 = ~x891 & n44816 ;
  assign n45105 = n45103 | n45104 ;
  assign n45106 = x1101 & ~n44816 ;
  assign n45107 = ~x892 & n44816 ;
  assign n45108 = n45106 | n45107 ;
  assign n45109 = x1119 & ~n44816 ;
  assign n45110 = ~x894 & n44816 ;
  assign n45111 = n45109 | n45110 ;
  assign n45112 = x1113 & ~n44816 ;
  assign n45113 = ~x895 & n44816 ;
  assign n45114 = n45112 | n45113 ;
  assign n45115 = x1118 & ~n44816 ;
  assign n45116 = ~x896 & n44816 ;
  assign n45117 = n45115 | n45116 ;
  assign n45118 = x1129 & ~n44816 ;
  assign n45119 = ~x898 & n44816 ;
  assign n45120 = n45118 | n45119 ;
  assign n45121 = ~x899 & n44816 ;
  assign n45122 = n44883 | n45121 ;
  assign n45123 = x1110 & ~n44816 ;
  assign n45124 = ~x900 & n44816 ;
  assign n45125 = n45123 | n45124 ;
  assign n45126 = x1111 & ~n44816 ;
  assign n45127 = ~x902 & n44816 ;
  assign n45128 = n45126 | n45127 ;
  assign n45129 = x1121 & ~n44816 ;
  assign n45130 = ~x903 & n44816 ;
  assign n45131 = n45129 | n45130 ;
  assign n45132 = ~x904 & n44816 ;
  assign n45133 = n44818 | n45132 ;
  assign n45134 = ~x905 & n44816 ;
  assign n45135 = n44817 | n45134 ;
  assign n45136 = x1128 & ~n44816 ;
  assign n45137 = ~x906 & n44816 ;
  assign n45138 = n45136 | n45137 ;
  assign n45139 = x782 | x907 ;
  assign n45140 = ( x598 & x782 ) | ( x598 & ~x979 ) | ( x782 & ~x979 ) ;
  assign n45141 = ( x624 & x782 ) | ( x624 & x979 ) | ( x782 & x979 ) ;
  assign n45142 = n45140 & n45141 ;
  assign n45143 = n45139 & ~n45142 ;
  assign n45144 = ( x615 & x782 ) | ( x615 & ~x979 ) | ( x782 & ~x979 ) ;
  assign n45145 = ( ~x604 & x782 ) | ( ~x604 & x979 ) | ( x782 & x979 ) ;
  assign n45146 = n45144 & n45145 ;
  assign n45147 = n45143 & ~n45146 ;
  assign n45148 = ~x908 & n44816 ;
  assign n45149 = n44840 | n45148 ;
  assign n45150 = x1105 & ~n44816 ;
  assign n45151 = ~x909 & n44816 ;
  assign n45152 = n45150 | n45151 ;
  assign n45153 = x1117 & ~n44816 ;
  assign n45154 = ~x910 & n44816 ;
  assign n45155 = n45153 | n45154 ;
  assign n45156 = x1130 & ~n44816 ;
  assign n45157 = ~x911 & n44816 ;
  assign n45158 = n45156 | n45157 ;
  assign n45159 = ~x912 & n44816 ;
  assign n45160 = n44884 | n45159 ;
  assign n45161 = x1106 & ~n44816 ;
  assign n45162 = ~x913 & n44816 ;
  assign n45163 = n45161 | n45162 ;
  assign n45164 = x280 & ~n43232 ;
  assign n45165 = n43233 | n45164 ;
  assign n45166 = x1108 & ~n44816 ;
  assign n45167 = ~x915 & n44816 ;
  assign n45168 = n45166 | n45167 ;
  assign n45169 = ~x916 & n44816 ;
  assign n45170 = n44839 | n45169 ;
  assign n45171 = x1112 & ~n44816 ;
  assign n45172 = ~x917 & n44816 ;
  assign n45173 = n45171 | n45172 ;
  assign n45174 = x1104 & ~n44816 ;
  assign n45175 = ~x918 & n44816 ;
  assign n45176 = n45174 | n45175 ;
  assign n45177 = x1102 & ~n44816 ;
  assign n45178 = ~x919 & n44816 ;
  assign n45179 = n45177 | n45178 ;
  assign n45180 = x1093 & x1139 ;
  assign n45181 = x920 & ~x1093 ;
  assign n45182 = n45180 | n45181 ;
  assign n45183 = x921 & ~x1093 ;
  assign n45184 = n45017 | n45183 ;
  assign n45185 = x922 | x1093 ;
  assign n45186 = x1093 & ~x1152 ;
  assign n45187 = n45185 & ~n45186 ;
  assign n45188 = x923 | x1093 ;
  assign n45189 = x1093 & ~x1154 ;
  assign n45190 = n45188 & ~n45189 ;
  assign n45191 = ~x300 & x301 ;
  assign n45192 = x311 & ~x312 ;
  assign n45193 = n45191 & n45192 ;
  assign n45194 = x925 | x1093 ;
  assign n45195 = x1093 & ~x1155 ;
  assign n45196 = n45194 & ~n45195 ;
  assign n45197 = x926 | x1093 ;
  assign n45198 = x1093 & ~x1157 ;
  assign n45199 = n45197 & ~n45198 ;
  assign n45200 = x927 | x1093 ;
  assign n45201 = x1093 & ~x1145 ;
  assign n45202 = n45200 & ~n45201 ;
  assign n45203 = x928 | x1093 ;
  assign n45204 = ~n45040 & n45203 ;
  assign n45205 = x929 | x1093 ;
  assign n45206 = x1093 & ~x1144 ;
  assign n45207 = n45205 & ~n45206 ;
  assign n45208 = x930 | x1093 ;
  assign n45209 = x1093 & ~x1134 ;
  assign n45210 = n45208 & ~n45209 ;
  assign n45211 = x931 | x1093 ;
  assign n45212 = x1093 & ~x1150 ;
  assign n45213 = n45211 & ~n45212 ;
  assign n45214 = x932 & ~x1093 ;
  assign n45215 = n39417 | n45214 ;
  assign n45216 = x933 & ~x1093 ;
  assign n45217 = n45059 | n45216 ;
  assign n45218 = x934 | x1093 ;
  assign n45219 = x1093 & ~x1147 ;
  assign n45220 = n45218 & ~n45219 ;
  assign n45221 = x935 & ~x1093 ;
  assign n45222 = n44988 | n45221 ;
  assign n45223 = x936 | x1093 ;
  assign n45224 = x1093 & ~x1149 ;
  assign n45225 = n45223 & ~n45224 ;
  assign n45226 = x937 | x1093 ;
  assign n45227 = x1093 & ~x1148 ;
  assign n45228 = n45226 & ~n45227 ;
  assign n45229 = x938 & ~x1093 ;
  assign n45230 = n45067 | n45229 ;
  assign n45231 = x939 | x1093 ;
  assign n45232 = x1093 & ~x1146 ;
  assign n45233 = n45231 & ~n45232 ;
  assign n45234 = x940 & ~x1093 ;
  assign n45235 = n45051 | n45234 ;
  assign n45236 = x941 | x1093 ;
  assign n45237 = x1093 & ~x1153 ;
  assign n45238 = n45236 & ~n45237 ;
  assign n45239 = x942 | x1093 ;
  assign n45240 = x1093 & ~x1156 ;
  assign n45241 = n45239 & ~n45240 ;
  assign n45242 = x943 | x1093 ;
  assign n45243 = x1093 & ~x1151 ;
  assign n45244 = n45242 & ~n45243 ;
  assign n45245 = x1093 & x1143 ;
  assign n45246 = x944 & ~x1093 ;
  assign n45247 = n45245 | n45246 ;
  assign n45248 = x230 & n1290 ;
  assign n45249 = ~x782 & x947 ;
  assign n45250 = n45142 | n45249 ;
  assign n45251 = x266 | x992 ;
  assign n45252 = ~n43232 & n45251 ;
  assign n45253 = x313 | x954 ;
  assign n45254 = x949 & x954 ;
  assign n45255 = n45253 & ~n45254 ;
  assign n45256 = ~n5995 & n12221 ;
  assign n45257 = x957 & x1092 ;
  assign n45258 = x31 | n45257 ;
  assign n45259 = ~x782 & x960 ;
  assign n45260 = ~x230 & x961 ;
  assign n45261 = ~x782 & x963 ;
  assign n45262 = ~x230 & x967 ;
  assign n45263 = ~x230 & x969 ;
  assign n45264 = ~x782 & x970 ;
  assign n45265 = ~x230 & x971 ;
  assign n45266 = ~x782 & x972 ;
  assign n45267 = ~x230 & x974 ;
  assign n45268 = ~x782 & x975 ;
  assign n45269 = ~x230 & x977 ;
  assign n45270 = ~x782 & x978 ;
  assign n45271 = ~x598 & x615 ;
  assign n45272 = x824 & x1092 ;
  assign n45273 = x604 | x624 ;
  assign y0 = x668 ;
  assign y1 = x672 ;
  assign y2 = x664 ;
  assign y3 = x667 ;
  assign y4 = x676 ;
  assign y5 = x673 ;
  assign y6 = x675 ;
  assign y7 = x666 ;
  assign y8 = x679 ;
  assign y9 = x674 ;
  assign y10 = x663 ;
  assign y11 = x670 ;
  assign y12 = x677 ;
  assign y13 = x682 ;
  assign y14 = x671 ;
  assign y15 = x678 ;
  assign y16 = x718 ;
  assign y17 = x707 ;
  assign y18 = x708 ;
  assign y19 = x713 ;
  assign y20 = x711 ;
  assign y21 = x716 ;
  assign y22 = x733 ;
  assign y23 = x712 ;
  assign y24 = x689 ;
  assign y25 = x717 ;
  assign y26 = x692 ;
  assign y27 = x719 ;
  assign y28 = x722 ;
  assign y29 = x714 ;
  assign y30 = x720 ;
  assign y31 = x685 ;
  assign y32 = x837 ;
  assign y33 = x850 ;
  assign y34 = x872 ;
  assign y35 = x871 ;
  assign y36 = x881 ;
  assign y37 = x866 ;
  assign y38 = x876 ;
  assign y39 = x873 ;
  assign y40 = x874 ;
  assign y41 = x859 ;
  assign y42 = x855 ;
  assign y43 = x852 ;
  assign y44 = x870 ;
  assign y45 = x848 ;
  assign y46 = x865 ;
  assign y47 = x856 ;
  assign y48 = x853 ;
  assign y49 = x847 ;
  assign y50 = x857 ;
  assign y51 = x854 ;
  assign y52 = x858 ;
  assign y53 = x845 ;
  assign y54 = x838 ;
  assign y55 = x842 ;
  assign y56 = x843 ;
  assign y57 = x839 ;
  assign y58 = x844 ;
  assign y59 = x868 ;
  assign y60 = x851 ;
  assign y61 = x867 ;
  assign y62 = x880 ;
  assign y63 = x860 ;
  assign y64 = x1030 ;
  assign y65 = x1034 ;
  assign y66 = x1015 ;
  assign y67 = x1020 ;
  assign y68 = x1025 ;
  assign y69 = x1005 ;
  assign y70 = x996 ;
  assign y71 = x1012 ;
  assign y72 = x993 ;
  assign y73 = x1016 ;
  assign y74 = x1021 ;
  assign y75 = x1010 ;
  assign y76 = x1027 ;
  assign y77 = x1018 ;
  assign y78 = x1017 ;
  assign y79 = x1024 ;
  assign y80 = x1009 ;
  assign y81 = x1032 ;
  assign y82 = x1003 ;
  assign y83 = x997 ;
  assign y84 = x1013 ;
  assign y85 = x1011 ;
  assign y86 = x1008 ;
  assign y87 = x1019 ;
  assign y88 = x1031 ;
  assign y89 = x1022 ;
  assign y90 = x1000 ;
  assign y91 = x1023 ;
  assign y92 = x1002 ;
  assign y93 = x1026 ;
  assign y94 = x1006 ;
  assign y95 = x998 ;
  assign y96 = x31 ;
  assign y97 = x80 ;
  assign y98 = x893 ;
  assign y99 = x467 ;
  assign y100 = x78 ;
  assign y101 = x112 ;
  assign y102 = x13 ;
  assign y103 = x25 ;
  assign y104 = x226 ;
  assign y105 = x127 ;
  assign y106 = x822 ;
  assign y107 = x808 ;
  assign y108 = x227 ;
  assign y109 = x477 ;
  assign y110 = x834 ;
  assign y111 = x229 ;
  assign y112 = x12 ;
  assign y113 = x11 ;
  assign y114 = x10 ;
  assign y115 = x9 ;
  assign y116 = x8 ;
  assign y117 = x7 ;
  assign y118 = x6 ;
  assign y119 = x5 ;
  assign y120 = x4 ;
  assign y121 = x3 ;
  assign y122 = x0 ;
  assign y123 = x2 ;
  assign y124 = x1 ;
  assign y125 = x310 ;
  assign y126 = x302 ;
  assign y127 = x475 ;
  assign y128 = x474 ;
  assign y129 = x466 ;
  assign y130 = x473 ;
  assign y131 = x471 ;
  assign y132 = x472 ;
  assign y133 = x470 ;
  assign y134 = x469 ;
  assign y135 = x465 ;
  assign y136 = x1028 ;
  assign y137 = x1033 ;
  assign y138 = x995 ;
  assign y139 = x994 ;
  assign y140 = x28 ;
  assign y141 = x27 ;
  assign y142 = x26 ;
  assign y143 = x29 ;
  assign y144 = x15 ;
  assign y145 = x14 ;
  assign y146 = x21 ;
  assign y147 = x20 ;
  assign y148 = x19 ;
  assign y149 = x18 ;
  assign y150 = x17 ;
  assign y151 = x16 ;
  assign y152 = x1096 ;
  assign y153 = n2067 ;
  assign y154 = n2292 ;
  assign y155 = n2453 ;
  assign y156 = ~n2665 ;
  assign y157 = ~n2874 ;
  assign y158 = n3077 ;
  assign y159 = n3280 ;
  assign y160 = n3490 ;
  assign y161 = n3692 ;
  assign y162 = n3894 ;
  assign y163 = n4107 ;
  assign y164 = n4320 ;
  assign y165 = n4647 ;
  assign y166 = ~1'b0 ;
  assign y167 = n4830 ;
  assign y168 = x228 ;
  assign y169 = x22 ;
  assign y170 = ~x1090 ;
  assign y171 = ~n5092 ;
  assign y172 = ~n5207 ;
  assign y173 = ~n5326 ;
  assign y174 = ~n5413 ;
  assign y175 = ~n5500 ;
  assign y176 = ~n5587 ;
  assign y177 = ~n5674 ;
  assign y178 = ~n5757 ;
  assign y179 = x1089 ;
  assign y180 = x23 ;
  assign y181 = n4830 ;
  assign y182 = n5810 ;
  assign y183 = n5859 ;
  assign y184 = ~n5864 ;
  assign y185 = ~n5866 ;
  assign y186 = ~n5868 ;
  assign y187 = ~n5870 ;
  assign y188 = x37 ;
  assign y189 = n7110 ;
  assign y190 = n7203 ;
  assign y191 = n7892 ;
  assign y192 = n8237 ;
  assign y193 = n8312 ;
  assign y194 = n8334 ;
  assign y195 = n5807 ;
  assign y196 = n8365 ;
  assign y197 = n8447 ;
  assign y198 = n8465 ;
  assign y199 = n8651 ;
  assign y200 = n8893 ;
  assign y201 = n9067 ;
  assign y202 = n9137 ;
  assign y203 = n9141 ;
  assign y204 = n9161 ;
  assign y205 = n9208 ;
  assign y206 = n9214 ;
  assign y207 = n9232 ;
  assign y208 = n9258 ;
  assign y209 = n9266 ;
  assign y210 = n9404 ;
  assign y211 = n9416 ;
  assign y212 = n9435 ;
  assign y213 = n9449 ;
  assign y214 = n9457 ;
  assign y215 = n9466 ;
  assign y216 = n9469 ;
  assign y217 = n9473 ;
  assign y218 = n9481 ;
  assign y219 = n9486 ;
  assign y220 = n9489 ;
  assign y221 = n9495 ;
  assign y222 = n9504 ;
  assign y223 = n9508 ;
  assign y224 = n9524 ;
  assign y225 = n9529 ;
  assign y226 = n9537 ;
  assign y227 = n9550 ;
  assign y228 = n9570 ;
  assign y229 = n9591 ;
  assign y230 = n9608 ;
  assign y231 = n9619 ;
  assign y232 = n9634 ;
  assign y233 = n9643 ;
  assign y234 = n9787 ;
  assign y235 = n9796 ;
  assign y236 = n9798 ;
  assign y237 = n10285 ;
  assign y238 = n11069 ;
  assign y239 = n11079 ;
  assign y240 = n11089 ;
  assign y241 = n11102 ;
  assign y242 = n11108 ;
  assign y243 = n11113 ;
  assign y244 = n11117 ;
  assign y245 = n11121 ;
  assign y246 = n11139 ;
  assign y247 = n11149 ;
  assign y248 = n11154 ;
  assign y249 = n11166 ;
  assign y250 = n11178 ;
  assign y251 = n11184 ;
  assign y252 = n11199 ;
  assign y253 = n11215 ;
  assign y254 = n11226 ;
  assign y255 = n11236 ;
  assign y256 = n11241 ;
  assign y257 = n11313 ;
  assign y258 = n11329 ;
  assign y259 = n11403 ;
  assign y260 = n11405 ;
  assign y261 = n11412 ;
  assign y262 = n11429 ;
  assign y263 = x117 ;
  assign y264 = n11439 ;
  assign y265 = n11441 ;
  assign y266 = n11458 ;
  assign y267 = n11460 ;
  assign y268 = n11470 ;
  assign y269 = n11476 ;
  assign y270 = ~n11477 ;
  assign y271 = n11525 ;
  assign y272 = n11567 ;
  assign y273 = n11608 ;
  assign y274 = n11658 ;
  assign y275 = n11673 ;
  assign y276 = n11956 ;
  assign y277 = n12009 ;
  assign y278 = n12390 ;
  assign y279 = n12791 ;
  assign y280 = n12798 ;
  assign y281 = ~n12850 ;
  assign y282 = n13232 ;
  assign y283 = n13508 ;
  assign y284 = n13595 ;
  assign y285 = x131 ;
  assign y286 = n13619 ;
  assign y287 = n13743 ;
  assign y288 = n13751 ;
  assign y289 = n13950 ;
  assign y290 = n14006 ;
  assign y291 = n14116 ;
  assign y292 = n14227 ;
  assign y293 = n14309 ;
  assign y294 = n14322 ;
  assign y295 = n14400 ;
  assign y296 = n14449 ;
  assign y297 = ~n16238 ;
  assign y298 = ~n16700 ;
  assign y299 = n17407 ;
  assign y300 = ~n17872 ;
  assign y301 = n18477 ;
  assign y302 = ~n18908 ;
  assign y303 = n18985 ;
  assign y304 = ~n19133 ;
  assign y305 = ~n19195 ;
  assign y306 = ~n19249 ;
  assign y307 = ~n19299 ;
  assign y308 = ~n19374 ;
  assign y309 = n19475 ;
  assign y310 = ~n19556 ;
  assign y311 = ~n19604 ;
  assign y312 = ~n19641 ;
  assign y313 = ~n19668 ;
  assign y314 = ~n19720 ;
  assign y315 = ~n19770 ;
  assign y316 = ~n19820 ;
  assign y317 = ~n19873 ;
  assign y318 = n19964 ;
  assign y319 = ~n20014 ;
  assign y320 = ~n20067 ;
  assign y321 = ~n20103 ;
  assign y322 = ~n20139 ;
  assign y323 = n20232 ;
  assign y324 = ~n20271 ;
  assign y325 = ~n20352 ;
  assign y326 = ~n20433 ;
  assign y327 = ~n20513 ;
  assign y328 = ~n20594 ;
  assign y329 = ~n20674 ;
  assign y330 = ~n21098 ;
  assign y331 = n21743 ;
  assign y332 = ~n22178 ;
  assign y333 = ~n22585 ;
  assign y334 = ~n23017 ;
  assign y335 = ~n23444 ;
  assign y336 = ~n23876 ;
  assign y337 = ~n24309 ;
  assign y338 = ~n24742 ;
  assign y339 = ~n25169 ;
  assign y340 = ~n25596 ;
  assign y341 = ~n26023 ;
  assign y342 = ~n26456 ;
  assign y343 = ~n26881 ;
  assign y344 = ~n27306 ;
  assign y345 = ~n27731 ;
  assign y346 = n28157 ;
  assign y347 = ~n28591 ;
  assign y348 = ~n29025 ;
  assign y349 = ~n29459 ;
  assign y350 = ~n29887 ;
  assign y351 = ~n30304 ;
  assign y352 = n30351 ;
  assign y353 = n30414 ;
  assign y354 = ~n30469 ;
  assign y355 = n31060 ;
  assign y356 = n31314 ;
  assign y357 = n31562 ;
  assign y358 = ~n31742 ;
  assign y359 = ~n31749 ;
  assign y360 = ~n31756 ;
  assign y361 = ~n31858 ;
  assign y362 = ~n31864 ;
  assign y363 = ~n31871 ;
  assign y364 = ~n32325 ;
  assign y365 = ~n32388 ;
  assign y366 = ~n32536 ;
  assign y367 = n32654 ;
  assign y368 = n32678 ;
  assign y369 = ~n32696 ;
  assign y370 = ~n32714 ;
  assign y371 = ~n32732 ;
  assign y372 = n32844 ;
  assign y373 = n32946 ;
  assign y374 = ~n32962 ;
  assign y375 = ~n32968 ;
  assign y376 = n32986 ;
  assign y377 = ~n32992 ;
  assign y378 = n33097 ;
  assign y379 = n33677 ;
  assign y380 = n34213 ;
  assign y381 = n34752 ;
  assign y382 = n34869 ;
  assign y383 = n34918 ;
  assign y384 = ~n34948 ;
  assign y385 = n34959 ;
  assign y386 = x232 ;
  assign y387 = n35040 ;
  assign y388 = x236 ;
  assign y389 = n35098 ;
  assign y390 = ~n35503 ;
  assign y391 = n35824 ;
  assign y392 = n36013 ;
  assign y393 = n36025 ;
  assign y394 = ~n36275 ;
  assign y395 = n36608 ;
  assign y396 = n36695 ;
  assign y397 = n37099 ;
  assign y398 = n37379 ;
  assign y399 = n37463 ;
  assign y400 = ~n37764 ;
  assign y401 = n37814 ;
  assign y402 = n38055 ;
  assign y403 = n38310 ;
  assign y404 = n38535 ;
  assign y405 = n38692 ;
  assign y406 = n38869 ;
  assign y407 = n38877 ;
  assign y408 = n38886 ;
  assign y409 = n38926 ;
  assign y410 = n39156 ;
  assign y411 = n39374 ;
  assign y412 = n39380 ;
  assign y413 = n39386 ;
  assign y414 = n39392 ;
  assign y415 = n39398 ;
  assign y416 = n39404 ;
  assign y417 = n39410 ;
  assign y418 = n39416 ;
  assign y419 = ~n39448 ;
  assign y420 = ~n39647 ;
  assign y421 = ~n39686 ;
  assign y422 = ~n39722 ;
  assign y423 = n39785 ;
  assign y424 = n39982 ;
  assign y425 = n40128 ;
  assign y426 = ~n40170 ;
  assign y427 = ~n40210 ;
  assign y428 = n40258 ;
  assign y429 = n40353 ;
  assign y430 = n40416 ;
  assign y431 = ~n40452 ;
  assign y432 = n40524 ;
  assign y433 = n40551 ;
  assign y434 = ~n40588 ;
  assign y435 = n40655 ;
  assign y436 = n40709 ;
  assign y437 = ~n40750 ;
  assign y438 = ~n40786 ;
  assign y439 = ~n40821 ;
  assign y440 = n40872 ;
  assign y441 = ~n40876 ;
  assign y442 = n40893 ;
  assign y443 = n40909 ;
  assign y444 = ~n40911 ;
  assign y445 = n40917 ;
  assign y446 = n40929 ;
  assign y447 = n40932 ;
  assign y448 = n40935 ;
  assign y449 = n40938 ;
  assign y450 = n40941 ;
  assign y451 = n40944 ;
  assign y452 = n40947 ;
  assign y453 = n40950 ;
  assign y454 = n40953 ;
  assign y455 = n40956 ;
  assign y456 = n40964 ;
  assign y457 = n40971 ;
  assign y458 = ~n40975 ;
  assign y459 = ~n40997 ;
  assign y460 = n41000 ;
  assign y461 = n41003 ;
  assign y462 = n41006 ;
  assign y463 = n41009 ;
  assign y464 = n41012 ;
  assign y465 = n41015 ;
  assign y466 = n41018 ;
  assign y467 = ~n41045 ;
  assign y468 = ~n41049 ;
  assign y469 = n41052 ;
  assign y470 = n41059 ;
  assign y471 = ~n41070 ;
  assign y472 = n41075 ;
  assign y473 = n41078 ;
  assign y474 = n41082 ;
  assign y475 = n41087 ;
  assign y476 = n41090 ;
  assign y477 = n41093 ;
  assign y478 = n41096 ;
  assign y479 = n41099 ;
  assign y480 = n41102 ;
  assign y481 = n41105 ;
  assign y482 = n41108 ;
  assign y483 = n41111 ;
  assign y484 = n41114 ;
  assign y485 = n41117 ;
  assign y486 = n41120 ;
  assign y487 = n41128 ;
  assign y488 = n41133 ;
  assign y489 = n41143 ;
  assign y490 = n41146 ;
  assign y491 = n41149 ;
  assign y492 = n41152 ;
  assign y493 = n41155 ;
  assign y494 = n41158 ;
  assign y495 = n41161 ;
  assign y496 = n41164 ;
  assign y497 = ~n41170 ;
  assign y498 = n41173 ;
  assign y499 = n41176 ;
  assign y500 = n41179 ;
  assign y501 = n41182 ;
  assign y502 = n41185 ;
  assign y503 = n41188 ;
  assign y504 = n41191 ;
  assign y505 = n41194 ;
  assign y506 = n41197 ;
  assign y507 = n41200 ;
  assign y508 = n41203 ;
  assign y509 = n41206 ;
  assign y510 = n41209 ;
  assign y511 = n41212 ;
  assign y512 = n41215 ;
  assign y513 = n41218 ;
  assign y514 = n41221 ;
  assign y515 = n41224 ;
  assign y516 = n41227 ;
  assign y517 = n41230 ;
  assign y518 = n41233 ;
  assign y519 = n41236 ;
  assign y520 = n41239 ;
  assign y521 = n41242 ;
  assign y522 = n41245 ;
  assign y523 = n41248 ;
  assign y524 = n41251 ;
  assign y525 = n41254 ;
  assign y526 = n41257 ;
  assign y527 = n41260 ;
  assign y528 = n41263 ;
  assign y529 = n41266 ;
  assign y530 = n41269 ;
  assign y531 = n41272 ;
  assign y532 = n41275 ;
  assign y533 = n41278 ;
  assign y534 = n41281 ;
  assign y535 = n41284 ;
  assign y536 = n41287 ;
  assign y537 = n41290 ;
  assign y538 = n41293 ;
  assign y539 = n41296 ;
  assign y540 = n41299 ;
  assign y541 = n41302 ;
  assign y542 = n41305 ;
  assign y543 = n41308 ;
  assign y544 = n41311 ;
  assign y545 = n41314 ;
  assign y546 = n41317 ;
  assign y547 = n41320 ;
  assign y548 = n41323 ;
  assign y549 = n41326 ;
  assign y550 = n41329 ;
  assign y551 = n41332 ;
  assign y552 = n41335 ;
  assign y553 = n41338 ;
  assign y554 = n41341 ;
  assign y555 = n41344 ;
  assign y556 = n41347 ;
  assign y557 = n41350 ;
  assign y558 = n41353 ;
  assign y559 = n41356 ;
  assign y560 = n41359 ;
  assign y561 = n41362 ;
  assign y562 = n41365 ;
  assign y563 = n41368 ;
  assign y564 = n41371 ;
  assign y565 = n41374 ;
  assign y566 = n41377 ;
  assign y567 = n41380 ;
  assign y568 = n41383 ;
  assign y569 = n41386 ;
  assign y570 = n41389 ;
  assign y571 = n41393 ;
  assign y572 = n41396 ;
  assign y573 = n41399 ;
  assign y574 = n41402 ;
  assign y575 = n41405 ;
  assign y576 = n41408 ;
  assign y577 = n41411 ;
  assign y578 = n41414 ;
  assign y579 = n41417 ;
  assign y580 = n41420 ;
  assign y581 = n41423 ;
  assign y582 = n41426 ;
  assign y583 = n41429 ;
  assign y584 = n41432 ;
  assign y585 = n41435 ;
  assign y586 = n41438 ;
  assign y587 = n41441 ;
  assign y588 = n41444 ;
  assign y589 = n41447 ;
  assign y590 = n41450 ;
  assign y591 = n41453 ;
  assign y592 = n41456 ;
  assign y593 = n41459 ;
  assign y594 = n41462 ;
  assign y595 = n41465 ;
  assign y596 = n41468 ;
  assign y597 = n41471 ;
  assign y598 = n41474 ;
  assign y599 = n41477 ;
  assign y600 = n41480 ;
  assign y601 = n41483 ;
  assign y602 = n41486 ;
  assign y603 = n41489 ;
  assign y604 = n41492 ;
  assign y605 = n41495 ;
  assign y606 = n41498 ;
  assign y607 = n41501 ;
  assign y608 = n41504 ;
  assign y609 = n41507 ;
  assign y610 = n41510 ;
  assign y611 = n41513 ;
  assign y612 = n41516 ;
  assign y613 = n41519 ;
  assign y614 = n41543 ;
  assign y615 = n41546 ;
  assign y616 = n41549 ;
  assign y617 = n41552 ;
  assign y618 = n41555 ;
  assign y619 = n41558 ;
  assign y620 = n41561 ;
  assign y621 = n41564 ;
  assign y622 = n41588 ;
  assign y623 = n41606 ;
  assign y624 = n41634 ;
  assign y625 = n41639 ;
  assign y626 = n41658 ;
  assign y627 = n41677 ;
  assign y628 = n41696 ;
  assign y629 = n41714 ;
  assign y630 = n41725 ;
  assign y631 = n41736 ;
  assign y632 = n41747 ;
  assign y633 = n41759 ;
  assign y634 = ~n41056 ;
  assign y635 = n41760 ;
  assign y636 = x583 ;
  assign y637 = n40912 ;
  assign y638 = n41763 ;
  assign y639 = n41766 ;
  assign y640 = n41769 ;
  assign y641 = n41772 ;
  assign y642 = n41775 ;
  assign y643 = n41778 ;
  assign y644 = n41781 ;
  assign y645 = ~n41784 ;
  assign y646 = n41787 ;
  assign y647 = n41790 ;
  assign y648 = n41793 ;
  assign y649 = n41796 ;
  assign y650 = n41799 ;
  assign y651 = ~n41802 ;
  assign y652 = n41805 ;
  assign y653 = n41808 ;
  assign y654 = ~n41811 ;
  assign y655 = n41814 ;
  assign y656 = n41817 ;
  assign y657 = n41820 ;
  assign y658 = n41823 ;
  assign y659 = n41826 ;
  assign y660 = n41829 ;
  assign y661 = n41832 ;
  assign y662 = n41840 ;
  assign y663 = n41843 ;
  assign y664 = n41846 ;
  assign y665 = n41849 ;
  assign y666 = n41852 ;
  assign y667 = n41855 ;
  assign y668 = n41861 ;
  assign y669 = n41864 ;
  assign y670 = n41867 ;
  assign y671 = n41870 ;
  assign y672 = n41873 ;
  assign y673 = n41876 ;
  assign y674 = n41879 ;
  assign y675 = n41885 ;
  assign y676 = ~n41888 ;
  assign y677 = n41891 ;
  assign y678 = n41894 ;
  assign y679 = n41897 ;
  assign y680 = n41902 ;
  assign y681 = ~n41905 ;
  assign y682 = n41908 ;
  assign y683 = n41911 ;
  assign y684 = n41914 ;
  assign y685 = n41917 ;
  assign y686 = n41920 ;
  assign y687 = n41923 ;
  assign y688 = n41926 ;
  assign y689 = n41929 ;
  assign y690 = n41932 ;
  assign y691 = ~n41935 ;
  assign y692 = n41938 ;
  assign y693 = n41941 ;
  assign y694 = n41944 ;
  assign y695 = n41947 ;
  assign y696 = n41950 ;
  assign y697 = n41953 ;
  assign y698 = n41956 ;
  assign y699 = n41959 ;
  assign y700 = n41962 ;
  assign y701 = n41967 ;
  assign y702 = n41970 ;
  assign y703 = n41973 ;
  assign y704 = n41976 ;
  assign y705 = n41979 ;
  assign y706 = n41982 ;
  assign y707 = ~n41985 ;
  assign y708 = n41988 ;
  assign y709 = n41991 ;
  assign y710 = n41994 ;
  assign y711 = n41997 ;
  assign y712 = n42000 ;
  assign y713 = n42003 ;
  assign y714 = n42008 ;
  assign y715 = n42011 ;
  assign y716 = n42014 ;
  assign y717 = n42017 ;
  assign y718 = n42020 ;
  assign y719 = n42023 ;
  assign y720 = n42026 ;
  assign y721 = n42029 ;
  assign y722 = n42032 ;
  assign y723 = n42035 ;
  assign y724 = n42139 ;
  assign y725 = n42142 ;
  assign y726 = ~n42145 ;
  assign y727 = n42150 ;
  assign y728 = n42153 ;
  assign y729 = n42156 ;
  assign y730 = n42159 ;
  assign y731 = n42162 ;
  assign y732 = n42165 ;
  assign y733 = n42168 ;
  assign y734 = n42171 ;
  assign y735 = n42174 ;
  assign y736 = n42177 ;
  assign y737 = n42180 ;
  assign y738 = n42183 ;
  assign y739 = n42186 ;
  assign y740 = n4800 ;
  assign y741 = n42189 ;
  assign y742 = n42192 ;
  assign y743 = n42195 ;
  assign y744 = n42202 ;
  assign y745 = n42206 ;
  assign y746 = n42227 ;
  assign y747 = ~n42230 ;
  assign y748 = n42233 ;
  assign y749 = n42236 ;
  assign y750 = n42985 ;
  assign y751 = n42992 ;
  assign y752 = n42997 ;
  assign y753 = n43003 ;
  assign y754 = n43006 ;
  assign y755 = n43012 ;
  assign y756 = n43016 ;
  assign y757 = n43019 ;
  assign y758 = n43022 ;
  assign y759 = n43032 ;
  assign y760 = n43046 ;
  assign y761 = n43053 ;
  assign y762 = ~n43056 ;
  assign y763 = n43061 ;
  assign y764 = n43064 ;
  assign y765 = n43067 ;
  assign y766 = n43070 ;
  assign y767 = n43073 ;
  assign y768 = n43076 ;
  assign y769 = n43079 ;
  assign y770 = n43082 ;
  assign y771 = n43086 ;
  assign y772 = ~n43091 ;
  assign y773 = n43095 ;
  assign y774 = n43100 ;
  assign y775 = n43103 ;
  assign y776 = n43106 ;
  assign y777 = n43109 ;
  assign y778 = n43112 ;
  assign y779 = n43115 ;
  assign y780 = n43118 ;
  assign y781 = n43124 ;
  assign y782 = n43132 ;
  assign y783 = n43135 ;
  assign y784 = n43138 ;
  assign y785 = n43141 ;
  assign y786 = n43144 ;
  assign y787 = n43147 ;
  assign y788 = ~n43150 ;
  assign y789 = ~n43153 ;
  assign y790 = n43156 ;
  assign y791 = n43159 ;
  assign y792 = ~n43162 ;
  assign y793 = n43165 ;
  assign y794 = n43168 ;
  assign y795 = n43171 ;
  assign y796 = n43174 ;
  assign y797 = n43177 ;
  assign y798 = n43180 ;
  assign y799 = n43183 ;
  assign y800 = n43186 ;
  assign y801 = n43189 ;
  assign y802 = n43192 ;
  assign y803 = ~n43195 ;
  assign y804 = n43198 ;
  assign y805 = n43201 ;
  assign y806 = ~n43204 ;
  assign y807 = ~n43207 ;
  assign y808 = n43210 ;
  assign y809 = n43213 ;
  assign y810 = n43216 ;
  assign y811 = ~n43219 ;
  assign y812 = ~n43222 ;
  assign y813 = n43225 ;
  assign y814 = ~n43228 ;
  assign y815 = n43231 ;
  assign y816 = ~n43243 ;
  assign y817 = n43246 ;
  assign y818 = n43249 ;
  assign y819 = n43252 ;
  assign y820 = n43298 ;
  assign y821 = n43334 ;
  assign y822 = n43337 ;
  assign y823 = n43369 ;
  assign y824 = n43401 ;
  assign y825 = n43433 ;
  assign y826 = ~n43436 ;
  assign y827 = n43467 ;
  assign y828 = n43497 ;
  assign y829 = n43529 ;
  assign y830 = n43561 ;
  assign y831 = n43595 ;
  assign y832 = n43628 ;
  assign y833 = n43660 ;
  assign y834 = n43690 ;
  assign y835 = n43720 ;
  assign y836 = n43754 ;
  assign y837 = n43757 ;
  assign y838 = n43760 ;
  assign y839 = n43790 ;
  assign y840 = n7136 ;
  assign y841 = ~n43794 ;
  assign y842 = n43831 ;
  assign y843 = ~n43834 ;
  assign y844 = n43837 ;
  assign y845 = ~n43840 ;
  assign y846 = n43872 ;
  assign y847 = n43875 ;
  assign y848 = n43878 ;
  assign y849 = n43910 ;
  assign y850 = ~n43913 ;
  assign y851 = ~n43916 ;
  assign y852 = ~n43919 ;
  assign y853 = n43922 ;
  assign y854 = ~n43925 ;
  assign y855 = ~n43928 ;
  assign y856 = n43931 ;
  assign y857 = n43934 ;
  assign y858 = ~n43937 ;
  assign y859 = ~n43940 ;
  assign y860 = n43943 ;
  assign y861 = ~n43946 ;
  assign y862 = n43949 ;
  assign y863 = n43952 ;
  assign y864 = n43986 ;
  assign y865 = n44024 ;
  assign y866 = ~n44027 ;
  assign y867 = n44030 ;
  assign y868 = n44062 ;
  assign y869 = n44096 ;
  assign y870 = n44128 ;
  assign y871 = n44161 ;
  assign y872 = n44164 ;
  assign y873 = n44198 ;
  assign y874 = n44230 ;
  assign y875 = n44264 ;
  assign y876 = n44296 ;
  assign y877 = n44329 ;
  assign y878 = n44383 ;
  assign y879 = n44413 ;
  assign y880 = ~n44416 ;
  assign y881 = ~n44419 ;
  assign y882 = ~n44422 ;
  assign y883 = n44425 ;
  assign y884 = n44428 ;
  assign y885 = ~n44431 ;
  assign y886 = n44434 ;
  assign y887 = n44437 ;
  assign y888 = n44453 ;
  assign y889 = ~n44456 ;
  assign y890 = n44490 ;
  assign y891 = ~n44493 ;
  assign y892 = n44496 ;
  assign y893 = n44499 ;
  assign y894 = ~n44502 ;
  assign y895 = ~n44505 ;
  assign y896 = n44511 ;
  assign y897 = n43037 ;
  assign y898 = ~n44514 ;
  assign y899 = ~n44517 ;
  assign y900 = n44520 ;
  assign y901 = ~n44523 ;
  assign y902 = ~n44526 ;
  assign y903 = n44529 ;
  assign y904 = n44541 ;
  assign y905 = n44544 ;
  assign y906 = n44547 ;
  assign y907 = ~n44550 ;
  assign y908 = ~n44553 ;
  assign y909 = ~n44556 ;
  assign y910 = ~n44559 ;
  assign y911 = ~n44562 ;
  assign y912 = ~n44565 ;
  assign y913 = ~n44568 ;
  assign y914 = ~n44571 ;
  assign y915 = n44574 ;
  assign y916 = n44578 ;
  assign y917 = ~n44581 ;
  assign y918 = ~n44584 ;
  assign y919 = ~n44587 ;
  assign y920 = n44590 ;
  assign y921 = n44593 ;
  assign y922 = ~n44616 ;
  assign y923 = n44619 ;
  assign y924 = ~n44622 ;
  assign y925 = ~n44625 ;
  assign y926 = n44640 ;
  assign y927 = ~n44643 ;
  assign y928 = n44653 ;
  assign y929 = n44656 ;
  assign y930 = n44664 ;
  assign y931 = ~n44667 ;
  assign y932 = n44683 ;
  assign y933 = ~n44686 ;
  assign y934 = ~n44689 ;
  assign y935 = n44697 ;
  assign y936 = ~n44698 ;
  assign y937 = ~n44699 ;
  assign y938 = n44702 ;
  assign y939 = ~n44704 ;
  assign y940 = n44707 ;
  assign y941 = n44710 ;
  assign y942 = n44713 ;
  assign y943 = ~n44716 ;
  assign y944 = n44719 ;
  assign y945 = n44722 ;
  assign y946 = n44725 ;
  assign y947 = n44728 ;
  assign y948 = n44731 ;
  assign y949 = n44734 ;
  assign y950 = ~n35076 ;
  assign y951 = n44738 ;
  assign y952 = n44741 ;
  assign y953 = ~n44750 ;
  assign y954 = n43129 ;
  assign y955 = n44753 ;
  assign y956 = ~n44756 ;
  assign y957 = n44759 ;
  assign y958 = n44762 ;
  assign y959 = n43241 ;
  assign y960 = ~n44765 ;
  assign y961 = n44768 ;
  assign y962 = ~n44772 ;
  assign y963 = n44648 ;
  assign y964 = n44775 ;
  assign y965 = n44778 ;
  assign y966 = ~n44781 ;
  assign y967 = n44784 ;
  assign y968 = n44787 ;
  assign y969 = ~n44790 ;
  assign y970 = n44793 ;
  assign y971 = ~n44796 ;
  assign y972 = n44799 ;
  assign y973 = n44802 ;
  assign y974 = ~n44804 ;
  assign y975 = n44806 ;
  assign y976 = ~n44808 ;
  assign y977 = ~n44810 ;
  assign y978 = ~n44594 ;
  assign y979 = ~n44811 ;
  assign y980 = n43791 ;
  assign y981 = n44815 ;
  assign y982 = n44838 ;
  assign y983 = n44860 ;
  assign y984 = n44882 ;
  assign y985 = n44904 ;
  assign y986 = n44907 ;
  assign y987 = ~n44909 ;
  assign y988 = n44508 ;
  assign y989 = n44912 ;
  assign y990 = n44914 ;
  assign y991 = n44915 ;
  assign y992 = ~n44917 ;
  assign y993 = n44920 ;
  assign y994 = n44923 ;
  assign y995 = n44926 ;
  assign y996 = n44929 ;
  assign y997 = ~n44930 ;
  assign y998 = n44933 ;
  assign y999 = n44936 ;
  assign y1000 = n44939 ;
  assign y1001 = n44942 ;
  assign y1002 = n44945 ;
  assign y1003 = n44948 ;
  assign y1004 = n44951 ;
  assign y1005 = n44954 ;
  assign y1006 = n44957 ;
  assign y1007 = n44960 ;
  assign y1008 = n44963 ;
  assign y1009 = n44966 ;
  assign y1010 = n44969 ;
  assign y1011 = n44972 ;
  assign y1012 = n44975 ;
  assign y1013 = n44978 ;
  assign y1014 = n44981 ;
  assign y1015 = n44984 ;
  assign y1016 = n44987 ;
  assign y1017 = n44995 ;
  assign y1018 = n44998 ;
  assign y1019 = n45001 ;
  assign y1020 = n45004 ;
  assign y1021 = n45007 ;
  assign y1022 = n45010 ;
  assign y1023 = n45013 ;
  assign y1024 = n45016 ;
  assign y1025 = n45024 ;
  assign y1026 = n45027 ;
  assign y1027 = n45030 ;
  assign y1028 = n45033 ;
  assign y1029 = n45036 ;
  assign y1030 = n45039 ;
  assign y1031 = n45047 ;
  assign y1032 = n45050 ;
  assign y1033 = n45058 ;
  assign y1034 = n45066 ;
  assign y1035 = n45074 ;
  assign y1036 = n45077 ;
  assign y1037 = n45080 ;
  assign y1038 = n6785 ;
  assign y1039 = n45082 ;
  assign y1040 = n45085 ;
  assign y1041 = n45088 ;
  assign y1042 = n45091 ;
  assign y1043 = n45093 ;
  assign y1044 = n45096 ;
  assign y1045 = n45099 ;
  assign y1046 = n45102 ;
  assign y1047 = n45105 ;
  assign y1048 = n45108 ;
  assign y1049 = n4862 ;
  assign y1050 = n45111 ;
  assign y1051 = n45114 ;
  assign y1052 = n45117 ;
  assign y1053 = x67 ;
  assign y1054 = n45120 ;
  assign y1055 = n45122 ;
  assign y1056 = n45125 ;
  assign y1057 = n4795 ;
  assign y1058 = n45128 ;
  assign y1059 = n45131 ;
  assign y1060 = n45133 ;
  assign y1061 = n45135 ;
  assign y1062 = n45138 ;
  assign y1063 = n45147 ;
  assign y1064 = n45149 ;
  assign y1065 = n45152 ;
  assign y1066 = n45155 ;
  assign y1067 = n45158 ;
  assign y1068 = n45160 ;
  assign y1069 = n45163 ;
  assign y1070 = ~n45165 ;
  assign y1071 = n45168 ;
  assign y1072 = n45170 ;
  assign y1073 = n45173 ;
  assign y1074 = n45176 ;
  assign y1075 = n45179 ;
  assign y1076 = n45182 ;
  assign y1077 = n45184 ;
  assign y1078 = n45187 ;
  assign y1079 = n45190 ;
  assign y1080 = n45193 ;
  assign y1081 = n45196 ;
  assign y1082 = n45199 ;
  assign y1083 = n45202 ;
  assign y1084 = n45204 ;
  assign y1085 = n45207 ;
  assign y1086 = n45210 ;
  assign y1087 = n45213 ;
  assign y1088 = n45215 ;
  assign y1089 = n45217 ;
  assign y1090 = n45220 ;
  assign y1091 = n45222 ;
  assign y1092 = n45225 ;
  assign y1093 = n45228 ;
  assign y1094 = n45230 ;
  assign y1095 = n45233 ;
  assign y1096 = n45235 ;
  assign y1097 = n45238 ;
  assign y1098 = n45241 ;
  assign y1099 = n45244 ;
  assign y1100 = n45247 ;
  assign y1101 = n4712 ;
  assign y1102 = n45248 ;
  assign y1103 = n45250 ;
  assign y1104 = n45252 ;
  assign y1105 = ~n45255 ;
  assign y1106 = n14746 ;
  assign y1107 = n45256 ;
  assign y1108 = x1134 ;
  assign y1109 = x964 ;
  assign y1110 = ~x954 ;
  assign y1111 = x965 ;
  assign y1112 = n45258 ;
  assign y1113 = x991 ;
  assign y1114 = x985 ;
  assign y1115 = n45259 ;
  assign y1116 = n45260 ;
  assign y1117 = x1014 ;
  assign y1118 = n45261 ;
  assign y1119 = x1029 ;
  assign y1120 = x1004 ;
  assign y1121 = x1007 ;
  assign y1122 = n45262 ;
  assign y1123 = x1135 ;
  assign y1124 = n45263 ;
  assign y1125 = n45264 ;
  assign y1126 = n45265 ;
  assign y1127 = n45266 ;
  assign y1128 = n45267 ;
  assign y1129 = n45268 ;
  assign y1130 = ~x278 ;
  assign y1131 = n45269 ;
  assign y1132 = n45270 ;
  assign y1133 = ~n45271 ;
  assign y1134 = x1064 ;
  assign y1135 = n45272 ;
  assign y1136 = x299 ;
  assign y1137 = n45273 ;
  assign y1138 = x1075 ;
  assign y1139 = x1052 ;
  assign y1140 = x771 ;
  assign y1141 = x765 ;
  assign y1142 = x605 ;
  assign y1143 = x601 ;
  assign y1144 = x278 ;
  assign y1145 = x279 ;
  assign y1146 = ~x915 ;
  assign y1147 = ~x825 ;
  assign y1148 = ~x826 ;
  assign y1149 = ~x913 ;
  assign y1150 = ~x894 ;
  assign y1151 = ~x905 ;
  assign y1152 = x1095 ;
  assign y1153 = ~x890 ;
  assign y1154 = x1094 ;
  assign y1155 = ~x906 ;
  assign y1156 = ~x896 ;
  assign y1157 = ~x909 ;
  assign y1158 = ~x911 ;
  assign y1159 = ~x908 ;
  assign y1160 = ~x891 ;
  assign y1161 = ~x902 ;
  assign y1162 = ~x903 ;
  assign y1163 = ~x883 ;
  assign y1164 = ~x888 ;
  assign y1165 = ~x919 ;
  assign y1166 = ~x886 ;
  assign y1167 = ~x912 ;
  assign y1168 = ~x895 ;
  assign y1169 = ~x916 ;
  assign y1170 = ~x889 ;
  assign y1171 = ~x900 ;
  assign y1172 = ~x885 ;
  assign y1173 = ~x904 ;
  assign y1174 = ~x899 ;
  assign y1175 = ~x918 ;
  assign y1176 = ~x898 ;
  assign y1177 = ~x917 ;
  assign y1178 = ~x827 ;
  assign y1179 = ~x887 ;
  assign y1180 = ~x884 ;
  assign y1181 = ~x910 ;
  assign y1182 = ~x828 ;
  assign y1183 = ~x892 ;
  assign y1184 = x1187 ;
  assign y1185 = x1172 ;
  assign y1186 = x1170 ;
  assign y1187 = x1138 ;
  assign y1188 = x1177 ;
  assign y1189 = x1178 ;
  assign y1190 = x863 ;
  assign y1191 = x1203 ;
  assign y1192 = x1185 ;
  assign y1193 = x1171 ;
  assign y1194 = x1192 ;
  assign y1195 = x1137 ;
  assign y1196 = x1186 ;
  assign y1197 = x1165 ;
  assign y1198 = x1164 ;
  assign y1199 = x1098 ;
  assign y1200 = x1183 ;
  assign y1201 = x230 ;
  assign y1202 = x1169 ;
  assign y1203 = x1136 ;
  assign y1204 = x1181 ;
  assign y1205 = x849 ;
  assign y1206 = x1193 ;
  assign y1207 = x1182 ;
  assign y1208 = x1168 ;
  assign y1209 = x1175 ;
  assign y1210 = x1191 ;
  assign y1211 = x1099 ;
  assign y1212 = x1174 ;
  assign y1213 = x1179 ;
  assign y1214 = x1202 ;
  assign y1215 = x1176 ;
  assign y1216 = x1173 ;
  assign y1217 = x1201 ;
  assign y1218 = x1167 ;
  assign y1219 = x840 ;
  assign y1220 = x1189 ;
  assign y1221 = x1195 ;
  assign y1222 = x864 ;
  assign y1223 = x1190 ;
  assign y1224 = x1188 ;
  assign y1225 = x1180 ;
  assign y1226 = x1194 ;
  assign y1227 = x1097 ;
  assign y1228 = x1166 ;
  assign y1229 = x1200 ;
  assign y1230 = x1184 ;
endmodule
