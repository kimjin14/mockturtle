//Written by the Majority Logic Package Fri Nov 14 23:20:52 2014
module top (
            b255, a255, a254, b254, a253, b253, a252, b252, a251, b251, a250, b250, a249, b249, a248, b248, a247, b247, a246, b246, a245, b245, a244, b244, a243, b243, a242, b242, a241, b241, a240, b240, a239, b239, a238, b238, a237, b237, a236, b236, a235, b235, a234, b234, a233, b233, a232, b232, a231, b231, a230, b230, a229, b229, a228, b228, a227, b227, a226, b226, a225, b225, a224, b224, a223, b223, a222, b222, a221, b221, a220, b220, a219, b219, a218, b218, a217, b217, a216, b216, a215, b215, a214, b214, a213, b213, a212, b212, a211, b211, a210, b210, a209, b209, a208, b208, a207, b207, a206, b206, a205, b205, a204, b204, a203, b203, a202, b202, a201, b201, a200, b200, a199, b199, a198, b198, a197, b197, a196, b196, a195, b195, a194, b194, a193, b193, a192, b192, a191, b191, a190, b190, a189, b189, a188, b188, a187, b187, a186, b186, a185, b185, a184, b184, a183, b183, a182, b182, a181, b181, a180, b180, a179, b179, a178, b178, a177, b177, a176, b176, a175, b175, a174, b174, a173, b173, a172, b172, a171, b171, a170, b170, a169, b169, a168, b168, a167, b167, a166, b166, a165, b165, a164, b164, a163, b163, a162, b162, a161, b161, a160, b160, a159, b159, a158, b158, a157, b157, a156, b156, a155, b155, a154, b154, a153, b153, a152, b152, a151, b151, a150, b150, a149, b149, a148, b148, a147, b147, a146, b146, a145, b145, a144, b144, a143, b143, a142, b142, a141, b141, a140, b140, a139, b139, a138, b138, a137, b137, a136, b136, a135, b135, a134, b134, a133, b133, a132, b132, a131, b131, a130, b130, a129, b129, a128, b128, a127, b127, a126, b126, a125, b125, a124, b124, a123, b123, a122, b122, a121, b121, a120, b120, a119, b119, a118, b118, a117, b117, a116, b116, a115, b115, a114, b114, a113, b113, a112, b112, a111, b111, a110, b110, a109, b109, a108, b108, a107, b107, a106, b106, a105, b105, a104, b104, a103, b103, a102, b102, a101, b101, a100, b100, a99, b99, a98, b98, a97, b97, a96, b96, a95, b95, a94, b94, a93, b93, a92, b92, a91, b91, a90, b90, a89, b89, a88, b88, a87, b87, a86, b86, a85, b85, a84, b84, a83, b83, a82, b82, a81, b81, a80, b80, a79, b79, a78, b78, a77, b77, a76, b76, a75, b75, a74, b74, a73, b73, a72, b72, a71, b71, a70, b70, a69, b69, a68, b68, a67, b67, a66, b66, a65, b65, a64, b64, a63, b63, a62, b62, a61, b61, a60, b60, a59, b59, a58, b58, a57, b57, a56, b56, a55, b55, a54, b54, a53, b53, a52, b52, a51, b51, a50, b50, a49, b49, a48, b48, a47, b47, a46, b46, a45, b45, a44, b44, a43, b43, a42, b42, a41, b41, a40, b40, a39, b39, a38, b38, a37, b37, a36, b36, a35, b35, a34, b34, a33, b33, a32, b32, a31, b31, a30, b30, a29, b29, a28, b28, a27, b27, a26, b26, a25, b25, a24, b24, a23, b23, a22, b22, a21, b21, a20, b20, a19, b19, a18, b18, a17, b17, a16, b16, a15, b15, a14, b14, a13, b13, a12, b12, a11, b11, a10, b10, a9, b9, a8, b8, a7, b7, a6, b6, a5, b5, a4, b4, a3, b3, a2, b2, a1, b1, b0, cin, a0, 
            s0, s1, s2, s3, s4, s5, s6, s7, s8, s9, s10, s11, s12, s13, s14, s15, s16, s17, s18, s19, s20, s21, s22, s23, s24, s25, s26, s27, s28, s29, s30, s31, s32, s33, s34, s35, s36, s37, s38, s39, s40, s41, s42, s43, s44, s45, s46, s47, s48, s49, s50, s51, s52, s53, s54, s55, s56, s57, s58, s59, s60, s61, s62, s63, s64, s65, s66, s67, s68, s69, s70, s71, s72, s73, s74, s75, s76, s77, s78, s79, s80, s81, s82, s83, s84, s85, s86, s87, s88, s89, s90, s91, s92, s93, s94, s95, s96, s97, s98, s99, s100, s101, s102, s103, s104, s105, s106, s107, s108, s109, s110, s111, s112, s113, s114, s115, s116, s117, s118, s119, s120, s121, s122, s123, s124, s125, s126, s127, s128, s129, s130, s131, s132, s133, s134, s135, s136, s137, s138, s139, s140, s141, s142, s143, s144, s145, s146, s147, s148, s149, s150, s151, s152, s153, s154, s155, s156, s157, s158, s159, s160, s161, s162, s163, s164, s165, s166, s167, s168, s169, s170, s171, s172, s173, s174, s175, s176, s177, s178, s179, s180, s181, s182, s183, s184, s185, s186, s187, s188, s189, s190, s191, s192, s193, s194, s195, s196, s197, s198, s199, s200, s201, s202, s203, s204, s205, s206, s207, s208, s209, s210, s211, s212, s213, s214, s215, s216, s217, s218, s219, s220, s221, s222, s223, s224, s225, s226, s227, s228, s229, s230, s231, s232, s233, s234, s235, s236, s237, s238, s239, s240, s241, s242, s243, s244, s245, s246, s247, s248, s249, s250, s251, s252, s253, s254, s255, s256);
input b255, a255, a254, b254, a253, b253, a252, b252, a251, b251, a250, b250, a249, b249, a248, b248, a247, b247, a246, b246, a245, b245, a244, b244, a243, b243, a242, b242, a241, b241, a240, b240, a239, b239, a238, b238, a237, b237, a236, b236, a235, b235, a234, b234, a233, b233, a232, b232, a231, b231, a230, b230, a229, b229, a228, b228, a227, b227, a226, b226, a225, b225, a224, b224, a223, b223, a222, b222, a221, b221, a220, b220, a219, b219, a218, b218, a217, b217, a216, b216, a215, b215, a214, b214, a213, b213, a212, b212, a211, b211, a210, b210, a209, b209, a208, b208, a207, b207, a206, b206, a205, b205, a204, b204, a203, b203, a202, b202, a201, b201, a200, b200, a199, b199, a198, b198, a197, b197, a196, b196, a195, b195, a194, b194, a193, b193, a192, b192, a191, b191, a190, b190, a189, b189, a188, b188, a187, b187, a186, b186, a185, b185, a184, b184, a183, b183, a182, b182, a181, b181, a180, b180, a179, b179, a178, b178, a177, b177, a176, b176, a175, b175, a174, b174, a173, b173, a172, b172, a171, b171, a170, b170, a169, b169, a168, b168, a167, b167, a166, b166, a165, b165, a164, b164, a163, b163, a162, b162, a161, b161, a160, b160, a159, b159, a158, b158, a157, b157, a156, b156, a155, b155, a154, b154, a153, b153, a152, b152, a151, b151, a150, b150, a149, b149, a148, b148, a147, b147, a146, b146, a145, b145, a144, b144, a143, b143, a142, b142, a141, b141, a140, b140, a139, b139, a138, b138, a137, b137, a136, b136, a135, b135, a134, b134, a133, b133, a132, b132, a131, b131, a130, b130, a129, b129, a128, b128, a127, b127, a126, b126, a125, b125, a124, b124, a123, b123, a122, b122, a121, b121, a120, b120, a119, b119, a118, b118, a117, b117, a116, b116, a115, b115, a114, b114, a113, b113, a112, b112, a111, b111, a110, b110, a109, b109, a108, b108, a107, b107, a106, b106, a105, b105, a104, b104, a103, b103, a102, b102, a101, b101, a100, b100, a99, b99, a98, b98, a97, b97, a96, b96, a95, b95, a94, b94, a93, b93, a92, b92, a91, b91, a90, b90, a89, b89, a88, b88, a87, b87, a86, b86, a85, b85, a84, b84, a83, b83, a82, b82, a81, b81, a80, b80, a79, b79, a78, b78, a77, b77, a76, b76, a75, b75, a74, b74, a73, b73, a72, b72, a71, b71, a70, b70, a69, b69, a68, b68, a67, b67, a66, b66, a65, b65, a64, b64, a63, b63, a62, b62, a61, b61, a60, b60, a59, b59, a58, b58, a57, b57, a56, b56, a55, b55, a54, b54, a53, b53, a52, b52, a51, b51, a50, b50, a49, b49, a48, b48, a47, b47, a46, b46, a45, b45, a44, b44, a43, b43, a42, b42, a41, b41, a40, b40, a39, b39, a38, b38, a37, b37, a36, b36, a35, b35, a34, b34, a33, b33, a32, b32, a31, b31, a30, b30, a29, b29, a28, b28, a27, b27, a26, b26, a25, b25, a24, b24, a23, b23, a22, b22, a21, b21, a20, b20, a19, b19, a18, b18, a17, b17, a16, b16, a15, b15, a14, b14, a13, b13, a12, b12, a11, b11, a10, b10, a9, b9, a8, b8, a7, b7, a6, b6, a5, b5, a4, b4, a3, b3, a2, b2, a1, b1, b0, cin, a0;
output s0, s1, s2, s3, s4, s5, s6, s7, s8, s9, s10, s11, s12, s13, s14, s15, s16, s17, s18, s19, s20, s21, s22, s23, s24, s25, s26, s27, s28, s29, s30, s31, s32, s33, s34, s35, s36, s37, s38, s39, s40, s41, s42, s43, s44, s45, s46, s47, s48, s49, s50, s51, s52, s53, s54, s55, s56, s57, s58, s59, s60, s61, s62, s63, s64, s65, s66, s67, s68, s69, s70, s71, s72, s73, s74, s75, s76, s77, s78, s79, s80, s81, s82, s83, s84, s85, s86, s87, s88, s89, s90, s91, s92, s93, s94, s95, s96, s97, s98, s99, s100, s101, s102, s103, s104, s105, s106, s107, s108, s109, s110, s111, s112, s113, s114, s115, s116, s117, s118, s119, s120, s121, s122, s123, s124, s125, s126, s127, s128, s129, s130, s131, s132, s133, s134, s135, s136, s137, s138, s139, s140, s141, s142, s143, s144, s145, s146, s147, s148, s149, s150, s151, s152, s153, s154, s155, s156, s157, s158, s159, s160, s161, s162, s163, s164, s165, s166, s167, s168, s169, s170, s171, s172, s173, s174, s175, s176, s177, s178, s179, s180, s181, s182, s183, s184, s185, s186, s187, s188, s189, s190, s191, s192, s193, s194, s195, s196, s197, s198, s199, s200, s201, s202, s203, s204, s205, s206, s207, s208, s209, s210, s211, s212, s213, s214, s215, s216, s217, s218, s219, s220, s221, s222, s223, s224, s225, s226, s227, s228, s229, s230, s231, s232, s233, s234, s235, s236, s237, s238, s239, s240, s241, s242, s243, s244, s245, s246, s247, s248, s249, s250, s251, s252, s253, s254, s255, s256;
wire one, w0, w1, w2, w3, w4, w5, w6, w7, w8, w9, w10, w11, w12, w13, w14, w15, w16, w17, w18, w19, w20, w21, w22, w23, w24, w25, w26, w27, w28, w29, w30, w31, w32, w33, w34, w35, w36, w37, w38, w39, w40, w41, w42, w43, w44, w45, w46, w47, w48, w49, w50, w51, w52, w53, w54, w55, w56, w57, w58, w59, w60, w61, w62, w63, w64, w65, w66, w67, w68, w69, w70, w71, w72, w73, w74, w75, w76, w77, w78, w79, w80, w81, w82, w83, w84, w85, w86, w87, w88, w89, w90, w91, w92, w93, w94, w95, w96, w97, w98, w99, w100, w101, w102, w103, w104, w105, w106, w107, w108, w109, w110, w111, w112, w113, w114, w115, w116, w117, w118, w119, w120, w121, w122, w123, w124, w125, w126, w127, w128, w129, w130, w131, w132, w133, w134, w135, w136, w137, w138, w139, w140, w141, w142, w143, w144, w145, w146, w147, w148, w149, w150, w151, w152, w153, w154, w155, w156, w157, w158, w159, w160, w161, w162, w163, w164, w165, w166, w167, w168, w169, w170, w171, w172, w173, w174, w175, w176, w177, w178, w179, w180, w181, w182, w183, w184, w185, w186, w187, w188, w189, w190, w191, w192, w193, w194, w195, w196, w197, w198, w199, w200, w201, w202, w203, w204, w205, w206, w207, w208, w209, w210, w211, w212, w213, w214, w215, w216, w217, w218, w219, w220, w221, w222, w223, w224, w225, w226, w227, w228, w229, w230, w231, w232, w233, w234, w235, w236, w237, w238, w239, w240, w241, w242, w243, w244, w245, w246, w247, w248, w249, w250, w251, w252, w253, w254, w255, w256, w257, w258, w259, w260, w261, w262, w263, w264, w265, w266, w267, w268, w269, w270, w271, w272, w273, w274, w275, w276, w277, w278, w279, w280, w281, w282, w283, w284, w285, w286, w287, w288, w289, w290, w291, w292, w293, w294, w295, w296, w297, w298, w299, w300, w301, w302, w303, w304, w305, w306, w307, w308, w309, w310, w311, w312, w313, w314, w315, w316, w317, w318, w319, w320, w321, w322, w323, w324, w325, w326, w327, w328, w329, w330, w331, w332, w333, w334, w335, w336, w337, w338, w339, w340, w341, w342, w343, w344, w345, w346, w347, w348, w349, w350, w351, w352, w353, w354, w355, w356, w357, w358, w359, w360, w361, w362, w363, w364, w365, w366, w367, w368, w369, w370, w371, w372, w373, w374, w375, w376, w377, w378, w379, w380, w381, w382, w383, w384, w385, w386, w387, w388, w389, w390, w391, w392, w393, w394, w395, w396, w397, w398, w399, w400, w401, w402, w403, w404, w405, w406, w407, w408, w409, w410, w411, w412, w413, w414, w415, w416, w417, w418, w419, w420, w421, w422, w423, w424, w425, w426, w427, w428, w429, w430, w431, w432, w433, w434, w435, w436, w437, w438, w439, w440, w441, w442, w443, w444, w445, w446, w447, w448, w449, w450, w451, w452, w453, w454, w455, w456, w457, w458, w459, w460, w461, w462, w463, w464, w465, w466, w467, w468, w469, w470, w471, w472, w473, w474, w475, w476, w477, w478, w479, w480, w481, w482, w483, w484, w485, w486, w487, w488, w489, w490, w491, w492, w493, w494, w495, w496, w497, w498, w499, w500, w501, w502, w503, w504, w505, w506, w507, w508, w509, w510, w511, w512, w513, w514, w515, w516, w517, w518, w519, w520, w521, w522, w523, w524, w525, w526, w527, w528, w529, w530, w531, w532, w533, w534, w535, w536, w537, w538, w539, w540, w541, w542, w543, w544, w545, w546, w547, w548, w549, w550, w551, w552, w553, w554, w555, w556, w557, w558, w559, w560, w561, w562, w563, w564, w565, w566, w567, w568, w569, w570, w571, w572, w573, w574, w575, w576, w577, w578, w579, w580, w581, w582, w583, w584, w585, w586, w587, w588, w589, w590, w591, w592, w593, w594, w595, w596, w597, w598, w599, w600, w601, w602, w603, w604, w605, w606, w607, w608, w609, w610, w611, w612, w613, w614, w615, w616, w617, w618, w619, w620, w621, w622, w623, w624, w625, w626, w627, w628, w629, w630, w631, w632, w633, w634, w635, w636, w637, w638, w639, w640, w641, w642, w643, w644, w645, w646, w647, w648, w649, w650, w651, w652, w653, w654, w655, w656, w657, w658, w659, w660, w661, w662, w663, w664, w665, w666, w667, w668, w669, w670, w671, w672, w673, w674, w675, w676, w677, w678, w679, w680, w681, w682, w683, w684, w685, w686, w687, w688, w689, w690, w691, w692, w693, w694, w695, w696, w697, w698, w699, w700, w701, w702, w703, w704, w705, w706, w707, w708, w709, w710, w711, w712, w713, w714, w715, w716, w717, w718, w719, w720, w721, w722, w723, w724, w725, w726, w727, w728, w729, w730, w731, w732, w733, w734, w735, w736, w737, w738, w739, w740, w741, w742, w743, w744, w745, w746, w747, w748, w749, w750, w751, w752, w753, w754, w755, w756, w757, w758, w759, w760, w761, w762, w763, w764, w765, w766, w767, w768, w769, w770, w771, w772, w773, w774, w775, w776, w777, w778, w779, w780, w781, w782, w783, w784, w785, w786, w787, w788, w789, w790, w791, w792, w793, w794, w795, w796, w797, w798, w799, w800, w801, w802, w803, w804, w805, w806, w807, w808, w809, w810, w811, w812, w813, w814, w815, w816, w817, w818, w819, w820, w821, w822, w823, w824, w825, w826, w827, w828, w829, w830, w831, w832, w833, w834, w835, w836, w837, w838, w839, w840, w841, w842, w843, w844, w845, w846, w847, w848, w849, w850, w851, w852, w853, w854, w855, w856, w857, w858, w859, w860, w861, w862, w863, w864, w865, w866, w867, w868, w869, w870, w871, w872, w873, w874, w875, w876, w877, w878, w879, w880, w881, w882, w883, w884, w885, w886, w887, w888, w889, w890, w891, w892, w893, w894, w895, w896, w897, w898, w899, w900, w901, w902, w903, w904, w905, w906, w907, w908, w909, w910, w911, w912, w913, w914, w915, w916, w917, w918, w919, w920, w921, w922, w923, w924, w925, w926, w927, w928, w929, w930, w931, w932, w933, w934, w935, w936, w937, w938, w939, w940, w941, w942, w943, w944, w945, w946, w947, w948, w949, w950, w951, w952, w953, w954, w955, w956, w957, w958, w959, w960, w961, w962, w963, w964, w965, w966, w967, w968, w969, w970, w971, w972, w973, w974, w975, w976, w977, w978, w979, w980, w981, w982, w983, w984, w985, w986, w987, w988, w989, w990, w991, w992, w993, w994, w995, w996, w997, w998, w999, w1000, w1001, w1002, w1003, w1004, w1005, w1006, w1007, w1008, w1009, w1010, w1011, w1012, w1013, w1014, w1015, w1016, w1017, w1018, w1019, w1020, w1021, w1022, w1023, w1024, w1025, w1026, w1027, w1028, w1029, w1030, w1031, w1032, w1033, w1034, w1035, w1036, w1037, w1038, w1039, w1040, w1041, w1042, w1043, w1044, w1045, w1046, w1047, w1048, w1049, w1050, w1051, w1052, w1053, w1054, w1055, w1056, w1057, w1058, w1059, w1060, w1061, w1062, w1063, w1064, w1065, w1066, w1067, w1068, w1069, w1070, w1071, w1072, w1073, w1074, w1075, w1076, w1077, w1078, w1079, w1080, w1081, w1082, w1083, w1084, w1085, w1086, w1087, w1088, w1089, w1090, w1091, w1092, w1093, w1094, w1095, w1096, w1097, w1098, w1099, w1100, w1101, w1102, w1103, w1104, w1105, w1106, w1107, w1108, w1109, w1110, w1111, w1112, w1113, w1114, w1115, w1116, w1117, w1118, w1119, w1120, w1121, w1122, w1123, w1124, w1125, w1126, w1127, w1128, w1129, w1130, w1131, w1132, w1133, w1134, w1135, w1136, w1137, w1138, w1139, w1140, w1141, w1142, w1143, w1144, w1145, w1146, w1147, w1148, w1149, w1150, w1151, w1152, w1153, w1154, w1155, w1156, w1157, w1158, w1159, w1160, w1161, w1162, w1163, w1164, w1165, w1166, w1167, w1168, w1169, w1170, w1171, w1172, w1173, w1174, w1175, w1176, w1177, w1178, w1179, w1180, w1181, w1182, w1183, w1184, w1185, w1186, w1187, w1188, w1189, w1190, w1191, w1192, w1193, w1194, w1195, w1196, w1197, w1198, w1199, w1200, w1201, w1202, w1203, w1204, w1205, w1206, w1207, w1208, w1209, w1210, w1211, w1212, w1213, w1214, w1215, w1216, w1217, w1218, w1219, w1220, w1221, w1222, w1223, w1224, w1225, w1226, w1227, w1228, w1229, w1230, w1231, w1232, w1233, w1234, w1235, w1236, w1237, w1238, w1239, w1240, w1241, w1242, w1243, w1244, w1245, w1246, w1247, w1248, w1249, w1250, w1251, w1252, w1253, w1254, w1255, w1256, w1257, w1258, w1259, w1260, w1261, w1262, w1263, w1264, w1265, w1266, w1267, w1268, w1269, w1270, w1271, w1272, w1273, w1274, w1275, w1276, w1277, w1278, w1279, w1280, w1281, w1282, w1283, w1284, w1285, w1286, w1287, w1288, w1289, w1290, w1291, w1292, w1293, w1294, w1295, w1296, w1297, w1298, w1299, w1300, w1301, w1302, w1303, w1304, w1305, w1306, w1307, w1308, w1309, w1310, w1311, w1312, w1313, w1314, w1315, w1316, w1317, w1318, w1319, w1320, w1321, w1322, w1323, w1324, w1325, w1326, w1327, w1328, w1329, w1330, w1331, w1332, w1333, w1334, w1335, w1336, w1337, w1338, w1339, w1340, w1341, w1342, w1343, w1344, w1345, w1346, w1347, w1348, w1349, w1350, w1351, w1352, w1353, w1354, w1355, w1356, w1357, w1358, w1359, w1360, w1361, w1362, w1363, w1364, w1365, w1366, w1367, w1368, w1369, w1370, w1371, w1372, w1373, w1374, w1375, w1376, w1377, w1378, w1379, w1380, w1381, w1382, w1383, w1384, w1385, w1386, w1387, w1388, w1389, w1390, w1391, w1392, w1393, w1394, w1395, w1396, w1397, w1398, w1399, w1400, w1401, w1402, w1403, w1404, w1405, w1406, w1407, w1408, w1409, w1410, w1411, w1412, w1413, w1414, w1415, w1416, w1417, w1418, w1419, w1420, w1421, w1422, w1423, w1424, w1425, w1426, w1427, w1428, w1429, w1430, w1431, w1432, w1433, w1434, w1435, w1436, w1437, w1438, w1439, w1440, w1441, w1442, w1443, w1444, w1445, w1446, w1447, w1448, w1449, w1450, w1451, w1452, w1453, w1454, w1455, w1456, w1457, w1458, w1459, w1460, w1461, w1462, w1463, w1464, w1465, w1466, w1467, w1468, w1469, w1470, w1471, w1472, w1473, w1474, w1475, w1476, w1477, w1478, w1479, w1480, w1481, w1482, w1483, w1484, w1485, w1486, w1487, w1488, w1489, w1490, w1491, w1492, w1493, w1494, w1495, w1496, w1497, w1498, w1499, w1500, w1501, w1502, w1503, w1504, w1505, w1506, w1507, w1508, w1509, w1510, w1511, w1512, w1513, w1514, w1515, w1516, w1517, w1518, w1519, w1520, w1521, w1522, w1523, w1524, w1525, w1526, w1527, w1528, w1529, w1530, w1531, w1532, w1533, w1534, w1535, w1536, w1537, w1538, w1539, w1540, w1541, w1542, w1543, w1544, w1545, w1546, w1547, w1548, w1549, w1550, w1551, w1552, w1553, w1554, w1555, w1556, w1557, w1558, w1559, w1560, w1561, w1562, w1563, w1564, w1565, w1566, w1567, w1568, w1569, w1570, w1571, w1572, w1573, w1574, w1575, w1576, w1577, w1578, w1579, w1580, w1581, w1582, w1583, w1584, w1585, w1586, w1587, w1588, w1589, w1590, w1591, w1592, w1593, w1594, w1595, w1596, w1597, w1598, w1599, w1600, w1601, w1602, w1603, w1604, w1605, w1606, w1607, w1608, w1609, w1610, w1611, w1612, w1613, w1614, w1615, w1616, w1617, w1618, w1619, w1620, w1621, w1622, w1623, w1624, w1625, w1626, w1627, w1628, w1629, w1630, w1631, w1632, w1633, w1634, w1635, w1636, w1637, w1638, w1639, w1640, w1641, w1642, w1643, w1644, w1645, w1646, w1647, w1648, w1649, w1650, w1651, w1652, w1653, w1654, w1655, w1656, w1657, w1658, w1659, w1660, w1661, w1662, w1663, w1664, w1665, w1666, w1667, w1668, w1669, w1670, w1671, w1672, w1673, w1674, w1675, w1676, w1677, w1678, w1679, w1680, w1681, w1682, w1683, w1684, w1685, w1686, w1687, w1688, w1689, w1690, w1691, w1692, w1693, w1694, w1695, w1696, w1697, w1698, w1699, w1700, w1701, w1702, w1703, w1704, w1705, w1706, w1707, w1708, w1709, w1710, w1711, w1712, w1713, w1714, w1715, w1716, w1717, w1718, w1719, w1720, w1721, w1722, w1723, w1724, w1725, w1726, w1727, w1728, w1729, w1730, w1731, w1732, w1733, w1734, w1735, w1736, w1737, w1738, w1739, w1740, w1741, w1742, w1743, w1744, w1745, w1746, w1747, w1748, w1749, w1750, w1751, w1752, w1753, w1754, w1755, w1756, w1757, w1758, w1759, w1760, w1761, w1762, w1763, w1764, w1765, w1766, w1767, w1768, w1769, w1770, w1771, w1772, w1773, w1774, w1775, w1776, w1777, w1778, w1779, w1780, w1781, w1782, w1783, w1784, w1785, w1786, w1787, w1788, w1789, w1790, w1791, w1792, w1793, w1794, w1795, w1796, w1797, w1798, w1799, w1800, w1801, w1802, w1803, w1804, w1805, w1806, w1807, w1808, w1809, w1810, w1811, w1812, w1813, w1814, w1815, w1816, w1817, w1818, w1819, w1820, w1821, w1822, w1823, w1824, w1825, w1826, w1827, w1828, w1829, w1830, w1831, w1832, w1833, w1834, w1835, w1836, w1837, w1838, w1839, w1840, w1841, w1842, w1843, w1844, w1845, w1846, w1847, w1848, w1849, w1850, w1851, w1852, w1853, w1854, w1855, w1856, w1857, w1858, w1859, w1860, w1861, w1862, w1863, w1864, w1865, w1866, w1867, w1868, w1869, w1870, w1871, w1872, w1873, w1874, w1875, w1876, w1877, w1878, w1879, w1880, w1881, w1882, w1883, w1884, w1885, w1886, w1887, w1888, w1889, w1890, w1891, w1892, w1893, w1894, w1895, w1896, w1897, w1898, w1899, w1900, w1901, w1902, w1903, w1904, w1905, w1906, w1907, w1908, w1909, w1910, w1911, w1912, w1913, w1914, w1915, w1916, w1917, w1918, w1919, w1920, w1921, w1922, w1923, w1924, w1925, w1926, w1927, w1928, w1929, w1930, w1931, w1932, w1933, w1934, w1935, w1936, w1937, w1938, w1939, w1940, w1941, w1942, w1943, w1944, w1945, w1946, w1947, w1948, w1949, w1950, w1951, w1952, w1953, w1954, w1955, w1956, w1957, w1958, w1959, w1960, w1961, w1962, w1963, w1964, w1965, w1966, w1967, w1968, w1969, w1970, w1971, w1972, w1973, w1974, w1975, w1976, w1977, w1978, w1979, w1980, w1981, w1982, w1983, w1984, w1985, w1986, w1987, w1988, w1989, w1990, w1991, w1992, w1993, w1994, w1995, w1996, w1997, w1998, w1999, w2000, w2001, w2002, w2003, w2004, w2005, w2006, w2007, w2008, w2009, w2010, w2011, w2012, w2013, w2014, w2015, w2016, w2017, w2018, w2019, w2020, w2021, w2022, w2023, w2024, w2025, w2026, w2027, w2028, w2029, w2030, w2031, w2032, w2033, w2034, w2035, w2036, w2037, w2038, w2039, w2040, w2041, w2042, w2043, w2044, w2045, w2046, w2047, w2048, w2049, w2050, w2051, w2052, w2053, w2054, w2055, w2056, w2057, w2058, w2059, w2060, w2061, w2062, w2063, w2064, w2065, w2066, w2067, w2068, w2069, w2070, w2071, w2072, w2073, w2074, w2075, w2076, w2077, w2078, w2079, w2080, w2081, w2082, w2083, w2084, w2085, w2086, w2087, w2088, w2089, w2090, w2091, w2092, w2093, w2094, w2095, w2096, w2097, w2098, w2099, w2100, w2101, w2102, w2103, w2104, w2105, w2106, w2107, w2108, w2109, w2110, w2111, w2112, w2113, w2114, w2115, w2116, w2117, w2118, w2119, w2120, w2121, w2122, w2123, w2124, w2125, w2126, w2127, w2128, w2129, w2130, w2131, w2132, w2133, w2134, w2135, w2136, w2137, w2138, w2139, w2140, w2141, w2142, w2143, w2144, w2145, w2146, w2147, w2148, w2149, w2150, w2151, w2152, w2153, w2154, w2155, w2156, w2157, w2158, w2159, w2160, w2161, w2162, w2163, w2164, w2165, w2166, w2167, w2168, w2169, w2170, w2171, w2172, w2173, w2174, w2175, w2176, w2177, w2178, w2179, w2180, w2181, w2182, w2183, w2184, w2185, w2186, w2187, w2188, w2189, w2190, w2191, w2192, w2193, w2194, w2195, w2196, w2197, w2198, w2199, w2200, w2201, w2202, w2203, w2204, w2205, w2206, w2207, w2208, w2209, w2210, w2211, w2212, w2213, w2214, w2215, w2216, w2217, w2218, w2219, w2220, w2221, w2222, w2223, w2224, w2225, w2226, w2227, w2228, w2229, w2230, w2231, w2232, w2233, w2234, w2235, w2236, w2237, w2238, w2239, w2240, w2241, w2242, w2243, w2244, w2245, w2246, w2247, w2248, w2249, w2250, w2251, w2252, w2253, w2254, w2255, w2256, w2257, w2258, w2259, w2260, w2261, w2262, w2263, w2264, w2265, w2266, w2267, w2268, w2269, w2270, w2271, w2272, w2273, w2274, w2275, w2276, w2277, w2278, w2279, w2280, w2281, w2282, w2283, w2284, w2285, w2286, w2287, w2288, w2289, w2290, w2291, w2292, w2293, w2294, w2295, w2296, w2297, w2298, w2299, w2300, w2301, w2302, w2303, w2304, w2305, w2306, w2307, w2308, w2309, w2310, w2311, w2312, w2313, w2314, w2315, w2316, w2317, w2318, w2319, w2320, w2321, w2322, w2323, w2324, w2325, w2326, w2327, w2328, w2329, w2330, w2331, w2332, w2333, w2334, w2335, w2336, w2337, w2338, w2339, w2340, w2341, w2342, w2343, w2344, w2345, w2346, w2347, w2348, w2349, w2350, w2351, w2352, w2353, w2354, w2355, w2356, w2357, w2358, w2359, w2360, w2361, w2362, w2363, w2364, w2365, w2366, w2367, w2368, w2369, w2370, w2371, w2372, w2373, w2374, w2375, w2376, w2377, w2378, w2379, w2380, w2381, w2382, w2383, w2384, w2385, w2386, w2387, w2388, w2389, w2390, w2391, w2392, w2393, w2394, w2395, w2396, w2397, w2398, w2399, w2400, w2401, w2402, w2403, w2404, w2405, w2406, w2407, w2408, w2409, w2410, w2411, w2412, w2413, w2414, w2415, w2416, w2417, w2418, w2419, w2420, w2421, w2422, w2423, w2424, w2425, w2426, w2427, w2428, w2429, w2430, w2431, w2432, w2433, w2434, w2435, w2436, w2437, w2438, w2439, w2440, w2441, w2442, w2443, w2444, w2445, w2446, w2447, w2448, w2449, w2450, w2451, w2452, w2453, w2454, w2455, w2456, w2457, w2458, w2459, w2460, w2461, w2462, w2463, w2464, w2465, w2466, w2467, w2468, w2469, w2470, w2471, w2472, w2473, w2474, w2475, w2476, w2477, w2478, w2479, w2480, w2481, w2482, w2483, w2484, w2485, w2486, w2487, w2488, w2489, w2490, w2491, w2492, w2493, w2494, w2495, w2496, w2497, w2498, w2499, w2500, w2501, w2502, w2503, w2504, w2505, w2506, w2507, w2508, w2509, w2510, w2511, w2512, w2513, w2514, w2515, w2516, w2517, w2518, w2519, w2520, w2521, w2522, w2523, w2524, w2525, w2526, w2527, w2528, w2529, w2530, w2531, w2532, w2533, w2534, w2535, w2536, w2537, w2538, w2539, w2540, w2541, w2542, w2543, w2544, w2545, w2546, w2547, w2548, w2549, w2550, w2551, w2552, w2553, w2554, w2555, w2556, w2557, w2558, w2559, w2560, w2561, w2562, w2563, w2564, w2565, w2566, w2567, w2568, w2569, w2570, w2571, w2572, w2573, w2574, w2575, w2576, w2577, w2578, w2579, w2580, w2581, w2582, w2583, w2584, w2585, w2586, w2587, w2588, w2589, w2590, w2591, w2592, w2593, w2594, w2595, w2596, w2597, w2598, w2599, w2600, w2601, w2602, w2603, w2604, w2605, w2606, w2607, w2608, w2609, w2610, w2611, w2612, w2613, w2614, w2615, w2616, w2617, w2618, w2619, w2620, w2621, w2622, w2623, w2624, w2625, w2626, w2627, w2628, w2629, w2630, w2631, w2632, w2633, w2634, w2635, w2636, w2637, w2638, w2639, w2640, w2641, w2642, w2643, w2644, w2645, w2646, w2647, w2648, w2649, w2650, w2651, w2652, w2653, w2654, w2655, w2656, w2657, w2658, w2659, w2660, w2661, w2662, w2663, w2664, w2665, w2666, w2667, w2668, w2669, w2670, w2671, w2672, w2673, w2674, w2675, w2676, w2677, w2678, w2679, w2680, w2681, w2682, w2683, w2684, w2685, w2686, w2687, w2688, w2689, w2690, w2691, w2692, w2693, w2694, w2695, w2696, w2697, w2698, w2699, w2700, w2701, w2702, w2703, w2704, w2705, w2706, w2707, w2708, w2709, w2710, w2711, w2712, w2713, w2714, w2715, w2716, w2717, w2718, w2719, w2720, w2721, w2722, w2723, w2724, w2725, w2726, w2727, w2728, w2729, w2730, w2731, w2732, w2733, w2734, w2735, w2736, w2737, w2738, w2739, w2740, w2741, w2742, w2743, w2744, w2745, w2746, w2747, w2748, w2749, w2750, w2751, w2752, w2753, w2754, w2755, w2756, w2757, w2758, w2759, w2760, w2761, w2762, w2763, w2764, w2765, w2766, w2767, w2768, w2769, w2770, w2771, w2772, w2773, w2774, w2775, w2776, w2777, w2778, w2779, w2780, w2781, w2782, w2783, w2784, w2785, w2786, w2787, w2788, w2789, w2790, w2791, w2792, w2793, w2794, w2795, w2796, w2797, w2798, w2799, w2800, w2801, w2802, w2803, w2804, w2805, w2806, w2807, w2808, w2809, w2810, w2811, w2812, w2813, w2814, w2815, w2816, w2817, w2818, w2819, w2820, w2821, w2822, w2823, w2824, w2825, w2826, w2827, w2828, w2829, w2830, w2831, w2832, w2833, w2834, w2835, w2836, w2837, w2838, w2839, w2840, w2841, w2842, w2843, w2844, w2845, w2846, w2847, w2848, w2849, w2850, w2851, w2852, w2853, w2854, w2855, w2856, w2857, w2858, w2859, w2860, w2861, w2862, w2863, w2864, w2865, w2866, w2867, w2868, w2869, w2870, w2871, w2872, w2873, w2874, w2875, w2876, w2877, w2878, w2879, w2880, w2881, w2882, w2883, w2884, w2885, w2886, w2887, w2888, w2889, w2890, w2891, w2892, w2893, w2894, w2895, w2896, w2897, w2898, w2899, w2900, w2901, w2902, w2903, w2904, w2905, w2906, w2907, w2908, w2909, w2910, w2911, w2912, w2913, w2914, w2915, w2916, w2917, w2918, w2919, w2920, w2921, w2922, w2923, w2924, w2925, w2926, w2927, w2928, w2929, w2930, w2931, w2932, w2933, w2934, w2935, w2936, w2937, w2938, w2939, w2940, w2941, w2942, w2943, w2944, w2945, w2946, w2947, w2948, w2949, w2950, w2951, w2952, w2953, w2954, w2955, w2956, w2957, w2958, w2959, w2960, w2961, w2962, w2963, w2964, w2965, w2966, w2967, w2968, w2969, w2970, w2971, w2972, w2973, w2974, w2975, w2976, w2977, w2978, w2979, w2980, w2981, w2982, w2983, w2984, w2985, w2986, w2987, w2988, w2989, w2990, w2991, w2992, w2993, w2994, w2995, w2996, w2997, w2998, w2999, w3000, w3001, w3002, w3003, w3004, w3005, w3006, w3007, w3008, w3009, w3010, w3011, w3012, w3013, w3014, w3015, w3016, w3017, w3018, w3019, w3020, w3021, w3022, w3023, w3024, w3025, w3026, w3027, w3028, w3029, w3030, w3031, w3032, w3033, w3034, w3035, w3036, w3037, w3038, w3039, w3040, w3041, w3042, w3043, w3044, w3045, w3046, w3047, w3048, w3049, w3050, w3051, w3052, w3053, w3054, w3055, w3056, w3057, w3058, w3059, w3060, w3061, w3062, w3063, w3064, w3065, w3066, w3067, w3068, w3069, w3070, w3071, w3072, w3073, w3074, w3075, w3076, w3077, w3078, w3079, w3080, w3081, w3082, w3083, w3084, w3085, w3086, w3087, w3088, w3089, w3090, w3091, w3092, w3093, w3094, w3095, w3096, w3097, w3098, w3099, w3100, w3101, w3102, w3103, w3104, w3105, w3106, w3107, w3108, w3109, w3110, w3111, w3112, w3113, w3114, w3115, w3116, w3117, w3118, w3119, w3120, w3121, w3122, w3123, w3124, w3125, w3126, w3127, w3128, w3129, w3130, w3131, w3132, w3133, w3134, w3135, w3136, w3137, w3138, w3139, w3140, w3141, w3142, w3143, w3144, w3145, w3146, w3147, w3148, w3149, w3150, w3151, w3152, w3153, w3154, w3155, w3156, w3157, w3158, w3159, w3160, w3161, w3162, w3163, w3164, w3165, w3166, w3167, w3168, w3169, w3170, w3171, w3172, w3173, w3174, w3175, w3176, w3177, w3178, w3179, w3180, w3181, w3182, w3183, w3184, w3185, w3186, w3187, w3188, w3189, w3190, w3191, w3192, w3193, w3194, w3195, w3196, w3197, w3198, w3199, w3200, w3201, w3202, w3203, w3204, w3205, w3206, w3207, w3208, w3209, w3210, w3211, w3212, w3213, w3214, w3215, w3216, w3217, w3218, w3219, w3220, w3221, w3222, w3223, w3224, w3225, w3226, w3227, w3228, w3229, w3230, w3231, w3232, w3233, w3234, w3235, w3236, w3237, w3238, w3239, w3240, w3241, w3242, w3243, w3244, w3245, w3246, w3247, w3248, w3249, w3250, w3251, w3252, w3253, w3254, w3255, w3256, w3257, w3258, w3259, w3260, w3261, w3262, w3263, w3264, w3265, w3266, w3267, w3268, w3269, w3270, w3271, w3272, w3273, w3274, w3275, w3276, w3277, w3278, w3279, w3280, w3281, w3282, w3283, w3284, w3285, w3286, w3287, w3288, w3289, w3290, w3291, w3292, w3293, w3294, w3295, w3296, w3297, w3298, w3299, w3300, w3301, w3302, w3303, w3304, w3305, w3306, w3307, w3308, w3309, w3310, w3311, w3312, w3313, w3314, w3315, w3316, w3317, w3318, w3319, w3320, w3321, w3322, w3323, w3324, w3325, w3326, w3327, w3328, w3329, w3330, w3331, w3332, w3333, w3334, w3335, w3336, w3337, w3338, w3339, w3340, w3341, w3342, w3343, w3344, w3345, w3346, w3347, w3348, w3349, w3350, w3351, w3352, w3353, w3354, w3355, w3356, w3357, w3358, w3359, w3360, w3361, w3362, w3363, w3364, w3365, w3366, w3367, w3368, w3369, w3370, w3371, w3372, w3373, w3374, w3375, w3376, w3377, w3378, w3379, w3380, w3381, w3382, w3383, w3384, w3385, w3386, w3387, w3388, w3389, w3390, w3391, w3392, w3393, w3394, w3395, w3396, w3397, w3398, w3399, w3400, w3401, w3402, w3403, w3404, w3405, w3406, w3407, w3408, w3409, w3410, w3411, w3412, w3413, w3414, w3415, w3416, w3417, w3418, w3419, w3420, w3421, w3422, w3423, w3424, w3425, w3426, w3427, w3428, w3429, w3430, w3431, w3432, w3433, w3434, w3435, w3436, w3437, w3438, w3439, w3440, w3441, w3442, w3443, w3444, w3445, w3446, w3447, w3448, w3449, w3450, w3451, w3452, w3453, w3454, w3455, w3456, w3457, w3458, w3459, w3460, w3461, w3462, w3463, w3464, w3465, w3466, w3467, w3468, w3469, w3470, w3471, w3472, w3473, w3474, w3475, w3476, w3477, w3478, w3479, w3480, w3481, w3482, w3483, w3484, w3485, w3486, w3487, w3488, w3489, w3490, w3491, w3492, w3493, w3494, w3495, w3496, w3497, w3498, w3499, w3500, w3501, w3502, w3503, w3504, w3505, w3506, w3507, w3508, w3509, w3510, w3511, w3512, w3513, w3514, w3515, w3516, w3517, w3518, w3519, w3520, w3521, w3522, w3523, w3524, w3525, w3526, w3527, w3528, w3529, w3530, w3531, w3532, w3533, w3534, w3535, w3536, w3537, w3538, w3539, w3540, w3541, w3542, w3543, w3544, w3545, w3546, w3547, w3548, w3549, w3550, w3551, w3552, w3553, w3554, w3555, w3556, w3557, w3558, w3559, w3560, w3561, w3562, w3563, w3564, w3565, w3566, w3567, w3568, w3569, w3570, w3571, w3572, w3573, w3574, w3575, w3576, w3577, w3578, w3579, w3580, w3581, w3582, w3583, w3584, w3585, w3586, w3587, w3588, w3589, w3590, w3591, w3592, w3593, w3594, w3595, w3596, w3597, w3598, w3599, w3600, w3601, w3602, w3603, w3604, w3605, w3606, w3607, w3608, w3609, w3610, w3611, w3612, w3613, w3614, w3615, w3616, w3617, w3618, w3619, w3620, w3621, w3622, w3623, w3624, w3625, w3626, w3627, w3628, w3629, w3630, w3631, w3632, w3633, w3634, w3635, w3636, w3637, w3638, w3639, w3640, w3641, w3642, w3643, w3644, w3645, w3646, w3647, w3648, w3649, w3650, w3651, w3652, w3653, w3654, w3655, w3656, w3657, w3658, w3659, w3660, w3661, w3662, w3663, w3664, w3665, w3666, w3667, w3668, w3669, w3670, w3671, w3672, w3673, w3674, w3675, w3676, w3677, w3678, w3679, w3680, w3681, w3682, w3683, w3684, w3685, w3686, w3687, w3688, w3689, w3690, w3691, w3692, w3693, w3694, w3695, w3696, w3697, w3698, w3699, w3700, w3701, w3702, w3703, w3704, w3705, w3706, w3707, w3708, w3709, w3710, w3711, w3712, w3713, w3714, w3715, w3716, w3717, w3718, w3719, w3720, w3721, w3722, w3723, w3724, w3725, w3726, w3727, w3728, w3729, w3730, w3731, w3732, w3733, w3734, w3735, w3736, w3737, w3738, w3739, w3740, w3741, w3742, w3743, w3744, w3745, w3746, w3747, w3748, w3749, w3750, w3751, w3752, w3753, w3754, w3755, w3756, w3757, w3758, w3759, w3760, w3761, w3762, w3763, w3764, w3765, w3766, w3767, w3768, w3769, w3770, w3771, w3772, w3773, w3774, w3775, w3776, w3777, w3778, w3779, w3780, w3781, w3782, w3783, w3784, w3785, w3786, w3787, w3788, w3789, w3790, w3791, w3792, w3793, w3794, w3795, w3796, w3797, w3798, w3799, w3800, w3801, w3802, w3803, w3804, w3805, w3806, w3807, w3808, w3809, w3810, w3811, w3812, w3813, w3814, w3815, w3816, w3817, w3818, w3819, w3820, w3821, w3822, w3823, w3824, w3825, w3826, w3827, w3828, w3829, w3830, w3831, w3832, w3833, w3834, w3835, w3836, w3837, w3838, w3839, w3840, w3841, w3842, w3843, w3844, w3845, w3846, w3847, w3848, w3849, w3850, w3851, w3852, w3853, w3854, w3855, w3856, w3857, w3858, w3859, w3860, w3861, w3862, w3863, w3864, w3865, w3866, w3867, w3868, w3869, w3870, w3871, w3872, w3873, w3874, w3875, w3876, w3877, w3878, w3879, w3880, w3881, w3882, w3883, w3884, w3885, w3886, w3887, w3888, w3889, w3890, w3891, w3892, w3893, w3894, w3895, w3896, w3897, w3898, w3899, w3900, w3901, w3902, w3903, w3904, w3905, w3906, w3907, w3908, w3909, w3910, w3911, w3912, w3913, w3914, w3915, w3916, w3917, w3918, w3919, w3920, w3921, w3922, w3923, w3924, w3925, w3926, w3927, w3928, w3929, w3930, w3931, w3932, w3933, w3934, w3935, w3936, w3937, w3938, w3939, w3940, w3941, w3942, w3943, w3944, w3945, w3946, w3947, w3948, w3949, w3950, w3951, w3952, w3953, w3954, w3955, w3956, w3957, w3958, w3959, w3960, w3961, w3962, w3963, w3964, w3965, w3966, w3967, w3968, w3969, w3970, w3971, w3972, w3973, w3974, w3975, w3976, w3977, w3978, w3979, w3980, w3981, w3982, w3983, w3984, w3985, w3986, w3987, w3988, w3989, w3990, w3991, w3992, w3993, w3994, w3995, w3996, w3997, w3998, w3999, w4000, w4001, w4002, w4003, w4004, w4005, w4006, w4007, w4008, w4009, w4010, w4011, w4012, w4013, w4014, w4015, w4016, w4017, w4018, w4019, w4020, w4021, w4022, w4023, w4024, w4025, w4026, w4027, w4028, w4029, w4030, w4031, w4032, w4033, w4034, w4035, w4036, w4037, w4038, w4039, w4040, w4041, w4042, w4043, w4044, w4045, w4046, w4047, w4048, w4049, w4050, w4051, w4052, w4053, w4054, w4055, w4056, w4057, w4058, w4059, w4060, w4061, w4062, w4063, w4064, w4065, w4066, w4067, w4068, w4069, w4070, w4071, w4072, w4073, w4074, w4075, w4076, w4077, w4078, w4079, w4080, w4081, w4082, w4083, w4084, w4085, w4086, w4087, w4088, w4089, w4090, w4091, w4092, w4093, w4094, w4095, w4096, w4097, w4098, w4099, w4100, w4101, w4102, w4103, w4104, w4105, w4106, w4107, w4108, w4109, w4110, w4111, w4112, w4113, w4114, w4115, w4116, w4117, w4118, w4119, w4120, w4121, w4122, w4123, w4124, w4125, w4126, w4127, w4128, w4129, w4130, w4131, w4132, w4133, w4134, w4135, w4136, w4137, w4138, w4139, w4140, w4141, w4142, w4143, w4144, w4145, w4146, w4147, w4148, w4149, w4150, w4151, w4152, w4153, w4154, w4155, w4156, w4157, w4158, w4159, w4160, w4161, w4162, w4163, w4164, w4165, w4166, w4167, w4168, w4169, w4170, w4171, w4172, w4173, w4174, w4175, w4176, w4177, w4178, w4179, w4180, w4181, w4182, w4183, w4184, w4185, w4186, w4187, w4188, w4189, w4190, w4191, w4192, w4193, w4194, w4195, w4196, w4197, w4198, w4199, w4200, w4201, w4202, w4203, w4204, w4205, w4206, w4207, w4208, w4209, w4210, w4211, w4212, w4213, w4214, w4215, w4216, w4217, w4218, w4219, w4220, w4221, w4222, w4223, w4224, w4225, w4226, w4227, w4228, w4229, w4230, w4231, w4232, w4233, w4234, w4235, w4236, w4237, w4238, w4239, w4240, w4241, w4242, w4243, w4244, w4245, w4246, w4247, w4248, w4249, w4250, w4251, w4252, w4253, w4254, w4255, w4256, w4257, w4258, w4259, w4260, w4261, w4262, w4263, w4264, w4265, w4266, w4267, w4268, w4269, w4270, w4271, w4272, w4273, w4274, w4275, w4276, w4277, w4278, w4279, w4280, w4281, w4282, w4283, w4284, w4285, w4286, w4287, w4288, w4289, w4290, w4291, w4292, w4293, w4294, w4295, w4296, w4297, w4298, w4299, w4300, w4301, w4302, w4303, w4304, w4305, w4306, w4307, w4308, w4309, w4310, w4311, w4312, w4313, w4314, w4315, w4316, w4317, w4318, w4319, w4320, w4321, w4322, w4323, w4324, w4325, w4326, w4327, w4328, w4329, w4330, w4331, w4332, w4333, w4334, w4335, w4336, w4337, w4338, w4339, w4340, w4341, w4342, w4343, w4344, w4345, w4346, w4347, w4348, w4349, w4350, w4351, w4352, w4353, w4354, w4355, w4356, w4357, w4358, w4359, w4360, w4361, w4362, w4363, w4364, w4365, w4366, w4367, w4368, w4369, w4370, w4371, w4372, w4373, w4374, w4375, w4376, w4377, w4378, w4379, w4380, w4381, w4382, w4383, w4384, w4385, w4386, w4387, w4388, w4389, w4390, w4391, w4392, w4393, w4394, w4395, w4396, w4397, w4398, w4399, w4400, w4401, w4402, w4403, w4404, w4405, w4406, w4407, w4408, w4409, w4410, w4411, w4412, w4413, w4414, w4415, w4416, w4417, w4418, w4419, w4420, w4421, w4422, w4423, w4424, w4425, w4426, w4427, w4428, w4429, w4430, w4431, w4432, w4433, w4434, w4435, w4436, w4437, w4438, w4439, w4440, w4441, w4442, w4443, w4444, w4445, w4446, w4447, w4448, w4449, w4450, w4451, w4452, w4453, w4454, w4455, w4456, w4457, w4458, w4459, w4460, w4461, w4462, w4463, w4464, w4465, w4466, w4467, w4468, w4469, w4470, w4471, w4472, w4473, w4474, w4475, w4476, w4477, w4478, w4479, w4480, w4481, w4482, w4483, w4484, w4485, w4486, w4487, w4488, w4489, w4490, w4491, w4492, w4493, w4494, w4495, w4496, w4497, w4498, w4499, w4500, w4501, w4502, w4503, w4504, w4505, w4506, w4507, w4508, w4509, w4510, w4511, w4512, w4513, w4514, w4515, w4516, w4517, w4518, w4519, w4520, w4521, w4522, w4523, w4524, w4525, w4526, w4527, w4528, w4529, w4530, w4531, w4532, w4533, w4534, w4535, w4536, w4537, w4538, w4539, w4540, w4541, w4542, w4543, w4544, w4545, w4546, w4547, w4548, w4549, w4550, w4551, w4552, w4553, w4554, w4555, w4556, w4557, w4558, w4559, w4560, w4561, w4562, w4563, w4564, w4565, w4566, w4567, w4568, w4569, w4570, w4571, w4572, w4573, w4574, w4575, w4576, w4577, w4578, w4579, w4580, w4581, w4582, w4583, w4584, w4585, w4586, w4587, w4588, w4589, w4590, w4591, w4592, w4593, w4594, w4595, w4596, w4597, w4598, w4599, w4600, w4601, w4602, w4603, w4604, w4605, w4606, w4607, w4608, w4609, w4610, w4611, w4612, w4613, w4614, w4615, w4616, w4617, w4618, w4619, w4620, w4621, w4622, w4623, w4624, w4625, w4626, w4627, w4628, w4629, w4630, w4631, w4632, w4633, w4634, w4635, w4636, w4637, w4638, w4639, w4640, w4641, w4642, w4643, w4644, w4645, w4646, w4647, w4648, w4649, w4650, w4651, w4652, w4653, w4654, w4655, w4656, w4657, w4658, w4659, w4660, w4661, w4662, w4663, w4664, w4665, w4666, w4667, w4668, w4669, w4670, w4671, w4672, w4673, w4674, w4675, w4676, w4677, w4678, w4679, w4680, w4681, w4682, w4683, w4684, w4685, w4686, w4687, w4688, w4689, w4690, w4691, w4692, w4693, w4694, w4695, w4696, w4697, w4698, w4699, w4700, w4701, w4702, w4703, w4704, w4705, w4706, w4707, w4708, w4709, w4710, w4711, w4712, w4713, w4714, w4715, w4716, w4717, w4718, w4719, w4720, w4721, w4722, w4723, w4724, w4725, w4726, w4727, w4728, w4729, w4730, w4731, w4732, w4733, w4734, w4735, w4736, w4737, w4738, w4739, w4740, w4741, w4742, w4743, w4744, w4745, w4746, w4747, w4748, w4749, w4750, w4751, w4752, w4753, w4754, w4755, w4756, w4757, w4758, w4759, w4760, w4761, w4762, w4763, w4764, w4765, w4766, w4767, w4768, w4769, w4770, w4771, w4772, w4773, w4774, w4775, w4776, w4777, w4778, w4779, w4780, w4781, w4782, w4783, w4784, w4785, w4786, w4787, w4788, w4789, w4790, w4791, w4792, w4793, w4794, w4795, w4796, w4797, w4798, w4799, w4800, w4801, w4802, w4803, w4804, w4805, w4806, w4807, w4808, w4809, w4810, w4811, w4812, w4813, w4814, w4815, w4816, w4817, w4818, w4819, w4820, w4821, w4822, w4823, w4824, w4825, w4826, w4827, w4828, w4829, w4830, w4831, w4832, w4833, w4834, w4835, w4836, w4837, w4838, w4839, w4840, w4841, w4842, w4843, w4844, w4845, w4846, w4847, w4848, w4849, w4850, w4851, w4852, w4853, w4854, w4855, w4856, w4857, w4858, w4859, w4860, w4861, w4862, w4863, w4864, w4865, w4866, w4867, w4868, w4869, w4870, w4871, w4872, w4873, w4874, w4875, w4876, w4877, w4878, w4879, w4880, w4881, w4882, w4883, w4884, w4885, w4886, w4887, w4888, w4889, w4890, w4891, w4892, w4893, w4894, w4895, w4896, w4897, w4898, w4899, w4900, w4901, w4902, w4903, w4904, w4905, w4906, w4907, w4908, w4909, w4910, w4911, w4912, w4913, w4914, w4915, w4916, w4917, w4918, w4919, w4920, w4921, w4922, w4923, w4924, w4925, w4926, w4927, w4928, w4929, w4930, w4931, w4932, w4933, w4934, w4935, w4936, w4937, w4938, w4939, w4940, w4941, w4942, w4943, w4944, w4945, w4946, w4947, w4948, w4949, w4950, w4951, w4952, w4953, w4954, w4955, w4956, w4957, w4958, w4959, w4960, w4961, w4962, w4963, w4964, w4965, w4966, w4967, w4968, w4969, w4970, w4971, w4972, w4973, w4974, w4975, w4976, w4977, w4978, w4979, w4980, w4981, w4982, w4983, w4984, w4985, w4986, w4987, w4988, w4989, w4990, w4991, w4992, w4993, w4994, w4995, w4996, w4997, w4998, w4999, w5000, w5001, w5002, w5003, w5004, w5005, w5006, w5007, w5008, w5009, w5010, w5011, w5012, w5013, w5014, w5015, w5016, w5017, w5018, w5019, w5020, w5021, w5022, w5023, w5024, w5025, w5026, w5027, w5028, w5029, w5030, w5031, w5032, w5033, w5034, w5035, w5036, w5037, w5038, w5039, w5040, w5041, w5042, w5043, w5044, w5045, w5046, w5047, w5048, w5049, w5050, w5051, w5052, w5053, w5054, w5055, w5056, w5057, w5058, w5059, w5060, w5061, w5062, w5063, w5064, w5065, w5066, w5067, w5068, w5069, w5070, w5071, w5072, w5073, w5074, w5075, w5076, w5077, w5078, w5079, w5080, w5081, w5082, w5083, w5084, w5085, w5086, w5087, w5088, w5089, w5090, w5091, w5092, w5093, w5094, w5095, w5096, w5097, w5098, w5099, w5100, w5101, w5102, w5103, w5104, w5105, w5106, w5107, w5108, w5109, w5110, w5111, w5112, w5113, w5114, w5115, w5116, w5117, w5118, w5119, w5120, w5121, w5122, w5123, w5124, w5125, w5126, w5127, w5128, w5129, w5130, w5131, w5132, w5133, w5134, w5135, w5136, w5137, w5138, w5139, w5140, w5141, w5142, w5143, w5144, w5145, w5146, w5147, w5148, w5149, w5150, w5151, w5152, w5153, w5154, w5155, w5156, w5157, w5158, w5159, w5160, w5161, w5162, w5163, w5164, w5165, w5166, w5167, w5168, w5169, w5170, w5171, w5172, w5173, w5174, w5175, w5176, w5177, w5178, w5179, w5180, w5181, w5182, w5183, w5184, w5185, w5186, w5187, w5188, w5189, w5190, w5191, w5192, w5193, w5194, w5195, w5196, w5197, w5198, w5199, w5200, w5201, w5202, w5203, w5204, w5205, w5206, w5207, w5208, w5209, w5210, w5211, w5212, w5213, w5214, w5215, w5216, w5217, w5218, w5219, w5220, w5221, w5222, w5223, w5224, w5225, w5226, w5227, w5228, w5229, w5230, w5231, w5232, w5233, w5234, w5235, w5236, w5237, w5238, w5239, w5240, w5241, w5242, w5243, w5244, w5245, w5246, w5247, w5248, w5249, w5250, w5251, w5252, w5253, w5254, w5255, w5256, w5257, w5258, w5259, w5260, w5261, w5262, w5263, w5264, w5265, w5266, w5267, w5268, w5269, w5270, w5271, w5272, w5273, w5274, w5275, w5276, w5277, w5278, w5279, w5280, w5281, w5282, w5283, w5284, w5285, w5286, w5287, w5288, w5289, w5290, w5291, w5292, w5293, w5294, w5295, w5296, w5297, w5298, w5299, w5300, w5301, w5302, w5303, w5304, w5305, w5306, w5307, w5308, w5309, w5310, w5311, w5312, w5313, w5314, w5315, w5316, w5317, w5318, w5319, w5320, w5321, w5322, w5323, w5324, w5325, w5326, w5327, w5328, w5329, w5330, w5331, w5332, w5333, w5334, w5335, w5336, w5337, w5338, w5339, w5340, w5341, w5342, w5343, w5344, w5345, w5346, w5347, w5348, w5349, w5350, w5351, w5352, w5353, w5354, w5355, w5356, w5357, w5358, w5359, w5360, w5361, w5362, w5363, w5364, w5365, w5366, w5367, w5368, w5369, w5370, w5371, w5372, w5373, w5374, w5375, w5376, w5377, w5378, w5379, w5380, w5381, w5382, w5383, w5384, w5385, w5386, w5387, w5388, w5389, w5390, w5391, w5392, w5393, w5394, w5395, w5396, w5397, w5398, w5399, w5400, w5401, w5402, w5403, w5404, w5405, w5406, w5407, w5408, w5409, w5410, w5411, w5412, w5413, w5414, w5415, w5416, w5417, w5418, w5419, w5420, w5421, w5422, w5423, w5424, w5425, w5426, w5427, w5428, w5429, w5430, w5431, w5432, w5433, w5434, w5435, w5436, w5437, w5438, w5439, w5440, w5441, w5442, w5443, w5444, w5445, w5446, w5447, w5448, w5449, w5450, w5451, w5452, w5453, w5454, w5455, w5456, w5457, w5458, w5459, w5460, w5461, w5462, w5463, w5464, w5465, w5466, w5467, w5468, w5469, w5470, w5471, w5472, w5473, w5474, w5475, w5476, w5477, w5478, w5479, w5480, w5481, w5482, w5483, w5484, w5485, w5486, w5487, w5488, w5489, w5490, w5491, w5492, w5493, w5494, w5495, w5496, w5497, w5498, w5499, w5500, w5501, w5502, w5503, w5504, w5505, w5506, w5507, w5508, w5509, w5510, w5511, w5512, w5513, w5514, w5515, w5516, w5517, w5518, w5519, w5520, w5521, w5522, w5523, w5524, w5525, w5526, w5527, w5528, w5529, w5530, w5531, w5532, w5533, w5534, w5535, w5536, w5537, w5538, w5539, w5540, w5541, w5542, w5543, w5544, w5545, w5546, w5547, w5548, w5549, w5550, w5551, w5552, w5553, w5554, w5555, w5556, w5557, w5558, w5559, w5560, w5561, w5562, w5563, w5564, w5565, w5566, w5567, w5568, w5569, w5570, w5571, w5572, w5573, w5574, w5575, w5576, w5577, w5578, w5579, w5580, w5581, w5582, w5583, w5584, w5585, w5586, w5587, w5588, w5589, w5590, w5591, w5592, w5593, w5594, w5595, w5596, w5597, w5598, w5599, w5600, w5601, w5602, w5603, w5604, w5605, w5606, w5607, w5608, w5609, w5610, w5611, w5612, w5613, w5614, w5615, w5616, w5617, w5618, w5619, w5620, w5621, w5622, w5623, w5624, w5625, w5626, w5627, w5628, w5629, w5630, w5631, w5632, w5633, w5634, w5635, w5636, w5637, w5638, w5639, w5640, w5641, w5642, w5643, w5644, w5645, w5646, w5647, w5648, w5649, w5650, w5651, w5652, w5653, w5654, w5655, w5656, w5657, w5658, w5659, w5660, w5661, w5662, w5663, w5664, w5665, w5666, w5667, w5668, w5669, w5670, w5671, w5672, w5673, w5674, w5675, w5676, w5677, w5678, w5679, w5680, w5681, w5682, w5683, w5684, w5685, w5686, w5687, w5688, w5689, w5690, w5691, w5692, w5693, w5694, w5695, w5696, w5697, w5698, w5699, w5700, w5701, w5702, w5703, w5704, w5705, w5706, w5707, w5708, w5709, w5710, w5711, w5712, w5713, w5714, w5715, w5716, w5717, w5718, w5719, w5720, w5721, w5722, w5723, w5724, w5725, w5726, w5727, w5728, w5729, w5730, w5731, w5732, w5733, w5734, w5735, w5736, w5737, w5738, w5739, w5740, w5741, w5742, w5743, w5744, w5745, w5746, w5747, w5748, w5749, w5750, w5751, w5752, w5753, w5754, w5755, w5756, w5757, w5758, w5759, w5760, w5761, w5762, w5763, w5764, w5765, w5766, w5767, w5768, w5769, w5770, w5771, w5772, w5773, w5774, w5775, w5776, w5777, w5778, w5779, w5780, w5781, w5782, w5783, w5784, w5785, w5786, w5787, w5788, w5789, w5790, w5791, w5792, w5793, w5794, w5795, w5796, w5797, w5798, w5799, w5800, w5801, w5802, w5803, w5804, w5805, w5806, w5807, w5808, w5809, w5810, w5811, w5812, w5813, w5814, w5815, w5816, w5817, w5818, w5819, w5820, w5821, w5822, w5823, w5824, w5825, w5826, w5827, w5828, w5829, w5830, w5831, w5832, w5833, w5834, w5835, w5836, w5837, w5838, w5839, w5840, w5841, w5842, w5843, w5844, w5845, w5846, w5847, w5848, w5849, w5850, w5851, w5852, w5853, w5854, w5855, w5856, w5857, w5858, w5859, w5860, w5861, w5862, w5863, w5864, w5865, w5866, w5867, w5868, w5869, w5870, w5871, w5872, w5873, w5874, w5875, w5876, w5877, w5878, w5879, w5880, w5881, w5882, w5883, w5884, w5885, w5886, w5887, w5888, w5889, w5890, w5891, w5892, w5893, w5894, w5895, w5896, w5897, w5898, w5899, w5900, w5901, w5902, w5903, w5904, w5905, w5906, w5907, w5908, w5909, w5910, w5911, w5912, w5913, w5914, w5915, w5916, w5917, w5918, w5919, w5920, w5921, w5922, w5923, w5924, w5925, w5926, w5927, w5928, w5929, w5930, w5931, w5932, w5933, w5934, w5935, w5936, w5937, w5938, w5939, w5940, w5941, w5942, w5943, w5944, w5945, w5946, w5947, w5948, w5949, w5950, w5951, w5952, w5953, w5954, w5955, w5956, w5957, w5958, w5959, w5960, w5961, w5962, w5963, w5964, w5965, w5966, w5967, w5968, w5969, w5970, w5971, w5972, w5973, w5974, w5975, w5976, w5977, w5978, w5979, w5980, w5981, w5982, w5983, w5984, w5985, w5986, w5987, w5988, w5989, w5990, w5991, w5992, w5993, w5994, w5995, w5996, w5997, w5998, w5999, w6000, w6001, w6002, w6003, w6004, w6005, w6006, w6007, w6008, w6009, w6010, w6011, w6012, w6013, w6014, w6015, w6016, w6017, w6018, w6019, w6020, w6021, w6022, w6023, w6024, w6025, w6026, w6027, w6028, w6029, w6030, w6031, w6032, w6033, w6034, w6035, w6036, w6037, w6038, w6039, w6040, w6041, w6042, w6043, w6044, w6045, w6046, w6047, w6048, w6049, w6050, w6051, w6052, w6053, w6054, w6055, w6056, w6057, w6058, w6059, w6060, w6061, w6062, w6063, w6064, w6065, w6066, w6067, w6068, w6069, w6070, w6071, w6072, w6073, w6074, w6075, w6076, w6077, w6078, w6079, w6080, w6081, w6082, w6083, w6084, w6085, w6086, w6087, w6088, w6089, w6090, w6091, w6092, w6093, w6094, w6095, w6096, w6097, w6098, w6099, w6100, w6101, w6102, w6103, w6104, w6105, w6106, w6107, w6108, w6109, w6110, w6111, w6112, w6113, w6114, w6115, w6116, w6117, w6118, w6119, w6120, w6121, w6122, w6123, w6124, w6125, w6126, w6127, w6128, w6129, w6130, w6131, w6132, w6133, w6134, w6135, w6136, w6137, w6138, w6139, w6140, w6141, w6142, w6143, w6144, w6145, w6146, w6147, w6148, w6149, w6150, w6151, w6152, w6153, w6154, w6155, w6156, w6157, w6158, w6159, w6160, w6161, w6162, w6163, w6164, w6165, w6166, w6167, w6168, w6169, w6170, w6171, w6172, w6173, w6174, w6175, w6176, w6177, w6178, w6179, w6180, w6181, w6182, w6183, w6184, w6185, w6186, w6187, w6188, w6189, w6190, w6191, w6192, w6193, w6194, w6195, w6196, w6197, w6198, w6199, w6200, w6201, w6202, w6203, w6204, w6205, w6206, w6207, w6208, w6209, w6210, w6211, w6212, w6213, w6214, w6215, w6216, w6217, w6218, w6219, w6220, w6221, w6222, w6223, w6224, w6225, w6226, w6227, w6228, w6229, w6230, w6231, w6232, w6233, w6234, w6235, w6236, w6237, w6238, w6239, w6240, w6241, w6242, w6243, w6244, w6245, w6246, w6247, w6248, w6249, w6250, w6251, w6252, w6253, w6254, w6255, w6256, w6257, w6258, w6259, w6260, w6261, w6262, w6263, w6264, w6265, w6266, w6267, w6268, w6269, w6270, w6271, w6272, w6273, w6274, w6275, w6276, w6277, w6278, w6279, w6280, w6281, w6282, w6283, w6284, w6285, w6286, w6287, w6288, w6289, w6290, w6291, w6292, w6293, w6294, w6295, w6296, w6297, w6298, w6299, w6300, w6301, w6302, w6303, w6304, w6305, w6306, w6307, w6308, w6309, w6310, w6311, w6312, w6313, w6314, w6315, w6316, w6317, w6318, w6319, w6320, w6321, w6322, w6323, w6324, w6325, w6326, w6327, w6328, w6329, w6330, w6331, w6332, w6333, w6334, w6335, w6336, w6337, w6338, w6339, w6340, w6341, w6342, w6343, w6344, w6345, w6346, w6347, w6348, w6349, w6350, w6351, w6352, w6353, w6354, w6355, w6356, w6357, w6358, w6359, w6360, w6361, w6362, w6363, w6364, w6365, w6366, w6367, w6368, w6369, w6370, w6371, w6372, w6373, w6374, w6375, w6376, w6377, w6378, w6379, w6380, w6381, w6382, w6383, w6384, w6385, w6386, w6387, w6388, w6389, w6390, w6391, w6392, w6393, w6394, w6395, w6396, w6397, w6398, w6399, w6400, w6401, w6402, w6403, w6404, w6405, w6406, w6407, w6408, w6409, w6410, w6411, w6412, w6413, w6414, w6415, w6416, w6417, w6418, w6419, w6420, w6421, w6422, w6423, w6424, w6425, w6426, w6427, w6428, w6429, w6430, w6431, w6432, w6433, w6434, w6435, w6436, w6437, w6438, w6439, w6440, w6441, w6442, w6443, w6444, w6445, w6446, w6447, w6448, w6449, w6450, w6451, w6452, w6453, w6454, w6455, w6456, w6457, w6458, w6459, w6460, w6461, w6462, w6463, w6464, w6465, w6466, w6467, w6468, w6469, w6470, w6471, w6472, w6473, w6474, w6475, w6476, w6477, w6478, w6479, w6480, w6481, w6482, w6483, w6484, w6485, w6486, w6487, w6488, w6489, w6490, w6491, w6492, w6493, w6494, w6495, w6496, w6497, w6498, w6499, w6500, w6501, w6502, w6503, w6504, w6505, w6506, w6507, w6508, w6509, w6510, w6511, w6512, w6513, w6514, w6515, w6516, w6517, w6518, w6519, w6520, w6521, w6522, w6523, w6524, w6525, w6526, w6527, w6528, w6529, w6530, w6531, w6532, w6533, w6534, w6535, w6536, w6537, w6538, w6539, w6540, w6541, w6542, w6543, w6544, w6545, w6546, w6547, w6548, w6549, w6550, w6551, w6552, w6553, w6554, w6555, w6556, w6557, w6558, w6559, w6560, w6561, w6562, w6563, w6564, w6565, w6566, w6567, w6568, w6569, w6570, w6571, w6572, w6573, w6574, w6575, w6576, w6577, w6578, w6579, w6580, w6581, w6582, w6583, w6584, w6585, w6586, w6587, w6588, w6589, w6590, w6591, w6592, w6593, w6594, w6595, w6596, w6597, w6598, w6599, w6600, w6601, w6602, w6603, w6604, w6605, w6606, w6607, w6608, w6609, w6610, w6611, w6612, w6613, w6614, w6615, w6616, w6617, w6618, w6619, w6620, w6621, w6622, w6623, w6624, w6625, w6626, w6627, w6628, w6629, w6630, w6631, w6632, w6633, w6634, w6635, w6636, w6637, w6638, w6639, w6640, w6641, w6642, w6643, w6644, w6645, w6646, w6647, w6648, w6649, w6650, w6651, w6652, w6653, w6654, w6655, w6656, w6657, w6658, w6659, w6660, w6661, w6662, w6663, w6664, w6665, w6666, w6667, w6668, w6669, w6670, w6671, w6672, w6673, w6674, w6675, w6676, w6677, w6678, w6679, w6680, w6681, w6682, w6683, w6684, w6685, w6686, w6687, w6688, w6689, w6690, w6691, w6692, w6693, w6694, w6695, w6696, w6697, w6698, w6699, w6700, w6701, w6702, w6703, w6704, w6705, w6706, w6707, w6708, w6709, w6710, w6711, w6712, w6713, w6714, w6715, w6716, w6717, w6718, w6719, w6720, w6721, w6722, w6723, w6724, w6725, w6726, w6727, w6728, w6729, w6730, w6731, w6732, w6733, w6734, w6735, w6736, w6737, w6738, w6739, w6740, w6741, w6742, w6743, w6744, w6745, w6746, w6747, w6748, w6749, w6750, w6751, w6752, w6753, w6754, w6755, w6756, w6757, w6758, w6759, w6760, w6761, w6762, w6763, w6764, w6765, w6766, w6767, w6768, w6769, w6770, w6771, w6772, w6773, w6774, w6775, w6776, w6777, w6778, w6779, w6780, w6781, w6782, w6783, w6784, w6785, w6786, w6787, w6788, w6789, w6790, w6791, w6792, w6793, w6794, w6795, w6796, w6797, w6798, w6799, w6800, w6801, w6802, w6803, w6804, w6805, w6806, w6807, w6808, w6809, w6810, w6811, w6812, w6813, w6814, w6815, w6816, w6817, w6818, w6819, w6820, w6821, w6822, w6823, w6824, w6825, w6826, w6827, w6828, w6829, w6830, w6831, w6832, w6833, w6834, w6835, w6836, w6837, w6838, w6839, w6840, w6841, w6842, w6843, w6844, w6845, w6846, w6847, w6848, w6849, w6850, w6851, w6852, w6853, w6854, w6855, w6856, w6857, w6858, w6859, w6860, w6861, w6862, w6863, w6864, w6865, w6866, w6867, w6868, w6869, w6870, w6871, w6872, w6873, w6874, w6875, w6876, w6877, w6878, w6879, w6880, w6881, w6882, w6883, w6884, w6885, w6886, w6887, w6888, w6889, w6890, w6891, w6892, w6893, w6894, w6895, w6896, w6897, w6898, w6899, w6900, w6901, w6902, w6903, w6904, w6905, w6906, w6907, w6908, w6909, w6910, w6911, w6912, w6913, w6914, w6915, w6916, w6917, w6918, w6919, w6920, w6921, w6922, w6923, w6924, w6925, w6926, w6927, w6928, w6929, w6930, w6931, w6932, w6933, w6934, w6935, w6936, w6937, w6938, w6939, w6940, w6941, w6942, w6943, w6944, w6945, w6946, w6947, w6948, w6949, w6950, w6951, w6952, w6953, w6954, w6955, w6956, w6957, w6958, w6959, w6960, w6961, w6962, w6963, w6964, w6965, w6966, w6967, w6968, w6969, w6970, w6971, w6972, w6973, w6974, w6975, w6976, w6977, w6978, w6979, w6980, w6981, w6982, w6983, w6984, w6985, w6986, w6987, w6988, w6989, w6990, w6991, w6992, w6993, w6994, w6995, w6996, w6997, w6998, w6999, w7000, w7001, w7002, w7003, w7004, w7005, w7006, w7007, w7008, w7009, w7010, w7011, w7012, w7013, w7014, w7015, w7016, w7017, w7018, w7019, w7020, w7021, w7022, w7023, w7024, w7025, w7026, w7027, w7028, w7029, w7030, w7031, w7032, w7033, w7034, w7035, w7036, w7037, w7038, w7039, w7040, w7041, w7042, w7043, w7044, w7045, w7046, w7047, w7048, w7049, w7050, w7051, w7052, w7053, w7054, w7055, w7056, w7057, w7058, w7059, w7060, w7061, w7062, w7063, w7064, w7065, w7066, w7067, w7068, w7069, w7070, w7071, w7072, w7073, w7074, w7075, w7076, w7077, w7078, w7079, w7080, w7081, w7082, w7083, w7084, w7085, w7086, w7087, w7088, w7089, w7090, w7091, w7092, w7093, w7094, w7095, w7096, w7097, w7098, w7099, w7100, w7101, w7102, w7103, w7104, w7105, w7106, w7107, w7108, w7109, w7110, w7111, w7112, w7113, w7114, w7115, w7116, w7117, w7118, w7119, w7120, w7121, w7122, w7123, w7124, w7125, w7126, w7127, w7128, w7129, w7130, w7131, w7132, w7133, w7134, w7135, w7136, w7137, w7138, w7139, w7140, w7141, w7142, w7143, w7144, w7145, w7146, w7147, w7148, w7149, w7150, w7151, w7152, w7153, w7154, w7155, w7156, w7157, w7158, w7159, w7160, w7161, w7162, w7163, w7164, w7165, w7166, w7167, w7168, w7169, w7170, w7171, w7172, w7173, w7174, w7175, w7176, w7177, w7178, w7179, w7180, w7181, w7182, w7183, w7184, w7185, w7186, w7187, w7188, w7189, w7190, w7191, w7192, w7193, w7194, w7195, w7196, w7197, w7198, w7199, w7200, w7201, w7202, w7203, w7204, w7205, w7206, w7207, w7208, w7209, w7210, w7211, w7212, w7213, w7214, w7215, w7216, w7217, w7218, w7219, w7220, w7221, w7222, w7223, w7224, w7225, w7226, w7227, w7228, w7229, w7230, w7231, w7232, w7233, w7234, w7235, w7236, w7237, w7238, w7239, w7240, w7241, w7242, w7243, w7244, w7245, w7246, w7247, w7248, w7249, w7250, w7251, w7252, w7253, w7254, w7255, w7256, w7257, w7258, w7259, w7260, w7261, w7262, w7263, w7264, w7265, w7266, w7267, w7268, w7269, w7270, w7271, w7272, w7273, w7274, w7275, w7276, w7277, w7278, w7279, w7280, w7281, w7282, w7283, w7284, w7285, w7286, w7287, w7288, w7289, w7290, w7291, w7292, w7293, w7294, w7295, w7296, w7297, w7298, w7299, w7300, w7301, w7302, w7303, w7304, w7305, w7306, w7307, w7308, w7309, w7310, w7311, w7312, w7313, w7314, w7315, w7316, w7317, w7318, w7319, w7320, w7321, w7322, w7323, w7324, w7325, w7326, w7327, w7328, w7329, w7330, w7331, w7332, w7333, w7334, w7335, w7336, w7337, w7338, w7339, w7340, w7341, w7342, w7343, w7344, w7345, w7346, w7347, w7348, w7349, w7350, w7351, w7352, w7353, w7354, w7355, w7356, w7357, w7358, w7359, w7360, w7361, w7362, w7363, w7364, w7365, w7366, w7367, w7368, w7369, w7370, w7371, w7372, w7373, w7374, w7375, w7376, w7377, w7378, w7379, w7380, w7381, w7382, w7383, w7384, w7385, w7386, w7387, w7388, w7389, w7390, w7391, w7392, w7393, w7394, w7395, w7396, w7397, w7398, w7399, w7400, w7401, w7402, w7403, w7404, w7405, w7406, w7407, w7408, w7409, w7410, w7411, w7412, w7413, w7414, w7415, w7416, w7417, w7418, w7419, w7420, w7421, w7422, w7423, w7424, w7425, w7426, w7427, w7428, w7429, w7430, w7431, w7432, w7433, w7434, w7435, w7436, w7437, w7438, w7439, w7440, w7441, w7442, w7443, w7444, w7445, w7446, w7447, w7448, w7449, w7450, w7451, w7452, w7453, w7454, w7455, w7456, w7457, w7458, w7459, w7460, w7461, w7462, w7463, w7464, w7465, w7466, w7467, w7468, w7469, w7470, w7471, w7472, w7473, w7474, w7475, w7476, w7477, w7478, w7479, w7480, w7481, w7482, w7483, w7484, w7485, w7486, w7487, w7488, w7489, w7490, w7491, w7492, w7493, w7494, w7495, w7496, w7497, w7498, w7499, w7500, w7501, w7502, w7503, w7504, w7505, w7506, w7507, w7508, w7509, w7510, w7511, w7512, w7513, w7514, w7515, w7516, w7517, w7518, w7519, w7520, w7521, w7522, w7523, w7524, w7525, w7526, w7527, w7528, w7529, w7530, w7531, w7532, w7533, w7534, w7535, w7536, w7537, w7538, w7539, w7540, w7541, w7542, w7543, w7544, w7545, w7546, w7547, w7548, w7549, w7550, w7551, w7552, w7553, w7554, w7555, w7556, w7557, w7558, w7559, w7560, w7561, w7562, w7563, w7564, w7565, w7566, w7567, w7568, w7569, w7570, w7571, w7572, w7573, w7574, w7575, w7576, w7577, w7578, w7579, w7580, w7581, w7582, w7583, w7584, w7585, w7586, w7587, w7588, w7589, w7590, w7591, w7592, w7593, w7594, w7595, w7596, w7597, w7598, w7599, w7600, w7601, w7602, w7603, w7604, w7605, w7606, w7607, w7608, w7609, w7610, w7611, w7612, w7613, w7614, w7615, w7616, w7617, w7618, w7619, w7620, w7621, w7622, w7623, w7624, w7625, w7626, w7627, w7628, w7629, w7630, w7631, w7632, w7633, w7634, w7635, w7636, w7637, w7638, w7639, w7640, w7641, w7642, w7643, w7644, w7645, w7646, w7647, w7648, w7649;
assign w0 = ~w6920 & w2327;
assign w1 = (w6386 & w3843) | (w6386 & w4430) | (w3843 & w4430);
assign w2 = ~w7345 & w422;
assign w3 = (w1559 & w1340) | (w1559 & w7124) | (w1340 & w7124);
assign w4 = ~w4337 & w6220;
assign w5 = (w5178 & w132) | (w5178 & w5070) | (w132 & w5070);
assign w6 = (~w4647 & w4009) | (~w4647 & w1551) | (w4009 & w1551);
assign w7 = ~w7363 & w4457;
assign w8 = w3048 & ~w5007;
assign w9 = ~w640 & ~w3167;
assign w10 = (~w6594 & w1728) | (~w6594 & w6956) | (w1728 & w6956);
assign w11 = ~w6870 & w7399;
assign w12 = (w6661 & w1461) | (w6661 & w6461) | (w1461 & w6461);
assign w13 = ~a137 & ~b137;
assign w14 = (w5178 & w3801) | (w5178 & w6880) | (w3801 & w6880);
assign w15 = (~w1813 & w3636) | (~w1813 & w3116) | (w3636 & w3116);
assign w16 = (w442 & w5126) | (w442 & w2965) | (w5126 & w2965);
assign w17 = w7150 & ~w1346;
assign w18 = (~w3774 & w1372) | (~w3774 & w5131) | (w1372 & w5131);
assign w19 = (~w5528 & w5091) | (~w5528 & w368) | (w5091 & w368);
assign w20 = ~w3017 & w983;
assign w21 = (~w1598 & w4014) | (~w1598 & w2302) | (w4014 & w2302);
assign w22 = (~w6100 & w4053) | (~w6100 & w4073) | (w4053 & w4073);
assign w23 = w912 & w4893;
assign w24 = (~w909 & w6061) | (~w909 & ~w5042) | (w6061 & ~w5042);
assign w25 = (w5030 & w2047) | (w5030 & w6714) | (w2047 & w6714);
assign w26 = (~w5178 & w3299) | (~w5178 & w695) | (w3299 & w695);
assign w27 = ~w1379 & w3823;
assign w28 = (w5054 & w823) | (w5054 & ~w2279) | (w823 & ~w2279);
assign w29 = (w5528 & w23) | (w5528 & w6550) | (w23 & w6550);
assign w30 = ~w6104 & ~w4010;
assign w31 = (~w5834 & w7479) | (~w5834 & w7241) | (w7479 & w7241);
assign w32 = w5058 & w3314;
assign w33 = w4002 & ~w2077;
assign w34 = ~w3212 & ~w1371;
assign w35 = w6352 | w4202;
assign w36 = (~w195 & w6462) | (~w195 & w1743) | (w6462 & w1743);
assign w37 = (w6100 & w5405) | (w6100 & w7470) | (w5405 & w7470);
assign w38 = (w1555 & ~w5970) | (w1555 & w6687) | (~w5970 & w6687);
assign w39 = (w6748 & w7372) | (w6748 & w2601) | (w7372 & w2601);
assign w40 = w2441 & ~w6222;
assign w41 = (~w2456 & w5249) | (~w2456 & w2113) | (w5249 & w2113);
assign w42 = ~w2724 & ~w3691;
assign w43 = (w5257 & w5728) | (w5257 & w49) | (w5728 & w49);
assign w44 = w6634 & w1479;
assign w45 = ~w3023 & w6635;
assign w46 = ~w4306 & ~w3990;
assign w47 = w2108 & ~w1532;
assign w48 = w994 & ~w1470;
assign w49 = w3247 & w6833;
assign w50 = ~w4139 & ~w3982;
assign w51 = ~a57 & ~b57;
assign w52 = (~w3122 & ~w2210) | (~w3122 & w2274) | (~w2210 & w2274);
assign w53 = w3105 & ~w3804;
assign w54 = a186 & b186;
assign w55 = (w3427 & w1687) | (w3427 & w5611) | (w1687 & w5611);
assign w56 = ~w5983 & ~w5069;
assign w57 = a221 & b221;
assign w58 = w1692 & ~w4132;
assign w59 = (~w6467 & w402) | (~w6467 & w7593) | (w402 & w7593);
assign w60 = a15 & b15;
assign w61 = (w2910 & w175) | (w2910 & ~w6894) | (w175 & ~w6894);
assign w62 = ~w7385 & w1187;
assign w63 = ~a86 & ~b86;
assign w64 = ~w3855 & ~w6811;
assign w65 = w4066 & ~w3123;
assign w66 = ~w3097 & ~w3522;
assign w67 = (~w887 & w3953) | (~w887 & w2919) | (w3953 & w2919);
assign w68 = w5259 & w71;
assign w69 = ~w5242 & ~w5926;
assign w70 = w5385 & w320;
assign w71 = w2798 & w4480;
assign w72 = w5922 & w1791;
assign w73 = w3061 & w7238;
assign w74 = (w5834 & w2547) | (w5834 & w3322) | (w2547 & w3322);
assign w75 = ~w5599 & ~w960;
assign w76 = ~w3893 & ~w1085;
assign w77 = ~w3989 & w4378;
assign w78 = (~w5078 & w4980) | (~w5078 & w3763) | (w4980 & w3763);
assign w79 = ~w1080 & ~w4121;
assign w80 = (w4787 & w4273) | (w4787 & ~w3533) | (w4273 & ~w3533);
assign w81 = w701 & ~w1383;
assign w82 = w3729 & w3011;
assign w83 = (w1104 & w4157) | (w1104 & w3202) | (w4157 & w3202);
assign w84 = w3706 & ~w3289;
assign w85 = (w3318 & w5283) | (w3318 & w2075) | (w5283 & w2075);
assign w86 = ~w5555 & ~w860;
assign w87 = (w1161 & w3967) | (w1161 & w3050) | (w3967 & w3050);
assign w88 = ~w813 & w4250;
assign w89 = (w5655 & w3143) | (w5655 & w793) | (w3143 & w793);
assign w90 = (w3057 & w186) | (w3057 & w1016) | (w186 & w1016);
assign w91 = (~w2084 & w2365) | (~w2084 & w2093) | (w2365 & w2093);
assign w92 = ~w7011 & w4946;
assign w93 = (~w5178 & w6416) | (~w5178 & w1835) | (w6416 & w1835);
assign w94 = w455 & w699;
assign w95 = w6757 & ~w6884;
assign w96 = (~w488 & w3067) | (~w488 & w5544) | (w3067 & w5544);
assign w97 = w1105 & ~w6161;
assign w98 = (~w3840 & w2975) | (~w3840 & w3616) | (w2975 & w3616);
assign w99 = ~w3570 & w5152;
assign w100 = ~w5802 & w2230;
assign w101 = ~a118 & ~b118;
assign w102 = w593 & ~w1938;
assign w103 = (w2297 & w3119) | (w2297 & w5938) | (w3119 & w5938);
assign w104 = (w3852 & w5523) | (w3852 & w6959) | (w5523 & w6959);
assign w105 = (~w3318 & w1781) | (~w3318 & w3752) | (w1781 & w3752);
assign w106 = ~w6510 & ~w4366;
assign w107 = (~w4203 & w5298) | (~w4203 & w6599) | (w5298 & w6599);
assign w108 = w4384 & ~w2950;
assign w109 = ~w2671 & w1327;
assign w110 = w7187 & w3467;
assign w111 = ~w3001 & w4709;
assign w112 = ~w6994 & ~w2435;
assign w113 = (~w3774 & w6736) | (~w3774 & w7071) | (w6736 & w7071);
assign w114 = w2007 & ~w3358;
assign w115 = (w5871 & w7055) | (w5871 & w4311) | (w7055 & w4311);
assign w116 = (w2874 & w4226) | (w2874 & w5540) | (w4226 & w5540);
assign w117 = ~w6008 & ~w37;
assign w118 = w7630 & ~w980;
assign w119 = w456 & ~w6986;
assign w120 = (w5178 & w6941) | (w5178 & w7367) | (w6941 & w7367);
assign w121 = ~w5059 & w2384;
assign w122 = w4323 & ~w4898;
assign w123 = (w5178 & w669) | (w5178 & w219) | (w669 & w219);
assign w124 = ~w2634 & w4725;
assign w125 = ~w471 & ~w7614;
assign w126 = ~w384 & w3323;
assign w127 = (w6100 & w5459) | (w6100 & w4443) | (w5459 & w4443);
assign w128 = ~w3057 & w6268;
assign w129 = ~w1085 & ~w7373;
assign w130 = (w155 & w6775) | (w155 & w5291) | (w6775 & w5291);
assign w131 = (~w1575 & w2483) | (~w1575 & w5774) | (w2483 & w5774);
assign w132 = (w3737 & w6997) | (w3737 & w4315) | (w6997 & w4315);
assign w133 = (w4118 & w1015) | (w4118 & w7503) | (w1015 & w7503);
assign w134 = ~w336 & w2749;
assign w135 = (~w444 & w687) | (~w444 & w7212) | (w687 & w7212);
assign w136 = (w5419 & w3955) | (w5419 & w5310) | (w3955 & w5310);
assign w137 = (~w5734 & w3489) | (~w5734 & ~w2965) | (w3489 & ~w2965);
assign w138 = ~w5073 & w4310;
assign w139 = ~w7372 & w4079;
assign w140 = (~w693 & w2110) | (~w693 & ~w3580) | (w2110 & ~w3580);
assign w141 = ~w2259 & ~w525;
assign w142 = a130 & b130;
assign w143 = a121 & b121;
assign w144 = ~w7528 & w6044;
assign w145 = ~w4392 & w322;
assign w146 = (~w1071 & w3572) | (~w1071 & w2080) | (w3572 & w2080);
assign w147 = w3101 & ~w1057;
assign w148 = ~w3199 & w286;
assign w149 = ~w3836 & ~w3905;
assign w150 = (~w5178 & w5867) | (~w5178 & w5607) | (w5867 & w5607);
assign w151 = ~w5430 & w2342;
assign w152 = ~w1151 & ~w1778;
assign w153 = (w1868 & w5634) | (w1868 & w5099) | (w5634 & w5099);
assign w154 = ~w1141 & w7067;
assign w155 = (w6906 & w3018) | (w6906 & w4199) | (w3018 & w4199);
assign w156 = w4998 & ~w7256;
assign w157 = ~w2255 & w6448;
assign w158 = (w200 & w2777) | (w200 & w6606) | (w2777 & w6606);
assign w159 = ~w4261 & w3473;
assign w160 = (w7513 & w1557) | (w7513 & w5532) | (w1557 & w5532);
assign w161 = w7000 & ~w6772;
assign w162 = ~w1080 & ~w384;
assign w163 = ~w6920 & w193;
assign w164 = ~a131 & ~b131;
assign w165 = w4651 & w4328;
assign w166 = w2203 & ~w4236;
assign w167 = (~w2199 & w1608) | (~w2199 & ~w3119) | (w1608 & ~w3119);
assign w168 = (~w7322 & w4319) | (~w7322 & w4793) | (w4319 & w4793);
assign w169 = ~w6981 & w7563;
assign w170 = (w3819 & w6596) | (w3819 & w1224) | (w6596 & w1224);
assign w171 = ~w234 & w5860;
assign w172 = (~w5257 & w3590) | (~w5257 & w3829) | (w3590 & w3829);
assign w173 = (w1168 & w3077) | (w1168 & w2453) | (w3077 & w2453);
assign w174 = w2339 & w872;
assign w175 = (w7072 & w1708) | (w7072 & w4131) | (w1708 & w4131);
assign w176 = w6354 & ~w7480;
assign w177 = ~w6594 & w6100;
assign w178 = (w3284 & w2694) | (w3284 & w2002) | (w2694 & w2002);
assign w179 = w2108 & w5807;
assign w180 = w2613 & ~w6490;
assign w181 = w95 & w3821;
assign w182 = ~a35 & ~b35;
assign w183 = (w7418 & w2859) | (w7418 & ~w6174) | (w2859 & ~w6174);
assign w184 = (w4251 & w846) | (w4251 & ~w3819) | (w846 & ~w3819);
assign w185 = w1555 & ~w5961;
assign w186 = w4906 & w1508;
assign w187 = ~w5295 & w1098;
assign w188 = ~w2735 & w5478;
assign w189 = ~w2847 & w2473;
assign w190 = (~w3033 & w2220) | (~w3033 & w4807) | (w2220 & w4807);
assign w191 = ~w6340 & ~w6487;
assign w192 = (~w7300 & w6853) | (~w7300 & w5609) | (w6853 & w5609);
assign w193 = ~w6147 & w2142;
assign w194 = ~w6760 & ~w2124;
assign w195 = ~a205 & ~b205;
assign w196 = (~w6100 & w5443) | (~w6100 & w3367) | (w5443 & w3367);
assign w197 = ~w3816 & ~w7088;
assign w198 = ~w3989 & ~w1369;
assign w199 = w3141 & ~w2081;
assign w200 = w5641 & ~w2996;
assign w201 = ~w3919 & ~w5;
assign w202 = ~w887 & ~w4742;
assign w203 = (w7346 & w3232) | (w7346 & w1544) | (w3232 & w1544);
assign w204 = ~w2691 & ~w5566;
assign w205 = ~w7044 & ~w2005;
assign w206 = w1377 & ~w4940;
assign w207 = (w7330 & w5016) | (w7330 & w7015) | (w5016 & w7015);
assign w208 = ~w7294 & w5785;
assign w209 = (w2517 & w4714) | (w2517 & w1037) | (w4714 & w1037);
assign w210 = (w6100 & w967) | (w6100 & w1202) | (w967 & w1202);
assign w211 = (w3852 & w3966) | (w3852 & w6856) | (w3966 & w6856);
assign w212 = ~w1635 & ~w731;
assign w213 = (w6214 & w4773) | (w6214 & ~w3679) | (w4773 & ~w3679);
assign w214 = ~w3561 & ~w5788;
assign w215 = ~w638 & ~w3712;
assign w216 = a89 & b89;
assign w217 = ~w5402 & w4917;
assign w218 = (w5178 & w3545) | (w5178 & w5876) | (w3545 & w5876);
assign w219 = (w5325 & w1459) | (w5325 & w4996) | (w1459 & w4996);
assign w220 = ~w4412 & ~w6992;
assign w221 = (w5128 & w4475) | (w5128 & w2411) | (w4475 & w2411);
assign w222 = ~w4148 & w7510;
assign w223 = ~w2150 & ~w3460;
assign w224 = ~w6366 & ~w5773;
assign w225 = ~w1283 & w7447;
assign w226 = a156 & b156;
assign w227 = (w7437 & w4873) | (w7437 & w5325) | (w4873 & w5325);
assign w228 = (w1878 & ~w5948) | (w1878 & w4718) | (~w5948 & w4718);
assign w229 = w5423 & w3133;
assign w230 = w5111 & ~w3476;
assign w231 = w139 & w5572;
assign w232 = (w6166 & w3540) | (w6166 & w632) | (w3540 & w632);
assign w233 = w7231 & ~w424;
assign w234 = a225 & b225;
assign w235 = ~w1485 & ~w4168;
assign w236 = w139 & w6633;
assign w237 = (w1324 & w1232) | (w1324 & w1936) | (w1232 & w1936);
assign w238 = w1622 & ~w1804;
assign w239 = (w5774 & ~w5259) | (w5774 & w2985) | (~w5259 & w2985);
assign w240 = (w5807 & w179) | (w5807 & w3046) | (w179 & w3046);
assign w241 = (w4549 & w552) | (w4549 & w2784) | (w552 & w2784);
assign w242 = w3451 & ~w4687;
assign w243 = ~w4348 & w5032;
assign w244 = (~w2052 & w6402) | (~w2052 & w6205) | (w6402 & w6205);
assign w245 = ~w6025 & ~w1083;
assign w246 = w1756 & ~w5998;
assign w247 = ~a210 & ~b210;
assign w248 = w5629 & w6733;
assign w249 = w6640 & w4648;
assign w250 = w2965 & w1523;
assign w251 = (w1048 & w5308) | (w1048 & ~w6100) | (w5308 & ~w6100);
assign w252 = w5170 & ~w3336;
assign w253 = ~w7279 & w7255;
assign w254 = (w4647 & w2911) | (w4647 & w5271) | (w2911 & w5271);
assign w255 = (w4647 & w1637) | (w4647 & w2348) | (w1637 & w2348);
assign w256 = (w7300 & w565) | (w7300 & w4776) | (w565 & w4776);
assign w257 = (w1922 & w6555) | (w1922 & w5220) | (w6555 & w5220);
assign w258 = (w1774 & w5026) | (w1774 & w6100) | (w5026 & w6100);
assign w259 = ~w2735 & ~w727;
assign w260 = w2740 & w6614;
assign w261 = ~w2295 & ~w1610;
assign w262 = w2515 & ~w3217;
assign w263 = (~w3811 & ~w6723) | (~w3811 & ~w472) | (~w6723 & ~w472);
assign w264 = ~w1607 & w7462;
assign w265 = (w544 & w1586) | (w544 & ~w6100) | (w1586 & ~w6100);
assign w266 = (~w909 & w6061) | (~w909 & w7610) | (w6061 & w7610);
assign w267 = (~w1420 & w2050) | (~w1420 & w5420) | (w2050 & w5420);
assign w268 = (w6770 & w464) | (w6770 & w5395) | (w464 & w5395);
assign w269 = (~w5344 & w7) | (~w5344 & w2276) | (w7 & w2276);
assign w270 = (~w6966 & w5017) | (~w6966 & w2403) | (w5017 & w2403);
assign w271 = (~w5257 & w5677) | (~w5257 & w5897) | (w5677 & w5897);
assign w272 = w5939 & w5497;
assign w273 = w2353 & ~w6094;
assign w274 = ~w1485 & ~w554;
assign w275 = ~w4082 & w6680;
assign w276 = (~w3612 & w2456) | (~w3612 & w1081) | (w2456 & w1081);
assign w277 = (~w2199 & w6704) | (~w2199 & w6780) | (w6704 & w6780);
assign w278 = a56 & b56;
assign w279 = ~w3512 & w3758;
assign w280 = (w6557 & w5844) | (w6557 & w3983) | (w5844 & w3983);
assign w281 = (w2773 & w6715) | (w2773 & ~w1730) | (w6715 & ~w1730);
assign w282 = (~w5424 & w394) | (~w5424 & ~w593) | (w394 & ~w593);
assign w283 = w2062 & w740;
assign w284 = ~w2496 & ~w3007;
assign w285 = ~w2838 | w3841;
assign w286 = ~w3945 & ~w5115;
assign w287 = ~w4165 & w2948;
assign w288 = (~w215 & w634) | (~w215 & w3051) | (w634 & w3051);
assign w289 = ~w212 & ~w1295;
assign w290 = a5 & b5;
assign w291 = ~w2027 & w2650;
assign w292 = ~w3700 & w5541;
assign w293 = (w5178 & w1090) | (w5178 & w5533) | (w1090 & w5533);
assign w294 = w2238 & w6158;
assign w295 = (w5655 & w7433) | (w5655 & w5887) | (w7433 & w5887);
assign w296 = w2769 & w2969;
assign w297 = ~w5357 & w6327;
assign w298 = ~w4614 & w7566;
assign w299 = (~w7604 & w478) | (~w7604 & w6779) | (w478 & w6779);
assign w300 = w7544 & ~w681;
assign w301 = ~a182 & ~b182;
assign w302 = (~w5178 & w1653) | (~w5178 & w7109) | (w1653 & w7109);
assign w303 = (w4562 & w3737) | (w4562 & ~w2965) | (w3737 & ~w2965);
assign w304 = ~w1304 & w4961;
assign w305 = (w5178 & w5943) | (w5178 & w672) | (w5943 & w672);
assign w306 = (w7626 & w285) | (w7626 & w3271) | (w285 & w3271);
assign w307 = (w4296 & w449) | (w4296 & w6755) | (w449 & w6755);
assign w308 = w1315 & w4811;
assign w309 = (w472 & w3946) | (w472 & w3781) | (w3946 & w3781);
assign w310 = (w6217 & w7288) | (w6217 & w5778) | (w7288 & w5778);
assign w311 = (w3734 & w5189) | (w3734 & w641) | (w5189 & w641);
assign w312 = (w1365 & w1301) | (w1365 & ~w6174) | (w1301 & ~w6174);
assign w313 = (w6966 & w2040) | (w6966 & w886) | (w2040 & w886);
assign w314 = ~w7575 & w1554;
assign w315 = (~w2847 & w2395) | (~w2847 & w2330) | (w2395 & w2330);
assign w316 = w855 & w5685;
assign w317 = w6757 & w7563;
assign w318 = ~w6304 & ~w2450;
assign w319 = w234 & ~w7012;
assign w320 = (w679 & w559) | (w679 & w6267) | (w559 & w6267);
assign w321 = ~w4010 & w5751;
assign w322 = ~w7391 & w4271;
assign w323 = ~w3420 & ~w5100;
assign w324 = ~w3193 & ~w6996;
assign w325 = w6709 & ~w6981;
assign w326 = (~w3433 & w7222) | (~w3433 & w5681) | (w7222 & w5681);
assign w327 = w6138 & w7519;
assign w328 = (w1284 & ~w5445) | (w1284 & w5822) | (~w5445 & w5822);
assign w329 = (w4962 & w2417) | (w4962 & ~w5629) | (w2417 & ~w5629);
assign w330 = ~w2836 & ~w2203;
assign w331 = ~w7530 & ~w6463;
assign w332 = w5808 & ~w7265;
assign w333 = (~w7300 & w7237) | (~w7300 & w5609) | (w7237 & w5609);
assign w334 = ~w6170 & w4692;
assign w335 = ~a105 & ~b105;
assign w336 = a64 & b64;
assign w337 = (~w5834 & w4729) | (~w5834 & w7025) | (w4729 & w7025);
assign w338 = (w236 & w1225) | (w236 & w4324) | (w1225 & w4324);
assign w339 = (w3624 & w3694) | (w3624 & w5655) | (w3694 & w5655);
assign w340 = (~w2901 & w1727) | (~w2901 & w1130) | (w1727 & w1130);
assign w341 = (w4609 & w2146) | (w4609 & ~w6174) | (w2146 & ~w6174);
assign w342 = (~w5056 & w7616) | (~w5056 & ~w6656) | (w7616 & ~w6656);
assign w343 = ~w5368 & w3679;
assign w344 = ~w7042 & w950;
assign w345 = ~w6516 & ~w4566;
assign w346 = (w3188 & w668) | (w3188 & ~w471) | (w668 & ~w471);
assign w347 = ~w3168 & ~w5622;
assign w348 = ~w2913 & w1033;
assign w349 = ~w85 & ~w1209;
assign w350 = w6517 & w5345;
assign w351 = a158 & b158;
assign w352 = (w5059 & ~w664) | (w5059 & ~w4337) | (~w664 & ~w4337);
assign w353 = w1259 & ~w7555;
assign w354 = w5259 & w2557;
assign w355 = ~w6481 & ~w1898;
assign w356 = (w6100 & w915) | (w6100 & w2932) | (w915 & w2932);
assign w357 = (w3110 & w1018) | (w3110 & ~w3014) | (w1018 & ~w3014);
assign w358 = (w6688 & w5162) | (w6688 & w3584) | (w5162 & w3584);
assign w359 = ~w6374 & ~w465;
assign w360 = w3267 & w6112;
assign w361 = (w1346 & w3345) | (w1346 & ~w1678) | (w3345 & ~w1678);
assign w362 = w5555 & ~w5966;
assign w363 = ~w4132 & w6431;
assign w364 = w5573 & ~w6690;
assign w365 = ~w1485 & w7526;
assign w366 = (w4182 & w6961) | (w4182 & w7649) | (w6961 & w7649);
assign w367 = ~w1608 & w7072;
assign w368 = (w4638 & w2338) | (w4638 & w261) | (w2338 & w261);
assign w369 = w157 & w4101;
assign w370 = (w5828 & w7063) | (w5828 & w4394) | (w7063 & w4394);
assign w371 = (w5847 & w3008) | (w5847 & w1469) | (w3008 & w1469);
assign w372 = (w3422 & w7143) | (w3422 & w5403) | (w7143 & w5403);
assign w373 = (w6127 & w6923) | (w6127 & w6323) | (w6923 & w6323);
assign w374 = (w5178 & w6456) | (w5178 & w4411) | (w6456 & w4411);
assign w375 = w5596 & ~w3631;
assign w376 = (w6082 & w6433) | (w6082 & w4805) | (w6433 & w4805);
assign w377 = w242 & ~w563;
assign w378 = (w5655 & w6196) | (w5655 & w7415) | (w6196 & w7415);
assign w379 = w151 & w2678;
assign w380 = (~w6184 & w5564) | (~w6184 & ~w512) | (w5564 & ~w512);
assign w381 = w5248 & ~w6552;
assign w382 = ~w1164 & w1654;
assign w383 = (w3842 & w2339) | (w3842 & w961) | (w2339 & w961);
assign w384 = w4550 | w1621;
assign w385 = ~a222 & ~b222;
assign w386 = ~w3917 & w4126;
assign w387 = (w5516 & w7260) | (w5516 & w2929) | (w7260 & w2929);
assign w388 = w1751 & ~w6286;
assign w389 = ~w2433 & w3173;
assign w390 = ~a52 & ~b52;
assign w391 = ~a176 & ~b176;
assign w392 = (~w6100 & w3376) | (~w6100 & w209) | (w3376 & w209);
assign w393 = (~w1328 & w1138) | (~w1328 & w87) | (w1138 & w87);
assign w394 = w790 & ~w5424;
assign w395 = (~w5703 & w3885) | (~w5703 & w3214) | (w3885 & w3214);
assign w396 = ~w1756 & ~w7397;
assign w397 = w6031 & w7336;
assign w398 = w4151 | w6512;
assign w399 = ~w6553 & ~w5888;
assign w400 = w3514 & w6999;
assign w401 = w4203 & ~w5745;
assign w402 = (w200 & w2777) | (w200 & w7199) | (w2777 & w7199);
assign w403 = (~w5674 & w5438) | (~w5674 & w5688) | (w5438 & w5688);
assign w404 = (~w471 & w1066) | (~w471 & w5275) | (w1066 & w5275);
assign w405 = (w1559 & w1340) | (w1559 & w632) | (w1340 & w632);
assign w406 = (w1272 & ~w1974) | (w1272 & w6504) | (~w1974 & w6504);
assign w407 = ~w4325 & ~w1205;
assign w408 = (w1890 & w4141) | (w1890 & w6501) | (w4141 & w6501);
assign w409 = (~w6451 & w7534) | (~w6451 & w3508) | (w7534 & w3508);
assign w410 = w6353 & w1204;
assign w411 = ~w84 & w6625;
assign w412 = (~w4811 & w3396) | (~w4811 & w6019) | (w3396 & w6019);
assign w413 = (w3421 & w3185) | (w3421 & w2361) | (w3185 & w2361);
assign w414 = w4084 & w3162;
assign w415 = w2257 & w139;
assign w416 = (w488 & w6205) | (w488 & w5028) | (w6205 & w5028);
assign w417 = (w4337 & w3126) | (w4337 & w3529) | (w3126 & w3529);
assign w418 = (~w2123 & w1417) | (~w2123 & w2577) | (w1417 & w2577);
assign w419 = (w5257 & w3637) | (w5257 & w6794) | (w3637 & w6794);
assign w420 = ~w693 & w1709;
assign w421 = (w3200 & w7015) | (w3200 & w5264) | (w7015 & w5264);
assign w422 = ~w6450 & ~w7005;
assign w423 = (w3278 & w3226) | (w3278 & w5871) | (w3226 & w5871);
assign w424 = w7027 & ~w6791;
assign w425 = ~w5905 & w2321;
assign w426 = a37 & b37;
assign w427 = w5699 & ~w7026;
assign w428 = (w4161 & w705) | (w4161 & w5839) | (w705 & w5839);
assign w429 = (w1023 & w3986) | (w1023 & w2277) | (w3986 & w2277);
assign w430 = (w7197 & w3002) | (w7197 & w2227) | (w3002 & w2227);
assign w431 = ~w5782 & w6032;
assign w432 = ~w2714 & ~w3455;
assign w433 = (w6100 & w3479) | (w6100 & w1115) | (w3479 & w1115);
assign w434 = ~a232 & ~b232;
assign w435 = w4969 & w1642;
assign w436 = w4637 & w5870;
assign w437 = w2011 & ~w5416;
assign w438 = ~w3587 & w1250;
assign w439 = (~w5178 & w557) | (~w5178 & w1867) | (w557 & w1867);
assign w440 = ~w5555 & w2380;
assign w441 = ~w2261 & w7151;
assign w442 = (~w3267 & w2847) | (~w3267 & w5301) | (w2847 & w5301);
assign w443 = ~w1622 & w5423;
assign w444 = ~a141 & ~b141;
assign w445 = ~w1071 & ~w2215;
assign w446 = (w4926 & w5462) | (w4926 & ~w4867) | (w5462 & ~w4867);
assign w447 = (w6680 & w2351) | (w6680 & w5158) | (w2351 & w5158);
assign w448 = ~w5403 & ~w1071;
assign w449 = (w2534 & w6311) | (w2534 & ~w1544) | (w6311 & ~w1544);
assign w450 = ~w1697 & ~w4971;
assign w451 = (~w6467 & w6160) | (~w6467 & w1396) | (w6160 & w1396);
assign w452 = (w912 & w874) | (w912 & w4867) | (w874 & w4867);
assign w453 = ~w4747 & w1098;
assign w454 = a13 & b13;
assign w455 = ~w3202 & w699;
assign w456 = w6924 & w5485;
assign w457 = ~w3503 & w3137;
assign w458 = (w5834 & w5626) | (w5834 & w3307) | (w5626 & w3307);
assign w459 = (~w6100 & w237) | (~w6100 & w2180) | (w237 & w2180);
assign w460 = (~w7108 & w2026) | (~w7108 & w5740) | (w2026 & w5740);
assign w461 = w2600 & ~w1831;
assign w462 = (w5834 & w6322) | (w5834 & w3310) | (w6322 & w3310);
assign w463 = w5423 & ~w1153;
assign w464 = (~w6451 & w6608) | (~w6451 & w4531) | (w6608 & w4531);
assign w465 = (~w6100 & w1671) | (~w6100 & w2921) | (w1671 & w2921);
assign w466 = w3119 & w6051;
assign w467 = ~w4208 & w1105;
assign w468 = ~w6776 & ~w4193;
assign w469 = (~w5325 & w6505) | (~w5325 & w1657) | (w6505 & w1657);
assign w470 = (w1062 & w6773) | (w1062 & ~w2429) | (w6773 & ~w2429);
assign w471 = ~a54 & ~b54;
assign w472 = (~w676 & w109) | (~w676 & w2967) | (w109 & w2967);
assign w473 = (~w5259 & w2186) | (~w5259 & w4439) | (w2186 & w4439);
assign w474 = (w6989 & w1210) | (w6989 & w5430) | (w1210 & w5430);
assign w475 = w4415 & w7486;
assign w476 = w7113 & w2343;
assign w477 = w2496 & w3007;
assign w478 = ~w7158 & w2971;
assign w479 = w4448 & ~w7491;
assign w480 = (~w6966 & w6817) | (~w6966 & w1388) | (w6817 & w1388);
assign w481 = (w4044 & w1707) | (w4044 & w6100) | (w1707 & w6100);
assign w482 = w7257 | ~w3490;
assign w483 = ~w161 & ~w7414;
assign w484 = w813 & ~w5196;
assign w485 = (w2285 & w1785) | (w2285 & ~w3819) | (w1785 & ~w3819);
assign w486 = ~w13 & ~w792;
assign w487 = (~w6254 & w4613) | (~w6254 & w3265) | (w4613 & w3265);
assign w488 = w1796 & w7378;
assign w489 = ~w726 & ~w3652;
assign w490 = w2566 & w263;
assign w491 = w5163 & ~w2707;
assign w492 = w2726 | w1863;
assign w493 = (w5965 & ~w5032) | (w5965 & w6554) | (~w5032 & w6554);
assign w494 = (w4392 & w1201) | (w4392 & w5151) | (w1201 & w5151);
assign w495 = w1527 & w7394;
assign w496 = w338 | w3301;
assign w497 = w5858 & w1292;
assign w498 = w4222 & ~w472;
assign w499 = ~w6979 & w7228;
assign w500 = (~w1954 & w6329) | (~w1954 & w317) | (w6329 & w317);
assign w501 = (~w236 & w4865) | (~w236 & w4973) | (w4865 & w4973);
assign w502 = ~w3462 & ~w6147;
assign w503 = (w7 & w4106) | (w7 & ~w145) | (w4106 & ~w145);
assign w504 = ~w6685 & w1292;
assign w505 = ~a178 & ~b178;
assign w506 = (w1316 & w6829) | (w1316 & w730) | (w6829 & w730);
assign w507 = w1485 & w554;
assign w508 = w7363 & ~w4467;
assign w509 = w3333 & ~w1053;
assign w510 = (~w2046 & w3907) | (~w2046 & w1766) | (w3907 & w1766);
assign w511 = (w6100 & w2528) | (w6100 & w5327) | (w2528 & w5327);
assign w512 = ~w5402 & w4844;
assign w513 = w4747 & ~w6504;
assign w514 = ~w2822 & ~w6826;
assign w515 = (w8 & w7382) | (w8 & w2157) | (w7382 & w2157);
assign w516 = a183 & b183;
assign w517 = (~w3359 & ~w6002) | (~w3359 & w7314) | (~w6002 & w7314);
assign w518 = ~w4035 & w4300;
assign w519 = (~w6966 & w4939) | (~w6966 & w4489) | (w4939 & w4489);
assign w520 = ~w7150 & w3345;
assign w521 = ~w523 & ~w5025;
assign w522 = (w1515 & w4320) | (w1515 & ~w2997) | (w4320 & ~w2997);
assign w523 = ~w3732 & ~w57;
assign w524 = w3369 & w398;
assign w525 = (w5834 & w1948) | (w5834 & w3316) | (w1948 & w3316);
assign w526 = (w60 & ~w2096) | (w60 & ~w7385) | (~w2096 & ~w7385);
assign w527 = ~w3455 & ~w7278;
assign w528 = ~w7647 & w833;
assign w529 = w5106 & w2095;
assign w530 = w1260 & w1535;
assign w531 = ~w7546 & ~w3096;
assign w532 = (~w757 & w5944) | (~w757 & w5329) | (w5944 & w5329);
assign w533 = ~w4254 & ~w1874;
assign w534 = w4511 & ~w2122;
assign w535 = (w4825 & w376) | (w4825 & w7236) | (w376 & w7236);
assign w536 = w548 | w5776;
assign w537 = (w2169 & w6379) | (w2169 & ~w139) | (w6379 & ~w139);
assign w538 = (w5655 & w2390) | (w5655 & w3594) | (w2390 & w3594);
assign w539 = w7278 & ~w5777;
assign w540 = w5015 & w5556;
assign w541 = w4336 & ~w2386;
assign w542 = (w5699 & w2407) | (w5699 & w427) | (w2407 & w427);
assign w543 = ~w6252 & ~w2728;
assign w544 = ~w5588 & ~w226;
assign w545 = (w6781 & w2940) | (w6781 & ~w5291) | (w2940 & ~w5291);
assign w546 = (~w5777 & w6564) | (~w5777 & w5617) | (w6564 & w5617);
assign w547 = ~w7641 & ~w4107;
assign w548 = (~w523 & ~w5484) | (~w523 & w4841) | (~w5484 & w4841);
assign w549 = w3933 & w5995;
assign w550 = w6423 & w7187;
assign w551 = (w6649 & w6532) | (w6649 & ~w5870) | (w6532 & ~w5870);
assign w552 = w306 & w4102;
assign w553 = (w4187 & w5391) | (w4187 & w6976) | (w5391 & w6976);
assign w554 = ~w5147 & ~w2954;
assign w555 = w125 & ~w7204;
assign w556 = w649 & ~w6626;
assign w557 = (~w3952 & w7440) | (~w3952 & w2044) | (w7440 & w2044);
assign w558 = ~w6450 & ~w2080;
assign w559 = ~w1692 & w4132;
assign w560 = (w5178 & w6160) | (w5178 & w451) | (w6160 & w451);
assign w561 = w1004 & ~w5525;
assign w562 = (w1005 & w5043) | (w1005 & ~w5403) | (w5043 & ~w5403);
assign w563 = (w2928 & w5344) | (w2928 & w6731) | (w5344 & w6731);
assign w564 = (w2969 & w296) | (w2969 & ~w5576) | (w296 & ~w5576);
assign w565 = w6954 & w3246;
assign w566 = (w3737 & w2701) | (w3737 & w4264) | (w2701 & w4264);
assign w567 = w3478 & w1856;
assign w568 = w4384 & ~w1793;
assign w569 = a43 & b43;
assign w570 = w1288 & w646;
assign w571 = w5965 & ~w243;
assign w572 = ~w6343 & w6479;
assign w573 = (~w1071 & w3572) | (~w1071 & ~w5930) | (w3572 & ~w5930);
assign w574 = (w5178 & w6273) | (w5178 & w2397) | (w6273 & w2397);
assign w575 = (w4320 & w1133) | (w4320 & w4540) | (w1133 & w4540);
assign w576 = a124 & b124;
assign w577 = ~w6643 & ~w1463;
assign w578 = w1455 & ~w7106;
assign w579 = (w1598 & w2925) | (w1598 & w4932) | (w2925 & w4932);
assign w580 = w1447 & w353;
assign w581 = ~w1426 & ~w1664;
assign w582 = ~w6640 & ~w4648;
assign w583 = ~w5480 & ~w3462;
assign w584 = (w6100 & w7054) | (w6100 & w3613) | (w7054 & w3613);
assign w585 = ~w7113 & w3808;
assign w586 = w1574 & w3546;
assign w587 = w4759 & ~w426;
assign w588 = ~w1205 & ~w6760;
assign w589 = (w1457 & w4187) | (w1457 & w5448) | (w4187 & w5448);
assign w590 = w2410 & w2625;
assign w591 = ~w6935 & w5464;
assign w592 = (w6246 & w1044) | (w6246 & w4786) | (w1044 & w4786);
assign w593 = ~a160 & ~b160;
assign w594 = (w4671 & w2551) | (w4671 & w6687) | (w2551 & w6687);
assign w595 = ~w2448 & ~w6056;
assign w596 = (~w5178 & w7639) | (~w5178 & w1934) | (w7639 & w1934);
assign w597 = (~w2104 & w4074) | (~w2104 & w1792) | (w4074 & w1792);
assign w598 = (w5196 & w5945) | (w5196 & w1289) | (w5945 & w1289);
assign w599 = w7243 & w4915;
assign w600 = (w5178 & w1106) | (w5178 & w6975) | (w1106 & w6975);
assign w601 = ~w5364 & ~w2631;
assign w602 = (w5178 & w4291) | (w5178 & w6970) | (w4291 & w6970);
assign w603 = (w7197 & w3536) | (w7197 & w1984) | (w3536 & w1984);
assign w604 = a52 & b52;
assign w605 = ~w1851 & ~w5437;
assign w606 = (~w3737 & w3674) | (~w3737 & w6947) | (w3674 & w6947);
assign w607 = ~w6002 & ~w3359;
assign w608 = w2406 & ~w3150;
assign w609 = w4706 & w3647;
assign w610 = (~w3852 & w1679) | (~w3852 & w7248) | (w1679 & w7248);
assign w611 = (~w5178 & w6627) | (~w5178 & w3182) | (w6627 & w3182);
assign w612 = ~w7027 & w6033;
assign w613 = (~w6233 & w1206) | (~w6233 & w3899) | (w1206 & w3899);
assign w614 = w4428 & ~w4401;
assign w615 = (~w390 & w1206) | (~w390 & w1472) | (w1206 & w1472);
assign w616 = w3896 & ~w4505;
assign w617 = ~w3461 & w3916;
assign w618 = ~a81 & ~b81;
assign w619 = (w2627 & w7335) | (w2627 & w881) | (w7335 & w881);
assign w620 = w2261 & ~w3319;
assign w621 = ~w157 & w1266;
assign w622 = w222 & ~w343;
assign w623 = w757 & w329;
assign w624 = a53 & b53;
assign w625 = a75 & b75;
assign w626 = (w550 & w3414) | (w550 & w6942) | (w3414 & w6942);
assign w627 = (w2417 & w4962) | (w2417 & w1020) | (w4962 & w1020);
assign w628 = ~w5951 & w7403;
assign w629 = (w4130 & w1168) | (w4130 & w2453) | (w1168 & w2453);
assign w630 = (~w2627 & w3870) | (~w2627 & w6153) | (w3870 & w6153);
assign w631 = (~w860 & w7372) | (~w860 & w2160) | (w7372 & w2160);
assign w632 = ~w1607 & w4132;
assign w633 = w1621 & ~w618;
assign w634 = w4146 & ~w215;
assign w635 = (~w3947 & w1875) | (~w3947 & w473) | (w1875 & w473);
assign w636 = ~w441 & w5374;
assign w637 = w7118 & w228;
assign w638 = ~a224 & ~b224;
assign w639 = ~w990 & w4966;
assign w640 = ~a6 & ~b6;
assign w641 = ~w4036 & w587;
assign w642 = w1601 & ~w3075;
assign w643 = ~w4601 & ~w2927;
assign w644 = (w5178 & w7298) | (w5178 & w2350) | (w7298 & w2350);
assign w645 = (~w5257 & w3263) | (~w5257 & w7343) | (w3263 & w7343);
assign w646 = ~w3855 & w3052;
assign w647 = w5217 & ~w3444;
assign w648 = (w3984 & w2222) | (w3984 & w3914) | (w2222 & w3914);
assign w649 = ~w6526 & ~w2597;
assign w650 = w4890 & w1982;
assign w651 = a93 & b93;
assign w652 = w5484 & w1008;
assign w653 = ~w6540 & ~w6312;
assign w654 = (w2021 & w6727) | (w2021 & w7416) | (w6727 & w7416);
assign w655 = ~w4496 & w4418;
assign w656 = ~a159 & ~b159;
assign w657 = w7365 & w527;
assign w658 = (w5257 & w963) | (w5257 & w1695) | (w963 & w1695);
assign w659 = (w1880 & w3641) | (w1880 & w563) | (w3641 & w563);
assign w660 = ~w7647 & w5404;
assign w661 = (w1814 & w3089) | (w1814 & w3029) | (w3089 & w3029);
assign w662 = w2863 & ~w269;
assign w663 = w2173 & ~w6524;
assign w664 = w2005 & ~w5059;
assign w665 = ~w6331 & ~w2648;
assign w666 = ~w5510 & ~w2567;
assign w667 = (w3070 & ~w3212) | (w3070 & w1888) | (~w3212 & w1888);
assign w668 = ~w2197 & w3669;
assign w669 = (w4354 & w1459) | (w4354 & w7045) | (w1459 & w7045);
assign w670 = ~w5178 & w250;
assign w671 = (w4132 & w7462) | (w4132 & ~w3847) | (w7462 & ~w3847);
assign w672 = (w7587 & w5458) | (w7587 & w4104) | (w5458 & w4104);
assign w673 = (w3528 & w1723) | (w3528 & w1595) | (w1723 & w1595);
assign w674 = ~w2768 & ~w5515;
assign w675 = w336 & ~w1851;
assign w676 = w1485 & w7420;
assign w677 = (w1458 & w1956) | (w1458 & ~w4867) | (w1956 & ~w4867);
assign w678 = (w6945 & w1947) | (w6945 & w251) | (w1947 & w251);
assign w679 = ~w4167 & w4132;
assign w680 = (~w794 & w1905) | (~w794 & w6702) | (w1905 & w6702);
assign w681 = ~w5950 & ~w6181;
assign w682 = (~w1851 & w675) | (~w1851 & ~w2749) | (w675 & ~w2749);
assign w683 = (~w7187 & w1035) | (~w7187 & w3863) | (w1035 & w3863);
assign w684 = (~w5178 & w6696) | (~w5178 & w2372) | (w6696 & w2372);
assign w685 = (~w526 & w7192) | (~w526 & ~w3056) | (w7192 & ~w3056);
assign w686 = (w6353 & w2309) | (w6353 & w2879) | (w2309 & w2879);
assign w687 = ~w6426 & ~w3252;
assign w688 = ~w4182 | ~w7292;
assign w689 = w272 & ~w5228;
assign w690 = w1311 & w808;
assign w691 = (~w3774 & w5186) | (~w3774 & w3718) | (w5186 & w3718);
assign w692 = ~w234 & w385;
assign w693 = a244 & b244;
assign w694 = (w4753 & w18) | (w4753 & w6100) | (w18 & w6100);
assign w695 = (~w5325 & w7416) | (~w5325 & w654) | (w7416 & w654);
assign w696 = (w1168 & w5824) | (w1168 & w4210) | (w5824 & w4210);
assign w697 = (w1678 & w4768) | (w1678 & w759) | (w4768 & w759);
assign w698 = a206 & b206;
assign w699 = ~w1923 & w1158;
assign w700 = (~w5827 & w1437) | (~w5827 & w2697) | (w1437 & w2697);
assign w701 = ~w5170 & w3336;
assign w702 = ~w4638 & w5927;
assign w703 = ~w1431 & ~w3096;
assign w704 = (~w5257 & w5358) | (~w5257 & w985) | (w5358 & w985);
assign w705 = ~w314 & w3258;
assign w706 = a71 & b71;
assign w707 = (~w7097 & w6965) | (~w7097 & ~w4922) | (w6965 & ~w4922);
assign w708 = w5219 | w3212;
assign w709 = w6228 & w2782;
assign w710 = ~w5178 & w4098;
assign w711 = ~w554 & w235;
assign w712 = (w6904 & w2232) | (w6904 & w4521) | (w2232 & w4521);
assign w713 = ~w4191 & w3754;
assign w714 = ~w5676 & w3384;
assign w715 = (~w5178 & w1437) | (~w5178 & w700) | (w1437 & w700);
assign w716 = (w6746 & w2956) | (w6746 & w5727) | (w2956 & w5727);
assign w717 = (w4521 & w7446) | (w4521 & w6968) | (w7446 & w6968);
assign w718 = (~w714 & ~w2083) | (~w714 & ~w3533) | (~w2083 & ~w3533);
assign w719 = ~w5951 & w743;
assign w720 = (~w7172 & w6285) | (~w7172 & ~w6228) | (w6285 & ~w6228);
assign w721 = (~w2596 & w1263) | (~w2596 & w1352) | (w1263 & w1352);
assign w722 = (~w6922 & w2603) | (~w6922 & w5713) | (w2603 & w5713);
assign w723 = ~w5772 & ~w2295;
assign w724 = w1929 & ~w7204;
assign w725 = (w902 & w7513) | (w902 & w1673) | (w7513 & w1673);
assign w726 = (~w5178 & w4817) | (~w5178 & w1060) | (w4817 & w1060);
assign w727 = ~a158 & ~b158;
assign w728 = ~a106 & ~b106;
assign w729 = ~w6872 & w2311;
assign w730 = (~w2707 & w5391) | (~w2707 & w2647) | (w5391 & w2647);
assign w731 = ~w3033 & ~w4788;
assign w732 = ~w656 & ~w7634;
assign w733 = w3424 & ~w6361;
assign w734 = ~w6222 & ~w741;
assign w735 = ~w5345 & ~w6517;
assign w736 = ~a23 & ~b23;
assign w737 = (w101 & ~w2818) | (w101 & ~w1728) | (~w2818 & ~w1728);
assign w738 = ~w1285 & w1860;
assign w739 = w5009 & w5323;
assign w740 = ~w3176 & ~w3450;
assign w741 = w3173 & w3751;
assign w742 = (w716 & w6929) | (w716 & w2456) | (w6929 & w2456);
assign w743 = w3353 & ~w7506;
assign w744 = ~w4275 & ~w2725;
assign w745 = (w699 & w455) | (w699 & w3888) | (w455 & w3888);
assign w746 = (~w2123 & w2470) | (~w2123 & w1943) | (w2470 & w1943);
assign w747 = ~w6935 & ~w5778;
assign w748 = w2777 & w200;
assign w749 = w2288 & ~w6367;
assign w750 = ~w3989 & ~w6520;
assign w751 = (~w4251 & w478) | (~w4251 & w1442) | (w478 & w1442);
assign w752 = ~w3183 & w3974;
assign w753 = (~w6614 & w708) | (~w6614 & w2977) | (w708 & w2977);
assign w754 = w1058 & w7583;
assign w755 = ~w2586 & ~w4530;
assign w756 = (w1542 & w5347) | (w1542 & w4623) | (w5347 & w4623);
assign w757 = ~w6209 & ~w693;
assign w758 = ~w390 & ~w95;
assign w759 = ~w6628 & w6860;
assign w760 = (w5559 & w2900) | (w5559 & ~w553) | (w2900 & ~w553);
assign w761 = ~w3471 & ~w2435;
assign w762 = (w7168 & w1402) | (w7168 & w563) | (w1402 & w563);
assign w763 = ~w2011 & w5428;
assign w764 = ~w1581 & w5832;
assign w765 = ~w2742 & ~w2306;
assign w766 = ~w5760 & ~w6226;
assign w767 = ~w5762 & w9;
assign w768 = (w1168 & w2656) | (w1168 & w5824) | (w2656 & w5824);
assign w769 = ~w3019 & ~w651;
assign w770 = (~w6451 & w3022) | (~w6451 & w361) | (w3022 & w361);
assign w771 = w3523 & ~w1730;
assign w772 = ~w644 & ~w93;
assign w773 = (~w5178 & w5563) | (~w5178 & w7039) | (w5563 & w7039);
assign w774 = (w3318 & w447) | (w3318 & w6477) | (w447 & w6477);
assign w775 = ~w6630 & w1570;
assign w776 = ~w1486 & ~w3606;
assign w777 = (w4647 & w981) | (w4647 & w307) | (w981 & w307);
assign w778 = ~w5118 & ~w5119;
assign w779 = ~w3745 & w6871;
assign w780 = (~w1923 & w1903) | (~w1923 & w4252) | (w1903 & w4252);
assign w781 = (~w6177 & w6119) | (~w6177 & w3554) | (w6119 & w3554);
assign w782 = (w4251 & w846) | (w4251 & ~w7187) | (w846 & ~w7187);
assign w783 = (w5346 & w2603) | (w5346 & w2809) | (w2603 & w2809);
assign w784 = (w3863 & w6749) | (w3863 & w5562) | (w6749 & w5562);
assign w785 = ~w5309 & ~w3537;
assign w786 = ~w5597 & w888;
assign w787 = ~w147 & ~w7292;
assign w788 = ~w2644 & ~w6279;
assign w789 = (w5725 & w5320) | (w5725 & w2876) | (w5320 & w2876);
assign w790 = a160 & b160;
assign w791 = (~w5178 & w5265) | (~w5178 & w2743) | (w5265 & w2743);
assign w792 = a137 & b137;
assign w793 = (w2598 & w7008) | (w2598 & w4381) | (w7008 & w4381);
assign w794 = ~w2124 & w3731;
assign w795 = (~w7575 & w5977) | (~w7575 & w766) | (w5977 & w766);
assign w796 = (~w5178 & w4491) | (~w5178 & w733) | (w4491 & w733);
assign w797 = ~w4045 & w1740;
assign w798 = w5643 & ~w831;
assign w799 = w5622 & w2563;
assign w800 = (~w5788 & w2254) | (~w5788 & ~w2090) | (w2254 & ~w2090);
assign w801 = ~w1917 & ~w6218;
assign w802 = w3503 & w2272;
assign w803 = (w6100 & w6067) | (w6100 & w764) | (w6067 & w764);
assign w804 = ~a213 & ~b213;
assign w805 = w3828 & w7174;
assign w806 = w4778 & ~w749;
assign w807 = (w6027 & w3708) | (w6027 & w1706) | (w3708 & w1706);
assign w808 = ~w4616 & ~w2632;
assign w809 = w3391 & w3719;
assign w810 = ~w2279 & ~w1279;
assign w811 = (w2843 & w5974) | (w2843 & ~w6633) | (w5974 & ~w6633);
assign w812 = ~a150 & ~b150;
assign w813 = ~w4669 & w3273;
assign w814 = ~w2984 & ~w3682;
assign w815 = w7310 & ~w3051;
assign w816 = (w5871 & w2581) | (w5871 & w3998) | (w2581 & w3998);
assign w817 = ~w2631 & ~w7299;
assign w818 = w5640 & w4728;
assign w819 = w2299 & ~w164;
assign w820 = w4811 & ~w6252;
assign w821 = (w1863 & w2726) | (w1863 & ~w6174) | (w2726 & ~w6174);
assign w822 = (~w6738 & w1293) | (~w6738 & w5527) | (w1293 & w5527);
assign w823 = w7350 & w5054;
assign w824 = w420 & ~w6239;
assign w825 = w7405 & ~w6702;
assign w826 = (~w3989 & w1763) | (~w3989 & w4245) | (w1763 & w4245);
assign w827 = (w6966 & w6740) | (w6966 & w7040) | (w6740 & w7040);
assign w828 = ~w1321 & w6215;
assign w829 = (~w6082 & w7038) | (~w6082 & w7532) | (w7038 & w7532);
assign w830 = w4257 & w1886;
assign w831 = ~w6656 & w2274;
assign w832 = ~a51 & ~b51;
assign w833 = ~w143 & ~w5573;
assign w834 = (w3952 & w2114) | (w3952 & w6011) | (w2114 & w6011);
assign w835 = (w5395 & w6601) | (w5395 & w6199) | (w6601 & w6199);
assign w836 = ~w2991 & ~w6065;
assign w837 = (~w3947 & w1710) | (~w3947 & w718) | (w1710 & w718);
assign w838 = ~w2450 & ~w3328;
assign w839 = (~w5993 & w1713) | (~w5993 & w2785) | (w1713 & w2785);
assign w840 = (w7414 & w2741) | (w7414 & w3568) | (w2741 & w3568);
assign w841 = a175 & b175;
assign w842 = ~w3933 & ~w5995;
assign w843 = ~w5015 & ~w5556;
assign w844 = (w680 & w5306) | (w680 & w2125) | (w5306 & w2125);
assign w845 = (w6630 & w1355) | (w6630 & w6015) | (w1355 & w6015);
assign w846 = w4251 & ~w4697;
assign w847 = (~w5961 & w7401) | (~w5961 & w38) | (w7401 & w38);
assign w848 = ~w6451 & w6806;
assign w849 = (w918 & w387) | (w918 & ~w2876) | (w387 & ~w2876);
assign w850 = (~w7390 & w1352) | (~w7390 & w6250) | (w1352 & w6250);
assign w851 = (w5501 & w5093) | (w5501 & w5291) | (w5093 & w5291);
assign w852 = w2847 | w6949;
assign w853 = w6467 & w5431;
assign w854 = (w5739 & w367) | (w5739 & w2456) | (w367 & w2456);
assign w855 = ~w7528 & w7279;
assign w856 = (~w7345 & ~w2884) | (~w7345 & w5174) | (~w2884 & w5174);
assign w857 = w4167 & w5235;
assign w858 = ~w51 & w388;
assign w859 = (~w4884 & w5346) | (~w4884 & w6356) | (w5346 & w6356);
assign w860 = ~w4784 & ~w5966;
assign w861 = ~w478 & w4599;
assign w862 = (~w1328 & w5689) | (~w1328 & w6762) | (w5689 & w6762);
assign w863 = (w2123 & w5179) | (w2123 & w6168) | (w5179 & w6168);
assign w864 = (~w3318 & w1223) | (~w3318 & w3577) | (w1223 & w3577);
assign w865 = (w2179 & ~w1574) | (w2179 & w3164) | (~w1574 & w3164);
assign w866 = (~w7350 & w2533) | (~w7350 & w1279) | (w2533 & w1279);
assign w867 = (~w3986 & w3623) | (~w3986 & w6798) | (w3623 & w6798);
assign w868 = ~w7147 & w5797;
assign w869 = a44 & b44;
assign w870 = w4206 & w685;
assign w871 = (w3000 & w6261) | (w3000 & w3194) | (w6261 & w3194);
assign w872 = ~w1550 & ~w3689;
assign w873 = w1860 & w4504;
assign w874 = (w4893 & w3465) | (w4893 & w5528) | (w3465 & w5528);
assign w875 = ~w2229 & ~w4176;
assign w876 = (w1515 & w1133) | (w1515 & w522) | (w1133 & w522);
assign w877 = ~w4965 & ~w4212;
assign w878 = a240 & b240;
assign w879 = (~w5871 & w2395) | (~w5871 & w315) | (w2395 & w315);
assign w880 = ~w1649 & w5411;
assign w881 = (w3852 & w2936) | (w3852 & w2505) | (w2936 & w2505);
assign w882 = (~w236 & w6085) | (~w236 & w5712) | (w6085 & w5712);
assign w883 = ~w6935 & ~w1424;
assign w884 = ~w2515 & ~w1883;
assign w885 = ~w5347 & w3525;
assign w886 = w5980 & ~w4640;
assign w887 = ~w434 & ~w6630;
assign w888 = ~w3665 & ~w3083;
assign w889 = (w4045 & w1858) | (w4045 & ~w2885) | (w1858 & ~w2885);
assign w890 = ~w3750 & ~w2298;
assign w891 = (w7644 & w1353) | (w7644 & w129) | (w1353 & w129);
assign w892 = w3217 & ~w4060;
assign w893 = ~w5915 & ~w516;
assign w894 = ~w7538 & ~w5542;
assign w895 = (~w5178 & w3084) | (~w5178 & w4586) | (w3084 & w4586);
assign w896 = w19 | w4726;
assign w897 = ~w6549 & w3526;
assign w898 = w6553 & w1587;
assign w899 = (w7269 & w3005) | (w7269 & w7015) | (w3005 & w7015);
assign w900 = (~w5121 & w7513) | (~w5121 & w1398) | (w7513 & w1398);
assign w901 = w2630 & ~w759;
assign w902 = ~w2769 & w5849;
assign w903 = (~w2112 & w4171) | (~w2112 & w798) | (w4171 & w798);
assign w904 = ~w5120 & ~w6581;
assign w905 = ~w1541 & w2885;
assign w906 = ~w6643 & w2739;
assign w907 = ~w6272 & w6599;
assign w908 = a2 & b2;
assign w909 = ~w1580 & ~w6994;
assign w910 = ~w5486 & ~w4166;
assign w911 = (w5345 & w1334) | (w5345 & w6566) | (w1334 & w6566);
assign w912 = (w4893 & w3465) | (w4893 & w3473) | (w3465 & w3473);
assign w913 = ~w2515 & w972;
assign w914 = (w2334 & w5498) | (w2334 & ~w6174) | (w5498 & ~w6174);
assign w915 = (w1224 & w1185) | (w1224 & w4308) | (w1185 & w4308);
assign w916 = (w3104 & w704) | (w3104 & w5611) | (w704 & w5611);
assign w917 = ~w5608 & w294;
assign w918 = w2259 & w7448;
assign w919 = ~w3959 & ~w3580;
assign w920 = w3864 & w5013;
assign w921 = w5593 & w4440;
assign w922 = w4 & w6189;
assign w923 = w3774 & w1076;
assign w924 = (~w4350 & ~w5555) | (~w4350 & w7629) | (~w5555 & w7629);
assign w925 = ~w1760 & ~w2209;
assign w926 = ~w6658 & ~w6936;
assign w927 = (~w625 & w5555) | (~w625 & w5561) | (w5555 & w5561);
assign w928 = (~w2985 & w1951) | (~w2985 & w622) | (w1951 & w622);
assign w929 = w5998 & w1368;
assign w930 = (~w3318 & w4263) | (~w3318 & w1045) | (w4263 & w1045);
assign w931 = ~w4297 & ~w1712;
assign w932 = (~w5325 & w3539) | (~w5325 & w5845) | (w3539 & w5845);
assign w933 = w5751 & w7421;
assign w934 = (w5776 & w548) | (w5776 & w3248) | (w548 & w3248);
assign w935 = (w5572 & ~w3819) | (w5572 & w231) | (~w3819 & w231);
assign w936 = (~w5655 & w691) | (~w5655 & w2292) | (w691 & w2292);
assign w937 = ~a246 & ~b246;
assign w938 = w1039 & w1794;
assign w939 = (~w3847 & w2139) | (~w3847 & ~w3119) | (w2139 & ~w3119);
assign w940 = w7634 & ~w1878;
assign w941 = (~w5655 & w5154) | (~w5655 & w1318) | (w5154 & w1318);
assign w942 = (~w4651 & w5553) | (~w4651 & w1736) | (w5553 & w1736);
assign w943 = ~w948 & ~w2430;
assign w944 = ~w343 & w6877;
assign w945 = (~w5834 & w5339) | (~w5834 & w5610) | (w5339 & w5610);
assign w946 = ~w7216 & ~w3205;
assign w947 = (~w7302 & w4030) | (~w7302 & ~w6860) | (w4030 & ~w6860);
assign w948 = (w6100 & w6485) | (w6100 & w5095) | (w6485 & w5095);
assign w949 = (~w2985 & w213) | (~w2985 & w4981) | (w213 & w4981);
assign w950 = ~w4325 & ~w973;
assign w951 = ~w5721 & ~w5655;
assign w952 = (w5178 & w1054) | (w5178 & w6172) | (w1054 & w6172);
assign w953 = (~w3108 & w2078) | (~w3108 & w303) | (w2078 & w303);
assign w954 = w147 & ~w5277;
assign w955 = (w4202 & w6352) | (w4202 & ~w1649) | (w6352 & ~w1649);
assign w956 = ~w1851 & ~w134;
assign w957 = w4545 & ~w2749;
assign w958 = (~w3688 & w417) | (~w3688 & w1180) | (w417 & w1180);
assign w959 = (w6803 & w3323) | (w6803 & w162) | (w3323 & w162);
assign w960 = ~a253 & ~b253;
assign w961 = ~w2379 & w3035;
assign w962 = ~w5066 & w2666;
assign w963 = w6763 & w5567;
assign w964 = w4950 & w512;
assign w965 = w1287 & ~w3553;
assign w966 = (~w4521 & w2088) | (~w4521 & w5649) | (w2088 & w5649);
assign w967 = ~w4251 & w7351;
assign w968 = ~w5863 & ~w3092;
assign w969 = w7231 & ~w7047;
assign w970 = w5298 & ~w4203;
assign w971 = w505 & ~w2632;
assign w972 = a76 & b76;
assign w973 = a194 & b194;
assign w974 = (~w3953 & w3728) | (~w3953 & w3071) | (w3728 & w3071);
assign w975 = ~w2751 & ~w4179;
assign w976 = ~w331 & ~w4521;
assign w977 = (~w5655 & w2738) | (~w5655 & w3171) | (w2738 & w3171);
assign w978 = ~w2090 & w5469;
assign w979 = ~w6054 & ~w400;
assign w980 = ~w689 & w5838;
assign w981 = (~w1611 & w5531) | (~w1611 & w1014) | (w5531 & w1014);
assign w982 = ~w3561 & w2254;
assign w983 = ~w7190 & w7000;
assign w984 = ~w2435 & ~w792;
assign w985 = (w2686 & w3104) | (w2686 & w4657) | (w3104 & w4657);
assign w986 = w6512 & ~w3206;
assign w987 = (w3843 & w7481) | (w3843 & ~w1315) | (w7481 & ~w1315);
assign w988 = (w5231 & w6967) | (w5231 & w5403) | (w6967 & w5403);
assign w989 = (~w3892 & w6270) | (~w3892 & w1808) | (w6270 & w1808);
assign w990 = ~a72 & ~b72;
assign w991 = ~w5364 & w817;
assign w992 = (w3105 & w4190) | (w3105 & ~w3894) | (w4190 & ~w3894);
assign w993 = (w2124 & w5188) | (w2124 & w3575) | (w5188 & w3575);
assign w994 = w6562 & w6296;
assign w995 = (w4260 & ~w400) | (w4260 & w4781) | (~w400 & w4781);
assign w996 = (w2285 & w1785) | (w2285 & ~w7187) | (w1785 & ~w7187);
assign w997 = w5782 & ~w6032;
assign w998 = w4419 & ~w3173;
assign w999 = ~a127 & ~b127;
assign w1000 = (w6451 & w4509) | (w6451 & w697) | (w4509 & w697);
assign w1001 = ~w1954 & ~w5305;
assign w1002 = a78 & b78;
assign w1003 = ~w7328 & ~w4829;
assign w1004 = ~a211 & ~b211;
assign w1005 = ~w1822 & w4523;
assign w1006 = ~w5830 & w157;
assign w1007 = ~a129 & ~b129;
assign w1008 = w4811 & w543;
assign w1009 = (w6805 & w1235) | (w6805 & ~w1607) | (w1235 & ~w1607);
assign w1010 = ~w5054 & w5426;
assign w1011 = (w3831 & w233) | (w3831 & ~w2993) | (w233 & ~w2993);
assign w1012 = w4190 & w3105;
assign w1013 = w5616 & ~w6526;
assign w1014 = (w2534 & w6311) | (w2534 & ~w2966) | (w6311 & ~w2966);
assign w1015 = (w7414 & w5359) | (w7414 & w5203) | (w5359 & w5203);
assign w1016 = (w1888 & w7570) | (w1888 & w2661) | (w7570 & w2661);
assign w1017 = (~w686 & w2839) | (~w686 & w224) | (w2839 & w224);
assign w1018 = ~w4 & w3110;
assign w1019 = ~w5851 | w5702;
assign w1020 = w2417 | w632;
assign w1021 = w7391 & ~w3840;
assign w1022 = ~w3503 & ~w6270;
assign w1023 = ~w3019 & ~w2407;
assign w1024 = (~w6424 & w1522) | (~w6424 & w7419) | (w1522 & w7419);
assign w1025 = w1864 & w148;
assign w1026 = ~a71 & ~b71;
assign w1027 = (w7162 & w1513) | (w7162 & w3334) | (w1513 & w3334);
assign w1028 = (w4143 & w5521) | (w4143 & w2251) | (w5521 & w2251);
assign w1029 = w7010 & ~w2453;
assign w1030 = ~w4333 & w3821;
assign w1031 = (w1272 & ~w1974) | (w1272 & w1544) | (~w1974 & w1544);
assign w1032 = (w777 & w2858) | (w777 & w717) | (w2858 & w717);
assign w1033 = ~w7213 & ~w1137;
assign w1034 = w6753 & ~w1371;
assign w1035 = (w3863 & w7060) | (w3863 & w6749) | (w7060 & w6749);
assign w1036 = ~w3836 & ~w6572;
assign w1037 = (w7273 & w3755) | (w7273 & ~w7187) | (w3755 & ~w7187);
assign w1038 = w5250 & ~w1621;
assign w1039 = (~w502 & w1536) | (~w502 & w868) | (w1536 & w868);
assign w1040 = (~w5325 & w2992) | (~w5325 & w61) | (w2992 & w61);
assign w1041 = (~w1791 & w7444) | (~w1791 & w6675) | (w7444 & w6675);
assign w1042 = w5242 & ~w7552;
assign w1043 = w388 & w3254;
assign w1044 = w5005 & w6246;
assign w1045 = (w5344 & w1714) | (w5344 & w7556) | (w1714 & w7556);
assign w1046 = (~w1053 & w5229) | (~w1053 & w2029) | (w5229 & w2029);
assign w1047 = (~w5568 & ~w5803) | (~w5568 & w3333) | (~w5803 & w3333);
assign w1048 = (~w7513 & w3412) | (~w7513 & w2682) | (w3412 & w2682);
assign w1049 = ~w7210 & ~w2918;
assign w1050 = (~w4651 & w5553) | (~w4651 & w4999) | (w5553 & w4999);
assign w1051 = (w4932 & w2499) | (w4932 & ~w5484) | (w2499 & ~w5484);
assign w1052 = (w7168 & w1402) | (w7168 & w5291) | (w1402 & w5291);
assign w1053 = ~w4169 & ~w569;
assign w1054 = (w5007 & w2789) | (w5007 & w6639) | (w2789 & w6639);
assign w1055 = (w5178 & w4326) | (w5178 & w3098) | (w4326 & w3098);
assign w1056 = w2853 & w1356;
assign w1057 = a203 & b203;
assign w1058 = (w517 & w5912) | (w517 & w3074) | (w5912 & w3074);
assign w1059 = (~w4265 & w4209) | (~w4265 & w2876) | (w4209 & w2876);
assign w1060 = w3631 & w6235;
assign w1061 = (w3119 & w241) | (w3119 & w5319) | (w241 & w5319);
assign w1062 = w5604 & ~w1085;
assign w1063 = w1873 & w6174;
assign w1064 = (~w6325 & w686) | (~w6325 & w6475) | (w686 & w6475);
assign w1065 = (w7409 & w903) | (w7409 & ~w52) | (w903 & ~w52);
assign w1066 = w624 & ~w3312;
assign w1067 = ~w3896 & ~w7147;
assign w1068 = (w4574 & w713) | (w4574 & w6742) | (w713 & w6742);
assign w1069 = (w2627 & w3341) | (w2627 & w6068) | (w3341 & w6068);
assign w1070 = w6718 & w5337;
assign w1071 = ~w6392 & ~w7005;
assign w1072 = w4921 & w1732;
assign w1073 = ~w2119 & w1739;
assign w1074 = (~w1722 & w4287) | (~w1722 & w3748) | (w4287 & w3748);
assign w1075 = w6009 & ~w6816;
assign w1076 = ~w7513 & w6137;
assign w1077 = w5759 & ~w3741;
assign w1078 = (~w1427 & w4522) | (~w1427 & w3939) | (w4522 & w3939);
assign w1079 = (w1692 & w1262) | (w1692 & w2456) | (w1262 & w2456);
assign w1080 = ~w618 & ~w3064;
assign w1081 = ~w2339 & ~w3612;
assign w1082 = (w2563 & w799) | (w2563 & w6709) | (w799 & w6709);
assign w1083 = ~a63 & ~b63;
assign w1084 = (w3100 & w5189) | (w3100 & w641) | (w5189 & w641);
assign w1085 = a30 & b30;
assign w1086 = (~w6791 & w424) | (~w6791 & w3719) | (w424 & w3719);
assign w1087 = (~w5296 & w1373) | (~w5296 & w1905) | (w1373 & w1905);
assign w1088 = (~w1847 & w3793) | (~w1847 & w1850) | (w3793 & w1850);
assign w1089 = (~w4169 & w5594) | (~w4169 & ~w4768) | (w5594 & ~w4768);
assign w1090 = (~w3866 & w570) | (~w3866 & w3937) | (w570 & w3937);
assign w1091 = (w2806 & w5132) | (w2806 & w4144) | (w5132 & w4144);
assign w1092 = ~w7283 & ~w4061;
assign w1093 = ~w1565 & w4614;
assign w1094 = ~w4901 & w3292;
assign w1095 = (w2843 & w5974) | (w2843 & w3819) | (w5974 & w3819);
assign w1096 = w6965 & ~w7097;
assign w1097 = ~w3865 & ~w4752;
assign w1098 = ~w3167 & ~w4632;
assign w1099 = w2863 & ~w503;
assign w1100 = w273 & w681;
assign w1101 = w1230 | w1369;
assign w1102 = w1072 & w1732;
assign w1103 = (w6174 & w7226) | (w6174 & w3398) | (w7226 & w3398);
assign w1104 = (w3774 & w6030) | (w3774 & w7467) | (w6030 & w7467);
assign w1105 = ~w6683 & ~w1283;
assign w1106 = (~w7637 & w2550) | (~w7637 & w6370) | (w2550 & w6370);
assign w1107 = (w384 & ~w4346) | (w384 & ~w1868) | (~w4346 & ~w1868);
assign w1108 = (w5178 & w5245) | (w5178 & w5019) | (w5245 & w5019);
assign w1109 = ~w5987 & w3039;
assign w1110 = (~w2407 & w2141) | (~w2407 & w4958) | (w2141 & w4958);
assign w1111 = w6870 & ~w7399;
assign w1112 = (~w5325 & w7531) | (~w5325 & w5085) | (w7531 & w5085);
assign w1113 = ~w7635 & ~w6139;
assign w1114 = ~w1369 & w144;
assign w1115 = (w6593 & w2776) | (w6593 & ~w5098) | (w2776 & ~w5098);
assign w1116 = w1338 & ~w3953;
assign w1117 = (w3201 & w5619) | (w3201 & ~w6688) | (w5619 & ~w6688);
assign w1118 = ~w4906 & ~w5851;
assign w1119 = (w4926 & w5462) | (w4926 & ~w2013) | (w5462 & ~w2013);
assign w1120 = ~w7027 & ~w2993;
assign w1121 = w5395 & w5204;
assign w1122 = (w5974 & w7187) | (w5974 & w3767) | (w7187 & w3767);
assign w1123 = w3561 & w5788;
assign w1124 = w7566 & w5441;
assign w1125 = ~w6630 & ~w2519;
assign w1126 = (w5178 & w5157) | (w5178 & w4160) | (w5157 & w4160);
assign w1127 = (~w7216 & w5123) | (~w7216 & w4635) | (w5123 & w4635);
assign w1128 = (w4199 & w7238) | (w4199 & w5291) | (w7238 & w5291);
assign w1129 = ~w4967 & w2242;
assign w1130 = ~w2899 & ~w2901;
assign w1131 = ~w3669 & ~w278;
assign w1132 = ~w713 & w1643;
assign w1133 = (~w1925 & w1731) | (~w1925 & w1383) | (w1731 & w1383);
assign w1134 = (~w1463 & w3838) | (~w1463 & w7412) | (w3838 & w7412);
assign w1135 = ~w4788 & ~w1635;
assign w1136 = ~w2798 & w5223;
assign w1137 = ~a33 & ~b33;
assign w1138 = (w1161 & w3967) | (w1161 & ~w5759) | (w3967 & ~w5759);
assign w1139 = (~w3471 & w2641) | (~w3471 & w1182) | (w2641 & w1182);
assign w1140 = ~w2880 & ~w2611;
assign w1141 = (w4966 & w6525) | (w4966 & w1514) | (w6525 & w1514);
assign w1142 = ~w2728 & w2087;
assign w1143 = ~w5005 & ~w1837;
assign w1144 = w887 & ~w4564;
assign w1145 = ~w7219 & ~w5808;
assign w1146 = (~w1760 & w4634) | (~w1760 & ~w2209) | (w4634 & ~w2209);
assign w1147 = ~w7177 & w2393;
assign w1148 = (~w5178 & w2048) | (~w5178 & w16) | (w2048 & w16);
assign w1149 = ~w6836 & w1800;
assign w1150 = (w264 & w2653) | (w264 & w5583) | (w2653 & w5583);
assign w1151 = (~w6100 & w2640) | (~w6100 & w1711) | (w2640 & w1711);
assign w1152 = w3604 & ~w1884;
assign w1153 = w1622 & ~w505;
assign w1154 = (~w5178 & w4404) | (~w5178 & w4636) | (w4404 & w4636);
assign w1155 = (w3040 & w7286) | (w3040 & w3686) | (w7286 & w3686);
assign w1156 = (~w1722 & w7562) | (~w1722 & w3491) | (w7562 & w3491);
assign w1157 = ~w3312 & ~w3136;
assign w1158 = ~w1256 & ~w5287;
assign w1159 = ~w3928 & ~w5156;
assign w1160 = ~w381 & w6341;
assign w1161 = (~w7647 & w5404) | (~w7647 & w528) | (w5404 & w528);
assign w1162 = ~w6510 & ~w7188;
assign w1163 = (w6851 & w4529) | (w6851 & w5037) | (w4529 & w5037);
assign w1164 = w1555 & ~w1652;
assign w1165 = ~w3306 & w7216;
assign w1166 = (~w7205 & w6061) | (~w7205 & w266) | (w6061 & w266);
assign w1167 = (~w4337 & w3511) | (~w4337 & w2307) | (w3511 & w2307);
assign w1168 = (~w3490 & w2086) | (~w3490 & w4116) | (w2086 & w4116);
assign w1169 = ~w6643 & w3289;
assign w1170 = w1204 & ~w7493;
assign w1171 = ~w2127 & ~w5486;
assign w1172 = (w867 & w3103) | (w867 & w5917) | (w3103 & w5917);
assign w1173 = (w632 & w2417) | (w632 & w329) | (w2417 & w329);
assign w1174 = (~w2513 & w6668) | (~w2513 & w1879) | (w6668 & w1879);
assign w1175 = (w6151 & w646) | (w6151 & w5476) | (w646 & w5476);
assign w1176 = ~w3905 & ~w3392;
assign w1177 = w4697 & w7187;
assign w1178 = (~w1847 & w6759) | (~w1847 & w6874) | (w6759 & w6874);
assign w1179 = (w6945 & w2670) | (w6945 & w4460) | (w2670 & w4460);
assign w1180 = (~w2649 & w7031) | (~w2649 & ~w5403) | (w7031 & ~w5403);
assign w1181 = w2368 & ~w6654;
assign w1182 = ~w112 & ~w3471;
assign w1183 = ~w6354 & ~w3480;
assign w1184 = (~w5178 & w1669) | (~w5178 & w4766) | (w1669 & w4766);
assign w1185 = ~w7604 & w3819;
assign w1186 = (w7322 & w7340) | (w7322 & w4362) | (w7340 & w4362);
assign w1187 = ~w2671 & ~w4222;
assign w1188 = ~w6902 & ~w6204;
assign w1189 = w5665 & w5972;
assign w1190 = w3903 & w3203;
assign w1191 = (~w5178 & w1988) | (~w5178 & w6280) | (w1988 & w6280);
assign w1192 = w1576 & w7002;
assign w1193 = w3883 & ~w3819;
assign w1194 = ~w6437 & ~w5861;
assign w1195 = ~w6558 & ~w5862;
assign w1196 = a82 & b82;
assign w1197 = (~w1435 & w5819) | (~w1435 & ~w3105) | (w5819 & ~w3105);
assign w1198 = ~w5042 & w5627;
assign w1199 = (w5178 & w1688) | (w5178 & w5720) | (w1688 & w5720);
assign w1200 = ~w7137 & ~w5863;
assign w1201 = w4458 & ~w4759;
assign w1202 = w4697 & w3085;
assign w1203 = ~w7538 & ~w1171;
assign w1204 = ~w6054 & ~w1007;
assign w1205 = ~a195 & ~b195;
assign w1206 = ~w95 & w6708;
assign w1207 = (w1473 & w6179) | (w1473 & w1029) | (w6179 & w1029);
assign w1208 = ~w1588 & ~w6690;
assign w1209 = (w4892 & w6827) | (w4892 & w6177) | (w6827 & w6177);
assign w1210 = ~w5512 & w2105;
assign w1211 = (~w385 & w6211) | (~w385 & w2595) | (w6211 & w2595);
assign w1212 = (w2545 & ~w4102) | (w2545 & w5302) | (~w4102 & w5302);
assign w1213 = w1162 & ~w6324;
assign w1214 = w7310 & ~w5240;
assign w1215 = ~w7633 & w1435;
assign w1216 = a49 & b49;
assign w1217 = (~w7491 & w479) | (~w7491 & w5391) | (w479 & w5391);
assign w1218 = (w3104 & w704) | (w3104 & ~w6100) | (w704 & ~w6100);
assign w1219 = (w4889 & w6733) | (w4889 & w4868) | (w6733 & w4868);
assign w1220 = w2598 & ~w3058;
assign w1221 = ~w965 & w3505;
assign w1222 = w3924 & ~w3354;
assign w1223 = (w7542 & w549) | (w7542 & w563) | (w549 & w563);
assign w1224 = (~w7604 & w299) | (~w7604 & ~w139) | (w299 & ~w139);
assign w1225 = (w5222 & w3301) | (w5222 & w6633) | (w3301 & w6633);
assign w1226 = ~w7575 & w6486;
assign w1227 = ~w7142 & ~w3997;
assign w1228 = ~w999 & ~w6342;
assign w1229 = (w5554 & w7528) | (w5554 & w2485) | (w7528 & w2485);
assign w1230 = w6520 & w1369;
assign w1231 = w1204 & ~w13;
assign w1232 = ~w5674 & w1324;
assign w1233 = (~w6149 & w6254) | (~w6149 & w1546) | (w6254 & w1546);
assign w1234 = ~w3266 & ~w5950;
assign w1235 = (w6614 & w7570) | (w6614 & w2661) | (w7570 & w2661);
assign w1236 = (~w303 & w4913) | (~w303 & w1087) | (w4913 & w1087);
assign w1237 = w1937 & ~w6685;
assign w1238 = (w6018 & w1091) | (w6018 & w3119) | (w1091 & w3119);
assign w1239 = w4777 & w4905;
assign w1240 = w2311 & w2324;
assign w1241 = ~a13 & ~b13;
assign w1242 = (~w5257 & w7094) | (~w5257 & w5311) | (w7094 & w5311);
assign w1243 = (w5655 & w4559) | (w5655 & w83) | (w4559 & w83);
assign w1244 = ~w4994 & ~w7589;
assign w1245 = w6281 & ~w390;
assign w1246 = (w7414 & ~w2526) | (w7414 & w840) | (~w2526 & w840);
assign w1247 = ~w6766 & ~w3934;
assign w1248 = ~w4242 & w7305;
assign w1249 = (w5146 & w6275) | (w5146 & w484) | (w6275 & w484);
assign w1250 = ~w3248 & ~w57;
assign w1251 = (~w3014 & w2830) | (~w3014 & ~w3903) | (w2830 & ~w3903);
assign w1252 = ~a245 & ~b245;
assign w1253 = ~w1491 & ~w2554;
assign w1254 = w3556 & ~w3224;
assign w1255 = ~w2506 & w7273;
assign w1256 = ~a155 & ~b155;
assign w1257 = (w6253 & w2161) | (w6253 & w5391) | (w2161 & w5391);
assign w1258 = w1831 & w6225;
assign w1259 = (w3821 & w169) | (w3821 & w181) | (w169 & w181);
assign w1260 = ~w4545 & w4884;
assign w1261 = w3880 & w4790;
assign w1262 = (w1692 & w5575) | (w1692 & ~w5385) | (w5575 & ~w5385);
assign w1263 = ~w60 & ~w6463;
assign w1264 = w1743 | w3989;
assign w1265 = w2216 & ~w5350;
assign w1266 = ~w3591 & w926;
assign w1267 = ~w1632 & ~w3285;
assign w1268 = ~w600 & ~w3764;
assign w1269 = (~w3461 & w6579) | (~w3461 & w5452) | (w6579 & w5452);
assign w1270 = ~w757 & ~w1468;
assign w1271 = ~w7634 & w3430;
assign w1272 = w2803 & ~w1974;
assign w1273 = (~w6100 & w4100) | (~w6100 & w6543) | (w4100 & w6543);
assign w1274 = (w5178 & w6782) | (w5178 & w1702) | (w6782 & w1702);
assign w1275 = ~w7453 & w5394;
assign w1276 = ~w3207 & w4717;
assign w1277 = (w3472 & w2886) | (w3472 & w5325) | (w2886 & w5325);
assign w1278 = w5385 & w5200;
assign w1279 = a84 & b84;
assign w1280 = w7506 & w4132;
assign w1281 = ~w4457 & w1655;
assign w1282 = (~w523 & w1456) | (~w523 & w2006) | (w1456 & w2006);
assign w1283 = ~w5743 & ~w4174;
assign w1284 = ~w804 & ~w2005;
assign w1285 = a68 & b68;
assign w1286 = (w5178 & w2181) | (w5178 & w6934) | (w2181 & w6934);
assign w1287 = w4347 & w4237;
assign w1288 = ~w7219 & ~w6811;
assign w1289 = (w5963 & w1502) | (w5963 & ~w813) | (w1502 & ~w813);
assign w1290 = w1196 & ~w5881;
assign w1291 = (~w2996 & w2727) | (~w2996 & w6606) | (w2727 & w6606);
assign w1292 = ~w6994 & w984;
assign w1293 = w7225 & w1834;
assign w1294 = w1018 & w3110;
assign w1295 = w3282 & ~w5781;
assign w1296 = (w3060 & w5312) | (w3060 & w2456) | (w5312 & w2456);
assign w1297 = w5767 & w7364;
assign w1298 = ~w2453 & ~w435;
assign w1299 = w7150 & ~w3345;
assign w1300 = a66 & b66;
assign w1301 = ~w3045 & w3805;
assign w1302 = ~w706 & ~w4149;
assign w1303 = ~w6849 & w169;
assign w1304 = ~w7527 & ~w1285;
assign w1305 = (w3727 & w6410) | (w3727 & w5304) | (w6410 & w5304);
assign w1306 = w6994 & ~w761;
assign w1307 = ~w3706 & ~w2872;
assign w1308 = ~w1266 & w4101;
assign w1309 = ~w6181 & ~w4400;
assign w1310 = (w1155 & w2510) | (w1155 & ~w7383) | (w2510 & ~w7383);
assign w1311 = ~w1443 & w808;
assign w1312 = (w1284 & w6537) | (w1284 & ~w512) | (w6537 & ~w512);
assign w1313 = (~w5066 & w2178) | (~w5066 & w1607) | (w2178 & w1607);
assign w1314 = w5948 & w3370;
assign w1315 = ~w2124 & w7329;
assign w1316 = (~w6626 & ~w2333) | (~w6626 & w1615) | (~w2333 & w1615);
assign w1317 = (w6499 & w2810) | (w6499 & w5511) | (w2810 & w5511);
assign w1318 = ~w1878 & ~w7008;
assign w1319 = (w5225 & w3410) | (w5225 & ~w7015) | (w3410 & ~w7015);
assign w1320 = ~w6999 & w1973;
assign w1321 = ~w4967 & w5362;
assign w1322 = w5066 & w3122;
assign w1323 = ~w6304 & w6922;
assign w1324 = ~w2914 & w1682;
assign w1325 = (w5871 & w579) | (w5871 & w1051) | (w579 & w1051);
assign w1326 = ~w2872 & w6184;
assign w1327 = a14 & b14;
assign w1328 = ~w3514 & w1093;
assign w1329 = (~w5881 & w1290) | (~w5881 & w6237) | (w1290 & w6237);
assign w1330 = w5756 & w3570;
assign w1331 = w6415 & w3321;
assign w1332 = (w3490 & w4956) | (w3490 & w6345) | (w4956 & w6345);
assign w1333 = (w5972 & w453) | (w5972 & w1189) | (w453 & w1189);
assign w1334 = ~w443 & w5345;
assign w1335 = (w3284 & w2694) | (w3284 & w7637) | (w2694 & w7637);
assign w1336 = (~w5944 & w5022) | (~w5944 & w824) | (w5022 & w824);
assign w1337 = (~w1936 & w2167) | (~w1936 & w7557) | (w2167 & w7557);
assign w1338 = (~w2112 & w1322) | (~w2112 & w3436) | (w1322 & w3436);
assign w1339 = w7024 & w2097;
assign w1340 = (w3057 & w768) | (w3057 & w696) | (w768 & w696);
assign w1341 = (w927 & w3365) | (w927 & w4894) | (w3365 & w4894);
assign w1342 = (w808 & w7442) | (w808 & w1129) | (w7442 & w1129);
assign w1343 = ~w5926 & ~w6839;
assign w1344 = w1759 & ~w1554;
assign w1345 = ~a1 & ~b1;
assign w1346 = ~w2913 & w3616;
assign w1347 = (~w7268 & w2418) | (~w7268 & w4106) | (w2418 & w4106);
assign w1348 = ~w2471 & ~w36;
assign w1349 = ~w790 & w593;
assign w1350 = w70 & w6894;
assign w1351 = w6704 & ~w2199;
assign w1352 = ~w2596 & w7530;
assign w1353 = w1601 & w7644;
assign w1354 = ~w1759 & w3062;
assign w1355 = (w6872 & w1856) | (w6872 & w4122) | (w1856 & w4122);
assign w1356 = w7188 & ~w6571;
assign w1357 = (w3681 & w3555) | (w3681 & w5655) | (w3555 & w5655);
assign w1358 = (~w5178 & w2323) | (~w5178 & w5957) | (w2323 & w5957);
assign w1359 = (w5659 & w5672) | (w5659 & w5637) | (w5672 & w5637);
assign w1360 = ~w4918 & ~w7424;
assign w1361 = (w2660 & w5661) | (w2660 & ~w139) | (w5661 & ~w139);
assign w1362 = (w5325 & w6576) | (w5325 & w2231) | (w6576 & w2231);
assign w1363 = w2078 & ~w3108;
assign w1364 = ~w3551 & w4651;
assign w1365 = w6353 & w2082;
assign w1366 = w2210 & w4090;
assign w1367 = (~w5442 & w6451) | (~w5442 & w1678) | (w6451 & w1678);
assign w1368 = ~w4967 & w1819;
assign w1369 = ~w195 & ~w2888;
assign w1370 = (w5325 & w4316) | (w5325 & w3635) | (w4316 & w3635);
assign w1371 = a239 & b239;
assign w1372 = ~w7471 & ~w6876;
assign w1373 = w2880 & ~w5296;
assign w1374 = w1587 & w2388;
assign w1375 = (w2123 & w4792) | (w2123 & w1178) | (w4792 & w1178);
assign w1376 = (w303 & w4181) | (w303 & w7009) | (w4181 & w7009);
assign w1377 = w4185 & ~w4940;
assign w1378 = ~w6791 & w814;
assign w1379 = (~w618 & w4550) | (~w618 & w633) | (w4550 & w633);
assign w1380 = ~w2978 & ~w3140;
assign w1381 = w3660 & ~w461;
assign w1382 = ~w356 & ~w4026;
assign w1383 = w1377 | ~w4940;
assign w1384 = ~w6169 & ~w5864;
assign w1385 = ~w756 & ~w5105;
assign w1386 = ~a174 & ~b174;
assign w1387 = w5930 & ~w7005;
assign w1388 = w4145 & ~w7520;
assign w1389 = ~w1901 & ~w3256;
assign w1390 = w7500 & ~w7414;
assign w1391 = (w2123 & w2060) | (w2123 & w5125) | (w2060 & w5125);
assign w1392 = (~w729 & w466) | (~w729 & w3504) | (w466 & w3504);
assign w1393 = (~w5655 & w244) | (~w5655 & w416) | (w244 & w416);
assign w1394 = ~w7631 & ~w7317;
assign w1395 = (~w3774 & w7476) | (~w3774 & w920) | (w7476 & w920);
assign w1396 = w6151 & w865;
assign w1397 = ~w1570 & ~w2376;
assign w1398 = w2216 & ~w5121;
assign w1399 = (~w5888 & ~w1587) | (~w5888 & w399) | (~w1587 & w399);
assign w1400 = (~w5362 & w6852) | (~w5362 & w3139) | (w6852 & w3139);
assign w1401 = (w2097 & w2857) | (w2097 & w108) | (w2857 & w108);
assign w1402 = (w6535 & w1674) | (w6535 & w4199) | (w1674 & w4199);
assign w1403 = (~w4286 & w6734) | (~w4286 & w6595) | (w6734 & w6595);
assign w1404 = ~w3597 & w5189;
assign w1405 = ~w1660 & w3291;
assign w1406 = (~w3989 & w3848) | (~w3989 & w577) | (w3848 & w577);
assign w1407 = (w4433 & w4164) | (w4433 & w4400) | (w4164 & w4400);
assign w1408 = (w681 & w5800) | (w681 & w1321) | (w5800 & w1321);
assign w1409 = w3044 & ~w4388;
assign w1410 = (w1254 & ~w7197) | (w1254 & w3556) | (~w7197 & w3556);
assign w1411 = w1364 & ~w4999;
assign w1412 = w6760 & ~w3267;
assign w1413 = w1080 & w1107;
assign w1414 = ~w6181 & ~w7575;
assign w1415 = (w5298 & w6052) | (w5298 & ~w2453) | (w6052 & ~w2453);
assign w1416 = (w3318 & w4983) | (w3318 & w4676) | (w4983 & w4676);
assign w1417 = (w1097 & w1872) | (w1097 & w3330) | (w1872 & w3330);
assign w1418 = (w76 & w7646) | (w76 & ~w6216) | (w7646 & ~w6216);
assign w1419 = (~w625 & w6844) | (~w625 & w927) | (w6844 & w927);
assign w1420 = ~w5480 & ~w5467;
assign w1421 = w3107 & w3157;
assign w1422 = (w2285 & w1785) | (w2285 & w3644) | (w1785 & w3644);
assign w1423 = (w3447 & w7281) | (w3447 & w4050) | (w7281 & w4050);
assign w1424 = (~w2515 & w7629) | (~w2515 & w913) | (w7629 & w913);
assign w1425 = (w7647 & w1518) | (w7647 & w1985) | (w1518 & w1985);
assign w1426 = (w777 & w2733) | (w777 & w3295) | (w2733 & w3295);
assign w1427 = ~w5059 & ~w2066;
assign w1428 = ~w4474 & w3720;
assign w1429 = ~w6169 & ~w6571;
assign w1430 = ~w3009 & w7034;
assign w1431 = ~a17 & ~b17;
assign w1432 = w4428 & w3144;
assign w1433 = (~w777 & w5023) | (~w777 & w6665) | (w5023 & w6665);
assign w1434 = w4843 & w931;
assign w1435 = ~w3932 & ~w3689;
assign w1436 = ~w4872 & ~w4371;
assign w1437 = w3664 & w6857;
assign w1438 = w2506 & ~w7273;
assign w1439 = (~w5178 & w4821) | (~w5178 & w2665) | (w4821 & w2665);
assign w1440 = ~w261 & ~w960;
assign w1441 = ~a28 & ~b28;
assign w1442 = ~w4922 & ~w4251;
assign w1443 = a178 & b178;
assign w1444 = w4966 & ~w5194;
assign w1445 = (w5178 & w2422) | (w5178 & w3794) | (w2422 & w3794);
assign w1446 = w3119 & w448;
assign w1447 = w4963 & w1907;
assign w1448 = ~w1288 & ~w1175;
assign w1449 = (w1736 & w3224) | (w1736 & w5678) | (w3224 & w5678);
assign w1450 = (w5257 & w6464) | (w5257 & w15) | (w6464 & w15);
assign w1451 = w351 & ~w656;
assign w1452 = ~w385 & ~w1591;
assign w1453 = (w7506 & w3057) | (w7506 & w4925) | (w3057 & w4925);
assign w1454 = w6990 & w7344;
assign w1455 = ~w2 & ~w7408;
assign w1456 = w3248 & ~w523;
assign w1457 = w651 & ~w1143;
assign w1458 = ~w723 & w6224;
assign w1459 = (w3929 & w1822) | (w3929 & ~w3868) | (w1822 & ~w3868);
assign w1460 = ~w3753 & ~w1583;
assign w1461 = ~w6100 & w5967;
assign w1462 = (w1076 & w923) | (w1076 & w6501) | (w923 & w6501);
assign w1463 = a208 & b208;
assign w1464 = (w777 & w3030) | (w777 & w3261) | (w3030 & w3261);
assign w1465 = (w735 & w5750) | (w735 & ~w5430) | (w5750 & ~w5430);
assign w1466 = ~w6103 & ~w2233;
assign w1467 = (~w3771 & ~w2409) | (~w3771 & w5871) | (~w2409 & w5871);
assign w1468 = (w3057 & w1173) | (w3057 & w627) | (w1173 & w627);
assign w1469 = (w632 & w568) | (w632 & w5258) | (w568 & w5258);
assign w1470 = ~w6200 & w50;
assign w1471 = a47 & b47;
assign w1472 = ~w390 & ~w7020;
assign w1473 = (~w1343 & w907) | (~w1343 & w6600) | (w907 & w6600);
assign w1474 = (~w3760 & w2287) | (~w3760 & w5618) | (w2287 & w5618);
assign w1475 = w4074 & ~w2104;
assign w1476 = (~w1135 & w5456) | (~w1135 & w1775) | (w5456 & w1775);
assign w1477 = w5241 & ~w6656;
assign w1478 = (w3658 & w591) | (w3658 & w883) | (w591 & w883);
assign w1479 = ~w2127 & ~w7265;
assign w1480 = (w550 & w3414) | (w550 & w6148) | (w3414 & w6148);
assign w1481 = (w4283 & w6269) | (w4283 & ~w563) | (w6269 & ~w563);
assign w1482 = (w6942 & w6148) | (w6942 & w4290) | (w6148 & w4290);
assign w1483 = (w2142 & w4602) | (w2142 & w6547) | (w4602 & w6547);
assign w1484 = (~w7197 & w165) | (~w7197 & w6338) | (w165 & w6338);
assign w1485 = w2803 & ~w3607;
assign w1486 = (w2683 & w3445) | (w2683 & w6957) | (w3445 & w6957);
assign w1487 = w4025 & ~w5914;
assign w1488 = w5600 & ~w2243;
assign w1489 = ~w937 & ~w4898;
assign w1490 = w1751 & w3488;
assign w1491 = (w6100 & w6130) | (w6100 & w4406) | (w6130 & w4406);
assign w1492 = ~w7291 & w1208;
assign w1493 = w2995 & w6174;
assign w1494 = w320 & w1892;
assign w1495 = (~w6450 & w6592) | (~w6450 & w4675) | (w6592 & w4675);
assign w1496 = (w5520 & w1690) | (w5520 & w6873) | (w1690 & w6873);
assign w1497 = ~w3212 & ~w5219;
assign w1498 = cin & ~w4606;
assign w1499 = (~w4033 & w4068) | (~w4033 & w2710) | (w4068 & w2710);
assign w1500 = ~w7566 & w1328;
assign w1501 = w1827 & ~w1722;
assign w1502 = (~w2603 & w2553) | (~w2603 & w889) | (w2553 & w889);
assign w1503 = ~w5965 & w5447;
assign w1504 = (w5089 & w6434) | (w5089 & w4862) | (w6434 & w4862);
assign w1505 = w4271 & w1762;
assign w1506 = w3062 & ~w3139;
assign w1507 = w1892 & w320;
assign w1508 = (w3070 & ~w3212) | (w3070 & ~w4123) | (~w3212 & ~w4123);
assign w1509 = (w2792 & w3986) | (w2792 & w1593) | (w3986 & w1593);
assign w1510 = (~w665 & w4551) | (~w665 & w6955) | (w4551 & w6955);
assign w1511 = ~w2173 & ~w3771;
assign w1512 = ~w2740 & w1939;
assign w1513 = ~w6927 & w2998;
assign w1514 = ~w5555 & w5778;
assign w1515 = ~w6992 & ~w2880;
assign w1516 = w4901 & ~w5770;
assign w1517 = ~w1416 & ~w3833;
assign w1518 = (w1328 & w7483) | (w1328 & w4299) | (w7483 & w4299);
assign w1519 = (~w2913 & w6608) | (~w2913 & w1346) | (w6608 & w1346);
assign w1520 = w1455 & w7266;
assign w1521 = w3210 & w2712;
assign w1522 = (w1724 & w419) | (w1724 & ~w5611) | (w419 & ~w5611);
assign w1523 = w2116 & ~w7161;
assign w1524 = (~w5178 & w5280) | (~w5178 & w515) | (w5280 & w515);
assign w1525 = (w3467 & w478) | (w3467 & w3943) | (w478 & w3943);
assign w1526 = w54 & ~w2179;
assign w1527 = w6458 & w7394;
assign w1528 = w5259 & w3449;
assign w1529 = ~w4976 & w1760;
assign w1530 = ~w478 & w7267;
assign w1531 = (w144 & w2087) | (w144 & w316) | (w2087 & w316);
assign w1532 = a27 & b27;
assign w1533 = w3840 & ~w7391;
assign w1534 = (~w1463 & w2820) | (~w1463 & w1632) | (w2820 & w1632);
assign w1535 = (w5196 & w1699) | (w5196 & w1970) | (w1699 & w1970);
assign w1536 = ~w4806 & ~w502;
assign w1537 = w1937 & ~w7512;
assign w1538 = (w3774 & w5124) | (w3774 & w1623) | (w5124 & w1623);
assign w1539 = w3045 & ~w3805;
assign w1540 = ~w4143 & w1507;
assign w1541 = w6458 & ~w3328;
assign w1542 = ~w7137 & w968;
assign w1543 = (w3909 & ~w3730) | (w3909 & ~w100) | (~w3730 & ~w100);
assign w1544 = ~a9 & ~b9;
assign w1545 = ~w2836 & w3306;
assign w1546 = (~w6149 & w6046) | (~w6149 & w3142) | (w6046 & w3142);
assign w1547 = w6500 & w4196;
assign w1548 = (~w3176 & w850) | (~w3176 & w2511) | (w850 & w2511);
assign w1549 = ~w931 & ~w5760;
assign w1550 = a226 & b226;
assign w1551 = (~w4296 & w203) | (~w4296 & w2702) | (w203 & w2702);
assign w1552 = w5478 & w5628;
assign w1553 = (w629 & w7252) | (w629 & w5208) | (w7252 & w5208);
assign w1554 = ~w6181 & w2654;
assign w1555 = ~w5525 & w1833;
assign w1556 = w7493 & ~w2648;
assign w1557 = w6244 & ~w2718;
assign w1558 = ~w1798 & w3582;
assign w1559 = (w4969 & w4243) | (w4969 & w2656) | (w4243 & w2656);
assign w1560 = ~w2353 & w7073;
assign w1561 = (w2123 & w6229) | (w2123 & w1088) | (w6229 & w1088);
assign w1562 = ~w2329 & ~w6387;
assign w1563 = a133 & b133;
assign w1564 = (w401 & w5761) | (w401 & w2097) | (w5761 & w2097);
assign w1565 = ~w1728 & w2463;
assign w1566 = (w1774 & w5026) | (w1774 & ~w4258) | (w5026 & ~w4258);
assign w1567 = (w5178 & w1597) | (w5178 & w6306) | (w1597 & w6306);
assign w1568 = (w3318 & w4391) | (w3318 & w1806) | (w4391 & w1806);
assign w1569 = (~w3318 & w1744) | (~w3318 & w1404) | (w1744 & w1404);
assign w1570 = ~w5557 & ~w2519;
assign w1571 = (~w7291 & w7147) | (~w7291 & w5738) | (w7147 & w5738);
assign w1572 = (w5325 & w41) | (w5325 & w2331) | (w41 & w2331);
assign w1573 = (w639 & w3871) | (w639 & w5724) | (w3871 & w5724);
assign w1574 = (~w5416 & w4533) | (~w5416 & w4761) | (w4533 & w4761);
assign w1575 = ~w3092 & ~w1200;
assign w1576 = ~w3007 & w6427;
assign w1577 = w6706 & ~w6257;
assign w1578 = (w6372 & w1844) | (w6372 & ~w4521) | (w1844 & ~w4521);
assign w1579 = (~w5178 & w5079) | (~w5178 & w606) | (w5079 & w606);
assign w1580 = ~a135 & ~b135;
assign w1581 = w5058 & w5934;
assign w1582 = (w6100 & w3220) | (w6100 & w1172) | (w3220 & w1172);
assign w1583 = (~w5178 & w5650) | (~w5178 & w1686) | (w5650 & w1686);
assign w1584 = w929 | w3431;
assign w1585 = (~w3318 & w6135) | (~w3318 & w2198) | (w6135 & w2198);
assign w1586 = (w3774 & w3121) | (w3774 & w4137) | (w3121 & w4137);
assign w1587 = w1131 & w2129;
assign w1588 = ~a122 & ~b122;
assign w1589 = ~w5721 & ~w5996;
assign w1590 = w4132 & ~w4123;
assign w1591 = a222 & b222;
assign w1592 = (~w6353 & w6364) | (~w6353 & w2383) | (w6364 & w2383);
assign w1593 = (w2792 & w4393) | (w2792 & ~w7187) | (w4393 & ~w7187);
assign w1594 = ~w4330 & ~w4530;
assign w1595 = w3437 & w3528;
assign w1596 = w5026 | w1774;
assign w1597 = (~w588 & w4125) | (~w588 & w7468) | (w4125 & w7468);
assign w1598 = ~w5402 & w4430;
assign w1599 = ~w210 & ~w3326;
assign w1600 = (w1936 & w4109) | (w1936 & w3563) | (w4109 & w3563);
assign w1601 = ~a31 & ~b31;
assign w1602 = ~w4045 & w2536;
assign w1603 = (~w6450 & w6592) | (~w6450 & w856) | (w6592 & w856);
assign w1604 = (~w3868 & w4451) | (~w3868 & ~w3396) | (w4451 & ~w3396);
assign w1605 = ~w6331 & ~w1580;
assign w1606 = ~w504 & w2819;
assign w1607 = ~w5958 & w1455;
assign w1608 = ~w1607 & ~w3953;
assign w1609 = (~w6714 & ~w4479) | (~w6714 & w3642) | (~w4479 & w3642);
assign w1610 = a253 & b253;
assign w1611 = (~w4191 & w6819) | (~w4191 & w2498) | (w6819 & w2498);
assign w1612 = (~w3113 & w5830) | (~w3113 & w3468) | (w5830 & w3468);
assign w1613 = (w5257 & w3588) | (w5257 & w292) | (w3588 & w292);
assign w1614 = w390 & ~w624;
assign w1615 = w5163 & ~w6626;
assign w1616 = (w7397 & w3951) | (w7397 & w4224) | (w3951 & w4224);
assign w1617 = ~w7137 & w468;
assign w1618 = w6640 & ~w5172;
assign w1619 = (w409 & w4213) | (w409 & w1770) | (w4213 & w1770);
assign w1620 = w3219 & ~w7592;
assign w1621 = a80 & b80;
assign w1622 = a177 & b177;
assign w1623 = (~w2985 & w1803) | (~w2985 & w5351) | (w1803 & w5351);
assign w1624 = (~w6082 & w862) | (~w6082 & w3592) | (w862 & w3592);
assign w1625 = (~w7205 & w1237) | (~w7205 & w3605) | (w1237 & w3605);
assign w1626 = (w7158 & w2708) | (w7158 & w2396) | (w2708 & w2396);
assign w1627 = ~w2969 & w6251;
assign w1628 = (w3719 & ~w7576) | (w3719 & w809) | (~w7576 & w809);
assign w1629 = ~w1792 & ~w3587;
assign w1630 = ~w5005 & ~w6246;
assign w1631 = ~w2090 & w3063;
assign w1632 = ~a207 & ~b207;
assign w1633 = (~w5344 & w2248) | (~w5344 & w2544) | (w2248 & w2544);
assign w1634 = ~w998 & w4266;
assign w1635 = a242 & b242;
assign w1636 = w3512 & ~w3758;
assign w1637 = ~w3152 & w2850;
assign w1638 = (w6082 & w6234) | (w6082 & w6778) | (w6234 & w6778);
assign w1639 = ~w4681 & w2503;
assign w1640 = (~w1670 & w6652) | (~w1670 & w2031) | (w6652 & w2031);
assign w1641 = ~w444 & w6879;
assign w1642 = w4130 & ~w2582;
assign w1643 = ~w7271 & ~w4574;
assign w1644 = w1044 | w6246;
assign w1645 = ~w4698 & ~w4944;
assign w1646 = (w2563 & w3268) | (w2563 & ~w5962) | (w3268 & ~w5962);
assign w1647 = ~w4843 & w1723;
assign w1648 = (~w2124 & w1363) | (~w2124 & w1968) | (w1363 & w1968);
assign w1649 = (w506 & w830) | (w506 & w3470) | (w830 & w3470);
assign w1650 = (~w6032 & w7063) | (~w6032 & w997) | (w7063 & w997);
assign w1651 = ~w7371 & w340;
assign w1652 = ~w3014 & ~w247;
assign w1653 = (w3939 & w7131) | (w3939 & ~w5403) | (w7131 & ~w5403);
assign w1654 = w121 & w5192;
assign w1655 = ~w6087 & ~w4467;
assign w1656 = ~a243 & ~b243;
assign w1657 = (w412 & w4666) | (w412 & w430) | (w4666 & w430);
assign w1658 = ~w4107 & ~w2261;
assign w1659 = w7342 & ~w6965;
assign w1660 = ~w4602 & w3880;
assign w1661 = a176 & b176;
assign w1662 = w1630 & ~w6580;
assign w1663 = (~w3113 & w5830) | (~w3113 & w4175) | (w5830 & w4175);
assign w1664 = (~w777 & w3621) | (~w777 & w6930) | (w3621 & w6930);
assign w1665 = w7283 & ~w1389;
assign w1666 = (w500 & w7079) | (w500 & w6016) | (w7079 & w6016);
assign w1667 = (w6100 & w589) | (w6100 & w3305) | (w589 & w3305);
assign w1668 = ~w4526 & ~w4875;
assign w1669 = (w4143 & w5224) | (w4143 & w871) | (w5224 & w871);
assign w1670 = ~w3669 & ~w2990;
assign w1671 = (w3986 & w1146) | (w3986 & w6266) | (w1146 & w6266);
assign w1672 = (~w2065 & w3579) | (~w2065 & w7359) | (w3579 & w7359);
assign w1673 = ~w3240 & w902;
assign w1674 = ~w2990 & w4437;
assign w1675 = ~w3679 & w3384;
assign w1676 = w4598 & w5408;
assign w1677 = w7222 & ~w3433;
assign w1678 = (~w5442 & w642) | (~w5442 & w2479) | (w642 & w2479);
assign w1679 = w3573 & ~w1532;
assign w1680 = (~w4510 & w5521) | (~w4510 & w7377) | (w5521 & w7377);
assign w1681 = (w1886 & w4453) | (w1886 & w6048) | (w4453 & w6048);
assign w1682 = ~w3137 & ~w7522;
assign w1683 = (~w5404 & w5821) | (~w5404 & w4299) | (w5821 & w4299);
assign w1684 = w3277 | w6248;
assign w1685 = (~w7183 & w2407) | (~w7183 & w2192) | (w2407 & w2192);
assign w1686 = (w5895 & w1908) | (w5895 & ~w5325) | (w1908 & ~w5325);
assign w1687 = (~w5257 & w5976) | (~w5257 & w3898) | (w5976 & w3898);
assign w1688 = (~w2548 & ~w103) | (~w2548 & w2061) | (~w103 & w2061);
assign w1689 = (w2456 & w4836) | (w2456 & w6321) | (w4836 & w6321);
assign w1690 = (~w3953 & w5520) | (~w3953 & w4851) | (w5520 & w4851);
assign w1691 = w6779 & ~w7604;
assign w1692 = ~w937 & ~w5745;
assign w1693 = (w2104 & ~w4074) | (w2104 & ~w3736) | (~w4074 & ~w3736);
assign w1694 = (w5655 & w3698) | (w5655 & w7119) | (w3698 & w7119);
assign w1695 = (w5567 & w6763) | (w5567 & w3391) | (w6763 & w3391);
assign w1696 = (w5528 & w6403) | (w5528 & w2477) | (w6403 & w2477);
assign w1697 = (w6100 & w631) | (w6100 & w6598) | (w631 & w6598);
assign w1698 = (~w3224 & ~w7197) | (~w3224 & w6645) | (~w7197 & w6645);
assign w1699 = ~w783 | ~w5346;
assign w1700 = (w3727 & w6410) | (w3727 & w6152) | (w6410 & w6152);
assign w1701 = ~w2221 & w2343;
assign w1702 = (w3952 & w2252) | (w3952 & w5518) | (w2252 & w5518);
assign w1703 = (~w7491 & w479) | (~w7491 & w6385) | (w479 & w6385);
assign w1704 = ~w2124 & w3047;
assign w1705 = ~w1148 & ~w2015;
assign w1706 = w2420 & w1006;
assign w1707 = (w686 & w3958) | (w686 & w4044) | (w3958 & w4044);
assign w1708 = w7013 & w342;
assign w1709 = ~w1252 & ~w6774;
assign w1710 = (~w714 & ~w2083) | (~w714 & ~w5368) | (~w2083 & ~w5368);
assign w1711 = (w7529 & w1659) | (w7529 & ~w3303) | (w1659 & ~w3303);
assign w1712 = a173 & b173;
assign w1713 = ~w5783 & w2617;
assign w1714 = w4503 & ~w4457;
assign w1715 = w7327 & ~w5223;
assign w1716 = w6381 & w3440;
assign w1717 = (~w4169 & w5594) | (~w4169 & ~w6577) | (w5594 & ~w6577);
assign w1718 = ~w5759 & w833;
assign w1719 = (~w2471 & ~w6462) | (~w2471 & w1763) | (~w6462 & w1763);
assign w1720 = ~w4906 & ~w671;
assign w1721 = w6255 & ~w6716;
assign w1722 = ~w3869 & ~w2751;
assign w1723 = ~w226 & w6582;
assign w1724 = ~w6354 & w7480;
assign w1725 = ~w6520 & ~w2888;
assign w1726 = w4747 & ~w2966;
assign w1727 = ~w5783 & w1769;
assign w1728 = ~w6375 & w3426;
assign w1729 = ~w1498 & ~w2058;
assign w1730 = (w3063 & w1631) | (w3063 & w7015) | (w1631 & w7015);
assign w1731 = w5170 & ~w1925;
assign w1732 = ~w4238 & ~w4377;
assign w1733 = (w2123 & w1920) | (w2123 & w7515) | (w1920 & w7515);
assign w1734 = w7294 & ~w5635;
assign w1735 = ~w5496 & w7214;
assign w1736 = w7044 & ~w2725;
assign w1737 = w313 & ~w32;
assign w1738 = ~w6117 & ~w4602;
assign w1739 = ~w1866 & ~w2253;
assign w1740 = ~w1541 & ~w6025;
assign w1741 = w2104 & ~w57;
assign w1742 = w2861 & w5778;
assign w1743 = ~w147 & w1247;
assign w1744 = (w2399 & w311) | (w2399 & w1084) | (w311 & w1084);
assign w1745 = w601 & ~w5879;
assign w1746 = w360 | w4517;
assign w1747 = ~w757 & ~w2097;
assign w1748 = w984 & ~w806;
assign w1749 = (w1355 & ~w5325) | (w1355 & w1916) | (~w5325 & w1916);
assign w1750 = (w5178 & w4683) | (w5178 & w6175) | (w4683 & w6175);
assign w1751 = ~w4669 & w4895;
assign w1752 = w681 & w4341;
assign w1753 = ~a56 & ~b56;
assign w1754 = ~w6683 & ~w4174;
assign w1755 = (w5078 & w4290) | (w5078 & w6913) | (w4290 & w6913);
assign w1756 = a168 & b168;
assign w1757 = ~w5937 & w437;
assign w1758 = ~w1455 & w7106;
assign w1759 = ~w3192 & ~w4297;
assign w1760 = ~w4242 & ~w4448;
assign w1761 = (~w2273 & w5409) | (~w2273 & w3038) | (w5409 & w3038);
assign w1762 = (~w4458 & w1281) | (~w4458 & w6406) | (w1281 & w6406);
assign w1763 = w195 & ~w2471;
assign w1764 = ~w4143 & w4313;
assign w1765 = ~w3223 & ~w998;
assign w1766 = (~w2909 & w6931) | (~w2909 & w4820) | (w6931 & w4820);
assign w1767 = (~w2847 & w3760) | (~w2847 & w6411) | (w3760 & w6411);
assign w1768 = ~w6114 & w518;
assign w1769 = w1757 & ~w2590;
assign w1770 = (w2429 & w1516) | (w2429 & w3983) | (w1516 & w3983);
assign w1771 = (w409 & w4213) | (w409 & w5395) | (w4213 & w5395);
assign w1772 = ~w1832 & ~w3978;
assign w1773 = (w3444 & w2226) | (w3444 & w7581) | (w2226 & w7581);
assign w1774 = w1796 & w4866;
assign w1775 = (~w5007 & w1219) | (~w5007 & w6212) | (w1219 & w6212);
assign w1776 = (w4340 & w5196) | (w4340 & w5892) | (w5196 & w5892);
assign w1777 = (w544 & w1586) | (w544 & w1942) | (w1586 & w1942);
assign w1778 = (w6100 & w3347) | (w6100 & w2135) | (w3347 & w2135);
assign w1779 = (~w693 & w2110) | (~w693 & w329) | (w2110 & w329);
assign w1780 = (~w1878 & ~w7118) | (~w1878 & w5492) | (~w7118 & w5492);
assign w1781 = (w2399 & w6988) | (w2399 & w7193) | (w6988 & w7193);
assign w1782 = (~w1847 & w477) | (~w1847 & w4763) | (w477 & w4763);
assign w1783 = ~w656 & ~w593;
assign w1784 = (w900 & w7036) | (w900 & ~w6501) | (w7036 & ~w6501);
assign w1785 = w6979 & w2285;
assign w1786 = ~w1345 & ~w6138;
assign w1787 = (~w2081 & w3141) | (~w2081 & w6028) | (w3141 & w6028);
assign w1788 = w1718 & ~w2811;
assign w1789 = ~w6991 & w6386;
assign w1790 = (~w3892 & w7077) | (~w3892 & w4413) | (w7077 & w4413);
assign w1791 = ~w3682 & ~w7027;
assign w1792 = ~w7215 & w6513;
assign w1793 = (w4323 & w2950) | (w4323 & ~w2453) | (w2950 & ~w2453);
assign w1794 = (~w1796 & ~w502) | (~w1796 & w1869) | (~w502 & w1869);
assign w1795 = (w615 & w1157) | (w615 & w4382) | (w1157 & w4382);
assign w1796 = ~w1565 & ~w7381;
assign w1797 = (w6180 & ~w268) | (w6180 & ~w2627) | (~w268 & ~w2627);
assign w1798 = w6031 & w1321;
assign w1799 = a169 & b169;
assign w1800 = w2099 & w124;
assign w1801 = ~w4496 & ~w1544;
assign w1802 = (w6323 & w6429) | (w6323 & w1743) | (w6429 & w1743);
assign w1803 = ~w1877 & w1575;
assign w1804 = ~w505 & ~w1443;
assign w1805 = ~w5368 & ~w2346;
assign w1806 = (~w7268 & w2418) | (~w7268 & w269) | (w2418 & w269);
assign w1807 = (w500 & w7079) | (w500 & ~w6981) | (w7079 & ~w6981);
assign w1808 = (~w3137 & w6270) | (~w3137 & w5674) | (w6270 & w5674);
assign w1809 = (w7174 & w3828) | (w7174 & ~w1632) | (w3828 & ~w1632);
assign w1810 = w2513 & w856;
assign w1811 = (w6082 & w6741) | (w6082 & w7318) | (w6741 & w7318);
assign w1812 = (w3391 & ~w5259) | (w3391 & w7030) | (~w5259 & w7030);
assign w1813 = ~w3480 & ~w6104;
assign w1814 = (w2847 & w688) | (w2847 & w3812) | (w688 & w3812);
assign w1815 = w719 | w5595;
assign w1816 = (~w2876 & w3980) | (~w2876 & w3125) | (w3980 & w3125);
assign w1817 = ~w2644 & w3349;
assign w1818 = w6383 & w730;
assign w1819 = w396 & ~w5223;
assign w1820 = (w5178 & w2322) | (w5178 & w6236) | (w2322 & w6236);
assign w1821 = ~w3855 & w1288;
assign w1822 = ~w4337 & w6539;
assign w1823 = w1929 & ~w5560;
assign w1824 = (w3327 & w6565) | (w3327 & w7560) | (w6565 & w7560);
assign w1825 = (w3728 & w974) | (w3728 & ~w3953) | (w974 & ~w3953);
assign w1826 = (~w4768 & ~w759) | (~w4768 & w5442) | (~w759 & w5442);
assign w1827 = a249 & b249;
assign w1828 = (w1598 & w2915) | (w1598 & w4604) | (w2915 & w4604);
assign w1829 = w322 & w4768;
assign w1830 = w113 & w6100;
assign w1831 = ~a70 & ~b70;
assign w1832 = ~w6510 & ~w3450;
assign w1833 = ~w6252 & ~w3320;
assign w1834 = (~w2624 & w6307) | (~w2624 & w5352) | (w6307 & w5352);
assign w1835 = (w3491 & w1834) | (w3491 & w7225) | (w1834 & w7225);
assign w1836 = (w6082 & w492) | (w6082 & w5709) | (w492 & w5709);
assign w1837 = a94 & b94;
assign w1838 = (~w788 & w4567) | (~w788 & ~w4966) | (w4567 & ~w4966);
assign w1839 = ~a8 & ~b8;
assign w1840 = w5042 & w5752;
assign w1841 = (w2123 & w3049) | (w2123 & w1782) | (w3049 & w1782);
assign w1842 = (~w4089 & w2753) | (~w4089 & w1406) | (w2753 & w1406);
assign w1843 = ~w3997 & ~w6386;
assign w1844 = (w7294 & w850) | (w7294 & w5020) | (w850 & w5020);
assign w1845 = w5284 & ~w7043;
assign w1846 = w6209 & ~w6774;
assign w1847 = (w5257 & w428) | (w5257 & w1924) | (w428 & w1924);
assign w1848 = a193 & b193;
assign w1849 = ~a130 & ~b130;
assign w1850 = (w2721 & w6686) | (w2721 & ~w5430) | (w6686 & ~w5430);
assign w1851 = ~w2636 & ~w5193;
assign w1852 = (w1765 & w1490) | (w1765 & w1634) | (w1490 & w1634);
assign w1853 = (w7437 & w4873) | (w7437 & w5403) | (w4873 & w5403);
assign w1854 = (~w5178 & w1392) | (~w5178 & w4312) | (w1392 & w4312);
assign w1855 = w1758 & w7547;
assign w1856 = ~w1570 & ~w3728;
assign w1857 = ~w7332 & w1110;
assign w1858 = w1541 & w4045;
assign w1859 = w7553 & ~w1227;
assign w1860 = ~a66 & ~b66;
assign w1861 = ~w7634 & w1878;
assign w1862 = w287 & ~w4639;
assign w1863 = (w488 & w7029) | (w488 & w7046) | (w7029 & w7046);
assign w1864 = w910 & w4548;
assign w1865 = (~w777 & w966) | (~w777 & w490) | (w966 & w490);
assign w1866 = ~a164 & ~b164;
assign w1867 = (w2301 & w7006) | (w2301 & w3491) | (w7006 & w3491);
assign w1868 = ~w1002 & ~w7372;
assign w1869 = (~w502 & w1536) | (~w502 & ~w7378) | (w1536 & ~w7378);
assign w1870 = (w681 & w1100) | (w681 & ~w3515) | (w1100 & ~w3515);
assign w1871 = ~w1847 & w752;
assign w1872 = ~w2131 & w1097;
assign w1873 = ~w6046 & ~w4918;
assign w1874 = (~w5178 & w5682) | (~w5178 & w460) | (w5682 & w460);
assign w1875 = w2483 & w3916;
assign w1876 = (w3318 & w3419) | (w3318 & w1633) | (w3419 & w1633);
assign w1877 = ~w812 & ~w4148;
assign w1878 = ~w593 & ~w790;
assign w1879 = ~w5732 & w2884;
assign w1880 = (w5995 & w5234) | (w5995 & w1001) | (w5234 & w1001);
assign w1881 = (~w6439 & w472) | (~w6439 & w3914) | (w472 & w3914);
assign w1882 = ~w999 & w583;
assign w1883 = ~a77 & ~b77;
assign w1884 = w7364 & ~w664;
assign w1885 = (~w783 & w7594) | (~w783 & w4845) | (w7594 & w4845);
assign w1886 = ~w5901 & w2906;
assign w1887 = (w6254 & w647) | (w6254 & w6107) | (w647 & w6107);
assign w1888 = (~w4123 & ~w5629) | (~w4123 & w1590) | (~w5629 & w1590);
assign w1889 = (~w7302 & w4030) | (~w7302 & ~w7567) | (w4030 & ~w7567);
assign w1890 = w6325 & ~w5499;
assign w1891 = ~w2751 & ~w3817;
assign w1892 = ~w2456 & w5385;
assign w1893 = (w550 & w7423) | (w550 & w3198) | (w7423 & w3198);
assign w1894 = w5799 | w3609;
assign w1895 = (~w5178 & w469) | (~w5178 & w1996) | (w469 & w1996);
assign w1896 = (~w1611 & w5833) | (~w1611 & w3941) | (w5833 & w3941);
assign w1897 = w1195 & ~w1265;
assign w1898 = (w1723 & ~w5257) | (w1723 & w3280) | (~w5257 & w3280);
assign w1899 = (~w7592 & w3099) | (~w7592 & w1620) | (w3099 & w1620);
assign w1900 = ~w6697 & ~w5073;
assign w1901 = a104 & b104;
assign w1902 = (w1365 & w1301) | (w1365 & ~w5098) | (w1301 & ~w5098);
assign w1903 = ~w714 & w3888;
assign w1904 = (w5083 & ~w2152) | (w5083 & ~w7108) | (~w2152 & ~w7108);
assign w1905 = w220 & ~w5493;
assign w1906 = w144 & ~w7481;
assign w1907 = w1131 & ~w1977;
assign w1908 = w5723 & ~w3640;
assign w1909 = (w5511 & w2857) | (w5511 & w108) | (w2857 & w108);
assign w1910 = (~w4822 & w6839) | (~w4822 & w6544) | (w6839 & w6544);
assign w1911 = ~w1799 & ~w6094;
assign w1912 = ~w4993 & ~w378;
assign w1913 = w5399 & ~w608;
assign w1914 = w3467 & w3819;
assign w1915 = (~w3336 & w252) | (~w3336 & ~w4940) | (w252 & ~w4940);
assign w1916 = w6015 | w1355;
assign w1917 = (w2897 & w2549) | (w2897 & w5655) | (w2549 & w5655);
assign w1918 = ~w3947 & w239;
assign w1919 = (~w5344 & w6835) | (~w5344 & w1961) | (w6835 & w1961);
assign w1920 = (~w4833 & ~w4685) | (~w4833 & w5490) | (~w4685 & w5490);
assign w1921 = ~w2024 & w1797;
assign w1922 = (~w4648 & w3163) | (~w4648 & ~w6174) | (w3163 & ~w6174);
assign w1923 = ~a154 & ~b154;
assign w1924 = (w4161 & w705) | (w4161 & w2835) | (w705 & w2835);
assign w1925 = a198 & b198;
assign w1926 = w3238 & w7187;
assign w1927 = (~w6149 & w6082) | (~w6149 & w1233) | (w6082 & w1233);
assign w1928 = (w5069 & w5841) | (w5069 & w7312) | (w5841 & w7312);
assign w1929 = ~w471 & w6516;
assign w1930 = w991 & w2971;
assign w1931 = ~w7450 & w3238;
assign w1932 = (~w6100 & w6185) | (~w6100 & w4112) | (w6185 & w4112);
assign w1933 = (w6324 & w5920) | (w6324 & w6313) | (w5920 & w6313);
assign w1934 = (w2952 & w7263) | (w2952 & w3491) | (w7263 & w3491);
assign w1935 = (~w5178 & w3725) | (~w5178 & w5975) | (w3725 & w5975);
assign w1936 = w5058 & w3197;
assign w1937 = ~w6994 & w761;
assign w1938 = a161 & b161;
assign w1939 = (~w671 & w4256) | (~w671 & w4172) | (w4256 & w4172);
assign w1940 = (w2367 & w3276) | (w2367 & ~w4199) | (w3276 & ~w4199);
assign w1941 = (~w978 & w3542) | (~w978 & w7358) | (w3542 & w7358);
assign w1942 = ~w6082 & w2695;
assign w1943 = (w1847 & w2374) | (w1847 & w5701) | (w2374 & w5701);
assign w1944 = ~w1812 & w7118;
assign w1945 = w7138 & w906;
assign w1946 = ~w3014 & w4102;
assign w1947 = (w1048 & w5308) | (w1048 & w6501) | (w5308 & w6501);
assign w1948 = (w7448 & w5165) | (w7448 & ~w1730) | (w5165 & ~w1730);
assign w1949 = w4130 & w1295;
assign w1950 = w6162 & w433;
assign w1951 = ~w3679 & w222;
assign w1952 = ~w3813 & w4336;
assign w1953 = (~w4296 & w5481) | (~w4296 & w6371) | (w5481 & w6371);
assign w1954 = ~w832 & ~w6281;
assign w1955 = (w3062 & w3286) | (w3062 & w2903) | (w3286 & w2903);
assign w1956 = (~w723 & w4665) | (~w723 & w1458) | (w4665 & w1458);
assign w1957 = w3480 & ~w3618;
assign w1958 = w5230 & ~w7614;
assign w1959 = w5399 & w5071;
assign w1960 = w5251 & ~w3262;
assign w1961 = w4672 & ~w2315;
assign w1962 = (~w4287 & w4732) | (~w4287 & w6447) | (w4732 & w6447);
assign w1963 = w2203 & ~w1545;
assign w1964 = ~w995 & w5556;
assign w1965 = w547 & ~w6984;
assign w1966 = (w6053 & w1347) | (w6053 & ~w145) | (w1347 & ~w145);
assign w1967 = a218 & b218;
assign w1968 = (~w3108 & w2078) | (~w3108 & w3731) | (w2078 & w3731);
assign w1969 = (~w4875 & ~w2981) | (~w4875 & w5669) | (~w2981 & w5669);
assign w1970 = (~w5346 & ~w783) | (~w5346 & ~w813) | (~w783 & ~w813);
assign w1971 = (~w5961 & w6807) | (~w5961 & w594) | (w6807 & w594);
assign w1972 = ~w1831 & ~w1026;
assign w1973 = ~w163 & ~w2917;
assign w1974 = a10 & b10;
assign w1975 = w6924 & ~w721;
assign w1976 = (~w6524 & w663) | (~w6524 & ~w3989) | (w663 & ~w3989);
assign w1977 = w3911 & ~w4831;
assign w1978 = (w2969 & w296) | (w2969 & w2718) | (w296 & w2718);
assign w1979 = (w912 & w874) | (w912 & w2013) | (w874 & w2013);
assign w1980 = ~a218 & ~b218;
assign w1981 = ~w1754 & ~w5743;
assign w1982 = (~w13 & ~w5627) | (~w13 & w3593) | (~w5627 & w3593);
assign w1983 = ~w2037 & w3851;
assign w1984 = ~w4651 & ~w6141;
assign w1985 = (w5821 & w3484) | (w5821 & w5454) | (w3484 & w5454);
assign w1986 = w3965 & ~w4911;
assign w1987 = (w6122 & ~w3854) | (w6122 & w3666) | (~w3854 & w3666);
assign w1988 = (~w7108 & w5090) | (~w7108 & w1118) | (w5090 & w1118);
assign w1989 = (w2006 & w536) | (w2006 & w934) | (w536 & w934);
assign w1990 = ~w990 & w788;
assign w1991 = ~w3306 & ~w2836;
assign w1992 = (w3387 & ~w857) | (w3387 & w3810) | (~w857 & w3810);
assign w1993 = w125 & ~w5560;
assign w1994 = (~w2985 & w6768) | (~w2985 & w3649) | (w6768 & w3649);
assign w1995 = ~w4368 & w3169;
assign w1996 = (~w5027 & w603) | (~w5027 & w4799) | (w603 & w4799);
assign w1997 = ~w3040 & w4389;
assign w1998 = w3474 & ~w6239;
assign w1999 = ~a50 & ~b50;
assign w2000 = ~w7553 & w1227;
assign w2001 = ~w1241 & ~w454;
assign w2002 = (~w5325 & ~w6468) | (~w5325 & ~w6142) | (~w6468 & ~w6142);
assign w2003 = (w3774 & w2700) | (w3774 & w5812) | (w2700 & w5812);
assign w2004 = (w3045 & ~w6353) | (w3045 & w6389) | (~w6353 & w6389);
assign w2005 = a213 & b213;
assign w2006 = (w2021 & w6449) | (w2021 & ~w1693) | (w6449 & ~w1693);
assign w2007 = w5292 & ~w2744;
assign w2008 = w1785 & w2285;
assign w2009 = w3281 & w4924;
assign w2010 = w3106 & w2978;
assign w2011 = ~w301 & ~w5915;
assign w2012 = (~w6945 & w5218) | (~w6945 & w694) | (w5218 & w694);
assign w2013 = w4867 & ~w2453;
assign w2014 = (~w5106 & w4716) | (~w5106 & w5391) | (w4716 & w5391);
assign w2015 = (w5178 & w1746) | (w5178 & w6825) | (w1746 & w6825);
assign w2016 = (w961 & w3565) | (w961 & w5403) | (w3565 & w5403);
assign w2017 = ~w385 & w3087;
assign w2018 = w4990 & w1547;
assign w2019 = a9 & b9;
assign w2020 = ~w6037 & w379;
assign w2021 = (w6019 & w3078) | (w6019 & w4522) | (w3078 & w4522);
assign w2022 = (w6649 & w519) | (w6649 & w7624) | (w519 & w7624);
assign w2023 = (~w4329 & ~w6324) | (~w4329 & w4521) | (~w6324 & w4521);
assign w2024 = ~w2913 & ~w3616;
assign w2025 = ~w1132 & ~w1068;
assign w2026 = (w719 & ~w671) | (w719 & w2788) | (~w671 & w2788);
assign w2027 = a42 & b42;
assign w2028 = (w4011 & w2847) | (w4011 & w5941) | (w2847 & w5941);
assign w2029 = w2027 & ~w1053;
assign w2030 = (w887 & ~w6688) | (w887 & w7393) | (~w6688 & w7393);
assign w2031 = (w3942 & w5388) | (w3942 & w346) | (w5388 & w346);
assign w2032 = w3894 & w4069;
assign w2033 = (~w5178 & w6509) | (~w5178 & w1992) | (w6509 & w1992);
assign w2034 = ~w7023 & ~w7620;
assign w2035 = (~w5257 & w7376) | (~w5257 & w3586) | (w7376 & w3586);
assign w2036 = w5848 | ~w651;
assign w2037 = (w6100 & w6197) | (w6100 & w4240) | (w6197 & w4240);
assign w2038 = (w343 & w3915) | (w343 & w609) | (w3915 & w609);
assign w2039 = ~w4018 & ~w7033;
assign w2040 = w5980 & ~w6397;
assign w2041 = (~w7564 & w4970) | (~w7564 & w5543) | (w4970 & w5543);
assign w2042 = (~w5478 & w3957) | (~w5478 & w4216) | (w3957 & w4216);
assign w2043 = ~w3093 & w1959;
assign w2044 = (~w3057 & w4405) | (~w3057 & w4390) | (w4405 & w4390);
assign w2045 = ~w4180 & ~w4564;
assign w2046 = (w3407 & w5471) | (w3407 & w5007) | (w5471 & w5007);
assign w2047 = (~w3947 & w7465) | (~w3947 & w80) | (w7465 & w80);
assign w2048 = w5126 & w442;
assign w2049 = w5616 & ~w3269;
assign w2050 = w576 & ~w1420;
assign w2051 = (~w1193 & w537) | (~w1193 & w3777) | (w537 & w3777);
assign w2052 = (w868 & ~w488) | (w868 & w4188) | (~w488 & w4188);
assign w2053 = (w3318 & w4608) | (w3318 & w5378) | (w4608 & w5378);
assign w2054 = w2853 & ~w6571;
assign w2055 = w4833 & ~w6013;
assign w2056 = (w5178 & w3783) | (w5178 & w6521) | (w3783 & w6521);
assign w2057 = ~w230 & w3118;
assign w2058 = ~cin & w4606;
assign w2059 = w2644 & ~w6279;
assign w2060 = (w735 & w5750) | (w735 & ~w3330) | (w5750 & ~w3330);
assign w2061 = w7124 & ~w2548;
assign w2062 = (~w7035 & w7218) | (~w7035 & w7445) | (w7218 & w7445);
assign w2063 = ~w4527 & ~w5195;
assign w2064 = ~w1860 & w978;
assign w2065 = (w4187 & w5321) | (w4187 & w4302) | (w5321 & w4302);
assign w2066 = a214 & b214;
assign w2067 = ~w1002 & w860;
assign w2068 = ~w7493 & ~w1563;
assign w2069 = ~w1143 & ~w5848;
assign w2070 = (w6100 & w1337) | (w6100 & w5495) | (w1337 & w5495);
assign w2071 = w1395 & w6100;
assign w2072 = w960 & ~w7536;
assign w2073 = ~w103 & ~w2548;
assign w2074 = ~w651 & ~w1837;
assign w2075 = (~w5291 & w4244) | (~w5291 & w2149) | (w4244 & w2149);
assign w2076 = (~w2453 & ~w632) | (~w2453 & ~w6738) | (~w632 & ~w6738);
assign w2077 = ~w6426 & ~w6939;
assign w2078 = w4185 & ~w3108;
assign w2079 = (w7409 & w903) | (w7409 & w5076) | (w903 & w5076);
assign w2080 = w7345 & ~w5930;
assign w2081 = ~w4468 & ~w5425;
assign w2082 = ~w6054 & ~w3045;
assign w2083 = ~w3679 & w714;
assign w2084 = ~a114 & ~b114;
assign w2085 = ~w314 & w7290;
assign w2086 = ~w2582 & w1295;
assign w2087 = (~w3078 & w6350) | (~w3078 & w7347) | (w6350 & w7347);
assign w2088 = w2566 & w7530;
assign w2089 = ~w1288 & ~w646;
assign w2090 = ~w2603 & w1421;
assign w2091 = (w7118 & w4381) | (w7118 & w4359) | (w4381 & w4359);
assign w2092 = (w6534 & w4469) | (w6534 & w5417) | (w4469 & w5417);
assign w2093 = w7127 & ~w2084;
assign w2094 = ~w6854 & w6594;
assign w2095 = ~w4306 & w4499;
assign w2096 = w2671 & ~w60;
assign w2097 = ~w5871 & w7124;
assign w2098 = (w5178 & w2646) | (w5178 & w2893) | (w2646 & w2893);
assign w2099 = ~w4218 & w1432;
assign w2100 = (w2627 & w104) | (w2627 & w3026) | (w104 & w3026);
assign w2101 = ~w5871 & w6508;
assign w2102 = (w6190 & w4650) | (w6190 & ~w3852) | (w4650 & ~w3852);
assign w2103 = (w7 & w4106) | (w7 & w3332) | (w4106 & w3332);
assign w2104 = ~a220 & ~b220;
assign w2105 = ~w2131 & w527;
assign w2106 = (w5178 & w6131) | (w5178 & w5335) | (w6131 & w5335);
assign w2107 = ~w2605 & ~w2636;
assign w2108 = w3905 & ~w3135;
assign w2109 = w7405 & ~w1905;
assign w2110 = ~w693 & w6209;
assign w2111 = (w7418 & w2859) | (w7418 & ~w5098) | (w2859 & ~w5098);
assign w2112 = ~w6492 & ~w2210;
assign w2113 = (~w7626 & w288) | (~w7626 & w2183) | (w288 & w2183);
assign w2114 = (w1458 & w1956) | (w1458 & ~w2013) | (w1956 & ~w2013);
assign w2115 = w4990 & ~w6621;
assign w2116 = (w144 & w5905) | (w144 & w1114) | (w5905 & w1114);
assign w2117 = (~w978 & w6865) | (~w978 & w2228) | (w6865 & w2228);
assign w2118 = w6805 & w7570;
assign w2119 = w6791 & ~w6243;
assign w2120 = (~w1141 & w7067) | (~w1141 & w2781) | (w7067 & w2781);
assign w2121 = w2975 | ~w3840;
assign w2122 = ~w1753 & ~w51;
assign w2123 = w2903 & w5655;
assign w2124 = w6991 & ~w4000;
assign w2125 = (w1474 & w2847) | (w1474 & w1373) | (w2847 & w1373);
assign w2126 = w1765 & ~w5046;
assign w2127 = a190 & b190;
assign w2128 = (~w2847 & w1363) | (~w2847 & w1648) | (w1363 & w1648);
assign w2129 = ~w5230 & ~w6281;
assign w2130 = (w3311 & w4423) | (w3311 & w7454) | (w4423 & w7454);
assign w2131 = w5423 & w5136;
assign w2132 = (~w3471 & w1182) | (~w3471 & w7512) | (w1182 & w7512);
assign w2133 = (w1692 & w4167) | (w1692 & w58) | (w4167 & w58);
assign w2134 = w1453 & w6359;
assign w2135 = (w1755 & w5332) | (w1755 & w3034) | (w5332 & w3034);
assign w2136 = ~w4082 & ~w5803;
assign w2137 = (w5655 & w6921) | (w5655 & w1955) | (w6921 & w1955);
assign w2138 = (w4687 & w2268) | (w4687 & w5291) | (w2268 & w5291);
assign w2139 = (~w3847 & ~w2456) | (~w3847 & ~w4286) | (~w2456 & ~w4286);
assign w2140 = ~w145 & w3333;
assign w2141 = ~w2688 & w7026;
assign w2142 = ~w6342 & ~w7525;
assign w2143 = ~w2011 & w64;
assign w2144 = (~w732 & w1898) | (~w732 & w2772) | (w1898 & w2772);
assign w2145 = w1247 & w1945;
assign w2146 = ~w7291 & ~w2797;
assign w2147 = (w4537 & w5270) | (w4537 & ~w5098) | (w5270 & ~w5098);
assign w2148 = ~w6193 & ~w2895;
assign w2149 = (w3899 & w613) | (w3899 & ~w7238) | (w613 & ~w7238);
assign w2150 = (~w5834 & w6672) | (~w5834 & w6305) | (w6672 & w6305);
assign w2151 = ~w425 & w4646;
assign w2152 = ~w6022 & ~w3043;
assign w2153 = w3152 & w1272;
assign w2154 = (w6966 & w6059) | (w6966 & w5116) | (w6059 & w5116);
assign w2155 = (w3301 & w338) | (w3301 & ~w7187) | (w338 & ~w7187);
assign w2156 = ~w2257 & w1279;
assign w2157 = (~w4415 & w2745) | (~w4415 & ~w2097) | (w2745 & ~w2097);
assign w2158 = (w599 & w5468) | (w599 & w4528) | (w5468 & w4528);
assign w2159 = (~w7238 & w6730) | (~w7238 & w1795) | (w6730 & w1795);
assign w2160 = w1002 & ~w860;
assign w2161 = (w4187 & w1703) | (w4187 & w1217) | (w1703 & w1217);
assign w2162 = (w4609 & w2146) | (w4609 & w6254) | (w2146 & w6254);
assign w2163 = w4975 & ~w5782;
assign w2164 = (w176 & w271) | (w176 & ~w6100) | (w271 & ~w6100);
assign w2165 = (~w5325 & w6527) | (~w5325 & w6368) | (w6527 & w6368);
assign w2166 = (w3444 & w2226) | (w3444 & ~w5432) | (w2226 & ~w5432);
assign w2167 = w7307 & ~w1682;
assign w2168 = (w6600 & w1473) | (w6600 & ~w2097) | (w1473 & ~w2097);
assign w2169 = w6965 | ~w7097;
assign w2170 = (w2874 & w4226) | (w2874 & w7199) | (w4226 & w7199);
assign w2171 = w1754 & ~w3075;
assign w2172 = ~w3719 & w612;
assign w2173 = ~a206 & ~b206;
assign w2174 = ~w1854 & ~w5145;
assign w2175 = w3430 & ~w3058;
assign w2176 = ~w3693 & w4081;
assign w2177 = ~w2317 & w2018;
assign w2178 = (w2112 & w3557) | (w2112 & w2666) | (w3557 & w2666);
assign w2179 = ~w3052 & ~w3855;
assign w2180 = (w1324 & w1232) | (w1324 & w3892) | (w1232 & w3892);
assign w2181 = (w7409 & w903) | (w7409 & ~w3576) | (w903 & ~w3576);
assign w2182 = ~w1723 & w5948;
assign w2183 = (~w215 & w634) | (~w215 & w5240) | (w634 & w5240);
assign w2184 = (w7015 & w2848) | (w7015 & w4052) | (w2848 & w4052);
assign w2185 = (~w5834 & w3510) | (~w5834 & w3935) | (w3510 & w3935);
assign w2186 = (w5774 & w3916) | (w5774 & w3615) | (w3916 & w3615);
assign w2187 = w3132 & w690;
assign w2188 = ~w4185 & w3108;
assign w2189 = w2981 & w4749;
assign w2190 = w2600 & ~w4265;
assign w2191 = (~w3312 & w615) | (~w3312 & w1066) | (w615 & w1066);
assign w2192 = w3019 & ~w7183;
assign w2193 = w2829 & w2267;
assign w2194 = (~w3819 & w1857) | (~w3819 & w2442) | (w1857 & w2442);
assign w2195 = ~w3086 & ~w4436;
assign w2196 = (~w5178 & w1476) | (~w5178 & w4937) | (w1476 & w4937);
assign w2197 = ~w1753 & ~w278;
assign w2198 = (w3242 & w6523) | (w3242 & w5291) | (w6523 & w5291);
assign w2199 = (w2456 & w3953) | (w2456 & w7091) | (w3953 & w7091);
assign w2200 = (~w1143 & w2069) | (~w1143 & ~w6633) | (w2069 & ~w6633);
assign w2201 = (~w5202 & w2827) | (~w5202 & w1181) | (w2827 & w1181);
assign w2202 = ~w6444 & ~w1588;
assign w2203 = ~w7641 & ~w3799;
assign w2204 = ~w7523 & ~w4957;
assign w2205 = w394 & ~w5424;
assign w2206 = ~w583 & ~w6147;
assign w2207 = (w3354 & w1644) | (w3354 & w592) | (w1644 & w592);
assign w2208 = (~w6353 & w3605) | (~w6353 & w1537) | (w3605 & w1537);
assign w2209 = (w4187 & w4065) | (w4187 & w2764) | (w4065 & w2764);
assign w2210 = ~w2519 & ~w6484;
assign w2211 = w3690 & ~w6099;
assign w2212 = (~w5178 & w562) | (~w5178 & w6441) | (w562 & w6441);
assign w2213 = ~w2098 & ~w6083;
assign w2214 = (~w3264 & ~w2382) | (~w3264 & w990) | (~w2382 & w990);
assign w2215 = (w4995 & w1603) | (w4995 & w1495) | (w1603 & w1495);
assign w2216 = a141 & b141;
assign w2217 = (w7625 & w438) | (w7625 & w3765) | (w438 & w3765);
assign w2218 = ~w6335 & ~w2084;
assign w2219 = (w6460 & w4738) | (w6460 & w4199) | (w4738 & w4199);
assign w2220 = (w3490 & w7032) | (w3490 & w4105) | (w7032 & w4105);
assign w2221 = ~w3382 & w7396;
assign w2222 = ~w1431 & ~w1352;
assign w2223 = (w2332 & w1043) | (w2332 & ~w7238) | (w1043 & ~w7238);
assign w2224 = (w1868 & w126) | (w1868 & w959) | (w126 & w959);
assign w2225 = (~w7106 & w578) | (~w7106 & w3847) | (w578 & w3847);
assign w2226 = w6375 & w3444;
assign w2227 = (~w4651 & w5553) | (~w4651 & w5836) | (w5553 & w5836);
assign w2228 = (w493 & w6542) | (w493 & w738) | (w6542 & w738);
assign w2229 = w2945 & ~w5676;
assign w2230 = ~w5999 & ~w5598;
assign w2231 = (w3496 & w2389) | (w3496 & ~w3119) | (w2389 & ~w3119);
assign w2232 = ~w7546 & ~w850;
assign w2233 = (w2627 & w280) | (w2627 & w6925) | (w280 & w6925);
assign w2234 = (~w1367 & w6145) | (~w1367 & w2552) | (w6145 & w2552);
assign w2235 = (~w761 & w1306) | (~w761 & w7512) | (w1306 & w7512);
assign w2236 = ~w4976 & w1529;
assign w2237 = w5330 & ~w968;
assign w2238 = ~w1441 & w6122;
assign w2239 = (w1609 & w2778) | (w1609 & ~w3679) | (w2778 & ~w3679);
assign w2240 = (w6738 & w4020) | (w6738 & w446) | (w4020 & w446);
assign w2241 = (w5648 & w858) | (w5648 & w1732) | (w858 & w1732);
assign w2242 = ~w7397 & w2440;
assign w2243 = ~a82 & ~b82;
assign w2244 = ~w7572 & ~w2591;
assign w2245 = w5762 & ~w9;
assign w2246 = ~w5510 & w6656;
assign w2247 = w4867 & ~w2097;
assign w2248 = ~w4503 & w4457;
assign w2249 = ~w3294 & ~w234;
assign w2250 = (~w2740 & ~w1888) | (~w2740 & w7062) | (~w1888 & w7062);
assign w2251 = (w1150 & w6646) | (w1150 & ~w1892) | (w6646 & ~w1892);
assign w2252 = (w5921 & w5290) | (w5921 & ~w2013) | (w5290 & ~w2013);
assign w2253 = ~a165 & ~b165;
assign w2254 = (~w5788 & w2452) | (~w5788 & w2258) | (w2452 & w2258);
assign w2255 = a105 & b105;
assign w2256 = (~w6746 & w1065) | (~w6746 & w2614) | (w1065 & w2614);
assign w2257 = ~w7350 & ~w2279;
assign w2258 = ~w4488 & ~w5788;
assign w2259 = ~w5464 & ~w5570;
assign w2260 = ~a104 & ~b104;
assign w2261 = a111 & b111;
assign w2262 = (w7018 & w5001) | (w7018 & w277) | (w5001 & w277);
assign w2263 = w577 & ~w4089;
assign w2264 = (~w3888 & w4777) | (~w3888 & w949) | (w4777 & w949);
assign w2265 = w6257 & ~w4296;
assign w2266 = (w412 & w1294) | (w412 & w357) | (w1294 & w357);
assign w2267 = (~w226 & ~w5257) | (~w226 & w5694) | (~w5257 & w5694);
assign w2268 = ~w3451 & w4687;
assign w2269 = (w5961 & w2581) | (w5961 & w3998) | (w2581 & w3998);
assign w2270 = ~w1371 & ~w6729;
assign w2271 = ~w161 & w468;
assign w2272 = (~w1936 & w6270) | (~w1936 & w1808) | (w6270 & w1808);
assign w2273 = ~w6181 & ~w2849;
assign w2274 = w5241 & ~w3122;
assign w2275 = (w2766 & w5297) | (w2766 & w5695) | (w5297 & w5695);
assign w2276 = ~w7363 & ~w2315;
assign w2277 = (~w3019 & w1023) | (~w3019 & ~w7187) | (w1023 & ~w7187);
assign w2278 = a182 & b182;
assign w2279 = a85 & b85;
assign w2280 = (w5257 & w5586) | (w5257 & w5918) | (w5586 & w5918);
assign w2281 = w7622 & ~w4765;
assign w2282 = (w5257 & w7459) | (w5257 & w3844) | (w7459 & w3844);
assign w2283 = a100 & b100;
assign w2284 = ~w1991 & w7216;
assign w2285 = ~w2658 & ~w216;
assign w2286 = w7614 & ~w3669;
assign w2287 = w1373 & ~w5296;
assign w2288 = ~w1563 & ~w2648;
assign w2289 = ~w4843 & ~w226;
assign w2290 = (~w1467 & w2359) | (~w1467 & w6584) | (w2359 & w6584);
assign w2291 = w4271 & w6682;
assign w2292 = (w837 & w94) | (w837 & w745) | (w94 & w745);
assign w2293 = w3911 & w758;
assign w2294 = ~w1137 & ~w5442;
assign w2295 = a252 & b252;
assign w2296 = ~w2066 & ~w664;
assign w2297 = (~w3932 & ~w4995) | (~w3932 & w2884) | (~w4995 & w2884);
assign w2298 = (w777 & w6578) | (w777 & w309) | (w6578 & w309);
assign w2299 = ~w3262 & ~w7493;
assign w2300 = w995 & ~w5556;
assign w2301 = ~w3643 & ~w7227;
assign w2302 = (~w5277 & ~w2588) | (~w5277 & w954) | (~w2588 & w954);
assign w2303 = (w2393 & w1147) | (w2393 & w1936) | (w1147 & w1936);
assign w2304 = ~w331 & w6439;
assign w2305 = w2197 & w2286;
assign w2306 = ~w5178 & w3645;
assign w2307 = w6063 & ~w664;
assign w2308 = (~w6718 & w6023) | (~w6718 & w3971) | (w6023 & w3971);
assign w2309 = w1606 & ~w5627;
assign w2310 = (~w4759 & w4458) | (~w4759 & w2405) | (w4458 & w2405);
assign w2311 = (~w7091 & w6182) | (~w7091 & w3531) | (w6182 & w3531);
assign w2312 = w1617 & w6863;
assign w2313 = ~w7566 | w5537;
assign w2314 = w3587 & ~w3331;
assign w2315 = (~w4457 & w145) | (~w4457 & w2720) | (w145 & w2720);
assign w2316 = (~w6016 & w6698) | (~w6016 & w7458) | (w6698 & w7458);
assign w2317 = w3028 & ~w917;
assign w2318 = (~w736 & ~w1384) | (~w736 & w3459) | (~w1384 & w3459);
assign w2319 = (w3066 & w676) | (w3066 & w5589) | (w676 & w5589);
assign w2320 = ~w2849 & w6486;
assign w2321 = (w2847 & w5878) | (w2847 & w5413) | (w5878 & w5413);
assign w2322 = (w834 & ~w3491) | (w834 & w1458) | (~w3491 & w1458);
assign w2323 = (~w1698 & w2805) | (~w1698 & w4441) | (w2805 & w4441);
assign w2324 = (~w1607 & w2030) | (~w1607 & w7645) | (w2030 & w7645);
assign w2325 = w3823 & ~w6744;
assign w2326 = ~w182 & ~w2521;
assign w2327 = ~w6147 & ~w6342;
assign w2328 = (w2985 & w3552) | (w2985 & w2009) | (w3552 & w2009);
assign w2329 = ~w7215 & ~w1980;
assign w2330 = (w1227 & w3408) | (w1227 & w1315) | (w3408 & w1315);
assign w2331 = (w6894 & w5249) | (w6894 & w2113) | (w5249 & w2113);
assign w2332 = w1751 & w2681;
assign w2333 = ~w5616 & w4084;
assign w2334 = (~w4505 & w488) | (~w4505 & w7638) | (w488 & w7638);
assign w2335 = (w3078 & w411) | (w3078 & w6788) | (w411 & w6788);
assign w2336 = ~w5665 & ~w1098;
assign w2337 = w5498 | w2334;
assign w2338 = w960 & w4638;
assign w2339 = (~w7626 & w6409) | (~w7626 & w4951) | (w6409 & w4951);
assign w2340 = ~w1304 & w4468;
assign w2341 = w188 & ~w4216;
assign w2342 = w229 & w5136;
assign w2343 = ~w651 & w5176;
assign w2344 = (~w2123 & w4255) | (~w2123 & w2532) | (w4255 & w2532);
assign w2345 = ~w6039 & ~w4494;
assign w2346 = w7137 & ~w3092;
assign w2347 = ~w5066 | w3557;
assign w2348 = (w4296 & w5890) | (w4296 & w3625) | (w5890 & w3625);
assign w2349 = (~w6467 & w4582) | (~w6467 & w7128) | (w4582 & w7128);
assign w2350 = (w6106 & w6585) | (w6106 & w5313) | (w6585 & w5313);
assign w2351 = (w5708 & w4030) | (w5708 & w3148) | (w4030 & w3148);
assign w2352 = ~w5863 & ~w2945;
assign w2353 = ~a169 & ~b169;
assign w2354 = ~w1216 & w3210;
assign w2355 = (w5834 & w3506) | (w5834 & w4809) | (w3506 & w4809);
assign w2356 = w7141 | w6071;
assign w2357 = ~w3353 & w7506;
assign w2358 = w222 & ~w3936;
assign w2359 = (~w5526 & w5460) | (~w5526 & w3434) | (w5460 & w3434);
assign w2360 = ~w4415 & ~w7486;
assign w2361 = w931 & w4078;
assign w2362 = (w1369 & w3989) | (w1369 & w1230) | (w3989 & w1230);
assign w2363 = ~w596 & ~w1820;
assign w2364 = (~w7317 & w7198) | (~w7317 & w1394) | (w7198 & w1394);
assign w2365 = ~w7399 & ~w6335;
assign w2366 = (w6100 & w802) | (w6100 & w7301) | (w802 & w7301);
assign w2367 = (~w7490 & w5275) | (~w7490 & w4566) | (w5275 & w4566);
assign w2368 = ~w7596 & w5360;
assign w2369 = w6969 & w7413;
assign w2370 = w5655 & w397;
assign w2371 = ~w3654 & ~w6981;
assign w2372 = ~w3737 & w2421;
assign w2373 = (w4251 & w846) | (w4251 & w6633) | (w846 & w6633);
assign w2374 = ~w5361 & w4833;
assign w2375 = w4890 & w3886;
assign w2376 = (w5385 & w3383) | (w5385 & w1825) | (w3383 & w1825);
assign w2377 = (~w5998 & w5806) | (~w5998 & w4560) | (w5806 & w4560);
assign w2378 = w1140 & w4570;
assign w2379 = ~w7633 & w4387;
assign w2380 = (~w4060 & w884) | (~w4060 & w892) | (w884 & w892);
assign w2381 = ~w602 & ~w7274;
assign w2382 = (w7629 & w924) | (w7629 & ~w5464) | (w924 & ~w5464);
assign w2383 = (w5556 & w6814) | (w5556 & ~w3886) | (w6814 & ~w3886);
assign w2384 = ~w4987 & ~w804;
assign w2385 = ~w3634 & w2953;
assign w2386 = w1125 & ~w4247;
assign w2387 = (w1123 & w6764) | (w1123 & ~w1730) | (w6764 & ~w1730);
assign w2388 = w6553 & w5888;
assign w2389 = (~w2806 & w7064) | (~w2806 & w6556) | (w7064 & w6556);
assign w2390 = (~w5257 & w1894) | (~w5257 & w5758) | (w1894 & w5758);
assign w2391 = ~w3631 | w5596;
assign w2392 = (w445 & w4871) | (w445 & w3119) | (w4871 & w3119);
assign w2393 = ~w2597 & ~w2914;
assign w2394 = ~w6791 & ~w5466;
assign w2395 = w3408 & w1227;
assign w2396 = ~w991 & w7158;
assign w2397 = (w3952 & w7144) | (w3952 & w2826) | (w7144 & w2826);
assign w2398 = (w4357 & w1240) | (w4357 & ~w5417) | (w1240 & ~w5417);
assign w2399 = (~w5522 & w6860) | (~w5522 & w7567) | (w6860 & w7567);
assign w2400 = ~w6254 & w5435;
assign w2401 = ~w4967 & w4791;
assign w2402 = (w728 & ~w5830) | (w728 & w4019) | (~w5830 & w4019);
assign w2403 = (w1658 & w4640) | (w1658 & w4700) | (w4640 & w4700);
assign w2404 = w2011 & ~w3128;
assign w2405 = w4392 & ~w759;
assign w2406 = ~w2997 & ~w4940;
assign w2407 = ~w5279 & w2612;
assign w2408 = (w2343 & w5901) | (w2343 & w1701) | (w5901 & w1701);
assign w2409 = (~w698 & w1725) | (~w698 & w3771) | (w1725 & w3771);
assign w2410 = ~w1883 & ~w4060;
assign w2411 = (~w4825 & w1624) | (~w4825 & w4645) | (w1624 & w4645);
assign w2412 = (w5513 & w4272) | (w5513 & ~w4143) | (w4272 & ~w4143);
assign w2413 = w6935 & w913;
assign w2414 = (~w3491 & w4732) | (~w3491 & w1962) | (w4732 & w1962);
assign w2415 = w5297 & ~w3819;
assign w2416 = (w472 & w3056) | (w472 & w648) | (w3056 & w648);
assign w2417 = ~w3580 & ~w5944;
assign w2418 = w6087 & ~w7268;
assign w2419 = ~w478 & w7246;
assign w2420 = ~w5883 & ~w478;
assign w2421 = (w2188 & w2847) | (w2188 & w2866) | (w2847 & w2866);
assign w2422 = (w5007 & w371) | (w5007 & w3839) | (w371 & w3839);
assign w2423 = (w5325 & w6089) | (w5325 & w4008) | (w6089 & w4008);
assign w2424 = (w3986 & w760) | (w3986 & w3954) | (w760 & w3954);
assign w2425 = w649 & w1886;
assign w2426 = ~w6713 & w3528;
assign w2427 = w3152 & w406;
assign w2428 = (~w2627 & w6432) | (~w2627 & w610) | (w6432 & w610);
assign w2429 = (w4901 & ~w47) | (w4901 & w6123) | (~w47 & w6123);
assign w2430 = (~w6100 & w2325) | (~w6100 & w5552) | (w2325 & w5552);
assign w2431 = (~w478 & w2008) | (~w478 & w1422) | (w2008 & w1422);
assign w2432 = ~w6630 & ~w4247;
assign w2433 = ~w6222 & ~w2441;
assign w2434 = ~w6162 & ~w1738;
assign w2435 = a136 & b136;
assign w2436 = w4151 & w6512;
assign w2437 = w7362 & ~w5600;
assign w2438 = (w6031 & w5799) | (w6031 & w1408) | (w5799 & w1408);
assign w2439 = (w6100 & w7374) | (w6100 & w1790) | (w7374 & w1790);
assign w2440 = w7078 & w1554;
assign w2441 = a59 & b59;
assign w2442 = (~w7332 & w1110) | (~w7332 & w4239) | (w1110 & w4239);
assign w2443 = (~w3774 & w617) | (~w3774 & w4439) | (w617 & w4439);
assign w2444 = (~w632 & w1332) | (~w632 & w5814) | (w1332 & w5814);
assign w2445 = ~w3106 & ~w3304;
assign w2446 = (w3063 & w214) | (w3063 & w982) | (w214 & w982);
assign w2447 = w5042 & w6685;
assign w2448 = (~w5178 & w6110) | (~w5178 & w1112) | (w6110 & w1112);
assign w2449 = w2368 & ~w5755;
assign w2450 = a61 & b61;
assign w2451 = ~w6195 & w6754;
assign w2452 = ~w4348 & w2981;
assign w2453 = (~w3490 & w1949) | (~w3490 & w5534) | (w1949 & w5534);
assign w2454 = (w6353 & w4124) | (w6353 & w3006) | (w4124 & w3006);
assign w2455 = (w931 & w5140) | (w931 & ~w6206) | (w5140 & ~w6206);
assign w2456 = w4102 & ~w3894;
assign w2457 = ~w2568 & ~w3452;
assign w2458 = ~w4759 & w2326;
assign w2459 = (w3808 & ~w3986) | (w3808 & w585) | (~w3986 & w585);
assign w2460 = ~w3909 & ~w3782;
assign w2461 = (w4687 & w2268) | (w4687 & w563) | (w2268 & w563);
assign w2462 = ~w6397 & w6415;
assign w2463 = ~w6854 & w1594;
assign w2464 = w7279 & w344;
assign w2465 = ~a4 & ~b4;
assign w2466 = (w5648 & w858) | (w5648 & w1072) | (w858 & w1072);
assign w2467 = (~w837 & w5041) | (~w837 & w4724) | (w5041 & w4724);
assign w2468 = w3117 | w5921;
assign w2469 = ~w4520 & ~w6050;
assign w2470 = ~w5361 & w2055;
assign w2471 = ~w2173 & ~w698;
assign w2472 = (~w2353 & w5806) | (~w2353 & w5567) | (w5806 & w5567);
assign w2473 = w1315 & w3534;
assign w2474 = ~w1452 & ~w7626;
assign w2475 = (w4392 & w1021) | (w4392 & w2121) | (w1021 & w2121);
assign w2476 = ~w6640 & w5172;
assign w2477 = ~w4638 & w1440;
assign w2478 = (~w7283 & ~w4061) | (~w7283 & w6887) | (~w4061 & w6887);
assign w2479 = w7213 & ~w5442;
assign w2480 = (~w7510 & w4923) | (~w7510 & w3936) | (w4923 & w3936);
assign w2481 = (w7081 & w3708) | (w7081 & w5317) | (w3708 & w5317);
assign w2482 = w4003 & w6414;
assign w2483 = ~w5368 & ~w1575;
assign w2484 = (~w4647 & w5746) | (~w4647 & w1953) | (w5746 & w1953);
assign w2485 = ~w7279 & w5554;
assign w2486 = ~w4123 & w34;
assign w2487 = ~w941 & ~w1694;
assign w2488 = w194 & ~w144;
assign w2489 = (w4440 & w5593) | (w4440 & w5526) | (w5593 & w5526);
assign w2490 = w1326 & ~w3014;
assign w2491 = (w5725 & w5320) | (w5725 & w1730) | (w5320 & w1730);
assign w2492 = (~w6387 & w4771) | (~w6387 & w5403) | (w4771 & w5403);
assign w2493 = w2978 & w3140;
assign w2494 = ~w48 & w4538;
assign w2495 = w2971 & w440;
assign w2496 = ~w391 & ~w1661;
assign w2497 = w1321 & w7327;
assign w2498 = (~w3602 & w7048) | (~w3602 & w3754) | (w7048 & w3754);
assign w2499 = (w1598 & w2862) | (w1598 & w4932) | (w2862 & w4932);
assign w2500 = ~w6558 & ~w1265;
assign w2501 = ~w1032 & ~w1865;
assign w2502 = (w4966 & w3796) | (w4966 & w5984) | (w3796 & w5984);
assign w2503 = (~w6844 & w7629) | (~w6844 & w5959) | (w7629 & w5959);
assign w2504 = (~w5178 & w958) | (~w5178 & w6559) | (w958 & w6559);
assign w2505 = (w1516 & w3401) | (w1516 & w6801) | (w3401 & w6801);
assign w2506 = ~w3382 & ~w3207;
assign w2507 = (~w6526 & ~w4084) | (~w6526 & w1013) | (~w4084 & w1013);
assign w2508 = ~w196 & ~w3021;
assign w2509 = (w7041 & ~w837) | (w7041 & w4041) | (~w837 & w4041);
assign w2510 = w3040 & ~w7323;
assign w2511 = ~w531 & ~w3176;
assign w2512 = ~w6047 & ~w6611;
assign w2513 = ~w5930 & ~w6450;
assign w2514 = ~w101 & w3426;
assign w2515 = ~a76 & ~b76;
assign w2516 = w2329 & w6387;
assign w2517 = (w236 & w1530) | (w236 & w4659) | (w1530 & w4659);
assign w2518 = (w4182 & w1719) | (w4182 & w1348) | (w1719 & w1348);
assign w2519 = a233 & b233;
assign w2520 = (w4250 & w5196) | (w4250 & w88) | (w5196 & w88);
assign w2521 = ~a36 & ~b36;
assign w2522 = ~w1550 & ~w319;
assign w2523 = ~w1288 & ~w7051;
assign w2524 = (~w5007 & w2076) | (~w5007 & w5873) | (w2076 & w5873);
assign w2525 = (~w1499 & w2867) | (~w1499 & w2234) | (w2867 & w2234);
assign w2526 = ~w2557 & ~w6776;
assign w2527 = (~w7172 & w6285) | (~w7172 & ~w3114) | (w6285 & ~w3114);
assign w2528 = (w5422 & w3617) | (w5422 & ~w6174) | (w3617 & ~w6174);
assign w2529 = (w3116 & w1450) | (w3116 & ~w5611) | (w1450 & ~w5611);
assign w2530 = ~w936 & ~w1243;
assign w2531 = w7177 & ~w2393;
assign w2532 = w6517 & w6636;
assign w2533 = ~w7350 & w2279;
assign w2534 = ~w4168 & ~w5147;
assign w2535 = (~w6394 & w1160) | (~w6394 & w2821) | (w1160 & w2821);
assign w2536 = (w2603 & w1740) | (w2603 & w905) | (w1740 & w905);
assign w2537 = (w7414 & w2741) | (w7414 & w4835) | (w2741 & w4835);
assign w2538 = w238 & ~w1804;
assign w2539 = (~w5178 & w510) | (~w5178 & w4853) | (w510 & w4853);
assign w2540 = ~w5759 & ~w143;
assign w2541 = (~w1133 & w2287) | (~w1133 & w5618) | (w2287 & w5618);
assign w2542 = ~w6054 & ~w7525;
assign w2543 = (w2952 & w7263) | (w2952 & w2013) | (w7263 & w2013);
assign w2544 = ~w4503 & ~w2315;
assign w2545 = (~w7626 & w3051) | (~w7626 & w5240) | (w3051 & w5240);
assign w2546 = ~w2976 & ~w6824;
assign w2547 = (w6334 & w1885) | (w6334 & ~w484) | (w1885 & ~w484);
assign w2548 = ~w5732 & ~w7345;
assign w2549 = ~w7205 & w1405;
assign w2550 = w2522 & ~w1435;
assign w2551 = (~w3078 & w328) | (~w3078 & w1312) | (w328 & w1312);
assign w2552 = (~w322 & w3878) | (~w322 & w1089) | (w3878 & w1089);
assign w2553 = (w4045 & w1858) | (w4045 & w6025) | (w1858 & w6025);
assign w2554 = (~w6100 & w5232) | (~w6100 & w1504) | (w5232 & w1504);
assign w2555 = (~w3986 & w7099) | (~w3986 & w3956) | (w7099 & w3956);
assign w2556 = ~w5382 & ~w6247;
assign w2557 = ~w7513 & w3181;
assign w2558 = ~w6964 & w5792;
assign w2559 = ~w3953 & w7157;
assign w2560 = ~w812 & w2352;
assign w2561 = (~w3669 & w2286) | (~w3669 & w471) | (w2286 & w471);
assign w2562 = (w6501 & w33) | (w6501 & w4723) | (w33 & w4723);
assign w2563 = ~w6455 & ~w6981;
assign w2564 = ~w7372 & w7296;
assign w2565 = (~w3224 & w4328) | (~w3224 & w6141) | (w4328 & w6141);
assign w2566 = ~w1431 & ~w2596;
assign w2567 = a236 & b236;
assign w2568 = (~w5178 & w6157) | (~w5178 & w373) | (w6157 & w373);
assign w2569 = w1221 & w3466;
assign w2570 = ~w1515 & w5104;
assign w2571 = ~w6632 & ~w1108;
assign w2572 = ~w2749 & w245;
assign w2573 = (w7450 & w683) | (w7450 & w1035) | (w683 & w1035);
assign w2574 = (w3843 & w1598) | (w3843 & w3059) | (w1598 & w3059);
assign w2575 = (w728 & ~w4142) | (w728 & ~w5830) | (~w4142 & ~w5830);
assign w2576 = w72 & ~w6675;
assign w2577 = (w1847 & w7623) | (w1847 & w5907) | (w7623 & w5907);
assign w2578 = w7032 & ~w7056;
assign w2579 = w3158 & w129;
assign w2580 = (~w4066 & w5068) | (~w4066 & w7279) | (w5068 & w7279);
assign w2581 = (~w1004 & w2335) | (~w1004 & w3998) | (w2335 & w3998);
assign w2582 = (~w7486 & w6729) | (~w7486 & w7349) | (w6729 & w7349);
assign w2583 = (w3335 & w4450) | (w3335 & ~w7238) | (w4450 & ~w7238);
assign w2584 = ~w5792 & w1281;
assign w2585 = (~w6046 & w249) | (~w6046 & w1618) | (w249 & w1618);
assign w2586 = ~a119 & ~b119;
assign w2587 = ~w2012 & ~w678;
assign w2588 = (~w6766 & ~w4692) | (~w6766 & w3756) | (~w4692 & w3756);
assign w2589 = (w4187 & w1457) | (w4187 & w2069) | (w1457 & w2069);
assign w2590 = ~w6811 & ~w4970;
assign w2591 = a185 & b185;
assign w2592 = (w6770 & w3053) | (w6770 & w2475) | (w3053 & w2475);
assign w2593 = (w5834 & w3300) | (w5834 & w2689) | (w3300 & w2689);
assign w2594 = w5284 & ~w4803;
assign w2595 = w57 & ~w385;
assign w2596 = a17 & b17;
assign w2597 = ~a102 & ~b102;
assign w2598 = ~w790 & w5424;
assign w2599 = (~w1608 & w5272) | (~w1608 & w2972) | (w5272 & w2972);
assign w2600 = a69 & b69;
assign w2601 = ~w5250 & w6748;
assign w2602 = (~w5424 & w394) | (~w5424 & w3058) | (w394 & w3058);
assign w2603 = ~w4511 & w6113;
assign w2604 = (w7028 & w5011) | (w7028 & w1892) | (w5011 & w1892);
assign w2605 = w2749 & ~w5193;
assign w2606 = (w6885 & w7058) | (w6885 & w5250) | (w7058 & w5250);
assign w2607 = ~w1611 & w279;
assign w2608 = (w6664 & w1646) | (w6664 & w5291) | (w1646 & w5291);
assign w2609 = ~w4169 & ~w508;
assign w2610 = (~w777 & w1578) | (~w777 & w7573) | (w1578 & w7573);
assign w2611 = a200 & b200;
assign w2612 = ~w2658 & ~w5687;
assign w2613 = ~w3618 & ~w4847;
assign w2614 = (w7409 & w903) | (w7409 & ~w3953) | (w903 & ~w3953);
assign w2615 = (w5178 & w6711) | (w5178 & w2290) | (w6711 & w2290);
assign w2616 = ~w2829 & ~w2289;
assign w2617 = w2011 & ~w5937;
assign w2618 = (~w3364 & w2902) | (~w3364 & w3815) | (w2902 & w3815);
assign w2619 = ~w6985 & w3156;
assign w2620 = w7006 & w2301;
assign w2621 = ~w3887 & ~w4830;
assign w2622 = w4806 & w502;
assign w2623 = ~w5170 & w4940;
assign w2624 = ~w4830 & ~w3235;
assign w2625 = (w3011 & w4682) | (w3011 & w82) | (w4682 & w82);
assign w2626 = (w2083 & w6569) | (w2083 & w2762) | (w6569 & w2762);
assign w2627 = (w777 & w5810) | (w777 & w7508) | (w5810 & w7508);
assign w2628 = ~w516 & ~w5581;
assign w2629 = w1901 & ~w335;
assign w2630 = ~w182 & ~w4885;
assign w2631 = ~a83 & ~b83;
assign w2632 = a179 & b179;
assign w2633 = w6390 & w6792;
assign w2634 = w1864 & ~w818;
assign w2635 = w2863 & w6860;
assign w2636 = ~a65 & ~b65;
assign w2637 = ~w7010 & w2453;
assign w2638 = ~w6481 & ~w1647;
assign w2639 = (w2871 & w5282) | (w2871 & w4007) | (w5282 & w4007);
assign w2640 = (~w550 & w78) | (~w550 & w3964) | (w78 & w3964);
assign w2641 = (w6685 & w1660) | (w6685 & w4470) | (w1660 & w4470);
assign w2642 = ~w3789 & ~w4625;
assign w2643 = w1923 & ~w5287;
assign w2644 = ~a73 & ~b73;
assign w2645 = w4849 & ~w590;
assign w2646 = (w3640 & w4093) | (w3640 & w2492) | (w4093 & w2492);
assign w2647 = ~w3524 & ~w2707;
assign w2648 = a134 & b134;
assign w2649 = ~w4275 & ~w3965;
assign w2650 = ~w569 & ~w869;
assign w2651 = (w2969 & w2003) | (w2969 & w7571) | (w2003 & w7571);
assign w2652 = ~w7089 & ~w7125;
assign w2653 = (w632 & w482) | (w632 & w6431) | (w482 & w6431);
assign w2654 = ~w5760 & ~w1712;
assign w2655 = ~w4094 & ~w3739;
assign w2656 = (w401 & w5761) | (w401 & w4130) | (w5761 & w4130);
assign w2657 = ~w4430 & w334;
assign w2658 = ~a89 & ~b89;
assign w2659 = ~w4496 & ~w2966;
assign w2660 = w2049 | ~w3269;
assign w2661 = w4906 & w3070;
assign w2662 = (~w1063 & w1927) | (~w1063 & w3530) | (w1927 & w3530);
assign w2663 = ~w3312 & ~w471;
assign w2664 = ~w336 & w1851;
assign w2665 = (w5735 & w2489) | (w5735 & w5386) | (w2489 & w5386);
assign w2666 = ~w5066 & w2274;
assign w2667 = ~w2343 & ~w3469;
assign w2668 = (w7383 & w7323) | (w7383 & w4689) | (w7323 & w4689);
assign w2669 = w4688 & ~w6100;
assign w2670 = (w6501 & w224) | (w6501 & w1017) | (w224 & w1017);
assign w2671 = ~a14 & ~b14;
assign w2672 = ~w3782 & w3909;
assign w2673 = w4393 | w2792;
assign w2674 = (w7506 & w4177) | (w7506 & ~w3847) | (w4177 & ~w3847);
assign w2675 = (w6106 & w3859) | (w6106 & w3317) | (w3859 & w3317);
assign w2676 = (~w2806 & w3236) | (~w2806 & w6207) | (w3236 & w6207);
assign w2677 = (w6851 & w4529) | (w6851 & w1000) | (w4529 & w1000);
assign w2678 = w3128 & ~w2706;
assign w2679 = w4272 | w5513;
assign w2680 = (w1609 & w2626) | (w1609 & w3533) | (w2626 & w3533);
assign w2681 = w3488 & w4419;
assign w2682 = w4317 & ~w1265;
assign w2683 = (w1683 & w1518) | (w1683 & ~w6174) | (w1518 & ~w6174);
assign w2684 = ~w7218 & w2808;
assign w2685 = ~w4038 & ~w6551;
assign w2686 = ~w3391 & w4480;
assign w2687 = ~w6647 & ~w541;
assign w2688 = a91 & b91;
assign w2689 = w4375 & w1543;
assign w2690 = w5559 & ~w867;
assign w2691 = (w6100 & w2527) | (w6100 & w720) | (w2527 & w720);
assign w2692 = ~w7647 & ~w4299;
assign w2693 = ~w7137 & ~w3351;
assign w2694 = ~w2522 & w1435;
assign w2695 = w5259 & w7209;
assign w2696 = ~w2774 & ~w2860;
assign w2697 = (w6857 & w3664) | (w6857 & w2988) | (w3664 & w2988);
assign w2698 = (w2267 & w3432) | (w2267 & w7568) | (w3432 & w7568);
assign w2699 = ~w3306 & ~w728;
assign w2700 = w2969 & ~w6251;
assign w2701 = (~w3336 & w252) | (~w3336 & w1383) | (w252 & w1383);
assign w2702 = (w7346 & w3232) | (w7346 & ~w4418) | (w3232 & ~w4418);
assign w2703 = w2107 & ~w4802;
assign w2704 = ~w2513 & ~w2676;
assign w2705 = ~w331 & ~w3914;
assign w2706 = ~w5428 & ~w5937;
assign w2707 = w4499 & ~w3990;
assign w2708 = ~w1379 & w6834;
assign w2709 = ~w2566 & w3811;
assign w2710 = ~w5229 & w5683;
assign w2711 = (~w5325 & w742) | (~w5325 & w6075) | (w742 & w6075);
assign w2712 = ~w1216 & w6757;
assign w2713 = w3915 & w4071;
assign w2714 = ~w7365 & ~w7278;
assign w2715 = ~w991 & ~w1279;
assign w2716 = (w3461 & w4235) | (w3461 & w2239) | (w4235 & w2239);
assign w2717 = ~w6656 & ~w3122;
assign w2718 = ~a143 & ~b143;
assign w2719 = (w4145 & w480) | (w4145 & w7624) | (w480 & w7624);
assign w2720 = ~w2558 & ~w4457;
assign w2721 = ~w6564 & w7022;
assign w2722 = ~w2257 & ~w6099;
assign w2723 = (w699 & w455) | (w699 & ~w6152) | (w455 & ~w6152);
assign w2724 = ~b0 & ~a0;
assign w2725 = ~a217 & ~b217;
assign w2726 = (~w2052 & w7129) | (~w2052 & w7029) | (w7129 & w7029);
assign w2727 = ~w2041 & ~w2996;
assign w2728 = ~w1004 & ~w3320;
assign w2729 = (~w3852 & w4117) | (~w3852 & w1418) | (w4117 & w1418);
assign w2730 = ~w1921 & ~w5455;
assign w2731 = (w6225 & w5278) | (w6225 & w1258) | (w5278 & w1258);
assign w2732 = (~w6566 & w4855) | (~w6566 & w5916) | (w4855 & w5916);
assign w2733 = ~w2001 & w2954;
assign w2734 = w3933 & ~w6981;
assign w2735 = ~a157 & ~b157;
assign w2736 = (w3736 & w5606) | (w3736 & w6903) | (w5606 & w6903);
assign w2737 = (~w1779 & w6095) | (~w1779 & w4984) | (w6095 & w4984);
assign w2738 = (w5257 & w4205) | (w5257 & w5221) | (w4205 & w5221);
assign w2739 = ~w2173 & ~w1632;
assign w2740 = ~w6753 & ~w3212;
assign w2741 = ~w902 & w3298;
assign w2742 = (w5178 & w6950) | (w5178 & w137) | (w6950 & w137);
assign w2743 = (~w5325 & w4186) | (~w5325 & w1238) | (w4186 & w1238);
assign w2744 = w7350 & ~w7622;
assign w2745 = (w3490 & w2360) | (w3490 & w4099) | (w2360 & w4099);
assign w2746 = (~w651 & w5848) | (~w651 & ~w2221) | (w5848 & ~w2221);
assign w2747 = ~w257 & ~w5829;
assign w2748 = (~w2179 & w3866) | (~w2179 & w1526) | (w3866 & w1526);
assign w2749 = ~a64 & ~b64;
assign w2750 = ~w4775 & ~w6964;
assign w2751 = a250 & b250;
assign w2752 = (~w3640 & w1018) | (~w3640 & w3628) | (w1018 & w3628);
assign w2753 = w3848 & ~w3989;
assign w2754 = ~w1950 & ~w339;
assign w2755 = (w702 & w1696) | (w702 & w2013) | (w1696 & w2013);
assign w2756 = (w4092 & w1936) | (w4092 & w7258) | (w1936 & w7258);
assign w2757 = w2497 & ~w5057;
assign w2758 = ~w1895 & ~w1055;
assign w2759 = ~w1384 & ~w736;
assign w2760 = (w6657 & w2159) | (w6657 & ~w563) | (w2159 & ~w563);
assign w2761 = (~w6738 & w7263) | (~w6738 & w4452) | (w7263 & w4452);
assign w2762 = (~w6714 & w3642) | (~w6714 & w4176) | (w3642 & w4176);
assign w2763 = ~w2600 & ~w4402;
assign w2764 = ~w4976 & ~w476;
assign w2765 = w4778 & ~w6339;
assign w2766 = w3197 & w1006;
assign w2767 = ~w1601 & ~w129;
assign w2768 = (w3318 & w2760) | (w3318 & w3346) | (w2760 & w3346);
assign w2769 = w5350 & ~w5862;
assign w2770 = ~w3654 & w169;
assign w2771 = (w2985 & w3544) | (w2985 & w5488) | (w3544 & w5488);
assign w2772 = w6481 & ~w732;
assign w2773 = (w6844 & w2845) | (w6844 & w1341) | (w2845 & w1341);
assign w2774 = ~w2394 & ~w295;
assign w2775 = w1296 & w3060;
assign w2776 = (w3805 & w4751) | (w3805 & w1738) | (w4751 & w1738);
assign w2777 = ~w2041 & w200;
assign w2778 = ~w6714 & ~w875;
assign w2779 = ~w7618 & ~w1667;
assign w2780 = (w4385 & w1918) | (w4385 & ~w5098) | (w1918 & ~w5098);
assign w2781 = (~w4875 & ~w4598) | (~w4875 & w1969) | (~w4598 & w1969);
assign w2782 = ~w4438 & w7172;
assign w2783 = ~w7167 & ~w5741;
assign w2784 = w306 & w6800;
assign w2785 = ~w2678 & ~w5993;
assign w2786 = ~w787 & ~w5383;
assign w2787 = w813 & ~w6286;
assign w2788 = w1607 & w719;
assign w2789 = (w7024 & w7443) | (w7024 & w632) | (w7443 & w632);
assign w2790 = ~w5783 & w2937;
assign w2791 = (w5217 & w4986) | (w5217 & ~w6174) | (w4986 & ~w6174);
assign w2792 = (w5986 & w5901) | (w5986 & w7133) | (w5901 & w7133);
assign w2793 = ~w5759 & w3741;
assign w2794 = (w856 & w4610) | (w856 & w3201) | (w4610 & w3201);
assign w2795 = (~w4123 & w6614) | (~w4123 & ~w3847) | (w6614 & ~w3847);
assign w2796 = ~w2708 & w1745;
assign w2797 = (w1067 & ~w488) | (w1067 & w6093) | (~w488 & w6093);
assign w2798 = w2557 & w944;
assign w2799 = ~w7427 & w2145;
assign w2800 = ~w1176 & ~w3854;
assign w2801 = w3656 & ~w5859;
assign w2802 = (~w7199 & w7569) | (~w7199 & w6316) | (w7569 & w6316);
assign w2803 = ~a10 & ~b10;
assign w2804 = (w3201 & w5619) | (w3201 & ~w2456) | (w5619 & ~w2456);
assign w2805 = (~w3903 & w7197) | (~w3903 & w6134) | (w7197 & w6134);
assign w2806 = ~w174 & w6688;
assign w2807 = (w6600 & w1473) | (w6600 & ~w5511) | (w1473 & ~w5511);
assign w2808 = w5686 & ~w5807;
assign w2809 = ~w3107 & w5346;
assign w2810 = ~w4867 & w6499;
assign w2811 = ~w2586 & ~w4891;
assign w2812 = ~w3229 & ~w6797;
assign w2813 = ~w2108 & w5912;
assign w2814 = ~w57 & ~w6211;
assign w2815 = (~w5466 & ~w424) | (~w5466 & w5996) | (~w424 & w5996);
assign w2816 = ~w1739 & w321;
assign w2817 = ~w3950 & ~w6474;
assign w2818 = w6854 & ~w101;
assign w2819 = ~w5015 & w3745;
assign w2820 = w6643 & ~w1463;
assign w2821 = w6684 & ~w6394;
assign w2822 = (w5655 & w4502) | (w5655 & w5450) | (w4502 & w5450);
assign w2823 = (~w1877 & ~w2483) | (~w1877 & w1803) | (~w2483 & w1803);
assign w2824 = w3003 & w91;
assign w2825 = (w2570 & w7179) | (w2570 & ~w206) | (w7179 & ~w206);
assign w2826 = (w6499 & w6738) | (w6499 & w2810) | (w6738 & w2810);
assign w2827 = (w4828 & w2449) | (w4828 & w4276) | (w2449 & w4276);
assign w2828 = (~w7493 & w7205) | (~w7493 & w4124) | (w7205 & w4124);
assign w2829 = ~w2735 & ~w3482;
assign w2830 = (~w3903 & w3224) | (~w3903 & w6134) | (w3224 & w6134);
assign w2831 = (w829 & w7334) | (w829 & w5390) | (w7334 & w5390);
assign w2832 = ~w118 & w2494;
assign w2833 = w4749 & ~w4681;
assign w2834 = w5368 & ~w2985;
assign w2835 = (~w1321 & ~w2401) | (~w1321 & w3391) | (~w2401 & w3391);
assign w2836 = a109 & b109;
assign w2837 = (~w3336 & w252) | (~w3336 & w1377) | (w252 & w1377);
assign w2838 = ~w4146 & ~w4881;
assign w2839 = ~w6366 & w4147;
assign w2840 = ~w1831 & w6898;
assign w2841 = w2869 & ~w4867;
assign w2842 = (w1419 & w7180) | (w1419 & w4064) | (w7180 & w4064);
assign w2843 = (w7332 & w3767) | (w7332 & w542) | (w3767 & w542);
assign w2844 = w2609 & w7092;
assign w2845 = (w7429 & w5646) | (w7429 & w3365) | (w5646 & w3365);
assign w2846 = ~a80 & ~b80;
assign w2847 = ~w4803 & w144;
assign w2848 = (~w1851 & ~w6518) | (~w1851 & w675) | (~w6518 & w675);
assign w2849 = (w4327 & w4485) | (w4327 & w1558) | (w4485 & w1558);
assign w2850 = (~w406 & w7019) | (~w406 & ~w1611) | (w7019 & ~w1611);
assign w2851 = (~w6100 & w7430) | (~w6100 & w7254) | (w7430 & w7254);
assign w2852 = ~w2 & ~w1387;
assign w2853 = ~w3665 & ~w6169;
assign w2854 = (w7394 & w1527) | (w7394 & w318) | (w1527 & w318);
assign w2855 = ~w3351 & ~w3092;
assign w2856 = w2057 & w2687;
assign w2857 = w4384 & ~w4323;
assign w2858 = (w472 & w2709) | (w472 & w6445) | (w2709 & w6445);
assign w2859 = (~w2068 & w7205) | (~w2068 & w5050) | (w7205 & w5050);
assign w2860 = (w5655 & w2035) | (w5655 & w4557) | (w2035 & w4557);
assign w2861 = ~w5555 & w4875;
assign w2862 = ~w147 & ~w6766;
assign w2863 = ~w6087 & w7268;
assign w2864 = (~w5259 & w131) | (~w5259 & w2922) | (w131 & w2922);
assign w2865 = (~w1791 & w7444) | (~w1791 & w7576) | (w7444 & w7576);
assign w2866 = (w2188 & w2124) | (w2188 & w3648) | (w2124 & w3648);
assign w2867 = (w5229 & w3878) | (w5229 & w3862) | (w3878 & w3862);
assign w2868 = (~w1435 & w5819) | (~w1435 & ~w4190) | (w5819 & ~w4190);
assign w2869 = ~w5837 & w2624;
assign w2870 = (w6112 & w575) | (w6112 & w6641) | (w575 & w6641);
assign w2871 = ~w4680 & w6028;
assign w2872 = w6643 & ~w6609;
assign w2873 = ~w3909 & w2230;
assign w2874 = w7538 & w1171;
assign w2875 = ~w5622 & ~w6709;
assign w2876 = (w3063 & w1631) | (w3063 & w484) | (w1631 & w484);
assign w2877 = w666 & w3122;
assign w2878 = ~w7372 & w2067;
assign w2879 = w1606 & ~w1198;
assign w2880 = a199 & b199;
assign w2881 = w4036 & w426;
assign w2882 = w344 & ~w6301;
assign w2883 = ~w5557 & ~w6656;
assign w2884 = w3689 & ~w3932;
assign w2885 = (~w6025 & ~w318) | (~w6025 & w4163) | (~w318 & w4163);
assign w2886 = (~w412 & w5473) | (~w412 & w1410) | (w5473 & w1410);
assign w2887 = ~w1831 & ~w6225;
assign w2888 = a205 & b205;
assign w2889 = (w1555 & w6722) | (w1555 & w3014) | (w6722 & w3014);
assign w2890 = ~w4665 & w5352;
assign w2891 = w7461 & ~w3974;
assign w2892 = w6444 & ~w5573;
assign w2893 = (w5325 & w4093) | (w5325 & w4178) | (w4093 & w4178);
assign w2894 = w5403 & ~w6872;
assign w2895 = (~w2627 & w4483) | (~w2627 & w4032) | (w4483 & w4032);
assign w2896 = (~w2590 & w3866) | (~w2590 & w6514) | (w3866 & w6514);
assign w2897 = (~w6353 & w1405) | (~w6353 & w2369) | (w1405 & w2369);
assign w2898 = w1798 & w5655;
assign w2899 = w6545 & ~w2896;
assign w2900 = (~w4187 & w6365) | (~w4187 & w4361) | (w6365 & w4361);
assign w2901 = ~w6545 & w2896;
assign w2902 = w3677 & w1534;
assign w2903 = w6031 & w1129;
assign w2904 = w7162 & w4523;
assign w2905 = w3446 & w1252;
assign w2906 = w2221 & w6385;
assign w2907 = ~w576 & ~w5467;
assign w2908 = ~w2607 & ~w5769;
assign w2909 = (w3057 & w6831) | (w3057 & w329) | (w6831 & w329);
assign w2910 = (w6746 & w5898) | (w6746 & w6001) | (w5898 & w6001);
assign w2911 = (~w1611 & w5406) | (~w1611 & w2659) | (w5406 & w2659);
assign w2912 = (w6206 & ~w6226) | (w6206 & ~w7575) | (~w6226 & ~w7575);
assign w2913 = ~a34 & ~b34;
assign w2914 = a102 & b102;
assign w2915 = w5277 & w2862;
assign w2916 = ~w2185 & ~w7186;
assign w2917 = w999 & ~w7525;
assign w2918 = (~w7003 & w5024) | (~w7003 & w2071) | (w5024 & w2071);
assign w2919 = (w1455 & w6575) | (w1455 & w202) | (w6575 & w202);
assign w2920 = (w173 & w7252) | (w173 & w5208) | (w7252 & w5208);
assign w2921 = (~w7187 & w4634) | (~w7187 & w5160) | (w4634 & w5160);
assign w2922 = (~w1575 & w2483) | (~w1575 & w2985) | (w2483 & w2985);
assign w2923 = (w6353 & w4127) | (w6353 & w2235) | (w4127 & w2235);
assign w2924 = (w6419 & w5657) | (w6419 & ~w2641) | (w5657 & ~w2641);
assign w2925 = w4932 | w2862;
assign w2926 = (w90 & w4914) | (w90 & w1892) | (w4914 & w1892);
assign w2927 = (~w2627 & w4108) | (~w2627 & w4345) | (w4108 & w4345);
assign w2928 = ~w5229 & w291;
assign w2929 = w6689 & ~w4838;
assign w2930 = (~w6100 & w2022) | (~w6100 & w6014) | (w2022 & w6014);
assign w2931 = (w6633 & w1857) | (w6633 & w2442) | (w1857 & w2442);
assign w2932 = (~w7604 & w170) | (~w7604 & w7187) | (w170 & w7187);
assign w2933 = (w4075 & w5363) | (w4075 & w484) | (w5363 & w484);
assign w2934 = (w3892 & w2478) | (w3892 & w6812) | (w2478 & w6812);
assign w2935 = w7576 & ~w3391;
assign w2936 = (w2429 & w3401) | (w2429 & w6801) | (w3401 & w6801);
assign w2937 = ~w5937 & w2404;
assign w2938 = ~w6912 & ~w7384;
assign w2939 = (~w6614 & ~w1888) | (~w6614 & w2456) | (~w1888 & w2456);
assign w2940 = w347 & w3177;
assign w2941 = (~w6082 & w4086) | (~w6082 & w168) | (w4086 & w168);
assign w2942 = w2740 & w2795;
assign w2943 = (w5545 & w3532) | (w5545 & w3533) | (w3532 & w3533);
assign w2944 = (~w5522 & w3209) | (~w5522 & w1299) | (w3209 & w1299);
assign w2945 = ~a151 & ~b151;
assign w2946 = (w1074 & w5840) | (w1074 & ~w629) | (w5840 & ~w629);
assign w2947 = ~w990 & ~w2644;
assign w2948 = ~w4140 & ~w7097;
assign w2949 = (~w4296 & w6917) | (~w4296 & w6590) | (w6917 & w6590);
assign w2950 = (~w6272 & w122) | (~w6272 & w3830) | (w122 & w3830);
assign w2951 = ~w4578 & ~w305;
assign w2952 = w723 & ~w6224;
assign w2953 = ~w6064 & ~w1307;
assign w2954 = a12 & b12;
assign w2955 = w4505 & w2797;
assign w2956 = (~w5066 & w2178) | (~w5066 & w52) | (w2178 & w52);
assign w2957 = (w4825 & w5377) | (w4825 & w5243) | (w5377 & w5243);
assign w2958 = ~w4906 & w708;
assign w2959 = (~w6147 & w6259) | (~w6147 & w2206) | (w6259 & w2206);
assign w2960 = (~w3057 & w7617) | (~w3057 & w2980) | (w7617 & w2980);
assign w2961 = w106 & ~w4329;
assign w2962 = ~w628 & w7024;
assign w2963 = w3235 & ~w3869;
assign w2964 = w5555 & w860;
assign w2965 = ~w5827 & w2988;
assign w2966 = ~w6114 & w6504;
assign w2967 = ~w2671 & ~w3313;
assign w2968 = ~w3507 & w6528;
assign w2969 = ~w5239 & ~w5348;
assign w2970 = ~w1607 & w4660;
assign w2971 = (~w4765 & w4403) | (~w4765 & w2281) | (w4403 & w2281);
assign w2972 = (~w887 & ~w2339) | (~w887 & w6132) | (~w2339 & w6132);
assign w2973 = ~w1241 & ~w3066;
assign w2974 = (w2627 & w5748) | (w2627 & w3124) | (w5748 & w3124);
assign w2975 = ~w3840 & ~w6682;
assign w2976 = (~w6100 & w2756) | (~w6100 & w3287) | (w2756 & w3287);
assign w2977 = ~w1497 | ~w3070;
assign w2978 = ~w1656 & ~w3580;
assign w2979 = (w2103 & w6662) | (w2103 & w4292) | (w6662 & w4292);
assign w2980 = (w6600 & w1473) | (w6600 & ~w629) | (w1473 & ~w629);
assign w2981 = ~w4321 & w6898;
assign w2982 = (~w3774 & w1627) | (~w3774 & w160) | (w1627 & w160);
assign w2983 = (~w4710 & ~w6435) | (~w4710 & w4158) | (~w6435 & w4158);
assign w2984 = ~a161 & ~b161;
assign w2985 = ~w2557 & w5774;
assign w2986 = w1759 | w1344;
assign w2987 = ~w1241 & w2534;
assign w2988 = ~w5783 & w1757;
assign w2989 = (~w5056 & w7616) | (~w5056 & w831) | (w7616 & w831);
assign w2990 = (w615 & w1993) | (w615 & w555) | (w1993 & w555);
assign w2991 = (w821 & w7087) | (w821 & w3856) | (w7087 & w3856);
assign w2992 = (w2910 & w175) | (w2910 & w2456) | (w175 & w2456);
assign w2993 = (w3719 & w2182) | (w3719 & w6971) | (w2182 & w6971);
assign w2994 = w2257 & ~w1279;
assign w2995 = w5259 & w5288;
assign w2996 = a189 & b189;
assign w2997 = a196 & b196;
assign w2998 = w3868 & ~w3014;
assign w2999 = (w3784 & w2502) | (w3784 & w1730) | (w2502 & w1730);
assign w3000 = (~w5385 & w3483) | (~w5385 & w2939) | (w3483 & w2939);
assign w3001 = (w2678 & w5178) | (w2678 & w2020) | (w5178 & w2020);
assign w3002 = (~w4651 & w5553) | (~w4651 & w4152) | (w5553 & w4152);
assign w3003 = ~w7308 & w547;
assign w3004 = ~w6206 & w1234;
assign w3005 = (w978 & w6230) | (w978 & w4506) | (w6230 & w4506);
assign w3006 = (~w7493 & ~w6969) | (~w7493 & w4882) | (~w6969 & w4882);
assign w3007 = ~a175 & ~b175;
assign w3008 = (w632 & w568) | (w632 & w3057) | (w568 & w3057);
assign w3009 = (w6397 & ~w6966) | (w6397 & w4640) | (~w6966 & w4640);
assign w3010 = (w101 & ~w1728) | (w101 & w3655) | (~w1728 & w3655);
assign w3011 = w6883 & w7311;
assign w3012 = w242 & ~w5291;
assign w3013 = w3231 & ~w1886;
assign w3014 = ~a209 & ~b209;
assign w3015 = ~w7010 & w1343;
assign w3016 = ~w101 & ~w4648;
assign w3017 = ~w6776 & ~w6772;
assign w3018 = (~w615 & w4815) | (~w615 & w6642) | (w4815 & w6642);
assign w3019 = a90 & b90;
assign w3020 = (~w2068 & ~w6969) | (~w2068 & w1261) | (~w6969 & w1261);
assign w3021 = (w6100 & w4869) | (w6100 & w6615) | (w4869 & w6615);
assign w3022 = (w1346 & w3345) | (w1346 & w5442) | (w3345 & w5442);
assign w3023 = (~w5655 & w658) | (~w5655 & w3650) | (w658 & w3650);
assign w3024 = w3391 & w5806;
assign w3025 = w5403 & w1212;
assign w3026 = (w3983 & w5523) | (w3983 & w6959) | (w5523 & w6959);
assign w3027 = (w3472 & w5403) | (w3472 & ~w7197) | (w5403 & ~w7197);
assign w3028 = ~w6161 & w3994;
assign w3029 = (w3657 & w5587) | (w3657 & w1743) | (w5587 & w1743);
assign w3030 = ~w4206 & w2416;
assign w3031 = (w7383 & w6905) | (w7383 & w2800) | (w6905 & w2800);
assign w3032 = ~w3802 & ~w2643;
assign w3033 = ~a241 & ~b241;
assign w3034 = (w6942 & w6148) | (w6942 & ~w7450) | (w6148 & ~w7450);
assign w3035 = ~w234 & w3842;
assign w3036 = (w6217 & w7288) | (w6217 & ~w5464) | (w7288 & ~w5464);
assign w3037 = w1260 & ~w5346;
assign w3038 = ~w4991 & ~w5655;
assign w3039 = ~w5699 & w6351;
assign w3040 = ~w3359 & ~w3135;
assign w3041 = (~w5178 & w661) | (~w5178 & w6263) | (w661 & w6263);
assign w3042 = (w6467 & w5866) | (w6467 & w2802) | (w5866 & w2802);
assign w3043 = (~w3304 & ~w248) | (~w3304 & w2445) | (~w248 & w2445);
assign w3044 = w2560 & w6747;
assign w3045 = ~w1007 & ~w5782;
assign w3046 = (~w517 & ~w5912) | (~w517 & ~w7383) | (~w5912 & ~w7383);
assign w3047 = ~w6760 & w3267;
assign w3048 = w628 & w6733;
assign w3049 = (w2496 & ~w5392) | (w2496 & w477) | (~w5392 & w477);
assign w3050 = ~w5759 & w4891;
assign w3051 = ~w4881 & w385;
assign w3052 = ~a187 & ~b187;
assign w3053 = (w4392 & w1021) | (w4392 & w98) | (w1021 & w98);
assign w3054 = ~w2542 & w6202;
assign w3055 = ~w1849 & ~w164;
assign w3056 = (w3984 & w2222) | (w3984 & ~w6439) | (w2222 & ~w6439);
assign w3057 = ~w1607 & w671;
assign w3058 = w7634 & ~w593;
assign w3059 = w3843 | w6386;
assign w3060 = w2249 & w6512;
assign w3061 = ~w4921 & ~w1732;
assign w3062 = ~w1386 & ~w3183;
assign w3063 = w4598 & w2189;
assign w3064 = a81 & b81;
assign w3065 = w1661 & ~w4587;
assign w3066 = ~w2671 & ~w1327;
assign w3067 = ~w6920 & w4444;
assign w3068 = (w6738 & w6457) | (w6738 & w4701) | (w6457 & w4701);
assign w3069 = (w3952 & w3581) | (w3952 & w3068) | (w3581 & w3068);
assign w3070 = w6753 & ~w3212;
assign w3071 = (~w1455 & w2432) | (~w1455 & w6587) | (w2432 & w6587);
assign w3072 = a38 & b38;
assign w3073 = ~a69 & ~b69;
assign w3074 = (w5686 & ~w1356) | (w5686 & w6407) | (~w1356 & w6407);
assign w3075 = a32 & b32;
assign w3076 = (w7269 & w3005) | (w7269 & w484) | (w3005 & w484);
assign w3077 = (w4130 & w5951) | (w4130 & w4285) | (w5951 & w4285);
assign w3078 = ~w4811 & ~w3014;
assign w3079 = ~w7243 & w2294;
assign w3080 = ~w54 & w2179;
assign w3081 = (~w2179 & ~w6151) | (~w2179 & w586) | (~w6151 & w586);
assign w3082 = ~w7360 & w6454;
assign w3083 = ~w736 & ~w5864;
assign w3084 = (w4143 & w1692) | (w4143 & w6079) | (w1692 & w6079);
assign w3085 = (~w236 & w751) | (~w236 & w6998) | (w751 & w6998);
assign w3086 = (~w6100 & w2303) | (~w6100 & w3373) | (w2303 & w3373);
assign w3087 = ~w3732 & ~w4146;
assign w3088 = (w7028 & w5011) | (w7028 & w5385) | (w5011 & w5385);
assign w3089 = w5587 & w3657;
assign w3090 = (~w2081 & w3141) | (~w2081 & ~w1860) | (w3141 & ~w1860);
assign w3091 = (w7409 & w903) | (w7409 & ~w2456) | (w903 & ~w2456);
assign w3092 = a149 & b149;
assign w3093 = ~w7316 & ~w6842;
assign w3094 = w2872 & ~w6184;
assign w3095 = (~w5056 & w7616) | (~w5056 & w2717) | (w7616 & w2717);
assign w3096 = ~a19 & ~b19;
assign w3097 = (w2627 & w4779) | (w2627 & w754) | (w4779 & w754);
assign w3098 = (w1484 & w5150) | (w1484 & w5325) | (w5150 & w5325);
assign w3099 = (w5834 & w281) | (w5834 & w4782) | (w281 & w4782);
assign w3100 = ~w7391 & ~w4392;
assign w3101 = ~a202 & ~b202;
assign w3102 = w5445 & ~w1284;
assign w3103 = (~w5106 & w4716) | (~w5106 & ~w4499) | (w4716 & ~w4499);
assign w3104 = w1813 & ~w4010;
assign w3105 = ~w7012 & w4387;
assign w3106 = w2582 & ~w212;
assign w3107 = w318 & ~w3328;
assign w3108 = ~w5170 & ~w4940;
assign w3109 = ~w6561 & ~w5103;
assign w3110 = ~w6265 & w2516;
assign w3111 = w2861 & ~w5464;
assign w3112 = (w5054 & w823) | (w5054 & w6099) | (w823 & w6099);
assign w3113 = ~w728 & ~w4438;
assign w3114 = (w1936 & w2402) | (w1936 & w4856) | (w2402 & w4856);
assign w3115 = (w1609 & w2626) | (w1609 & w5368) | (w2626 & w5368);
assign w3116 = ~w1813 & w4010;
assign w3117 = ~w2295 & ~w4893;
assign w3118 = w1998 & w666;
assign w3119 = w412 & w1946;
assign w3120 = ~w4370 & ~w3589;
assign w3121 = (w544 & w5625) | (w544 & w5376) | (w5625 & w5376);
assign w3122 = ~a234 & ~b234;
assign w3123 = a192 & b192;
assign w3124 = ~w2853 & ~w1356;
assign w3125 = w4681 & w3519;
assign w3126 = (~w2649 & w7031) | (~w2649 & ~w5059) | (w7031 & ~w5059);
assign w3127 = w5111 & ~w1034;
assign w3128 = ~w5416 & ~w54;
assign w3129 = ~w3248 & w523;
assign w3130 = (w4537 & w5270) | (w4537 & ~w6174) | (w5270 & ~w6174);
assign w3131 = w649 & ~w2333;
assign w3132 = (~w5430 & w3832) | (~w5430 & w7511) | (w3832 & w7511);
assign w3133 = ~w7278 & ~w2278;
assign w3134 = ~w4306 & w5106;
assign w3135 = a26 & b26;
assign w3136 = ~w471 & ~w5230;
assign w3137 = ~a103 & ~b103;
assign w3138 = ~w3266 & ~w6094;
assign w3139 = ~w314 & w1344;
assign w3140 = (w3490 & w289) | (w3490 & w4534) | (w289 & w4534);
assign w3141 = w1300 & ~w2081;
assign w3142 = w4918 & ~w6149;
assign w3143 = (~w5257 & w6369) | (~w5257 & w2091) | (w6369 & w2091);
assign w3144 = w3082 & w2017;
assign w3145 = w4448 & ~w4499;
assign w3146 = w6558 & ~w7471;
assign w3147 = w1338 & ~w3576;
assign w3148 = w6452 & ~w7302;
assign w3149 = (w65 & w4938) | (w65 & w4803) | (w4938 & w4803);
assign w3150 = w6760 & ~w4185;
assign w3151 = (w2849 & w2455) | (w2849 & w6511) | (w2455 & w6511);
assign w3152 = ~w4168 & ~w3607;
assign w3153 = (~w6922 & w7154) | (~w6922 & w813) | (w7154 & w813);
assign w3154 = (w639 & w3036) | (w639 & w310) | (w3036 & w310);
assign w3155 = w6415 & w3819;
assign w3156 = w7319 & w2832;
assign w3157 = ~w4545 & w5349;
assign w3158 = w1441 & ~w4174;
assign w3159 = w270 & w1658;
assign w3160 = ~w6539 & ~w6927;
assign w3161 = w174 & w2970;
assign w3162 = ~w1862 & w7007;
assign w3163 = (~w4648 & w6046) | (~w4648 & w5172) | (w6046 & w5172);
assign w3164 = ~w2011 & w2179;
assign w3165 = ~w7408 & w6712;
assign w3166 = a24 & b24;
assign w3167 = a6 & b6;
assign w3168 = ~w100 & w1030;
assign w3169 = ~w1142 & ~w4492;
assign w3170 = (~w4647 & w3639) | (~w4647 & w2949) | (w3639 & w2949);
assign w3171 = (w4327 & w4560) | (w4327 & w2377) | (w4560 & w2377);
assign w3172 = ~w3007 & ~w391;
assign w3173 = ~w4921 & ~w4377;
assign w3174 = (w2627 & w211) | (w2627 & w5869) | (w211 & w5869);
assign w3175 = (~w5914 & w4025) | (~w5914 & w1379) | (w4025 & w1379);
assign w3176 = a19 & b19;
assign w3177 = ~w1030 & w3922;
assign w3178 = w5555 & w6357;
assign w3179 = w301 & w893;
assign w3180 = ~w3744 & ~w5994;
assign w3181 = w3240 & w3298;
assign w3182 = (~w5325 & w1296) | (~w5325 & w6034) | (w1296 & w6034);
assign w3183 = a174 & b174;
assign w3184 = (~w5484 & w4493) | (~w5484 & w7410) | (w4493 & w7410);
assign w3185 = w5948 & w1434;
assign w3186 = ~w4863 & w7200;
assign w3187 = (~w3471 & w6685) | (~w3471 & w1182) | (w6685 & w1182);
assign w3188 = ~w2197 & ~w2286;
assign w3189 = w3288 & w2085;
assign w3190 = (~w5834 & w6907) | (~w5834 & w1640) | (w6907 & w1640);
assign w3191 = (~w1103 & w1811) | (~w1103 & w177) | (w1811 & w177);
assign w3192 = w6206 & ~w1712;
assign w3193 = w5933 & w5843;
assign w3194 = (~w2740 & ~w671) | (~w2740 & w3653) | (~w671 & w3653);
assign w3195 = ~w2645 & w5882;
assign w3196 = w2049 & ~w3269;
assign w3197 = w4459 & ~w7187;
assign w3198 = (~w1193 & w1361) | (~w1193 & w5315) | (w1361 & w5315);
assign w3199 = w7365 & ~w3455;
assign w3200 = ~w6458 & ~w7394;
assign w3201 = w1071 & w6592;
assign w3202 = ~w6713 & ~w7146;
assign w3203 = ~w7044 & w3014;
assign w3204 = w3547 & w2572;
assign w3205 = (w1266 & w5830) | (w1266 & w621) | (w5830 & w621);
assign w3206 = ~w3712 & w3051;
assign w3207 = ~a92 & ~b92;
assign w3208 = (w2037 & w7085) | (w2037 & w7250) | (w7085 & w7250);
assign w3209 = w7150 & ~w1519;
assign w3210 = ~w1999 & ~w6884;
assign w3211 = (~w5655 & w2923) | (~w5655 & w3325) | (w2923 & w3325);
assign w3212 = a238 & b238;
assign w3213 = w4754 & w994;
assign w3214 = (~w788 & w4567) | (~w788 & ~w6129) | (w4567 & ~w6129);
assign w3215 = ~w2836 & ~w3799;
assign w3216 = (w5506 & w96) | (w5506 & w5655) | (w96 & w5655);
assign w3217 = a77 & b77;
assign w3218 = (~w6966 & w7068) | (~w6966 & w3270) | (w7068 & w3270);
assign w3219 = ~w3217 & ~w884;
assign w3220 = (w501 & w3806) | (w501 & w4356) | (w3806 & w4356);
assign w3221 = w3152 & ~w1974;
assign w3222 = (w2627 & w6074) | (w2627 & w6750) | (w6074 & w6750);
assign w3223 = w4238 & ~w2433;
assign w3224 = (~w4911 & w5503) | (~w4911 & w1986) | (w5503 & w1986);
assign w3225 = (~w2456 & w4233) | (~w2456 & w4955) | (w4233 & w4955);
assign w3226 = ~w5403 & w3278;
assign w3227 = ~w4797 & ~w3308;
assign w3228 = w4510 & w5747;
assign w3229 = ~w2033 & w895;
assign w3230 = (w6106 & w1564) | (w6106 & w6993) | (w1564 & w6993);
assign w3231 = ~w5616 & w3269;
assign w3232 = w2803 & w7346;
assign w3233 = ~w676 & w2973;
assign w3234 = (w7330 & w5016) | (w7330 & w484) | (w5016 & w484);
assign w3235 = b255 & a255;
assign w3236 = (w4995 & w4675) | (w4995 & w856) | (w4675 & w856);
assign w3237 = (w5655 & w645) | (w5655 & w2193) | (w645 & w2193);
assign w3238 = (w1886 & w7070) | (w1886 & w1818) | (w7070 & w1818);
assign w3239 = w3158 & ~w1085;
assign w3240 = ~w2216 & w1195;
assign w3241 = ~w535 & ~w221;
assign w3242 = w2460 & ~w4333;
assign w3243 = (~w6100 & w2690) | (~w6100 & w2424) | (w2690 & w2424);
assign w3244 = a202 & b202;
assign w3245 = (w1338 & ~w7072) | (w1338 & w6617) | (~w7072 & w6617);
assign w3246 = (w1751 & w7195) | (w1751 & w7163) | (w7195 & w7163);
assign w3247 = ~w1866 & ~w4480;
assign w3248 = a220 & b220;
assign w3249 = w4637 & w2482;
assign w3250 = (w3074 & w6905) | (w3074 & w2800) | (w6905 & w2800);
assign w3251 = (w972 & ~w7429) | (w972 & ~w927) | (~w7429 & ~w927);
assign w3252 = ~a140 & ~b140;
assign w3253 = w2286 | ~w3669;
assign w3254 = w2433 & w7417;
assign w3255 = w1364 & ~w1449;
assign w3256 = ~w3137 & ~w2260;
assign w3257 = w3888 & w837;
assign w3258 = ~w3192 & w6427;
assign w3259 = (~w1722 & w7562) | (~w1722 & w2013) | (w7562 & w2013);
assign w3260 = (w777 & w6309) | (w777 & w62) | (w6309 & w62);
assign w3261 = (w4521 & w6442) | (w4521 & w5414) | (w6442 & w5414);
assign w3262 = ~a132 & ~b132;
assign w3263 = w2829 & ~w226;
assign w3264 = (w7629 & w924) | (w7629 & w5778) | (w924 & w5778);
assign w3265 = w2094 & ~w7453;
assign w3266 = ~a170 & ~b170;
assign w3267 = ~w4185 & ~w2997;
assign w3268 = (w2563 & w3168) | (w2563 & w799) | (w3168 & w799);
assign w3269 = ~w7097 & ~w2283;
assign w3270 = (w3306 & ~w1165) | (w3306 & ~w7520) | (~w1165 & ~w7520);
assign w3271 = ~w2838 | w5636;
assign w3272 = w3558 & w819;
assign w3273 = w7565 & w6113;
assign w3274 = (w5655 & w172) | (w5655 & w1041) | (w172 & w1041);
assign w3275 = ~w684 & ~w5539;
assign w3276 = (w615 & w4566) | (w615 & w404) | (w4566 & w404);
assign w3277 = w4991 & w6071;
assign w3278 = (w3078 & w5149) | (w3078 & w964) | (w5149 & w964);
assign w3279 = (~w5178 & w3226) | (~w5178 & w423) | (w3226 & w423);
assign w3280 = ~w5281 & w1723;
assign w3281 = (~w4176 & w4479) | (~w4176 & w3679) | (w4479 & w3679);
assign w3282 = ~w4808 & ~w1635;
assign w3283 = w1770 & w5204;
assign w3284 = (w1435 & ~w2522) | (w1435 & w1215) | (~w2522 & w1215);
assign w3285 = w2173 & ~w7648;
assign w3286 = (~w5257 & w5868) | (~w5257 & w5494) | (w5868 & w5494);
assign w3287 = w3113 & w5517;
assign w3288 = (w1759 & w1344) | (w1759 & ~w2401) | (w1344 & ~w2401);
assign w3289 = ~w3771 & w2739;
assign w3290 = ~w2914 & ~w7522;
assign w3291 = ~w5463 & w2068;
assign w3292 = ~w3075 & w129;
assign w3293 = (w3491 & w4539) | (w3491 & w4893) | (w4539 & w4893);
assign w3294 = ~a225 & ~b225;
assign w3295 = ~w2001 & ~w7407;
assign w3296 = (w3511 & w1167) | (w3511 & w6645) | (w1167 & w6645);
assign w3297 = w5370 & ~w615;
assign w3298 = ~w5348 & w4741;
assign w3299 = (~w372 & w7416) | (~w372 & w4686) | (w7416 & w4686);
assign w3300 = w4375 & ~w3730;
assign w3301 = ~w2407 & w5222;
assign w3302 = ~w2173 & w6524;
assign w3303 = ~w7450 & w6423;
assign w3304 = ~w2493 & ~w1380;
assign w3305 = (~w3986 & w4628) | (~w3986 & w4221) | (w4628 & w4221);
assign w3306 = ~a109 & ~b109;
assign w3307 = (w2842 & w7331) | (w2842 & ~w2876) | (w7331 & ~w2876);
assign w3308 = (~w5178 & w4541) | (~w5178 & w2711) | (w4541 & w2711);
assign w3309 = (w5672 & ~w6846) | (w5672 & ~w4647) | (~w6846 & ~w4647);
assign w3310 = (w7394 & w1527) | (w7394 & w2520) | (w1527 & w2520);
assign w3311 = ~w6444 & ~w5128;
assign w3312 = ~a53 & ~b53;
assign w3313 = w1241 & ~w1327;
assign w3314 = w4459 & w6397;
assign w3315 = (w7506 & w4177) | (w7506 & w632) | (w4177 & w632);
assign w3316 = (w7448 & w5165) | (w7448 & ~w2876) | (w5165 & ~w2876);
assign w3317 = (w2097 & w7252) | (w2097 & w5208) | (w7252 & w5208);
assign w3318 = (w2627 & w1770) | (w2627 & w5395) | (w1770 & w5395);
assign w3319 = ~w7399 & ~w5693;
assign w3320 = a211 & b211;
assign w3321 = w91 & w4257;
assign w3322 = (w6334 & w1885) | (w6334 & ~w7015) | (w1885 & ~w7015);
assign w3323 = ~w1621 & ~w1080;
assign w3324 = w3843 & w6386;
assign w3325 = (w7205 & w3550) | (w7205 & w4127) | (w3550 & w4127);
assign w3326 = (~w6100 & w5096) | (~w6100 & w6287) | (w5096 & w6287);
assign w3327 = w4188 & w6174;
assign w3328 = a62 & b62;
assign w3329 = (~w6594 & w6956) | (~w6594 & w7453) | (w6956 & w7453);
assign w3330 = w5430 & w6566;
assign w3331 = ~w2104 & ~w3248;
assign w3332 = ~w2291 & ~w145;
assign w3333 = w2558 & w6804;
assign w3334 = (w3868 & ~w6927) | (w3868 & w2998) | (~w6927 & w2998);
assign w3335 = (w615 & w1823) | (w615 & w724) | (w1823 & w724);
assign w3336 = ~w4412 & ~w1925;
assign w3337 = w1452 & w7626;
assign w3338 = (~w5325 & w2736) | (~w5325 & w1282) | (w2736 & w1282);
assign w3339 = (~w887 & w6872) | (~w887 & w5899) | (w6872 & w5899);
assign w3340 = (w6140 & w4410) | (w6140 & ~w6633) | (w4410 & ~w6633);
assign w3341 = w2318 & w1036;
assign w3342 = (w1843 & w5402) | (w1843 & w4380) | (w5402 & w4380);
assign w3343 = (w1458 & w4665) | (w1458 & ~w723) | (w4665 & ~w723);
assign w3344 = w3365 & ~w3264;
assign w3345 = ~w2913 & ~w6860;
assign w3346 = (w6657 & w2159) | (w6657 & ~w5291) | (w2159 & ~w5291);
assign w3347 = (w2051 & w626) | (w2051 & w1480) | (w626 & w1480);
assign w3348 = (w334 & w5402) | (w334 & w2657) | (w5402 & w2657);
assign w3349 = ~w990 & w4149;
assign w3350 = w4688 & ~w5420;
assign w3351 = a148 & b148;
assign w3352 = w56 & ~w5198;
assign w3353 = ~w5496 & ~w7289;
assign w3354 = ~w1837 & w6096;
assign w3355 = (w6100 & w6502) | (w6100 & w6077) | (w6502 & w6077);
assign w3356 = w5122 & w3706;
assign w3357 = ~w2750 & w5035;
assign w3358 = w7158 & ~w817;
assign w3359 = ~a26 & ~b26;
assign w3360 = w5965 & ~w5032;
assign w3361 = (w6475 & w1064) | (w6475 & ~w6501) | (w1064 & ~w6501);
assign w3362 = ~w6210 & ~w3052;
assign w3363 = (w5808 & ~w5486) | (w5808 & ~w2041) | (~w5486 & ~w2041);
assign w3364 = (w7648 & ~w3285) | (w7648 & ~w2409) | (~w3285 & ~w2409);
assign w3365 = ~w972 & ~w3217;
assign w3366 = w7291 & ~w5467;
assign w3367 = (w3218 & w5307) | (w3218 & w5094) | (w5307 & w5094);
assign w3368 = (w5834 & w4192) | (w5834 & w4649) | (w4192 & w4649);
assign w3369 = (w4102 & w2436) | (w4102 & w5209) | (w2436 & w5209);
assign w3370 = w4843 & ~w593;
assign w3371 = (w5834 & w333) | (w5834 & w192) | (w333 & w192);
assign w3372 = (~w6100 & w6815) | (~w6100 & w5904) | (w6815 & w5904);
assign w3373 = (w2393 & w1147) | (w2393 & w3892) | (w1147 & w3892);
assign w3374 = ~w2456 | ~w3847;
assign w3375 = ~w5295 & w453;
assign w3376 = (w3986 & w4714) | (w3986 & w5546) | (w4714 & w5546);
assign w3377 = (w1834 & w7225) | (w1834 & w2013) | (w7225 & w2013);
assign w3378 = (w7346 & w3232) | (w7346 & w6504) | (w3232 & w6504);
assign w3379 = (~w3444 & w4986) | (~w3444 & w647) | (w4986 & w647);
assign w3380 = (w3848 & w2263) | (w3848 & ~w5871) | (w2263 & ~w5871);
assign w3381 = w6366 & w5773;
assign w3382 = w7026 & ~w5289;
assign w3383 = (w3728 & w974) | (w3728 & ~w1607) | (w974 & ~w1607);
assign w3384 = ~w4148 & ~w6319;
assign w3385 = (w2686 & w30) | (w2686 & w4572) | (w30 & w4572);
assign w3386 = ~w208 & ~w2610;
assign w3387 = (~w248 & w4331) | (~w248 & w6471) | (w4331 & w6471);
assign w3388 = (w7346 & w3232) | (w7346 & w2966) | (w3232 & w2966);
assign w3389 = w6422 & ~w7355;
assign w3390 = ~w4253 & ~w4810;
assign w3391 = w4843 & w5948;
assign w3392 = a25 & b25;
assign w3393 = w4988 & w414;
assign w3394 = w5958 & w887;
assign w3395 = ~w5717 & ~w1983;
assign w3396 = ~w84 & w7016;
assign w3397 = w1792 & w1211;
assign w3398 = ~w6854 & ~w7453;
assign w3399 = ~w2172 & w1073;
assign w3400 = ~w1199 & ~w7533;
assign w3401 = w5236 & ~w129;
assign w3402 = (~w3461 & ~w5371) | (~w3461 & ~w6152) | (~w5371 & ~w6152);
assign w3403 = (w5257 & w4129) | (w5257 & w2341) | (w4129 & w2341);
assign w3404 = ~w1876 & ~w930;
assign w3405 = ~w6265 & w4376;
assign w3406 = w2254 & ~w5788;
assign w3407 = (~w5944 & w2110) | (~w5944 & w5565) | (w2110 & w5565);
assign w3408 = (w1227 & w5402) | (w1227 & w2000) | (w5402 & w2000);
assign w3409 = ~w2295 & w4661;
assign w3410 = w4802 & ~w978;
assign w3411 = w2596 & ~w1431;
assign w3412 = w7471 & w6876;
assign w3413 = w3421 & w2361;
assign w3414 = (w5078 & w1482) | (w5078 & w1681) | (w1482 & w1681);
assign w3415 = ~w332 & ~w4677;
assign w3416 = (~w6100 & w3705) | (~w6100 & w5114) | (w3705 & w5114);
assign w3417 = w666 & ~w2274;
assign w3418 = ~a180 & ~b180;
assign w3419 = (w6680 & w2248) | (w6680 & w4571) | (w2248 & w4571);
assign w3420 = (w6100 & w5973) | (w6100 & w5956) | (w5973 & w5956);
assign w3421 = (~w766 & ~w795) | (~w766 & ~w2401) | (~w795 & ~w2401);
assign w3422 = (~w3587 & w6265) | (~w3587 & w1629) | (w6265 & w1629);
assign w3423 = ~w2836 & w3218;
assign w3424 = w6960 & w588;
assign w3425 = ~w6473 & ~w6926;
assign w3426 = ~w7581 & ~w7221;
assign w3427 = ~w2253 & ~w4010;
assign w3428 = (w5178 & w6699) | (w5178 & w3230) | (w6699 & w3230);
assign w3429 = (w2627 & w5300) | (w2627 & w1997) | (w5300 & w1997);
assign w3430 = ~w790 & ~w1938;
assign w3431 = ~w4967 & w6893;
assign w3432 = w3957 & ~w5478;
assign w3433 = ~w164 & ~w5251;
assign w3434 = (~w6524 & w2409) | (~w6524 & w663) | (w2409 & w663);
assign w3435 = w54 & ~w3052;
assign w3436 = w5066 & ~w2274;
assign w3437 = w2735 & ~w351;
assign w3438 = (w1332 & ~w3057) | (w1332 & w3779) | (~w3057 & w3779);
assign w3439 = ~w5177 & ~w7609;
assign w3440 = w6033 & ~w4618;
assign w3441 = ~w3488 & w3061;
assign w3442 = (~w2603 & w495) | (~w2603 & w2854) | (w495 & w2854);
assign w3443 = (w4222 & w7385) | (w4222 & w6678) | (w7385 & w6678);
assign w3444 = ~w7221 & ~w6854;
assign w3445 = (w6082 & w3827) | (w6082 & w1425) | (w3827 & w1425);
assign w3446 = w4898 & ~w5926;
assign w3447 = (~w2849 & w5977) | (~w2849 & w766) | (w5977 & w766);
assign w3448 = w2471 & w6462;
assign w3449 = w2557 & ~w6254;
assign w3450 = a20 & b20;
assign w3451 = ~w5999 & ~w5802;
assign w3452 = (w5178 & w6546) | (w5178 & w4627) | (w6546 & w4627);
assign w3453 = (~w3292 & ~w6451) | (~w3292 & w1516) | (~w6451 & w1516);
assign w3454 = (~w2123 & w3814) | (~w2123 & w4277) | (w3814 & w4277);
assign w3455 = ~a181 & ~b181;
assign w3456 = ~w5972 & w2336;
assign w3457 = ~w5992 & ~w1433;
assign w3458 = w2819 & w135;
assign w3459 = w6571 & ~w736;
assign w3460 = (w5834 & w598) | (w5834 & w6823) | (w598 & w6823);
assign w3461 = (w5368 & w2741) | (w5368 & w3749) | (w2741 & w3749);
assign w3462 = ~a126 & ~b126;
assign w3463 = ~w6376 & ~w3874;
assign w3464 = ~w3190 & ~w4879;
assign w3465 = w2295 & w4893;
assign w3466 = w5333 & w6692;
assign w3467 = ~w6979 & ~w2285;
assign w3468 = w4175 & ~w3113;
assign w3469 = w5005 & ~w7632;
assign w3470 = w4257 & w4280;
assign w3471 = ~a136 & ~b136;
assign w3472 = ~w7197 & w3556;
assign w3473 = (~w5772 & w5633) | (~w5772 & w7456) | (w5633 & w7456);
assign w3474 = ~w693 & ~w6774;
assign w3475 = ~w3191 & ~w12;
assign w3476 = w3282 & ~w3963;
assign w3477 = (~w7008 & w2205) | (~w7008 & w282) | (w2205 & w282);
assign w3478 = (w1455 & w4556) | (w1455 & w3968) | (w4556 & w3968);
assign w3479 = (w6593 & w2776) | (w6593 & ~w6174) | (w2776 & ~w6174);
assign w3480 = ~a166 & ~b166;
assign w3481 = w2171 & ~w2767;
assign w3482 = a157 & b157;
assign w3483 = ~w6614 | ~w1888;
assign w3484 = w7647 & ~w5404;
assign w3485 = (w6053 & w1347) | (w6053 & w3332) | (w1347 & w3332);
assign w3486 = ~w1709 & ~w5565;
assign w3487 = w6714 & w1269;
assign w3488 = (~w51 & ~w1587) | (~w51 & w3497) | (~w1587 & w3497);
assign w3489 = (~w144 & w5946) | (~w144 & w852) | (w5946 & w852);
assign w3490 = ~w2486 & ~w2270;
assign w3491 = (~w6106 & w4663) | (~w6106 & w2247) | (w4663 & w2247);
assign w3492 = ~w4289 & ~w7399;
assign w3493 = w2513 & w4675;
assign w3494 = (w1076 & w923) | (w1076 & ~w6100) | (w923 & ~w6100);
assign w3495 = ~w1569 & ~w5817;
assign w3496 = (w4995 & w1810) | (w4995 & w3493) | (w1810 & w3493);
assign w3497 = ~w6553 & ~w51;
assign w3498 = w2146 | w4609;
assign w3499 = (w4726 & w19) | (w4726 & ~w2013) | (w19 & ~w2013);
assign w3500 = ~w625 & w3365;
assign w3501 = ~w1563 & w665;
assign w3502 = (w304 & w1941) | (w304 & ~w484) | (w1941 & ~w484);
assign w3503 = ~w2260 & ~w1901;
assign w3504 = (~w887 & w6872) | (~w887 & w67) | (w6872 & w67);
assign w3505 = (~w5698 & w3500) | (~w5698 & w6767) | (w3500 & w6767);
assign w3506 = w5380 & ~w1730;
assign w3507 = w6426 & ~w7384;
assign w3508 = w4088 & ~w1678;
assign w3509 = w1954 & ~w7563;
assign w3510 = w1304 & w899;
assign w3511 = w2649 & w4204;
assign w3512 = ~a3 & ~b3;
assign w3513 = (w236 & w2931) | (w236 & w2194) | (w2931 & w2194);
assign w3514 = ~w6046 & w4594;
assign w3515 = (~w3266 & ~w1911) | (~w3266 & w7338) | (~w1911 & w7338);
assign w3516 = (~w6019 & w6412) | (~w6019 & w4076) | (w6412 & w4076);
assign w3517 = w4795 & ~w2097;
assign w3518 = (w4966 & ~w5190) | (w4966 & ~w2214) | (~w5190 & ~w2214);
assign w3519 = (~w4966 & w5190) | (~w4966 & w2214) | (w5190 & w2214);
assign w3520 = (w935 & w2008) | (w935 & w996) | (w2008 & w996);
assign w3521 = (~w3138 & w3023) | (~w3138 & w4119) | (w3023 & w4119);
assign w3522 = (~w2627 & w240) | (~w2627 & w6737) | (w240 & w6737);
assign w3523 = ~w2452 & w2763;
assign w3524 = ~w4448 & w46;
assign w3525 = ~w4004 & w2693;
assign w3526 = (~w5178 & w7380) | (~w5178 & w4814) | (w7380 & w4814);
assign w3527 = w5058 & w2766;
assign w3528 = ~w7146 & ~w5287;
assign w3529 = (~w2649 & w7031) | (~w2649 & w664) | (w7031 & w664);
assign w3530 = ~w6149 & w6100;
assign w3531 = ~w4564 & ~w2456;
assign w3532 = (~w1158 & w6299) | (~w1158 & ~w1903) | (w6299 & ~w1903);
assign w3533 = (w5259 & w3461) | (w5259 & w2834) | (w3461 & w2834);
assign w3534 = ~w3989 & w4478;
assign w3535 = ~w3415 & ~w4710;
assign w3536 = ~w4651 & ~w4328;
assign w3537 = (w4840 & w1111) | (w4840 & w7333) | (w1111 & w7333);
assign w3538 = ~w2613 & ~w321;
assign w3539 = w6186 & w2225;
assign w3540 = (w3057 & w2920) | (w3057 & w1553) | (w2920 & w1553);
assign w3541 = (w5655 & w2208) | (w5655 & w1625) | (w2208 & w1625);
assign w3542 = (~w1304 & w2340) | (~w1304 & w4504) | (w2340 & w4504);
assign w3543 = w5827 & w2899;
assign w3544 = (w1903 & w4518) | (w1903 & w7061) | (w4518 & w7061);
assign w3545 = (~w4143 & w7478) | (~w4143 & w2604) | (w7478 & w2604);
assign w3546 = w2011 & ~w2179;
assign w3547 = ~w6222 & ~w4612;
assign w3548 = ~w6375 & w5432;
assign w3549 = w2793 & ~w7454;
assign w3550 = (~w761 & w1306) | (~w761 & w6685) | (w1306 & w6685);
assign w3551 = a217 & b217;
assign w3552 = w6714 & w3614;
assign w3553 = ~w4028 & w4941;
assign w3554 = ~w5370 & w615;
assign w3555 = (~w6046 & w1773) | (~w6046 & w2166) | (w1773 & w2166);
assign w3556 = ~w7044 & w3903;
assign w3557 = ~w5066 & ~w3122;
assign w3558 = ~w4848 & w2765;
assign w3559 = (~w5655 & w2282) | (~w5655 & w3477) | (w2282 & w3477);
assign w3560 = (~w2871 & w3360) | (~w2871 & w571) | (w3360 & w571);
assign w3561 = ~w990 & ~w4149;
assign w3562 = (~w5257 & w6021) | (~w5257 & w6855) | (w6021 & w6855);
assign w3563 = (w6887 & w4398) | (w6887 & ~w5674) | (w4398 & ~w5674);
assign w3564 = (~w1936 & w1612) | (~w1936 & w5700) | (w1612 & w5700);
assign w3565 = (~w2456 & w961) | (~w2456 & w383) | (w961 & w383);
assign w3566 = (w918 & w387) | (w918 & ~w1730) | (w387 & ~w1730);
assign w3567 = ~w5820 & ~w4822;
assign w3568 = w161 & w7414;
assign w3569 = w1447 & ~w3873;
assign w3570 = ~w4765 & ~w5883;
assign w3571 = w2420 & w5297;
assign w3572 = w6450 & ~w1071;
assign w3573 = ~w1441 & ~w6683;
assign w3574 = (~w7391 & ~w4392) | (~w7391 & w5482) | (~w4392 & w5482);
assign w3575 = w701 & ~w206;
assign w3576 = (w4143 & w5880) | (w4143 & w854) | (w5880 & w854);
assign w3577 = (w7542 & w549) | (w7542 & w5291) | (w549 & w5291);
assign w3578 = ~w2957 & ~w4854;
assign w3579 = w3134 & ~w6017;
assign w3580 = a243 & b243;
assign w3581 = (w4732 & w1962) | (w4732 & ~w2013) | (w1962 & ~w2013);
assign w3582 = w7575 & ~w2401;
assign w3583 = (w6904 & w2232) | (w6904 & w1881) | (w2232 & w1881);
assign w3584 = ~w1071 & ~w558;
assign w3585 = ~w5958 & ~w1709;
assign w3586 = w6681 & ~w1628;
assign w3587 = a219 & b219;
assign w3588 = (w3636 & w5541) | (w3636 & w4223) | (w5541 & w4223);
assign w3589 = (w518 & w1611) | (w518 & w1768) | (w1611 & w1768);
assign w3590 = (w2935 & w2865) | (w2935 & ~w1791) | (w2865 & ~w1791);
assign w3591 = w728 & ~w4643;
assign w3592 = (~w7322 & w6762) | (~w7322 & w6136) | (w6762 & w6136);
assign w3593 = w3880 & w1231;
assign w3594 = (~w4327 & w2438) | (~w4327 & w6653) | (w2438 & w6653);
assign w3595 = w516 & w5581;
assign w3596 = ~w5871 & ~w189;
assign w3597 = (~w1367 & w2310) | (~w1367 & w494) | (w2310 & w494);
assign w3598 = (~w3741 & w1077) | (~w3741 & w6660) | (w1077 & w6660);
assign w3599 = w2471 & w36;
assign w3600 = w6415 & ~w2420;
assign w3601 = (~w6 & w4040) | (~w6 & w119) | (w4040 & w119);
assign w3602 = a3 & b3;
assign w3603 = (~w6945 & w4576) | (~w6945 & w481) | (w4576 & w481);
assign w3604 = ~w4911 & w744;
assign w3605 = w1937 & ~w2641;
assign w3606 = (w5000 & w393) | (w5000 & w5655) | (w393 & w5655);
assign w3607 = a11 & b11;
assign w3608 = w990 & w6195;
assign w3609 = (w681 & w2401) | (w681 & w5254) | (w2401 & w5254);
assign w3610 = (w4675 & w4610) | (w4675 & w3201) | (w4610 & w3201);
assign w3611 = (~w5257 & w1584) | (~w5257 & w3976) | (w1584 & w3976);
assign w3612 = ~w234 & ~w2379;
assign w3613 = w2796 & ~w7554;
assign w3614 = (w343 & w875) | (w343 & w4787) | (w875 & w4787);
assign w3615 = w1877 & w2483;
assign w3616 = a34 & b34;
assign w3617 = (w7205 & w3187) | (w7205 & w1139) | (w3187 & w1139);
assign w3618 = a167 & b167;
assign w3619 = w6994 & ~w3471;
assign w3620 = (w5581 & w3595) | (w5581 & w2011) | (w3595 & w2011);
assign w3621 = w2001 & ~w2954;
assign w3622 = (~w6162 & w4848) | (~w6162 & w6097) | (w4848 & w6097);
assign w3623 = (w7187 & w6798) | (w7187 & w553) | (w6798 & w553);
assign w3624 = (~w6353 & w2434) | (~w6353 & w3622) | (w2434 & w3622);
assign w3625 = ~w3152 & w7348;
assign w3626 = (~w6467 & w3761) | (~w6467 & w6867) | (w3761 & w6867);
assign w3627 = ~w3174 & ~w630;
assign w3628 = w3110 & ~w5403;
assign w3629 = ~w7471 & ~w2500;
assign w3630 = w5348 & ~w7000;
assign w3631 = ~w4987 & ~w5525;
assign w3632 = w2988 & w144;
assign w3633 = (~w5106 & w4716) | (~w5106 & w2221) | (w4716 & w2221);
assign w3634 = ~w5122 & w1169;
assign w3635 = (w5045 & w3245) | (w5045 & w6894) | (w3245 & w6894);
assign w3636 = w3399 & ~w4480;
assign w3637 = (w3636 & w1183) | (w3636 & w1724) | (w1183 & w1724);
assign w3638 = (w5173 & w3562) | (w5173 & ~w6100) | (w3562 & ~w6100);
assign w3639 = (w1611 & w2427) | (w1611 & w5387) | (w2427 & w5387);
assign w3640 = ~w2021 & w4;
assign w3641 = (~w5419 & w1807) | (~w5419 & w1666) | (w1807 & w1666);
assign w3642 = w2229 & ~w6714;
assign w3643 = ~w5599 & ~w4179;
assign w3644 = ~w5883 & ~w5923;
assign w3645 = ~w5827 & w5835;
assign w3646 = ~w1550 & w7012;
assign w3647 = ~w3384 & ~w2945;
assign w3648 = ~w3731 & w2188;
assign w3649 = (~w343 & w7588) | (~w343 & w3889) | (w7588 & w3889);
assign w3650 = (w4327 & w5567) | (w4327 & w2472) | (w5567 & w2472);
assign w3651 = (w1074 & w5840) | (w1074 & ~w173) | (w5840 & ~w173);
assign w3652 = (w5178 & w5318) | (w5178 & w6651) | (w5318 & w6651);
assign w3653 = w1455 & w5801;
assign w3654 = w6849 & ~w6709;
assign w3655 = ~w2818 & w101;
assign w3656 = ~w5999 & ~w869;
assign w3657 = ~w2409 & w3302;
assign w3658 = (w2515 & ~w913) | (w2515 & ~w924) | (~w913 & ~w924);
assign w3659 = ~w4034 & ~w74;
assign w3660 = ~w4402 & ~w706;
assign w3661 = ~w488 & w7608;
assign w3662 = w5348 & ~w5813;
assign w3663 = (~w5178 & w7253) | (~w5178 & w4774) | (w7253 & w4774);
assign w3664 = ~w4803 & w6857;
assign w3665 = ~a22 & ~b22;
assign w3666 = ~w6002 & w6122;
assign w3667 = (~w7187 & w4958) | (~w7187 & w1110) | (w4958 & w1110);
assign w3668 = (~w1420 & w2050) | (~w1420 & w6100) | (w2050 & w6100);
assign w3669 = a55 & b55;
assign w3670 = ~w3429 & ~w6232;
assign w3671 = ~w4082 & ~w5568;
assign w3672 = ~w504 & w3458;
assign w3673 = (~w3947 & w3687) | (~w3947 & w5502) | (w3687 & w5502);
assign w3674 = (w2570 & w7179) | (w2570 & ~w1383) | (w7179 & ~w1383);
assign w3675 = ~w5044 & ~w7428;
assign w3676 = (~w1143 & w2069) | (~w1143 & w3819) | (w2069 & w3819);
assign w3677 = ~w3014 & ~w6609;
assign w3678 = (w922 & w5067) | (w922 & w5403) | (w5067 & w5403);
assign w3679 = (~w812 & w1200) | (~w812 & w5582) | (w1200 & w5582);
assign w3680 = (~w4143 & w6780) | (~w4143 & w1351) | (w6780 & w1351);
assign w3681 = w3444 & ~w5217;
assign w3682 = ~a162 & ~b162;
assign w3683 = (~w1427 & w3078) | (~w1427 & w3939) | (w3078 & w3939);
assign w3684 = (~w6254 & ~w6966) | (~w6254 & w4355) | (~w6966 & w4355);
assign w3685 = (w3119 & w524) | (w3119 & w7004) | (w524 & w7004);
assign w3686 = w3905 & w3040;
assign w3687 = (w3647 & w4897) | (w3647 & ~w5368) | (w4897 & ~w5368);
assign w3688 = (w5059 & w352) | (w5059 & ~w2021) | (w352 & ~w2021);
assign w3689 = a227 & b227;
assign w3690 = ~w7350 & ~w5054;
assign w3691 = ~cin & ~w6548;
assign w3692 = ~a138 & ~b138;
assign w3693 = ~w1718 & ~w2892;
assign w3694 = (~w3805 & w5491) | (~w3805 & w6277) | (w5491 & w6277);
assign w3695 = (~w5655 & w4916) | (~w5655 & w4546) | (w4916 & w4546);
assign w3696 = w3835 & w6553;
assign w3697 = (w686 & w7601) | (w686 & w3381) | (w7601 & w3381);
assign w3698 = (~w5257 & w5075) | (~w5257 & w637) | (w5075 & w637);
assign w3699 = (~w7510 & w4923) | (~w7510 & w3679) | (w4923 & w3679);
assign w3700 = (w2686 & w321) | (w2686 & w933) | (w321 & w933);
assign w3701 = ~w2872 & ~w247;
assign w3702 = w3507 & ~w3619;
assign w3703 = ~w5803 | ~w5568;
assign w3704 = w2838 & w385;
assign w3705 = (~w550 & w5893) | (~w550 & w5536) | (w5893 & w5536);
assign w3706 = ~w7648 & w4422;
assign w3707 = ~w453 & w7392;
assign w3708 = w139 & w2420;
assign w3709 = (w3062 & w314) | (w3062 & w1354) | (w314 & w1354);
assign w3710 = w6503 & ~w5658;
assign w3711 = ~w7076 & ~w1357;
assign w3712 = a224 & b224;
assign w3713 = ~w1723 & ~w3437;
assign w3714 = ~w1761 & ~w3715;
assign w3715 = (w5655 & w4051) | (w5655 & w2320) | (w4051 & w2320);
assign w3716 = ~w4616 & ~w3418;
assign w3717 = w4167 & ~w2453;
assign w3718 = (w2985 & w6496) | (w2985 & w2723) | (w6496 & w2723);
assign w3719 = ~w102 & w814;
assign w3720 = ~w5416 & w3362;
assign w3721 = (w5834 & w6020) | (w5834 & w6629) | (w6020 & w6629);
assign w3722 = ~w1805 & ~w7484;
assign w3723 = ~w3057 & w1815;
assign w3724 = (~w3455 & w6564) | (~w3455 & w432) | (w6564 & w432);
assign w3725 = (w3866 & w2089) | (w3866 & w2523) | (w2089 & w2523);
assign w3726 = w2486 & ~w7214;
assign w3727 = (~w1158 & w6299) | (~w1158 & w3202) | (w6299 & w3202);
assign w3728 = ~w6630 & w434;
assign w3729 = ~w2515 & w6754;
assign w3730 = ~w3909 & w4333;
assign w3731 = ~w6760 & ~w2997;
assign w3732 = ~a221 & ~b221;
assign w3733 = w4305 & w6203;
assign w3734 = (~w7391 & ~w4392) | (~w7391 & w6682) | (~w4392 & w6682);
assign w3735 = ~a192 & ~b192;
assign w3736 = ~w4 & w6718;
assign w3737 = ~w2997 & w6112;
assign w3738 = (w5178 & w1540) | (w5178 & w4736) | (w1540 & w4736);
assign w3739 = w2112 & ~w4090;
assign w3740 = (w7145 & w4446) | (w7145 & ~w5291) | (w4446 & ~w5291);
assign w3741 = ~w6444 & ~w143;
assign w3742 = ~w6450 & w4827;
assign w3743 = w5385 & w6894;
assign w3744 = (~w5672 & w7606) | (~w5672 & w5440) | (w7606 & w5440);
assign w3745 = ~w13 & ~w3692;
assign w3746 = ~w1196 & w2243;
assign w3747 = (w6246 & w1044) | (w6246 & w6580) | (w1044 & w6580);
assign w3748 = w1501 & ~w1722;
assign w3749 = ~w2271 & w5368;
assign w3750 = (~w777 & w976) | (~w777 & w4349) | (w976 & w4349);
assign w3751 = ~w2441 & w51;
assign w3752 = w3840 & w6789;
assign w3753 = (w5178 & w3678) | (w5178 & w7636) | (w3678 & w7636);
assign w3754 = ~w6138 & ~w908;
assign w3755 = (w7273 & w5901) | (w7273 & w1255) | (w5901 & w1255);
assign w3756 = w1057 & ~w6766;
assign w3757 = (w6359 & w1453) | (w6359 & w1892) | (w1453 & w1892);
assign w3758 = ~w2465 & ~w4035;
assign w3759 = (w7145 & w4446) | (w7145 & ~w563) | (w4446 & ~w563);
assign w3760 = (~w1925 & w1731) | (~w1925 & w206) | (w1731 & w206);
assign w3761 = (w7199 & w1171) | (w7199 & w5542) | (w1171 & w5542);
assign w3762 = w6683 & w1283;
assign w3763 = (w7529 & w1659) | (w7529 & ~w1886) | (w1659 & ~w1886);
assign w3764 = (~w5178 & w1335) | (~w5178 & w178) | (w1335 & w178);
assign w3765 = w1741 & w7625;
assign w3766 = w1053 & w7489;
assign w3767 = w2688 & w7332;
assign w3768 = w4812 | ~w6184;
assign w3769 = (w5703 & w2446) | (w5703 & w7434) | (w2446 & w7434);
assign w3770 = (~w4468 & w6230) | (~w4468 & w6028) | (w6230 & w6028);
assign w3771 = w195 & ~w698;
assign w3772 = w1560 & w3004;
assign w3773 = ~w7475 & ~w864;
assign w3774 = (~w4494 & ~w6353) | (~w4494 & w2345) | (~w6353 & w2345);
assign w3775 = ~w7190 & ~w3017;
assign w3776 = w1321 & w6637;
assign w3777 = (w2169 & w6379) | (w2169 & ~w3883) | (w6379 & ~w3883);
assign w3778 = (w4385 & w1918) | (w4385 & ~w6174) | (w1918 & ~w6174);
assign w3779 = (w1332 & w5814) | (w1332 & ~w632) | (w5814 & ~w632);
assign w3780 = w3523 & ~w2876;
assign w3781 = w331 & w3914;
assign w3782 = a46 & b46;
assign w3783 = ~w652 | w4757;
assign w3784 = ~w6844 & w7165;
assign w3785 = (w6649 & w6532) | (w6649 & ~w2482) | (w6532 & ~w2482);
assign w3786 = w6872 & w5212;
assign w3787 = w2119 & w3427;
assign w3788 = (w5427 & w6896) | (w5427 & w6328) | (w6896 & w6328);
assign w3789 = (w5237 & w3257) | (w5237 & w6294) | (w3257 & w6294);
assign w3790 = (~w236 & w3340) | (~w236 & w5716) | (w3340 & w5716);
assign w3791 = w2915 | w4604;
assign w3792 = (w5257 & w5784) | (w5257 & w2638) | (w5784 & w2638);
assign w3793 = (w2721 & w6686) | (w2721 & ~w6566) | (w6686 & ~w6566);
assign w3794 = (w6106 & w1909) | (w6106 & w1401) | (w1909 & w1401);
assign w3795 = ~w7027 & ~w1628;
assign w3796 = w3111 & w1742;
assign w3797 = w99 & w4989;
assign w3798 = w1457 & ~w1143;
assign w3799 = a110 & b110;
assign w3800 = w4036 & w5979;
assign w3801 = (w7386 & ~w2021) | (w7386 & w4655) | (~w2021 & w4655);
assign w3802 = ~w3888 & w2426;
assign w3803 = (w5178 & w2412) | (w5178 & w4229) | (w2412 & w4229);
assign w3804 = w5860 & ~w6848;
assign w3805 = w6353 & w979;
assign w3806 = (w2065 & w4668) | (w2065 & w7595) | (w4668 & w7595);
assign w3807 = w5484 & w820;
assign w3808 = ~w5901 & w1438;
assign w3809 = (~w6100 & w2719) | (~w6100 & w5227) | (w2719 & w5227);
assign w3810 = (~w5325 & ~w1892) | (~w5325 & ~w3743) | (~w1892 & ~w3743);
assign w3811 = (~w7530 & w6705) | (~w7530 & w3914) | (w6705 & w3914);
assign w3812 = (~w7292 & ~w4182) | (~w7292 & ~w1315) | (~w4182 & ~w1315);
assign w3813 = w2 & ~w6712;
assign w3814 = (w5430 & w2538) | (w5430 & w4085) | (w2538 & w4085);
assign w3815 = w3677 & w5161;
assign w3816 = (~w5178 & w3184) | (~w5178 & w5434) | (w3184 & w5434);
assign w3817 = w1827 & ~w3869;
assign w3818 = w6718 & w5929;
assign w3819 = ~w2708 & w1930;
assign w3820 = (~w3952 & w532) | (~w3952 & w6828) | (w532 & w6828);
assign w3821 = ~w3782 & ~w1471;
assign w3822 = ~w2831 & ~w4949;
assign w3823 = ~w3064 & w5914;
assign w3824 = (w6353 & w3886) | (w6353 & w1982) | (w3886 & w1982);
assign w3825 = ~w791 & ~w5613;
assign w3826 = w5333 & ~w3195;
assign w3827 = (w1518 & w5340) | (w1518 & w1985) | (w5340 & w1985);
assign w3828 = ~w3677 & w1463;
assign w3829 = (w2935 & w2865) | (w2935 & w7444) | (w2865 & w7444);
assign w3830 = (~w4898 & w4323) | (~w4898 & w6599) | (w4323 & w6599);
assign w3831 = w5721 & w5996;
assign w3832 = ~w1153 | w505;
assign w3833 = (~w3318 & w5786) | (~w3318 & w3766) | (w5786 & w3766);
assign w3834 = (~w3210 & w4611) | (~w3210 & ~w6757) | (w4611 & ~w6757);
assign w3835 = ~w5230 & w1131;
assign w3836 = w3665 & ~w5864;
assign w3837 = ~w1568 & ~w5874;
assign w3838 = (~w7648 & w3771) | (~w7648 & w3285) | (w3771 & w3285);
assign w3839 = (w568 & w6943) | (w568 & w7124) | (w6943 & w7124);
assign w3840 = ~w4759 & ~w426;
assign w3841 = ~w2838 & w7352;
assign w3842 = ~w7012 & ~w1550;
assign w3843 = w6386 & w3997;
assign w3844 = (~w7118 & w282) | (~w7118 & w5063) | (w282 & w5063);
assign w3845 = (w5178 & w2414) | (w5178 & w3069) | (w2414 & w3069);
assign w3846 = (w5257 & w6493) | (w5257 & w4516) | (w6493 & w4516);
assign w3847 = (~w4995 & w3165) | (~w4995 & w6362) | (w3165 & w6362);
assign w3848 = (w577 & w3838) | (w577 & w3872) | (w3838 & w3872);
assign w3849 = (w1155 & w2510) | (w1155 & ~w3074) | (w2510 & ~w3074);
assign w3850 = ~w1935 & ~w293;
assign w3851 = ~w5348 & w5813;
assign w3852 = (w1987 & w6081) | (w1987 & w3074) | (w6081 & w3074);
assign w3853 = ~w127 & ~w3243;
assign w3854 = w3836 & ~w3166;
assign w3855 = a187 & b187;
assign w3856 = w2542 & w6100;
assign w3857 = w3119 & w5779;
assign w3858 = (w3061 & ~w1751) | (w3061 & w3441) | (~w1751 & w3441);
assign w3859 = (w5511 & w7252) | (w5511 & w5208) | (w7252 & w5208);
assign w3860 = w4923 & ~w7510;
assign w3861 = (w4337 & w6604) | (w4337 & w5955) | (w6604 & w5955);
assign w3862 = (~w4169 & w5594) | (~w4169 & w2027) | (w5594 & w2027);
assign w3863 = ~w4165 & ~w5616;
assign w3864 = ~w3802 & w6891;
assign w3865 = ~w6990 & ~w6989;
assign w3866 = ~w5428 & w1574;
assign w3867 = (~w2335 & w5596) | (~w2335 & w4049) | (w5596 & w4049);
assign w3868 = ~w4911 & ~w7044;
assign w3869 = ~a250 & ~b250;
assign w3870 = (~w3983 & w470) | (~w3983 & w4846) | (w470 & w4846);
assign w3871 = ~w4681 & w3264;
assign w3872 = w1632 & w577;
assign w3873 = ~w1303 & w7152;
assign w3874 = (w5181 & w2370) | (w5181 & w7494) | (w2370 & w7494);
assign w3875 = (w4812 & w5331) | (w4812 & ~w5871) | (w5331 & ~w5871);
assign w3876 = ~w1544 & ~w4780;
assign w3877 = ~w105 & ~w3222;
assign w3878 = w5594 | ~w4169;
assign w3879 = (w5257 & w3413) | (w5257 & w413) | (w3413 & w413);
assign w3880 = (~w3262 & w3055) | (~w3262 & w1960) | (w3055 & w1960);
assign w3881 = (w5178 & w1853) | (w5178 & w227) | (w1853 & w227);
assign w3882 = (~w7372 & w5634) | (~w7372 & w2606) | (w5634 & w2606);
assign w3883 = ~w5391 & w6751;
assign w3884 = w139 & w861;
assign w3885 = (~w3063 & w5711) | (~w3063 & w1838) | (w5711 & w1838);
assign w3886 = ~w13 & ~w5627;
assign w3887 = ~a254 & ~b254;
assign w3888 = ~w2229 & w7201;
assign w3889 = ~w4706 & ~w3647;
assign w3890 = (w5257 & w5924) | (w5257 & w2616) | (w5924 & w2616);
assign w3891 = (w4604 & w1598) | (w4604 & w3791) | (w1598 & w3791);
assign w3892 = w5058 & w4459;
assign w3893 = ~a30 & ~b30;
assign w3894 = ~w4337 & w1297;
assign w3895 = (~w2693 & w5347) | (~w2693 & w4431) | (w5347 & w4431);
assign w3896 = a123 & b123;
assign w3897 = (w185 & w6249) | (w185 & w4270) | (w6249 & w4270);
assign w3898 = (w3427 & w7600) | (w3427 & ~w3247) | (w7600 & ~w3247);
assign w3899 = ~w6233 & w6281;
assign w3900 = ~w4484 & ~w574;
assign w3901 = ~w3158 & ~w76;
assign w3902 = (w6038 & w3973) | (w6038 & w5579) | (w3973 & w5579);
assign w3903 = ~w2725 & ~w3551;
assign w3904 = (~w6100 & w6288) | (~w6100 & w5704) | (w6288 & w5704);
assign w3905 = ~a25 & ~b25;
assign w3906 = ~w6507 & w839;
assign w3907 = ~w1709 & ~w2097;
assign w3908 = (w6082 & w3379) | (w6082 & w1887) | (w3379 & w1887);
assign w3909 = ~a46 & ~b46;
assign w3910 = (w5441 & w5805) | (w5441 & ~w6254) | (w5805 & ~w6254);
assign w3911 = ~w7614 & w2663;
assign w3912 = w7187 & w3808;
assign w3913 = w3007 & ~w1661;
assign w3914 = ~w6439 & w60;
assign w3915 = w4706 & ~w2945;
assign w3916 = w1877 & ~w1575;
assign w3917 = w4988 & ~w5034;
assign w3918 = ~a167 & ~b167;
assign w3919 = (~w5178 & w5592) | (~w5178 & w1236) | (w5592 & w1236);
assign w3920 = (~w6127 & w1763) | (~w6127 & w4245) | (w1763 & w4245);
assign w3921 = (w342 & w7013) | (w342 & w3576) | (w7013 & w3576);
assign w3922 = ~w6709 & ~w2563;
assign w3923 = w2047 & w5030;
assign w3924 = ~w4786 & w1630;
assign w3925 = (w410 & w5167) | (w410 & ~w6174) | (w5167 & ~w6174);
assign w3926 = (w3737 & w7160) | (w3737 & w2128) | (w7160 & w2128);
assign w3927 = ~w3573 & ~w47;
assign w3928 = (~w5178 & w6605) | (~w5178 & w4153) | (w6605 & w4153);
assign w3929 = w6927 & ~w3868;
assign w3930 = (w3381 & w3697) | (w3381 & w6100) | (w3697 & w6100);
assign w3931 = w2110 | ~w693;
assign w3932 = ~a227 & ~b227;
assign w3933 = ~w6757 & ~w1216;
assign w3934 = ~a204 & ~b204;
assign w3935 = w1304 & w3076;
assign w3936 = (~w3947 & w343) | (~w3947 & w4929) | (w343 & w4929);
assign w3937 = w1821 & ~w3435;
assign w3938 = (w7453 & w6732) | (w7453 & w4369) | (w6732 & w4369);
assign w3939 = (~w1427 & w4337) | (~w1427 & w5504) | (w4337 & w5504);
assign w3940 = w3565 | w961;
assign w3941 = w767 & ~w2966;
assign w3942 = (w5230 & ~w5560) | (w5230 & ~w7490) | (~w5560 & ~w7490);
assign w3943 = ~w3644 & w3467;
assign w3944 = (w5068 & w6918) | (w5068 & ~w7043) | (w6918 & ~w7043);
assign w3945 = w7002 & ~w463;
assign w3946 = w331 & ~w6439;
assign w3947 = w3774 & w2557;
assign w3948 = ~w1813 & ~w7421;
assign w3949 = ~w1002 & ~w5600;
assign w3950 = (~w5178 & w5164) | (~w5178 & w1904) | (w5164 & w1904);
assign w3951 = ~w3266 & ~w273;
assign w3952 = (w632 & w5007) | (w632 & w7124) | (w5007 & w7124);
assign w3953 = (~w4995 & w5602) | (~w4995 & w6610) | (w5602 & w6610);
assign w3954 = (w5559 & w2900) | (w5559 & ~w6798) | (w2900 & ~w6798);
assign w3955 = ~w3933 & w6981;
assign w3956 = ~w2408 & w2236;
assign w3957 = w2735 & ~w5478;
assign w3958 = ~w4002 & ~w6426;
assign w3959 = (~w1656 & w731) | (~w1656 & w5645) | (w731 & w5645);
assign w3960 = ~w2100 & ~w4553;
assign w3961 = (w5178 & w3149) | (w5178 & w4133) | (w3149 & w4133);
assign w3962 = w628 & ~w632;
assign w3963 = w878 & ~w3033;
assign w3964 = (w7529 & w1659) | (w7529 & w7450) | (w1659 & w7450);
assign w3965 = a215 & b215;
assign w3966 = (w2429 & w5142) | (w2429 & w4472) | (w5142 & w4472);
assign w3967 = w5404 & ~w7647;
assign w3968 = ~w1570 & ~w2432;
assign w3969 = w4905 & w6214;
assign w3970 = (~w4884 & w783) | (~w4884 & w6356) | (w783 & w6356);
assign w3971 = w3129 & ~w4074;
assign w3972 = w1080 & w4121;
assign w3973 = w6125 & w7187;
assign w3974 = ~w3007 & ~w841;
assign w3975 = (w3057 & w4542) | (w3057 & w5591) | (w4542 & w5591);
assign w3976 = (w3431 & w929) | (w3431 & ~w3391) | (w929 & ~w3391);
assign w3977 = (w1692 & w1262) | (w1692 & ~w6894) | (w1262 & ~w6894);
assign w3978 = (~w777 & w6116) | (~w777 & w5638) | (w6116 & w5638);
assign w3979 = (~w5672 & w3456) | (~w5672 & w3707) | (w3456 & w3707);
assign w3980 = w4681 & ~w2503;
assign w3981 = ~w6706 & w6257;
assign w3982 = w3004 & ~w7304;
assign w3983 = (w1987 & w6081) | (w1987 & w7383) | (w6081 & w7383);
assign w3984 = (~w1431 & w6705) | (~w1431 & w3411) | (w6705 & w3411);
assign w3985 = ~w2515 & ~w7429;
assign w3986 = (w6633 & ~w3819) | (w6633 & w236) | (~w3819 & w236);
assign w3987 = w386 & w7630;
assign w3988 = (w6424 & w55) | (w6424 & w7217) | (w55 & w7217);
assign w3989 = ~w7292 & w1743;
assign w3990 = a98 & b98;
assign w3991 = (~w5178 & w5632) | (~w5178 & w6090) | (w5632 & w6090);
assign w3992 = (~w5834 & w2999) | (~w5834 & w7086) | (w2999 & w7086);
assign w3993 = w2630 & ~w5397;
assign w3994 = ~w6890 & w3481;
assign w3995 = ~w6757 & ~w1999;
assign w3996 = (~w5196 & w722) | (~w5196 & w3153) | (w722 & w3153);
assign w3997 = a201 & b201;
assign w3998 = ~w1833 & ~w1004;
assign w3999 = ~w6660 & w2540;
assign w4000 = ~w973 & w6301;
assign w4001 = ~w2724 & ~w1345;
assign w4002 = ~w3252 & ~w7384;
assign w4003 = (~w335 & w3256) | (~w335 & w2629) | (w3256 & w2629);
assign w4004 = a147 & b147;
assign w4005 = (~w7205 & w5780) | (~w7205 & w2924) | (w5780 & w2924);
assign w4006 = (w1367 & w17) | (w1367 & w1299) | (w17 & w1299);
assign w4007 = ~w5965 & w243;
assign w4008 = w4069 & w6894;
assign w4009 = (w1611 & w3378) | (w1611 & w3388) | (w3378 & w3388);
assign w4010 = a165 & b165;
assign w4011 = ~w5402 & w1859;
assign w4012 = ~w5170 & ~w4412;
assign w4013 = (w6126 & w5155) | (w6126 & w3391) | (w5155 & w3391);
assign w4014 = ~w5277 & ~w2862;
assign w4015 = w4871 & w445;
assign w4016 = ~w5474 & ~w6790;
assign w4017 = (w5752 & ~w7610) | (w5752 & w1840) | (~w7610 & w1840);
assign w4018 = (w5178 & w566) | (w5178 & w5137) | (w566 & w5137);
assign w4019 = ~w4142 | w728;
assign w4020 = w5462 | w4926;
assign w4021 = (~w736 & ~w1356) | (~w736 & w2759) | (~w1356 & w2759);
assign w4022 = w1260 & ~w783;
assign w4023 = (w6100 & w312) | (w6100 & w1902) | (w312 & w1902);
assign w4024 = (~w5672 & w711) | (~w5672 & w5401) | (w711 & w5401);
assign w4025 = w3064 & ~w5914;
assign w4026 = (w5415 & ~w6100) | (w5415 & w6188) | (~w6100 & w6188);
assign w4027 = ~w7424 & ~w6810;
assign w4028 = w2572 & ~w5696;
assign w4029 = ~w7332 & ~w3819;
assign w4030 = ~w1655 & ~w7302;
assign w4031 = (w4323 & w2950) | (w4323 & ~w2097) | (w2950 & ~w2097);
assign w4032 = (w3083 & w5597) | (w3083 & w5718) | (w5597 & w5718);
assign w4033 = ~w145 & w2558;
assign w4034 = (~w5834 & w2184) | (~w5834 & w6932) | (w2184 & w6932);
assign w4035 = a4 & b4;
assign w4036 = ~w4775 & ~w3072;
assign w4037 = (w4036 & w3597) | (w4036 & w2881) | (w3597 & w2881);
assign w4038 = (w1493 & w2651) | (w1493 & w5574) | (w2651 & w5574);
assign w4039 = (w777 & w7487) | (w777 & w6440) | (w7487 & w6440);
assign w4040 = w456 & ~w7385;
assign w4041 = (w3774 & w5714) | (w3774 & w3969) | (w5714 & w3969);
assign w4042 = (w6467 & w4785) | (w6467 & w3620) | (w4785 & w3620);
assign w4043 = ~w486 & w3471;
assign w4044 = ~w4002 & w2077;
assign w4045 = ~w1083 & ~w4545;
assign w4046 = (~w6413 & w5520) | (~w6413 & w6982) | (w5520 & w6982);
assign w4047 = (w2004 & w1539) | (w2004 & w5655) | (w1539 & w5655);
assign w4048 = w3677 & w7473;
assign w4049 = ~w3631 & ~w3998;
assign w4050 = ~w931 & w5655;
assign w4051 = (~w5257 & w1684) | (~w5257 & w7130) | (w1684 & w7130);
assign w4052 = (w783 & w956) | (w783 & w605) | (w956 & w605);
assign w4053 = w5435 & w6174;
assign w4054 = (w5262 & w556) | (w5262 & w3131) | (w556 & w3131);
assign w4055 = (~w6738 & w1415) | (~w6738 & w4583) | (w1415 & w4583);
assign w4056 = (w6541 & w1670) | (w6541 & w7238) | (w1670 & w7238);
assign w4057 = ~w2127 & w7538;
assign w4058 = (w412 & w7602) | (w412 & w6821) | (w7602 & w6821);
assign w4059 = ~w3083 & w6679;
assign w4060 = ~a78 & ~b78;
assign w4061 = ~w5118 & ~w1389;
assign w4062 = (w136 & w842) | (w136 & ~w563) | (w842 & ~w563);
assign w4063 = ~w4731 & ~w2053;
assign w4064 = ~w6935 & ~w3985;
assign w4065 = ~w4976 & ~w2343;
assign w4066 = ~w7042 & ~w1848;
assign w4067 = w7114 & ~w3272;
assign w4068 = ~w5229 & ~w2027;
assign w4069 = (~w7626 & w3704) | (~w7626 & w6808) | (w3704 & w6808);
assign w4070 = ~w2158 & ~w7135;
assign w4071 = (~w3947 & w7389) | (~w3947 & w5129) | (w7389 & w5129);
assign w4072 = ~w7345 & w2513;
assign w4073 = ~w6082 & w2400;
assign w4074 = w3587 & ~w2104;
assign w4075 = (~w4680 & w199) | (~w4680 & w1787) | (w199 & w1787);
assign w4076 = (w1190 & w3556) | (w1190 & ~w3396) | (w3556 & ~w3396);
assign w4077 = w5370 & ~w1472;
assign w4078 = (w4967 & w4796) | (w4967 & w1407) | (w4796 & w1407);
assign w4079 = w7296 & w6357;
assign w4080 = ~w2127 & w7521;
assign w4081 = w1594 & ~w2818;
assign w4082 = ~w5622 & ~w1471;
assign w4083 = ~w1913 & w2786;
assign w4084 = ~w2283 & ~w5276;
assign w4085 = (~w1804 & w238) | (~w1804 & w6566) | (w238 & w6566);
assign w4086 = (~w1328 & w3549) | (~w1328 & w4319) | (w3549 & w4319);
assign w4087 = w6354 & w3480;
assign w4088 = w2024 & ~w1137;
assign w4089 = (~w2409 & w5384) | (~w2409 & w1267) | (w5384 & w1267);
assign w4090 = ~w3122 & ~w5241;
assign w4091 = (w4889 & w4372) | (w4889 & w6733) | (w4372 & w6733);
assign w4092 = ~w5830 & w6219;
assign w4093 = (~w6387 & w4771) | (~w6387 & w4) | (w4771 & w4);
assign w4094 = ~w2112 & w4090;
assign w4095 = (w681 & w1100) | (w681 & w3266) | (w1100 & w3266);
assign w4096 = w5823 | w3434;
assign w4097 = (w3060 & w1296) | (w3060 & ~w5403) | (w1296 & ~w5403);
assign w4098 = w2965 & w1531;
assign w4099 = ~w4415 & w5781;
assign w4100 = (w3892 & w7496) | (w3892 & w6838) | (w7496 & w6838);
assign w4101 = ~w7216 & w3215;
assign w4102 = ~w6265 & w3397;
assign w4103 = (~w1655 & ~w7302) | (~w1655 & w1919) | (~w7302 & w1919);
assign w4104 = (w632 & w5007) | (w632 & w2097) | (w5007 & w2097);
assign w4105 = ~w3033 & w5781;
assign w4106 = (~w7363 & w2558) | (~w7363 & w7) | (w2558 & w7);
assign w4107 = ~a111 & ~b111;
assign w4108 = (w1163 & w2677) | (w1163 & ~w5395) | (w2677 & ~w5395);
assign w4109 = w4398 | w6887;
assign w4110 = w5433 & ~w3062;
assign w4111 = ~w5082 & ~w3371;
assign w4112 = (w5879 & w5252) | (w5879 & w7554) | (w5252 & w7554);
assign w4113 = (w900 & w7036) | (w900 & w6100) | (w7036 & w6100);
assign w4114 = (~w4940 & w1377) | (~w4940 & w3731) | (w1377 & w3731);
assign w4115 = w5248 & w3567;
assign w4116 = ~w2582 & w7354;
assign w4117 = (w76 & w7646) | (w76 & ~w4764) | (w7646 & ~w4764);
assign w4118 = w354 & w6174;
assign w4119 = w1799 & ~w3138;
assign w4120 = (w5702 & ~w5851) | (w5702 & ~w1892) | (~w5851 & ~w1892);
assign w4121 = (w384 & w7372) | (w384 & w5004) | (w7372 & w5004);
assign w4122 = (w3847 & w567) | (w3847 & w4819) | (w567 & w4819);
assign w4123 = a237 & b237;
assign w4124 = (~w7493 & w1660) | (~w7493 & w6367) | (w1660 & w6367);
assign w4125 = ~w6960 & ~w588;
assign w4126 = w272 & w6315;
assign w4127 = (~w761 & w1306) | (~w761 & w2641) | (w1306 & w2641);
assign w4128 = (w6257 & w3375) | (w6257 & w3981) | (w3375 & w3981);
assign w4129 = w188 & ~w7574;
assign w4130 = ~w3580 & w3474;
assign w4131 = (w3953 & w5991) | (w3953 & w6574) | (w5991 & w6574);
assign w4132 = w6492 & w5197;
assign w4133 = (~w6467 & w3149) | (~w6467 & w6618) | (w3149 & w6618);
assign w4134 = ~w4832 & ~w3237;
assign w4135 = w1176 & w3854;
assign w4136 = ~w6628 & ~w5442;
assign w4137 = (w544 & w5625) | (w544 & ~w5013) | (w5625 & ~w5013);
assign w4138 = ~w4143 & w1892;
assign w4139 = ~w6013 & ~w3913;
assign w4140 = ~a98 & ~b98;
assign w4141 = ~w686 & w1890;
assign w4142 = w2255 & ~w728;
assign w4143 = w3119 & ~w5403;
assign w4144 = (~w2513 & w6668) | (~w2513 & w2456) | (w6668 & w2456);
assign w4145 = w1991 & ~w7216;
assign w4146 = ~a223 & ~b223;
assign w4147 = ~w7384 & ~w687;
assign w4148 = a150 & b150;
assign w4149 = a72 & b72;
assign w4150 = (~w6716 & w1721) | (~w6716 & w441) | (w1721 & w441);
assign w4151 = (w7626 & w7518) | (w7626 & w986) | (w7518 & w986);
assign w4152 = (w1736 & w3224) | (w1736 & w5040) | (w3224 & w5040);
assign w4153 = (w702 & w1696) | (w702 & w3491) | (w1696 & w3491);
assign w4154 = (w5323 & w3713) | (w5323 & w739) | (w3713 & w739);
assign w4155 = (w426 & ~w587) | (w426 & w7391) | (~w587 & w7391);
assign w4156 = (~w6222 & ~w3173) | (~w6222 & w40) | (~w3173 & w40);
assign w4157 = (w3947 & w6098) | (w3947 & w2943) | (w6098 & w2943);
assign w4158 = (~w4710 & w7528) | (~w4710 & w3535) | (w7528 & w3535);
assign w4159 = (w4995 & w3742) | (w4995 & w4573) | (w3742 & w4573);
assign w4160 = (w5325 & w1855) | (w5325 & w4927) | (w1855 & w4927);
assign w4161 = ~w1386 & w3139;
assign w4162 = w1455 & w3585;
assign w4163 = w3328 & ~w6025;
assign w4164 = ~w5977 | w5760;
assign w4165 = ~a99 & ~b99;
assign w4166 = w5640 & ~w6612;
assign w4167 = ~w6272 & w5436;
assign w4168 = ~a11 & ~b11;
assign w4169 = ~a43 & ~b43;
assign w4170 = ~w6516 & ~w404;
assign w4171 = w5643 & ~w2717;
assign w4172 = (w4123 & ~w6614) | (w4123 & w1607) | (~w6614 & w1607);
assign w4173 = w1276 & w287;
assign w4174 = a29 & b29;
assign w4175 = w2255 & ~w3113;
assign w4176 = ~a152 & ~b152;
assign w4177 = (w7506 & ~w4284) | (w7506 & w1280) | (~w4284 & w1280);
assign w4178 = (~w2021 & w6318) | (~w2021 & w4093) | (w6318 & w4093);
assign w4179 = a251 & b251;
assign w4180 = (~w5958 & w4933) | (~w5958 & w5964) | (w4933 & w5964);
assign w4181 = (w1515 & w4320) | (w1515 & w5493) | (w4320 & w5493);
assign w4182 = (w7292 & w5402) | (w7292 & w4486) | (w5402 & w4486);
assign w4183 = ~w2221 & w2074;
assign w4184 = (~w3461 & w3860) | (~w3461 & w3699) | (w3860 & w3699);
assign w4185 = ~a196 & ~b196;
assign w4186 = w1091 & w6018;
assign w4187 = ~w5901 & w2221;
assign w4188 = w3514 & w868;
assign w4189 = (~w6878 & w6847) | (~w6878 & w2618) | (w6847 & w2618);
assign w4190 = (w7626 & w5336) | (w7626 & w7578) | (w5336 & w7578);
assign w4191 = ~w3691 & w4001;
assign w4192 = (~w858 & w73) | (~w858 & w3858) | (w73 & w3858);
assign w4193 = ~a147 & ~b147;
assign w4194 = (w4357 & w1240) | (w4357 & ~w4143) | (w1240 & ~w4143);
assign w4195 = w1607 & w5212;
assign w4196 = w348 & ~w1094;
assign w4197 = (w8 & w190) | (w8 & w7293) | (w190 & w7293);
assign w4198 = (~w4333 & w6648) | (~w4333 & w5341) | (w6648 & w5341);
assign w4199 = (w169 & w3168) | (w169 & w2770) | (w3168 & w2770);
assign w4200 = (~w1925 & w1731) | (~w1925 & ~w4940) | (w1731 & ~w4940);
assign w4201 = ~w2542 & w999;
assign w4202 = w7172 & w6974;
assign w4203 = ~w4898 & ~w5242;
assign w4204 = ~w2066 & w5059;
assign w4205 = w5107 & w4560;
assign w4206 = ~w7546 & ~w7390;
assign w4207 = ~w7522 & ~w1901;
assign w4208 = (~w1441 & ~w2108) | (~w1441 & w6161) | (~w2108 & w6161);
assign w4209 = (~w4265 & w2452) | (~w4265 & w2190) | (w2452 & w2190);
assign w4210 = (w401 & w5761) | (w401 & w3077) | (w5761 & w3077);
assign w4211 = w1073 & w4249;
assign w4212 = (w5834 & w1776) | (w5834 & w7164) | (w1776 & w7164);
assign w4213 = (w5522 & w4088) | (w5522 & w7534) | (w4088 & w7534);
assign w4214 = ~w4976 & ~w2408;
assign w4215 = w7111 & w5143;
assign w4216 = ~w4843 & w7574;
assign w4217 = (w5178 & w5919) | (w5178 & w1277) | (w5919 & w1277);
assign w4218 = w7181 & ~w382;
assign w4219 = (w6071 & w7141) | (w6071 & ~w3391) | (w7141 & ~w3391);
assign w4220 = ~w4811 & ~w4651;
assign w4221 = (w4628 & w7187) | (w4628 & w2589) | (w7187 & w2589);
assign w4222 = ~w6439 & ~w60;
assign w4223 = w6490 & w3538;
assign w4224 = ~w273 & w3515;
assign w4225 = (w5655 & w1592) | (w5655 & w4740) | (w1592 & w4740);
assign w4226 = w3363 & w4057;
assign w4227 = (~w6614 & w2958) | (~w6614 & w5326) | (w2958 & w5326);
assign w4228 = w5259 & w6469;
assign w4229 = (w5325 & w2679) | (w5325 & w4365) | (w2679 & w4365);
assign w4230 = ~w3192 & w6566;
assign w4231 = (~w7552 & w1042) | (~w7552 & w2950) | (w1042 & w2950);
assign w4232 = (~w6252 & w2872) | (~w6252 & w4617) | (w2872 & w4617);
assign w4233 = ~w2249 & ~w6512;
assign w4234 = w788 & w3349;
assign w4235 = w2778 | w1609;
assign w4236 = ~w2836 & ~w1165;
assign w4237 = ~w4321 & w2840;
assign w4238 = ~a58 & ~b58;
assign w4239 = w4958 & ~w7332;
assign w4240 = (w7095 & w572) | (w7095 & ~w5098) | (w572 & ~w5098);
assign w4241 = (~w3318 & w2461) | (~w3318 & w2138) | (w2461 & w2138);
assign w4242 = ~a96 & ~b96;
assign w4243 = w5761 & w401;
assign w4244 = (w3899 & w613) | (w3899 & ~w4199) | (w613 & ~w4199);
assign w4245 = ~w2471 & ~w6462;
assign w4246 = (~w2542 & w4201) | (~w2542 & w2327) | (w4201 & w2327);
assign w4247 = w4564 & ~w434;
assign w4248 = ~w3057 & w7551;
assign w4249 = (~w4409 & w4847) | (~w4409 & w5285) | (w4847 & w5285);
assign w4250 = ~w2603 & w318;
assign w4251 = ~w5687 & ~w3019;
assign w4252 = w6713 & ~w1923;
assign w4253 = (w5997 & w7134) | (w5997 & w4024) | (w7134 & w4024);
assign w4254 = (w5178 & w5375) | (w5178 & w4748) | (w5375 & w4748);
assign w4255 = (w3330 & w350) | (w3330 & w5255) | (w350 & w5255);
assign w4256 = ~w6614 | w4123;
assign w4257 = w649 & w4003;
assign w4258 = w4188 & ~w6254;
assign w4259 = ~w2294 & w5522;
assign w4260 = ~w504 & ~w5015;
assign w4261 = ~w1827 & w975;
assign w4262 = ~w3333 & w4068;
assign w4263 = (~w6680 & w1714) | (~w6680 & w7356) | (w1714 & w7356);
assign w4264 = (~w2847 & w7121) | (~w2847 & w5670) | (w7121 & w5670);
assign w4265 = ~w1831 & ~w4402;
assign w4266 = ~w3223 & ~w389;
assign w4267 = (w5204 & w1770) | (w5204 & ~w7150) | (w1770 & ~w7150);
assign w4268 = (~w5178 & w7249) | (~w5178 & w4386) | (w7249 & w4386);
assign w4269 = (w7644 & w1353) | (w7644 & w2579) | (w1353 & w2579);
assign w4270 = (w1284 & w6537) | (w1284 & w7401) | (w6537 & w7401);
assign w4271 = ~w426 & ~w3072;
assign w4272 = (~w2806 & w1117) | (~w2806 & w2804) | (w1117 & w2804);
assign w4273 = ~w2083 & w875;
assign w4274 = (~w5998 & w7397) | (~w5998 & w246) | (w7397 & w246);
assign w4275 = ~a215 & ~b215;
assign w4276 = w2368 & w4959;
assign w4277 = (w1847 & w4085) | (w1847 & w6928) | (w4085 & w6928);
assign w4278 = (w893 & ~w6467) | (w893 & w3179) | (~w6467 & w3179);
assign w4279 = (~w3631 & w5596) | (~w3631 & w1833) | (w5596 & w1833);
assign w4280 = (~w6626 & ~w2333) | (~w6626 & w5262) | (~w2333 & w5262);
assign w4281 = (w2453 & w632) | (w2453 & w629) | (w632 & w629);
assign w4282 = ~w7000 & w5849;
assign w4283 = (w5419 & w7259) | (w5419 & w2316) | (w7259 & w2316);
assign w4284 = ~w5951 & w3353;
assign w4285 = ~w1735 & w4130;
assign w4286 = ~w174 & w3847;
assign w4287 = ~w4596 & w1910;
assign w4288 = w3365 & w5464;
assign w4289 = ~w2261 & ~w5693;
assign w4290 = (w6965 & ~w7097) | (w6965 & w491) | (~w7097 & w491);
assign w4291 = (w5484 & w2302) | (w5484 & w21) | (w2302 & w21);
assign w4292 = (~w7302 & w4030) | (~w7302 & w503) | (w4030 & w503);
assign w4293 = (~w5881 & w1290) | (~w5881 & w1488) | (w1290 & w1488);
assign w4294 = ~w2439 & ~w5660;
assign w4295 = ~w319 & w872;
assign w4296 = w6706 & ~w187;
assign w4297 = ~a173 & ~b173;
assign w4298 = (~w5178 & w6631) | (~w5178 & w6333) | (w6631 & w6333);
assign w4299 = ~w1718 & ~w5404;
assign w4300 = ~w5762 & ~w290;
assign w4301 = (~w5178 & w3921) | (~w5178 & w1040) | (w3921 & w1040);
assign w4302 = (~w4499 & w3145) | (~w4499 & w5391) | (w3145 & w5391);
assign w4303 = w1321 & w5639;
assign w4304 = (w7238 & w5014) | (w7238 & w7140) | (w5014 & w7140);
assign w4305 = (~w6844 & w6183) | (~w6844 & w3251) | (w6183 & w3251);
assign w4306 = a97 & b97;
assign w4307 = (~w6177 & w2241) | (~w6177 & w2466) | (w2241 & w2466);
assign w4308 = ~w7604 & w6596;
assign w4309 = (~w3989 & w1134) | (~w3989 & ~w1463) | (w1134 & ~w1463);
assign w4310 = ~w6697 & ~w334;
assign w4311 = (w138 & w4622) | (w138 & ~w5484) | (w4622 & ~w5484);
assign w4312 = (w5417 & w3339) | (w5417 & w4673) | (w3339 & w4673);
assign w4313 = w1892 & w5749;
assign w4314 = (w2417 & w2909) | (w2417 & w5007) | (w2909 & w5007);
assign w4315 = (~w2847 & w2633) | (~w2847 & w6391) | (w2633 & w6391);
assign w4316 = (w5045 & w3245) | (w5045 & ~w2456) | (w3245 & ~w2456);
assign w4317 = ~w6558 & w7471;
assign w4318 = (w7024 & w2962) | (w7024 & ~w3847) | (w2962 & ~w3847);
assign w4319 = (w2793 & w1565) | (w2793 & w7233) | (w1565 & w7233);
assign w4320 = w4412 & w1515;
assign w4321 = w4468 & ~w1285;
assign w4322 = (w6748 & ~w1868) | (w6748 & w6832) | (~w1868 & w6832);
assign w4323 = ~w4898 & w5745;
assign w4324 = (w5222 & w3301) | (w5222 & ~w3819) | (w3301 & ~w3819);
assign w4325 = ~a194 & ~b194;
assign w4326 = (w5403 & w1484) | (w5403 & w5150) | (w1484 & w5150);
assign w4327 = w5257 & w3391;
assign w4328 = ~w3551 & w2725;
assign w4329 = (w740 & w850) | (w740 & w4699) | (w850 & w4699);
assign w4330 = a118 & b118;
assign w4331 = ~w4132 & ~w3717;
assign w4332 = (w1609 & w2778) | (w1609 & ~w343) | (w2778 & ~w343);
assign w4333 = a45 & b45;
assign w4334 = (~w5834 & w421) | (~w5834 & w7065) | (w421 & w7065);
assign w4335 = (w6945 & w1462) | (w6945 & w3494) | (w1462 & w3494);
assign w4336 = ~w3122 & w2883;
assign w4337 = ~w1555 & w5842;
assign w4338 = (w860 & ~w2380) | (w860 & w2964) | (~w2380 & w2964);
assign w4339 = w6966 & w1331;
assign w4340 = ~w2603 & w1323;
assign w4341 = (~w7397 & w4095) | (~w7397 & w1870) | (w4095 & w1870);
assign w4342 = (~w6252 & w84) | (~w6252 & w4232) | (w84 & w4232);
assign w4343 = (w5069 & w5841) | (w5069 & w5198) | (w5841 & w5198);
assign w4344 = w6002 & ~w3166;
assign w4345 = (w1163 & w2677) | (w1163 & ~w1770) | (w2677 & ~w1770);
assign w4346 = (~w1621 & ~w384) | (~w1621 & w6803) | (~w384 & w6803);
assign w4347 = ~w7053 & w5519;
assign w4348 = ~w1285 & w4504;
assign w4349 = (~w472 & w2304) | (~w472 & w2705) | (w2304 & w2705);
assign w4350 = ~a75 & ~b75;
assign w4351 = (w4149 & ~w5194) | (w4149 & ~w4488) | (~w5194 & ~w4488);
assign w4352 = ~w6344 & ~w1841;
assign w4353 = w6452 & w4030;
assign w4354 = (~w6019 & w4544) | (~w6019 & w1604) | (w4544 & w1604);
assign w4355 = ~w4912 & ~w6254;
assign w4356 = (w2065 & w4668) | (w2065 & w2014) | (w4668 & w2014);
assign w4357 = w4442 & w6873;
assign w4358 = w6429 & w6323;
assign w4359 = w2598 & ~w1314;
assign w4360 = (w4962 & w3931) | (w4962 & w7315) | (w3931 & w7315);
assign w4361 = w5559 & ~w5391;
assign w4362 = (~w3741 & w1077) | (~w3741 & w6254) | (w1077 & w6254);
assign w4363 = (w681 & w1100) | (w681 & w6671) | (w1100 & w6671);
assign w4364 = ~w1179 & ~w7387;
assign w4365 = (w5513 & w4272) | (w5513 & ~w3119) | (w4272 & ~w3119);
assign w4366 = ~a21 & ~b21;
assign w4367 = w4496 & w2966;
assign w4368 = w6588 & ~w3807;
assign w4369 = (w755 & w6042) | (w755 & w2818) | (w6042 & w2818);
assign w4370 = (~w1611 & w6674) | (~w1611 & w4878) | (w6674 & w4878);
assign w4371 = (~w4840 & w1721) | (~w4840 & w4150) | (w1721 & w4150);
assign w4372 = (~w3033 & w2220) | (~w3033 & w628) | (w2220 & w628);
assign w4373 = (~w5325 & w276) | (~w5325 & w5601) | (w276 & w5601);
assign w4374 = ~w123 & ~w2212;
assign w4375 = ~w3782 & w4082;
assign w4376 = w1792 & ~w2814;
assign w4377 = a58 & b58;
assign w4378 = ~w1743 & ~w6520;
assign w4379 = w2011 & ~w3052;
assign w4380 = ~w4430 & w1843;
assign w4381 = w5424 & w1349;
assign w4382 = ~w3136 & w1066;
assign w4383 = (w1847 & ~w5655) | (w1847 & w6710) | (~w5655 & w6710);
assign w4384 = ~w5242 & w7552;
assign w4385 = (w5774 & ~w3774) | (w5774 & w2985) | (~w3774 & w2985);
assign w4386 = (~w5325 & w4015) | (~w5325 & w2392) | (w4015 & w2392);
assign w4387 = ~w638 & ~w3294;
assign w4388 = ~w5875 & w3722;
assign w4389 = (w3074 & w7323) | (w3074 & w4689) | (w7323 & w4689);
assign w4390 = (w5910 & w2620) | (w5910 & ~w629) | (w2620 & ~w629);
assign w4391 = (~w2399 & w1966) | (~w2399 & w3485) | (w1966 & w3485);
assign w4392 = ~w4885 & w2326;
assign w4393 = w1143 & w6096;
assign w4394 = ~w5681 & w5828;
assign w4395 = (w961 & w3565) | (w961 & ~w3119) | (w3565 & ~w3119);
assign w4396 = w5972 & ~w2336;
assign w4397 = (w3318 & w5811) | (w3318 & w545) | (w5811 & w545);
assign w4398 = (~w7283 & w6887) | (~w7283 & w5118) | (w6887 & w5118);
assign w4399 = (w5178 & w6693) | (w5178 & w4416) | (w6693 & w4416);
assign w4400 = (w7575 & w7397) | (w7575 & w4801) | (w7397 & w4801);
assign w4401 = ~w2852 & w6260;
assign w4402 = a70 & b70;
assign w4403 = ~w7350 & ~w63;
assign w4404 = (~w7199 & w1203) | (~w7199 & w894) | (w1203 & w894);
assign w4405 = (w5910 & w2620) | (w5910 & ~w173) | (w2620 & ~w173);
assign w4406 = (~w5089 & w4293) | (~w5089 & w1329) | (w4293 & w1329);
assign w4407 = (~w6100 & w5931) | (~w6100 & w4772) | (w5931 & w4772);
assign w4408 = (w410 & w5167) | (w410 & ~w5098) | (w5167 & ~w5098);
assign w4409 = ~a168 & ~b168;
assign w4410 = w1685 & w3019;
assign w4411 = (w1496 & w4046) | (w1496 & ~w5417) | (w4046 & ~w5417);
assign w4412 = ~a198 & ~b198;
assign w4413 = (w1665 & w6399) | (w1665 & w5674) | (w6399 & w5674);
assign w4414 = ~w3260 & ~w6915;
assign w4415 = ~w3033 & ~w4808;
assign w4416 = (w5325 & w3225) | (w5325 & w5356) | (w3225 & w5356);
assign w4417 = ~w4543 & ~w3208;
assign w4418 = w2019 & ~w1544;
assign w4419 = ~w4238 & w2433;
assign w4420 = w4716 & ~w5106;
assign w4421 = ~w931 & w766;
assign w4422 = ~w1463 & ~w6609;
assign w4423 = ~w2540 & w3311;
assign w4424 = w6299 | ~w1158;
assign w4425 = ~w2597 & ~w3137;
assign w4426 = (~w6100 & w79) | (~w6100 & w2224) | (w79 & w2224);
assign w4427 = (w632 & w3407) | (w632 & ~w693) | (w3407 & ~w693);
assign w4428 = w1952 & w6187;
assign w4429 = (w1252 & w4596) | (w1252 & w2905) | (w4596 & w2905);
assign w4430 = ~w6703 & w5960;
assign w4431 = w4004 & ~w2693;
assign w4432 = (w2628 & ~w6467) | (w2628 & w6173) | (~w6467 & w6173);
assign w4433 = (w5760 & ~w5977) | (w5760 & w6181) | (~w5977 & w6181);
assign w4434 = (w7626 & w815) | (w7626 & w1214) | (w815 & w1214);
assign w4435 = (w5834 & w2219) | (w5834 & w5187) | (w2219 & w5187);
assign w4436 = (w6100 & w6086) | (w6100 & w7543) | (w6086 & w7543);
assign w4437 = w2197 & ~w3669;
assign w4438 = a106 & b106;
assign w4439 = (w2985 & w3916) | (w2985 & w3615) | (w3916 & w3615);
assign w4440 = (w3364 & w805) | (w3364 & w1809) | (w805 & w1809);
assign w4441 = (~w3903 & w6134) | (~w3903 & ~w5403) | (w6134 & ~w5403);
assign w4442 = ~w3953 & w6192;
assign w4443 = (w501 & w1257) | (w501 & w6563) | (w1257 & w6563);
assign w4444 = w1228 & ~w6147;
assign w4445 = ~w5033 & ~w2731;
assign w4446 = (~w2460 & w100) | (~w2460 & w7145) | (w100 & w7145);
assign w4447 = w2451 & w6754;
assign w4448 = a96 & b96;
assign w4449 = ~w6330 & ~w3988;
assign w4450 = w3942 & w1929;
assign w4451 = (~w3868 & w6927) | (~w3868 & w6881) | (w6927 & w6881);
assign w4452 = (w2952 & w7263) | (w2952 & w4867) | (w7263 & w4867);
assign w4453 = (w6942 & w6148) | (w6942 & ~w7097) | (w6148 & ~w7097);
assign w4454 = (w4011 & w5871) | (w4011 & w2028) | (w5871 & w2028);
assign w4455 = w6758 & w5080;
assign w4456 = (w4006 & w2944) | (w4006 & ~w1770) | (w2944 & ~w1770);
assign w4457 = a39 & b39;
assign w4458 = w7391 & ~w4759;
assign w4459 = w3883 & w5507;
assign w4460 = (~w6100 & w224) | (~w6100 & w1017) | (w224 & w1017);
assign w4461 = ~w3070 & ~w4906;
assign w4462 = ~w4900 & w7103;
assign w4463 = (w6572 & w4621) | (w6572 & ~w2318) | (w4621 & ~w2318);
assign w4464 = (w6415 & ~w4459) | (w6415 & w2462) | (~w4459 & w2462);
assign w4465 = ~w84 & w3701;
assign w4466 = w887 & w4742;
assign w4467 = a41 & b41;
assign w4468 = ~a67 & ~b67;
assign w4469 = (w5212 & w3786) | (w5212 & w2199) | (w3786 & w2199);
assign w4470 = ~w5858 & w6685;
assign w4471 = w5629 & w2010;
assign w4472 = ~w5604 & ~w3239;
assign w4473 = w833 & w3050;
assign w4474 = w5983 & ~w2591;
assign w4475 = w6444 & w5128;
assign w4476 = ~a42 & ~b42;
assign w4477 = (w6100 & w1893) | (w6100 & w6910) | (w1893 & w6910);
assign w4478 = ~w6520 & ~w1369;
assign w4479 = (~w4176 & ~w3384) | (~w4176 & w6530) | (~w3384 & w6530);
assign w4480 = ~w2182 & w5729;
assign w4481 = (~w5178 & w2028) | (~w5178 & w4454) | (w2028 & w4454);
assign w4482 = ~w5018 & ~w133;
assign w4483 = w3083 & ~w6679;
assign w4484 = (~w5178 & w5855) | (~w5178 & w1156) | (w5855 & w1156);
assign w4485 = (w6215 & ~w6031) | (w6215 & w828) | (~w6031 & w828);
assign w4486 = ~w4430 & w7292;
assign w4487 = (w1489 & w230) | (w1489 & w7472) | (w230 & w7472);
assign w4488 = w3660 & ~w2600;
assign w4489 = (w1006 & w4656) | (w1006 & w3785) | (w4656 & w3785);
assign w4490 = (w6100 & w6478) | (w6100 & w7395) | (w6478 & w7395);
assign w4491 = w3424 & ~w7468;
assign w4492 = ~w2056 & ~w710;
assign w4493 = (w3989 & w5483) | (w3989 & w3448) | (w5483 & w3448);
assign w4494 = ~w5627 & w3672;
assign w4495 = (w4855 & w5916) | (w4855 & ~w5430) | (w5916 & ~w5430);
assign w4496 = ~w2803 & ~w1974;
assign w4497 = ~a93 & ~b93;
assign w4498 = ~w7590 & ~w7621;
assign w4499 = ~a97 & ~b97;
assign w4500 = ~w6208 & ~w5884;
assign w4501 = (~w236 & w811) | (~w236 & w1095) | (w811 & w1095);
assign w4502 = (w3774 & w4590) | (w3774 & w1994) | (w4590 & w1994);
assign w4503 = ~w7363 & ~w6087;
assign w4504 = ~w1300 & ~w5425;
assign w4505 = ~w7291 & ~w576;
assign w4506 = (~w4468 & ~w4504) | (~w4468 & w5794) | (~w4504 & w5794);
assign w4507 = (~w7471 & w3146) | (~w7471 & w1265) | (w3146 & w1265);
assign w4508 = ~w3183 & ~w841;
assign w4509 = (w6860 & w4136) | (w6860 & w4768) | (w4136 & w4768);
assign w4510 = (~w2456 & w5325) | (~w2456 & w6894) | (w5325 & w6894);
assign w4511 = ~w2441 & w3173;
assign w4512 = w1821 & ~w4745;
assign w4513 = ~w2127 & w7166;
assign w4514 = ~w7044 & w7625;
assign w4515 = ~w2070 & ~w459;
assign w4516 = (w1628 & w1589) | (w1628 & w5233) | (w1589 & w5233);
assign w4517 = ~w2847 & w1704;
assign w4518 = (~w6911 & w6271) | (~w6911 & w3679) | (w6271 & w3679);
assign w4519 = ~w2496 & w5392;
assign w4520 = (w6100 & w1010) | (w6100 & w6623) | (w1010 & w6623);
assign w4521 = (~w7385 & w3914) | (~w7385 & w7509) | (w3914 & w7509);
assign w4522 = ~w3014 & w3396;
assign w4523 = ~w6927 & w3868;
assign w4524 = (~w5325 & w1018) | (~w5325 & w2266) | (w1018 & w2266);
assign w4525 = w7010 & w2960;
assign w4526 = ~w5464 & ~w5555;
assign w4527 = (~w6100 & w4589) | (~w6100 & w2573) | (w4589 & w2573);
assign w4528 = (w2627 & w5065) | (w2627 & ~w2294) | (w5065 & ~w2294);
assign w4529 = ~w2630 & w6851;
assign w4530 = a119 & b119;
assign w4531 = ~w1137 & ~w1678;
assign w4532 = ~w3342 & ~w765;
assign w4533 = ~w5983 & ~w6210;
assign w4534 = ~w212 & ~w7354;
assign w4535 = (w5178 & w6850) | (w5178 & w7098) | (w6850 & w7098);
assign w4536 = w1338 & ~w52;
assign w4537 = (w6353 & w650) | (w6353 & w2375) | (w650 & w2375);
assign w4538 = w3133 & w1025;
assign w4539 = (~w3952 & w1979) | (~w3952 & w6506) | (w1979 & w6506);
assign w4540 = w4320 & w1515;
assign w4541 = (~w5066 & w2178) | (~w5066 & w3576) | (w2178 & w3576);
assign w4542 = (w5022 & w420) | (w5022 & w329) | (w420 & w329);
assign w4543 = (~w2037 & w20) | (~w2037 & w4943) | (w20 & w4943);
assign w4544 = (~w3868 & w4451) | (~w3868 & w4811) | (w4451 & w4811);
assign w4545 = a63 & b63;
assign w4546 = (w5752 & w7205) | (w5752 & w5846) | (w7205 & w5846);
assign w4547 = (w3774 & w5211) | (w3774 & w928) | (w5211 & w928);
assign w4548 = (w1479 & w4000) | (w1479 & w44) | (w4000 & w44);
assign w4549 = (~w2838 & w7582) | (~w2838 & ~w3894) | (w7582 & ~w3894);
assign w4550 = ~w4784 & ~w2846;
assign w4551 = (w6100 & w6156) | (w6100 & w7230) | (w6156 & w7230);
assign w4552 = (w2627 & w5407) | (w2627 & w5048) | (w5407 & w5048);
assign w4553 = (~w2627 & w6622) | (~w2627 & w2729) | (w6622 & w2729);
assign w4554 = (w1515 & w1133) | (w1515 & w4540) | (w1133 & w4540);
assign w4555 = ~w2005 & w1427;
assign w4556 = ~w1570 & ~w6587;
assign w4557 = (w6681 & w6675) | (w6681 & w6958) | (w6675 & w6958);
assign w4558 = (w236 & w2419) | (w236 & w4029) | (w2419 & w4029);
assign w4559 = w4157 & w1104;
assign w4560 = (~w5998 & w4967) | (~w5998 & w4274) | (w4967 & w4274);
assign w4561 = (w6570 & w6787) | (w6570 & ~w3391) | (w6787 & ~w3391);
assign w4562 = ~w2847 & w794;
assign w4563 = ~w945 & ~w458;
assign w4564 = a231 & b231;
assign w4565 = (~w3986 & w4953) | (~w3986 & w1222) | (w4953 & w1222);
assign w4566 = ~w471 & ~w5560;
assign w4567 = w990 & ~w788;
assign w4568 = (w5672 & w4396) | (w5672 & w1333) | (w4396 & w1333);
assign w4569 = ~w7391 & ~w2405;
assign w4570 = ~w1925 & ~w6760;
assign w4571 = (~w4503 & w2558) | (~w4503 & w2248) | (w2558 & w2248);
assign w4572 = ~w6104 & w7421;
assign w4573 = (~w1879 & w6592) | (~w1879 & w558) | (w6592 & w558);
assign w4574 = ~w3512 & ~w3602;
assign w4575 = ~w3333 & w2928;
assign w4576 = (w4044 & w1707) | (w4044 & ~w6501) | (w1707 & ~w6501);
assign w4577 = (w5655 & w4547) | (w5655 & w2358) | (w4547 & w2358);
assign w4578 = (~w5178 & w3820) | (~w5178 & w7191) | (w3820 & w7191);
assign w4579 = w1832 & w1548;
assign w4580 = (~w1053 & ~w4068) | (~w1053 & w509) | (~w4068 & w509);
assign w4581 = (~w5834 & w2933) | (~w5834 & w5913) | (w2933 & w5913);
assign w4582 = (w7255 & w5850) | (w7255 & w4803) | (w5850 & w4803);
assign w4583 = (w5298 & w6052) | (w5298 & ~w632) | (w6052 & ~w632);
assign w4584 = ~a27 & ~b27;
assign w4585 = ~w2798 & w4843;
assign w4586 = (~w5325 & w1079) | (~w5325 & w3977) | (w1079 & w3977);
assign w4587 = ~a177 & ~b177;
assign w4588 = ~w4690 & w1728;
assign w4589 = (w1035 & w7450) | (w1035 & w784) | (w7450 & w784);
assign w4590 = (w3461 & w3889) | (w3461 & w6768) | (w3889 & w6768);
assign w4591 = ~w7460 & w2177;
assign w4592 = (w6151 & w2727) | (w6151 & w1291) | (w2727 & w1291);
assign w4593 = ~w3368 & ~w4307;
assign w4594 = w4690 & w2463;
assign w4595 = (w5054 & w823) | (w5054 & w810) | (w823 & w810);
assign w4596 = ~w5745 & w69;
assign w4597 = ~w6791 & ~w727;
assign w4598 = ~w4680 & ~w2605;
assign w4599 = ~w5883 & w7604;
assign w4600 = (~w968 & w5330) | (~w968 & w6310) | (w5330 & w6310);
assign w4601 = ~w6851 & w6221;
assign w4602 = ~w5782 & w7111;
assign w4603 = ~w3735 & ~w4677;
assign w4604 = w2588 & w6813;
assign w4605 = w6304 & ~w6458;
assign w4606 = ~w2724 & ~w6548;
assign w4607 = ~w4737 & ~w5603;
assign w4608 = (~w563 & w7176) | (~w563 & w2583) | (w7176 & w2583);
assign w4609 = (~w7291 & w488) | (~w7291 & w1571) | (w488 & w1571);
assign w4610 = w1071 & ~w6450;
assign w4611 = w1216 & ~w3210;
assign w4612 = ~a60 & ~b60;
assign w4613 = ~w1728 & w2094;
assign w4614 = ~w7381 & ~w2586;
assign w4615 = w4850 & w5421;
assign w4616 = ~a179 & ~b179;
assign w4617 = w247 & ~w6252;
assign w4618 = w1378 & ~w2175;
assign w4619 = w6805 & w2661;
assign w4620 = ~w5466 & ~w424;
assign w4621 = w3836 & w6572;
assign w4622 = w1900 & ~w3348;
assign w4623 = ~w6310 & w1542;
assign w4624 = w6633 & w3883;
assign w4625 = (w5655 & w2509) | (w5655 & w2467) | (w2509 & w2467);
assign w4626 = (w7599 & w6265) | (w7599 & w5902) | (w6265 & w5902);
assign w4627 = (~w5735 & w5690) | (~w5735 & w3380) | (w5690 & w3380);
assign w4628 = (~w5901 & w3798) | (~w5901 & w4902) | (w3798 & w4902);
assign w4629 = (w1328 & w5982) | (w1328 & w7340) | (w5982 & w7340);
assign w4630 = ~w1393 & ~w3216;
assign w4631 = (w5655 & w1538) | (w5655 & w5988) | (w1538 & w5988);
assign w4632 = a7 & b7;
assign w4633 = (w6395 & w7524) | (w6395 & w3800) | (w7524 & w3800);
assign w4634 = (~w1760 & w2408) | (~w1760 & w5184) | (w2408 & w5184);
assign w4635 = w5058 & w6396;
assign w4636 = ~w7538 & ~w3626;
assign w4637 = ~w3591 & ~w6649;
assign w4638 = ~w3887 & ~w7536;
assign w4639 = w46 & ~w3145;
assign w4640 = ~w4257 & w6397;
assign w4641 = w5816 & w2578;
assign w4642 = (w4182 & w4096) | (w4182 & w5969) | (w4096 & w5969);
assign w4643 = a107 & b107;
assign w4644 = ~w2930 & ~w5742;
assign w4645 = w2540 & ~w6100;
assign w4646 = (~w7161 & w6060) | (~w7161 & w670) | (w6060 & w670);
assign w4647 = (~w3375 & w4418) | (~w3375 & w3876) | (w4418 & w3876);
assign w4648 = ~a115 & ~b115;
assign w4649 = (~w858 & w6837) | (~w858 & w3858) | (w6837 & w3858);
assign w4650 = (~w1516 & w891) | (~w1516 & w4269) | (w891 & w4269);
assign w4651 = ~w1980 & ~w1967;
assign w4652 = w1751 & w1399;
assign w4653 = (w5178 & w2983) | (w5178 & w4794) | (w2983 & w4794);
assign w4654 = ~w3695 & ~w7642;
assign w4655 = w7386 & w5403;
assign w4656 = (w6649 & w6532) | (w6649 & w6658) | (w6532 & w6658);
assign w4657 = w1813 & w7421;
assign w4658 = w1868 & w4338;
assign w4659 = w7113 & ~w3819;
assign w4660 = w4132 & ~w3490;
assign w4661 = ~w1610 & ~w7536;
assign w4662 = (~w9 & w2245) | (~w9 & w2966) | (w2245 & w2966);
assign w4663 = w4867 & ~w5511;
assign w4664 = (w4102 & w6800) | (w4102 & w4549) | (w6800 & w4549);
assign w4665 = ~w4287 & w4261;
assign w4666 = (w7197 & w6337) | (w7197 & w1050) | (w6337 & w1050);
assign w4667 = (w6082 & w1596) | (w6082 & w1566) | (w1596 & w1566);
assign w4668 = (~w5106 & w4716) | (~w5106 & w6017) | (w4716 & w6017);
assign w4669 = w3835 & ~w7404;
assign w4670 = ~w6293 & ~w2355;
assign w4671 = (w1284 & w6537) | (w1284 & w1555) | (w6537 & w1555);
assign w4672 = ~w7302 & ~w7363;
assign w4673 = (~w887 & w2599) | (~w887 & ~w2311) | (w2599 & ~w2311);
assign w4674 = ~a237 & ~b237;
assign w4675 = ~w7345 & ~w6712;
assign w4676 = ~w1053 & ~w7489;
assign w4677 = ~a191 & ~b191;
assign w4678 = ~w3603 & ~w6314;
assign w4679 = ~w931 & w5977;
assign w4680 = ~w5346 & w3157;
assign w4681 = ~w2515 & ~w972;
assign w4682 = ~w3500 & ~w262;
assign w4683 = (w1336 & w3975) | (w1336 & w3952) | (w3975 & w3952);
assign w4684 = (~w1866 & ~w4480) | (~w1866 & w5201) | (~w4480 & w5201);
assign w4685 = ~w6013 & ~w5361;
assign w4686 = ~w3331 & w2021;
assign w4687 = ~w5598 & ~w4333;
assign w4688 = ~w576 & w1420;
assign w4689 = ~w3905 & ~w7286;
assign w4690 = ~w4918 & w4027;
assign w4691 = ~w3235 & ~w5051;
assign w4692 = ~w3997 & ~w3244;
assign w4693 = (w3496 & w2389) | (w3496 & ~w4143) | (w2389 & ~w4143);
assign w4694 = (w1279 & ~w139) | (w1279 & ~w6099) | (~w139 & ~w6099);
assign w4695 = (w5178 & w2170) | (w5178 & w5865) | (w2170 & w5865);
assign w4696 = (~w1367 & w4876) | (~w1367 & w6529) | (w4876 & w6529);
assign w4697 = ~w5279 & ~w2658;
assign w4698 = (w6100 & w1662) | (w6100 & w4565) | (w1662 & w4565);
assign w4699 = w7546 & w740;
assign w4700 = (w1658 & w1308) | (w1658 & w7498) | (w1308 & w7498);
assign w4701 = (w4732 & w1962) | (w4732 & ~w4867) | (w1962 & ~w4867);
assign w4702 = w4190 | w3105;
assign w4703 = (w304 & w1941) | (w304 & ~w7015) | (w1941 & ~w7015);
assign w4704 = (w1770 & w6601) | (w1770 & w6199) | (w6601 & w6199);
assign w4705 = (w3570 & ~w5152) | (w3570 & w1330) | (~w5152 & w1330);
assign w4706 = ~w4176 & ~w5676;
assign w4707 = (w3986 & w592) | (w3986 & w2207) | (w592 & w2207);
assign w4708 = ~w4918 & w6149;
assign w4709 = (w839 & w5178) | (w839 & w3906) | (w5178 & w3906);
assign w4710 = ~w3735 & ~w3123;
assign w4711 = w113 & ~w5203;
assign w4712 = (w2985 & w5621) | (w2985 & w2038) | (w5621 & w2038);
assign w4713 = ~w1632 & ~w6643;
assign w4714 = w3755 & w7273;
assign w4715 = (~w6945 & w3361) | (~w6945 & w5509) | (w3361 & w5509);
assign w4716 = w4306 & ~w5106;
assign w4717 = ~w4497 & ~w5005;
assign w4718 = ~w4843 & w1878;
assign w4719 = (w5204 & w5395) | (w5204 & ~w7150) | (w5395 & ~w7150);
assign w4720 = ~w808 & ~w4855;
assign w4721 = ~w318 & w3200;
assign w4722 = ~w314 & w2986;
assign w4723 = (~w686 & w7368) | (~w686 & w33) | (w7368 & w33);
assign w4724 = (w3774 & w2264) | (w3774 & w7464) | (w2264 & w7464);
assign w4725 = w2799 & w2043;
assign w4726 = w4638 & ~w5927;
assign w4727 = (w287 & w2667) | (w287 & w4173) | (w2667 & w4173);
assign w4728 = ~w763 & w1428;
assign w4729 = (w2639 & w5097) | (w2639 & w484) | (w5097 & w484);
assign w4730 = w807 & w4459;
assign w4731 = (~w3318 & w7295) | (~w3318 & w6494) | (w7295 & w6494);
assign w4732 = w3643 & w7227;
assign w4733 = (~w434 & ~w2311) | (~w434 & w6413) | (~w2311 & w6413);
assign w4734 = (w5146 & w6275) | (w5146 & w7015) | (w6275 & w7015);
assign w4735 = (~w6184 & w3094) | (~w6184 & w3014) | (w3094 & w3014);
assign w4736 = (w5325 & w1494) | (w5325 & w1350) | (w1494 & w1350);
assign w4737 = ~w441 & ~w6984;
assign w4738 = w5888 & ~w388;
assign w4739 = (~w215 & w634) | (~w215 & w5479) | (w634 & w5479);
assign w4740 = (w5556 & ~w3824) | (w5556 & w1964) | (~w3824 & w1964);
assign w4741 = ~w7190 & ~w6772;
assign w4742 = w5958 & ~w4564;
assign w4743 = w5881 & w3746;
assign w4744 = ~w2829 & ~w2267;
assign w4745 = w1574 & w4379;
assign w4746 = ~a153 & ~b153;
assign w4747 = ~w5762 & ~w640;
assign w4748 = (~w4143 & w2134) | (~w4143 & w3757) | (w2134 & w3757);
assign w4749 = ~w2636 & ~w1860;
assign w4750 = w2766 & w6421;
assign w4751 = ~w6117 & ~w4215;
assign w4752 = ~w3455 & w546;
assign w4753 = (w7513 & w5985) | (w7513 & w4507) | (w5985 & w4507);
assign w4754 = ~w1957 & w6619;
assign w4755 = (w5501 & w5093) | (w5501 & w563) | (w5093 & w563);
assign w4756 = ~w6516 & ~w1940;
assign w4757 = (~w144 & ~w5484) | (~w144 & w6721) | (~w5484 & w6721);
assign w4758 = (w5178 & w1376) | (w5178 & w5668) | (w1376 & w5668);
assign w4759 = ~a37 & ~b37;
assign w4760 = (w752 & w2123) | (w752 & w1871) | (w2123 & w1871);
assign w4761 = w2591 & ~w5416;
assign w4762 = ~w5182 & ~w2882;
assign w4763 = w2496 & ~w5392;
assign w4764 = (~w5743 & ~w1754) | (~w5743 & w5263) | (~w1754 & w5263);
assign w4765 = ~a87 & ~b87;
assign w4766 = (~w7108 & w6143) | (~w7108 & w1512) | (w6143 & w1512);
assign w4767 = w3365 & ~w7629;
assign w4768 = ~w3616 & ~w6628;
assign w4769 = ~w4435 & ~w31;
assign w4770 = ~w1315 & w1598;
assign w4771 = (~w6387 & w6265) | (~w6387 & w1562) | (w6265 & w1562);
assign w4772 = (w4908 & w3159) | (w4908 & w3197) | (w3159 & w3197);
assign w4773 = w4777 & ~w1903;
assign w4774 = (~w3952 & w1207) | (~w3952 & w4525) | (w1207 & w4525);
assign w4775 = ~a38 & ~b38;
assign w4776 = w6954 & ~w4199;
assign w4777 = ~w6713 & w6911;
assign w4778 = ~w3471 & w1605;
assign w4779 = (w2813 & w2684) | (w2813 & w4857) | (w2684 & w4857);
assign w4780 = (~w2019 & w7196) | (~w2019 & w4859) | (w7196 & w4859);
assign w4781 = ~w5627 & w4260;
assign w4782 = (w2773 & w6715) | (w2773 & ~w2876) | (w6715 & ~w2876);
assign w4783 = (w7126 & w5909) | (w7126 & ~w1770) | (w5909 & ~w1770);
assign w4784 = ~a79 & ~b79;
assign w4785 = w3595 & w5581;
assign w4786 = (w2074 & w5901) | (w2074 & w4183) | (w5901 & w4183);
assign w4787 = ~w2229 & w4479;
assign w4788 = ~a242 & ~b242;
assign w4789 = ~w5159 & ~w3992;
assign w4790 = w1204 & ~w2068;
assign w4791 = w5362 & ~w5223;
assign w4792 = (w5266 & ~w5430) | (w5266 & w6759) | (~w5430 & w6759);
assign w4793 = w2793 & ~w6254;
assign w4794 = (~w2965 & w4158) | (~w2965 & w5166) | (w4158 & w5166);
assign w4795 = w103 & w2548;
assign w4796 = (w4433 & w4164) | (w4433 & w7575) | (w4164 & w7575);
assign w4797 = (w5178 & w3147) | (w5178 & w1370) | (w3147 & w1370);
assign w4798 = (w4392 & w4155) | (w4392 & ~w587) | (w4155 & ~w587);
assign w4799 = (~w4651 & ~w5484) | (~w4651 & w4220) | (~w5484 & w4220);
assign w4800 = (w2985 & w3699) | (w2985 & w7612) | (w3699 & w7612);
assign w4801 = ~w7078 & w7575;
assign w4802 = ~w1860 & ~w1300;
assign w4803 = ~w3866 & w4615;
assign w4804 = (w4824 & ~w3119) | (w4824 & w7402) | (~w3119 & w7402);
assign w4805 = (w7322 & w5268) | (w7322 & w7280) | (w5268 & w7280);
assign w4806 = ~w5480 & ~w3366;
assign w4807 = ~w3057 & w3962;
assign w4808 = a241 & b241;
assign w4809 = w5380 & ~w2876;
assign w4810 = (w5590 & w6868) | (w5590 & w3309) | (w6868 & w3309);
assign w4811 = ~w3989 & w3356;
assign w4812 = (~w3078 & w5942) | (~w3078 & w380) | (w5942 & w380);
assign w4813 = (~w3318 & w659) | (~w3318 & w5047) | (w659 & w5047);
assign w4814 = w4762 & ~w2349;
assign w4815 = w3136 & w3312;
assign w4816 = (w770 & w1121) | (w770 & w4719) | (w1121 & w4719);
assign w4817 = w3631 & w2269;
assign w4818 = w103 & w6163;
assign w4819 = (w1856 & w3478) | (w1856 & ~w5958) | (w3478 & ~w5958);
assign w4820 = ~w1709 & ~w4427;
assign w4821 = (w1814 & w921) | (w1814 & w6676) | (w921 & w6676);
assign w4822 = ~a249 & ~b249;
assign w4823 = w823 & w5054;
assign w4824 = (w4069 & ~w4102) | (w4069 & w2032) | (~w4102 & w2032);
assign w4825 = (w5821 & w7322) | (w5821 & ~w6174) | (w7322 & ~w6174);
assign w4826 = (w1123 & w6764) | (w1123 & ~w2876) | (w6764 & ~w2876);
assign w4827 = (w5930 & ~w2080) | (w5930 & ~w6712) | (~w2080 & ~w6712);
assign w4828 = w2569 & ~w4934;
assign w4829 = ~w4840 & w5666;
assign w4830 = ~b255 & ~a255;
assign w4831 = w6553 & ~w1245;
assign w4832 = (~w5655 & w3890) | (~w5655 & w4744) | (w3890 & w4744);
assign w4833 = ~w4587 & ~w1622;
assign w4834 = (~w6467 & w1928) | (~w6467 & w4343) | (w1928 & w4343);
assign w4835 = ~w7500 & w7414;
assign w4836 = (~w3842 & w2379) | (~w3842 & w6446) | (w2379 & w6446);
assign w4837 = ~w3656 & w5859;
assign w4838 = ~w5194 & w2947;
assign w4839 = ~w3769 & ~w7096;
assign w4840 = (w6100 & w1430) | (w6100 & w7584) | (w1430 & w7584);
assign w4841 = ~w4811 & ~w523;
assign w4842 = (~w4265 & w4209) | (~w4265 & w1730) | (w4209 & w1730);
assign w4843 = ~w1256 & ~w5588;
assign w4844 = w4430 & w1743;
assign w4845 = w2664 & ~w957;
assign w4846 = (w1062 & w6773) | (w1062 & ~w1516) | (w6773 & ~w1516);
assign w4847 = ~w3480 & ~w3918;
assign w4848 = w4602 & ~w1204;
assign w4849 = w4016 & w4455;
assign w4850 = ~w54 & w64;
assign w4851 = (~w1455 & w6761) | (~w1455 & w6388) | (w6761 & w6388);
assign w4852 = (~w6690 & w2202) | (~w6690 & w364) | (w2202 & w364);
assign w4853 = (~w3952 & w4930) | (~w3952 & w2737) | (w4930 & w2737);
assign w4854 = (~w4825 & w2941) | (~w4825 & w6201) | (w2941 & w6201);
assign w4855 = ~w1443 & w505;
assign w4856 = (w728 & w2575) | (w728 & ~w1649) | (w2575 & ~w1649);
assign w4857 = w517 & w7583;
assign w4858 = (w1631 & w1639) | (w1631 & w1573) | (w1639 & w1573);
assign w4859 = w1839 & ~w2019;
assign w4860 = (w1847 & w5856) | (w1847 & w7052) | (w5856 & w7052);
assign w4861 = (w7554 & w4595) | (w7554 & w6213) | (w4595 & w6213);
assign w4862 = w7362 & ~w6237;
assign w4863 = (~w5178 & w7585) | (~w5178 & w7207) | (w7585 & w7207);
assign w4864 = w1176 & ~w3166;
assign w4865 = (w6385 & w6976) | (w6385 & ~w6633) | (w6976 & ~w6633);
assign w4866 = w7378 & w2622;
assign w4867 = ~w6272 & w7541;
assign w4868 = (w4889 & w4372) | (w4889 & ~w632) | (w4372 & ~w632);
assign w4869 = (w166 & w2154) | (w166 & ~w4635) | (w2154 & ~w4635);
assign w4870 = ~w2898 & w300;
assign w4871 = (w2806 & w358) | (w2806 & w5060) | (w358 & w5060);
assign w4872 = (w5374 & w4840) | (w5374 & w636) | (w4840 & w636);
assign w4873 = (~w2021 & w2308) | (~w2021 & w7437) | (w2308 & w7437);
assign w4874 = (w2225 & w6186) | (w2225 & w4143) | (w6186 & w4143);
assign w4875 = ~w4350 & ~w625;
assign w4876 = ~w145 & ~w7132;
assign w4877 = ~w6398 & ~w4481;
assign w4878 = (~w4300 & w6843) | (~w4300 & w6114) | (w6843 & w6114);
assign w4879 = (~w3318 & w762) | (~w3318 & w1052) | (w762 & w1052);
assign w4880 = w6954 & ~w7238;
assign w4881 = a223 & b223;
assign w4882 = w3880 & w1170;
assign w4883 = ~w6533 & ~w4225;
assign w4884 = ~w2749 & ~w336;
assign w4885 = w2913 & ~w6628;
assign w4886 = ~w4681 & w7629;
assign w4887 = ~w3979 & ~w4568;
assign w4888 = w1162 & ~w4329;
assign w4889 = (w3490 & w6049) | (w3490 & w4105) | (w6049 & w4105);
assign w4890 = ~w504 & w843;
assign w4891 = ~a120 & ~b120;
assign w4892 = w6233 & ~w6281;
assign w4893 = ~w960 & ~w1610;
assign w4894 = ~w3217 & w7429;
assign w4895 = ~w5183 & ~w1753;
assign w4896 = (~w5881 & w1290) | (~w5881 & w5600) | (w1290 & w5600);
assign w4897 = (~w2945 & w3647) | (~w2945 & w3679) | (w3647 & w3679);
assign w4898 = ~a247 & ~b247;
assign w4899 = (~w3292 & ~w6451) | (~w3292 & w2429) | (~w6451 & w2429);
assign w4900 = (w2899 & w5178) | (w2899 & w3543) | (w5178 & w3543);
assign w4901 = ~w5743 & ~w3893;
assign w4902 = (~w1143 & w1457) | (~w1143 & w2221) | (w1457 & w2221);
assign w4903 = ~w2344 & ~w1391;
assign w4904 = w5119 & ~w6965;
assign w4905 = (w3461 & w5371) | (w3461 & w6152) | (w5371 & w6152);
assign w4906 = ~w7056 & ~w1371;
assign w4907 = (~w7106 & w578) | (~w7106 & w2456) | (w578 & w2456);
assign w4908 = (w1658 & w270) | (w1658 & w2481) | (w270 & w2481);
assign w4909 = (w341 & w267) | (w341 & w3668) | (w267 & w3668);
assign w4910 = (~w303 & w7411) | (~w303 & w7169) | (w7411 & w7169);
assign w4911 = ~a216 & ~b216;
assign w4912 = w1331 & w7187;
assign w4913 = (~w5296 & w1373) | (~w5296 & w6702) | (w1373 & w6702);
assign w4914 = (w671 & w7514) | (w671 & w1009) | (w7514 & w1009);
assign w4915 = (w3852 & w4899) | (w3852 & w3453) | (w4899 & w3453);
assign w4916 = (w6353 & w5846) | (w6353 & w4017) | (w5846 & w4017);
assign w4917 = w4430 & w7439;
assign w4918 = a114 & b114;
assign w4919 = (~w5257 & w7105) | (~w5257 & w2042) | (w7105 & w2042);
assign w4920 = (w5178 & w5369) | (w5178 & w3875) | (w5369 & w3875);
assign w4921 = a57 & b57;
assign w4922 = w3644 & ~w216;
assign w4923 = w4148 & ~w7510;
assign w4924 = ~w2229 & w6714;
assign w4925 = w6560 & w7506;
assign w4926 = w2869 & ~w5352;
assign w4927 = w1758 & w939;
assign w4928 = (~w3774 & w4184) | (~w3774 & w4800) | (w4184 & w4800);
assign w4929 = w3679 & ~w3533;
assign w4930 = (w5944 & w6796) | (w5944 & w3486) | (w6796 & w3486);
assign w4931 = ~w2974 & ~w5342;
assign w4932 = ~w147 & w2588;
assign w4933 = ~w5930 & ~w6392;
assign w4934 = ~w5908 & w7202;
assign w4935 = ~w6682 | ~w6860;
assign w4936 = ~w7159 & ~w370;
assign w4937 = (~w1135 & w5456) | (~w1135 & w4197) | (w5456 & w4197);
assign w4938 = (w65 & w7528) | (w65 & w7406) | (w7528 & w7406);
assign w4939 = (~w5830 & w4656) | (~w5830 & w551) | (w4656 & w551);
assign w4940 = a197 & b197;
assign w4941 = w4348 & ~w7320;
assign w4942 = ~w1308 & w2824;
assign w4943 = w3775 & ~w3630;
assign w4944 = (~w6100 & w3747) | (~w6100 & w4707) | (w3747 & w4707);
assign w4945 = (w2112 & w7558) | (w2112 & w2347) | (w7558 & w2347);
assign w4946 = (w1852 & w7517) | (w1852 & ~w6177) | (w7517 & ~w6177);
assign w4947 = ~w746 & ~w1733;
assign w4948 = (~w7026 & w2407) | (~w7026 & w5699) | (w2407 & w5699);
assign w4949 = (w6100 & w7229) | (w6100 & w1638) | (w7229 & w1638);
assign w4950 = ~w84 & w1326;
assign w4951 = w171 & ~w7352;
assign w4952 = (~w2627 & w6624) | (~w2627 & w4456) | (w6624 & w4456);
assign w4953 = w3924 & ~w4786;
assign w4954 = (~w2203 & w5297) | (~w2203 & w2420) | (w5297 & w2420);
assign w4955 = ~w2249 & ~w4151;
assign w4956 = ~w4415 & w4099;
assign w4957 = ~w5178 & w853;
assign w4958 = ~w2688 & ~w5699;
assign w4959 = w3466 & w5418;
assign w4960 = ~w1632 & ~w577;
assign w4961 = (w4680 & w5549) | (w4680 & ~w3770) | (w5549 & ~w3770);
assign w4962 = (w4969 & w919) | (w4969 & w6869) | (w919 & w6869);
assign w4963 = (~w1958 & w4511) | (~w1958 & w6256) | (w4511 & w6256);
assign w4964 = (~w2401 & w6852) | (~w2401 & w3139) | (w6852 & w3139);
assign w4965 = (~w5834 & w3996) | (~w5834 & w5825) | (w3996 & w5825);
assign w4966 = (w2452 & w5580) | (w2452 & w4351) | (w5580 & w4351);
assign w4967 = ~w4480 & w5223;
assign w4968 = (w632 & w5138) | (w632 & w260) | (w5138 & w260);
assign w4969 = (~w3490 & w7354) | (~w3490 & w1295) | (w7354 & w1295);
assign w4970 = ~w3052 & ~w7219;
assign w4971 = (~w6100 & w2878) | (~w6100 & w4658) | (w2878 & w4658);
assign w4972 = (~w5178 & w3338) | (~w5178 & w1989) | (w3338 & w1989);
assign w4973 = (w6385 & w6976) | (w6385 & w3819) | (w6976 & w3819);
assign w4974 = ~w3454 & ~w1375;
assign w4975 = ~w6162 & w7111;
assign w4976 = ~w7632 & ~w5077;
assign w4977 = w4843 & ~w1878;
assign w4978 = ~w4972 & ~w3881;
assign w4979 = (w5007 & w232) | (w5007 & w5990) | (w232 & w5990);
assign w4980 = (w7529 & w1659) | (w7529 & ~w491) | (w1659 & ~w491);
assign w4981 = (w6214 & w4773) | (w6214 & ~w343) | (w4773 & ~w343);
assign w4982 = (w1847 & w284) | (w1847 & w4519) | (w284 & w4519);
assign w4983 = (w6680 & w1046) | (w6680 & w4580) | (w1046 & w4580);
assign w4984 = (~w1709 & ~w671) | (~w1709 & w4162) | (~w671 & w4162);
assign w4985 = (w5921 & ~w5528) | (w5921 & w2468) | (~w5528 & w2468);
assign w4986 = (w6046 & w5217) | (w6046 & w3548) | (w5217 & w3548);
assign w4987 = ~a212 & ~b212;
assign w4988 = w5514 & w4607;
assign w4989 = ~w3570 & ~w5756;
assign w4990 = ~w2584 & w2844;
assign w4991 = ~w6206 & ~w5760;
assign w4992 = ~w26 & ~w5505;
assign w4993 = (~w7628 & w3846) | (~w7628 & w951) | (w3846 & w951);
assign w4994 = (~w6424 & w7244) | (~w6424 & w6165) | (w7244 & w6165);
assign w4995 = (~w2379 & w3646) | (~w2379 & w2522) | (w3646 & w2522);
assign w4996 = (w3929 & w1822) | (w3929 & w4354) | (w1822 & w4354);
assign w4997 = ~w7101 & w3213;
assign w4998 = w4238 & ~w2441;
assign w4999 = (~w2725 & w3224) | (~w2725 & w5678) | (w3224 & w5678);
assign w5000 = (~w5821 & w660) | (~w5821 & w2692) | (w660 & w2692);
assign w5001 = ~w5871 & w2894;
assign w5002 = w4206 & ~w2416;
assign w5003 = (~w5834 & w1249) | (~w5834 & w4734) | (w1249 & w4734);
assign w5004 = ~w1038 & w384;
assign w5005 = ~a94 & ~b94;
assign w5006 = (~w2456 & w6592) | (~w2456 & w558) | (w6592 & w558);
assign w5007 = ~w3119 & w5343;
assign w5008 = ~w5665 & ~w4632;
assign w5009 = ~w2735 & w4843;
assign w5010 = ~w6476 & ~w5355;
assign w5011 = (w264 & w4968) | (w264 & w2942) | (w4968 & w2942);
assign w5012 = ~w1736 & ~w1152;
assign w5013 = ~w2798 & ~w5376;
assign w5014 = (~w6516 & ~w3942) | (~w6516 & w5705) | (~w3942 & w5705);
assign w5015 = w3471 & ~w792;
assign w5016 = ~w4802 & w978;
assign w5017 = w1658 & ~w2040;
assign w5018 = (~w4118 & w4711) | (~w4118 & w1830) | (w4711 & w1830);
assign w5019 = (w5325 & w3940) | (w5325 & w4395) | (w3940 & w4395);
assign w5020 = w7294 & w7546;
assign w5021 = (~w6100 & w33) | (~w6100 & w4723) | (w33 & w4723);
assign w5022 = w1709 & w2110;
assign w5023 = (w7379 & w1933) | (w7379 & ~w4521) | (w1933 & ~w4521);
assign w5024 = w1395 & ~w1942;
assign w5025 = ~w3248 & ~w4074;
assign w5026 = w2622 & ~w868;
assign w5027 = (~w2021 & w2565) | (~w2021 & w7337) | (w2565 & w7337);
assign w5028 = (~w1228 & w6402) | (~w1228 & w6889) | (w6402 & w6889);
assign w5029 = (w3318 & w5081) | (w3318 & w6769) | (w5081 & w6769);
assign w5030 = (~w3774 & w2328) | (~w3774 & w3487) | (w2328 & w3487);
assign w5031 = (w3953 & w4945) | (w3953 & w1313) | (w4945 & w1313);
assign w5032 = ~w7527 & ~w4321;
assign w5033 = ~w5278 & w2887;
assign w5034 = w5036 & w7123;
assign w5035 = ~w5900 & ~w4457;
assign w5036 = ~w2260 & ~w335;
assign w5037 = (~w5522 & w759) | (~w5522 & w5397) | (w759 & w5397);
assign w5038 = (w7015 & w859) | (w7015 & w3970) | (w859 & w3970);
assign w5039 = ~w1073 & ~w4010;
assign w5040 = w1736 & ~w2725;
assign w5041 = (w3774 & w5064) | (w3774 & w4777) | (w5064 & w4777);
assign w5042 = w1204 & w3880;
assign w5043 = (w412 & w2904) | (w412 & w1027) | (w2904 & w1027);
assign w5044 = (w777 & w5324) | (w777 & w3233) | (w5324 & w3233);
assign w5045 = (~w6746 & w4536) | (~w6746 & w1116) | (w4536 & w1116);
assign w5046 = w51 & w389;
assign w5047 = (w1880 & w3641) | (w1880 & w5291) | (w3641 & w5291);
assign w5048 = (w3852 & w5644) | (w3852 & w3927) | (w5644 & w3927);
assign w5049 = ~w1579 & ~w4758;
assign w5050 = (~w2068 & w1660) | (~w2068 & w6495) | (w1660 & w6495);
assign w5051 = w2295 & ~w960;
assign w5052 = (w4864 & w4135) | (w4864 & ~w7383) | (w4135 & ~w7383);
assign w5053 = a83 & b83;
assign w5054 = ~w63 & ~w7622;
assign w5055 = (~w341 & w3350) | (~w341 & w2669) | (w3350 & w2669);
assign w5056 = ~w7289 & ~w2567;
assign w5057 = w5257 & w3024;
assign w5058 = (w2420 & ~w3819) | (w2420 & w3708) | (~w3819 & w3708);
assign w5059 = ~a214 & ~b214;
assign w5060 = (w2456 & w573) | (w2456 & w146) | (w573 & w146);
assign w5061 = (~w2456 & w1197) | (~w2456 & w2868) | (w1197 & w2868);
assign w5062 = ~w439 & ~w3845;
assign w5063 = (~w5424 & w394) | (~w5424 & w1314) | (w394 & w1314);
assign w5064 = w4777 | w949;
assign w5065 = (w1770 & w4259) | (w1770 & w848) | (w4259 & w848);
assign w5066 = ~w6656 & ~w5510;
assign w5067 = ~w2021 & w922;
assign w5068 = ~w4066 & w3123;
assign w5069 = ~w6210 & ~w2591;
assign w5070 = (w303 & w825) | (w303 & w2109) | (w825 & w2109);
assign w5071 = ~w4185 & w407;
assign w5072 = (~w4103 & ~w2979) | (~w4103 & ~w3318) | (~w2979 & ~w3318);
assign w5073 = w7439 & ~w4692;
assign w5074 = ~w1650 & ~w7422;
assign w5075 = ~w2182 & w1861;
assign w5076 = (~w5739 & ~w367) | (~w5739 & w6894) | (~w367 & w6894);
assign w5077 = ~w5005 & ~w6346;
assign w5078 = w5163 & w730;
assign w5079 = (~w303 & w6290) | (~w303 & w5906) | (w6290 & w5906);
assign w5080 = (~w5600 & ~w3011) | (~w5600 & w3949) | (~w3011 & w3949);
assign w5081 = (~w563 & w3671) | (~w563 & w2136) | (w3671 & w2136);
assign w5082 = (~w5834 & w256) | (~w5834 & w6908) | (w256 & w6908);
assign w5083 = (~w4132 & w3043) | (~w4132 & w128) | (w3043 & w128);
assign w5084 = (~w3852 & w225) | (~w3852 & w467) | (w225 & w467);
assign w5085 = (w7310 & w4434) | (w7310 & ~w6894) | (w4434 & ~w6894);
assign w5086 = w3066 & ~w7326;
assign w5087 = ~w4143 & w1278;
assign w5088 = (~w5995 & w7591) | (~w5995 & w3834) | (w7591 & w3834);
assign w5089 = w1868 & w6070;
assign w5090 = (w5141 & w1720) | (w5141 & w4227) | (w1720 & w4227);
assign w5091 = w2338 & w4638;
assign w5092 = (w5173 & w3562) | (w5173 & w5611) | (w3562 & w5611);
assign w5093 = w2354 & ~w6882;
assign w5094 = w330 & w4635;
assign w5095 = (~w5089 & w1487) | (~w5089 & w3175) | (w1487 & w3175);
assign w5096 = (w236 & w2373) | (w236 & w184) | (w2373 & w184);
assign w5097 = (w978 & w4007) | (w978 & w1503) | (w4007 & w1503);
assign w5098 = ~w6082 & ~w6254;
assign w5099 = (w6885 & w7058) | (w6885 & w6803) | (w7058 & w6803);
assign w5100 = (~w6100 & w6666) | (~w6100 & w3520) | (w6666 & w3520);
assign w5101 = ~w392 & ~w5932;
assign w5102 = w3933 & w6016;
assign w5103 = ~w5461 & ~w3425;
assign w5104 = ~w4412 & w1925;
assign w5105 = (~w5347 & w2237) | (~w5347 & w4600) | (w2237 & w4600);
assign w5106 = ~w4140 & ~w3990;
assign w5107 = ~w5998 & ~w1368;
assign w5108 = w2522 & w5061;
assign w5109 = ~w3312 & ~w7490;
assign w5110 = ~w2366 & ~w1273;
assign w5111 = ~w1656 & w6291;
assign w5112 = ~w1206 & ~w6281;
assign w5113 = w5042 & ~w400;
assign w5114 = w3231 & ~w3303;
assign w5115 = ~w5428 & ~w4474;
assign w5116 = (w7520 & w1963) | (w7520 & w166) | (w1963 & w166);
assign w5117 = ~w5400 & ~w374;
assign w5118 = ~w2914 & w4207;
assign w5119 = w3137 & ~w1901;
assign w5120 = ~w1786 & ~w42;
assign w5121 = ~w5350 & ~w6558;
assign w5122 = ~w698 & w1725;
assign w5123 = (~w6966 & w946) | (~w6966 & w6101) | (w946 & w6101);
assign w5124 = (~w1877 & w3461) | (~w1877 & w1803) | (w3461 & w1803);
assign w5125 = (~w1847 & w5134) | (~w1847 & w1465) | (w5134 & w1465);
assign w5126 = ~w3267 & ~w6112;
assign w5127 = w72 & ~w7576;
assign w5128 = ~w1588 & ~w5573;
assign w5129 = (~w3384 & ~w1675) | (~w3384 & ~w3533) | (~w1675 & ~w3533);
assign w5130 = (~w6647 & w4429) | (~w6647 & ~w1489) | (w4429 & ~w1489);
assign w5131 = (w7513 & w1372) | (w7513 & w3629) | (w1372 & w3629);
assign w5132 = (~w4995 & w6919) | (~w4995 & w1174) | (w6919 & w1174);
assign w5133 = (~w2065 & w3579) | (~w2065 & w5853) | (w3579 & w5853);
assign w5134 = (w735 & w5750) | (w735 & ~w6566) | (w5750 & ~w6566);
assign w5135 = w3032 & ~w5376;
assign w5136 = ~w1622 & ~w7365;
assign w5137 = (w303 & w1915) | (w303 & w2837) | (w1915 & w2837);
assign w5138 = w2740 & ~w4123;
assign w5139 = (w7126 & w5909) | (w7126 & ~w5395) | (w5909 & ~w5395);
assign w5140 = w5760 & w931;
assign w5141 = (~w1497 & w5475) | (~w1497 & w1607) | (w5475 & w1607);
assign w5142 = ~w5604 & w1085;
assign w5143 = ~w5782 & w1007;
assign w5144 = (w3119 & w6515) | (w3119 & w5530) | (w6515 & w5530);
assign w5145 = (w5178 & w4194) | (w5178 & w2398) | (w4194 & w2398);
assign w5146 = (w7239 & w5551) | (w7239 & w3063) | (w5551 & w3063);
assign w5147 = ~a12 & ~b12;
assign w5148 = w5191 & w7083;
assign w5149 = ~w84 & w2490;
assign w5150 = (~w412 & w6284) | (~w412 & w6613) | (w6284 & w6613);
assign w5151 = (~w4759 & w4458) | (~w4759 & ~w4768) | (w4458 & ~w4768);
assign w5152 = ~w7158 & ~w5756;
assign w5153 = ~w999 & ~w2959;
assign w5154 = (w5257 & w6223) | (w5257 & w1780) | (w6223 & w1780);
assign w5155 = (w4967 & w3951) | (w4967 & w1616) | (w3951 & w1616);
assign w5156 = (w5178 & w6735) | (w5178 & w6691) | (w6735 & w6691);
assign w5157 = (~w4143 & w6734) | (~w4143 & w1403) | (w6734 & w1403);
assign w5158 = (w4106 & w3148) | (w4106 & w4353) | (w3148 & w4353);
assign w5159 = (~w5703 & w5981) | (~w5703 & w2120) | (w5981 & w2120);
assign w5160 = (w3986 & w925) | (w3986 & w4634) | (w925 & w4634);
assign w5161 = w2820 | ~w1463;
assign w5162 = ~w1071 & ~w6592;
assign w5163 = ~w4140 & ~w4165;
assign w5164 = (w5083 & ~w2152) | (w5083 & ~w4138) | (~w2152 & ~w4138);
assign w5165 = (w5516 & w7398) | (w5516 & w7448) | (w7398 & w7448);
assign w5166 = ~w4710 & ~w6435;
assign w5167 = ~w1007 & w3805;
assign w5168 = (w3947 & w3115) | (w3947 & w2680) | (w3115 & w2680);
assign w5169 = ~w1024 & ~w7184;
assign w5170 = ~a197 & ~b197;
assign w5171 = (w6100 & w7182) | (w6100 & w5793) | (w7182 & w5793);
assign w5172 = ~w1360 & ~w4648;
assign w5173 = ~w6490 & ~w3538;
assign w5174 = w5732 & ~w7345;
assign w5175 = w2110 & ~w693;
assign w5176 = ~w1837 & ~w7632;
assign w5177 = w732 & w7375;
assign w5178 = (w5655 & w7297) | (w5655 & w2757) | (w7297 & w2757);
assign w5179 = w6198 | w1454;
assign w5180 = (~w5178 & w2748) | (~w5178 & w5754) | (w2748 & w5754);
assign w5181 = (~w1847 & w2732) | (~w1847 & w4495) | (w2732 & w4495);
assign w5182 = w7042 & ~w950;
assign w5183 = w7614 & ~w278;
assign w5184 = w4976 & ~w1760;
assign w5185 = w4257 & w1266;
assign w5186 = (w699 & w455) | (w699 & ~w4905) | (w455 & ~w4905);
assign w5187 = (w6460 & w4738) | (w6460 & w7238) | (w4738 & w7238);
assign w5188 = w701 & ~w4114;
assign w5189 = ~w4036 & ~w426;
assign w5190 = ~w2382 | ~w3264;
assign w5191 = w4347 & w5663;
assign w5192 = ~w561 & w3604;
assign w5193 = a65 & b65;
assign w5194 = ~w1972 & w1302;
assign w5195 = (w6100 & w1931) | (w6100 & w6076) | (w1931 & w6076);
assign w5196 = (w898 & w6286) | (w898 & w4199) | (w6286 & w4199);
assign w5197 = w666 & ~w5241;
assign w5198 = ~w2011 & w7312;
assign w5199 = w6304 & ~w6922;
assign w5200 = ~w2456 & w4660;
assign w5201 = w5948 & w7361;
assign w5202 = w1149 & ~w2619;
assign w5203 = ~w6082 & w1528;
assign w5204 = (w5522 & w7194) | (w5522 & w520) | (w7194 & w520);
assign w5205 = ~w6331 & ~w1556;
assign w5206 = ~w6818 & ~w5353;
assign w5207 = (w4702 & w6875) | (w4702 & ~w5403) | (w6875 & ~w5403);
assign w5208 = (~w907 & w3015) | (~w907 & w7252) | (w3015 & w7252);
assign w5209 = (w6512 & w4151) | (w6512 & ~w3894) | (w4151 & ~w3894);
assign w5210 = (w6754 & w2451) | (w6754 & ~w990) | (w2451 & ~w990);
assign w5211 = (w222 & w3461) | (w222 & w1951) | (w3461 & w1951);
assign w5212 = ~w1366 & ~w6336;
assign w5213 = ~w5180 & ~w560;
assign w5214 = ~w2615 & ~w3041;
assign w5215 = (~w3269 & w2049) | (~w3269 & w1886) | (w2049 & w1886);
assign w5216 = (w2871 & w2064) | (w2871 & w484) | (w2064 & w484);
assign w5217 = ~w6375 & ~w7581;
assign w5218 = (w4753 & w18) | (w4753 & ~w6501) | (w18 & ~w6501);
assign w5219 = ~w6753 & w4123;
assign w5220 = ~w6640 & w6100;
assign w5221 = (w4560 & w5107) | (w4560 & w3391) | (w5107 & w3391);
assign w5222 = w7183 & ~w3019;
assign w5223 = ~w2172 & w4211;
assign w5224 = (~w3057 & w6261) | (~w3057 & w2250) | (w6261 & w2250);
assign w5225 = (w4802 & w4680) | (w4802 & w5631) | (w4680 & w5631);
assign w5226 = ~w4366 & ~w6571;
assign w5227 = (w4145 & w480) | (w4145 & w4730) | (w480 & w4730);
assign w5228 = w2176 & w5947;
assign w5229 = w6804 & ~w1281;
assign w5230 = a54 & b54;
assign w5231 = w7599 & ~w3736;
assign w5232 = (~w6744 & w4743) | (~w6744 & w2437) | (w4743 & w2437);
assign w5233 = ~w5721 & ~w4620;
assign w5234 = ~w1954 & ~w6191;
assign w5235 = (~w3057 & w1298) | (~w3057 & w7224) | (w1298 & w7224);
assign w5236 = ~w1601 & ~w7644;
assign w5237 = (~w3774 & w6489) | (~w3774 & w2771) | (w6489 & w2771);
assign w5238 = w3161 & w6894;
assign w5239 = ~a144 & ~b144;
assign w5240 = ~w4881 & ~w7352;
assign w5241 = a234 & b234;
assign w5242 = a247 & b247;
assign w5243 = (~w3741 & w1077) | (~w3741 & w6100) | (w1077 & w6100);
assign w5244 = ~w2838 & w3841;
assign w5245 = (~w3119 & w3940) | (~w3119 & w2016) | (w3940 & w2016);
assign w5246 = ~w1999 & w1954;
assign w5247 = (w3330 & w4720) | (w3330 & w6428) | (w4720 & w6428);
assign w5248 = ~w5772 & w75;
assign w5249 = w634 & ~w215;
assign w5250 = ~w1002 & ~w5966;
assign w5251 = a131 & b131;
assign w5252 = (w5879 & w2708) | (w5879 & w5253) | (w2708 & w5253);
assign w5253 = ~w601 & w5879;
assign w5254 = ~w3951 & w681;
assign w5255 = w6517 & w1334;
assign w5256 = ~w6488 & ~w1896;
assign w5257 = (~w3774 & w5135) | (~w3774 & w6078) | (w5135 & w6078);
assign w5258 = (w173 & w2857) | (w173 & w108) | (w2857 & w108);
assign w5259 = w400 & ~w4494;
assign w5260 = ~w7278 & w5777;
assign w5261 = (~w2103 & w7245) | (~w2103 & w1099) | (w7245 & w1099);
assign w5262 = w1615 & ~w2707;
assign w5263 = w1532 & ~w5743;
assign w5264 = (w3200 & w2603) | (w3200 & w4721) | (w2603 & w4721);
assign w5265 = (w4143 & w6018) | (w4143 & w2704) | (w6018 & w2704);
assign w5266 = ~w1622 & w1804;
assign w5267 = ~w434 & ~w4742;
assign w5268 = (w3311 & w4423) | (w3311 & w5821) | (w4423 & w5821);
assign w5269 = (~w3869 & w2621) | (~w3869 & w2963) | (w2621 & w2963);
assign w5270 = w3824 & w2300;
assign w5271 = (w4296 & w1801) | (w4296 & w655) | (w1801 & w655);
assign w5272 = w1455 & w7082;
assign w5273 = ~w4587 & ~w505;
assign w5274 = (~w3318 & w5524) | (~w3318 & w2608) | (w5524 & w2608);
assign w5275 = ~w471 & w5230;
assign w5276 = a101 & b101;
assign w5277 = ~w3934 & ~w6520;
assign w5278 = (w5834 & w771) | (w5834 & w3780) | (w771 & w3780);
assign w5279 = w6979 & ~w216;
assign w5280 = (~w5007 & w3438) | (~w5007 & w5953) | (w3438 & w5953);
assign w5281 = (w4843 & ~w5259) | (w4843 & w4585) | (~w5259 & w4585);
assign w5282 = ~w5965 & w5032;
assign w5283 = (~w563 & w4244) | (~w563 & w2149) | (w4244 & w2149);
assign w5284 = ~w7528 & w2464;
assign w5285 = w3618 & ~w4409;
assign w5286 = w1716 & ~w780;
assign w5287 = a155 & b155;
assign w5288 = ~w7513 & w3240;
assign w5289 = a92 & b92;
assign w5290 = w3117 & ~w5528;
assign w5291 = (w2928 & ~w6680) | (w2928 & w4575) | (~w6680 & w4575);
assign w5292 = ~w7026 & w2612;
assign w5293 = ~w1069 & ~w5457;
assign w5294 = w1364 & ~w5836;
assign w5295 = a8 & b8;
assign w5296 = ~w6980 & ~w2611;
assign w5297 = w4236 & ~w2203;
assign w5298 = ~w4203 & w5745;
assign w5299 = w5519 & ~w1381;
assign w5300 = ~w3040 & w2668;
assign w5301 = (~w3267 & w2124) | (~w3267 & w1412) | (w2124 & w1412);
assign w5302 = w3894 & w2545;
assign w5303 = w5381 & w2218;
assign w5304 = (~w3888 & ~w1903) | (~w3888 & ~w343) | (~w1903 & ~w343);
assign w5305 = ~w1999 & ~w7563;
assign w5306 = (w1474 & w2847) | (w1474 & ~w5296) | (w2847 & ~w5296);
assign w5307 = w330 & ~w1165;
assign w5308 = (w3774 & w3412) | (w3774 & w1048) | (w3412 & w1048);
assign w5309 = (~w4840 & w11) | (~w4840 & w5671) | (w11 & w5671);
assign w5310 = ~w3933 & ~w6016;
assign w5311 = (~w732 & w1647) | (~w732 & w2772) | (w1647 & w2772);
assign w5312 = ~w5818 & w3060;
assign w5313 = (w5462 & w5790) | (w5462 & w2097) | (w5790 & w2097);
assign w5314 = ~w4833 & ~w4685;
assign w5315 = (w2660 & w5661) | (w2660 & ~w3883) | (w5661 & ~w3883);
assign w5316 = (~w2353 & w7397) | (~w2353 & w7049) | (w7397 & w7049);
assign w5317 = w2420 & w6397;
assign w5318 = (w7449 & w6118) | (w7449 & w5439) | (w6118 & w5439);
assign w5319 = (w306 & w4664) | (w306 & ~w5403) | (w4664 & ~w5403);
assign w5320 = (w4966 & w4447) | (w4966 & w5210) | (w4447 & w5210);
assign w5321 = (~w4499 & w3145) | (~w4499 & w6385) | (w3145 & w6385);
assign w5322 = (~w7552 & w1042) | (~w7552 & w4323) | (w1042 & w4323);
assign w5323 = w814 & w4597;
assign w5324 = ~w3066 & w7326;
assign w5325 = ~w5871 & w5403;
assign w5326 = (~w4906 & ~w1497) | (~w4906 & w4461) | (~w1497 & w4461);
assign w5327 = (w5422 & w3617) | (w5422 & ~w5098) | (w3617 & ~w5098);
assign w5328 = ~w7352 & w5860;
assign w5329 = w3580 & ~w757;
assign w5330 = w7137 & ~w968;
assign w5331 = (~w6184 & w5403) | (~w6184 & w4812) | (w5403 & w4812);
assign w5332 = (w6942 & w6148) | (w6942 & w1096) | (w6148 & w1096);
assign w5333 = ~w3389 & w3393;
assign w5334 = ~w302 & ~w14;
assign w5335 = (w1167 & w3296) | (w1167 & w5325) | (w3296 & w5325);
assign w5336 = w3105 & ~w5328;
assign w5337 = w1211 & w7275;
assign w5338 = (~w3269 & w2049) | (~w3269 & w491) | (w2049 & w491);
assign w5339 = (w3733 & w3154) | (w3733 & w1730) | (w3154 & w1730);
assign w5340 = w7647 & w6254;
assign w5341 = ~w2230 & ~w4333;
assign w5342 = (~w2627 & w2054) | (~w2627 & w1056) | (w2054 & w1056);
assign w5343 = ~w2456 & w6536;
assign w5344 = (w1367 & w1829) | (w1367 & w7132) | (w1829 & w7132);
assign w5345 = ~w4616 & ~w971;
assign w5346 = ~w1541 & w245;
assign w5347 = (w6100 & w3778) | (w6100 & w2780) | (w3778 & w2780);
assign w5348 = a144 & b144;
assign w5349 = ~w336 & ~w5193;
assign w5350 = ~a142 & ~b142;
assign w5351 = ~w1877 & ~w2483;
assign w5352 = w3473 & w7539;
assign w5353 = (w3661 & w2955) | (w3661 & w5655) | (w2955 & w5655);
assign w5354 = (w5178 & w4979) | (w5178 & w2675) | (w4979 & w2675);
assign w5355 = (w5655 & w7001) | (w5655 & w5168) | (w7001 & w5168);
assign w5356 = (w6894 & w4233) | (w6894 & w4955) | (w4233 & w4955);
assign w5357 = (w3984 & w531) | (w3984 & w5679) | (w531 & w5679);
assign w5358 = ~w3636 & w3104;
assign w5359 = (w3774 & w2537) | (w3774 & w1246) | (w2537 & w1246);
assign w5360 = w5787 & ~w614;
assign w5361 = ~w1661 & ~w3172;
assign w5362 = ~w7397 & w7078;
assign w5363 = (w978 & w199) | (w978 & w3090) | (w199 & w3090);
assign w5364 = w2243 & ~w5053;
assign w5365 = w2655 & w1608;
assign w5366 = ~w5373 & w6317;
assign w5367 = w3102 & w5871;
assign w5368 = ~w4004 & w2855;
assign w5369 = (w5403 & w3768) | (w5403 & w4812) | (w3768 & w4812);
assign w5370 = ~w3312 & ~w624;
assign w5371 = ~w1903 | ~w3888;
assign w5372 = (w2334 & w5498) | (w2334 & w6254) | (w5498 & w6254);
assign w5373 = w2799 & ~w4083;
assign w5374 = ~w6255 & w6716;
assign w5375 = (w6359 & w1453) | (w6359 & w7108) | (w1453 & w7108);
assign w5376 = w944 & ~w7321;
assign w5377 = (w6082 & w4629) | (w6082 & w1186) | (w4629 & w1186);
assign w5378 = (~w5291 & w7176) | (~w5291 & w2583) | (w7176 & w2583);
assign w5379 = ~w2513 & ~w4675;
assign w5380 = ~w2452 & w6777;
assign w5381 = w3426 & w3016;
assign w5382 = w486 & w511;
assign w5383 = ~w5809 & ~w6703;
assign w5384 = ~w1632 & w7648;
assign w5385 = w174 & ~w1607;
assign w5386 = (w4440 & w5593) | (w4440 & w5871) | (w5593 & w5871);
assign w5387 = (w2966 & w3221) | (w2966 & w2153) | (w3221 & w2153);
assign w5388 = w668 & w3188;
assign w5389 = ~w1377 & w4012;
assign w5390 = (w6418 & w5529) | (w6418 & w6620) | (w5529 & w6620);
assign w5391 = ~w2343 & w6385;
assign w5392 = ~w4508 & ~w3007;
assign w5393 = ~w4837 & ~w2801;
assign w5394 = w2094 & w4613;
assign w5395 = (w2429 & w1516) | (w2429 & w3852) | (w1516 & w3852);
assign w5396 = (w6534 & w4469) | (w6534 & w4143) | (w4469 & w4143);
assign w5397 = ~w6608 & w4768;
assign w5398 = ~w6983 & w4768;
assign w5399 = ~w6992 & w4012;
assign w5400 = (~w5178 & w7501) | (~w5178 & w6938) | (w7501 & w6938);
assign w5401 = w7526 & w274;
assign w5402 = w5809 & ~w5389;
assign w5403 = ~w2847 & w308;
assign w5404 = ~w5573 & ~w2202;
assign w5405 = (w5537 & w1500) | (w5537 & ~w6174) | (w1500 & ~w6174);
assign w5406 = ~w4496 & ~w6504;
assign w5407 = (w3983 & w5644) | (w3983 & w3927) | (w5644 & w3927);
assign w5408 = w2981 & w2833;
assign w5409 = ~w4991 & ~w5584;
assign w5410 = (~w1158 & w6299) | (~w1158 & ~w3888) | (w6299 & ~w3888);
assign w5411 = ~w2255 & ~w5830;
assign w5412 = ~w2119 & ~w3427;
assign w5413 = (w1369 & w2362) | (w1369 & ~w1315) | (w2362 & ~w1315);
assign w5414 = ~w4206 & w2222;
assign w5415 = (w861 & ~w3819) | (w861 & w3884) | (~w3819 & w3884);
assign w5416 = ~a186 & ~b186;
assign w5417 = w3119 & ~w5325;
assign w5418 = w1221 & ~w7202;
assign w5419 = ~w3168 & w6849;
assign w5420 = (w6082 & w3498) | (w6082 & w2162) | (w3498 & w2162);
assign w5421 = ~w2996 & w1479;
assign w5422 = (w6353 & w1139) | (w6353 & w2132) | (w1139 & w2132);
assign w5423 = ~w1443 & ~w2632;
assign w5424 = ~w2984 & ~w1938;
assign w5425 = a67 & b67;
assign w5426 = (~w7554 & w866) | (~w7554 & w5651) | (w866 & w5651);
assign w5427 = (~w6451 & w1826) | (~w6451 & ~w697) | (w1826 & ~w697);
assign w5428 = ~w516 & w2244;
assign w5429 = w813 & ~w898;
assign w5430 = w6566 & ~w6013;
assign w5431 = ~w301 & ~w893;
assign w5432 = (~w7581 & ~w4027) | (~w7581 & w6866) | (~w4027 & w6866);
assign w5433 = (w5257 & w3189) | (w5257 & w6295) | (w3189 & w6295);
assign w5434 = (w6127 & w5483) | (w6127 & w3448) | (w5483 & w3448);
assign w5435 = ~w6046 & w4708;
assign w5436 = ~w1846 & ~w1252;
assign w5437 = ~w336 & ~w957;
assign w5438 = w457 & ~w3503;
assign w5439 = (w5596 & ~w2335) | (w5596 & w6072) | (~w2335 & w6072);
assign w5440 = w1577 & ~w3375;
assign w5441 = (w7566 & w1565) | (w7566 & w298) | (w1565 & w298);
assign w5442 = a33 & b33;
assign w5443 = (w3423 & w4750) | (w3423 & w2275) | (w4750 & w2275);
assign w5444 = ~w5664 & ~w4241;
assign w5445 = ~w4987 & ~w561;
assign w5446 = w2875 & ~w2563;
assign w5447 = w5032 & ~w7549;
assign w5448 = (~w236 & w2200) | (~w236 & w3676) | (w2200 & w3676);
assign w5449 = ~w1204 & w2068;
assign w5450 = ~w4706 & ~w3673;
assign w5451 = (w5834 & w3566) | (w5834 & w849) | (w3566 & w849);
assign w5452 = w4479 & w875;
assign w5453 = ~w1026 & ~w2644;
assign w5454 = w7647 & w4299;
assign w5455 = (w2627 & w1771) | (w2627 & w1619) | (w1771 & w1619);
assign w5456 = w4808 & ~w1135;
assign w5457 = (~w2627 & w4463) | (~w2627 & w7499) | (w4463 & w7499);
assign w5458 = (w3057 & w623) | (w3057 & w7285) | (w623 & w7285);
assign w5459 = (~w7491 & w479) | (~w7491 & w867) | (w479 & w867);
assign w5460 = (~w6524 & w663) | (~w6524 & w3771) | (w663 & w3771);
assign w5461 = ~w7486 & ~w878;
assign w5462 = w2869 & ~w2890;
assign w5463 = a132 & b132;
assign w5464 = ~a74 & ~b74;
assign w5465 = ~w781 & ~w7115;
assign w5466 = a163 & b163;
assign w5467 = a125 & b125;
assign w5468 = w5065 & w2627;
assign w5469 = ~w4680 & w2107;
assign w5470 = (w5871 & w3891) | (w5871 & w6302) | (w3891 & w6302);
assign w5471 = (w3057 & w1779) | (w3057 & w4360) | (w1779 & w4360);
assign w5472 = ~w395 & ~w5003;
assign w5473 = (w1254 & ~w7197) | (w1254 & w1190) | (~w7197 & w1190);
assign w5474 = ~w7158 & ~w2744;
assign w5475 = (w3212 & ~w3070) | (w3212 & ~w6614) | (~w3070 & ~w6614);
assign w5476 = ~w3855 & ~w4745;
assign w5477 = w2027 & ~w4169;
assign w5478 = ~w727 & ~w351;
assign w5479 = (w1212 & ~w3119) | (w1212 & w3025) | (~w3119 & w3025);
assign w5480 = ~a125 & ~b125;
assign w5481 = w4496 & w1544;
assign w5482 = w4768 & ~w7391;
assign w5483 = w2471 & ~w195;
assign w5484 = ~w2847 & w1315;
assign w5485 = w6785 & ~w2671;
assign w5486 = w2996 & ~w5808;
assign w5487 = ~w6757 & ~w6016;
assign w5488 = (~w6911 & w6271) | (~w6911 & ~w5304) | (w6271 & ~w5304);
assign w5489 = ~w314 & w4230;
assign w5490 = ~w4833 & w5361;
assign w5491 = (~w6162 & w6117) | (~w6162 & w7173) | (w6117 & w7173);
assign w5492 = w5948 & w4977;
assign w5493 = (~w1925 & w1731) | (~w1925 & w1377) | (w1731 & w1377);
assign w5494 = (w3709 & w1506) | (w3709 & ~w2835) | (w1506 & ~w2835);
assign w5495 = (~w3892 & w2167) | (~w3892 & w7557) | (w2167 & w7557);
assign w5496 = w6656 & ~w2567;
assign w5497 = w1492 & ~w2892;
assign w5498 = ~w4505 & ~w2797;
assign w5499 = a138 & b138;
assign w5500 = (w5554 & w1229) | (w5554 & w7043) | (w1229 & w7043);
assign w5501 = (w2354 & w5995) | (w2354 & w1521) | (w5995 & w1521);
assign w5502 = (w3647 & w4897) | (w3647 & ~w3533) | (w4897 & ~w3533);
assign w5503 = ~w5059 & ~w4275;
assign w5504 = w2005 & ~w1427;
assign w5505 = (w5178 & w988) | (w5178 & w6405) | (w988 & w6405);
assign w5506 = (w2052 & w4444) | (w2052 & w3067) | (w4444 & w3067);
assign w5507 = w6503 & w2333;
assign w5508 = (w1794 & w1039) | (w1794 & w4258) | (w1039 & w4258);
assign w5509 = (w6475 & w1064) | (w6475 & w6100) | (w1064 & w6100);
assign w5510 = a235 & b235;
assign w5511 = (w3057 & w6453) | (w3057 & w4281) | (w6453 & w4281);
assign w5512 = ~w7365 & ~w6564;
assign w5513 = (w4995 & w2794) | (w4995 & w3610) | (w2794 & w3610);
assign w5514 = ~w7425 & ~w5577;
assign w5515 = (~w3318 & w6726) | (~w3318 & w130) | (w6726 & w130);
assign w5516 = ~w2452 & w4488;
assign w5517 = (w5411 & w3892) | (w5411 & w880) | (w3892 & w880);
assign w5518 = (w6738 & w4985) | (w6738 & w7431) | (w4985 & w7431);
assign w5519 = ~w990 & w5453;
assign w5520 = w1570 & w3728;
assign w5521 = w6646 | w1150;
assign w5522 = w7243 & ~w3292;
assign w5523 = w3901 & w4764;
assign w5524 = (w6664 & w1646) | (w6664 & w563) | (w1646 & w563);
assign w5525 = a212 & b212;
assign w5526 = (w3989 & ~w4182) | (w3989 & w1264) | (~w4182 & w1264);
assign w5527 = (w1834 & w7225) | (w1834 & w4867) | (w7225 & w4867);
assign w5528 = (w3473 & w4287) | (w3473 & w159) | (w4287 & w159);
assign w5529 = w6620 & ~w6100;
assign w5530 = (w4836 & w1689) | (w4836 & ~w5403) | (w1689 & ~w5403);
assign w5531 = (w2534 & w6311) | (w2534 & ~w6504) | (w6311 & ~w6504);
assign w5532 = w6244 & w5576;
assign w5533 = (~w6467 & w1090) | (~w6467 & w5623) | (w1090 & w5623);
assign w5534 = w4130 & w7354;
assign w5535 = w4914 & w90;
assign w5536 = w3231 & w7450;
assign w5537 = ~w1565 & w6430;
assign w5538 = w1783 & w4154;
assign w5539 = (w5178 & w953) | (w5178 & w3926) | (w953 & w3926);
assign w5540 = w6151 & w6606;
assign w5541 = w6490 & ~w2613;
assign w5542 = (~w2041 & w7093) | (~w2041 & w1171) | (w7093 & w1171);
assign w5543 = w6811 & ~w7564;
assign w5544 = w4444 & ~w6889;
assign w5545 = (w2083 & w4424) | (w2083 & w5410) | (w4424 & w5410);
assign w5546 = (w7273 & w3755) | (w7273 & w7113) | (w3755 & w7113);
assign w5547 = ~w2123 & w4110;
assign w5548 = w43 & w6100;
assign w5549 = w4504 | w4468;
assign w5550 = w6002 & ~w6963;
assign w5551 = (~w5516 & w4234) | (~w5516 & w7239) | (w4234 & w7239);
assign w5552 = (w3823 & w5089) | (w3823 & w27) | (w5089 & w27);
assign w5553 = w3551 & ~w4651;
assign w5554 = w7577 & ~w3123;
assign w5555 = w2644 & ~w5570;
assign w5556 = ~w3692 & ~w5499;
assign w5557 = ~a233 & ~b233;
assign w5558 = ~w1899 & ~w5630;
assign w5559 = ~w4448 & w7491;
assign w5560 = w3312 & ~w5230;
assign w5561 = w5464 & ~w625;
assign w5562 = w7060 | w3863;
assign w5563 = (w5298 & w6052) | (w5298 & w2524) | (w6052 & w2524);
assign w5564 = (~w6184 & w84) | (~w6184 & w3094) | (w84 & w3094);
assign w5565 = ~w693 & ~w6239;
assign w5566 = (~w6100 & w709) | (~w6100 & w6363) | (w709 & w6363);
assign w5567 = (~w2353 & w4967) | (~w2353 & w5316) | (w4967 & w5316);
assign w5568 = ~w3782 & ~w3730;
assign w5569 = ~w1812 & w7576;
assign w5570 = a74 & b74;
assign w5571 = w7632 & ~w4242;
assign w5572 = ~w478 & w3644;
assign w5573 = a122 & b122;
assign w5574 = (w2969 & w2003) | (w2969 & ~w6100) | (w2003 & ~w6100);
assign w5575 = (~w2453 & w58) | (~w2453 & w2133) | (w58 & w2133);
assign w5576 = (~w2718 & ~w1195) | (~w2718 & w7178) | (~w1195 & w7178);
assign w5577 = ~w6448 & w6522;
assign w5578 = (w6680 & w4696) | (w6680 & w5395) | (w4696 & w5395);
assign w5579 = (w7187 & w6125) | (w7187 & w1760) | (w6125 & w1760);
assign w5580 = ~w5194 | w4149;
assign w5581 = ~w5983 & ~w7572;
assign w5582 = w3092 & ~w812;
assign w5583 = (~w3847 & w482) | (~w3847 & w6431) | (w482 & w6431);
assign w5584 = (~w5257 & w2356) | (~w5257 & w4219) | (w2356 & w4219);
assign w5585 = ~w3701 & w1555;
assign w5586 = w5127 & ~w2935;
assign w5587 = w6524 & w1511;
assign w5588 = ~a156 & ~b156;
assign w5589 = w1241 & w3066;
assign w5590 = (w554 & ~w7526) | (w554 & w507) | (~w7526 & w507);
assign w5591 = (w5022 & w420) | (w5022 & w6831) | (w420 & w6831);
assign w5592 = (~w3737 & w2541) | (~w3737 & w844) | (w2541 & w844);
assign w5593 = ~w3677 & ~w1134;
assign w5594 = w569 & ~w4169;
assign w5595 = w719 & ~w4132;
assign w5596 = ~w3631 & w1004;
assign w5597 = w7188 & w1429;
assign w5598 = ~a45 & ~b45;
assign w5599 = ~a251 & ~b251;
assign w5600 = w3064 & ~w2243;
assign w5601 = (~w3612 & w276) | (~w3612 & w3119) | (w276 & w3119);
assign w5602 = w4180 & w6712;
assign w5603 = w2255 & w6644;
assign w5604 = ~w1601 & ~w7373;
assign w5605 = (w3318 & w3759) | (w3318 & w3740) | (w3759 & w3740);
assign w5606 = (~w523 & w1456) | (~w523 & ~w2104) | (w1456 & ~w2104);
assign w5607 = (w6467 & w5867) | (w6467 & w3944) | (w5867 & w3944);
assign w5608 = ~w106 & w7218;
assign w5609 = (~w7256 & w156) | (~w7256 & ~w3246) | (w156 & ~w3246);
assign w5610 = (w3733 & w3154) | (w3733 & w2876) | (w3154 & w2876);
assign w5611 = ~w6082 & w6384;
assign w5612 = (w5178 & w3897) | (w5178 & w1971) | (w3897 & w1971);
assign w5613 = (w5178 & w4693) | (w5178 & w1362) | (w4693 & w1362);
assign w5614 = w1696 & w702;
assign w5615 = ~w1274 & ~w6146;
assign w5616 = a99 & b99;
assign w5617 = w7365 & ~w5777;
assign w5618 = (~w5296 & w1373) | (~w5296 & w220) | (w1373 & w220);
assign w5619 = w4610 & ~w2080;
assign w5620 = (~w6984 & ~w441) | (~w6984 & w1965) | (~w441 & w1965);
assign w5621 = w4706 & w4897;
assign w5622 = ~a47 & ~b47;
assign w5623 = (w6151 & w570) | (w6151 & w4512) | (w570 & w4512);
assign w5624 = w4282 & w1641;
assign w5625 = (w544 & w3802) | (w544 & w6144) | (w3802 & w6144);
assign w5626 = (w2842 & w7331) | (w2842 & ~w1730) | (w7331 & ~w1730);
assign w5627 = ~w1660 & w497;
assign w5628 = ~w2735 & w3482;
assign w5629 = ~w5951 & w1735;
assign w5630 = ~w3099 & w7185;
assign w5631 = ~w2107 & w4802;
assign w5632 = (~w7552 & w1042) | (~w7552 & w6120) | (w1042 & w6120);
assign w5633 = ~w3869 & ~w5599;
assign w5634 = w7058 & w6885;
assign w5635 = w7390 & ~w7546;
assign w5636 = ~w2838 & ~w385;
assign w5637 = ~w4747 & w5659;
assign w5638 = (w1548 & w7220) | (w1548 & ~w1881) | (w7220 & ~w1881);
assign w5639 = w7327 | w1715;
assign w5640 = ~w7564 & w1145;
assign w5641 = ~w5808 & ~w2127;
assign w5642 = (w3063 & w3406) | (w3063 & w800) | (w3406 & w800);
assign w5643 = ~w5510 & w5056;
assign w5644 = ~w3573 & w1532;
assign w5645 = w1635 & ~w1656;
assign w5646 = ~w3217 & ~w625;
assign w5647 = ~w6909 & ~w4581;
assign w5648 = (w1751 & w1102) | (w1751 & w7353) | (w1102 & w7353);
assign w5649 = w2566 & ~w6705;
assign w5650 = (w5895 & w1908) | (w5895 & ~w5403) | (w1908 & ~w5403);
assign w5651 = (~w7350 & w2533) | (~w7350 & ~w6099) | (w2533 & ~w6099);
assign w5652 = ~w7183 & ~w429;
assign w5653 = ~w1772 & ~w6289;
assign w5654 = (~w1851 & w675) | (~w1851 & w957) | (w675 & w957);
assign w5655 = (w5098 & ~w6100) | (w5098 & w6174) | (~w6100 & w6174);
assign w5656 = w7131 | w3939;
assign w5657 = w4043 & ~w486;
assign w5658 = w5883 & ~w6979;
assign w5659 = ~w3167 & w5008;
assign w5660 = (~w6100 & w2934) | (~w6100 & w1600) | (w2934 & w1600);
assign w5661 = (w478 & w2660) | (w478 & w7235) | (w2660 & w7235);
assign w5662 = w5797 & w193;
assign w5663 = w4237 & w6802;
assign w5664 = (w3318 & w377) | (w3318 & w3012) | (w377 & w3012);
assign w5665 = ~a7 & ~b7;
assign w5666 = ~w2261 & w3319;
assign w5667 = (w4726 & w19) | (w4726 & ~w4867) | (w19 & ~w4867);
assign w5668 = (w1767 & w6262) | (w1767 & w2870) | (w6262 & w2870);
assign w5669 = ~w4749 & ~w4875;
assign w5670 = (w2837 & w1915) | (w2837 & w794) | (w1915 & w794);
assign w5671 = ~w6870 & ~w3492;
assign w5672 = (w6504 & w1611) | (w6504 & w2966) | (w1611 & w2966);
assign w5673 = (w6100 & w4501) | (w6100 & w7050) | (w4501 & w7050);
assign w5674 = (w506 & w2425) | (w506 & w4054) | (w2425 & w4054);
assign w5675 = w1483 & ~w5153;
assign w5676 = a152 & b152;
assign w5677 = (~w3636 & w4087) | (~w3636 & w176) | (w4087 & w176);
assign w5678 = (~w2725 & w1736) | (~w2725 & ~w3014) | (w1736 & ~w3014);
assign w5679 = ~w3096 & w5635;
assign w5680 = ~w3444 & w6100;
assign w5681 = ~w5782 & ~w142;
assign w5682 = (w4143 & w3723) | (w4143 & w4248) | (w3723 & w4248);
assign w5683 = ~w2027 & ~w6804;
assign w5684 = (w3831 & w233) | (w3831 & ~w1628) | (w233 & ~w1628);
assign w5685 = w6991 & ~w2728;
assign w5686 = ~w736 & ~w7452;
assign w5687 = ~a90 & ~b90;
assign w5688 = (~w3503 & w457) | (~w3503 & w3290) | (w457 & w3290);
assign w5689 = w2540 & ~w7454;
assign w5690 = (w3848 & w2263) | (w3848 & ~w5526) | (w2263 & ~w5526);
assign w5691 = ~w4027 & w2514;
assign w5692 = ~w6682 | ~w7567;
assign w5693 = a112 & b112;
assign w5694 = ~w5281 & ~w226;
assign w5695 = (w3708 & w4954) | (w3708 & w6109) | (w4954 & w6109);
assign w5696 = ~w4605 & w838;
assign w5697 = (~w3892 & w1612) | (~w3892 & w5700) | (w1612 & w5700);
assign w5698 = w4149 & ~w2644;
assign w5699 = w3019 & ~w7026;
assign w5700 = (~w3113 & w1663) | (~w3113 & w1649) | (w1663 & w1649);
assign w5701 = w4833 & w4685;
assign w5702 = (~w671 & w753) | (~w671 & w5141) | (w753 & w5141);
assign w5703 = (w3318 & w6227) | (w3318 & w7155) | (w6227 & w7155);
assign w5704 = (~w867 & w529) | (~w867 & w6012) | (w529 & w6012);
assign w5705 = w471 & ~w6516;
assign w5706 = ~w2838 & w5636;
assign w5707 = (w6738 & w896) | (w6738 & w5667) | (w896 & w5667);
assign w5708 = w6452 & w7;
assign w5709 = (w1863 & w2726) | (w1863 & w6254) | (w2726 & w6254);
assign w5710 = w5068 & ~w4066;
assign w5711 = (~w788 & w4567) | (~w788 & w5194) | (w4567 & w5194);
assign w5712 = (w5699 & w4948) | (w5699 & w3819) | (w4948 & w3819);
assign w5713 = w5199 & ~w6922;
assign w5714 = ~w3888 & w949;
assign w5715 = ~w2947 & ~w6279;
assign w5716 = (w6140 & w4410) | (w6140 & w3819) | (w4410 & w3819);
assign w5717 = (~w5813 & w2037) | (~w5813 & w3662) | (w2037 & w3662);
assign w5718 = w3665 & w3083;
assign w5719 = ~w6035 & ~w5673;
assign w5720 = (~w2548 & w2097) | (~w2548 & w2073) | (w2097 & w2073);
assign w5721 = ~w1866 & ~w6243;
assign w5722 = w6452 & ~w1655;
assign w5723 = ~w3818 & ~w7627;
assign w5724 = (w924 & w5771) | (w924 & w4886) | (w5771 & w4886);
assign w5725 = w6754 & ~w6844;
assign w5726 = ~w2741 & w483;
assign w5727 = (~w5066 & w2178) | (~w5066 & w3953) | (w2178 & w3953);
assign w5728 = w4684 & w6833;
assign w5729 = w1271 & w612;
assign w5730 = ~w1932 & ~w584;
assign w5731 = ~w4870 & ~w538;
assign w5732 = ~a228 & ~b228;
assign w5733 = ~w5171 & ~w3372;
assign w5734 = ~w2847 & w6108;
assign w5735 = w1743 & w1814;
assign w5736 = ~w6164 & ~w4952;
assign w5737 = ~w1582 & ~w3904;
assign w5738 = w3896 & ~w7291;
assign w5739 = (w52 & w3953) | (w52 & w6746) | (w3953 & w6746);
assign w5740 = ~w3057 & w5595;
assign w5741 = (w5178 & w402) | (w5178 & w59) | (w402 & w59);
assign w5742 = (w6100 & w6159) | (w6100 & w6978) | (w6159 & w6978);
assign w5743 = ~a29 & ~b29;
assign w5744 = ~w1756 & w5998;
assign w5745 = a246 & b246;
assign w5746 = (w1611 & w7324) | (w1611 & w4367) | (w7324 & w4367);
assign w5747 = w5385 & w5749;
assign w5748 = ~w2853 & w6571;
assign w5749 = w4132 & ~w3304;
assign w5750 = (~w6517 & w735) | (~w6517 & w443) | (w735 & w443);
assign w5751 = ~w6104 & ~w3618;
assign w5752 = w5205 & w909;
assign w5753 = (w5298 & w6052) | (w5298 & ~w2097) | (w6052 & ~w2097);
assign w5754 = (w6467 & w2748) | (w6467 & w3081) | (w2748 & w3081);
assign w5755 = (w2177 & w3601) | (w2177 & w4591) | (w3601 & w4591);
assign w5756 = ~w7622 & ~w4403;
assign w5757 = (w6415 & ~w5934) | (w6415 & w6717) | (~w5934 & w6717);
assign w5758 = (w3609 & w5799) | (w3609 & ~w3391) | (w5799 & ~w3391);
assign w5759 = a120 & b120;
assign w5760 = a172 & b172;
assign w5761 = (w401 & w6272) | (w401 & w7607) | (w6272 & w7607);
assign w5762 = ~a5 & ~b5;
assign w5763 = ~w1991 & ~w5123;
assign w5764 = ~w1191 & ~w120;
assign w5765 = (w101 & ~w2818) | (w101 & ~w7453) | (~w2818 & ~w7453);
assign w5766 = (w7067 & ~w1141) | (w7067 & ~w4875) | (~w1141 & ~w4875);
assign w5767 = w7625 & w205;
assign w5768 = (w3518 & w1639) | (w3518 & w1676) | (w1639 & w1676);
assign w5769 = (~w3758 & w1611) | (~w3758 & w1636) | (w1611 & w1636);
assign w5770 = w1754 & ~w1532;
assign w5771 = ~w4681 & ~w5464;
assign w5772 = ~a252 & ~b252;
assign w5773 = ~w4147 & ~w6871;
assign w5774 = ~w2741 & w2271;
assign w5775 = ~w6040 & ~w4760;
assign w5776 = (w3736 & w7309) | (w3736 & w521) | (w7309 & w521);
assign w5777 = ~w301 & ~w2278;
assign w5778 = ~w6195 & ~w5464;
assign w5779 = ~w5403 & ~w1570;
assign w5780 = (w6419 & w5657) | (w6419 & ~w6685) | (w5657 & ~w6685);
assign w5781 = w878 & ~w7486;
assign w5782 = a129 & b129;
assign w5783 = ~w2278 & ~w3724;
assign w5784 = ~w6481 & ~w1723;
assign w5785 = (w777 & w712) | (w777 & w3583) | (w712 & w3583);
assign w5786 = w1053 & w6577;
assign w5787 = w2856 & w6283;
assign w5788 = ~w706 & ~w1972;
assign w5789 = w2271 & w3679;
assign w5790 = (~w2890 & w4926) | (~w2890 & w2841) | (w4926 & w2841);
assign w5791 = (w4383 & w6348) | (w4383 & w474) | (w6348 & w474);
assign w5792 = ~w4775 & ~w5900;
assign w5793 = (~w7554 & w2156) | (~w7554 & w2722) | (w2156 & w2722);
assign w5794 = ~w1860 & ~w4468;
assign w5795 = (~w3989 & w1134) | (~w3989 & w2820) | (w1134 & w2820);
assign w5796 = (w6254 & w582) | (w6254 & w6482) | (w582 & w6482);
assign w5797 = ~w3896 & w2907;
assign w5798 = w1077 & ~w3741;
assign w5799 = (~w4967 & w4363) | (~w4967 & w1752) | (w4363 & w1752);
assign w5800 = (~w4967 & w4095) | (~w4967 & w4341) | (w4095 & w4341);
assign w5801 = ~w5958 & ~w2740;
assign w5802 = w4169 & ~w869;
assign w5803 = (~w100 & w2672) | (~w100 & w5568) | (w2672 & w5568);
assign w5804 = (w3658 & w747) | (w3658 & w883) | (w747 & w883);
assign w5805 = w7566 & ~w1328;
assign w5806 = (w5223 & ~w5259) | (w5223 & w1136) | (~w5259 & w1136);
assign w5807 = ~w4584 & ~w1532;
assign w5808 = ~a190 & ~b190;
assign w5809 = ~w1925 & w1140;
assign w5810 = (w6274 & w2961) | (w6274 & w4521) | (w2961 & w4521);
assign w5811 = (w6781 & w2940) | (w6781 & ~w563) | (w2940 & ~w563);
assign w5812 = (~w7513 & w1978) | (~w7513 & w564) | (w1978 & w564);
assign w5813 = ~w7000 & ~w7190;
assign w5814 = (~w4415 & w2745) | (~w4415 & w628) | (w2745 & w628);
assign w5815 = (w6084 & w4595) | (w6084 & w3112) | (w4595 & w3112);
assign w5816 = ~w3726 & w3127;
assign w5817 = (w3318 & w4633) | (w3318 & w4037) | (w4633 & w4037);
assign w5818 = (~w7626 & w3206) | (~w7626 & w5328) | (w3206 & w5328);
assign w5819 = w7633 & ~w1435;
assign w5820 = ~a248 & ~b248;
assign w5821 = ~w1565 & w6660;
assign w5822 = w1284 & w3014;
assign w5823 = ~w6524 & ~w1511;
assign w5824 = (w401 & w5761) | (w401 & w2453) | (w5761 & w2453);
assign w5825 = (~w6922 & w7154) | (~w6922 & w7015) | (w7154 & w7015);
assign w5826 = w2131 & ~w527;
assign w5827 = w151 & ~w6037;
assign w5828 = ~w1849 & w3433;
assign w5829 = (w5655 & w249) | (w5655 & w2585) | (w249 & w2585);
assign w5830 = ~w5118 & w4003;
assign w5831 = (~w5178 & w4785) | (~w5178 & w4042) | (w4785 & w4042);
assign w5832 = w313 & ~w1658;
assign w5833 = w767 & ~w6504;
assign w5834 = (~w3318 & w5291) | (~w3318 & w563) | (w5291 & w563);
assign w5835 = w2988 & w1906;
assign w5836 = (~w2725 & w3224) | (~w2725 & w5040) | (w3224 & w5040);
assign w5837 = ~w3409 & w7539;
assign w5838 = w7114 & w5675;
assign w5839 = ~w2401 & ~w1321;
assign w5840 = (~w1722 & w7562) | (~w1722 & w4867) | (w7562 & w4867);
assign w5841 = w5983 & w5069;
assign w5842 = ~w561 & w2384;
assign w5843 = w2750 & ~w5035;
assign w5844 = w1283 & ~w7447;
assign w5845 = (w2225 & w6186) | (w2225 & w3119) | (w6186 & w3119);
assign w5846 = w5752 & ~w7610;
assign w5847 = (w629 & w2857) | (w629 & w108) | (w2857 & w108);
assign w5848 = w6351 & w769;
assign w5849 = ~w2718 & ~w5239;
assign w5850 = (w7255 & w7528) | (w7255 & w253) | (w7528 & w253);
assign w5851 = (w3057 & w1508) | (w3057 & w667) | (w1508 & w667);
assign w5852 = w1364 & ~w4152;
assign w5853 = w3134 & ~w5391;
assign w5854 = (~w4327 & w3431) | (~w4327 & w6799) | (w3431 & w6799);
assign w5855 = (~w3952 & w3259) | (~w3952 & w6745) | (w3259 & w6745);
assign w5856 = ~w808 & ~w2732;
assign w5857 = (~w6647 & w4429) | (~w6647 & ~w4487) | (w4429 & ~w4487);
assign w5858 = ~w5463 & w2288;
assign w5859 = (w3318 & w1717) | (w3318 & w2525) | (w1717 & w2525);
assign w5860 = ~w4881 & ~w3712;
assign w5861 = (w5834 & w530) | (w5834 & w7170) | (w530 & w7170);
assign w5862 = a143 & b143;
assign w5863 = ~a149 & ~b149;
assign w5864 = a23 & b23;
assign w5865 = (~w6467 & w2170) | (~w6467 & w116) | (w2170 & w116);
assign w5866 = ~w5641 & ~w4592;
assign w5867 = (w5068 & w6918) | (w5068 & ~w4803) | (w6918 & ~w4803);
assign w5868 = (w3709 & w1506) | (w3709 & ~w5839) | (w1506 & ~w5839);
assign w5869 = (w3983 & w3966) | (w3983 & w6856) | (w3966 & w6856);
assign w5870 = (~w6658 & ~w6448) | (~w6658 & w7537) | (~w6448 & w7537);
assign w5871 = ~w5827 & w3632;
assign w5872 = (w5345 & w1334) | (w5345 & w5430) | (w1334 & w5430);
assign w5873 = (~w2453 & ~w6738) | (~w2453 & ~w7124) | (~w6738 & ~w7124);
assign w5874 = (~w3318 & w5261) | (~w3318 & w662) | (w5261 & w662);
assign w5875 = w4282 & ~w1897;
assign w5876 = (w4510 & w7478) | (w4510 & w3088) | (w7478 & w3088);
assign w5877 = ~w1038 & w1379;
assign w5878 = (w1369 & w3989) | (w1369 & w1101) | (w3989 & w1101);
assign w5879 = ~w7299 & ~w1279;
assign w5880 = w367 | w5739;
assign w5881 = ~w2631 & ~w5053;
assign w5882 = w6422 & w6586;
assign w5883 = a87 & b87;
assign w5884 = (w5655 & w4919) | (w5655 & w2698) | (w4919 & w2698);
assign w5885 = (w1555 & w6722) | (w1555 & ~w512) | (w6722 & ~w512);
assign w5886 = (~w2928 & w3671) | (~w2928 & w2136) | (w3671 & w2136);
assign w5887 = (~w7027 & w6675) | (~w7027 & w6607) | (w6675 & w6607);
assign w5888 = ~w51 & ~w4921;
assign w5889 = ~w4047 & ~w4023;
assign w5890 = ~w3152 & ~w1031;
assign w5891 = (~w2627 & w2102) | (~w2627 & w7441) | (w2102 & w7441);
assign w5892 = ~w813 & w4340;
assign w5893 = (~w5078 & w7559) | (~w5078 & w3013) | (w7559 & w3013);
assign w5894 = (~w6082 & w6568) | (~w6082 & w3910) | (w6568 & w3910);
assign w5895 = ~w7627 & w6073;
assign w5896 = (w5834 & w6417) | (w5834 & w1816) | (w6417 & w1816);
assign w5897 = (w6354 & w3385) | (w6354 & w4087) | (w3385 & w4087);
assign w5898 = (w342 & w7013) | (w342 & w52) | (w7013 & w52);
assign w5899 = ~w887 & ~w2559;
assign w5900 = ~a39 & ~b39;
assign w5901 = ~w2407 & w7113;
assign w5902 = ~w1792 & w7599;
assign w5903 = (~w1925 & w1731) | (~w1925 & w4114) | (w1731 & w4114);
assign w5904 = (w7554 & w2994) | (w7554 & w6944) | (w2994 & w6944);
assign w5905 = (~w1598 & w750) | (~w1598 & w77) | (w750 & w77);
assign w5906 = w5978 & ~w4200;
assign w5907 = (w1097 & w1872) | (w1097 & w5430) | (w1872 & w5430);
assign w5908 = w580 & ~w2115;
assign w5909 = w2294 & ~w5522;
assign w5910 = (w2301 & w7006) | (w2301 & w4867) | (w7006 & w4867);
assign w5911 = (~w924 & w4288) | (~w924 & w4767) | (w4288 & w4767);
assign w5912 = (~w3359 & ~w3854) | (~w3359 & w607) | (~w3854 & w607);
assign w5913 = (w4075 & w5363) | (w4075 & w7015) | (w5363 & w7015);
assign w5914 = ~w2243 & ~w1196;
assign w5915 = ~a183 & ~b183;
assign w5916 = ~w1443 & ~w1153;
assign w5917 = (~w5106 & w4716) | (~w5106 & w3145) | (w4716 & w3145);
assign w5918 = (~w2935 & w5127) | (~w2935 & w72) | (w5127 & w72);
assign w5919 = (w3516 & w7643) | (w3516 & w3027) | (w7643 & w3027);
assign w5920 = w6466 | w5226;
assign w5921 = w3117 & ~w3473;
assign w5922 = ~w2984 & ~w102;
assign w5923 = a88 & b88;
assign w5924 = ~w2829 & w226;
assign w5925 = ~w2021 & w7386;
assign w5926 = a248 & b248;
assign w5927 = (~w960 & w3473) | (~w960 & w1440) | (w3473 & w1440);
assign w5928 = (w5325 & w6583) | (w5325 & w5238) | (w6583 & w5238);
assign w5929 = ~w2814 & w1452;
assign w5930 = ~a229 & ~b229;
assign w5931 = (w4908 & w3159) | (w4908 & w4459) | (w3159 & w4459);
assign w5932 = (w6100 & w2459) | (w6100 & w7021) | (w2459 & w7021);
assign w5933 = (w2627 & w5578) | (w2627 & w6007) | (w5578 & w6007);
assign w5934 = w3197 & w6397;
assign w5935 = w2863 & w7567;
assign w5936 = (w6100 & w3972) | (w6100 & w1413) | (w3972 & w1413);
assign w5937 = ~w2591 & ~w4533;
assign w5938 = (w2297 & w2456) | (w2297 & w7122) | (w2456 & w7122);
assign w5939 = ~w1788 & w1882;
assign w5940 = ~w3279 & ~w4920;
assign w5941 = ~w1315 & w4011;
assign w5942 = (~w6184 & w84) | (~w6184 & w4735) | (w84 & w4735);
assign w5943 = (w7587 & w5458) | (w7587 & w3952) | (w5458 & w3952);
assign w5944 = (w3490 & w6026) | (w3490 & w6669) | (w6026 & w6669);
assign w5945 = w1502 | w5963;
assign w5946 = (w6386 & ~w855) | (w6386 & w1789) | (~w855 & w1789);
assign w5947 = ~w5691 & ~w6010;
assign w5948 = (~w656 & w259) | (~w656 & w1451) | (w259 & w1451);
assign w5949 = ~w2539 & ~w1750;
assign w5950 = ~a171 & ~b171;
assign w5951 = (w2210 & w2877) | (w2210 & w3417) | (w2877 & w3417);
assign w5952 = (~w5655 & w2443) | (~w5655 & w635) | (w2443 & w635);
assign w5953 = (w1332 & w6326) | (w1332 & ~w7124) | (w6326 & ~w7124);
assign w5954 = w5246 & w3509;
assign w5955 = ~w2649 & ~w2296;
assign w5956 = (w3467 & ~w935) | (w3467 & w110) | (~w935 & w110);
assign w5957 = (~w5325 & w2805) | (~w5325 & w4058) | (w2805 & w4058);
assign w5958 = ~a231 & ~b231;
assign w5959 = ~w4350 & ~w927;
assign w5960 = ~w6980 & ~w7142;
assign w5961 = ~w5403 & w2335;
assign w5962 = ~w1030 & ~w6709;
assign w5963 = w4045 & ~w1740;
assign w5964 = w7005 & ~w5958;
assign w5965 = ~w3073 & ~w2600;
assign w5966 = a79 & b79;
assign w5967 = (~w6082 & w1275) | (~w6082 & w487) | (w1275 & w487);
assign w5968 = ~w1423 & ~w6987;
assign w5969 = (w3434 & w5823) | (w3434 & ~w1743) | (w5823 & ~w1743);
assign w5970 = (~w3014 & w512) | (~w3014 & w3078) | (w512 & w3078);
assign w5971 = ~w1358 & ~w4217;
assign w5972 = ~w1839 & ~w5295;
assign w5973 = (~w231 & w1525) | (~w231 & w1914) | (w1525 & w1914);
assign w5974 = (w7332 & w4948) | (w7332 & w3767) | (w4948 & w3767);
assign w5975 = (w6467 & w1448) | (w6467 & w3725) | (w1448 & w3725);
assign w5976 = (w3427 & w7600) | (w3427 & ~w4684) | (w7600 & ~w4684);
assign w5977 = w6206 & ~w5760;
assign w5978 = ~w4412 & ~w1515;
assign w5979 = (w4392 & w4155) | (w4392 & w426) | (w4155 & w426);
assign w5980 = ~w1308 & w6861;
assign w5981 = (~w1631 & w154) | (~w1631 & w5766) | (w154 & w5766);
assign w5982 = (~w3741 & w1077) | (~w3741 & w7454) | (w1077 & w7454);
assign w5983 = ~a184 & ~b184;
assign w5984 = (w1742 & w3111) | (w1742 & ~w990) | (w3111 & ~w990);
assign w5985 = (~w7471 & w3146) | (~w7471 & ~w5350) | (w3146 & ~w5350);
assign w5986 = ~w651 & w1143;
assign w5987 = w5292 & ~w3710;
assign w5988 = (w3947 & w2823) | (w3947 & w6888) | (w2823 & w6888);
assign w5989 = ~w1439 & ~w6864;
assign w5990 = (w6166 & w3540) | (w6166 & w7124) | (w3540 & w7124);
assign w5991 = w7013 | w342;
assign w5992 = ~w5226 & w4039;
assign w5993 = ~w3128 & w2706;
assign w5994 = (w5672 & w2265) | (w5672 & w4128) | (w2265 & w4128);
assign w5995 = (~w6981 & w3168) | (~w6981 & w2371) | (w3168 & w2371);
assign w5996 = ~w5466 & w6791;
assign w5997 = (w6846 & w235) | (w6846 & w365) | (w235 & w365);
assign w5998 = ~w2353 & ~w1799;
assign w5999 = ~a44 & ~b44;
assign w6000 = (w5262 & w6080) | (w5262 & w2507) | (w6080 & w2507);
assign w6001 = (w342 & w7013) | (w342 & w3953) | (w7013 & w3953);
assign w6002 = ~w3392 & ~w3135;
assign w6003 = ~w977 & ~w7436;
assign w6004 = w740 & ~w5635;
assign w6005 = ~w5888 & w388;
assign w6006 = ~w2364 & ~w2201;
assign w6007 = (w6680 & w4696) | (w6680 & w1770) | (w4696 & w1770);
assign w6008 = (~w6100 & w6150) | (~w6100 & w5894) | (w6150 & w5894);
assign w6009 = ~w1300 & w2081;
assign w6010 = w4918 & w5381;
assign w6011 = (w6738 & w3343) | (w6738 & w677) | (w3343 & w677);
assign w6012 = w3134 & ~w3145;
assign w6013 = ~w3183 & w7438;
assign w6014 = (w6649 & w519) | (w6649 & w4730) | (w519 & w4730);
assign w6015 = w412 & w1070;
assign w6016 = (~w6981 & w1030) | (~w6981 & w325) | (w1030 & w325);
assign w6017 = w3145 & ~w4499;
assign w6018 = (~w4995 & w7366) | (~w4995 & w5379) | (w7366 & w5379);
assign w6019 = w3396 & w512;
assign w6020 = (w3560 & w2117) | (w3560 & ~w484) | (w2117 & ~w484);
assign w6021 = (~w3636 & w180) | (~w3636 & w5173) | (w180 & w5173);
assign w6022 = w4471 & w6733;
assign w6023 = w523 & w7451;
assign w6024 = ~w6254 & w7102;
assign w6025 = ~a62 & ~b62;
assign w6026 = w3959 & ~w1295;
assign w6027 = w1006 & ~w3819;
assign w6028 = ~w2605 & w4749;
assign w6029 = ~w7272 & ~w6404;
assign w6030 = (~w2985 & w1305) | (~w2985 & w1700) | (w1305 & w1700);
assign w6031 = w5259 & w2798;
assign w6032 = ~w1849 & ~w142;
assign w6033 = ~w5466 & ~w6243;
assign w6034 = (w3060 & w5312) | (w3060 & ~w6894) | (w5312 & ~w6894);
assign w6035 = (~w6100 & w6786) | (~w6100 & w3513) | (w6786 & w3513);
assign w6036 = (~w3974 & w7461) | (~w3974 & w1847) | (w7461 & w1847);
assign w6037 = w6427 & w5489;
assign w6038 = (~w3986 & w4214) | (~w3986 & w2209) | (w4214 & w2209);
assign w6039 = w5042 & w3672;
assign w6040 = (~w2123 & w2891) | (~w2123 & w6036) | (w2891 & w6036);
assign w6041 = ~w2279 & ~w7622;
assign w6042 = w4330 & w755;
assign w6043 = ~w1252 & ~w937;
assign w6044 = w7279 & w6991;
assign w6045 = (w887 & ~w1455) | (w887 & w3394) | (~w1455 & w3394);
assign w6046 = w91 & ~w441;
assign w6047 = (w5834 & w7136) | (w5834 & w1319) | (w7136 & w1319);
assign w6048 = (w6942 & w6148) | (w6942 & w6965) | (w6148 & w6965);
assign w6049 = ~w3033 & w7032;
assign w6050 = (~w6100 & w4861) | (~w6100 & w5815) | (w4861 & w5815);
assign w6051 = ~w5403 & ~w887;
assign w6052 = (~w6272 & w970) | (~w6272 & w107) | (w970 & w107);
assign w6053 = (~w7268 & w2418) | (~w7268 & w7) | (w2418 & w7);
assign w6054 = ~a128 & ~b128;
assign w6055 = (w6031 & w2187) | (w6031 & w1342) | (w2187 & w1342);
assign w6056 = (w5178 & w4739) | (w5178 & w1572) | (w4739 & w1572);
assign w6057 = ~w4808 & w1135;
assign w6058 = ~w434 & w6597;
assign w6059 = (w3205 & w1963) | (w3205 & w166) | (w1963 & w166);
assign w6060 = (~w189 & w5178) | (~w189 & w3596) | (w5178 & w3596);
assign w6061 = ~w5205 & ~w909;
assign w6062 = w2380 & w86;
assign w6063 = ~w2066 & w2649;
assign w6064 = ~w561 & ~w1555;
assign w6065 = (w3054 & w6105) | (w3054 & w5655) | (w6105 & w5655);
assign w6066 = (w3473 & w5528) | (w3473 & ~w5178) | (w5528 & ~w5178);
assign w6067 = ~w1658 & w1737;
assign w6068 = w4021 & w1036;
assign w6069 = ~w7495 & ~w6783;
assign w6070 = w6803 & ~w1621;
assign w6071 = (~w4967 & w1414) | (~w4967 & w1309) | (w1414 & w1309);
assign w6072 = w4049 | w5596;
assign w6073 = ~w3818 & ~w4;
assign w6074 = (w3788 & w2592) | (w3788 & w5395) | (w2592 & w5395);
assign w6075 = (w716 & w6929) | (w716 & ~w6894) | (w6929 & ~w6894);
assign w6076 = (~w7450 & w1926) | (~w7450 & w3238) | (w1926 & w3238);
assign w6077 = ~w1991 & ~w1127;
assign w6078 = w3032 & w5013;
assign w6079 = (w1692 & w5575) | (w1692 & ~w1892) | (w5575 & ~w1892);
assign w6080 = ~w6526 & ~w6626;
assign w6081 = w6122 & ~w4344;
assign w6082 = ~w3892 & w4339;
assign w6083 = (~w5178 & w2752) | (~w5178 & w4524) | (w2752 & w4524);
assign w6084 = ~w2279 & w139;
assign w6085 = (w5699 & w4948) | (w5699 & ~w6633) | (w4948 & ~w6633);
assign w6086 = ~w3892 & w2531;
assign w6087 = a40 & b40;
assign w6088 = (w632 & w3407) | (w632 & w2110) | (w3407 & w2110);
assign w6089 = w4069 & ~w2456;
assign w6090 = (w2524 & w5322) | (w2524 & w4231) | (w5322 & w4231);
assign w6091 = (w4989 & w99) | (w4989 & w6663) | (w99 & w6663);
assign w6092 = ~w5791 & ~w1561;
assign w6093 = w3514 & w1067;
assign w6094 = a170 & b170;
assign w6095 = ~w1709 & ~w4360;
assign w6096 = (w5901 & w2036) | (w5901 & w2746) | (w2036 & w2746);
assign w6097 = w6117 & ~w6162;
assign w6098 = (w5545 & w3532) | (w5545 & w5368) | (w3532 & w5368);
assign w6099 = (~w1279 & w2708) | (~w1279 & w2715) | (w2708 & w2715);
assign w6100 = (~w5834 & w2491) | (~w5834 & w789) | (w2491 & w789);
assign w6101 = ~w7216 & ~w7520;
assign w6102 = (w297 & w4579) | (w297 & ~w1881) | (w4579 & ~w1881);
assign w6103 = (~w2627 & w5084) | (~w2627 & w6240) | (w5084 & w6240);
assign w6104 = a166 & b166;
assign w6105 = (w2052 & w4246) | (w2052 & w7240) | (w4246 & w7240);
assign w6106 = (w2453 & w6738) | (w2453 & w5007) | (w6738 & w5007);
assign w6107 = ~w3444 & w4986;
assign w6108 = w1315 & w1843;
assign w6109 = (~w2203 & w5297) | (~w2203 & ~w3819) | (w5297 & ~w3819);
assign w6110 = w7310 & ~w5479;
assign w6111 = (~w2818 & ~w1728) | (~w2818 & w3655) | (~w1728 & w3655);
assign w6112 = ~w2847 & w2488;
assign w6113 = ~w4998 & w3547;
assign w6114 = ~w3512 & ~w2465;
assign w6115 = (~w5008 & w7469) | (~w5008 & w6977) | (w7469 & w6977);
assign w6116 = (w1548 & w7220) | (w1548 & ~w4521) | (w7220 & ~w4521);
assign w6117 = ~w5251 & ~w3055;
assign w6118 = (~w2335 & w2391) | (~w2335 & ~w3631) | (w2391 & ~w3631);
assign w6119 = ~w5370 & w1472;
assign w6120 = (~w6106 & w7084) | (~w6106 & w4031) | (w7084 & w4031);
assign w6121 = (w1890 & w4141) | (w1890 & ~w6100) | (w4141 & ~w6100);
assign w6122 = ~w3359 & ~w4584;
assign w6123 = ~w1754 & w4901;
assign w6124 = ~w4813 & ~w7540;
assign w6125 = ~w2408 & w1529;
assign w6126 = ~w2401 & w3951;
assign w6127 = (w5871 & w5526) | (w5871 & w5735) | (w5526 & w5735);
assign w6128 = ~w3895 & ~w885;
assign w6129 = (w3063 & w1444) | (w3063 & w6194) | (w1444 & w6194);
assign w6130 = (w6744 & w6425) | (w6744 & w4896) | (w6425 & w4896);
assign w6131 = (w1167 & w3296) | (w1167 & w5403) | (w3296 & w5403);
assign w6132 = ~w872 & ~w887;
assign w6133 = ~w254 & ~w2484;
assign w6134 = w7044 & ~w3903;
assign w6135 = (w3242 & w6523) | (w3242 & w563) | (w6523 & w563);
assign w6136 = w2540 & ~w6254;
assign w6137 = ~w2216 & w5121;
assign w6138 = a1 & b1;
assign w6139 = (~w2627 & w6655) | (~w2627 & w5052) | (w6655 & w5052);
assign w6140 = w1685 & ~w1023;
assign w6141 = ~w3551 & ~w1736;
assign w6142 = (~w3105 & ~w4190) | (~w3105 & w6894) | (~w4190 & w6894);
assign w6143 = (~w3057 & w6261) | (~w3057 & w7037) | (w6261 & w7037);
assign w6144 = ~w6465 & w544;
assign w6145 = (~w4169 & w5594) | (~w4169 & ~w7132) | (w5594 & ~w7132);
assign w6146 = (w6066 & w3293) | (w6066 & w6382) | (w3293 & w6382);
assign w6147 = a126 & b126;
assign w6148 = w2283 & w6942;
assign w6149 = ~w4648 & ~w7424;
assign w6150 = (w5441 & w5805) | (w5441 & w6174) | (w5805 & w6174);
assign w6151 = ~w54 & ~w3866;
assign w6152 = (~w3888 & ~w1903) | (~w3888 & ~w3679) | (~w1903 & ~w3679);
assign w6153 = (~w3852 & w470) | (~w3852 & w4846) | (w470 & w4846);
assign w6154 = ~w1510 & ~w6897;
assign w6155 = w2131 & w6990;
assign w6156 = (w2454 & w2828) | (w2454 & ~w6174) | (w2828 & ~w6174);
assign w6157 = (w1814 & w4358) | (w1814 & w1802) | (w4358 & w1802);
assign w6158 = w5686 & w149;
assign w6159 = w827 & ~w4635;
assign w6160 = ~w3866 & w3080;
assign w6161 = w1532 & ~w1441;
assign w6162 = ~w3262 & ~w5463;
assign w6163 = w2548 & ~w7124;
assign w6164 = (w2627 & w4816) | (w2627 & w7057) | (w4816 & w7057);
assign w6165 = (w4223 & w1613) | (w4223 & w6100) | (w1613 & w6100);
assign w6166 = (~w1473 & w7252) | (~w1473 & w2637) | (w7252 & w2637);
assign w6167 = (~w3327 & w258) | (~w3327 & w4667) | (w258 & w4667);
assign w6168 = (w1454 & w6198) | (w1454 & ~w1847) | (w6198 & ~w1847);
assign w6169 = a22 & b22;
assign w6170 = ~w6766 & ~w1057;
assign w6171 = ~w2662 & ~w22;
assign w6172 = (~w8 & w6360) | (~w8 & w1339) | (w6360 & w1339);
assign w6173 = ~w2011 & w2628;
assign w6174 = ~w6082 & w3684;
assign w6175 = (w1336 & w3975) | (w1336 & w4104) | (w3975 & w4104);
assign w6176 = (w3848 & w2263) | (w3848 & ~w6878) | (w2263 & ~w6878);
assign w6177 = (~w3318 & w7303) | (~w3318 & w1128) | (w7303 & w1128);
assign w6178 = ~w2428 & ~w4552;
assign w6179 = w7010 & w6600;
assign w6180 = (~w6770 & ~w464) | (~w6770 & ~w1770) | (~w464 & ~w1770);
assign w6181 = a171 & b171;
assign w6182 = (~w4564 & ~w6688) | (~w4564 & w2045) | (~w6688 & w2045);
assign w6183 = (w972 & ~w7429) | (w972 & w625) | (~w7429 & w625);
assign w6184 = ~w247 & ~w6252;
assign w6185 = (w5879 & w5252) | (w5879 & w139) | (w5252 & w139);
assign w6186 = (w4286 & w2225) | (w4286 & w4907) | (w2225 & w4907);
assign w6187 = w6058 & ~w1387;
assign w6188 = ~w7187 & w5415;
assign w6189 = ~w2474 & ~w3337;
assign w6190 = (~w2429 & w891) | (~w2429 & w4269) | (w891 & w4269);
assign w6191 = (~w1999 & ~w7563) | (~w1999 & w3995) | (~w7563 & w3995);
assign w6192 = (~w1455 & w1144) | (~w1455 & w4466) | (w1144 & w4466);
assign w6193 = (w2627 & w4059) | (w2627 & w786) | (w4059 & w786);
assign w6194 = (~w5194 & w4966) | (~w5194 & ~w2090) | (w4966 & ~w2090);
assign w6195 = ~w6279 & ~w5570;
assign w6196 = (~w5257 & w1011) | (~w5257 & w5684) | (w1011 & w5684);
assign w6197 = (w7095 & w572) | (w7095 & ~w6174) | (w572 & ~w6174);
assign w6198 = w6155 & ~w5430;
assign w6199 = (w5522 & w3993) | (w5522 & w901) | (w3993 & w901);
assign w6200 = ~w1554 & ~w3192;
assign w6201 = w2793 & ~w6100;
assign w6202 = (~w488 & ~w7029) | (~w488 & ~w7046) | (~w7029 & ~w7046);
assign w6203 = w6935 & ~w2515;
assign w6204 = (w6424 & w916) | (w6424 & w1218) | (w916 & w1218);
assign w6205 = (~w1228 & w6920) | (~w1228 & w6402) | (w6920 & w6402);
assign w6206 = ~a172 & ~b172;
assign w6207 = ~w7345 & ~w2456;
assign w6208 = (~w5655 & w3403) | (~w5655 & w7370) | (w3403 & w7370);
assign w6209 = ~a244 & ~b244;
assign w6210 = ~a185 & ~b185;
assign w6211 = ~w2104 & ~w3732;
assign w6212 = (w4889 & w4091) | (w4889 & ~w7124) | (w4091 & ~w7124);
assign w6213 = (w6099 & w4823) | (w6099 & w28) | (w4823 & w28);
assign w6214 = w4777 & ~w3888;
assign w6215 = (w7575 & w4967) | (w7575 & w4400) | (w4967 & w4400);
assign w6216 = (~w5743 & ~w47) | (~w5743 & w1981) | (~w47 & w1981);
assign w6217 = (w924 & w6203) | (w924 & w2413) | (w6203 & w2413);
assign w6218 = (w6100 & w183) | (w6100 & w2111) | (w183 & w2111);
assign w6219 = ~w2255 & w3113;
assign w6220 = w6539 & w4514;
assign w6221 = (w2627 & w4704) | (w2627 & w835) | (w4704 & w835);
assign w6222 = ~a59 & ~b59;
assign w6223 = (~w1878 & w2182) | (~w1878 & w940) | (w2182 & w940);
assign w6224 = ~w4179 & ~w5633;
assign w6225 = ~w1026 & ~w706;
assign w6226 = w6181 & ~w6206;
assign w6227 = (w484 & w7015) | (w484 & ~w563) | (w7015 & ~w563);
assign w6228 = (w3892 & w2402) | (w3892 & w4856) | (w2402 & w4856);
assign w6229 = (w2721 & w6686) | (w2721 & ~w3330) | (w6686 & ~w3330);
assign w6230 = ~w4504 & ~w4468;
assign w6231 = w3570 & ~w5152;
assign w6232 = (~w2627 & w3849) | (~w2627 & w1310) | (w3849 & w1310);
assign w6233 = ~w390 & ~w604;
assign w6234 = w3938 | w6724;
assign w6235 = (w5961 & w7325) | (w5961 & w816) | (w7325 & w816);
assign w6236 = (w834 & ~w3491) | (w834 & w1956) | (~w3491 & w1956);
assign w6237 = (~w2243 & w5600) | (~w2243 & w1379) | (w5600 & w1379);
assign w6238 = (w5537 & w1500) | (w5537 & w6254) | (w1500 & w6254);
assign w6239 = w3580 & ~w6209;
assign w6240 = (~w3983 & w97) | (~w3983 & w467) | (w97 & w467);
assign w6241 = ~w4909 & ~w5055;
assign w6242 = (~w6252 & w4232) | (~w6252 & w3014) | (w4232 & w3014);
assign w6243 = a164 & b164;
assign w6244 = ~w2769 & ~w2969;
assign w6245 = ~w3991 & ~w1445;
assign w6246 = ~w6346 & ~w7632;
assign w6247 = (w6438 & w4005) | (w6438 & w5655) | (w4005 & w5655);
assign w6248 = (w2401 & w6486) | (w2401 & w1226) | (w6486 & w1226);
assign w6249 = (w1284 & w6537) | (w1284 & ~w5871) | (w6537 & ~w5871);
assign w6250 = w1431 & ~w7390;
assign w6251 = ~w2769 & ~w2718;
assign w6252 = a210 & b210;
assign w6253 = w479 & ~w7491;
assign w6254 = ~w6397 & w4942;
assign w6255 = ~w7127 & ~w2365;
assign w6256 = w4998 & ~w1958;
assign w6257 = ~w1544 & ~w2019;
assign w6258 = (w297 & w4579) | (w297 & ~w4521) | (w4579 & ~w4521);
assign w6259 = w2907 & ~w5738;
assign w6260 = ~w53 & w4295;
assign w6261 = ~w2740 & w4123;
assign w6262 = (w6112 & w4554) | (w6112 & w876) | (w4554 & w876);
assign w6263 = (w3657 & w5587) | (w3657 & w6127) | (w5587 & w6127);
assign w6264 = ~w6757 & w6981;
assign w6265 = ~w3224 & w4514;
assign w6266 = (~w1760 & w4634) | (~w1760 & ~w4214) | (w4634 & ~w4214);
assign w6267 = ~w1692 & w2453;
assign w6268 = w4471 & ~w4132;
assign w6269 = (~w5995 & w5954) | (~w5995 & w6739) | (w5954 & w6739);
assign w6270 = ~w3290 & ~w3137;
assign w6271 = w6713 & ~w6911;
assign w6272 = ~w3959 & w4130;
assign w6273 = (w6106 & w1317) | (w6106 & w7400) | (w1317 & w7400);
assign w6274 = w106 & ~w6324;
assign w6275 = (w7239 & w5551) | (w7239 & w1631) | (w5551 & w1631);
assign w6276 = w2782 & ~w4142;
assign w6277 = (~w6162 & w6117) | (~w6162 & w2163) | (w6117 & w2163);
assign w6278 = (w3434 & w5823) | (w3434 & ~w3989) | (w5823 & ~w3989);
assign w6279 = a73 & b73;
assign w6280 = ~w4906 & w6951;
assign w6281 = a51 & b51;
assign w6282 = (~w3210 & w4611) | (~w3210 & w6882) | (w4611 & w6882);
assign w6283 = ~w1477 & w2535;
assign w6284 = (~w7197 & w3255) | (~w7197 & w1411) | (w3255 & w1411);
assign w6285 = w4438 & ~w7172;
assign w6286 = w5112 & w3696;
assign w6287 = (w846 & w3986) | (w846 & w782) | (w3986 & w782);
assign w6288 = (~w501 & w1672) | (~w501 & w5133) | (w1672 & w5133);
assign w6289 = (~w777 & w6258) | (~w777 & w6102) | (w6258 & w6102);
assign w6290 = w5978 & ~w5493;
assign w6291 = ~w4788 & ~w6209;
assign w6292 = w6195 & ~w5299;
assign w6293 = (~w5834 & w4842) | (~w5834 & w1059) | (w4842 & w1059);
assign w6294 = (~w6911 & w6271) | (~w6911 & ~w5655) | (w6271 & ~w5655);
assign w6295 = (w4964 & w7290) | (w4964 & w3391) | (w7290 & w3391);
assign w6296 = (w7002 & w4139) | (w7002 & w1192) | (w4139 & w1192);
assign w6297 = ~w1827 & w1722;
assign w6298 = (~w3619 & w6871) | (~w3619 & w3702) | (w6871 & w3702);
assign w6299 = w1923 & ~w1158;
assign w6300 = w5155 & w6126;
assign w6301 = ~w3123 & ~w1848;
assign w6302 = (w4604 & w1828) | (w4604 & ~w5484) | (w1828 & ~w5484);
assign w6303 = ~w6452 & w5072;
assign w6304 = a60 & b60;
assign w6305 = (w484 & w797) | (w484 & w1602) | (w797 & w1602);
assign w6306 = (~w588 & w4125) | (~w588 & w6361) | (w4125 & w6361);
assign w6307 = w5837 & ~w2624;
assign w6308 = ~w7597 & w4532;
assign w6309 = ~w4222 & w472;
assign w6310 = ~w4004 & ~w3351;
assign w6311 = ~w7346 & w2534;
assign w6312 = (~w6100 & w3882) | (~w6100 & w153) | (w3882 & w153);
assign w6313 = (w5226 & w6466) | (w5226 & w6510) | (w6466 & w6510);
assign w6314 = (w6945 & w2562) | (w6945 & w5021) | (w2562 & w5021);
assign w6315 = w5620 & w5303;
assign w6316 = (~w5641 & w2041) | (~w5641 & w7569) | (w2041 & w7569);
assign w6317 = w2385 & w7181;
assign w6318 = w4771 & ~w6387;
assign w6319 = a151 & b151;
assign w6320 = ~w4399 & ~w611;
assign w6321 = ~w2339 & w4836;
assign w6322 = (~w7015 & w495) | (~w7015 & w3442) | (w495 & w3442);
assign w6323 = ~w3838 & w4960;
assign w6324 = (~w3984 & w4699) | (~w3984 & w6004) | (w4699 & w6004);
assign w6325 = ~w6426 & ~w6912;
assign w6326 = (~w3057 & w1332) | (~w3057 & w5814) | (w1332 & w5814);
assign w6327 = ~w3176 & w1832;
assign w6328 = (~w3840 & w1021) | (~w3840 & w4392) | (w1021 & w4392);
assign w6329 = w1999 & ~w1954;
assign w6330 = (~w6424 & w6841) | (~w6424 & w5548) | (w6841 & w5548);
assign w6331 = ~a134 & ~b134;
assign w6332 = (w2847 & w3575) | (w2847 & w993) | (w3575 & w993);
assign w6333 = (~w185 & w7477) | (~w185 & w5367) | (w7477 & w5367);
assign w6334 = w6518 & w2664;
assign w6335 = ~a113 & ~b113;
assign w6336 = ~w2210 & ~w4090;
assign w6337 = (~w4651 & w5553) | (~w4651 & w1449) | (w5553 & w1449);
assign w6338 = w1364 & ~w1736;
assign w6339 = w1849 & ~w5251;
assign w6340 = (w5178 & w3680) | (w5178 & w2262) | (w3680 & w2262);
assign w6341 = w4661 & w4691;
assign w6342 = a127 & b127;
assign w6343 = w3774 & w5288;
assign w6344 = (~w2123 & w4519) | (~w2123 & w4982) | (w4519 & w4982);
assign w6345 = ~w4415 & w2360;
assign w6346 = ~a95 & ~b95;
assign w6347 = w6787 | w6570;
assign w6348 = (w6989 & w1210) | (w6989 & w6566) | (w1210 & w6566);
assign w6349 = ~w2504 & ~w2106;
assign w6350 = (~w6252 & w84) | (~w6252 & w6242) | (w84 & w6242);
assign w6351 = ~w2688 & ~w5289;
assign w6352 = (~w5830 & w4202) | (~w5830 & w6276) | (w4202 & w6276);
assign w6353 = (w1973 & w488) | (w1973 & w1320) | (w488 & w1320);
assign w6354 = ~w3918 & ~w3618;
assign w6355 = (w7563 & w317) | (w7563 & ~w6981) | (w317 & ~w6981);
assign w6356 = w4545 & ~w4884;
assign w6357 = ~w5966 & ~w1621;
assign w6358 = ~w6167 & ~w1824;
assign w6359 = (w264 & w3315) | (w264 & w2674) | (w3315 & w2674);
assign w6360 = w7024 & ~w4807;
assign w6361 = (~w6467 & w7468) | (~w6467 & w5500) | (w7468 & w5500);
assign w6362 = ~w7408 & w1879;
assign w6363 = (w1936 & w35) | (w1936 & w955) | (w35 & w955);
assign w6364 = (w5556 & w6814) | (w5556 & ~w1982) | (w6814 & ~w1982);
assign w6365 = w5559 & ~w6385;
assign w6366 = ~w444 & ~w2216;
assign w6367 = w5463 & ~w7493;
assign w6368 = (~w2838 & w7582) | (~w2838 & ~w6894) | (w7582 & ~w6894);
assign w6369 = (~w2182 & w4381) | (~w2182 & w1220) | (w4381 & w1220);
assign w6370 = w2522 & w5819;
assign w6371 = w4496 & ~w4418;
assign w6372 = (~w3984 & w5020) | (~w3984 & w1734) | (w5020 & w1734);
assign w6373 = ~w5797 & w6920;
assign w6374 = (w6100 & w2555) | (w6100 & w3902) | (w2555 & w3902);
assign w6375 = w4648 & ~w6810;
assign w6376 = (~w2123 & w5247) | (~w2123 & w4860) | (w5247 & w4860);
assign w6377 = w4415 & ~w5781;
assign w6378 = w3690 & ~w810;
assign w6379 = (w478 & w2169) | (w478 & w707) | (w2169 & w707);
assign w6380 = ~w7153 & ~w1126;
assign w6381 = (~w424 & w321) | (~w424 & w7313) | (w321 & w7313);
assign w6382 = (w3491 & w4539) | (w3491 & w3465) | (w4539 & w3465);
assign w6383 = ~w4140 & ~w3863;
assign w6384 = ~w6254 & w68;
assign w6385 = (~w4242 & w5077) | (~w4242 & w5571) | (w5077 & w5571);
assign w6386 = ~w3101 & ~w3244;
assign w6387 = ~w7507 & ~w3587;
assign w6388 = w775 & ~w5267;
assign w6389 = w6054 & w3045;
assign w6390 = (w7405 & w6497) | (w7405 & w5493) | (w6497 & w5493);
assign w6391 = (w6792 & w6390) | (w6792 & w794) | (w6390 & w794);
assign w6392 = ~a230 & ~b230;
assign w6393 = ~w3663 & ~w5354;
assign w6394 = ~w2486 & ~w1034;
assign w6395 = (w5522 & w4935) | (w5522 & w5692) | (w4935 & w5692);
assign w6396 = w4459 & w1006;
assign w6397 = ~w5830 & w369;
assign w6398 = (w5178 & w315) | (w5178 & w879) | (w315 & w879);
assign w6399 = w7283 & w4061;
assign w6400 = (~w5291 & w5088) | (~w5291 & w6282) | (w5088 & w6282);
assign w6401 = ~w1162 & w5226;
assign w6402 = ~w1228 & w6147;
assign w6403 = ~w4638 & ~w960;
assign w6404 = (w7519 & w4191) | (w7519 & w327) | (w4191 & w327);
assign w6405 = (w5231 & w6967) | (w5231 & w5325) | (w6967 & w5325);
assign w6406 = w508 & ~w4458;
assign w6407 = ~w1384 & w5686;
assign w6408 = (w6357 & ~w2380) | (w6357 & w3178) | (~w2380 & w3178);
assign w6409 = w5860 & w692;
assign w6410 = w6299 & ~w1158;
assign w6411 = (~w2124 & w5903) | (~w2124 & w3760) | (w5903 & w3760);
assign w6412 = (w1190 & w3556) | (w1190 & w4811) | (w3556 & w4811);
assign w6413 = (w1607 & w6830) | (w1607 & w6972) | (w6830 & w6972);
assign w6414 = w649 & ~w6658;
assign w6415 = ~w1308 & w3003;
assign w6416 = (~w3952 & w3377) | (~w3952 & w822) | (w3377 & w822);
assign w6417 = (~w1730 & w3980) | (~w1730 & w3125) | (w3980 & w3125);
assign w6418 = (w6174 & w737) | (w6174 & w5765) | (w737 & w5765);
assign w6419 = (~w486 & w4043) | (~w486 & w112) | (w4043 & w112);
assign w6420 = ~w6630 & ~w4733;
assign w6421 = (w2415 & w3571) | (w2415 & w3708) | (w3571 & w3708);
assign w6422 = w1248 & w4727;
assign w6423 = (w1886 & w491) | (w1886 & w5078) | (w491 & w5078);
assign w6424 = w68 & w6174;
assign w6425 = (~w5881 & w1290) | (~w5881 & ~w2243) | (w1290 & ~w2243);
assign w6426 = ~a139 & ~b139;
assign w6427 = ~w4297 & ~w1386;
assign w6428 = ~w808 & ~w5916;
assign w6429 = w4960 & w3364;
assign w6430 = w4614 & ~w7566;
assign w6431 = (~w3490 & w7257) | (~w3490 & ~w5629) | (w7257 & ~w5629);
assign w6432 = (~w3983 & w1679) | (~w3983 & w7248) | (w1679 & w7248);
assign w6433 = (w1328 & w2130) | (w1328 & w5268) | (w2130 & w5268);
assign w6434 = w7362 & ~w1488;
assign w6435 = ~w4803 & w6436;
assign w6436 = ~w7528 & w3415;
assign w6437 = (~w5834 & w5038) | (~w5834 & w6670) | (w5038 & w6670);
assign w6438 = ~w486 & ~w5422;
assign w6439 = ~a15 & ~b15;
assign w6440 = (w1881 & w4888) | (w1881 & w1213) | (w4888 & w1213);
assign w6441 = (w1005 & w5043) | (w1005 & ~w5325) | (w5043 & ~w5325);
assign w6442 = ~w4206 & w3984;
assign w6443 = ~w5962 & w169;
assign w6444 = ~a121 & ~b121;
assign w6445 = ~w2566 & w6723;
assign w6446 = w234 & ~w3842;
assign w6447 = w3643 & w1891;
assign w6448 = ~w4438 & ~w4643;
assign w6449 = (~w6265 & w1475) | (~w6265 & w597) | (w1475 & w597);
assign w6450 = a229 & b229;
assign w6451 = ~w3075 & w2579;
assign w6452 = ~w4476 & ~w2027;
assign w6453 = (w2453 & w632) | (w2453 & w173) | (w632 & w173);
assign w6454 = w3105 & ~w1741;
assign w6455 = ~a48 & ~b48;
assign w6456 = (w1496 & w4046) | (w1496 & ~w4143) | (w4046 & ~w4143);
assign w6457 = w1962 | w4732;
assign w6458 = ~a61 & ~b61;
assign w6459 = (~w6520 & w4378) | (~w6520 & ~w1598) | (w4378 & ~w1598);
assign w6460 = (w5888 & ~w1751) | (w5888 & w1374) | (~w1751 & w1374);
assign w6461 = (w5967 & ~w6100) | (w5967 & w2094) | (~w6100 & w2094);
assign w6462 = ~w1725 & ~w195;
assign w6463 = a16 & b16;
assign w6464 = (~w2686 & w3116) | (~w2686 & w3948) | (w3116 & w3948);
assign w6465 = ~w1256 & ~w2643;
assign w6466 = w7188 & w5226;
assign w6467 = (~w5783 & w6037) | (~w5783 & w7223) | (w6037 & w7223);
assign w6468 = (~w3105 & ~w4190) | (~w3105 & ~w2456) | (~w4190 & ~w2456);
assign w6469 = w5288 & ~w6254;
assign w6470 = (w7024 & w2962) | (w7024 & w632) | (w2962 & w632);
assign w6471 = (~w4132 & w435) | (~w4132 & w7603) | (w435 & w7603);
assign w6472 = w3840 & w6682;
assign w6473 = (~w5178 & w1028) | (~w5178 & w1680) | (w1028 & w1680);
assign w6474 = (w5178 & w1764) | (w5178 & w3228) | (w1764 & w3228);
assign w6475 = ~w6325 & w5499;
assign w6476 = (~w5655 & w3923) | (~w5655 & w25) | (w3923 & w25);
assign w6477 = (w1919 & w3148) | (w1919 & w5722) | (w3148 & w5722);
assign w6478 = (~w7554 & w3797) | (~w7554 & w6091) | (w3797 & w6091);
assign w6479 = (w902 & ~w5259) | (w902 & w725) | (~w5259 & w725);
assign w6480 = (w6894 & w1197) | (w6894 & w2868) | (w1197 & w2868);
assign w6481 = ~w351 & ~w259;
assign w6482 = (w6046 & w582) | (w6046 & w2476) | (w582 & w2476);
assign w6483 = ~w4298 & ~w5612;
assign w6484 = ~w434 & ~w5557;
assign w6485 = (~w5914 & w4025) | (~w5914 & w6744) | (w4025 & w6744);
assign w6486 = ~w6181 & w4991;
assign w6487 = (~w5178 & w5396) | (~w5178 & w2092) | (w5396 & w2092);
assign w6488 = (w1611 & w7435) | (w1611 & w4662) | (w7435 & w4662);
assign w6489 = (~w6911 & w6271) | (~w6911 & w3402) | (w6271 & w3402);
assign w6490 = ~w4409 & ~w1756;
assign w6491 = (~w6127 & w6847) | (~w6127 & w2618) | (w6847 & w2618);
assign w6492 = ~w4564 & w1125;
assign w6493 = (w2993 & w1589) | (w2993 & w5233) | (w1589 & w5233);
assign w6494 = (w4756 & w4304) | (w4756 & w5291) | (w4304 & w5291);
assign w6495 = w5463 & ~w2068;
assign w6496 = (w699 & w455) | (w699 & ~w5304) | (w455 & ~w5304);
assign w6497 = ~w220 & w7405;
assign w6498 = (w702 & w1696) | (w702 & w4867) | (w1696 & w4867);
assign w6499 = ~w4287 & w6297;
assign w6500 = ~w642 & w2458;
assign w6501 = ~w6082 & w6024;
assign w6502 = (~w3527 & w2284) | (~w3527 & w5763) | (w2284 & w5763);
assign w6503 = ~w5923 & ~w216;
assign w6504 = ~w4035 & ~w290;
assign w6505 = (w7197 & w7234) | (w7197 & w942) | (w7234 & w942);
assign w6506 = (~w6738 & w29) | (~w6738 & w452) | (w29 & w452);
assign w6507 = ~w5827 & w2790;
assign w6508 = w5403 & w2522;
assign w6509 = (w3387 & ~w857) | (w3387 & ~w4138) | (~w857 & ~w4138);
assign w6510 = ~a20 & ~b20;
assign w6511 = (w931 & w5140) | (w931 & w6226) | (w5140 & w6226);
assign w6512 = ~w7633 & ~w638;
assign w6513 = ~w1980 & ~w7507;
assign w6514 = ~w4850 & ~w2590;
assign w6515 = w1689 & w4836;
assign w6516 = ~w7614 & ~w3669;
assign w6517 = ~w3418 & ~w7365;
assign w6518 = (w2749 & ~w957) | (w2749 & ~w5346) | (~w957 & ~w5346);
assign w6519 = ~w3521 & ~w45;
assign w6520 = a204 & b204;
assign w6521 = (w4757 & ~w652) | (w4757 & ~w2965) | (~w652 & ~w2965);
assign w6522 = ~w3306 & w926;
assign w6523 = ~w100 & w3242;
assign w6524 = ~w1632 & ~w7648;
assign w6525 = ~w5555 & w7112;
assign w6526 = ~a101 & ~b101;
assign w6527 = (~w2838 & w7582) | (~w2838 & w2456) | (w7582 & w2456);
assign w6528 = ~w779 & w5624;
assign w6529 = ~w145 & ~w1829;
assign w6530 = w5676 & ~w4176;
assign w6531 = (w6467 & w2594) | (w6467 & w1845) | (w2594 & w1845);
assign w6532 = w3591 & w6649;
assign w6533 = (w6100 & w3130) | (w6100 & w2147) | (w3130 & w2147);
assign w6534 = (w5212 & w6872) | (w5212 & w7264) | (w6872 & w7264);
assign w6535 = (~w2367 & w4437) | (~w2367 & w2305) | (w4437 & w2305);
assign w6536 = w174 & w632;
assign w6537 = ~w5445 & w1284;
assign w6538 = ~w4577 & ~w7388;
assign w6539 = ~w2005 & w7364;
assign w6540 = (w6100 & w39) | (w6100 & w4322) | (w39 & w4322);
assign w6541 = (~w3942 & w3253) | (~w3942 & w2561) | (w3253 & w2561);
assign w6542 = ~w5032 & w5965;
assign w6543 = (w1936 & w5688) | (w1936 & w403) | (w5688 & w403);
assign w6544 = w5926 & ~w4822;
assign w6545 = ~w7564 & ~w2996;
assign w6546 = (w5484 & w1842) | (w5484 & w6176) | (w1842 & w6176);
assign w6547 = w6339 & w2142;
assign w6548 = b0 & a0;
assign w6549 = (~w5178 & w2594) | (~w5178 & w6531) | (w2594 & w6531);
assign w6550 = w912 & w3465;
assign w6551 = (~w1493 & w7492) | (~w1493 & w7502) | (w7492 & w7502);
assign w6552 = w975 & ~w3817;
assign w6553 = ~w604 & ~w624;
assign w6554 = w5965 & w4504;
assign w6555 = (w6082 & w582) | (w6082 & w5796) | (w582 & w5796);
assign w6556 = w4072 & ~w2456;
assign w6557 = (w1283 & w4208) | (w1283 & w3762) | (w4208 & w3762);
assign w6558 = a142 & b142;
assign w6559 = (~w5325 & w3861) | (~w5325 & w7505) | (w3861 & w7505);
assign w6560 = (w7506 & w5951) | (w7506 & w2357) | (w5951 & w2357);
assign w6561 = w5461 & w3425;
assign w6562 = ~w391 & w5273;
assign w6563 = (w6253 & w2161) | (w6253 & w4187) | (w2161 & w4187);
assign w6564 = ~w971 & w3716;
assign w6565 = (w1794 & w1039) | (w1794 & ~w6100) | (w1039 & ~w6100);
assign w6566 = (~w4587 & w3172) | (~w4587 & w3065) | (w3172 & w3065);
assign w6567 = ~w141 & ~w5451;
assign w6568 = ~w1328 & w1124;
assign w6569 = w3642 | ~w6714;
assign w6570 = (w6071 & w1549) | (w6071 & w4679) | (w1549 & w4679);
assign w6571 = a21 & b21;
assign w6572 = ~w7452 & ~w3166;
assign w6573 = (~w6663 & w1330) | (~w6663 & w6231) | (w1330 & w6231);
assign w6574 = (w342 & w7013) | (w342 & w1607) | (w7013 & w1607);
assign w6575 = ~w887 & w4564;
assign w6576 = w2389 | w3496;
assign w6577 = (w4068 & ~w6680) | (w4068 & w4262) | (~w6680 & w4262);
assign w6578 = w331 & w4521;
assign w6579 = ~w2229 & w3281;
assign w6580 = (w3986 & w4786) | (w3986 & w7276) | (w4786 & w7276);
assign w6581 = w1786 & w42;
assign w6582 = ~w3482 & ~w351;
assign w6583 = w3161 & ~w2456;
assign w6584 = (w5484 & w1976) | (w5484 & w366) | (w1976 & w366);
assign w6585 = (w5462 & w5790) | (w5462 & w5511) | (w5790 & w5511);
assign w6586 = w499 & w114;
assign w6587 = (~w6630 & w4742) | (~w6630 & w3728) | (w4742 & w3728);
assign w6588 = w2728 & ~w2087;
assign w6589 = (w176 & w271) | (w176 & w5611) | (w271 & w5611);
assign w6590 = w3152 & ~w7348;
assign w6591 = (~w777 & w870) | (~w777 & w5002) | (w870 & w5002);
assign w6592 = w5930 & ~w6450;
assign w6593 = (w6353 & w1738) | (w6353 & w6752) | (w1738 & w6752);
assign w6594 = ~w101 & ~w4330;
assign w6595 = w1758 & ~w2456;
assign w6596 = (~w7604 & w478) | (~w7604 & w1691) | (w478 & w1691);
assign w6597 = ~w6392 & ~w5958;
assign w6598 = (~w860 & ~w1868) | (~w860 & w6062) | (~w1868 & w6062);
assign w6599 = ~w1846 & w6043;
assign w6600 = ~w1343 & ~w4596;
assign w6601 = w2630 & ~w1000;
assign w6602 = (~w2928 & w3703) | (~w2928 & w1047) | (w3703 & w1047);
assign w6603 = (w3116 & w1450) | (w3116 & w6100) | (w1450 & w6100);
assign w6604 = ~w2649 & ~w4204;
assign w6605 = (~w3952 & w2755) | (~w3952 & w7548) | (w2755 & w7548);
assign w6606 = (w64 & ~w1574) | (w64 & w2143) | (~w1574 & w2143);
assign w6607 = ~w3719 & ~w7027;
assign w6608 = w5442 & ~w1137;
assign w6609 = a209 & b209;
assign w6610 = w4180 & w1879;
assign w6611 = (~w5834 & w3234) | (~w5834 & w207) | (w3234 & w207);
assign w6612 = w64 & ~w3435;
assign w6613 = (~w7197 & w5852) | (~w7197 & w5294) | (w5852 & w5294);
assign w6614 = (~w4123 & w5951) | (~w4123 & w7341) | (w5951 & w7341);
assign w6615 = (w166 & w2154) | (w166 & ~w3527) | (w2154 & ~w3527);
assign w6616 = (~w3014 & w2830) | (~w3014 & w6134) | (w2830 & w6134);
assign w6617 = w1608 & w1338;
assign w6618 = (w65 & w4938) | (w65 & w7043) | (w4938 & w7043);
assign w6619 = ~w2816 & w3772;
assign w6620 = ~w4330 & ~w755;
assign w6621 = ~w7598 & w1505;
assign w6622 = (~w3983 & w4117) | (~w3983 & w1418) | (w4117 & w1418);
assign w6623 = (~w6084 & w6378) | (~w6084 & w2211) | (w6378 & w2211);
assign w6624 = (w4006 & w2944) | (w4006 & ~w5395) | (w2944 & ~w5395);
assign w6625 = ~w2872 & w1652;
assign w6626 = w7097 & ~w5276;
assign w6627 = (w3119 & w2775) | (w3119 & w4097) | (w2775 & w4097);
assign w6628 = a35 & b35;
assign w6629 = (w3560 & w2117) | (w3560 & ~w7015) | (w2117 & ~w7015);
assign w6630 = a232 & b232;
assign w6631 = w3102 & ~w847;
assign w6632 = (~w5178 & w5144) | (~w5178 & w6638) | (w5144 & w6638);
assign w6633 = ~w478 & w4922;
assign w6634 = w7042 & ~w973;
assign w6635 = ~w1799 & w3138;
assign w6636 = (w1847 & w911) | (w1847 & w5872) | (w911 & w5872);
assign w6637 = (w1715 & w7327) | (w1715 & ~w3391) | (w7327 & ~w3391);
assign w6638 = ~w3842 & w4373;
assign w6639 = (w7024 & w7443) | (w7024 & w7124) | (w7443 & w7124);
assign w6640 = ~w7581 & ~w6810;
assign w6641 = (w4320 & w1133) | (w4320 & w522) | (w1133 & w522);
assign w6642 = w3136 & ~w1066;
assign w6643 = ~a208 & ~b208;
assign w6644 = w926 & w2699;
assign w6645 = (~w6019 & ~w3078) | (~w6019 & ~w4522) | (~w3078 & ~w4522);
assign w6646 = (w3057 & w6695) | (w3057 & w363) | (w6695 & w363);
assign w6647 = ~w4596 & ~w3446;
assign w6648 = w2650 & ~w5477;
assign w6649 = ~w6936 & ~w7216;
assign w6650 = w5421 & ~w7120;
assign w6651 = (w3867 & w6701) | (w3867 & ~w5871) | (w6701 & ~w5871);
assign w6652 = ~w2197 & ~w4199;
assign w6653 = (w681 & w1798) | (w681 & w3609) | (w1798 & w3609);
assign w6654 = w1149 & ~w3156;
assign w6655 = (w4864 & w4135) | (w4864 & ~w3074) | (w4135 & ~w3074);
assign w6656 = ~a235 & ~b235;
assign w6657 = ~w3136 & w6771;
assign w6658 = ~a107 & ~b107;
assign w6659 = (~w6353 & w266) | (~w6353 & w7066) | (w266 & w7066);
assign w6660 = ~w7381 & w2811;
assign w6661 = (~w1728 & ~w7453) | (~w1728 & w6174) | (~w7453 & w6174);
assign w6662 = (w5522 & w947) | (w5522 & w1889) | (w947 & w1889);
assign w6663 = ~w2708 & w991;
assign w6664 = (w2563 & w3168) | (w2563 & w1082) | (w3168 & w1082);
assign w6665 = (w7379 & w1933) | (w7379 & ~w1881) | (w1933 & ~w1881);
assign w6666 = (w231 & w2431) | (w231 & w485) | (w2431 & w485);
assign w6667 = (w3381 & w3697) | (w3381 & ~w6501) | (w3697 & ~w6501);
assign w6668 = w7345 & ~w2513;
assign w6669 = w3959 & ~w7354;
assign w6670 = (~w4884 & ~w1535) | (~w4884 & w6356) | (~w1535 & w6356);
assign w6671 = w681 & w3266;
assign w6672 = (w7015 & w797) | (w7015 & w1602) | (w797 & w1602);
assign w6673 = ~w3064 & ~w1002;
assign w6674 = w6843 & ~w4300;
assign w6675 = (w7576 & ~w5257) | (w7576 & w5569) | (~w5257 & w5569);
assign w6676 = (w4440 & w5593) | (w4440 & w1743) | (w5593 & w1743);
assign w6677 = (w90 & w4914) | (w90 & w5385) | (w4914 & w5385);
assign w6678 = w2671 & w4222;
assign w6679 = ~w3665 & ~w1429;
assign w6680 = (~w145 & ~w2399) | (~w145 & w3332) | (~w2399 & w3332);
assign w6681 = ~w7027 & w2394;
assign w6682 = ~w6628 & ~w7391;
assign w6683 = a28 & b28;
assign w6684 = ~w3235 & ~w2621;
assign w6685 = ~w1556 & w1605;
assign w6686 = (~w527 & w5512) | (~w527 & w5826) | (w5512 & w5826);
assign w6687 = w6722 | w1555;
assign w6688 = (~w4995 & w6712) | (~w4995 & w1879) | (w6712 & w1879);
assign w6689 = ~w6279 & w2259;
assign w6690 = ~a123 & ~b123;
assign w6691 = (w3952 & w3499) | (w3952 & w5707) | (w3499 & w5707);
assign w6692 = w4849 & w6292;
assign w6693 = ~w2249 & ~w3685;
assign w6694 = (~w3737 & w81) | (~w3737 & w6332) | (w81 & w6332);
assign w6695 = ~w3490 & ~w4132;
assign w6696 = w2188 & ~w303;
assign w6697 = w3101 & ~w6170;
assign w6698 = w5246 & ~w7563;
assign w6699 = (w5007 & w405) | (w5007 & w3) | (w405 & w3);
assign w6700 = ~w1464 & ~w6591;
assign w6701 = (~w5961 & w375) | (~w5961 & w4279) | (w375 & w4279);
assign w6702 = w220 & ~w4200;
assign w6703 = w6992 & ~w2611;
assign w6704 = w2655 & ~w6872;
assign w6705 = w6463 & ~w7530;
assign w6706 = ~w1839 & ~w7196;
assign w6707 = w6009 & ~w5216;
assign w6708 = ~w1999 & ~w832;
assign w6709 = w3909 & ~w1471;
assign w6710 = ~w2903 & w1847;
assign w6711 = (w5484 & w6278) | (w5484 & w4642) | (w6278 & w4642);
assign w6712 = ~w3932 & ~w5732;
assign w6713 = a153 & b153;
assign w6714 = ~w4746 & ~w6713;
assign w6715 = (~w639 & w3344) | (~w639 & w5911) | (w3344 & w5911);
assign w6716 = ~w2084 & ~w4918;
assign w6717 = (~w3708 & w3600) | (~w3708 & w3155) | (w3600 & w3155);
assign w6718 = ~w6265 & w1792;
assign w6719 = ~w6138 & ~w7519;
assign w6720 = ~w4301 & ~w1286;
assign w6721 = ~w1008 & ~w144;
assign w6722 = (w1555 & w84) | (w1555 & w5585) | (w84 & w5585);
assign w6723 = (~w7530 & w6705) | (~w7530 & ~w6439) | (w6705 & ~w6439);
assign w6724 = (w755 & ~w737) | (w755 & w6042) | (~w737 & w6042);
assign w6725 = (w2570 & w7179) | (w2570 & ~w7074) | (w7179 & ~w7074);
assign w6726 = (w155 & w6775) | (w155 & w563) | (w6775 & w563);
assign w6727 = ~w3331 & ~w3422;
assign w6728 = ~w5547 & ~w2137;
assign w6729 = ~w6753 & ~w7056;
assign w6730 = ~w7490 & w1157;
assign w6731 = ~w2140 & w2928;
assign w6732 = (w755 & w6042) | (w755 & ~w101) | (w6042 & ~w101);
assign w6733 = (~w632 & w3847) | (~w632 & ~w264) | (w3847 & ~w264);
assign w6734 = w1758 & ~w3847;
assign w6735 = (w4726 & w19) | (w4726 & ~w3491) | (w19 & ~w3491);
assign w6736 = ~w2741 & w1390;
assign w6737 = (w5807 & w179) | (w5807 & ~w1058) | (w179 & ~w1058);
assign w6738 = (w3057 & w629) | (w3057 & w173) | (w629 & w173);
assign w6739 = (w3509 & w5246) | (w3509 & w3995) | (w5246 & w3995);
assign w6740 = (w5830 & w6862) | (w5830 & w436) | (w6862 & w436);
assign w6741 = (~w6594 & w7453) | (~w6594 & w10) | (w7453 & w10);
assign w6742 = w7271 & w4574;
assign w6743 = (~w3774 & w7561) | (~w3774 & w4712) | (w7561 & w4712);
assign w6744 = (w1379 & w7372) | (w1379 & w5877) | (w7372 & w5877);
assign w6745 = (~w3057 & w3651) | (~w3057 & w2946) | (w3651 & w2946);
assign w6746 = w1607 & w52;
assign w6747 = (w6863 & w1805) | (w6863 & w2312) | (w1805 & w2312);
assign w6748 = ~w4784 & ~w6885;
assign w6749 = (w2707 & ~w730) | (w2707 & ~w1886) | (~w730 & ~w1886);
assign w6750 = (w3788 & w2592) | (w3788 & w1770) | (w2592 & w1770);
assign w6751 = w3524 & w7113;
assign w6752 = ~w6117 & ~w4848;
assign w6753 = ~a238 & ~b238;
assign w6754 = ~w5464 & ~w4350;
assign w6755 = (w2534 & w6311) | (w2534 & w4418) | (w6311 & w4418);
assign w6756 = ~w619 & ~w5891;
assign w6757 = ~a49 & ~b49;
assign w6758 = ~w1196 & ~w5053;
assign w6759 = w5266 & ~w6566;
assign w6760 = a195 & b195;
assign w6761 = w775 & ~w4247;
assign w6762 = (w2540 & w1565) | (w2540 & w3999) | (w1565 & w3999);
assign w6763 = ~w2353 & ~w1368;
assign w6764 = (w3561 & w5516) | (w3561 & w1123) | (w5516 & w1123);
assign w6765 = ~w1154 & ~w4695;
assign w6766 = ~a203 & ~b203;
assign w6767 = w262 & ~w5698;
assign w6768 = ~w4706 & ~w4897;
assign w6769 = (w6602 & w275) | (w6602 & w5886) | (w275 & w5886);
assign w6770 = (~w1137 & w5522) | (~w1137 & w6608) | (w5522 & w6608);
assign w6771 = (w5109 & w2191) | (w5109 & ~w4199) | (w2191 & ~w4199);
assign w6772 = a146 & b146;
assign w6773 = w5604 & w3239;
assign w6774 = a245 & b245;
assign w6775 = (w6906 & w3018) | (w6906 & w7238) | (w3018 & w7238);
assign w6776 = ~a146 & ~b146;
assign w6777 = ~w2600 & w4265;
assign w6778 = (w6724 & w3938) | (w6724 & w6254) | (w3938 & w6254);
assign w6779 = w5883 & ~w7604;
assign w6780 = ~w6872 & w5365;
assign w6781 = ~w3168 & w5446;
assign w6782 = (~w3491 & w5921) | (~w3491 & w5290) | (w5921 & w5290);
assign w6783 = (~w6100 & w496) | (~w6100 & w2155) | (w496 & w2155);
assign w6784 = (~w5655 & w2280) | (~w5655 & w2576) | (w2280 & w2576);
assign w6785 = ~w6439 & ~w7530;
assign w6786 = (w3667 & w1857) | (w3667 & w4558) | (w1857 & w4558);
assign w6787 = (w2401 & w4421) | (w2401 & w6962) | (w4421 & w6962);
assign w6788 = w4465 & w512;
assign w6789 = (w1367 & w4569) | (w1367 & w3574) | (w4569 & w3574);
assign w6790 = ~w6357 & w6953;
assign w6791 = ~a163 & ~b163;
assign w6792 = (w7405 & w6497) | (w7405 & w4200) | (w6497 & w4200);
assign w6793 = (w4283 & w6269) | (w4283 & ~w5291) | (w6269 & ~w5291);
assign w6794 = ~w3385 & w1183;
assign w6795 = ~w6933 & ~w5831;
assign w6796 = ~w1709 & ~w2110;
assign w6797 = (~w1692 & w2033) | (~w1692 & w3738) | (w2033 & w3738);
assign w6798 = (w6385 & w4187) | (w6385 & w5391) | (w4187 & w5391);
assign w6799 = ~w5806 & w3431;
assign w6800 = (w7626 & w5244) | (w7626 & w5706) | (w5244 & w5706);
assign w6801 = w5236 & ~w2579;
assign w6802 = ~w4998 & ~w6458;
assign w6803 = (~w5966 & ~w2380) | (~w5966 & w362) | (~w2380 & w362);
assign w6804 = ~w508 & w7357;
assign w6805 = w4906 & w1497;
assign w6806 = w7243 & ~w2294;
assign w6807 = (w4671 & w2551) | (w4671 & w6722) | (w2551 & w6722);
assign w6808 = w2838 & ~w7352;
assign w6809 = (~w6106 & w2807) | (~w6106 & w2168) | (w2807 & w2168);
assign w6810 = a116 & b116;
assign w6811 = a188 & b188;
assign w6812 = (~w5674 & w6887) | (~w5674 & w1092) | (w6887 & w1092);
assign w6813 = ~w147 & w5277;
assign w6814 = (w5556 & w504) | (w5556 & w540) | (w504 & w540);
assign w6815 = (w6099 & w2994) | (w6099 & w415) | (w2994 & w415);
assign w6816 = (w2871 & w2064) | (w2871 & w7015) | (w2064 & w7015);
assign w6817 = w4145 & ~w3205;
assign w6818 = (w6100 & w914) | (w6100 & w7116) | (w914 & w7116);
assign w6819 = w7048 & ~w3602;
assign w6820 = ~w4477 & ~w3416;
assign w6821 = (w7197 & w1251) | (w7197 & w6616) | (w1251 & w6616);
assign w6822 = ~w3392 & ~w3166;
assign w6823 = (w5963 & w1502) | (w5963 & ~w7015) | (w1502 & ~w7015);
assign w6824 = (w6100 & w5697) | (w6100 & w3564) | (w5697 & w3564);
assign w6825 = (w4517 & w360) | (w4517 & ~w2965) | (w360 & ~w2965);
assign w6826 = (~w5655 & w6743) | (~w5655 & w2713) | (w6743 & w2713);
assign w6827 = ~w1206 & w4892;
assign w6828 = ~w757 & ~w2909;
assign w6829 = ~w6626 & ~w2333;
assign w6830 = w6688 & w7107;
assign w6831 = w2417 | w4962;
assign w6832 = ~w6803 & w6748;
assign w6833 = ~w2172 & w5412;
assign w6834 = ~w3064 & w6758;
assign w6835 = w4672 & w4457;
assign w6836 = w2494 & ~w4997;
assign w6837 = w3061 & w4199;
assign w6838 = (~w5674 & w457) | (~w5674 & w1022) | (w457 & w1022);
assign w6839 = ~w4898 & ~w5820;
assign w6840 = (w1598 & w2847) | (w1598 & w4770) | (w2847 & w4770);
assign w6841 = w43 & ~w5611;
assign w6842 = ~w6634 & w4603;
assign w6843 = w4035 & ~w4300;
assign w6844 = (w6195 & w5194) | (w6195 & w3608) | (w5194 & w3608);
assign w6845 = (~w7158 & ~w139) | (~w7158 & ~w1626) | (~w139 & ~w1626);
assign w6846 = (~w1544 & w4296) | (~w1544 & w4418) | (w4296 & w4418);
assign w6847 = w3677 & w1134;
assign w6848 = w1591 & ~w4146;
assign w6849 = ~w5622 & ~w6455;
assign w6850 = w6057 & ~w1775;
assign w6851 = ~w2521 & ~w7391;
assign w6852 = ~w314 & w1759;
assign w6853 = (~w7256 & w156) | (~w7256 & w4199) | (w156 & w4199);
assign w6854 = a117 & b117;
assign w6855 = (~w6490 & w3700) | (~w6490 & w180) | (w3700 & w180);
assign w6856 = (w1516 & w5142) | (w1516 & w4472) | (w5142 & w4472);
assign w6857 = ~w7528 & w7605;
assign w6858 = (~w5325 & w7284) | (~w5325 & w845) | (w7284 & w845);
assign w6859 = ~w4715 & ~w7206;
assign w6860 = ~w3616 & w1137;
assign w6861 = ~w7308 & ~w7641;
assign w6862 = w4637 & ~w6658;
assign w6863 = ~w1923 & w7201;
assign w6864 = (w5178 & w7261) | (w5178 & w6491) | (w7261 & w6491);
assign w6865 = (w493 & w6542) | (w493 & ~w1285) | (w6542 & ~w1285);
assign w6866 = w4918 & ~w7581;
assign w6867 = (w6151 & w4080) | (w6151 & w4513) | (w4080 & w4513);
assign w6868 = w554 & ~w235;
assign w6869 = (~w3580 & w919) | (~w3580 & ~w2582) | (w919 & ~w2582);
assign w6870 = ~w6335 & ~w7127;
assign w6871 = ~w5499 & w2938;
assign w6872 = (w1607 & ~w174) | (w1607 & ~w1608) | (~w174 & ~w1608);
assign w6873 = (~w1607 & w174) | (~w1607 & w1608) | (w174 & w1608);
assign w6874 = w5266 & ~w5430;
assign w6875 = (w4102 & w1012) | (w4102 & w992) | (w1012 & w992);
assign w6876 = ~w6558 & w5350;
assign w6877 = w714 & w2426;
assign w6878 = w1743 & ~w4182;
assign w6879 = ~w3252 & ~w5350;
assign w6880 = (w7386 & w5925) | (w7386 & w5325) | (w5925 & w5325);
assign w6881 = ~w3868 & w3014;
assign w6882 = (w5419 & w6264) | (w5419 & w5487) | (w6264 & w5487);
assign w6883 = ~w2846 & ~w2243;
assign w6884 = a50 & b50;
assign w6885 = ~w2846 & ~w1621;
assign w6886 = ~w6526 & w1886;
assign w6887 = w1389 & ~w7283;
assign w6888 = ~w1877 & ~w2864;
assign w6889 = (w6920 & w7147) | (w6920 & w6373) | (w7147 & w6373);
assign w6890 = w2238 & ~w5550;
assign w6891 = w6465 & ~w544;
assign w6892 = ~w5464 & ~w990;
assign w6893 = ~w7397 & w5744;
assign w6894 = (~w2456 & ~w412) | (~w2456 & w7474) | (~w412 & w7474);
assign w6895 = w3044 & w2968;
assign w6896 = w1021 & ~w3840;
assign w6897 = ~w4551 & w3501;
assign w6898 = ~w7527 & ~w3073;
assign w6899 = ~w4335 & ~w6995;
assign w6900 = w7242 & w6644;
assign w6901 = w2740 & w1888;
assign w6902 = (~w6424 & w2529) | (~w6424 & w6603) | (w2529 & w6603);
assign w6903 = (~w523 & w1456) | (~w523 & w4074) | (w1456 & w4074);
assign w6904 = (~w7546 & w3984) | (~w7546 & w5635) | (w3984 & w5635);
assign w6905 = ~w1176 & w3166;
assign w6906 = (w3136 & w7490) | (w3136 & w4815) | (w7490 & w4815);
assign w6907 = ~w2197 & ~w4056;
assign w6908 = (w7300 & w565) | (w7300 & w4880) | (w565 & w4880);
assign w6909 = (w5834 & w1075) | (w5834 & w6707) | (w1075 & w6707);
assign w6910 = (~w7450 & w3196) | (~w7450 & w7423) | (w3196 & w7423);
assign w6911 = ~w1923 & ~w7146;
assign w6912 = a139 & b139;
assign w6913 = (~w7097 & w6965) | (~w7097 & w1886) | (w6965 & w1886);
assign w6914 = (w5537 & w1328) | (w5537 & w2313) | (w1328 & w2313);
assign w6915 = (~w777 & w3443) | (~w777 & w498) | (w3443 & w498);
assign w6916 = (w5703 & w4858) | (w5703 & w5768) | (w4858 & w5768);
assign w6917 = w3152 & w1031;
assign w6918 = (~w7528 & w5710) | (~w7528 & w2580) | (w5710 & w2580);
assign w6919 = (~w2513 & w6668) | (~w2513 & w6712) | (w6668 & w6712);
assign w6920 = ~w3366 & w583;
assign w6921 = w3286 & w3062;
assign w6922 = ~w6458 & ~w2450;
assign w6923 = ~w577 & w4089;
assign w6924 = ~w7546 & w703;
assign w6925 = (w6557 & w5844) | (w6557 & w3852) | (w5844 & w3852);
assign w6926 = (w5178 & w5087) | (w5178 & w5928) | (w5087 & w5928);
assign w6927 = ~w3965 & ~w5503;
assign w6928 = (~w1804 & w238) | (~w1804 & w5430) | (w238 & w5430);
assign w6929 = (w7072 & w7148) | (w7072 & w5031) | (w7148 & w5031);
assign w6930 = w2001 & w7407;
assign w6931 = ~w1709 & ~w6088;
assign w6932 = (~w1535 & w682) | (~w1535 & w5654) | (w682 & w5654);
assign w6933 = (w2628 & w5178) | (w2628 & w4432) | (w5178 & w4432);
assign w6934 = (w5325 & w7117) | (w5325 & w2079) | (w7117 & w2079);
assign w6935 = ~w1883 & ~w3217;
assign w6936 = ~a108 & ~b108;
assign w6937 = w2830 & ~w3903;
assign w6938 = (~w6420 & w3857) | (~w6420 & w1397) | (w3857 & w1397);
assign w6939 = ~w6912 & ~w5499;
assign w6940 = ~w5605 & ~w1585;
assign w6941 = (~w4143 & w5535) | (~w4143 & w2926) | (w5535 & w2926);
assign w6942 = ~w6526 & ~w5276;
assign w6943 = (w3057 & w5258) | (w3057 & w5847) | (w5258 & w5847);
assign w6944 = w2257 & w6099;
assign w6945 = w7102 & w6174;
assign w6946 = ~w5029 & ~w2593;
assign w6947 = (w2847 & w2825) | (w2847 & w6725) | (w2825 & w6725);
assign w6948 = (w2332 & w1043) | (w2332 & ~w4199) | (w1043 & ~w4199);
assign w6949 = ~w1315 | w3997;
assign w6950 = w3489 | ~w5734;
assign w6951 = (w4143 & w1019) | (w4143 & w4120) | (w1019 & w4120);
assign w6952 = ~w2196 & ~w4535;
assign w6953 = ~w618 & w6883;
assign w6954 = ~w4998 & w7256;
assign w6955 = w1563 & ~w665;
assign w6956 = w6854 & ~w6594;
assign w6957 = w7647 & w6100;
assign w6958 = ~w3719 & w6681;
assign w6959 = w3901 & w6216;
assign w6960 = ~w4325 & ~w6634;
assign w6961 = w663 | ~w6524;
assign w6962 = w2912 & w1549;
assign w6963 = w3166 & ~w3905;
assign w6964 = w4759 & ~w3072;
assign w6965 = w5616 & ~w7097;
assign w6966 = (w1886 & w4280) | (w1886 & w506) | (w4280 & w506);
assign w6967 = (~w2021 & w4626) | (~w2021 & w5231) | (w4626 & w5231);
assign w6968 = ~w2566 & w6705;
assign w6969 = ~w5463 & ~w1660;
assign w6970 = ~w5277 & ~w1325;
assign w6971 = ~w1271 & w3719;
assign w6972 = (~w434 & ~w174) | (~w434 & w1520) | (~w174 & w1520);
assign w6973 = ~w3428 & ~w773;
assign w6974 = ~w4438 & w728;
assign w6975 = (w6480 & w5108) | (w6480 & w2101) | (w5108 & w2101);
assign w6976 = w6385 & ~w476;
assign w6977 = w3167 & ~w5008;
assign w6978 = w827 & ~w3527;
assign w6979 = ~a88 & ~b88;
assign w6980 = ~a200 & ~b200;
assign w6981 = a48 & b48;
assign w6982 = w775 & w2311;
assign w6983 = w5442 & ~w2913;
assign w6984 = w7399 & ~w7127;
assign w6985 = ~w3826 & w3987;
assign w6986 = ~w2987 & w7385;
assign w6987 = (~w5655 & w3879) | (~w5655 & w3151) | (w3879 & w3151);
assign w6988 = (~w4392 & w1533) | (~w4392 & w6472) | (w1533 & w6472);
assign w6989 = (w527 & w6564) | (w527 & w657) | (w6564 & w657);
assign w6990 = ~w539 & ~w5260;
assign w6991 = ~w6634 & w407;
assign w6992 = ~a199 & ~b199;
assign w6993 = (w401 & w5761) | (w401 & w5511) | (w5761 & w5511);
assign w6994 = a135 & b135;
assign w6995 = (~w6945 & w1784) | (~w6945 & w4113) | (w1784 & w4113);
assign w6996 = (w5035 & ~w5933) | (w5035 & w3357) | (~w5933 & w3357);
assign w6997 = (w7405 & w6497) | (w7405 & w1133) | (w6497 & w1133);
assign w6998 = ~w4251 & w3819;
assign w6999 = ~w7147 & w5662;
assign w7000 = ~a145 & ~b145;
assign w7001 = (w3774 & w2716) | (w3774 & w7619) | (w2716 & w7619);
assign w7002 = ~w3455 & w3716;
assign w7003 = w6031 & w6174;
assign w7004 = (w398 & w3369) | (w398 & ~w5403) | (w3369 & ~w5403);
assign w7005 = a230 & b230;
assign w7006 = (w4287 & w2301) | (w4287 & w7339) | (w2301 & w7339);
assign w7007 = (~w6965 & w5118) | (~w6965 & w4904) | (w5118 & w4904);
assign w7008 = (w7118 & ~w5257) | (w7118 & w1944) | (~w5257 & w1944);
assign w7009 = (w1515 & w4320) | (w1515 & w4200) | (w4320 & w4200);
assign w7010 = ~w4822 & ~w1827;
assign w7011 = (~w5834 & w6948) | (~w5834 & w2223) | (w6948 & w2223);
assign w7012 = ~a226 & ~b226;
assign w7013 = (w2112 & w3095) | (w2112 & w2989) | (w3095 & w2989);
assign w7014 = ~w6545 & w1727;
assign w7015 = (~w7238 & w5429) | (~w7238 & w2787) | (w5429 & w2787);
assign w7016 = w3701 & w5842;
assign w7017 = w56 & ~w7312;
assign w7018 = w2655 & w167;
assign w7019 = (~w1272 & w1974) | (~w1272 & ~w2966) | (w1974 & ~w2966);
assign w7020 = ~w604 & ~w6281;
assign w7021 = (w3808 & ~w2517) | (w3808 & w3912) | (~w2517 & w3912);
assign w7022 = ~w7365 & ~w527;
assign w7023 = (~w5178 & w7017) | (~w5178 & w7282) | (w7017 & w7282);
assign w7024 = (~w3490 & w475) | (~w3490 & w6377) | (w475 & w6377);
assign w7025 = (w2639 & w5097) | (w2639 & w7015) | (w5097 & w7015);
assign w7026 = ~a91 & ~b91;
assign w7027 = a162 & b162;
assign w7028 = (w3057 & w5138) | (w3057 & w6901) | (w5138 & w6901);
assign w7029 = (~w999 & w6920) | (~w999 & w7129) | (w6920 & w7129);
assign w7030 = ~w2798 & w3391;
assign w7031 = w2066 & ~w2649;
assign w7032 = ~w7486 & ~w3033;
assign w7033 = (~w5178 & w6694) | (~w5178 & w4910) | (w6694 & w4910);
assign w7034 = (w6415 & ~w5058) | (w6415 & w4464) | (~w5058 & w4464);
assign w7035 = w7390 & ~w3096;
assign w7036 = (~w5121 & ~w3774) | (~w5121 & w900) | (~w3774 & w900);
assign w7037 = ~w2740 & ~w1888;
assign w7038 = (~w7453 & w3010) | (~w7453 & w6111) | (w3010 & w6111);
assign w7039 = (~w6106 & w5753) | (~w6106 & w4055) | (w5753 & w4055);
assign w7040 = (~w1006 & w6862) | (~w1006 & w3249) | (w6862 & w3249);
assign w7041 = (w3774 & w1239) | (w3774 & w949) | (w1239 & w949);
assign w7042 = ~a193 & ~b193;
assign w7043 = w7199 & w6650;
assign w7044 = a216 & b216;
assign w7045 = (w3929 & w1822) | (w3929 & w5403) | (w1822 & w5403);
assign w7046 = (~w999 & w7129) | (~w999 & w6889) | (w7129 & w6889);
assign w7047 = w424 & ~w6791;
assign w7048 = w7271 & ~w3602;
assign w7049 = w1756 & ~w2353;
assign w7050 = (w882 & w7189) | (w882 & w1122) | (w7189 & w1122);
assign w7051 = ~w3855 & ~w3435;
assign w7052 = (w5430 & w4720) | (w5430 & w6428) | (w4720 & w6428);
assign w7053 = w4348 & ~w4749;
assign w7054 = w2796 & ~w139;
assign w7055 = w4622 | w138;
assign w7056 = ~a239 & ~b239;
assign w7057 = (w770 & w3283) | (w770 & w4267) | (w3283 & w4267);
assign w7058 = w4784 & w6885;
assign w7059 = ~w1524 & ~w952;
assign w7060 = w4140 & w3863;
assign w7061 = (~w6911 & w6271) | (~w6911 & w3888) | (w6271 & w3888);
assign w7062 = ~w6614 & ~w2740;
assign w7063 = (w6100 & w3925) | (w6100 & w4408) | (w3925 & w4408);
assign w7064 = (w4995 & w7175) | (w4995 & w7463) | (w7175 & w7463);
assign w7065 = w3200 & ~w2520;
assign w7066 = (w6061 & w7610) | (w6061 & w24) | (w7610 & w24);
assign w7067 = (~w4875 & w6844) | (~w4875 & w1668) | (w6844 & w1668);
assign w7068 = (w3306 & ~w1165) | (w3306 & ~w3205) | (~w1165 & ~w3205);
assign w7069 = ~w3559 & ~w89;
assign w7070 = w6383 & ~w2707;
assign w7071 = w2526 & w5726;
assign w7072 = (w52 & ~w174) | (w52 & w6746) | (~w174 & w6746);
assign w7073 = ~w3918 & ~w4409;
assign w7074 = (~w2124 & w206) | (~w2124 & w4114) | (w206 & w4114);
assign w7075 = ~w4334 & ~w462;
assign w7076 = (w2791 & w3908) | (w2791 & w5680) | (w3908 & w5680);
assign w7077 = w6399 & w1665;
assign w7078 = ~w1756 & w1911;
assign w7079 = (~w1954 & w6329) | (~w1954 & w7563) | (w6329 & w7563);
assign w7080 = ~w6539 & w3224;
assign w7081 = w6397 & ~w3819;
assign w7082 = ~w5958 & ~w887;
assign w7083 = ~w534 & w3204;
assign w7084 = (w4323 & w2950) | (w4323 & ~w5511) | (w2950 & ~w5511);
assign w7085 = (w3017 & w7100) | (w3017 & ~w7000) | (w7100 & ~w7000);
assign w7086 = (w3784 & w2502) | (w3784 & w2876) | (w2502 & w2876);
assign w7087 = w2542 & w1836;
assign w7088 = (w5178 & w7488) | (w5178 & w3920) | (w7488 & w3920);
assign w7089 = (w3318 & w7287) | (w3318 & w6400) | (w7287 & w6400);
assign w7090 = ~w2456 & w174;
assign w7091 = w1607 & w2456;
assign w7092 = w7357 & w2873;
assign w7093 = ~w2127 & w5808;
assign w7094 = ~w732 & ~w5784;
assign w7095 = (w902 & ~w3774) | (w902 & w725) | (~w3774 & w725);
assign w7096 = (w5834 & w2387) | (w5834 & w4826) | (w2387 & w4826);
assign w7097 = ~a100 & ~b100;
assign w7098 = w6057 & ~w4197;
assign w7099 = w6125 & w2209;
assign w7100 = w7190 & w3017;
assign w7101 = w1716 & ~w5538;
assign w7102 = w400 & w5627;
assign w7103 = (w340 & w5178) | (w340 & w1651) | (w5178 & w1651);
assign w7104 = ~w4426 & ~w5936;
assign w7105 = (~w5478 & w3957) | (~w5478 & w7574) | (w3957 & w7574);
assign w7106 = ~w5958 & ~w4564;
assign w7107 = w4180 & ~w434;
assign w7108 = (w5325 & w1892) | (w5325 & w3743) | (w1892 & w3743);
assign w7109 = (w5871 & w5656) | (w5871 & w1653) | (w5656 & w1653);
assign w7110 = ~w5066 & w3557;
assign w7111 = ~w142 & ~w5251;
assign w7112 = (~w5464 & ~w6195) | (~w5464 & w6892) | (~w6195 & w6892);
assign w7113 = ~w3019 & w6351;
assign w7114 = w6298 & w1748;
assign w7115 = (w6177 & w4077) | (w6177 & w3297) | (w4077 & w3297);
assign w7116 = (w6082 & w2337) | (w6082 & w5372) | (w2337 & w5372);
assign w7117 = (~w367 & w3091) | (~w367 & w2256) | (w3091 & w2256);
assign w7118 = ~w7634 & ~w2182;
assign w7119 = w1878 & w7008;
assign w7120 = w2011 & w1574;
assign w7121 = w1915 & w2837;
assign w7122 = ~w174 & w2297;
assign w7123 = (w6644 & w778) | (w6644 & w6900) | (w778 & w6900);
assign w7124 = w5403 & w7090;
assign w7125 = (~w3318 & w4755) | (~w3318 & w851) | (w4755 & w851);
assign w7126 = (w2294 & w6451) | (w2294 & w3079) | (w6451 & w3079);
assign w7127 = a113 & b113;
assign w7128 = (w7255 & w5850) | (w7255 & w7043) | (w5850 & w7043);
assign w7129 = ~w2327 & ~w999;
assign w7130 = (w6248 & w3277) | (w6248 & ~w3391) | (w3277 & ~w3391);
assign w7131 = (w6019 & w3683) | (w6019 & w1078) | (w3683 & w1078);
assign w7132 = w322 & w759;
assign w7133 = ~w2221 & w5986;
assign w7134 = ~w554 & w4647;
assign w7135 = (~w2627 & w5139) | (~w2627 & w4783) | (w5139 & w4783);
assign w7136 = (w5225 & w3410) | (w5225 & ~w484) | (w3410 & ~w484);
assign w7137 = ~a148 & ~b148;
assign w7138 = ~w147 & ~w195;
assign w7139 = ~w6303 & ~w774;
assign w7140 = (~w615 & w4170) | (~w615 & w345) | (w4170 & w345);
assign w7141 = (~w6181 & w2401) | (~w6181 & w1414) | (w2401 & w1414);
assign w7142 = ~a201 & ~b201;
assign w7143 = ~w3587 & ~w3736;
assign w7144 = w6499 & ~w2013;
assign w7145 = ~w2460 & w4333;
assign w7146 = a154 & b154;
assign w7147 = ~w1718 & w4852;
assign w7148 = (w2112 & w962) | (w2112 & w7110) | (w962 & w7110);
assign w7149 = ~w6916 & ~w5896;
assign w7150 = ~w182 & ~w6628;
assign w7151 = ~w5693 & ~w7127;
assign w7152 = w6708 & w2293;
assign w7153 = (~w5178 & w4874) | (~w5178 & w932) | (w4874 & w932);
assign w7154 = (~w6922 & w2603) | (~w6922 & w5199) | (w2603 & w5199);
assign w7155 = (w484 & w7015) | (w484 & ~w5291) | (w7015 & ~w5291);
assign w7156 = w6660 | ~w4891;
assign w7157 = (~w4564 & ~w1455) | (~w4564 & w4742) | (~w1455 & w4742);
assign w7158 = ~w1279 & w6041;
assign w7159 = (~w7063 & w1677) | (~w7063 & w326) | (w1677 & w326);
assign w7160 = w2078 | ~w3108;
assign w7161 = w6459 & w198;
assign w7162 = (~w6927 & w4337) | (~w6927 & w3160) | (w4337 & w3160);
assign w7163 = (~w6222 & w4156) | (~w6222 & w3488) | (w4156 & w3488);
assign w7164 = w4340 & ~w7015;
assign w7165 = w4526 & w4875;
assign w7166 = (~w5486 & w3363) | (~w5486 & w6606) | (w3363 & w6606);
assign w7167 = (~w5178 & w2802) | (~w5178 & w3042) | (w2802 & w3042);
assign w7168 = (w6535 & w1674) | (w6535 & w7238) | (w1674 & w7238);
assign w7169 = w701 & ~w1377;
assign w7170 = (~w7015 & w3037) | (~w7015 & w4022) | (w3037 & w4022);
assign w7171 = (w2792 & w3986) | (w2792 & w2673) | (w3986 & w2673);
assign w7172 = ~w6658 & ~w4643;
assign w7173 = w4975 & w5143;
assign w7174 = ~w3677 & ~w2820;
assign w7175 = w4072 & ~w6712;
assign w7176 = (w3335 & w4450) | (w3335 & ~w4199) | (w4450 & ~w4199);
assign w7177 = (w506 & w6886) | (w506 & w6000) | (w6886 & w6000);
assign w7178 = w2216 & ~w2718;
assign w7179 = w5978 & ~w1731;
assign w7180 = ~w6935 & ~w913;
assign w7181 = w5012 & w2217;
assign w7182 = ~w2257 & w4694;
assign w7183 = ~w7026 & ~w2688;
assign w7184 = (w6424 & w6589) | (w6424 & w2164) | (w6589 & w2164);
assign w7185 = ~w3219 & w7592;
assign w7186 = (w5834 & w3502) | (w5834 & w4703) | (w3502 & w4703);
assign w7187 = w6663 & w2495;
assign w7188 = w3096 & ~w3450;
assign w7189 = (w5974 & w7187) | (w5974 & w7332) | (w7187 & w7332);
assign w7190 = a145 & b145;
assign w7191 = (~w4314 & w1747) | (~w4314 & w1270) | (w1747 & w1270);
assign w7192 = ~w2222 | ~w3984;
assign w7193 = ~w4392 & w1533;
assign w7194 = ~w7150 & w1519;
assign w7195 = w4156 & ~w6222;
assign w7196 = w5665 & ~w5295;
assign w7197 = (w3224 & w4337) | (w3224 & w7080) | (w4337 & w7080);
assign w7198 = (~w4641 & w5130) | (~w4641 & w5857) | (w5130 & w5857);
assign w7199 = ~w3866 & w4850;
assign w7200 = (~w5178 & w4311) | (~w5178 & w115) | (w4311 & w115);
assign w7201 = ~w4176 & ~w4746;
assign w7202 = ~w3569 & w5148;
assign w7203 = w3994 & w7262;
assign w7204 = ~w5230 & ~w1066;
assign w7205 = w6353 & w5113;
assign w7206 = (w6945 & w408) | (w6945 & w6121) | (w408 & w6121);
assign w7207 = (w5871 & w217) | (w5871 & w7585) | (w217 & w7585);
assign w7208 = ~w255 & ~w3170;
assign w7209 = w2798 & ~w6254;
assign w7210 = (w7003 & w1777) | (w7003 & w265) | (w1777 & w265);
assign w7211 = ~w1184 & ~w218;
assign w7212 = w7384 & ~w444;
assign w7213 = ~a32 & ~b32;
assign w7214 = ~w7289 & ~w4674;
assign w7215 = w2725 & ~w1967;
assign w7216 = a108 & b108;
assign w7217 = (w3427 & w1687) | (w3427 & ~w6100) | (w1687 & ~w6100);
assign w7218 = ~w6571 & w1384;
assign w7219 = ~a188 & ~b188;
assign w7220 = ~w3176 & ~w5357;
assign w7221 = ~a117 & ~b117;
assign w7222 = w1849 & ~w3433;
assign w7223 = ~w151 & ~w5783;
assign w7224 = (~w435 & ~w2453) | (~w435 & w5629) | (~w2453 & w5629);
assign w7225 = (~w2624 & w6307) | (~w2624 & w2890) | (w6307 & w2890);
assign w7226 = ~w1728 & ~w6854;
assign w7227 = ~w2751 & w3869;
assign w7228 = ~w63 & ~w4765;
assign w7229 = (w6724 & w3938) | (w6724 & ~w6174) | (w3938 & ~w6174);
assign w7230 = (w2454 & w2828) | (w2454 & ~w5098) | (w2828 & ~w5098);
assign w7231 = ~w5466 & w5721;
assign w7232 = ~w5486 & w5808;
assign w7233 = ~w6660 & w2793;
assign w7234 = (~w4651 & w5553) | (~w4651 & ~w2725) | (w5553 & ~w2725);
assign w7235 = (~w3269 & w2049) | (~w3269 & ~w4922) | (w2049 & ~w4922);
assign w7236 = (w3311 & w4423) | (w3311 & w6100) | (w4423 & w6100);
assign w7237 = (~w7256 & w156) | (~w7256 & w7238) | (w156 & w7238);
assign w7238 = (w169 & ~w5419) | (w169 & w6443) | (~w5419 & w6443);
assign w7239 = ~w5194 & w1990;
assign w7240 = (~w2542 & w4201) | (~w2542 & w0) | (w4201 & w0);
assign w7241 = (w4652 & w6005) | (w4652 & ~w7238) | (w6005 & ~w7238);
assign w7242 = ~w6526 & w4425;
assign w7243 = ~w7213 & ~w642;
assign w7244 = (w4223 & w1613) | (w4223 & ~w5611) | (w1613 & ~w5611);
assign w7245 = (~w5522 & w2635) | (~w5522 & w5935) | (w2635 & w5935);
assign w7246 = w4922 & ~w7332;
assign w7247 = ~w803 & ~w4407;
assign w7248 = w3573 & w47;
assign w7249 = (~w7306 & w445) | (~w7306 & w1446) | (w445 & w1446);
assign w7250 = (w3017 & w7100) | (w3017 & w3630) | (w7100 & w3630);
assign w7251 = ~w796 & ~w1567;
assign w7252 = ~w7010 & ~w6600;
assign w7253 = w7010 & w6809;
assign w7254 = (w7554 & w4705) | (w7554 & w6573) | (w4705 & w6573);
assign w7255 = ~w950 & w6301;
assign w7256 = ~w4612 & ~w6304;
assign w7257 = w2270 & ~w3490;
assign w7258 = ~w1649 & w4092;
assign w7259 = w5246 & ~w6355;
assign w7260 = w6689 & ~w1817;
assign w7261 = (w5484 & w4048) | (w5484 & w4189) | (w4048 & w4189);
assign w7262 = ~w6161 & ~w1975;
assign w7263 = ~w4665 & w2952;
assign w7264 = (w5212 & w3953) | (w5212 & w4195) | (w3953 & w4195);
assign w7265 = a191 & b191;
assign w7266 = ~w5958 & ~w434;
assign w7267 = w4922 & w7113;
assign w7268 = ~w7302 & ~w4467;
assign w7269 = (~w4680 & w6230) | (~w4680 & w3770) | (w6230 & w3770);
assign w7270 = ~w4268 & ~w3803;
assign w7271 = ~a2 & ~b2;
assign w7272 = ~w4191 & w6719;
assign w7273 = ~w4497 & ~w651;
assign w7274 = (~w5178 & w6302) | (~w5178 & w5470) | (w6302 & w5470);
assign w7275 = ~w1570 & ~w3014;
assign w7276 = (w4786 & ~w7187) | (w4786 & w3354) | (~w7187 & w3354);
assign w7277 = ~w2221 & w3134;
assign w7278 = a181 & b181;
assign w7279 = ~w332 & w4603;
assign w7280 = (w3311 & w4423) | (w3311 & w6254) | (w4423 & w6254);
assign w7281 = (~w5257 & w6347) | (~w5257 & w4561) | (w6347 & w4561);
assign w7282 = (w6467 & w7017) | (w6467 & w3352) | (w7017 & w3352);
assign w7283 = ~w335 & ~w2255;
assign w7284 = w1355 & w6630;
assign w7285 = w757 & w6831;
assign w7286 = w3836 & w6822;
assign w7287 = (~w563 & w5088) | (~w563 & w6282) | (w5088 & w6282);
assign w7288 = w6935 & w1424;
assign w7289 = ~a236 & ~b236;
assign w7290 = (w4967 & w4722) | (w4967 & w1400) | (w4722 & w1400);
assign w7291 = ~a124 & ~b124;
assign w7292 = ~w1057 & w4692;
assign w7293 = (~w3033 & w2220) | (~w3033 & ~w2097) | (w2220 & ~w2097);
assign w7294 = ~w3096 & ~w3176;
assign w7295 = (w4756 & w4304) | (w4756 & w563) | (w4304 & w563);
assign w7296 = w6758 & w6673;
assign w7297 = (~w5257 & w4303) | (~w5257 & w3776) | (w4303 & w3776);
assign w7298 = (w3952 & w1119) | (w3952 & w2240) | (w1119 & w2240);
assign w7299 = ~a84 & ~b84;
assign w7300 = (w388 & w734) | (w388 & w4156) | (w734 & w4156);
assign w7301 = w3503 & w989;
assign w7302 = ~a41 & ~b41;
assign w7303 = (w4199 & w7238) | (w4199 & w563) | (w7238 & w563);
assign w7304 = w1911 & ~w7049;
assign w7305 = ~w6346 & ~w4499;
assign w7306 = (~w2806 & w4159) | (~w2806 & w5006) | (w4159 & w5006);
assign w7307 = w2914 & ~w1682;
assign w7308 = w3306 & ~w3799;
assign w7309 = ~w523 & ~w7451;
assign w7310 = ~w4146 & w215;
assign w7311 = ~w618 & ~w4784;
assign w7312 = ~w516 & ~w7572;
assign w7313 = w1957 & ~w424;
assign w7314 = w3166 & ~w3359;
assign w7315 = (~w5944 & w5175) | (~w5944 & w140) | (w5175 & w140);
assign w7316 = ~w6634 & ~w4000;
assign w7317 = ~w1160 & ~w6684;
assign w7318 = (w6254 & w10) | (w6254 & w3329) | (w10 & w3329);
assign w7319 = w7432 & w673;
assign w7320 = ~w3157 & ~w2605;
assign w7321 = ~w2741 & w5789;
assign w7322 = ~w4891 & w1328;
assign w7323 = ~w3905 & ~w6822;
assign w7324 = w4496 & w6504;
assign w7325 = (w5871 & w2581) | (w5871 & ~w1004) | (w2581 & ~w1004);
assign w7326 = ~w1241 & ~w7420;
assign w7327 = w1554 & w151;
assign w7328 = (~w3319 & w4840) | (~w3319 & w620) | (w4840 & w620);
assign w7329 = w2378 & w2406;
assign w7330 = ~w4680 & w2703;
assign w7331 = (~w639 & w5804) | (~w639 & w1478) | (w5804 & w1478);
assign w7332 = ~w3207 & ~w5289;
assign w7333 = w6870 & w3492;
assign w7334 = w5529 & w6418;
assign w7335 = (w3983 & w2936) | (w3983 & w2505) | (w2936 & w2505);
assign w7336 = w1129 & w7442;
assign w7337 = (~w7197 & w4328) | (~w7197 & w6141) | (w4328 & w6141);
assign w7338 = w1756 & ~w3266;
assign w7339 = ~w3643 & ~w1891;
assign w7340 = (~w1565 & w5798) | (~w1565 & w3598) | (w5798 & w3598);
assign w7341 = ~w1735 & ~w4123;
assign w7342 = ~w2283 & ~w6942;
assign w7343 = w2829 & w2289;
assign w7344 = w2131 & ~w6566;
assign w7345 = a228 & b228;
assign w7346 = ~w1974 & ~w3607;
assign w7347 = (~w6252 & w4342) | (~w6252 & ~w512) | (w4342 & ~w512);
assign w7348 = (~w1272 & w1974) | (~w1272 & w4418) | (w1974 & w4418);
assign w7349 = w1371 & ~w7486;
assign w7350 = ~a85 & ~b85;
assign w7351 = (w4697 & ~w3986) | (w4697 & w1177) | (~w3986 & w1177);
assign w7352 = w1591 & ~w385;
assign w7353 = (w1732 & w1072) | (w1732 & w3488) | (w1072 & w3488);
assign w7354 = w3282 & w7486;
assign w7355 = ~w2667 & w1109;
assign w7356 = ~w2558 & w1714;
assign w7357 = ~w7302 & ~w4476;
assign w7358 = (~w1304 & w2340) | (~w1304 & w873) | (w2340 & w873);
assign w7359 = (w3134 & w5901) | (w3134 & w7277) | (w5901 & w7277);
assign w7360 = w438 & ~w6513;
assign w7361 = w4843 & ~w1866;
assign w7362 = ~w1196 & w5881;
assign w7363 = ~a40 & ~b40;
assign w7364 = ~w2066 & ~w3965;
assign w7365 = a180 & b180;
assign w7366 = ~w2513 & ~w856;
assign w7367 = (w4510 & w5535) | (w4510 & w6677) | (w5535 & w6677);
assign w7368 = w4002 & w6426;
assign w7369 = (~w3719 & w5996) | (~w3719 & w4620) | (w5996 & w4620);
assign w7370 = (~w2267 & w188) | (~w2267 & w1552) | (w188 & w1552);
assign w7371 = ~w5827 & w7014;
assign w7372 = w2380 & ~w3500;
assign w7373 = a31 & b31;
assign w7374 = (~w1936 & w7077) | (~w1936 & w4413) | (w7077 & w4413);
assign w7375 = (~w5655 & w3792) | (~w5655 & w355) | (w3792 & w355);
assign w7376 = w6681 & ~w2993;
assign w7377 = (w6646 & w1150) | (w6646 & ~w5385) | (w1150 & ~w5385);
assign w7378 = w2811 & w4852;
assign w7379 = (w5226 & w4329) | (w5226 & w6401) | (w4329 & w6401);
assign w7380 = w4762 & ~w4582;
assign w7381 = w101 & ~w4530;
assign w7382 = (~w3057 & w1332) | (~w3057 & w2444) | (w1332 & w2444);
assign w7383 = w5686 & ~w7218;
assign w7384 = a140 & b140;
assign w7385 = (~w1327 & w7420) | (~w1327 & w3313) | (w7420 & w3313);
assign w7386 = ~w4337 & w4555;
assign w7387 = (~w6945 & w6667) | (~w6945 & w3930) | (w6667 & w3930);
assign w7388 = (~w5655 & w4928) | (~w5655 & w2480) | (w4928 & w2480);
assign w7389 = (~w3384 & ~w1675) | (~w3384 & ~w5368) | (~w1675 & ~w5368);
assign w7390 = a18 & b18;
assign w7391 = a36 & b36;
assign w7392 = ~w5665 & ~w5972;
assign w7393 = ~w4180 & w887;
assign w7394 = ~w6025 & ~w3328;
assign w7395 = w6845 & w4989;
assign w7396 = ~w3207 & ~w4497;
assign w7397 = w4249 & ~w321;
assign w7398 = (~w6279 & ~w3349) | (~w6279 & w2059) | (~w3349 & w2059);
assign w7399 = ~a112 & ~b112;
assign w7400 = (w6499 & w2810) | (w6499 & w2097) | (w2810 & w2097);
assign w7401 = (~w3078 & w2889) | (~w3078 & w5885) | (w2889 & w5885);
assign w7402 = w5403 & w4824;
assign w7403 = w1735 & w2582;
assign w7404 = ~w1614 & w2663;
assign w7405 = ~w2880 & w5296;
assign w7406 = ~w7279 & w65;
assign w7407 = w1485 & ~w2954;
assign w7408 = ~w7005 & ~w4933;
assign w7409 = w5056 & w2246;
assign w7410 = (~w4182 & w3448) | (~w4182 & w3599) | (w3448 & w3599);
assign w7411 = w3336 & w2623;
assign w7412 = ~w4713 & ~w1463;
assign w7413 = (w2068 & ~w3880) | (w2068 & w5449) | (~w3880 & w5449);
assign w7414 = ~w4193 & ~w4004;
assign w7415 = (w6675 & w969) | (w6675 & w7615) | (w969 & w7615);
assign w7416 = (~w3331 & w3736) | (~w3331 & w2314) | (w3736 & w2314);
assign w7417 = ~w4238 & ~w51;
assign w7418 = (w6353 & w5050) | (w6353 & w3020) | (w5050 & w3020);
assign w7419 = (w1724 & w419) | (w1724 & w6100) | (w419 & w6100);
assign w7420 = ~w2954 & ~w454;
assign w7421 = (~w4010 & w2172) | (~w4010 & w5039) | (w2172 & w5039);
assign w7422 = ~w7063 & w431;
assign w7423 = (w5078 & w5338) | (w5078 & w5215) | (w5338 & w5215);
assign w7424 = a115 & b115;
assign w7425 = ~w4101 & ~w7308;
assign w7426 = ~w4397 & ~w5274;
assign w7427 = w7292 & ~w5960;
assign w7428 = (~w777 & w5086) | (~w777 & w2319) | (w5086 & w2319);
assign w7429 = w4350 & ~w972;
assign w7430 = (w3570 & ~w6845) | (w3570 & w1330) | (~w6845 & w1330);
assign w7431 = (w5921 & w5290) | (w5921 & ~w4867) | (w5290 & ~w4867);
assign w7432 = ~w1409 & w5286;
assign w7433 = (~w5257 & w1120) | (~w5257 & w3795) | (w1120 & w3795);
assign w7434 = ~w3561 & w5642;
assign w7435 = (~w9 & w2245) | (~w9 & w6504) | (w2245 & w6504);
assign w7436 = (w5655 & w3611) | (w5655 & w5854) | (w3611 & w5854);
assign w7437 = (~w3736 & w6023) | (~w3736 & w3971) | (w6023 & w3971);
assign w7438 = ~w841 & ~w1661;
assign w7439 = ~w3101 & w6170;
assign w7440 = (w2301 & w7006) | (w2301 & w2013) | (w7006 & w2013);
assign w7441 = (w6190 & w4650) | (w6190 & ~w3983) | (w4650 & ~w3983);
assign w7442 = w3132 & w1311;
assign w7443 = (w264 & w6470) | (w264 & w4318) | (w6470 & w4318);
assign w7444 = ~w5922 & ~w1791;
assign w7445 = w3836 & ~w7035;
assign w7446 = ~w2566 & ~w7530;
assign w7447 = ~w6683 & ~w6161;
assign w7448 = (~w6279 & w5194) | (~w6279 & w5715) | (w5194 & w5715);
assign w7449 = w1833 & ~w5961;
assign w7450 = (w1193 & w236) | (w1193 & w4624) | (w236 & w4624);
assign w7451 = ~w3248 & w2104;
assign w7452 = ~a24 & ~b24;
assign w7453 = (w1728 & w6046) | (w1728 & w4588) | (w6046 & w4588);
assign w7454 = (~w4891 & ~w1565) | (~w4891 & w7156) | (~w1565 & w7156);
assign w7455 = ~w337 & ~w3721;
assign w7456 = w4179 & ~w5772;
assign w7457 = ~w3355 & ~w3809;
assign w7458 = w5246 & ~w317;
assign w7459 = (w2182 & w282) | (w2182 & w2602) | (w282 & w2602);
assign w7460 = w7203 & w283;
assign w7461 = w3183 & ~w3974;
assign w7462 = w4132 & w5958;
assign w7463 = w4072 & ~w1879;
assign w7464 = (w4777 & w4905) | (w4777 & w6214) | (w4905 & w6214);
assign w7465 = (w4787 & w4273) | (w4787 & ~w5368) | (w4273 & ~w5368);
assign w7466 = ~w4490 & ~w2851;
assign w7467 = (w4905 & w6410) | (w4905 & w3727) | (w6410 & w3727);
assign w7468 = (w5554 & w1229) | (w5554 & w4803) | (w1229 & w4803);
assign w7469 = (~w1611 & w513) | (~w1611 & w1726) | (w513 & w1726);
assign w7470 = (w6082 & w6914) | (w6082 & w6238) | (w6914 & w6238);
assign w7471 = ~w2718 & ~w5862;
assign w7472 = ~w1998 & w1489;
assign w7473 = (~w4089 & w4309) | (~w4089 & w5795) | (w4309 & w5795);
assign w7474 = ~w1946 & ~w2456;
assign w7475 = (w3318 & w4062) | (w3318 & w7586) | (w4062 & w7586);
assign w7476 = w3864 & ~w5376;
assign w7477 = w3102 & ~w7401;
assign w7478 = w5011 & w7028;
assign w7479 = (w4652 & w6005) | (w4652 & ~w4199) | (w6005 & ~w4199);
assign w7480 = ~w3480 & ~w30;
assign w7481 = (~w5402 & w3324) | (~w5402 & w1) | (w3324 & w1);
assign w7482 = ~w4653 & ~w715;
assign w7483 = ~w5404 & ~w4473;
assign w7484 = ~w3298 & ~w161;
assign w7485 = (w719 & w5595) | (w719 & w2456) | (w5595 & w2456);
assign w7486 = ~a240 & ~b240;
assign w7487 = w1162 & w2023;
assign w7488 = (w5484 & w826) | (w5484 & w2518) | (w826 & w2518);
assign w7489 = (w5344 & w4068) | (w5344 & w1499) | (w4068 & w1499);
assign w7490 = (~w624 & w7020) | (~w624 & w1614) | (w7020 & w1614);
assign w7491 = ~w4499 & ~w4306;
assign w7492 = w2982 & ~w7571;
assign w7493 = ~a133 & ~b133;
assign w7494 = (w5655 & w2187) | (w5655 & w6055) | (w2187 & w6055);
assign w7495 = (w6100 & w5652) | (w6100 & w3790) | (w5652 & w3790);
assign w7496 = (~w3503 & ~w6270) | (~w3503 & w457) | (~w6270 & w457);
assign w7497 = ~w863 & ~w418;
assign w7498 = ~w6861 & w1658;
assign w7499 = (w6572 & w4621) | (w6572 & ~w4021) | (w4621 & ~w4021);
assign w7500 = ~w161 & ~w6776;
assign w7501 = (w4733 & w1749) | (w4733 & w6858) | (w1749 & w6858);
assign w7502 = w2982 & w6100;
assign w7503 = (w7414 & w5359) | (w7414 & ~w6100) | (w5359 & ~w6100);
assign w7504 = ~w5952 & ~w4631;
assign w7505 = (w2021 & w6604) | (w2021 & w3861) | (w6604 & w3861);
assign w7506 = ~w4674 & ~w4123;
assign w7507 = ~a219 & ~b219;
assign w7508 = (w6274 & w2961) | (w6274 & w1881) | (w2961 & w1881);
assign w7509 = ~w6439 & ~w2096;
assign w7510 = ~w2945 & ~w6319;
assign w7511 = (w505 & ~w1153) | (w505 & ~w6566) | (~w1153 & ~w6566);
assign w7512 = (w6685 & ~w7610) | (w6685 & w2447) | (~w7610 & w2447);
assign w7513 = w135 & ~w6871;
assign w7514 = (w6614 & w4619) | (w6614 & w2118) | (w4619 & w2118);
assign w7515 = (~w1847 & w5490) | (~w1847 & w5314) | (w5490 & w5314);
assign w7516 = w2830 & w6134;
assign w7517 = (w388 & w1634) | (w388 & w2126) | (w1634 & w2126);
assign w7518 = w6512 & ~w5328;
assign w7519 = ~w7271 & ~w908;
assign w7520 = (w1266 & ~w1006) | (w1266 & w5185) | (~w1006 & w5185);
assign w7521 = (~w5486 & ~w2041) | (~w5486 & w7232) | (~w2041 & w7232);
assign w7522 = a103 & b103;
assign w7523 = (w893 & w5178) | (w893 & w4278) | (w5178 & w4278);
assign w7524 = w4036 & w4798;
assign w7525 = a128 & b128;
assign w7526 = ~w7346 & ~w4168;
assign w7527 = ~a68 & ~b68;
assign w7528 = ~w2041 & w5421;
assign w7529 = ~w6942 & w7640;
assign w7530 = ~a16 & ~b16;
assign w7531 = (w7310 & w4434) | (w7310 & w2456) | (w4434 & w2456);
assign w7532 = (w737 & w5765) | (w737 & ~w6254) | (w5765 & ~w6254);
assign w7533 = (~w5178 & w4818) | (~w5178 & w3517) | (w4818 & w3517);
assign w7534 = w2024 & w6608;
assign w7535 = ~w3896 & w4505;
assign w7536 = a254 & b254;
assign w7537 = w2255 & ~w6658;
assign w7538 = ~w4677 & ~w7265;
assign w7539 = ~w3887 & ~w2072;
assign w7540 = (w3318 & w1481) | (w3318 & w6793) | (w1481 & w6793);
assign w7541 = w6599 & w1910;
assign w7542 = (~w5419 & w2734) | (~w5419 & w5102) | (w2734 & w5102);
assign w7543 = ~w1936 & w2531;
assign w7544 = (w5257 & w6300) | (w5257 & w4013) | (w6300 & w4013);
assign w7545 = ~w3580 & w757;
assign w7546 = ~a18 & ~b18;
assign w7547 = (~w3847 & ~w4286) | (~w3847 & w3374) | (~w4286 & w3374);
assign w7548 = (~w6738 & w5614) | (~w6738 & w6498) | (w5614 & w6498);
assign w7549 = w4504 & w738;
assign w7550 = ~w3961 & ~w150;
assign w7551 = (~w5385 & w1815) | (~w5385 & w7485) | (w1815 & w7485);
assign w7552 = ~w5820 & ~w5926;
assign w7553 = ~w6703 & ~w6980;
assign w7554 = w2564 & w6408;
assign w7555 = ~w3909 & ~w4198;
assign w7556 = w4503 & w2315;
assign w7557 = (~w1682 & w7307) | (~w1682 & w5674) | (w7307 & w5674);
assign w7558 = ~w5066 | w2666;
assign w7559 = w3231 & ~w491;
assign w7560 = (~w6082 & w938) | (~w6082 & w5508) | (w938 & w5508);
assign w7561 = (~w3461 & w609) | (~w3461 & w5621) | (w609 & w5621);
assign w7562 = (~w1722 & w4287) | (~w1722 & w1501) | (w4287 & w1501);
assign w7563 = ~w1216 & ~w6884;
assign w7564 = ~a189 & ~b189;
assign w7565 = ~w5183 & w2122;
assign w7566 = ~w4891 & ~w5759;
assign w7567 = ~w3616 & ~w6608;
assign w7568 = (~w5478 & w3957) | (~w5478 & ~w3482) | (w3957 & ~w3482);
assign w7569 = ~w5641 & w2996;
assign w7570 = w4906 & ~w3212;
assign w7571 = ~w6082 & w4228;
assign w7572 = a184 & b184;
assign w7573 = (w6372 & w1844) | (w6372 & ~w1881) | (w1844 & ~w1881);
assign w7574 = ~w3482 & ~w226;
assign w7575 = ~w273 & w1234;
assign w7576 = ~w2182 & w1271;
assign w7577 = ~w1848 & ~w973;
assign w7578 = w3105 & ~w3206;
assign w7579 = ~w6784 & ~w3274;
assign w7580 = w6875 & w4702;
assign w7581 = ~a116 & ~b116;
assign w7582 = (w7626 & w5636) | (w7626 & w3841) | (w5636 & w3841);
assign w7583 = ~w2108 & ~w5807;
assign w7584 = ~w3009 & w5757;
assign w7585 = w7439 & w6840;
assign w7586 = (w136 & w842) | (w136 & ~w5291) | (w842 & ~w5291);
assign w7587 = ~w5944 & w7545;
assign w7588 = ~w4706 & w2945;
assign w7589 = (w6424 & w5092) | (w6424 & w3638) | (w5092 & w3638);
assign w7590 = (~w5178 & w1061) | (~w5178 & w2165) | (w1061 & w2165);
assign w7591 = w4611 & ~w3210;
assign w7592 = ~w4060 & ~w1002;
assign w7593 = (w6151 & w748) | (w6151 & w158) | (w748 & w158);
assign w7594 = w1851 & w134;
assign w7595 = (~w5901 & w4420) | (~w5901 & w3633) | (w4420 & w3633);
assign w7596 = w2099 & ~w5366;
assign w7597 = (w2847 & w2574) | (w2847 & w987) | (w2574 & w987);
assign w7598 = w2458 & ~w5398;
assign w7599 = ~w3587 & w3331;
assign w7600 = (w3427 & w2172) | (w3427 & w3787) | (w2172 & w3787);
assign w7601 = w6366 & ~w4147;
assign w7602 = (w7197 & w6937) | (w7197 & w7516) | (w6937 & w7516);
assign w7603 = ~w4167 & ~w4132;
assign w7604 = ~w6979 & ~w5923;
assign w7605 = w3415 & w4710;
assign w7606 = w1577 & ~w187;
assign w7607 = ~w6599 & w401;
assign w7608 = ~w7147 & w7535;
assign w7609 = (w5655 & w1242) | (w5655 & w2144) | (w1242 & w2144);
assign w7610 = ~w1660 & w5858;
assign w7611 = ~w3211 & ~w3541;
assign w7612 = (~w7510 & w4923) | (~w7510 & w343) | (w4923 & w343);
assign w7613 = ~w6115 & ~w1359;
assign w7614 = ~a55 & ~b55;
assign w7615 = w7231 & ~w1086;
assign w7616 = w5510 & ~w5056;
assign w7617 = (w6600 & w1473) | (w6600 & ~w173) | (w1473 & ~w173);
assign w7618 = (~w6100 & w1509) | (~w6100 & w7171) | (w1509 & w7171);
assign w7619 = (~w2985 & w2239) | (~w2985 & w4332) | (w2239 & w4332);
assign w7620 = (w5178 & w1928) | (w5178 & w4834) | (w1928 & w4834);
assign w7621 = (w5178 & w4804) | (w5178 & w2423) | (w4804 & w2423);
assign w7622 = a86 & b86;
assign w7623 = (w1097 & w1872) | (w1097 & w6566) | (w1872 & w6566);
assign w7624 = w807 & w3197;
assign w7625 = ~w3551 & ~w1967;
assign w7626 = ~w438 & ~w2814;
assign w7627 = ~w6189 & ~w3405;
assign w7628 = (w6675 & w2815) | (w6675 & w7369) | (w2815 & w7369);
assign w7629 = ~w4350 & w625;
assign w7630 = ~w4067 & w6895;
assign w7631 = w4115 & w5269;
assign w7632 = a95 & b95;
assign w7633 = w4146 & ~w3712;
assign w7634 = a159 & b159;
assign w7635 = (w2627 & w3031) | (w2627 & w3250) | (w3031 & w3250);
assign w7636 = (w922 & w5067) | (w922 & w5325) | (w5067 & w5325);
assign w7637 = (w3119 & w7580) | (w3119 & w5207) | (w7580 & w5207);
assign w7638 = (~w4505 & w7147) | (~w4505 & w616) | (w7147 & w616);
assign w7639 = (~w3952 & w2543) | (~w3952 & w2761) | (w2543 & w2761);
assign w7640 = ~w2283 & w7097;
assign w7641 = ~a110 & ~b110;
assign w7642 = (w5655 & w6659) | (w5655 & w1166) | (w6659 & w1166);
assign w7643 = (w3472 & w5403) | (w3472 & w1254) | (w5403 & w1254);
assign w7644 = ~w7213 & ~w3075;
assign w7645 = w174 & w6045;
assign w7646 = w3158 & w76;
assign w7647 = ~w6690 & ~w3896;
assign w7648 = a207 & b207;
assign w7649 = (~w6524 & w663) | (~w6524 & ~w1743) | (w663 & ~w1743);
assign one = 1;
assign s0 = ~w1729;// level 4
assign s1 = w904;// level 5
assign s2 = w6029;// level 5
assign s3 = ~w2025;// level 6
assign s4 = w2908;// level 6
assign s5 = ~w3120;// level 6
assign s6 = w5256;// level 6
assign s7 = ~w7613;// level 7
assign s8 = ~w4887;// level 7
assign s9 = ~w3180;// level 7
assign s10 = ~w6133;// level 7
assign s11 = ~w7208;// level 8
assign s12 = ~w3390;// level 8
assign s13 = ~w581;// level 8
assign s14 = ~w3675;// level 8
assign s15 = ~w4414;// level 8
assign s16 = w890;// level 8
assign s17 = ~w2501;// level 8
assign s18 = ~w6700;// level 8
assign s19 = ~w3386;// level 9
assign s20 = ~w5653;// level 9
assign s21 = ~w3457;// level 9
assign s22 = ~w4931;// level 9
assign s23 = ~w2148;// level 9
assign s24 = ~w5293;// level 9
assign s25 = ~w1113;// level 9
assign s26 = ~w3670;// level 9
assign s27 = ~w66;// level 9
assign s28 = ~w6178;// level 9
assign s29 = w1466;// level 9
assign s30 = ~w3960;// level 9
assign s31 = ~w3627;// level 9
assign s32 = ~w6756;// level 9
assign s33 = ~w4070;// level 10
assign s34 = w2730;// level 10
assign s35 = ~w5736;// level 10
assign s36 = ~w643;// level 10
assign s37 = ~w3877;// level 10
assign s38 = w3495;// level 10
assign s39 = ~w324;// level 10
assign s40 = ~w3404;// level 10
assign s41 = ~w3837;// level 10
assign s42 = w7139;// level 11
assign s43 = ~w1517;// level 10
assign s44 = ~w5393;// level 11
assign s45 = ~w5444;// level 10
assign s46 = ~w6940;// level 10
assign s47 = ~w6946;// level 11
assign s48 = ~w7426;// level 10
assign s49 = ~w3773;// level 10
assign s50 = ~w2652;// level 10
assign s51 = w6124;// level 10
assign s52 = ~w349;// level 11
assign s53 = ~w5465;// level 11
assign s54 = ~w674;// level 10
assign s55 = w4063;// level 10
assign s56 = ~w3464;// level 11
assign s57 = ~w4769;// level 11
assign s58 = w4593;// level 11
assign s59 = w92;// level 11
assign s60 = w4111;// level 11
assign s61 = ~w877;// level 11
assign s62 = ~w7075;// level 11
assign s63 = ~w223;// level 11
assign s64 = ~w1194;// level 11
assign s65 = ~w3659;// level 11
assign s66 = ~w2512;// level 11
assign s67 = ~w5647;// level 11
assign s68 = w2916;// level 11
assign s69 = ~w7455;// level 11
assign s70 = ~w4670;// level 11
assign s71 = ~w4445;// level 12
assign s72 = ~w4839;// level 11
assign s73 = w5472;// level 11
assign s74 = ~w6567;// level 12
assign s75 = w4789;// level 11
assign s76 = ~w7149;// level 11
assign s77 = w4563;// level 11
assign s78 = w5558;// level 12
assign s79 = ~w450;// level 12
assign s80 = ~w653;// level 12
assign s81 = w7104;// level 12
assign s82 = ~w943;// level 12
assign s83 = ~w1253;// level 12
assign s84 = ~w5730;// level 12
assign s85 = ~w5733;// level 12
assign s86 = ~w2469;// level 12
assign s87 = ~w7466;// level 12
assign s88 = ~w1382;// level 12
assign s89 = ~w323;// level 12
assign s90 = ~w1599;// level 12
assign s91 = ~w6069;// level 12
assign s92 = w5719;// level 12
assign s93 = ~w5101;// level 12
assign s94 = ~w2779;// level 12
assign s95 = ~w1645;// level 12
assign s96 = w359;// level 12
assign s97 = ~w3853;// level 12
assign s98 = ~w5737;// level 12
assign s99 = ~w2063;// level 12
assign s100 = ~w6820;// level 12
assign s101 = w152;// level 12
assign s102 = ~w2195;// level 12
assign s103 = ~w4515;// level 12
assign s104 = w5110;// level 12
assign s105 = w4294;// level 12
assign s106 = ~w2546;// level 12
assign s107 = ~w204;// level 12
assign s108 = ~w4644;// level 12
assign s109 = ~w7457;// level 12
assign s110 = w2508;// level 12
assign s111 = ~w7247;// level 12
assign s112 = ~w1003;// level 13
assign s113 = w785;// level 13
assign s114 = w1436;// level 13
assign s115 = ~w6171;// level 13
assign s116 = ~w2747;// level 13
assign s117 = ~w3711;// level 13
assign s118 = ~w3475;// level 13
assign s119 = w3822;// level 14
assign s120 = ~w117;// level 13
assign s121 = ~w3578;// level 13
assign s122 = ~w3241;// level 14
assign s123 = w776;// level 13
assign s124 = ~w5206;// level 13
assign s125 = ~w6241;// level 13
assign s126 = w6358;// level 13
assign s127 = ~w4630;// level 13
assign s128 = w836;// level 13
assign s129 = ~w5889;// level 13
assign s130 = ~w5074;// level 14
assign s131 = w4936;// level 14
assign s132 = w2754;// level 14
assign s133 = ~w801;// level 13
assign s134 = ~w6154;// level 14
assign s135 = w4654;// level 13
assign s136 = ~w7611;// level 13
assign s137 = w2556;// level 14
assign s138 = ~w4883;// level 13
assign s139 = ~w6859;// level 13
assign s140 = ~w4678;// level 13
assign s141 = w4364;// level 13
assign s142 = ~w6899;// level 13
assign s143 = ~w2587;// level 13
assign s144 = ~w2685;// level 13
assign s145 = ~w3395;// level 14
assign s146 = w4417;// level 14
assign s147 = ~w4482;// level 13
assign s148 = ~w6128;// level 14
assign s149 = w1385;// level 14
assign s150 = w7504;// level 13
assign s151 = ~w6538;// level 13
assign s152 = w514;// level 13
assign s153 = w5010;// level 13
assign s154 = ~w2642;// level 14
assign s155 = w2530;// level 13
assign s156 = ~w1049;// level 13
assign s157 = ~w4134;// level 13
assign s158 = w4500;// level 13
assign s159 = w3439;// level 14
assign s160 = ~w2487;// level 13
assign s161 = ~w7069;// level 13
assign s162 = w7579;// level 13
assign s163 = ~w2696;// level 14
assign s164 = ~w1912;// level 14
assign s165 = ~w4449;// level 13
assign s166 = ~w1188;// level 13
assign s167 = ~w5169;// level 13
assign s168 = w1244;// level 13
assign s169 = ~w6003;// level 13
assign s170 = ~w6519;// level 14
assign s171 = ~w5731;// level 14
assign s172 = ~w3714;// level 14
assign s173 = w5968;// level 14
assign s174 = ~w6728;// level 14
assign s175 = ~w5775;// level 14
assign s176 = ~w4352;// level 14
assign s177 = w4947;// level 14
assign s178 = ~w4974;// level 14
assign s179 = ~w3463;// level 14
assign s180 = w4903;// level 14
assign s181 = w6092;// level 14
assign s182 = w7497;// level 14
assign s183 = ~w2204;// level 14
assign s184 = w6795;// level 14
assign s185 = ~w2034;// level 14
assign s186 = ~w111;// level 14
assign s187 = ~w5213;// level 14
assign s188 = ~w3850;// level 14
assign s189 = ~w4462;// level 14
assign s190 = ~w2783;// level 14
assign s191 = ~w6765;// level 14
assign s192 = w7482;// level 14
assign s193 = ~w7550;// level 14
assign s194 = w897;// level 14
assign s195 = w7251;// level 14
assign s196 = ~w1705;// level 14
assign s197 = w3275;// level 14
assign s198 = w2039;// level 14
assign s199 = ~w5049;// level 14
assign s200 = ~w201;// level 14
assign s201 = ~w4877;// level 14
assign s202 = w6308;// level 16
assign s203 = w3186;// level 14
assign s204 = w2381;// level 14
assign s205 = w2151;// level 15
assign s206 = w197;// level 14
assign s207 = w5214;// level 14
assign s208 = ~w2457;// level 14
assign s209 = ~w5989;// level 14
assign s210 = w5940;// level 14
assign s211 = w1995;// level 16
assign s212 = w489;// level 14
assign s213 = ~w6483;// level 14
assign s214 = ~w5334;// level 14
assign s215 = ~w6349;// level 14
assign s216 = w4374;// level 14
assign s217 = ~w5971;// level 14
assign s218 = ~w2758;// level 14
assign s219 = w2213;// level 14
assign s220 = ~w4992;// level 14
assign s221 = ~w4978;// level 14
assign s222 = ~w1460;// level 14
assign s223 = ~w4498;// level 14
assign s224 = w595;// level 14
assign s225 = w6320;// level 14
assign s226 = ~w2571;// level 14
assign s227 = w1268;// level 14
assign s228 = w3400;// level 14
assign s229 = ~w3825;// level 14
assign s230 = ~w7270;// level 14
assign s231 = ~w6380;// level 14
assign s232 = ~w2174;// level 14
assign s233 = ~w5117;// level 14
assign s234 = w191;// level 14
assign s235 = ~w3227;// level 14
assign s236 = ~w6720;// level 14
assign s237 = ~w533;// level 14
assign s238 = ~w7211;// level 14
assign s239 = ~w5764;// level 14
assign s240 = w3109;// level 16
assign s241 = ~w7059;// level 14
assign s242 = ~w6952;// level 14
assign s243 = w2817;// level 14
assign s244 = ~w2951;// level 14
assign s245 = ~w5949;// level 14
assign s246 = w2812;// level 15
assign s247 = ~w6973;// level 14
assign s248 = ~w6245;// level 14
assign s249 = w6393;// level 14
assign s250 = ~w3900;// level 14
assign s251 = ~w5062;// level 14
assign s252 = w2363;// level 14
assign s253 = w5615;// level 15
assign s254 = ~w1159;// level 14
assign s255 = ~w772;// level 14
assign s256 = w6006;// level 15
endmodule
