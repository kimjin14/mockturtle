module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 ;
  wire n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , n3931 , n3932 , n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , n3940 , n3941 , n3942 , n3943 , n3944 , n3945 , n3946 , n3947 , n3948 , n3949 , n3950 , n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , n3970 , n3971 , n3972 , n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , n3980 , n3981 , n3982 , n3983 , n3984 , n3985 , n3986 , n3987 , n3988 , n3989 , n3990 , n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , n4000 , n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , n4009 , n4010 , n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , n4019 , n4020 , n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , n4029 , n4030 , n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , n4039 , n4040 , n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4049 , n4050 , n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , n4059 , n4060 , n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , n4070 , n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , n4079 , n4080 , n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , n4089 , n4090 , n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , n4097 , n4098 , n4099 , n4100 , n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , n4109 , n4110 , n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , n4119 , n4120 , n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , n4129 , n4130 , n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , n4139 , n4140 , n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , n4150 , n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , n4159 , n4160 , n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , n4169 , n4170 , n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , n4179 , n4180 , n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , n4189 , n4190 , n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , n4197 , n4198 , n4199 , n4200 , n4201 , n4202 , n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , n4209 , n4210 , n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , n4217 , n4218 , n4219 , n4220 , n4221 , n4222 , n4223 , n4224 , n4225 , n4226 , n4227 , n4228 , n4229 , n4230 , n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , n4237 , n4238 , n4239 , n4240 , n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , n4247 , n4248 , n4249 , n4250 , n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , n4259 , n4260 , n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , n4269 , n4270 , n4271 , n4272 , n4273 , n4274 , n4275 , n4276 , n4277 , n4278 , n4279 , n4280 , n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , n4289 , n4290 , n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , n4299 , n4300 , n4301 , n4302 , n4303 , n4304 , n4305 , n4306 , n4307 , n4308 , n4309 , n4310 , n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , n4319 , n4320 , n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , n4329 , n4330 , n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , n4340 , n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , n4349 , n4350 , n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , n4360 , n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , n4370 , n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , n4380 , n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , n4390 , n4391 , n4392 , n4393 , n4394 , n4395 , n4396 , n4397 , n4398 , n4399 , n4400 , n4401 , n4402 , n4403 , n4404 , n4405 , n4406 , n4407 , n4408 , n4409 , n4410 , n4411 , n4412 , n4413 , n4414 , n4415 , n4416 , n4417 , n4418 , n4419 , n4420 , n4421 , n4422 , n4423 , n4424 , n4425 , n4426 , n4427 , n4428 , n4429 , n4430 , n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , n4437 , n4438 , n4439 , n4440 , n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , n4449 , n4450 , n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , n4459 , n4460 , n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , n4469 , n4470 , n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , n4479 , n4480 , n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , n4487 , n4488 , n4489 , n4490 , n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , n4497 , n4498 , n4499 , n4500 , n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , n4509 , n4510 , n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , n4519 , n4520 , n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , n4529 , n4530 , n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , n4537 , n4538 , n4539 , n4540 , n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , n4547 , n4548 , n4549 , n4550 , n4551 , n4552 , n4553 , n4554 , n4555 , n4556 , n4557 , n4558 , n4559 , n4560 , n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , n4567 , n4568 , n4569 , n4570 , n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , n4579 , n4580 , n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , n4589 , n4590 , n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , n4597 , n4598 , n4599 , n4600 , n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , n4607 , n4608 , n4609 , n4610 , n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , n4617 , n4618 , n4619 , n4620 , n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , n4627 , n4628 , n4629 , n4630 , n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , n4637 , n4638 , n4639 , n4640 , n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , n4647 , n4648 , n4649 , n4650 , n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , n4657 , n4658 , n4659 , n4660 , n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , n4669 , n4670 , n4671 , n4672 , n4673 , n4674 , n4675 , n4676 , n4677 , n4678 , n4679 , n4680 , n4681 , n4682 , n4683 , n4684 , n4685 , n4686 , n4687 , n4688 , n4689 , n4690 , n4691 , n4692 , n4693 , n4694 , n4695 , n4696 , n4697 , n4698 , n4699 , n4700 , n4701 , n4702 , n4703 , n4704 , n4705 , n4706 , n4707 , n4708 , n4709 , n4710 , n4711 , n4712 , n4713 , n4714 , n4715 , n4716 , n4717 , n4718 , n4719 , n4720 , n4721 , n4722 , n4723 , n4724 , n4725 , n4726 , n4727 , n4728 , n4729 , n4730 , n4731 , n4732 , n4733 , n4734 , n4735 , n4736 , n4737 , n4738 , n4739 , n4740 , n4741 , n4742 , n4743 , n4744 , n4745 , n4746 , n4747 , n4748 , n4749 , n4750 , n4751 , n4752 , n4753 , n4754 , n4755 , n4756 , n4757 , n4758 , n4759 , n4760 , n4761 , n4762 , n4763 , n4764 , n4765 , n4766 , n4767 , n4768 , n4769 , n4770 , n4771 , n4772 , n4773 , n4774 , n4775 , n4776 , n4777 , n4778 , n4779 , n4780 , n4781 , n4782 , n4783 , n4784 , n4785 , n4786 , n4787 , n4788 , n4789 , n4790 , n4791 , n4792 , n4793 , n4794 , n4795 , n4796 , n4797 , n4798 , n4799 , n4800 , n4801 , n4802 , n4803 , n4804 , n4805 , n4806 , n4807 , n4808 , n4809 , n4810 , n4811 , n4812 , n4813 , n4814 , n4815 , n4816 , n4817 , n4818 , n4819 , n4820 , n4821 , n4822 , n4823 , n4824 , n4825 , n4826 , n4827 , n4828 , n4829 , n4830 , n4831 , n4832 , n4833 , n4834 , n4835 , n4836 , n4837 , n4838 , n4839 , n4840 , n4841 , n4842 , n4843 , n4844 , n4845 , n4846 , n4847 , n4848 , n4849 , n4850 , n4851 , n4852 , n4853 , n4854 , n4855 , n4856 , n4857 , n4858 , n4859 , n4860 , n4861 , n4862 , n4863 , n4864 , n4865 , n4866 , n4867 , n4868 , n4869 , n4870 , n4871 , n4872 , n4873 , n4874 , n4875 , n4876 , n4877 , n4878 , n4879 , n4880 , n4881 , n4882 , n4883 , n4884 , n4885 , n4886 , n4887 , n4888 , n4889 , n4890 , n4891 , n4892 , n4893 , n4894 , n4895 , n4896 , n4897 , n4898 , n4899 , n4900 , n4901 , n4902 , n4903 , n4904 , n4905 , n4906 , n4907 , n4908 , n4909 , n4910 , n4911 , n4912 , n4913 , n4914 , n4915 , n4916 , n4917 , n4918 , n4919 , n4920 , n4921 , n4922 , n4923 , n4924 , n4925 , n4926 , n4927 , n4928 , n4929 , n4930 , n4931 , n4932 , n4933 , n4934 , n4935 , n4936 , n4937 , n4938 , n4939 , n4940 , n4941 , n4942 , n4943 , n4944 , n4945 , n4946 , n4947 , n4948 , n4949 , n4950 , n4951 , n4952 , n4953 , n4954 , n4955 , n4956 , n4957 , n4958 , n4959 , n4960 , n4961 , n4962 , n4963 , n4964 , n4965 , n4966 , n4967 , n4968 , n4969 , n4970 , n4971 , n4972 , n4973 , n4974 , n4975 , n4976 , n4977 , n4978 , n4979 , n4980 , n4981 , n4982 , n4983 , n4984 , n4985 , n4986 , n4987 , n4988 , n4989 , n4990 , n4991 , n4992 , n4993 , n4994 , n4995 , n4996 , n4997 , n4998 , n4999 , n5000 , n5001 , n5002 , n5003 , n5004 , n5005 , n5006 , n5007 , n5008 , n5009 , n5010 , n5011 , n5012 , n5013 , n5014 , n5015 , n5016 , n5017 , n5018 , n5019 , n5020 , n5021 , n5022 , n5023 , n5024 , n5025 , n5026 , n5027 , n5028 , n5029 , n5030 , n5031 , n5032 , n5033 , n5034 , n5035 , n5036 , n5037 , n5038 , n5039 , n5040 , n5041 , n5042 , n5043 , n5044 , n5045 , n5046 , n5047 , n5048 , n5049 , n5050 , n5051 , n5052 , n5053 , n5054 , n5055 , n5056 , n5057 , n5058 , n5059 , n5060 , n5061 , n5062 , n5063 , n5064 , n5065 , n5066 , n5067 , n5068 , n5069 , n5070 , n5071 , n5072 , n5073 , n5074 , n5075 , n5076 , n5077 , n5078 , n5079 , n5080 , n5081 , n5082 , n5083 , n5084 , n5085 , n5086 , n5087 , n5088 , n5089 , n5090 , n5091 , n5092 , n5093 , n5094 , n5095 , n5096 , n5097 , n5098 , n5099 , n5100 , n5101 , n5102 , n5103 , n5104 , n5105 , n5106 , n5107 , n5108 , n5109 , n5110 , n5111 , n5112 , n5113 , n5114 , n5115 , n5116 , n5117 , n5118 , n5119 , n5120 , n5121 , n5122 , n5123 , n5124 , n5125 , n5126 , n5127 , n5128 , n5129 , n5130 , n5131 , n5132 , n5133 , n5134 , n5135 , n5136 , n5137 , n5138 , n5139 , n5140 , n5141 , n5142 , n5143 , n5144 , n5145 , n5146 , n5147 , n5148 , n5149 , n5150 , n5151 , n5152 , n5153 , n5154 , n5155 , n5156 , n5157 , n5158 , n5159 , n5160 , n5161 , n5162 , n5163 , n5164 , n5165 , n5166 , n5167 , n5168 , n5169 , n5170 , n5171 , n5172 , n5173 , n5174 , n5175 , n5176 , n5177 , n5178 , n5179 , n5180 , n5181 , n5182 , n5183 , n5184 , n5185 , n5186 , n5187 , n5188 , n5189 , n5190 , n5191 , n5192 , n5193 , n5194 , n5195 , n5196 , n5197 , n5198 , n5199 , n5200 , n5201 , n5202 , n5203 , n5204 , n5205 , n5206 , n5207 , n5208 , n5209 , n5210 , n5211 , n5212 , n5213 , n5214 , n5215 , n5216 , n5217 , n5218 , n5219 , n5220 , n5221 , n5222 , n5223 , n5224 , n5225 , n5226 , n5227 , n5228 , n5229 , n5230 , n5231 , n5232 , n5233 , n5234 , n5235 , n5236 , n5237 , n5238 , n5239 , n5240 , n5241 , n5242 , n5243 , n5244 , n5245 , n5246 , n5247 , n5248 , n5249 , n5250 , n5251 , n5252 , n5253 , n5254 , n5255 , n5256 , n5257 , n5258 , n5259 , n5260 , n5261 , n5262 , n5263 , n5264 , n5265 , n5266 , n5267 , n5268 , n5269 , n5270 , n5271 , n5272 , n5273 , n5274 , n5275 , n5276 , n5277 , n5278 , n5279 , n5280 , n5281 , n5282 , n5283 , n5284 , n5285 , n5286 , n5287 , n5288 , n5289 , n5290 , n5291 , n5292 , n5293 , n5294 , n5295 , n5296 , n5297 , n5298 , n5299 , n5300 , n5301 , n5302 , n5303 , n5304 , n5305 , n5306 , n5307 , n5308 , n5309 , n5310 , n5311 , n5312 , n5313 , n5314 , n5315 , n5316 , n5317 , n5318 , n5319 , n5320 , n5321 , n5322 , n5323 , n5324 , n5325 , n5326 , n5327 , n5328 , n5329 , n5330 , n5331 , n5332 , n5333 , n5334 , n5335 , n5336 , n5337 , n5338 , n5339 , n5340 , n5341 , n5342 , n5343 , n5344 , n5345 , n5346 , n5347 , n5348 , n5349 , n5350 , n5351 , n5352 , n5353 , n5354 , n5355 , n5356 , n5357 , n5358 , n5359 , n5360 , n5361 , n5362 , n5363 , n5364 , n5365 , n5366 , n5367 , n5368 , n5369 , n5370 ;
  assign n25 = x1 | x2 ;
  assign n26 = x0 | x3 ;
  assign n27 = n25 | n26 ;
  assign n28 = ~x22 & n27 ;
  assign n29 = ( x4 & ~x22 ) | ( x4 & n28 ) | ( ~x22 & n28 ) ;
  assign n30 = ~x5 & n29 ;
  assign n31 = x5 | n30 ;
  assign n32 = ( ~n29 & n30 ) | ( ~n29 & n31 ) | ( n30 & n31 ) ;
  assign n33 = x21 & x22 ;
  assign n34 = x4 | x5 ;
  assign n35 = x6 | n34 ;
  assign n36 = n27 | n35 ;
  assign n37 = x7 | x8 ;
  assign n38 = x9 | x10 ;
  assign n39 = n37 | n38 ;
  assign n40 = n36 | n39 ;
  assign n41 = x11 | x12 ;
  assign n42 = x13 | x14 ;
  assign n43 = n41 | n42 ;
  assign n44 = x15 | n43 ;
  assign n45 = n40 | n44 ;
  assign n46 = x16 | x17 ;
  assign n47 = x18 | x19 ;
  assign n48 = n46 | n47 ;
  assign n49 = x20 | n48 ;
  assign n50 = x21 & n49 ;
  assign n51 = ( x21 & n45 ) | ( x21 & n50 ) | ( n45 & n50 ) ;
  assign n52 = x20 | x21 ;
  assign n53 = ( ~n45 & n48 ) | ( ~n45 & n52 ) | ( n48 & n52 ) ;
  assign n54 = n45 | n53 ;
  assign n55 = ~n51 & n54 ;
  assign n56 = x22 & ~n33 ;
  assign n57 = ( n33 & n55 ) | ( n33 & ~n56 ) | ( n55 & ~n56 ) ;
  assign n58 = n40 | n48 ;
  assign n59 = ( ~x22 & n44 ) | ( ~x22 & n58 ) | ( n44 & n58 ) ;
  assign n60 = ( ~x20 & x22 ) | ( ~x20 & n59 ) | ( x22 & n59 ) ;
  assign n61 = n59 & ~n60 ;
  assign n62 = ~x22 & n60 ;
  assign n63 = ( x20 & ~n61 ) | ( x20 & n62 ) | ( ~n61 & n62 ) ;
  assign n64 = n57 | n63 ;
  assign n65 = ( ~x22 & n40 ) | ( ~x22 & n43 ) | ( n40 & n43 ) ;
  assign n66 = ( ~x15 & x22 ) | ( ~x15 & n65 ) | ( x22 & n65 ) ;
  assign n67 = n65 & ~n66 ;
  assign n68 = ~x22 & n66 ;
  assign n69 = ( x15 & ~n67 ) | ( x15 & n68 ) | ( ~n67 & n68 ) ;
  assign n70 = ~n64 & n69 ;
  assign n71 = x18 & ~x22 ;
  assign n72 = ( ~x22 & n46 ) | ( ~x22 & n71 ) | ( n46 & n71 ) ;
  assign n73 = x19 & ~n72 ;
  assign n74 = x19 & x22 ;
  assign n75 = ( ~n45 & n73 ) | ( ~n45 & n74 ) | ( n73 & n74 ) ;
  assign n76 = ( ~x22 & n40 ) | ( ~x22 & n44 ) | ( n40 & n44 ) ;
  assign n77 = ( ~x22 & n72 ) | ( ~x22 & n76 ) | ( n72 & n76 ) ;
  assign n78 = ( ~x19 & n74 ) | ( ~x19 & n77 ) | ( n74 & n77 ) ;
  assign n79 = n75 | n78 ;
  assign n80 = x18 & x22 ;
  assign n81 = n44 | n46 ;
  assign n82 = x18 & n40 ;
  assign n83 = ( x18 & n81 ) | ( x18 & n82 ) | ( n81 & n82 ) ;
  assign n84 = n77 & ~n83 ;
  assign n85 = n80 | n84 ;
  assign n86 = n79 | n85 ;
  assign n87 = ( ~x16 & x22 ) | ( ~x16 & n76 ) | ( x22 & n76 ) ;
  assign n88 = n76 & ~n87 ;
  assign n89 = ~x22 & n87 ;
  assign n90 = ( x16 & ~n88 ) | ( x16 & n89 ) | ( ~n88 & n89 ) ;
  assign n91 = ( x16 & ~x22 ) | ( x16 & n89 ) | ( ~x22 & n89 ) ;
  assign n92 = ~x17 & n91 ;
  assign n93 = x17 | n92 ;
  assign n94 = ( ~n91 & n92 ) | ( ~n91 & n93 ) | ( n92 & n93 ) ;
  assign n95 = ~n90 & n94 ;
  assign n96 = ~n86 & n95 ;
  assign n97 = n70 & n96 ;
  assign n98 = n64 | n69 ;
  assign n99 = ~n79 & n85 ;
  assign n100 = n95 & n99 ;
  assign n101 = ~n98 & n100 ;
  assign n102 = n97 | n101 ;
  assign n103 = n57 & ~n63 ;
  assign n104 = ~n69 & n103 ;
  assign n105 = n90 | n94 ;
  assign n106 = n79 & ~n85 ;
  assign n107 = ~n105 & n106 ;
  assign n108 = n104 & n107 ;
  assign n109 = n79 & n85 ;
  assign n110 = n95 & n109 ;
  assign n111 = n69 & n103 ;
  assign n112 = n110 & n111 ;
  assign n113 = n108 | n112 ;
  assign n114 = ~n57 & n63 ;
  assign n115 = ~n69 & n114 ;
  assign n116 = n110 & n115 ;
  assign n117 = n69 & n114 ;
  assign n118 = n90 & ~n94 ;
  assign n119 = n99 & n118 ;
  assign n120 = n117 & n119 ;
  assign n121 = n116 | n120 ;
  assign n122 = n113 | n121 ;
  assign n123 = n102 | n122 ;
  assign n124 = n86 | n105 ;
  assign n125 = n117 & ~n124 ;
  assign n126 = n99 & ~n105 ;
  assign n127 = n111 & n126 ;
  assign n128 = n111 & n119 ;
  assign n129 = n127 | n128 ;
  assign n130 = n125 | n129 ;
  assign n131 = ~n86 & n118 ;
  assign n132 = n115 & n131 ;
  assign n133 = n100 & n104 ;
  assign n134 = n117 & n131 ;
  assign n135 = n133 | n134 ;
  assign n136 = n132 | n135 ;
  assign n137 = n130 | n136 ;
  assign n138 = n123 | n137 ;
  assign n139 = n57 & n63 ;
  assign n140 = ~n69 & n139 ;
  assign n141 = n110 & n140 ;
  assign n142 = ~n105 & n109 ;
  assign n143 = n140 & n142 ;
  assign n144 = n141 | n143 ;
  assign n145 = n90 & n94 ;
  assign n146 = n109 & n145 ;
  assign n147 = n140 & n146 ;
  assign n148 = n109 & n118 ;
  assign n149 = n117 & n148 ;
  assign n150 = n147 | n149 ;
  assign n151 = n144 | n150 ;
  assign n152 = n115 & ~n124 ;
  assign n153 = n69 & n139 ;
  assign n154 = ~n124 & n153 ;
  assign n155 = n119 & n140 ;
  assign n156 = n154 | n155 ;
  assign n157 = n117 & n142 ;
  assign n158 = ~n124 & n140 ;
  assign n159 = n157 | n158 ;
  assign n160 = n156 | n159 ;
  assign n161 = n152 | n160 ;
  assign n162 = n151 | n161 ;
  assign n163 = n138 | n162 ;
  assign n164 = n107 & n117 ;
  assign n165 = n70 & n100 ;
  assign n166 = n164 | n165 ;
  assign n167 = n99 & n145 ;
  assign n168 = n70 & n167 ;
  assign n169 = n166 | n168 ;
  assign n170 = n163 | n169 ;
  assign n171 = n111 & n142 ;
  assign n172 = n106 & n118 ;
  assign n173 = n117 & n172 ;
  assign n174 = n171 | n173 ;
  assign n175 = n115 & n146 ;
  assign n176 = n70 & n172 ;
  assign n177 = n175 | n176 ;
  assign n178 = n174 | n177 ;
  assign n179 = n111 & n131 ;
  assign n180 = n104 & n172 ;
  assign n181 = n100 & n140 ;
  assign n182 = n180 | n181 ;
  assign n183 = n179 | n182 ;
  assign n184 = n178 | n183 ;
  assign n185 = n96 & ~n98 ;
  assign n186 = n115 & n119 ;
  assign n187 = n115 & n167 ;
  assign n188 = n186 | n187 ;
  assign n189 = n185 | n188 ;
  assign n190 = n184 | n189 ;
  assign n191 = n153 & n167 ;
  assign n192 = n111 & n167 ;
  assign n193 = n191 | n192 ;
  assign n194 = ~n86 & n145 ;
  assign n195 = n115 & n194 ;
  assign n196 = n106 & n145 ;
  assign n197 = n117 & n196 ;
  assign n198 = n195 | n197 ;
  assign n199 = n193 | n198 ;
  assign n200 = n70 & n146 ;
  assign n201 = ~n98 & n196 ;
  assign n202 = n200 | n201 ;
  assign n203 = n199 | n202 ;
  assign n204 = n104 & n167 ;
  assign n205 = n100 & n111 ;
  assign n206 = n204 | n205 ;
  assign n207 = n140 & n196 ;
  assign n208 = n95 & n106 ;
  assign n209 = n140 & n208 ;
  assign n210 = n207 | n209 ;
  assign n211 = n107 & n111 ;
  assign n212 = n140 & n148 ;
  assign n213 = n211 | n212 ;
  assign n214 = n210 | n213 ;
  assign n215 = n206 | n214 ;
  assign n216 = n203 | n215 ;
  assign n217 = n190 | n216 ;
  assign n218 = n70 & n131 ;
  assign n219 = n115 & n196 ;
  assign n220 = ~n98 & n194 ;
  assign n221 = n219 | n220 ;
  assign n222 = n218 | n221 ;
  assign n223 = n104 & n142 ;
  assign n224 = n104 & n110 ;
  assign n225 = n223 | n224 ;
  assign n226 = n111 & n196 ;
  assign n227 = n96 & n117 ;
  assign n228 = n226 | n227 ;
  assign n229 = n225 | n228 ;
  assign n230 = n222 | n229 ;
  assign n231 = ~n98 & n148 ;
  assign n232 = n117 & n146 ;
  assign n233 = n231 | n232 ;
  assign n234 = n70 & n142 ;
  assign n235 = n104 & n131 ;
  assign n236 = n104 & n119 ;
  assign n237 = n235 | n236 ;
  assign n238 = ~n98 & n119 ;
  assign n239 = n96 & n115 ;
  assign n240 = n238 | n239 ;
  assign n241 = n237 | n240 ;
  assign n242 = n234 | n241 ;
  assign n243 = n233 | n242 ;
  assign n244 = n230 | n243 ;
  assign n245 = n217 | n244 ;
  assign n246 = n170 | n245 ;
  assign n247 = n70 & n126 ;
  assign n248 = ~n98 & n146 ;
  assign n249 = n153 & n194 ;
  assign n250 = n96 & n140 ;
  assign n251 = n249 | n250 ;
  assign n252 = n70 & n107 ;
  assign n253 = n153 & n172 ;
  assign n254 = n252 | n253 ;
  assign n255 = n251 | n254 ;
  assign n256 = n117 & n167 ;
  assign n257 = n104 & n126 ;
  assign n258 = n107 & n153 ;
  assign n259 = n257 | n258 ;
  assign n260 = n256 | n259 ;
  assign n261 = n255 | n260 ;
  assign n262 = n248 | n261 ;
  assign n263 = n247 | n262 ;
  assign n264 = n246 | n263 ;
  assign n265 = n104 & n194 ;
  assign n266 = n235 | n265 ;
  assign n267 = n117 & n208 ;
  assign n268 = n232 | n267 ;
  assign n269 = n266 | n268 ;
  assign n270 = n116 | n269 ;
  assign n271 = n96 & n111 ;
  assign n272 = n179 | n271 ;
  assign n273 = n96 & n104 ;
  assign n274 = n111 & n194 ;
  assign n275 = n273 | n274 ;
  assign n276 = n133 | n175 ;
  assign n277 = n275 | n276 ;
  assign n278 = n272 | n277 ;
  assign n279 = n270 | n278 ;
  assign n280 = n104 & ~n124 ;
  assign n281 = n115 & n148 ;
  assign n282 = n149 | n157 ;
  assign n283 = n281 | n282 ;
  assign n284 = n110 & n117 ;
  assign n285 = n197 | n219 ;
  assign n286 = n284 | n285 ;
  assign n287 = n283 | n286 ;
  assign n288 = n280 | n287 ;
  assign n289 = n279 | n288 ;
  assign n290 = n111 & ~n124 ;
  assign n291 = n115 & n142 ;
  assign n292 = n290 | n291 ;
  assign n293 = n100 & n115 ;
  assign n294 = n120 | n187 ;
  assign n295 = n293 | n294 ;
  assign n296 = n100 & n117 ;
  assign n297 = n115 & n208 ;
  assign n298 = n256 | n297 ;
  assign n299 = n296 | n298 ;
  assign n300 = n295 | n299 ;
  assign n301 = ( n107 & n114 ) | ( n107 & n172 ) | ( n114 & n172 ) ;
  assign n302 = n300 | n301 ;
  assign n303 = n292 | n302 ;
  assign n304 = n289 | n303 ;
  assign n305 = n117 & n126 ;
  assign n306 = n132 | n305 ;
  assign n307 = n134 | n239 ;
  assign n308 = n306 | n307 ;
  assign n309 = ( n114 & n194 ) | ( n114 & n227 ) | ( n194 & n227 ) ;
  assign n310 = n308 | n309 ;
  assign n311 = n115 & n126 ;
  assign n312 = n236 | n257 ;
  assign n313 = n129 | n312 ;
  assign n314 = n311 | n313 ;
  assign n315 = n310 | n314 ;
  assign n316 = n186 | n315 ;
  assign n317 = n304 | n316 ;
  assign n318 = n289 | n292 ;
  assign n319 = n70 & n110 ;
  assign n320 = n152 | n319 ;
  assign n321 = n70 & n148 ;
  assign n322 = n234 | n321 ;
  assign n323 = n320 | n322 ;
  assign n324 = n130 | n323 ;
  assign n325 = ~n98 & n110 ;
  assign n326 = n248 | n325 ;
  assign n327 = n312 | n326 ;
  assign n328 = n324 | n327 ;
  assign n329 = n70 & n196 ;
  assign n330 = n200 | n231 ;
  assign n331 = ~n98 & n142 ;
  assign n332 = n201 | n331 ;
  assign n333 = n330 | n332 ;
  assign n334 = n329 | n333 ;
  assign n335 = n328 | n334 ;
  assign n336 = n70 & n208 ;
  assign n337 = n252 | n336 ;
  assign n338 = ~n98 & n208 ;
  assign n339 = ( ~n64 & n172 ) | ( ~n64 & n338 ) | ( n172 & n338 ) ;
  assign n340 = ( ~n335 & n337 ) | ( ~n335 & n339 ) | ( n337 & n339 ) ;
  assign n341 = n335 | n340 ;
  assign n342 = n318 | n341 ;
  assign n343 = n317 | n342 ;
  assign n344 = ~n342 & n343 ;
  assign n345 = ( ~n317 & n343 ) | ( ~n317 & n344 ) | ( n343 & n344 ) ;
  assign n346 = n108 | n191 ;
  assign n347 = n211 | n346 ;
  assign n348 = n140 & n167 ;
  assign n349 = n126 & n140 ;
  assign n350 = n348 | n349 ;
  assign n351 = n100 & n153 ;
  assign n352 = n180 | n351 ;
  assign n353 = n350 | n352 ;
  assign n354 = n347 | n353 ;
  assign n355 = n126 & n153 ;
  assign n356 = n111 & n172 ;
  assign n357 = n355 | n356 ;
  assign n358 = n354 | n357 ;
  assign n359 = n140 & n194 ;
  assign n360 = n171 | n359 ;
  assign n361 = n210 | n360 ;
  assign n362 = n111 & n148 ;
  assign n363 = n153 & n208 ;
  assign n364 = n249 | n363 ;
  assign n365 = n362 | n364 ;
  assign n366 = n361 | n365 ;
  assign n367 = n111 & n146 ;
  assign n368 = n158 | n367 ;
  assign n369 = n104 & n148 ;
  assign n370 = n223 | n369 ;
  assign n371 = n368 | n370 ;
  assign n372 = n366 | n371 ;
  assign n373 = n358 | n372 ;
  assign n374 = n154 | n253 ;
  assign n375 = n131 & n140 ;
  assign n376 = ( n64 & n141 ) | ( n64 & n375 ) | ( n141 & n375 ) ;
  assign n377 = ( n139 & n148 ) | ( n139 & n376 ) | ( n148 & n376 ) ;
  assign n378 = n374 | n377 ;
  assign n379 = n373 | n378 ;
  assign n380 = n107 & n140 ;
  assign n381 = n104 & n196 ;
  assign n382 = n380 | n381 ;
  assign n383 = n206 | n382 ;
  assign n384 = n119 & n153 ;
  assign n385 = n192 | n384 ;
  assign n386 = n140 & n172 ;
  assign n387 = n181 | n386 ;
  assign n388 = n385 | n387 ;
  assign n389 = n383 | n388 ;
  assign n390 = n104 & n208 ;
  assign n391 = n111 & n208 ;
  assign n392 = n390 | n391 ;
  assign n393 = n155 | n258 ;
  assign n394 = n392 | n393 ;
  assign n395 = n226 | n394 ;
  assign n396 = n389 | n395 ;
  assign n397 = n153 & n196 ;
  assign n398 = n143 | n397 ;
  assign n399 = n104 & n146 ;
  assign n400 = n142 & n153 ;
  assign n401 = n399 | n400 ;
  assign n402 = n398 | n401 ;
  assign n403 = n112 | n224 ;
  assign n404 = n110 & n153 ;
  assign n405 = n131 & n153 ;
  assign n406 = n404 | n405 ;
  assign n407 = n403 | n406 ;
  assign n408 = n402 | n407 ;
  assign n409 = n250 | n408 ;
  assign n410 = n396 | n409 ;
  assign n411 = n96 & n153 ;
  assign n412 = ( n139 & n146 ) | ( n139 & n411 ) | ( n146 & n411 ) ;
  assign n413 = n410 | n412 ;
  assign n414 = n379 | n413 ;
  assign n415 = n343 & ~n414 ;
  assign n416 = n345 & ~n415 ;
  assign n417 = ( ~n342 & n414 ) | ( ~n342 & n416 ) | ( n414 & n416 ) ;
  assign n418 = n345 | n417 ;
  assign n419 = x4 & n28 ;
  assign n420 = x4 & ~n419 ;
  assign n421 = ( n28 & ~n419 ) | ( n28 & n420 ) | ( ~n419 & n420 ) ;
  assign n422 = n418 | n421 ;
  assign n423 = n345 | n415 ;
  assign n424 = n421 & ~n423 ;
  assign n425 = n422 & ~n424 ;
  assign n426 = ( n32 & n416 ) | ( n32 & ~n425 ) | ( n416 & ~n425 ) ;
  assign n427 = n345 & ~n417 ;
  assign n428 = ( n32 & n425 ) | ( n32 & ~n427 ) | ( n425 & ~n427 ) ;
  assign n429 = ~n426 & n428 ;
  assign n430 = x0 & ~x22 ;
  assign n431 = ( ~x22 & n25 ) | ( ~x22 & n430 ) | ( n25 & n430 ) ;
  assign n432 = x3 & ~n431 ;
  assign n433 = ~x3 & n431 ;
  assign n434 = n432 | n433 ;
  assign n435 = n416 & n434 ;
  assign n436 = n223 | n265 ;
  assign n437 = n149 | n236 ;
  assign n438 = n436 | n437 ;
  assign n439 = n406 | n438 ;
  assign n440 = n351 | n390 ;
  assign n441 = n195 | n440 ;
  assign n442 = n113 | n441 ;
  assign n443 = n439 | n442 ;
  assign n444 = n231 | n280 ;
  assign n445 = n154 | n380 ;
  assign n446 = n444 | n445 ;
  assign n447 = n369 | n446 ;
  assign n448 = n443 | n447 ;
  assign n449 = n98 | n124 ;
  assign n450 = ~n274 & n449 ;
  assign n451 = n125 | n290 ;
  assign n452 = n450 & ~n451 ;
  assign n453 = n115 & n172 ;
  assign n454 = n152 | n453 ;
  assign n455 = n297 | n454 ;
  assign n456 = n452 & ~n455 ;
  assign n457 = n117 & n194 ;
  assign n458 = n248 | n457 ;
  assign n459 = n247 | n325 ;
  assign n460 = n168 | n234 ;
  assign n461 = n459 | n460 ;
  assign n462 = n458 | n461 ;
  assign n463 = n456 & ~n462 ;
  assign n464 = ~n448 & n463 ;
  assign n465 = n179 | n220 ;
  assign n466 = n381 | n384 ;
  assign n467 = n465 | n466 ;
  assign n468 = n271 | n356 ;
  assign n469 = n232 | n468 ;
  assign n470 = n467 | n469 ;
  assign n471 = ~n98 & n167 ;
  assign n472 = n175 | n471 ;
  assign n473 = n185 | n472 ;
  assign n474 = n470 | n473 ;
  assign n475 = n143 | n366 ;
  assign n476 = n474 | n475 ;
  assign n477 = n70 & n119 ;
  assign n478 = ~n98 & n126 ;
  assign n479 = n477 | n478 ;
  assign n480 = n155 | n305 ;
  assign n481 = ~n98 & n131 ;
  assign n482 = n120 | n481 ;
  assign n483 = n480 | n482 ;
  assign n484 = n479 | n483 ;
  assign n485 = n476 | n484 ;
  assign n486 = n464 & ~n485 ;
  assign n487 = x13 | x22 ;
  assign n488 = n41 & ~n487 ;
  assign n489 = ( n40 & ~n487 ) | ( n40 & n488 ) | ( ~n487 & n488 ) ;
  assign n490 = ~x22 & n40 ;
  assign n491 = ( ~x22 & n41 ) | ( ~x22 & n490 ) | ( n41 & n490 ) ;
  assign n492 = ( x13 & n488 ) | ( x13 & ~n491 ) | ( n488 & ~n491 ) ;
  assign n493 = n489 | n492 ;
  assign n494 = n112 | n227 ;
  assign n495 = n281 | n471 ;
  assign n496 = n494 | n495 ;
  assign n497 = ~n493 & n496 ;
  assign n498 = ~n356 & n449 ;
  assign n499 = n155 | n384 ;
  assign n500 = n102 | n499 ;
  assign n501 = n248 | n500 ;
  assign n502 = n355 | n411 ;
  assign n503 = n176 | n478 ;
  assign n504 = n181 | n211 ;
  assign n505 = n503 | n504 ;
  assign n506 = n502 | n505 ;
  assign n507 = n501 | n506 ;
  assign n508 = n498 & ~n507 ;
  assign n509 = n305 | n319 ;
  assign n510 = n392 | n509 ;
  assign n511 = n267 | n285 ;
  assign n512 = n510 | n511 ;
  assign n513 = n148 & n153 ;
  assign n514 = n252 | n513 ;
  assign n515 = n275 | n514 ;
  assign n516 = n154 | n223 ;
  assign n517 = n256 | n516 ;
  assign n518 = n515 | n517 ;
  assign n519 = n70 & ~n124 ;
  assign n520 = n239 | n519 ;
  assign n521 = n518 | n520 ;
  assign n522 = n512 | n521 ;
  assign n523 = n508 & ~n522 ;
  assign n524 = n291 | n296 ;
  assign n525 = n143 | n257 ;
  assign n526 = n524 | n525 ;
  assign n527 = n271 | n477 ;
  assign n528 = n191 | n527 ;
  assign n529 = n526 | n528 ;
  assign n530 = n127 | n180 ;
  assign n531 = n157 | n164 ;
  assign n532 = n530 | n531 ;
  assign n533 = n329 | n532 ;
  assign n534 = n529 | n533 ;
  assign n535 = n523 & ~n534 ;
  assign n536 = n224 | n290 ;
  assign n537 = n185 | n536 ;
  assign n538 = n265 | n400 ;
  assign n539 = n231 | n453 ;
  assign n540 = n538 | n539 ;
  assign n541 = n537 | n540 ;
  assign n542 = n136 | n541 ;
  assign n543 = n349 | n375 ;
  assign n544 = n146 & n153 ;
  assign n545 = n258 | n544 ;
  assign n546 = n543 | n545 ;
  assign n547 = n369 | n546 ;
  assign n548 = n186 | n284 ;
  assign n549 = n147 | n204 ;
  assign n550 = n232 | n336 ;
  assign n551 = n549 | n550 ;
  assign n552 = ( ~n547 & n548 ) | ( ~n547 & n551 ) | ( n548 & n551 ) ;
  assign n553 = n547 | n552 ;
  assign n554 = n542 | n553 ;
  assign n555 = n359 | n554 ;
  assign n556 = n535 & ~n555 ;
  assign n557 = ( n493 & ~n497 ) | ( n493 & n556 ) | ( ~n497 & n556 ) ;
  assign n558 = n486 & ~n557 ;
  assign n559 = x14 & x22 ;
  assign n560 = x22 & ~n559 ;
  assign n561 = x13 & x14 ;
  assign n562 = ( x14 & n41 ) | ( x14 & n561 ) | ( n41 & n561 ) ;
  assign n563 = ( x14 & n40 ) | ( x14 & n562 ) | ( n40 & n562 ) ;
  assign n564 = n43 & ~n563 ;
  assign n565 = ( n40 & ~n563 ) | ( n40 & n564 ) | ( ~n563 & n564 ) ;
  assign n566 = ( n559 & ~n560 ) | ( n559 & n565 ) | ( ~n560 & n565 ) ;
  assign n567 = n496 | n555 ;
  assign n568 = n535 & ~n567 ;
  assign n569 = n566 & ~n568 ;
  assign n570 = ( n486 & ~n566 ) | ( n486 & n568 ) | ( ~n566 & n568 ) ;
  assign n571 = ( ~n558 & n569 ) | ( ~n558 & n570 ) | ( n569 & n570 ) ;
  assign n572 = n417 & ~n571 ;
  assign n573 = ~n435 & n572 ;
  assign n574 = n429 & n573 ;
  assign n575 = n429 | n573 ;
  assign n576 = ~n574 & n575 ;
  assign n577 = n70 & n194 ;
  assign n578 = n257 | n477 ;
  assign n579 = n247 | n578 ;
  assign n580 = n233 | n579 ;
  assign n581 = n258 | n348 ;
  assign n582 = n133 | n390 ;
  assign n583 = n581 | n582 ;
  assign n584 = n186 | n223 ;
  assign n585 = n583 | n584 ;
  assign n586 = n580 | n585 ;
  assign n587 = n108 | n359 ;
  assign n588 = n166 | n587 ;
  assign n589 = n116 | n588 ;
  assign n590 = n586 | n589 ;
  assign n591 = n154 | n355 ;
  assign n592 = n296 | n591 ;
  assign n593 = n235 | n271 ;
  assign n594 = n362 | n593 ;
  assign n595 = n592 | n594 ;
  assign n596 = n203 | n595 ;
  assign n597 = ~n98 & n172 ;
  assign n598 = n471 | n597 ;
  assign n599 = n596 | n598 ;
  assign n600 = n590 | n599 ;
  assign n601 = n134 | n380 ;
  assign n602 = n293 | n453 ;
  assign n603 = n601 | n602 ;
  assign n604 = ~n98 & n107 ;
  assign n605 = n319 | n604 ;
  assign n606 = n603 | n605 ;
  assign n607 = n226 | n356 ;
  assign n608 = n218 | n297 ;
  assign n609 = n607 | n608 ;
  assign n610 = n130 | n609 ;
  assign n611 = n606 | n610 ;
  assign n612 = n256 | n386 ;
  assign n613 = n157 | n227 ;
  assign n614 = n612 | n613 ;
  assign n615 = n325 | n614 ;
  assign n616 = n97 | n615 ;
  assign n617 = n611 | n616 ;
  assign n618 = n158 | n375 ;
  assign n619 = n249 | n311 ;
  assign n620 = n618 | n619 ;
  assign n621 = n281 | n331 ;
  assign n622 = n338 | n621 ;
  assign n623 = n620 | n622 ;
  assign n624 = n349 | n519 ;
  assign n625 = ( ~n403 & n623 ) | ( ~n403 & n624 ) | ( n623 & n624 ) ;
  assign n626 = n403 | n625 ;
  assign n627 = n617 | n626 ;
  assign n628 = n600 | n627 ;
  assign n629 = n577 | n628 ;
  assign n630 = n465 | n527 ;
  assign n631 = n481 | n548 ;
  assign n632 = n630 | n631 ;
  assign n633 = n157 | n338 ;
  assign n634 = n227 | n633 ;
  assign n635 = n604 | n634 ;
  assign n636 = n632 | n635 ;
  assign n637 = n213 | n636 ;
  assign n638 = n320 | n502 ;
  assign n639 = n133 | n236 ;
  assign n640 = n397 | n639 ;
  assign n641 = n638 | n640 ;
  assign n642 = n168 | n641 ;
  assign n643 = n210 | n406 ;
  assign n644 = n298 | n349 ;
  assign n645 = n643 | n644 ;
  assign n646 = n141 | n359 ;
  assign n647 = n128 | n187 ;
  assign n648 = n646 | n647 ;
  assign n649 = n238 | n648 ;
  assign n650 = n544 | n649 ;
  assign n651 = n645 | n650 ;
  assign n652 = n642 | n651 ;
  assign n653 = n637 | n652 ;
  assign n654 = n356 | n400 ;
  assign n655 = n180 | n362 ;
  assign n656 = n654 | n655 ;
  assign n657 = n291 | n513 ;
  assign n658 = n331 | n657 ;
  assign n659 = n143 | n253 ;
  assign n660 = n232 | n659 ;
  assign n661 = n658 | n660 ;
  assign n662 = n250 | n363 ;
  assign n663 = n273 | n662 ;
  assign n664 = n178 | n663 ;
  assign n665 = n661 | n664 ;
  assign n666 = n249 | n390 ;
  assign n667 = n112 | n369 ;
  assign n668 = n666 | n667 ;
  assign n669 = n195 | n668 ;
  assign n670 = n665 | n669 ;
  assign n671 = n325 | n670 ;
  assign n672 = n656 | n671 ;
  assign n673 = n653 | n672 ;
  assign n674 = n224 | n281 ;
  assign n675 = n321 | n577 ;
  assign n676 = n674 | n675 ;
  assign n677 = n147 | n305 ;
  assign n678 = n125 | n677 ;
  assign n679 = n676 | n678 ;
  assign n680 = n218 | n329 ;
  assign n681 = n239 | n680 ;
  assign n682 = n679 | n681 ;
  assign n683 = n673 | n682 ;
  assign n684 = n629 | n683 ;
  assign n685 = ~n683 & n684 ;
  assign n686 = ( ~n629 & n684 ) | ( ~n629 & n685 ) | ( n684 & n685 ) ;
  assign n687 = n232 | n274 ;
  assign n688 = n331 | n687 ;
  assign n689 = n226 | n351 ;
  assign n690 = n127 | n689 ;
  assign n691 = n380 | n690 ;
  assign n692 = n688 | n691 ;
  assign n693 = n168 | n404 ;
  assign n694 = n210 | n693 ;
  assign n695 = n116 | n212 ;
  assign n696 = n548 | n695 ;
  assign n697 = n694 | n696 ;
  assign n698 = ( n139 & n167 ) | ( n139 & n387 ) | ( n167 & n387 ) ;
  assign n699 = n697 | n698 ;
  assign n700 = n112 | n253 ;
  assign n701 = n165 | n700 ;
  assign n702 = n258 | n701 ;
  assign n703 = n311 | n702 ;
  assign n704 = n699 | n703 ;
  assign n705 = n107 & n115 ;
  assign n706 = n453 | n705 ;
  assign n707 = n677 | n706 ;
  assign n708 = n336 | n707 ;
  assign n709 = n164 | n175 ;
  assign n710 = n152 | n709 ;
  assign n711 = n171 | n220 ;
  assign n712 = n710 | n711 ;
  assign n713 = n438 | n712 ;
  assign n714 = n708 | n713 ;
  assign n715 = n704 | n714 ;
  assign n716 = n692 | n715 ;
  assign n717 = n362 | n369 ;
  assign n718 = n329 | n717 ;
  assign n719 = n397 | n544 ;
  assign n720 = n363 | n719 ;
  assign n721 = n319 | n457 ;
  assign n722 = n97 | n577 ;
  assign n723 = n721 | n722 ;
  assign n724 = ( n90 & n200 ) | ( n90 & n723 ) | ( n200 & n723 ) ;
  assign n725 = n720 | n724 ;
  assign n726 = n718 | n725 ;
  assign n727 = n501 | n726 ;
  assign n728 = n133 | n185 ;
  assign n729 = n400 | n513 ;
  assign n730 = n525 | n729 ;
  assign n731 = n125 | n381 ;
  assign n732 = n173 | n731 ;
  assign n733 = n730 | n732 ;
  assign n734 = n201 | n733 ;
  assign n735 = n141 | n734 ;
  assign n736 = n728 | n735 ;
  assign n737 = n727 | n736 ;
  assign n738 = n471 | n604 ;
  assign n739 = n224 | n391 ;
  assign n740 = n128 | n604 ;
  assign n741 = n739 | n740 ;
  assign n742 = n297 | n741 ;
  assign n743 = ( ~n604 & n738 ) | ( ~n604 & n742 ) | ( n738 & n742 ) ;
  assign n744 = n737 | n743 ;
  assign n745 = n716 | n744 ;
  assign n746 = ( ~n629 & n685 ) | ( ~n629 & n745 ) | ( n685 & n745 ) ;
  assign n747 = n686 & ~n746 ;
  assign n748 = ( x7 & ~x22 ) | ( x7 & n36 ) | ( ~x22 & n36 ) ;
  assign n749 = ( x8 & x22 ) | ( x8 & n748 ) | ( x22 & n748 ) ;
  assign n750 = n748 & ~n749 ;
  assign n751 = ~x22 & n749 ;
  assign n752 = ( x8 & n750 ) | ( x8 & ~n751 ) | ( n750 & ~n751 ) ;
  assign n753 = ~x22 & n36 ;
  assign n754 = x7 & n753 ;
  assign n755 = x7 & ~n754 ;
  assign n756 = ( n753 & ~n754 ) | ( n753 & n755 ) | ( ~n754 & n755 ) ;
  assign n757 = n686 | n746 ;
  assign n758 = n756 | n757 ;
  assign n759 = n684 & ~n745 ;
  assign n760 = n686 | n759 ;
  assign n761 = n756 & ~n760 ;
  assign n762 = n758 & ~n761 ;
  assign n763 = ( ~n747 & n752 ) | ( ~n747 & n762 ) | ( n752 & n762 ) ;
  assign n764 = n686 & ~n759 ;
  assign n765 = ( n752 & ~n762 ) | ( n752 & n764 ) | ( ~n762 & n764 ) ;
  assign n766 = n763 & ~n765 ;
  assign n767 = n387 | n459 ;
  assign n768 = n125 | n351 ;
  assign n769 = ( n69 & n253 ) | ( n69 & n768 ) | ( n253 & n768 ) ;
  assign n770 = n767 | n769 ;
  assign n771 = n164 | n293 ;
  assign n772 = n101 | n771 ;
  assign n773 = n770 | n772 ;
  assign n774 = n375 | n380 ;
  assign n775 = n705 | n774 ;
  assign n776 = n173 | n191 ;
  assign n777 = n156 | n776 ;
  assign n778 = n234 | n265 ;
  assign n779 = n604 | n778 ;
  assign n780 = n777 | n779 ;
  assign n781 = n775 | n780 ;
  assign n782 = n773 | n781 ;
  assign n783 = n652 | n782 ;
  assign n784 = n235 | n367 ;
  assign n785 = n212 | n784 ;
  assign n786 = n663 | n785 ;
  assign n787 = n200 | n384 ;
  assign n788 = n165 | n787 ;
  assign n789 = n249 | n788 ;
  assign n790 = n786 | n789 ;
  assign n791 = n321 | n581 ;
  assign n792 = n179 | n525 ;
  assign n793 = n791 | n792 ;
  assign n794 = n444 | n793 ;
  assign n795 = n790 | n794 ;
  assign n796 = n453 | n513 ;
  assign n797 = n158 | n399 ;
  assign n798 = n796 | n797 ;
  assign n799 = n147 | n400 ;
  assign n800 = n271 | n799 ;
  assign n801 = n798 | n800 ;
  assign n802 = n296 | n801 ;
  assign n803 = n127 | n290 ;
  assign n804 = n479 | n803 ;
  assign n805 = n802 | n804 ;
  assign n806 = n795 | n805 ;
  assign n807 = n783 | n806 ;
  assign n808 = n120 | n274 ;
  assign n809 = n248 | n471 ;
  assign n810 = n808 | n809 ;
  assign n811 = n807 | n810 ;
  assign n812 = n745 & n811 ;
  assign n813 = n342 & ~n812 ;
  assign n814 = n745 | n811 ;
  assign n815 = ~n811 & n814 ;
  assign n816 = ( ~n745 & n814 ) | ( ~n745 & n815 ) | ( n814 & n815 ) ;
  assign n817 = ~n813 & n816 ;
  assign n818 = ( ~x22 & n27 ) | ( ~x22 & n34 ) | ( n27 & n34 ) ;
  assign n819 = ( ~x6 & x22 ) | ( ~x6 & n818 ) | ( x22 & n818 ) ;
  assign n820 = n818 & ~n819 ;
  assign n821 = ~x22 & n819 ;
  assign n822 = ( x6 & ~n820 ) | ( x6 & n821 ) | ( ~n820 & n821 ) ;
  assign n823 = n813 | n816 ;
  assign n824 = n32 | n823 ;
  assign n825 = ~n342 & n814 ;
  assign n826 = n816 | n825 ;
  assign n827 = n32 & ~n826 ;
  assign n828 = n824 & ~n827 ;
  assign n829 = ( ~n817 & n822 ) | ( ~n817 & n828 ) | ( n822 & n828 ) ;
  assign n830 = n816 & ~n825 ;
  assign n831 = ( n822 & ~n828 ) | ( n822 & n830 ) | ( ~n828 & n830 ) ;
  assign n832 = n829 & ~n831 ;
  assign n833 = n306 | n690 ;
  assign n834 = n355 | n404 ;
  assign n835 = n604 | n834 ;
  assign n836 = n219 | n544 ;
  assign n837 = n319 | n836 ;
  assign n838 = n835 | n837 ;
  assign n839 = n833 | n838 ;
  assign n840 = n112 | n218 ;
  assign n841 = n234 | n840 ;
  assign n842 = ( n257 & n391 ) | ( n257 & ~n516 ) | ( n391 & ~n516 ) ;
  assign n843 = n516 | n842 ;
  assign n844 = n841 | n843 ;
  assign n845 = n498 & ~n844 ;
  assign n846 = ~n839 & n845 ;
  assign n847 = n204 | n386 ;
  assign n848 = n796 | n847 ;
  assign n849 = n724 | n848 ;
  assign n850 = n220 | n297 ;
  assign n851 = n248 | n850 ;
  assign n852 = ( ~n347 & n363 ) | ( ~n347 & n851 ) | ( n363 & n851 ) ;
  assign n853 = n347 | n852 ;
  assign n854 = n849 | n853 ;
  assign n855 = n252 | n273 ;
  assign n856 = n175 | n597 ;
  assign n857 = n855 | n856 ;
  assign n858 = n180 | n249 ;
  assign n859 = n857 | n858 ;
  assign n860 = n186 | n859 ;
  assign n861 = n854 | n860 ;
  assign n862 = n846 & ~n861 ;
  assign n863 = n141 | n411 ;
  assign n864 = n205 | n863 ;
  assign n865 = n195 | n705 ;
  assign n866 = n385 | n865 ;
  assign n867 = n864 | n866 ;
  assign n868 = n232 | n399 ;
  assign n869 = n867 | n868 ;
  assign n870 = n281 | n290 ;
  assign n871 = n695 | n870 ;
  assign n872 = n97 | n471 ;
  assign n873 = n329 | n872 ;
  assign n874 = n871 | n873 ;
  assign n875 = n331 | n381 ;
  assign n876 = n375 | n390 ;
  assign n877 = n875 | n876 ;
  assign n878 = n519 | n524 ;
  assign n879 = n877 | n878 ;
  assign n880 = n874 | n879 ;
  assign n881 = n869 | n880 ;
  assign n882 = n147 | n207 ;
  assign n883 = n171 | n256 ;
  assign n884 = n882 | n883 ;
  assign n885 = n134 | n168 ;
  assign n886 = n884 | n885 ;
  assign n887 = n881 | n886 ;
  assign n888 = n271 | n887 ;
  assign n889 = n862 & ~n888 ;
  assign n890 = n367 | n481 ;
  assign n891 = n185 | n890 ;
  assign n892 = n889 & ~n891 ;
  assign n893 = n113 | n338 ;
  assign n894 = n200 | n336 ;
  assign n895 = n212 | n894 ;
  assign n896 = n893 | n895 ;
  assign n897 = n204 | n290 ;
  assign n898 = n195 | n897 ;
  assign n899 = n896 | n898 ;
  assign n900 = n219 | n296 ;
  assign n901 = n127 | n381 ;
  assign n902 = n900 | n901 ;
  assign n903 = n201 | n738 ;
  assign n904 = n902 | n903 ;
  assign n905 = n387 | n904 ;
  assign n906 = n899 | n905 ;
  assign n907 = n151 | n784 ;
  assign n908 = n547 | n907 ;
  assign n909 = n250 | n513 ;
  assign n910 = n857 | n909 ;
  assign n911 = n674 | n768 ;
  assign n912 = n176 | n380 ;
  assign n913 = n400 | n912 ;
  assign n914 = n911 | n913 ;
  assign n915 = n910 | n914 ;
  assign n916 = n908 | n915 ;
  assign n917 = n906 | n916 ;
  assign n918 = n223 | n390 ;
  assign n919 = n457 | n918 ;
  assign n920 = n173 | n197 ;
  assign n921 = ( n69 & n274 ) | ( n69 & n920 ) | ( n274 & n920 ) ;
  assign n922 = n404 | n921 ;
  assign n923 = n919 | n922 ;
  assign n924 = n187 | n311 ;
  assign n925 = n923 | n924 ;
  assign n926 = n642 | n925 ;
  assign n927 = n180 | n453 ;
  assign n928 = n926 | n927 ;
  assign n929 = n917 | n928 ;
  assign n930 = n248 | n929 ;
  assign n931 = n892 & ~n930 ;
  assign n932 = n930 | n931 ;
  assign n933 = ( ~n892 & n931 ) | ( ~n892 & n932 ) | ( n931 & n932 ) ;
  assign n934 = n629 | n931 ;
  assign n935 = ~n933 & n934 ;
  assign n936 = ( n629 & n892 ) | ( n629 & n935 ) | ( n892 & n935 ) ;
  assign n937 = n933 | n936 ;
  assign n938 = x10 & x22 ;
  assign n939 = x10 & ~n938 ;
  assign n940 = ( x9 & n37 ) | ( x9 & n939 ) | ( n37 & n939 ) ;
  assign n941 = n939 & n940 ;
  assign n942 = ( n36 & n939 ) | ( n36 & n941 ) | ( n939 & n941 ) ;
  assign n943 = ( n490 & n938 ) | ( n490 & ~n942 ) | ( n938 & ~n942 ) ;
  assign n944 = ( ~x22 & n36 ) | ( ~x22 & n37 ) | ( n36 & n37 ) ;
  assign n945 = ( ~x9 & x22 ) | ( ~x9 & n944 ) | ( x22 & n944 ) ;
  assign n946 = n944 & ~n945 ;
  assign n947 = ~x22 & n945 ;
  assign n948 = ( x9 & ~n946 ) | ( x9 & n947 ) | ( ~n946 & n947 ) ;
  assign n949 = n933 & ~n936 ;
  assign n950 = ~n948 & n949 ;
  assign n951 = n933 & n934 ;
  assign n952 = n948 & n951 ;
  assign n953 = n950 | n952 ;
  assign n954 = ( n937 & n943 ) | ( n937 & ~n953 ) | ( n943 & ~n953 ) ;
  assign n955 = ( n935 & n943 ) | ( n935 & n953 ) | ( n943 & n953 ) ;
  assign n956 = n954 & ~n955 ;
  assign n957 = ( n766 & n832 ) | ( n766 & n956 ) | ( n832 & n956 ) ;
  assign n958 = n576 & n957 ;
  assign n959 = n576 | n957 ;
  assign n960 = ~n958 & n959 ;
  assign n961 = ~n752 & n949 ;
  assign n962 = n752 & n951 ;
  assign n963 = n961 | n962 ;
  assign n964 = ( n937 & n948 ) | ( n937 & ~n963 ) | ( n948 & ~n963 ) ;
  assign n965 = ( n935 & n948 ) | ( n935 & n963 ) | ( n948 & n963 ) ;
  assign n966 = n964 & ~n965 ;
  assign n967 = n757 | n822 ;
  assign n968 = ~n760 & n822 ;
  assign n969 = n967 & ~n968 ;
  assign n970 = ( ~n747 & n756 ) | ( ~n747 & n969 ) | ( n756 & n969 ) ;
  assign n971 = ( n756 & n764 ) | ( n756 & ~n969 ) | ( n764 & ~n969 ) ;
  assign n972 = n970 & ~n971 ;
  assign n973 = ( ~x22 & n36 ) | ( ~x22 & n39 ) | ( n36 & n39 ) ;
  assign n974 = ( ~x11 & x22 ) | ( ~x11 & n973 ) | ( x22 & n973 ) ;
  assign n975 = n973 & ~n974 ;
  assign n976 = ~x22 & n974 ;
  assign n977 = ( x11 & ~n975 ) | ( x11 & n976 ) | ( ~n975 & n976 ) ;
  assign n978 = n496 & ~n977 ;
  assign n979 = ( n556 & n977 ) | ( n556 & ~n978 ) | ( n977 & ~n978 ) ;
  assign n980 = n486 & n979 ;
  assign n981 = x12 & x22 ;
  assign n982 = ( x11 & x12 ) | ( x11 & ~n41 ) | ( x12 & ~n41 ) ;
  assign n983 = ( x12 & n40 ) | ( x12 & n982 ) | ( n40 & n982 ) ;
  assign n984 = n491 & ~n983 ;
  assign n985 = n981 | n984 ;
  assign n986 = ( ~n486 & n568 ) | ( ~n486 & n985 ) | ( n568 & n985 ) ;
  assign n987 = n568 & n985 ;
  assign n988 = ( n980 & n986 ) | ( n980 & ~n987 ) | ( n986 & ~n987 ) ;
  assign n989 = n813 & ~n988 ;
  assign n990 = n434 & n816 ;
  assign n991 = n989 & ~n990 ;
  assign n992 = ( n966 & n972 ) | ( n966 & n991 ) | ( n972 & n991 ) ;
  assign n993 = n496 & ~n985 ;
  assign n994 = ( n556 & n985 ) | ( n556 & ~n993 ) | ( n985 & ~n993 ) ;
  assign n995 = n486 & n994 ;
  assign n996 = ( ~n486 & n493 ) | ( ~n486 & n568 ) | ( n493 & n568 ) ;
  assign n997 = n493 & n568 ;
  assign n998 = ( n995 & n996 ) | ( n995 & ~n997 ) | ( n996 & ~n997 ) ;
  assign n999 = n718 | n893 ;
  assign n1000 = n449 & ~n999 ;
  assign n1001 = n797 | n875 ;
  assign n1002 = n154 | n405 ;
  assign n1003 = n133 | n1002 ;
  assign n1004 = n1001 | n1003 ;
  assign n1005 = n180 | n471 ;
  assign n1006 = n218 | n1005 ;
  assign n1007 = n1004 | n1006 ;
  assign n1008 = n1000 & ~n1007 ;
  assign n1009 = n211 | n226 ;
  assign n1010 = n129 | n1009 ;
  assign n1011 = n481 | n519 ;
  assign n1012 = n1010 | n1011 ;
  assign n1013 = n1008 & ~n1012 ;
  assign n1014 = n155 | n349 ;
  assign n1015 = n116 | n291 ;
  assign n1016 = n1014 | n1015 ;
  assign n1017 = n233 | n1016 ;
  assign n1018 = n283 | n298 ;
  assign n1019 = n1017 | n1018 ;
  assign n1020 = n168 | n247 ;
  assign n1021 = n239 | n311 ;
  assign n1022 = n808 | n1021 ;
  assign n1023 = n152 | n187 ;
  assign n1024 = n1022 | n1023 ;
  assign n1025 = n387 | n1024 ;
  assign n1026 = n1020 | n1025 ;
  assign n1027 = n1019 | n1026 ;
  assign n1028 = n1013 & ~n1027 ;
  assign n1029 = n207 | n249 ;
  assign n1030 = n132 | n1029 ;
  assign n1031 = n791 | n835 ;
  assign n1032 = n385 | n1031 ;
  assign n1033 = n512 | n1032 ;
  assign n1034 = n147 | n209 ;
  assign n1035 = n173 | n280 ;
  assign n1036 = n1034 | n1035 ;
  assign n1037 = n195 | n238 ;
  assign n1038 = n1036 | n1037 ;
  assign n1039 = n272 | n503 ;
  assign n1040 = n351 | n654 ;
  assign n1041 = n1039 | n1040 ;
  assign n1042 = n544 | n1041 ;
  assign n1043 = n141 | n1042 ;
  assign n1044 = n1038 | n1043 ;
  assign n1045 = n1033 | n1044 ;
  assign n1046 = n1030 | n1045 ;
  assign n1047 = n1028 & ~n1046 ;
  assign n1048 = n568 & n1047 ;
  assign n1049 = n568 & ~n1048 ;
  assign n1050 = ( n1047 & ~n1048 ) | ( n1047 & n1049 ) | ( ~n1048 & n1049 ) ;
  assign n1051 = n892 & ~n1048 ;
  assign n1052 = n1050 & ~n1051 ;
  assign n1053 = ( n568 & ~n892 ) | ( n568 & n1052 ) | ( ~n892 & n1052 ) ;
  assign n1054 = n1050 & ~n1053 ;
  assign n1055 = n1050 | n1053 ;
  assign n1056 = n943 | n1055 ;
  assign n1057 = n1050 | n1051 ;
  assign n1058 = n943 & ~n1057 ;
  assign n1059 = n1056 & ~n1058 ;
  assign n1060 = ( n977 & ~n1054 ) | ( n977 & n1059 ) | ( ~n1054 & n1059 ) ;
  assign n1061 = ( n977 & n1052 ) | ( n977 & ~n1059 ) | ( n1052 & ~n1059 ) ;
  assign n1062 = n1060 & ~n1061 ;
  assign n1063 = n421 | n823 ;
  assign n1064 = n421 & ~n826 ;
  assign n1065 = n1063 & ~n1064 ;
  assign n1066 = ( n32 & ~n817 ) | ( n32 & n1065 ) | ( ~n817 & n1065 ) ;
  assign n1067 = ( n32 & n830 ) | ( n32 & ~n1065 ) | ( n830 & ~n1065 ) ;
  assign n1068 = n1066 & ~n1067 ;
  assign n1069 = ( ~n998 & n1062 ) | ( ~n998 & n1068 ) | ( n1062 & n1068 ) ;
  assign n1070 = ( n766 & n956 ) | ( n766 & ~n957 ) | ( n956 & ~n957 ) ;
  assign n1071 = ( n832 & ~n957 ) | ( n832 & n1070 ) | ( ~n957 & n1070 ) ;
  assign n1072 = ( n992 & n1069 ) | ( n992 & n1071 ) | ( n1069 & n1071 ) ;
  assign n1073 = n960 & n1072 ;
  assign n1074 = n960 | n1072 ;
  assign n1075 = ~n1073 & n1074 ;
  assign n1076 = ~n943 & n949 ;
  assign n1077 = n943 & n951 ;
  assign n1078 = n1076 | n1077 ;
  assign n1079 = ( n937 & n977 ) | ( n937 & ~n1078 ) | ( n977 & ~n1078 ) ;
  assign n1080 = ( n935 & n977 ) | ( n935 & n1078 ) | ( n977 & n1078 ) ;
  assign n1081 = n1079 & ~n1080 ;
  assign n1082 = n752 | n757 ;
  assign n1083 = n752 & ~n760 ;
  assign n1084 = n1082 & ~n1083 ;
  assign n1085 = ( n764 & n948 ) | ( n764 & ~n1084 ) | ( n948 & ~n1084 ) ;
  assign n1086 = ( ~n747 & n948 ) | ( ~n747 & n1084 ) | ( n948 & n1084 ) ;
  assign n1087 = ~n1085 & n1086 ;
  assign n1088 = n822 | n823 ;
  assign n1089 = n822 & ~n826 ;
  assign n1090 = n1088 & ~n1089 ;
  assign n1091 = ( n756 & n830 ) | ( n756 & ~n1090 ) | ( n830 & ~n1090 ) ;
  assign n1092 = ( n756 & ~n817 ) | ( n756 & n1090 ) | ( ~n817 & n1090 ) ;
  assign n1093 = ~n1091 & n1092 ;
  assign n1094 = ( n1081 & n1087 ) | ( n1081 & n1093 ) | ( n1087 & n1093 ) ;
  assign n1095 = ( n1087 & n1093 ) | ( n1087 & ~n1094 ) | ( n1093 & ~n1094 ) ;
  assign n1096 = ( n1081 & ~n1094 ) | ( n1081 & n1095 ) | ( ~n1094 & n1095 ) ;
  assign n1097 = ~n484 & n566 ;
  assign n1098 = ~n476 & n1097 ;
  assign n1099 = n464 & n1098 ;
  assign n1100 = n412 & n434 ;
  assign n1101 = ( n414 & n434 ) | ( n414 & n1100 ) | ( n434 & n1100 ) ;
  assign n1102 = ~n1099 & n1101 ;
  assign n1103 = ~n568 & n1102 ;
  assign n1104 = n1099 & ~n1101 ;
  assign n1105 = ( n568 & ~n1101 ) | ( n568 & n1104 ) | ( ~n1101 & n1104 ) ;
  assign n1106 = n1103 | n1105 ;
  assign n1107 = n985 | n1055 ;
  assign n1108 = n985 & ~n1057 ;
  assign n1109 = n1107 & ~n1108 ;
  assign n1110 = ( n493 & n1052 ) | ( n493 & ~n1109 ) | ( n1052 & ~n1109 ) ;
  assign n1111 = ( n493 & ~n1054 ) | ( n493 & n1109 ) | ( ~n1054 & n1109 ) ;
  assign n1112 = ~n1110 & n1111 ;
  assign n1113 = ~n1106 & n1112 ;
  assign n1114 = n1106 & ~n1112 ;
  assign n1115 = n1113 | n1114 ;
  assign n1116 = ( ~n417 & n435 ) | ( ~n417 & n571 ) | ( n435 & n571 ) ;
  assign n1117 = n573 | n1116 ;
  assign n1118 = n977 | n1055 ;
  assign n1119 = n977 & ~n1057 ;
  assign n1120 = n1118 & ~n1119 ;
  assign n1121 = ( n985 & ~n1054 ) | ( n985 & n1120 ) | ( ~n1054 & n1120 ) ;
  assign n1122 = ( n985 & n1052 ) | ( n985 & ~n1120 ) | ( n1052 & ~n1120 ) ;
  assign n1123 = n1121 & ~n1122 ;
  assign n1124 = n418 | n434 ;
  assign n1125 = ~n423 & n434 ;
  assign n1126 = n1124 & ~n1125 ;
  assign n1127 = ( n416 & n421 ) | ( n416 & ~n1126 ) | ( n421 & ~n1126 ) ;
  assign n1128 = ( n421 & ~n427 ) | ( n421 & n1126 ) | ( ~n427 & n1126 ) ;
  assign n1129 = ~n1127 & n1128 ;
  assign n1130 = ( ~n1117 & n1123 ) | ( ~n1117 & n1129 ) | ( n1123 & n1129 ) ;
  assign n1131 = ~n1115 & n1130 ;
  assign n1132 = n1115 & ~n1130 ;
  assign n1133 = n1131 | n1132 ;
  assign n1134 = n1096 & ~n1133 ;
  assign n1135 = n1133 | n1134 ;
  assign n1136 = ( ~n1096 & n1134 ) | ( ~n1096 & n1135 ) | ( n1134 & n1135 ) ;
  assign n1137 = n1075 & ~n1136 ;
  assign n1138 = ~n1075 & n1136 ;
  assign n1139 = n1137 | n1138 ;
  assign n1140 = ( n345 & n434 ) | ( n345 & n435 ) | ( n434 & n435 ) ;
  assign n1141 = n948 | n1055 ;
  assign n1142 = n948 & ~n1057 ;
  assign n1143 = n1141 & ~n1142 ;
  assign n1144 = ( n943 & ~n1054 ) | ( n943 & n1143 ) | ( ~n1054 & n1143 ) ;
  assign n1145 = ( n943 & n1052 ) | ( n943 & ~n1143 ) | ( n1052 & ~n1143 ) ;
  assign n1146 = n1144 & ~n1145 ;
  assign n1147 = n32 | n757 ;
  assign n1148 = n32 & ~n760 ;
  assign n1149 = n1147 & ~n1148 ;
  assign n1150 = ( ~n747 & n822 ) | ( ~n747 & n1149 ) | ( n822 & n1149 ) ;
  assign n1151 = ( n764 & n822 ) | ( n764 & ~n1149 ) | ( n822 & ~n1149 ) ;
  assign n1152 = n1150 & ~n1151 ;
  assign n1153 = ~n756 & n949 ;
  assign n1154 = n756 & n951 ;
  assign n1155 = n1153 | n1154 ;
  assign n1156 = ( n752 & n937 ) | ( n752 & ~n1155 ) | ( n937 & ~n1155 ) ;
  assign n1157 = ( n752 & n935 ) | ( n752 & n1155 ) | ( n935 & n1155 ) ;
  assign n1158 = n1156 & ~n1157 ;
  assign n1159 = ( n1146 & n1152 ) | ( n1146 & n1158 ) | ( n1152 & n1158 ) ;
  assign n1160 = n1140 & n1159 ;
  assign n1161 = ( n972 & n991 ) | ( n972 & ~n992 ) | ( n991 & ~n992 ) ;
  assign n1162 = ( n966 & ~n992 ) | ( n966 & n1161 ) | ( ~n992 & n1161 ) ;
  assign n1163 = n1140 & ~n1160 ;
  assign n1164 = ( n1159 & ~n1160 ) | ( n1159 & n1163 ) | ( ~n1160 & n1163 ) ;
  assign n1165 = n1162 & n1164 ;
  assign n1166 = n1160 | n1165 ;
  assign n1167 = ( n992 & ~n1069 ) | ( n992 & n1071 ) | ( ~n1069 & n1071 ) ;
  assign n1168 = ( ~n992 & n1069 ) | ( ~n992 & n1167 ) | ( n1069 & n1167 ) ;
  assign n1169 = ( ~n1071 & n1167 ) | ( ~n1071 & n1168 ) | ( n1167 & n1168 ) ;
  assign n1170 = ( n1117 & ~n1123 ) | ( n1117 & n1130 ) | ( ~n1123 & n1130 ) ;
  assign n1171 = ( ~n1129 & n1130 ) | ( ~n1129 & n1170 ) | ( n1130 & n1170 ) ;
  assign n1172 = ( n1166 & n1169 ) | ( n1166 & ~n1171 ) | ( n1169 & ~n1171 ) ;
  assign n1173 = ~n1139 & n1172 ;
  assign n1174 = n1139 & ~n1172 ;
  assign n1175 = n1173 | n1174 ;
  assign n1176 = ( n434 & n813 ) | ( n434 & n823 ) | ( n813 & n823 ) ;
  assign n1177 = ( n988 & n990 ) | ( n988 & ~n1176 ) | ( n990 & ~n1176 ) ;
  assign n1178 = n991 | n1177 ;
  assign n1179 = n434 | n823 ;
  assign n1180 = n434 & ~n826 ;
  assign n1181 = n1179 & ~n1180 ;
  assign n1182 = ( n421 & ~n817 ) | ( n421 & n1181 ) | ( ~n817 & n1181 ) ;
  assign n1183 = ( n421 & n830 ) | ( n421 & ~n1181 ) | ( n830 & ~n1181 ) ;
  assign n1184 = n1182 & ~n1183 ;
  assign n1185 = n568 | n943 ;
  assign n1186 = n486 & n1185 ;
  assign n1187 = ( ~n486 & n568 ) | ( ~n486 & n977 ) | ( n568 & n977 ) ;
  assign n1188 = n568 & n977 ;
  assign n1189 = ( n1186 & n1187 ) | ( n1186 & ~n1188 ) | ( n1187 & ~n1188 ) ;
  assign n1190 = n752 | n1055 ;
  assign n1191 = n752 & ~n1057 ;
  assign n1192 = n1190 & ~n1191 ;
  assign n1193 = ( n948 & ~n1054 ) | ( n948 & n1192 ) | ( ~n1054 & n1192 ) ;
  assign n1194 = ( n948 & n1052 ) | ( n948 & ~n1192 ) | ( n1052 & ~n1192 ) ;
  assign n1195 = n1193 & ~n1194 ;
  assign n1196 = ~n822 & n949 ;
  assign n1197 = n822 & n951 ;
  assign n1198 = n1196 | n1197 ;
  assign n1199 = ( n756 & n935 ) | ( n756 & n1198 ) | ( n935 & n1198 ) ;
  assign n1200 = ( n756 & n937 ) | ( n756 & ~n1198 ) | ( n937 & ~n1198 ) ;
  assign n1201 = ~n1199 & n1200 ;
  assign n1202 = ( ~n1189 & n1195 ) | ( ~n1189 & n1201 ) | ( n1195 & n1201 ) ;
  assign n1203 = ( ~n1178 & n1184 ) | ( ~n1178 & n1202 ) | ( n1184 & n1202 ) ;
  assign n1204 = ( n998 & ~n1062 ) | ( n998 & n1069 ) | ( ~n1062 & n1069 ) ;
  assign n1205 = ( ~n1068 & n1069 ) | ( ~n1068 & n1204 ) | ( n1069 & n1204 ) ;
  assign n1206 = n1203 & ~n1205 ;
  assign n1207 = n1162 | n1164 ;
  assign n1208 = ~n1165 & n1207 ;
  assign n1209 = n1205 | n1206 ;
  assign n1210 = ( ~n1203 & n1206 ) | ( ~n1203 & n1209 ) | ( n1206 & n1209 ) ;
  assign n1211 = n1208 & ~n1210 ;
  assign n1212 = n1206 | n1211 ;
  assign n1213 = n421 | n757 ;
  assign n1214 = n421 & ~n760 ;
  assign n1215 = n1213 & ~n1214 ;
  assign n1216 = ( n32 & ~n747 ) | ( n32 & n1215 ) | ( ~n747 & n1215 ) ;
  assign n1217 = ( n32 & n764 ) | ( n32 & ~n1215 ) | ( n764 & ~n1215 ) ;
  assign n1218 = n1216 & ~n1217 ;
  assign n1219 = n568 | n948 ;
  assign n1220 = n486 & n1219 ;
  assign n1221 = ( n486 & n568 ) | ( n486 & n943 ) | ( n568 & n943 ) ;
  assign n1222 = ( n1185 & n1220 ) | ( n1185 & ~n1221 ) | ( n1220 & ~n1221 ) ;
  assign n1223 = n434 & n764 ;
  assign n1224 = ( n434 & n746 ) | ( n434 & n757 ) | ( n746 & n757 ) ;
  assign n1225 = ~n1223 & n1224 ;
  assign n1226 = n746 & n1225 ;
  assign n1227 = n1222 & ~n1226 ;
  assign n1228 = ( ~n1222 & n1226 ) | ( ~n1222 & n1227 ) | ( n1226 & n1227 ) ;
  assign n1229 = ( n990 & n1218 ) | ( n990 & n1228 ) | ( n1218 & n1228 ) ;
  assign n1230 = ( n1146 & n1158 ) | ( n1146 & ~n1159 ) | ( n1158 & ~n1159 ) ;
  assign n1231 = ( n1152 & ~n1159 ) | ( n1152 & n1230 ) | ( ~n1159 & n1230 ) ;
  assign n1232 = ( n1178 & ~n1202 ) | ( n1178 & n1203 ) | ( ~n1202 & n1203 ) ;
  assign n1233 = ( ~n1184 & n1203 ) | ( ~n1184 & n1232 ) | ( n1203 & n1232 ) ;
  assign n1234 = ( n1229 & n1231 ) | ( n1229 & ~n1233 ) | ( n1231 & ~n1233 ) ;
  assign n1235 = n756 | n1055 ;
  assign n1236 = n756 & ~n1057 ;
  assign n1237 = n1235 & ~n1236 ;
  assign n1238 = ( n752 & ~n1054 ) | ( n752 & n1237 ) | ( ~n1054 & n1237 ) ;
  assign n1239 = ( n752 & n1052 ) | ( n752 & ~n1237 ) | ( n1052 & ~n1237 ) ;
  assign n1240 = n1238 & ~n1239 ;
  assign n1241 = ~n32 & n949 ;
  assign n1242 = n32 & n951 ;
  assign n1243 = n1241 | n1242 ;
  assign n1244 = ( n822 & n935 ) | ( n822 & n1243 ) | ( n935 & n1243 ) ;
  assign n1245 = ( n822 & n937 ) | ( n822 & ~n1243 ) | ( n937 & ~n1243 ) ;
  assign n1246 = ~n1244 & n1245 ;
  assign n1247 = n434 | n757 ;
  assign n1248 = n434 & ~n760 ;
  assign n1249 = n1247 & ~n1248 ;
  assign n1250 = ( n421 & ~n747 ) | ( n421 & n1249 ) | ( ~n747 & n1249 ) ;
  assign n1251 = ( n421 & n764 ) | ( n421 & ~n1249 ) | ( n764 & ~n1249 ) ;
  assign n1252 = n1250 & ~n1251 ;
  assign n1253 = ( n1240 & n1246 ) | ( n1240 & n1252 ) | ( n1246 & n1252 ) ;
  assign n1254 = ( n1189 & ~n1195 ) | ( n1189 & n1202 ) | ( ~n1195 & n1202 ) ;
  assign n1255 = ( ~n1201 & n1202 ) | ( ~n1201 & n1254 ) | ( n1202 & n1254 ) ;
  assign n1256 = n1253 & ~n1255 ;
  assign n1257 = n1255 | n1256 ;
  assign n1258 = n1253 & n1255 ;
  assign n1259 = ( n990 & n1228 ) | ( n990 & ~n1229 ) | ( n1228 & ~n1229 ) ;
  assign n1260 = ( n1218 & ~n1229 ) | ( n1218 & n1259 ) | ( ~n1229 & n1259 ) ;
  assign n1261 = ( ~n1257 & n1258 ) | ( ~n1257 & n1260 ) | ( n1258 & n1260 ) ;
  assign n1262 = n1256 | n1261 ;
  assign n1263 = n1227 | n1228 ;
  assign n1264 = n568 | n752 ;
  assign n1265 = n486 & n1264 ;
  assign n1266 = ( n486 & n568 ) | ( n486 & n948 ) | ( n568 & n948 ) ;
  assign n1267 = ( n1219 & n1265 ) | ( n1219 & ~n1266 ) | ( n1265 & ~n1266 ) ;
  assign n1268 = n822 | n1055 ;
  assign n1269 = n822 & ~n1057 ;
  assign n1270 = n1268 & ~n1269 ;
  assign n1271 = ( n756 & ~n1054 ) | ( n756 & n1270 ) | ( ~n1054 & n1270 ) ;
  assign n1272 = ( n756 & n1052 ) | ( n756 & ~n1270 ) | ( n1052 & ~n1270 ) ;
  assign n1273 = n1271 & ~n1272 ;
  assign n1274 = ~n421 & n949 ;
  assign n1275 = n421 & n951 ;
  assign n1276 = n1274 | n1275 ;
  assign n1277 = ( n32 & n935 ) | ( n32 & n1276 ) | ( n935 & n1276 ) ;
  assign n1278 = ( n32 & n937 ) | ( n32 & ~n1276 ) | ( n937 & ~n1276 ) ;
  assign n1279 = ~n1277 & n1278 ;
  assign n1280 = ( ~n1267 & n1273 ) | ( ~n1267 & n1279 ) | ( n1273 & n1279 ) ;
  assign n1281 = ~n1263 & n1280 ;
  assign n1282 = n1263 & ~n1280 ;
  assign n1283 = n1281 | n1282 ;
  assign n1284 = ( n1240 & n1252 ) | ( n1240 & ~n1253 ) | ( n1252 & ~n1253 ) ;
  assign n1285 = ( n1246 & ~n1253 ) | ( n1246 & n1284 ) | ( ~n1253 & n1284 ) ;
  assign n1286 = ~n1283 & n1285 ;
  assign n1287 = n1281 | n1286 ;
  assign n1288 = n568 | n756 ;
  assign n1289 = n486 & n1288 ;
  assign n1290 = ( n486 & n568 ) | ( n486 & n752 ) | ( n568 & n752 ) ;
  assign n1291 = ( n1264 & n1289 ) | ( n1264 & ~n1290 ) | ( n1289 & ~n1290 ) ;
  assign n1292 = n936 & ~n1291 ;
  assign n1293 = n434 & ~n933 ;
  assign n1294 = n1292 & ~n1293 ;
  assign n1295 = ( n746 & ~n1225 ) | ( n746 & n1294 ) | ( ~n1225 & n1294 ) ;
  assign n1296 = ( ~n746 & n1225 ) | ( ~n746 & n1295 ) | ( n1225 & n1295 ) ;
  assign n1297 = ( ~n1294 & n1295 ) | ( ~n1294 & n1296 ) | ( n1295 & n1296 ) ;
  assign n1298 = ( n937 & ~n949 ) | ( n937 & n1293 ) | ( ~n949 & n1293 ) ;
  assign n1299 = ( n1291 & n1293 ) | ( n1291 & ~n1298 ) | ( n1293 & ~n1298 ) ;
  assign n1300 = n1294 | n1299 ;
  assign n1301 = n32 | n1055 ;
  assign n1302 = n32 & ~n1057 ;
  assign n1303 = n1301 & ~n1302 ;
  assign n1304 = ( n822 & ~n1054 ) | ( n822 & n1303 ) | ( ~n1054 & n1303 ) ;
  assign n1305 = ( n822 & n1052 ) | ( n822 & ~n1303 ) | ( n1052 & ~n1303 ) ;
  assign n1306 = n1304 & ~n1305 ;
  assign n1307 = ~n434 & n949 ;
  assign n1308 = n434 & n951 ;
  assign n1309 = n1307 | n1308 ;
  assign n1310 = ( n421 & n937 ) | ( n421 & ~n1309 ) | ( n937 & ~n1309 ) ;
  assign n1311 = ( n421 & n935 ) | ( n421 & n1309 ) | ( n935 & n1309 ) ;
  assign n1312 = n1310 & ~n1311 ;
  assign n1313 = ( ~n1300 & n1306 ) | ( ~n1300 & n1312 ) | ( n1306 & n1312 ) ;
  assign n1314 = n1297 & n1313 ;
  assign n1315 = n1297 & ~n1314 ;
  assign n1316 = ~n1297 & n1313 ;
  assign n1317 = n1315 | n1316 ;
  assign n1318 = ( n1300 & ~n1306 ) | ( n1300 & n1313 ) | ( ~n1306 & n1313 ) ;
  assign n1319 = ( ~n1312 & n1313 ) | ( ~n1312 & n1318 ) | ( n1313 & n1318 ) ;
  assign n1320 = n434 | n1055 ;
  assign n1321 = n434 & n1052 ;
  assign n1322 = ( n434 & n1053 ) | ( n434 & n1055 ) | ( n1053 & n1055 ) ;
  assign n1323 = ~n1321 & n1322 ;
  assign n1324 = n32 | n568 ;
  assign n1325 = n486 & n1324 ;
  assign n1326 = ( n486 & n568 ) | ( n486 & n822 ) | ( n568 & n822 ) ;
  assign n1327 = n496 & ~n822 ;
  assign n1328 = ( n556 & n822 ) | ( n556 & ~n1327 ) | ( n822 & ~n1327 ) ;
  assign n1329 = ( n1325 & ~n1326 ) | ( n1325 & n1328 ) | ( ~n1326 & n1328 ) ;
  assign n1330 = ~n1053 & n1329 ;
  assign n1331 = ( ~n1323 & n1329 ) | ( ~n1323 & n1330 ) | ( n1329 & n1330 ) ;
  assign n1332 = n1053 & n1323 ;
  assign n1333 = ( ~n1329 & n1330 ) | ( ~n1329 & n1332 ) | ( n1330 & n1332 ) ;
  assign n1334 = n1331 | n1333 ;
  assign n1335 = n1320 & ~n1334 ;
  assign n1336 = n421 & ~n464 ;
  assign n1337 = ( n421 & n485 ) | ( n421 & n1336 ) | ( n485 & n1336 ) ;
  assign n1338 = n434 | n568 ;
  assign n1339 = n1337 | n1338 ;
  assign n1340 = n421 | n486 ;
  assign n1341 = ( n421 & n568 ) | ( n421 & n1340 ) | ( n568 & n1340 ) ;
  assign n1342 = ~n1337 & n1341 ;
  assign n1343 = ( n32 & n486 ) | ( n32 & n568 ) | ( n486 & n568 ) ;
  assign n1344 = ( n1324 & n1342 ) | ( n1324 & ~n1343 ) | ( n1342 & ~n1343 ) ;
  assign n1345 = n1322 & ~n1332 ;
  assign n1346 = ( n1339 & n1344 ) | ( n1339 & ~n1345 ) | ( n1344 & ~n1345 ) ;
  assign n1347 = ( n1320 & n1335 ) | ( n1320 & ~n1346 ) | ( n1335 & ~n1346 ) ;
  assign n1348 = n434 & ~n1057 ;
  assign n1349 = ( n421 & n1052 ) | ( n421 & n1348 ) | ( n1052 & n1348 ) ;
  assign n1350 = ( ~n421 & n1054 ) | ( ~n421 & n1348 ) | ( n1054 & n1348 ) ;
  assign n1351 = n1349 | n1350 ;
  assign n1352 = n1347 & ~n1351 ;
  assign n1353 = n1293 & ~n1334 ;
  assign n1354 = ~n1346 & n1353 ;
  assign n1355 = ( n1293 & n1352 ) | ( n1293 & n1354 ) | ( n1352 & n1354 ) ;
  assign n1356 = ~n1319 & n1355 ;
  assign n1357 = ~n1293 & n1334 ;
  assign n1358 = ( ~n1293 & n1346 ) | ( ~n1293 & n1357 ) | ( n1346 & n1357 ) ;
  assign n1359 = ~n1352 & n1358 ;
  assign n1360 = n421 | n1055 ;
  assign n1361 = n421 & ~n1057 ;
  assign n1362 = n1360 & ~n1361 ;
  assign n1363 = ( n32 & ~n1054 ) | ( n32 & n1362 ) | ( ~n1054 & n1362 ) ;
  assign n1364 = ( n32 & n1052 ) | ( n32 & ~n1362 ) | ( n1052 & ~n1362 ) ;
  assign n1365 = n1363 & ~n1364 ;
  assign n1366 = n486 & n1328 ;
  assign n1367 = ( n486 & n568 ) | ( n486 & n756 ) | ( n568 & n756 ) ;
  assign n1368 = ( n1288 & n1366 ) | ( n1288 & ~n1367 ) | ( n1366 & ~n1367 ) ;
  assign n1369 = ( n1333 & n1365 ) | ( n1333 & ~n1368 ) | ( n1365 & ~n1368 ) ;
  assign n1370 = ( ~n1333 & n1365 ) | ( ~n1333 & n1368 ) | ( n1365 & n1368 ) ;
  assign n1371 = ( ~n1365 & n1369 ) | ( ~n1365 & n1370 ) | ( n1369 & n1370 ) ;
  assign n1372 = n1359 | n1371 ;
  assign n1373 = ( n1319 & ~n1356 ) | ( n1319 & n1372 ) | ( ~n1356 & n1372 ) ;
  assign n1374 = n1317 & ~n1373 ;
  assign n1375 = n1319 & ~n1355 ;
  assign n1376 = n1372 & n1375 ;
  assign n1377 = n1369 & ~n1376 ;
  assign n1378 = ( n1317 & n1374 ) | ( n1317 & n1377 ) | ( n1374 & n1377 ) ;
  assign n1379 = ( n1294 & n1314 ) | ( n1294 & ~n1315 ) | ( n1314 & ~n1315 ) ;
  assign n1380 = ( n1223 & n1296 ) | ( n1223 & n1379 ) | ( n1296 & n1379 ) ;
  assign n1381 = n1378 | n1380 ;
  assign n1382 = ~n1317 & n1373 ;
  assign n1383 = ~n1377 & n1382 ;
  assign n1384 = ( n1267 & ~n1273 ) | ( n1267 & n1279 ) | ( ~n1273 & n1279 ) ;
  assign n1385 = ( ~n1279 & n1280 ) | ( ~n1279 & n1384 ) | ( n1280 & n1384 ) ;
  assign n1386 = n1383 | n1385 ;
  assign n1387 = ~n1381 & n1386 ;
  assign n1388 = ( n1283 & ~n1285 ) | ( n1283 & n1387 ) | ( ~n1285 & n1387 ) ;
  assign n1389 = n1286 | n1388 ;
  assign n1390 = n1378 & n1380 ;
  assign n1391 = ( n1380 & ~n1386 ) | ( n1380 & n1390 ) | ( ~n1386 & n1390 ) ;
  assign n1392 = n1287 & n1391 ;
  assign n1393 = ( n1287 & ~n1389 ) | ( n1287 & n1392 ) | ( ~n1389 & n1392 ) ;
  assign n1394 = n1262 & n1393 ;
  assign n1395 = n1287 | n1391 ;
  assign n1396 = n1389 & ~n1395 ;
  assign n1397 = n1257 & ~n1258 ;
  assign n1398 = ( ~n1260 & n1396 ) | ( ~n1260 & n1397 ) | ( n1396 & n1397 ) ;
  assign n1399 = n1261 | n1398 ;
  assign n1400 = ( n1262 & n1394 ) | ( n1262 & ~n1399 ) | ( n1394 & ~n1399 ) ;
  assign n1401 = n1234 & n1400 ;
  assign n1402 = n1229 & n1231 ;
  assign n1403 = n1229 | n1231 ;
  assign n1404 = ~n1402 & n1403 ;
  assign n1405 = n1233 | n1404 ;
  assign n1406 = n1262 | n1393 ;
  assign n1407 = n1399 & ~n1406 ;
  assign n1408 = ( ~n1404 & n1405 ) | ( ~n1404 & n1407 ) | ( n1405 & n1407 ) ;
  assign n1409 = ( ~n1233 & n1405 ) | ( ~n1233 & n1408 ) | ( n1405 & n1408 ) ;
  assign n1410 = ( n1234 & n1401 ) | ( n1234 & ~n1409 ) | ( n1401 & ~n1409 ) ;
  assign n1411 = n1212 & n1410 ;
  assign n1412 = n1234 | n1400 ;
  assign n1413 = n1409 & ~n1412 ;
  assign n1414 = ( ~n1208 & n1210 ) | ( ~n1208 & n1413 ) | ( n1210 & n1413 ) ;
  assign n1415 = n1211 | n1414 ;
  assign n1416 = ( n1212 & n1411 ) | ( n1212 & ~n1415 ) | ( n1411 & ~n1415 ) ;
  assign n1417 = ( n1160 & n1165 ) | ( n1160 & n1171 ) | ( n1165 & n1171 ) ;
  assign n1418 = n1166 | n1171 ;
  assign n1419 = ~n1417 & n1418 ;
  assign n1420 = ~n1169 & n1419 ;
  assign n1421 = n1212 | n1410 ;
  assign n1422 = n1415 & ~n1421 ;
  assign n1423 = ( n1169 & ~n1419 ) | ( n1169 & n1422 ) | ( ~n1419 & n1422 ) ;
  assign n1424 = ( ~n1416 & n1420 ) | ( ~n1416 & n1423 ) | ( n1420 & n1423 ) ;
  assign n1425 = n1175 | n1424 ;
  assign n1426 = n566 & n951 ;
  assign n1427 = ( n566 & n936 ) | ( n566 & n937 ) | ( n936 & n937 ) ;
  assign n1428 = ~n1426 & n1427 ;
  assign n1429 = n412 & n756 ;
  assign n1430 = ( ~n379 & n410 ) | ( ~n379 & n1429 ) | ( n410 & n1429 ) ;
  assign n1431 = ( n379 & n756 ) | ( n379 & n1430 ) | ( n756 & n1430 ) ;
  assign n1432 = n1428 & ~n1431 ;
  assign n1433 = ~n1428 & n1431 ;
  assign n1434 = n1432 | n1433 ;
  assign n1435 = n757 | n985 ;
  assign n1436 = ~n760 & n985 ;
  assign n1437 = n1435 & ~n1436 ;
  assign n1438 = ( n493 & ~n747 ) | ( n493 & n1437 ) | ( ~n747 & n1437 ) ;
  assign n1439 = ( n493 & n764 ) | ( n493 & ~n1437 ) | ( n764 & ~n1437 ) ;
  assign n1440 = n1438 & ~n1439 ;
  assign n1441 = ~n1434 & n1440 ;
  assign n1442 = n1434 & ~n1440 ;
  assign n1443 = n1441 | n1442 ;
  assign n1444 = n823 | n948 ;
  assign n1445 = ~n826 & n948 ;
  assign n1446 = n1444 & ~n1445 ;
  assign n1447 = ( ~n817 & n943 ) | ( ~n817 & n1446 ) | ( n943 & n1446 ) ;
  assign n1448 = ( n830 & n943 ) | ( n830 & ~n1446 ) | ( n943 & ~n1446 ) ;
  assign n1449 = n1447 & ~n1448 ;
  assign n1450 = n418 | n756 ;
  assign n1451 = ~n423 & n756 ;
  assign n1452 = n1450 & ~n1451 ;
  assign n1453 = ( ~n427 & n752 ) | ( ~n427 & n1452 ) | ( n752 & n1452 ) ;
  assign n1454 = ( n416 & n752 ) | ( n416 & ~n1452 ) | ( n752 & ~n1452 ) ;
  assign n1455 = n1453 & ~n1454 ;
  assign n1456 = ~n493 & n949 ;
  assign n1457 = n493 & n951 ;
  assign n1458 = n1456 | n1457 ;
  assign n1459 = ( n566 & n937 ) | ( n566 & ~n1458 ) | ( n937 & ~n1458 ) ;
  assign n1460 = ( n566 & n935 ) | ( n566 & n1458 ) | ( n935 & n1458 ) ;
  assign n1461 = n1459 & ~n1460 ;
  assign n1462 = ( n1449 & n1455 ) | ( n1449 & n1461 ) | ( n1455 & n1461 ) ;
  assign n1463 = ~n1443 & n1462 ;
  assign n1464 = n1462 & ~n1463 ;
  assign n1465 = n1443 | n1463 ;
  assign n1466 = ~n1464 & n1465 ;
  assign n1467 = n418 | n752 ;
  assign n1468 = ~n423 & n752 ;
  assign n1469 = n1467 & ~n1468 ;
  assign n1470 = ( ~n427 & n948 ) | ( ~n427 & n1469 ) | ( n948 & n1469 ) ;
  assign n1471 = ( n416 & n948 ) | ( n416 & ~n1469 ) | ( n948 & ~n1469 ) ;
  assign n1472 = n1470 & ~n1471 ;
  assign n1473 = n823 | n943 ;
  assign n1474 = ~n826 & n943 ;
  assign n1475 = n1473 & ~n1474 ;
  assign n1476 = ( ~n817 & n977 ) | ( ~n817 & n1475 ) | ( n977 & n1475 ) ;
  assign n1477 = ( n830 & n977 ) | ( n830 & ~n1475 ) | ( n977 & ~n1475 ) ;
  assign n1478 = n1476 & ~n1477 ;
  assign n1479 = ~n568 & n1053 ;
  assign n1480 = ( n568 & n892 ) | ( n568 & n1479 ) | ( n892 & n1479 ) ;
  assign n1481 = n412 & n822 ;
  assign n1482 = ( ~n379 & n410 ) | ( ~n379 & n1481 ) | ( n410 & n1481 ) ;
  assign n1483 = ( n379 & n822 ) | ( n379 & n1482 ) | ( n822 & n1482 ) ;
  assign n1484 = ( ~n1479 & n1480 ) | ( ~n1479 & n1483 ) | ( n1480 & n1483 ) ;
  assign n1485 = ( n1472 & n1478 ) | ( n1472 & n1484 ) | ( n1478 & n1484 ) ;
  assign n1486 = ( n1478 & n1484 ) | ( n1478 & ~n1485 ) | ( n1484 & ~n1485 ) ;
  assign n1487 = ( n1472 & ~n1485 ) | ( n1472 & n1486 ) | ( ~n1485 & n1486 ) ;
  assign n1488 = n1466 | n1487 ;
  assign n1489 = ( n1463 & ~n1466 ) | ( n1463 & n1488 ) | ( ~n1466 & n1488 ) ;
  assign n1490 = n823 | n977 ;
  assign n1491 = ~n826 & n977 ;
  assign n1492 = n1490 & ~n1491 ;
  assign n1493 = ( ~n817 & n985 ) | ( ~n817 & n1492 ) | ( n985 & n1492 ) ;
  assign n1494 = ( n830 & n985 ) | ( n830 & ~n1492 ) | ( n985 & ~n1492 ) ;
  assign n1495 = n1493 & ~n1494 ;
  assign n1496 = n493 | n757 ;
  assign n1497 = n493 & ~n760 ;
  assign n1498 = n1496 & ~n1497 ;
  assign n1499 = ( n566 & ~n747 ) | ( n566 & n1498 ) | ( ~n747 & n1498 ) ;
  assign n1500 = ( n566 & n764 ) | ( n566 & ~n1498 ) | ( n764 & ~n1498 ) ;
  assign n1501 = n1499 & ~n1500 ;
  assign n1502 = n418 | n948 ;
  assign n1503 = ~n423 & n948 ;
  assign n1504 = n1502 & ~n1503 ;
  assign n1505 = ( ~n427 & n943 ) | ( ~n427 & n1504 ) | ( n943 & n1504 ) ;
  assign n1506 = ( n416 & n943 ) | ( n416 & ~n1504 ) | ( n943 & ~n1504 ) ;
  assign n1507 = n1505 & ~n1506 ;
  assign n1508 = ( n1495 & n1501 ) | ( n1495 & n1507 ) | ( n1501 & n1507 ) ;
  assign n1509 = ( n1501 & n1507 ) | ( n1501 & ~n1508 ) | ( n1507 & ~n1508 ) ;
  assign n1510 = ( n1495 & ~n1508 ) | ( n1495 & n1509 ) | ( ~n1508 & n1509 ) ;
  assign n1511 = n1489 & n1510 ;
  assign n1512 = n1489 | n1510 ;
  assign n1513 = ~n1511 & n1512 ;
  assign n1514 = n414 & n752 ;
  assign n1515 = ( n936 & ~n1431 ) | ( n936 & n1514 ) | ( ~n1431 & n1514 ) ;
  assign n1516 = ( ~n936 & n1431 ) | ( ~n936 & n1515 ) | ( n1431 & n1515 ) ;
  assign n1517 = ( ~n1514 & n1515 ) | ( ~n1514 & n1516 ) | ( n1515 & n1516 ) ;
  assign n1518 = n1432 | n1441 ;
  assign n1519 = ( n1485 & n1517 ) | ( n1485 & ~n1518 ) | ( n1517 & ~n1518 ) ;
  assign n1520 = ( ~n1485 & n1518 ) | ( ~n1485 & n1519 ) | ( n1518 & n1519 ) ;
  assign n1521 = ( ~n1517 & n1519 ) | ( ~n1517 & n1520 ) | ( n1519 & n1520 ) ;
  assign n1522 = n1513 & n1521 ;
  assign n1523 = n1513 | n1521 ;
  assign n1524 = ~n1522 & n1523 ;
  assign n1525 = n1479 | n1484 ;
  assign n1526 = ( n1479 & n1480 ) | ( n1479 & n1483 ) | ( n1480 & n1483 ) ;
  assign n1527 = n1525 & ~n1526 ;
  assign n1528 = n757 | n977 ;
  assign n1529 = ~n760 & n977 ;
  assign n1530 = n1528 & ~n1529 ;
  assign n1531 = ( ~n747 & n985 ) | ( ~n747 & n1530 ) | ( n985 & n1530 ) ;
  assign n1532 = ( n764 & n985 ) | ( n764 & ~n1530 ) | ( n985 & ~n1530 ) ;
  assign n1533 = n1531 & ~n1532 ;
  assign n1534 = ~n1527 & n1533 ;
  assign n1535 = n1527 & ~n1533 ;
  assign n1536 = n1534 | n1535 ;
  assign n1537 = n32 & n379 ;
  assign n1538 = ( n32 & n413 ) | ( n32 & n1537 ) | ( n413 & n1537 ) ;
  assign n1539 = ~n568 & n1538 ;
  assign n1540 = n568 & ~n1538 ;
  assign n1541 = n1539 | n1540 ;
  assign n1542 = n566 & ~n1057 ;
  assign n1543 = ( n566 & n1053 ) | ( n566 & ~n1054 ) | ( n1053 & ~n1054 ) ;
  assign n1544 = ~n1542 & n1543 ;
  assign n1545 = ~n1541 & n1544 ;
  assign n1546 = n1539 | n1545 ;
  assign n1547 = ~n1536 & n1546 ;
  assign n1548 = n1534 | n1547 ;
  assign n1549 = n949 & ~n985 ;
  assign n1550 = n951 & n985 ;
  assign n1551 = n1549 | n1550 ;
  assign n1552 = ( n493 & n937 ) | ( n493 & ~n1551 ) | ( n937 & ~n1551 ) ;
  assign n1553 = ( n493 & n935 ) | ( n493 & n1551 ) | ( n935 & n1551 ) ;
  assign n1554 = n1552 & ~n1553 ;
  assign n1555 = n757 | n943 ;
  assign n1556 = ~n760 & n943 ;
  assign n1557 = n1555 & ~n1556 ;
  assign n1558 = ( ~n747 & n977 ) | ( ~n747 & n1557 ) | ( n977 & n1557 ) ;
  assign n1559 = ( n764 & n977 ) | ( n764 & ~n1557 ) | ( n977 & ~n1557 ) ;
  assign n1560 = n1558 & ~n1559 ;
  assign n1561 = n752 | n823 ;
  assign n1562 = n752 & ~n826 ;
  assign n1563 = n1561 & ~n1562 ;
  assign n1564 = ( ~n817 & n948 ) | ( ~n817 & n1563 ) | ( n948 & n1563 ) ;
  assign n1565 = ( n830 & n948 ) | ( n830 & ~n1563 ) | ( n948 & ~n1563 ) ;
  assign n1566 = n1564 & ~n1565 ;
  assign n1567 = ( n1554 & n1560 ) | ( n1554 & n1566 ) | ( n1560 & n1566 ) ;
  assign n1568 = ( n1449 & n1461 ) | ( n1449 & ~n1462 ) | ( n1461 & ~n1462 ) ;
  assign n1569 = ( n1455 & ~n1462 ) | ( n1455 & n1568 ) | ( ~n1462 & n1568 ) ;
  assign n1570 = n1567 & n1569 ;
  assign n1571 = n1567 | n1569 ;
  assign n1572 = ~n1570 & n1571 ;
  assign n1573 = n418 | n822 ;
  assign n1574 = ~n423 & n822 ;
  assign n1575 = n1573 & ~n1574 ;
  assign n1576 = ( ~n427 & n756 ) | ( ~n427 & n1575 ) | ( n756 & n1575 ) ;
  assign n1577 = ( n416 & n756 ) | ( n416 & ~n1575 ) | ( n756 & ~n1575 ) ;
  assign n1578 = n1576 & ~n1577 ;
  assign n1579 = n412 & n421 ;
  assign n1580 = ( ~n379 & n410 ) | ( ~n379 & n1579 ) | ( n410 & n1579 ) ;
  assign n1581 = ( n379 & n421 ) | ( n379 & n1580 ) | ( n421 & n1580 ) ;
  assign n1582 = ~n568 & n1581 ;
  assign n1583 = n568 & ~n1581 ;
  assign n1584 = n493 | n1055 ;
  assign n1585 = n493 & ~n1057 ;
  assign n1586 = n1584 & ~n1585 ;
  assign n1587 = ( n566 & ~n1054 ) | ( n566 & n1586 ) | ( ~n1054 & n1586 ) ;
  assign n1588 = ( n566 & n1052 ) | ( n566 & ~n1586 ) | ( n1052 & ~n1586 ) ;
  assign n1589 = n1587 & ~n1588 ;
  assign n1590 = ( n1582 & ~n1583 ) | ( n1582 & n1589 ) | ( ~n1583 & n1589 ) ;
  assign n1591 = n1578 & n1590 ;
  assign n1592 = n1578 | n1590 ;
  assign n1593 = ~n1591 & n1592 ;
  assign n1594 = n757 | n948 ;
  assign n1595 = ~n760 & n948 ;
  assign n1596 = n1594 & ~n1595 ;
  assign n1597 = ( ~n747 & n943 ) | ( ~n747 & n1596 ) | ( n943 & n1596 ) ;
  assign n1598 = ( n764 & n943 ) | ( n764 & ~n1596 ) | ( n943 & ~n1596 ) ;
  assign n1599 = n1597 & ~n1598 ;
  assign n1600 = n949 & ~n977 ;
  assign n1601 = n951 & n977 ;
  assign n1602 = n1600 | n1601 ;
  assign n1603 = ( n937 & n985 ) | ( n937 & ~n1602 ) | ( n985 & ~n1602 ) ;
  assign n1604 = ( n935 & n985 ) | ( n935 & n1602 ) | ( n985 & n1602 ) ;
  assign n1605 = n1603 & ~n1604 ;
  assign n1606 = n756 | n823 ;
  assign n1607 = n756 & ~n826 ;
  assign n1608 = n1606 & ~n1607 ;
  assign n1609 = ( n752 & ~n817 ) | ( n752 & n1608 ) | ( ~n817 & n1608 ) ;
  assign n1610 = ( n752 & n830 ) | ( n752 & ~n1608 ) | ( n830 & ~n1608 ) ;
  assign n1611 = n1609 & ~n1610 ;
  assign n1612 = ( n1599 & n1605 ) | ( n1599 & n1611 ) | ( n1605 & n1611 ) ;
  assign n1613 = n1593 & n1612 ;
  assign n1614 = n1591 | n1613 ;
  assign n1615 = n1572 & n1614 ;
  assign n1616 = n1570 | n1615 ;
  assign n1617 = n1466 & n1487 ;
  assign n1618 = n1488 & ~n1617 ;
  assign n1619 = ( n1548 & n1616 ) | ( n1548 & ~n1618 ) | ( n1616 & ~n1618 ) ;
  assign n1620 = ~n1524 & n1619 ;
  assign n1621 = n1524 & ~n1619 ;
  assign n1622 = n1620 | n1621 ;
  assign n1623 = n1548 & ~n1616 ;
  assign n1624 = ~n1548 & n1616 ;
  assign n1625 = n1623 | n1624 ;
  assign n1626 = n1536 & ~n1546 ;
  assign n1627 = n1547 | n1626 ;
  assign n1628 = n1541 | n1545 ;
  assign n1629 = ( ~n1544 & n1545 ) | ( ~n1544 & n1628 ) | ( n1545 & n1628 ) ;
  assign n1630 = ( n1554 & n1566 ) | ( n1554 & ~n1567 ) | ( n1566 & ~n1567 ) ;
  assign n1631 = ( n1560 & ~n1567 ) | ( n1560 & n1630 ) | ( ~n1567 & n1630 ) ;
  assign n1632 = ~n1629 & n1631 ;
  assign n1633 = n32 | n418 ;
  assign n1634 = n32 & ~n423 ;
  assign n1635 = n1633 & ~n1634 ;
  assign n1636 = ( ~n427 & n822 ) | ( ~n427 & n1635 ) | ( n822 & n1635 ) ;
  assign n1637 = ( n416 & n822 ) | ( n416 & ~n1635 ) | ( n822 & ~n1635 ) ;
  assign n1638 = n1636 & ~n1637 ;
  assign n1639 = ( n1103 & n1113 ) | ( n1103 & n1638 ) | ( n1113 & n1638 ) ;
  assign n1640 = ( n1103 & ~n1105 ) | ( n1103 & n1112 ) | ( ~n1105 & n1112 ) ;
  assign n1641 = n1638 | n1640 ;
  assign n1642 = ~n1639 & n1641 ;
  assign n1643 = n1094 & n1642 ;
  assign n1644 = n1639 | n1643 ;
  assign n1645 = n1629 & ~n1631 ;
  assign n1646 = n1632 | n1645 ;
  assign n1647 = n1644 & ~n1646 ;
  assign n1648 = ( ~n1627 & n1632 ) | ( ~n1627 & n1647 ) | ( n1632 & n1647 ) ;
  assign n1649 = n1627 & ~n1632 ;
  assign n1650 = ~n1647 & n1649 ;
  assign n1651 = n1648 | n1650 ;
  assign n1652 = n1572 | n1614 ;
  assign n1653 = ~n1615 & n1652 ;
  assign n1654 = ~n1651 & n1653 ;
  assign n1655 = n1648 | n1654 ;
  assign n1656 = ( ~n1618 & n1625 ) | ( ~n1618 & n1655 ) | ( n1625 & n1655 ) ;
  assign n1657 = ( n1618 & ~n1625 ) | ( n1618 & n1656 ) | ( ~n1625 & n1656 ) ;
  assign n1658 = n1656 & n1657 ;
  assign n1659 = ~n1622 & n1658 ;
  assign n1660 = ( ~n1655 & n1656 ) | ( ~n1655 & n1657 ) | ( n1656 & n1657 ) ;
  assign n1661 = n1593 | n1612 ;
  assign n1662 = ~n1613 & n1661 ;
  assign n1663 = ( n568 & ~n1581 ) | ( n568 & n1589 ) | ( ~n1581 & n1589 ) ;
  assign n1664 = ( ~n1589 & n1590 ) | ( ~n1589 & n1663 ) | ( n1590 & n1663 ) ;
  assign n1665 = ( n1599 & n1611 ) | ( n1599 & ~n1612 ) | ( n1611 & ~n1612 ) ;
  assign n1666 = ( n1605 & ~n1612 ) | ( n1605 & n1665 ) | ( ~n1612 & n1665 ) ;
  assign n1667 = n574 | n958 ;
  assign n1668 = ( n1664 & ~n1666 ) | ( n1664 & n1667 ) | ( ~n1666 & n1667 ) ;
  assign n1669 = ( ~n1664 & n1666 ) | ( ~n1664 & n1668 ) | ( n1666 & n1668 ) ;
  assign n1670 = n1662 & n1669 ;
  assign n1671 = n1644 & n1646 ;
  assign n1672 = n1644 | n1646 ;
  assign n1673 = ~n1671 & n1672 ;
  assign n1674 = n1662 | n1669 ;
  assign n1675 = ~n1670 & n1674 ;
  assign n1676 = ~n1673 & n1675 ;
  assign n1677 = n1670 | n1676 ;
  assign n1678 = n1651 & ~n1653 ;
  assign n1679 = n1654 | n1678 ;
  assign n1680 = n1677 & ~n1679 ;
  assign n1681 = ~n1660 & n1680 ;
  assign n1682 = ~n1677 & n1679 ;
  assign n1683 = n1660 | n1682 ;
  assign n1684 = n1094 | n1642 ;
  assign n1685 = ~n1643 & n1684 ;
  assign n1686 = ( n1131 & n1134 ) | ( n1131 & n1685 ) | ( n1134 & n1685 ) ;
  assign n1687 = ( ~n1132 & n1135 ) | ( ~n1132 & n1685 ) | ( n1135 & n1685 ) ;
  assign n1688 = ~n1686 & n1687 ;
  assign n1689 = ( ~n1667 & n1668 ) | ( ~n1667 & n1669 ) | ( n1668 & n1669 ) ;
  assign n1690 = n1688 & ~n1689 ;
  assign n1691 = n1686 | n1690 ;
  assign n1692 = n1673 & ~n1675 ;
  assign n1693 = n1676 | n1692 ;
  assign n1694 = ~n1688 & n1689 ;
  assign n1695 = n1690 | n1694 ;
  assign n1696 = n1073 | n1137 ;
  assign n1697 = ~n1695 & n1696 ;
  assign n1698 = n1695 & ~n1696 ;
  assign n1699 = n1697 | n1698 ;
  assign n1700 = n1173 & ~n1699 ;
  assign n1701 = n1697 | n1700 ;
  assign n1702 = ( n1691 & ~n1693 ) | ( n1691 & n1701 ) | ( ~n1693 & n1701 ) ;
  assign n1703 = ( n1681 & ~n1683 ) | ( n1681 & n1702 ) | ( ~n1683 & n1702 ) ;
  assign n1704 = ( ~n1622 & n1659 ) | ( ~n1622 & n1703 ) | ( n1659 & n1703 ) ;
  assign n1705 = n493 | n823 ;
  assign n1706 = n493 & ~n826 ;
  assign n1707 = n1705 & ~n1706 ;
  assign n1708 = ( n566 & ~n817 ) | ( n566 & n1707 ) | ( ~n817 & n1707 ) ;
  assign n1709 = ( n566 & n830 ) | ( n566 & ~n1707 ) | ( n830 & ~n1707 ) ;
  assign n1710 = n1708 & ~n1709 ;
  assign n1711 = n418 | n977 ;
  assign n1712 = ~n423 & n977 ;
  assign n1713 = n1711 & ~n1712 ;
  assign n1714 = ( ~n427 & n985 ) | ( ~n427 & n1713 ) | ( n985 & n1713 ) ;
  assign n1715 = ( n416 & n985 ) | ( n416 & ~n1713 ) | ( n985 & ~n1713 ) ;
  assign n1716 = n1714 & ~n1715 ;
  assign n1717 = n1710 & n1716 ;
  assign n1718 = n1710 | n1716 ;
  assign n1719 = ~n1717 & n1718 ;
  assign n1720 = n412 & n948 ;
  assign n1721 = ( ~n379 & n410 ) | ( ~n379 & n1720 ) | ( n410 & n1720 ) ;
  assign n1722 = ( n379 & n948 ) | ( n379 & n1721 ) | ( n948 & n1721 ) ;
  assign n1723 = ( n566 & n747 ) | ( n566 & ~n760 ) | ( n747 & ~n760 ) ;
  assign n1724 = ( n566 & n746 ) | ( n566 & ~n747 ) | ( n746 & ~n747 ) ;
  assign n1725 = ~n1723 & n1724 ;
  assign n1726 = ~n1722 & n1725 ;
  assign n1727 = n1722 & ~n1725 ;
  assign n1728 = n1726 | n1727 ;
  assign n1729 = n823 | n985 ;
  assign n1730 = ~n826 & n985 ;
  assign n1731 = n1729 & ~n1730 ;
  assign n1732 = ( n493 & ~n817 ) | ( n493 & n1731 ) | ( ~n817 & n1731 ) ;
  assign n1733 = ( n493 & n830 ) | ( n493 & ~n1731 ) | ( n830 & ~n1731 ) ;
  assign n1734 = n1732 & ~n1733 ;
  assign n1735 = ~n1728 & n1734 ;
  assign n1736 = n1726 | n1735 ;
  assign n1737 = n1719 & n1736 ;
  assign n1738 = ~n746 & n1722 ;
  assign n1739 = ( n746 & ~n1722 ) | ( n746 & n1738 ) | ( ~n1722 & n1738 ) ;
  assign n1740 = n1738 | n1739 ;
  assign n1741 = n379 & n943 ;
  assign n1742 = ( n413 & n943 ) | ( n413 & n1741 ) | ( n943 & n1741 ) ;
  assign n1743 = ~n1740 & n1742 ;
  assign n1744 = n1738 | n1743 ;
  assign n1745 = n1716 & n1744 ;
  assign n1746 = n1710 & n1745 ;
  assign n1747 = ( n1737 & n1744 ) | ( n1737 & n1746 ) | ( n1744 & n1746 ) ;
  assign n1748 = ( n566 & n817 ) | ( n566 & ~n826 ) | ( n817 & ~n826 ) ;
  assign n1749 = ( n566 & n813 ) | ( n566 & ~n817 ) | ( n813 & ~n817 ) ;
  assign n1750 = ~n1748 & n1749 ;
  assign n1751 = n379 & n977 ;
  assign n1752 = ( n413 & n977 ) | ( n413 & n1751 ) | ( n977 & n1751 ) ;
  assign n1753 = n1750 & ~n1752 ;
  assign n1754 = ~n1750 & n1752 ;
  assign n1755 = n1753 | n1754 ;
  assign n1756 = n418 | n985 ;
  assign n1757 = ~n423 & n985 ;
  assign n1758 = n1756 & ~n1757 ;
  assign n1759 = ( ~n427 & n493 ) | ( ~n427 & n1758 ) | ( n493 & n1758 ) ;
  assign n1760 = ( n416 & n493 ) | ( n416 & ~n1758 ) | ( n493 & ~n1758 ) ;
  assign n1761 = n1759 & ~n1760 ;
  assign n1762 = ~n1755 & n1761 ;
  assign n1763 = n1755 & ~n1761 ;
  assign n1764 = n1762 | n1763 ;
  assign n1765 = n1744 & ~n1746 ;
  assign n1766 = ~n1737 & n1765 ;
  assign n1767 = ( n1717 & n1737 ) | ( n1717 & ~n1747 ) | ( n1737 & ~n1747 ) ;
  assign n1768 = n1766 | n1767 ;
  assign n1769 = ~n1764 & n1768 ;
  assign n1770 = n1747 | n1769 ;
  assign n1771 = n418 | n493 ;
  assign n1772 = ~n423 & n493 ;
  assign n1773 = n1771 & ~n1772 ;
  assign n1774 = ( ~n427 & n566 ) | ( ~n427 & n1773 ) | ( n566 & n1773 ) ;
  assign n1775 = ( n416 & n566 ) | ( n416 & ~n1773 ) | ( n566 & ~n1773 ) ;
  assign n1776 = n1774 & ~n1775 ;
  assign n1777 = n1753 | n1762 ;
  assign n1778 = n1776 & n1777 ;
  assign n1779 = n1776 | n1777 ;
  assign n1780 = ~n1778 & n1779 ;
  assign n1781 = n379 & n985 ;
  assign n1782 = ( n413 & n985 ) | ( n413 & n1781 ) | ( n985 & n1781 ) ;
  assign n1783 = ( n813 & n1752 ) | ( n813 & n1782 ) | ( n1752 & n1782 ) ;
  assign n1784 = ( n813 & n1782 ) | ( n813 & ~n1783 ) | ( n1782 & ~n1783 ) ;
  assign n1785 = ( n1752 & ~n1783 ) | ( n1752 & n1784 ) | ( ~n1783 & n1784 ) ;
  assign n1786 = n1780 & ~n1785 ;
  assign n1787 = ~n1780 & n1785 ;
  assign n1788 = n1786 | n1787 ;
  assign n1789 = n1770 & ~n1788 ;
  assign n1790 = ~n1770 & n1788 ;
  assign n1791 = n1789 | n1790 ;
  assign n1792 = n1764 & ~n1768 ;
  assign n1793 = n1769 | n1792 ;
  assign n1794 = n1740 & ~n1742 ;
  assign n1795 = n1743 | n1794 ;
  assign n1796 = n418 | n943 ;
  assign n1797 = ~n423 & n943 ;
  assign n1798 = n1796 & ~n1797 ;
  assign n1799 = ( ~n427 & n977 ) | ( ~n427 & n1798 ) | ( n977 & n1798 ) ;
  assign n1800 = ( n416 & n977 ) | ( n416 & ~n1798 ) | ( n977 & ~n1798 ) ;
  assign n1801 = n1799 & ~n1800 ;
  assign n1802 = ( n1508 & n1516 ) | ( n1508 & n1801 ) | ( n1516 & n1801 ) ;
  assign n1803 = ~n1795 & n1802 ;
  assign n1804 = n1795 & ~n1802 ;
  assign n1805 = n1803 | n1804 ;
  assign n1806 = n1719 | n1736 ;
  assign n1807 = ~n1737 & n1806 ;
  assign n1808 = ~n1805 & n1807 ;
  assign n1809 = n1803 | n1808 ;
  assign n1810 = n1805 & ~n1807 ;
  assign n1811 = n1808 | n1810 ;
  assign n1812 = n1485 & n1518 ;
  assign n1813 = n1728 & ~n1734 ;
  assign n1814 = n1735 | n1813 ;
  assign n1815 = ( n1485 & ~n1517 ) | ( n1485 & n1518 ) | ( ~n1517 & n1518 ) ;
  assign n1816 = ~n1812 & n1815 ;
  assign n1817 = ( n1812 & ~n1814 ) | ( n1812 & n1816 ) | ( ~n1814 & n1816 ) ;
  assign n1818 = ( n1508 & ~n1516 ) | ( n1508 & n1801 ) | ( ~n1516 & n1801 ) ;
  assign n1819 = ( n1516 & ~n1801 ) | ( n1516 & n1818 ) | ( ~n1801 & n1818 ) ;
  assign n1820 = ( ~n1508 & n1818 ) | ( ~n1508 & n1819 ) | ( n1818 & n1819 ) ;
  assign n1821 = ~n1812 & n1814 ;
  assign n1822 = ~n1816 & n1821 ;
  assign n1823 = n1817 | n1822 ;
  assign n1824 = n1820 | n1823 ;
  assign n1825 = ~n1820 & n1824 ;
  assign n1826 = ( ~n1823 & n1824 ) | ( ~n1823 & n1825 ) | ( n1824 & n1825 ) ;
  assign n1827 = ( n1817 & n1820 ) | ( n1817 & n1826 ) | ( n1820 & n1826 ) ;
  assign n1828 = ~n1811 & n1827 ;
  assign n1829 = ( n1511 & n1513 ) | ( n1511 & ~n1522 ) | ( n1513 & ~n1522 ) ;
  assign n1830 = ~n1826 & n1829 ;
  assign n1831 = n1826 | n1830 ;
  assign n1832 = n1826 & n1829 ;
  assign n1833 = n1831 & ~n1832 ;
  assign n1834 = n1620 & ~n1833 ;
  assign n1835 = n1811 & ~n1827 ;
  assign n1836 = n1828 | n1835 ;
  assign n1837 = ( n1830 & n1834 ) | ( n1830 & ~n1836 ) | ( n1834 & ~n1836 ) ;
  assign n1838 = n1828 | n1837 ;
  assign n1839 = ( ~n1793 & n1809 ) | ( ~n1793 & n1838 ) | ( n1809 & n1838 ) ;
  assign n1840 = ~n1791 & n1839 ;
  assign n1841 = n1789 | n1840 ;
  assign n1842 = n1793 & n1809 ;
  assign n1843 = n1793 | n1809 ;
  assign n1844 = ~n1842 & n1843 ;
  assign n1845 = n1835 | n1844 ;
  assign n1846 = ~n1830 & n1833 ;
  assign n1847 = n1836 & n1846 ;
  assign n1848 = ( n1845 & n1846 ) | ( n1845 & ~n1847 ) | ( n1846 & ~n1847 ) ;
  assign n1849 = ~n1793 & n1809 ;
  assign n1850 = n1848 & ~n1849 ;
  assign n1851 = n1791 | n1850 ;
  assign n1852 = ~n1789 & n1851 ;
  assign n1853 = ( n1704 & n1841 ) | ( n1704 & ~n1852 ) | ( n1841 & ~n1852 ) ;
  assign n1854 = n1680 | n1682 ;
  assign n1855 = n1691 & ~n1693 ;
  assign n1856 = ~n1691 & n1693 ;
  assign n1857 = n1855 | n1856 ;
  assign n1858 = n1698 | n1857 ;
  assign n1859 = ( n1854 & ~n1855 ) | ( n1854 & n1858 ) | ( ~n1855 & n1858 ) ;
  assign n1860 = ( n1660 & ~n1681 ) | ( n1660 & n1859 ) | ( ~n1681 & n1859 ) ;
  assign n1861 = ( n1622 & ~n1659 ) | ( n1622 & n1860 ) | ( ~n1659 & n1860 ) ;
  assign n1862 = ( ~n1841 & n1852 ) | ( ~n1841 & n1861 ) | ( n1852 & n1861 ) ;
  assign n1863 = ( n1425 & ~n1853 ) | ( n1425 & n1862 ) | ( ~n1853 & n1862 ) ;
  assign n1864 = ( n1776 & n1777 ) | ( n1776 & n1786 ) | ( n1777 & n1786 ) ;
  assign n1865 = ( ~n423 & n427 ) | ( ~n423 & n566 ) | ( n427 & n566 ) ;
  assign n1866 = ( n417 & ~n427 ) | ( n417 & n566 ) | ( ~n427 & n566 ) ;
  assign n1867 = ~n1865 & n1866 ;
  assign n1868 = n379 & n493 ;
  assign n1869 = ( n413 & n493 ) | ( n413 & n1868 ) | ( n493 & n1868 ) ;
  assign n1870 = ~n1867 & n1869 ;
  assign n1871 = ( ~n813 & n1752 ) | ( ~n813 & n1782 ) | ( n1752 & n1782 ) ;
  assign n1872 = ( n1867 & ~n1869 ) | ( n1867 & n1871 ) | ( ~n1869 & n1871 ) ;
  assign n1873 = n1870 | n1872 ;
  assign n1874 = n1867 & ~n1869 ;
  assign n1875 = ( n1870 & n1871 ) | ( n1870 & n1874 ) | ( n1871 & n1874 ) ;
  assign n1876 = n1873 & ~n1875 ;
  assign n1877 = ~n1864 & n1876 ;
  assign n1878 = n1876 & ~n1877 ;
  assign n1879 = ( n1864 & n1877 ) | ( n1864 & ~n1878 ) | ( n1877 & ~n1878 ) ;
  assign n1880 = n1863 & ~n1879 ;
  assign n1881 = n1879 | n1880 ;
  assign n1882 = ( ~n1863 & n1880 ) | ( ~n1863 & n1881 ) | ( n1880 & n1881 ) ;
  assign n1883 = n264 & ~n1882 ;
  assign n1884 = ( ~n1840 & n1851 ) | ( ~n1840 & n1861 ) | ( n1851 & n1861 ) ;
  assign n1885 = ( n1704 & n1840 ) | ( n1704 & ~n1851 ) | ( n1840 & ~n1851 ) ;
  assign n1886 = ( n1425 & n1884 ) | ( n1425 & ~n1885 ) | ( n1884 & ~n1885 ) ;
  assign n1887 = n1791 & n1850 ;
  assign n1888 = n1791 & ~n1839 ;
  assign n1889 = ( n1861 & n1887 ) | ( n1861 & n1888 ) | ( n1887 & n1888 ) ;
  assign n1890 = ( ~n1704 & n1887 ) | ( ~n1704 & n1888 ) | ( n1887 & n1888 ) ;
  assign n1891 = ( n1425 & n1889 ) | ( n1425 & n1890 ) | ( n1889 & n1890 ) ;
  assign n1892 = n1886 & ~n1891 ;
  assign n1893 = n658 | n695 ;
  assign n1894 = n320 | n864 ;
  assign n1895 = n1893 | n1894 ;
  assign n1896 = n609 | n797 ;
  assign n1897 = n1895 | n1896 ;
  assign n1898 = n773 | n925 ;
  assign n1899 = n1897 | n1898 ;
  assign n1900 = n157 | n179 ;
  assign n1901 = n201 | n239 ;
  assign n1902 = n1900 | n1901 ;
  assign n1903 = n577 | n1902 ;
  assign n1904 = n554 | n1903 ;
  assign n1905 = n1899 | n1904 ;
  assign n1906 = n1892 & ~n1905 ;
  assign n1907 = ~n264 & n1882 ;
  assign n1908 = ( ~n1883 & n1906 ) | ( ~n1883 & n1907 ) | ( n1906 & n1907 ) ;
  assign n1909 = n1864 & ~n1876 ;
  assign n1910 = ~n1872 & n1909 ;
  assign n1911 = ( n1872 & n1879 ) | ( n1872 & ~n1910 ) | ( n1879 & ~n1910 ) ;
  assign n1912 = ( n1853 & n1910 ) | ( n1853 & ~n1911 ) | ( n1910 & ~n1911 ) ;
  assign n1913 = ( n1862 & ~n1910 ) | ( n1862 & n1911 ) | ( ~n1910 & n1911 ) ;
  assign n1914 = ( n1425 & ~n1912 ) | ( n1425 & n1913 ) | ( ~n1912 & n1913 ) ;
  assign n1915 = n1872 & ~n1909 ;
  assign n1916 = n1879 & n1915 ;
  assign n1917 = ( ~n1853 & n1915 ) | ( ~n1853 & n1916 ) | ( n1915 & n1916 ) ;
  assign n1918 = ( n1862 & n1915 ) | ( n1862 & n1916 ) | ( n1915 & n1916 ) ;
  assign n1919 = ( n1425 & n1917 ) | ( n1425 & n1918 ) | ( n1917 & n1918 ) ;
  assign n1920 = n1914 & ~n1919 ;
  assign n1921 = ~n493 & n566 ;
  assign n1922 = n493 & ~n566 ;
  assign n1923 = n1921 | n1922 ;
  assign n1924 = n317 & n342 ;
  assign n1925 = n1923 & ~n1924 ;
  assign n1926 = ( n414 & n1923 ) | ( n414 & ~n1924 ) | ( n1923 & ~n1924 ) ;
  assign n1927 = ~n1925 & n1926 ;
  assign n1928 = n1920 & n1927 ;
  assign n1929 = n1920 | n1927 ;
  assign n1930 = ~n1928 & n1929 ;
  assign n1931 = n338 | n363 ;
  assign n1932 = n248 | n273 ;
  assign n1933 = n1931 | n1932 ;
  assign n1934 = n459 | n1933 ;
  assign n1935 = n1024 | n1934 ;
  assign n1936 = n381 | n742 ;
  assign n1937 = n1935 | n1936 ;
  assign n1938 = n112 | n284 ;
  assign n1939 = n176 | n1938 ;
  assign n1940 = n390 | n693 ;
  assign n1941 = n1939 | n1940 ;
  assign n1942 = n276 | n1941 ;
  assign n1943 = n1937 | n1942 ;
  assign n1944 = n359 | n380 ;
  assign n1945 = n211 | n400 ;
  assign n1946 = n1944 | n1945 ;
  assign n1947 = n132 | n1946 ;
  assign n1948 = n108 | n481 ;
  assign n1949 = n209 | n519 ;
  assign n1950 = n1948 | n1949 ;
  assign n1951 = n778 | n1950 ;
  assign n1952 = n1947 | n1951 ;
  assign n1953 = n236 | n250 ;
  assign n1954 = n204 | n367 ;
  assign n1955 = n1953 | n1954 ;
  assign n1956 = n201 | n238 ;
  assign n1957 = n1955 | n1956 ;
  assign n1958 = n498 & ~n1957 ;
  assign n1959 = ~n1952 & n1958 ;
  assign n1960 = ~n1943 & n1959 ;
  assign n1961 = n534 | n869 ;
  assign n1962 = n155 | n1961 ;
  assign n1963 = n253 | n1962 ;
  assign n1964 = n1960 & ~n1963 ;
  assign n1965 = n1930 | n1964 ;
  assign n1966 = n101 | n471 ;
  assign n1967 = n176 | n1966 ;
  assign n1968 = n359 | n397 ;
  assign n1969 = n381 | n1968 ;
  assign n1970 = n349 | n660 ;
  assign n1971 = n1969 | n1970 ;
  assign n1972 = n338 | n1971 ;
  assign n1973 = n524 | n847 ;
  assign n1974 = n579 | n1973 ;
  assign n1975 = n173 | n705 ;
  assign n1976 = n238 | n336 ;
  assign n1977 = n1975 | n1976 ;
  assign n1978 = n1974 | n1977 ;
  assign n1979 = n136 | n322 ;
  assign n1980 = n1978 | n1979 ;
  assign n1981 = n1972 | n1980 ;
  assign n1982 = n447 | n458 ;
  assign n1983 = n443 | n1982 ;
  assign n1984 = n548 | n788 ;
  assign n1985 = n786 | n1984 ;
  assign n1986 = n180 | n836 ;
  assign n1987 = n1985 | n1986 ;
  assign n1988 = n1983 | n1987 ;
  assign n1989 = n1981 | n1988 ;
  assign n1990 = n1967 | n1989 ;
  assign n1991 = n1965 & ~n1990 ;
  assign n1992 = n1930 & n1964 ;
  assign n1993 = n1965 & ~n1992 ;
  assign n1994 = n1991 & ~n1993 ;
  assign n1995 = ( n1908 & n1991 ) | ( n1908 & n1994 ) | ( n1991 & n1994 ) ;
  assign n1996 = n1838 & ~n1844 ;
  assign n1997 = ( n1848 & n1861 ) | ( n1848 & ~n1996 ) | ( n1861 & ~n1996 ) ;
  assign n1998 = ( n1704 & ~n1848 ) | ( n1704 & n1996 ) | ( ~n1848 & n1996 ) ;
  assign n1999 = ( n1425 & n1997 ) | ( n1425 & ~n1998 ) | ( n1997 & ~n1998 ) ;
  assign n2000 = ~n1838 & n1844 ;
  assign n2001 = ( ~n1828 & n1835 ) | ( ~n1828 & n1846 ) | ( n1835 & n1846 ) ;
  assign n2002 = n1844 & n2001 ;
  assign n2003 = ( n1861 & n2000 ) | ( n1861 & n2002 ) | ( n2000 & n2002 ) ;
  assign n2004 = ( ~n1704 & n2000 ) | ( ~n1704 & n2002 ) | ( n2000 & n2002 ) ;
  assign n2005 = ( n1425 & n2003 ) | ( n1425 & n2004 ) | ( n2003 & n2004 ) ;
  assign n2006 = n1999 & ~n2005 ;
  assign n2007 = n708 | n777 ;
  assign n2008 = n197 | n235 ;
  assign n2009 = n870 | n2008 ;
  assign n2010 = n186 | n291 ;
  assign n2011 = n97 | n2010 ;
  assign n2012 = n2009 | n2011 ;
  assign n2013 = n397 | n2012 ;
  assign n2014 = n2007 | n2013 ;
  assign n2015 = n356 | n369 ;
  assign n2016 = n218 | n2015 ;
  assign n2017 = n2014 | n2016 ;
  assign n2018 = n192 | n296 ;
  assign n2019 = n597 | n2018 ;
  assign n2020 = n322 | n2019 ;
  assign n2021 = n143 | n293 ;
  assign n2022 = n200 | n2021 ;
  assign n2023 = n693 | n2022 ;
  assign n2024 = n2020 | n2023 ;
  assign n2025 = n444 | n692 ;
  assign n2026 = n2024 | n2025 ;
  assign n2027 = n2017 | n2026 ;
  assign n2028 = n101 | n211 ;
  assign n2029 = n367 | n1953 ;
  assign n2030 = n122 | n2029 ;
  assign n2031 = n527 | n721 ;
  assign n2032 = n797 | n2031 ;
  assign n2033 = n2030 | n2032 ;
  assign n2034 = n249 | n254 ;
  assign n2035 = n742 | n2034 ;
  assign n2036 = n2033 | n2035 ;
  assign n2037 = n384 | n544 ;
  assign n2038 = n227 | n362 ;
  assign n2039 = n2037 | n2038 ;
  assign n2040 = n411 | n2039 ;
  assign n2041 = n2036 | n2040 ;
  assign n2042 = n2028 | n2041 ;
  assign n2043 = n2027 | n2042 ;
  assign n2044 = ~n2006 & n2043 ;
  assign n2045 = ( ~n1892 & n1905 ) | ( ~n1892 & n2044 ) | ( n1905 & n2044 ) ;
  assign n2046 = ( n1883 & ~n1907 ) | ( n1883 & n2045 ) | ( ~n1907 & n2045 ) ;
  assign n2047 = ( n1991 & n1994 ) | ( n1991 & ~n2046 ) | ( n1994 & ~n2046 ) ;
  assign n2048 = n2006 & ~n2043 ;
  assign n2049 = n2044 | n2048 ;
  assign n2050 = n1836 | n1846 ;
  assign n2051 = ( ~n1837 & n1861 ) | ( ~n1837 & n2050 ) | ( n1861 & n2050 ) ;
  assign n2052 = ( n1704 & n1837 ) | ( n1704 & ~n2050 ) | ( n1837 & ~n2050 ) ;
  assign n2053 = ( n1425 & n2051 ) | ( n1425 & ~n2052 ) | ( n2051 & ~n2052 ) ;
  assign n2054 = ~n1830 & n1836 ;
  assign n2055 = ~n1834 & n2054 ;
  assign n2056 = ( n1847 & n1861 ) | ( n1847 & n2055 ) | ( n1861 & n2055 ) ;
  assign n2057 = ( ~n1704 & n1847 ) | ( ~n1704 & n2055 ) | ( n1847 & n2055 ) ;
  assign n2058 = ( n1425 & n2056 ) | ( n1425 & n2057 ) | ( n2056 & n2057 ) ;
  assign n2059 = n2053 & ~n2058 ;
  assign n2060 = n207 | n329 ;
  assign n2061 = n2039 | n2060 ;
  assign n2062 = n2036 | n2061 ;
  assign n2063 = n197 | n471 ;
  assign n2064 = n577 | n2063 ;
  assign n2065 = ( n247 & ~n441 ) | ( n247 & n2064 ) | ( ~n441 & n2064 ) ;
  assign n2066 = n441 | n2065 ;
  assign n2067 = n498 & ~n2066 ;
  assign n2068 = ~n190 & n2067 ;
  assign n2069 = ~n2062 & n2068 ;
  assign n2070 = n382 | n2022 ;
  assign n2071 = n283 | n386 ;
  assign n2072 = n2070 | n2071 ;
  assign n2073 = n132 | n311 ;
  assign n2074 = n646 | n2073 ;
  assign n2075 = n248 | n2074 ;
  assign n2076 = n478 | n2075 ;
  assign n2077 = n2072 | n2076 ;
  assign n2078 = n543 | n2077 ;
  assign n2079 = n265 | n274 ;
  assign n2080 = ( n64 & n226 ) | ( n64 & n2079 ) | ( n226 & n2079 ) ;
  assign n2081 = ( n57 & n513 ) | ( n57 & n2080 ) | ( n513 & n2080 ) ;
  assign n2082 = n192 | n2081 ;
  assign n2083 = n2078 | n2082 ;
  assign n2084 = n2069 & ~n2083 ;
  assign n2085 = n2059 | n2084 ;
  assign n2086 = ( n1833 & ~n1834 ) | ( n1833 & n1861 ) | ( ~n1834 & n1861 ) ;
  assign n2087 = ( n1704 & ~n1833 ) | ( n1704 & n1834 ) | ( ~n1833 & n1834 ) ;
  assign n2088 = ( n1425 & n2086 ) | ( n1425 & ~n2087 ) | ( n2086 & ~n2087 ) ;
  assign n2089 = ( n1425 & ~n1704 ) | ( n1425 & n1861 ) | ( ~n1704 & n1861 ) ;
  assign n2090 = ~n1620 & n1833 ;
  assign n2091 = n2089 & n2090 ;
  assign n2092 = n2088 & ~n2091 ;
  assign n2093 = n348 | n397 ;
  assign n2094 = n125 | n356 ;
  assign n2095 = n2093 | n2094 ;
  assign n2096 = n187 | n457 ;
  assign n2097 = n297 | n2096 ;
  assign n2098 = n2095 | n2097 ;
  assign n2099 = n201 | n2098 ;
  assign n2100 = n387 | n503 ;
  assign n2101 = n444 | n2100 ;
  assign n2102 = n844 | n2101 ;
  assign n2103 = n179 | n380 ;
  assign n2104 = n1931 | n2103 ;
  assign n2105 = n197 | n2104 ;
  assign n2106 = n2102 | n2105 ;
  assign n2107 = n175 | n2106 ;
  assign n2108 = n2099 | n2107 ;
  assign n2109 = n128 | n258 ;
  assign n2110 = n284 | n477 ;
  assign n2111 = n2109 | n2110 ;
  assign n2112 = n238 | n325 ;
  assign n2113 = n336 | n2112 ;
  assign n2114 = ( ~n887 & n2111 ) | ( ~n887 & n2113 ) | ( n2111 & n2113 ) ;
  assign n2115 = n887 | n2114 ;
  assign n2116 = n2108 | n2115 ;
  assign n2117 = n164 | n282 ;
  assign n2118 = ( n64 & n251 ) | ( n64 & n405 ) | ( n251 & n405 ) ;
  assign n2119 = ( n57 & n349 ) | ( n57 & n2118 ) | ( n349 & n2118 ) ;
  assign n2120 = n2117 | n2119 ;
  assign n2121 = n597 | n2120 ;
  assign n2122 = n2116 | n2121 ;
  assign n2123 = ~n2092 & n2122 ;
  assign n2124 = n2059 & n2084 ;
  assign n2125 = n2085 & ~n2124 ;
  assign n2126 = n2123 & n2125 ;
  assign n2127 = n2085 & ~n2126 ;
  assign n2128 = n2049 | n2127 ;
  assign n2129 = n2049 | n2124 ;
  assign n2130 = n2092 | n2123 ;
  assign n2131 = n2092 & n2122 ;
  assign n2132 = n2130 & ~n2131 ;
  assign n2133 = ( n1425 & ~n1703 ) | ( n1425 & n1860 ) | ( ~n1703 & n1860 ) ;
  assign n2134 = n1622 & ~n1658 ;
  assign n2135 = n2133 & n2134 ;
  assign n2136 = n2089 & ~n2135 ;
  assign n2137 = n133 | n325 ;
  assign n2138 = n97 | n2137 ;
  assign n2139 = n284 | n348 ;
  assign n2140 = n406 | n2139 ;
  assign n2141 = n2138 | n2140 ;
  assign n2142 = n510 | n778 ;
  assign n2143 = n2141 | n2142 ;
  assign n2144 = n385 | n2143 ;
  assign n2145 = n1978 | n2144 ;
  assign n2146 = n176 | n911 ;
  assign n2147 = n910 | n2146 ;
  assign n2148 = n908 | n2147 ;
  assign n2149 = n218 | n519 ;
  assign n2150 = n280 | n295 ;
  assign n2151 = n2149 | n2150 ;
  assign n2152 = n853 | n2151 ;
  assign n2153 = n128 | n207 ;
  assign n2154 = n134 | n2153 ;
  assign n2155 = n2152 | n2154 ;
  assign n2156 = n2148 | n2155 ;
  assign n2157 = n2145 | n2156 ;
  assign n2158 = n2136 & ~n2157 ;
  assign n2159 = n2132 | n2158 ;
  assign n2160 = n1660 & n1682 ;
  assign n2161 = n1660 & ~n1680 ;
  assign n2162 = ( ~n1702 & n2160 ) | ( ~n1702 & n2161 ) | ( n2160 & n2161 ) ;
  assign n2163 = n1859 & n2161 ;
  assign n2164 = ( n1425 & n2162 ) | ( n1425 & n2163 ) | ( n2162 & n2163 ) ;
  assign n2165 = n2133 & ~n2164 ;
  assign n2166 = n285 | n1941 ;
  assign n2167 = n1937 | n2166 ;
  assign n2168 = n369 | n399 ;
  assign n2169 = n387 | n2168 ;
  assign n2170 = n192 | n267 ;
  assign n2171 = n185 | n2170 ;
  assign n2172 = n2169 | n2171 ;
  assign n2173 = n166 | n319 ;
  assign n2174 = n147 | n2173 ;
  assign n2175 = n2172 | n2174 ;
  assign n2176 = n384 | n2175 ;
  assign n2177 = n149 | n367 ;
  assign n2178 = n101 | n2177 ;
  assign n2179 = n405 | n577 ;
  assign n2180 = n2178 | n2179 ;
  assign n2181 = n874 | n2180 ;
  assign n2182 = n204 | n359 ;
  assign n2183 = n639 | n2182 ;
  assign n2184 = n127 | n2183 ;
  assign n2185 = n453 | n2184 ;
  assign n2186 = n2181 | n2185 ;
  assign n2187 = n2176 | n2186 ;
  assign n2188 = n2167 | n2187 ;
  assign n2189 = n226 | n544 ;
  assign n2190 = n175 | n231 ;
  assign n2191 = n2189 | n2190 ;
  assign n2192 = n2188 | n2191 ;
  assign n2193 = ~n2165 & n2192 ;
  assign n2194 = ( ~n2136 & n2157 ) | ( ~n2136 & n2193 ) | ( n2157 & n2193 ) ;
  assign n2195 = ~n2132 & n2194 ;
  assign n2196 = n2165 & ~n2192 ;
  assign n2197 = n2193 | n2196 ;
  assign n2198 = n1702 & ~n1854 ;
  assign n2199 = ( n1425 & n1859 ) | ( n1425 & ~n2198 ) | ( n1859 & ~n2198 ) ;
  assign n2200 = ~n1702 & n1854 ;
  assign n2201 = n1854 & ~n1855 ;
  assign n2202 = n1858 & n2201 ;
  assign n2203 = ( n1425 & n2200 ) | ( n1425 & n2202 ) | ( n2200 & n2202 ) ;
  assign n2204 = n2199 & ~n2203 ;
  assign n2205 = n457 | n481 ;
  assign n2206 = n101 | n234 ;
  assign n2207 = n2205 | n2206 ;
  assign n2208 = n329 | n2207 ;
  assign n2209 = n720 | n2019 ;
  assign n2210 = n353 | n870 ;
  assign n2211 = n2209 | n2210 ;
  assign n2212 = n274 | n705 ;
  assign n2213 = n176 | n238 ;
  assign n2214 = n2212 | n2213 ;
  assign n2215 = n2211 | n2214 ;
  assign n2216 = n312 | n368 ;
  assign n2217 = n164 | n305 ;
  assign n2218 = n267 | n2217 ;
  assign n2219 = n2216 | n2218 ;
  assign n2220 = n248 | n2219 ;
  assign n2221 = n711 | n2220 ;
  assign n2222 = n2215 | n2221 ;
  assign n2223 = n258 | n548 ;
  assign n2224 = n151 | n2223 ;
  assign n2225 = n224 | n249 ;
  assign n2226 = n211 | n2225 ;
  assign n2227 = n2224 | n2226 ;
  assign n2228 = n617 | n2227 ;
  assign n2229 = n2222 | n2228 ;
  assign n2230 = n2208 | n2229 ;
  assign n2231 = n382 | n655 ;
  assign n2232 = n256 | n604 ;
  assign n2233 = n498 & ~n2232 ;
  assign n2234 = ~n2231 & n2233 ;
  assign n2235 = ~n2220 & n2234 ;
  assign n2236 = n547 | n869 ;
  assign n2237 = n2235 & ~n2236 ;
  assign n2238 = n698 | n701 ;
  assign n2239 = n697 | n2238 ;
  assign n2240 = n2237 & ~n2239 ;
  assign n2241 = n185 | n478 ;
  assign n2242 = n132 | n291 ;
  assign n2243 = n2241 | n2242 ;
  assign n2244 = n321 | n2243 ;
  assign n2245 = n149 | n329 ;
  assign n2246 = n894 | n2245 ;
  assign n2247 = n2064 | n2246 ;
  assign n2248 = n2244 | n2247 ;
  assign n2249 = n231 | n1021 ;
  assign n2250 = n857 | n2249 ;
  assign n2251 = n459 | n2151 ;
  assign n2252 = n2250 | n2251 ;
  assign n2253 = n2248 | n2252 ;
  assign n2254 = n176 | n2253 ;
  assign n2255 = n154 | n250 ;
  assign n2256 = n108 | n274 ;
  assign n2257 = n2255 | n2256 ;
  assign n2258 = n97 | n2257 ;
  assign n2259 = n2254 | n2258 ;
  assign n2260 = n2240 & ~n2259 ;
  assign n2261 = ( n1425 & n1698 ) | ( n1425 & ~n1701 ) | ( n1698 & ~n1701 ) ;
  assign n2262 = n1857 & n2261 ;
  assign n2263 = n1857 & ~n2262 ;
  assign n2264 = ( n2261 & ~n2262 ) | ( n2261 & n2263 ) | ( ~n2262 & n2263 ) ;
  assign n2265 = ( n1425 & n1699 ) | ( n1425 & ~n1700 ) | ( n1699 & ~n1700 ) ;
  assign n2266 = ~n1173 & n1699 ;
  assign n2267 = n1425 & n2266 ;
  assign n2268 = n2265 & ~n2267 ;
  assign n2269 = n784 | n2245 ;
  assign n2270 = n320 | n2269 ;
  assign n2271 = n1978 | n2270 ;
  assign n2272 = n399 | n513 ;
  assign n2273 = n120 | n273 ;
  assign n2274 = n2272 | n2273 ;
  assign n2275 = n165 | n2274 ;
  assign n2276 = n207 | n397 ;
  assign n2277 = n504 | n2276 ;
  assign n2278 = n101 | n175 ;
  assign n2279 = n2277 | n2278 ;
  assign n2280 = n2275 | n2279 ;
  assign n2281 = n179 | n265 ;
  assign n2282 = n311 | n471 ;
  assign n2283 = n2281 | n2282 ;
  assign n2284 = n168 | n2283 ;
  assign n2285 = n2280 | n2284 ;
  assign n2286 = n2271 | n2285 ;
  assign n2287 = n155 | n380 ;
  assign n2288 = n253 | n2287 ;
  assign n2289 = n676 | n2288 ;
  assign n2290 = n391 | n2289 ;
  assign n2291 = n267 | n356 ;
  assign n2292 = n187 | n597 ;
  assign n2293 = n2291 | n2292 ;
  assign n2294 = n2290 | n2293 ;
  assign n2295 = n2286 | n2294 ;
  assign n2296 = n519 | n877 ;
  assign n2297 = n540 | n594 ;
  assign n2298 = n2296 | n2297 ;
  assign n2299 = n459 | n2298 ;
  assign n2300 = n2215 | n2299 ;
  assign n2301 = n609 | n2300 ;
  assign n2302 = n239 | n391 ;
  assign n2303 = n219 | n478 ;
  assign n2304 = n2302 | n2303 ;
  assign n2305 = n170 | n369 ;
  assign n2306 = n2304 | n2305 ;
  assign n2307 = n2301 | n2306 ;
  assign n2308 = n1175 & n1424 ;
  assign n2309 = n1425 & ~n2308 ;
  assign n2310 = ~n2307 & n2309 ;
  assign n2311 = ( n2268 & ~n2295 ) | ( n2268 & n2310 ) | ( ~n2295 & n2310 ) ;
  assign n2312 = ( n2260 & n2264 ) | ( n2260 & n2311 ) | ( n2264 & n2311 ) ;
  assign n2313 = ( n2204 & ~n2230 ) | ( n2204 & n2312 ) | ( ~n2230 & n2312 ) ;
  assign n2314 = n2197 | n2313 ;
  assign n2315 = ( n2159 & ~n2195 ) | ( n2159 & n2314 ) | ( ~n2195 & n2314 ) ;
  assign n2316 = ( n2128 & n2129 ) | ( n2128 & n2315 ) | ( n2129 & n2315 ) ;
  assign n2317 = ( n1995 & n2047 ) | ( n1995 & n2316 ) | ( n2047 & n2316 ) ;
  assign n2318 = n120 | n290 ;
  assign n2319 = n321 | n2318 ;
  assign n2320 = n693 | n2178 ;
  assign n2321 = n606 | n2320 ;
  assign n2322 = n598 | n2321 ;
  assign n2323 = n590 | n2322 ;
  assign n2324 = n351 | n513 ;
  assign n2325 = n397 | n2324 ;
  assign n2326 = n155 | n205 ;
  assign n2327 = n227 | n2326 ;
  assign n2328 = n209 | n2327 ;
  assign n2329 = n2325 | n2328 ;
  assign n2330 = n171 | n2329 ;
  assign n2331 = n147 | n405 ;
  assign n2332 = n127 | n391 ;
  assign n2333 = n2331 | n2332 ;
  assign n2334 = n219 | n2333 ;
  assign n2335 = n238 | n271 ;
  assign n2336 = n213 | n2335 ;
  assign n2337 = n2034 | n2336 ;
  assign n2338 = n2334 | n2337 ;
  assign n2339 = n158 | n224 ;
  assign n2340 = n273 | n280 ;
  assign n2341 = n2339 | n2340 ;
  assign n2342 = n197 | n2341 ;
  assign n2343 = n132 | n705 ;
  assign n2344 = n239 | n325 ;
  assign n2345 = n2343 | n2344 ;
  assign n2346 = n234 | n2345 ;
  assign n2347 = n2342 | n2346 ;
  assign n2348 = n2338 | n2347 ;
  assign n2349 = n2330 | n2348 ;
  assign n2350 = n2323 | n2349 ;
  assign n2351 = n2319 | n2350 ;
  assign n2352 = n2317 | n2351 ;
  assign n2353 = n2317 & n2351 ;
  assign n2354 = n2352 & ~n2353 ;
  assign n2355 = ~n32 & n421 ;
  assign n2356 = n32 & ~n421 ;
  assign n2357 = n2355 | n2356 ;
  assign n2358 = x2 & x22 ;
  assign n2359 = x0 | x1 ;
  assign n2360 = x2 & n2359 ;
  assign n2361 = n431 & ~n2360 ;
  assign n2362 = n2358 | n2361 ;
  assign n2363 = ~n434 & n2362 ;
  assign n2364 = n434 & ~n2362 ;
  assign n2365 = n2363 | n2364 ;
  assign n2366 = ~n2357 & n2365 ;
  assign n2367 = n2354 & n2366 ;
  assign n2368 = ~n1964 & n1990 ;
  assign n2369 = ~n1930 & n2368 ;
  assign n2370 = ( n1990 & n1993 ) | ( n1990 & n2369 ) | ( n1993 & n2369 ) ;
  assign n2371 = ( ~n1908 & n2369 ) | ( ~n1908 & n2370 ) | ( n2369 & n2370 ) ;
  assign n2372 = ( n2046 & n2369 ) | ( n2046 & n2370 ) | ( n2369 & n2370 ) ;
  assign n2373 = ( ~n2316 & n2371 ) | ( ~n2316 & n2372 ) | ( n2371 & n2372 ) ;
  assign n2374 = n2317 | n2373 ;
  assign n2375 = n421 & ~n434 ;
  assign n2376 = ~n421 & n434 ;
  assign n2377 = n2375 | n2376 ;
  assign n2378 = ~n2365 & n2377 ;
  assign n2379 = n2374 & n2378 ;
  assign n2380 = n2357 & ~n2365 ;
  assign n2381 = ~n2377 & n2380 ;
  assign n2382 = ( n1908 & ~n2046 ) | ( n1908 & n2316 ) | ( ~n2046 & n2316 ) ;
  assign n2383 = n1993 | n2382 ;
  assign n2384 = n1993 & n2382 ;
  assign n2385 = ( n2381 & ~n2383 ) | ( n2381 & n2384 ) | ( ~n2383 & n2384 ) ;
  assign n2386 = n2379 | n2385 ;
  assign n2387 = n2367 | n2386 ;
  assign n2388 = n2357 & n2365 ;
  assign n2389 = n32 & n2388 ;
  assign n2390 = n2049 & n2127 ;
  assign n2391 = n2049 & n2124 ;
  assign n2392 = ( n2315 & n2390 ) | ( n2315 & n2391 ) | ( n2390 & n2391 ) ;
  assign n2393 = n2316 & ~n2392 ;
  assign n2394 = ~n2124 & n2127 ;
  assign n2395 = n2315 & n2394 ;
  assign n2396 = ~n2123 & n2315 ;
  assign n2397 = n2125 | n2396 ;
  assign n2398 = ~n2395 & n2397 ;
  assign n2399 = ~n2393 & n2398 ;
  assign n2400 = ( n2158 & ~n2194 ) | ( n2158 & n2314 ) | ( ~n2194 & n2314 ) ;
  assign n2401 = n2132 & ~n2400 ;
  assign n2402 = ~n2132 & n2315 ;
  assign n2403 = n2401 | n2402 ;
  assign n2404 = n2158 | n2194 ;
  assign n2405 = n2314 & ~n2404 ;
  assign n2406 = ~n2136 & n2157 ;
  assign n2407 = ~n2193 & n2314 ;
  assign n2408 = n2158 & ~n2407 ;
  assign n2409 = ( n2406 & ~n2407 ) | ( n2406 & n2408 ) | ( ~n2407 & n2408 ) ;
  assign n2410 = n2405 | n2409 ;
  assign n2411 = n2403 & n2410 ;
  assign n2412 = n2403 | n2410 ;
  assign n2413 = ~n2411 & n2412 ;
  assign n2414 = n2197 & n2313 ;
  assign n2415 = n2314 & ~n2414 ;
  assign n2416 = n2410 & n2415 ;
  assign n2417 = n2413 & n2416 ;
  assign n2418 = n2405 | n2415 ;
  assign n2419 = n2409 | n2418 ;
  assign n2420 = ~n2416 & n2419 ;
  assign n2421 = ( ~n2204 & n2230 ) | ( ~n2204 & n2313 ) | ( n2230 & n2313 ) ;
  assign n2422 = ( ~n2312 & n2313 ) | ( ~n2312 & n2421 ) | ( n2313 & n2421 ) ;
  assign n2423 = n2415 & n2422 ;
  assign n2424 = ( n2260 & n2311 ) | ( n2260 & ~n2312 ) | ( n2311 & ~n2312 ) ;
  assign n2425 = ( n2264 & ~n2312 ) | ( n2264 & n2424 ) | ( ~n2312 & n2424 ) ;
  assign n2426 = n2422 & ~n2425 ;
  assign n2427 = ~n2422 & n2425 ;
  assign n2428 = n2426 | n2427 ;
  assign n2429 = n2268 & ~n2295 ;
  assign n2430 = n2311 & ~n2429 ;
  assign n2431 = ~n2268 & n2295 ;
  assign n2432 = ( ~n2310 & n2429 ) | ( ~n2310 & n2431 ) | ( n2429 & n2431 ) ;
  assign n2433 = n2430 | n2432 ;
  assign n2434 = n2307 & ~n2309 ;
  assign n2435 = n2310 | n2434 ;
  assign n2436 = n2433 & ~n2435 ;
  assign n2437 = ~n2425 & n2436 ;
  assign n2438 = ( n2433 & n2435 ) | ( n2433 & n2437 ) | ( n2435 & n2437 ) ;
  assign n2439 = ~n2428 & n2438 ;
  assign n2440 = n2415 | n2422 ;
  assign n2441 = ~n2423 & n2440 ;
  assign n2442 = ( n2426 & n2439 ) | ( n2426 & n2441 ) | ( n2439 & n2441 ) ;
  assign n2443 = ( n2420 & n2423 ) | ( n2420 & n2442 ) | ( n2423 & n2442 ) ;
  assign n2444 = ( n2413 & n2417 ) | ( n2413 & n2443 ) | ( n2417 & n2443 ) ;
  assign n2445 = ~n2398 & n2403 ;
  assign n2446 = n2398 & ~n2403 ;
  assign n2447 = n2445 | n2446 ;
  assign n2448 = ( n2411 & n2444 ) | ( n2411 & ~n2447 ) | ( n2444 & ~n2447 ) ;
  assign n2449 = ( n2393 & ~n2398 ) | ( n2393 & n2445 ) | ( ~n2398 & n2445 ) ;
  assign n2450 = ( ~n2399 & n2448 ) | ( ~n2399 & n2449 ) | ( n2448 & n2449 ) ;
  assign n2451 = n1906 | n2045 ;
  assign n2452 = n2316 & ~n2451 ;
  assign n2453 = ~n2044 & n2316 ;
  assign n2454 = ~n1892 & n1905 ;
  assign n2455 = ~n2453 & n2454 ;
  assign n2456 = ( n1906 & ~n2453 ) | ( n1906 & n2455 ) | ( ~n2453 & n2455 ) ;
  assign n2457 = n2452 | n2456 ;
  assign n2458 = ( n1906 & ~n2045 ) | ( n1906 & n2316 ) | ( ~n2045 & n2316 ) ;
  assign n2459 = ( n264 & ~n1882 ) | ( n264 & n2458 ) | ( ~n1882 & n2458 ) ;
  assign n2460 = ( ~n264 & n1882 ) | ( ~n264 & n2459 ) | ( n1882 & n2459 ) ;
  assign n2461 = ( ~n2458 & n2459 ) | ( ~n2458 & n2460 ) | ( n2459 & n2460 ) ;
  assign n2462 = n2393 | n2452 ;
  assign n2463 = n2456 | n2462 ;
  assign n2464 = ( n2457 & n2461 ) | ( n2457 & n2463 ) | ( n2461 & n2463 ) ;
  assign n2465 = n2393 & n2457 ;
  assign n2466 = ( n2457 & n2461 ) | ( n2457 & n2465 ) | ( n2461 & n2465 ) ;
  assign n2467 = ( n2450 & n2464 ) | ( n2450 & n2466 ) | ( n2464 & n2466 ) ;
  assign n2468 = n2383 & ~n2384 ;
  assign n2469 = ~n2461 & n2468 ;
  assign n2470 = ~n2374 & n2468 ;
  assign n2471 = ( n2383 & n2469 ) | ( n2383 & n2470 ) | ( n2469 & n2470 ) ;
  assign n2472 = n2374 & ~n2468 ;
  assign n2473 = n2461 & ~n2468 ;
  assign n2474 = n2472 | n2473 ;
  assign n2475 = ( n2467 & ~n2471 ) | ( n2467 & n2474 ) | ( ~n2471 & n2474 ) ;
  assign n2476 = ( n2354 & ~n2374 ) | ( n2354 & n2475 ) | ( ~n2374 & n2475 ) ;
  assign n2477 = ( ~n2354 & n2374 ) | ( ~n2354 & n2476 ) | ( n2374 & n2476 ) ;
  assign n2478 = ( ~n2475 & n2476 ) | ( ~n2475 & n2477 ) | ( n2476 & n2477 ) ;
  assign n2479 = n2389 & n2478 ;
  assign n2480 = ( n32 & n2387 ) | ( n32 & n2479 ) | ( n2387 & n2479 ) ;
  assign n2481 = n32 | n2388 ;
  assign n2482 = ( n32 & n2478 ) | ( n32 & n2481 ) | ( n2478 & n2481 ) ;
  assign n2483 = n2387 | n2482 ;
  assign n2484 = ~n2480 & n2483 ;
  assign n2485 = n566 & n2435 ;
  assign n2486 = ~n977 & n985 ;
  assign n2487 = n977 & ~n985 ;
  assign n2488 = n2486 | n2487 ;
  assign n2489 = n2435 & n2488 ;
  assign n2490 = n566 & ~n2489 ;
  assign n2491 = n1923 & n2488 ;
  assign n2492 = ~n2432 & n2435 ;
  assign n2493 = ~n2430 & n2492 ;
  assign n2494 = n2436 | n2493 ;
  assign n2495 = n2491 & n2494 ;
  assign n2496 = ~n493 & n985 ;
  assign n2497 = n493 & ~n985 ;
  assign n2498 = n2496 | n2497 ;
  assign n2499 = ~n2488 & n2498 ;
  assign n2500 = n2435 & n2499 ;
  assign n2501 = ~n1923 & n2488 ;
  assign n2502 = n2433 & n2501 ;
  assign n2503 = n2500 | n2502 ;
  assign n2504 = n2495 | n2503 ;
  assign n2505 = ~n566 & n2504 ;
  assign n2506 = n566 & ~n2504 ;
  assign n2507 = ( n2490 & n2505 ) | ( n2490 & n2506 ) | ( n2505 & n2506 ) ;
  assign n2508 = ~n2425 & n2501 ;
  assign n2509 = n2425 & ~n2436 ;
  assign n2510 = n2437 | n2509 ;
  assign n2511 = n1923 & ~n2488 ;
  assign n2512 = ~n2498 & n2511 ;
  assign n2513 = n2435 & n2512 ;
  assign n2514 = n2433 & n2499 ;
  assign n2515 = n2513 | n2514 ;
  assign n2516 = n2508 | n2515 ;
  assign n2517 = n2510 & ~n2516 ;
  assign n2518 = n2491 | n2515 ;
  assign n2519 = ( n2508 & ~n2517 ) | ( n2508 & n2518 ) | ( ~n2517 & n2518 ) ;
  assign n2520 = ( ~n566 & n2517 ) | ( ~n566 & n2519 ) | ( n2517 & n2519 ) ;
  assign n2521 = n2519 & ~n2520 ;
  assign n2522 = ~n2517 & n2520 ;
  assign n2523 = ( n566 & ~n2521 ) | ( n566 & n2522 ) | ( ~n2521 & n2522 ) ;
  assign n2524 = n2507 & n2523 ;
  assign n2525 = n2485 | n2524 ;
  assign n2526 = n2485 & n2524 ;
  assign n2527 = n2525 & ~n2526 ;
  assign n2528 = n2438 & ~n2439 ;
  assign n2529 = n2428 | n2439 ;
  assign n2530 = ~n2528 & n2529 ;
  assign n2531 = ~n2425 & n2499 ;
  assign n2532 = n2433 & n2512 ;
  assign n2533 = n2501 | n2532 ;
  assign n2534 = ( n2422 & n2532 ) | ( n2422 & n2533 ) | ( n2532 & n2533 ) ;
  assign n2535 = n2531 | n2534 ;
  assign n2536 = ( n2491 & ~n2530 ) | ( n2491 & n2535 ) | ( ~n2530 & n2535 ) ;
  assign n2537 = ( n566 & n2535 ) | ( n566 & ~n2536 ) | ( n2535 & ~n2536 ) ;
  assign n2538 = n2536 | n2537 ;
  assign n2539 = ~n2535 & n2537 ;
  assign n2540 = ( ~n566 & n2538 ) | ( ~n566 & n2539 ) | ( n2538 & n2539 ) ;
  assign n2541 = n2527 & ~n2540 ;
  assign n2542 = ~n2527 & n2540 ;
  assign n2543 = n2541 | n2542 ;
  assign n2544 = n2413 | n2416 ;
  assign n2545 = n2443 | n2544 ;
  assign n2546 = ~n2444 & n2545 ;
  assign n2547 = n752 & ~n948 ;
  assign n2548 = ~n752 & n948 ;
  assign n2549 = n2547 | n2548 ;
  assign n2550 = n943 & ~n977 ;
  assign n2551 = ~n943 & n977 ;
  assign n2552 = n2550 | n2551 ;
  assign n2553 = n943 & ~n948 ;
  assign n2554 = ~n943 & n948 ;
  assign n2555 = n2553 | n2554 ;
  assign n2556 = n2552 & ~n2555 ;
  assign n2557 = ~n2549 & n2556 ;
  assign n2558 = n2415 & n2557 ;
  assign n2559 = ~n2549 & n2555 ;
  assign n2560 = ( n2405 & n2409 ) | ( n2405 & n2559 ) | ( n2409 & n2559 ) ;
  assign n2561 = n2558 | n2560 ;
  assign n2562 = n2549 & n2552 ;
  assign n2563 = n2549 & ~n2552 ;
  assign n2564 = n2403 & n2563 ;
  assign n2565 = n2562 | n2564 ;
  assign n2566 = n2561 | n2565 ;
  assign n2567 = n977 & n2566 ;
  assign n2568 = n977 & n2564 ;
  assign n2569 = ( n977 & n2561 ) | ( n977 & n2568 ) | ( n2561 & n2568 ) ;
  assign n2570 = ( n2546 & n2567 ) | ( n2546 & n2569 ) | ( n2567 & n2569 ) ;
  assign n2571 = n977 | n2566 ;
  assign n2572 = n977 | n2564 ;
  assign n2573 = n2561 | n2572 ;
  assign n2574 = ( n2546 & n2571 ) | ( n2546 & n2573 ) | ( n2571 & n2573 ) ;
  assign n2575 = ~n2570 & n2574 ;
  assign n2576 = n2543 & n2575 ;
  assign n2577 = n2543 & ~n2576 ;
  assign n2578 = n2422 & n2557 ;
  assign n2579 = n2415 & n2559 ;
  assign n2580 = n2578 | n2579 ;
  assign n2581 = ( n2405 & n2409 ) | ( n2405 & n2563 ) | ( n2409 & n2563 ) ;
  assign n2582 = n2580 | n2581 ;
  assign n2583 = n2420 | n2423 ;
  assign n2584 = n2442 | n2583 ;
  assign n2585 = ~n2443 & n2584 ;
  assign n2586 = n977 & n2562 ;
  assign n2587 = n2585 & n2586 ;
  assign n2588 = ( n977 & n2582 ) | ( n977 & n2587 ) | ( n2582 & n2587 ) ;
  assign n2589 = n977 | n2562 ;
  assign n2590 = ( n977 & n2585 ) | ( n977 & n2589 ) | ( n2585 & n2589 ) ;
  assign n2591 = n2582 | n2590 ;
  assign n2592 = ~n2588 & n2591 ;
  assign n2593 = n2507 | n2523 ;
  assign n2594 = ~n2524 & n2593 ;
  assign n2595 = n2592 & n2594 ;
  assign n2596 = n2592 | n2594 ;
  assign n2597 = ~n2595 & n2596 ;
  assign n2598 = n2490 | n2506 ;
  assign n2599 = n2505 | n2598 ;
  assign n2600 = ~n2507 & n2599 ;
  assign n2601 = n2422 & n2559 ;
  assign n2602 = n2415 & n2563 ;
  assign n2603 = n2601 | n2602 ;
  assign n2604 = ~n2425 & n2557 ;
  assign n2605 = n2603 | n2604 ;
  assign n2606 = n2426 | n2439 ;
  assign n2607 = n2441 | n2606 ;
  assign n2608 = ~n2442 & n2607 ;
  assign n2609 = n2562 | n2605 ;
  assign n2610 = ( n2605 & n2608 ) | ( n2605 & n2609 ) | ( n2608 & n2609 ) ;
  assign n2611 = n977 & n2610 ;
  assign n2612 = n977 & ~n2611 ;
  assign n2613 = ( n2610 & ~n2611 ) | ( n2610 & n2612 ) | ( ~n2611 & n2612 ) ;
  assign n2614 = n2600 & n2613 ;
  assign n2615 = n2600 | n2613 ;
  assign n2616 = ~n2614 & n2615 ;
  assign n2617 = ~n2425 & n2563 ;
  assign n2618 = n2435 & n2557 ;
  assign n2619 = n2433 & n2559 ;
  assign n2620 = n2618 | n2619 ;
  assign n2621 = n2617 | n2620 ;
  assign n2622 = n2510 & ~n2621 ;
  assign n2623 = n2562 | n2620 ;
  assign n2624 = ( n2617 & ~n2622 ) | ( n2617 & n2623 ) | ( ~n2622 & n2623 ) ;
  assign n2625 = ( ~n977 & n2622 ) | ( ~n977 & n2624 ) | ( n2622 & n2624 ) ;
  assign n2626 = n2624 & ~n2625 ;
  assign n2627 = ~n2622 & n2625 ;
  assign n2628 = ( n977 & ~n2626 ) | ( n977 & n2627 ) | ( ~n2626 & n2627 ) ;
  assign n2629 = n2435 & n2549 ;
  assign n2630 = n977 & ~n2629 ;
  assign n2631 = n2494 & n2562 ;
  assign n2632 = n2435 & n2559 ;
  assign n2633 = n2631 | n2632 ;
  assign n2634 = n2433 & n2563 ;
  assign n2635 = ~n2633 & n2634 ;
  assign n2636 = ( n977 & ~n2633 ) | ( n977 & n2635 ) | ( ~n2633 & n2635 ) ;
  assign n2637 = ( n977 & n2635 ) | ( n977 & ~n2636 ) | ( n2635 & ~n2636 ) ;
  assign n2638 = ( n2633 & n2636 ) | ( n2633 & ~n2637 ) | ( n2636 & ~n2637 ) ;
  assign n2639 = n2630 & n2638 ;
  assign n2640 = n2489 & n2639 ;
  assign n2641 = n2628 & n2640 ;
  assign n2642 = ~n2425 & n2559 ;
  assign n2643 = n2433 & n2557 ;
  assign n2644 = n2563 | n2643 ;
  assign n2645 = ( n2422 & n2643 ) | ( n2422 & n2644 ) | ( n2643 & n2644 ) ;
  assign n2646 = n2642 | n2645 ;
  assign n2647 = ~n2530 & n2586 ;
  assign n2648 = ( n977 & n2646 ) | ( n977 & n2647 ) | ( n2646 & n2647 ) ;
  assign n2649 = ( n977 & ~n2530 ) | ( n977 & n2589 ) | ( ~n2530 & n2589 ) ;
  assign n2650 = n2646 | n2649 ;
  assign n2651 = ~n2648 & n2650 ;
  assign n2652 = n2628 & n2639 ;
  assign n2653 = n2489 | n2652 ;
  assign n2654 = ~n2641 & n2653 ;
  assign n2655 = n2651 & n2654 ;
  assign n2656 = n2641 | n2655 ;
  assign n2657 = n2616 & n2656 ;
  assign n2658 = n2614 | n2657 ;
  assign n2659 = n2597 & n2658 ;
  assign n2660 = n2595 | n2659 ;
  assign n2661 = ~n2541 & n2575 ;
  assign n2662 = ~n2542 & n2661 ;
  assign n2663 = n2660 | n2662 ;
  assign n2664 = n2577 | n2663 ;
  assign n2665 = ( n2577 & n2660 ) | ( n2577 & n2662 ) | ( n2660 & n2662 ) ;
  assign n2666 = n2664 & ~n2665 ;
  assign n2667 = ~n32 & n822 ;
  assign n2668 = n32 & ~n822 ;
  assign n2669 = n2667 | n2668 ;
  assign n2670 = ~n756 & n822 ;
  assign n2671 = n756 & ~n822 ;
  assign n2672 = n2670 | n2671 ;
  assign n2673 = ~n2669 & n2672 ;
  assign n2674 = n2393 & n2673 ;
  assign n2675 = n752 & ~n756 ;
  assign n2676 = ~n752 & n756 ;
  assign n2677 = n2675 | n2676 ;
  assign n2678 = n2669 | n2672 ;
  assign n2679 = n2677 & ~n2678 ;
  assign n2680 = ~n2398 & n2679 ;
  assign n2681 = n2674 | n2680 ;
  assign n2682 = n2669 & ~n2677 ;
  assign n2683 = ( n2452 & n2456 ) | ( n2452 & n2682 ) | ( n2456 & n2682 ) ;
  assign n2684 = n2681 | n2683 ;
  assign n2685 = n752 | n2684 ;
  assign n2686 = n2669 & n2677 ;
  assign n2687 = ( n2393 & n2450 ) | ( n2393 & ~n2457 ) | ( n2450 & ~n2457 ) ;
  assign n2688 = ( ~n2450 & n2457 ) | ( ~n2450 & n2687 ) | ( n2457 & n2687 ) ;
  assign n2689 = ( ~n2393 & n2687 ) | ( ~n2393 & n2688 ) | ( n2687 & n2688 ) ;
  assign n2690 = ( n2685 & n2686 ) | ( n2685 & n2689 ) | ( n2686 & n2689 ) ;
  assign n2691 = n2685 | n2690 ;
  assign n2692 = n752 & n2686 ;
  assign n2693 = n2689 & n2692 ;
  assign n2694 = ( n752 & n2684 ) | ( n752 & n2693 ) | ( n2684 & n2693 ) ;
  assign n2695 = n2691 & ~n2694 ;
  assign n2696 = n2666 & n2695 ;
  assign n2697 = n2666 & ~n2696 ;
  assign n2698 = ( n2695 & ~n2696 ) | ( n2695 & n2697 ) | ( ~n2696 & n2697 ) ;
  assign n2699 = n2597 | n2658 ;
  assign n2700 = ~n2659 & n2699 ;
  assign n2701 = n2403 & n2673 ;
  assign n2702 = ( n2405 & n2409 ) | ( n2405 & n2679 ) | ( n2409 & n2679 ) ;
  assign n2703 = n2701 | n2702 ;
  assign n2704 = ~n2398 & n2682 ;
  assign n2705 = n2703 | n2704 ;
  assign n2706 = ~n2411 & n2447 ;
  assign n2707 = ~n2444 & n2706 ;
  assign n2708 = n2448 | n2707 ;
  assign n2709 = n2686 | n2705 ;
  assign n2710 = ( n2705 & ~n2708 ) | ( n2705 & n2709 ) | ( ~n2708 & n2709 ) ;
  assign n2711 = ~n752 & n2710 ;
  assign n2712 = n752 & ~n2710 ;
  assign n2713 = n2711 | n2712 ;
  assign n2714 = n2616 | n2656 ;
  assign n2715 = ~n2657 & n2714 ;
  assign n2716 = n2415 & n2679 ;
  assign n2717 = ( n2405 & n2409 ) | ( n2405 & n2673 ) | ( n2409 & n2673 ) ;
  assign n2718 = n2716 | n2717 ;
  assign n2719 = n2403 & n2682 ;
  assign n2720 = n2718 | n2719 ;
  assign n2721 = n2686 | n2720 ;
  assign n2722 = ( n2546 & n2720 ) | ( n2546 & n2721 ) | ( n2720 & n2721 ) ;
  assign n2723 = n752 & n2722 ;
  assign n2724 = n752 & ~n2723 ;
  assign n2725 = ( n2722 & ~n2723 ) | ( n2722 & n2724 ) | ( ~n2723 & n2724 ) ;
  assign n2726 = n2654 & ~n2655 ;
  assign n2727 = ( n2651 & ~n2655 ) | ( n2651 & n2726 ) | ( ~n2655 & n2726 ) ;
  assign n2728 = n2725 & n2727 ;
  assign n2729 = n2725 | n2727 ;
  assign n2730 = ~n2728 & n2729 ;
  assign n2731 = n2628 | n2639 ;
  assign n2732 = ~n2652 & n2731 ;
  assign n2733 = n2422 & n2679 ;
  assign n2734 = n2415 & n2673 ;
  assign n2735 = n2733 | n2734 ;
  assign n2736 = ( n2405 & n2409 ) | ( n2405 & n2682 ) | ( n2409 & n2682 ) ;
  assign n2737 = n2735 | n2736 ;
  assign n2738 = ( n2585 & n2686 ) | ( n2585 & n2737 ) | ( n2686 & n2737 ) ;
  assign n2739 = ( n752 & ~n2737 ) | ( n752 & n2738 ) | ( ~n2737 & n2738 ) ;
  assign n2740 = ~n2738 & n2739 ;
  assign n2741 = n2737 | n2739 ;
  assign n2742 = ( ~n752 & n2740 ) | ( ~n752 & n2741 ) | ( n2740 & n2741 ) ;
  assign n2743 = n2732 | n2742 ;
  assign n2744 = n2630 | n2638 ;
  assign n2745 = ~n2639 & n2744 ;
  assign n2746 = n2422 & n2673 ;
  assign n2747 = n2415 & n2682 ;
  assign n2748 = n2746 | n2747 ;
  assign n2749 = ~n2425 & n2679 ;
  assign n2750 = n2748 | n2749 ;
  assign n2751 = n2686 | n2750 ;
  assign n2752 = ( n2608 & n2750 ) | ( n2608 & n2751 ) | ( n2750 & n2751 ) ;
  assign n2753 = n752 & n2752 ;
  assign n2754 = n752 & ~n2753 ;
  assign n2755 = ( n2752 & ~n2753 ) | ( n2752 & n2754 ) | ( ~n2753 & n2754 ) ;
  assign n2756 = n2745 & n2755 ;
  assign n2757 = n2745 | n2755 ;
  assign n2758 = ~n2756 & n2757 ;
  assign n2759 = n2435 & n2669 ;
  assign n2760 = n752 & ~n2759 ;
  assign n2761 = n2494 & n2686 ;
  assign n2762 = n2435 & n2673 ;
  assign n2763 = n2433 & n2682 ;
  assign n2764 = n2762 | n2763 ;
  assign n2765 = n2761 | n2764 ;
  assign n2766 = ~n752 & n2765 ;
  assign n2767 = n752 & ~n2765 ;
  assign n2768 = ( n2760 & n2766 ) | ( n2760 & n2767 ) | ( n2766 & n2767 ) ;
  assign n2769 = ~n2425 & n2682 ;
  assign n2770 = n2435 & n2679 ;
  assign n2771 = n2433 & n2673 ;
  assign n2772 = n2770 | n2771 ;
  assign n2773 = n2769 | n2772 ;
  assign n2774 = n2510 & ~n2773 ;
  assign n2775 = n2686 | n2772 ;
  assign n2776 = ( n2769 & ~n2774 ) | ( n2769 & n2775 ) | ( ~n2774 & n2775 ) ;
  assign n2777 = ( ~n752 & n2774 ) | ( ~n752 & n2776 ) | ( n2774 & n2776 ) ;
  assign n2778 = n2776 & ~n2777 ;
  assign n2779 = ~n2774 & n2777 ;
  assign n2780 = ( n752 & ~n2778 ) | ( n752 & n2779 ) | ( ~n2778 & n2779 ) ;
  assign n2781 = n2768 & n2780 ;
  assign n2782 = n2629 & n2781 ;
  assign n2783 = n2781 & ~n2782 ;
  assign n2784 = n2629 & ~n2781 ;
  assign n2785 = n2783 | n2784 ;
  assign n2786 = ~n2425 & n2673 ;
  assign n2787 = n2433 & n2679 ;
  assign n2788 = n2682 | n2787 ;
  assign n2789 = ( n2422 & n2787 ) | ( n2422 & n2788 ) | ( n2787 & n2788 ) ;
  assign n2790 = n2786 | n2789 ;
  assign n2791 = n752 & ~n2692 ;
  assign n2792 = ( n752 & n2530 ) | ( n752 & n2791 ) | ( n2530 & n2791 ) ;
  assign n2793 = ~n2790 & n2792 ;
  assign n2794 = n2686 | n2790 ;
  assign n2795 = ( ~n2530 & n2790 ) | ( ~n2530 & n2794 ) | ( n2790 & n2794 ) ;
  assign n2796 = ~n752 & n2795 ;
  assign n2797 = n2793 | n2796 ;
  assign n2798 = n2785 & ~n2797 ;
  assign n2799 = ( n2782 & n2785 ) | ( n2782 & ~n2798 ) | ( n2785 & ~n2798 ) ;
  assign n2800 = n2758 & n2799 ;
  assign n2801 = n2756 | n2800 ;
  assign n2802 = ( n2732 & ~n2742 ) | ( n2732 & n2801 ) | ( ~n2742 & n2801 ) ;
  assign n2803 = ( ~n2732 & n2742 ) | ( ~n2732 & n2802 ) | ( n2742 & n2802 ) ;
  assign n2804 = ( ~n2801 & n2802 ) | ( ~n2801 & n2803 ) | ( n2802 & n2803 ) ;
  assign n2805 = ( n2743 & n2801 ) | ( n2743 & ~n2804 ) | ( n2801 & ~n2804 ) ;
  assign n2806 = n2730 & n2805 ;
  assign n2807 = n2728 | n2806 ;
  assign n2808 = ( n2713 & n2715 ) | ( n2713 & n2807 ) | ( n2715 & n2807 ) ;
  assign n2809 = n2393 & ~n2398 ;
  assign n2810 = n2399 | n2809 ;
  assign n2811 = ~n2445 & n2810 ;
  assign n2812 = ~n2448 & n2811 ;
  assign n2813 = ( n2445 & n2448 ) | ( n2445 & ~n2810 ) | ( n2448 & ~n2810 ) ;
  assign n2814 = n2812 | n2813 ;
  assign n2815 = ~n2398 & n2673 ;
  assign n2816 = n2403 & n2679 ;
  assign n2817 = n2815 | n2816 ;
  assign n2818 = ( n2393 & n2669 ) | ( n2393 & n2686 ) | ( n2669 & n2686 ) ;
  assign n2819 = n2817 | n2818 ;
  assign n2820 = ( ~n2677 & n2817 ) | ( ~n2677 & n2819 ) | ( n2817 & n2819 ) ;
  assign n2821 = ( ~n2814 & n2819 ) | ( ~n2814 & n2820 ) | ( n2819 & n2820 ) ;
  assign n2822 = ~n752 & n2821 ;
  assign n2823 = n752 | n2822 ;
  assign n2824 = ( ~n2821 & n2822 ) | ( ~n2821 & n2823 ) | ( n2822 & n2823 ) ;
  assign n2825 = ( n2700 & n2808 ) | ( n2700 & n2824 ) | ( n2808 & n2824 ) ;
  assign n2826 = n2698 & n2825 ;
  assign n2827 = n2696 | n2826 ;
  assign n2828 = n2403 & n2559 ;
  assign n2829 = ( n2405 & n2409 ) | ( n2405 & n2557 ) | ( n2409 & n2557 ) ;
  assign n2830 = n2828 | n2829 ;
  assign n2831 = ~n2398 & n2563 ;
  assign n2832 = n2562 | n2831 ;
  assign n2833 = n2830 | n2832 ;
  assign n2834 = n977 & n2833 ;
  assign n2835 = n977 & n2831 ;
  assign n2836 = ( n977 & n2830 ) | ( n977 & n2835 ) | ( n2830 & n2835 ) ;
  assign n2837 = ( ~n2708 & n2834 ) | ( ~n2708 & n2836 ) | ( n2834 & n2836 ) ;
  assign n2838 = n977 | n2833 ;
  assign n2839 = n977 | n2831 ;
  assign n2840 = n2830 | n2839 ;
  assign n2841 = ( ~n2708 & n2838 ) | ( ~n2708 & n2840 ) | ( n2838 & n2840 ) ;
  assign n2842 = ~n2837 & n2841 ;
  assign n2843 = ( n2485 & n2524 ) | ( n2485 & n2540 ) | ( n2524 & n2540 ) ;
  assign n2844 = n2422 & n2499 ;
  assign n2845 = n2415 & n2501 ;
  assign n2846 = n2844 | n2845 ;
  assign n2847 = ~n2425 & n2512 ;
  assign n2848 = n2491 | n2847 ;
  assign n2849 = n2846 | n2848 ;
  assign n2850 = n566 | n2849 ;
  assign n2851 = n566 | n2847 ;
  assign n2852 = n2846 | n2851 ;
  assign n2853 = ( n2608 & n2850 ) | ( n2608 & n2852 ) | ( n2850 & n2852 ) ;
  assign n2854 = n566 & n2847 ;
  assign n2855 = ( n566 & n2846 ) | ( n566 & n2854 ) | ( n2846 & n2854 ) ;
  assign n2856 = ( n2608 & n2849 ) | ( n2608 & n2855 ) | ( n2849 & n2855 ) ;
  assign n2857 = ( n566 & n2854 ) | ( n566 & n2856 ) | ( n2854 & n2856 ) ;
  assign n2858 = n2853 & ~n2857 ;
  assign n2859 = n566 & n2433 ;
  assign n2860 = ~n2856 & n2859 ;
  assign n2861 = n2859 & ~n2860 ;
  assign n2862 = ( n2858 & ~n2860 ) | ( n2858 & n2861 ) | ( ~n2860 & n2861 ) ;
  assign n2863 = n2843 & n2862 ;
  assign n2864 = n2862 & ~n2863 ;
  assign n2865 = ( n2843 & ~n2863 ) | ( n2843 & n2864 ) | ( ~n2863 & n2864 ) ;
  assign n2866 = n2842 & n2865 ;
  assign n2867 = n2865 & ~n2866 ;
  assign n2868 = ( n2842 & ~n2866 ) | ( n2842 & n2867 ) | ( ~n2866 & n2867 ) ;
  assign n2869 = n2576 | n2665 ;
  assign n2870 = ~n2868 & n2869 ;
  assign n2871 = n2868 & ~n2869 ;
  assign n2872 = n2870 | n2871 ;
  assign n2873 = n2393 & n2679 ;
  assign n2874 = ( n2452 & n2456 ) | ( n2452 & n2673 ) | ( n2456 & n2673 ) ;
  assign n2875 = n2873 | n2874 ;
  assign n2876 = ( n2461 & n2669 ) | ( n2461 & n2686 ) | ( n2669 & n2686 ) ;
  assign n2877 = n2875 | n2876 ;
  assign n2878 = ( n2682 & n2875 ) | ( n2682 & n2877 ) | ( n2875 & n2877 ) ;
  assign n2879 = ( n2450 & n2463 ) | ( n2450 & n2465 ) | ( n2463 & n2465 ) ;
  assign n2880 = ( n2457 & ~n2461 ) | ( n2457 & n2879 ) | ( ~n2461 & n2879 ) ;
  assign n2881 = ( ~n2457 & n2461 ) | ( ~n2457 & n2880 ) | ( n2461 & n2880 ) ;
  assign n2882 = ( ~n2879 & n2880 ) | ( ~n2879 & n2881 ) | ( n2880 & n2881 ) ;
  assign n2883 = ( n2877 & n2878 ) | ( n2877 & n2882 ) | ( n2878 & n2882 ) ;
  assign n2884 = n752 & n2883 ;
  assign n2885 = n752 & ~n2884 ;
  assign n2886 = ( n2883 & ~n2884 ) | ( n2883 & n2885 ) | ( ~n2884 & n2885 ) ;
  assign n2887 = n2872 & n2886 ;
  assign n2888 = n2872 | n2886 ;
  assign n2889 = ~n2887 & n2888 ;
  assign n2890 = n2827 & n2889 ;
  assign n2891 = n2827 | n2889 ;
  assign n2892 = ~n2890 & n2891 ;
  assign n2893 = n2484 & n2892 ;
  assign n2894 = n2484 | n2892 ;
  assign n2895 = ~n2893 & n2894 ;
  assign n2896 = n2381 & n2461 ;
  assign n2897 = ( n2378 & ~n2383 ) | ( n2378 & n2384 ) | ( ~n2383 & n2384 ) ;
  assign n2898 = n2896 | n2897 ;
  assign n2899 = n2366 & n2374 ;
  assign n2900 = n2388 | n2899 ;
  assign n2901 = n2898 | n2900 ;
  assign n2902 = n32 & n2901 ;
  assign n2903 = n32 & n2899 ;
  assign n2904 = ( n32 & n2898 ) | ( n32 & n2903 ) | ( n2898 & n2903 ) ;
  assign n2905 = ( n2467 & ~n2469 ) | ( n2467 & n2473 ) | ( ~n2469 & n2473 ) ;
  assign n2906 = ( n2374 & ~n2468 ) | ( n2374 & n2905 ) | ( ~n2468 & n2905 ) ;
  assign n2907 = ( ~n2374 & n2468 ) | ( ~n2374 & n2906 ) | ( n2468 & n2906 ) ;
  assign n2908 = ( ~n2905 & n2906 ) | ( ~n2905 & n2907 ) | ( n2906 & n2907 ) ;
  assign n2909 = ( n2902 & n2904 ) | ( n2902 & ~n2908 ) | ( n2904 & ~n2908 ) ;
  assign n2910 = n32 | n2901 ;
  assign n2911 = n32 | n2899 ;
  assign n2912 = n2898 | n2911 ;
  assign n2913 = ( ~n2908 & n2910 ) | ( ~n2908 & n2912 ) | ( n2910 & n2912 ) ;
  assign n2914 = ~n2909 & n2913 ;
  assign n2915 = n2698 & ~n2826 ;
  assign n2916 = ( n2825 & ~n2826 ) | ( n2825 & n2915 ) | ( ~n2826 & n2915 ) ;
  assign n2917 = n2914 & n2916 ;
  assign n2918 = n2916 & ~n2917 ;
  assign n2919 = n2914 & ~n2916 ;
  assign n2920 = n2918 | n2919 ;
  assign n2921 = n2469 | n2473 ;
  assign n2922 = n2467 & ~n2921 ;
  assign n2923 = ~n2467 & n2921 ;
  assign n2924 = n2922 | n2923 ;
  assign n2925 = n2378 & n2461 ;
  assign n2926 = ( n2381 & n2452 ) | ( n2381 & n2456 ) | ( n2452 & n2456 ) ;
  assign n2927 = n2925 | n2926 ;
  assign n2928 = ( n2366 & ~n2383 ) | ( n2366 & n2384 ) | ( ~n2383 & n2384 ) ;
  assign n2929 = n2388 | n2928 ;
  assign n2930 = n2927 | n2929 ;
  assign n2931 = n32 & n2930 ;
  assign n2932 = n32 & n2928 ;
  assign n2933 = ( n32 & n2927 ) | ( n32 & n2932 ) | ( n2927 & n2932 ) ;
  assign n2934 = ( ~n2924 & n2931 ) | ( ~n2924 & n2933 ) | ( n2931 & n2933 ) ;
  assign n2935 = n32 | n2930 ;
  assign n2936 = n32 | n2928 ;
  assign n2937 = n2927 | n2936 ;
  assign n2938 = ( ~n2924 & n2935 ) | ( ~n2924 & n2937 ) | ( n2935 & n2937 ) ;
  assign n2939 = ~n2934 & n2938 ;
  assign n2940 = n2378 & n2393 ;
  assign n2941 = n2381 & ~n2398 ;
  assign n2942 = n2940 | n2941 ;
  assign n2943 = ( n2366 & n2452 ) | ( n2366 & n2456 ) | ( n2452 & n2456 ) ;
  assign n2944 = n2942 | n2943 ;
  assign n2945 = ( n2388 & n2689 ) | ( n2388 & n2944 ) | ( n2689 & n2944 ) ;
  assign n2946 = ( n32 & ~n2944 ) | ( n32 & n2945 ) | ( ~n2944 & n2945 ) ;
  assign n2947 = ~n2945 & n2946 ;
  assign n2948 = n2944 | n2946 ;
  assign n2949 = ( ~n32 & n2947 ) | ( ~n32 & n2948 ) | ( n2947 & n2948 ) ;
  assign n2950 = n2378 & ~n2398 ;
  assign n2951 = n2381 & n2403 ;
  assign n2952 = n2950 | n2951 ;
  assign n2953 = ( n2365 & n2388 ) | ( n2365 & n2393 ) | ( n2388 & n2393 ) ;
  assign n2954 = n2952 | n2953 ;
  assign n2955 = ( ~n2357 & n2952 ) | ( ~n2357 & n2954 ) | ( n2952 & n2954 ) ;
  assign n2956 = ( ~n2814 & n2954 ) | ( ~n2814 & n2955 ) | ( n2954 & n2955 ) ;
  assign n2957 = ~n32 & n2956 ;
  assign n2958 = n32 | n2957 ;
  assign n2959 = ( ~n2956 & n2957 ) | ( ~n2956 & n2958 ) | ( n2957 & n2958 ) ;
  assign n2960 = n2378 & n2403 ;
  assign n2961 = ( n2381 & n2405 ) | ( n2381 & n2409 ) | ( n2405 & n2409 ) ;
  assign n2962 = n2960 | n2961 ;
  assign n2963 = n2366 & ~n2398 ;
  assign n2964 = n2388 | n2963 ;
  assign n2965 = n2962 | n2964 ;
  assign n2966 = n32 & n2965 ;
  assign n2967 = n32 & n2963 ;
  assign n2968 = ( n32 & n2962 ) | ( n32 & n2967 ) | ( n2962 & n2967 ) ;
  assign n2969 = ( ~n2708 & n2966 ) | ( ~n2708 & n2968 ) | ( n2966 & n2968 ) ;
  assign n2970 = n32 | n2965 ;
  assign n2971 = n32 | n2963 ;
  assign n2972 = n2962 | n2971 ;
  assign n2973 = ( ~n2708 & n2970 ) | ( ~n2708 & n2972 ) | ( n2970 & n2972 ) ;
  assign n2974 = ~n2969 & n2973 ;
  assign n2975 = n2758 | n2799 ;
  assign n2976 = ~n2800 & n2975 ;
  assign n2977 = n2974 | n2976 ;
  assign n2978 = ~n2785 & n2797 ;
  assign n2979 = n2798 | n2978 ;
  assign n2980 = n2381 & n2415 ;
  assign n2981 = ( n2378 & n2405 ) | ( n2378 & n2409 ) | ( n2405 & n2409 ) ;
  assign n2982 = n2980 | n2981 ;
  assign n2983 = n2366 & n2403 ;
  assign n2984 = n2982 | n2983 ;
  assign n2985 = n2388 | n2984 ;
  assign n2986 = ( n2546 & n2984 ) | ( n2546 & n2985 ) | ( n2984 & n2985 ) ;
  assign n2987 = n32 & n2986 ;
  assign n2988 = n32 & ~n2987 ;
  assign n2989 = ( n2986 & ~n2987 ) | ( n2986 & n2988 ) | ( ~n2987 & n2988 ) ;
  assign n2990 = n2979 & n2989 ;
  assign n2991 = n2979 | n2989 ;
  assign n2992 = ~n2990 & n2991 ;
  assign n2993 = n2381 & n2422 ;
  assign n2994 = n2378 & n2415 ;
  assign n2995 = n2993 | n2994 ;
  assign n2996 = ( n2366 & n2405 ) | ( n2366 & n2409 ) | ( n2405 & n2409 ) ;
  assign n2997 = n2995 | n2996 ;
  assign n2998 = n2389 & n2585 ;
  assign n2999 = ( n32 & n2997 ) | ( n32 & n2998 ) | ( n2997 & n2998 ) ;
  assign n3000 = ( n32 & n2481 ) | ( n32 & n2585 ) | ( n2481 & n2585 ) ;
  assign n3001 = n2997 | n3000 ;
  assign n3002 = ~n2999 & n3001 ;
  assign n3003 = n2768 | n2780 ;
  assign n3004 = ~n2781 & n3003 ;
  assign n3005 = n3002 & n3004 ;
  assign n3006 = n3002 | n3004 ;
  assign n3007 = ~n3005 & n3006 ;
  assign n3008 = n2760 | n2767 ;
  assign n3009 = n2766 | n3008 ;
  assign n3010 = ~n2768 & n3009 ;
  assign n3011 = n2366 & ~n2425 ;
  assign n3012 = n2381 & n2435 ;
  assign n3013 = n2378 & n2433 ;
  assign n3014 = n3012 | n3013 ;
  assign n3015 = n3011 | n3014 ;
  assign n3016 = n2510 & ~n3015 ;
  assign n3017 = n2388 | n3014 ;
  assign n3018 = ( n3011 & ~n3016 ) | ( n3011 & n3017 ) | ( ~n3016 & n3017 ) ;
  assign n3019 = ( ~n32 & n3016 ) | ( ~n32 & n3018 ) | ( n3016 & n3018 ) ;
  assign n3020 = n3018 & ~n3019 ;
  assign n3021 = ~n3016 & n3019 ;
  assign n3022 = ( n32 & ~n3020 ) | ( n32 & n3021 ) | ( ~n3020 & n3021 ) ;
  assign n3023 = n2365 & n2435 ;
  assign n3024 = n32 & ~n3023 ;
  assign n3025 = n2388 & n2494 ;
  assign n3026 = n2378 & n2435 ;
  assign n3027 = n3025 | n3026 ;
  assign n3028 = n2366 & n2433 ;
  assign n3029 = ~n3027 & n3028 ;
  assign n3030 = ( n32 & ~n3027 ) | ( n32 & n3029 ) | ( ~n3027 & n3029 ) ;
  assign n3031 = ( n32 & n3029 ) | ( n32 & ~n3030 ) | ( n3029 & ~n3030 ) ;
  assign n3032 = ( n3027 & n3030 ) | ( n3027 & ~n3031 ) | ( n3030 & ~n3031 ) ;
  assign n3033 = n3024 & n3032 ;
  assign n3034 = n2759 & n3033 ;
  assign n3035 = n3022 & n3034 ;
  assign n3036 = n2378 & ~n2425 ;
  assign n3037 = n2381 & n2433 ;
  assign n3038 = n2366 | n3037 ;
  assign n3039 = ( n2422 & n3037 ) | ( n2422 & n3038 ) | ( n3037 & n3038 ) ;
  assign n3040 = n3036 | n3039 ;
  assign n3041 = n2389 & ~n2530 ;
  assign n3042 = ( n32 & n3040 ) | ( n32 & n3041 ) | ( n3040 & n3041 ) ;
  assign n3043 = ( n32 & n2481 ) | ( n32 & ~n2530 ) | ( n2481 & ~n2530 ) ;
  assign n3044 = n3040 | n3043 ;
  assign n3045 = ~n3042 & n3044 ;
  assign n3046 = n3022 & n3033 ;
  assign n3047 = n2759 | n3046 ;
  assign n3048 = ~n3035 & n3047 ;
  assign n3049 = n3045 & n3048 ;
  assign n3050 = n3035 | n3049 ;
  assign n3051 = n2378 & n2422 ;
  assign n3052 = n2366 & n2415 ;
  assign n3053 = n3051 | n3052 ;
  assign n3054 = n2381 & ~n2425 ;
  assign n3055 = n3053 | n3054 ;
  assign n3056 = n2388 | n3055 ;
  assign n3057 = ( n2608 & n3055 ) | ( n2608 & n3056 ) | ( n3055 & n3056 ) ;
  assign n3058 = n32 & n3057 ;
  assign n3059 = n32 & ~n3058 ;
  assign n3060 = ( n3057 & ~n3058 ) | ( n3057 & n3059 ) | ( ~n3058 & n3059 ) ;
  assign n3061 = ( n3010 & n3050 ) | ( n3010 & n3060 ) | ( n3050 & n3060 ) ;
  assign n3062 = n3007 & n3061 ;
  assign n3063 = n3005 | n3062 ;
  assign n3064 = n2992 & n3063 ;
  assign n3065 = n2990 | n3064 ;
  assign n3066 = ( n2974 & ~n2976 ) | ( n2974 & n3065 ) | ( ~n2976 & n3065 ) ;
  assign n3067 = ( ~n2974 & n2976 ) | ( ~n2974 & n3066 ) | ( n2976 & n3066 ) ;
  assign n3068 = ( ~n3065 & n3066 ) | ( ~n3065 & n3067 ) | ( n3066 & n3067 ) ;
  assign n3069 = ( n2977 & n3065 ) | ( n2977 & ~n3068 ) | ( n3065 & ~n3068 ) ;
  assign n3070 = ( n2804 & n2959 ) | ( n2804 & n3069 ) | ( n2959 & n3069 ) ;
  assign n3071 = n2805 & ~n2806 ;
  assign n3072 = ( n2730 & ~n2806 ) | ( n2730 & n3071 ) | ( ~n2806 & n3071 ) ;
  assign n3073 = ( n2949 & n3070 ) | ( n2949 & n3072 ) | ( n3070 & n3072 ) ;
  assign n3074 = ( n2713 & ~n2715 ) | ( n2713 & n2807 ) | ( ~n2715 & n2807 ) ;
  assign n3075 = ( ~n2713 & n2715 ) | ( ~n2713 & n3074 ) | ( n2715 & n3074 ) ;
  assign n3076 = ( ~n2807 & n3074 ) | ( ~n2807 & n3075 ) | ( n3074 & n3075 ) ;
  assign n3077 = n2381 & n2393 ;
  assign n3078 = ( n2378 & n2452 ) | ( n2378 & n2456 ) | ( n2452 & n2456 ) ;
  assign n3079 = n3077 | n3078 ;
  assign n3080 = ( n2365 & n2388 ) | ( n2365 & n2461 ) | ( n2388 & n2461 ) ;
  assign n3081 = n3079 | n3080 ;
  assign n3082 = ( n2366 & n3079 ) | ( n2366 & n3081 ) | ( n3079 & n3081 ) ;
  assign n3083 = ( n2882 & n3081 ) | ( n2882 & n3082 ) | ( n3081 & n3082 ) ;
  assign n3084 = n32 & n3083 ;
  assign n3085 = n32 & ~n3084 ;
  assign n3086 = ( n3083 & ~n3084 ) | ( n3083 & n3085 ) | ( ~n3084 & n3085 ) ;
  assign n3087 = ( n3073 & n3076 ) | ( n3073 & n3086 ) | ( n3076 & n3086 ) ;
  assign n3088 = ~n2700 & n2824 ;
  assign n3089 = n2700 & ~n2824 ;
  assign n3090 = n3088 | n3089 ;
  assign n3091 = ( n2808 & n2939 ) | ( n2808 & ~n3090 ) | ( n2939 & ~n3090 ) ;
  assign n3092 = ( ~n2808 & n3090 ) | ( ~n2808 & n3091 ) | ( n3090 & n3091 ) ;
  assign n3093 = ( ~n2939 & n3091 ) | ( ~n2939 & n3092 ) | ( n3091 & n3092 ) ;
  assign n3094 = n3087 & n3093 ;
  assign n3095 = n3087 | n3093 ;
  assign n3096 = ~n3094 & n3095 ;
  assign n3097 = ( n2939 & n3087 ) | ( n2939 & ~n3096 ) | ( n3087 & ~n3096 ) ;
  assign n3098 = n2920 & n3097 ;
  assign n3099 = n2917 | n3098 ;
  assign n3100 = n2895 & n3099 ;
  assign n3101 = n2895 | n3099 ;
  assign n3102 = ~n3100 & n3101 ;
  assign n3103 = n232 | n481 ;
  assign n3104 = n577 | n3103 ;
  assign n3105 = n449 & ~n465 ;
  assign n3106 = ~n330 & n3105 ;
  assign n3107 = ~n2012 & n3106 ;
  assign n3108 = ~n328 & n3107 ;
  assign n3109 = n256 | n900 ;
  assign n3110 = n157 | n3109 ;
  assign n3111 = n2151 | n2241 ;
  assign n3112 = n3110 | n3111 ;
  assign n3113 = n3108 & ~n3112 ;
  assign n3114 = ~n379 & n3113 ;
  assign n3115 = ~n3104 & n3114 ;
  assign n3116 = ~n2351 & n3115 ;
  assign n3117 = n2317 & n3116 ;
  assign n3118 = ( n2317 & ~n2353 ) | ( n2317 & n3115 ) | ( ~n2353 & n3115 ) ;
  assign n3119 = ~n3117 & n3118 ;
  assign n3120 = x1 & ~n430 ;
  assign n3121 = ~x1 & n430 ;
  assign n3122 = n3120 | n3121 ;
  assign n3123 = n2362 & ~n3122 ;
  assign n3124 = ~n2362 & n3122 ;
  assign n3125 = n3123 | n3124 ;
  assign n3126 = ~n2359 & n3125 ;
  assign n3127 = ~n3119 & n3126 ;
  assign n3128 = ~x0 & n3122 ;
  assign n3129 = n310 | n311 ;
  assign n3130 = n327 | n330 ;
  assign n3131 = n324 | n3130 ;
  assign n3132 = n3129 | n3131 ;
  assign n3133 = n276 | n370 ;
  assign n3134 = n1016 | n3133 ;
  assign n3135 = n366 | n3134 ;
  assign n3136 = n206 | n403 ;
  assign n3137 = n402 | n3136 ;
  assign n3138 = n385 | n3137 ;
  assign n3139 = n3135 | n3138 ;
  assign n3140 = n3132 | n3139 ;
  assign n3141 = n253 | n355 ;
  assign n3142 = n181 | n3141 ;
  assign n3143 = n287 | n3142 ;
  assign n3144 = n3140 | n3143 ;
  assign n3145 = n3117 & n3144 ;
  assign n3146 = n3144 & ~n3145 ;
  assign n3147 = ( n3117 & ~n3145 ) | ( n3117 & n3146 ) | ( ~n3145 & n3146 ) ;
  assign n3148 = n3128 & n3147 ;
  assign n3149 = n3127 | n3148 ;
  assign n3150 = n133 | n311 ;
  assign n3151 = n186 | n3150 ;
  assign n3152 = n310 | n3151 ;
  assign n3153 = n302 | n3152 ;
  assign n3154 = n3131 | n3153 ;
  assign n3155 = n358 | n396 ;
  assign n3156 = n359 | n3155 ;
  assign n3157 = n3154 | n3156 ;
  assign n3158 = n249 | n267 ;
  assign n3159 = n3157 | n3158 ;
  assign n3160 = ( n3117 & n3145 ) | ( n3117 & n3159 ) | ( n3145 & n3159 ) ;
  assign n3161 = ( n3145 & n3159 ) | ( n3145 & ~n3160 ) | ( n3159 & ~n3160 ) ;
  assign n3162 = ( n3117 & ~n3160 ) | ( n3117 & n3161 ) | ( ~n3160 & n3161 ) ;
  assign n3163 = x0 & n3125 ;
  assign n3164 = ( x0 & n3162 ) | ( x0 & n3163 ) | ( n3162 & n3163 ) ;
  assign n3165 = n3149 | n3164 ;
  assign n3166 = x0 & ~n3125 ;
  assign n3167 = ( n3149 & n3165 ) | ( n3149 & n3166 ) | ( n3165 & n3166 ) ;
  assign n3168 = ~n3119 & n3147 ;
  assign n3169 = n3119 & ~n3147 ;
  assign n3170 = n2354 & ~n3119 ;
  assign n3171 = n2354 | n2374 ;
  assign n3172 = ~n2354 & n3119 ;
  assign n3173 = n3170 | n3172 ;
  assign n3174 = n3171 & ~n3173 ;
  assign n3175 = n2354 & n2374 ;
  assign n3176 = ~n3173 & n3175 ;
  assign n3177 = ( n2475 & n3174 ) | ( n2475 & n3176 ) | ( n3174 & n3176 ) ;
  assign n3178 = n3170 | n3177 ;
  assign n3179 = ( n3168 & ~n3169 ) | ( n3168 & n3178 ) | ( ~n3169 & n3178 ) ;
  assign n3180 = ( n3147 & ~n3162 ) | ( n3147 & n3179 ) | ( ~n3162 & n3179 ) ;
  assign n3181 = ( ~n3147 & n3162 ) | ( ~n3147 & n3180 ) | ( n3162 & n3180 ) ;
  assign n3182 = ( ~n3179 & n3180 ) | ( ~n3179 & n3181 ) | ( n3180 & n3181 ) ;
  assign n3183 = ( n3165 & n3167 ) | ( n3165 & n3182 ) | ( n3167 & n3182 ) ;
  assign n3184 = n2362 & n3183 ;
  assign n3185 = n2362 & ~n3184 ;
  assign n3186 = ( n3183 & ~n3184 ) | ( n3183 & n3185 ) | ( ~n3184 & n3185 ) ;
  assign n3187 = n3102 & n3186 ;
  assign n3188 = n3102 | n3186 ;
  assign n3189 = ~n3187 & n3188 ;
  assign n3190 = n2920 | n3097 ;
  assign n3191 = ~n3098 & n3190 ;
  assign n3192 = ~n3171 & n3173 ;
  assign n3193 = n3173 & ~n3175 ;
  assign n3194 = ( n2471 & n3192 ) | ( n2471 & n3193 ) | ( n3192 & n3193 ) ;
  assign n3195 = ( ~n2474 & n3192 ) | ( ~n2474 & n3193 ) | ( n3192 & n3193 ) ;
  assign n3196 = ( ~n2467 & n3194 ) | ( ~n2467 & n3195 ) | ( n3194 & n3195 ) ;
  assign n3197 = n3177 | n3196 ;
  assign n3198 = n2374 & n3126 ;
  assign n3199 = n2354 & n3128 ;
  assign n3200 = n3198 | n3199 ;
  assign n3201 = ( x0 & ~n3119 ) | ( x0 & n3163 ) | ( ~n3119 & n3163 ) ;
  assign n3202 = n3200 | n3201 ;
  assign n3203 = ( n3166 & n3200 ) | ( n3166 & n3202 ) | ( n3200 & n3202 ) ;
  assign n3204 = ( ~n3197 & n3202 ) | ( ~n3197 & n3203 ) | ( n3202 & n3203 ) ;
  assign n3205 = ~n2362 & n3204 ;
  assign n3206 = n2362 | n3205 ;
  assign n3207 = ( ~n3204 & n3205 ) | ( ~n3204 & n3206 ) | ( n3205 & n3206 ) ;
  assign n3208 = n3096 & n3207 ;
  assign n3209 = n3096 & ~n3208 ;
  assign n3210 = ( n3207 & ~n3208 ) | ( n3207 & n3209 ) | ( ~n3208 & n3209 ) ;
  assign n3211 = n2461 & n3126 ;
  assign n3212 = ( ~n2383 & n2384 ) | ( ~n2383 & n3128 ) | ( n2384 & n3128 ) ;
  assign n3213 = n3211 | n3212 ;
  assign n3214 = n2374 & n3166 ;
  assign n3215 = n3163 | n3214 ;
  assign n3216 = n3213 | n3215 ;
  assign n3217 = n2362 & n3216 ;
  assign n3218 = n2362 & n3214 ;
  assign n3219 = ( n2362 & n3213 ) | ( n2362 & n3218 ) | ( n3213 & n3218 ) ;
  assign n3220 = ( ~n2908 & n3217 ) | ( ~n2908 & n3219 ) | ( n3217 & n3219 ) ;
  assign n3221 = n2362 | n3216 ;
  assign n3222 = n2362 | n3214 ;
  assign n3223 = n3213 | n3222 ;
  assign n3224 = ( ~n2908 & n3221 ) | ( ~n2908 & n3223 ) | ( n3221 & n3223 ) ;
  assign n3225 = ~n3220 & n3224 ;
  assign n3226 = n2461 & n3128 ;
  assign n3227 = ( n2452 & n2456 ) | ( n2452 & n3126 ) | ( n2456 & n3126 ) ;
  assign n3228 = n3226 | n3227 ;
  assign n3229 = ( ~n2383 & n2384 ) | ( ~n2383 & n3166 ) | ( n2384 & n3166 ) ;
  assign n3230 = n3163 | n3229 ;
  assign n3231 = n3228 | n3230 ;
  assign n3232 = ~n2362 & n3231 ;
  assign n3233 = ~n2362 & n3229 ;
  assign n3234 = ( ~n2362 & n3228 ) | ( ~n2362 & n3233 ) | ( n3228 & n3233 ) ;
  assign n3235 = ( ~n2924 & n3232 ) | ( ~n2924 & n3234 ) | ( n3232 & n3234 ) ;
  assign n3236 = n2362 & ~n3231 ;
  assign n3237 = n2362 & ~n3229 ;
  assign n3238 = ~n3228 & n3237 ;
  assign n3239 = ( n2924 & n3236 ) | ( n2924 & n3238 ) | ( n3236 & n3238 ) ;
  assign n3240 = n3235 | n3239 ;
  assign n3241 = n3007 | n3061 ;
  assign n3242 = ~n3062 & n3241 ;
  assign n3243 = n2422 & n3126 ;
  assign n3244 = n2415 & n3128 ;
  assign n3245 = n3243 | n3244 ;
  assign n3246 = ( n2405 & n2409 ) | ( n2405 & n3166 ) | ( n2409 & n3166 ) ;
  assign n3247 = n3245 | n3246 ;
  assign n3248 = n3163 | n3247 ;
  assign n3249 = ( n2585 & n3247 ) | ( n2585 & n3248 ) | ( n3247 & n3248 ) ;
  assign n3250 = ( x0 & n3123 ) | ( x0 & n3128 ) | ( n3123 & n3128 ) ;
  assign n3251 = n2585 & n3250 ;
  assign n3252 = ( n2362 & n3247 ) | ( n2362 & n3251 ) | ( n3247 & n3251 ) ;
  assign n3253 = n3249 & ~n3252 ;
  assign n3254 = n2362 & ~n3250 ;
  assign n3255 = ( n2362 & ~n2585 ) | ( n2362 & n3254 ) | ( ~n2585 & n3254 ) ;
  assign n3256 = ~n3247 & n3255 ;
  assign n3257 = n3253 | n3256 ;
  assign n3258 = n3024 | n3032 ;
  assign n3259 = ~n3033 & n3258 ;
  assign n3260 = ~n2425 & n3128 ;
  assign n3261 = n2433 & n3126 ;
  assign n3262 = n3166 | n3261 ;
  assign n3263 = ( n2422 & n3261 ) | ( n2422 & n3262 ) | ( n3261 & n3262 ) ;
  assign n3264 = n3260 | n3263 ;
  assign n3265 = ~n2530 & n3250 ;
  assign n3266 = ( n2362 & n3264 ) | ( n2362 & n3265 ) | ( n3264 & n3265 ) ;
  assign n3267 = n2362 | n3163 ;
  assign n3268 = ( n2362 & ~n2530 ) | ( n2362 & n3267 ) | ( ~n2530 & n3267 ) ;
  assign n3269 = n3264 | n3268 ;
  assign n3270 = ~n3266 & n3269 ;
  assign n3271 = ~n2510 & n3250 ;
  assign n3272 = n2494 & n3250 ;
  assign n3273 = n2362 & ~n3128 ;
  assign n3274 = ( n2362 & ~n2435 ) | ( n2362 & n3273 ) | ( ~n2435 & n3273 ) ;
  assign n3275 = n2433 & n3166 ;
  assign n3276 = n3274 & ~n3275 ;
  assign n3277 = ~n3272 & n3276 ;
  assign n3278 = ~n2425 & n3166 ;
  assign n3279 = n2433 & n3128 ;
  assign n3280 = n2435 & n3126 ;
  assign n3281 = ( n2362 & n3279 ) | ( n2362 & n3280 ) | ( n3279 & n3280 ) ;
  assign n3282 = ( n2362 & n3278 ) | ( n2362 & n3281 ) | ( n3278 & n3281 ) ;
  assign n3283 = n3277 & ~n3282 ;
  assign n3284 = ~n3271 & n3283 ;
  assign n3285 = x0 & n2435 ;
  assign n3286 = n3284 & ~n3285 ;
  assign n3287 = ( n3023 & n3270 ) | ( n3023 & n3286 ) | ( n3270 & n3286 ) ;
  assign n3288 = n2608 & n3250 ;
  assign n3289 = n2422 & n3128 ;
  assign n3290 = n2415 & n3166 ;
  assign n3291 = n3289 | n3290 ;
  assign n3292 = ~n2425 & n3126 ;
  assign n3293 = n2362 | n3292 ;
  assign n3294 = n3291 | n3293 ;
  assign n3295 = ( ~n3267 & n3291 ) | ( ~n3267 & n3292 ) | ( n3291 & n3292 ) ;
  assign n3296 = n3267 | n3295 ;
  assign n3297 = ( n2608 & n3294 ) | ( n2608 & n3296 ) | ( n3294 & n3296 ) ;
  assign n3298 = ~n3288 & n3297 ;
  assign n3299 = ( n2362 & n3291 ) | ( n2362 & n3292 ) | ( n3291 & n3292 ) ;
  assign n3300 = n3298 & ~n3299 ;
  assign n3301 = ( n3259 & n3287 ) | ( n3259 & n3300 ) | ( n3287 & n3300 ) ;
  assign n3302 = n3257 & n3301 ;
  assign n3303 = n3048 & ~n3049 ;
  assign n3304 = ( n3045 & ~n3049 ) | ( n3045 & n3303 ) | ( ~n3049 & n3303 ) ;
  assign n3305 = n3302 | n3304 ;
  assign n3306 = n2546 & n3250 ;
  assign n3307 = n2415 & n3126 ;
  assign n3308 = ( n2405 & n2409 ) | ( n2405 & n3128 ) | ( n2409 & n3128 ) ;
  assign n3309 = n3307 | n3308 ;
  assign n3310 = n2403 & n3166 ;
  assign n3311 = n2362 | n3310 ;
  assign n3312 = n3309 | n3311 ;
  assign n3313 = ( ~n3267 & n3309 ) | ( ~n3267 & n3310 ) | ( n3309 & n3310 ) ;
  assign n3314 = n3267 | n3313 ;
  assign n3315 = ( n2546 & n3312 ) | ( n2546 & n3314 ) | ( n3312 & n3314 ) ;
  assign n3316 = ~n3306 & n3315 ;
  assign n3317 = n2362 & n3310 ;
  assign n3318 = ( n2362 & n3309 ) | ( n2362 & n3317 ) | ( n3309 & n3317 ) ;
  assign n3319 = n3316 & ~n3318 ;
  assign n3320 = n3022 | n3033 ;
  assign n3321 = ~n3046 & n3257 ;
  assign n3322 = ( ~n3046 & n3301 ) | ( ~n3046 & n3321 ) | ( n3301 & n3321 ) ;
  assign n3323 = n3320 & n3322 ;
  assign n3324 = n3319 & n3323 ;
  assign n3325 = ( n3305 & n3319 ) | ( n3305 & n3324 ) | ( n3319 & n3324 ) ;
  assign n3326 = n2403 & n3128 ;
  assign n3327 = ( n2405 & n2409 ) | ( n2405 & n3126 ) | ( n2409 & n3126 ) ;
  assign n3328 = n3326 | n3327 ;
  assign n3329 = ~n2398 & n3166 ;
  assign n3330 = n3328 | n3329 ;
  assign n3331 = n3163 | n3330 ;
  assign n3332 = ( ~n2708 & n3330 ) | ( ~n2708 & n3331 ) | ( n3330 & n3331 ) ;
  assign n3333 = ~n2362 & n3332 ;
  assign n3334 = n2362 & ~n3332 ;
  assign n3335 = n3333 | n3334 ;
  assign n3336 = n3302 & n3304 ;
  assign n3337 = ( n3304 & n3323 ) | ( n3304 & n3336 ) | ( n3323 & n3336 ) ;
  assign n3338 = n3335 & n3337 ;
  assign n3339 = ( n3325 & n3335 ) | ( n3325 & n3338 ) | ( n3335 & n3338 ) ;
  assign n3340 = n3242 | n3339 ;
  assign n3341 = n3335 | n3337 ;
  assign n3342 = n3325 | n3341 ;
  assign n3343 = ( ~n3010 & n3050 ) | ( ~n3010 & n3060 ) | ( n3050 & n3060 ) ;
  assign n3344 = ( n3010 & n3050 ) | ( n3010 & ~n3060 ) | ( n3050 & ~n3060 ) ;
  assign n3345 = ( ~n3050 & n3343 ) | ( ~n3050 & n3344 ) | ( n3343 & n3344 ) ;
  assign n3346 = n3342 & n3345 ;
  assign n3347 = n3340 | n3346 ;
  assign n3348 = ~n2398 & n3128 ;
  assign n3349 = n2403 & n3126 ;
  assign n3350 = n3348 | n3349 ;
  assign n3351 = n2362 & n3166 ;
  assign n3352 = n2393 & n3351 ;
  assign n3353 = ( n2362 & n3350 ) | ( n2362 & n3352 ) | ( n3350 & n3352 ) ;
  assign n3354 = ~n2814 & n3250 ;
  assign n3355 = n2393 & n3166 ;
  assign n3356 = n2362 | n3355 ;
  assign n3357 = n3350 | n3356 ;
  assign n3358 = ( ~n3267 & n3350 ) | ( ~n3267 & n3355 ) | ( n3350 & n3355 ) ;
  assign n3359 = n3267 | n3358 ;
  assign n3360 = ( ~n2814 & n3357 ) | ( ~n2814 & n3359 ) | ( n3357 & n3359 ) ;
  assign n3361 = ~n3354 & n3360 ;
  assign n3362 = ~n3353 & n3361 ;
  assign n3363 = n3347 & n3362 ;
  assign n3364 = n2992 & ~n3064 ;
  assign n3365 = ~n2992 & n3063 ;
  assign n3366 = n3364 | n3365 ;
  assign n3367 = n3242 & n3339 ;
  assign n3368 = ( n3242 & n3346 ) | ( n3242 & n3367 ) | ( n3346 & n3367 ) ;
  assign n3369 = n3366 | n3368 ;
  assign n3370 = n3363 | n3369 ;
  assign n3371 = n2393 & n3128 ;
  assign n3372 = ~n2398 & n3126 ;
  assign n3373 = n3371 | n3372 ;
  assign n3374 = ( n2452 & n2456 ) | ( n2452 & n3166 ) | ( n2456 & n3166 ) ;
  assign n3375 = n3373 | n3374 ;
  assign n3376 = n2689 & n3250 ;
  assign n3377 = ( n2362 & n2689 ) | ( n2362 & n3267 ) | ( n2689 & n3267 ) ;
  assign n3378 = ( n3375 & ~n3376 ) | ( n3375 & n3377 ) | ( ~n3376 & n3377 ) ;
  assign n3379 = ( n2362 & n3375 ) | ( n2362 & n3376 ) | ( n3375 & n3376 ) ;
  assign n3380 = n3378 & ~n3379 ;
  assign n3381 = n3370 & n3380 ;
  assign n3382 = n3366 & n3368 ;
  assign n3383 = ( n3363 & n3366 ) | ( n3363 & n3382 ) | ( n3366 & n3382 ) ;
  assign n3384 = n3068 | n3383 ;
  assign n3385 = n3381 | n3384 ;
  assign n3386 = n2393 & n3126 ;
  assign n3387 = ( n2452 & n2456 ) | ( n2452 & n3128 ) | ( n2456 & n3128 ) ;
  assign n3388 = n3386 | n3387 ;
  assign n3389 = n2461 & n3351 ;
  assign n3390 = ( n2362 & n3388 ) | ( n2362 & n3389 ) | ( n3388 & n3389 ) ;
  assign n3391 = n2882 & n3250 ;
  assign n3392 = n2461 & n3166 ;
  assign n3393 = n2362 | n3392 ;
  assign n3394 = n3388 | n3393 ;
  assign n3395 = ( ~n3267 & n3388 ) | ( ~n3267 & n3392 ) | ( n3388 & n3392 ) ;
  assign n3396 = n3267 | n3395 ;
  assign n3397 = ( n2882 & n3394 ) | ( n2882 & n3396 ) | ( n3394 & n3396 ) ;
  assign n3398 = ~n3391 & n3397 ;
  assign n3399 = ~n3390 & n3398 ;
  assign n3400 = n3385 & n3399 ;
  assign n3401 = ( n2804 & ~n2959 ) | ( n2804 & n3069 ) | ( ~n2959 & n3069 ) ;
  assign n3402 = ( ~n2804 & n2959 ) | ( ~n2804 & n3401 ) | ( n2959 & n3401 ) ;
  assign n3403 = ( ~n3069 & n3401 ) | ( ~n3069 & n3402 ) | ( n3401 & n3402 ) ;
  assign n3404 = n3068 & n3383 ;
  assign n3405 = ( n3068 & n3381 ) | ( n3068 & n3404 ) | ( n3381 & n3404 ) ;
  assign n3406 = n3403 & n3405 ;
  assign n3407 = ( n3400 & n3403 ) | ( n3400 & n3406 ) | ( n3403 & n3406 ) ;
  assign n3408 = n3240 | n3407 ;
  assign n3409 = ( ~n2949 & n3070 ) | ( ~n2949 & n3072 ) | ( n3070 & n3072 ) ;
  assign n3410 = ( n2949 & ~n3072 ) | ( n2949 & n3409 ) | ( ~n3072 & n3409 ) ;
  assign n3411 = ( ~n3070 & n3409 ) | ( ~n3070 & n3410 ) | ( n3409 & n3410 ) ;
  assign n3412 = n3403 | n3405 ;
  assign n3413 = n3400 | n3412 ;
  assign n3414 = n3411 | n3413 ;
  assign n3415 = ( n3408 & n3411 ) | ( n3408 & n3414 ) | ( n3411 & n3414 ) ;
  assign n3416 = n3225 & n3415 ;
  assign n3417 = n2354 & n3166 ;
  assign n3418 = n2374 & n3128 ;
  assign n3419 = ( ~n2383 & n2384 ) | ( ~n2383 & n3126 ) | ( n2384 & n3126 ) ;
  assign n3420 = n3418 | n3419 ;
  assign n3421 = n3417 | n3420 ;
  assign n3422 = ( n2478 & n3163 ) | ( n2478 & n3421 ) | ( n3163 & n3421 ) ;
  assign n3423 = ( n2362 & ~n3421 ) | ( n2362 & n3422 ) | ( ~n3421 & n3422 ) ;
  assign n3424 = ~n3422 & n3423 ;
  assign n3425 = n3421 | n3423 ;
  assign n3426 = ( ~n2362 & n3424 ) | ( ~n2362 & n3425 ) | ( n3424 & n3425 ) ;
  assign n3427 = n3411 & n3413 ;
  assign n3428 = n3408 & n3427 ;
  assign n3429 = n3426 & n3428 ;
  assign n3430 = ( n3416 & n3426 ) | ( n3416 & n3429 ) | ( n3426 & n3429 ) ;
  assign n3431 = n3210 & n3430 ;
  assign n3432 = n3426 | n3428 ;
  assign n3433 = n3416 | n3432 ;
  assign n3434 = ( n3073 & ~n3076 ) | ( n3073 & n3086 ) | ( ~n3076 & n3086 ) ;
  assign n3435 = ( n3073 & n3076 ) | ( n3073 & ~n3086 ) | ( n3076 & ~n3086 ) ;
  assign n3436 = ( ~n3073 & n3434 ) | ( ~n3073 & n3435 ) | ( n3434 & n3435 ) ;
  assign n3437 = n3433 & n3436 ;
  assign n3438 = ( n3210 & n3431 ) | ( n3210 & n3437 ) | ( n3431 & n3437 ) ;
  assign n3439 = n3208 | n3438 ;
  assign n3440 = n2354 & n3126 ;
  assign n3441 = ~n3119 & n3128 ;
  assign n3442 = n3440 | n3441 ;
  assign n3443 = ( x0 & n3147 ) | ( x0 & n3163 ) | ( n3147 & n3163 ) ;
  assign n3444 = n3442 | n3443 ;
  assign n3445 = ( n3166 & n3442 ) | ( n3166 & n3444 ) | ( n3442 & n3444 ) ;
  assign n3446 = ( n3119 & ~n3147 ) | ( n3119 & n3178 ) | ( ~n3147 & n3178 ) ;
  assign n3447 = ( ~n3178 & n3179 ) | ( ~n3178 & n3446 ) | ( n3179 & n3446 ) ;
  assign n3448 = ( n3444 & n3445 ) | ( n3444 & ~n3447 ) | ( n3445 & ~n3447 ) ;
  assign n3449 = ~n2362 & n3448 ;
  assign n3450 = n2362 | n3449 ;
  assign n3451 = ( ~n3448 & n3449 ) | ( ~n3448 & n3450 ) | ( n3449 & n3450 ) ;
  assign n3452 = ( n3191 & n3439 ) | ( n3191 & n3451 ) | ( n3439 & n3451 ) ;
  assign n3453 = n3189 | n3452 ;
  assign n3454 = n3189 & n3452 ;
  assign n3455 = n3453 & ~n3454 ;
  assign n3456 = n784 | n1948 ;
  assign n3457 = n2327 | n3456 ;
  assign n3458 = n258 | n397 ;
  assign n3459 = n224 | n362 ;
  assign n3460 = n3458 | n3459 ;
  assign n3461 = n176 | n267 ;
  assign n3462 = n3460 | n3461 ;
  assign n3463 = n375 | n723 ;
  assign n3464 = n3462 | n3463 ;
  assign n3465 = n351 | n384 ;
  assign n3466 = n223 | n249 ;
  assign n3467 = n3465 | n3466 ;
  assign n3468 = n128 | n3467 ;
  assign n3469 = n247 | n297 ;
  assign n3470 = n3468 | n3469 ;
  assign n3471 = n3464 | n3470 ;
  assign n3472 = n154 | n280 ;
  assign n3473 = n232 | n477 ;
  assign n3474 = ( ~n3471 & n3472 ) | ( ~n3471 & n3473 ) | ( n3472 & n3473 ) ;
  assign n3475 = n3471 | n3474 ;
  assign n3476 = n3457 | n3475 ;
  assign n3477 = n360 | n2334 ;
  assign n3478 = n226 | n3477 ;
  assign n3479 = n734 | n3478 ;
  assign n3480 = n281 | n2239 ;
  assign n3481 = n3479 | n3480 ;
  assign n3482 = n3476 | n3481 ;
  assign n3483 = n141 | n363 ;
  assign n3484 = n305 | n356 ;
  assign n3485 = n3483 | n3484 ;
  assign n3486 = n291 | n705 ;
  assign n3487 = n325 | n3486 ;
  assign n3488 = n3485 | n3487 ;
  assign n3489 = n3482 | n3488 ;
  assign n3490 = n3455 & n3489 ;
  assign n3491 = n3455 & ~n3490 ;
  assign n3492 = ~n3455 & n3489 ;
  assign n3493 = n3491 | n3492 ;
  assign n3494 = n3210 | n3430 ;
  assign n3495 = n3437 | n3494 ;
  assign n3496 = ~n3438 & n3495 ;
  assign n3497 = n321 | n454 ;
  assign n3498 = n206 | n212 ;
  assign n3499 = n2064 | n3498 ;
  assign n3500 = n3497 | n3499 ;
  assign n3501 = n2099 | n3500 ;
  assign n3502 = n158 | n319 ;
  assign n3503 = n209 | n3502 ;
  assign n3504 = n411 | n3503 ;
  assign n3505 = n2172 | n3504 ;
  assign n3506 = n3501 | n3505 ;
  assign n3507 = n338 | n632 ;
  assign n3508 = n191 | n1947 ;
  assign n3509 = n3507 | n3508 ;
  assign n3510 = n404 | n3509 ;
  assign n3511 = n275 | n2245 ;
  assign n3512 = n778 | n2232 ;
  assign n3513 = ( ~n3510 & n3511 ) | ( ~n3510 & n3512 ) | ( n3511 & n3512 ) ;
  assign n3514 = n3510 | n3513 ;
  assign n3515 = n3506 | n3514 ;
  assign n3516 = ( n296 & n381 ) | ( n296 & ~n3466 ) | ( n381 & ~n3466 ) ;
  assign n3517 = n3466 | n3516 ;
  assign n3518 = n3515 | n3517 ;
  assign n3519 = n3496 & n3518 ;
  assign n3520 = n164 | n369 ;
  assign n3521 = n676 | n3520 ;
  assign n3522 = n2279 | n3521 ;
  assign n3523 = n293 | n705 ;
  assign n3524 = n680 | n3523 ;
  assign n3525 = n168 | n655 ;
  assign n3526 = n3524 | n3525 ;
  assign n3527 = n209 | n386 ;
  assign n3528 = n171 | n192 ;
  assign n3529 = n3527 | n3528 ;
  assign n3530 = n112 | n311 ;
  assign n3531 = n116 | n325 ;
  assign n3532 = n3530 | n3531 ;
  assign n3533 = n3529 | n3532 ;
  assign n3534 = n3526 | n3533 ;
  assign n3535 = n3522 | n3534 ;
  assign n3536 = n128 | n298 ;
  assign n3537 = n1933 | n3536 ;
  assign n3538 = n134 | n367 ;
  assign n3539 = n185 | n597 ;
  assign n3540 = n3538 | n3539 ;
  assign n3541 = n200 | n247 ;
  assign n3542 = n3540 | n3541 ;
  assign n3543 = n3537 | n3542 ;
  assign n3544 = n1042 | n3543 ;
  assign n3545 = n3535 | n3544 ;
  assign n3546 = n191 | n235 ;
  assign n3547 = n543 | n3546 ;
  assign n3548 = n284 | n897 ;
  assign n3549 = n3547 | n3548 ;
  assign n3550 = n157 | n3549 ;
  assign n3551 = n132 | n331 ;
  assign n3552 = n234 | n3551 ;
  assign n3553 = n3550 | n3552 ;
  assign n3554 = n3545 | n3553 ;
  assign n3555 = ( n3191 & ~n3439 ) | ( n3191 & n3451 ) | ( ~n3439 & n3451 ) ;
  assign n3556 = ( n3439 & ~n3451 ) | ( n3439 & n3555 ) | ( ~n3451 & n3555 ) ;
  assign n3557 = ( ~n3191 & n3555 ) | ( ~n3191 & n3556 ) | ( n3555 & n3556 ) ;
  assign n3558 = ( n3519 & n3554 ) | ( n3519 & n3557 ) | ( n3554 & n3557 ) ;
  assign n3559 = n3493 & n3558 ;
  assign n3560 = n3493 | n3558 ;
  assign n3561 = ~n3559 & n3560 ;
  assign n3562 = n3490 | n3559 ;
  assign n3563 = n3144 | n3159 ;
  assign n3564 = n3116 & ~n3563 ;
  assign n3565 = n2317 & n3564 ;
  assign n3566 = n165 | n176 ;
  assign n3567 = n711 | n722 ;
  assign n3568 = n356 | n390 ;
  assign n3569 = n192 | n3568 ;
  assign n3570 = n3567 | n3569 ;
  assign n3571 = n205 | n597 ;
  assign n3572 = n336 | n3571 ;
  assign n3573 = n3570 | n3572 ;
  assign n3574 = n252 | n604 ;
  assign n3575 = n739 | n3574 ;
  assign n3576 = n1020 | n3575 ;
  assign n3577 = n1957 | n3576 ;
  assign n3578 = n3573 | n3577 ;
  assign n3579 = n375 | n411 ;
  assign n3580 = n2241 | n3579 ;
  assign n3581 = n223 | n257 ;
  assign n3582 = n101 | n3581 ;
  assign n3583 = n3580 | n3582 ;
  assign n3584 = n477 | n3583 ;
  assign n3585 = n3578 | n3584 ;
  assign n3586 = n1013 & ~n3585 ;
  assign n3587 = ~n3566 & n3586 ;
  assign n3588 = n3565 & ~n3587 ;
  assign n3589 = n3587 | n3588 ;
  assign n3590 = ( ~n3565 & n3588 ) | ( ~n3565 & n3589 ) | ( n3588 & n3589 ) ;
  assign n3591 = n3166 & ~n3590 ;
  assign n3592 = n3126 & n3147 ;
  assign n3593 = n3128 & n3162 ;
  assign n3594 = n3592 | n3593 ;
  assign n3595 = n3591 | n3594 ;
  assign n3596 = ~n3162 & n3590 ;
  assign n3597 = n3162 & ~n3590 ;
  assign n3598 = n3596 | n3597 ;
  assign n3599 = n3147 | n3162 ;
  assign n3600 = ( ~n3169 & n3564 ) | ( ~n3169 & n3599 ) | ( n3564 & n3599 ) ;
  assign n3601 = ~n3598 & n3600 ;
  assign n3602 = ( n3147 & n3159 ) | ( n3147 & n3168 ) | ( n3159 & n3168 ) ;
  assign n3603 = ~n3598 & n3602 ;
  assign n3604 = ( n3178 & n3601 ) | ( n3178 & n3603 ) | ( n3601 & n3603 ) ;
  assign n3605 = ( n3178 & n3600 ) | ( n3178 & n3602 ) | ( n3600 & n3602 ) ;
  assign n3606 = n3598 & ~n3605 ;
  assign n3607 = n3604 | n3606 ;
  assign n3608 = n3163 | n3595 ;
  assign n3609 = ( n3595 & ~n3607 ) | ( n3595 & n3608 ) | ( ~n3607 & n3608 ) ;
  assign n3610 = ~n2362 & n3609 ;
  assign n3611 = n2362 & ~n3609 ;
  assign n3612 = n3610 | n3611 ;
  assign n3613 = n2374 & n2381 ;
  assign n3614 = n2354 & n2378 ;
  assign n3615 = n3613 | n3614 ;
  assign n3616 = ( n2365 & n2388 ) | ( n2365 & ~n3119 ) | ( n2388 & ~n3119 ) ;
  assign n3617 = n3615 | n3616 ;
  assign n3618 = ( n2366 & n3615 ) | ( n2366 & n3617 ) | ( n3615 & n3617 ) ;
  assign n3619 = ( ~n3197 & n3617 ) | ( ~n3197 & n3618 ) | ( n3617 & n3618 ) ;
  assign n3620 = ~n32 & n3619 ;
  assign n3621 = n32 | n3620 ;
  assign n3622 = ( ~n3619 & n3620 ) | ( ~n3619 & n3621 ) | ( n3620 & n3621 ) ;
  assign n3623 = n2461 & n2673 ;
  assign n3624 = ( n2452 & n2456 ) | ( n2452 & n2679 ) | ( n2456 & n2679 ) ;
  assign n3625 = n3623 | n3624 ;
  assign n3626 = ( ~n2383 & n2384 ) | ( ~n2383 & n2682 ) | ( n2384 & n2682 ) ;
  assign n3627 = n3625 | n3626 ;
  assign n3628 = n2686 | n3627 ;
  assign n3629 = ( ~n2924 & n3627 ) | ( ~n2924 & n3628 ) | ( n3627 & n3628 ) ;
  assign n3630 = ~n752 & n3629 ;
  assign n3631 = n752 & ~n3629 ;
  assign n3632 = n3630 | n3631 ;
  assign n3633 = n2860 | n2863 ;
  assign n3634 = n566 & n2425 ;
  assign n3635 = n2422 & n2512 ;
  assign n3636 = n2415 & n2499 ;
  assign n3637 = n3635 | n3636 ;
  assign n3638 = ( n2405 & n2409 ) | ( n2405 & n2501 ) | ( n2409 & n2501 ) ;
  assign n3639 = n3637 | n3638 ;
  assign n3640 = ( n2491 & n2585 ) | ( n2491 & n3639 ) | ( n2585 & n3639 ) ;
  assign n3641 = ( n3634 & ~n3639 ) | ( n3634 & n3640 ) | ( ~n3639 & n3640 ) ;
  assign n3642 = ~n3640 & n3641 ;
  assign n3643 = n3639 | n3641 ;
  assign n3644 = ( ~n3634 & n3642 ) | ( ~n3634 & n3643 ) | ( n3642 & n3643 ) ;
  assign n3645 = n3633 | n3644 ;
  assign n3646 = ~n3644 & n3645 ;
  assign n3647 = ( ~n3633 & n3645 ) | ( ~n3633 & n3646 ) | ( n3645 & n3646 ) ;
  assign n3648 = ~n2398 & n2559 ;
  assign n3649 = n2403 & n2557 ;
  assign n3650 = n3648 | n3649 ;
  assign n3651 = ( n2393 & n2549 ) | ( n2393 & n2562 ) | ( n2549 & n2562 ) ;
  assign n3652 = n3650 | n3651 ;
  assign n3653 = ( ~n2552 & n3650 ) | ( ~n2552 & n3652 ) | ( n3650 & n3652 ) ;
  assign n3654 = ( ~n2814 & n3652 ) | ( ~n2814 & n3653 ) | ( n3652 & n3653 ) ;
  assign n3655 = ~n977 & n3654 ;
  assign n3656 = n977 | n3655 ;
  assign n3657 = ( ~n3654 & n3655 ) | ( ~n3654 & n3656 ) | ( n3655 & n3656 ) ;
  assign n3658 = ~n3647 & n3657 ;
  assign n3659 = n3647 & ~n3657 ;
  assign n3660 = n3658 | n3659 ;
  assign n3661 = ( n2866 & n2868 ) | ( n2866 & ~n2871 ) | ( n2868 & ~n2871 ) ;
  assign n3662 = ( n3632 & n3660 ) | ( n3632 & ~n3661 ) | ( n3660 & ~n3661 ) ;
  assign n3663 = ( ~n3660 & n3661 ) | ( ~n3660 & n3662 ) | ( n3661 & n3662 ) ;
  assign n3664 = ( ~n3632 & n3662 ) | ( ~n3632 & n3663 ) | ( n3662 & n3663 ) ;
  assign n3665 = n2887 | n2890 ;
  assign n3666 = n3664 | n3665 ;
  assign n3667 = n3664 & n3665 ;
  assign n3668 = n3666 & ~n3667 ;
  assign n3669 = n3622 & n3668 ;
  assign n3670 = n3668 & ~n3669 ;
  assign n3671 = ( n3622 & ~n3669 ) | ( n3622 & n3670 ) | ( ~n3669 & n3670 ) ;
  assign n3672 = n2893 | n3100 ;
  assign n3673 = ~n3671 & n3672 ;
  assign n3674 = n3671 & ~n3672 ;
  assign n3675 = n3673 | n3674 ;
  assign n3676 = n3612 & n3675 ;
  assign n3677 = n3612 | n3675 ;
  assign n3678 = ~n3676 & n3677 ;
  assign n3679 = n3187 | n3454 ;
  assign n3680 = n3678 | n3679 ;
  assign n3681 = n3678 & n3679 ;
  assign n3682 = n3680 & ~n3681 ;
  assign n3683 = n645 | n649 ;
  assign n3684 = n642 | n3683 ;
  assign n3685 = n2327 | n3684 ;
  assign n3686 = n655 | n722 ;
  assign n3687 = n537 | n3686 ;
  assign n3688 = n175 | n441 ;
  assign n3689 = n3687 | n3688 ;
  assign n3690 = n802 | n3689 ;
  assign n3691 = n2106 | n3690 ;
  assign n3692 = n3685 | n3691 ;
  assign n3693 = n186 | n367 ;
  assign n3694 = n519 | n3693 ;
  assign n3695 = n3692 | n3694 ;
  assign n3696 = n3682 | n3695 ;
  assign n3697 = n3682 & n3695 ;
  assign n3698 = n3696 & ~n3697 ;
  assign n3699 = n3562 & n3698 ;
  assign n3700 = n3562 | n3698 ;
  assign n3701 = ~n3699 & n3700 ;
  assign n3702 = n3561 & n3701 ;
  assign n3703 = n3701 & ~n3702 ;
  assign n3704 = ( n3561 & ~n3702 ) | ( n3561 & n3703 ) | ( ~n3702 & n3703 ) ;
  assign n3705 = n3676 | n3681 ;
  assign n3706 = n2317 & n3587 ;
  assign n3707 = n456 & ~n460 ;
  assign n3708 = n102 | n865 ;
  assign n3709 = n634 | n3708 ;
  assign n3710 = n632 | n3709 ;
  assign n3711 = n3707 & ~n3710 ;
  assign n3712 = n721 | n2232 ;
  assign n3713 = n166 | n3712 ;
  assign n3714 = n270 | n3713 ;
  assign n3715 = n173 | n305 ;
  assign n3716 = n201 | n281 ;
  assign n3717 = n3715 | n3716 ;
  assign n3718 = n3714 | n3717 ;
  assign n3719 = n3711 & ~n3718 ;
  assign n3720 = ~n900 & n3719 ;
  assign n3721 = n134 | n331 ;
  assign n3722 = n238 | n248 ;
  assign n3723 = n3721 | n3722 ;
  assign n3724 = n2254 | n3723 ;
  assign n3725 = n3720 & ~n3724 ;
  assign n3726 = ~n3564 & n3706 ;
  assign n3727 = ( n3706 & n3725 ) | ( n3706 & n3726 ) | ( n3725 & n3726 ) ;
  assign n3728 = ( n3725 & n3726 ) | ( n3725 & ~n3727 ) | ( n3726 & ~n3727 ) ;
  assign n3729 = ( n3706 & ~n3727 ) | ( n3706 & n3728 ) | ( ~n3727 & n3728 ) ;
  assign n3730 = n3166 & ~n3729 ;
  assign n3731 = n3126 & n3162 ;
  assign n3732 = n3128 & ~n3590 ;
  assign n3733 = n3731 | n3732 ;
  assign n3734 = n3730 | n3733 ;
  assign n3735 = n3590 & n3729 ;
  assign n3736 = n3590 | n3729 ;
  assign n3737 = ~n3735 & n3736 ;
  assign n3738 = n3597 | n3737 ;
  assign n3739 = n3604 | n3738 ;
  assign n3740 = n3597 & n3737 ;
  assign n3741 = ( n3604 & n3737 ) | ( n3604 & n3740 ) | ( n3737 & n3740 ) ;
  assign n3742 = n3739 & ~n3741 ;
  assign n3743 = n3163 | n3734 ;
  assign n3744 = ( n3734 & n3742 ) | ( n3734 & n3743 ) | ( n3742 & n3743 ) ;
  assign n3745 = ~n2362 & n3744 ;
  assign n3746 = n2362 & ~n3744 ;
  assign n3747 = n3745 | n3746 ;
  assign n3748 = n2354 & n2381 ;
  assign n3749 = n2378 & ~n3119 ;
  assign n3750 = n3748 | n3749 ;
  assign n3751 = ( n2365 & n2388 ) | ( n2365 & n3147 ) | ( n2388 & n3147 ) ;
  assign n3752 = n3750 | n3751 ;
  assign n3753 = ( n2366 & n3750 ) | ( n2366 & n3752 ) | ( n3750 & n3752 ) ;
  assign n3754 = ( ~n3447 & n3752 ) | ( ~n3447 & n3753 ) | ( n3752 & n3753 ) ;
  assign n3755 = ~n32 & n3754 ;
  assign n3756 = n32 | n3755 ;
  assign n3757 = ( ~n3754 & n3755 ) | ( ~n3754 & n3756 ) | ( n3755 & n3756 ) ;
  assign n3758 = ( n3647 & n3657 ) | ( n3647 & n3661 ) | ( n3657 & n3661 ) ;
  assign n3759 = n2374 & n2682 ;
  assign n3760 = n2461 & n2679 ;
  assign n3761 = ( ~n2383 & n2384 ) | ( ~n2383 & n2673 ) | ( n2384 & n2673 ) ;
  assign n3762 = n3760 | n3761 ;
  assign n3763 = n3759 | n3762 ;
  assign n3764 = n2686 | n3763 ;
  assign n3765 = ( ~n2908 & n3763 ) | ( ~n2908 & n3764 ) | ( n3763 & n3764 ) ;
  assign n3766 = ~n752 & n3765 ;
  assign n3767 = n752 & ~n3765 ;
  assign n3768 = n3766 | n3767 ;
  assign n3769 = n2393 & n2559 ;
  assign n3770 = ~n2398 & n2557 ;
  assign n3771 = n3769 | n3770 ;
  assign n3772 = ( n2452 & n2456 ) | ( n2452 & n2563 ) | ( n2456 & n2563 ) ;
  assign n3773 = n3771 | n3772 ;
  assign n3774 = ( n2562 & n2689 ) | ( n2562 & n3773 ) | ( n2689 & n3773 ) ;
  assign n3775 = ( n977 & ~n3773 ) | ( n977 & n3774 ) | ( ~n3773 & n3774 ) ;
  assign n3776 = ~n3774 & n3775 ;
  assign n3777 = n3773 | n3775 ;
  assign n3778 = ( ~n977 & n3776 ) | ( ~n977 & n3777 ) | ( n3776 & n3777 ) ;
  assign n3779 = n566 & ~n2425 ;
  assign n3780 = ~n3639 & n3779 ;
  assign n3781 = ~n2491 & n3780 ;
  assign n3782 = ( ~n2585 & n3780 ) | ( ~n2585 & n3781 ) | ( n3780 & n3781 ) ;
  assign n3783 = n3644 | n3782 ;
  assign n3784 = ( n2860 & n3782 ) | ( n2860 & n3783 ) | ( n3782 & n3783 ) ;
  assign n3785 = ( n2863 & n3783 ) | ( n2863 & n3784 ) | ( n3783 & n3784 ) ;
  assign n3786 = n566 & ~n2422 ;
  assign n3787 = n2415 & n2512 ;
  assign n3788 = ( n2405 & n2409 ) | ( n2405 & n2499 ) | ( n2409 & n2499 ) ;
  assign n3789 = n3787 | n3788 ;
  assign n3790 = n2403 & n2501 ;
  assign n3791 = n2491 | n3790 ;
  assign n3792 = n3789 | n3791 ;
  assign n3793 = n3786 & n3792 ;
  assign n3794 = n3786 & n3790 ;
  assign n3795 = ( n3786 & n3789 ) | ( n3786 & n3794 ) | ( n3789 & n3794 ) ;
  assign n3796 = ( n2546 & n3793 ) | ( n2546 & n3795 ) | ( n3793 & n3795 ) ;
  assign n3797 = n3786 | n3792 ;
  assign n3798 = n3786 | n3790 ;
  assign n3799 = n3789 | n3798 ;
  assign n3800 = ( n2546 & n3797 ) | ( n2546 & n3799 ) | ( n3797 & n3799 ) ;
  assign n3801 = ~n3796 & n3800 ;
  assign n3802 = n3785 & n3801 ;
  assign n3803 = n3785 | n3801 ;
  assign n3804 = ~n3802 & n3803 ;
  assign n3805 = n3778 & n3804 ;
  assign n3806 = n3804 & ~n3805 ;
  assign n3807 = ( n3778 & ~n3805 ) | ( n3778 & n3806 ) | ( ~n3805 & n3806 ) ;
  assign n3808 = ( n3758 & n3768 ) | ( n3758 & ~n3807 ) | ( n3768 & ~n3807 ) ;
  assign n3809 = ( ~n3768 & n3807 ) | ( ~n3768 & n3808 ) | ( n3807 & n3808 ) ;
  assign n3810 = ( ~n3758 & n3808 ) | ( ~n3758 & n3809 ) | ( n3808 & n3809 ) ;
  assign n3811 = n3660 & n3661 ;
  assign n3812 = ( n3632 & n3660 ) | ( n3632 & n3661 ) | ( n3660 & n3661 ) ;
  assign n3813 = ( n3667 & ~n3811 ) | ( n3667 & n3812 ) | ( ~n3811 & n3812 ) ;
  assign n3814 = n3810 | n3813 ;
  assign n3815 = n3810 & n3813 ;
  assign n3816 = n3814 & ~n3815 ;
  assign n3817 = n3757 & n3816 ;
  assign n3818 = n3816 & ~n3817 ;
  assign n3819 = ( n3757 & ~n3817 ) | ( n3757 & n3818 ) | ( ~n3817 & n3818 ) ;
  assign n3820 = ( n3669 & n3671 ) | ( n3669 & ~n3674 ) | ( n3671 & ~n3674 ) ;
  assign n3821 = ~n3819 & n3820 ;
  assign n3822 = n3819 & ~n3820 ;
  assign n3823 = n3821 | n3822 ;
  assign n3824 = n3747 & n3823 ;
  assign n3825 = n3747 | n3823 ;
  assign n3826 = ~n3824 & n3825 ;
  assign n3827 = n3705 | n3826 ;
  assign n3828 = n3705 & n3826 ;
  assign n3829 = n3827 & ~n3828 ;
  assign n3830 = n797 | n2139 ;
  assign n3831 = n478 | n3830 ;
  assign n3832 = n2075 | n3831 ;
  assign n3833 = n2072 | n3832 ;
  assign n3834 = n3471 | n3833 ;
  assign n3835 = n181 | n355 ;
  assign n3836 = n482 | n3835 ;
  assign n3837 = n166 | n3836 ;
  assign n3838 = n2327 | n2336 ;
  assign n3839 = n3837 | n3838 ;
  assign n3840 = n400 | n404 ;
  assign n3841 = n3839 | n3840 ;
  assign n3842 = n127 | n204 ;
  assign n3843 = n305 | n597 ;
  assign n3844 = n3842 | n3843 ;
  assign n3845 = n3841 | n3844 ;
  assign n3846 = n3834 | n3845 ;
  assign n3847 = n3829 | n3846 ;
  assign n3848 = n3829 & n3846 ;
  assign n3849 = n3847 & ~n3848 ;
  assign n3850 = n3697 | n3699 ;
  assign n3851 = n3849 & n3850 ;
  assign n3852 = n3849 | n3850 ;
  assign n3853 = ~n3851 & n3852 ;
  assign n3854 = n3702 & n3853 ;
  assign n3855 = n3702 | n3853 ;
  assign n3856 = ~n3854 & n3855 ;
  assign n3857 = x22 & ~x23 ;
  assign n3858 = ~x22 & x23 ;
  assign n3859 = n3857 | n3858 ;
  assign n3860 = n3704 & n3859 ;
  assign n3861 = ~n3856 & n3860 ;
  assign n3862 = n3856 & ~n3860 ;
  assign n3863 = n3861 | n3862 ;
  assign n3864 = n3824 | n3828 ;
  assign n3865 = n3126 & ~n3590 ;
  assign n3866 = n3128 & ~n3729 ;
  assign n3867 = n3865 | n3866 ;
  assign n3868 = ( ~n3601 & n3729 ) | ( ~n3601 & n3736 ) | ( n3729 & n3736 ) ;
  assign n3869 = ( ~n3603 & n3729 ) | ( ~n3603 & n3736 ) | ( n3729 & n3736 ) ;
  assign n3870 = ( ~n3178 & n3868 ) | ( ~n3178 & n3869 ) | ( n3868 & n3869 ) ;
  assign n3871 = n3729 & ~n3740 ;
  assign n3872 = ( ~n3601 & n3735 ) | ( ~n3601 & n3871 ) | ( n3735 & n3871 ) ;
  assign n3873 = ( ~n3603 & n3735 ) | ( ~n3603 & n3871 ) | ( n3735 & n3871 ) ;
  assign n3874 = ( ~n3178 & n3872 ) | ( ~n3178 & n3873 ) | ( n3872 & n3873 ) ;
  assign n3875 = n3870 & ~n3874 ;
  assign n3876 = n3163 | n3867 ;
  assign n3877 = ( n3867 & n3875 ) | ( n3867 & n3876 ) | ( n3875 & n3876 ) ;
  assign n3878 = n3250 & n3875 ;
  assign n3879 = ( n2362 & n3867 ) | ( n2362 & n3878 ) | ( n3867 & n3878 ) ;
  assign n3880 = n3877 & ~n3879 ;
  assign n3881 = ( n2362 & n3254 ) | ( n2362 & ~n3875 ) | ( n3254 & ~n3875 ) ;
  assign n3882 = ~n3867 & n3881 ;
  assign n3883 = n3880 | n3882 ;
  assign n3884 = n2381 & ~n3119 ;
  assign n3885 = n2378 & n3147 ;
  assign n3886 = n3884 | n3885 ;
  assign n3887 = ( n2365 & n2388 ) | ( n2365 & n3162 ) | ( n2388 & n3162 ) ;
  assign n3888 = n3886 | n3887 ;
  assign n3889 = ( n2366 & n3886 ) | ( n2366 & n3888 ) | ( n3886 & n3888 ) ;
  assign n3890 = ( n3182 & n3888 ) | ( n3182 & n3889 ) | ( n3888 & n3889 ) ;
  assign n3891 = n32 & n3890 ;
  assign n3892 = n32 & ~n3891 ;
  assign n3893 = ( n3890 & ~n3891 ) | ( n3890 & n3892 ) | ( ~n3891 & n3892 ) ;
  assign n3894 = n2354 & n2682 ;
  assign n3895 = n2374 & n2673 ;
  assign n3896 = ( ~n2383 & n2384 ) | ( ~n2383 & n2679 ) | ( n2384 & n2679 ) ;
  assign n3897 = n3895 | n3896 ;
  assign n3898 = n3894 | n3897 ;
  assign n3899 = ( n2478 & n2686 ) | ( n2478 & n3898 ) | ( n2686 & n3898 ) ;
  assign n3900 = ( n752 & ~n3898 ) | ( n752 & n3899 ) | ( ~n3898 & n3899 ) ;
  assign n3901 = ~n3899 & n3900 ;
  assign n3902 = n3898 | n3900 ;
  assign n3903 = ( ~n752 & n3901 ) | ( ~n752 & n3902 ) | ( n3901 & n3902 ) ;
  assign n3904 = n566 & ~n2415 ;
  assign n3905 = n2403 & n2499 ;
  assign n3906 = ( n2405 & n2409 ) | ( n2405 & n2512 ) | ( n2409 & n2512 ) ;
  assign n3907 = n3905 | n3906 ;
  assign n3908 = ~n2398 & n2501 ;
  assign n3909 = n2491 | n3908 ;
  assign n3910 = n3907 | n3909 ;
  assign n3911 = n3904 & n3910 ;
  assign n3912 = n3904 & n3908 ;
  assign n3913 = ( n3904 & n3907 ) | ( n3904 & n3912 ) | ( n3907 & n3912 ) ;
  assign n3914 = ( ~n2708 & n3911 ) | ( ~n2708 & n3913 ) | ( n3911 & n3913 ) ;
  assign n3915 = n3904 | n3910 ;
  assign n3916 = n3904 | n3908 ;
  assign n3917 = n3907 | n3916 ;
  assign n3918 = ( ~n2708 & n3915 ) | ( ~n2708 & n3917 ) | ( n3915 & n3917 ) ;
  assign n3919 = ~n3914 & n3918 ;
  assign n3920 = n566 & n2422 ;
  assign n3921 = ( n3789 & n3790 ) | ( n3789 & n3920 ) | ( n3790 & n3920 ) ;
  assign n3922 = ( n2546 & n3792 ) | ( n2546 & n3921 ) | ( n3792 & n3921 ) ;
  assign n3923 = n3920 & ~n3922 ;
  assign n3924 = n3802 | n3923 ;
  assign n3925 = n2393 & n2557 ;
  assign n3926 = ( n2452 & n2456 ) | ( n2452 & n2559 ) | ( n2456 & n2559 ) ;
  assign n3927 = n3925 | n3926 ;
  assign n3928 = ( n2461 & n2549 ) | ( n2461 & n2562 ) | ( n2549 & n2562 ) ;
  assign n3929 = n3927 | n3928 ;
  assign n3930 = ( n2563 & n3927 ) | ( n2563 & n3929 ) | ( n3927 & n3929 ) ;
  assign n3931 = ( n2882 & n3929 ) | ( n2882 & n3930 ) | ( n3929 & n3930 ) ;
  assign n3932 = n977 & n3931 ;
  assign n3933 = n977 & ~n3932 ;
  assign n3934 = ( n3931 & ~n3932 ) | ( n3931 & n3933 ) | ( ~n3932 & n3933 ) ;
  assign n3935 = ( n3919 & ~n3924 ) | ( n3919 & n3934 ) | ( ~n3924 & n3934 ) ;
  assign n3936 = ( n3924 & ~n3934 ) | ( n3924 & n3935 ) | ( ~n3934 & n3935 ) ;
  assign n3937 = ( ~n3919 & n3935 ) | ( ~n3919 & n3936 ) | ( n3935 & n3936 ) ;
  assign n3938 = n3758 & ~n3807 ;
  assign n3939 = ( n3758 & n3805 ) | ( n3758 & ~n3938 ) | ( n3805 & ~n3938 ) ;
  assign n3940 = ~n3937 & n3939 ;
  assign n3941 = n3937 & ~n3939 ;
  assign n3942 = n3940 | n3941 ;
  assign n3943 = ( n3768 & ~n3808 ) | ( n3768 & n3938 ) | ( ~n3808 & n3938 ) ;
  assign n3944 = n3815 | n3943 ;
  assign n3945 = ( n3903 & ~n3942 ) | ( n3903 & n3944 ) | ( ~n3942 & n3944 ) ;
  assign n3946 = ( n3942 & ~n3944 ) | ( n3942 & n3945 ) | ( ~n3944 & n3945 ) ;
  assign n3947 = ( ~n3903 & n3945 ) | ( ~n3903 & n3946 ) | ( n3945 & n3946 ) ;
  assign n3948 = n3893 & n3947 ;
  assign n3949 = n3947 & ~n3948 ;
  assign n3950 = ( n3893 & ~n3948 ) | ( n3893 & n3949 ) | ( ~n3948 & n3949 ) ;
  assign n3951 = ( n3817 & n3819 ) | ( n3817 & ~n3822 ) | ( n3819 & ~n3822 ) ;
  assign n3952 = ( n3883 & n3950 ) | ( n3883 & ~n3951 ) | ( n3950 & ~n3951 ) ;
  assign n3953 = ( ~n3950 & n3951 ) | ( ~n3950 & n3952 ) | ( n3951 & n3952 ) ;
  assign n3954 = ( ~n3883 & n3952 ) | ( ~n3883 & n3953 ) | ( n3952 & n3953 ) ;
  assign n3955 = n3864 & ~n3954 ;
  assign n3956 = ~n3864 & n3954 ;
  assign n3957 = n3955 | n3956 ;
  assign n3958 = n141 | n349 ;
  assign n3959 = n1949 | n3958 ;
  assign n3960 = n116 | n258 ;
  assign n3961 = n165 | n3960 ;
  assign n3962 = n3959 | n3961 ;
  assign n3963 = n325 | n368 ;
  assign n3964 = n775 | n3963 ;
  assign n3965 = n3962 | n3964 ;
  assign n3966 = n670 | n3965 ;
  assign n3967 = n179 | n192 ;
  assign n3968 = n164 | n256 ;
  assign n3969 = n3967 | n3968 ;
  assign n3970 = n284 | n293 ;
  assign n3971 = n238 | n3970 ;
  assign n3972 = n3969 | n3971 ;
  assign n3973 = n3501 | n3972 ;
  assign n3974 = n3966 | n3973 ;
  assign n3975 = n3957 & n3974 ;
  assign n3976 = n3957 | n3974 ;
  assign n3977 = ~n3975 & n3976 ;
  assign n3978 = n3848 | n3851 ;
  assign n3979 = n3977 & n3978 ;
  assign n3980 = n3978 & ~n3979 ;
  assign n3981 = ( n3977 & ~n3979 ) | ( n3977 & n3980 ) | ( ~n3979 & n3980 ) ;
  assign n3982 = n3854 | n3981 ;
  assign n3983 = n3854 & n3981 ;
  assign n3984 = n3982 & ~n3983 ;
  assign n3985 = n3704 | n3856 ;
  assign n3986 = n3859 & n3985 ;
  assign n3987 = ~n3984 & n3986 ;
  assign n3988 = n3984 & ~n3986 ;
  assign n3989 = n3987 | n3988 ;
  assign n3990 = n3984 | n3985 ;
  assign n3991 = n3859 & n3990 ;
  assign n3992 = n3975 | n3979 ;
  assign n3993 = n3903 & n3942 ;
  assign n3994 = n3903 | n3942 ;
  assign n3995 = ( n3944 & n3993 ) | ( n3944 & n3994 ) | ( n3993 & n3994 ) ;
  assign n3996 = ~n2398 & n2499 ;
  assign n3997 = n2403 & n2512 ;
  assign n3998 = n3996 | n3997 ;
  assign n3999 = n2393 & n2501 ;
  assign n4000 = n2491 | n3999 ;
  assign n4001 = n3998 | n4000 ;
  assign n4002 = n566 & n2415 ;
  assign n4003 = ( ~n2410 & n3904 ) | ( ~n2410 & n4002 ) | ( n3904 & n4002 ) ;
  assign n4004 = n4001 & n4003 ;
  assign n4005 = n3999 & n4003 ;
  assign n4006 = ( n3998 & n4003 ) | ( n3998 & n4005 ) | ( n4003 & n4005 ) ;
  assign n4007 = ( ~n2814 & n4004 ) | ( ~n2814 & n4006 ) | ( n4004 & n4006 ) ;
  assign n4008 = n4001 | n4003 ;
  assign n4009 = n3999 | n4003 ;
  assign n4010 = n3998 | n4009 ;
  assign n4011 = ( ~n2814 & n4008 ) | ( ~n2814 & n4010 ) | ( n4008 & n4010 ) ;
  assign n4012 = ~n4007 & n4011 ;
  assign n4013 = ( n3907 & n3908 ) | ( n3907 & n4002 ) | ( n3908 & n4002 ) ;
  assign n4014 = ( ~n2708 & n3910 ) | ( ~n2708 & n4013 ) | ( n3910 & n4013 ) ;
  assign n4015 = n4002 & ~n4014 ;
  assign n4016 = n3919 & n3924 ;
  assign n4017 = n4015 | n4016 ;
  assign n4018 = ~n4012 & n4017 ;
  assign n4019 = n4012 & ~n4017 ;
  assign n4020 = n2461 & n2559 ;
  assign n4021 = ( n2452 & n2456 ) | ( n2452 & n2557 ) | ( n2456 & n2557 ) ;
  assign n4022 = n4020 | n4021 ;
  assign n4023 = ( ~n2383 & n2384 ) | ( ~n2383 & n2563 ) | ( n2384 & n2563 ) ;
  assign n4024 = n4022 | n4023 ;
  assign n4025 = n2562 | n4024 ;
  assign n4026 = ( ~n2924 & n4024 ) | ( ~n2924 & n4025 ) | ( n4024 & n4025 ) ;
  assign n4027 = ~n977 & n4026 ;
  assign n4028 = n977 | n4027 ;
  assign n4029 = ( ~n4026 & n4027 ) | ( ~n4026 & n4028 ) | ( n4027 & n4028 ) ;
  assign n4030 = n4019 | n4029 ;
  assign n4031 = n4018 | n4030 ;
  assign n4032 = ( n4018 & n4019 ) | ( n4018 & n4029 ) | ( n4019 & n4029 ) ;
  assign n4033 = n4031 & ~n4032 ;
  assign n4034 = ( n3919 & n3924 ) | ( n3919 & n3934 ) | ( n3924 & n3934 ) ;
  assign n4035 = ~n4016 & n4034 ;
  assign n4036 = ( n3939 & ~n3940 ) | ( n3939 & n4035 ) | ( ~n3940 & n4035 ) ;
  assign n4037 = n4033 & n4036 ;
  assign n4038 = n4033 | n4036 ;
  assign n4039 = ~n4037 & n4038 ;
  assign n4040 = n2682 & ~n3119 ;
  assign n4041 = n2374 & n2679 ;
  assign n4042 = n2354 & n2673 ;
  assign n4043 = n4041 | n4042 ;
  assign n4044 = n4040 | n4043 ;
  assign n4045 = n2686 | n4044 ;
  assign n4046 = ( ~n3197 & n4044 ) | ( ~n3197 & n4045 ) | ( n4044 & n4045 ) ;
  assign n4047 = ~n752 & n4046 ;
  assign n4048 = n752 & ~n4046 ;
  assign n4049 = n4047 | n4048 ;
  assign n4050 = n4039 & n4049 ;
  assign n4051 = n4039 & ~n4050 ;
  assign n4052 = ~n4039 & n4049 ;
  assign n4053 = n4051 | n4052 ;
  assign n4054 = n3995 & n4053 ;
  assign n4055 = n4053 & ~n4054 ;
  assign n4056 = ( n3995 & ~n4054 ) | ( n3995 & n4055 ) | ( ~n4054 & n4055 ) ;
  assign n4057 = n3126 & ~n3729 ;
  assign n4058 = n3163 & ~n3729 ;
  assign n4059 = n4057 | n4058 ;
  assign n4060 = ( ~n3590 & n4057 ) | ( ~n3590 & n4059 ) | ( n4057 & n4059 ) ;
  assign n4061 = ( n3604 & n4059 ) | ( n3604 & n4060 ) | ( n4059 & n4060 ) ;
  assign n4062 = n2362 & ~n4061 ;
  assign n4063 = ~n2362 & n4061 ;
  assign n4064 = n4062 | n4063 ;
  assign n4065 = n2381 & n3147 ;
  assign n4066 = n2378 & n3162 ;
  assign n4067 = n4065 | n4066 ;
  assign n4068 = ( n2365 & n2388 ) | ( n2365 & ~n3590 ) | ( n2388 & ~n3590 ) ;
  assign n4069 = n4067 | n4068 ;
  assign n4070 = ( n2366 & n4067 ) | ( n2366 & n4069 ) | ( n4067 & n4069 ) ;
  assign n4071 = ( ~n3607 & n4069 ) | ( ~n3607 & n4070 ) | ( n4069 & n4070 ) ;
  assign n4072 = ~n32 & n4071 ;
  assign n4073 = n32 | n4072 ;
  assign n4074 = ( ~n4071 & n4072 ) | ( ~n4071 & n4073 ) | ( n4072 & n4073 ) ;
  assign n4075 = ( n4056 & n4064 ) | ( n4056 & ~n4074 ) | ( n4064 & ~n4074 ) ;
  assign n4076 = ( ~n4064 & n4074 ) | ( ~n4064 & n4075 ) | ( n4074 & n4075 ) ;
  assign n4077 = ( ~n4056 & n4075 ) | ( ~n4056 & n4076 ) | ( n4075 & n4076 ) ;
  assign n4078 = ( n3893 & n3947 ) | ( n3893 & n3951 ) | ( n3947 & n3951 ) ;
  assign n4079 = n4077 & n4078 ;
  assign n4080 = n4077 | n4078 ;
  assign n4081 = ~n4079 & n4080 ;
  assign n4082 = n3883 & ~n3953 ;
  assign n4083 = ( n3883 & ~n3952 ) | ( n3883 & n4082 ) | ( ~n3952 & n4082 ) ;
  assign n4084 = ( n3864 & n3954 ) | ( n3864 & n4083 ) | ( n3954 & n4083 ) ;
  assign n4085 = ( n4081 & ~n4083 ) | ( n4081 & n4084 ) | ( ~n4083 & n4084 ) ;
  assign n4086 = ~n4084 & n4085 ;
  assign n4087 = n4083 | n4085 ;
  assign n4088 = ( ~n4081 & n4086 ) | ( ~n4081 & n4087 ) | ( n4086 & n4087 ) ;
  assign n4089 = n97 | n481 ;
  assign n4090 = n519 | n623 ;
  assign n4091 = n168 | n2139 ;
  assign n4092 = n3524 | n4091 ;
  assign n4093 = n206 | n837 ;
  assign n4094 = n4092 | n4093 ;
  assign n4095 = n190 | n4094 ;
  assign n4096 = n4090 | n4095 ;
  assign n4097 = n297 | n411 ;
  assign n4098 = n400 | n4097 ;
  assign n4099 = n741 | n4098 ;
  assign n4100 = n273 | n291 ;
  assign n4101 = n4099 | n4100 ;
  assign n4102 = n1983 | n4101 ;
  assign n4103 = n4096 | n4102 ;
  assign n4104 = n4089 | n4103 ;
  assign n4105 = n4088 & n4104 ;
  assign n4106 = n4104 & ~n4105 ;
  assign n4107 = ( n4088 & ~n4105 ) | ( n4088 & n4106 ) | ( ~n4105 & n4106 ) ;
  assign n4108 = n3992 & n4107 ;
  assign n4109 = n3992 | n4107 ;
  assign n4110 = ~n4108 & n4109 ;
  assign n4111 = n3983 & n4110 ;
  assign n4112 = n3983 & ~n4111 ;
  assign n4113 = ( n4110 & ~n4111 ) | ( n4110 & n4112 ) | ( ~n4111 & n4112 ) ;
  assign n4114 = n3991 & n4113 ;
  assign n4115 = n3991 | n4113 ;
  assign n4116 = ~n4114 & n4115 ;
  assign n4117 = n2682 & n3147 ;
  assign n4118 = n2354 & n2679 ;
  assign n4119 = n2673 & ~n3119 ;
  assign n4120 = n4118 | n4119 ;
  assign n4121 = n4117 | n4120 ;
  assign n4122 = n2686 | n4121 ;
  assign n4123 = ( ~n3447 & n4121 ) | ( ~n3447 & n4122 ) | ( n4121 & n4122 ) ;
  assign n4124 = ~n752 & n4123 ;
  assign n4125 = n752 & ~n4123 ;
  assign n4126 = n4124 | n4125 ;
  assign n4127 = n4032 | n4037 ;
  assign n4128 = n4012 & n4017 ;
  assign n4129 = ( n566 & n2405 ) | ( n566 & n2409 ) | ( n2405 & n2409 ) ;
  assign n4130 = ~n4001 & n4129 ;
  assign n4131 = ~n3999 & n4129 ;
  assign n4132 = ~n3998 & n4131 ;
  assign n4133 = ( n2814 & n4130 ) | ( n2814 & n4132 ) | ( n4130 & n4132 ) ;
  assign n4134 = n4128 | n4133 ;
  assign n4135 = n2393 & n2499 ;
  assign n4136 = ~n2398 & n2512 ;
  assign n4137 = n4135 | n4136 ;
  assign n4138 = ( n2452 & n2456 ) | ( n2452 & n2501 ) | ( n2456 & n2501 ) ;
  assign n4139 = n4137 | n4138 ;
  assign n4140 = n566 & ~n4139 ;
  assign n4141 = n566 & n2491 ;
  assign n4142 = ( n2689 & ~n4140 ) | ( n2689 & n4141 ) | ( ~n4140 & n4141 ) ;
  assign n4143 = n4140 & ~n4142 ;
  assign n4144 = n566 & n2362 ;
  assign n4145 = n2403 & n4144 ;
  assign n4146 = n566 & n2403 ;
  assign n4147 = n2362 & ~n4145 ;
  assign n4148 = ( ~n4145 & n4146 ) | ( ~n4145 & n4147 ) | ( n4146 & n4147 ) ;
  assign n4149 = n2491 | n4139 ;
  assign n4150 = ( n2689 & n4139 ) | ( n2689 & n4149 ) | ( n4139 & n4149 ) ;
  assign n4151 = ~n566 & n4150 ;
  assign n4152 = ( ~n4143 & n4148 ) | ( ~n4143 & n4151 ) | ( n4148 & n4151 ) ;
  assign n4153 = n4143 | n4152 ;
  assign n4154 = ( n4143 & n4148 ) | ( n4143 & n4151 ) | ( n4148 & n4151 ) ;
  assign n4155 = n4153 & ~n4154 ;
  assign n4156 = n2461 & n2557 ;
  assign n4157 = ( ~n2383 & n2384 ) | ( ~n2383 & n2559 ) | ( n2384 & n2559 ) ;
  assign n4158 = n4156 | n4157 ;
  assign n4159 = n2374 & n2563 ;
  assign n4160 = n2562 | n4159 ;
  assign n4161 = n4158 | n4160 ;
  assign n4162 = n977 & n4161 ;
  assign n4163 = n977 & n4159 ;
  assign n4164 = ( n977 & n4158 ) | ( n977 & n4163 ) | ( n4158 & n4163 ) ;
  assign n4165 = ( ~n2908 & n4162 ) | ( ~n2908 & n4164 ) | ( n4162 & n4164 ) ;
  assign n4166 = n977 | n4161 ;
  assign n4167 = n977 | n4159 ;
  assign n4168 = n4158 | n4167 ;
  assign n4169 = ( ~n2908 & n4166 ) | ( ~n2908 & n4168 ) | ( n4166 & n4168 ) ;
  assign n4170 = ~n4165 & n4169 ;
  assign n4171 = ( n4134 & n4155 ) | ( n4134 & n4170 ) | ( n4155 & n4170 ) ;
  assign n4172 = ( n4155 & n4170 ) | ( n4155 & ~n4171 ) | ( n4170 & ~n4171 ) ;
  assign n4173 = ( n4134 & ~n4171 ) | ( n4134 & n4172 ) | ( ~n4171 & n4172 ) ;
  assign n4174 = ( n4126 & n4127 ) | ( n4126 & ~n4173 ) | ( n4127 & ~n4173 ) ;
  assign n4175 = ( ~n4127 & n4173 ) | ( ~n4127 & n4174 ) | ( n4173 & n4174 ) ;
  assign n4176 = ( ~n4126 & n4174 ) | ( ~n4126 & n4175 ) | ( n4174 & n4175 ) ;
  assign n4177 = n4050 | n4054 ;
  assign n4178 = n4176 & n4177 ;
  assign n4179 = n4176 | n4177 ;
  assign n4180 = ~n4178 & n4179 ;
  assign n4181 = n2381 & n3162 ;
  assign n4182 = n2378 & ~n3590 ;
  assign n4183 = n4181 | n4182 ;
  assign n4184 = n2366 & ~n3729 ;
  assign n4185 = n2388 | n4184 ;
  assign n4186 = n4183 | n4185 ;
  assign n4187 = n32 & n4186 ;
  assign n4188 = n32 & n4184 ;
  assign n4189 = ( n32 & n4183 ) | ( n32 & n4188 ) | ( n4183 & n4188 ) ;
  assign n4190 = ( n3742 & n4187 ) | ( n3742 & n4189 ) | ( n4187 & n4189 ) ;
  assign n4191 = n32 | n4186 ;
  assign n4192 = n32 | n4184 ;
  assign n4193 = n4183 | n4192 ;
  assign n4194 = ( n3742 & n4191 ) | ( n3742 & n4193 ) | ( n4191 & n4193 ) ;
  assign n4195 = ~n4190 & n4194 ;
  assign n4196 = n4180 & n4195 ;
  assign n4197 = n4180 | n4195 ;
  assign n4198 = ~n4196 & n4197 ;
  assign n4199 = ( n4056 & n4064 ) | ( n4056 & n4074 ) | ( n4064 & n4074 ) ;
  assign n4200 = n4198 | n4199 ;
  assign n4201 = n4198 & n4199 ;
  assign n4202 = n4200 & ~n4201 ;
  assign n4203 = n4079 | n4202 ;
  assign n4204 = n3864 & n3954 ;
  assign n4205 = ( n4081 & n4083 ) | ( n4081 & n4204 ) | ( n4083 & n4204 ) ;
  assign n4206 = n4203 | n4205 ;
  assign n4207 = ( n4079 & n4202 ) | ( n4079 & n4205 ) | ( n4202 & n4205 ) ;
  assign n4208 = n4206 & ~n4207 ;
  assign n4209 = n306 | n1949 ;
  assign n4210 = n527 | n4209 ;
  assign n4211 = n899 | n4210 ;
  assign n4212 = n2285 | n4211 ;
  assign n4213 = n444 | n2241 ;
  assign n4214 = n143 | n405 ;
  assign n4215 = n220 | n4214 ;
  assign n4216 = n4213 | n4215 ;
  assign n4217 = n617 | n4216 ;
  assign n4218 = n4212 | n4217 ;
  assign n4219 = n4105 | n4108 ;
  assign n4220 = ( n4208 & n4218 ) | ( n4208 & ~n4219 ) | ( n4218 & ~n4219 ) ;
  assign n4221 = ( ~n4218 & n4219 ) | ( ~n4218 & n4220 ) | ( n4219 & n4220 ) ;
  assign n4222 = ( ~n4208 & n4220 ) | ( ~n4208 & n4221 ) | ( n4220 & n4221 ) ;
  assign n4223 = n4111 | n4222 ;
  assign n4224 = n4111 & n4222 ;
  assign n4225 = n4223 & ~n4224 ;
  assign n4226 = n3990 | n4113 ;
  assign n4227 = n3859 & n4226 ;
  assign n4228 = ~n4225 & n4227 ;
  assign n4229 = n4225 & ~n4227 ;
  assign n4230 = n4228 | n4229 ;
  assign n4315 = ( n4208 & n4218 ) | ( n4208 & n4219 ) | ( n4218 & n4219 ) ;
  assign n4231 = n2381 & ~n3590 ;
  assign n4232 = n2378 & ~n3729 ;
  assign n4233 = n4231 | n4232 ;
  assign n4234 = n2389 & n3875 ;
  assign n4235 = ( n32 & n4233 ) | ( n32 & n4234 ) | ( n4233 & n4234 ) ;
  assign n4236 = ( n32 & n2481 ) | ( n32 & n3875 ) | ( n2481 & n3875 ) ;
  assign n4237 = n4233 | n4236 ;
  assign n4238 = ~n4235 & n4237 ;
  assign n4239 = n2682 & n3162 ;
  assign n4240 = n2679 & ~n3119 ;
  assign n4241 = n2673 & n3147 ;
  assign n4242 = n4240 | n4241 ;
  assign n4243 = n4239 | n4242 ;
  assign n4244 = n2686 | n4243 ;
  assign n4245 = ( n3182 & n4243 ) | ( n3182 & n4244 ) | ( n4243 & n4244 ) ;
  assign n4246 = ~n752 & n4245 ;
  assign n4247 = n752 & ~n4245 ;
  assign n4248 = n4246 | n4247 ;
  assign n4249 = n4145 | n4154 ;
  assign n4250 = ~n2398 & n4144 ;
  assign n4251 = n2362 | n2398 ;
  assign n4252 = n566 & ~n4251 ;
  assign n4253 = ( n2362 & ~n4250 ) | ( n2362 & n4252 ) | ( ~n4250 & n4252 ) ;
  assign n4254 = n4249 | n4253 ;
  assign n4255 = ~n4253 & n4254 ;
  assign n4256 = ( ~n4249 & n4254 ) | ( ~n4249 & n4255 ) | ( n4254 & n4255 ) ;
  assign n4257 = n2393 & n2512 ;
  assign n4258 = ( n2452 & n2456 ) | ( n2452 & n2499 ) | ( n2456 & n2499 ) ;
  assign n4259 = n4257 | n4258 ;
  assign n4260 = ( n2461 & n2488 ) | ( n2461 & n2491 ) | ( n2488 & n2491 ) ;
  assign n4261 = n4259 | n4260 ;
  assign n4262 = ( n2501 & n4259 ) | ( n2501 & n4261 ) | ( n4259 & n4261 ) ;
  assign n4263 = ( n2882 & n4261 ) | ( n2882 & n4262 ) | ( n4261 & n4262 ) ;
  assign n4264 = n566 & n4263 ;
  assign n4265 = n566 & ~n4264 ;
  assign n4266 = ( n4263 & ~n4264 ) | ( n4263 & n4265 ) | ( ~n4264 & n4265 ) ;
  assign n4267 = n4256 & n4266 ;
  assign n4268 = n4256 & ~n4267 ;
  assign n4269 = n2354 & n2563 ;
  assign n4270 = n2374 & n2559 ;
  assign n4271 = ( ~n2383 & n2384 ) | ( ~n2383 & n2557 ) | ( n2384 & n2557 ) ;
  assign n4272 = n4270 | n4271 ;
  assign n4273 = n4269 | n4272 ;
  assign n4274 = n2478 & n2586 ;
  assign n4275 = ( n977 & n4273 ) | ( n977 & n4274 ) | ( n4273 & n4274 ) ;
  assign n4276 = ( n977 & n2478 ) | ( n977 & n2589 ) | ( n2478 & n2589 ) ;
  assign n4277 = n4273 | n4276 ;
  assign n4278 = ~n4275 & n4277 ;
  assign n4279 = n4266 & ~n4267 ;
  assign n4280 = n4278 | n4279 ;
  assign n4281 = n4268 | n4280 ;
  assign n4282 = ( n4268 & n4278 ) | ( n4268 & n4279 ) | ( n4278 & n4279 ) ;
  assign n4283 = n4281 & ~n4282 ;
  assign n4284 = ( ~n4171 & n4248 ) | ( ~n4171 & n4283 ) | ( n4248 & n4283 ) ;
  assign n4285 = ( n4171 & ~n4283 ) | ( n4171 & n4284 ) | ( ~n4283 & n4284 ) ;
  assign n4286 = ( ~n4248 & n4284 ) | ( ~n4248 & n4285 ) | ( n4284 & n4285 ) ;
  assign n4287 = ( n4126 & n4127 ) | ( n4126 & n4173 ) | ( n4127 & n4173 ) ;
  assign n4288 = ( n4238 & n4286 ) | ( n4238 & ~n4287 ) | ( n4286 & ~n4287 ) ;
  assign n4289 = ( ~n4286 & n4287 ) | ( ~n4286 & n4288 ) | ( n4287 & n4288 ) ;
  assign n4290 = ( ~n4238 & n4288 ) | ( ~n4238 & n4289 ) | ( n4288 & n4289 ) ;
  assign n4291 = n4178 | n4196 ;
  assign n4292 = n4290 & n4291 ;
  assign n4293 = n4290 | n4291 ;
  assign n4294 = ~n4292 & n4293 ;
  assign n4295 = n4201 & n4294 ;
  assign n4296 = ( n4207 & n4294 ) | ( n4207 & n4295 ) | ( n4294 & n4295 ) ;
  assign n4297 = n4201 | n4294 ;
  assign n4298 = n4207 | n4297 ;
  assign n4299 = ~n4296 & n4298 ;
  assign n4300 = n336 | n2111 ;
  assign n4301 = n311 | n411 ;
  assign n4302 = n231 | n4301 ;
  assign n4303 = n360 | n654 ;
  assign n4304 = n4302 | n4303 ;
  assign n4305 = n4300 | n4304 ;
  assign n4306 = n385 | n4305 ;
  assign n4307 = n3718 | n4306 ;
  assign n4308 = n143 | n1931 ;
  assign n4309 = n3836 | n4308 ;
  assign n4310 = n180 | n369 ;
  assign n4311 = n577 | n4310 ;
  assign n4312 = n4309 | n4311 ;
  assign n4313 = n2348 | n4312 ;
  assign n4314 = n4307 | n4313 ;
  assign n4316 = ( n4299 & ~n4314 ) | ( n4299 & n4315 ) | ( ~n4314 & n4315 ) ;
  assign n4317 = ( ~n4299 & n4314 ) | ( ~n4299 & n4316 ) | ( n4314 & n4316 ) ;
  assign n4318 = ( ~n4315 & n4316 ) | ( ~n4315 & n4317 ) | ( n4316 & n4317 ) ;
  assign n4319 = n4224 | n4318 ;
  assign n4320 = n4224 & n4318 ;
  assign n4321 = n4319 & ~n4320 ;
  assign n4322 = n4225 | n4226 ;
  assign n4323 = n3859 & n4322 ;
  assign n4324 = ~n4321 & n4323 ;
  assign n4325 = n4321 & ~n4323 ;
  assign n4326 = n4324 | n4325 ;
  assign n4327 = n2381 & ~n3729 ;
  assign n4328 = n2388 & ~n3729 ;
  assign n4329 = n4327 | n4328 ;
  assign n4330 = ( ~n3590 & n4327 ) | ( ~n3590 & n4329 ) | ( n4327 & n4329 ) ;
  assign n4331 = ( n3604 & n4329 ) | ( n3604 & n4330 ) | ( n4329 & n4330 ) ;
  assign n4332 = ~n32 & n4331 ;
  assign n4333 = n32 & ~n4331 ;
  assign n4334 = n4332 | n4333 ;
  assign n4335 = n4171 & n4281 ;
  assign n4336 = ~n4282 & n4335 ;
  assign n4337 = n4283 & ~n4336 ;
  assign n4338 = n4171 & ~n4336 ;
  assign n4339 = n4337 | n4338 ;
  assign n4340 = n4248 | n4336 ;
  assign n4341 = ( n4336 & n4339 ) | ( n4336 & n4340 ) | ( n4339 & n4340 ) ;
  assign n4342 = n4334 | n4341 ;
  assign n4343 = n4334 & n4340 ;
  assign n4344 = ( n4336 & n4339 ) | ( n4336 & n4343 ) | ( n4339 & n4343 ) ;
  assign n4345 = n4342 & ~n4344 ;
  assign n4346 = n4267 | n4282 ;
  assign n4347 = n2362 & ~n4144 ;
  assign n4348 = ( n2362 & ~n2393 ) | ( n2362 & n4347 ) | ( ~n2393 & n4347 ) ;
  assign n4349 = n2393 & n4144 ;
  assign n4350 = n566 & n2393 ;
  assign n4351 = ~n4349 & n4350 ;
  assign n4352 = n4348 | n4351 ;
  assign n4353 = n4250 | n4253 ;
  assign n4354 = n4145 | n4250 ;
  assign n4355 = ( n4154 & n4353 ) | ( n4154 & n4354 ) | ( n4353 & n4354 ) ;
  assign n4356 = ~n4352 & n4355 ;
  assign n4357 = n4352 & ~n4355 ;
  assign n4358 = n4356 | n4357 ;
  assign n4359 = n2461 & n2499 ;
  assign n4360 = ( n2452 & n2456 ) | ( n2452 & n2512 ) | ( n2456 & n2512 ) ;
  assign n4361 = n4359 | n4360 ;
  assign n4362 = ( ~n2383 & n2384 ) | ( ~n2383 & n2501 ) | ( n2384 & n2501 ) ;
  assign n4363 = n4361 | n4362 ;
  assign n4364 = n2491 | n4363 ;
  assign n4365 = ( ~n2924 & n4363 ) | ( ~n2924 & n4364 ) | ( n4363 & n4364 ) ;
  assign n4366 = ~n566 & n4365 ;
  assign n4367 = n566 | n4366 ;
  assign n4368 = ( ~n4365 & n4366 ) | ( ~n4365 & n4367 ) | ( n4366 & n4367 ) ;
  assign n4369 = n4358 & n4368 ;
  assign n4370 = n4358 & ~n4369 ;
  assign n4371 = n4368 & ~n4369 ;
  assign n4372 = n2374 & n2557 ;
  assign n4373 = n2354 & n2559 ;
  assign n4374 = n4372 | n4373 ;
  assign n4375 = n2563 & ~n3119 ;
  assign n4376 = n2562 | n4375 ;
  assign n4377 = n4374 | n4376 ;
  assign n4378 = n977 & n4377 ;
  assign n4379 = n977 & n4375 ;
  assign n4380 = ( n977 & n4374 ) | ( n977 & n4379 ) | ( n4374 & n4379 ) ;
  assign n4381 = ( ~n3197 & n4378 ) | ( ~n3197 & n4380 ) | ( n4378 & n4380 ) ;
  assign n4382 = n977 | n4377 ;
  assign n4383 = n977 | n4375 ;
  assign n4384 = n4374 | n4383 ;
  assign n4385 = ( ~n3197 & n4382 ) | ( ~n3197 & n4384 ) | ( n4382 & n4384 ) ;
  assign n4386 = ~n4381 & n4385 ;
  assign n4387 = n4371 | n4386 ;
  assign n4388 = n4370 | n4387 ;
  assign n4389 = ( n4370 & n4371 ) | ( n4370 & n4386 ) | ( n4371 & n4386 ) ;
  assign n4390 = n4388 & ~n4389 ;
  assign n4391 = n2682 & ~n3590 ;
  assign n4392 = n2679 & n3147 ;
  assign n4393 = n2673 & n3162 ;
  assign n4394 = n4392 | n4393 ;
  assign n4395 = n4391 | n4394 ;
  assign n4396 = n2686 | n4395 ;
  assign n4397 = ( ~n3607 & n4395 ) | ( ~n3607 & n4396 ) | ( n4395 & n4396 ) ;
  assign n4398 = ~n752 & n4397 ;
  assign n4399 = n752 & ~n4397 ;
  assign n4400 = n4398 | n4399 ;
  assign n4401 = ( n4346 & n4390 ) | ( n4346 & n4400 ) | ( n4390 & n4400 ) ;
  assign n4402 = ( n4390 & n4400 ) | ( n4390 & ~n4401 ) | ( n4400 & ~n4401 ) ;
  assign n4403 = ( n4346 & ~n4401 ) | ( n4346 & n4402 ) | ( ~n4401 & n4402 ) ;
  assign n4404 = n4345 & n4403 ;
  assign n4405 = n4345 | n4403 ;
  assign n4406 = ~n4404 & n4405 ;
  assign n4407 = ( n4238 & n4286 ) | ( n4238 & n4287 ) | ( n4286 & n4287 ) ;
  assign n4408 = n4406 | n4407 ;
  assign n4409 = n4406 & n4407 ;
  assign n4410 = n4408 & ~n4409 ;
  assign n4411 = n4292 & n4410 ;
  assign n4412 = ( n4295 & n4410 ) | ( n4295 & n4411 ) | ( n4410 & n4411 ) ;
  assign n4413 = ( n4294 & n4410 ) | ( n4294 & n4411 ) | ( n4410 & n4411 ) ;
  assign n4414 = ( n4207 & n4412 ) | ( n4207 & n4413 ) | ( n4412 & n4413 ) ;
  assign n4415 = n4292 | n4410 ;
  assign n4416 = n4296 | n4415 ;
  assign n4417 = ~n4414 & n4416 ;
  assign n4418 = n165 | n894 ;
  assign n4419 = n2274 | n4418 ;
  assign n4420 = n3141 | n4419 ;
  assign n4421 = n3475 | n4420 ;
  assign n4422 = n504 | n865 ;
  assign n4423 = n710 | n4422 ;
  assign n4424 = n2244 | n4423 ;
  assign n4425 = n693 | n2139 ;
  assign n4426 = n900 | n1931 ;
  assign n4427 = n4425 | n4426 ;
  assign n4428 = n187 | n4427 ;
  assign n4429 = n4424 | n4428 ;
  assign n4430 = n380 | n4429 ;
  assign n4431 = n4421 | n4430 ;
  assign n4432 = n125 | n209 ;
  assign n4433 = n920 | n4432 ;
  assign n4434 = n186 | n4433 ;
  assign n4435 = n4431 | n4434 ;
  assign n4436 = n4417 | n4435 ;
  assign n4437 = n4417 & n4435 ;
  assign n4438 = n4436 & ~n4437 ;
  assign n4439 = n4299 | n4314 ;
  assign n4440 = n4299 & n4314 ;
  assign n4441 = ( n4315 & n4439 ) | ( n4315 & n4440 ) | ( n4439 & n4440 ) ;
  assign n4442 = n4438 & n4441 ;
  assign n4443 = n4438 | n4441 ;
  assign n4444 = ~n4442 & n4443 ;
  assign n4445 = n4318 & n4444 ;
  assign n4446 = n4224 & n4445 ;
  assign n4447 = n4320 | n4444 ;
  assign n4448 = ~n4446 & n4447 ;
  assign n4449 = ( n3859 & n4321 ) | ( n3859 & n4323 ) | ( n4321 & n4323 ) ;
  assign n4450 = ~n4448 & n4449 ;
  assign n4451 = n4448 & ~n4449 ;
  assign n4452 = n4450 | n4451 ;
  assign n4453 = n191 | n405 ;
  assign n4454 = n223 | n4453 ;
  assign n4455 = n135 | n201 ;
  assign n4456 = n4454 | n4455 ;
  assign n4457 = n597 | n4456 ;
  assign n4458 = n141 | n4429 ;
  assign n4459 = n247 | n847 ;
  assign n4460 = n4302 | n4459 ;
  assign n4461 = n465 | n4460 ;
  assign n4462 = ( ~n2062 & n4458 ) | ( ~n2062 & n4461 ) | ( n4458 & n4461 ) ;
  assign n4463 = n2062 | n4462 ;
  assign n4464 = n4457 | n4463 ;
  assign n4465 = n4437 | n4442 ;
  assign n4466 = n4344 | n4404 ;
  assign n4467 = n2679 & n3162 ;
  assign n4468 = n2673 & ~n3590 ;
  assign n4469 = n4467 | n4468 ;
  assign n4470 = ( n2669 & n2686 ) | ( n2669 & ~n3729 ) | ( n2686 & ~n3729 ) ;
  assign n4471 = n4469 | n4470 ;
  assign n4472 = ( n2682 & n4469 ) | ( n2682 & n4471 ) | ( n4469 & n4471 ) ;
  assign n4473 = ( n3742 & n4471 ) | ( n3742 & n4472 ) | ( n4471 & n4472 ) ;
  assign n4474 = n752 & n4473 ;
  assign n4475 = n752 & ~n4474 ;
  assign n4476 = ( n4473 & ~n4474 ) | ( n4473 & n4475 ) | ( ~n4474 & n4475 ) ;
  assign n4477 = n4401 & n4476 ;
  assign n4478 = n4401 | n4476 ;
  assign n4479 = ~n4477 & n4478 ;
  assign n4480 = n4369 | n4389 ;
  assign n4481 = n2374 & n2501 ;
  assign n4482 = n2461 & n2512 ;
  assign n4483 = ( ~n2383 & n2384 ) | ( ~n2383 & n2499 ) | ( n2384 & n2499 ) ;
  assign n4484 = n4482 | n4483 ;
  assign n4485 = n4481 | n4484 ;
  assign n4486 = n2491 | n4485 ;
  assign n4487 = ( ~n2908 & n4485 ) | ( ~n2908 & n4486 ) | ( n4485 & n4486 ) ;
  assign n4488 = ~n566 & n4487 ;
  assign n4489 = n566 & n2452 ;
  assign n4490 = ( n566 & n2456 ) | ( n566 & n4489 ) | ( n2456 & n4489 ) ;
  assign n4491 = ( n32 & ~n2362 ) | ( n32 & n4490 ) | ( ~n2362 & n4490 ) ;
  assign n4492 = ( ~n32 & n2362 ) | ( ~n32 & n4491 ) | ( n2362 & n4491 ) ;
  assign n4493 = ( ~n4490 & n4491 ) | ( ~n4490 & n4492 ) | ( n4491 & n4492 ) ;
  assign n4494 = n566 & ~n4487 ;
  assign n4495 = n4493 & ~n4494 ;
  assign n4496 = ~n4488 & n4495 ;
  assign n4497 = ( n4488 & ~n4493 ) | ( n4488 & n4494 ) | ( ~n4493 & n4494 ) ;
  assign n4498 = n4496 | n4497 ;
  assign n4499 = n4352 & n4354 ;
  assign n4500 = n4352 & n4353 ;
  assign n4501 = ( n4154 & n4499 ) | ( n4154 & n4500 ) | ( n4499 & n4500 ) ;
  assign n4502 = n4349 | n4501 ;
  assign n4503 = n4498 | n4502 ;
  assign n4504 = ~n4502 & n4503 ;
  assign n4505 = ( ~n4498 & n4503 ) | ( ~n4498 & n4504 ) | ( n4503 & n4504 ) ;
  assign n4506 = n2354 & n2557 ;
  assign n4507 = n2559 & ~n3119 ;
  assign n4508 = n4506 | n4507 ;
  assign n4509 = ( n2549 & n2562 ) | ( n2549 & n3147 ) | ( n2562 & n3147 ) ;
  assign n4510 = n4508 | n4509 ;
  assign n4511 = ( n2563 & n4508 ) | ( n2563 & n4510 ) | ( n4508 & n4510 ) ;
  assign n4512 = ( ~n3447 & n4510 ) | ( ~n3447 & n4511 ) | ( n4510 & n4511 ) ;
  assign n4513 = ~n977 & n4512 ;
  assign n4514 = n977 | n4513 ;
  assign n4515 = ( ~n4512 & n4513 ) | ( ~n4512 & n4514 ) | ( n4513 & n4514 ) ;
  assign n4516 = n4505 & n4515 ;
  assign n4517 = n4515 & ~n4516 ;
  assign n4518 = ( n4505 & ~n4516 ) | ( n4505 & n4517 ) | ( ~n4516 & n4517 ) ;
  assign n4519 = n4480 & n4518 ;
  assign n4520 = n4480 | n4518 ;
  assign n4521 = ~n4519 & n4520 ;
  assign n4522 = ( n4466 & n4479 ) | ( n4466 & ~n4521 ) | ( n4479 & ~n4521 ) ;
  assign n4523 = ( ~n4479 & n4521 ) | ( ~n4479 & n4522 ) | ( n4521 & n4522 ) ;
  assign n4524 = ( ~n4466 & n4522 ) | ( ~n4466 & n4523 ) | ( n4522 & n4523 ) ;
  assign n4525 = n4409 | n4412 ;
  assign n4526 = n4524 & n4525 ;
  assign n4527 = ( n4409 & n4413 ) | ( n4409 & n4524 ) | ( n4413 & n4524 ) ;
  assign n4528 = ( n4207 & n4526 ) | ( n4207 & n4527 ) | ( n4526 & n4527 ) ;
  assign n4529 = n4524 | n4525 ;
  assign n4530 = n4409 | n4524 ;
  assign n4531 = n4413 | n4530 ;
  assign n4532 = ( n4207 & n4529 ) | ( n4207 & n4531 ) | ( n4529 & n4531 ) ;
  assign n4533 = ~n4528 & n4532 ;
  assign n4534 = ( n4464 & n4465 ) | ( n4464 & ~n4533 ) | ( n4465 & ~n4533 ) ;
  assign n4535 = ( ~n4465 & n4533 ) | ( ~n4465 & n4534 ) | ( n4533 & n4534 ) ;
  assign n4536 = ( ~n4464 & n4534 ) | ( ~n4464 & n4535 ) | ( n4534 & n4535 ) ;
  assign n4537 = n4446 & n4536 ;
  assign n4538 = n4446 | n4536 ;
  assign n4539 = ~n4537 & n4538 ;
  assign n4540 = n4321 | n4448 ;
  assign n4541 = n4322 | n4540 ;
  assign n4542 = n3859 & n4541 ;
  assign n4543 = ~n4539 & n4542 ;
  assign n4544 = n4539 & ~n4542 ;
  assign n4545 = n4543 | n4544 ;
  assign n4546 = n201 | n902 ;
  assign n4547 = n921 | n2138 ;
  assign n4548 = n4546 | n4547 ;
  assign n4549 = n3521 | n4548 ;
  assign n4550 = n3544 | n4549 ;
  assign n4551 = n161 | n502 ;
  assign n4552 = n701 | n4551 ;
  assign n4553 = n699 | n4552 ;
  assign n4554 = n249 | n384 ;
  assign n4555 = n226 | n362 ;
  assign n4556 = n4554 | n4555 ;
  assign n4557 = n292 | n4556 ;
  assign n4558 = n477 | n4557 ;
  assign n4559 = n4553 | n4558 ;
  assign n4560 = n4550 | n4559 ;
  assign n4561 = n108 | n349 ;
  assign n4562 = n120 | n205 ;
  assign n4563 = n4561 | n4562 ;
  assign n4564 = n267 | n1976 ;
  assign n4565 = n4563 | n4564 ;
  assign n4566 = n4560 | n4565 ;
  assign n4567 = n4479 & n4521 ;
  assign n4568 = n4479 & ~n4567 ;
  assign n4569 = ( n4466 & ~n4522 ) | ( n4466 & n4568 ) | ( ~n4522 & n4568 ) ;
  assign n4570 = n4527 | n4569 ;
  assign n4571 = ( n4525 & n4569 ) | ( n4525 & n4570 ) | ( n4569 & n4570 ) ;
  assign n4572 = ( n4207 & n4570 ) | ( n4207 & n4571 ) | ( n4570 & n4571 ) ;
  assign n4573 = n4477 | n4567 ;
  assign n4574 = ( n4493 & n4497 ) | ( n4493 & ~n4504 ) | ( n4497 & ~n4504 ) ;
  assign n4575 = n2354 & n2501 ;
  assign n4576 = n2374 & n2499 ;
  assign n4577 = ( ~n2383 & n2384 ) | ( ~n2383 & n2512 ) | ( n2384 & n2512 ) ;
  assign n4578 = n4576 | n4577 ;
  assign n4579 = n4575 | n4578 ;
  assign n4580 = n566 | n4579 ;
  assign n4581 = ( n2478 & n2491 ) | ( n2478 & n4580 ) | ( n2491 & n4580 ) ;
  assign n4582 = n4580 | n4581 ;
  assign n4583 = n2478 & n4141 ;
  assign n4584 = ( n566 & n4579 ) | ( n566 & n4583 ) | ( n4579 & n4583 ) ;
  assign n4585 = n4582 & ~n4584 ;
  assign n4586 = n32 | n2362 ;
  assign n4587 = n32 & n2362 ;
  assign n4588 = ( ~n4489 & n4586 ) | ( ~n4489 & n4587 ) | ( n4586 & n4587 ) ;
  assign n4589 = ( ~n566 & n4586 ) | ( ~n566 & n4587 ) | ( n4586 & n4587 ) ;
  assign n4590 = ( ~n2456 & n4588 ) | ( ~n2456 & n4589 ) | ( n4588 & n4589 ) ;
  assign n4591 = n566 & n2461 ;
  assign n4592 = ( n4585 & n4590 ) | ( n4585 & ~n4591 ) | ( n4590 & ~n4591 ) ;
  assign n4593 = ( ~n4590 & n4591 ) | ( ~n4590 & n4592 ) | ( n4591 & n4592 ) ;
  assign n4594 = ( ~n4585 & n4592 ) | ( ~n4585 & n4593 ) | ( n4592 & n4593 ) ;
  assign n4595 = n4574 & n4594 ;
  assign n4596 = n4574 & ~n4595 ;
  assign n4597 = n2557 & ~n3119 ;
  assign n4598 = n2559 & n3147 ;
  assign n4599 = n4597 | n4598 ;
  assign n4600 = n2563 & n3162 ;
  assign n4601 = n2562 | n4600 ;
  assign n4602 = n4599 | n4601 ;
  assign n4603 = n977 & n4602 ;
  assign n4604 = n977 & n4600 ;
  assign n4605 = ( n977 & n4599 ) | ( n977 & n4604 ) | ( n4599 & n4604 ) ;
  assign n4606 = ( n3182 & n4603 ) | ( n3182 & n4605 ) | ( n4603 & n4605 ) ;
  assign n4607 = n977 | n4602 ;
  assign n4608 = n977 | n4600 ;
  assign n4609 = n4599 | n4608 ;
  assign n4610 = ( n3182 & n4607 ) | ( n3182 & n4609 ) | ( n4607 & n4609 ) ;
  assign n4611 = ~n4606 & n4610 ;
  assign n4612 = ~n4574 & n4594 ;
  assign n4613 = n4611 | n4612 ;
  assign n4614 = n4596 | n4613 ;
  assign n4615 = ( n4596 & n4611 ) | ( n4596 & n4612 ) | ( n4611 & n4612 ) ;
  assign n4616 = n4614 & ~n4615 ;
  assign n4617 = n2679 & ~n3590 ;
  assign n4618 = n2673 & ~n3729 ;
  assign n4619 = n4617 | n4618 ;
  assign n4620 = ( n752 & n2791 ) | ( n752 & ~n3875 ) | ( n2791 & ~n3875 ) ;
  assign n4621 = ~n4619 & n4620 ;
  assign n4622 = n2686 | n4619 ;
  assign n4623 = ( n3875 & n4619 ) | ( n3875 & n4622 ) | ( n4619 & n4622 ) ;
  assign n4624 = ~n752 & n4623 ;
  assign n4625 = n4621 | n4624 ;
  assign n4626 = n4516 | n4519 ;
  assign n4627 = ( n4616 & n4625 ) | ( n4616 & ~n4626 ) | ( n4625 & ~n4626 ) ;
  assign n4628 = ( ~n4625 & n4626 ) | ( ~n4625 & n4627 ) | ( n4626 & n4627 ) ;
  assign n4629 = ( ~n4616 & n4627 ) | ( ~n4616 & n4628 ) | ( n4627 & n4628 ) ;
  assign n4630 = n4573 & n4629 ;
  assign n4631 = n4573 | n4629 ;
  assign n4632 = ~n4630 & n4631 ;
  assign n4633 = n4572 & n4632 ;
  assign n4634 = n4632 & ~n4633 ;
  assign n4635 = ( n4572 & ~n4633 ) | ( n4572 & n4634 ) | ( ~n4633 & n4634 ) ;
  assign n4636 = n4566 | n4635 ;
  assign n4637 = n4566 & n4635 ;
  assign n4638 = n4636 & ~n4637 ;
  assign n4639 = n4464 | n4533 ;
  assign n4640 = ( n4437 & n4464 ) | ( n4437 & n4533 ) | ( n4464 & n4533 ) ;
  assign n4641 = ( n4442 & n4639 ) | ( n4442 & n4640 ) | ( n4639 & n4640 ) ;
  assign n4642 = n4638 | n4641 ;
  assign n4643 = n4638 & n4641 ;
  assign n4644 = n4642 & ~n4643 ;
  assign n4645 = n4536 & n4644 ;
  assign n4646 = n4446 & n4645 ;
  assign n4647 = n4537 | n4644 ;
  assign n4648 = ~n4646 & n4647 ;
  assign n4649 = ( n3859 & n4539 ) | ( n3859 & n4542 ) | ( n4539 & n4542 ) ;
  assign n4650 = ~n4648 & n4649 ;
  assign n4651 = n4648 & ~n4649 ;
  assign n4652 = n4650 | n4651 ;
  assign n4653 = n2679 & ~n3729 ;
  assign n4654 = n2686 & ~n3729 ;
  assign n4655 = n4653 | n4654 ;
  assign n4656 = ( ~n3590 & n4653 ) | ( ~n3590 & n4655 ) | ( n4653 & n4655 ) ;
  assign n4657 = ( n3604 & n4655 ) | ( n3604 & n4656 ) | ( n4655 & n4656 ) ;
  assign n4658 = n752 & ~n4657 ;
  assign n4659 = ~n752 & n4657 ;
  assign n4660 = n4658 | n4659 ;
  assign n4661 = n4595 | n4660 ;
  assign n4662 = n4615 | n4661 ;
  assign n4663 = ( n4595 & n4615 ) | ( n4595 & n4660 ) | ( n4615 & n4660 ) ;
  assign n4664 = n4662 & ~n4663 ;
  assign n4665 = n2557 & n3147 ;
  assign n4666 = n2559 & n3162 ;
  assign n4667 = n4665 | n4666 ;
  assign n4668 = n2563 & ~n3590 ;
  assign n4669 = n2562 | n4668 ;
  assign n4670 = n4667 | n4669 ;
  assign n4671 = n977 & n4670 ;
  assign n4672 = n977 & n4668 ;
  assign n4673 = ( n977 & n4667 ) | ( n977 & n4672 ) | ( n4667 & n4672 ) ;
  assign n4674 = ( ~n3607 & n4671 ) | ( ~n3607 & n4673 ) | ( n4671 & n4673 ) ;
  assign n4675 = n977 | n4670 ;
  assign n4676 = n977 | n4668 ;
  assign n4677 = n4667 | n4676 ;
  assign n4678 = ( ~n3607 & n4675 ) | ( ~n3607 & n4677 ) | ( n4675 & n4677 ) ;
  assign n4679 = ~n4674 & n4678 ;
  assign n4680 = ( ~n4585 & n4590 ) | ( ~n4585 & n4591 ) | ( n4590 & n4591 ) ;
  assign n4681 = n566 & ~n2921 ;
  assign n4682 = n2501 & ~n3119 ;
  assign n4683 = n2374 & n2512 ;
  assign n4684 = n2354 & n2499 ;
  assign n4685 = n4683 | n4684 ;
  assign n4686 = n4682 | n4685 ;
  assign n4687 = n2491 | n4686 ;
  assign n4688 = ( ~n3197 & n4686 ) | ( ~n3197 & n4687 ) | ( n4686 & n4687 ) ;
  assign n4689 = n566 & ~n4688 ;
  assign n4690 = ~n4681 & n4689 ;
  assign n4691 = ~n566 & n4688 ;
  assign n4692 = ( ~n4681 & n4690 ) | ( ~n4681 & n4691 ) | ( n4690 & n4691 ) ;
  assign n4693 = ( ~n2921 & n4688 ) | ( ~n2921 & n4692 ) | ( n4688 & n4692 ) ;
  assign n4694 = ( n566 & n4692 ) | ( n566 & n4693 ) | ( n4692 & n4693 ) ;
  assign n4695 = ( n4679 & ~n4680 ) | ( n4679 & n4694 ) | ( ~n4680 & n4694 ) ;
  assign n4696 = ( n4680 & ~n4694 ) | ( n4680 & n4695 ) | ( ~n4694 & n4695 ) ;
  assign n4697 = ( ~n4679 & n4695 ) | ( ~n4679 & n4696 ) | ( n4695 & n4696 ) ;
  assign n4698 = n4664 & ~n4697 ;
  assign n4699 = n4697 | n4698 ;
  assign n4700 = ( ~n4664 & n4698 ) | ( ~n4664 & n4699 ) | ( n4698 & n4699 ) ;
  assign n4701 = ( n4616 & n4625 ) | ( n4616 & n4626 ) | ( n4625 & n4626 ) ;
  assign n4702 = n4700 & n4701 ;
  assign n4703 = n4701 & ~n4702 ;
  assign n4704 = ( n4700 & ~n4702 ) | ( n4700 & n4703 ) | ( ~n4702 & n4703 ) ;
  assign n4705 = n4630 & n4704 ;
  assign n4706 = ( n4632 & n4704 ) | ( n4632 & n4705 ) | ( n4704 & n4705 ) ;
  assign n4707 = ( n4572 & n4705 ) | ( n4572 & n4706 ) | ( n4705 & n4706 ) ;
  assign n4708 = n4630 | n4704 ;
  assign n4709 = n4633 | n4708 ;
  assign n4710 = ~n4707 & n4709 ;
  assign n4711 = n281 | n2336 ;
  assign n4712 = n465 | n585 ;
  assign n4713 = n4711 | n4712 ;
  assign n4714 = n3141 | n4713 ;
  assign n4715 = n3479 | n4714 ;
  assign n4716 = n2254 | n4715 ;
  assign n4717 = n204 | n380 ;
  assign n4718 = n112 | n362 ;
  assign n4719 = n4717 | n4718 ;
  assign n4720 = n152 | n457 ;
  assign n4721 = n297 | n4720 ;
  assign n4722 = n4719 | n4721 ;
  assign n4723 = n4716 | n4722 ;
  assign n4724 = n4710 | n4723 ;
  assign n4725 = n4710 & n4723 ;
  assign n4726 = n4724 & ~n4725 ;
  assign n4727 = n4637 | n4726 ;
  assign n4728 = n4643 | n4727 ;
  assign n4729 = n4637 & n4726 ;
  assign n4730 = ( n4643 & n4726 ) | ( n4643 & n4729 ) | ( n4726 & n4729 ) ;
  assign n4731 = n4728 & ~n4730 ;
  assign n4732 = n4646 | n4731 ;
  assign n4733 = n4646 & n4731 ;
  assign n4734 = n4732 & ~n4733 ;
  assign n4735 = n4539 | n4648 ;
  assign n4736 = n4541 | n4735 ;
  assign n4737 = n3859 & n4736 ;
  assign n4738 = ~n4734 & n4737 ;
  assign n4739 = n4734 & ~n4737 ;
  assign n4740 = n4738 | n4739 ;
  assign n4741 = ( ~n4679 & n4680 ) | ( ~n4679 & n4694 ) | ( n4680 & n4694 ) ;
  assign n4742 = n2557 & n3162 ;
  assign n4743 = n2559 & ~n3590 ;
  assign n4744 = n4742 | n4743 ;
  assign n4745 = ( n2549 & n2562 ) | ( n2549 & ~n3729 ) | ( n2562 & ~n3729 ) ;
  assign n4746 = n4744 | n4745 ;
  assign n4747 = ( n2563 & n4744 ) | ( n2563 & n4746 ) | ( n4744 & n4746 ) ;
  assign n4748 = ( n3742 & n4746 ) | ( n3742 & n4747 ) | ( n4746 & n4747 ) ;
  assign n4749 = n977 & n4748 ;
  assign n4750 = n977 & ~n4749 ;
  assign n4751 = ( n4748 & ~n4749 ) | ( n4748 & n4750 ) | ( ~n4749 & n4750 ) ;
  assign n4752 = ~n4741 & n4751 ;
  assign n4753 = n4741 | n4752 ;
  assign n4754 = n4741 & n4751 ;
  assign n4755 = n2501 & n3147 ;
  assign n4756 = n2354 & n2512 ;
  assign n4757 = n2499 & ~n3119 ;
  assign n4758 = n4756 | n4757 ;
  assign n4759 = n4755 | n4758 ;
  assign n4760 = n2491 | n4759 ;
  assign n4761 = ( ~n3447 & n4759 ) | ( ~n3447 & n4760 ) | ( n4759 & n4760 ) ;
  assign n4762 = ~n566 & n4761 ;
  assign n4763 = n566 & ~n4761 ;
  assign n4764 = n4762 | n4763 ;
  assign n4765 = ~n566 & n752 ;
  assign n4766 = ( n752 & ~n2374 ) | ( n752 & n4765 ) | ( ~n2374 & n4765 ) ;
  assign n4767 = n566 & ~n752 ;
  assign n4768 = n2374 & n4767 ;
  assign n4769 = ( n4591 & ~n4766 ) | ( n4591 & n4768 ) | ( ~n4766 & n4768 ) ;
  assign n4770 = n4766 | n4769 ;
  assign n4771 = ( n4591 & n4766 ) | ( n4591 & n4768 ) | ( n4766 & n4768 ) ;
  assign n4772 = n4770 & ~n4771 ;
  assign n4773 = ~n2468 & n4681 ;
  assign n4774 = ~n4772 & n4773 ;
  assign n4775 = n4772 | n4774 ;
  assign n4776 = n4692 | n4775 ;
  assign n4777 = ( n4692 & n4772 ) | ( n4692 & n4773 ) | ( n4772 & n4773 ) ;
  assign n4778 = n4776 & ~n4777 ;
  assign n4779 = n4764 | n4778 ;
  assign n4780 = ( n4764 & ~n4776 ) | ( n4764 & n4777 ) | ( ~n4776 & n4777 ) ;
  assign n4781 = ( ~n4764 & n4779 ) | ( ~n4764 & n4780 ) | ( n4779 & n4780 ) ;
  assign n4782 = ~n4754 & n4781 ;
  assign n4783 = n4753 & n4782 ;
  assign n4784 = ( n4753 & ~n4754 ) | ( n4753 & n4781 ) | ( ~n4754 & n4781 ) ;
  assign n4785 = ~n4783 & n4784 ;
  assign n4786 = ( n4662 & n4663 ) | ( n4662 & n4697 ) | ( n4663 & n4697 ) ;
  assign n4787 = n4785 & n4786 ;
  assign n4788 = n4785 | n4786 ;
  assign n4789 = ~n4787 & n4788 ;
  assign n4790 = n4702 & n4789 ;
  assign n4791 = ( n4706 & n4789 ) | ( n4706 & n4790 ) | ( n4789 & n4790 ) ;
  assign n4792 = ( n4705 & n4789 ) | ( n4705 & n4790 ) | ( n4789 & n4790 ) ;
  assign n4793 = ( n4572 & n4791 ) | ( n4572 & n4792 ) | ( n4791 & n4792 ) ;
  assign n4794 = n4702 | n4789 ;
  assign n4795 = n4707 | n4794 ;
  assign n4796 = ~n4793 & n4795 ;
  assign n4797 = n554 | n3141 ;
  assign n4798 = n179 | n1948 ;
  assign n4799 = n130 | n4798 ;
  assign n4800 = n298 | n4799 ;
  assign n4801 = n790 | n4800 ;
  assign n4802 = n2327 | n3534 ;
  assign n4803 = n4801 | n4802 ;
  assign n4804 = n4797 | n4803 ;
  assign n4805 = n381 | n399 ;
  assign n4806 = n900 | n4805 ;
  assign n4807 = n195 | n391 ;
  assign n4808 = n4806 | n4807 ;
  assign n4809 = n4804 | n4808 ;
  assign n4810 = n4796 | n4809 ;
  assign n4811 = n4796 & n4809 ;
  assign n4812 = n4810 & ~n4811 ;
  assign n4813 = n4725 | n4729 ;
  assign n4814 = ( n4643 & n4724 ) | ( n4643 & n4813 ) | ( n4724 & n4813 ) ;
  assign n4815 = n4812 & n4814 ;
  assign n4816 = n4812 | n4814 ;
  assign n4817 = ~n4815 & n4816 ;
  assign n4818 = n4731 & n4817 ;
  assign n4819 = n4646 & n4818 ;
  assign n4820 = n4733 | n4817 ;
  assign n4821 = ~n4819 & n4820 ;
  assign n4822 = ( n3859 & n4734 ) | ( n3859 & n4737 ) | ( n4734 & n4737 ) ;
  assign n4823 = ~n4821 & n4822 ;
  assign n4824 = n4821 & ~n4822 ;
  assign n4825 = n4823 | n4824 ;
  assign n4826 = n4734 | n4821 ;
  assign n4827 = n4736 | n4826 ;
  assign n4828 = n3859 & n4827 ;
  assign n4829 = n4787 | n4790 ;
  assign n4830 = ( n4705 & n4788 ) | ( n4705 & n4829 ) | ( n4788 & n4829 ) ;
  assign n4831 = ( n4706 & n4788 ) | ( n4706 & n4829 ) | ( n4788 & n4829 ) ;
  assign n4832 = ( n4572 & n4830 ) | ( n4572 & n4831 ) | ( n4830 & n4831 ) ;
  assign n4833 = ~n4752 & n4784 ;
  assign n4834 = n2557 & ~n3590 ;
  assign n4835 = n2559 & ~n3729 ;
  assign n4836 = n4834 | n4835 ;
  assign n4837 = n2586 & n3875 ;
  assign n4838 = ( n977 & n4836 ) | ( n977 & n4837 ) | ( n4836 & n4837 ) ;
  assign n4839 = ( n977 & n2589 ) | ( n977 & n3875 ) | ( n2589 & n3875 ) ;
  assign n4840 = n4836 | n4839 ;
  assign n4841 = ~n4838 & n4840 ;
  assign n4842 = n566 & n2354 ;
  assign n4843 = n4769 & ~n4842 ;
  assign n4844 = ( ~n4769 & n4842 ) | ( ~n4769 & n4843 ) | ( n4842 & n4843 ) ;
  assign n4845 = ( n566 & n4843 ) | ( n566 & n4844 ) | ( n4843 & n4844 ) ;
  assign n4846 = n2512 & ~n3119 ;
  assign n4847 = n2499 & n3147 ;
  assign n4848 = n4846 | n4847 ;
  assign n4849 = ( n2488 & n2491 ) | ( n2488 & n3162 ) | ( n2491 & n3162 ) ;
  assign n4850 = n4848 | n4849 ;
  assign n4851 = ( n2501 & n4848 ) | ( n2501 & n4850 ) | ( n4848 & n4850 ) ;
  assign n4852 = ( n3182 & n4850 ) | ( n3182 & n4851 ) | ( n4850 & n4851 ) ;
  assign n4853 = n566 & n4852 ;
  assign n4854 = n566 & ~n4853 ;
  assign n4855 = ( n4852 & ~n4853 ) | ( n4852 & n4854 ) | ( ~n4853 & n4854 ) ;
  assign n4856 = ~n4845 & n4855 ;
  assign n4857 = n4845 & ~n4855 ;
  assign n4858 = n4856 | n4857 ;
  assign n4859 = ( n4691 & ~n4772 ) | ( n4691 & n4778 ) | ( ~n4772 & n4778 ) ;
  assign n4860 = n4780 | n4859 ;
  assign n4861 = ( n4841 & n4858 ) | ( n4841 & ~n4860 ) | ( n4858 & ~n4860 ) ;
  assign n4862 = ( ~n4858 & n4860 ) | ( ~n4858 & n4861 ) | ( n4860 & n4861 ) ;
  assign n4863 = ( ~n4841 & n4861 ) | ( ~n4841 & n4862 ) | ( n4861 & n4862 ) ;
  assign n4864 = n4833 | n4863 ;
  assign n4865 = n4833 & n4863 ;
  assign n4866 = n4864 & ~n4865 ;
  assign n4867 = n4832 & n4866 ;
  assign n4868 = n4866 & ~n4867 ;
  assign n4869 = ( n4832 & ~n4867 ) | ( n4832 & n4868 ) | ( ~n4867 & n4868 ) ;
  assign n4870 = n4811 | n4815 ;
  assign n4871 = n195 | n308 ;
  assign n4872 = n875 | n893 ;
  assign n4873 = n4871 | n4872 ;
  assign n4874 = n3573 | n4873 ;
  assign n4875 = n287 | n804 ;
  assign n4876 = n4874 | n4875 ;
  assign n4877 = n783 | n4876 ;
  assign n4878 = n211 | n4877 ;
  assign n4879 = ( n4869 & n4870 ) | ( n4869 & ~n4878 ) | ( n4870 & ~n4878 ) ;
  assign n4880 = ( ~n4870 & n4878 ) | ( ~n4870 & n4879 ) | ( n4878 & n4879 ) ;
  assign n4881 = ( ~n4869 & n4879 ) | ( ~n4869 & n4880 ) | ( n4879 & n4880 ) ;
  assign n4882 = n4819 & ~n4881 ;
  assign n4883 = n4881 | n4882 ;
  assign n4884 = ( ~n4819 & n4882 ) | ( ~n4819 & n4883 ) | ( n4882 & n4883 ) ;
  assign n4885 = n4828 & ~n4884 ;
  assign n4886 = ~n4828 & n4884 ;
  assign n4887 = n4885 | n4886 ;
  assign n4888 = n171 | n257 ;
  assign n4889 = n205 | n457 ;
  assign n4890 = n4888 | n4889 ;
  assign n4891 = n132 | n2179 ;
  assign n4892 = n4890 | n4891 ;
  assign n4893 = n837 | n4892 ;
  assign n4894 = n3962 | n4893 ;
  assign n4895 = n2017 | n4894 ;
  assign n4896 = n1936 | n1939 ;
  assign n4897 = n1935 | n4896 ;
  assign n4898 = n386 | n4897 ;
  assign n4899 = n253 | n477 ;
  assign n4900 = n4898 | n4899 ;
  assign n4901 = n4895 | n4900 ;
  assign n4902 = n4869 | n4878 ;
  assign n4903 = ( n4811 & n4869 ) | ( n4811 & n4878 ) | ( n4869 & n4878 ) ;
  assign n4904 = ( n4815 & n4902 ) | ( n4815 & n4903 ) | ( n4902 & n4903 ) ;
  assign n4905 = n4831 & n4866 ;
  assign n4906 = n566 & ~n3119 ;
  assign n4907 = ~n4842 & n4906 ;
  assign n4908 = n4842 & ~n4906 ;
  assign n4909 = ( n4856 & n4907 ) | ( n4856 & n4908 ) | ( n4907 & n4908 ) ;
  assign n4910 = ( n4769 & n4907 ) | ( n4769 & n4909 ) | ( n4907 & n4909 ) ;
  assign n4911 = n4907 | n4908 ;
  assign n4912 = ( n4769 & ~n4906 ) | ( n4769 & n4908 ) | ( ~n4906 & n4908 ) ;
  assign n4913 = ( n4844 & n4907 ) | ( n4844 & ~n4908 ) | ( n4907 & ~n4908 ) ;
  assign n4914 = ( n4855 & n4912 ) | ( n4855 & ~n4913 ) | ( n4912 & ~n4913 ) ;
  assign n4915 = n4911 | n4914 ;
  assign n4916 = ~n4910 & n4915 ;
  assign n4917 = n2501 & ~n3590 ;
  assign n4918 = n2512 & n3147 ;
  assign n4919 = n2499 & n3162 ;
  assign n4920 = n4918 | n4919 ;
  assign n4921 = n4917 | n4920 ;
  assign n4922 = n2491 | n4921 ;
  assign n4923 = ( ~n3607 & n4921 ) | ( ~n3607 & n4922 ) | ( n4921 & n4922 ) ;
  assign n4924 = ~n566 & n4923 ;
  assign n4925 = n566 & ~n4923 ;
  assign n4926 = n4924 | n4925 ;
  assign n4927 = n2557 & ~n3729 ;
  assign n4928 = n2562 & ~n3729 ;
  assign n4929 = n4927 | n4928 ;
  assign n4930 = ( ~n3590 & n4927 ) | ( ~n3590 & n4929 ) | ( n4927 & n4929 ) ;
  assign n4931 = ( n3604 & n4929 ) | ( n3604 & n4930 ) | ( n4929 & n4930 ) ;
  assign n4932 = n977 & n4931 ;
  assign n4933 = n977 | n4931 ;
  assign n4934 = ~n4932 & n4933 ;
  assign n4935 = n4926 | n4934 ;
  assign n4936 = ~n4934 & n4935 ;
  assign n4937 = ( ~n4926 & n4935 ) | ( ~n4926 & n4936 ) | ( n4935 & n4936 ) ;
  assign n4938 = n4916 & n4937 ;
  assign n4939 = n4916 | n4937 ;
  assign n4940 = ~n4938 & n4939 ;
  assign n4941 = n4862 & ~n4940 ;
  assign n4942 = ~n4862 & n4940 ;
  assign n4943 = n4941 | n4942 ;
  assign n4944 = n4864 | n4943 ;
  assign n4945 = ( ~n4905 & n4943 ) | ( ~n4905 & n4944 ) | ( n4943 & n4944 ) ;
  assign n4946 = n4865 | n4943 ;
  assign n4947 = ( ~n4830 & n4944 ) | ( ~n4830 & n4946 ) | ( n4944 & n4946 ) ;
  assign n4948 = ( ~n4572 & n4945 ) | ( ~n4572 & n4947 ) | ( n4945 & n4947 ) ;
  assign n4949 = n4864 & n4943 ;
  assign n4950 = ~n4905 & n4949 ;
  assign n4951 = n4865 & n4943 ;
  assign n4952 = ( ~n4830 & n4949 ) | ( ~n4830 & n4951 ) | ( n4949 & n4951 ) ;
  assign n4953 = ( ~n4572 & n4950 ) | ( ~n4572 & n4952 ) | ( n4950 & n4952 ) ;
  assign n4954 = ( n4950 & n4952 ) | ( n4950 & n4953 ) | ( n4952 & n4953 ) ;
  assign n4955 = n4948 & ~n4954 ;
  assign n4956 = ( n4901 & n4904 ) | ( n4901 & ~n4955 ) | ( n4904 & ~n4955 ) ;
  assign n4957 = ( ~n4904 & n4955 ) | ( ~n4904 & n4956 ) | ( n4955 & n4956 ) ;
  assign n4958 = ( ~n4901 & n4956 ) | ( ~n4901 & n4957 ) | ( n4956 & n4957 ) ;
  assign n4959 = n4881 & n4958 ;
  assign n4960 = n4819 & n4959 ;
  assign n4961 = ( n4819 & ~n4882 ) | ( n4819 & n4958 ) | ( ~n4882 & n4958 ) ;
  assign n4962 = ~n4960 & n4961 ;
  assign n4963 = ( n3859 & n4828 ) | ( n3859 & n4884 ) | ( n4828 & n4884 ) ;
  assign n4964 = ~n4962 & n4963 ;
  assign n4965 = n4962 & ~n4963 ;
  assign n4966 = n4964 | n4965 ;
  assign n4967 = n405 | n544 ;
  assign n4968 = n274 | n367 ;
  assign n4969 = n4967 | n4968 ;
  assign n4970 = n305 | n693 ;
  assign n4971 = n4969 | n4970 ;
  assign n4972 = n3836 | n4971 ;
  assign n4973 = n534 | n4972 ;
  assign n4974 = n244 | n543 ;
  assign n4975 = n4973 | n4974 ;
  assign n4976 = n147 | n3501 ;
  assign n4977 = n4975 | n4976 ;
  assign n4978 = n108 | n265 ;
  assign n4979 = n116 | n173 ;
  assign n4980 = n4978 | n4979 ;
  assign n4981 = n331 | n604 ;
  assign n4982 = n4980 | n4981 ;
  assign n4983 = n4977 | n4982 ;
  assign n4984 = n4901 | n4955 ;
  assign n4985 = n4901 & n4955 ;
  assign n4986 = ( n4903 & n4984 ) | ( n4903 & n4985 ) | ( n4984 & n4985 ) ;
  assign n4987 = ( n4902 & n4984 ) | ( n4902 & n4985 ) | ( n4984 & n4985 ) ;
  assign n4988 = ( n4815 & n4986 ) | ( n4815 & n4987 ) | ( n4986 & n4987 ) ;
  assign n4989 = n566 & ~n977 ;
  assign n4990 = ~n3119 & n4989 ;
  assign n4991 = n977 & ~n4906 ;
  assign n4992 = n4990 | n4991 ;
  assign n4993 = n566 & n3147 ;
  assign n4994 = ~n4992 & n4993 ;
  assign n4995 = n4992 & ~n4993 ;
  assign n4996 = n4994 | n4995 ;
  assign n4997 = n2501 & ~n3729 ;
  assign n4998 = n2512 & n3162 ;
  assign n4999 = n2499 & ~n3590 ;
  assign n5000 = n4998 | n4999 ;
  assign n5001 = n4997 | n5000 ;
  assign n5002 = n2491 | n5001 ;
  assign n5003 = ( n3742 & n5001 ) | ( n3742 & n5002 ) | ( n5001 & n5002 ) ;
  assign n5004 = ~n566 & n5003 ;
  assign n5005 = n566 & ~n5003 ;
  assign n5006 = ( n4996 & n5004 ) | ( n4996 & n5005 ) | ( n5004 & n5005 ) ;
  assign n5007 = n5004 | n5005 ;
  assign n5008 = n4996 | n5007 ;
  assign n5009 = ~n5006 & n5008 ;
  assign n5010 = n4914 & n5009 ;
  assign n5011 = n4914 & ~n5010 ;
  assign n5012 = ( n5009 & ~n5010 ) | ( n5009 & n5011 ) | ( ~n5010 & n5011 ) ;
  assign n5013 = n4926 & n4934 ;
  assign n5014 = ( n4937 & ~n4938 ) | ( n4937 & n5013 ) | ( ~n4938 & n5013 ) ;
  assign n5015 = ~n5012 & n5014 ;
  assign n5016 = n5012 & ~n5014 ;
  assign n5017 = n5015 | n5016 ;
  assign n5018 = ~n4941 & n4944 ;
  assign n5019 = n5017 | n5018 ;
  assign n5020 = n4942 | n5017 ;
  assign n5021 = ( ~n4905 & n5019 ) | ( ~n4905 & n5020 ) | ( n5019 & n5020 ) ;
  assign n5022 = ~n4941 & n4946 ;
  assign n5023 = n5017 | n5022 ;
  assign n5024 = ( ~n4830 & n5019 ) | ( ~n4830 & n5023 ) | ( n5019 & n5023 ) ;
  assign n5025 = ( ~n4572 & n5021 ) | ( ~n4572 & n5024 ) | ( n5021 & n5024 ) ;
  assign n5026 = n5017 & n5018 ;
  assign n5027 = n4942 & n5017 ;
  assign n5028 = ( ~n4905 & n5026 ) | ( ~n4905 & n5027 ) | ( n5026 & n5027 ) ;
  assign n5029 = n5017 & n5022 ;
  assign n5030 = ( ~n4830 & n5026 ) | ( ~n4830 & n5029 ) | ( n5026 & n5029 ) ;
  assign n5031 = ( ~n4572 & n5028 ) | ( ~n4572 & n5030 ) | ( n5028 & n5030 ) ;
  assign n5032 = ( n5028 & n5030 ) | ( n5028 & n5031 ) | ( n5030 & n5031 ) ;
  assign n5033 = n5025 & ~n5032 ;
  assign n5034 = ( n4983 & n4988 ) | ( n4983 & ~n5033 ) | ( n4988 & ~n5033 ) ;
  assign n5035 = ( ~n4988 & n5033 ) | ( ~n4988 & n5034 ) | ( n5033 & n5034 ) ;
  assign n5036 = ( ~n4983 & n5034 ) | ( ~n4983 & n5035 ) | ( n5034 & n5035 ) ;
  assign n5037 = n4959 & n5036 ;
  assign n5038 = n4819 & n5037 ;
  assign n5039 = n4960 | n5036 ;
  assign n5040 = ~n5038 & n5039 ;
  assign n5041 = n4884 | n4962 ;
  assign n5042 = n4827 | n5041 ;
  assign n5043 = n3859 & n5042 ;
  assign n5044 = ~n5040 & n5043 ;
  assign n5045 = n5040 & ~n5043 ;
  assign n5046 = n5044 | n5045 ;
  assign n5047 = n4983 | n5033 ;
  assign n5048 = n2179 | n2232 ;
  assign n5049 = n312 | n5048 ;
  assign n5050 = n925 | n5049 ;
  assign n5051 = n474 | n5050 ;
  assign n5052 = n170 | n5051 ;
  assign n5053 = n265 | n273 ;
  assign n5054 = n211 | n293 ;
  assign n5055 = n5053 | n5054 ;
  assign n5056 = n348 | n513 ;
  assign n5057 = n363 | n5056 ;
  assign n5058 = ( ~n547 & n3141 ) | ( ~n547 & n5057 ) | ( n3141 & n5057 ) ;
  assign n5059 = n547 | n5058 ;
  assign n5060 = n5055 | n5059 ;
  assign n5061 = n5052 | n5060 ;
  assign n5062 = ~n5015 & n5024 ;
  assign n5063 = ~n5015 & n5021 ;
  assign n5064 = ( ~n4571 & n5062 ) | ( ~n4571 & n5063 ) | ( n5062 & n5063 ) ;
  assign n5065 = ( ~n4570 & n5062 ) | ( ~n4570 & n5063 ) | ( n5062 & n5063 ) ;
  assign n5066 = ( ~n4207 & n5064 ) | ( ~n4207 & n5065 ) | ( n5064 & n5065 ) ;
  assign n5067 = ( ~n4996 & n5008 ) | ( ~n4996 & n5011 ) | ( n5008 & n5011 ) ;
  assign n5068 = n4990 | n4994 ;
  assign n5069 = n2512 & ~n3590 ;
  assign n5070 = n2499 & ~n3729 ;
  assign n5071 = n5069 | n5070 ;
  assign n5072 = ( n2491 & n3875 ) | ( n2491 & n5071 ) | ( n3875 & n5071 ) ;
  assign n5073 = ( n566 & ~n5071 ) | ( n566 & n5072 ) | ( ~n5071 & n5072 ) ;
  assign n5074 = ~n5072 & n5073 ;
  assign n5075 = n5071 | n5073 ;
  assign n5076 = ( ~n566 & n5074 ) | ( ~n566 & n5075 ) | ( n5074 & n5075 ) ;
  assign n5077 = ( ~n3162 & n5068 ) | ( ~n3162 & n5076 ) | ( n5068 & n5076 ) ;
  assign n5078 = n566 & ~n5068 ;
  assign n5079 = ( ~n3162 & n5076 ) | ( ~n3162 & n5078 ) | ( n5076 & n5078 ) ;
  assign n5080 = ( ~n5068 & n5076 ) | ( ~n5068 & n5078 ) | ( n5076 & n5078 ) ;
  assign n5081 = ( n5077 & ~n5079 ) | ( n5077 & n5080 ) | ( ~n5079 & n5080 ) ;
  assign n5082 = n5067 & ~n5081 ;
  assign n5083 = ~n5067 & n5081 ;
  assign n5084 = n5082 | n5083 ;
  assign n5085 = n5066 & n5084 ;
  assign n5086 = n5084 & ~n5085 ;
  assign n5087 = ( n5066 & ~n5085 ) | ( n5066 & n5086 ) | ( ~n5085 & n5086 ) ;
  assign n5088 = n5061 | n5087 ;
  assign n5089 = n5061 & n5087 ;
  assign n5090 = n5088 & ~n5089 ;
  assign n5091 = n5047 & n5090 ;
  assign n5092 = n4983 & n5033 ;
  assign n5093 = n5090 & n5092 ;
  assign n5094 = ( n4987 & n5091 ) | ( n4987 & n5093 ) | ( n5091 & n5093 ) ;
  assign n5095 = ( n4986 & n5091 ) | ( n4986 & n5093 ) | ( n5091 & n5093 ) ;
  assign n5096 = ( n4815 & n5094 ) | ( n4815 & n5095 ) | ( n5094 & n5095 ) ;
  assign n5097 = n5047 | n5090 ;
  assign n5098 = n5090 | n5092 ;
  assign n5099 = ( n4987 & n5097 ) | ( n4987 & n5098 ) | ( n5097 & n5098 ) ;
  assign n5100 = ( n4986 & n5097 ) | ( n4986 & n5098 ) | ( n5097 & n5098 ) ;
  assign n5101 = ( n4815 & n5099 ) | ( n4815 & n5100 ) | ( n5099 & n5100 ) ;
  assign n5102 = ~n5096 & n5101 ;
  assign n5103 = n5038 | n5102 ;
  assign n5104 = n5038 & n5102 ;
  assign n5105 = n5103 & ~n5104 ;
  assign n5106 = n5040 | n5042 ;
  assign n5107 = n3859 & n5106 ;
  assign n5108 = ~n5105 & n5107 ;
  assign n5109 = n5105 & ~n5107 ;
  assign n5110 = n5108 | n5109 ;
  assign n5111 = n566 & n3162 ;
  assign n5112 = ( n5068 & n5076 ) | ( n5068 & ~n5111 ) | ( n5076 & ~n5111 ) ;
  assign n5113 = n2512 & ~n3729 ;
  assign n5114 = n2491 & ~n3729 ;
  assign n5115 = n5113 | n5114 ;
  assign n5116 = ( ~n3590 & n5113 ) | ( ~n3590 & n5115 ) | ( n5113 & n5115 ) ;
  assign n5117 = ( n3604 & n5115 ) | ( n3604 & n5116 ) | ( n5115 & n5116 ) ;
  assign n5118 = ~n566 & n5117 ;
  assign n5119 = n566 & ~n3598 ;
  assign n5120 = ( n5117 & ~n5118 ) | ( n5117 & n5119 ) | ( ~n5118 & n5119 ) ;
  assign n5121 = ( n566 & n5118 ) | ( n566 & ~n5120 ) | ( n5118 & ~n5120 ) ;
  assign n5122 = ( ~n3598 & n5117 ) | ( ~n3598 & n5121 ) | ( n5117 & n5121 ) ;
  assign n5123 = ( n566 & n5121 ) | ( n566 & n5122 ) | ( n5121 & n5122 ) ;
  assign n5124 = ~n5112 & n5123 ;
  assign n5125 = n5112 & ~n5123 ;
  assign n5126 = n5124 | n5125 ;
  assign n5127 = n5082 & ~n5126 ;
  assign n5128 = ( n5084 & n5126 ) | ( n5084 & ~n5127 ) | ( n5126 & ~n5127 ) ;
  assign n5129 = ( n5066 & ~n5127 ) | ( n5066 & n5128 ) | ( ~n5127 & n5128 ) ;
  assign n5130 = ~n5082 & n5126 ;
  assign n5131 = ( n5066 & n5086 ) | ( n5066 & n5130 ) | ( n5086 & n5130 ) ;
  assign n5132 = n5129 & ~n5131 ;
  assign n5133 = n132 | n4890 ;
  assign n5134 = n235 | n250 ;
  assign n5135 = n894 | n5134 ;
  assign n5136 = n778 | n5135 ;
  assign n5137 = n5133 | n5136 ;
  assign n5138 = n2186 | n5137 ;
  assign n5139 = n380 | n1044 ;
  assign n5140 = n1033 | n5139 ;
  assign n5141 = n5138 | n5140 ;
  assign n5142 = n218 | n293 ;
  assign n5143 = n363 | n520 ;
  assign n5144 = n224 | n5143 ;
  assign n5145 = n518 | n5144 ;
  assign n5146 = n128 | n152 ;
  assign n5147 = n5145 | n5146 ;
  assign n5148 = n5142 | n5147 ;
  assign n5149 = n5141 | n5148 ;
  assign n5150 = n5132 & n5149 ;
  assign n5151 = n5132 | n5149 ;
  assign n5152 = ~n5150 & n5151 ;
  assign n5153 = n5089 | n5093 ;
  assign n5154 = n5089 | n5091 ;
  assign n5155 = ( n4988 & n5153 ) | ( n4988 & n5154 ) | ( n5153 & n5154 ) ;
  assign n5156 = n5152 | n5155 ;
  assign n5157 = n5152 & n5155 ;
  assign n5158 = n5156 & ~n5157 ;
  assign n5159 = n5102 & n5158 ;
  assign n5160 = n5038 & n5159 ;
  assign n5161 = n5104 | n5158 ;
  assign n5162 = ~n5160 & n5161 ;
  assign n5163 = ( n3859 & n5105 ) | ( n3859 & n5107 ) | ( n5105 & n5107 ) ;
  assign n5164 = ~n5162 & n5163 ;
  assign n5165 = n5162 & ~n5163 ;
  assign n5166 = n5164 | n5165 ;
  assign n5167 = n5105 | n5162 ;
  assign n5168 = n5106 | n5167 ;
  assign n5169 = n3859 & n5168 ;
  assign n5170 = n305 | n4969 ;
  assign n5171 = n796 | n2112 ;
  assign n5172 = n2022 | n5171 ;
  assign n5173 = n5170 | n5172 ;
  assign n5174 = n129 | n3462 ;
  assign n5175 = n5173 | n5174 ;
  assign n5176 = n887 | n5175 ;
  assign n5177 = n155 | n3510 ;
  assign n5178 = n197 | n321 ;
  assign n5179 = n5177 | n5178 ;
  assign n5180 = n5176 | n5179 ;
  assign n5181 = ~n5111 & n5119 ;
  assign n5182 = n5121 | n5181 ;
  assign n5183 = n5125 & ~n5182 ;
  assign n5184 = ( n5128 & n5182 ) | ( n5128 & ~n5183 ) | ( n5182 & ~n5183 ) ;
  assign n5185 = ( n5127 & ~n5182 ) | ( n5127 & n5183 ) | ( ~n5182 & n5183 ) ;
  assign n5186 = ( n5064 & n5184 ) | ( n5064 & ~n5185 ) | ( n5184 & ~n5185 ) ;
  assign n5187 = ( n5065 & n5184 ) | ( n5065 & ~n5185 ) | ( n5184 & ~n5185 ) ;
  assign n5188 = ( ~n4207 & n5186 ) | ( ~n4207 & n5187 ) | ( n5186 & n5187 ) ;
  assign n5189 = ~n5125 & n5182 ;
  assign n5190 = n5129 & n5189 ;
  assign n5191 = n5188 & ~n5190 ;
  assign n5192 = ( n3729 & n5111 ) | ( n3729 & n5191 ) | ( n5111 & n5191 ) ;
  assign n5193 = n566 & n5192 ;
  assign n5194 = ( n3729 & n5111 ) | ( n3729 & ~n5192 ) | ( n5111 & ~n5192 ) ;
  assign n5195 = n566 & n5194 ;
  assign n5196 = ( n5191 & ~n5193 ) | ( n5191 & n5195 ) | ( ~n5193 & n5195 ) ;
  assign n5197 = n5180 & n5196 ;
  assign n5198 = n5180 | n5196 ;
  assign n5199 = ~n5197 & n5198 ;
  assign n5200 = n5150 & n5199 ;
  assign n5201 = ( n5157 & n5199 ) | ( n5157 & n5200 ) | ( n5199 & n5200 ) ;
  assign n5202 = ( ~n5150 & n5157 ) | ( ~n5150 & n5199 ) | ( n5157 & n5199 ) ;
  assign n5203 = n5150 | n5202 ;
  assign n5204 = ~n5201 & n5203 ;
  assign n5205 = n5160 & n5204 ;
  assign n5206 = n5160 & ~n5205 ;
  assign n5207 = ( n5204 & ~n5205 ) | ( n5204 & n5206 ) | ( ~n5205 & n5206 ) ;
  assign n5208 = n5169 & ~n5207 ;
  assign n5209 = ~n5169 & n5207 ;
  assign n5210 = n5208 | n5209 ;
  assign n5211 = n548 | n694 ;
  assign n5212 = n592 | n870 ;
  assign n5213 = n5211 | n5212 ;
  assign n5214 = n1948 | n5213 ;
  assign n5215 = n2348 | n5214 ;
  assign n5216 = n737 | n5215 ;
  assign n5217 = n205 | n386 ;
  assign n5218 = n543 | n5217 ;
  assign n5219 = n247 | n633 ;
  assign n5220 = n5218 | n5219 ;
  assign n5221 = n5216 | n5220 ;
  assign n5222 = n5197 & n5221 ;
  assign n5223 = ( n5200 & n5221 ) | ( n5200 & n5222 ) | ( n5221 & n5222 ) ;
  assign n5224 = ( n5199 & n5221 ) | ( n5199 & n5222 ) | ( n5221 & n5222 ) ;
  assign n5225 = ( n5157 & n5223 ) | ( n5157 & n5224 ) | ( n5223 & n5224 ) ;
  assign n5226 = n5197 | n5221 ;
  assign n5227 = n5201 | n5226 ;
  assign n5228 = ~n5225 & n5227 ;
  assign n5229 = n5205 & ~n5228 ;
  assign n5230 = n5228 | n5229 ;
  assign n5231 = ( ~n5205 & n5229 ) | ( ~n5205 & n5230 ) | ( n5229 & n5230 ) ;
  assign n5232 = ( n3859 & n5169 ) | ( n3859 & n5207 ) | ( n5169 & n5207 ) ;
  assign n5233 = n5231 & n5232 ;
  assign n5234 = n5231 | n5232 ;
  assign n5235 = ~n5233 & n5234 ;
  assign n5236 = n5207 | n5231 ;
  assign n5237 = ( n3859 & n5169 ) | ( n3859 & n5236 ) | ( n5169 & n5236 ) ;
  assign n5238 = n242 | n775 ;
  assign n5239 = n1007 | n5238 ;
  assign n5240 = n704 | n5239 ;
  assign n5241 = n151 | n512 ;
  assign n5242 = n5240 | n5241 ;
  assign n5243 = n513 | n3544 ;
  assign n5244 = n205 | n397 ;
  assign n5245 = n97 | n187 ;
  assign n5246 = n5244 | n5245 ;
  assign n5247 = n5243 | n5246 ;
  assign n5248 = n5242 | n5247 ;
  assign n5249 = n5204 & n5228 ;
  assign n5250 = n5160 & n5249 ;
  assign n5251 = ( n5225 & ~n5248 ) | ( n5225 & n5250 ) | ( ~n5248 & n5250 ) ;
  assign n5252 = ( n5225 & n5248 ) | ( n5225 & ~n5250 ) | ( n5248 & ~n5250 ) ;
  assign n5253 = ( ~n5225 & n5251 ) | ( ~n5225 & n5252 ) | ( n5251 & n5252 ) ;
  assign n5254 = n5237 & ~n5253 ;
  assign n5255 = ~n5237 & n5253 ;
  assign n5256 = n5254 | n5255 ;
  assign n5257 = n459 | n5134 ;
  assign n5258 = n4302 | n5257 ;
  assign n5259 = n1972 | n5258 ;
  assign n5260 = n861 | n5259 ;
  assign n5261 = n5140 | n5260 ;
  assign n5262 = n207 | n212 ;
  assign n5263 = n155 | n181 ;
  assign n5264 = n5262 | n5263 ;
  assign n5265 = n164 | n290 ;
  assign n5266 = n227 | n5265 ;
  assign n5267 = n5264 | n5266 ;
  assign n5268 = n5261 | n5267 ;
  assign n5269 = n5248 | n5268 ;
  assign n5270 = ( n5224 & n5268 ) | ( n5224 & n5269 ) | ( n5268 & n5269 ) ;
  assign n5271 = ( n5223 & n5268 ) | ( n5223 & n5269 ) | ( n5268 & n5269 ) ;
  assign n5272 = ( n5157 & n5270 ) | ( n5157 & n5271 ) | ( n5270 & n5271 ) ;
  assign n5273 = n5248 & n5268 ;
  assign n5274 = n5225 & n5273 ;
  assign n5275 = n5272 & ~n5274 ;
  assign n5276 = n5225 | n5248 ;
  assign n5277 = n5250 & ~n5276 ;
  assign n5278 = ( n5250 & n5275 ) | ( n5250 & n5277 ) | ( n5275 & n5277 ) ;
  assign n5279 = ( n5275 & n5277 ) | ( n5275 & ~n5278 ) | ( n5277 & ~n5278 ) ;
  assign n5280 = ( n5250 & ~n5278 ) | ( n5250 & n5279 ) | ( ~n5278 & n5279 ) ;
  assign n5281 = ( n3859 & n5237 ) | ( n3859 & n5253 ) | ( n5237 & n5253 ) ;
  assign n5282 = ~n5280 & n5281 ;
  assign n5283 = n5280 & ~n5281 ;
  assign n5284 = n5282 | n5283 ;
  assign n5285 = n5168 | n5236 ;
  assign n5286 = ( n5253 & n5280 ) | ( n5253 & ~n5285 ) | ( n5280 & ~n5285 ) ;
  assign n5287 = n5285 | n5286 ;
  assign n5288 = n3859 & n5287 ;
  assign n5289 = n5249 & n5276 ;
  assign n5290 = n272 | n360 ;
  assign n5291 = n738 | n5290 ;
  assign n5292 = n3129 | n5291 ;
  assign n5293 = n916 | n5292 ;
  assign n5294 = n4559 | n5293 ;
  assign n5295 = n397 | n405 ;
  assign n5296 = n1931 | n5295 ;
  assign n5297 = n223 | n399 ;
  assign n5298 = n280 | n5297 ;
  assign n5299 = n5296 | n5298 ;
  assign n5300 = n101 | n232 ;
  assign n5301 = n5299 | n5300 ;
  assign n5302 = n5294 | n5301 ;
  assign n5303 = n5273 | n5302 ;
  assign n5304 = ( n5224 & n5302 ) | ( n5224 & n5303 ) | ( n5302 & n5303 ) ;
  assign n5305 = ( n5223 & n5302 ) | ( n5223 & n5303 ) | ( n5302 & n5303 ) ;
  assign n5306 = ( n5157 & n5304 ) | ( n5157 & n5305 ) | ( n5304 & n5305 ) ;
  assign n5307 = ( n5275 & ~n5289 ) | ( n5275 & n5306 ) | ( ~n5289 & n5306 ) ;
  assign n5308 = n5289 & n5307 ;
  assign n5309 = n5160 & n5308 ;
  assign n5310 = n5273 & n5302 ;
  assign n5311 = n5225 & n5310 ;
  assign n5312 = n5306 & ~n5311 ;
  assign n5313 = ( ~n5277 & n5278 ) | ( ~n5277 & n5312 ) | ( n5278 & n5312 ) ;
  assign n5314 = ~n5309 & n5313 ;
  assign n5315 = n5288 & ~n5314 ;
  assign n5316 = ~n5288 & n5314 ;
  assign n5317 = n5315 | n5316 ;
  assign n5318 = n336 | n3152 ;
  assign n5319 = n412 | n5318 ;
  assign n5320 = n335 | n5319 ;
  assign n5321 = n2079 | n5320 ;
  assign n5322 = n414 | n5321 ;
  assign n5323 = n5310 | n5322 ;
  assign n5324 = ( n5224 & n5322 ) | ( n5224 & n5323 ) | ( n5322 & n5323 ) ;
  assign n5325 = ( n5223 & n5322 ) | ( n5223 & n5323 ) | ( n5322 & n5323 ) ;
  assign n5326 = ( n5157 & n5324 ) | ( n5157 & n5325 ) | ( n5324 & n5325 ) ;
  assign n5327 = n5302 & n5322 ;
  assign n5328 = n5273 & n5327 ;
  assign n5329 = n5225 & n5328 ;
  assign n5330 = n5326 & ~n5329 ;
  assign n5331 = n5309 | n5330 ;
  assign n5332 = n5309 & n5330 ;
  assign n5333 = n5331 & ~n5332 ;
  assign n5334 = ( n3859 & n5288 ) | ( n3859 & n5314 ) | ( n5288 & n5314 ) ;
  assign n5335 = ~n5333 & n5334 ;
  assign n5336 = n5333 & ~n5334 ;
  assign n5337 = n5335 | n5336 ;
  assign n5338 = ( ~n304 & n313 ) | ( ~n304 & n414 ) | ( n313 & n414 ) ;
  assign n5339 = n304 | n5338 ;
  assign n5340 = n5328 | n5339 ;
  assign n5341 = ( n5224 & n5339 ) | ( n5224 & n5340 ) | ( n5339 & n5340 ) ;
  assign n5342 = ( n5223 & n5339 ) | ( n5223 & n5340 ) | ( n5339 & n5340 ) ;
  assign n5343 = ( n5157 & n5341 ) | ( n5157 & n5342 ) | ( n5341 & n5342 ) ;
  assign n5344 = n5328 & n5339 ;
  assign n5345 = n5225 & n5344 ;
  assign n5346 = n5343 & ~n5345 ;
  assign n5347 = n5332 | n5346 ;
  assign n5348 = ~n5343 & n5347 ;
  assign n5349 = ( ~n5332 & n5347 ) | ( ~n5332 & n5348 ) | ( n5347 & n5348 ) ;
  assign n5350 = ( n3859 & n5333 ) | ( n3859 & n5334 ) | ( n5333 & n5334 ) ;
  assign n5351 = ~n5349 & n5350 ;
  assign n5352 = n5349 & ~n5350 ;
  assign n5353 = n5351 | n5352 ;
  assign n5354 = ( n3859 & n5349 ) | ( n3859 & n5350 ) | ( n5349 & n5350 ) ;
  assign n5355 = ( ~n5332 & n5343 ) | ( ~n5332 & n5345 ) | ( n5343 & n5345 ) ;
  assign n5356 = n5332 & n5355 ;
  assign n5357 = ( n5332 & n5343 ) | ( n5332 & n5345 ) | ( n5343 & n5345 ) ;
  assign n5358 = ~n5356 & n5357 ;
  assign n5359 = n5354 | n5358 ;
  assign n5360 = x22 | n54 ;
  assign n5361 = ( n5358 & ~n5359 ) | ( n5358 & n5360 ) | ( ~n5359 & n5360 ) ;
  assign n5362 = ( n5354 & ~n5359 ) | ( n5354 & n5361 ) | ( ~n5359 & n5361 ) ;
  assign n5363 = n5314 | n5333 ;
  assign n5364 = n5349 | n5363 ;
  assign n5365 = n5287 | n5364 ;
  assign n5366 = n5357 & ~n5365 ;
  assign n5367 = ~n5356 & n5365 ;
  assign n5368 = n5366 | n5367 ;
  assign n5369 = n3859 & ~n5360 ;
  assign n5370 = ( n3859 & n5368 ) | ( n3859 & n5369 ) | ( n5368 & n5369 ) ;
  assign y0 = n3704 ;
  assign y1 = n3863 ;
  assign y2 = n3989 ;
  assign y3 = n4116 ;
  assign y4 = n4230 ;
  assign y5 = n4326 ;
  assign y6 = n4452 ;
  assign y7 = n4545 ;
  assign y8 = n4652 ;
  assign y9 = n4740 ;
  assign y10 = n4825 ;
  assign y11 = n4887 ;
  assign y12 = n4966 ;
  assign y13 = n5046 ;
  assign y14 = n5110 ;
  assign y15 = n5166 ;
  assign y16 = n5210 ;
  assign y17 = n5235 ;
  assign y18 = n5256 ;
  assign y19 = n5284 ;
  assign y20 = n5317 ;
  assign y21 = n5337 ;
  assign y22 = n5353 ;
  assign y23 = ~n5362 ;
  assign y24 = n5370 ;
endmodule
