//Written by the Majority Logic Package Fri Nov 14 23:12:53 2014
module top (
            b0, a0, cin, b1, a1, b10, b9, b8, b7, b6, b5, b4, b3, b2, a2, a3, a4, a5, a6, a7, a8, a9, a10, b11, a11, b12, a12, b13, a13, b14, a14, b15, a15, b16, a16, b17, a17, b18, a18, b19, a19, b20, a20, b21, a21, b22, a22, b23, a23, b24, a24, b25, a25, b26, a26, b27, a27, b28, a28, b29, a29, b30, a30, b31, a31, b32, a32, b33, a33, b34, a34, b35, a35, b36, a36, b37, a37, b38, a38, b39, a39, b40, a40, b41, a41, b42, a42, b43, a43, b44, a44, b45, a45, b46, a46, b47, a47, b48, a48, b49, a49, b50, a50, b51, a51, b52, a52, b53, a53, b54, a54, b55, a55, b56, a56, b57, a57, b58, a58, b59, a59, b60, a60, b61, a61, b62, a62, a63, b63, 
            s0, s1, s10, s11, s12, s13, s14, s15, s16, s17, s18, s19, s2, s20, s21, s22, s23, s24, s25, s26, s27, s28, s29, s3, s30, s31, s32, s33, s34, s35, s36, s37, s38, s39, s4, s40, s41, s42, s43, s44, s45, s46, s47, s48, s49, s5, s50, s51, s52, s53, s54, s55, s56, s57, s58, s59, s6, s60, s61, s62, s63, s64, s7, s8, s9);
input b0, a0, cin, b1, a1, b10, b9, b8, b7, b6, b5, b4, b3, b2, a2, a3, a4, a5, a6, a7, a8, a9, a10, b11, a11, b12, a12, b13, a13, b14, a14, b15, a15, b16, a16, b17, a17, b18, a18, b19, a19, b20, a20, b21, a21, b22, a22, b23, a23, b24, a24, b25, a25, b26, a26, b27, a27, b28, a28, b29, a29, b30, a30, b31, a31, b32, a32, b33, a33, b34, a34, b35, a35, b36, a36, b37, a37, b38, a38, b39, a39, b40, a40, b41, a41, b42, a42, b43, a43, b44, a44, b45, a45, b46, a46, b47, a47, b48, a48, b49, a49, b50, a50, b51, a51, b52, a52, b53, a53, b54, a54, b55, a55, b56, a56, b57, a57, b58, a58, b59, a59, b60, a60, b61, a61, b62, a62, a63, b63;
output s0, s1, s10, s11, s12, s13, s14, s15, s16, s17, s18, s19, s2, s20, s21, s22, s23, s24, s25, s26, s27, s28, s29, s3, s30, s31, s32, s33, s34, s35, s36, s37, s38, s39, s4, s40, s41, s42, s43, s44, s45, s46, s47, s48, s49, s5, s50, s51, s52, s53, s54, s55, s56, s57, s58, s59, s6, s60, s61, s62, s63, s64, s7, s8, s9;
wire one, w0, w1, w2, w3, w4, w5, w6, w7, w8, w9, w10, w11, w12, w13, w14, w15, w16, w17, w18, w19, w20, w21, w22, w23, w24, w25, w26, w27, w28, w29, w30, w31, w32, w33, w34, w35, w36, w37, w38, w39, w40, w41, w42, w43, w44, w45, w46, w47, w48, w49, w50, w51, w52, w53, w54, w55, w56, w57, w58, w59, w60, w61, w62, w63, w64, w65, w66, w67, w68, w69, w70, w71, w72, w73, w74, w75, w76, w77, w78, w79, w80, w81, w82, w83, w84, w85, w86, w87, w88, w89, w90, w91, w92, w93, w94, w95, w96, w97, w98, w99, w100, w101, w102, w103, w104, w105, w106, w107, w108, w109, w110, w111, w112, w113, w114, w115, w116, w117, w118, w119, w120, w121, w122, w123, w124, w125, w126, w127, w128, w129, w130, w131, w132, w133, w134, w135, w136, w137, w138, w139, w140, w141, w142, w143, w144, w145, w146, w147, w148, w149, w150, w151, w152, w153, w154, w155, w156, w157, w158, w159, w160, w161, w162, w163, w164, w165, w166, w167, w168, w169, w170, w171, w172, w173, w174, w175, w176, w177, w178, w179, w180, w181, w182, w183, w184, w185, w186, w187, w188, w189, w190, w191, w192, w193, w194, w195, w196, w197, w198, w199, w200, w201, w202, w203, w204, w205, w206, w207, w208, w209, w210, w211, w212, w213, w214, w215, w216, w217, w218, w219, w220, w221, w222, w223, w224, w225, w226, w227, w228, w229, w230, w231, w232, w233, w234, w235, w236, w237, w238, w239, w240, w241, w242, w243, w244, w245, w246, w247, w248, w249, w250, w251, w252, w253, w254, w255, w256, w257, w258, w259, w260, w261, w262, w263, w264, w265, w266, w267, w268, w269, w270, w271, w272, w273, w274, w275, w276, w277, w278, w279, w280, w281, w282, w283, w284, w285, w286, w287, w288, w289, w290, w291, w292, w293, w294, w295, w296, w297, w298, w299, w300, w301, w302, w303, w304, w305, w306, w307, w308, w309, w310, w311, w312, w313, w314, w315, w316, w317, w318, w319, w320, w321, w322, w323, w324, w325, w326, w327, w328, w329, w330, w331, w332, w333, w334, w335, w336, w337, w338, w339, w340, w341, w342, w343, w344, w345, w346, w347, w348, w349, w350, w351, w352, w353, w354, w355, w356, w357, w358, w359, w360, w361, w362, w363, w364, w365, w366, w367, w368, w369, w370, w371, w372, w373, w374, w375, w376, w377, w378, w379, w380, w381, w382, w383, w384, w385, w386, w387, w388, w389, w390, w391, w392, w393, w394, w395, w396, w397, w398, w399, w400, w401, w402, w403, w404, w405, w406, w407, w408, w409, w410, w411, w412, w413, w414, w415, w416, w417, w418, w419, w420, w421, w422, w423, w424, w425, w426, w427, w428, w429, w430, w431, w432, w433, w434, w435, w436, w437, w438, w439, w440, w441, w442, w443, w444, w445, w446, w447, w448, w449, w450, w451, w452, w453, w454, w455, w456, w457, w458, w459, w460, w461, w462, w463, w464, w465, w466, w467, w468, w469, w470, w471, w472, w473, w474, w475, w476, w477, w478, w479, w480, w481, w482, w483, w484, w485, w486, w487, w488, w489, w490, w491, w492, w493, w494, w495, w496, w497, w498, w499, w500, w501, w502, w503, w504, w505, w506, w507, w508, w509, w510, w511, w512, w513, w514, w515, w516, w517, w518, w519, w520, w521, w522, w523, w524, w525, w526, w527, w528, w529, w530, w531, w532, w533, w534, w535, w536, w537, w538, w539, w540, w541, w542, w543, w544, w545, w546, w547, w548, w549, w550, w551, w552, w553, w554, w555, w556, w557, w558, w559, w560, w561, w562, w563, w564, w565, w566, w567, w568, w569, w570, w571, w572, w573, w574, w575, w576, w577, w578, w579, w580, w581, w582, w583, w584, w585, w586, w587, w588, w589, w590, w591, w592, w593, w594, w595, w596, w597, w598, w599, w600, w601, w602, w603, w604, w605, w606, w607, w608, w609, w610, w611, w612, w613, w614, w615, w616, w617, w618, w619, w620, w621, w622, w623, w624, w625, w626, w627, w628, w629, w630, w631, w632, w633, w634, w635, w636, w637, w638, w639, w640, w641, w642, w643, w644, w645, w646, w647, w648, w649, w650, w651, w652, w653, w654, w655, w656, w657, w658, w659, w660, w661, w662, w663, w664, w665, w666, w667, w668, w669, w670, w671, w672, w673, w674, w675, w676, w677, w678, w679, w680, w681, w682, w683, w684, w685, w686, w687, w688, w689, w690, w691, w692, w693, w694, w695, w696, w697, w698, w699, w700, w701, w702, w703, w704, w705, w706, w707, w708, w709, w710, w711, w712, w713, w714, w715, w716, w717, w718, w719, w720, w721, w722, w723, w724, w725, w726, w727, w728, w729, w730, w731, w732, w733, w734, w735, w736, w737, w738, w739, w740, w741, w742, w743, w744, w745, w746, w747, w748, w749, w750, w751, w752, w753, w754, w755, w756, w757, w758, w759, w760, w761, w762, w763, w764, w765, w766, w767, w768, w769, w770, w771, w772, w773, w774, w775, w776, w777, w778, w779, w780, w781, w782, w783, w784, w785, w786, w787, w788, w789, w790, w791, w792, w793, w794, w795, w796, w797, w798, w799, w800, w801, w802, w803, w804, w805, w806, w807, w808, w809, w810, w811, w812, w813, w814, w815, w816, w817, w818, w819, w820, w821, w822, w823, w824, w825, w826, w827, w828, w829, w830, w831, w832, w833, w834, w835, w836, w837, w838, w839, w840, w841, w842, w843, w844, w845, w846, w847, w848, w849, w850, w851, w852, w853, w854, w855, w856, w857, w858, w859, w860, w861, w862, w863, w864, w865, w866, w867, w868, w869, w870, w871, w872, w873, w874, w875, w876, w877, w878, w879, w880, w881, w882, w883, w884, w885, w886, w887, w888, w889, w890, w891, w892, w893, w894, w895, w896, w897, w898, w899, w900, w901, w902, w903, w904, w905, w906, w907, w908, w909, w910, w911, w912, w913, w914, w915, w916, w917, w918, w919, w920, w921, w922, w923, w924, w925, w926, w927, w928, w929, w930, w931, w932, w933, w934, w935, w936, w937, w938, w939, w940, w941, w942, w943, w944, w945, w946, w947, w948, w949, w950, w951, w952, w953, w954, w955, w956, w957, w958, w959, w960, w961, w962, w963, w964, w965, w966, w967, w968, w969, w970, w971, w972, w973, w974, w975, w976, w977, w978, w979, w980, w981, w982, w983, w984, w985, w986, w987, w988, w989, w990, w991, w992, w993, w994, w995, w996, w997, w998, w999, w1000, w1001, w1002, w1003, w1004, w1005, w1006, w1007, w1008, w1009, w1010, w1011, w1012, w1013, w1014, w1015, w1016, w1017, w1018, w1019, w1020, w1021, w1022, w1023, w1024, w1025, w1026, w1027, w1028, w1029, w1030, w1031, w1032, w1033, w1034, w1035, w1036, w1037, w1038, w1039, w1040, w1041, w1042, w1043, w1044, w1045, w1046, w1047, w1048, w1049, w1050, w1051, w1052, w1053, w1054, w1055, w1056, w1057, w1058, w1059, w1060, w1061, w1062, w1063, w1064, w1065, w1066, w1067, w1068, w1069, w1070, w1071, w1072, w1073, w1074, w1075, w1076, w1077, w1078, w1079, w1080, w1081, w1082, w1083, w1084, w1085, w1086, w1087, w1088, w1089, w1090, w1091, w1092, w1093, w1094, w1095, w1096, w1097, w1098, w1099, w1100, w1101, w1102, w1103, w1104, w1105, w1106, w1107, w1108, w1109, w1110, w1111, w1112, w1113, w1114, w1115, w1116, w1117, w1118, w1119, w1120, w1121, w1122, w1123, w1124, w1125, w1126, w1127, w1128, w1129, w1130, w1131, w1132, w1133, w1134, w1135, w1136, w1137, w1138, w1139, w1140, w1141, w1142, w1143, w1144, w1145, w1146, w1147, w1148, w1149, w1150, w1151, w1152, w1153, w1154, w1155, w1156, w1157, w1158;
assign w0 = b20 & a20;
assign w1 = ~b28 & ~a28;
assign w2 = w1123 & w821;
assign w3 = (w958 & w295) | (w958 & w91) | (w295 & w91);
assign w4 = ~w924 & ~w408;
assign w5 = (w77 & w99) | (w77 & w1045) | (w99 & w1045);
assign w6 = (w262 & w125) | (w262 & ~w1101) | (w125 & ~w1101);
assign w7 = w1138 & w610;
assign w8 = ~w1131 & ~w848;
assign w9 = (w294 & w846) | (w294 & w264) | (w846 & w264);
assign w10 = w709 & w329;
assign w11 = ~w165 & ~w327;
assign w12 = ~w953 & ~w495;
assign w13 = ~w592 & w434;
assign w14 = ~w123 & w2;
assign w15 = ~w551 & ~w248;
assign w16 = (w381 & w768) | (w381 & w956) | (w768 & w956);
assign w17 = ~w448 & w1134;
assign w18 = ~w115 & w1120;
assign w19 = ~w861 & w298;
assign w20 = w532 & w90;
assign w21 = ~w690 & ~w640;
assign w22 = (w958 & w295) | (w958 & w898) | (w295 & w898);
assign w23 = (w80 & w926) | (w80 & w1053) | (w926 & w1053);
assign w24 = b7 & a7;
assign w25 = w194 & w672;
assign w26 = w191 & ~w1060;
assign w27 = ~w317 & ~w445;
assign w28 = (~w898 & w110) | (~w898 & w86) | (w110 & w86);
assign w29 = (w829 & w75) | (w829 & w527) | (w75 & w527);
assign w30 = b0 & a0;
assign w31 = ~w1131 & ~w303;
assign w32 = w202 & w677;
assign w33 = ~w1100 & ~w634;
assign w34 = w346 & w77;
assign w35 = b2 & a2;
assign w36 = ~w1155 & w637;
assign w37 = (~w742 & w626) | (~w742 & w245) | (w626 & w245);
assign w38 = (w387 & w822) | (w387 & w365) | (w822 & w365);
assign w39 = ~w84 & ~w403;
assign w40 = w349 & w269;
assign w41 = (w692 & w1096) | (w692 & w584) | (w1096 & w584);
assign w42 = ~w843 & ~w33;
assign w43 = w55 & ~w1019;
assign w44 = (w28 & w177) | (w28 & ~w1101) | (w177 & ~w1101);
assign w45 = ~w228 & ~w1119;
assign w46 = (~w518 & w660) | (~w518 & w200) | (w660 & w200);
assign w47 = ~w492 & ~w76;
assign w48 = w700 & w684;
assign w49 = (w170 & w884) | (w170 & w77) | (w884 & w77);
assign w50 = ~w35 & ~w509;
assign w51 = w361 & ~w627;
assign w52 = (w89 & w337) | (w89 & w856) | (w337 & w856);
assign w53 = ~w930 & ~w324;
assign w54 = w1100 & w653;
assign w55 = ~w728 & w793;
assign w56 = (~w733 & w1015) | (~w733 & w1149) | (w1015 & w1149);
assign w57 = (~w531 & w773) | (~w531 & w840) | (w773 & w840);
assign w58 = ~w423 & ~w994;
assign w59 = (~w263 & w526) | (~w263 & w687) | (w526 & w687);
assign w60 = w1062 & w795;
assign w61 = w346 & ~w183;
assign w62 = ~w778 & ~w1156;
assign w63 = (w916 & ~w913) | (w916 & w1098) | (~w913 & w1098);
assign w64 = (w88 & w1075) | (w88 & ~w83) | (w1075 & ~w83);
assign w65 = w661 & w593;
assign w66 = ~w287 & ~w783;
assign w67 = w689 & w284;
assign w68 = (~w658 & w254) | (~w658 & w237) | (w254 & w237);
assign w69 = w1109 & ~w673;
assign w70 = w154 & w706;
assign w71 = (~w531 & w1041) | (~w531 & w435) | (w1041 & w435);
assign w72 = (w718 & w1000) | (w718 & w59) | (w1000 & w59);
assign w73 = (w552 & w742) | (w552 & w833) | (w742 & w833);
assign w74 = b49 & a49;
assign w75 = (w593 & w65) | (w593 & ~w461) | (w65 & ~w461);
assign w76 = (~w658 & w268) | (~w658 & w438) | (w268 & w438);
assign w77 = ~w671 & w395;
assign w78 = w1024 & ~w337;
assign w79 = w223 & w559;
assign w80 = ~w656 & ~w636;
assign w81 = ~w384 & w338;
assign w82 = (w854 & ~w1012) | (w854 & ~w83) | (~w1012 & ~w83);
assign w83 = w672 & w236;
assign w84 = (~w1034 & w600) | (~w1034 & w937) | (w600 & w937);
assign w85 = w991 & w550;
assign w86 = (~w115 & w291) | (~w115 & w110) | (w291 & w110);
assign w87 = (w658 & w770) | (w658 & w145) | (w770 & w145);
assign w88 = w222 & ~w726;
assign w89 = ~w528 & w523;
assign w90 = ~w557 & ~w35;
assign w91 = (w904 & ~w17) | (w904 & w1142) | (~w17 & w1142);
assign w92 = (~w898 & w852) | (~w898 & w1110) | (w852 & w1110);
assign w93 = ~w1109 & w683;
assign w94 = (~w1101 & w1051) | (~w1101 & w1157) | (w1051 & w1157);
assign w95 = ~w138 & w717;
assign w96 = ~w286 & w979;
assign w97 = ~w753 & ~w959;
assign w98 = w202 & w361;
assign w99 = (w388 & w1088) | (w388 & w613) | (w1088 & w613);
assign w100 = (w1008 & w570) | (w1008 & w810) | (w570 & w810);
assign w101 = (w529 & w149) | (w529 & w278) | (w149 & w278);
assign w102 = (w533 & w301) | (w533 & ~w1101) | (w301 & ~w1101);
assign w103 = (w658 & w393) | (w658 & w246) | (w393 & w246);
assign w104 = ~b10 & ~a10;
assign w105 = ~b24 & ~a24;
assign w106 = ~w104 & ~w279;
assign w107 = ~w1109 & ~w431;
assign w108 = (w718 & w1000) | (w718 & w857) | (w1000 & w857);
assign w109 = (~w531 & w204) | (~w531 & w409) | (w204 & w409);
assign w110 = ~w115 & ~w7;
assign w111 = ~w1018 & ~w0;
assign w112 = ~w1133 & w454;
assign w113 = ~w893 & ~w536;
assign w114 = (w283 & w219) | (w283 & w1008) | (w219 & w1008);
assign w115 = w1128 & w1138;
assign w116 = b43 & a43;
assign w117 = (w91 & w898) | (w91 & w769) | (w898 & w769);
assign w118 = ~w474 & ~w930;
assign w119 = ~w756 & ~w1068;
assign w120 = ~w164 & w1042;
assign w121 = (w284 & w689) | (w284 & w55) | (w689 & w55);
assign w122 = w225 & ~w83;
assign w123 = ~w317 & w269;
assign w124 = b38 & a38;
assign w125 = (~w898 & w972) | (~w898 & w990) | (w972 & w990);
assign w126 = ~w154 & ~w706;
assign w127 = w563 & ~w106;
assign w128 = (w1081 & w574) | (w1081 & ~w278) | (w574 & ~w278);
assign w129 = ~w844 & ~w854;
assign w130 = w474 & w53;
assign w131 = (~w298 & w729) | (~w298 & w599) | (w729 & w599);
assign w132 = ~w55 & w710;
assign w133 = (~w1103 & ~w1019) | (~w1103 & ~w752) | (~w1019 & ~w752);
assign w134 = w402 & ~w901;
assign w135 = ~w819 & ~w1146;
assign w136 = ~w733 & w446;
assign w137 = ~w201 & ~w467;
assign w138 = w796 & w223;
assign w139 = w79 & w323;
assign w140 = ~w13 & w1095;
assign w141 = (~w829 & w1090) | (~w829 & w738) | (w1090 & w738);
assign w142 = ~b38 & ~a38;
assign w143 = ~b16 & ~a16;
assign w144 = (~w1101 & w88) | (~w1101 & w1075) | (w88 & w1075);
assign w145 = (~w996 & w1021) | (~w996 & w612) | (w1021 & w612);
assign w146 = ~w476 & ~w663;
assign w147 = ~w784 & ~w954;
assign w148 = ~w248 & ~w1056;
assign w149 = w881 & w400;
assign w150 = (~w509 & ~w552) | (~w509 & w50) | (~w552 & w50);
assign w151 = ~w349 & ~w984;
assign w152 = (w692 & w308) | (w692 & w422) | (w308 & w422);
assign w153 = ~w279 & ~w624;
assign w154 = ~b30 & ~a30;
assign w155 = (w540 & w518) | (w540 & w416) | (w518 & w416);
assign w156 = (~w77 & w856) | (~w77 & w52) | (w856 & w52);
assign w157 = ~w74 & ~w239;
assign w158 = (w531 & w213) | (w531 & w155) | (w213 & w155);
assign w159 = (~w531 & w537) | (~w531 & w1117) | (w537 & w1117);
assign w160 = (~w683 & ~w381) | (~w683 & ~w830) | (~w381 & ~w830);
assign w161 = (w531 & w730) | (w531 & w1017) | (w730 & w1017);
assign w162 = ~w594 & ~w488;
assign w163 = w581 & w981;
assign w164 = ~w664 & ~w623;
assign w165 = (w531 & w561) | (w531 & w1001) | (w561 & w1001);
assign w166 = (w987 & w841) | (w987 & ~w769) | (w841 & ~w769);
assign w167 = (w938 & w732) | (w938 & w805) | (w732 & w805);
assign w168 = w500 & ~w898;
assign w169 = (w17 & w716) | (w17 & w465) | (w716 & w465);
assign w170 = ~w485 & ~w303;
assign w171 = w286 & ~w568;
assign w172 = w1036 & ~w582;
assign w173 = (w133 & w1096) | (w133 & w584) | (w1096 & w584);
assign w174 = ~w298 & w803;
assign w175 = ~w235 & ~w531;
assign w176 = ~w1029 & ~w444;
assign w177 = ~w115 & ~w410;
assign w178 = w202 & w373;
assign w179 = (w653 & ~w1102) | (w653 & w54) | (~w1102 & w54);
assign w180 = (w749 & w762) | (w749 & w278) | (w762 & w278);
assign w181 = w382 & ~w642;
assign w182 = b36 & a36;
assign w183 = (w31 & w733) | (w31 & w771) | (w733 & w771);
assign w184 = ~w862 & ~w24;
assign w185 = (w53 & w130) | (w53 & ~w79) | (w130 & ~w79);
assign w186 = (~w824 & w740) | (~w824 & w1085) | (w740 & w1085);
assign w187 = ~b60 & ~a60;
assign w188 = (w482 & w316) | (w482 & ~w531) | (w316 & ~w531);
assign w189 = b46 & a46;
assign w190 = (w82 & ~w379) | (w82 & ~w518) | (~w379 & ~w518);
assign w191 = ~w296 & w535;
assign w192 = (w731 & w592) | (w731 & w813) | (w592 & w813);
assign w193 = ~w582 & ~w581;
assign w194 = ~b35 & ~a35;
assign w195 = ~w991 & ~w550;
assign w196 = (w531 & w977) | (w531 & w1057) | (w977 & w1057);
assign w197 = ~w661 & ~w719;
assign w198 = w1130 & ~w510;
assign w199 = (w329 & ~w1015) | (w329 & w10) | (~w1015 & w10);
assign w200 = (w533 & w301) | (w533 & ~w505) | (w301 & ~w505);
assign w201 = (w711 & w658) | (w711 & w974) | (w658 & w974);
assign w202 = ~w247 & ~w620;
assign w203 = w709 & w1140;
assign w204 = (~w534 & w621) | (~w534 & w249) | (w621 & w249);
assign w205 = ~w646 & ~w80;
assign w206 = ~w806 & ~w818;
assign w207 = ~b8 & ~a8;
assign w208 = b53 & a53;
assign w209 = (w876 & w596) | (w876 & ~w278) | (w596 & ~w278);
assign w210 = ~w495 & ~w1099;
assign w211 = b60 & a60;
assign w212 = (~w528 & w867) | (~w528 & w655) | (w867 & w655);
assign w213 = (w540 & w824) | (w540 & w416) | (w824 & w416);
assign w214 = ~w1133 & w493;
assign w215 = w1140 & ~w1015;
assign w216 = ~w25 & ~w83;
assign w217 = ~w17 & w904;
assign w218 = w844 & w190;
assign w219 = w74 & w283;
assign w220 = (~w759 & ~w981) | (~w759 & w807) | (~w981 & w807);
assign w221 = (w195 & w458) | (w195 & w278) | (w458 & w278);
assign w222 = ~w142 & ~w62;
assign w223 = ~w154 & ~w811;
assign w224 = ~w597 & ~w952;
assign w225 = w1155 & ~w637;
assign w226 = (w531 & w426) | (w531 & w1040) | (w426 & w1040);
assign w227 = (w1042 & w816) | (w1042 & w120) | (w816 & w120);
assign w228 = (w77 & w1027) | (w77 & w590) | (w1027 & w590);
assign w229 = (w981 & w163) | (w981 & ~w582) | (w163 & ~w582);
assign w230 = w307 & w1118;
assign w231 = ~w498 & ~w161;
assign w232 = ~w105 & ~w315;
assign w233 = ~w292 & ~w723;
assign w234 = (w663 & w866) | (w663 & w17) | (w866 & w17);
assign w235 = w485 & w433;
assign w236 = ~w875 & ~w897;
assign w237 = w32 & ~w675;
assign w238 = (w118 & ~w95) | (w118 & w603) | (~w95 & w603);
assign w239 = ~b49 & ~a49;
assign w240 = w519 & w345;
assign w241 = w131 & ~w746;
assign w242 = ~w156 & ~w1028;
assign w243 = ~w693 & ~w938;
assign w244 = (w67 & w121) | (w67 & ~w1019) | (w121 & ~w1019);
assign w245 = w713 & ~w370;
assign w246 = (~w365 & w272) | (~w365 & w320) | (w272 & w320);
assign w247 = b58 & a58;
assign w248 = ~b18 & ~a18;
assign w249 = (w760 & w828) | (w760 & w291) | (w828 & w291);
assign w250 = ~w745 & ~w456;
assign w251 = ~w178 & w1005;
assign w252 = w900 & ~w568;
assign w253 = w1102 & w695;
assign w254 = w32 & ~w568;
assign w255 = ~b15 & ~a15;
assign w256 = (~w77 & w1038) | (~w77 & w579) | (w1038 & w579);
assign w257 = (~w582 & w528) | (~w582 & w172) | (w528 & w172);
assign w258 = ~w843 & ~w1100;
assign w259 = (w257 & w868) | (w257 & w460) | (w868 & w460);
assign w260 = ~w743 & ~w269;
assign w261 = ~w324 & ~w560;
assign w262 = ~w410 & w1064;
assign w263 = b12 & a12;
assign w264 = ~w95 & w294;
assign w265 = ~w507 & ~w207;
assign w266 = ~w906 & ~w618;
assign w267 = w382 & ~w559;
assign w268 = (w829 & w515) | (w829 & w802) | (w515 & w802);
assign w269 = b5 & a5;
assign w270 = b21 & a21;
assign w271 = ~w951 & ~w736;
assign w272 = w907 & ~w731;
assign w273 = (~w518 & w740) | (~w518 & w1085) | (w740 & w1085);
assign w274 = (~w85 & w881) | (~w85 & w613) | (w881 & w613);
assign w275 = ~b40 & ~a40;
assign w276 = w378 & w961;
assign w277 = ~w380 & w726;
assign w278 = ~w89 & w613;
assign w279 = b10 & a10;
assign w280 = w1137 & ~w1069;
assign w281 = (w987 & w841) | (w987 & ~w1101) | (w841 & ~w1101);
assign w282 = w519 & w461;
assign w283 = ~w843 & ~w496;
assign w284 = ~w767 & ~w620;
assign w285 = ~w962 & w27;
assign w286 = w373 & w98;
assign w287 = ~w761 & ~w861;
assign w288 = (w150 & w493) | (w150 & ~w742) | (w493 & ~w742);
assign w289 = w250 & w754;
assign w290 = ~w847 & ~w1080;
assign w291 = ~w296 & w210;
assign w292 = (~w658 & w696) | (~w658 & w735) | (w696 & w735);
assign w293 = ~w547 & ~w196;
assign w294 = ~w474 & ~w53;
assign w295 = ~w421 & w958;
assign w296 = w953 & w520;
assign w297 = w710 & w1103;
assign w298 = ~w513 & ~w927;
assign w299 = ~w74 & ~w283;
assign w300 = (~w1080 & ~w1112) | (~w1080 & w616) | (~w1112 & w616);
assign w301 = (~w448 & w314) | (~w448 & w533) | (w314 & w533);
assign w302 = ~w349 & ~w269;
assign w303 = b26 & a26;
assign w304 = b17 & a17;
assign w305 = ~w485 & ~w786;
assign w306 = w184 & w469;
assign w307 = w62 & w726;
assign w308 = w206 & ~w818;
assign w309 = w993 & w250;
assign w310 = w807 & w582;
assign w311 = (~w531 & w464) | (~w531 & w942) | (w464 & w942);
assign w312 = (~w531 & w44) | (~w531 & w791) | (w44 & w791);
assign w313 = (~w518 & w122) | (~w518 & w1007) | (w122 & w1007);
assign w314 = ~w25 & w380;
assign w315 = b24 & a24;
assign w316 = (~w769 & w1151) | (~w769 & w966) | (w1151 & w966);
assign w317 = ~b6 & ~a6;
assign w318 = b18 & a18;
assign w319 = ~w851 & ~w1093;
assign w320 = w907 & ~w192;
assign w321 = w175 & ~w376;
assign w322 = (~w786 & ~w433) | (~w786 & w305) | (~w433 & w305);
assign w323 = w560 & w118;
assign w324 = ~b32 & ~a32;
assign w325 = (w569 & w824) | (w569 & w895) | (w824 & w895);
assign w326 = w767 & ~w677;
assign w327 = (~w531 & w436) | (~w531 & w313) | (w436 & w313);
assign w328 = (~w752 & w461) | (~w752 & w345) | (w461 & w345);
assign w329 = ~w940 & ~w737;
assign w330 = w286 & ~w675;
assign w331 = w1020 & ~w59;
assign w332 = ~w860 & ~w68;
assign w333 = ~w783 & ~w861;
assign w334 = ~w287 & w720;
assign w335 = ~w754 & w888;
assign w336 = ~w77 & w853;
assign w337 = ~w1018 & ~w1056;
assign w338 = ~w940 & ~w575;
assign w339 = (~w278 & w555) | (~w278 & w356) | (w555 & w356);
assign w340 = w989 & ~w998;
assign w341 = (w77 & w483) | (w77 & w980) | (w483 & w980);
assign w342 = ~w189 & ~w711;
assign w343 = ~w361 & w627;
assign w344 = (w952 & ~w312) | (w952 & w1115) | (~w312 & w1115);
assign w345 = (~w728 & w1053) | (~w728 & w461) | (w1053 & w461);
assign w346 = ~w485 & ~w433;
assign w347 = (w726 & w25) | (w726 & w277) | (w25 & w277);
assign w348 = (w236 & w957) | (w236 & w643) | (w957 & w643);
assign w349 = ~w743 & ~w317;
assign w350 = ~w509 & w588;
assign w351 = ~w207 & ~w862;
assign w352 = (~w531 & w983) | (~w531 & w705) | (w983 & w705);
assign w353 = (~w752 & w1090) | (~w752 & w738) | (w1090 & w738);
assign w354 = w18 & ~w410;
assign w355 = (~w658 & w702) | (~w658 & w29) | (w702 & w29);
assign w356 = (w31 & w183) | (w31 & w215) | (w183 & w215);
assign w357 = w909 & w153;
assign w358 = w747 & ~w569;
assign w359 = (~w742 & w429) | (~w742 & w214) | (w429 & w214);
assign w360 = (w658 & w141) | (w658 & w353) | (w141 & w353);
assign w361 = ~w783 & ~w939;
assign w362 = ~w693 & ~w304;
assign w363 = (w742 & w306) | (w742 & w1116) | (w306 & w1116);
assign w364 = ~a1 & ~w608;
assign w365 = (w1076 & ~w1008) | (w1076 & w870) | (~w1008 & w870);
assign w366 = w136 & ~w215;
assign w367 = (w864 & w309) | (w864 & w992) | (w309 & w992);
assign w368 = (w1140 & ~w1015) | (w1140 & w203) | (~w1015 & w203);
assign w369 = ~w708 & w148;
assign w370 = w1133 & ~w493;
assign w371 = ~w1132 & w559;
assign w372 = ~w993 & ~w745;
assign w373 = ~w767 & w677;
assign w374 = (w883 & w93) | (w883 & w925) | (w93 & w925);
assign w375 = w792 & w455;
assign w376 = (~w339 & w34) | (~w339 & w669) | (w34 & w669);
assign w377 = w583 & ~w8;
assign w378 = ~w693 & ~w143;
assign w379 = (~w854 & w1012) | (~w854 & w505) | (w1012 & w505);
assign w380 = ~w453 & ~w1044;
assign w381 = (~w743 & w666) | (~w743 & ~w984) | (w666 & ~w984);
assign w382 = ~w796 & ~w223;
assign w383 = (w976 & w1039) | (w976 & ~w1101) | (w1039 & ~w1101);
assign w384 = (w77 & w1124) | (w77 & w963) | (w1124 & w963);
assign w385 = (w329 & w85) | (w329 & w614) | (w85 & w614);
assign w386 = ~w915 & ~w525;
assign w387 = ~w617 & ~w662;
assign w388 = ~w991 & ~w0;
assign w389 = w311 & ~w1006;
assign w390 = (w288 & w964) | (w288 & w685) | (w964 & w685);
assign w391 = w1133 & ~w150;
assign w392 = (w195 & w458) | (w195 & w613) | (w458 & w613);
assign w393 = (~w996 & w272) | (~w996 & w320) | (w272 & w320);
assign w394 = w1136 & ~w622;
assign w395 = ~w450 & w842;
assign w396 = (w913 & w838) | (w913 & w1025) | (w838 & w1025);
assign w397 = (~w439 & w449) | (~w439 & w63) | (w449 & w63);
assign w398 = (w692 & w549) | (w692 & w511) | (w549 & w511);
assign w399 = (w984 & w1122) | (w984 & w391) | (w1122 & w391);
assign w400 = ~w1062 & ~w795;
assign w401 = (w637 & w36) | (w637 & w505) | (w36 & w505);
assign w402 = (~w309 & w658) | (~w309 & w670) | (w658 & w670);
assign w403 = (w654 & w16) | (w654 & w1065) | (w16 & w1065);
assign w404 = ~w1113 & ~w918;
assign w405 = w349 & w984;
assign w406 = b41 & a41;
assign w407 = (~w518 & w64) | (~w518 & w517) | (w64 & w517);
assign w408 = (~w658 & w252) | (~w658 & w1114) | (w252 & w1114);
assign w409 = (~w769 & w577) | (~w769 & w1135) | (w577 & w1135);
assign w410 = (w7 & w91) | (w7 & w727) | (w91 & w727);
assign w411 = (~w257 & w751) | (~w257 & w459) | (w751 & w459);
assign w412 = w929 & w909;
assign w413 = ~w484 & ~w81;
assign w414 = w1030 & ~w886;
assign w415 = ~w1036 & ~w581;
assign w416 = ~w750 & w540;
assign w417 = (w77 & w633) | (w77 & w595) | (w633 & w595);
assign w418 = (w205 & w985) | (w205 & w752) | (w985 & w752);
assign w419 = (~w531 & w441) | (~w531 & w591) | (w441 & w591);
assign w420 = (w77 & w274) | (w77 & w1154) | (w274 & w1154);
assign w421 = (~w495 & ~w520) | (~w495 & w12) | (~w520 & w12);
assign w422 = (~w818 & w206) | (~w818 & w55) | (w206 & w55);
assign w423 = (~w658 & w179) | (~w658 & w859) | (w179 & w859);
assign w424 = (w146 & w494) | (w146 & w686) | (w494 & w686);
assign w425 = w126 & w942;
assign w426 = (w932 & w424) | (w932 & w1101) | (w424 & w1101);
assign w427 = w875 & w645;
assign w428 = (w387 & w822) | (w387 & w996) | (w822 & w996);
assign w429 = ~w1133 & w150;
assign w430 = ~w847 & w651;
assign w431 = (~w673 & ~w883) | (~w673 & ~w381) | (~w883 & ~w381);
assign w432 = ~w583 & w8;
assign w433 = ~w786 & ~w530;
assign w434 = ~w1100 & ~w1139;
assign w435 = ~w957 & ~w518;
assign w436 = w225 & ~w1101;
assign w437 = ~w546 & ~w232;
assign w438 = w710 & ~w675;
assign w439 = (w278 & w790) | (w278 & w366) | (w790 & w366);
assign w440 = ~w624 & w104;
assign w441 = (w169 & w615) | (w169 & ~w1101) | (w615 & ~w1101);
assign w442 = (~w829 & w797) | (~w829 & w23) | (w797 & w23);
assign w443 = (w133 & w308) | (w133 & w422) | (w308 & w422);
assign w444 = ~b13 & ~a13;
assign w445 = ~b4 & ~a4;
assign w446 = ~w105 & ~w848;
assign w447 = ~w194 & ~w453;
assign w448 = w142 & w62;
assign w449 = w916 & ~w77;
assign w450 = w14 & ~w1066;
assign w451 = (w133 & w48) | (w133 & w631) | (w48 & w631);
assign w452 = ~w945 & ~w894;
assign w453 = ~b36 & ~a36;
assign w454 = ~w971 & ~w269;
assign w455 = b28 & a28;
assign w456 = b48 & a48;
assign w457 = w1026 & ~w440;
assign w458 = ~w111 & w195;
assign w459 = w243 & ~w805;
assign w460 = (w805 & w290) | (w805 & w668) | (w290 & w668);
assign w461 = ~w728 & ~w1103;
assign w462 = (~w24 & w679) | (~w24 & w683) | (w679 & w683);
assign w463 = b47 & a47;
assign w464 = ~w138 & ~w79;
assign w465 = (w663 & w866) | (w663 & ~w307) | (w866 & ~w307);
assign w466 = (w77 & w229) | (w77 & w933) | (w229 & w933);
assign w467 = ~w658 & w342;
assign w468 = (w284 & w689) | (w284 & w568) | (w689 & w568);
assign w469 = (~w683 & ~w381) | (~w683 & ~w629) | (~w381 & ~w629);
assign w470 = (w531 & w548) | (w531 & w1052) | (w548 & w1052);
assign w471 = w14 & w350;
assign w472 = (w1012 & w1010) | (w1012 & w978) | (w1010 & w978);
assign w473 = (~w1100 & ~w33) | (~w1100 & w258) | (~w33 & w258);
assign w474 = b31 & a31;
assign w475 = ~b0 & ~a0;
assign w476 = b40 & a40;
assign w477 = ~w1062 & ~w845;
assign w478 = w289 & w299;
assign w479 = ~w476 & ~w275;
assign w480 = (~w1080 & ~w1112) | (~w1080 & ~w582) | (~w1112 & ~w582);
assign w481 = ~w571 & ~w887;
assign w482 = (~w610 & ~w801) | (~w610 & ~w534) | (~w801 & ~w534);
assign w483 = ~w708 & ~w414;
assign w484 = (w575 & w384) | (w575 & w567) | (w384 & w567);
assign w485 = ~b26 & ~a26;
assign w486 = ~w646 & ~w623;
assign w487 = ~w563 & w106;
assign w488 = (w563 & w457) | (w563 & w923) | (w457 & w923);
assign w489 = ~b46 & ~a46;
assign w490 = ~w269 & ~w984;
assign w491 = ~w1132 & ~w455;
assign w492 = (w658 & w468) | (w658 & w973) | (w468 & w973);
assign w493 = ~w509 & ~w552;
assign w494 = ~w314 & w307;
assign w495 = ~b42 & ~a42;
assign w496 = b50 & a50;
assign w497 = ~w106 & ~w104;
assign w498 = (~w531 & w375) | (~w531 & w1121) | (w375 & w1121);
assign w499 = ~w578 & ~w37;
assign w500 = w421 & ~w958;
assign w501 = w261 & ~w522;
assign w502 = ~w109 & ~w1077;
assign w503 = ~w210 & w610;
assign w504 = (~w654 & w630) | (~w654 & w798) | (w630 & w798);
assign w505 = ~w750 & w83;
assign w506 = ~cin & ~w30;
assign w507 = b8 & a8;
assign w508 = ~b58 & ~a58;
assign w509 = b3 & a3;
assign w510 = (w658 & w678) | (w658 & w647) | (w678 & w647);
assign w511 = (w979 & w96) | (w979 & w55) | (w96 & w55);
assign w512 = (~w518 & w216) | (~w518 & w982) | (w216 & w982);
assign w513 = ~a63 & ~b63;
assign w514 = (~w531 & w102) | (~w531 & w46) | (w102 & w46);
assign w515 = (w710 & ~w55) | (w710 & w297) | (~w55 & w297);
assign w516 = (w133 & w549) | (w133 & w511) | (w549 & w511);
assign w517 = (w88 & w1075) | (w88 & ~w505) | (w1075 & ~w505);
assign w518 = (w323 & w846) | (w323 & w812) | (w846 & w812);
assign w519 = ~w661 & ~w593;
assign w520 = ~w495 & ~w850;
assign w521 = ~w89 & w911;
assign w522 = (w118 & w138) | (w118 & w688) | (w138 & w688);
assign w523 = w1030 & w809;
assign w524 = (w563 & w855) | (w563 & w331) | (w855 & w331);
assign w525 = ~w703 & w602;
assign w526 = w929 & ~w263;
assign w527 = (w593 & w65) | (w593 & ~w345) | (w65 & ~w345);
assign w528 = w611 & ~w357;
assign w529 = ~w795 & w878;
assign w530 = b27 & a27;
assign w531 = (~w77 & w1105) | (~w77 & w128) | (w1105 & w128);
assign w532 = (~b1 & w506) | (~b1 & w598) | (w506 & w598);
assign w533 = ~w448 & ~w307;
assign w534 = (w91 & w898) | (w91 & w1101) | (w898 & w1101);
assign w535 = (~w531 & ~w534) | (~w531 & ~w117) | (~w534 & ~w117);
assign w536 = (~w531 & w652) | (~w531 & w425) | (w652 & w425);
assign w537 = (w1125 & w1108) | (w1125 & ~w824) | (w1108 & ~w824);
assign w538 = (w658 & w674) | (w658 & w914) | (w674 & w914);
assign w539 = w287 & w783;
assign w540 = ~w875 & ~w645;
assign w541 = w157 & ~w943;
assign w542 = ~w380 & ~w854;
assign w543 = w589 & ~w360;
assign w544 = ~w581 & ~w981;
assign w545 = ~w709 & w1015;
assign w546 = ~b23 & ~a23;
assign w547 = (~w531 & w607) | (~w531 & w218) | (w607 & w218);
assign w548 = (w958 & w295) | (w958 & w534) | (w295 & w534);
assign w549 = w96 & w979;
assign w550 = ~w1062 & ~w270;
assign w551 = ~b17 & ~a17;
assign w552 = ~w1061 & ~w509;
assign w553 = (~w752 & w282) | (~w752 & w240) | (w282 & w240);
assign w554 = ~w745 & ~w239;
assign w555 = (w31 & w183) | (w31 & w368) | (w183 & w368);
assign w556 = w701 & w286;
assign w557 = ~b2 & ~a2;
assign w558 = (~w269 & ~w984) | (~w269 & w454) | (~w984 & w454);
assign w559 = ~w455 & ~w1082;
assign w560 = ~w756 & ~w1106;
assign w561 = (w637 & w36) | (w637 & w1101) | (w36 & w1101);
assign w562 = b44 & a44;
assign w563 = w763 & ~w671;
assign w564 = (w909 & w412) | (w909 & w440) | (w412 & w440);
assign w565 = ~w1144 & ~w524;
assign w566 = ~w778 & ~w479;
assign w567 = w940 & w575;
assign w568 = (~w829 & w912) | (~w829 & w43) | (w912 & w43);
assign w569 = ~w875 & ~w1068;
assign w570 = w219 & w283;
assign w571 = (w531 & w1013) | (w531 & w1037) | (w1013 & w1037);
assign w572 = w514 & ~w1092;
assign w573 = (w938 & w732) | (w938 & ~w582) | (w732 & ~w582);
assign w574 = (w779 & w215) | (w779 & w814) | (w215 & w814);
assign w575 = ~w546 & ~w737;
assign w576 = ~w693 & w582;
assign w577 = (w621 & w249) | (w621 & ~w91) | (w249 & ~w91);
assign w578 = (w742 & w399) | (w742 & w1047) | (w399 & w1047);
assign w579 = w934 & ~w278;
assign w580 = w778 & w479;
assign w581 = b14 & a14;
assign w582 = ~b14 & ~a14;
assign w583 = (w77 & w920) | (w77 & w180) | (w920 & w180);
assign w584 = (w1005 & w251) | (w1005 & w55) | (w251 & w55);
assign w585 = ~w733 & ~w368;
assign w586 = w670 & w772;
assign w587 = (~w752 & w797) | (~w752 & w23) | (w797 & w23);
assign w588 = ~w971 & ~w35;
assign w589 = (w658 & w891) | (w658 & w328) | (w891 & w328);
assign w590 = (w257 & w755) | (w257 & w167) | (w755 & w167);
assign w591 = (w169 & w615) | (w169 & ~w769) | (w615 & ~w769);
assign w592 = w843 & w33;
assign w593 = ~w247 & ~w508;
assign w594 = (~w563 & w564) | (~w563 & w1091) | (w564 & w1091);
assign w595 = (w278 & w837) | (w278 & w1016) | (w837 & w1016);
assign w596 = (w795 & ~w881) | (w795 & w60) | (~w881 & w60);
assign w597 = ~b45 & ~a45;
assign w598 = w475 & ~b1;
assign w599 = w861 & ~w298;
assign w600 = w265 & w24;
assign w601 = ~w800 & ~w336;
assign w602 = ~w532 & ~w90;
assign w603 = w79 & w118;
assign w604 = w844 & ~w1012;
assign w605 = ~w104 & w611;
assign w606 = (w654 & w107) | (w654 & w374) | (w107 & w374);
assign w607 = (~w1101 & w776) | (~w1101 & w604) | (w776 & w604);
assign w608 = ~w997 & ~w532;
assign w609 = (w151 & w302) | (w151 & w629) | (w302 & w629);
assign w610 = ~w116 & ~w562;
assign w611 = ~w526 & w176;
assign w612 = (w662 & w1094) | (w662 & w13) | (w1094 & w13);
assign w613 = w369 & ~w414;
assign w614 = ~w477 & w329;
assign w615 = (~w494 & w716) | (~w494 & w234) | (w716 & w234);
assign w616 = (~w143 & w981) | (~w143 & w1127) | (w981 & w1127);
assign w617 = b52 & a52;
assign w618 = (w658 & w41) | (w658 & w173) | (w41 & w173);
assign w619 = ~w743 & ~w184;
assign w620 = b59 & a59;
assign w621 = w828 & w760;
assign w622 = (~w531 & w186) | (~w531 & w273) | (w186 & w273);
assign w623 = ~b55 & ~a55;
assign w624 = b11 & a11;
assign w625 = w1109 & ~w683;
assign w626 = w713 & ~w391;
assign w627 = (~w211 & ~w677) | (~w211 & w787) | (~w677 & w787);
assign w628 = (w479 & w580) | (w479 & ~w533) | (w580 & ~w533);
assign w629 = (w454 & w493) | (w454 & w112) | (w493 & w112);
assign w630 = (~w883 & w625) | (~w883 & w69) | (w625 & w69);
assign w631 = (w684 & w700) | (w684 & w55) | (w700 & w55);
assign w632 = ~w116 & ~w760;
assign w633 = w437 & w1011;
assign w634 = b51 & a51;
assign w635 = ~w35 & ~w552;
assign w636 = ~b56 & ~a56;
assign w637 = ~w854 & ~w1044;
assign w638 = (w56 & w585) | (w56 & w278) | (w585 & w278);
assign w639 = ~w1086 & ~w104;
assign w640 = (w77 & w276) | (w77 & w947) | (w276 & w947);
assign w641 = (w77 & w430) | (w77 & w259) | (w430 & w259);
assign w642 = (w559 & w235) | (w559 & w371) | (w235 & w371);
assign w643 = ~w119 & w236;
assign w644 = b54 & a54;
assign w645 = ~w194 & ~w897;
assign w646 = b55 & a55;
assign w647 = (w692 & w241) | (w692 & w908) | (w241 & w908);
assign w648 = w1036 & w193;
assign w649 = ~w355 & ~w766;
assign w650 = (w299 & ~w1008) | (w299 & w478) | (~w1008 & w478);
assign w651 = (w805 & w480) | (w805 & w300) | (w480 & w300);
assign w652 = w126 & w464;
assign w653 = ~w617 & ~w1139;
assign w654 = (~w742 & w830) | (~w742 & w629) | (w830 & w629);
assign w655 = w544 & ~w172;
assign w656 = b56 & a56;
assign w657 = w694 & w188;
assign w658 = (~w531 & w1145) | (~w531 & w1049) | (w1145 & w1049);
assign w659 = w420 & ~w1059;
assign w660 = (w533 & w301) | (w533 & ~w83) | (w301 & ~w83);
assign w661 = ~b57 & ~a57;
assign w662 = ~w872 & ~w208;
assign w663 = ~w953 & ~w406;
assign w664 = ~b54 & ~a54;
assign w665 = (w1003 & w168) | (w1003 & ~w1101) | (w168 & ~w1101);
assign w666 = ~w349 & ~w743;
assign w667 = w1123 & ~w351;
assign w668 = ~w847 & ~w1112;
assign w669 = (w913 & w1031) | (w913 & w61) | (w1031 & w61);
assign w670 = ~w289 & ~w309;
assign w671 = ~w742 & w471;
assign w672 = ~w453 & ~w182;
assign w673 = (~w507 & ~w265) | (~w507 & w1147) | (~w265 & w1147);
assign w674 = ~w816 & ~w829;
assign w675 = (~w752 & w912) | (~w752 & w43) | (w912 & w43);
assign w676 = ~w184 & w683;
assign w677 = ~w211 & ~w187;
assign w678 = (w133 & w241) | (w133 & w908) | (w241 & w908);
assign w679 = ~w184 & ~w24;
assign w680 = ~w127 & ~w487;
assign w681 = (~w658 & w38) | (~w658 & w428) | (w38 & w428);
assign w682 = w807 & ~w172;
assign w683 = (~w743 & ~w349) | (~w743 & w260) | (~w349 & w260);
assign w684 = ~w373 & ~w326;
assign w685 = (w676 & w885) | (w676 & w112) | (w885 & w112);
assign w686 = ~w17 & w146;
assign w687 = (~w624 & w106) | (~w624 & w440) | (w106 & w440);
assign w688 = ~w717 & w118;
assign w689 = w247 & w284;
assign w690 = (~w77 & w865) | (~w77 & w890) | (w865 & w890);
assign w691 = ~w455 & ~w1;
assign w692 = (~w1103 & ~w1019) | (~w1103 & ~w829) | (~w1019 & ~w829);
assign w693 = b16 & a16;
assign w694 = ~w1128 & ~w1138;
assign w695 = ~w1100 & ~w653;
assign w696 = (w486 & w1079) | (w486 & w752) | (w1079 & w752);
assign w697 = (w981 & w163) | (w981 & w172) | (w163 & w172);
assign w698 = ~w1022 & ~w780;
assign w699 = (~w664 & ~w879) | (~w664 & w968) | (~w879 & w968);
assign w700 = ~w202 & w684;
assign w701 = (w627 & w66) | (w627 & w334) | (w66 & w334);
assign w702 = (w752 & w75) | (w752 & w527) | (w75 & w527);
assign w703 = ~a1 & ~w997;
assign w704 = (~w759 & ~w981) | (~w759 & w682) | (~w981 & w682);
assign w705 = w358 & ~w518;
assign w706 = ~w474 & ~w877;
assign w707 = ~w287 & w19;
assign w708 = w551 & w847;
assign w709 = w550 & w111;
assign w710 = ~w247 & ~w284;
assign w711 = ~w993 & ~w463;
assign w712 = (w151 & w302) | (w151 & w830) | (w302 & w830);
assign w713 = ~w971 & ~w984;
assign w714 = ~w752 & w1063;
assign w715 = ~w991 & ~w1062;
assign w716 = w866 & w663;
assign w717 = ~w154 & ~w877;
assign w718 = ~w1036 & ~w444;
assign w719 = b57 & a57;
assign w720 = w939 & ~w783;
assign w721 = w1067 & ~w417;
assign w722 = ~w324 & ~w756;
assign w723 = (w658 & w758) | (w658 & w714) | (w758 & w714);
assign w724 = w298 & w32;
assign w725 = ~w157 & w943;
assign w726 = ~w854 & ~w124;
assign w727 = ~w291 & w7;
assign w728 = w636 & w197;
assign w729 = (~w627 & w539) | (~w627 & w1058) | (w539 & w1058);
assign w730 = ~w792 & ~w455;
assign w731 = ~w617 & ~w208;
assign w732 = w693 & w938;
assign w733 = w546 & w232;
assign w734 = (w569 & w518) | (w569 & w895) | (w518 & w895);
assign w735 = (w486 & w1079) | (w486 & w829) | (w1079 & w829);
assign w736 = (w531 & w871) | (w531 & w9) | (w871 & w9);
assign w737 = b23 & a23;
assign w738 = w825 & ~w227;
assign w739 = (w1118 & ~w17) | (w1118 & w230) | (~w17 & w230);
assign w740 = w782 & ~w236;
assign w741 = (w976 & w1039) | (w976 & ~w769) | (w1039 & ~w769);
assign w742 = ~w703 & w950;
assign w743 = b6 & a6;
assign w744 = ~b9 & ~a9;
assign w745 = ~b48 & ~a48;
assign w746 = w32 & ~w174;
assign w747 = (~w756 & ~w560) | (~w756 & w722) | (~w560 & w722);
assign w748 = ~w475 & ~w30;
assign w749 = ~w368 & w1002;
assign w750 = ~w957 & w119;
assign w751 = w243 & ~w616;
assign w752 = (w1095 & w365) | (w1095 & w140) | (w365 & w140);
assign w753 = (w742 & w905) | (w742 & w1143) | (w905 & w1143);
assign w754 = ~w189 & ~w463;
assign w755 = (w938 & w732) | (w938 & w616) | (w732 & w616);
assign w756 = ~b33 & ~a33;
assign w757 = w745 & w157;
assign w758 = ~w829 & w1063;
assign w759 = b15 & a15;
assign w760 = ~w1128 & ~w562;
assign w761 = ~b62 & ~a62;
assign w762 = ~w105 & w56;
assign w763 = ~w450 & w1089;
assign w764 = ~w473 & w653;
assign w765 = (~w769 & w1051) | (~w769 & w1157) | (w1051 & w1157);
assign w766 = (w658 & w553) | (w658 & w1043) | (w553 & w1043);
assign w767 = ~b59 & ~a59;
assign w768 = ~w265 & ~w24;
assign w769 = (w83 & w518) | (w83 & w505) | (w518 & w505);
assign w770 = (~w365 & w1021) | (~w365 & w612) | (w1021 & w612);
assign w771 = ~w446 & w31;
assign w772 = ~w745 & ~w157;
assign w773 = w261 & ~w238;
assign w774 = (w262 & w125) | (w262 & ~w769) | (w125 & ~w769);
assign w775 = ~w944 & ~w364;
assign w776 = w844 & w854;
assign w777 = w307 & w146;
assign w778 = ~b39 & ~a39;
assign w779 = w433 & w31;
assign w780 = ~w531 & w832;
assign w781 = w71 & ~w57;
assign w782 = ~w194 & ~w672;
assign w783 = b61 & a61;
assign w784 = (w563 & w639) | (w563 & w995) | (w639 & w995);
assign w785 = ~w1036 & ~w193;
assign w786 = ~b27 & ~a27;
assign w787 = w767 & ~w211;
assign w788 = w312 & ~w657;
assign w789 = (w529 & w149) | (w529 & w613) | (w149 & w613);
assign w790 = w136 & ~w368;
assign w791 = (w28 & w177) | (w28 & ~w769) | (w177 & ~w769);
assign w792 = ~w796 & ~w1082;
assign w793 = ~w661 & ~w508;
assign w794 = ~w475 & b1;
assign w795 = ~w940 & ~w845;
assign w796 = ~b29 & ~a29;
assign w797 = w926 & w80;
assign w798 = w1109 & w431;
assign w799 = w538 & ~w103;
assign w800 = (w193 & w77) | (w193 & w1107) | (w77 & w1107);
assign w801 = (w610 & w296) | (w610 & w503) | (w296 & w503);
assign w802 = (w710 & w132) | (w710 & w1019) | (w132 & w1019);
assign w803 = ~w761 & ~w333;
assign w804 = ~w265 & ~w507;
assign w805 = ~w143 & ~w220;
assign w806 = ~w803 & w724;
assign w807 = ~w581 & ~w759;
assign w808 = ~w592 & ~w365;
assign w809 = w981 & w415;
assign w810 = (w283 & w219) | (w283 & ~w289) | (w219 & ~w289);
assign w811 = b30 & a30;
assign w812 = ~w95 & w323;
assign w813 = ~w434 & w731;
assign w814 = ~w136 & w779;
assign w815 = ~w344 & ~w1055;
assign w816 = w872 & w879;
assign w817 = ~w25 & ~w1101;
assign w818 = (w19 & ~w1104) | (w19 & w707) | (~w1104 & w707);
assign w819 = (w658 & w114) | (w658 & w100) | (w114 & w100);
assign w820 = (w95 & w931) | (w95 & w185) | (w931 & w185);
assign w821 = ~w743 & ~w24;
assign w822 = ~w13 & w387;
assign w823 = ~w466 & ~w986;
assign w824 = (w323 & ~w95) | (w323 & w139) | (~w95 & w139);
assign w825 = ~w636 & ~w197;
assign w826 = ~w73 & ~w1152;
assign w827 = (w53 & w130) | (w53 & w95) | (w130 & w95);
assign w828 = w116 & w760;
assign w829 = (w1095 & w996) | (w1095 & w140) | (w996 & w140);
assign w830 = (w454 & w150) | (w454 & w112) | (w150 & w112);
assign w831 = ~w938 & w576;
assign w832 = w322 & ~w691;
assign w833 = w35 & w552;
assign w834 = ~w159 & ~w158;
assign w835 = (w479 & w580) | (w479 & ~w301) | (w580 & ~w301);
assign w836 = (w439 & w49) | (w439 & w396) | (w49 & w396);
assign w837 = w437 & ~w385;
assign w838 = w884 & w170;
assign w839 = ~w581 & w582;
assign w840 = (~w846 & w874) | (~w846 & w501) | (w874 & w501);
assign w841 = w291 & ~w898;
assign w842 = w1089 & w605;
assign w843 = ~b50 & ~a50;
assign w844 = ~w142 & ~w124;
assign w845 = ~b22 & ~a22;
assign w846 = ~w921 & w79;
assign w847 = ~w248 & ~w318;
assign w848 = ~b25 & ~a25;
assign w849 = ~w432 & ~w377;
assign w850 = b42 & a42;
assign w851 = (~w658 & w541) | (~w658 & w902) | (w541 & w902);
assign w852 = w18 & ~w7;
assign w853 = ~w528 & w785;
assign w854 = b37 & a37;
assign w855 = w1020 & ~w857;
assign w856 = (w337 & w869) | (w337 & w414) | (w869 & w414);
assign w857 = (~w263 & w526) | (~w263 & w440) | (w526 & w440);
assign w858 = ~w1054 & ~w352;
assign w859 = (w653 & w365) | (w653 & w764) | (w365 & w764);
assign w860 = (w658 & w1129) | (w658 & w451) | (w1129 & w451);
assign w861 = b62 & a62;
assign w862 = ~b7 & ~a7;
assign w863 = (w505 & w129) | (w505 & w1035) | (w129 & w1035);
assign w864 = ~w74 & ~w496;
assign w865 = ~w378 & ~w961;
assign w866 = w476 & w663;
assign w867 = ~w981 & w839;
assign w868 = ~w847 & w300;
assign w869 = ~w1024 & w337;
assign w870 = w289 & w1076;
assign w871 = (w294 & ~w95) | (w294 & w1032) | (~w95 & w1032);
assign w872 = ~b53 & ~a53;
assign w873 = ~w87 & ~w681;
assign w874 = w261 & ~w118;
assign w875 = b34 & a34;
assign w876 = w795 & ~w878;
assign w877 = ~b31 & ~a31;
assign w878 = (~w1062 & ~w550) | (~w1062 & w715) | (~w550 & w715);
assign w879 = ~w664 & ~w644;
assign w880 = ~w365 & w1070;
assign w881 = ~w709 & ~w85;
assign w882 = (w864 & ~w1008) | (w864 & w1126) | (~w1008 & w1126);
assign w883 = (~w507 & w679) | (~w507 & w804) | (w679 & w804);
assign w884 = w1131 & w170;
assign w885 = (w1083 & w666) | (w1083 & w619) | (w666 & w619);
assign w886 = ~w1141 & w965;
assign w887 = (~w531 & w94) | (~w531 & w765) | (w94 & w765);
assign w888 = ~w993 & ~w250;
assign w889 = ~w1008 & w299;
assign w890 = ~w378 & w946;
assign w891 = (~w829 & w461) | (~w829 & w345) | (w461 & w345);
assign w892 = (w56 & w585) | (w56 & w613) | (w585 & w613);
assign w893 = (w531 & w1084) | (w531 & w1023) | (w1084 & w1023);
assign w894 = (~w658 & w418) | (~w658 & w1111) | (w418 & w1111);
assign w895 = ~w747 & w569;
assign w896 = (~w805 & w831) | (~w805 & w751) | (w831 & w751);
assign w897 = b35 & a35;
assign w898 = (w904 & w494) | (w904 & w217) | (w494 & w217);
assign w899 = ~w513 & w1130;
assign w900 = (w286 & w729) | (w286 & w556) | (w729 & w556);
assign w901 = (w888 & w658) | (w888 & w335) | (w658 & w335);
assign w902 = (w157 & ~w670) | (w157 & w757) | (~w670 & w757);
assign w903 = w42 & ~w882;
assign w904 = w520 & w1118;
assign w905 = (~w830 & w40) | (~w830 & w405) | (w40 & w405);
assign w906 = (~w658 & w171) | (~w658 & w330) | (w171 & w330);
assign w907 = ~w872 & ~w879;
assign w908 = w131 & ~w928;
assign w909 = ~w1029 & ~w263;
assign w910 = ~w504 & ~w606;
assign w911 = w78 & ~w414;
assign w912 = w55 & ~w1103;
assign w913 = (~w368 & ~w215) | (~w368 & w613) | (~w215 & w613);
assign w914 = ~w816 & ~w752;
assign w915 = (w90 & w703) | (w90 & w20) | (w703 & w20);
assign w916 = ~w1131 & ~w170;
assign w917 = ~w419 & ~w226;
assign w918 = (w77 & w789) | (w77 & w101) | (w789 & w101);
assign w919 = w1137 & ~w1118;
assign w920 = (w749 & w762) | (w749 & w613) | (w762 & w613);
assign w921 = ~w235 & w1132;
assign w922 = (w1003 & w168) | (w1003 & ~w769) | (w168 & ~w769);
assign w923 = w1026 & ~w687;
assign w924 = (w658 & w398) | (w658 & w516) | (w398 & w516);
assign w925 = ~w1109 & w673;
assign w926 = w646 & w80;
assign w927 = a63 & b63;
assign w928 = ~w55 & w746;
assign w929 = ~b11 & ~a11;
assign w930 = b32 & a32;
assign w931 = w130 & w53;
assign w932 = (w146 & ~w17) | (w146 & w777) | (~w17 & w777);
assign w933 = (w528 & w229) | (w528 & w697) | (w229 & w697);
assign w934 = ~w1018 & ~w388;
assign w935 = ~w322 & w691;
assign w936 = b45 & a45;
assign w937 = w265 & ~w679;
assign w938 = ~w551 & ~w304;
assign w939 = ~b61 & ~a61;
assign w940 = b22 & a22;
assign w941 = w349 & ~w558;
assign w942 = (~w138 & w921) | (~w138 & w464) | (w921 & w464);
assign w943 = (~w745 & ~w250) | (~w745 & w372) | (~w250 & w372);
assign w944 = a1 & w608;
assign w945 = (w658 & w587) | (w658 & w442) | (w587 & w442);
assign w946 = (~w528 & w704) | (~w528 & w967) | (w704 & w967);
assign w947 = w378 & ~w946;
assign w948 = (~w531 & w665) | (~w531 & w922) | (w665 & w922);
assign w949 = ~w836 & ~w397;
assign w950 = ~w532 & ~w557;
assign w951 = (~w531 & w820) | (~w531 & w1158) | (w820 & w1158);
assign w952 = ~w189 & ~w489;
assign w953 = ~b41 & ~a41;
assign w954 = (~w563 & w1050) | (~w563 & w960) | (w1050 & w960);
assign w955 = w341 & ~w641;
assign w956 = ~w265 & w679;
assign w957 = w324 & w560;
assign w958 = ~w116 & ~w1099;
assign w959 = (~w742 & w609) | (~w742 & w712) | (w609 & w712);
assign w960 = w1086 & ~w497;
assign w961 = (~w220 & ~w1087) | (~w220 & ~w582) | (~w1087 & ~w582);
assign w962 = ~b5 & ~a5;
assign w963 = (w1015 & w545) | (w1015 & w278) | (w545 & w278);
assign w964 = (w676 & w885) | (w676 & w454) | (w885 & w454);
assign w965 = ~w255 & ~w143;
assign w966 = (~w610 & ~w801) | (~w610 & ~w898) | (~w801 & ~w898);
assign w967 = (~w759 & ~w981) | (~w759 & w310) | (~w981 & w310);
assign w968 = ~w872 & ~w664;
assign w969 = (w742 & w370) | (w742 & w391) | (w370 & w391);
assign w970 = w42 & ~w367;
assign w971 = b4 & a4;
assign w972 = w224 & w110;
assign w973 = (~w752 & w1004) | (~w752 & w244) | (w1004 & w244);
assign w974 = w189 & w711;
assign w975 = b9 & a9;
assign w976 = (~w494 & w919) | (~w494 & w280) | (w919 & w280);
assign w977 = (w1101 & w129) | (w1101 & w1035) | (w129 & w1035);
assign w978 = (w83 & w129) | (w83 & ~w844) | (w129 & ~w844);
assign w979 = ~w701 & ~w729;
assign w980 = ~w89 & w483;
assign w981 = ~w255 & ~w759;
assign w982 = (~w25 & w750) | (~w25 & w216) | (w750 & w216);
assign w983 = w358 & ~w824;
assign w984 = ~w269 & ~w962;
assign w985 = ~w1053 & w205;
assign w986 = (~w77 & w867) | (~w77 & w212) | (w867 & w212);
assign w987 = w291 & ~w91;
assign w988 = ~w1134 & w1118;
assign w989 = (w658 & w1102) | (w658 & w808) | (w1102 & w808);
assign w990 = w224 & w86;
assign w991 = ~b20 & ~a20;
assign w992 = ~w554 & w864;
assign w993 = ~b47 & ~a47;
assign w994 = (w658 & w253) | (w658 & w880) | (w253 & w880);
assign w995 = ~w1086 & w497;
assign w996 = w1076 & ~w1008;
assign w997 = ~w506 & w794;
assign w998 = (w658 & w970) | (w658 & w903) | (w970 & w903);
assign w999 = ~w1076 & ~w592;
assign w1000 = w1029 & w718;
assign w1001 = (w518 & w1150) | (w518 & w401) | (w1150 & w401);
assign w1002 = (~w105 & ~w232) | (~w105 & w1009) | (~w232 & w1009);
assign w1003 = w500 & ~w91;
assign w1004 = (w67 & w121) | (w67 & ~w1103) | (w121 & ~w1103);
assign w1005 = ~w51 & ~w343;
assign w1006 = (~w531 & w267) | (~w531 & w181) | (w267 & w181);
assign w1007 = w225 & ~w505;
assign w1008 = ~w309 & w554;
assign w1009 = ~w546 & ~w105;
assign w1010 = w129 & w83;
assign w1011 = (~w385 & ~w199) | (~w385 & w613) | (~w199 & w613);
assign w1012 = (~w854 & w25) | (~w854 & w542) | (w25 & w542);
assign w1013 = (w1101 & w628) | (w1101 & w835) | (w628 & w835);
assign w1014 = ~w1078 & ~w1071;
assign w1015 = ~w85 & w477;
assign w1016 = w437 & ~w199;
assign w1017 = ~w792 & w1046;
assign w1018 = b19 & a19;
assign w1019 = ~w1053 & w1103;
assign w1020 = ~w1029 & ~w718;
assign w1021 = w1094 & w662;
assign w1022 = (w691 & w531) | (w691 & w935) | (w531 & w935);
assign w1023 = (w706 & ~w942) | (w706 & w70) | (~w942 & w70);
assign w1024 = (~w248 & ~w847) | (~w248 & w15) | (~w847 & w15);
assign w1025 = (w170 & w884) | (w170 & w136) | (w884 & w136);
assign w1026 = ~w929 & ~w909;
assign w1027 = (w805 & w573) | (w805 & w755) | (w573 & w755);
assign w1028 = (w77 & w911) | (w77 & w521) | (w911 & w521);
assign w1029 = ~b12 & ~a12;
assign w1030 = w847 & w362;
assign w1031 = w346 & ~w31;
assign w1032 = w79 & w294;
assign w1033 = w349 & ~w490;
assign w1034 = (~w742 & ~w469) | (~w742 & ~w160) | (~w469 & ~w160);
assign w1035 = ~w844 & w1012;
assign w1036 = b13 & a13;
assign w1037 = (w769 & w628) | (w769 & w835) | (w628 & w835);
assign w1038 = w934 & ~w613;
assign w1039 = w1137 & ~w739;
assign w1040 = (w932 & w424) | (w932 & w769) | (w424 & w769);
assign w1041 = ~w957 & ~w824;
assign w1042 = ~w646 & ~w656;
assign w1043 = (~w829 & w282) | (~w829 & w240) | (w282 & w240);
assign w1044 = ~b37 & ~a37;
assign w1045 = (w388 & w1088) | (w388 & w278) | (w1088 & w278);
assign w1046 = (~w455 & w235) | (~w455 & w491) | (w235 & w491);
assign w1047 = (w984 & w1122) | (w984 & w370) | (w1122 & w370);
assign w1048 = (w876 & w596) | (w876 & ~w613) | (w596 & ~w613);
assign w1049 = (w92 & w354) | (w92 & ~w769) | (w354 & ~w769);
assign w1050 = w1086 & w104;
assign w1051 = w566 & w533;
assign w1052 = (w769 & w3) | (w769 & w22) | (w3 & w22);
assign w1053 = ~w816 & w164;
assign w1054 = (w531 & w325) | (w531 & w734) | (w325 & w734);
assign w1055 = (~w531 & w6) | (~w531 & w774) | (w6 & w774);
assign w1056 = ~b19 & ~a19;
assign w1057 = (w518 & w472) | (w518 & w863) | (w472 & w863);
assign w1058 = w287 & ~w720;
assign w1059 = (w77 & w392) | (w77 & w221) | (w392 & w221);
assign w1060 = (~w531 & w383) | (~w531 & w741) | (w383 & w741);
assign w1061 = ~b3 & ~a3;
assign w1062 = ~b21 & ~a21;
assign w1063 = w699 & ~w486;
assign w1064 = ~w115 & w224;
assign w1065 = ~w265 & w462;
assign w1066 = ~w1074 & w285;
assign w1067 = (w77 & w892) | (w77 & w638) | (w892 & w638);
assign w1068 = ~b34 & ~a34;
assign w1069 = (w1118 & w448) | (w1118 & w988) | (w448 & w988);
assign w1070 = w473 & ~w653;
assign w1071 = ~cin & w748;
assign w1072 = ~w5 & ~w256;
assign w1073 = ~w470 & ~w948;
assign w1074 = ~w971 & w1061;
assign w1075 = w222 & ~w347;
assign w1076 = w33 & w864;
assign w1077 = ~w1097 & w632;
assign w1078 = cin & ~w748;
assign w1079 = ~w699 & w486;
assign w1080 = (~w304 & ~w938) | (~w304 & w362) | (~w938 & w362);
assign w1081 = (w779 & w368) | (w779 & w814) | (w368 & w814);
assign w1082 = b29 & a29;
assign w1083 = ~w184 & ~w984;
assign w1084 = (w706 & ~w464) | (w706 & w70) | (~w464 & w70);
assign w1085 = w782 & ~w348;
assign w1086 = ~w624 & ~w929;
assign w1087 = ~w759 & ~w981;
assign w1088 = w1018 & w388;
assign w1089 = ~w744 & ~w667;
assign w1090 = w825 & ~w1042;
assign w1091 = (w909 & w412) | (w909 & w687) | (w412 & w687);
assign w1092 = (~w531 & w407) | (~w531 & w144) | (w407 & w144);
assign w1093 = (w658 & w725) | (w658 & w586) | (w725 & w586);
assign w1094 = w617 & w662;
assign w1095 = w879 & w731;
assign w1096 = w251 & w1005;
assign w1097 = (~w531 & w281) | (~w531 & w166) | (w281 & w166);
assign w1098 = ~w136 & w916;
assign w1099 = ~b43 & ~a43;
assign w1100 = ~b51 & ~a51;
assign w1101 = (w83 & w824) | (w83 & w505) | (w824 & w505);
assign w1102 = (~w592 & w1008) | (~w592 & w999) | (w1008 & w999);
assign w1103 = w1042 & w197;
assign w1104 = (w783 & ~w720) | (w783 & ~w627) | (~w720 & ~w627);
assign w1105 = (w1081 & w574) | (w1081 & ~w613) | (w574 & ~w613);
assign w1106 = b33 & a33;
assign w1107 = (w193 & w528) | (w193 & w648) | (w528 & w648);
assign w1108 = (w645 & w427) | (w645 & w750) | (w427 & w750);
assign w1109 = ~w744 & ~w975;
assign w1110 = w18 & ~w727;
assign w1111 = (w205 & w985) | (w205 & w829) | (w985 & w829);
assign w1112 = ~w304 & ~w938;
assign w1113 = (~w77 & w1048) | (~w77 & w209) | (w1048 & w209);
assign w1114 = w900 & ~w675;
assign w1115 = w597 & w952;
assign w1116 = w184 & w160;
assign w1117 = (w1125 & w1108) | (w1125 & ~w518) | (w1108 & ~w518);
assign w1118 = ~w476 & ~w406;
assign w1119 = (~w77 & w896) | (~w77 & w411) | (w896 & w411);
assign w1120 = ~w597 & ~w489;
assign w1121 = w792 & ~w1046;
assign w1122 = w971 & w984;
assign w1123 = ~w975 & ~w507;
assign w1124 = (w1015 & w545) | (w1015 & w613) | (w545 & w613);
assign w1125 = w427 & w645;
assign w1126 = w289 & w864;
assign w1127 = w759 & ~w143;
assign w1128 = ~b44 & ~a44;
assign w1129 = (w692 & w48) | (w692 & w631) | (w48 & w631);
assign w1130 = (w658 & w152) | (w658 & w443) | (w152 & w443);
assign w1131 = b25 & a25;
assign w1132 = ~w786 & ~w1;
assign w1133 = ~w445 & ~w971;
assign w1134 = ~w778 & ~w275;
assign w1135 = (w621 & w249) | (w621 & ~w898) | (w249 & ~w898);
assign w1136 = (~w531 & w817) | (~w531 & w512) | (w817 & w512);
assign w1137 = ~w953 & ~w520;
assign w1138 = ~w597 & ~w936;
assign w1139 = ~b52 & ~a52;
assign w1140 = w232 & w329;
assign w1141 = w582 & ~w759;
assign w1142 = w307 & w904;
assign w1143 = (w370 & w941) | (w370 & w1033) | (w941 & w1033);
assign w1144 = (~w563 & w108) | (~w563 & w72) | (w108 & w72);
assign w1145 = (w92 & w354) | (w92 & ~w1101) | (w354 & ~w1101);
assign w1146 = (~w658 & w889) | (~w658 & w650) | (w889 & w650);
assign w1147 = ~w24 & ~w507;
assign w1148 = ~w969 & ~w359;
assign w1149 = ~w1140 & ~w733;
assign w1150 = (w637 & w36) | (w637 & w83) | (w36 & w83);
assign w1151 = (~w610 & ~w801) | (~w610 & ~w91) | (~w801 & ~w91);
assign w1152 = ~w742 & w635;
assign w1153 = ~w363 & ~w390;
assign w1154 = (~w85 & w881) | (~w85 & w278) | (w881 & w278);
assign w1155 = (~w453 & ~w672) | (~w453 & w447) | (~w672 & w447);
assign w1156 = b39 & a39;
assign w1157 = w566 & w301;
assign w1158 = (~w846 & w931) | (~w846 & w827) | (w931 & w827);
assign one = 1;
assign s0 = ~w1014;// level 4
assign s1 = w775;// level 6
assign s10 = ~w680;// level 9
assign s11 = ~w147;// level 9
assign s12 = ~w162;// level 9
assign s13 = ~w565;// level 9
assign s14 = w601;// level 9
assign s15 = w823;// level 9
assign s16 = w21;// level 9
assign s17 = w45;// level 9
assign s18 = ~w955;// level 9
assign s19 = ~w242;// level 9
assign s2 = ~w386;// level 6
assign s20 = w1072;// level 9
assign s21 = ~w659;// level 9
assign s22 = ~w404;// level 9
assign s23 = w413;// level 10
assign s24 = ~w721;// level 9
assign s25 = ~w849;// level 10
assign s26 = w949;// level 10
assign s27 = ~w321;// level 10
assign s28 = ~w698;// level 10
assign s29 = w231;// level 10
assign s3 = w826;// level 7
assign s30 = ~w389;// level 10
assign s31 = ~w113;// level 10
assign s32 = w271;// level 10
assign s33 = ~w781;// level 10
assign s34 = ~w858;// level 10
assign s35 = w834;// level 10
assign s36 = ~w394;// level 10
assign s37 = ~w11;// level 10
assign s38 = w293;// level 10
assign s39 = ~w572;// level 10
assign s4 = w1148;// level 7
assign s40 = ~w481;// level 10
assign s41 = w917;// level 10
assign s42 = ~w26;// level 11
assign s43 = ~w1073;// level 10
assign s44 = w502;// level 11
assign s45 = ~w788;// level 11
assign s46 = ~w815;// level 11
assign s47 = w137;// level 11
assign s48 = ~w134;// level 11
assign s49 = ~w319;// level 11
assign s5 = w499;// level 7
assign s50 = w135;// level 11
assign s51 = ~w340;// level 11
assign s52 = ~w58;// level 11
assign s53 = w873;// level 11
assign s54 = ~w799;// level 11
assign s55 = ~w233;// level 11
assign s56 = w452;// level 11
assign s57 = ~w543;// level 11
assign s58 = ~w649;// level 11
assign s59 = w47;// level 11
assign s6 = w97;// level 7
assign s60 = ~w332;// level 11
assign s61 = ~w266;// level 11
assign s62 = ~w4;// level 11
assign s63 = ~w198;// level 11
assign s64 = w899;// level 11
assign s7 = w1153;// level 8
assign s8 = w39;// level 8
assign s9 = w910;// level 8
endmodule
