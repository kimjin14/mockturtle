module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , y0 , y1 , y2 , y3 , y4 , y5 , y6 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 ;
  wire n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 ;
  assign n12 = x4 & x8 ;
  assign n13 = x6 | x7 ;
  assign n14 = x0 & ~x1 ;
  assign n15 = ( x0 & x1 ) | ( x0 & x4 ) | ( x1 & x4 ) ;
  assign n16 = x4 | x8 ;
  assign n17 = x0 & n16 ;
  assign n18 = ( n14 & n15 ) | ( n14 & ~n17 ) | ( n15 & ~n17 ) ;
  assign n19 = n12 | n18 ;
  assign n20 = ( n12 & ~n13 ) | ( n12 & n19 ) | ( ~n13 & n19 ) ;
  assign n21 = ~x5 & n20 ;
  assign n22 = x3 & ~x4 ;
  assign n23 = ( x3 & x4 ) | ( x3 & x7 ) | ( x4 & x7 ) ;
  assign n24 = x1 & ~x2 ;
  assign n25 = x5 & ~x7 ;
  assign n26 = n24 & n25 ;
  assign n27 = x3 & ~n26 ;
  assign n28 = ( n22 & n23 ) | ( n22 & ~n27 ) | ( n23 & ~n27 ) ;
  assign n29 = ~x8 & n28 ;
  assign n30 = ~x4 & x5 ;
  assign n31 = x8 | n29 ;
  assign n32 = ( n29 & n30 ) | ( n29 & n31 ) | ( n30 & n31 ) ;
  assign n33 = n21 | n32 ;
  assign n34 = ~x9 & n33 ;
  assign n35 = ~x5 & x6 ;
  assign n36 = x5 & ~x6 ;
  assign n37 = ~x1 & x2 ;
  assign n38 = x7 | x8 ;
  assign n39 = n37 & ~n38 ;
  assign n40 = x9 | n39 ;
  assign n41 = x4 & ~x8 ;
  assign n42 = ~x3 & n41 ;
  assign n43 = x4 | x7 ;
  assign n44 = ( n24 & n42 ) | ( n24 & ~n43 ) | ( n42 & ~n43 ) ;
  assign n45 = n24 & n44 ;
  assign n46 = ( n36 & n40 ) | ( n36 & n45 ) | ( n40 & n45 ) ;
  assign n47 = n36 & n46 ;
  assign n48 = x9 | n47 ;
  assign n49 = ( n35 & n47 ) | ( n35 & n48 ) | ( n47 & n48 ) ;
  assign n50 = n34 | n49 ;
  assign n51 = ~x10 & n50 ;
  assign n52 = x8 | x9 ;
  assign n53 = ~x2 & x3 ;
  assign n54 = x2 & ~x3 ;
  assign n55 = ( ~n52 & n53 ) | ( ~n52 & n54 ) | ( n53 & n54 ) ;
  assign n56 = ~n52 & n55 ;
  assign n57 = x10 | n56 ;
  assign n58 = ~x7 & n57 ;
  assign n59 = x9 & x10 ;
  assign n60 = x8 & n59 ;
  assign n61 = n58 | n60 ;
  assign n62 = x6 & n61 ;
  assign n63 = ~x6 & x10 ;
  assign n64 = x7 & n63 ;
  assign n65 = n62 | n64 ;
  assign n66 = n51 | n65 ;
  assign n67 = x4 | x9 ;
  assign n68 = x2 | x7 ;
  assign n69 = n67 & n68 ;
  assign n70 = x1 | n69 ;
  assign n71 = ( ~x0 & x2 ) | ( ~x0 & x7 ) | ( x2 & x7 ) ;
  assign n72 = x1 & x2 ;
  assign n73 = ( x0 & x7 ) | ( x0 & ~n72 ) | ( x7 & ~n72 ) ;
  assign n74 = n71 | n73 ;
  assign n75 = x4 & ~n74 ;
  assign n76 = x8 & ~x9 ;
  assign n77 = n75 | n76 ;
  assign n78 = n70 & ~n77 ;
  assign n79 = x6 | n78 ;
  assign n80 = ~x7 & x9 ;
  assign n81 = x3 & x4 ;
  assign n82 = x7 & ~n81 ;
  assign n83 = n80 | n82 ;
  assign n84 = ( ~n52 & n80 ) | ( ~n52 & n83 ) | ( n80 & n83 ) ;
  assign n85 = n79 & ~n84 ;
  assign n86 = ~x4 & n76 ;
  assign n87 = n80 | n86 ;
  assign n88 = ~x6 & n87 ;
  assign n89 = ( x5 & n85 ) | ( x5 & ~n88 ) | ( n85 & ~n88 ) ;
  assign n90 = x7 & ~x9 ;
  assign n91 = n41 & n90 ;
  assign n92 = x4 | n13 ;
  assign n93 = x9 & n92 ;
  assign n94 = ( ~n41 & n92 ) | ( ~n41 & n93 ) | ( n92 & n93 ) ;
  assign n95 = ~n91 & n94 ;
  assign n96 = ( n72 & n91 ) | ( n72 & ~n95 ) | ( n91 & ~n95 ) ;
  assign n97 = x3 & n96 ;
  assign n98 = x4 & n76 ;
  assign n99 = x7 & x9 ;
  assign n100 = n98 | n99 ;
  assign n101 = x6 & n100 ;
  assign n102 = n97 | n101 ;
  assign n103 = ( x5 & n88 ) | ( x5 & n102 ) | ( n88 & n102 ) ;
  assign n104 = n89 & ~n103 ;
  assign n105 = x10 | n104 ;
  assign n106 = x6 & ~x9 ;
  assign n107 = ~x4 & n106 ;
  assign n108 = ~x3 & n36 ;
  assign n109 = n107 | n108 ;
  assign n110 = ~x2 & n109 ;
  assign n111 = ~x1 & n36 ;
  assign n112 = n107 | n111 ;
  assign n113 = ~x3 & n112 ;
  assign n114 = x2 & x3 ;
  assign n115 = x4 & n106 ;
  assign n116 = n114 & n115 ;
  assign n117 = x10 | n116 ;
  assign n118 = n113 | n117 ;
  assign n119 = n110 | n118 ;
  assign n120 = ~x7 & n119 ;
  assign n121 = n63 | n120 ;
  assign n122 = ~x8 & n121 ;
  assign n123 = x6 & x7 ;
  assign n124 = ( x10 & n76 ) | ( x10 & ~n123 ) | ( n76 & ~n123 ) ;
  assign n125 = n123 & n124 ;
  assign n126 = n122 | n125 ;
  assign n127 = n105 & ~n126 ;
  assign n128 = x4 & ~x6 ;
  assign n129 = x0 & ~x3 ;
  assign n130 = n128 & n129 ;
  assign n131 = x3 & n30 ;
  assign n132 = n130 | n131 ;
  assign n133 = x1 & n132 ;
  assign n134 = x0 & x1 ;
  assign n135 = n81 & ~n134 ;
  assign n136 = x5 | x6 ;
  assign n137 = x4 | n136 ;
  assign n138 = ( x5 & ~n135 ) | ( x5 & n137 ) | ( ~n135 & n137 ) ;
  assign n139 = x2 & ~n138 ;
  assign n140 = ( x2 & n133 ) | ( x2 & n139 ) | ( n133 & n139 ) ;
  assign n141 = x2 & n35 ;
  assign n142 = n111 | n141 ;
  assign n143 = x5 & x6 ;
  assign n144 = ~n81 & n143 ;
  assign n145 = n81 | n144 ;
  assign n146 = ( n142 & n144 ) | ( n142 & n145 ) | ( n144 & n145 ) ;
  assign n147 = x3 & ~x6 ;
  assign n148 = ~x2 & n147 ;
  assign n149 = x4 & x5 ;
  assign n150 = ~x3 & n149 ;
  assign n151 = ( x4 & n148 ) | ( x4 & n150 ) | ( n148 & n150 ) ;
  assign n152 = ~x7 & n151 ;
  assign n153 = n146 | n152 ;
  assign n154 = x7 & ~n146 ;
  assign n155 = ( n140 & n153 ) | ( n140 & ~n154 ) | ( n153 & ~n154 ) ;
  assign n156 = ~x6 & x7 ;
  assign n157 = x3 & n156 ;
  assign n158 = x6 & ~x7 ;
  assign n159 = ~x2 & n158 ;
  assign n160 = n157 | n159 ;
  assign n161 = ( ~x5 & n30 ) | ( ~x5 & n123 ) | ( n30 & n123 ) ;
  assign n162 = ( x5 & ~n30 ) | ( x5 & n161 ) | ( ~n30 & n161 ) ;
  assign n163 = ( n160 & n161 ) | ( n160 & n162 ) | ( n161 & n162 ) ;
  assign n164 = x8 | n163 ;
  assign n165 = ( x9 & ~n163 ) | ( x9 & n164 ) | ( ~n163 & n164 ) ;
  assign n166 = ~x9 & n163 ;
  assign n167 = ( n155 & ~n165 ) | ( n155 & n166 ) | ( ~n165 & n166 ) ;
  assign n168 = x5 & x7 ;
  assign n169 = x8 | x10 ;
  assign n170 = ( x10 & ~n168 ) | ( x10 & n169 ) | ( ~n168 & n169 ) ;
  assign n171 = x9 & n170 ;
  assign n172 = ~x8 & x9 ;
  assign n173 = x5 & n172 ;
  assign n174 = x8 & x10 ;
  assign n175 = n123 & n174 ;
  assign n176 = ( n123 & n173 ) | ( n123 & n175 ) | ( n173 & n175 ) ;
  assign n177 = n171 | n176 ;
  assign n178 = x4 & x6 ;
  assign n179 = n25 & n178 ;
  assign n180 = x8 & n156 ;
  assign n181 = ( x8 & n179 ) | ( x8 & n180 ) | ( n179 & n180 ) ;
  assign n182 = x10 | n181 ;
  assign n183 = ( ~x10 & n177 ) | ( ~x10 & n182 ) | ( n177 & n182 ) ;
  assign n184 = x10 & ~n177 ;
  assign n185 = ( n167 & n183 ) | ( n167 & ~n184 ) | ( n183 & ~n184 ) ;
  assign n186 = x9 | x10 ;
  assign n187 = ~x2 & n123 ;
  assign n188 = x5 & n12 ;
  assign n189 = n187 & n188 ;
  assign n190 = x5 | n16 ;
  assign n191 = n13 | n190 ;
  assign n192 = ( n186 & ~n189 ) | ( n186 & n191 ) | ( ~n189 & n191 ) ;
  assign n193 = n186 | n192 ;
  assign n194 = x3 | n193 ;
  assign n195 = x4 | n158 ;
  assign n196 = x7 | n36 ;
  assign n197 = ~x3 & n196 ;
  assign n198 = x7 & ~n143 ;
  assign n199 = ~x9 & n72 ;
  assign n200 = ( x9 & n36 ) | ( x9 & ~n199 ) | ( n36 & ~n199 ) ;
  assign n201 = n198 | n200 ;
  assign n202 = n197 | n201 ;
  assign n203 = n195 & ~n202 ;
  assign n204 = x4 & ~x7 ;
  assign n205 = n143 & n204 ;
  assign n206 = n134 & ~n136 ;
  assign n207 = ( n114 & n205 ) | ( n114 & n206 ) | ( n205 & n206 ) ;
  assign n208 = n114 & n207 ;
  assign n209 = n203 & ~n208 ;
  assign n210 = x8 | n209 ;
  assign n211 = x4 & x7 ;
  assign n212 = x3 & x8 ;
  assign n213 = ( n54 & n143 ) | ( n54 & n212 ) | ( n143 & n212 ) ;
  assign n214 = n143 & n213 ;
  assign n215 = ( x9 & n211 ) | ( x9 & ~n214 ) | ( n211 & ~n214 ) ;
  assign n216 = n211 & ~n215 ;
  assign n217 = ( x9 & n80 ) | ( x9 & ~n143 ) | ( n80 & ~n143 ) ;
  assign n218 = n216 | n217 ;
  assign n219 = n210 & ~n218 ;
  assign n220 = x10 | n219 ;
  assign n221 = x8 & n168 ;
  assign n222 = x6 & n221 ;
  assign n223 = x5 | n38 ;
  assign n224 = ( ~x3 & n134 ) | ( ~x3 & n223 ) | ( n134 & n223 ) ;
  assign n225 = n134 & ~n224 ;
  assign n226 = n222 | n225 ;
  assign n227 = x2 & n226 ;
  assign n228 = x3 & x6 ;
  assign n229 = n221 & n228 ;
  assign n230 = n227 | n229 ;
  assign n231 = x4 & n230 ;
  assign n232 = n114 & n178 ;
  assign n233 = x5 & ~n232 ;
  assign n234 = ( n35 & ~n38 ) | ( n35 & n233 ) | ( ~n38 & n233 ) ;
  assign n235 = ~n38 & n234 ;
  assign n236 = n186 | n235 ;
  assign n237 = n231 | n236 ;
  assign n238 = x2 & n81 ;
  assign n239 = ( n143 & n186 ) | ( n143 & n238 ) | ( n186 & n238 ) ;
  assign n240 = n186 | n239 ;
  assign n241 = n38 | n240 ;
  assign y0 = n66 ;
  assign y1 = n127 ;
  assign y2 = n185 ;
  assign y3 = n194 ;
  assign y4 = n220 ;
  assign y5 = n237 ;
  assign y6 = n241 ;
endmodule
