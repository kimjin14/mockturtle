module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 ;
  wire n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , n3931 , n3932 , n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , n3940 , n3941 , n3942 , n3943 , n3944 , n3945 , n3946 , n3947 , n3948 , n3949 , n3950 , n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , n3970 , n3971 , n3972 , n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , n3980 , n3981 , n3982 , n3983 , n3984 , n3985 , n3986 , n3987 , n3988 , n3989 , n3990 , n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , n4000 , n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , n4009 , n4010 , n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , n4019 , n4020 , n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , n4029 , n4030 , n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , n4039 , n4040 , n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4049 , n4050 , n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , n4059 , n4060 , n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , n4070 , n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , n4079 , n4080 , n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , n4089 , n4090 , n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , n4097 , n4098 , n4099 , n4100 , n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , n4109 , n4110 , n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , n4119 , n4120 , n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , n4129 , n4130 , n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , n4139 , n4140 , n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , n4150 , n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , n4159 , n4160 , n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , n4169 , n4170 , n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , n4179 , n4180 , n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , n4189 , n4190 , n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , n4197 , n4198 , n4199 , n4200 , n4201 , n4202 , n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , n4209 , n4210 , n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , n4217 , n4218 , n4219 , n4220 , n4221 , n4222 , n4223 , n4224 , n4225 , n4226 , n4227 , n4228 , n4229 , n4230 , n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , n4237 , n4238 , n4239 , n4240 , n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , n4247 , n4248 , n4249 , n4250 , n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , n4259 , n4260 , n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , n4269 , n4270 , n4271 , n4272 , n4273 , n4274 , n4275 , n4276 , n4277 , n4278 , n4279 , n4280 , n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , n4289 , n4290 , n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , n4299 , n4300 , n4301 , n4302 , n4303 , n4304 , n4305 , n4306 , n4307 , n4308 , n4309 , n4310 , n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , n4319 , n4320 , n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , n4329 , n4330 , n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , n4340 , n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , n4349 , n4350 , n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , n4360 , n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , n4370 , n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , n4380 , n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , n4390 , n4391 , n4392 , n4393 , n4394 , n4395 , n4396 , n4397 , n4398 , n4399 , n4400 , n4401 , n4402 , n4403 , n4404 , n4405 , n4406 , n4407 , n4408 , n4409 , n4410 , n4411 , n4412 , n4413 , n4414 , n4415 , n4416 , n4417 , n4418 , n4419 , n4420 , n4421 , n4422 , n4423 , n4424 , n4425 , n4426 , n4427 , n4428 , n4429 , n4430 , n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , n4437 , n4438 , n4439 , n4440 , n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , n4449 , n4450 , n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , n4459 , n4460 , n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , n4469 , n4470 , n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , n4479 , n4480 , n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , n4487 , n4488 , n4489 , n4490 , n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , n4497 , n4498 , n4499 , n4500 , n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , n4509 , n4510 , n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , n4519 , n4520 , n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , n4529 , n4530 , n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , n4537 , n4538 , n4539 , n4540 , n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , n4547 , n4548 , n4549 , n4550 , n4551 , n4552 , n4553 , n4554 , n4555 , n4556 , n4557 , n4558 , n4559 , n4560 , n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , n4567 , n4568 , n4569 , n4570 , n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , n4579 , n4580 , n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , n4589 , n4590 , n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , n4597 , n4598 , n4599 , n4600 , n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , n4607 , n4608 , n4609 , n4610 , n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , n4617 , n4618 , n4619 , n4620 , n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , n4627 , n4628 , n4629 , n4630 , n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , n4637 , n4638 , n4639 , n4640 , n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , n4647 , n4648 , n4649 , n4650 , n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , n4657 , n4658 , n4659 , n4660 , n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , n4669 , n4670 , n4671 , n4672 , n4673 , n4674 , n4675 , n4676 , n4677 , n4678 , n4679 , n4680 , n4681 , n4682 , n4683 , n4684 , n4685 , n4686 , n4687 , n4688 , n4689 , n4690 , n4691 , n4692 , n4693 , n4694 , n4695 , n4696 , n4697 , n4698 , n4699 , n4700 , n4701 , n4702 , n4703 , n4704 , n4705 , n4706 , n4707 , n4708 , n4709 , n4710 , n4711 , n4712 , n4713 , n4714 , n4715 , n4716 , n4717 , n4718 , n4719 , n4720 , n4721 , n4722 , n4723 , n4724 , n4725 , n4726 , n4727 , n4728 , n4729 , n4730 , n4731 , n4732 , n4733 , n4734 , n4735 , n4736 , n4737 , n4738 , n4739 , n4740 , n4741 , n4742 , n4743 , n4744 , n4745 , n4746 , n4747 , n4748 , n4749 , n4750 , n4751 , n4752 , n4753 , n4754 , n4755 , n4756 , n4757 , n4758 , n4759 , n4760 , n4761 , n4762 , n4763 , n4764 , n4765 , n4766 , n4767 , n4768 , n4769 , n4770 , n4771 , n4772 , n4773 , n4774 , n4775 , n4776 , n4777 , n4778 , n4779 , n4780 , n4781 , n4782 , n4783 , n4784 , n4785 , n4786 , n4787 , n4788 , n4789 , n4790 , n4791 , n4792 , n4793 , n4794 , n4795 , n4796 , n4797 , n4798 , n4799 , n4800 , n4801 , n4802 , n4803 , n4804 , n4805 , n4806 , n4807 , n4808 , n4809 , n4810 , n4811 , n4812 , n4813 , n4814 , n4815 , n4816 , n4817 , n4818 , n4819 , n4820 , n4821 , n4822 , n4823 , n4824 , n4825 , n4826 , n4827 , n4828 , n4829 , n4830 , n4831 , n4832 , n4833 , n4834 , n4835 , n4836 , n4837 , n4838 , n4839 , n4840 , n4841 , n4842 , n4843 , n4844 , n4845 , n4846 , n4847 , n4848 , n4849 , n4850 , n4851 , n4852 , n4853 , n4854 , n4855 , n4856 , n4857 , n4858 , n4859 , n4860 , n4861 , n4862 , n4863 , n4864 , n4865 , n4866 , n4867 , n4868 , n4869 , n4870 , n4871 , n4872 , n4873 , n4874 , n4875 , n4876 , n4877 , n4878 , n4879 , n4880 , n4881 , n4882 , n4883 , n4884 , n4885 , n4886 , n4887 , n4888 , n4889 , n4890 , n4891 , n4892 , n4893 , n4894 , n4895 , n4896 , n4897 , n4898 , n4899 , n4900 , n4901 , n4902 , n4903 , n4904 , n4905 , n4906 , n4907 , n4908 , n4909 , n4910 , n4911 , n4912 , n4913 , n4914 , n4915 , n4916 , n4917 , n4918 , n4919 , n4920 , n4921 , n4922 , n4923 , n4924 , n4925 , n4926 , n4927 , n4928 , n4929 , n4930 , n4931 , n4932 , n4933 , n4934 , n4935 , n4936 , n4937 , n4938 , n4939 , n4940 , n4941 , n4942 , n4943 , n4944 , n4945 , n4946 , n4947 , n4948 , n4949 , n4950 , n4951 , n4952 , n4953 , n4954 , n4955 , n4956 , n4957 , n4958 , n4959 , n4960 , n4961 , n4962 , n4963 , n4964 , n4965 , n4966 , n4967 , n4968 , n4969 , n4970 , n4971 , n4972 , n4973 , n4974 , n4975 , n4976 , n4977 , n4978 , n4979 , n4980 , n4981 , n4982 , n4983 , n4984 , n4985 , n4986 , n4987 , n4988 , n4989 , n4990 , n4991 , n4992 , n4993 , n4994 , n4995 , n4996 , n4997 , n4998 , n4999 , n5000 , n5001 , n5002 , n5003 , n5004 , n5005 , n5006 , n5007 , n5008 , n5009 , n5010 , n5011 , n5012 , n5013 , n5014 , n5015 , n5016 , n5017 , n5018 , n5019 , n5020 , n5021 , n5022 , n5023 , n5024 , n5025 , n5026 , n5027 , n5028 , n5029 , n5030 , n5031 , n5032 , n5033 , n5034 , n5035 , n5036 , n5037 , n5038 , n5039 , n5040 , n5041 , n5042 , n5043 , n5044 , n5045 , n5046 , n5047 , n5048 , n5049 , n5050 , n5051 , n5052 , n5053 , n5054 , n5055 , n5056 , n5057 , n5058 , n5059 , n5060 , n5061 , n5062 , n5063 , n5064 , n5065 , n5066 , n5067 , n5068 , n5069 , n5070 , n5071 , n5072 , n5073 , n5074 , n5075 , n5076 , n5077 , n5078 , n5079 , n5080 , n5081 , n5082 , n5083 , n5084 , n5085 , n5086 , n5087 , n5088 , n5089 , n5090 , n5091 , n5092 , n5093 , n5094 , n5095 , n5096 , n5097 , n5098 , n5099 , n5100 , n5101 , n5102 , n5103 , n5104 , n5105 , n5106 , n5107 , n5108 , n5109 , n5110 , n5111 , n5112 , n5113 , n5114 , n5115 , n5116 , n5117 , n5118 , n5119 , n5120 , n5121 , n5122 , n5123 , n5124 , n5125 , n5126 , n5127 , n5128 , n5129 , n5130 , n5131 , n5132 , n5133 , n5134 , n5135 , n5136 , n5137 , n5138 , n5139 , n5140 , n5141 , n5142 , n5143 , n5144 , n5145 , n5146 , n5147 , n5148 , n5149 , n5150 , n5151 , n5152 , n5153 , n5154 , n5155 , n5156 , n5157 , n5158 , n5159 , n5160 , n5161 , n5162 , n5163 , n5164 , n5165 , n5166 , n5167 , n5168 , n5169 , n5170 , n5171 , n5172 , n5173 , n5174 , n5175 , n5176 , n5177 , n5178 , n5179 , n5180 , n5181 , n5182 , n5183 , n5184 , n5185 , n5186 , n5187 , n5188 , n5189 , n5190 , n5191 , n5192 , n5193 , n5194 , n5195 , n5196 , n5197 , n5198 , n5199 , n5200 , n5201 , n5202 , n5203 , n5204 , n5205 , n5206 , n5207 , n5208 , n5209 , n5210 , n5211 , n5212 , n5213 , n5214 , n5215 , n5216 , n5217 , n5218 , n5219 , n5220 , n5221 , n5222 , n5223 , n5224 , n5225 , n5226 , n5227 , n5228 , n5229 , n5230 , n5231 , n5232 , n5233 , n5234 , n5235 , n5236 , n5237 , n5238 , n5239 , n5240 , n5241 , n5242 , n5243 , n5244 , n5245 , n5246 , n5247 , n5248 , n5249 , n5250 , n5251 , n5252 , n5253 , n5254 , n5255 , n5256 , n5257 , n5258 , n5259 , n5260 , n5261 , n5262 , n5263 , n5264 , n5265 , n5266 , n5267 , n5268 , n5269 , n5270 , n5271 , n5272 , n5273 , n5274 , n5275 , n5276 , n5277 , n5278 , n5279 , n5280 , n5281 , n5282 , n5283 , n5284 , n5285 , n5286 , n5287 , n5288 , n5289 , n5290 , n5291 , n5292 , n5293 , n5294 , n5295 , n5296 , n5297 , n5298 , n5299 , n5300 , n5301 , n5302 , n5303 , n5304 , n5305 , n5306 , n5307 , n5308 , n5309 , n5310 , n5311 , n5312 , n5313 , n5314 , n5315 , n5316 , n5317 , n5318 , n5319 , n5320 , n5321 , n5322 , n5323 , n5324 , n5325 , n5326 , n5327 , n5328 , n5329 , n5330 , n5331 , n5332 , n5333 , n5334 , n5335 , n5336 , n5337 , n5338 , n5339 , n5340 , n5341 , n5342 , n5343 , n5344 , n5345 , n5346 , n5347 , n5348 , n5349 , n5350 , n5351 , n5352 , n5353 , n5354 , n5355 , n5356 , n5357 , n5358 , n5359 , n5360 , n5361 , n5362 , n5363 , n5364 , n5365 , n5366 , n5367 , n5368 , n5369 , n5370 , n5371 , n5372 , n5373 , n5374 , n5375 , n5376 , n5377 , n5378 , n5379 , n5380 , n5381 , n5382 , n5383 , n5384 , n5385 , n5386 , n5387 , n5388 , n5389 , n5390 , n5391 , n5392 , n5393 , n5394 , n5395 , n5396 , n5397 , n5398 , n5399 , n5400 , n5401 , n5402 , n5403 , n5404 , n5405 , n5406 , n5407 , n5408 , n5409 , n5410 , n5411 , n5412 , n5413 , n5414 , n5415 , n5416 , n5417 , n5418 , n5419 , n5420 , n5421 , n5422 , n5423 , n5424 , n5425 , n5426 , n5427 , n5428 , n5429 , n5430 , n5431 , n5432 , n5433 , n5434 , n5435 , n5436 , n5437 , n5438 , n5439 , n5440 , n5441 , n5442 , n5443 , n5444 , n5445 , n5446 , n5447 , n5448 , n5449 , n5450 , n5451 , n5452 , n5453 , n5454 , n5455 , n5456 , n5457 , n5458 , n5459 , n5460 , n5461 , n5462 , n5463 , n5464 , n5465 , n5466 , n5467 , n5468 , n5469 , n5470 , n5471 , n5472 , n5473 , n5474 , n5475 , n5476 , n5477 , n5478 , n5479 , n5480 , n5481 , n5482 , n5483 , n5484 , n5485 , n5486 , n5487 , n5488 , n5489 , n5490 , n5491 , n5492 , n5493 , n5494 , n5495 , n5496 , n5497 , n5498 , n5499 , n5500 , n5501 , n5502 , n5503 , n5504 , n5505 , n5506 , n5507 , n5508 , n5509 , n5510 , n5511 , n5512 , n5513 , n5514 , n5515 , n5516 , n5517 , n5518 , n5519 , n5520 , n5521 , n5522 , n5523 , n5524 , n5525 , n5526 , n5527 , n5528 , n5529 , n5530 , n5531 , n5532 , n5533 , n5534 , n5535 , n5536 , n5537 , n5538 , n5539 , n5540 , n5541 , n5542 , n5543 , n5544 , n5545 , n5546 , n5547 , n5548 , n5549 , n5550 , n5551 , n5552 , n5553 , n5554 , n5555 , n5556 , n5557 , n5558 , n5559 , n5560 , n5561 , n5562 , n5563 , n5564 , n5565 , n5566 , n5567 , n5568 , n5569 , n5570 , n5571 , n5572 , n5573 , n5574 , n5575 , n5576 , n5577 , n5578 , n5579 , n5580 , n5581 , n5582 , n5583 , n5584 , n5585 , n5586 , n5587 , n5588 , n5589 , n5590 , n5591 , n5592 , n5593 , n5594 , n5595 , n5596 , n5597 , n5598 , n5599 , n5600 , n5601 , n5602 , n5603 , n5604 , n5605 , n5606 , n5607 , n5608 , n5609 , n5610 , n5611 , n5612 , n5613 , n5614 , n5615 , n5616 , n5617 , n5618 , n5619 , n5620 , n5621 , n5622 , n5623 , n5624 , n5625 , n5626 , n5627 , n5628 , n5629 , n5630 , n5631 , n5632 , n5633 , n5634 , n5635 , n5636 , n5637 , n5638 , n5639 , n5640 , n5641 , n5642 , n5643 , n5644 , n5645 , n5646 , n5647 , n5648 , n5649 , n5650 , n5651 , n5652 , n5653 , n5654 , n5655 , n5656 , n5657 , n5658 , n5659 , n5660 , n5661 , n5662 , n5663 , n5664 , n5665 , n5666 , n5667 , n5668 , n5669 , n5670 , n5671 , n5672 , n5673 , n5674 , n5675 , n5676 , n5677 , n5678 , n5679 , n5680 , n5681 , n5682 , n5683 , n5684 , n5685 , n5686 , n5687 , n5688 , n5689 , n5690 , n5691 , n5692 , n5693 , n5694 , n5695 , n5696 , n5697 , n5698 , n5699 , n5700 , n5701 , n5702 , n5703 , n5704 , n5705 , n5706 , n5707 , n5708 , n5709 , n5710 , n5711 , n5712 , n5713 , n5714 , n5715 , n5716 , n5717 , n5718 , n5719 , n5720 , n5721 , n5722 , n5723 , n5724 , n5725 , n5726 , n5727 , n5728 , n5729 , n5730 , n5731 , n5732 , n5733 , n5734 , n5735 , n5736 , n5737 , n5738 , n5739 , n5740 , n5741 , n5742 , n5743 , n5744 , n5745 , n5746 , n5747 , n5748 , n5749 , n5750 , n5751 , n5752 , n5753 , n5754 , n5755 , n5756 , n5757 , n5758 , n5759 , n5760 , n5761 , n5762 , n5763 , n5764 , n5765 , n5766 , n5767 , n5768 , n5769 , n5770 , n5771 , n5772 , n5773 , n5774 , n5775 , n5776 , n5777 , n5778 , n5779 , n5780 , n5781 , n5782 , n5783 , n5784 , n5785 , n5786 , n5787 , n5788 , n5789 , n5790 , n5791 , n5792 , n5793 , n5794 , n5795 , n5796 , n5797 , n5798 , n5799 , n5800 , n5801 , n5802 , n5803 , n5804 , n5805 , n5806 , n5807 , n5808 , n5809 , n5810 , n5811 , n5812 , n5813 , n5814 , n5815 , n5816 , n5817 , n5818 , n5819 , n5820 , n5821 , n5822 , n5823 , n5824 , n5825 , n5826 , n5827 , n5828 , n5829 , n5830 , n5831 , n5832 , n5833 , n5834 , n5835 , n5836 , n5837 , n5838 , n5839 , n5840 , n5841 , n5842 , n5843 , n5844 , n5845 , n5846 , n5847 , n5848 , n5849 , n5850 , n5851 , n5852 , n5853 , n5854 , n5855 , n5856 , n5857 , n5858 , n5859 , n5860 , n5861 , n5862 , n5863 , n5864 , n5865 , n5866 , n5867 , n5868 , n5869 , n5870 , n5871 , n5872 , n5873 , n5874 , n5875 , n5876 , n5877 , n5878 , n5879 , n5880 , n5881 , n5882 , n5883 , n5884 , n5885 , n5886 , n5887 , n5888 , n5889 , n5890 , n5891 , n5892 , n5893 , n5894 , n5895 , n5896 , n5897 , n5898 , n5899 , n5900 , n5901 , n5902 , n5903 , n5904 , n5905 , n5906 , n5907 , n5908 , n5909 , n5910 , n5911 , n5912 , n5913 , n5914 , n5915 , n5916 , n5917 , n5918 , n5919 , n5920 , n5921 , n5922 , n5923 , n5924 , n5925 , n5926 , n5927 , n5928 , n5929 , n5930 , n5931 , n5932 , n5933 , n5934 , n5935 , n5936 , n5937 , n5938 , n5939 , n5940 , n5941 , n5942 , n5943 , n5944 , n5945 , n5946 , n5947 , n5948 , n5949 , n5950 , n5951 , n5952 , n5953 , n5954 , n5955 , n5956 , n5957 , n5958 , n5959 , n5960 , n5961 , n5962 , n5963 , n5964 , n5965 , n5966 , n5967 , n5968 , n5969 , n5970 , n5971 , n5972 , n5973 , n5974 , n5975 , n5976 , n5977 , n5978 , n5979 , n5980 , n5981 , n5982 , n5983 , n5984 , n5985 , n5986 , n5987 , n5988 , n5989 , n5990 , n5991 , n5992 , n5993 , n5994 , n5995 , n5996 , n5997 , n5998 , n5999 , n6000 , n6001 , n6002 , n6003 , n6004 , n6005 , n6006 , n6007 , n6008 , n6009 , n6010 , n6011 , n6012 , n6013 , n6014 , n6015 , n6016 , n6017 , n6018 , n6019 , n6020 , n6021 , n6022 , n6023 , n6024 , n6025 , n6026 , n6027 , n6028 , n6029 , n6030 , n6031 , n6032 , n6033 , n6034 , n6035 , n6036 , n6037 , n6038 , n6039 , n6040 , n6041 , n6042 , n6043 , n6044 , n6045 , n6046 , n6047 , n6048 , n6049 , n6050 , n6051 , n6052 , n6053 , n6054 , n6055 , n6056 , n6057 , n6058 , n6059 , n6060 , n6061 , n6062 , n6063 , n6064 , n6065 , n6066 , n6067 , n6068 , n6069 , n6070 , n6071 , n6072 , n6073 , n6074 , n6075 , n6076 , n6077 , n6078 , n6079 , n6080 , n6081 , n6082 , n6083 , n6084 , n6085 , n6086 , n6087 , n6088 , n6089 , n6090 , n6091 , n6092 , n6093 , n6094 , n6095 , n6096 , n6097 , n6098 , n6099 , n6100 , n6101 , n6102 , n6103 , n6104 , n6105 , n6106 , n6107 , n6108 , n6109 , n6110 , n6111 , n6112 , n6113 , n6114 , n6115 , n6116 , n6117 , n6118 , n6119 , n6120 , n6121 , n6122 , n6123 , n6124 , n6125 , n6126 , n6127 , n6128 , n6129 , n6130 , n6131 , n6132 , n6133 , n6134 , n6135 , n6136 , n6137 , n6138 , n6139 , n6140 , n6141 , n6142 , n6143 , n6144 , n6145 , n6146 , n6147 , n6148 , n6149 , n6150 , n6151 , n6152 , n6153 , n6154 , n6155 , n6156 , n6157 , n6158 , n6159 , n6160 , n6161 , n6162 , n6163 , n6164 , n6165 , n6166 , n6167 , n6168 , n6169 , n6170 , n6171 , n6172 , n6173 , n6174 , n6175 , n6176 , n6177 , n6178 , n6179 , n6180 , n6181 , n6182 , n6183 , n6184 , n6185 , n6186 , n6187 , n6188 , n6189 , n6190 , n6191 , n6192 , n6193 , n6194 , n6195 , n6196 , n6197 , n6198 , n6199 , n6200 , n6201 , n6202 , n6203 , n6204 , n6205 , n6206 , n6207 , n6208 , n6209 , n6210 , n6211 , n6212 , n6213 , n6214 , n6215 , n6216 , n6217 , n6218 , n6219 , n6220 , n6221 , n6222 , n6223 , n6224 , n6225 , n6226 , n6227 , n6228 , n6229 , n6230 , n6231 , n6232 , n6233 , n6234 , n6235 , n6236 , n6237 , n6238 , n6239 , n6240 , n6241 , n6242 , n6243 , n6244 , n6245 , n6246 , n6247 , n6248 , n6249 , n6250 , n6251 , n6252 , n6253 , n6254 , n6255 , n6256 , n6257 , n6258 , n6259 , n6260 , n6261 , n6262 , n6263 , n6264 , n6265 , n6266 , n6267 , n6268 , n6269 , n6270 , n6271 , n6272 , n6273 , n6274 , n6275 , n6276 , n6277 , n6278 , n6279 , n6280 , n6281 , n6282 , n6283 , n6284 , n6285 , n6286 , n6287 , n6288 , n6289 , n6290 , n6291 , n6292 , n6293 , n6294 , n6295 , n6296 , n6297 , n6298 , n6299 , n6300 , n6301 , n6302 , n6303 , n6304 , n6305 , n6306 , n6307 , n6308 , n6309 , n6310 , n6311 , n6312 , n6313 , n6314 , n6315 , n6316 , n6317 , n6318 , n6319 , n6320 , n6321 , n6322 , n6323 , n6324 , n6325 , n6326 , n6327 , n6328 , n6329 , n6330 , n6331 , n6332 , n6333 , n6334 , n6335 , n6336 , n6337 , n6338 , n6339 , n6340 , n6341 , n6342 , n6343 , n6344 , n6345 , n6346 , n6347 , n6348 , n6349 , n6350 , n6351 , n6352 , n6353 , n6354 , n6355 , n6356 , n6357 , n6358 , n6359 , n6360 , n6361 , n6362 , n6363 , n6364 , n6365 , n6366 , n6367 , n6368 , n6369 , n6370 , n6371 , n6372 , n6373 , n6374 , n6375 , n6376 , n6377 , n6378 , n6379 , n6380 , n6381 , n6382 , n6383 , n6384 , n6385 , n6386 , n6387 , n6388 , n6389 , n6390 , n6391 , n6392 , n6393 , n6394 , n6395 , n6396 , n6397 , n6398 , n6399 , n6400 , n6401 , n6402 , n6403 , n6404 , n6405 , n6406 , n6407 , n6408 , n6409 , n6410 , n6411 , n6412 , n6413 , n6414 , n6415 , n6416 , n6417 , n6418 , n6419 , n6420 , n6421 , n6422 , n6423 , n6424 , n6425 , n6426 , n6427 , n6428 , n6429 , n6430 , n6431 , n6432 , n6433 , n6434 , n6435 , n6436 , n6437 , n6438 , n6439 , n6440 , n6441 , n6442 , n6443 , n6444 , n6445 , n6446 , n6447 , n6448 , n6449 , n6450 , n6451 , n6452 , n6453 , n6454 , n6455 , n6456 , n6457 , n6458 , n6459 , n6460 , n6461 , n6462 , n6463 , n6464 , n6465 , n6466 , n6467 , n6468 , n6469 , n6470 , n6471 , n6472 , n6473 , n6474 , n6475 , n6476 , n6477 , n6478 , n6479 , n6480 , n6481 , n6482 , n6483 , n6484 , n6485 , n6486 , n6487 , n6488 , n6489 , n6490 , n6491 , n6492 , n6493 , n6494 , n6495 , n6496 , n6497 , n6498 , n6499 , n6500 , n6501 , n6502 , n6503 , n6504 , n6505 , n6506 , n6507 , n6508 , n6509 , n6510 , n6511 , n6512 , n6513 , n6514 , n6515 , n6516 , n6517 , n6518 , n6519 , n6520 , n6521 , n6522 , n6523 , n6524 , n6525 , n6526 , n6527 , n6528 , n6529 , n6530 , n6531 , n6532 , n6533 , n6534 , n6535 , n6536 , n6537 , n6538 , n6539 , n6540 , n6541 , n6542 , n6543 , n6544 , n6545 , n6546 , n6547 , n6548 , n6549 , n6550 , n6551 , n6552 , n6553 , n6554 , n6555 , n6556 , n6557 , n6558 , n6559 , n6560 , n6561 , n6562 , n6563 , n6564 , n6565 , n6566 , n6567 , n6568 , n6569 , n6570 , n6571 , n6572 , n6573 , n6574 , n6575 , n6576 , n6577 , n6578 , n6579 , n6580 , n6581 , n6582 , n6583 , n6584 , n6585 , n6586 , n6587 , n6588 , n6589 , n6590 , n6591 , n6592 , n6593 , n6594 , n6595 , n6596 , n6597 , n6598 , n6599 , n6600 , n6601 , n6602 , n6603 , n6604 , n6605 , n6606 , n6607 , n6608 , n6609 , n6610 , n6611 , n6612 , n6613 , n6614 , n6615 , n6616 , n6617 , n6618 , n6619 , n6620 , n6621 , n6622 , n6623 , n6624 , n6625 , n6626 , n6627 , n6628 , n6629 , n6630 , n6631 , n6632 , n6633 , n6634 , n6635 , n6636 , n6637 , n6638 , n6639 , n6640 , n6641 , n6642 , n6643 , n6644 , n6645 , n6646 , n6647 , n6648 , n6649 , n6650 , n6651 , n6652 , n6653 , n6654 , n6655 , n6656 , n6657 , n6658 , n6659 , n6660 , n6661 , n6662 , n6663 , n6664 , n6665 , n6666 , n6667 , n6668 , n6669 , n6670 , n6671 , n6672 , n6673 , n6674 , n6675 , n6676 , n6677 , n6678 , n6679 , n6680 , n6681 , n6682 , n6683 , n6684 , n6685 , n6686 , n6687 , n6688 , n6689 , n6690 , n6691 , n6692 , n6693 , n6694 , n6695 , n6696 , n6697 , n6698 , n6699 , n6700 , n6701 , n6702 , n6703 , n6704 , n6705 , n6706 , n6707 , n6708 , n6709 , n6710 , n6711 , n6712 , n6713 , n6714 , n6715 , n6716 , n6717 , n6718 , n6719 , n6720 , n6721 , n6722 , n6723 , n6724 , n6725 , n6726 , n6727 , n6728 , n6729 , n6730 , n6731 , n6732 , n6733 , n6734 , n6735 , n6736 , n6737 , n6738 , n6739 , n6740 , n6741 , n6742 , n6743 , n6744 , n6745 , n6746 , n6747 , n6748 , n6749 , n6750 , n6751 , n6752 , n6753 , n6754 , n6755 , n6756 , n6757 , n6758 , n6759 , n6760 , n6761 , n6762 , n6763 , n6764 , n6765 , n6766 , n6767 , n6768 , n6769 , n6770 , n6771 , n6772 , n6773 , n6774 , n6775 , n6776 , n6777 , n6778 , n6779 , n6780 , n6781 , n6782 , n6783 , n6784 , n6785 , n6786 , n6787 , n6788 , n6789 , n6790 , n6791 , n6792 , n6793 , n6794 , n6795 , n6796 , n6797 , n6798 , n6799 , n6800 , n6801 , n6802 , n6803 , n6804 , n6805 , n6806 , n6807 , n6808 , n6809 , n6810 , n6811 , n6812 , n6813 , n6814 , n6815 , n6816 , n6817 , n6818 , n6819 , n6820 , n6821 , n6822 , n6823 , n6824 , n6825 , n6826 , n6827 , n6828 , n6829 , n6830 , n6831 , n6832 , n6833 , n6834 , n6835 , n6836 , n6837 , n6838 , n6839 , n6840 , n6841 , n6842 , n6843 , n6844 , n6845 , n6846 , n6847 , n6848 , n6849 , n6850 , n6851 , n6852 , n6853 , n6854 , n6855 , n6856 , n6857 , n6858 , n6859 , n6860 , n6861 , n6862 , n6863 , n6864 , n6865 , n6866 , n6867 , n6868 , n6869 , n6870 , n6871 , n6872 , n6873 , n6874 , n6875 , n6876 , n6877 , n6878 , n6879 , n6880 , n6881 , n6882 , n6883 , n6884 , n6885 , n6886 , n6887 , n6888 , n6889 , n6890 , n6891 , n6892 , n6893 , n6894 , n6895 , n6896 , n6897 , n6898 , n6899 , n6900 , n6901 , n6902 , n6903 , n6904 , n6905 , n6906 , n6907 , n6908 , n6909 , n6910 , n6911 , n6912 , n6913 , n6914 , n6915 , n6916 , n6917 , n6918 , n6919 , n6920 , n6921 , n6922 , n6923 , n6924 , n6925 , n6926 , n6927 , n6928 , n6929 , n6930 , n6931 , n6932 , n6933 , n6934 , n6935 , n6936 , n6937 , n6938 , n6939 , n6940 , n6941 , n6942 , n6943 , n6944 , n6945 , n6946 , n6947 , n6948 , n6949 , n6950 , n6951 , n6952 , n6953 , n6954 , n6955 , n6956 , n6957 , n6958 , n6959 , n6960 , n6961 , n6962 , n6963 , n6964 , n6965 , n6966 , n6967 , n6968 , n6969 , n6970 , n6971 , n6972 , n6973 , n6974 , n6975 , n6976 , n6977 , n6978 , n6979 , n6980 , n6981 , n6982 , n6983 , n6984 , n6985 , n6986 , n6987 , n6988 , n6989 , n6990 , n6991 , n6992 , n6993 , n6994 , n6995 , n6996 , n6997 , n6998 , n6999 , n7000 , n7001 , n7002 , n7003 , n7004 , n7005 , n7006 , n7007 , n7008 , n7009 , n7010 , n7011 , n7012 , n7013 , n7014 , n7015 , n7016 , n7017 , n7018 , n7019 , n7020 , n7021 , n7022 , n7023 , n7024 , n7025 , n7026 , n7027 , n7028 , n7029 , n7030 , n7031 , n7032 , n7033 , n7034 , n7035 , n7036 , n7037 , n7038 , n7039 , n7040 , n7041 , n7042 , n7043 , n7044 , n7045 , n7046 , n7047 , n7048 , n7049 , n7050 , n7051 , n7052 , n7053 , n7054 , n7055 , n7056 , n7057 , n7058 , n7059 , n7060 , n7061 , n7062 , n7063 , n7064 , n7065 , n7066 , n7067 , n7068 , n7069 , n7070 , n7071 , n7072 , n7073 , n7074 , n7075 , n7076 , n7077 , n7078 , n7079 , n7080 , n7081 , n7082 , n7083 , n7084 , n7085 , n7086 , n7087 , n7088 , n7089 , n7090 , n7091 , n7092 , n7093 , n7094 , n7095 , n7096 , n7097 , n7098 , n7099 , n7100 , n7101 , n7102 , n7103 , n7104 , n7105 , n7106 , n7107 , n7108 , n7109 , n7110 , n7111 , n7112 , n7113 , n7114 , n7115 , n7116 , n7117 , n7118 , n7119 , n7120 , n7121 , n7122 , n7123 , n7124 , n7125 , n7126 , n7127 , n7128 , n7129 , n7130 , n7131 , n7132 , n7133 , n7134 , n7135 , n7136 , n7137 , n7138 , n7139 , n7140 , n7141 , n7142 , n7143 , n7144 , n7145 , n7146 , n7147 , n7148 , n7149 , n7150 , n7151 , n7152 , n7153 , n7154 , n7155 , n7156 , n7157 , n7158 , n7159 , n7160 , n7161 , n7162 , n7163 , n7164 , n7165 , n7166 , n7167 , n7168 , n7169 , n7170 , n7171 , n7172 , n7173 , n7174 , n7175 , n7176 , n7177 , n7178 , n7179 , n7180 , n7181 , n7182 , n7183 , n7184 , n7185 , n7186 , n7187 , n7188 , n7189 , n7190 , n7191 , n7192 , n7193 , n7194 , n7195 , n7196 , n7197 , n7198 , n7199 , n7200 , n7201 , n7202 , n7203 , n7204 , n7205 , n7206 , n7207 , n7208 , n7209 , n7210 , n7211 , n7212 , n7213 , n7214 , n7215 , n7216 , n7217 , n7218 , n7219 , n7220 , n7221 , n7222 , n7223 , n7224 , n7225 , n7226 , n7227 , n7228 , n7229 , n7230 , n7231 , n7232 , n7233 , n7234 , n7235 , n7236 , n7237 , n7238 , n7239 , n7240 , n7241 , n7242 , n7243 , n7244 , n7245 , n7246 , n7247 , n7248 , n7249 , n7250 , n7251 , n7252 , n7253 , n7254 , n7255 , n7256 , n7257 , n7258 , n7259 , n7260 , n7261 , n7262 , n7263 , n7264 , n7265 , n7266 , n7267 , n7268 , n7269 , n7270 , n7271 , n7272 , n7273 , n7274 , n7275 , n7276 , n7277 , n7278 , n7279 , n7280 , n7281 , n7282 , n7283 , n7284 , n7285 , n7286 , n7287 , n7288 , n7289 , n7290 , n7291 , n7292 , n7293 , n7294 , n7295 , n7296 , n7297 , n7298 , n7299 , n7300 , n7301 , n7302 , n7303 , n7304 , n7305 , n7306 , n7307 , n7308 , n7309 , n7310 , n7311 , n7312 , n7313 , n7314 , n7315 , n7316 , n7317 , n7318 , n7319 , n7320 , n7321 , n7322 , n7323 , n7324 , n7325 , n7326 , n7327 , n7328 , n7329 , n7330 , n7331 , n7332 , n7333 , n7334 , n7335 , n7336 , n7337 , n7338 , n7339 , n7340 , n7341 , n7342 , n7343 , n7344 , n7345 , n7346 , n7347 , n7348 , n7349 , n7350 , n7351 , n7352 , n7353 , n7354 , n7355 , n7356 , n7357 , n7358 , n7359 , n7360 , n7361 , n7362 , n7363 , n7364 , n7365 , n7366 , n7367 , n7368 , n7369 , n7370 , n7371 , n7372 , n7373 , n7374 , n7375 , n7376 , n7377 , n7378 , n7379 , n7380 , n7381 , n7382 , n7383 , n7384 , n7385 , n7386 , n7387 , n7388 , n7389 , n7390 , n7391 , n7392 , n7393 , n7394 , n7395 , n7396 , n7397 , n7398 , n7399 , n7400 , n7401 , n7402 , n7403 , n7404 , n7405 , n7406 , n7407 , n7408 , n7409 , n7410 , n7411 , n7412 , n7413 , n7414 , n7415 , n7416 , n7417 , n7418 , n7419 , n7420 , n7421 , n7422 , n7423 , n7424 , n7425 , n7426 , n7427 , n7428 , n7429 , n7430 , n7431 , n7432 , n7433 , n7434 , n7435 , n7436 , n7437 , n7438 , n7439 , n7440 , n7441 , n7442 , n7443 , n7444 , n7445 , n7446 , n7447 , n7448 , n7449 , n7450 , n7451 , n7452 , n7453 , n7454 , n7455 , n7456 , n7457 , n7458 , n7459 , n7460 , n7461 , n7462 , n7463 , n7464 , n7465 , n7466 , n7467 , n7468 , n7469 , n7470 , n7471 , n7472 , n7473 , n7474 , n7475 , n7476 , n7477 , n7478 , n7479 , n7480 , n7481 , n7482 , n7483 , n7484 , n7485 , n7486 , n7487 , n7488 , n7489 , n7490 , n7491 , n7492 , n7493 , n7494 , n7495 , n7496 , n7497 , n7498 , n7499 , n7500 , n7501 , n7502 , n7503 , n7504 , n7505 , n7506 , n7507 , n7508 , n7509 , n7510 , n7511 , n7512 , n7513 , n7514 , n7515 , n7516 , n7517 , n7518 , n7519 , n7520 , n7521 , n7522 , n7523 , n7524 , n7525 , n7526 , n7527 , n7528 , n7529 , n7530 , n7531 , n7532 , n7533 , n7534 , n7535 , n7536 , n7537 , n7538 , n7539 , n7540 , n7541 , n7542 , n7543 , n7544 , n7545 , n7546 , n7547 , n7548 , n7549 , n7550 , n7551 , n7552 , n7553 , n7554 , n7555 , n7556 , n7557 , n7558 , n7559 , n7560 , n7561 , n7562 , n7563 , n7564 , n7565 , n7566 , n7567 , n7568 , n7569 , n7570 , n7571 , n7572 , n7573 , n7574 , n7575 , n7576 , n7577 , n7578 , n7579 , n7580 , n7581 , n7582 , n7583 , n7584 , n7585 , n7586 , n7587 , n7588 , n7589 , n7590 , n7591 , n7592 , n7593 , n7594 , n7595 , n7596 , n7597 , n7598 , n7599 , n7600 , n7601 , n7602 , n7603 , n7604 , n7605 , n7606 , n7607 , n7608 , n7609 , n7610 , n7611 , n7612 , n7613 , n7614 , n7615 , n7616 , n7617 , n7618 , n7619 , n7620 , n7621 , n7622 , n7623 , n7624 , n7625 , n7626 , n7627 , n7628 , n7629 , n7630 , n7631 , n7632 , n7633 , n7634 , n7635 , n7636 , n7637 , n7638 , n7639 , n7640 , n7641 , n7642 , n7643 , n7644 , n7645 , n7646 , n7647 , n7648 , n7649 , n7650 , n7651 , n7652 , n7653 , n7654 , n7655 , n7656 , n7657 , n7658 , n7659 , n7660 , n7661 , n7662 , n7663 , n7664 , n7665 , n7666 , n7667 , n7668 , n7669 , n7670 , n7671 , n7672 , n7673 , n7674 , n7675 , n7676 , n7677 , n7678 , n7679 , n7680 , n7681 , n7682 , n7683 , n7684 , n7685 , n7686 , n7687 , n7688 , n7689 , n7690 , n7691 , n7692 , n7693 , n7694 , n7695 , n7696 , n7697 , n7698 , n7699 , n7700 , n7701 , n7702 , n7703 , n7704 , n7705 , n7706 , n7707 , n7708 , n7709 , n7710 , n7711 , n7712 , n7713 , n7714 , n7715 , n7716 , n7717 , n7718 , n7719 , n7720 , n7721 , n7722 , n7723 , n7724 , n7725 , n7726 , n7727 , n7728 , n7729 , n7730 , n7731 , n7732 , n7733 , n7734 , n7735 , n7736 , n7737 , n7738 , n7739 , n7740 , n7741 , n7742 , n7743 , n7744 , n7745 , n7746 , n7747 , n7748 , n7749 , n7750 , n7751 , n7752 , n7753 , n7754 , n7755 , n7756 , n7757 , n7758 , n7759 , n7760 , n7761 , n7762 , n7763 , n7764 , n7765 , n7766 , n7767 , n7768 , n7769 , n7770 , n7771 , n7772 , n7773 , n7774 , n7775 , n7776 , n7777 , n7778 , n7779 , n7780 , n7781 , n7782 , n7783 , n7784 , n7785 , n7786 , n7787 , n7788 , n7789 , n7790 , n7791 , n7792 , n7793 , n7794 , n7795 , n7796 , n7797 , n7798 , n7799 , n7800 , n7801 , n7802 , n7803 , n7804 , n7805 , n7806 , n7807 , n7808 , n7809 , n7810 , n7811 , n7812 , n7813 , n7814 , n7815 , n7816 , n7817 , n7818 , n7819 , n7820 , n7821 , n7822 , n7823 , n7824 , n7825 , n7826 , n7827 , n7828 , n7829 , n7830 , n7831 , n7832 , n7833 , n7834 , n7835 , n7836 , n7837 , n7838 , n7839 , n7840 , n7841 , n7842 , n7843 , n7844 , n7845 , n7846 , n7847 , n7848 , n7849 , n7850 , n7851 , n7852 , n7853 , n7854 , n7855 , n7856 , n7857 , n7858 , n7859 , n7860 , n7861 , n7862 , n7863 , n7864 , n7865 , n7866 , n7867 , n7868 , n7869 , n7870 , n7871 , n7872 , n7873 , n7874 , n7875 , n7876 , n7877 , n7878 , n7879 , n7880 , n7881 , n7882 , n7883 , n7884 , n7885 , n7886 , n7887 , n7888 , n7889 , n7890 , n7891 , n7892 , n7893 , n7894 , n7895 , n7896 , n7897 , n7898 , n7899 , n7900 , n7901 , n7902 , n7903 , n7904 , n7905 , n7906 , n7907 , n7908 , n7909 , n7910 , n7911 , n7912 , n7913 , n7914 , n7915 , n7916 , n7917 , n7918 , n7919 , n7920 , n7921 , n7922 , n7923 , n7924 , n7925 , n7926 , n7927 , n7928 , n7929 , n7930 , n7931 , n7932 , n7933 , n7934 , n7935 , n7936 , n7937 , n7938 , n7939 , n7940 , n7941 , n7942 , n7943 , n7944 , n7945 , n7946 , n7947 , n7948 , n7949 , n7950 , n7951 , n7952 , n7953 , n7954 , n7955 , n7956 , n7957 , n7958 , n7959 , n7960 , n7961 , n7962 , n7963 , n7964 , n7965 , n7966 , n7967 , n7968 , n7969 , n7970 , n7971 , n7972 , n7973 , n7974 , n7975 , n7976 , n7977 , n7978 , n7979 , n7980 , n7981 , n7982 , n7983 , n7984 , n7985 , n7986 , n7987 , n7988 , n7989 , n7990 , n7991 , n7992 , n7993 , n7994 , n7995 , n7996 , n7997 , n7998 , n7999 , n8000 , n8001 , n8002 , n8003 , n8004 , n8005 , n8006 , n8007 , n8008 , n8009 , n8010 , n8011 , n8012 , n8013 , n8014 , n8015 , n8016 , n8017 , n8018 , n8019 , n8020 , n8021 , n8022 , n8023 , n8024 , n8025 , n8026 , n8027 , n8028 , n8029 , n8030 , n8031 , n8032 , n8033 , n8034 , n8035 , n8036 , n8037 , n8038 , n8039 , n8040 , n8041 , n8042 , n8043 , n8044 , n8045 , n8046 , n8047 , n8048 , n8049 , n8050 , n8051 , n8052 , n8053 , n8054 , n8055 , n8056 , n8057 , n8058 , n8059 , n8060 , n8061 , n8062 , n8063 , n8064 , n8065 , n8066 , n8067 , n8068 , n8069 , n8070 , n8071 , n8072 , n8073 , n8074 , n8075 , n8076 , n8077 , n8078 , n8079 , n8080 , n8081 , n8082 , n8083 , n8084 , n8085 , n8086 , n8087 , n8088 , n8089 , n8090 , n8091 , n8092 , n8093 , n8094 , n8095 , n8096 , n8097 , n8098 , n8099 , n8100 , n8101 , n8102 , n8103 , n8104 , n8105 , n8106 , n8107 , n8108 , n8109 , n8110 , n8111 , n8112 , n8113 , n8114 , n8115 , n8116 , n8117 , n8118 , n8119 , n8120 , n8121 , n8122 , n8123 , n8124 , n8125 , n8126 , n8127 , n8128 , n8129 , n8130 , n8131 , n8132 , n8133 , n8134 , n8135 , n8136 , n8137 , n8138 , n8139 , n8140 , n8141 , n8142 , n8143 , n8144 , n8145 , n8146 , n8147 , n8148 , n8149 , n8150 , n8151 , n8152 , n8153 , n8154 , n8155 , n8156 , n8157 , n8158 , n8159 , n8160 , n8161 , n8162 , n8163 , n8164 , n8165 , n8166 , n8167 , n8168 , n8169 , n8170 , n8171 , n8172 , n8173 , n8174 , n8175 , n8176 , n8177 , n8178 , n8179 , n8180 , n8181 , n8182 , n8183 , n8184 , n8185 , n8186 , n8187 , n8188 , n8189 , n8190 , n8191 , n8192 , n8193 , n8194 , n8195 , n8196 , n8197 , n8198 , n8199 , n8200 , n8201 , n8202 , n8203 , n8204 , n8205 , n8206 , n8207 , n8208 , n8209 , n8210 , n8211 , n8212 , n8213 , n8214 , n8215 , n8216 , n8217 , n8218 , n8219 , n8220 , n8221 , n8222 , n8223 , n8224 , n8225 , n8226 , n8227 , n8228 , n8229 , n8230 , n8231 , n8232 , n8233 , n8234 , n8235 , n8236 , n8237 , n8238 , n8239 , n8240 , n8241 , n8242 , n8243 , n8244 , n8245 , n8246 , n8247 , n8248 , n8249 , n8250 , n8251 , n8252 , n8253 , n8254 , n8255 , n8256 , n8257 , n8258 , n8259 , n8260 , n8261 , n8262 , n8263 , n8264 , n8265 , n8266 , n8267 , n8268 , n8269 , n8270 , n8271 , n8272 , n8273 , n8274 , n8275 , n8276 , n8277 , n8278 , n8279 , n8280 , n8281 , n8282 , n8283 , n8284 , n8285 , n8286 , n8287 , n8288 , n8289 , n8290 , n8291 , n8292 , n8293 , n8294 , n8295 , n8296 , n8297 , n8298 , n8299 , n8300 , n8301 , n8302 , n8303 , n8304 , n8305 , n8306 , n8307 , n8308 , n8309 , n8310 , n8311 , n8312 , n8313 , n8314 , n8315 , n8316 , n8317 , n8318 , n8319 , n8320 , n8321 , n8322 , n8323 , n8324 , n8325 , n8326 , n8327 , n8328 , n8329 , n8330 , n8331 , n8332 , n8333 , n8334 , n8335 , n8336 , n8337 , n8338 , n8339 , n8340 , n8341 , n8342 , n8343 , n8344 , n8345 , n8346 , n8347 , n8348 , n8349 , n8350 , n8351 , n8352 , n8353 , n8354 , n8355 , n8356 , n8357 , n8358 , n8359 , n8360 , n8361 , n8362 , n8363 , n8364 , n8365 , n8366 , n8367 , n8368 , n8369 , n8370 , n8371 , n8372 , n8373 , n8374 , n8375 , n8376 , n8377 , n8378 , n8379 , n8380 , n8381 , n8382 , n8383 , n8384 , n8385 , n8386 , n8387 , n8388 , n8389 , n8390 , n8391 , n8392 , n8393 , n8394 , n8395 , n8396 , n8397 , n8398 , n8399 , n8400 , n8401 , n8402 , n8403 , n8404 , n8405 , n8406 , n8407 , n8408 , n8409 , n8410 , n8411 , n8412 , n8413 , n8414 , n8415 , n8416 , n8417 , n8418 , n8419 , n8420 , n8421 , n8422 , n8423 , n8424 , n8425 , n8426 , n8427 , n8428 , n8429 , n8430 , n8431 , n8432 , n8433 , n8434 , n8435 , n8436 , n8437 , n8438 , n8439 , n8440 , n8441 , n8442 , n8443 , n8444 , n8445 , n8446 , n8447 , n8448 , n8449 , n8450 , n8451 , n8452 , n8453 , n8454 , n8455 , n8456 , n8457 , n8458 , n8459 , n8460 , n8461 , n8462 , n8463 , n8464 , n8465 , n8466 , n8467 , n8468 , n8469 , n8470 , n8471 , n8472 , n8473 , n8474 , n8475 , n8476 , n8477 , n8478 , n8479 , n8480 , n8481 , n8482 , n8483 , n8484 , n8485 , n8486 , n8487 , n8488 , n8489 , n8490 , n8491 , n8492 , n8493 , n8494 , n8495 , n8496 , n8497 , n8498 , n8499 , n8500 , n8501 , n8502 , n8503 , n8504 , n8505 , n8506 , n8507 , n8508 , n8509 , n8510 , n8511 , n8512 , n8513 , n8514 , n8515 , n8516 , n8517 , n8518 , n8519 , n8520 , n8521 , n8522 , n8523 , n8524 , n8525 , n8526 , n8527 , n8528 , n8529 , n8530 , n8531 , n8532 , n8533 , n8534 , n8535 , n8536 , n8537 , n8538 , n8539 , n8540 , n8541 , n8542 , n8543 , n8544 , n8545 , n8546 , n8547 , n8548 , n8549 , n8550 , n8551 , n8552 , n8553 , n8554 , n8555 , n8556 , n8557 , n8558 , n8559 , n8560 , n8561 , n8562 , n8563 , n8564 , n8565 , n8566 , n8567 , n8568 , n8569 , n8570 , n8571 , n8572 , n8573 , n8574 , n8575 , n8576 , n8577 , n8578 , n8579 , n8580 , n8581 , n8582 , n8583 , n8584 , n8585 , n8586 , n8587 , n8588 , n8589 , n8590 , n8591 , n8592 , n8593 , n8594 , n8595 , n8596 , n8597 , n8598 , n8599 , n8600 , n8601 , n8602 , n8603 , n8604 , n8605 , n8606 , n8607 , n8608 , n8609 , n8610 , n8611 , n8612 , n8613 , n8614 , n8615 , n8616 , n8617 , n8618 , n8619 , n8620 , n8621 , n8622 , n8623 , n8624 , n8625 , n8626 , n8627 , n8628 , n8629 , n8630 , n8631 , n8632 , n8633 , n8634 , n8635 , n8636 , n8637 , n8638 , n8639 , n8640 , n8641 , n8642 , n8643 , n8644 , n8645 , n8646 , n8647 , n8648 , n8649 , n8650 , n8651 , n8652 , n8653 , n8654 , n8655 , n8656 , n8657 , n8658 , n8659 , n8660 , n8661 , n8662 , n8663 , n8664 , n8665 , n8666 , n8667 , n8668 , n8669 , n8670 , n8671 , n8672 , n8673 , n8674 , n8675 , n8676 , n8677 , n8678 , n8679 , n8680 , n8681 , n8682 , n8683 , n8684 , n8685 , n8686 , n8687 , n8688 , n8689 , n8690 , n8691 , n8692 , n8693 , n8694 , n8695 , n8696 , n8697 , n8698 , n8699 , n8700 , n8701 , n8702 , n8703 , n8704 , n8705 , n8706 , n8707 , n8708 , n8709 , n8710 , n8711 , n8712 , n8713 , n8714 , n8715 , n8716 , n8717 , n8718 , n8719 , n8720 , n8721 , n8722 , n8723 , n8724 , n8725 , n8726 , n8727 , n8728 , n8729 , n8730 , n8731 , n8732 , n8733 , n8734 , n8735 , n8736 , n8737 , n8738 , n8739 , n8740 , n8741 , n8742 , n8743 , n8744 , n8745 , n8746 , n8747 , n8748 , n8749 , n8750 , n8751 , n8752 , n8753 , n8754 , n8755 , n8756 , n8757 , n8758 , n8759 , n8760 , n8761 , n8762 , n8763 , n8764 , n8765 , n8766 , n8767 , n8768 , n8769 , n8770 , n8771 , n8772 , n8773 , n8774 , n8775 , n8776 , n8777 , n8778 , n8779 , n8780 , n8781 , n8782 , n8783 , n8784 , n8785 , n8786 , n8787 , n8788 , n8789 , n8790 , n8791 , n8792 , n8793 , n8794 , n8795 , n8796 , n8797 , n8798 , n8799 , n8800 , n8801 , n8802 , n8803 , n8804 , n8805 , n8806 , n8807 , n8808 , n8809 , n8810 , n8811 , n8812 , n8813 , n8814 , n8815 , n8816 , n8817 , n8818 , n8819 , n8820 , n8821 , n8822 , n8823 , n8824 , n8825 , n8826 , n8827 , n8828 , n8829 , n8830 , n8831 , n8832 , n8833 , n8834 , n8835 , n8836 , n8837 , n8838 , n8839 , n8840 , n8841 , n8842 , n8843 , n8844 , n8845 , n8846 , n8847 , n8848 , n8849 , n8850 , n8851 , n8852 , n8853 , n8854 , n8855 , n8856 , n8857 , n8858 , n8859 , n8860 , n8861 , n8862 , n8863 , n8864 , n8865 , n8866 , n8867 , n8868 , n8869 , n8870 , n8871 , n8872 , n8873 , n8874 , n8875 , n8876 , n8877 , n8878 , n8879 , n8880 , n8881 , n8882 , n8883 , n8884 , n8885 , n8886 , n8887 , n8888 , n8889 , n8890 , n8891 , n8892 , n8893 , n8894 , n8895 , n8896 , n8897 , n8898 , n8899 , n8900 , n8901 , n8902 , n8903 , n8904 , n8905 , n8906 , n8907 , n8908 , n8909 , n8910 , n8911 , n8912 , n8913 , n8914 , n8915 , n8916 , n8917 , n8918 , n8919 , n8920 , n8921 , n8922 , n8923 , n8924 , n8925 , n8926 , n8927 , n8928 , n8929 , n8930 , n8931 , n8932 , n8933 , n8934 , n8935 , n8936 , n8937 , n8938 , n8939 , n8940 , n8941 , n8942 , n8943 , n8944 , n8945 , n8946 , n8947 , n8948 , n8949 , n8950 , n8951 , n8952 , n8953 , n8954 , n8955 , n8956 , n8957 , n8958 , n8959 , n8960 , n8961 , n8962 , n8963 , n8964 , n8965 , n8966 , n8967 , n8968 , n8969 , n8970 , n8971 , n8972 , n8973 , n8974 , n8975 , n8976 , n8977 , n8978 , n8979 , n8980 , n8981 , n8982 , n8983 , n8984 , n8985 , n8986 , n8987 , n8988 , n8989 , n8990 , n8991 , n8992 , n8993 , n8994 , n8995 , n8996 , n8997 , n8998 , n8999 , n9000 , n9001 , n9002 , n9003 , n9004 , n9005 , n9006 , n9007 , n9008 , n9009 , n9010 , n9011 , n9012 , n9013 , n9014 , n9015 , n9016 , n9017 , n9018 , n9019 , n9020 , n9021 , n9022 , n9023 , n9024 , n9025 , n9026 , n9027 , n9028 , n9029 , n9030 , n9031 , n9032 , n9033 , n9034 , n9035 , n9036 , n9037 , n9038 , n9039 , n9040 , n9041 , n9042 , n9043 , n9044 , n9045 , n9046 , n9047 , n9048 , n9049 , n9050 , n9051 , n9052 , n9053 , n9054 , n9055 , n9056 , n9057 , n9058 , n9059 , n9060 , n9061 , n9062 , n9063 , n9064 , n9065 , n9066 , n9067 , n9068 , n9069 , n9070 , n9071 , n9072 , n9073 , n9074 , n9075 , n9076 , n9077 , n9078 , n9079 , n9080 , n9081 , n9082 , n9083 , n9084 , n9085 , n9086 , n9087 , n9088 , n9089 , n9090 , n9091 , n9092 , n9093 , n9094 , n9095 , n9096 , n9097 , n9098 , n9099 , n9100 , n9101 , n9102 , n9103 , n9104 , n9105 , n9106 , n9107 , n9108 , n9109 , n9110 , n9111 , n9112 , n9113 , n9114 , n9115 , n9116 , n9117 , n9118 , n9119 , n9120 , n9121 , n9122 , n9123 , n9124 , n9125 , n9126 , n9127 , n9128 , n9129 , n9130 , n9131 , n9132 , n9133 , n9134 , n9135 , n9136 , n9137 , n9138 , n9139 , n9140 , n9141 , n9142 , n9143 , n9144 , n9145 , n9146 , n9147 , n9148 , n9149 , n9150 , n9151 , n9152 , n9153 , n9154 , n9155 , n9156 , n9157 , n9158 , n9159 , n9160 , n9161 , n9162 , n9163 , n9164 , n9165 , n9166 , n9167 , n9168 , n9169 , n9170 , n9171 , n9172 , n9173 , n9174 , n9175 , n9176 , n9177 , n9178 , n9179 , n9180 , n9181 , n9182 , n9183 , n9184 , n9185 , n9186 , n9187 , n9188 , n9189 , n9190 , n9191 , n9192 , n9193 , n9194 , n9195 , n9196 , n9197 , n9198 , n9199 , n9200 , n9201 , n9202 , n9203 , n9204 , n9205 , n9206 , n9207 , n9208 , n9209 , n9210 , n9211 , n9212 , n9213 , n9214 , n9215 , n9216 , n9217 , n9218 , n9219 , n9220 , n9221 , n9222 , n9223 , n9224 , n9225 , n9226 , n9227 , n9228 , n9229 , n9230 , n9231 , n9232 , n9233 , n9234 , n9235 , n9236 , n9237 , n9238 , n9239 , n9240 , n9241 , n9242 , n9243 , n9244 , n9245 , n9246 , n9247 , n9248 , n9249 , n9250 , n9251 , n9252 , n9253 , n9254 , n9255 , n9256 , n9257 , n9258 , n9259 , n9260 , n9261 , n9262 , n9263 , n9264 , n9265 , n9266 , n9267 , n9268 , n9269 , n9270 , n9271 , n9272 , n9273 , n9274 , n9275 , n9276 , n9277 , n9278 , n9279 , n9280 , n9281 , n9282 , n9283 , n9284 , n9285 , n9286 , n9287 , n9288 , n9289 , n9290 , n9291 , n9292 , n9293 , n9294 , n9295 , n9296 , n9297 , n9298 , n9299 , n9300 , n9301 , n9302 , n9303 , n9304 , n9305 , n9306 , n9307 , n9308 , n9309 , n9310 , n9311 , n9312 , n9313 , n9314 , n9315 , n9316 , n9317 , n9318 , n9319 , n9320 , n9321 , n9322 , n9323 , n9324 , n9325 , n9326 , n9327 , n9328 , n9329 , n9330 , n9331 , n9332 , n9333 , n9334 , n9335 , n9336 , n9337 , n9338 , n9339 , n9340 , n9341 , n9342 , n9343 , n9344 , n9345 , n9346 , n9347 , n9348 , n9349 , n9350 , n9351 , n9352 , n9353 , n9354 , n9355 , n9356 , n9357 , n9358 , n9359 , n9360 , n9361 , n9362 , n9363 , n9364 , n9365 , n9366 , n9367 , n9368 , n9369 , n9370 , n9371 , n9372 , n9373 , n9374 , n9375 , n9376 , n9377 , n9378 , n9379 , n9380 , n9381 , n9382 , n9383 , n9384 , n9385 , n9386 , n9387 , n9388 , n9389 , n9390 , n9391 , n9392 , n9393 , n9394 , n9395 , n9396 , n9397 , n9398 , n9399 , n9400 , n9401 , n9402 , n9403 , n9404 , n9405 , n9406 , n9407 , n9408 , n9409 , n9410 , n9411 , n9412 , n9413 , n9414 , n9415 , n9416 , n9417 , n9418 , n9419 , n9420 , n9421 , n9422 , n9423 , n9424 , n9425 , n9426 , n9427 , n9428 , n9429 , n9430 , n9431 , n9432 , n9433 , n9434 , n9435 , n9436 , n9437 , n9438 , n9439 , n9440 , n9441 , n9442 , n9443 , n9444 , n9445 , n9446 , n9447 , n9448 , n9449 , n9450 , n9451 , n9452 , n9453 , n9454 , n9455 , n9456 , n9457 , n9458 , n9459 , n9460 , n9461 , n9462 , n9463 , n9464 , n9465 , n9466 , n9467 , n9468 , n9469 , n9470 , n9471 , n9472 , n9473 , n9474 , n9475 , n9476 , n9477 , n9478 , n9479 , n9480 , n9481 , n9482 , n9483 , n9484 , n9485 , n9486 , n9487 , n9488 , n9489 , n9490 , n9491 , n9492 , n9493 , n9494 , n9495 , n9496 , n9497 , n9498 , n9499 , n9500 , n9501 , n9502 , n9503 , n9504 , n9505 , n9506 , n9507 , n9508 , n9509 , n9510 , n9511 , n9512 , n9513 , n9514 , n9515 , n9516 , n9517 , n9518 , n9519 , n9520 , n9521 , n9522 , n9523 , n9524 , n9525 , n9526 , n9527 , n9528 , n9529 , n9530 , n9531 , n9532 , n9533 , n9534 , n9535 , n9536 , n9537 , n9538 , n9539 , n9540 , n9541 , n9542 , n9543 , n9544 , n9545 , n9546 , n9547 , n9548 , n9549 , n9550 , n9551 , n9552 , n9553 , n9554 , n9555 , n9556 , n9557 , n9558 , n9559 , n9560 , n9561 , n9562 , n9563 , n9564 , n9565 , n9566 , n9567 , n9568 , n9569 , n9570 , n9571 , n9572 , n9573 , n9574 , n9575 , n9576 , n9577 , n9578 , n9579 , n9580 , n9581 , n9582 , n9583 , n9584 , n9585 , n9586 , n9587 , n9588 , n9589 , n9590 , n9591 , n9592 , n9593 , n9594 , n9595 , n9596 , n9597 , n9598 , n9599 , n9600 , n9601 , n9602 , n9603 , n9604 , n9605 , n9606 , n9607 , n9608 , n9609 , n9610 , n9611 , n9612 , n9613 , n9614 , n9615 , n9616 , n9617 , n9618 , n9619 , n9620 , n9621 , n9622 , n9623 , n9624 , n9625 , n9626 , n9627 , n9628 , n9629 , n9630 , n9631 , n9632 , n9633 , n9634 , n9635 , n9636 , n9637 , n9638 , n9639 , n9640 , n9641 , n9642 , n9643 , n9644 , n9645 , n9646 , n9647 , n9648 , n9649 , n9650 , n9651 , n9652 , n9653 , n9654 , n9655 , n9656 , n9657 , n9658 , n9659 , n9660 , n9661 , n9662 , n9663 , n9664 , n9665 , n9666 , n9667 , n9668 , n9669 , n9670 , n9671 , n9672 , n9673 , n9674 , n9675 , n9676 , n9677 , n9678 , n9679 , n9680 , n9681 , n9682 , n9683 , n9684 , n9685 , n9686 , n9687 , n9688 , n9689 , n9690 , n9691 , n9692 , n9693 , n9694 , n9695 , n9696 , n9697 , n9698 , n9699 , n9700 , n9701 , n9702 , n9703 , n9704 , n9705 , n9706 , n9707 , n9708 , n9709 , n9710 , n9711 , n9712 , n9713 , n9714 , n9715 , n9716 , n9717 , n9718 , n9719 , n9720 , n9721 , n9722 , n9723 , n9724 , n9725 , n9726 , n9727 , n9728 , n9729 , n9730 , n9731 , n9732 , n9733 , n9734 , n9735 , n9736 , n9737 , n9738 , n9739 , n9740 , n9741 , n9742 , n9743 , n9744 , n9745 , n9746 , n9747 , n9748 , n9749 , n9750 , n9751 , n9752 , n9753 , n9754 , n9755 , n9756 , n9757 , n9758 , n9759 , n9760 , n9761 , n9762 , n9763 , n9764 , n9765 , n9766 , n9767 , n9768 , n9769 , n9770 , n9771 , n9772 , n9773 , n9774 , n9775 , n9776 , n9777 , n9778 , n9779 , n9780 , n9781 , n9782 , n9783 , n9784 , n9785 , n9786 , n9787 , n9788 , n9789 , n9790 , n9791 , n9792 , n9793 , n9794 , n9795 , n9796 , n9797 , n9798 , n9799 , n9800 , n9801 , n9802 , n9803 , n9804 , n9805 , n9806 , n9807 , n9808 , n9809 , n9810 , n9811 , n9812 , n9813 , n9814 , n9815 , n9816 , n9817 , n9818 , n9819 , n9820 , n9821 , n9822 , n9823 , n9824 , n9825 , n9826 , n9827 , n9828 , n9829 , n9830 , n9831 , n9832 , n9833 , n9834 , n9835 , n9836 , n9837 , n9838 , n9839 , n9840 , n9841 , n9842 , n9843 , n9844 , n9845 , n9846 , n9847 , n9848 , n9849 , n9850 , n9851 , n9852 , n9853 , n9854 , n9855 , n9856 , n9857 , n9858 , n9859 , n9860 , n9861 , n9862 , n9863 , n9864 , n9865 , n9866 , n9867 , n9868 , n9869 , n9870 , n9871 , n9872 , n9873 , n9874 , n9875 , n9876 , n9877 , n9878 , n9879 , n9880 , n9881 , n9882 , n9883 , n9884 , n9885 , n9886 , n9887 , n9888 , n9889 , n9890 , n9891 , n9892 , n9893 , n9894 , n9895 , n9896 , n9897 , n9898 , n9899 , n9900 , n9901 , n9902 , n9903 , n9904 , n9905 , n9906 , n9907 , n9908 , n9909 , n9910 , n9911 , n9912 , n9913 , n9914 , n9915 , n9916 , n9917 , n9918 , n9919 , n9920 , n9921 , n9922 , n9923 , n9924 , n9925 , n9926 , n9927 , n9928 , n9929 , n9930 , n9931 , n9932 , n9933 , n9934 , n9935 , n9936 , n9937 , n9938 , n9939 , n9940 , n9941 , n9942 , n9943 , n9944 , n9945 , n9946 , n9947 , n9948 , n9949 , n9950 , n9951 , n9952 , n9953 , n9954 , n9955 , n9956 , n9957 , n9958 , n9959 , n9960 , n9961 , n9962 , n9963 , n9964 , n9965 , n9966 , n9967 , n9968 , n9969 , n9970 , n9971 , n9972 , n9973 , n9974 , n9975 , n9976 , n9977 , n9978 , n9979 , n9980 , n9981 , n9982 , n9983 , n9984 , n9985 , n9986 , n9987 , n9988 , n9989 , n9990 , n9991 , n9992 , n9993 , n9994 , n9995 , n9996 , n9997 , n9998 , n9999 , n10000 , n10001 , n10002 , n10003 , n10004 , n10005 , n10006 , n10007 , n10008 , n10009 , n10010 , n10011 , n10012 , n10013 , n10014 , n10015 , n10016 , n10017 , n10018 , n10019 , n10020 , n10021 , n10022 , n10023 , n10024 , n10025 , n10026 , n10027 , n10028 , n10029 , n10030 , n10031 , n10032 , n10033 , n10034 , n10035 , n10036 , n10037 , n10038 , n10039 , n10040 , n10041 , n10042 , n10043 , n10044 , n10045 , n10046 , n10047 , n10048 , n10049 , n10050 , n10051 , n10052 , n10053 , n10054 , n10055 , n10056 , n10057 , n10058 , n10059 , n10060 , n10061 , n10062 , n10063 , n10064 , n10065 , n10066 , n10067 , n10068 , n10069 , n10070 , n10071 , n10072 , n10073 , n10074 , n10075 , n10076 , n10077 , n10078 , n10079 , n10080 , n10081 , n10082 , n10083 , n10084 , n10085 , n10086 , n10087 , n10088 , n10089 , n10090 , n10091 , n10092 , n10093 , n10094 , n10095 , n10096 , n10097 , n10098 , n10099 , n10100 , n10101 , n10102 , n10103 , n10104 , n10105 , n10106 , n10107 , n10108 , n10109 , n10110 , n10111 , n10112 , n10113 , n10114 , n10115 , n10116 , n10117 , n10118 , n10119 , n10120 , n10121 , n10122 , n10123 , n10124 , n10125 , n10126 , n10127 , n10128 , n10129 , n10130 , n10131 , n10132 , n10133 , n10134 , n10135 , n10136 , n10137 , n10138 , n10139 , n10140 , n10141 , n10142 , n10143 , n10144 , n10145 , n10146 , n10147 , n10148 , n10149 , n10150 , n10151 , n10152 , n10153 , n10154 , n10155 , n10156 , n10157 , n10158 , n10159 , n10160 , n10161 , n10162 , n10163 , n10164 , n10165 , n10166 , n10167 , n10168 , n10169 , n10170 , n10171 , n10172 , n10173 , n10174 , n10175 , n10176 , n10177 , n10178 , n10179 , n10180 , n10181 , n10182 , n10183 , n10184 , n10185 , n10186 , n10187 , n10188 , n10189 , n10190 , n10191 , n10192 , n10193 , n10194 , n10195 , n10196 , n10197 , n10198 , n10199 , n10200 , n10201 , n10202 , n10203 , n10204 , n10205 , n10206 , n10207 , n10208 , n10209 , n10210 , n10211 , n10212 , n10213 , n10214 , n10215 , n10216 , n10217 , n10218 , n10219 , n10220 , n10221 , n10222 , n10223 , n10224 , n10225 , n10226 , n10227 , n10228 , n10229 , n10230 , n10231 , n10232 , n10233 , n10234 , n10235 , n10236 , n10237 , n10238 , n10239 , n10240 , n10241 , n10242 , n10243 , n10244 , n10245 , n10246 , n10247 , n10248 , n10249 , n10250 , n10251 , n10252 , n10253 , n10254 , n10255 , n10256 , n10257 , n10258 , n10259 , n10260 , n10261 , n10262 , n10263 , n10264 , n10265 , n10266 , n10267 , n10268 , n10269 , n10270 , n10271 , n10272 , n10273 , n10274 , n10275 , n10276 , n10277 , n10278 , n10279 , n10280 , n10281 , n10282 , n10283 , n10284 , n10285 , n10286 , n10287 , n10288 , n10289 , n10290 , n10291 , n10292 , n10293 , n10294 , n10295 , n10296 , n10297 , n10298 , n10299 , n10300 , n10301 , n10302 , n10303 , n10304 , n10305 , n10306 , n10307 , n10308 , n10309 , n10310 , n10311 , n10312 , n10313 , n10314 , n10315 , n10316 , n10317 , n10318 , n10319 , n10320 , n10321 , n10322 , n10323 , n10324 , n10325 , n10326 , n10327 , n10328 , n10329 , n10330 , n10331 , n10332 , n10333 , n10334 , n10335 , n10336 , n10337 , n10338 , n10339 , n10340 , n10341 , n10342 , n10343 , n10344 , n10345 , n10346 , n10347 , n10348 , n10349 , n10350 , n10351 , n10352 , n10353 , n10354 , n10355 , n10356 , n10357 , n10358 , n10359 , n10360 , n10361 , n10362 , n10363 , n10364 , n10365 , n10366 , n10367 , n10368 , n10369 , n10370 , n10371 , n10372 , n10373 , n10374 , n10375 , n10376 , n10377 , n10378 , n10379 , n10380 , n10381 , n10382 , n10383 , n10384 , n10385 , n10386 , n10387 , n10388 , n10389 , n10390 , n10391 , n10392 , n10393 , n10394 , n10395 , n10396 , n10397 , n10398 , n10399 , n10400 , n10401 , n10402 , n10403 , n10404 , n10405 , n10406 , n10407 , n10408 , n10409 , n10410 , n10411 , n10412 , n10413 , n10414 , n10415 , n10416 , n10417 , n10418 , n10419 , n10420 , n10421 , n10422 , n10423 , n10424 , n10425 , n10426 , n10427 , n10428 , n10429 , n10430 , n10431 , n10432 , n10433 , n10434 , n10435 , n10436 , n10437 , n10438 , n10439 , n10440 , n10441 , n10442 , n10443 , n10444 , n10445 , n10446 , n10447 , n10448 , n10449 , n10450 , n10451 , n10452 , n10453 , n10454 , n10455 , n10456 , n10457 , n10458 , n10459 , n10460 , n10461 , n10462 , n10463 , n10464 , n10465 , n10466 , n10467 , n10468 , n10469 , n10470 , n10471 , n10472 , n10473 , n10474 , n10475 , n10476 , n10477 , n10478 , n10479 , n10480 , n10481 , n10482 , n10483 , n10484 , n10485 , n10486 , n10487 , n10488 , n10489 , n10490 , n10491 , n10492 , n10493 , n10494 , n10495 , n10496 , n10497 , n10498 , n10499 , n10500 , n10501 , n10502 , n10503 , n10504 , n10505 , n10506 , n10507 , n10508 , n10509 , n10510 , n10511 , n10512 , n10513 , n10514 , n10515 , n10516 , n10517 , n10518 , n10519 , n10520 , n10521 , n10522 , n10523 , n10524 , n10525 , n10526 , n10527 , n10528 , n10529 , n10530 , n10531 , n10532 , n10533 , n10534 , n10535 , n10536 , n10537 , n10538 , n10539 , n10540 , n10541 , n10542 , n10543 , n10544 , n10545 , n10546 , n10547 , n10548 , n10549 , n10550 , n10551 , n10552 , n10553 , n10554 , n10555 , n10556 , n10557 , n10558 , n10559 , n10560 , n10561 , n10562 , n10563 , n10564 , n10565 , n10566 , n10567 , n10568 , n10569 , n10570 , n10571 , n10572 , n10573 , n10574 , n10575 , n10576 , n10577 , n10578 , n10579 , n10580 , n10581 , n10582 , n10583 , n10584 , n10585 , n10586 , n10587 , n10588 , n10589 , n10590 , n10591 , n10592 , n10593 , n10594 , n10595 , n10596 , n10597 , n10598 , n10599 , n10600 , n10601 , n10602 , n10603 , n10604 , n10605 , n10606 , n10607 , n10608 , n10609 , n10610 , n10611 , n10612 , n10613 , n10614 , n10615 , n10616 , n10617 , n10618 , n10619 , n10620 , n10621 , n10622 , n10623 , n10624 , n10625 , n10626 , n10627 , n10628 , n10629 , n10630 , n10631 , n10632 , n10633 , n10634 , n10635 , n10636 , n10637 , n10638 , n10639 , n10640 , n10641 , n10642 , n10643 , n10644 , n10645 , n10646 , n10647 , n10648 , n10649 , n10650 , n10651 , n10652 , n10653 , n10654 , n10655 , n10656 , n10657 , n10658 , n10659 , n10660 , n10661 , n10662 , n10663 , n10664 , n10665 , n10666 , n10667 , n10668 , n10669 , n10670 , n10671 , n10672 , n10673 , n10674 , n10675 , n10676 , n10677 , n10678 , n10679 , n10680 , n10681 , n10682 , n10683 , n10684 , n10685 , n10686 , n10687 , n10688 , n10689 , n10690 , n10691 , n10692 , n10693 , n10694 , n10695 , n10696 , n10697 , n10698 , n10699 , n10700 , n10701 , n10702 , n10703 , n10704 , n10705 , n10706 , n10707 , n10708 , n10709 , n10710 , n10711 , n10712 , n10713 , n10714 , n10715 , n10716 , n10717 , n10718 , n10719 , n10720 , n10721 , n10722 , n10723 , n10724 , n10725 , n10726 , n10727 , n10728 , n10729 , n10730 , n10731 , n10732 , n10733 , n10734 , n10735 , n10736 , n10737 , n10738 , n10739 , n10740 , n10741 , n10742 , n10743 , n10744 , n10745 , n10746 , n10747 , n10748 , n10749 , n10750 , n10751 , n10752 , n10753 , n10754 , n10755 , n10756 , n10757 , n10758 , n10759 , n10760 , n10761 , n10762 , n10763 , n10764 , n10765 , n10766 , n10767 , n10768 , n10769 , n10770 , n10771 , n10772 , n10773 , n10774 , n10775 , n10776 , n10777 , n10778 , n10779 , n10780 , n10781 , n10782 , n10783 , n10784 , n10785 , n10786 , n10787 , n10788 , n10789 , n10790 , n10791 , n10792 , n10793 , n10794 , n10795 , n10796 , n10797 , n10798 , n10799 , n10800 , n10801 , n10802 , n10803 , n10804 , n10805 , n10806 , n10807 , n10808 , n10809 , n10810 , n10811 , n10812 , n10813 , n10814 , n10815 , n10816 , n10817 , n10818 , n10819 , n10820 , n10821 , n10822 , n10823 , n10824 , n10825 , n10826 , n10827 , n10828 , n10829 , n10830 , n10831 , n10832 , n10833 , n10834 , n10835 , n10836 , n10837 , n10838 , n10839 , n10840 , n10841 , n10842 , n10843 , n10844 , n10845 , n10846 , n10847 , n10848 , n10849 , n10850 , n10851 , n10852 , n10853 , n10854 , n10855 , n10856 , n10857 , n10858 , n10859 , n10860 , n10861 , n10862 , n10863 , n10864 , n10865 , n10866 , n10867 , n10868 , n10869 , n10870 , n10871 , n10872 , n10873 , n10874 , n10875 , n10876 , n10877 , n10878 , n10879 , n10880 , n10881 , n10882 , n10883 , n10884 , n10885 , n10886 , n10887 , n10888 , n10889 , n10890 , n10891 , n10892 , n10893 , n10894 , n10895 , n10896 , n10897 , n10898 , n10899 , n10900 , n10901 , n10902 , n10903 , n10904 , n10905 , n10906 , n10907 , n10908 , n10909 , n10910 , n10911 , n10912 , n10913 , n10914 , n10915 , n10916 , n10917 , n10918 , n10919 , n10920 , n10921 , n10922 , n10923 , n10924 , n10925 , n10926 , n10927 , n10928 , n10929 , n10930 , n10931 , n10932 , n10933 , n10934 , n10935 , n10936 , n10937 , n10938 , n10939 , n10940 , n10941 , n10942 , n10943 , n10944 , n10945 , n10946 , n10947 , n10948 , n10949 , n10950 , n10951 , n10952 , n10953 , n10954 , n10955 , n10956 , n10957 , n10958 , n10959 , n10960 , n10961 , n10962 , n10963 , n10964 , n10965 , n10966 , n10967 , n10968 , n10969 , n10970 , n10971 , n10972 , n10973 , n10974 , n10975 , n10976 , n10977 , n10978 , n10979 , n10980 , n10981 , n10982 , n10983 , n10984 , n10985 , n10986 , n10987 , n10988 , n10989 , n10990 , n10991 , n10992 , n10993 , n10994 , n10995 , n10996 , n10997 , n10998 , n10999 , n11000 , n11001 , n11002 , n11003 , n11004 , n11005 , n11006 , n11007 , n11008 , n11009 , n11010 , n11011 , n11012 , n11013 , n11014 , n11015 , n11016 , n11017 , n11018 , n11019 , n11020 , n11021 , n11022 , n11023 , n11024 , n11025 , n11026 , n11027 , n11028 , n11029 , n11030 , n11031 , n11032 , n11033 , n11034 , n11035 , n11036 , n11037 , n11038 , n11039 , n11040 , n11041 , n11042 , n11043 , n11044 , n11045 , n11046 , n11047 , n11048 , n11049 , n11050 , n11051 , n11052 , n11053 , n11054 , n11055 , n11056 , n11057 , n11058 , n11059 , n11060 , n11061 , n11062 , n11063 , n11064 , n11065 , n11066 , n11067 , n11068 , n11069 , n11070 , n11071 , n11072 , n11073 , n11074 , n11075 , n11076 , n11077 , n11078 , n11079 , n11080 , n11081 , n11082 , n11083 , n11084 , n11085 , n11086 , n11087 , n11088 , n11089 , n11090 , n11091 , n11092 , n11093 , n11094 , n11095 , n11096 , n11097 , n11098 , n11099 , n11100 , n11101 , n11102 , n11103 , n11104 , n11105 , n11106 , n11107 , n11108 , n11109 , n11110 , n11111 , n11112 , n11113 , n11114 , n11115 , n11116 , n11117 , n11118 , n11119 , n11120 , n11121 , n11122 , n11123 , n11124 , n11125 , n11126 , n11127 , n11128 , n11129 , n11130 , n11131 , n11132 , n11133 , n11134 , n11135 , n11136 , n11137 , n11138 , n11139 , n11140 , n11141 , n11142 , n11143 , n11144 , n11145 , n11146 , n11147 , n11148 , n11149 , n11150 , n11151 , n11152 , n11153 , n11154 , n11155 , n11156 , n11157 , n11158 , n11159 , n11160 , n11161 , n11162 , n11163 , n11164 , n11165 , n11166 , n11167 , n11168 , n11169 , n11170 , n11171 , n11172 , n11173 , n11174 , n11175 , n11176 , n11177 , n11178 , n11179 , n11180 , n11181 , n11182 , n11183 , n11184 , n11185 , n11186 , n11187 , n11188 , n11189 , n11190 , n11191 , n11192 , n11193 , n11194 , n11195 , n11196 , n11197 , n11198 , n11199 , n11200 , n11201 , n11202 , n11203 , n11204 , n11205 , n11206 , n11207 , n11208 , n11209 , n11210 , n11211 , n11212 , n11213 , n11214 , n11215 , n11216 , n11217 , n11218 , n11219 , n11220 , n11221 , n11222 , n11223 , n11224 , n11225 , n11226 , n11227 , n11228 , n11229 , n11230 , n11231 , n11232 , n11233 , n11234 , n11235 , n11236 , n11237 , n11238 , n11239 , n11240 , n11241 , n11242 , n11243 , n11244 , n11245 , n11246 , n11247 , n11248 , n11249 , n11250 , n11251 , n11252 , n11253 , n11254 , n11255 , n11256 , n11257 , n11258 , n11259 , n11260 , n11261 , n11262 , n11263 , n11264 , n11265 , n11266 , n11267 , n11268 , n11269 , n11270 , n11271 , n11272 , n11273 , n11274 , n11275 , n11276 , n11277 , n11278 , n11279 , n11280 , n11281 , n11282 , n11283 , n11284 , n11285 , n11286 , n11287 , n11288 , n11289 , n11290 , n11291 , n11292 , n11293 , n11294 , n11295 , n11296 , n11297 , n11298 , n11299 , n11300 , n11301 , n11302 , n11303 , n11304 , n11305 , n11306 , n11307 , n11308 , n11309 , n11310 , n11311 , n11312 , n11313 , n11314 , n11315 , n11316 , n11317 , n11318 , n11319 , n11320 , n11321 , n11322 , n11323 , n11324 , n11325 , n11326 , n11327 , n11328 , n11329 , n11330 , n11331 , n11332 , n11333 , n11334 , n11335 , n11336 , n11337 , n11338 , n11339 , n11340 , n11341 , n11342 , n11343 , n11344 , n11345 , n11346 , n11347 , n11348 , n11349 , n11350 , n11351 , n11352 , n11353 , n11354 , n11355 , n11356 , n11357 , n11358 , n11359 , n11360 , n11361 , n11362 , n11363 , n11364 , n11365 , n11366 , n11367 , n11368 , n11369 , n11370 , n11371 , n11372 , n11373 , n11374 , n11375 , n11376 , n11377 , n11378 , n11379 , n11380 , n11381 , n11382 , n11383 , n11384 , n11385 , n11386 , n11387 , n11388 , n11389 , n11390 , n11391 , n11392 , n11393 , n11394 , n11395 , n11396 , n11397 , n11398 , n11399 , n11400 , n11401 , n11402 , n11403 , n11404 , n11405 , n11406 , n11407 , n11408 , n11409 , n11410 , n11411 , n11412 , n11413 , n11414 , n11415 , n11416 , n11417 , n11418 , n11419 , n11420 , n11421 , n11422 , n11423 , n11424 , n11425 , n11426 , n11427 , n11428 , n11429 , n11430 , n11431 , n11432 , n11433 , n11434 , n11435 , n11436 , n11437 , n11438 , n11439 , n11440 , n11441 , n11442 , n11443 , n11444 , n11445 , n11446 , n11447 , n11448 , n11449 , n11450 , n11451 , n11452 , n11453 , n11454 , n11455 , n11456 , n11457 , n11458 , n11459 , n11460 , n11461 , n11462 , n11463 , n11464 , n11465 , n11466 , n11467 , n11468 , n11469 , n11470 , n11471 , n11472 , n11473 , n11474 , n11475 , n11476 , n11477 , n11478 , n11479 , n11480 , n11481 , n11482 , n11483 , n11484 , n11485 , n11486 , n11487 , n11488 , n11489 , n11490 , n11491 , n11492 , n11493 , n11494 , n11495 , n11496 , n11497 , n11498 , n11499 , n11500 , n11501 , n11502 , n11503 , n11504 , n11505 , n11506 , n11507 , n11508 , n11509 , n11510 , n11511 , n11512 , n11513 , n11514 , n11515 , n11516 , n11517 , n11518 , n11519 , n11520 , n11521 , n11522 , n11523 , n11524 , n11525 , n11526 , n11527 , n11528 , n11529 , n11530 , n11531 , n11532 , n11533 , n11534 , n11535 , n11536 , n11537 , n11538 , n11539 , n11540 , n11541 , n11542 , n11543 , n11544 , n11545 , n11546 , n11547 , n11548 , n11549 , n11550 , n11551 , n11552 , n11553 , n11554 , n11555 , n11556 , n11557 , n11558 , n11559 , n11560 , n11561 , n11562 , n11563 , n11564 , n11565 , n11566 , n11567 , n11568 , n11569 , n11570 , n11571 , n11572 , n11573 , n11574 , n11575 , n11576 , n11577 , n11578 , n11579 , n11580 , n11581 , n11582 , n11583 , n11584 , n11585 , n11586 , n11587 , n11588 , n11589 , n11590 , n11591 , n11592 , n11593 , n11594 , n11595 , n11596 , n11597 , n11598 , n11599 , n11600 , n11601 , n11602 , n11603 , n11604 , n11605 , n11606 , n11607 , n11608 , n11609 , n11610 , n11611 , n11612 , n11613 , n11614 , n11615 , n11616 , n11617 , n11618 , n11619 , n11620 , n11621 , n11622 , n11623 , n11624 , n11625 , n11626 , n11627 , n11628 , n11629 , n11630 , n11631 , n11632 , n11633 , n11634 , n11635 , n11636 , n11637 , n11638 , n11639 , n11640 , n11641 , n11642 , n11643 , n11644 , n11645 , n11646 , n11647 , n11648 , n11649 , n11650 , n11651 , n11652 , n11653 , n11654 , n11655 , n11656 , n11657 , n11658 , n11659 , n11660 , n11661 , n11662 , n11663 , n11664 , n11665 , n11666 , n11667 , n11668 , n11669 , n11670 , n11671 , n11672 , n11673 , n11674 , n11675 , n11676 , n11677 , n11678 , n11679 , n11680 , n11681 , n11682 , n11683 , n11684 , n11685 , n11686 , n11687 , n11688 , n11689 , n11690 , n11691 , n11692 , n11693 , n11694 , n11695 , n11696 , n11697 , n11698 , n11699 , n11700 , n11701 , n11702 , n11703 , n11704 , n11705 , n11706 , n11707 , n11708 , n11709 , n11710 , n11711 , n11712 , n11713 , n11714 , n11715 , n11716 , n11717 , n11718 , n11719 , n11720 , n11721 , n11722 , n11723 , n11724 , n11725 , n11726 , n11727 , n11728 , n11729 , n11730 , n11731 , n11732 , n11733 , n11734 , n11735 , n11736 , n11737 , n11738 , n11739 , n11740 , n11741 , n11742 , n11743 , n11744 , n11745 , n11746 , n11747 , n11748 , n11749 , n11750 , n11751 , n11752 , n11753 , n11754 , n11755 , n11756 , n11757 , n11758 , n11759 , n11760 , n11761 , n11762 , n11763 , n11764 , n11765 , n11766 , n11767 , n11768 , n11769 , n11770 , n11771 , n11772 , n11773 , n11774 , n11775 , n11776 , n11777 , n11778 , n11779 , n11780 , n11781 , n11782 , n11783 , n11784 , n11785 , n11786 , n11787 , n11788 , n11789 , n11790 , n11791 , n11792 , n11793 , n11794 , n11795 , n11796 , n11797 , n11798 , n11799 , n11800 , n11801 , n11802 , n11803 , n11804 , n11805 , n11806 , n11807 , n11808 , n11809 , n11810 , n11811 , n11812 , n11813 , n11814 , n11815 , n11816 , n11817 , n11818 , n11819 , n11820 , n11821 , n11822 , n11823 , n11824 , n11825 , n11826 , n11827 , n11828 , n11829 , n11830 , n11831 , n11832 , n11833 , n11834 , n11835 , n11836 , n11837 , n11838 , n11839 , n11840 , n11841 , n11842 , n11843 , n11844 , n11845 , n11846 , n11847 , n11848 , n11849 , n11850 , n11851 , n11852 , n11853 , n11854 , n11855 , n11856 , n11857 , n11858 , n11859 , n11860 , n11861 , n11862 , n11863 , n11864 , n11865 , n11866 , n11867 , n11868 , n11869 , n11870 , n11871 , n11872 , n11873 , n11874 , n11875 , n11876 , n11877 , n11878 , n11879 , n11880 , n11881 , n11882 , n11883 , n11884 , n11885 , n11886 , n11887 , n11888 , n11889 , n11890 , n11891 , n11892 , n11893 , n11894 , n11895 , n11896 , n11897 , n11898 , n11899 , n11900 , n11901 , n11902 , n11903 , n11904 , n11905 , n11906 , n11907 , n11908 , n11909 , n11910 , n11911 , n11912 , n11913 , n11914 , n11915 , n11916 , n11917 , n11918 , n11919 , n11920 , n11921 , n11922 , n11923 , n11924 , n11925 , n11926 , n11927 , n11928 , n11929 , n11930 , n11931 , n11932 , n11933 , n11934 , n11935 , n11936 , n11937 , n11938 , n11939 , n11940 , n11941 , n11942 , n11943 , n11944 , n11945 , n11946 , n11947 , n11948 , n11949 , n11950 , n11951 , n11952 , n11953 , n11954 , n11955 , n11956 , n11957 , n11958 , n11959 , n11960 , n11961 , n11962 , n11963 , n11964 , n11965 , n11966 , n11967 , n11968 , n11969 , n11970 , n11971 , n11972 , n11973 , n11974 , n11975 , n11976 , n11977 , n11978 , n11979 , n11980 , n11981 , n11982 , n11983 , n11984 , n11985 , n11986 , n11987 , n11988 , n11989 , n11990 , n11991 , n11992 , n11993 , n11994 , n11995 , n11996 , n11997 , n11998 , n11999 , n12000 , n12001 , n12002 , n12003 , n12004 , n12005 , n12006 , n12007 , n12008 , n12009 , n12010 , n12011 , n12012 , n12013 , n12014 , n12015 , n12016 , n12017 , n12018 , n12019 , n12020 , n12021 , n12022 , n12023 , n12024 , n12025 , n12026 , n12027 , n12028 , n12029 , n12030 , n12031 , n12032 , n12033 , n12034 , n12035 , n12036 , n12037 , n12038 , n12039 , n12040 , n12041 , n12042 , n12043 , n12044 , n12045 , n12046 , n12047 , n12048 , n12049 , n12050 , n12051 , n12052 , n12053 , n12054 , n12055 , n12056 , n12057 , n12058 , n12059 , n12060 , n12061 , n12062 , n12063 , n12064 , n12065 , n12066 , n12067 , n12068 , n12069 , n12070 , n12071 , n12072 , n12073 , n12074 , n12075 , n12076 , n12077 , n12078 , n12079 , n12080 , n12081 , n12082 , n12083 , n12084 , n12085 , n12086 , n12087 , n12088 , n12089 , n12090 , n12091 , n12092 , n12093 , n12094 , n12095 , n12096 , n12097 , n12098 , n12099 , n12100 , n12101 , n12102 , n12103 , n12104 , n12105 , n12106 , n12107 , n12108 , n12109 , n12110 , n12111 , n12112 , n12113 , n12114 , n12115 , n12116 , n12117 , n12118 , n12119 , n12120 , n12121 , n12122 , n12123 , n12124 , n12125 , n12126 , n12127 , n12128 , n12129 , n12130 , n12131 , n12132 , n12133 , n12134 , n12135 , n12136 , n12137 , n12138 , n12139 , n12140 , n12141 , n12142 , n12143 , n12144 , n12145 , n12146 , n12147 , n12148 , n12149 , n12150 , n12151 , n12152 , n12153 , n12154 , n12155 , n12156 , n12157 , n12158 , n12159 , n12160 , n12161 , n12162 , n12163 , n12164 , n12165 , n12166 , n12167 , n12168 , n12169 , n12170 , n12171 , n12172 , n12173 , n12174 , n12175 , n12176 , n12177 , n12178 , n12179 , n12180 , n12181 , n12182 , n12183 , n12184 , n12185 , n12186 , n12187 , n12188 , n12189 , n12190 , n12191 , n12192 , n12193 , n12194 , n12195 , n12196 , n12197 , n12198 , n12199 , n12200 , n12201 , n12202 , n12203 , n12204 , n12205 , n12206 , n12207 , n12208 , n12209 , n12210 , n12211 , n12212 , n12213 , n12214 , n12215 , n12216 , n12217 , n12218 , n12219 , n12220 , n12221 , n12222 , n12223 , n12224 , n12225 , n12226 , n12227 , n12228 , n12229 , n12230 , n12231 , n12232 , n12233 , n12234 , n12235 , n12236 , n12237 , n12238 , n12239 , n12240 , n12241 , n12242 , n12243 , n12244 , n12245 , n12246 , n12247 , n12248 , n12249 , n12250 , n12251 , n12252 , n12253 , n12254 , n12255 , n12256 , n12257 , n12258 , n12259 , n12260 , n12261 , n12262 , n12263 , n12264 , n12265 , n12266 , n12267 , n12268 , n12269 , n12270 , n12271 , n12272 , n12273 , n12274 , n12275 , n12276 , n12277 , n12278 , n12279 , n12280 , n12281 , n12282 , n12283 , n12284 , n12285 , n12286 , n12287 , n12288 , n12289 , n12290 , n12291 , n12292 , n12293 , n12294 , n12295 , n12296 , n12297 , n12298 , n12299 , n12300 , n12301 , n12302 , n12303 , n12304 , n12305 , n12306 , n12307 , n12308 , n12309 , n12310 , n12311 , n12312 , n12313 , n12314 , n12315 , n12316 , n12317 , n12318 , n12319 , n12320 , n12321 , n12322 , n12323 , n12324 , n12325 , n12326 , n12327 , n12328 , n12329 , n12330 , n12331 , n12332 , n12333 , n12334 , n12335 , n12336 , n12337 , n12338 , n12339 , n12340 , n12341 , n12342 , n12343 , n12344 , n12345 , n12346 , n12347 , n12348 , n12349 , n12350 , n12351 , n12352 , n12353 , n12354 , n12355 , n12356 , n12357 , n12358 , n12359 , n12360 , n12361 , n12362 , n12363 , n12364 , n12365 , n12366 , n12367 , n12368 , n12369 , n12370 , n12371 , n12372 , n12373 , n12374 , n12375 , n12376 , n12377 , n12378 , n12379 , n12380 , n12381 , n12382 , n12383 , n12384 , n12385 , n12386 , n12387 , n12388 , n12389 , n12390 , n12391 , n12392 , n12393 , n12394 , n12395 , n12396 , n12397 , n12398 , n12399 , n12400 , n12401 , n12402 , n12403 , n12404 , n12405 , n12406 , n12407 , n12408 , n12409 , n12410 , n12411 , n12412 , n12413 , n12414 , n12415 , n12416 , n12417 , n12418 , n12419 , n12420 , n12421 , n12422 , n12423 , n12424 , n12425 , n12426 , n12427 , n12428 , n12429 , n12430 , n12431 , n12432 , n12433 , n12434 , n12435 , n12436 , n12437 , n12438 , n12439 , n12440 , n12441 , n12442 , n12443 , n12444 , n12445 , n12446 , n12447 , n12448 , n12449 , n12450 , n12451 , n12452 , n12453 , n12454 , n12455 , n12456 , n12457 , n12458 , n12459 , n12460 , n12461 , n12462 , n12463 , n12464 , n12465 , n12466 , n12467 , n12468 , n12469 , n12470 , n12471 , n12472 , n12473 , n12474 , n12475 , n12476 , n12477 , n12478 , n12479 , n12480 , n12481 , n12482 , n12483 , n12484 , n12485 , n12486 , n12487 , n12488 , n12489 , n12490 , n12491 , n12492 , n12493 , n12494 , n12495 , n12496 , n12497 , n12498 , n12499 , n12500 , n12501 , n12502 , n12503 , n12504 , n12505 , n12506 , n12507 , n12508 , n12509 , n12510 , n12511 , n12512 , n12513 , n12514 , n12515 , n12516 , n12517 , n12518 , n12519 , n12520 , n12521 , n12522 , n12523 , n12524 , n12525 , n12526 , n12527 , n12528 , n12529 , n12530 , n12531 , n12532 , n12533 , n12534 , n12535 , n12536 , n12537 , n12538 , n12539 , n12540 , n12541 , n12542 , n12543 , n12544 , n12545 , n12546 , n12547 , n12548 , n12549 , n12550 , n12551 , n12552 , n12553 , n12554 , n12555 , n12556 , n12557 , n12558 , n12559 , n12560 , n12561 , n12562 , n12563 , n12564 , n12565 , n12566 , n12567 , n12568 , n12569 , n12570 , n12571 , n12572 , n12573 , n12574 , n12575 , n12576 , n12577 , n12578 , n12579 , n12580 , n12581 , n12582 , n12583 , n12584 , n12585 , n12586 , n12587 , n12588 , n12589 , n12590 , n12591 , n12592 , n12593 , n12594 , n12595 , n12596 , n12597 , n12598 , n12599 , n12600 , n12601 , n12602 , n12603 , n12604 , n12605 , n12606 , n12607 , n12608 , n12609 , n12610 , n12611 , n12612 , n12613 , n12614 , n12615 , n12616 , n12617 , n12618 , n12619 , n12620 , n12621 , n12622 , n12623 , n12624 , n12625 , n12626 , n12627 , n12628 , n12629 , n12630 , n12631 , n12632 , n12633 , n12634 , n12635 , n12636 , n12637 , n12638 , n12639 , n12640 , n12641 , n12642 , n12643 , n12644 , n12645 , n12646 , n12647 , n12648 , n12649 , n12650 , n12651 , n12652 , n12653 , n12654 , n12655 , n12656 , n12657 , n12658 , n12659 , n12660 , n12661 , n12662 , n12663 , n12664 , n12665 , n12666 , n12667 , n12668 , n12669 , n12670 , n12671 , n12672 , n12673 , n12674 , n12675 , n12676 , n12677 , n12678 , n12679 , n12680 , n12681 , n12682 , n12683 , n12684 , n12685 , n12686 , n12687 , n12688 , n12689 , n12690 , n12691 , n12692 , n12693 , n12694 , n12695 , n12696 , n12697 , n12698 , n12699 , n12700 , n12701 , n12702 , n12703 , n12704 , n12705 , n12706 , n12707 , n12708 , n12709 , n12710 , n12711 , n12712 , n12713 , n12714 , n12715 , n12716 , n12717 , n12718 , n12719 , n12720 , n12721 , n12722 , n12723 , n12724 , n12725 , n12726 , n12727 , n12728 , n12729 , n12730 , n12731 , n12732 , n12733 , n12734 , n12735 , n12736 , n12737 , n12738 , n12739 , n12740 , n12741 , n12742 , n12743 , n12744 , n12745 , n12746 , n12747 , n12748 , n12749 , n12750 , n12751 , n12752 , n12753 , n12754 , n12755 , n12756 , n12757 , n12758 , n12759 , n12760 , n12761 , n12762 , n12763 , n12764 , n12765 , n12766 , n12767 , n12768 , n12769 , n12770 , n12771 , n12772 , n12773 , n12774 , n12775 , n12776 , n12777 , n12778 , n12779 , n12780 , n12781 , n12782 , n12783 , n12784 , n12785 , n12786 , n12787 , n12788 , n12789 , n12790 , n12791 , n12792 , n12793 , n12794 , n12795 , n12796 , n12797 , n12798 , n12799 , n12800 , n12801 , n12802 , n12803 , n12804 , n12805 , n12806 , n12807 , n12808 , n12809 , n12810 , n12811 , n12812 , n12813 , n12814 , n12815 , n12816 , n12817 , n12818 , n12819 , n12820 , n12821 , n12822 , n12823 , n12824 , n12825 , n12826 , n12827 , n12828 , n12829 , n12830 , n12831 , n12832 , n12833 , n12834 , n12835 , n12836 , n12837 , n12838 , n12839 , n12840 , n12841 , n12842 , n12843 , n12844 , n12845 , n12846 , n12847 , n12848 , n12849 , n12850 , n12851 , n12852 , n12853 , n12854 , n12855 , n12856 , n12857 , n12858 , n12859 , n12860 , n12861 , n12862 , n12863 , n12864 , n12865 , n12866 , n12867 , n12868 , n12869 , n12870 , n12871 , n12872 , n12873 , n12874 , n12875 , n12876 , n12877 , n12878 , n12879 , n12880 , n12881 , n12882 , n12883 , n12884 , n12885 , n12886 , n12887 , n12888 , n12889 , n12890 , n12891 , n12892 , n12893 , n12894 , n12895 , n12896 , n12897 , n12898 , n12899 , n12900 , n12901 , n12902 , n12903 , n12904 , n12905 , n12906 , n12907 , n12908 , n12909 , n12910 , n12911 , n12912 , n12913 , n12914 , n12915 , n12916 , n12917 , n12918 , n12919 , n12920 , n12921 , n12922 , n12923 , n12924 , n12925 , n12926 , n12927 , n12928 , n12929 , n12930 , n12931 , n12932 , n12933 , n12934 , n12935 , n12936 , n12937 , n12938 , n12939 , n12940 , n12941 , n12942 , n12943 , n12944 , n12945 , n12946 , n12947 , n12948 , n12949 , n12950 , n12951 , n12952 , n12953 , n12954 , n12955 , n12956 , n12957 , n12958 , n12959 , n12960 , n12961 , n12962 , n12963 , n12964 , n12965 , n12966 , n12967 , n12968 , n12969 , n12970 , n12971 , n12972 , n12973 , n12974 , n12975 , n12976 , n12977 , n12978 , n12979 , n12980 , n12981 , n12982 , n12983 , n12984 , n12985 , n12986 , n12987 , n12988 , n12989 , n12990 , n12991 , n12992 , n12993 , n12994 , n12995 , n12996 , n12997 , n12998 , n12999 , n13000 , n13001 , n13002 , n13003 , n13004 , n13005 , n13006 , n13007 , n13008 , n13009 , n13010 , n13011 , n13012 , n13013 , n13014 , n13015 , n13016 , n13017 , n13018 , n13019 , n13020 , n13021 , n13022 , n13023 , n13024 , n13025 , n13026 , n13027 , n13028 , n13029 , n13030 , n13031 , n13032 , n13033 , n13034 , n13035 , n13036 , n13037 , n13038 , n13039 , n13040 , n13041 , n13042 , n13043 , n13044 , n13045 , n13046 , n13047 , n13048 , n13049 , n13050 , n13051 , n13052 , n13053 , n13054 , n13055 , n13056 , n13057 , n13058 , n13059 , n13060 , n13061 , n13062 , n13063 , n13064 , n13065 , n13066 , n13067 , n13068 , n13069 , n13070 , n13071 , n13072 , n13073 , n13074 , n13075 , n13076 , n13077 , n13078 , n13079 , n13080 , n13081 , n13082 , n13083 , n13084 , n13085 , n13086 , n13087 , n13088 , n13089 , n13090 , n13091 , n13092 , n13093 , n13094 , n13095 , n13096 , n13097 , n13098 , n13099 , n13100 , n13101 , n13102 , n13103 , n13104 , n13105 , n13106 , n13107 , n13108 , n13109 , n13110 , n13111 , n13112 , n13113 , n13114 , n13115 , n13116 , n13117 , n13118 , n13119 , n13120 , n13121 , n13122 , n13123 , n13124 , n13125 , n13126 , n13127 , n13128 , n13129 , n13130 , n13131 , n13132 , n13133 , n13134 , n13135 , n13136 , n13137 , n13138 , n13139 , n13140 , n13141 , n13142 , n13143 , n13144 , n13145 , n13146 , n13147 , n13148 , n13149 , n13150 , n13151 , n13152 , n13153 , n13154 , n13155 , n13156 , n13157 , n13158 , n13159 , n13160 , n13161 , n13162 , n13163 , n13164 , n13165 , n13166 , n13167 , n13168 , n13169 , n13170 , n13171 , n13172 , n13173 , n13174 , n13175 , n13176 , n13177 , n13178 , n13179 , n13180 , n13181 , n13182 , n13183 , n13184 , n13185 , n13186 , n13187 , n13188 , n13189 , n13190 , n13191 , n13192 , n13193 , n13194 , n13195 , n13196 , n13197 , n13198 , n13199 , n13200 , n13201 , n13202 , n13203 , n13204 , n13205 , n13206 , n13207 , n13208 , n13209 , n13210 , n13211 , n13212 , n13213 , n13214 , n13215 , n13216 , n13217 , n13218 , n13219 , n13220 , n13221 , n13222 , n13223 , n13224 , n13225 , n13226 , n13227 , n13228 , n13229 , n13230 , n13231 , n13232 , n13233 , n13234 , n13235 , n13236 , n13237 , n13238 , n13239 , n13240 , n13241 , n13242 , n13243 , n13244 , n13245 , n13246 , n13247 , n13248 , n13249 , n13250 , n13251 , n13252 , n13253 , n13254 , n13255 , n13256 , n13257 , n13258 , n13259 , n13260 , n13261 , n13262 , n13263 , n13264 , n13265 , n13266 , n13267 , n13268 , n13269 , n13270 , n13271 , n13272 , n13273 , n13274 , n13275 , n13276 , n13277 , n13278 , n13279 , n13280 , n13281 , n13282 , n13283 , n13284 , n13285 , n13286 , n13287 , n13288 , n13289 , n13290 , n13291 , n13292 , n13293 , n13294 , n13295 , n13296 , n13297 , n13298 , n13299 , n13300 , n13301 , n13302 , n13303 , n13304 , n13305 , n13306 , n13307 , n13308 , n13309 , n13310 , n13311 , n13312 , n13313 , n13314 , n13315 , n13316 , n13317 , n13318 , n13319 , n13320 , n13321 , n13322 , n13323 , n13324 , n13325 , n13326 , n13327 , n13328 , n13329 , n13330 , n13331 , n13332 , n13333 , n13334 , n13335 , n13336 , n13337 , n13338 , n13339 , n13340 , n13341 , n13342 , n13343 , n13344 , n13345 , n13346 , n13347 , n13348 , n13349 , n13350 , n13351 , n13352 , n13353 , n13354 , n13355 , n13356 , n13357 , n13358 , n13359 , n13360 , n13361 , n13362 , n13363 , n13364 , n13365 , n13366 , n13367 , n13368 , n13369 , n13370 , n13371 , n13372 , n13373 , n13374 , n13375 , n13376 , n13377 , n13378 , n13379 , n13380 , n13381 , n13382 , n13383 , n13384 , n13385 , n13386 , n13387 , n13388 , n13389 , n13390 , n13391 , n13392 , n13393 , n13394 , n13395 , n13396 , n13397 , n13398 , n13399 , n13400 , n13401 , n13402 , n13403 , n13404 , n13405 , n13406 , n13407 , n13408 , n13409 , n13410 , n13411 , n13412 , n13413 , n13414 , n13415 , n13416 , n13417 , n13418 , n13419 , n13420 , n13421 , n13422 , n13423 , n13424 , n13425 , n13426 , n13427 , n13428 , n13429 , n13430 , n13431 , n13432 , n13433 , n13434 , n13435 , n13436 , n13437 , n13438 , n13439 , n13440 , n13441 , n13442 , n13443 , n13444 , n13445 , n13446 , n13447 , n13448 , n13449 , n13450 , n13451 , n13452 , n13453 , n13454 , n13455 , n13456 , n13457 , n13458 , n13459 , n13460 , n13461 , n13462 , n13463 , n13464 , n13465 , n13466 , n13467 , n13468 , n13469 , n13470 , n13471 , n13472 , n13473 , n13474 , n13475 , n13476 , n13477 , n13478 , n13479 , n13480 , n13481 , n13482 , n13483 , n13484 , n13485 , n13486 , n13487 , n13488 , n13489 , n13490 , n13491 , n13492 , n13493 , n13494 , n13495 , n13496 , n13497 , n13498 , n13499 , n13500 , n13501 , n13502 , n13503 , n13504 , n13505 , n13506 , n13507 , n13508 , n13509 , n13510 , n13511 , n13512 , n13513 , n13514 , n13515 , n13516 , n13517 , n13518 , n13519 , n13520 , n13521 , n13522 , n13523 , n13524 , n13525 , n13526 , n13527 , n13528 , n13529 , n13530 , n13531 , n13532 , n13533 , n13534 , n13535 , n13536 , n13537 , n13538 , n13539 , n13540 , n13541 , n13542 , n13543 , n13544 , n13545 , n13546 , n13547 , n13548 , n13549 , n13550 , n13551 , n13552 , n13553 , n13554 , n13555 , n13556 , n13557 , n13558 , n13559 , n13560 , n13561 , n13562 , n13563 , n13564 , n13565 , n13566 , n13567 , n13568 , n13569 , n13570 , n13571 , n13572 , n13573 , n13574 , n13575 , n13576 , n13577 , n13578 , n13579 , n13580 , n13581 , n13582 , n13583 , n13584 , n13585 , n13586 , n13587 , n13588 , n13589 , n13590 , n13591 , n13592 , n13593 , n13594 , n13595 , n13596 , n13597 , n13598 , n13599 , n13600 , n13601 , n13602 , n13603 , n13604 , n13605 , n13606 , n13607 , n13608 , n13609 , n13610 , n13611 , n13612 , n13613 , n13614 , n13615 , n13616 , n13617 , n13618 , n13619 , n13620 , n13621 , n13622 , n13623 , n13624 , n13625 , n13626 , n13627 , n13628 , n13629 , n13630 , n13631 , n13632 , n13633 , n13634 , n13635 , n13636 , n13637 , n13638 , n13639 , n13640 , n13641 , n13642 , n13643 , n13644 , n13645 , n13646 , n13647 , n13648 , n13649 , n13650 , n13651 , n13652 , n13653 , n13654 , n13655 , n13656 , n13657 , n13658 , n13659 , n13660 , n13661 , n13662 , n13663 , n13664 , n13665 , n13666 , n13667 , n13668 , n13669 , n13670 , n13671 , n13672 , n13673 , n13674 , n13675 , n13676 , n13677 , n13678 , n13679 , n13680 , n13681 , n13682 , n13683 , n13684 , n13685 , n13686 , n13687 , n13688 , n13689 , n13690 , n13691 , n13692 , n13693 , n13694 , n13695 , n13696 , n13697 , n13698 , n13699 , n13700 , n13701 , n13702 , n13703 , n13704 , n13705 , n13706 , n13707 , n13708 , n13709 , n13710 , n13711 , n13712 , n13713 , n13714 , n13715 , n13716 , n13717 , n13718 , n13719 , n13720 , n13721 , n13722 , n13723 , n13724 , n13725 , n13726 , n13727 , n13728 , n13729 , n13730 , n13731 , n13732 , n13733 , n13734 , n13735 , n13736 , n13737 , n13738 , n13739 , n13740 , n13741 , n13742 , n13743 , n13744 , n13745 , n13746 , n13747 , n13748 , n13749 , n13750 , n13751 , n13752 , n13753 , n13754 , n13755 , n13756 , n13757 , n13758 , n13759 , n13760 , n13761 , n13762 , n13763 , n13764 , n13765 , n13766 , n13767 , n13768 , n13769 , n13770 , n13771 , n13772 , n13773 , n13774 , n13775 , n13776 , n13777 , n13778 , n13779 , n13780 , n13781 , n13782 , n13783 , n13784 , n13785 , n13786 , n13787 , n13788 , n13789 , n13790 , n13791 , n13792 , n13793 , n13794 , n13795 , n13796 , n13797 , n13798 , n13799 , n13800 , n13801 , n13802 , n13803 , n13804 , n13805 , n13806 , n13807 , n13808 , n13809 , n13810 , n13811 , n13812 , n13813 , n13814 , n13815 , n13816 , n13817 , n13818 , n13819 , n13820 , n13821 , n13822 , n13823 , n13824 , n13825 , n13826 , n13827 , n13828 , n13829 , n13830 , n13831 , n13832 , n13833 , n13834 , n13835 , n13836 , n13837 , n13838 , n13839 , n13840 , n13841 , n13842 , n13843 , n13844 , n13845 , n13846 , n13847 , n13848 , n13849 , n13850 , n13851 , n13852 , n13853 , n13854 , n13855 , n13856 , n13857 , n13858 , n13859 , n13860 , n13861 , n13862 , n13863 , n13864 , n13865 , n13866 , n13867 , n13868 , n13869 , n13870 , n13871 , n13872 , n13873 , n13874 , n13875 , n13876 , n13877 , n13878 , n13879 , n13880 , n13881 , n13882 , n13883 , n13884 , n13885 , n13886 , n13887 , n13888 , n13889 , n13890 , n13891 , n13892 , n13893 , n13894 , n13895 , n13896 , n13897 , n13898 , n13899 , n13900 , n13901 , n13902 , n13903 , n13904 , n13905 , n13906 , n13907 , n13908 , n13909 , n13910 , n13911 , n13912 , n13913 , n13914 , n13915 , n13916 , n13917 , n13918 , n13919 , n13920 , n13921 , n13922 , n13923 , n13924 , n13925 , n13926 , n13927 , n13928 , n13929 , n13930 , n13931 , n13932 , n13933 , n13934 , n13935 , n13936 , n13937 , n13938 , n13939 , n13940 , n13941 , n13942 , n13943 , n13944 , n13945 , n13946 , n13947 , n13948 , n13949 , n13950 , n13951 , n13952 , n13953 , n13954 , n13955 , n13956 , n13957 , n13958 , n13959 , n13960 , n13961 , n13962 , n13963 , n13964 , n13965 , n13966 , n13967 , n13968 , n13969 , n13970 , n13971 , n13972 , n13973 , n13974 , n13975 , n13976 , n13977 , n13978 , n13979 , n13980 , n13981 , n13982 , n13983 , n13984 , n13985 , n13986 , n13987 , n13988 , n13989 , n13990 , n13991 , n13992 , n13993 , n13994 , n13995 , n13996 , n13997 , n13998 , n13999 , n14000 , n14001 , n14002 , n14003 , n14004 , n14005 , n14006 , n14007 , n14008 , n14009 , n14010 , n14011 , n14012 , n14013 , n14014 , n14015 , n14016 , n14017 , n14018 , n14019 , n14020 , n14021 , n14022 , n14023 , n14024 , n14025 , n14026 , n14027 , n14028 , n14029 , n14030 , n14031 , n14032 , n14033 , n14034 , n14035 , n14036 , n14037 , n14038 , n14039 , n14040 , n14041 , n14042 , n14043 , n14044 , n14045 , n14046 , n14047 , n14048 , n14049 , n14050 , n14051 , n14052 , n14053 , n14054 , n14055 , n14056 , n14057 , n14058 , n14059 , n14060 , n14061 , n14062 , n14063 , n14064 , n14065 , n14066 , n14067 , n14068 , n14069 , n14070 , n14071 , n14072 , n14073 , n14074 , n14075 , n14076 , n14077 , n14078 , n14079 , n14080 , n14081 , n14082 , n14083 , n14084 , n14085 , n14086 , n14087 , n14088 , n14089 , n14090 , n14091 , n14092 , n14093 , n14094 , n14095 , n14096 , n14097 , n14098 , n14099 , n14100 , n14101 , n14102 , n14103 , n14104 , n14105 , n14106 , n14107 , n14108 , n14109 , n14110 , n14111 , n14112 , n14113 , n14114 , n14115 , n14116 , n14117 , n14118 , n14119 , n14120 , n14121 , n14122 , n14123 , n14124 , n14125 , n14126 , n14127 , n14128 , n14129 , n14130 , n14131 , n14132 , n14133 , n14134 , n14135 , n14136 , n14137 , n14138 , n14139 , n14140 , n14141 , n14142 , n14143 , n14144 , n14145 , n14146 , n14147 , n14148 , n14149 , n14150 , n14151 , n14152 , n14153 , n14154 , n14155 , n14156 , n14157 , n14158 , n14159 , n14160 , n14161 , n14162 , n14163 , n14164 , n14165 , n14166 , n14167 , n14168 , n14169 , n14170 , n14171 , n14172 , n14173 , n14174 , n14175 , n14176 , n14177 , n14178 , n14179 , n14180 , n14181 , n14182 , n14183 , n14184 , n14185 , n14186 , n14187 , n14188 , n14189 , n14190 , n14191 , n14192 , n14193 , n14194 , n14195 , n14196 , n14197 , n14198 , n14199 , n14200 , n14201 , n14202 , n14203 , n14204 , n14205 , n14206 , n14207 , n14208 , n14209 , n14210 , n14211 , n14212 , n14213 , n14214 , n14215 , n14216 , n14217 , n14218 , n14219 , n14220 , n14221 , n14222 , n14223 , n14224 , n14225 , n14226 , n14227 , n14228 , n14229 , n14230 , n14231 , n14232 , n14233 , n14234 , n14235 , n14236 , n14237 , n14238 , n14239 , n14240 , n14241 , n14242 , n14243 , n14244 , n14245 , n14246 , n14247 , n14248 , n14249 , n14250 , n14251 , n14252 , n14253 , n14254 , n14255 , n14256 , n14257 , n14258 , n14259 , n14260 , n14261 , n14262 , n14263 , n14264 , n14265 , n14266 , n14267 , n14268 , n14269 , n14270 , n14271 , n14272 , n14273 , n14274 , n14275 , n14276 , n14277 , n14278 , n14279 , n14280 , n14281 , n14282 , n14283 , n14284 , n14285 , n14286 , n14287 , n14288 , n14289 , n14290 , n14291 , n14292 , n14293 , n14294 , n14295 , n14296 , n14297 , n14298 , n14299 , n14300 , n14301 , n14302 , n14303 , n14304 , n14305 , n14306 , n14307 , n14308 , n14309 , n14310 , n14311 , n14312 , n14313 , n14314 , n14315 , n14316 , n14317 , n14318 , n14319 , n14320 , n14321 , n14322 , n14323 , n14324 , n14325 , n14326 , n14327 , n14328 , n14329 , n14330 , n14331 , n14332 , n14333 , n14334 , n14335 , n14336 , n14337 , n14338 , n14339 , n14340 , n14341 , n14342 , n14343 , n14344 , n14345 , n14346 , n14347 , n14348 , n14349 , n14350 , n14351 , n14352 , n14353 , n14354 , n14355 , n14356 , n14357 , n14358 , n14359 , n14360 , n14361 , n14362 , n14363 , n14364 , n14365 , n14366 , n14367 , n14368 , n14369 , n14370 , n14371 , n14372 , n14373 , n14374 , n14375 , n14376 , n14377 , n14378 , n14379 , n14380 , n14381 , n14382 , n14383 , n14384 , n14385 , n14386 , n14387 , n14388 , n14389 , n14390 , n14391 , n14392 , n14393 , n14394 , n14395 , n14396 , n14397 , n14398 , n14399 , n14400 , n14401 , n14402 , n14403 , n14404 , n14405 , n14406 , n14407 , n14408 , n14409 , n14410 , n14411 , n14412 , n14413 , n14414 , n14415 , n14416 , n14417 , n14418 , n14419 , n14420 , n14421 , n14422 , n14423 , n14424 , n14425 , n14426 , n14427 , n14428 , n14429 , n14430 , n14431 , n14432 , n14433 , n14434 , n14435 , n14436 , n14437 , n14438 , n14439 , n14440 , n14441 , n14442 , n14443 , n14444 , n14445 , n14446 , n14447 , n14448 , n14449 , n14450 , n14451 , n14452 , n14453 , n14454 , n14455 , n14456 , n14457 , n14458 , n14459 , n14460 , n14461 , n14462 , n14463 , n14464 , n14465 , n14466 , n14467 , n14468 , n14469 , n14470 , n14471 , n14472 , n14473 , n14474 , n14475 , n14476 , n14477 , n14478 , n14479 , n14480 , n14481 , n14482 , n14483 , n14484 , n14485 , n14486 , n14487 , n14488 , n14489 , n14490 , n14491 , n14492 , n14493 , n14494 , n14495 , n14496 , n14497 , n14498 , n14499 , n14500 , n14501 , n14502 , n14503 , n14504 , n14505 , n14506 , n14507 , n14508 , n14509 , n14510 , n14511 , n14512 , n14513 , n14514 , n14515 , n14516 , n14517 , n14518 , n14519 , n14520 , n14521 , n14522 , n14523 , n14524 , n14525 , n14526 , n14527 , n14528 , n14529 , n14530 , n14531 , n14532 , n14533 , n14534 , n14535 , n14536 , n14537 , n14538 , n14539 , n14540 , n14541 , n14542 , n14543 , n14544 , n14545 , n14546 , n14547 , n14548 , n14549 , n14550 , n14551 , n14552 , n14553 , n14554 , n14555 , n14556 , n14557 , n14558 , n14559 , n14560 , n14561 , n14562 , n14563 , n14564 , n14565 , n14566 , n14567 , n14568 , n14569 , n14570 , n14571 , n14572 , n14573 , n14574 , n14575 , n14576 , n14577 , n14578 , n14579 , n14580 , n14581 , n14582 , n14583 , n14584 , n14585 , n14586 , n14587 , n14588 , n14589 , n14590 , n14591 , n14592 , n14593 , n14594 , n14595 , n14596 , n14597 , n14598 , n14599 , n14600 , n14601 , n14602 , n14603 , n14604 , n14605 , n14606 , n14607 , n14608 , n14609 , n14610 , n14611 , n14612 , n14613 , n14614 , n14615 , n14616 , n14617 , n14618 , n14619 , n14620 , n14621 , n14622 , n14623 , n14624 , n14625 , n14626 , n14627 , n14628 , n14629 , n14630 , n14631 , n14632 , n14633 , n14634 , n14635 , n14636 , n14637 , n14638 , n14639 , n14640 , n14641 , n14642 , n14643 , n14644 , n14645 , n14646 , n14647 , n14648 , n14649 , n14650 , n14651 , n14652 , n14653 , n14654 , n14655 , n14656 , n14657 , n14658 , n14659 , n14660 , n14661 , n14662 , n14663 , n14664 , n14665 , n14666 , n14667 , n14668 , n14669 , n14670 , n14671 , n14672 , n14673 , n14674 , n14675 , n14676 , n14677 , n14678 , n14679 , n14680 , n14681 , n14682 , n14683 , n14684 , n14685 , n14686 , n14687 , n14688 , n14689 , n14690 , n14691 , n14692 , n14693 , n14694 , n14695 , n14696 , n14697 , n14698 , n14699 , n14700 , n14701 , n14702 , n14703 , n14704 , n14705 , n14706 , n14707 , n14708 , n14709 , n14710 , n14711 , n14712 , n14713 , n14714 , n14715 , n14716 , n14717 , n14718 , n14719 , n14720 , n14721 , n14722 , n14723 , n14724 , n14725 , n14726 , n14727 , n14728 , n14729 , n14730 , n14731 , n14732 , n14733 , n14734 , n14735 , n14736 , n14737 , n14738 , n14739 , n14740 , n14741 , n14742 , n14743 , n14744 , n14745 , n14746 , n14747 , n14748 , n14749 , n14750 , n14751 , n14752 , n14753 , n14754 , n14755 , n14756 , n14757 , n14758 , n14759 , n14760 , n14761 , n14762 , n14763 , n14764 , n14765 , n14766 , n14767 , n14768 , n14769 , n14770 , n14771 , n14772 , n14773 , n14774 , n14775 , n14776 , n14777 , n14778 , n14779 , n14780 , n14781 , n14782 , n14783 , n14784 , n14785 , n14786 , n14787 , n14788 , n14789 , n14790 , n14791 , n14792 , n14793 , n14794 , n14795 , n14796 , n14797 , n14798 , n14799 , n14800 , n14801 , n14802 , n14803 , n14804 , n14805 , n14806 , n14807 , n14808 , n14809 , n14810 , n14811 , n14812 , n14813 , n14814 , n14815 , n14816 , n14817 , n14818 , n14819 , n14820 , n14821 , n14822 , n14823 , n14824 , n14825 , n14826 , n14827 , n14828 , n14829 , n14830 , n14831 , n14832 , n14833 , n14834 , n14835 , n14836 , n14837 , n14838 , n14839 , n14840 , n14841 , n14842 , n14843 , n14844 , n14845 , n14846 , n14847 , n14848 , n14849 , n14850 , n14851 , n14852 , n14853 , n14854 , n14855 , n14856 , n14857 , n14858 , n14859 , n14860 , n14861 , n14862 , n14863 , n14864 , n14865 , n14866 , n14867 , n14868 , n14869 , n14870 , n14871 , n14872 , n14873 , n14874 , n14875 , n14876 , n14877 , n14878 , n14879 , n14880 , n14881 , n14882 , n14883 , n14884 , n14885 , n14886 , n14887 , n14888 , n14889 , n14890 , n14891 , n14892 , n14893 , n14894 , n14895 , n14896 , n14897 , n14898 , n14899 , n14900 , n14901 , n14902 , n14903 , n14904 , n14905 , n14906 , n14907 , n14908 , n14909 , n14910 , n14911 , n14912 , n14913 , n14914 , n14915 , n14916 , n14917 , n14918 , n14919 , n14920 , n14921 , n14922 , n14923 , n14924 , n14925 , n14926 , n14927 , n14928 , n14929 , n14930 , n14931 , n14932 , n14933 , n14934 , n14935 , n14936 , n14937 , n14938 , n14939 , n14940 , n14941 , n14942 , n14943 , n14944 , n14945 , n14946 , n14947 , n14948 , n14949 , n14950 , n14951 , n14952 , n14953 , n14954 , n14955 , n14956 , n14957 , n14958 , n14959 , n14960 , n14961 , n14962 , n14963 , n14964 , n14965 , n14966 , n14967 , n14968 , n14969 , n14970 , n14971 , n14972 , n14973 , n14974 , n14975 , n14976 , n14977 , n14978 , n14979 , n14980 , n14981 , n14982 , n14983 , n14984 , n14985 , n14986 , n14987 , n14988 , n14989 , n14990 , n14991 , n14992 , n14993 , n14994 , n14995 , n14996 , n14997 , n14998 , n14999 , n15000 , n15001 , n15002 , n15003 , n15004 , n15005 , n15006 , n15007 , n15008 , n15009 , n15010 , n15011 , n15012 , n15013 , n15014 , n15015 , n15016 , n15017 , n15018 , n15019 , n15020 , n15021 , n15022 , n15023 , n15024 , n15025 , n15026 , n15027 , n15028 , n15029 , n15030 , n15031 , n15032 , n15033 , n15034 , n15035 , n15036 , n15037 , n15038 , n15039 , n15040 , n15041 , n15042 , n15043 , n15044 , n15045 , n15046 , n15047 , n15048 , n15049 , n15050 , n15051 , n15052 , n15053 , n15054 , n15055 , n15056 , n15057 , n15058 , n15059 , n15060 , n15061 , n15062 , n15063 , n15064 , n15065 , n15066 , n15067 , n15068 , n15069 , n15070 , n15071 , n15072 , n15073 , n15074 , n15075 , n15076 , n15077 , n15078 , n15079 , n15080 , n15081 , n15082 , n15083 , n15084 , n15085 , n15086 , n15087 , n15088 , n15089 , n15090 , n15091 , n15092 , n15093 , n15094 , n15095 , n15096 , n15097 , n15098 , n15099 , n15100 , n15101 , n15102 , n15103 , n15104 , n15105 , n15106 , n15107 , n15108 , n15109 , n15110 , n15111 , n15112 , n15113 , n15114 , n15115 , n15116 , n15117 , n15118 , n15119 , n15120 , n15121 , n15122 , n15123 , n15124 , n15125 , n15126 , n15127 , n15128 , n15129 , n15130 , n15131 , n15132 , n15133 , n15134 , n15135 , n15136 , n15137 , n15138 , n15139 , n15140 , n15141 , n15142 , n15143 , n15144 , n15145 , n15146 , n15147 , n15148 , n15149 , n15150 , n15151 , n15152 , n15153 , n15154 , n15155 , n15156 , n15157 , n15158 , n15159 , n15160 , n15161 , n15162 , n15163 , n15164 , n15165 , n15166 , n15167 , n15168 , n15169 , n15170 , n15171 , n15172 , n15173 , n15174 , n15175 , n15176 , n15177 , n15178 , n15179 , n15180 , n15181 , n15182 , n15183 , n15184 , n15185 , n15186 , n15187 , n15188 , n15189 , n15190 , n15191 , n15192 , n15193 , n15194 , n15195 , n15196 , n15197 , n15198 , n15199 , n15200 , n15201 , n15202 , n15203 , n15204 , n15205 , n15206 , n15207 , n15208 , n15209 , n15210 , n15211 , n15212 , n15213 , n15214 , n15215 , n15216 , n15217 , n15218 , n15219 , n15220 , n15221 , n15222 , n15223 , n15224 , n15225 , n15226 , n15227 , n15228 , n15229 , n15230 , n15231 , n15232 , n15233 , n15234 , n15235 , n15236 , n15237 , n15238 , n15239 , n15240 , n15241 , n15242 , n15243 , n15244 , n15245 , n15246 , n15247 , n15248 , n15249 , n15250 , n15251 , n15252 , n15253 , n15254 , n15255 , n15256 , n15257 , n15258 , n15259 , n15260 , n15261 , n15262 , n15263 , n15264 , n15265 , n15266 , n15267 , n15268 , n15269 , n15270 , n15271 , n15272 , n15273 , n15274 , n15275 , n15276 , n15277 , n15278 , n15279 , n15280 , n15281 , n15282 , n15283 , n15284 , n15285 , n15286 , n15287 , n15288 , n15289 , n15290 , n15291 , n15292 , n15293 , n15294 , n15295 , n15296 , n15297 , n15298 , n15299 , n15300 , n15301 , n15302 , n15303 , n15304 , n15305 , n15306 , n15307 , n15308 , n15309 , n15310 , n15311 , n15312 , n15313 , n15314 , n15315 , n15316 , n15317 , n15318 , n15319 , n15320 , n15321 , n15322 , n15323 , n15324 , n15325 , n15326 , n15327 , n15328 , n15329 , n15330 , n15331 , n15332 , n15333 , n15334 , n15335 , n15336 , n15337 , n15338 , n15339 , n15340 , n15341 , n15342 , n15343 , n15344 , n15345 , n15346 , n15347 , n15348 , n15349 , n15350 , n15351 , n15352 , n15353 , n15354 , n15355 , n15356 , n15357 , n15358 , n15359 , n15360 , n15361 , n15362 , n15363 , n15364 , n15365 , n15366 , n15367 , n15368 , n15369 , n15370 , n15371 , n15372 , n15373 , n15374 , n15375 , n15376 , n15377 , n15378 , n15379 , n15380 , n15381 , n15382 , n15383 , n15384 , n15385 , n15386 , n15387 , n15388 , n15389 , n15390 , n15391 , n15392 , n15393 , n15394 , n15395 , n15396 , n15397 , n15398 , n15399 , n15400 , n15401 , n15402 , n15403 , n15404 , n15405 , n15406 , n15407 , n15408 , n15409 , n15410 , n15411 , n15412 , n15413 , n15414 , n15415 , n15416 , n15417 , n15418 , n15419 , n15420 , n15421 , n15422 , n15423 , n15424 , n15425 , n15426 , n15427 , n15428 , n15429 , n15430 , n15431 , n15432 , n15433 , n15434 , n15435 , n15436 , n15437 , n15438 , n15439 , n15440 , n15441 , n15442 , n15443 , n15444 , n15445 , n15446 , n15447 , n15448 , n15449 , n15450 , n15451 , n15452 , n15453 , n15454 , n15455 , n15456 , n15457 , n15458 , n15459 , n15460 , n15461 , n15462 , n15463 , n15464 , n15465 , n15466 , n15467 , n15468 , n15469 , n15470 , n15471 , n15472 , n15473 , n15474 , n15475 , n15476 , n15477 , n15478 , n15479 , n15480 , n15481 , n15482 , n15483 , n15484 , n15485 , n15486 , n15487 , n15488 , n15489 , n15490 , n15491 , n15492 , n15493 , n15494 , n15495 , n15496 , n15497 , n15498 , n15499 , n15500 , n15501 , n15502 , n15503 , n15504 , n15505 , n15506 , n15507 , n15508 , n15509 , n15510 , n15511 , n15512 , n15513 , n15514 , n15515 , n15516 , n15517 , n15518 , n15519 , n15520 , n15521 , n15522 , n15523 , n15524 , n15525 , n15526 , n15527 , n15528 , n15529 , n15530 , n15531 , n15532 , n15533 , n15534 , n15535 , n15536 , n15537 , n15538 , n15539 , n15540 , n15541 , n15542 , n15543 , n15544 , n15545 , n15546 , n15547 , n15548 , n15549 , n15550 , n15551 , n15552 , n15553 , n15554 , n15555 , n15556 , n15557 , n15558 , n15559 , n15560 , n15561 , n15562 , n15563 , n15564 , n15565 , n15566 , n15567 , n15568 , n15569 , n15570 , n15571 , n15572 , n15573 , n15574 , n15575 , n15576 , n15577 , n15578 , n15579 , n15580 , n15581 , n15582 , n15583 , n15584 , n15585 , n15586 , n15587 , n15588 , n15589 , n15590 , n15591 , n15592 , n15593 , n15594 , n15595 , n15596 , n15597 , n15598 , n15599 , n15600 , n15601 , n15602 , n15603 , n15604 , n15605 , n15606 , n15607 , n15608 , n15609 , n15610 , n15611 , n15612 , n15613 , n15614 , n15615 , n15616 , n15617 , n15618 , n15619 , n15620 , n15621 , n15622 , n15623 , n15624 , n15625 , n15626 , n15627 , n15628 , n15629 , n15630 , n15631 , n15632 , n15633 , n15634 , n15635 , n15636 , n15637 , n15638 , n15639 , n15640 , n15641 , n15642 , n15643 , n15644 , n15645 , n15646 , n15647 , n15648 , n15649 , n15650 , n15651 , n15652 , n15653 , n15654 , n15655 , n15656 , n15657 , n15658 , n15659 , n15660 , n15661 , n15662 , n15663 , n15664 , n15665 , n15666 , n15667 , n15668 , n15669 , n15670 , n15671 , n15672 , n15673 , n15674 , n15675 , n15676 , n15677 , n15678 , n15679 , n15680 , n15681 , n15682 , n15683 , n15684 , n15685 , n15686 , n15687 , n15688 , n15689 , n15690 , n15691 , n15692 , n15693 , n15694 , n15695 , n15696 , n15697 , n15698 , n15699 , n15700 , n15701 , n15702 , n15703 , n15704 , n15705 , n15706 , n15707 , n15708 , n15709 , n15710 , n15711 , n15712 , n15713 , n15714 , n15715 , n15716 , n15717 , n15718 , n15719 , n15720 , n15721 , n15722 , n15723 , n15724 , n15725 , n15726 , n15727 , n15728 , n15729 , n15730 , n15731 , n15732 , n15733 , n15734 , n15735 , n15736 , n15737 , n15738 , n15739 , n15740 , n15741 , n15742 , n15743 , n15744 , n15745 , n15746 , n15747 , n15748 , n15749 , n15750 , n15751 , n15752 , n15753 , n15754 , n15755 , n15756 , n15757 , n15758 , n15759 , n15760 , n15761 , n15762 , n15763 , n15764 , n15765 , n15766 , n15767 , n15768 , n15769 , n15770 , n15771 , n15772 , n15773 , n15774 , n15775 , n15776 , n15777 , n15778 , n15779 , n15780 , n15781 , n15782 , n15783 , n15784 , n15785 , n15786 , n15787 , n15788 , n15789 , n15790 , n15791 , n15792 , n15793 , n15794 , n15795 , n15796 , n15797 , n15798 , n15799 , n15800 , n15801 , n15802 , n15803 , n15804 , n15805 , n15806 , n15807 , n15808 , n15809 , n15810 , n15811 , n15812 , n15813 , n15814 , n15815 , n15816 , n15817 , n15818 , n15819 , n15820 , n15821 , n15822 , n15823 , n15824 , n15825 , n15826 , n15827 , n15828 , n15829 , n15830 , n15831 , n15832 , n15833 , n15834 , n15835 , n15836 , n15837 , n15838 , n15839 , n15840 , n15841 , n15842 , n15843 , n15844 , n15845 , n15846 , n15847 , n15848 , n15849 , n15850 , n15851 , n15852 , n15853 , n15854 , n15855 , n15856 , n15857 , n15858 , n15859 , n15860 , n15861 , n15862 , n15863 , n15864 , n15865 , n15866 , n15867 , n15868 , n15869 , n15870 , n15871 , n15872 , n15873 , n15874 , n15875 , n15876 , n15877 , n15878 , n15879 , n15880 , n15881 , n15882 , n15883 , n15884 , n15885 , n15886 , n15887 , n15888 , n15889 , n15890 , n15891 , n15892 , n15893 , n15894 , n15895 , n15896 , n15897 , n15898 , n15899 , n15900 , n15901 , n15902 , n15903 , n15904 , n15905 , n15906 , n15907 , n15908 , n15909 , n15910 , n15911 , n15912 , n15913 , n15914 , n15915 , n15916 , n15917 , n15918 , n15919 , n15920 , n15921 , n15922 , n15923 , n15924 , n15925 , n15926 , n15927 , n15928 , n15929 , n15930 , n15931 , n15932 , n15933 , n15934 , n15935 , n15936 , n15937 , n15938 , n15939 , n15940 , n15941 , n15942 , n15943 , n15944 , n15945 , n15946 , n15947 , n15948 , n15949 , n15950 , n15951 , n15952 , n15953 , n15954 , n15955 , n15956 , n15957 , n15958 , n15959 , n15960 , n15961 , n15962 , n15963 , n15964 , n15965 , n15966 , n15967 , n15968 , n15969 , n15970 , n15971 , n15972 , n15973 , n15974 , n15975 , n15976 , n15977 , n15978 , n15979 , n15980 , n15981 , n15982 , n15983 , n15984 , n15985 , n15986 , n15987 , n15988 , n15989 , n15990 , n15991 , n15992 , n15993 , n15994 , n15995 , n15996 , n15997 , n15998 , n15999 , n16000 , n16001 , n16002 , n16003 , n16004 , n16005 , n16006 , n16007 , n16008 , n16009 , n16010 , n16011 , n16012 , n16013 , n16014 , n16015 , n16016 , n16017 , n16018 , n16019 , n16020 , n16021 , n16022 , n16023 , n16024 , n16025 , n16026 , n16027 , n16028 , n16029 , n16030 , n16031 , n16032 , n16033 , n16034 , n16035 , n16036 , n16037 , n16038 , n16039 , n16040 , n16041 , n16042 , n16043 , n16044 , n16045 , n16046 , n16047 , n16048 , n16049 , n16050 , n16051 , n16052 , n16053 , n16054 , n16055 , n16056 , n16057 , n16058 , n16059 , n16060 , n16061 , n16062 , n16063 , n16064 , n16065 , n16066 , n16067 , n16068 , n16069 , n16070 , n16071 , n16072 , n16073 , n16074 , n16075 , n16076 , n16077 , n16078 , n16079 , n16080 , n16081 , n16082 , n16083 , n16084 , n16085 , n16086 , n16087 , n16088 , n16089 , n16090 , n16091 , n16092 , n16093 , n16094 , n16095 , n16096 , n16097 , n16098 , n16099 , n16100 , n16101 , n16102 , n16103 , n16104 , n16105 , n16106 , n16107 , n16108 , n16109 , n16110 , n16111 , n16112 , n16113 , n16114 , n16115 , n16116 , n16117 , n16118 , n16119 , n16120 , n16121 , n16122 , n16123 , n16124 , n16125 , n16126 , n16127 , n16128 , n16129 , n16130 , n16131 , n16132 , n16133 , n16134 , n16135 , n16136 , n16137 , n16138 , n16139 , n16140 , n16141 , n16142 , n16143 , n16144 , n16145 , n16146 , n16147 , n16148 , n16149 , n16150 , n16151 , n16152 , n16153 , n16154 , n16155 , n16156 , n16157 , n16158 , n16159 , n16160 , n16161 , n16162 , n16163 , n16164 , n16165 , n16166 , n16167 , n16168 , n16169 , n16170 , n16171 , n16172 , n16173 , n16174 , n16175 , n16176 , n16177 , n16178 , n16179 , n16180 , n16181 , n16182 , n16183 , n16184 , n16185 , n16186 , n16187 , n16188 , n16189 , n16190 , n16191 , n16192 , n16193 , n16194 , n16195 , n16196 , n16197 , n16198 , n16199 , n16200 , n16201 , n16202 , n16203 , n16204 , n16205 , n16206 , n16207 , n16208 , n16209 , n16210 , n16211 , n16212 , n16213 , n16214 , n16215 , n16216 , n16217 , n16218 , n16219 , n16220 , n16221 , n16222 , n16223 , n16224 , n16225 , n16226 , n16227 , n16228 , n16229 , n16230 , n16231 , n16232 , n16233 , n16234 , n16235 , n16236 , n16237 , n16238 , n16239 , n16240 , n16241 , n16242 , n16243 , n16244 , n16245 , n16246 , n16247 , n16248 , n16249 , n16250 , n16251 , n16252 , n16253 , n16254 , n16255 , n16256 , n16257 , n16258 , n16259 , n16260 , n16261 , n16262 , n16263 , n16264 , n16265 , n16266 , n16267 , n16268 , n16269 , n16270 , n16271 , n16272 , n16273 , n16274 , n16275 , n16276 , n16277 , n16278 , n16279 , n16280 , n16281 , n16282 , n16283 , n16284 , n16285 , n16286 , n16287 , n16288 , n16289 , n16290 , n16291 , n16292 , n16293 , n16294 , n16295 , n16296 , n16297 , n16298 , n16299 , n16300 , n16301 , n16302 , n16303 , n16304 , n16305 , n16306 , n16307 , n16308 , n16309 , n16310 , n16311 , n16312 , n16313 , n16314 , n16315 , n16316 , n16317 , n16318 , n16319 , n16320 , n16321 , n16322 , n16323 , n16324 , n16325 , n16326 , n16327 , n16328 , n16329 , n16330 , n16331 , n16332 , n16333 , n16334 , n16335 , n16336 , n16337 , n16338 , n16339 , n16340 , n16341 , n16342 , n16343 , n16344 , n16345 , n16346 , n16347 , n16348 , n16349 , n16350 , n16351 , n16352 , n16353 , n16354 , n16355 , n16356 , n16357 , n16358 , n16359 , n16360 , n16361 , n16362 , n16363 , n16364 , n16365 , n16366 , n16367 , n16368 , n16369 , n16370 , n16371 , n16372 , n16373 , n16374 , n16375 , n16376 , n16377 , n16378 , n16379 , n16380 , n16381 , n16382 , n16383 , n16384 , n16385 , n16386 , n16387 , n16388 , n16389 , n16390 , n16391 , n16392 , n16393 , n16394 , n16395 , n16396 , n16397 , n16398 , n16399 , n16400 , n16401 , n16402 , n16403 , n16404 , n16405 , n16406 , n16407 , n16408 , n16409 , n16410 , n16411 , n16412 , n16413 , n16414 , n16415 , n16416 , n16417 , n16418 , n16419 , n16420 , n16421 , n16422 , n16423 , n16424 , n16425 , n16426 , n16427 , n16428 , n16429 , n16430 , n16431 , n16432 , n16433 , n16434 , n16435 , n16436 , n16437 , n16438 , n16439 , n16440 , n16441 , n16442 , n16443 , n16444 , n16445 , n16446 , n16447 , n16448 , n16449 , n16450 , n16451 , n16452 , n16453 , n16454 , n16455 , n16456 , n16457 , n16458 , n16459 , n16460 , n16461 , n16462 , n16463 , n16464 , n16465 , n16466 , n16467 , n16468 , n16469 , n16470 , n16471 , n16472 , n16473 , n16474 , n16475 , n16476 , n16477 , n16478 , n16479 , n16480 , n16481 , n16482 , n16483 , n16484 , n16485 , n16486 , n16487 , n16488 , n16489 , n16490 , n16491 , n16492 , n16493 , n16494 , n16495 , n16496 , n16497 , n16498 , n16499 , n16500 , n16501 , n16502 , n16503 , n16504 , n16505 , n16506 , n16507 , n16508 , n16509 , n16510 , n16511 , n16512 , n16513 , n16514 , n16515 , n16516 , n16517 , n16518 , n16519 , n16520 , n16521 , n16522 , n16523 , n16524 , n16525 , n16526 , n16527 , n16528 , n16529 , n16530 , n16531 , n16532 , n16533 , n16534 , n16535 , n16536 , n16537 , n16538 , n16539 , n16540 , n16541 , n16542 , n16543 , n16544 , n16545 , n16546 , n16547 , n16548 , n16549 , n16550 , n16551 , n16552 , n16553 , n16554 , n16555 , n16556 , n16557 , n16558 , n16559 , n16560 , n16561 , n16562 , n16563 , n16564 , n16565 , n16566 , n16567 , n16568 , n16569 , n16570 , n16571 , n16572 , n16573 , n16574 , n16575 , n16576 , n16577 , n16578 , n16579 , n16580 , n16581 , n16582 , n16583 , n16584 , n16585 , n16586 , n16587 , n16588 , n16589 , n16590 , n16591 , n16592 , n16593 , n16594 , n16595 , n16596 , n16597 , n16598 , n16599 , n16600 , n16601 , n16602 , n16603 , n16604 , n16605 , n16606 , n16607 , n16608 , n16609 , n16610 , n16611 , n16612 , n16613 , n16614 , n16615 , n16616 , n16617 , n16618 , n16619 , n16620 , n16621 , n16622 , n16623 , n16624 , n16625 , n16626 , n16627 , n16628 , n16629 , n16630 , n16631 , n16632 , n16633 , n16634 , n16635 , n16636 , n16637 , n16638 , n16639 , n16640 , n16641 , n16642 , n16643 , n16644 , n16645 , n16646 , n16647 , n16648 , n16649 , n16650 , n16651 , n16652 , n16653 , n16654 , n16655 , n16656 , n16657 , n16658 , n16659 , n16660 , n16661 , n16662 , n16663 , n16664 , n16665 , n16666 , n16667 , n16668 , n16669 , n16670 , n16671 , n16672 , n16673 , n16674 , n16675 , n16676 , n16677 , n16678 , n16679 , n16680 , n16681 , n16682 , n16683 , n16684 , n16685 , n16686 , n16687 , n16688 , n16689 , n16690 , n16691 , n16692 , n16693 , n16694 , n16695 , n16696 , n16697 , n16698 , n16699 , n16700 , n16701 , n16702 , n16703 , n16704 , n16705 , n16706 , n16707 , n16708 , n16709 , n16710 , n16711 , n16712 , n16713 , n16714 , n16715 , n16716 , n16717 , n16718 , n16719 , n16720 , n16721 , n16722 , n16723 , n16724 , n16725 , n16726 , n16727 , n16728 , n16729 , n16730 , n16731 , n16732 , n16733 , n16734 , n16735 , n16736 , n16737 , n16738 , n16739 , n16740 , n16741 , n16742 , n16743 , n16744 , n16745 , n16746 , n16747 , n16748 , n16749 , n16750 , n16751 , n16752 , n16753 , n16754 , n16755 , n16756 , n16757 , n16758 , n16759 , n16760 , n16761 , n16762 , n16763 , n16764 , n16765 , n16766 , n16767 , n16768 , n16769 , n16770 , n16771 , n16772 , n16773 , n16774 , n16775 , n16776 , n16777 , n16778 , n16779 , n16780 , n16781 , n16782 , n16783 , n16784 , n16785 , n16786 , n16787 , n16788 , n16789 , n16790 , n16791 , n16792 , n16793 , n16794 , n16795 , n16796 , n16797 , n16798 , n16799 , n16800 , n16801 , n16802 , n16803 , n16804 , n16805 , n16806 , n16807 , n16808 , n16809 , n16810 , n16811 , n16812 , n16813 , n16814 , n16815 , n16816 , n16817 , n16818 , n16819 , n16820 , n16821 , n16822 , n16823 , n16824 , n16825 , n16826 , n16827 , n16828 , n16829 , n16830 , n16831 , n16832 , n16833 , n16834 , n16835 , n16836 , n16837 , n16838 , n16839 , n16840 , n16841 , n16842 , n16843 , n16844 , n16845 , n16846 , n16847 , n16848 , n16849 , n16850 , n16851 , n16852 , n16853 , n16854 , n16855 , n16856 , n16857 , n16858 , n16859 , n16860 , n16861 , n16862 , n16863 , n16864 , n16865 , n16866 , n16867 , n16868 , n16869 , n16870 , n16871 , n16872 , n16873 , n16874 , n16875 , n16876 , n16877 , n16878 , n16879 , n16880 , n16881 , n16882 , n16883 , n16884 , n16885 , n16886 , n16887 , n16888 , n16889 , n16890 , n16891 , n16892 , n16893 , n16894 , n16895 , n16896 , n16897 , n16898 , n16899 , n16900 , n16901 , n16902 , n16903 , n16904 , n16905 , n16906 , n16907 , n16908 , n16909 , n16910 , n16911 , n16912 , n16913 , n16914 , n16915 , n16916 , n16917 , n16918 , n16919 , n16920 , n16921 , n16922 , n16923 , n16924 , n16925 , n16926 , n16927 , n16928 , n16929 , n16930 , n16931 , n16932 , n16933 , n16934 , n16935 , n16936 , n16937 , n16938 , n16939 , n16940 , n16941 , n16942 , n16943 , n16944 , n16945 , n16946 , n16947 , n16948 , n16949 , n16950 , n16951 , n16952 , n16953 , n16954 , n16955 , n16956 , n16957 , n16958 , n16959 , n16960 , n16961 , n16962 , n16963 , n16964 , n16965 , n16966 , n16967 , n16968 , n16969 , n16970 , n16971 , n16972 , n16973 , n16974 , n16975 , n16976 , n16977 , n16978 , n16979 , n16980 , n16981 , n16982 , n16983 , n16984 , n16985 , n16986 , n16987 , n16988 , n16989 , n16990 , n16991 , n16992 , n16993 , n16994 , n16995 , n16996 , n16997 , n16998 , n16999 , n17000 , n17001 , n17002 , n17003 , n17004 , n17005 , n17006 , n17007 , n17008 , n17009 , n17010 , n17011 , n17012 , n17013 , n17014 , n17015 , n17016 , n17017 , n17018 , n17019 , n17020 , n17021 , n17022 , n17023 , n17024 , n17025 , n17026 , n17027 , n17028 , n17029 , n17030 , n17031 , n17032 , n17033 , n17034 , n17035 , n17036 , n17037 , n17038 , n17039 , n17040 , n17041 , n17042 , n17043 , n17044 , n17045 , n17046 , n17047 , n17048 , n17049 , n17050 , n17051 , n17052 , n17053 , n17054 , n17055 , n17056 , n17057 , n17058 , n17059 , n17060 , n17061 , n17062 , n17063 , n17064 , n17065 , n17066 , n17067 , n17068 , n17069 , n17070 , n17071 , n17072 , n17073 , n17074 , n17075 , n17076 , n17077 , n17078 , n17079 , n17080 , n17081 , n17082 , n17083 , n17084 , n17085 , n17086 , n17087 , n17088 , n17089 , n17090 , n17091 , n17092 , n17093 , n17094 , n17095 , n17096 , n17097 , n17098 , n17099 , n17100 , n17101 , n17102 , n17103 , n17104 , n17105 , n17106 , n17107 , n17108 , n17109 , n17110 , n17111 , n17112 , n17113 , n17114 , n17115 , n17116 , n17117 , n17118 , n17119 , n17120 , n17121 , n17122 , n17123 , n17124 , n17125 , n17126 , n17127 , n17128 , n17129 , n17130 , n17131 , n17132 , n17133 , n17134 , n17135 , n17136 , n17137 , n17138 , n17139 , n17140 , n17141 , n17142 , n17143 , n17144 , n17145 , n17146 , n17147 , n17148 , n17149 , n17150 , n17151 , n17152 , n17153 , n17154 , n17155 , n17156 , n17157 , n17158 , n17159 , n17160 , n17161 , n17162 , n17163 , n17164 , n17165 , n17166 , n17167 , n17168 , n17169 , n17170 , n17171 , n17172 , n17173 , n17174 , n17175 , n17176 , n17177 , n17178 , n17179 , n17180 , n17181 , n17182 , n17183 , n17184 , n17185 , n17186 , n17187 , n17188 , n17189 , n17190 , n17191 , n17192 , n17193 , n17194 , n17195 , n17196 , n17197 , n17198 , n17199 , n17200 , n17201 , n17202 , n17203 , n17204 , n17205 , n17206 , n17207 , n17208 , n17209 , n17210 , n17211 , n17212 , n17213 , n17214 , n17215 , n17216 , n17217 , n17218 , n17219 , n17220 , n17221 , n17222 , n17223 , n17224 , n17225 , n17226 , n17227 , n17228 , n17229 , n17230 , n17231 , n17232 , n17233 , n17234 , n17235 , n17236 , n17237 , n17238 , n17239 , n17240 , n17241 , n17242 , n17243 , n17244 , n17245 , n17246 , n17247 , n17248 , n17249 , n17250 , n17251 , n17252 , n17253 , n17254 , n17255 , n17256 , n17257 , n17258 , n17259 , n17260 , n17261 , n17262 , n17263 , n17264 , n17265 , n17266 , n17267 , n17268 , n17269 , n17270 , n17271 , n17272 , n17273 , n17274 , n17275 , n17276 , n17277 , n17278 , n17279 , n17280 , n17281 , n17282 , n17283 , n17284 , n17285 , n17286 , n17287 , n17288 , n17289 , n17290 , n17291 , n17292 , n17293 , n17294 , n17295 , n17296 , n17297 , n17298 , n17299 , n17300 , n17301 , n17302 , n17303 , n17304 , n17305 , n17306 , n17307 , n17308 , n17309 , n17310 , n17311 , n17312 , n17313 , n17314 , n17315 , n17316 , n17317 , n17318 , n17319 , n17320 , n17321 , n17322 , n17323 , n17324 , n17325 , n17326 , n17327 , n17328 , n17329 , n17330 , n17331 , n17332 , n17333 , n17334 , n17335 , n17336 , n17337 , n17338 , n17339 , n17340 , n17341 , n17342 , n17343 , n17344 , n17345 , n17346 , n17347 , n17348 , n17349 , n17350 , n17351 , n17352 , n17353 , n17354 , n17355 , n17356 , n17357 , n17358 , n17359 , n17360 , n17361 , n17362 , n17363 , n17364 , n17365 , n17366 , n17367 , n17368 , n17369 , n17370 , n17371 , n17372 , n17373 , n17374 , n17375 , n17376 , n17377 , n17378 , n17379 , n17380 , n17381 , n17382 , n17383 , n17384 , n17385 , n17386 , n17387 , n17388 , n17389 , n17390 , n17391 , n17392 , n17393 , n17394 , n17395 , n17396 , n17397 , n17398 , n17399 , n17400 , n17401 , n17402 , n17403 , n17404 , n17405 , n17406 , n17407 , n17408 , n17409 , n17410 , n17411 , n17412 , n17413 , n17414 , n17415 , n17416 , n17417 , n17418 , n17419 , n17420 , n17421 , n17422 , n17423 , n17424 , n17425 , n17426 , n17427 , n17428 , n17429 , n17430 , n17431 , n17432 , n17433 , n17434 , n17435 , n17436 , n17437 , n17438 , n17439 , n17440 , n17441 , n17442 , n17443 , n17444 , n17445 , n17446 , n17447 , n17448 , n17449 , n17450 , n17451 , n17452 , n17453 , n17454 , n17455 , n17456 , n17457 , n17458 , n17459 , n17460 , n17461 , n17462 , n17463 , n17464 , n17465 , n17466 , n17467 , n17468 , n17469 , n17470 , n17471 , n17472 , n17473 , n17474 , n17475 , n17476 , n17477 , n17478 , n17479 , n17480 , n17481 , n17482 , n17483 , n17484 , n17485 , n17486 , n17487 , n17488 , n17489 , n17490 , n17491 , n17492 , n17493 , n17494 , n17495 , n17496 , n17497 , n17498 , n17499 , n17500 , n17501 , n17502 , n17503 , n17504 , n17505 , n17506 , n17507 , n17508 , n17509 , n17510 , n17511 , n17512 , n17513 , n17514 , n17515 , n17516 , n17517 , n17518 , n17519 , n17520 , n17521 , n17522 , n17523 , n17524 , n17525 , n17526 , n17527 , n17528 , n17529 , n17530 , n17531 , n17532 , n17533 , n17534 , n17535 , n17536 , n17537 , n17538 , n17539 , n17540 , n17541 , n17542 , n17543 , n17544 , n17545 , n17546 , n17547 , n17548 , n17549 , n17550 , n17551 , n17552 , n17553 , n17554 , n17555 , n17556 , n17557 , n17558 , n17559 , n17560 , n17561 , n17562 , n17563 , n17564 , n17565 , n17566 , n17567 , n17568 , n17569 , n17570 , n17571 , n17572 , n17573 , n17574 , n17575 , n17576 , n17577 , n17578 , n17579 , n17580 , n17581 , n17582 , n17583 , n17584 , n17585 , n17586 , n17587 , n17588 , n17589 , n17590 , n17591 , n17592 , n17593 , n17594 , n17595 , n17596 , n17597 , n17598 , n17599 , n17600 , n17601 , n17602 , n17603 , n17604 , n17605 , n17606 , n17607 , n17608 , n17609 , n17610 , n17611 , n17612 , n17613 , n17614 , n17615 , n17616 , n17617 , n17618 , n17619 , n17620 , n17621 , n17622 , n17623 , n17624 , n17625 , n17626 , n17627 , n17628 , n17629 , n17630 , n17631 , n17632 , n17633 , n17634 , n17635 , n17636 , n17637 , n17638 , n17639 , n17640 , n17641 , n17642 , n17643 , n17644 , n17645 , n17646 , n17647 , n17648 , n17649 , n17650 , n17651 , n17652 , n17653 , n17654 , n17655 , n17656 , n17657 , n17658 , n17659 , n17660 , n17661 , n17662 , n17663 , n17664 , n17665 , n17666 , n17667 , n17668 , n17669 , n17670 , n17671 , n17672 , n17673 , n17674 , n17675 , n17676 , n17677 , n17678 , n17679 , n17680 , n17681 , n17682 , n17683 , n17684 , n17685 , n17686 , n17687 , n17688 , n17689 , n17690 , n17691 , n17692 , n17693 , n17694 , n17695 , n17696 , n17697 , n17698 , n17699 , n17700 , n17701 , n17702 , n17703 , n17704 , n17705 , n17706 , n17707 , n17708 , n17709 , n17710 , n17711 , n17712 , n17713 , n17714 , n17715 , n17716 , n17717 , n17718 , n17719 , n17720 , n17721 , n17722 , n17723 , n17724 , n17725 , n17726 , n17727 , n17728 , n17729 , n17730 , n17731 , n17732 , n17733 , n17734 , n17735 , n17736 , n17737 , n17738 , n17739 , n17740 , n17741 , n17742 , n17743 , n17744 , n17745 , n17746 , n17747 , n17748 , n17749 , n17750 , n17751 , n17752 , n17753 , n17754 , n17755 , n17756 , n17757 , n17758 , n17759 , n17760 , n17761 , n17762 , n17763 , n17764 , n17765 , n17766 , n17767 , n17768 , n17769 , n17770 , n17771 , n17772 , n17773 , n17774 , n17775 , n17776 , n17777 , n17778 , n17779 , n17780 , n17781 , n17782 , n17783 , n17784 , n17785 , n17786 , n17787 , n17788 , n17789 , n17790 , n17791 , n17792 , n17793 , n17794 , n17795 , n17796 , n17797 , n17798 , n17799 , n17800 , n17801 , n17802 , n17803 , n17804 , n17805 , n17806 , n17807 , n17808 , n17809 , n17810 , n17811 , n17812 , n17813 , n17814 , n17815 , n17816 , n17817 , n17818 , n17819 , n17820 , n17821 , n17822 , n17823 , n17824 , n17825 , n17826 , n17827 , n17828 , n17829 , n17830 , n17831 , n17832 , n17833 , n17834 , n17835 , n17836 , n17837 , n17838 , n17839 , n17840 , n17841 , n17842 , n17843 , n17844 , n17845 , n17846 , n17847 , n17848 , n17849 , n17850 , n17851 , n17852 , n17853 , n17854 , n17855 , n17856 , n17857 , n17858 , n17859 , n17860 , n17861 , n17862 , n17863 , n17864 , n17865 , n17866 , n17867 , n17868 , n17869 , n17870 , n17871 , n17872 , n17873 , n17874 , n17875 , n17876 , n17877 , n17878 , n17879 , n17880 , n17881 , n17882 , n17883 , n17884 , n17885 , n17886 , n17887 , n17888 , n17889 , n17890 , n17891 , n17892 , n17893 , n17894 , n17895 , n17896 , n17897 , n17898 , n17899 , n17900 , n17901 , n17902 , n17903 , n17904 , n17905 , n17906 , n17907 , n17908 , n17909 , n17910 , n17911 , n17912 , n17913 , n17914 , n17915 , n17916 , n17917 , n17918 , n17919 , n17920 , n17921 , n17922 , n17923 , n17924 , n17925 , n17926 , n17927 , n17928 , n17929 , n17930 , n17931 , n17932 , n17933 , n17934 , n17935 , n17936 , n17937 , n17938 , n17939 , n17940 , n17941 , n17942 , n17943 , n17944 , n17945 , n17946 , n17947 , n17948 , n17949 , n17950 , n17951 , n17952 , n17953 , n17954 , n17955 , n17956 , n17957 , n17958 , n17959 , n17960 , n17961 , n17962 , n17963 , n17964 , n17965 , n17966 , n17967 , n17968 , n17969 , n17970 , n17971 , n17972 , n17973 , n17974 , n17975 , n17976 , n17977 , n17978 , n17979 , n17980 , n17981 , n17982 , n17983 , n17984 , n17985 , n17986 , n17987 , n17988 , n17989 , n17990 , n17991 , n17992 , n17993 , n17994 , n17995 , n17996 , n17997 , n17998 , n17999 , n18000 , n18001 , n18002 , n18003 , n18004 , n18005 , n18006 , n18007 , n18008 , n18009 , n18010 , n18011 , n18012 , n18013 , n18014 , n18015 , n18016 , n18017 , n18018 , n18019 , n18020 , n18021 , n18022 , n18023 , n18024 , n18025 , n18026 , n18027 , n18028 , n18029 , n18030 , n18031 , n18032 , n18033 , n18034 , n18035 , n18036 , n18037 , n18038 , n18039 , n18040 , n18041 , n18042 , n18043 , n18044 , n18045 , n18046 , n18047 , n18048 , n18049 , n18050 , n18051 , n18052 , n18053 , n18054 , n18055 , n18056 , n18057 , n18058 , n18059 , n18060 , n18061 , n18062 , n18063 , n18064 , n18065 , n18066 , n18067 , n18068 , n18069 , n18070 , n18071 , n18072 , n18073 , n18074 , n18075 , n18076 , n18077 , n18078 , n18079 , n18080 , n18081 , n18082 , n18083 , n18084 , n18085 , n18086 , n18087 , n18088 , n18089 , n18090 , n18091 , n18092 , n18093 , n18094 , n18095 , n18096 , n18097 , n18098 , n18099 , n18100 , n18101 , n18102 , n18103 , n18104 , n18105 , n18106 , n18107 , n18108 , n18109 , n18110 , n18111 , n18112 , n18113 , n18114 , n18115 , n18116 , n18117 , n18118 , n18119 , n18120 , n18121 , n18122 , n18123 , n18124 , n18125 , n18126 , n18127 , n18128 , n18129 , n18130 , n18131 , n18132 , n18133 , n18134 , n18135 , n18136 , n18137 , n18138 , n18139 , n18140 , n18141 , n18142 , n18143 , n18144 , n18145 , n18146 , n18147 , n18148 , n18149 , n18150 , n18151 , n18152 , n18153 , n18154 , n18155 , n18156 , n18157 , n18158 , n18159 , n18160 , n18161 , n18162 , n18163 , n18164 , n18165 , n18166 , n18167 , n18168 , n18169 , n18170 , n18171 , n18172 , n18173 , n18174 , n18175 , n18176 , n18177 , n18178 , n18179 , n18180 , n18181 , n18182 , n18183 , n18184 , n18185 , n18186 , n18187 , n18188 , n18189 , n18190 , n18191 , n18192 , n18193 , n18194 , n18195 , n18196 , n18197 , n18198 , n18199 , n18200 , n18201 , n18202 , n18203 , n18204 , n18205 , n18206 , n18207 , n18208 , n18209 , n18210 , n18211 , n18212 , n18213 , n18214 , n18215 , n18216 , n18217 , n18218 , n18219 , n18220 , n18221 , n18222 , n18223 , n18224 , n18225 , n18226 , n18227 , n18228 , n18229 , n18230 , n18231 , n18232 , n18233 , n18234 , n18235 , n18236 , n18237 , n18238 , n18239 , n18240 , n18241 , n18242 , n18243 , n18244 , n18245 , n18246 , n18247 , n18248 , n18249 , n18250 , n18251 , n18252 , n18253 , n18254 , n18255 , n18256 , n18257 , n18258 , n18259 , n18260 , n18261 , n18262 , n18263 , n18264 , n18265 , n18266 , n18267 , n18268 , n18269 , n18270 , n18271 , n18272 , n18273 , n18274 , n18275 , n18276 , n18277 , n18278 , n18279 , n18280 , n18281 , n18282 , n18283 , n18284 , n18285 , n18286 , n18287 , n18288 , n18289 , n18290 , n18291 , n18292 , n18293 , n18294 , n18295 , n18296 , n18297 , n18298 , n18299 , n18300 , n18301 , n18302 , n18303 , n18304 , n18305 , n18306 , n18307 , n18308 , n18309 , n18310 , n18311 , n18312 , n18313 , n18314 , n18315 , n18316 , n18317 , n18318 , n18319 , n18320 , n18321 , n18322 , n18323 , n18324 , n18325 , n18326 , n18327 , n18328 , n18329 , n18330 , n18331 , n18332 , n18333 , n18334 , n18335 , n18336 , n18337 , n18338 , n18339 , n18340 , n18341 , n18342 , n18343 , n18344 , n18345 , n18346 , n18347 , n18348 , n18349 , n18350 , n18351 , n18352 , n18353 , n18354 , n18355 , n18356 , n18357 , n18358 , n18359 , n18360 , n18361 , n18362 , n18363 , n18364 , n18365 , n18366 , n18367 , n18368 , n18369 , n18370 , n18371 , n18372 , n18373 , n18374 , n18375 , n18376 , n18377 , n18378 , n18379 , n18380 , n18381 , n18382 , n18383 , n18384 , n18385 , n18386 , n18387 , n18388 , n18389 , n18390 , n18391 , n18392 , n18393 , n18394 , n18395 , n18396 , n18397 , n18398 , n18399 , n18400 , n18401 , n18402 , n18403 , n18404 , n18405 , n18406 , n18407 , n18408 , n18409 , n18410 , n18411 , n18412 , n18413 , n18414 , n18415 , n18416 , n18417 , n18418 , n18419 , n18420 , n18421 , n18422 , n18423 , n18424 , n18425 , n18426 , n18427 , n18428 , n18429 , n18430 , n18431 , n18432 , n18433 , n18434 , n18435 , n18436 , n18437 , n18438 , n18439 , n18440 , n18441 , n18442 , n18443 , n18444 , n18445 , n18446 , n18447 , n18448 , n18449 , n18450 , n18451 , n18452 , n18453 , n18454 , n18455 , n18456 , n18457 , n18458 , n18459 , n18460 , n18461 , n18462 , n18463 , n18464 , n18465 , n18466 , n18467 , n18468 , n18469 , n18470 , n18471 , n18472 , n18473 , n18474 , n18475 , n18476 , n18477 , n18478 , n18479 , n18480 , n18481 , n18482 , n18483 , n18484 , n18485 , n18486 , n18487 , n18488 , n18489 , n18490 , n18491 , n18492 , n18493 , n18494 , n18495 , n18496 , n18497 , n18498 , n18499 , n18500 , n18501 , n18502 , n18503 , n18504 , n18505 , n18506 , n18507 , n18508 , n18509 , n18510 , n18511 , n18512 , n18513 , n18514 , n18515 , n18516 , n18517 , n18518 , n18519 , n18520 , n18521 , n18522 , n18523 , n18524 , n18525 , n18526 , n18527 , n18528 , n18529 , n18530 , n18531 , n18532 , n18533 , n18534 , n18535 , n18536 , n18537 , n18538 , n18539 , n18540 , n18541 , n18542 , n18543 , n18544 , n18545 , n18546 , n18547 , n18548 , n18549 , n18550 , n18551 , n18552 , n18553 , n18554 , n18555 , n18556 , n18557 , n18558 , n18559 , n18560 , n18561 , n18562 , n18563 , n18564 , n18565 , n18566 , n18567 , n18568 , n18569 , n18570 , n18571 , n18572 , n18573 , n18574 , n18575 , n18576 , n18577 , n18578 , n18579 , n18580 , n18581 , n18582 , n18583 , n18584 , n18585 , n18586 , n18587 , n18588 , n18589 , n18590 , n18591 , n18592 , n18593 , n18594 , n18595 , n18596 , n18597 , n18598 , n18599 , n18600 , n18601 , n18602 , n18603 , n18604 , n18605 , n18606 , n18607 , n18608 , n18609 , n18610 , n18611 , n18612 , n18613 , n18614 , n18615 , n18616 , n18617 , n18618 , n18619 , n18620 , n18621 , n18622 , n18623 , n18624 , n18625 , n18626 , n18627 , n18628 , n18629 , n18630 , n18631 , n18632 , n18633 , n18634 , n18635 , n18636 , n18637 , n18638 , n18639 , n18640 , n18641 , n18642 , n18643 , n18644 , n18645 , n18646 , n18647 , n18648 , n18649 , n18650 , n18651 , n18652 , n18653 , n18654 , n18655 , n18656 , n18657 , n18658 , n18659 , n18660 , n18661 , n18662 , n18663 , n18664 , n18665 , n18666 , n18667 , n18668 , n18669 , n18670 , n18671 , n18672 , n18673 , n18674 , n18675 , n18676 , n18677 , n18678 , n18679 , n18680 , n18681 , n18682 , n18683 , n18684 , n18685 , n18686 , n18687 , n18688 , n18689 , n18690 , n18691 , n18692 , n18693 , n18694 , n18695 , n18696 , n18697 , n18698 , n18699 , n18700 , n18701 , n18702 , n18703 , n18704 , n18705 , n18706 , n18707 , n18708 , n18709 , n18710 , n18711 , n18712 , n18713 , n18714 , n18715 , n18716 , n18717 , n18718 , n18719 , n18720 , n18721 , n18722 , n18723 , n18724 , n18725 , n18726 , n18727 , n18728 , n18729 , n18730 , n18731 , n18732 , n18733 , n18734 , n18735 , n18736 , n18737 , n18738 , n18739 , n18740 , n18741 , n18742 , n18743 , n18744 , n18745 , n18746 , n18747 , n18748 , n18749 , n18750 , n18751 , n18752 , n18753 , n18754 , n18755 , n18756 , n18757 , n18758 , n18759 , n18760 , n18761 , n18762 , n18763 , n18764 , n18765 , n18766 , n18767 , n18768 , n18769 , n18770 , n18771 , n18772 , n18773 , n18774 , n18775 , n18776 , n18777 , n18778 , n18779 , n18780 , n18781 , n18782 , n18783 , n18784 , n18785 , n18786 , n18787 , n18788 , n18789 , n18790 , n18791 , n18792 , n18793 , n18794 , n18795 , n18796 , n18797 , n18798 , n18799 , n18800 , n18801 , n18802 , n18803 , n18804 , n18805 , n18806 , n18807 , n18808 , n18809 , n18810 , n18811 , n18812 , n18813 , n18814 , n18815 , n18816 , n18817 , n18818 , n18819 , n18820 , n18821 , n18822 , n18823 , n18824 , n18825 , n18826 , n18827 , n18828 , n18829 , n18830 , n18831 , n18832 , n18833 , n18834 , n18835 , n18836 , n18837 , n18838 , n18839 , n18840 , n18841 , n18842 , n18843 , n18844 , n18845 , n18846 , n18847 , n18848 , n18849 , n18850 , n18851 , n18852 , n18853 , n18854 , n18855 , n18856 , n18857 , n18858 , n18859 , n18860 , n18861 , n18862 , n18863 , n18864 , n18865 , n18866 , n18867 , n18868 , n18869 , n18870 , n18871 , n18872 , n18873 , n18874 , n18875 , n18876 , n18877 , n18878 , n18879 , n18880 , n18881 , n18882 , n18883 , n18884 , n18885 , n18886 , n18887 , n18888 , n18889 , n18890 , n18891 , n18892 , n18893 , n18894 , n18895 , n18896 , n18897 , n18898 , n18899 , n18900 , n18901 , n18902 , n18903 , n18904 , n18905 , n18906 , n18907 , n18908 , n18909 , n18910 , n18911 , n18912 , n18913 , n18914 , n18915 , n18916 , n18917 , n18918 , n18919 , n18920 , n18921 , n18922 , n18923 , n18924 , n18925 , n18926 , n18927 , n18928 , n18929 , n18930 , n18931 , n18932 , n18933 , n18934 , n18935 , n18936 , n18937 , n18938 , n18939 , n18940 , n18941 , n18942 , n18943 , n18944 , n18945 , n18946 , n18947 , n18948 , n18949 , n18950 , n18951 , n18952 , n18953 , n18954 , n18955 , n18956 , n18957 , n18958 , n18959 , n18960 , n18961 , n18962 , n18963 , n18964 , n18965 , n18966 , n18967 , n18968 , n18969 , n18970 , n18971 , n18972 , n18973 , n18974 , n18975 , n18976 , n18977 , n18978 , n18979 , n18980 , n18981 , n18982 , n18983 , n18984 , n18985 , n18986 , n18987 , n18988 , n18989 , n18990 , n18991 , n18992 , n18993 , n18994 , n18995 , n18996 , n18997 , n18998 , n18999 , n19000 , n19001 , n19002 , n19003 , n19004 , n19005 , n19006 , n19007 , n19008 , n19009 , n19010 , n19011 , n19012 , n19013 , n19014 , n19015 , n19016 , n19017 , n19018 , n19019 , n19020 , n19021 , n19022 , n19023 , n19024 , n19025 , n19026 , n19027 , n19028 , n19029 , n19030 , n19031 , n19032 , n19033 , n19034 , n19035 , n19036 , n19037 , n19038 , n19039 , n19040 , n19041 , n19042 , n19043 , n19044 , n19045 , n19046 , n19047 , n19048 , n19049 , n19050 , n19051 , n19052 , n19053 , n19054 , n19055 , n19056 , n19057 , n19058 , n19059 , n19060 , n19061 , n19062 , n19063 , n19064 , n19065 , n19066 , n19067 , n19068 , n19069 , n19070 , n19071 , n19072 , n19073 , n19074 , n19075 , n19076 , n19077 , n19078 , n19079 , n19080 , n19081 , n19082 , n19083 , n19084 , n19085 , n19086 , n19087 , n19088 , n19089 , n19090 , n19091 , n19092 , n19093 , n19094 , n19095 , n19096 , n19097 , n19098 , n19099 , n19100 , n19101 , n19102 , n19103 , n19104 , n19105 , n19106 , n19107 , n19108 , n19109 , n19110 , n19111 , n19112 , n19113 , n19114 , n19115 , n19116 , n19117 , n19118 , n19119 , n19120 , n19121 , n19122 , n19123 , n19124 , n19125 , n19126 , n19127 , n19128 , n19129 , n19130 , n19131 , n19132 , n19133 , n19134 , n19135 , n19136 , n19137 , n19138 , n19139 , n19140 , n19141 , n19142 , n19143 , n19144 , n19145 , n19146 , n19147 , n19148 , n19149 , n19150 , n19151 , n19152 , n19153 , n19154 , n19155 , n19156 , n19157 , n19158 , n19159 , n19160 , n19161 , n19162 , n19163 , n19164 , n19165 , n19166 , n19167 , n19168 , n19169 , n19170 , n19171 , n19172 , n19173 , n19174 , n19175 , n19176 , n19177 , n19178 , n19179 , n19180 , n19181 , n19182 , n19183 , n19184 , n19185 , n19186 , n19187 , n19188 , n19189 , n19190 , n19191 , n19192 , n19193 , n19194 , n19195 , n19196 , n19197 , n19198 , n19199 , n19200 , n19201 , n19202 , n19203 , n19204 , n19205 , n19206 , n19207 , n19208 , n19209 , n19210 , n19211 , n19212 , n19213 , n19214 , n19215 , n19216 , n19217 , n19218 , n19219 , n19220 , n19221 , n19222 , n19223 , n19224 , n19225 , n19226 , n19227 , n19228 , n19229 , n19230 , n19231 , n19232 , n19233 , n19234 , n19235 , n19236 , n19237 , n19238 , n19239 , n19240 , n19241 , n19242 , n19243 , n19244 , n19245 , n19246 , n19247 , n19248 , n19249 , n19250 , n19251 , n19252 , n19253 , n19254 , n19255 , n19256 , n19257 , n19258 , n19259 , n19260 , n19261 , n19262 , n19263 , n19264 , n19265 , n19266 , n19267 , n19268 , n19269 , n19270 , n19271 , n19272 , n19273 , n19274 , n19275 , n19276 , n19277 , n19278 , n19279 , n19280 , n19281 , n19282 , n19283 , n19284 , n19285 , n19286 , n19287 , n19288 , n19289 , n19290 , n19291 , n19292 , n19293 , n19294 , n19295 , n19296 , n19297 , n19298 , n19299 , n19300 , n19301 , n19302 , n19303 , n19304 , n19305 , n19306 , n19307 , n19308 , n19309 , n19310 , n19311 , n19312 , n19313 , n19314 , n19315 , n19316 , n19317 , n19318 , n19319 , n19320 , n19321 , n19322 , n19323 , n19324 , n19325 , n19326 , n19327 , n19328 , n19329 , n19330 , n19331 , n19332 , n19333 , n19334 , n19335 , n19336 , n19337 , n19338 , n19339 , n19340 , n19341 , n19342 , n19343 , n19344 , n19345 , n19346 , n19347 , n19348 , n19349 , n19350 , n19351 , n19352 , n19353 , n19354 , n19355 , n19356 , n19357 , n19358 , n19359 , n19360 , n19361 , n19362 , n19363 , n19364 , n19365 , n19366 , n19367 , n19368 , n19369 , n19370 , n19371 , n19372 , n19373 , n19374 , n19375 , n19376 , n19377 , n19378 , n19379 , n19380 , n19381 , n19382 , n19383 , n19384 , n19385 , n19386 , n19387 , n19388 , n19389 , n19390 , n19391 , n19392 , n19393 , n19394 , n19395 , n19396 , n19397 , n19398 , n19399 , n19400 , n19401 , n19402 , n19403 , n19404 , n19405 , n19406 , n19407 , n19408 , n19409 , n19410 , n19411 , n19412 , n19413 , n19414 , n19415 , n19416 , n19417 , n19418 , n19419 , n19420 , n19421 , n19422 , n19423 , n19424 , n19425 , n19426 , n19427 , n19428 , n19429 , n19430 , n19431 , n19432 , n19433 , n19434 , n19435 , n19436 , n19437 , n19438 , n19439 , n19440 , n19441 , n19442 , n19443 , n19444 , n19445 , n19446 , n19447 , n19448 , n19449 , n19450 , n19451 , n19452 , n19453 , n19454 , n19455 , n19456 , n19457 , n19458 , n19459 , n19460 , n19461 , n19462 , n19463 , n19464 , n19465 , n19466 , n19467 , n19468 , n19469 , n19470 , n19471 , n19472 , n19473 , n19474 , n19475 , n19476 , n19477 , n19478 , n19479 , n19480 , n19481 , n19482 , n19483 , n19484 , n19485 , n19486 , n19487 , n19488 , n19489 , n19490 , n19491 , n19492 , n19493 , n19494 , n19495 , n19496 , n19497 , n19498 , n19499 , n19500 , n19501 , n19502 , n19503 , n19504 , n19505 , n19506 , n19507 , n19508 , n19509 , n19510 , n19511 , n19512 , n19513 , n19514 , n19515 , n19516 , n19517 , n19518 , n19519 , n19520 , n19521 , n19522 , n19523 , n19524 , n19525 , n19526 , n19527 , n19528 , n19529 , n19530 , n19531 , n19532 , n19533 , n19534 , n19535 , n19536 , n19537 , n19538 , n19539 , n19540 , n19541 , n19542 , n19543 , n19544 , n19545 , n19546 , n19547 , n19548 , n19549 , n19550 , n19551 , n19552 , n19553 , n19554 , n19555 , n19556 , n19557 , n19558 , n19559 , n19560 , n19561 , n19562 , n19563 , n19564 , n19565 , n19566 , n19567 , n19568 , n19569 , n19570 , n19571 , n19572 , n19573 , n19574 , n19575 , n19576 , n19577 , n19578 , n19579 , n19580 , n19581 , n19582 , n19583 , n19584 , n19585 , n19586 , n19587 , n19588 , n19589 , n19590 , n19591 , n19592 , n19593 , n19594 , n19595 , n19596 , n19597 , n19598 , n19599 , n19600 , n19601 , n19602 , n19603 , n19604 , n19605 , n19606 , n19607 , n19608 , n19609 , n19610 , n19611 , n19612 , n19613 , n19614 , n19615 , n19616 , n19617 , n19618 , n19619 , n19620 , n19621 , n19622 , n19623 , n19624 , n19625 , n19626 , n19627 , n19628 , n19629 , n19630 , n19631 , n19632 , n19633 , n19634 , n19635 , n19636 , n19637 , n19638 , n19639 , n19640 , n19641 , n19642 , n19643 , n19644 , n19645 , n19646 , n19647 , n19648 , n19649 , n19650 , n19651 , n19652 , n19653 , n19654 , n19655 , n19656 , n19657 , n19658 , n19659 , n19660 , n19661 , n19662 , n19663 , n19664 , n19665 , n19666 , n19667 , n19668 , n19669 , n19670 , n19671 , n19672 , n19673 , n19674 , n19675 , n19676 , n19677 , n19678 , n19679 , n19680 , n19681 , n19682 , n19683 , n19684 , n19685 , n19686 , n19687 , n19688 , n19689 , n19690 , n19691 , n19692 , n19693 , n19694 , n19695 , n19696 , n19697 , n19698 , n19699 , n19700 , n19701 , n19702 , n19703 , n19704 , n19705 , n19706 , n19707 , n19708 , n19709 , n19710 , n19711 , n19712 , n19713 , n19714 , n19715 , n19716 , n19717 , n19718 , n19719 , n19720 , n19721 , n19722 , n19723 , n19724 , n19725 , n19726 , n19727 , n19728 , n19729 , n19730 , n19731 , n19732 , n19733 , n19734 , n19735 , n19736 , n19737 , n19738 , n19739 , n19740 , n19741 , n19742 , n19743 , n19744 , n19745 , n19746 , n19747 , n19748 , n19749 , n19750 , n19751 , n19752 , n19753 , n19754 , n19755 , n19756 , n19757 , n19758 , n19759 , n19760 , n19761 , n19762 , n19763 , n19764 , n19765 , n19766 , n19767 , n19768 , n19769 , n19770 , n19771 , n19772 , n19773 , n19774 , n19775 , n19776 , n19777 , n19778 , n19779 , n19780 , n19781 , n19782 , n19783 , n19784 , n19785 , n19786 , n19787 , n19788 , n19789 , n19790 , n19791 , n19792 , n19793 , n19794 , n19795 , n19796 , n19797 , n19798 , n19799 , n19800 , n19801 , n19802 , n19803 , n19804 , n19805 , n19806 , n19807 , n19808 , n19809 , n19810 , n19811 , n19812 , n19813 , n19814 , n19815 , n19816 , n19817 , n19818 , n19819 , n19820 , n19821 , n19822 , n19823 , n19824 , n19825 , n19826 , n19827 , n19828 , n19829 , n19830 , n19831 , n19832 , n19833 , n19834 , n19835 , n19836 , n19837 , n19838 , n19839 , n19840 , n19841 , n19842 , n19843 , n19844 , n19845 , n19846 , n19847 , n19848 , n19849 , n19850 , n19851 , n19852 , n19853 , n19854 , n19855 , n19856 , n19857 , n19858 , n19859 , n19860 , n19861 , n19862 , n19863 , n19864 , n19865 , n19866 , n19867 , n19868 , n19869 , n19870 , n19871 , n19872 , n19873 , n19874 , n19875 , n19876 , n19877 , n19878 , n19879 , n19880 , n19881 , n19882 , n19883 , n19884 , n19885 , n19886 , n19887 , n19888 , n19889 , n19890 , n19891 , n19892 , n19893 , n19894 , n19895 , n19896 , n19897 , n19898 , n19899 , n19900 , n19901 , n19902 , n19903 , n19904 , n19905 , n19906 , n19907 , n19908 , n19909 , n19910 , n19911 , n19912 , n19913 , n19914 , n19915 , n19916 , n19917 , n19918 , n19919 , n19920 , n19921 , n19922 , n19923 , n19924 , n19925 , n19926 , n19927 , n19928 , n19929 , n19930 , n19931 , n19932 , n19933 , n19934 , n19935 , n19936 , n19937 , n19938 , n19939 , n19940 , n19941 , n19942 , n19943 , n19944 , n19945 , n19946 , n19947 , n19948 , n19949 , n19950 , n19951 , n19952 , n19953 , n19954 , n19955 , n19956 , n19957 , n19958 , n19959 , n19960 , n19961 , n19962 , n19963 , n19964 , n19965 , n19966 , n19967 , n19968 , n19969 , n19970 , n19971 , n19972 , n19973 , n19974 , n19975 , n19976 , n19977 , n19978 , n19979 , n19980 , n19981 , n19982 , n19983 , n19984 , n19985 , n19986 , n19987 , n19988 , n19989 , n19990 , n19991 , n19992 , n19993 , n19994 , n19995 , n19996 , n19997 , n19998 , n19999 , n20000 , n20001 , n20002 , n20003 , n20004 , n20005 , n20006 , n20007 , n20008 , n20009 , n20010 , n20011 , n20012 , n20013 , n20014 , n20015 , n20016 , n20017 , n20018 , n20019 , n20020 , n20021 , n20022 , n20023 , n20024 , n20025 , n20026 , n20027 , n20028 , n20029 , n20030 , n20031 , n20032 , n20033 , n20034 , n20035 , n20036 , n20037 , n20038 , n20039 , n20040 , n20041 , n20042 , n20043 , n20044 , n20045 , n20046 , n20047 , n20048 , n20049 , n20050 , n20051 , n20052 , n20053 , n20054 , n20055 , n20056 , n20057 , n20058 , n20059 , n20060 , n20061 , n20062 , n20063 , n20064 , n20065 , n20066 , n20067 , n20068 , n20069 , n20070 , n20071 , n20072 , n20073 , n20074 , n20075 , n20076 , n20077 , n20078 , n20079 , n20080 , n20081 , n20082 , n20083 , n20084 , n20085 , n20086 , n20087 , n20088 , n20089 , n20090 , n20091 , n20092 , n20093 , n20094 , n20095 , n20096 , n20097 , n20098 , n20099 , n20100 , n20101 , n20102 , n20103 , n20104 , n20105 , n20106 , n20107 , n20108 , n20109 , n20110 , n20111 , n20112 , n20113 , n20114 , n20115 , n20116 , n20117 , n20118 , n20119 , n20120 , n20121 , n20122 , n20123 , n20124 , n20125 , n20126 , n20127 , n20128 , n20129 , n20130 , n20131 , n20132 , n20133 , n20134 , n20135 , n20136 , n20137 , n20138 , n20139 , n20140 , n20141 , n20142 , n20143 , n20144 , n20145 , n20146 , n20147 , n20148 , n20149 , n20150 , n20151 , n20152 , n20153 , n20154 , n20155 , n20156 , n20157 , n20158 , n20159 , n20160 , n20161 , n20162 , n20163 , n20164 , n20165 , n20166 , n20167 , n20168 , n20169 , n20170 , n20171 , n20172 , n20173 , n20174 , n20175 , n20176 , n20177 , n20178 , n20179 , n20180 , n20181 , n20182 , n20183 , n20184 , n20185 , n20186 , n20187 , n20188 , n20189 , n20190 , n20191 , n20192 , n20193 , n20194 , n20195 , n20196 , n20197 , n20198 , n20199 , n20200 , n20201 , n20202 , n20203 , n20204 , n20205 , n20206 , n20207 , n20208 , n20209 , n20210 , n20211 , n20212 , n20213 , n20214 , n20215 , n20216 , n20217 , n20218 , n20219 , n20220 , n20221 , n20222 , n20223 , n20224 , n20225 , n20226 , n20227 , n20228 , n20229 , n20230 , n20231 , n20232 , n20233 , n20234 , n20235 , n20236 , n20237 , n20238 , n20239 , n20240 , n20241 , n20242 , n20243 , n20244 , n20245 , n20246 , n20247 , n20248 , n20249 , n20250 , n20251 , n20252 , n20253 , n20254 , n20255 , n20256 , n20257 , n20258 , n20259 , n20260 , n20261 , n20262 , n20263 , n20264 , n20265 , n20266 , n20267 , n20268 , n20269 , n20270 , n20271 , n20272 , n20273 , n20274 , n20275 , n20276 , n20277 , n20278 , n20279 , n20280 , n20281 , n20282 , n20283 , n20284 , n20285 , n20286 , n20287 , n20288 , n20289 , n20290 , n20291 , n20292 , n20293 , n20294 , n20295 , n20296 , n20297 , n20298 , n20299 , n20300 , n20301 , n20302 , n20303 , n20304 , n20305 , n20306 , n20307 , n20308 , n20309 , n20310 , n20311 , n20312 , n20313 , n20314 , n20315 , n20316 , n20317 , n20318 , n20319 , n20320 , n20321 , n20322 , n20323 , n20324 , n20325 , n20326 , n20327 , n20328 , n20329 , n20330 , n20331 , n20332 , n20333 , n20334 , n20335 , n20336 , n20337 , n20338 , n20339 , n20340 , n20341 , n20342 , n20343 , n20344 , n20345 , n20346 , n20347 , n20348 , n20349 , n20350 , n20351 , n20352 , n20353 , n20354 , n20355 , n20356 , n20357 , n20358 , n20359 , n20360 , n20361 , n20362 , n20363 , n20364 , n20365 , n20366 , n20367 , n20368 , n20369 , n20370 , n20371 , n20372 , n20373 , n20374 , n20375 , n20376 , n20377 , n20378 , n20379 , n20380 , n20381 , n20382 , n20383 , n20384 , n20385 , n20386 , n20387 , n20388 , n20389 , n20390 , n20391 , n20392 , n20393 , n20394 , n20395 , n20396 , n20397 , n20398 , n20399 , n20400 , n20401 , n20402 , n20403 , n20404 , n20405 , n20406 , n20407 , n20408 , n20409 , n20410 , n20411 , n20412 , n20413 , n20414 , n20415 , n20416 , n20417 , n20418 , n20419 , n20420 , n20421 , n20422 , n20423 , n20424 , n20425 , n20426 , n20427 , n20428 , n20429 , n20430 , n20431 , n20432 , n20433 , n20434 , n20435 , n20436 , n20437 , n20438 , n20439 , n20440 , n20441 , n20442 , n20443 , n20444 , n20445 , n20446 , n20447 , n20448 , n20449 , n20450 , n20451 , n20452 , n20453 , n20454 , n20455 , n20456 , n20457 , n20458 , n20459 , n20460 , n20461 , n20462 , n20463 , n20464 , n20465 , n20466 , n20467 , n20468 , n20469 , n20470 , n20471 , n20472 , n20473 , n20474 , n20475 , n20476 , n20477 , n20478 , n20479 , n20480 , n20481 , n20482 , n20483 , n20484 , n20485 , n20486 , n20487 , n20488 , n20489 , n20490 , n20491 , n20492 , n20493 , n20494 , n20495 , n20496 , n20497 , n20498 , n20499 , n20500 , n20501 , n20502 , n20503 , n20504 , n20505 , n20506 , n20507 , n20508 , n20509 , n20510 , n20511 , n20512 , n20513 , n20514 , n20515 , n20516 , n20517 , n20518 , n20519 , n20520 , n20521 , n20522 , n20523 , n20524 , n20525 , n20526 , n20527 , n20528 , n20529 , n20530 , n20531 , n20532 , n20533 , n20534 , n20535 , n20536 , n20537 , n20538 , n20539 , n20540 , n20541 , n20542 , n20543 , n20544 , n20545 , n20546 , n20547 , n20548 , n20549 , n20550 , n20551 , n20552 , n20553 , n20554 , n20555 , n20556 , n20557 , n20558 , n20559 , n20560 , n20561 , n20562 , n20563 , n20564 , n20565 , n20566 , n20567 , n20568 , n20569 , n20570 , n20571 , n20572 , n20573 , n20574 , n20575 , n20576 , n20577 , n20578 , n20579 , n20580 , n20581 , n20582 , n20583 , n20584 , n20585 , n20586 , n20587 , n20588 , n20589 , n20590 , n20591 , n20592 , n20593 , n20594 , n20595 , n20596 , n20597 , n20598 , n20599 , n20600 , n20601 , n20602 , n20603 , n20604 , n20605 , n20606 , n20607 , n20608 , n20609 , n20610 , n20611 , n20612 , n20613 , n20614 , n20615 , n20616 , n20617 , n20618 , n20619 , n20620 , n20621 , n20622 , n20623 , n20624 , n20625 , n20626 , n20627 , n20628 , n20629 , n20630 , n20631 , n20632 , n20633 , n20634 , n20635 , n20636 , n20637 , n20638 , n20639 , n20640 , n20641 , n20642 , n20643 , n20644 , n20645 , n20646 , n20647 , n20648 , n20649 , n20650 , n20651 , n20652 , n20653 , n20654 , n20655 , n20656 , n20657 , n20658 , n20659 , n20660 , n20661 , n20662 , n20663 , n20664 , n20665 , n20666 , n20667 , n20668 , n20669 , n20670 , n20671 , n20672 , n20673 , n20674 , n20675 , n20676 , n20677 , n20678 , n20679 , n20680 , n20681 , n20682 , n20683 , n20684 , n20685 , n20686 , n20687 , n20688 , n20689 , n20690 , n20691 , n20692 , n20693 , n20694 , n20695 , n20696 , n20697 , n20698 , n20699 , n20700 , n20701 , n20702 , n20703 , n20704 , n20705 , n20706 , n20707 , n20708 , n20709 , n20710 , n20711 , n20712 , n20713 , n20714 , n20715 , n20716 , n20717 , n20718 , n20719 , n20720 , n20721 , n20722 , n20723 , n20724 , n20725 , n20726 , n20727 , n20728 , n20729 , n20730 , n20731 , n20732 , n20733 , n20734 , n20735 , n20736 , n20737 , n20738 , n20739 , n20740 , n20741 , n20742 , n20743 , n20744 , n20745 , n20746 , n20747 , n20748 , n20749 , n20750 , n20751 , n20752 , n20753 , n20754 , n20755 , n20756 , n20757 , n20758 , n20759 , n20760 , n20761 , n20762 , n20763 , n20764 , n20765 , n20766 , n20767 , n20768 , n20769 , n20770 , n20771 , n20772 , n20773 , n20774 , n20775 , n20776 , n20777 , n20778 , n20779 , n20780 , n20781 , n20782 , n20783 , n20784 , n20785 , n20786 , n20787 , n20788 , n20789 , n20790 , n20791 , n20792 , n20793 , n20794 , n20795 , n20796 , n20797 , n20798 , n20799 , n20800 , n20801 , n20802 , n20803 , n20804 , n20805 , n20806 , n20807 , n20808 , n20809 , n20810 , n20811 , n20812 , n20813 , n20814 , n20815 , n20816 , n20817 , n20818 , n20819 , n20820 , n20821 , n20822 , n20823 , n20824 , n20825 , n20826 , n20827 , n20828 , n20829 , n20830 , n20831 , n20832 , n20833 , n20834 , n20835 , n20836 , n20837 , n20838 , n20839 , n20840 , n20841 , n20842 , n20843 , n20844 , n20845 , n20846 , n20847 , n20848 , n20849 , n20850 , n20851 , n20852 , n20853 , n20854 , n20855 , n20856 , n20857 , n20858 , n20859 , n20860 , n20861 , n20862 , n20863 , n20864 , n20865 , n20866 , n20867 , n20868 , n20869 , n20870 , n20871 , n20872 , n20873 , n20874 , n20875 , n20876 , n20877 , n20878 , n20879 , n20880 , n20881 , n20882 , n20883 , n20884 , n20885 , n20886 , n20887 , n20888 , n20889 , n20890 , n20891 , n20892 , n20893 , n20894 , n20895 , n20896 , n20897 , n20898 , n20899 , n20900 , n20901 , n20902 , n20903 , n20904 , n20905 , n20906 , n20907 , n20908 , n20909 , n20910 , n20911 , n20912 , n20913 , n20914 , n20915 , n20916 , n20917 , n20918 , n20919 , n20920 , n20921 , n20922 , n20923 , n20924 , n20925 , n20926 , n20927 , n20928 , n20929 , n20930 , n20931 , n20932 , n20933 , n20934 , n20935 , n20936 , n20937 , n20938 , n20939 , n20940 , n20941 , n20942 , n20943 , n20944 , n20945 , n20946 , n20947 , n20948 , n20949 , n20950 , n20951 , n20952 , n20953 , n20954 , n20955 , n20956 , n20957 , n20958 , n20959 , n20960 , n20961 , n20962 , n20963 , n20964 , n20965 , n20966 , n20967 , n20968 , n20969 , n20970 , n20971 , n20972 , n20973 , n20974 , n20975 , n20976 , n20977 , n20978 , n20979 , n20980 , n20981 , n20982 , n20983 , n20984 , n20985 , n20986 , n20987 , n20988 , n20989 , n20990 , n20991 , n20992 , n20993 , n20994 , n20995 , n20996 , n20997 , n20998 , n20999 , n21000 , n21001 , n21002 , n21003 , n21004 , n21005 , n21006 , n21007 , n21008 , n21009 , n21010 , n21011 , n21012 , n21013 , n21014 , n21015 , n21016 , n21017 , n21018 , n21019 , n21020 , n21021 , n21022 , n21023 , n21024 , n21025 , n21026 , n21027 , n21028 , n21029 , n21030 , n21031 , n21032 , n21033 , n21034 , n21035 , n21036 , n21037 , n21038 , n21039 , n21040 , n21041 , n21042 , n21043 , n21044 , n21045 , n21046 , n21047 , n21048 , n21049 , n21050 , n21051 , n21052 , n21053 , n21054 , n21055 , n21056 , n21057 , n21058 , n21059 , n21060 , n21061 , n21062 , n21063 , n21064 , n21065 , n21066 , n21067 , n21068 , n21069 , n21070 , n21071 , n21072 , n21073 , n21074 , n21075 , n21076 , n21077 , n21078 , n21079 , n21080 , n21081 , n21082 , n21083 , n21084 ;
  assign n65 = x0 & x1 ;
  assign n66 = x1 & ~n65 ;
  assign n67 = x0 & x2 ;
  assign n68 = n65 & n67 ;
  assign n69 = n65 | n67 ;
  assign n70 = ~n68 & n69 ;
  assign n71 = x0 & x3 ;
  assign n72 = x1 & x2 ;
  assign n73 = x2 & ~n72 ;
  assign n74 = ( n68 & n71 ) | ( n68 & ~n73 ) | ( n71 & ~n73 ) ;
  assign n75 = ( ~n68 & n73 ) | ( ~n68 & n74 ) | ( n73 & n74 ) ;
  assign n76 = ( ~n71 & n74 ) | ( ~n71 & n75 ) | ( n74 & n75 ) ;
  assign n77 = x2 & x3 ;
  assign n78 = x0 & n77 ;
  assign n79 = x3 & x4 ;
  assign n80 = n65 & n79 ;
  assign n81 = x1 & x3 ;
  assign n82 = x0 & x4 ;
  assign n83 = n81 | n82 ;
  assign n84 = ~n80 & n83 ;
  assign n85 = ( n72 & n78 ) | ( n72 & ~n84 ) | ( n78 & ~n84 ) ;
  assign n86 = ( ~n72 & n84 ) | ( ~n72 & n85 ) | ( n84 & n85 ) ;
  assign n87 = ( ~n78 & n85 ) | ( ~n78 & n86 ) | ( n85 & n86 ) ;
  assign n88 = x1 & x4 ;
  assign n89 = x0 & x5 ;
  assign n90 = n88 | n89 ;
  assign n91 = x4 & x5 ;
  assign n92 = n65 & n91 ;
  assign n93 = n90 & ~n92 ;
  assign n94 = n80 | n92 ;
  assign n95 = ( n92 & n93 ) | ( n92 & n94 ) | ( n93 & n94 ) ;
  assign n96 = n90 & ~n95 ;
  assign n97 = x3 & ~n77 ;
  assign n98 = n80 & n97 ;
  assign n99 = ~n93 & n98 ;
  assign n100 = ( n96 & n97 ) | ( n96 & n99 ) | ( n97 & n99 ) ;
  assign n101 = n80 | n97 ;
  assign n102 = ( ~n93 & n97 ) | ( ~n93 & n101 ) | ( n97 & n101 ) ;
  assign n103 = n96 | n102 ;
  assign n104 = ~n100 & n103 ;
  assign n105 = n72 & n84 ;
  assign n106 = n72 & n78 ;
  assign n107 = ( n78 & n84 ) | ( n78 & n106 ) | ( n84 & n106 ) ;
  assign n108 = n105 | n107 ;
  assign n109 = n104 | n108 ;
  assign n110 = n104 & n108 ;
  assign n111 = n109 & ~n110 ;
  assign n112 = x0 & x6 ;
  assign n113 = n77 & n112 ;
  assign n114 = n77 & ~n113 ;
  assign n115 = n112 & ~n113 ;
  assign n116 = n114 | n115 ;
  assign n117 = n72 & n91 ;
  assign n118 = x1 & x5 ;
  assign n119 = x2 & x4 ;
  assign n120 = n118 | n119 ;
  assign n121 = ~n117 & n120 ;
  assign n122 = n116 | n121 ;
  assign n123 = n116 & n121 ;
  assign n124 = n122 & ~n123 ;
  assign n125 = n95 | n124 ;
  assign n126 = n95 & n124 ;
  assign n127 = n125 | n126 ;
  assign n128 = n103 & n108 ;
  assign n129 = n100 | n128 ;
  assign n130 = ( n126 & ~n127 ) | ( n126 & n129 ) | ( ~n127 & n129 ) ;
  assign n131 = ( n126 & n127 ) | ( n126 & n129 ) | ( n127 & n129 ) ;
  assign n132 = ( n127 & n130 ) | ( n127 & ~n131 ) | ( n130 & ~n131 ) ;
  assign n133 = x0 & x7 ;
  assign n134 = n79 & n133 ;
  assign n135 = x5 & x7 ;
  assign n136 = n67 & n135 ;
  assign n137 = n134 | n136 ;
  assign n138 = n77 & n91 ;
  assign n139 = n133 & n138 ;
  assign n140 = ( n133 & ~n137 ) | ( n133 & n139 ) | ( ~n137 & n139 ) ;
  assign n141 = n137 | n138 ;
  assign n142 = x2 & x5 ;
  assign n143 = ( n79 & ~n138 ) | ( n79 & n142 ) | ( ~n138 & n142 ) ;
  assign n144 = n79 & n142 ;
  assign n145 = ( ~n137 & n143 ) | ( ~n137 & n144 ) | ( n143 & n144 ) ;
  assign n146 = ~n141 & n145 ;
  assign n147 = n140 | n146 ;
  assign n148 = x1 & x6 ;
  assign n149 = n117 & ~n148 ;
  assign n150 = n117 & ~n149 ;
  assign n151 = x4 & n148 ;
  assign n152 = x4 | n148 ;
  assign n153 = ( ~n117 & n148 ) | ( ~n117 & n152 ) | ( n148 & n152 ) ;
  assign n154 = ( n150 & ~n151 ) | ( n150 & n153 ) | ( ~n151 & n153 ) ;
  assign n155 = n113 | n121 ;
  assign n156 = ( n113 & n116 ) | ( n113 & n155 ) | ( n116 & n155 ) ;
  assign n157 = n154 & n156 ;
  assign n158 = n154 | n156 ;
  assign n159 = ~n157 & n158 ;
  assign n160 = ( n131 & n147 ) | ( n131 & ~n159 ) | ( n147 & ~n159 ) ;
  assign n161 = ( ~n147 & n159 ) | ( ~n147 & n160 ) | ( n159 & n160 ) ;
  assign n162 = ( ~n131 & n160 ) | ( ~n131 & n161 ) | ( n160 & n161 ) ;
  assign n163 = n147 & n159 ;
  assign n164 = n147 | n159 ;
  assign n165 = n163 | n164 ;
  assign n166 = ( n131 & n163 ) | ( n131 & n165 ) | ( n163 & n165 ) ;
  assign n167 = n149 | n157 ;
  assign n168 = x1 & x7 ;
  assign n169 = x3 & x5 ;
  assign n170 = n168 & n169 ;
  assign n171 = n168 & ~n170 ;
  assign n172 = n169 & ~n170 ;
  assign n173 = n171 | n172 ;
  assign n174 = n141 & n173 ;
  assign n175 = n141 & ~n174 ;
  assign n176 = n173 & ~n174 ;
  assign n177 = n175 | n176 ;
  assign n178 = x0 & x8 ;
  assign n179 = x2 & x6 ;
  assign n180 = n178 | n179 ;
  assign n181 = x6 & x8 ;
  assign n182 = n67 & n181 ;
  assign n183 = n180 & ~n182 ;
  assign n184 = n151 | n182 ;
  assign n185 = ( n182 & n183 ) | ( n182 & n184 ) | ( n183 & n184 ) ;
  assign n186 = n180 & ~n185 ;
  assign n187 = n151 & ~n183 ;
  assign n188 = n186 | n187 ;
  assign n189 = n177 & n188 ;
  assign n190 = n177 | n188 ;
  assign n191 = ~n189 & n190 ;
  assign n192 = ( n166 & n167 ) | ( n166 & ~n191 ) | ( n167 & ~n191 ) ;
  assign n193 = ( ~n167 & n191 ) | ( ~n167 & n192 ) | ( n191 & n192 ) ;
  assign n194 = ( ~n166 & n192 ) | ( ~n166 & n193 ) | ( n192 & n193 ) ;
  assign n195 = n167 & n191 ;
  assign n196 = n167 | n191 ;
  assign n197 = n166 & n196 ;
  assign n198 = n195 | n197 ;
  assign n199 = n119 & n135 ;
  assign n200 = x6 & x7 ;
  assign n201 = n77 & n200 ;
  assign n202 = n199 | n201 ;
  assign n203 = x2 & x7 ;
  assign n204 = x5 & x6 ;
  assign n205 = n79 & n204 ;
  assign n206 = n203 & n205 ;
  assign n207 = ( ~n202 & n203 ) | ( ~n202 & n206 ) | ( n203 & n206 ) ;
  assign n208 = n202 | n205 ;
  assign n209 = x3 & x6 ;
  assign n210 = ( n91 & ~n205 ) | ( n91 & n209 ) | ( ~n205 & n209 ) ;
  assign n211 = n91 & n209 ;
  assign n212 = ( ~n202 & n210 ) | ( ~n202 & n211 ) | ( n210 & n211 ) ;
  assign n213 = ~n208 & n212 ;
  assign n214 = n207 | n213 ;
  assign n215 = n185 & n207 ;
  assign n216 = ( n185 & n213 ) | ( n185 & n215 ) | ( n213 & n215 ) ;
  assign n217 = n214 & ~n216 ;
  assign n218 = x0 & x9 ;
  assign n219 = n170 & ~n218 ;
  assign n220 = ~n170 & n218 ;
  assign n221 = n219 | n220 ;
  assign n222 = x5 & x8 ;
  assign n223 = x1 & x8 ;
  assign n224 = ~n222 & n223 ;
  assign n225 = ~x1 & x5 ;
  assign n226 = ( x5 & ~n222 ) | ( x5 & n225 ) | ( ~n222 & n225 ) ;
  assign n227 = n224 | n226 ;
  assign n228 = n221 & n227 ;
  assign n229 = n221 | n227 ;
  assign n230 = ~n228 & n229 ;
  assign n231 = n185 & ~n207 ;
  assign n232 = ~n213 & n231 ;
  assign n233 = n230 & n232 ;
  assign n234 = ( n217 & n230 ) | ( n217 & n233 ) | ( n230 & n233 ) ;
  assign n235 = n230 | n232 ;
  assign n236 = n217 | n235 ;
  assign n237 = ~n234 & n236 ;
  assign n238 = n174 | n188 ;
  assign n239 = ( n174 & n177 ) | ( n174 & n238 ) | ( n177 & n238 ) ;
  assign n240 = ( n198 & n237 ) | ( n198 & ~n239 ) | ( n237 & ~n239 ) ;
  assign n241 = ( ~n237 & n239 ) | ( ~n237 & n240 ) | ( n239 & n240 ) ;
  assign n242 = ( ~n198 & n240 ) | ( ~n198 & n241 ) | ( n240 & n241 ) ;
  assign n243 = n237 & n239 ;
  assign n244 = n237 | n239 ;
  assign n245 = n195 & n244 ;
  assign n246 = ( n197 & n244 ) | ( n197 & n245 ) | ( n244 & n245 ) ;
  assign n247 = n243 | n246 ;
  assign n248 = n216 | n234 ;
  assign n249 = x8 & x10 ;
  assign n250 = n67 & n249 ;
  assign n251 = x7 & x8 ;
  assign n252 = n77 & n251 ;
  assign n253 = n250 | n252 ;
  assign n254 = x0 & x10 ;
  assign n255 = x3 & x7 ;
  assign n256 = n254 & n255 ;
  assign n257 = x2 & n256 ;
  assign n258 = ( x2 & ~n253 ) | ( x2 & n257 ) | ( ~n253 & n257 ) ;
  assign n259 = x8 & n258 ;
  assign n260 = ( n170 & n218 ) | ( n170 & n227 ) | ( n218 & n227 ) ;
  assign n261 = ( ~n253 & n254 ) | ( ~n253 & n255 ) | ( n254 & n255 ) ;
  assign n262 = ~n260 & n261 ;
  assign n263 = n170 | n256 ;
  assign n264 = n218 | n256 ;
  assign n265 = ( n227 & n263 ) | ( n227 & n264 ) | ( n263 & n264 ) ;
  assign n266 = ( n259 & n262 ) | ( n259 & ~n265 ) | ( n262 & ~n265 ) ;
  assign n267 = n260 & ~n261 ;
  assign n268 = n170 & n256 ;
  assign n269 = n218 & n256 ;
  assign n270 = ( n227 & n268 ) | ( n227 & n269 ) | ( n268 & n269 ) ;
  assign n271 = ( ~n259 & n267 ) | ( ~n259 & n270 ) | ( n267 & n270 ) ;
  assign n272 = n266 | n271 ;
  assign n273 = x1 & x9 ;
  assign n274 = x4 & x6 ;
  assign n275 = n273 | n274 ;
  assign n276 = x4 & x9 ;
  assign n277 = n148 & n276 ;
  assign n278 = n275 & ~n277 ;
  assign n279 = x1 & n222 ;
  assign n280 = n278 & n279 ;
  assign n281 = n278 & ~n280 ;
  assign n282 = ~n278 & n279 ;
  assign n283 = n208 & n282 ;
  assign n284 = ( n208 & n281 ) | ( n208 & n283 ) | ( n281 & n283 ) ;
  assign n285 = n208 | n282 ;
  assign n286 = n281 | n285 ;
  assign n287 = ~n284 & n286 ;
  assign n288 = n272 & n287 ;
  assign n289 = n272 | n287 ;
  assign n290 = ~n288 & n289 ;
  assign n291 = n248 | n290 ;
  assign n292 = n248 & n290 ;
  assign n293 = n291 & ~n292 ;
  assign n294 = n247 | n293 ;
  assign n295 = n243 & n291 ;
  assign n296 = ( n246 & n291 ) | ( n246 & n295 ) | ( n291 & n295 ) ;
  assign n297 = ~n292 & n296 ;
  assign n298 = n294 & ~n297 ;
  assign n299 = n253 | n256 ;
  assign n300 = x1 & ~x10 ;
  assign n301 = ( x1 & ~n148 ) | ( x1 & n300 ) | ( ~n148 & n300 ) ;
  assign n302 = x10 & n301 ;
  assign n303 = x6 & ~x10 ;
  assign n304 = ( x6 & ~n148 ) | ( x6 & n303 ) | ( ~n148 & n303 ) ;
  assign n305 = n302 | n304 ;
  assign n306 = n299 & n305 ;
  assign n307 = n299 & ~n306 ;
  assign n308 = n305 & ~n306 ;
  assign n309 = n307 | n308 ;
  assign n310 = x2 & x9 ;
  assign n311 = x3 & x8 ;
  assign n312 = n310 | n311 ;
  assign n313 = x8 & x9 ;
  assign n314 = n77 & n313 ;
  assign n315 = n312 & ~n314 ;
  assign n316 = n277 | n314 ;
  assign n317 = ( n314 & n315 ) | ( n314 & n316 ) | ( n315 & n316 ) ;
  assign n318 = n312 & ~n317 ;
  assign n319 = n277 & ~n315 ;
  assign n320 = n318 | n319 ;
  assign n321 = ~n309 & n320 ;
  assign n322 = n309 & ~n320 ;
  assign n323 = n321 | n322 ;
  assign n324 = n280 | n284 ;
  assign n325 = x4 & x7 ;
  assign n326 = n204 | n325 ;
  assign n327 = n91 & n200 ;
  assign n328 = n326 & ~n327 ;
  assign n329 = x0 & x11 ;
  assign n330 = n327 | n329 ;
  assign n331 = ( n327 & n328 ) | ( n327 & n330 ) | ( n328 & n330 ) ;
  assign n332 = n326 & ~n331 ;
  assign n333 = ~n328 & n329 ;
  assign n334 = n332 | n333 ;
  assign n335 = n324 & n334 ;
  assign n336 = n324 & ~n335 ;
  assign n337 = ~n324 & n334 ;
  assign n338 = n336 | n337 ;
  assign n339 = n323 & n338 ;
  assign n340 = ( ~n323 & n336 ) | ( ~n323 & n337 ) | ( n336 & n337 ) ;
  assign n341 = n323 | n340 ;
  assign n342 = ~n339 & n341 ;
  assign n343 = ( ~n256 & n259 ) | ( ~n256 & n261 ) | ( n259 & n261 ) ;
  assign n344 = ( n260 & n287 ) | ( n260 & n343 ) | ( n287 & n343 ) ;
  assign n345 = n342 | n344 ;
  assign n346 = n342 & n344 ;
  assign n347 = n345 | n346 ;
  assign n348 = n292 | n295 ;
  assign n349 = n291 | n292 ;
  assign n350 = ( n246 & n348 ) | ( n246 & n349 ) | ( n348 & n349 ) ;
  assign n351 = ( n346 & ~n347 ) | ( n346 & n350 ) | ( ~n347 & n350 ) ;
  assign n352 = ( n342 & n344 ) | ( n342 & n350 ) | ( n344 & n350 ) ;
  assign n353 = ( n347 & n351 ) | ( n347 & ~n352 ) | ( n351 & ~n352 ) ;
  assign n354 = n317 | n331 ;
  assign n355 = n317 & n331 ;
  assign n356 = n354 & ~n355 ;
  assign n357 = x3 & x9 ;
  assign n358 = x0 & x12 ;
  assign n359 = n357 & n358 ;
  assign n360 = x9 & x10 ;
  assign n361 = n77 & n360 ;
  assign n362 = n359 | n361 ;
  assign n363 = x10 & x12 ;
  assign n364 = n67 & n363 ;
  assign n365 = n357 & n364 ;
  assign n366 = ( n357 & ~n362 ) | ( n357 & n365 ) | ( ~n362 & n365 ) ;
  assign n367 = n362 | n364 ;
  assign n368 = x2 & x10 ;
  assign n369 = ( n358 & ~n364 ) | ( n358 & n368 ) | ( ~n364 & n368 ) ;
  assign n370 = n358 & n368 ;
  assign n371 = ( ~n362 & n369 ) | ( ~n362 & n370 ) | ( n369 & n370 ) ;
  assign n372 = ~n367 & n371 ;
  assign n373 = n366 | n372 ;
  assign n374 = ~n356 & n373 ;
  assign n375 = n356 & ~n373 ;
  assign n376 = n374 | n375 ;
  assign n377 = x5 & x11 ;
  assign n378 = n168 & n377 ;
  assign n379 = x1 & x11 ;
  assign n380 = n135 | n379 ;
  assign n381 = ~n378 & n380 ;
  assign n382 = x10 & n148 ;
  assign n383 = x4 & x8 ;
  assign n384 = n382 & n383 ;
  assign n385 = n381 & ~n384 ;
  assign n386 = n382 | n383 ;
  assign n387 = n381 & ~n386 ;
  assign n388 = ( n381 & ~n385 ) | ( n381 & n387 ) | ( ~n385 & n387 ) ;
  assign n389 = ~n382 & n386 ;
  assign n390 = n382 & ~n383 ;
  assign n391 = ( ~n385 & n389 ) | ( ~n385 & n390 ) | ( n389 & n390 ) ;
  assign n392 = n388 | n391 ;
  assign n393 = n306 | n320 ;
  assign n394 = ( n306 & n309 ) | ( n306 & n393 ) | ( n309 & n393 ) ;
  assign n395 = n392 & n394 ;
  assign n396 = n392 | n394 ;
  assign n397 = ~n395 & n396 ;
  assign n398 = n376 & n397 ;
  assign n399 = n376 | n397 ;
  assign n400 = ~n398 & n399 ;
  assign n401 = n323 | n335 ;
  assign n402 = ( n335 & n338 ) | ( n335 & n401 ) | ( n338 & n401 ) ;
  assign n403 = ( n352 & ~n400 ) | ( n352 & n402 ) | ( ~n400 & n402 ) ;
  assign n404 = ( n400 & ~n402 ) | ( n400 & n403 ) | ( ~n402 & n403 ) ;
  assign n405 = ( ~n352 & n403 ) | ( ~n352 & n404 ) | ( n403 & n404 ) ;
  assign n406 = n400 & n402 ;
  assign n407 = n400 | n402 ;
  assign n408 = n406 | n407 ;
  assign n409 = ( n352 & n406 ) | ( n352 & n408 ) | ( n406 & n408 ) ;
  assign n410 = ( n382 & n383 ) | ( n382 & n385 ) | ( n383 & n385 ) ;
  assign n411 = n79 & n360 ;
  assign n412 = x3 & x13 ;
  assign n413 = n254 & n412 ;
  assign n414 = n411 | n413 ;
  assign n415 = x9 & x13 ;
  assign n416 = n82 & n415 ;
  assign n417 = x3 & n416 ;
  assign n418 = ( x3 & ~n414 ) | ( x3 & n417 ) | ( ~n414 & n417 ) ;
  assign n419 = x10 & n418 ;
  assign n420 = n414 | n416 ;
  assign n421 = x0 & x13 ;
  assign n422 = ( n276 & ~n416 ) | ( n276 & n421 ) | ( ~n416 & n421 ) ;
  assign n423 = n276 & n421 ;
  assign n424 = ( ~n414 & n422 ) | ( ~n414 & n423 ) | ( n422 & n423 ) ;
  assign n425 = ~n420 & n424 ;
  assign n426 = n419 | n425 ;
  assign n427 = ~n410 & n426 ;
  assign n428 = n410 & ~n426 ;
  assign n429 = n427 | n428 ;
  assign n430 = n200 | n222 ;
  assign n431 = n204 & n251 ;
  assign n432 = x2 & x11 ;
  assign n433 = ~n431 & n432 ;
  assign n434 = n430 | n431 ;
  assign n435 = ( n431 & n433 ) | ( n431 & n434 ) | ( n433 & n434 ) ;
  assign n436 = n430 & ~n435 ;
  assign n437 = ~n430 & n432 ;
  assign n438 = ( n432 & ~n433 ) | ( n432 & n437 ) | ( ~n433 & n437 ) ;
  assign n439 = n436 | n438 ;
  assign n440 = n429 & n439 ;
  assign n441 = n429 | n439 ;
  assign n442 = ~n440 & n441 ;
  assign n443 = ~x12 & n378 ;
  assign n444 = ( x1 & x12 ) | ( x1 & n378 ) | ( x12 & n378 ) ;
  assign n445 = ( x7 & n378 ) | ( x7 & ~n444 ) | ( n378 & ~n444 ) ;
  assign n446 = ~x7 & x12 ;
  assign n447 = x1 & ~x7 ;
  assign n448 = ( n378 & n446 ) | ( n378 & n447 ) | ( n446 & n447 ) ;
  assign n449 = ( ~n443 & n445 ) | ( ~n443 & n448 ) | ( n445 & n448 ) ;
  assign n450 = n367 & n449 ;
  assign n451 = n367 | n449 ;
  assign n452 = ~n450 & n451 ;
  assign n453 = n356 & n373 ;
  assign n454 = n355 | n453 ;
  assign n455 = n452 | n454 ;
  assign n456 = n452 & n454 ;
  assign n457 = n455 & ~n456 ;
  assign n458 = n376 | n395 ;
  assign n459 = ( n395 & n397 ) | ( n395 & n458 ) | ( n397 & n458 ) ;
  assign n460 = n457 | n459 ;
  assign n461 = n457 & n459 ;
  assign n462 = n460 & ~n461 ;
  assign n463 = ( n409 & n442 ) | ( n409 & ~n462 ) | ( n442 & ~n462 ) ;
  assign n464 = ( ~n442 & n462 ) | ( ~n442 & n463 ) | ( n462 & n463 ) ;
  assign n465 = ( ~n409 & n463 ) | ( ~n409 & n464 ) | ( n463 & n464 ) ;
  assign n466 = x1 & x13 ;
  assign n467 = n181 | n466 ;
  assign n468 = n181 & n466 ;
  assign n469 = n467 & ~n468 ;
  assign n470 = n435 & n469 ;
  assign n471 = n435 & ~n470 ;
  assign n472 = ( n469 & ~n470 ) | ( n469 & n471 ) | ( ~n470 & n471 ) ;
  assign n473 = ~n420 & n470 ;
  assign n474 = n420 | n469 ;
  assign n475 = ( n471 & ~n473 ) | ( n471 & n474 ) | ( ~n473 & n474 ) ;
  assign n476 = ~n472 & n475 ;
  assign n477 = ( n410 & n426 ) | ( n410 & n439 ) | ( n426 & n439 ) ;
  assign n478 = n475 | n477 ;
  assign n479 = n420 & ~n477 ;
  assign n480 = ( n476 & n478 ) | ( n476 & ~n479 ) | ( n478 & ~n479 ) ;
  assign n481 = n475 & n477 ;
  assign n482 = ~n420 & n477 ;
  assign n483 = ( n476 & n481 ) | ( n476 & n482 ) | ( n481 & n482 ) ;
  assign n484 = n480 & ~n483 ;
  assign n485 = x3 & x14 ;
  assign n486 = n329 & n485 ;
  assign n487 = x12 & x14 ;
  assign n488 = n67 & n487 ;
  assign n489 = n486 | n488 ;
  assign n490 = x11 & x12 ;
  assign n491 = n77 & n490 ;
  assign n492 = x14 & n491 ;
  assign n493 = ( x14 & ~n489 ) | ( x14 & n492 ) | ( ~n489 & n492 ) ;
  assign n494 = x0 & n493 ;
  assign n495 = n489 | n491 ;
  assign n496 = x2 & x12 ;
  assign n497 = x3 & x11 ;
  assign n498 = ( ~n491 & n496 ) | ( ~n491 & n497 ) | ( n496 & n497 ) ;
  assign n499 = n496 & n497 ;
  assign n500 = ( ~n489 & n498 ) | ( ~n489 & n499 ) | ( n498 & n499 ) ;
  assign n501 = ~n495 & n500 ;
  assign n502 = n494 | n501 ;
  assign n503 = x4 & x10 ;
  assign n504 = x5 & x9 ;
  assign n505 = n503 | n504 ;
  assign n506 = n91 & n360 ;
  assign n507 = n505 & ~n506 ;
  assign n508 = x12 & n168 ;
  assign n509 = n506 | n508 ;
  assign n510 = ( n506 & n507 ) | ( n506 & n509 ) | ( n507 & n509 ) ;
  assign n511 = n505 & ~n510 ;
  assign n512 = ~n507 & n508 ;
  assign n513 = n511 | n512 ;
  assign n514 = n502 & n513 ;
  assign n515 = n502 & ~n514 ;
  assign n516 = n513 & ~n514 ;
  assign n517 = n515 | n516 ;
  assign n518 = n367 | n443 ;
  assign n519 = ( n443 & n449 ) | ( n443 & n518 ) | ( n449 & n518 ) ;
  assign n520 = n517 | n519 ;
  assign n521 = n517 & n519 ;
  assign n522 = n520 & ~n521 ;
  assign n523 = n484 & ~n522 ;
  assign n524 = ~n484 & n522 ;
  assign n525 = n523 | n524 ;
  assign n526 = n456 | n457 ;
  assign n527 = ( n456 & n459 ) | ( n456 & n526 ) | ( n459 & n526 ) ;
  assign n528 = n525 & n527 ;
  assign n529 = n525 | n527 ;
  assign n530 = ~n528 & n529 ;
  assign n531 = n442 & n462 ;
  assign n532 = n442 | n462 ;
  assign n533 = n531 | n532 ;
  assign n534 = ( n409 & n531 ) | ( n409 & n533 ) | ( n531 & n533 ) ;
  assign n535 = n530 | n534 ;
  assign n536 = n529 & n534 ;
  assign n537 = ~n528 & n536 ;
  assign n538 = n535 & ~n537 ;
  assign n539 = x1 & x14 ;
  assign n540 = x8 & n539 ;
  assign n541 = x8 & ~n539 ;
  assign n542 = ( n539 & ~n540 ) | ( n539 & n541 ) | ( ~n540 & n541 ) ;
  assign n543 = x4 & x11 ;
  assign n544 = n468 & n543 ;
  assign n545 = n542 & ~n544 ;
  assign n546 = n468 | n543 ;
  assign n547 = n542 & ~n546 ;
  assign n548 = ( n542 & ~n545 ) | ( n542 & n547 ) | ( ~n545 & n547 ) ;
  assign n549 = ~n468 & n546 ;
  assign n550 = n468 & ~n543 ;
  assign n551 = ( ~n545 & n549 ) | ( ~n545 & n550 ) | ( n549 & n550 ) ;
  assign n552 = n548 | n551 ;
  assign n553 = x6 & x9 ;
  assign n554 = n251 | n553 ;
  assign n555 = x2 & x13 ;
  assign n556 = ( n251 & n553 ) | ( n251 & n555 ) | ( n553 & n555 ) ;
  assign n557 = n554 & ~n556 ;
  assign n558 = n251 & n553 ;
  assign n559 = n555 & ~n558 ;
  assign n560 = ~n554 & n555 ;
  assign n561 = ( n555 & ~n559 ) | ( n555 & n560 ) | ( ~n559 & n560 ) ;
  assign n562 = n557 | n561 ;
  assign n563 = n552 & n562 ;
  assign n564 = n552 & ~n563 ;
  assign n565 = n420 & ~n470 ;
  assign n566 = n420 & n469 ;
  assign n567 = ( n471 & n565 ) | ( n471 & n566 ) | ( n565 & n566 ) ;
  assign n568 = n470 | n567 ;
  assign n569 = ~n552 & n562 ;
  assign n570 = n568 & n569 ;
  assign n571 = ( n564 & n568 ) | ( n564 & n570 ) | ( n568 & n570 ) ;
  assign n572 = n568 | n569 ;
  assign n573 = n564 | n572 ;
  assign n574 = ~n571 & n573 ;
  assign n575 = n495 | n510 ;
  assign n576 = n495 & n510 ;
  assign n577 = n575 & ~n576 ;
  assign n578 = x0 & x15 ;
  assign n579 = x3 & x12 ;
  assign n580 = n578 & n579 ;
  assign n581 = x5 & x10 ;
  assign n582 = x10 & x15 ;
  assign n583 = x0 & n582 ;
  assign n584 = x3 & n363 ;
  assign n585 = n583 | n584 ;
  assign n586 = x5 & ~n580 ;
  assign n587 = n585 & n586 ;
  assign n588 = n581 & ~n587 ;
  assign n589 = ( n578 & n579 ) | ( n578 & ~n587 ) | ( n579 & ~n587 ) ;
  assign n590 = ( ~n580 & n588 ) | ( ~n580 & n589 ) | ( n588 & n589 ) ;
  assign n591 = n577 & n590 ;
  assign n592 = n577 & ~n591 ;
  assign n593 = n590 & ~n591 ;
  assign n594 = n592 | n593 ;
  assign n595 = n514 | n519 ;
  assign n596 = ( n514 & n517 ) | ( n514 & n595 ) | ( n517 & n595 ) ;
  assign n597 = n594 | n596 ;
  assign n598 = n594 & n596 ;
  assign n599 = n597 & ~n598 ;
  assign n600 = n574 & ~n599 ;
  assign n601 = ~n574 & n599 ;
  assign n602 = n600 | n601 ;
  assign n603 = ( ~n420 & n475 ) | ( ~n420 & n476 ) | ( n475 & n476 ) ;
  assign n604 = ( n477 & n522 ) | ( n477 & n603 ) | ( n522 & n603 ) ;
  assign n605 = n602 & n604 ;
  assign n606 = n602 | n604 ;
  assign n607 = ~n605 & n606 ;
  assign n608 = n528 | n529 ;
  assign n609 = ( n528 & n534 ) | ( n528 & n608 ) | ( n534 & n608 ) ;
  assign n610 = ~n607 & n609 ;
  assign n611 = n607 & ~n609 ;
  assign n612 = n610 | n611 ;
  assign n686 = ( n602 & n604 ) | ( n602 & n608 ) | ( n604 & n608 ) ;
  assign n687 = ( n528 & n602 ) | ( n528 & n604 ) | ( n602 & n604 ) ;
  assign n688 = ( n534 & n686 ) | ( n534 & n687 ) | ( n686 & n687 ) ;
  assign n613 = ( n468 & n543 ) | ( n468 & n545 ) | ( n543 & n545 ) ;
  assign n614 = n580 | n587 ;
  assign n615 = n613 | n614 ;
  assign n616 = n613 & n614 ;
  assign n617 = n615 & ~n616 ;
  assign n618 = x10 & x11 ;
  assign n619 = n204 & n618 ;
  assign n620 = x0 & x16 ;
  assign n621 = n377 & n620 ;
  assign n622 = n619 | n621 ;
  assign n623 = x6 & x16 ;
  assign n624 = n254 & n623 ;
  assign n625 = n377 & n624 ;
  assign n626 = ( n377 & ~n622 ) | ( n377 & n625 ) | ( ~n622 & n625 ) ;
  assign n627 = n622 | n624 ;
  assign n628 = x6 & x10 ;
  assign n629 = ( n620 & ~n624 ) | ( n620 & n628 ) | ( ~n624 & n628 ) ;
  assign n630 = n620 & n628 ;
  assign n631 = ( ~n622 & n629 ) | ( ~n622 & n630 ) | ( n629 & n630 ) ;
  assign n632 = ~n627 & n631 ;
  assign n633 = n626 | n632 ;
  assign n634 = ~n617 & n633 ;
  assign n635 = n616 | n633 ;
  assign n636 = n615 & ~n635 ;
  assign n637 = n634 | n636 ;
  assign n638 = n563 | n568 ;
  assign n639 = n563 | n564 ;
  assign n640 = ( n570 & n638 ) | ( n570 & n639 ) | ( n638 & n639 ) ;
  assign n641 = n637 | n640 ;
  assign n642 = n637 & n640 ;
  assign n643 = n641 & ~n642 ;
  assign n644 = n576 | n591 ;
  assign n645 = x4 & x12 ;
  assign n646 = n119 & n487 ;
  assign n647 = x12 & x13 ;
  assign n648 = n79 & n647 ;
  assign n649 = n646 | n648 ;
  assign n650 = x13 & x14 ;
  assign n651 = n77 & n650 ;
  assign n652 = n645 & n651 ;
  assign n653 = ( n645 & ~n649 ) | ( n645 & n652 ) | ( ~n649 & n652 ) ;
  assign n654 = n649 | n651 ;
  assign n655 = x2 & x14 ;
  assign n656 = ( n412 & ~n651 ) | ( n412 & n655 ) | ( ~n651 & n655 ) ;
  assign n657 = n412 & n655 ;
  assign n658 = ( ~n649 & n656 ) | ( ~n649 & n657 ) | ( n656 & n657 ) ;
  assign n659 = ~n654 & n658 ;
  assign n660 = n653 | n659 ;
  assign n661 = n576 & n660 ;
  assign n662 = ( n591 & n660 ) | ( n591 & n661 ) | ( n660 & n661 ) ;
  assign n663 = n644 & ~n662 ;
  assign n664 = n660 & ~n661 ;
  assign n665 = ~n591 & n664 ;
  assign n666 = n663 | n665 ;
  assign n667 = x7 & x9 ;
  assign n668 = x1 & x15 ;
  assign n669 = n667 & n668 ;
  assign n670 = n667 | n668 ;
  assign n671 = ~n669 & n670 ;
  assign n672 = ~n540 & n671 ;
  assign n673 = n540 & ~n671 ;
  assign n674 = n672 | n673 ;
  assign n675 = n556 & ~n674 ;
  assign n676 = n556 & n674 ;
  assign n677 = n674 & ~n676 ;
  assign n678 = n675 | n677 ;
  assign n679 = n666 & n678 ;
  assign n680 = n666 | n678 ;
  assign n681 = ~n679 & n680 ;
  assign n682 = n643 | n681 ;
  assign n683 = n643 & n681 ;
  assign n684 = n682 & ~n683 ;
  assign n685 = ( n574 & n594 ) | ( n574 & n596 ) | ( n594 & n596 ) ;
  assign n689 = ( n684 & ~n685 ) | ( n684 & n688 ) | ( ~n685 & n688 ) ;
  assign n690 = ( ~n684 & n685 ) | ( ~n684 & n689 ) | ( n685 & n689 ) ;
  assign n691 = ( ~n688 & n689 ) | ( ~n688 & n690 ) | ( n689 & n690 ) ;
  assign n692 = n684 & n685 ;
  assign n693 = n684 | n685 ;
  assign n694 = n692 | n693 ;
  assign n695 = ( n688 & n692 ) | ( n688 & n694 ) | ( n692 & n694 ) ;
  assign n696 = x7 & x10 ;
  assign n697 = n313 | n696 ;
  assign n698 = n251 & n360 ;
  assign n699 = n485 & ~n698 ;
  assign n700 = n697 | n698 ;
  assign n701 = ( n698 & n699 ) | ( n698 & n700 ) | ( n699 & n700 ) ;
  assign n702 = n697 & ~n701 ;
  assign n703 = n485 & ~n697 ;
  assign n704 = ( n485 & ~n699 ) | ( n485 & n703 ) | ( ~n699 & n703 ) ;
  assign n705 = n702 | n704 ;
  assign n706 = x5 & x12 ;
  assign n707 = x0 & x17 ;
  assign n708 = n706 | n707 ;
  assign n709 = ( n669 & n706 ) | ( n669 & n707 ) | ( n706 & n707 ) ;
  assign n710 = n708 & ~n709 ;
  assign n711 = n706 & n707 ;
  assign n712 = n708 & ~n711 ;
  assign n713 = n669 & ~n712 ;
  assign n714 = n710 | n713 ;
  assign n715 = n705 & n714 ;
  assign n716 = n705 & ~n715 ;
  assign n717 = x6 & x11 ;
  assign n718 = x11 & x15 ;
  assign n719 = x2 & n718 ;
  assign n720 = x11 & x13 ;
  assign n721 = x4 & n720 ;
  assign n722 = n719 | n721 ;
  assign n723 = x13 & x15 ;
  assign n724 = n119 & n723 ;
  assign n725 = x6 & ~n724 ;
  assign n726 = n722 & n725 ;
  assign n727 = n717 & ~n726 ;
  assign n728 = n724 | n726 ;
  assign n729 = x2 & x15 ;
  assign n730 = x4 & x13 ;
  assign n731 = ( ~n724 & n729 ) | ( ~n724 & n730 ) | ( n729 & n730 ) ;
  assign n732 = n729 & n730 ;
  assign n733 = ( ~n726 & n731 ) | ( ~n726 & n732 ) | ( n731 & n732 ) ;
  assign n734 = ~n728 & n733 ;
  assign n735 = n727 | n734 ;
  assign n736 = ~n705 & n714 ;
  assign n737 = n735 & ~n736 ;
  assign n738 = ~n716 & n737 ;
  assign n739 = ~n735 & n736 ;
  assign n740 = ( n716 & ~n735 ) | ( n716 & n739 ) | ( ~n735 & n739 ) ;
  assign n741 = n738 | n740 ;
  assign n742 = n662 | n678 ;
  assign n743 = ( n662 & n666 ) | ( n662 & n742 ) | ( n666 & n742 ) ;
  assign n744 = n741 | n743 ;
  assign n745 = n741 & n743 ;
  assign n746 = n744 & ~n745 ;
  assign n747 = ( n540 & n556 ) | ( n540 & n671 ) | ( n556 & n671 ) ;
  assign n748 = ( n616 & n617 ) | ( n616 & n635 ) | ( n617 & n635 ) ;
  assign n749 = n747 | n748 ;
  assign n750 = n747 & n748 ;
  assign n751 = n749 & ~n750 ;
  assign n752 = x1 & x16 ;
  assign n753 = x9 | n752 ;
  assign n754 = x9 & x16 ;
  assign n755 = x1 & n754 ;
  assign n756 = n651 & ~n755 ;
  assign n757 = ( n649 & ~n755 ) | ( n649 & n756 ) | ( ~n755 & n756 ) ;
  assign n758 = n753 & n757 ;
  assign n759 = n654 & ~n758 ;
  assign n760 = n753 & ~n755 ;
  assign n761 = ~n757 & n760 ;
  assign n762 = n627 & n761 ;
  assign n763 = ( n627 & n759 ) | ( n627 & n762 ) | ( n759 & n762 ) ;
  assign n764 = n627 | n761 ;
  assign n765 = n759 | n764 ;
  assign n766 = ~n763 & n765 ;
  assign n767 = n751 | n766 ;
  assign n768 = n751 & n766 ;
  assign n769 = n767 & ~n768 ;
  assign n770 = n746 & n769 ;
  assign n771 = n746 | n769 ;
  assign n772 = ~n770 & n771 ;
  assign n773 = n642 | n683 ;
  assign n774 = ( n695 & n772 ) | ( n695 & ~n773 ) | ( n772 & ~n773 ) ;
  assign n775 = ( ~n772 & n773 ) | ( ~n772 & n774 ) | ( n773 & n774 ) ;
  assign n776 = ( ~n695 & n774 ) | ( ~n695 & n775 ) | ( n774 & n775 ) ;
  assign n827 = n750 | n766 ;
  assign n828 = ( n750 & n751 ) | ( n750 & n827 ) | ( n751 & n827 ) ;
  assign n777 = x0 & x18 ;
  assign n778 = x5 & x13 ;
  assign n779 = n777 & n778 ;
  assign n780 = x7 & x18 ;
  assign n781 = n329 & n780 ;
  assign n782 = n135 & n720 ;
  assign n783 = n781 | n782 ;
  assign n784 = x11 & n779 ;
  assign n785 = ( x11 & ~n783 ) | ( x11 & n784 ) | ( ~n783 & n784 ) ;
  assign n786 = x7 & n785 ;
  assign n787 = ( n777 & n778 ) | ( n777 & ~n783 ) | ( n778 & ~n783 ) ;
  assign n788 = ( ~n779 & n786 ) | ( ~n779 & n787 ) | ( n786 & n787 ) ;
  assign n789 = x4 & x14 ;
  assign n790 = x14 & x16 ;
  assign n791 = n119 & n790 ;
  assign n792 = x14 & x15 ;
  assign n793 = n79 & n792 ;
  assign n794 = n791 | n793 ;
  assign n795 = x15 & x16 ;
  assign n796 = n77 & n795 ;
  assign n797 = n789 & n796 ;
  assign n798 = ( n789 & ~n794 ) | ( n789 & n797 ) | ( ~n794 & n797 ) ;
  assign n799 = n794 | n796 ;
  assign n800 = x3 & x15 ;
  assign n801 = x2 & x16 ;
  assign n802 = ( ~n796 & n800 ) | ( ~n796 & n801 ) | ( n800 & n801 ) ;
  assign n803 = n800 & n801 ;
  assign n804 = ( ~n794 & n802 ) | ( ~n794 & n803 ) | ( n802 & n803 ) ;
  assign n805 = ~n799 & n804 ;
  assign n806 = n798 | n805 ;
  assign n807 = n788 & n806 ;
  assign n808 = n788 & ~n807 ;
  assign n809 = x6 & x12 ;
  assign n810 = n755 | n809 ;
  assign n811 = n755 & n809 ;
  assign n812 = n810 & ~n811 ;
  assign n813 = x1 & x17 ;
  assign n814 = n249 & n813 ;
  assign n815 = n249 & ~n814 ;
  assign n816 = ~n249 & n813 ;
  assign n817 = n815 | n816 ;
  assign n818 = n812 & n817 ;
  assign n819 = n817 & ~n818 ;
  assign n820 = ( n812 & ~n818 ) | ( n812 & n819 ) | ( ~n818 & n819 ) ;
  assign n821 = ~n788 & n806 ;
  assign n822 = n820 & n821 ;
  assign n823 = ( n808 & n820 ) | ( n808 & n822 ) | ( n820 & n822 ) ;
  assign n824 = n820 | n821 ;
  assign n825 = n808 | n824 ;
  assign n826 = ~n823 & n825 ;
  assign n829 = n826 & n828 ;
  assign n830 = n828 & ~n829 ;
  assign n831 = n826 & ~n828 ;
  assign n832 = n830 | n831 ;
  assign n833 = n701 | n728 ;
  assign n834 = n701 & n728 ;
  assign n835 = n833 & ~n834 ;
  assign n836 = n709 | n835 ;
  assign n837 = n709 & n835 ;
  assign n838 = n836 & ~n837 ;
  assign n839 = n716 | n736 ;
  assign n840 = n758 | n763 ;
  assign n841 = n715 | n735 ;
  assign n842 = n840 & n841 ;
  assign n843 = n715 & n840 ;
  assign n844 = ( n839 & n842 ) | ( n839 & n843 ) | ( n842 & n843 ) ;
  assign n845 = n840 | n841 ;
  assign n846 = n715 | n840 ;
  assign n847 = ( n839 & n845 ) | ( n839 & n846 ) | ( n845 & n846 ) ;
  assign n848 = ~n844 & n847 ;
  assign n849 = n838 & n848 ;
  assign n850 = n838 | n848 ;
  assign n851 = ~n849 & n850 ;
  assign n852 = n832 & n851 ;
  assign n853 = n832 | n851 ;
  assign n854 = ~n852 & n853 ;
  assign n855 = n772 & n773 ;
  assign n856 = ~n692 & n693 ;
  assign n857 = n772 | n773 ;
  assign n858 = ( n692 & n856 ) | ( n692 & n857 ) | ( n856 & n857 ) ;
  assign n859 = n692 & n857 ;
  assign n860 = ( n688 & n858 ) | ( n688 & n859 ) | ( n858 & n859 ) ;
  assign n861 = n855 | n860 ;
  assign n862 = n745 | n769 ;
  assign n863 = ( n745 & n746 ) | ( n745 & n862 ) | ( n746 & n862 ) ;
  assign n864 = ( n854 & ~n861 ) | ( n854 & n863 ) | ( ~n861 & n863 ) ;
  assign n865 = ( n861 & ~n863 ) | ( n861 & n864 ) | ( ~n863 & n864 ) ;
  assign n866 = ( ~n854 & n864 ) | ( ~n854 & n865 ) | ( n864 & n865 ) ;
  assign n867 = n854 & n863 ;
  assign n868 = n854 | n863 ;
  assign n869 = n855 & n868 ;
  assign n870 = ( n860 & n868 ) | ( n860 & n869 ) | ( n868 & n869 ) ;
  assign n871 = n867 | n870 ;
  assign n872 = x1 & x18 ;
  assign n873 = n814 & ~n872 ;
  assign n874 = n814 & ~n873 ;
  assign n875 = x10 | n872 ;
  assign n876 = x10 & n872 ;
  assign n877 = n875 & ~n876 ;
  assign n878 = ~n873 & n877 ;
  assign n879 = n874 | n878 ;
  assign n880 = n799 | n879 ;
  assign n881 = ~n799 & n879 ;
  assign n882 = ( ~n879 & n880 ) | ( ~n879 & n881 ) | ( n880 & n881 ) ;
  assign n883 = n807 & n882 ;
  assign n884 = ( n823 & n882 ) | ( n823 & n883 ) | ( n882 & n883 ) ;
  assign n885 = n807 | n882 ;
  assign n886 = n823 | n885 ;
  assign n887 = ~n884 & n886 ;
  assign n888 = n779 | n783 ;
  assign n889 = n811 & n888 ;
  assign n890 = ( n818 & n888 ) | ( n818 & n889 ) | ( n888 & n889 ) ;
  assign n891 = n811 | n888 ;
  assign n892 = n818 | n891 ;
  assign n893 = ~n890 & n892 ;
  assign n894 = x8 & x11 ;
  assign n895 = n360 | n894 ;
  assign n896 = x3 & x16 ;
  assign n897 = ( n360 & n894 ) | ( n360 & n896 ) | ( n894 & n896 ) ;
  assign n898 = n895 & ~n897 ;
  assign n899 = n360 & n894 ;
  assign n900 = n896 & ~n899 ;
  assign n901 = ~n895 & n896 ;
  assign n902 = ( n896 & ~n900 ) | ( n896 & n901 ) | ( ~n900 & n901 ) ;
  assign n903 = n898 | n902 ;
  assign n904 = n893 & ~n903 ;
  assign n905 = n893 | n903 ;
  assign n906 = ( ~n893 & n904 ) | ( ~n893 & n905 ) | ( n904 & n905 ) ;
  assign n907 = n887 & n906 ;
  assign n908 = n887 | n906 ;
  assign n909 = ~n907 & n908 ;
  assign n910 = x15 & n82 ;
  assign n911 = x17 & n67 ;
  assign n912 = n910 | n911 ;
  assign n913 = x15 & x17 ;
  assign n914 = n119 & n913 ;
  assign n915 = x19 & ~n914 ;
  assign n916 = n912 & n915 ;
  assign n917 = x0 & x19 ;
  assign n918 = ~n916 & n917 ;
  assign n919 = n914 | n916 ;
  assign n920 = x2 & x17 ;
  assign n921 = x4 & x15 ;
  assign n922 = ( ~n914 & n920 ) | ( ~n914 & n921 ) | ( n920 & n921 ) ;
  assign n923 = n920 & n921 ;
  assign n924 = ( ~n916 & n922 ) | ( ~n916 & n923 ) | ( n922 & n923 ) ;
  assign n925 = ~n919 & n924 ;
  assign n926 = n918 | n925 ;
  assign n927 = n135 & n487 ;
  assign n928 = n204 & n650 ;
  assign n929 = n927 | n928 ;
  assign n930 = n200 & n647 ;
  assign n931 = x14 & n930 ;
  assign n932 = ( x14 & ~n929 ) | ( x14 & n931 ) | ( ~n929 & n931 ) ;
  assign n933 = x5 & n932 ;
  assign n934 = n929 | n930 ;
  assign n935 = x6 & x13 ;
  assign n936 = x7 & x12 ;
  assign n937 = ( ~n930 & n935 ) | ( ~n930 & n936 ) | ( n935 & n936 ) ;
  assign n938 = n935 & n936 ;
  assign n939 = ( ~n929 & n937 ) | ( ~n929 & n938 ) | ( n937 & n938 ) ;
  assign n940 = ~n934 & n939 ;
  assign n941 = n933 | n940 ;
  assign n942 = n926 & n941 ;
  assign n943 = n926 & ~n942 ;
  assign n944 = ( n701 & n709 ) | ( n701 & n728 ) | ( n709 & n728 ) ;
  assign n945 = n941 & n944 ;
  assign n946 = ~n926 & n945 ;
  assign n947 = ( n943 & n944 ) | ( n943 & n946 ) | ( n944 & n946 ) ;
  assign n948 = n941 | n944 ;
  assign n949 = ( ~n926 & n944 ) | ( ~n926 & n948 ) | ( n944 & n948 ) ;
  assign n950 = n943 | n949 ;
  assign n951 = ~n947 & n950 ;
  assign n952 = n838 | n844 ;
  assign n953 = ( n844 & n848 ) | ( n844 & n952 ) | ( n848 & n952 ) ;
  assign n954 = n951 & n953 ;
  assign n955 = n951 | n953 ;
  assign n956 = ~n954 & n955 ;
  assign n957 = n909 & n956 ;
  assign n958 = n909 | n956 ;
  assign n959 = ~n957 & n958 ;
  assign n960 = n829 | n851 ;
  assign n961 = ( n829 & n832 ) | ( n829 & n960 ) | ( n832 & n960 ) ;
  assign n962 = ( n871 & n959 ) | ( n871 & ~n961 ) | ( n959 & ~n961 ) ;
  assign n963 = ( ~n959 & n961 ) | ( ~n959 & n962 ) | ( n961 & n962 ) ;
  assign n964 = ( ~n871 & n962 ) | ( ~n871 & n963 ) | ( n962 & n963 ) ;
  assign n965 = n959 & n961 ;
  assign n966 = n959 | n961 ;
  assign n967 = n965 | n966 ;
  assign n968 = ( n871 & n965 ) | ( n871 & n967 ) | ( n965 & n967 ) ;
  assign n969 = x9 & x11 ;
  assign n970 = x1 & x19 ;
  assign n971 = n969 | n970 ;
  assign n972 = n969 & n970 ;
  assign n973 = n971 & ~n972 ;
  assign n974 = n897 & n973 ;
  assign n975 = n897 & ~n973 ;
  assign n976 = ( n973 & ~n974 ) | ( n973 & n975 ) | ( ~n974 & n975 ) ;
  assign n977 = n919 | n976 ;
  assign n978 = ~n976 & n977 ;
  assign n979 = ( ~n919 & n977 ) | ( ~n919 & n978 ) | ( n977 & n978 ) ;
  assign n980 = n942 & n979 ;
  assign n981 = ( n947 & n979 ) | ( n947 & n980 ) | ( n979 & n980 ) ;
  assign n982 = n942 | n979 ;
  assign n983 = n947 | n982 ;
  assign n984 = ~n981 & n983 ;
  assign n985 = x0 & x20 ;
  assign n986 = x7 & x13 ;
  assign n987 = n985 | n986 ;
  assign n988 = n985 & n986 ;
  assign n989 = n987 & ~n988 ;
  assign n990 = n876 & n989 ;
  assign n991 = n876 | n989 ;
  assign n992 = ~n990 & n991 ;
  assign n993 = n934 & n992 ;
  assign n994 = n934 | n992 ;
  assign n995 = ~n993 & n994 ;
  assign n996 = n181 & n487 ;
  assign n997 = x8 & x15 ;
  assign n998 = n706 & n997 ;
  assign n999 = n996 | n998 ;
  assign n1000 = n204 & n792 ;
  assign n1001 = x12 & n1000 ;
  assign n1002 = ( x12 & ~n999 ) | ( x12 & n1001 ) | ( ~n999 & n1001 ) ;
  assign n1003 = x8 & n1002 ;
  assign n1004 = n999 | n1000 ;
  assign n1005 = x5 & x15 ;
  assign n1006 = x6 & x14 ;
  assign n1007 = ( ~n1000 & n1005 ) | ( ~n1000 & n1006 ) | ( n1005 & n1006 ) ;
  assign n1008 = n1005 & n1006 ;
  assign n1009 = ( ~n999 & n1007 ) | ( ~n999 & n1008 ) | ( n1007 & n1008 ) ;
  assign n1010 = ~n1004 & n1009 ;
  assign n1011 = n1003 | n1010 ;
  assign n1012 = ~n995 & n1011 ;
  assign n1013 = n995 & ~n1011 ;
  assign n1014 = n1012 | n1013 ;
  assign n1015 = n984 & n1014 ;
  assign n1016 = n984 | n1014 ;
  assign n1017 = ~n1015 & n1016 ;
  assign n1036 = n799 | n873 ;
  assign n1037 = ( n873 & n879 ) | ( n873 & n1036 ) | ( n879 & n1036 ) ;
  assign n1018 = x16 & x18 ;
  assign n1019 = n119 & n1018 ;
  assign n1020 = x17 & x18 ;
  assign n1021 = n77 & n1020 ;
  assign n1022 = n1019 | n1021 ;
  assign n1023 = x16 & x17 ;
  assign n1024 = n79 & n1023 ;
  assign n1025 = x18 & n1024 ;
  assign n1026 = ( x18 & ~n1022 ) | ( x18 & n1025 ) | ( ~n1022 & n1025 ) ;
  assign n1027 = x2 & n1026 ;
  assign n1028 = n1022 | n1024 ;
  assign n1029 = x3 & x17 ;
  assign n1030 = x4 & x16 ;
  assign n1031 = ( ~n1024 & n1029 ) | ( ~n1024 & n1030 ) | ( n1029 & n1030 ) ;
  assign n1032 = n1029 & n1030 ;
  assign n1033 = ( ~n1022 & n1031 ) | ( ~n1022 & n1032 ) | ( n1031 & n1032 ) ;
  assign n1034 = ~n1028 & n1033 ;
  assign n1035 = n1027 | n1034 ;
  assign n1038 = n1035 & n1037 ;
  assign n1039 = n1037 & ~n1038 ;
  assign n1040 = n1035 & ~n1038 ;
  assign n1041 = n1039 | n1040 ;
  assign n1042 = n890 | n903 ;
  assign n1043 = ( n890 & n893 ) | ( n890 & n1042 ) | ( n893 & n1042 ) ;
  assign n1044 = n1041 | n1043 ;
  assign n1045 = n1041 & n1043 ;
  assign n1046 = n1044 & ~n1045 ;
  assign n1047 = n884 | n906 ;
  assign n1048 = ( n884 & n887 ) | ( n884 & n1047 ) | ( n887 & n1047 ) ;
  assign n1049 = n1046 | n1048 ;
  assign n1050 = n1046 & n1048 ;
  assign n1051 = n1049 & ~n1050 ;
  assign n1052 = n1017 & n1051 ;
  assign n1053 = n1051 & ~n1052 ;
  assign n1054 = ( n1017 & ~n1052 ) | ( n1017 & n1053 ) | ( ~n1052 & n1053 ) ;
  assign n1055 = n909 | n954 ;
  assign n1056 = ( n954 & n956 ) | ( n954 & n1055 ) | ( n956 & n1055 ) ;
  assign n1057 = ( n968 & n1054 ) | ( n968 & ~n1056 ) | ( n1054 & ~n1056 ) ;
  assign n1058 = ( ~n1054 & n1056 ) | ( ~n1054 & n1057 ) | ( n1056 & n1057 ) ;
  assign n1059 = ( ~n968 & n1057 ) | ( ~n968 & n1058 ) | ( n1057 & n1058 ) ;
  assign n1163 = n1052 & ~n1056 ;
  assign n1164 = n1017 | n1056 ;
  assign n1165 = ( n1053 & ~n1163 ) | ( n1053 & n1164 ) | ( ~n1163 & n1164 ) ;
  assign n1166 = n965 & n1165 ;
  assign n1167 = ~n1052 & n1056 ;
  assign n1168 = n1017 & n1056 ;
  assign n1169 = ( n1053 & n1167 ) | ( n1053 & n1168 ) | ( n1167 & n1168 ) ;
  assign n1170 = n1166 | n1169 ;
  assign n1171 = n1165 | n1169 ;
  assign n1172 = ( n967 & n1169 ) | ( n967 & n1171 ) | ( n1169 & n1171 ) ;
  assign n1173 = ( n871 & n1170 ) | ( n871 & n1172 ) | ( n1170 & n1172 ) ;
  assign n1060 = n1050 | n1052 ;
  assign n1061 = n1004 | n1028 ;
  assign n1062 = n1004 & n1028 ;
  assign n1063 = n1061 & ~n1062 ;
  assign n1064 = n876 | n988 ;
  assign n1065 = ( n988 & n989 ) | ( n988 & n1064 ) | ( n989 & n1064 ) ;
  assign n1066 = n1063 | n1065 ;
  assign n1067 = n1063 & n1065 ;
  assign n1068 = n1066 & ~n1067 ;
  assign n1069 = n1038 | n1043 ;
  assign n1070 = ( n1038 & n1041 ) | ( n1038 & n1069 ) | ( n1041 & n1069 ) ;
  assign n1071 = n1068 | n1070 ;
  assign n1072 = n1068 & n1070 ;
  assign n1073 = n1071 & ~n1072 ;
  assign n1074 = x19 & n801 ;
  assign n1075 = x3 & n1018 ;
  assign n1076 = n1074 | n1075 ;
  assign n1077 = x18 & x19 ;
  assign n1078 = n77 & n1077 ;
  assign n1079 = x5 & ~n1078 ;
  assign n1080 = n1076 & n1079 ;
  assign n1081 = x5 & x16 ;
  assign n1082 = ~n1080 & n1081 ;
  assign n1083 = n1078 | n1080 ;
  assign n1084 = x2 & x19 ;
  assign n1085 = x3 & x18 ;
  assign n1086 = ( ~n1078 & n1084 ) | ( ~n1078 & n1085 ) | ( n1084 & n1085 ) ;
  assign n1087 = n1084 & n1085 ;
  assign n1088 = ( ~n1080 & n1086 ) | ( ~n1080 & n1087 ) | ( n1086 & n1087 ) ;
  assign n1089 = ~n1083 & n1088 ;
  assign n1090 = n1082 | n1089 ;
  assign n1091 = n181 & n723 ;
  assign n1092 = n200 & n792 ;
  assign n1093 = n1091 | n1092 ;
  assign n1094 = n251 & n650 ;
  assign n1095 = x15 & n1094 ;
  assign n1096 = ( x15 & ~n1093 ) | ( x15 & n1095 ) | ( ~n1093 & n1095 ) ;
  assign n1097 = x6 & n1096 ;
  assign n1098 = n1093 | n1094 ;
  assign n1099 = x7 & x14 ;
  assign n1100 = x8 & x13 ;
  assign n1101 = ( ~n1094 & n1099 ) | ( ~n1094 & n1100 ) | ( n1099 & n1100 ) ;
  assign n1102 = n1099 & n1100 ;
  assign n1103 = ( ~n1093 & n1101 ) | ( ~n1093 & n1102 ) | ( n1101 & n1102 ) ;
  assign n1104 = ~n1098 & n1103 ;
  assign n1105 = n1097 | n1104 ;
  assign n1106 = n1090 & n1105 ;
  assign n1107 = n1090 & ~n1106 ;
  assign n1108 = x9 & x12 ;
  assign n1109 = n618 | n1108 ;
  assign n1110 = n360 & n490 ;
  assign n1111 = x4 & x17 ;
  assign n1112 = ~n1110 & n1111 ;
  assign n1113 = n1109 | n1110 ;
  assign n1114 = ( n1110 & n1112 ) | ( n1110 & n1113 ) | ( n1112 & n1113 ) ;
  assign n1115 = n1109 & ~n1114 ;
  assign n1116 = ~n1109 & n1111 ;
  assign n1117 = ( n1111 & ~n1112 ) | ( n1111 & n1116 ) | ( ~n1112 & n1116 ) ;
  assign n1118 = n1115 | n1117 ;
  assign n1119 = ~n1105 & n1118 ;
  assign n1120 = ( n1090 & n1118 ) | ( n1090 & n1119 ) | ( n1118 & n1119 ) ;
  assign n1121 = ~n1107 & n1120 ;
  assign n1122 = n1105 & ~n1118 ;
  assign n1123 = ~n1090 & n1122 ;
  assign n1124 = ( n1107 & ~n1118 ) | ( n1107 & n1123 ) | ( ~n1118 & n1123 ) ;
  assign n1125 = n1121 | n1124 ;
  assign n1126 = n1073 | n1125 ;
  assign n1127 = n1073 & n1125 ;
  assign n1128 = n1126 & ~n1127 ;
  assign n1129 = x0 & x21 ;
  assign n1130 = n972 & ~n1129 ;
  assign n1131 = ~n972 & n1129 ;
  assign n1132 = n1130 | n1131 ;
  assign n1133 = x1 & x20 ;
  assign n1134 = x11 & n1133 ;
  assign n1135 = x11 & ~n1133 ;
  assign n1136 = ( n1133 & ~n1134 ) | ( n1133 & n1135 ) | ( ~n1134 & n1135 ) ;
  assign n1137 = n1132 & n1136 ;
  assign n1138 = n1132 | n1136 ;
  assign n1139 = ~n1137 & n1138 ;
  assign n1140 = n919 | n974 ;
  assign n1141 = ( n974 & n976 ) | ( n974 & n1140 ) | ( n976 & n1140 ) ;
  assign n1142 = n1139 & n1141 ;
  assign n1143 = n1139 | n1141 ;
  assign n1144 = ~n1142 & n1143 ;
  assign n1145 = n993 | n1011 ;
  assign n1146 = ( n993 & n995 ) | ( n993 & n1145 ) | ( n995 & n1145 ) ;
  assign n1147 = n1144 | n1146 ;
  assign n1148 = n1144 & n1146 ;
  assign n1149 = n1147 & ~n1148 ;
  assign n1150 = n980 | n1014 ;
  assign n1151 = n979 | n1014 ;
  assign n1152 = ( n947 & n1150 ) | ( n947 & n1151 ) | ( n1150 & n1151 ) ;
  assign n1153 = n1149 & n1152 ;
  assign n1154 = n981 & n1149 ;
  assign n1155 = ( n984 & n1153 ) | ( n984 & n1154 ) | ( n1153 & n1154 ) ;
  assign n1156 = n1149 | n1152 ;
  assign n1157 = n981 | n1149 ;
  assign n1158 = ( n984 & n1156 ) | ( n984 & n1157 ) | ( n1156 & n1157 ) ;
  assign n1159 = ~n1155 & n1158 ;
  assign n1160 = n1128 & n1159 ;
  assign n1161 = n1128 | n1159 ;
  assign n1162 = ~n1160 & n1161 ;
  assign n1174 = ( n1060 & ~n1162 ) | ( n1060 & n1173 ) | ( ~n1162 & n1173 ) ;
  assign n1175 = ( ~n1060 & n1162 ) | ( ~n1060 & n1174 ) | ( n1162 & n1174 ) ;
  assign n1176 = ( ~n1173 & n1174 ) | ( ~n1173 & n1175 ) | ( n1174 & n1175 ) ;
  assign n1177 = n1083 | n1098 ;
  assign n1178 = n1083 & n1098 ;
  assign n1179 = n1177 & ~n1178 ;
  assign n1180 = ( n972 & n1129 ) | ( n972 & n1136 ) | ( n1129 & n1136 ) ;
  assign n1181 = n1179 | n1180 ;
  assign n1182 = n1179 & n1180 ;
  assign n1183 = n1181 & ~n1182 ;
  assign n1184 = n1142 | n1146 ;
  assign n1185 = ( n1142 & n1144 ) | ( n1142 & n1184 ) | ( n1144 & n1184 ) ;
  assign n1186 = n1183 | n1185 ;
  assign n1187 = n1183 & n1185 ;
  assign n1188 = n1186 & ~n1187 ;
  assign n1189 = x7 & x15 ;
  assign n1190 = x8 & x14 ;
  assign n1191 = n1189 | n1190 ;
  assign n1192 = n251 & n792 ;
  assign n1193 = n1191 | n1192 ;
  assign n1194 = x0 & x22 ;
  assign n1195 = ( ~n1192 & n1193 ) | ( ~n1192 & n1194 ) | ( n1193 & n1194 ) ;
  assign n1196 = ( n1192 & n1193 ) | ( n1192 & ~n1194 ) | ( n1193 & ~n1194 ) ;
  assign n1197 = ( ~n1193 & n1195 ) | ( ~n1193 & n1196 ) | ( n1195 & n1196 ) ;
  assign n1198 = x2 & x20 ;
  assign n1199 = n623 | n1198 ;
  assign n1200 = ( n415 & n623 ) | ( n415 & n1198 ) | ( n623 & n1198 ) ;
  assign n1201 = n1199 & ~n1200 ;
  assign n1202 = n623 & n1198 ;
  assign n1203 = n415 & ~n1202 ;
  assign n1204 = n415 & ~n1199 ;
  assign n1205 = ( n415 & ~n1203 ) | ( n415 & n1204 ) | ( ~n1203 & n1204 ) ;
  assign n1206 = n1201 | n1205 ;
  assign n1207 = n1197 & n1206 ;
  assign n1208 = n1197 & ~n1207 ;
  assign n1209 = n1206 & ~n1207 ;
  assign n1210 = n1208 | n1209 ;
  assign n1211 = x3 & x19 ;
  assign n1212 = n79 & n1077 ;
  assign n1213 = x5 & x17 ;
  assign n1214 = n1211 & n1213 ;
  assign n1215 = n1212 | n1214 ;
  assign n1216 = n91 & n1020 ;
  assign n1217 = n1211 & n1216 ;
  assign n1218 = ( n1211 & ~n1215 ) | ( n1211 & n1217 ) | ( ~n1215 & n1217 ) ;
  assign n1219 = n1215 | n1216 ;
  assign n1220 = x4 & x18 ;
  assign n1221 = ( n1213 & ~n1216 ) | ( n1213 & n1220 ) | ( ~n1216 & n1220 ) ;
  assign n1222 = n1213 & n1220 ;
  assign n1223 = ( ~n1215 & n1221 ) | ( ~n1215 & n1222 ) | ( n1221 & n1222 ) ;
  assign n1224 = ~n1219 & n1223 ;
  assign n1225 = n1218 | n1224 ;
  assign n1226 = ~n1210 & n1225 ;
  assign n1227 = n1210 & ~n1225 ;
  assign n1228 = n1226 | n1227 ;
  assign n1229 = n1188 | n1228 ;
  assign n1230 = n1188 & n1228 ;
  assign n1231 = n1229 & ~n1230 ;
  assign n1256 = n1072 | n1125 ;
  assign n1257 = ( n1072 & n1073 ) | ( n1072 & n1256 ) | ( n1073 & n1256 ) ;
  assign n1242 = n1062 | n1065 ;
  assign n1243 = ( n1062 & n1063 ) | ( n1062 & n1242 ) | ( n1063 & n1242 ) ;
  assign n1232 = x1 & x21 ;
  assign n1233 = n363 & n1232 ;
  assign n1234 = n363 | n1232 ;
  assign n1235 = ~n1233 & n1234 ;
  assign n1236 = n1134 & n1235 ;
  assign n1237 = n1134 | n1235 ;
  assign n1238 = ~n1236 & n1237 ;
  assign n1239 = n1114 & n1238 ;
  assign n1240 = n1114 | n1238 ;
  assign n1241 = ~n1239 & n1240 ;
  assign n1244 = n1241 & n1243 ;
  assign n1245 = n1243 & ~n1244 ;
  assign n1246 = n1241 & ~n1244 ;
  assign n1247 = n1245 | n1246 ;
  assign n1248 = n1105 & n1118 ;
  assign n1249 = ~n1090 & n1248 ;
  assign n1250 = n1106 | n1249 ;
  assign n1251 = n1106 | n1118 ;
  assign n1252 = ( n1107 & n1250 ) | ( n1107 & n1251 ) | ( n1250 & n1251 ) ;
  assign n1253 = n1247 & n1252 ;
  assign n1254 = n1247 | n1252 ;
  assign n1255 = ~n1253 & n1254 ;
  assign n1258 = n1255 & n1257 ;
  assign n1259 = n1257 & ~n1258 ;
  assign n1260 = n1255 & ~n1257 ;
  assign n1261 = n1231 & n1260 ;
  assign n1262 = ( n1231 & n1259 ) | ( n1231 & n1261 ) | ( n1259 & n1261 ) ;
  assign n1263 = n1231 | n1260 ;
  assign n1264 = n1259 | n1263 ;
  assign n1265 = ~n1262 & n1264 ;
  assign n1266 = n1128 | n1155 ;
  assign n1267 = ( n1155 & n1159 ) | ( n1155 & n1266 ) | ( n1159 & n1266 ) ;
  assign n1268 = n1265 & n1267 ;
  assign n1269 = n1265 | n1267 ;
  assign n1270 = ~n1268 & n1269 ;
  assign n1271 = n1060 & n1162 ;
  assign n1272 = n1060 | n1162 ;
  assign n1273 = n1271 | n1272 ;
  assign n1274 = ( n1173 & n1271 ) | ( n1173 & n1273 ) | ( n1271 & n1273 ) ;
  assign n1275 = n1270 | n1274 ;
  assign n1276 = n1269 & n1273 ;
  assign n1277 = n1269 & n1271 ;
  assign n1278 = ( n1173 & n1276 ) | ( n1173 & n1277 ) | ( n1276 & n1277 ) ;
  assign n1279 = ~n1268 & n1278 ;
  assign n1280 = n1275 & ~n1279 ;
  assign n1383 = n1268 | n1277 ;
  assign n1384 = n1268 | n1276 ;
  assign n1385 = ( n1173 & n1383 ) | ( n1173 & n1384 ) | ( n1383 & n1384 ) ;
  assign n1281 = x17 & x20 ;
  assign n1282 = n209 & n1281 ;
  assign n1283 = n204 & n1020 ;
  assign n1284 = n1282 | n1283 ;
  assign n1285 = x18 & x20 ;
  assign n1286 = n169 & n1285 ;
  assign n1287 = x17 & n1286 ;
  assign n1288 = ( x17 & ~n1284 ) | ( x17 & n1287 ) | ( ~n1284 & n1287 ) ;
  assign n1289 = x6 & n1288 ;
  assign n1290 = n1284 | n1286 ;
  assign n1291 = x3 & x20 ;
  assign n1292 = x5 & x18 ;
  assign n1293 = ( ~n1286 & n1291 ) | ( ~n1286 & n1292 ) | ( n1291 & n1292 ) ;
  assign n1294 = n1291 & n1292 ;
  assign n1295 = ( ~n1284 & n1293 ) | ( ~n1284 & n1294 ) | ( n1293 & n1294 ) ;
  assign n1296 = ~n1290 & n1295 ;
  assign n1297 = n1289 | n1296 ;
  assign n1298 = x10 & x13 ;
  assign n1299 = n490 | n1298 ;
  assign n1300 = n618 & n647 ;
  assign n1301 = x4 & x19 ;
  assign n1302 = ~n1300 & n1301 ;
  assign n1303 = n1299 | n1300 ;
  assign n1304 = ( n1300 & n1302 ) | ( n1300 & n1303 ) | ( n1302 & n1303 ) ;
  assign n1305 = n1299 & ~n1304 ;
  assign n1306 = ~n1299 & n1301 ;
  assign n1307 = ( n1301 & ~n1302 ) | ( n1301 & n1306 ) | ( ~n1302 & n1306 ) ;
  assign n1308 = n1305 | n1307 ;
  assign n1309 = n1297 & n1308 ;
  assign n1310 = n1297 & ~n1309 ;
  assign n1311 = n1308 & ~n1309 ;
  assign n1312 = n1310 | n1311 ;
  assign n1313 = n1114 | n1236 ;
  assign n1314 = ( n1236 & n1238 ) | ( n1236 & n1313 ) | ( n1238 & n1313 ) ;
  assign n1315 = n1312 | n1314 ;
  assign n1316 = n1312 & n1314 ;
  assign n1317 = n1315 & ~n1316 ;
  assign n1318 = n667 & n790 ;
  assign n1319 = n251 & n795 ;
  assign n1320 = n1318 | n1319 ;
  assign n1321 = n313 & n792 ;
  assign n1322 = x16 & n1321 ;
  assign n1323 = ( x16 & ~n1320 ) | ( x16 & n1322 ) | ( ~n1320 & n1322 ) ;
  assign n1324 = x7 & n1323 ;
  assign n1325 = n1320 | n1321 ;
  assign n1326 = x9 & x14 ;
  assign n1327 = ( n997 & ~n1321 ) | ( n997 & n1326 ) | ( ~n1321 & n1326 ) ;
  assign n1328 = n997 & n1326 ;
  assign n1329 = ( ~n1320 & n1327 ) | ( ~n1320 & n1328 ) | ( n1327 & n1328 ) ;
  assign n1330 = ~n1325 & n1329 ;
  assign n1331 = n1324 | n1330 ;
  assign n1332 = ~n1192 & n1194 ;
  assign n1333 = ( n1192 & n1193 ) | ( n1192 & n1332 ) | ( n1193 & n1332 ) ;
  assign n1334 = x0 & x23 ;
  assign n1335 = x2 & x21 ;
  assign n1336 = n1334 | n1335 ;
  assign n1337 = x21 & x23 ;
  assign n1338 = n67 & n1337 ;
  assign n1339 = n1336 & ~n1338 ;
  assign n1340 = ( ~n1233 & n1333 ) | ( ~n1233 & n1339 ) | ( n1333 & n1339 ) ;
  assign n1341 = ( n1233 & n1333 ) | ( n1233 & ~n1339 ) | ( n1333 & ~n1339 ) ;
  assign n1342 = ( ~n1333 & n1340 ) | ( ~n1333 & n1341 ) | ( n1340 & n1341 ) ;
  assign n1343 = n1331 & n1342 ;
  assign n1344 = n1331 | n1342 ;
  assign n1345 = ~n1343 & n1344 ;
  assign n1346 = n1317 | n1345 ;
  assign n1347 = n1317 & n1345 ;
  assign n1348 = n1346 & ~n1347 ;
  assign n1349 = n1244 | n1247 ;
  assign n1350 = ( n1244 & n1252 ) | ( n1244 & n1349 ) | ( n1252 & n1349 ) ;
  assign n1351 = n1348 & n1350 ;
  assign n1352 = n1348 | n1350 ;
  assign n1353 = ~n1351 & n1352 ;
  assign n1354 = n1207 | n1225 ;
  assign n1355 = ( n1207 & n1210 ) | ( n1207 & n1354 ) | ( n1210 & n1354 ) ;
  assign n1356 = n1098 | n1180 ;
  assign n1357 = ( n1083 & n1180 ) | ( n1083 & n1356 ) | ( n1180 & n1356 ) ;
  assign n1358 = ( n1178 & n1179 ) | ( n1178 & n1357 ) | ( n1179 & n1357 ) ;
  assign n1359 = n1355 & n1358 ;
  assign n1360 = n1355 | n1358 ;
  assign n1361 = ~n1359 & n1360 ;
  assign n1362 = x1 & x22 ;
  assign n1363 = x12 & n1362 ;
  assign n1364 = x12 | n1362 ;
  assign n1365 = ~n1363 & n1364 ;
  assign n1366 = n1219 | n1365 ;
  assign n1367 = n1219 & n1365 ;
  assign n1368 = n1366 & ~n1367 ;
  assign n1369 = n1200 | n1368 ;
  assign n1370 = n1200 & n1368 ;
  assign n1371 = n1369 & ~n1370 ;
  assign n1372 = n1361 & n1371 ;
  assign n1373 = n1361 | n1371 ;
  assign n1374 = ~n1372 & n1373 ;
  assign n1375 = n1187 | n1228 ;
  assign n1376 = ( n1187 & n1188 ) | ( n1187 & n1375 ) | ( n1188 & n1375 ) ;
  assign n1377 = n1374 & n1376 ;
  assign n1378 = n1374 | n1376 ;
  assign n1379 = ~n1377 & n1378 ;
  assign n1380 = n1353 & n1379 ;
  assign n1381 = n1353 | n1379 ;
  assign n1382 = ~n1380 & n1381 ;
  assign n1386 = n1259 | n1260 ;
  assign n1387 = n1231 | n1258 ;
  assign n1388 = ( n1258 & n1386 ) | ( n1258 & n1387 ) | ( n1386 & n1387 ) ;
  assign n1389 = ( n1382 & n1385 ) | ( n1382 & ~n1388 ) | ( n1385 & ~n1388 ) ;
  assign n1390 = ( ~n1382 & n1388 ) | ( ~n1382 & n1389 ) | ( n1388 & n1389 ) ;
  assign n1391 = ( ~n1385 & n1389 ) | ( ~n1385 & n1390 ) | ( n1389 & n1390 ) ;
  assign n1392 = x0 & x24 ;
  assign n1393 = n1363 & n1392 ;
  assign n1394 = n1363 & ~n1393 ;
  assign n1395 = ~n1363 & n1392 ;
  assign n1396 = n1394 | n1395 ;
  assign n1397 = x1 & x23 ;
  assign n1398 = n720 & n1397 ;
  assign n1399 = n1397 & ~n1398 ;
  assign n1400 = n720 & ~n1398 ;
  assign n1401 = n1399 | n1400 ;
  assign n1402 = ~n1396 & n1401 ;
  assign n1403 = n1396 & ~n1401 ;
  assign n1404 = n1402 | n1403 ;
  assign n1405 = x7 & x17 ;
  assign n1406 = n200 & n1020 ;
  assign n1407 = x2 & x22 ;
  assign n1408 = n1405 & n1407 ;
  assign n1409 = n1406 | n1408 ;
  assign n1410 = x18 & x22 ;
  assign n1411 = n179 & n1410 ;
  assign n1412 = n1405 & n1411 ;
  assign n1413 = ( n1405 & ~n1409 ) | ( n1405 & n1412 ) | ( ~n1409 & n1412 ) ;
  assign n1414 = n1409 | n1411 ;
  assign n1415 = x6 & x18 ;
  assign n1416 = ( n1407 & ~n1411 ) | ( n1407 & n1415 ) | ( ~n1411 & n1415 ) ;
  assign n1417 = n1407 & n1415 ;
  assign n1418 = ( ~n1409 & n1416 ) | ( ~n1409 & n1417 ) | ( n1416 & n1417 ) ;
  assign n1419 = ~n1414 & n1418 ;
  assign n1420 = n1413 | n1419 ;
  assign n1421 = n1404 & n1420 ;
  assign n1422 = n1404 | n1420 ;
  assign n1423 = ~n1421 & n1422 ;
  assign n1424 = n1200 | n1365 ;
  assign n1425 = ( n1200 & n1219 ) | ( n1200 & n1424 ) | ( n1219 & n1424 ) ;
  assign n1426 = ( n1367 & n1368 ) | ( n1367 & n1425 ) | ( n1368 & n1425 ) ;
  assign n1427 = n1423 | n1426 ;
  assign n1428 = n1423 & n1426 ;
  assign n1429 = n1427 & ~n1428 ;
  assign n1430 = n1233 | n1338 ;
  assign n1431 = ( n1338 & n1339 ) | ( n1338 & n1430 ) | ( n1339 & n1430 ) ;
  assign n1432 = x19 & x21 ;
  assign n1433 = n169 & n1432 ;
  assign n1434 = x20 & x21 ;
  assign n1435 = n79 & n1434 ;
  assign n1436 = n1433 | n1435 ;
  assign n1437 = x19 & x20 ;
  assign n1438 = n91 & n1437 ;
  assign n1439 = x3 & n1438 ;
  assign n1440 = ( x3 & ~n1436 ) | ( x3 & n1439 ) | ( ~n1436 & n1439 ) ;
  assign n1441 = x21 & n1440 ;
  assign n1442 = n1436 | n1438 ;
  assign n1443 = x4 & x20 ;
  assign n1444 = x5 & x19 ;
  assign n1445 = ( ~n1438 & n1443 ) | ( ~n1438 & n1444 ) | ( n1443 & n1444 ) ;
  assign n1446 = n1443 & n1444 ;
  assign n1447 = ( ~n1436 & n1445 ) | ( ~n1436 & n1446 ) | ( n1445 & n1446 ) ;
  assign n1448 = ~n1442 & n1447 ;
  assign n1449 = ~n1431 & n1448 ;
  assign n1450 = ( ~n1431 & n1441 ) | ( ~n1431 & n1449 ) | ( n1441 & n1449 ) ;
  assign n1451 = n1431 & ~n1448 ;
  assign n1452 = ~n1441 & n1451 ;
  assign n1453 = n1450 | n1452 ;
  assign n1454 = x8 & x16 ;
  assign n1455 = n249 & n790 ;
  assign n1456 = n313 & n795 ;
  assign n1457 = n1455 | n1456 ;
  assign n1458 = n360 & n792 ;
  assign n1459 = n1454 & n1458 ;
  assign n1460 = ( n1454 & ~n1457 ) | ( n1454 & n1459 ) | ( ~n1457 & n1459 ) ;
  assign n1461 = n1457 | n1458 ;
  assign n1462 = x9 & x15 ;
  assign n1463 = x10 & x14 ;
  assign n1464 = ( ~n1458 & n1462 ) | ( ~n1458 & n1463 ) | ( n1462 & n1463 ) ;
  assign n1465 = n1462 & n1463 ;
  assign n1466 = ( ~n1457 & n1464 ) | ( ~n1457 & n1465 ) | ( n1464 & n1465 ) ;
  assign n1467 = ~n1461 & n1466 ;
  assign n1468 = n1460 | n1467 ;
  assign n1469 = n1453 & n1468 ;
  assign n1470 = n1453 | n1468 ;
  assign n1471 = ~n1469 & n1470 ;
  assign n1472 = n1429 | n1471 ;
  assign n1473 = n1429 & n1471 ;
  assign n1474 = n1472 & ~n1473 ;
  assign n1475 = n1358 | n1371 ;
  assign n1476 = ( n1355 & n1371 ) | ( n1355 & n1475 ) | ( n1371 & n1475 ) ;
  assign n1477 = ( n1359 & n1361 ) | ( n1359 & n1476 ) | ( n1361 & n1476 ) ;
  assign n1478 = n1474 & n1477 ;
  assign n1479 = n1474 | n1477 ;
  assign n1480 = ~n1478 & n1479 ;
  assign n1503 = n1347 | n1350 ;
  assign n1504 = ( n1347 & n1348 ) | ( n1347 & n1503 ) | ( n1348 & n1503 ) ;
  assign n1481 = n1290 | n1304 ;
  assign n1482 = n1290 & n1304 ;
  assign n1483 = n1481 & ~n1482 ;
  assign n1484 = n1325 | n1483 ;
  assign n1485 = n1325 & n1483 ;
  assign n1486 = n1484 & ~n1485 ;
  assign n1487 = n1336 & ~n1431 ;
  assign n1488 = n1233 & ~n1339 ;
  assign n1489 = n1333 & n1488 ;
  assign n1490 = ( n1333 & n1487 ) | ( n1333 & n1489 ) | ( n1487 & n1489 ) ;
  assign n1491 = n1343 | n1490 ;
  assign n1492 = n1309 | n1314 ;
  assign n1493 = n1491 & n1492 ;
  assign n1494 = n1309 & n1491 ;
  assign n1495 = ( n1312 & n1493 ) | ( n1312 & n1494 ) | ( n1493 & n1494 ) ;
  assign n1496 = n1491 | n1492 ;
  assign n1497 = n1309 | n1491 ;
  assign n1498 = ( n1312 & n1496 ) | ( n1312 & n1497 ) | ( n1496 & n1497 ) ;
  assign n1499 = ~n1495 & n1498 ;
  assign n1500 = n1486 & n1499 ;
  assign n1501 = n1486 | n1499 ;
  assign n1502 = ~n1500 & n1501 ;
  assign n1505 = n1502 & n1504 ;
  assign n1506 = n1504 & ~n1505 ;
  assign n1507 = n1502 & ~n1504 ;
  assign n1508 = n1480 | n1507 ;
  assign n1509 = n1506 | n1508 ;
  assign n1510 = ~n1480 & n1509 ;
  assign n1511 = n1377 | n1380 ;
  assign n1512 = n1509 & n1511 ;
  assign n1513 = n1506 | n1507 ;
  assign n1514 = n1511 & ~n1513 ;
  assign n1515 = ( n1510 & n1512 ) | ( n1510 & n1514 ) | ( n1512 & n1514 ) ;
  assign n1516 = n1509 | n1511 ;
  assign n1517 = ~n1511 & n1513 ;
  assign n1518 = ( n1510 & n1516 ) | ( n1510 & ~n1517 ) | ( n1516 & ~n1517 ) ;
  assign n1519 = ~n1515 & n1518 ;
  assign n1520 = n1382 & n1388 ;
  assign n1521 = n1382 | n1388 ;
  assign n1522 = n1520 | n1521 ;
  assign n1523 = ( n1385 & n1520 ) | ( n1385 & n1522 ) | ( n1520 & n1522 ) ;
  assign n1524 = n1519 | n1523 ;
  assign n1525 = n1518 & n1522 ;
  assign n1526 = n1518 & n1520 ;
  assign n1527 = ( n1385 & n1525 ) | ( n1385 & n1526 ) | ( n1525 & n1526 ) ;
  assign n1528 = ~n1515 & n1527 ;
  assign n1529 = n1524 & ~n1528 ;
  assign n1651 = n1515 | n1526 ;
  assign n1652 = n1515 | n1525 ;
  assign n1653 = ( n1385 & n1651 ) | ( n1385 & n1652 ) | ( n1651 & n1652 ) ;
  assign n1548 = n1473 | n1477 ;
  assign n1549 = ( n1473 & n1474 ) | ( n1473 & n1548 ) | ( n1474 & n1548 ) ;
  assign n1530 = n1414 | n1461 ;
  assign n1531 = n1414 & n1461 ;
  assign n1532 = n1530 & ~n1531 ;
  assign n1533 = n1393 | n1401 ;
  assign n1534 = ( n1393 & n1396 ) | ( n1393 & n1533 ) | ( n1396 & n1533 ) ;
  assign n1535 = n1532 | n1534 ;
  assign n1536 = n1532 & n1534 ;
  assign n1537 = n1535 & ~n1536 ;
  assign n1538 = n1441 | n1448 ;
  assign n1539 = ( n1431 & n1468 ) | ( n1431 & n1538 ) | ( n1468 & n1538 ) ;
  assign n1540 = n1537 | n1539 ;
  assign n1541 = n1537 & n1539 ;
  assign n1542 = n1540 & ~n1541 ;
  assign n1543 = n1421 | n1426 ;
  assign n1544 = ( n1421 & n1423 ) | ( n1421 & n1543 ) | ( n1423 & n1543 ) ;
  assign n1545 = n1542 | n1544 ;
  assign n1546 = n1542 & n1544 ;
  assign n1547 = n1545 & ~n1546 ;
  assign n1550 = n1547 & n1549 ;
  assign n1551 = n1549 & ~n1550 ;
  assign n1552 = n1547 & ~n1549 ;
  assign n1553 = n1551 | n1552 ;
  assign n1604 = n1486 | n1495 ;
  assign n1605 = ( n1495 & n1499 ) | ( n1495 & n1604 ) | ( n1499 & n1604 ) ;
  assign n1554 = x0 & x25 ;
  assign n1555 = x2 & x23 ;
  assign n1556 = n1554 | n1555 ;
  assign n1557 = x23 & x25 ;
  assign n1558 = n67 & n1557 ;
  assign n1559 = n582 & ~n1558 ;
  assign n1560 = n1556 | n1558 ;
  assign n1561 = ( n1558 & n1559 ) | ( n1558 & n1560 ) | ( n1559 & n1560 ) ;
  assign n1562 = n1556 & ~n1561 ;
  assign n1563 = n582 & ~n1556 ;
  assign n1564 = ( n582 & ~n1559 ) | ( n582 & n1563 ) | ( ~n1559 & n1563 ) ;
  assign n1565 = n1562 | n1564 ;
  assign n1566 = n667 & n1018 ;
  assign n1567 = n251 & n1020 ;
  assign n1568 = n1566 | n1567 ;
  assign n1569 = n313 & n1023 ;
  assign n1570 = n780 & n1569 ;
  assign n1571 = ( n780 & ~n1568 ) | ( n780 & n1570 ) | ( ~n1568 & n1570 ) ;
  assign n1572 = n1568 | n1569 ;
  assign n1573 = x8 & x17 ;
  assign n1574 = ( n754 & ~n1569 ) | ( n754 & n1573 ) | ( ~n1569 & n1573 ) ;
  assign n1575 = n754 & n1573 ;
  assign n1576 = ( ~n1568 & n1574 ) | ( ~n1568 & n1575 ) | ( n1574 & n1575 ) ;
  assign n1577 = ~n1572 & n1576 ;
  assign n1578 = n1571 | n1577 ;
  assign n1579 = n1565 & n1578 ;
  assign n1580 = n1565 & ~n1579 ;
  assign n1581 = x6 & x19 ;
  assign n1582 = x22 & n1211 ;
  assign n1583 = x4 & n1432 ;
  assign n1584 = n1582 | n1583 ;
  assign n1585 = x21 & x22 ;
  assign n1586 = n79 & n1585 ;
  assign n1587 = x6 & ~n1586 ;
  assign n1588 = n1584 & n1587 ;
  assign n1589 = n1581 & ~n1588 ;
  assign n1590 = n1586 | n1588 ;
  assign n1591 = x3 & x22 ;
  assign n1592 = x4 & x21 ;
  assign n1593 = ( ~n1586 & n1591 ) | ( ~n1586 & n1592 ) | ( n1591 & n1592 ) ;
  assign n1594 = n1591 & n1592 ;
  assign n1595 = ( ~n1588 & n1593 ) | ( ~n1588 & n1594 ) | ( n1593 & n1594 ) ;
  assign n1596 = ~n1590 & n1595 ;
  assign n1597 = n1589 | n1596 ;
  assign n1598 = ~n1565 & n1578 ;
  assign n1599 = n1597 & n1598 ;
  assign n1600 = ( n1580 & n1597 ) | ( n1580 & n1599 ) | ( n1597 & n1599 ) ;
  assign n1601 = n1597 | n1598 ;
  assign n1602 = n1580 | n1601 ;
  assign n1603 = ~n1600 & n1602 ;
  assign n1606 = n1603 & n1605 ;
  assign n1607 = n1605 & ~n1606 ;
  assign n1608 = x1 & x24 ;
  assign n1609 = x13 & n1608 ;
  assign n1610 = x13 | n1608 ;
  assign n1611 = ~n1609 & n1610 ;
  assign n1612 = n1398 & n1611 ;
  assign n1613 = n1398 | n1611 ;
  assign n1614 = ~n1612 & n1613 ;
  assign n1615 = n1442 & n1614 ;
  assign n1616 = n1442 | n1614 ;
  assign n1617 = ~n1615 & n1616 ;
  assign n1628 = n1325 | n1482 ;
  assign n1629 = ( n1482 & n1483 ) | ( n1482 & n1628 ) | ( n1483 & n1628 ) ;
  assign n1618 = x11 & x14 ;
  assign n1619 = n647 | n1618 ;
  assign n1620 = x5 & x20 ;
  assign n1621 = ( n647 & n1618 ) | ( n647 & n1620 ) | ( n1618 & n1620 ) ;
  assign n1622 = n1619 & ~n1621 ;
  assign n1623 = n647 & n1618 ;
  assign n1624 = n1620 & ~n1623 ;
  assign n1625 = ~n1619 & n1620 ;
  assign n1626 = ( n1620 & ~n1624 ) | ( n1620 & n1625 ) | ( ~n1624 & n1625 ) ;
  assign n1627 = n1622 | n1626 ;
  assign n1630 = n1627 & n1629 ;
  assign n1631 = n1629 & ~n1630 ;
  assign n1632 = n1627 & ~n1629 ;
  assign n1633 = n1617 & n1632 ;
  assign n1634 = ( n1617 & n1631 ) | ( n1617 & n1633 ) | ( n1631 & n1633 ) ;
  assign n1635 = n1617 | n1632 ;
  assign n1636 = n1631 | n1635 ;
  assign n1637 = ~n1634 & n1636 ;
  assign n1638 = n1603 & n1637 ;
  assign n1639 = ~n1605 & n1638 ;
  assign n1640 = ( n1607 & n1637 ) | ( n1607 & n1639 ) | ( n1637 & n1639 ) ;
  assign n1641 = n1603 | n1637 ;
  assign n1642 = ( ~n1605 & n1637 ) | ( ~n1605 & n1641 ) | ( n1637 & n1641 ) ;
  assign n1643 = n1607 | n1642 ;
  assign n1644 = ~n1640 & n1643 ;
  assign n1645 = n1553 & n1644 ;
  assign n1646 = n1553 | n1644 ;
  assign n1647 = ~n1645 & n1646 ;
  assign n1648 = n1480 & n1507 ;
  assign n1649 = ( n1480 & n1506 ) | ( n1480 & n1648 ) | ( n1506 & n1648 ) ;
  assign n1650 = n1505 | n1649 ;
  assign n1654 = ( n1647 & ~n1650 ) | ( n1647 & n1653 ) | ( ~n1650 & n1653 ) ;
  assign n1655 = ( ~n1647 & n1650 ) | ( ~n1647 & n1654 ) | ( n1650 & n1654 ) ;
  assign n1656 = ( ~n1653 & n1654 ) | ( ~n1653 & n1655 ) | ( n1654 & n1655 ) ;
  assign n1769 = n1647 & n1650 ;
  assign n1770 = n1647 | n1650 ;
  assign n1771 = n1769 | n1770 ;
  assign n1772 = ( n1652 & n1769 ) | ( n1652 & n1771 ) | ( n1769 & n1771 ) ;
  assign n1773 = ( n1651 & n1769 ) | ( n1651 & n1771 ) | ( n1769 & n1771 ) ;
  assign n1774 = ( n1385 & n1772 ) | ( n1385 & n1773 ) | ( n1772 & n1773 ) ;
  assign n1657 = n1630 | n1634 ;
  assign n1658 = x1 & x25 ;
  assign n1659 = n487 | n1658 ;
  assign n1660 = n487 & n1658 ;
  assign n1661 = n1659 & ~n1660 ;
  assign n1662 = ~n1621 & n1661 ;
  assign n1663 = n1621 & ~n1661 ;
  assign n1664 = n1662 | n1663 ;
  assign n1665 = n1590 & n1664 ;
  assign n1666 = n1590 | n1664 ;
  assign n1667 = ~n1665 & n1666 ;
  assign n1668 = n1579 & n1667 ;
  assign n1669 = ( n1600 & n1667 ) | ( n1600 & n1668 ) | ( n1667 & n1668 ) ;
  assign n1670 = n1579 | n1667 ;
  assign n1671 = n1600 | n1670 ;
  assign n1672 = ~n1669 & n1671 ;
  assign n1673 = n1657 & n1672 ;
  assign n1674 = n1657 | n1672 ;
  assign n1675 = ~n1673 & n1674 ;
  assign n1676 = n1606 & n1675 ;
  assign n1677 = ( n1640 & n1675 ) | ( n1640 & n1676 ) | ( n1675 & n1676 ) ;
  assign n1678 = n1606 | n1675 ;
  assign n1679 = n1640 | n1678 ;
  assign n1680 = ~n1677 & n1679 ;
  assign n1681 = x3 & x23 ;
  assign n1682 = x7 & x19 ;
  assign n1683 = n1681 & n1682 ;
  assign n1684 = x19 & x24 ;
  assign n1685 = n203 & n1684 ;
  assign n1686 = x23 & x24 ;
  assign n1687 = n77 & n1686 ;
  assign n1688 = n1685 | n1687 ;
  assign n1689 = x24 & n1683 ;
  assign n1690 = ( x24 & ~n1688 ) | ( x24 & n1689 ) | ( ~n1688 & n1689 ) ;
  assign n1691 = x2 & n1690 ;
  assign n1692 = ( n1681 & n1682 ) | ( n1681 & ~n1688 ) | ( n1682 & ~n1688 ) ;
  assign n1693 = ( ~n1683 & n1691 ) | ( ~n1683 & n1692 ) | ( n1691 & n1692 ) ;
  assign n1694 = x9 & x17 ;
  assign n1695 = n718 & n1694 ;
  assign n1696 = n360 & n1023 ;
  assign n1697 = n1695 | n1696 ;
  assign n1698 = n618 & n795 ;
  assign n1699 = n1694 & n1698 ;
  assign n1700 = ( n1694 & ~n1697 ) | ( n1694 & n1699 ) | ( ~n1697 & n1699 ) ;
  assign n1701 = n1697 | n1698 ;
  assign n1702 = x10 & x16 ;
  assign n1703 = ( n718 & ~n1698 ) | ( n718 & n1702 ) | ( ~n1698 & n1702 ) ;
  assign n1704 = n718 & n1702 ;
  assign n1705 = ( ~n1697 & n1703 ) | ( ~n1697 & n1704 ) | ( n1703 & n1704 ) ;
  assign n1706 = ~n1701 & n1705 ;
  assign n1707 = n1700 | n1706 ;
  assign n1708 = n1693 & n1707 ;
  assign n1709 = n1693 & ~n1708 ;
  assign n1710 = x20 & x22 ;
  assign n1711 = n274 & n1710 ;
  assign n1712 = n91 & n1585 ;
  assign n1713 = n1711 | n1712 ;
  assign n1714 = n204 & n1434 ;
  assign n1715 = x22 & n1714 ;
  assign n1716 = ( x22 & ~n1713 ) | ( x22 & n1715 ) | ( ~n1713 & n1715 ) ;
  assign n1717 = x4 & n1716 ;
  assign n1718 = n1713 | n1714 ;
  assign n1719 = x5 & x21 ;
  assign n1720 = x6 & x20 ;
  assign n1721 = ( ~n1714 & n1719 ) | ( ~n1714 & n1720 ) | ( n1719 & n1720 ) ;
  assign n1722 = n1719 & n1720 ;
  assign n1723 = ( ~n1713 & n1721 ) | ( ~n1713 & n1722 ) | ( n1721 & n1722 ) ;
  assign n1724 = ~n1718 & n1723 ;
  assign n1725 = n1717 | n1724 ;
  assign n1726 = ~n1693 & n1707 ;
  assign n1727 = n1725 & n1726 ;
  assign n1728 = ( n1709 & n1725 ) | ( n1709 & n1727 ) | ( n1725 & n1727 ) ;
  assign n1729 = n1725 | n1726 ;
  assign n1730 = n1709 | n1729 ;
  assign n1731 = ~n1728 & n1730 ;
  assign n1732 = n1541 | n1731 ;
  assign n1733 = n1546 | n1732 ;
  assign n1734 = n1541 & n1731 ;
  assign n1735 = ( n1546 & n1731 ) | ( n1546 & n1734 ) | ( n1731 & n1734 ) ;
  assign n1736 = n1733 & ~n1735 ;
  assign n1737 = n1442 | n1612 ;
  assign n1738 = ( n1612 & n1614 ) | ( n1612 & n1737 ) | ( n1614 & n1737 ) ;
  assign n1739 = n1531 & n1738 ;
  assign n1740 = ( n1536 & n1738 ) | ( n1536 & n1739 ) | ( n1738 & n1739 ) ;
  assign n1741 = n1531 | n1738 ;
  assign n1742 = n1536 | n1741 ;
  assign n1743 = ~n1740 & n1742 ;
  assign n1744 = n1561 | n1572 ;
  assign n1745 = n1561 & n1572 ;
  assign n1746 = n1744 & ~n1745 ;
  assign n1747 = x0 & x26 ;
  assign n1748 = x8 & x18 ;
  assign n1749 = n1747 | n1748 ;
  assign n1750 = ( n1609 & n1747 ) | ( n1609 & n1748 ) | ( n1747 & n1748 ) ;
  assign n1751 = n1749 & ~n1750 ;
  assign n1752 = n1747 & n1748 ;
  assign n1753 = n1749 & ~n1752 ;
  assign n1754 = n1609 & ~n1753 ;
  assign n1755 = n1751 | n1754 ;
  assign n1756 = n1746 & n1755 ;
  assign n1757 = n1746 & ~n1756 ;
  assign n1758 = ~n1746 & n1755 ;
  assign n1759 = n1757 | n1758 ;
  assign n1760 = n1743 & n1759 ;
  assign n1761 = n1743 | n1759 ;
  assign n1762 = ~n1760 & n1761 ;
  assign n1763 = ~n1736 & n1762 ;
  assign n1764 = n1736 & ~n1762 ;
  assign n1765 = n1763 | n1764 ;
  assign n1766 = n1680 & n1765 ;
  assign n1767 = ~n1680 & n1765 ;
  assign n1768 = ( n1680 & ~n1766 ) | ( n1680 & n1767 ) | ( ~n1766 & n1767 ) ;
  assign n1775 = n1550 | n1644 ;
  assign n1776 = ( n1550 & n1553 ) | ( n1550 & n1775 ) | ( n1553 & n1775 ) ;
  assign n1777 = ( n1768 & n1774 ) | ( n1768 & ~n1776 ) | ( n1774 & ~n1776 ) ;
  assign n1778 = ( ~n1768 & n1776 ) | ( ~n1768 & n1777 ) | ( n1776 & n1777 ) ;
  assign n1779 = ( ~n1774 & n1777 ) | ( ~n1774 & n1778 ) | ( n1777 & n1778 ) ;
  assign n1780 = n1768 & n1776 ;
  assign n1781 = n1768 | n1776 ;
  assign n1782 = n1774 & n1781 ;
  assign n1783 = n1780 | n1782 ;
  assign n1784 = x4 & x23 ;
  assign n1785 = x6 & x21 ;
  assign n1786 = n1784 & n1785 ;
  assign n1787 = x21 & x24 ;
  assign n1788 = n209 & n1787 ;
  assign n1789 = n79 & n1686 ;
  assign n1790 = n1788 | n1789 ;
  assign n1791 = x24 & n1786 ;
  assign n1792 = ( x24 & ~n1790 ) | ( x24 & n1791 ) | ( ~n1790 & n1791 ) ;
  assign n1793 = x3 & n1792 ;
  assign n1794 = ( n1784 & n1785 ) | ( n1784 & ~n1790 ) | ( n1785 & ~n1790 ) ;
  assign n1795 = ( ~n1786 & n1793 ) | ( ~n1786 & n1794 ) | ( n1793 & n1794 ) ;
  assign n1796 = x12 & x15 ;
  assign n1797 = n650 | n1796 ;
  assign n1798 = n647 & n792 ;
  assign n1799 = x5 & x22 ;
  assign n1800 = ~n1798 & n1799 ;
  assign n1801 = n1797 | n1798 ;
  assign n1802 = ( n1798 & n1800 ) | ( n1798 & n1801 ) | ( n1800 & n1801 ) ;
  assign n1803 = n1797 & ~n1802 ;
  assign n1804 = ( ~n1797 & n1798 ) | ( ~n1797 & n1799 ) | ( n1798 & n1799 ) ;
  assign n1805 = n1799 & n1804 ;
  assign n1806 = n1803 | n1805 ;
  assign n1807 = n1795 & n1806 ;
  assign n1808 = n1795 & ~n1807 ;
  assign n1809 = n1806 & ~n1807 ;
  assign n1810 = n1808 | n1809 ;
  assign n1811 = x0 & x27 ;
  assign n1812 = n1660 & ~n1811 ;
  assign n1813 = ~n1660 & n1811 ;
  assign n1814 = n1812 | n1813 ;
  assign n1815 = x1 & ~x26 ;
  assign n1816 = ( x1 & ~n539 ) | ( x1 & n1815 ) | ( ~n539 & n1815 ) ;
  assign n1817 = x26 & n1816 ;
  assign n1818 = x14 & ~x26 ;
  assign n1819 = ( x14 & ~n539 ) | ( x14 & n1818 ) | ( ~n539 & n1818 ) ;
  assign n1820 = n1817 | n1819 ;
  assign n1821 = n1814 & n1820 ;
  assign n1822 = n1814 | n1820 ;
  assign n1823 = ~n1821 & n1822 ;
  assign n1824 = ~n1810 & n1823 ;
  assign n1825 = n1810 & ~n1823 ;
  assign n1826 = n1824 | n1825 ;
  assign n1827 = n1701 | n1718 ;
  assign n1828 = n1701 & n1718 ;
  assign n1829 = n1827 & ~n1828 ;
  assign n1830 = n1683 | n1688 ;
  assign n1831 = n1829 | n1830 ;
  assign n1832 = n1829 & n1830 ;
  assign n1833 = n1831 & ~n1832 ;
  assign n1834 = n1740 | n1833 ;
  assign n1835 = n1760 | n1834 ;
  assign n1836 = ( n1740 & n1760 ) | ( n1740 & n1833 ) | ( n1760 & n1833 ) ;
  assign n1837 = n1835 & ~n1836 ;
  assign n1838 = n1826 & n1837 ;
  assign n1839 = n1826 | n1837 ;
  assign n1840 = ~n1838 & n1839 ;
  assign n1841 = n1541 | n1546 ;
  assign n1842 = ( n1731 & n1762 ) | ( n1731 & n1841 ) | ( n1762 & n1841 ) ;
  assign n1843 = n1840 | n1842 ;
  assign n1844 = n1840 & n1842 ;
  assign n1845 = n1843 & ~n1844 ;
  assign n1846 = x11 & x16 ;
  assign n1847 = x20 & x25 ;
  assign n1848 = n203 & n1847 ;
  assign n1849 = x2 & x25 ;
  assign n1850 = x7 & x20 ;
  assign n1851 = n1849 | n1850 ;
  assign n1852 = ~n1848 & n1851 ;
  assign n1853 = n1846 | n1852 ;
  assign n1854 = n1846 & n1852 ;
  assign n1855 = n1853 & ~n1854 ;
  assign n1856 = n1750 | n1855 ;
  assign n1857 = n1750 & n1855 ;
  assign n1858 = n1856 & ~n1857 ;
  assign n1859 = x8 & x19 ;
  assign n1860 = x10 & x17 ;
  assign n1861 = n1859 & n1860 ;
  assign n1862 = n313 & n1077 ;
  assign n1863 = n1861 | n1862 ;
  assign n1864 = n360 & n1020 ;
  assign n1865 = n1859 & n1864 ;
  assign n1866 = ( n1859 & ~n1863 ) | ( n1859 & n1865 ) | ( ~n1863 & n1865 ) ;
  assign n1867 = n1863 | n1864 ;
  assign n1868 = x9 & x18 ;
  assign n1869 = ( n1860 & ~n1864 ) | ( n1860 & n1868 ) | ( ~n1864 & n1868 ) ;
  assign n1870 = n1860 & n1868 ;
  assign n1871 = ( ~n1863 & n1869 ) | ( ~n1863 & n1870 ) | ( n1869 & n1870 ) ;
  assign n1872 = ~n1867 & n1871 ;
  assign n1873 = n1866 | n1872 ;
  assign n1874 = ~n1858 & n1873 ;
  assign n1875 = n1858 & ~n1873 ;
  assign n1876 = n1874 | n1875 ;
  assign n1877 = n1669 | n1876 ;
  assign n1878 = n1673 | n1877 ;
  assign n1879 = n1669 & n1876 ;
  assign n1880 = ( n1673 & n1876 ) | ( n1673 & n1879 ) | ( n1876 & n1879 ) ;
  assign n1881 = n1878 & ~n1880 ;
  assign n1882 = n1621 & n1661 ;
  assign n1883 = n1665 | n1882 ;
  assign n1884 = n1745 | n1755 ;
  assign n1885 = ( n1745 & n1746 ) | ( n1745 & n1884 ) | ( n1746 & n1884 ) ;
  assign n1886 = n1883 | n1885 ;
  assign n1887 = n1883 & n1885 ;
  assign n1888 = n1886 & ~n1887 ;
  assign n1889 = n1708 | n1728 ;
  assign n1890 = n1888 | n1889 ;
  assign n1891 = n1888 & n1889 ;
  assign n1892 = n1890 & ~n1891 ;
  assign n1893 = n1881 & n1892 ;
  assign n1894 = n1881 | n1892 ;
  assign n1895 = ~n1893 & n1894 ;
  assign n1896 = n1845 & n1895 ;
  assign n1897 = n1845 | n1895 ;
  assign n1898 = ~n1896 & n1897 ;
  assign n1899 = n1677 | n1765 ;
  assign n1900 = ( n1677 & n1680 ) | ( n1677 & n1899 ) | ( n1680 & n1899 ) ;
  assign n1901 = ( n1783 & ~n1898 ) | ( n1783 & n1900 ) | ( ~n1898 & n1900 ) ;
  assign n1902 = ( n1898 & ~n1900 ) | ( n1898 & n1901 ) | ( ~n1900 & n1901 ) ;
  assign n1903 = ( ~n1783 & n1901 ) | ( ~n1783 & n1902 ) | ( n1901 & n1902 ) ;
  assign n1904 = n1898 & n1900 ;
  assign n1905 = n1898 | n1900 ;
  assign n1906 = n1904 | n1905 ;
  assign n1907 = ( n1780 & n1904 ) | ( n1780 & n1906 ) | ( n1904 & n1906 ) ;
  assign n1908 = ( n1782 & n1906 ) | ( n1782 & n1907 ) | ( n1906 & n1907 ) ;
  assign n1909 = x3 & x25 ;
  assign n1910 = x4 & x24 ;
  assign n1911 = n1909 | n1910 ;
  assign n1912 = x24 & x25 ;
  assign n1913 = n79 & n1912 ;
  assign n1914 = x8 & x20 ;
  assign n1915 = ~n1913 & n1914 ;
  assign n1916 = n1911 | n1913 ;
  assign n1917 = ( n1913 & n1915 ) | ( n1913 & n1916 ) | ( n1915 & n1916 ) ;
  assign n1918 = n1911 & ~n1917 ;
  assign n1919 = ( n1660 & n1811 ) | ( n1660 & n1819 ) | ( n1811 & n1819 ) ;
  assign n1920 = n1660 | n1811 ;
  assign n1921 = ( n1817 & n1919 ) | ( n1817 & n1920 ) | ( n1919 & n1920 ) ;
  assign n1922 = ( ~n1911 & n1913 ) | ( ~n1911 & n1914 ) | ( n1913 & n1914 ) ;
  assign n1923 = n1914 & n1922 ;
  assign n1924 = ~n1921 & n1923 ;
  assign n1925 = ( n1918 & ~n1921 ) | ( n1918 & n1924 ) | ( ~n1921 & n1924 ) ;
  assign n1926 = n1921 & ~n1923 ;
  assign n1927 = ~n1918 & n1926 ;
  assign n1928 = n1925 | n1927 ;
  assign n1929 = n135 & n1337 ;
  assign n1930 = n200 & n1585 ;
  assign n1931 = n1929 | n1930 ;
  assign n1932 = x22 & x23 ;
  assign n1933 = n204 & n1932 ;
  assign n1934 = x21 & n1933 ;
  assign n1935 = ( x21 & ~n1931 ) | ( x21 & n1934 ) | ( ~n1931 & n1934 ) ;
  assign n1936 = x7 & n1935 ;
  assign n1937 = n1931 | n1933 ;
  assign n1938 = x5 & x23 ;
  assign n1939 = x6 & x22 ;
  assign n1940 = ( ~n1933 & n1938 ) | ( ~n1933 & n1939 ) | ( n1938 & n1939 ) ;
  assign n1941 = n1938 & n1939 ;
  assign n1942 = ( ~n1931 & n1940 ) | ( ~n1931 & n1941 ) | ( n1940 & n1941 ) ;
  assign n1943 = ~n1937 & n1942 ;
  assign n1944 = n1936 | n1943 ;
  assign n1945 = n1928 & n1944 ;
  assign n1946 = n1928 | n1944 ;
  assign n1947 = ~n1945 & n1946 ;
  assign n1948 = n1826 | n1836 ;
  assign n1949 = ( n1836 & n1837 ) | ( n1836 & n1948 ) | ( n1837 & n1948 ) ;
  assign n1950 = n1947 | n1949 ;
  assign n1951 = n1947 & n1949 ;
  assign n1952 = n1950 & ~n1951 ;
  assign n1953 = x26 & n539 ;
  assign n1954 = x1 & x27 ;
  assign n1955 = n723 & n1954 ;
  assign n1956 = n723 | n1954 ;
  assign n1957 = ~n1955 & n1956 ;
  assign n1958 = ~n1953 & n1957 ;
  assign n1959 = n1953 & ~n1957 ;
  assign n1960 = n1958 | n1959 ;
  assign n1961 = n1802 & n1960 ;
  assign n1962 = n1802 | n1960 ;
  assign n1963 = ~n1961 & n1962 ;
  assign n1964 = n1857 | n1873 ;
  assign n1965 = ( n1857 & n1858 ) | ( n1857 & n1964 ) | ( n1858 & n1964 ) ;
  assign n1966 = n1963 & n1965 ;
  assign n1967 = n1963 | n1965 ;
  assign n1968 = ~n1966 & n1967 ;
  assign n1969 = ( n1795 & n1806 ) | ( n1795 & n1823 ) | ( n1806 & n1823 ) ;
  assign n1970 = n1968 | n1969 ;
  assign n1971 = n1968 & n1969 ;
  assign n1972 = n1970 & ~n1971 ;
  assign n1973 = n1952 & n1972 ;
  assign n1974 = n1952 | n1972 ;
  assign n1975 = ~n1973 & n1974 ;
  assign n1976 = n1786 | n1790 ;
  assign n1977 = n1867 | n1976 ;
  assign n1978 = n1867 & n1976 ;
  assign n1979 = n1977 & ~n1978 ;
  assign n1980 = n1846 | n1848 ;
  assign n1981 = ( n1848 & n1852 ) | ( n1848 & n1980 ) | ( n1852 & n1980 ) ;
  assign n1982 = n1979 | n1981 ;
  assign n1983 = n1979 & n1981 ;
  assign n1984 = n1982 & ~n1983 ;
  assign n1985 = n1887 & n1984 ;
  assign n1986 = ( n1888 & n1984 ) | ( n1888 & n1985 ) | ( n1984 & n1985 ) ;
  assign n1987 = n1984 & n1985 ;
  assign n1988 = ( n1889 & n1986 ) | ( n1889 & n1987 ) | ( n1986 & n1987 ) ;
  assign n1989 = n1887 | n1984 ;
  assign n1990 = n1888 | n1989 ;
  assign n1991 = ( n1889 & n1989 ) | ( n1889 & n1990 ) | ( n1989 & n1990 ) ;
  assign n1992 = ~n1988 & n1991 ;
  assign n1993 = x0 & x28 ;
  assign n1994 = x12 & x16 ;
  assign n1995 = n1993 & n1994 ;
  assign n1996 = x11 & x28 ;
  assign n1997 = n707 & n1996 ;
  assign n1998 = n490 & n1023 ;
  assign n1999 = n1997 | n1998 ;
  assign n2000 = x17 & n1995 ;
  assign n2001 = ( x17 & ~n1999 ) | ( x17 & n2000 ) | ( ~n1999 & n2000 ) ;
  assign n2002 = x11 & n2001 ;
  assign n2003 = ( n1993 & n1994 ) | ( n1993 & ~n1999 ) | ( n1994 & ~n1999 ) ;
  assign n2004 = ( ~n1995 & n2002 ) | ( ~n1995 & n2003 ) | ( n2002 & n2003 ) ;
  assign n2005 = x9 & x19 ;
  assign n2006 = x10 & x18 ;
  assign n2007 = n2005 | n2006 ;
  assign n2008 = n360 & n1077 ;
  assign n2009 = x2 & x26 ;
  assign n2010 = ~n2008 & n2009 ;
  assign n2011 = n2007 | n2008 ;
  assign n2012 = ( n2008 & n2010 ) | ( n2008 & n2011 ) | ( n2010 & n2011 ) ;
  assign n2013 = n2007 & ~n2012 ;
  assign n2014 = ~n2007 & n2009 ;
  assign n2015 = ( n2009 & ~n2010 ) | ( n2009 & n2014 ) | ( ~n2010 & n2014 ) ;
  assign n2016 = n2013 | n2015 ;
  assign n2017 = n2004 & n2016 ;
  assign n2018 = n2004 & ~n2017 ;
  assign n2019 = n2016 & ~n2017 ;
  assign n2020 = n2018 | n2019 ;
  assign n2021 = n1828 | n1830 ;
  assign n2022 = ( n1828 & n1829 ) | ( n1828 & n2021 ) | ( n1829 & n2021 ) ;
  assign n2023 = n2020 | n2022 ;
  assign n2024 = n2020 & n2022 ;
  assign n2025 = n2023 & ~n2024 ;
  assign n2026 = n1992 & n2025 ;
  assign n2027 = n1992 | n2025 ;
  assign n2028 = ~n2026 & n2027 ;
  assign n2029 = n1669 | n1673 ;
  assign n2030 = ( n1876 & n1892 ) | ( n1876 & n2029 ) | ( n1892 & n2029 ) ;
  assign n2031 = n2028 | n2030 ;
  assign n2032 = n2028 & n2030 ;
  assign n2033 = n2031 & ~n2032 ;
  assign n2034 = n1844 & n2033 ;
  assign n2035 = ( n1896 & n2033 ) | ( n1896 & n2034 ) | ( n2033 & n2034 ) ;
  assign n2036 = n1844 | n2033 ;
  assign n2037 = n1896 | n2036 ;
  assign n2038 = ~n2035 & n2037 ;
  assign n2039 = ( n1908 & n1975 ) | ( n1908 & ~n2038 ) | ( n1975 & ~n2038 ) ;
  assign n2040 = ( ~n1975 & n2038 ) | ( ~n1975 & n2039 ) | ( n2038 & n2039 ) ;
  assign n2041 = ( ~n1908 & n2039 ) | ( ~n1908 & n2040 ) | ( n2039 & n2040 ) ;
  assign n2042 = n1975 & n2038 ;
  assign n2043 = n1975 | n2038 ;
  assign n2044 = n1906 & n2043 ;
  assign n2045 = n1907 & n2043 ;
  assign n2046 = ( n1781 & n2044 ) | ( n1781 & n2045 ) | ( n2044 & n2045 ) ;
  assign n2047 = n2044 & n2045 ;
  assign n2048 = ( n1774 & n2046 ) | ( n1774 & n2047 ) | ( n2046 & n2047 ) ;
  assign n2049 = n2042 | n2048 ;
  assign n2050 = n1963 | n1969 ;
  assign n2051 = ( n1965 & n1969 ) | ( n1965 & n2050 ) | ( n1969 & n2050 ) ;
  assign n2052 = ( n1966 & n1968 ) | ( n1966 & n2051 ) | ( n1968 & n2051 ) ;
  assign n2053 = n1988 | n2025 ;
  assign n2054 = ( n1988 & n1992 ) | ( n1988 & n2053 ) | ( n1992 & n2053 ) ;
  assign n2055 = n2052 | n2054 ;
  assign n2056 = n2052 & n2054 ;
  assign n2057 = n2055 & ~n2056 ;
  assign n2058 = n1918 | n1923 ;
  assign n2059 = ( n1921 & n1944 ) | ( n1921 & n2058 ) | ( n1944 & n2058 ) ;
  assign n2060 = n2017 | n2022 ;
  assign n2061 = n2059 | n2060 ;
  assign n2062 = n2017 | n2059 ;
  assign n2063 = ( n2020 & n2061 ) | ( n2020 & n2062 ) | ( n2061 & n2062 ) ;
  assign n2064 = n2059 & n2060 ;
  assign n2065 = n2017 & n2059 ;
  assign n2066 = ( n2020 & n2064 ) | ( n2020 & n2065 ) | ( n2064 & n2065 ) ;
  assign n2067 = n2063 & ~n2066 ;
  assign n2068 = n1995 | n1999 ;
  assign n2069 = n2012 | n2068 ;
  assign n2070 = n2012 & n2068 ;
  assign n2071 = n2069 & ~n2070 ;
  assign n2072 = x0 & x29 ;
  assign n2073 = x2 & x27 ;
  assign n2074 = n2072 | n2073 ;
  assign n2075 = x27 & x29 ;
  assign n2076 = n67 & n2075 ;
  assign n2077 = n2074 & ~n2076 ;
  assign n2078 = n1955 | n2076 ;
  assign n2079 = ( n2076 & n2077 ) | ( n2076 & n2078 ) | ( n2077 & n2078 ) ;
  assign n2080 = n2074 & ~n2079 ;
  assign n2081 = n1955 & ~n2077 ;
  assign n2082 = n2080 | n2081 ;
  assign n2083 = n2071 & n2082 ;
  assign n2084 = n2071 & ~n2083 ;
  assign n2085 = n2082 & ~n2083 ;
  assign n2086 = n2084 | n2085 ;
  assign n2087 = n2067 & n2086 ;
  assign n2088 = n2067 | n2086 ;
  assign n2089 = ~n2087 & n2088 ;
  assign n2090 = ~n2057 & n2089 ;
  assign n2091 = n2057 & ~n2089 ;
  assign n2092 = n2090 | n2091 ;
  assign n2093 = ( n1947 & n1949 ) | ( n1947 & n1972 ) | ( n1949 & n1972 ) ;
  assign n2094 = ( n1802 & n1953 ) | ( n1802 & n1957 ) | ( n1953 & n1957 ) ;
  assign n2095 = x13 & x16 ;
  assign n2096 = n792 | n2095 ;
  assign n2097 = x6 & x23 ;
  assign n2098 = ( n792 & n2095 ) | ( n792 & n2097 ) | ( n2095 & n2097 ) ;
  assign n2099 = n2096 & ~n2098 ;
  assign n2100 = n792 & n2095 ;
  assign n2101 = n2097 & ~n2100 ;
  assign n2102 = ~n2096 & n2097 ;
  assign n2103 = ( n2097 & ~n2101 ) | ( n2097 & n2102 ) | ( ~n2101 & n2102 ) ;
  assign n2104 = n2099 | n2103 ;
  assign n2105 = n2094 & n2104 ;
  assign n2106 = n2094 & ~n2105 ;
  assign n2107 = n2104 & ~n2105 ;
  assign n2108 = n2106 | n2107 ;
  assign n2109 = n1978 | n1981 ;
  assign n2110 = ( n1978 & n1979 ) | ( n1978 & n2109 ) | ( n1979 & n2109 ) ;
  assign n2111 = n2108 | n2110 ;
  assign n2112 = n2108 & n2110 ;
  assign n2113 = n2111 & ~n2112 ;
  assign n2114 = n969 & n1285 ;
  assign n2115 = n360 & n1437 ;
  assign n2116 = n2114 | n2115 ;
  assign n2117 = n618 & n1077 ;
  assign n2118 = x20 & n2117 ;
  assign n2119 = ( x20 & ~n2116 ) | ( x20 & n2118 ) | ( ~n2116 & n2118 ) ;
  assign n2120 = x9 & n2119 ;
  assign n2121 = n2116 | n2117 ;
  assign n2122 = x10 & x19 ;
  assign n2123 = x11 & x18 ;
  assign n2124 = ( ~n2117 & n2122 ) | ( ~n2117 & n2123 ) | ( n2122 & n2123 ) ;
  assign n2125 = n2122 & n2123 ;
  assign n2126 = ( ~n2116 & n2124 ) | ( ~n2116 & n2125 ) | ( n2124 & n2125 ) ;
  assign n2127 = ~n2121 & n2126 ;
  assign n2128 = n2120 | n2127 ;
  assign n2129 = x3 & x26 ;
  assign n2130 = x8 & x21 ;
  assign n2131 = n2129 | n2130 ;
  assign n2132 = x21 & x26 ;
  assign n2133 = n311 & n2132 ;
  assign n2134 = n2131 | n2133 ;
  assign n2135 = x12 & x17 ;
  assign n2136 = ( ~n2133 & n2134 ) | ( ~n2133 & n2135 ) | ( n2134 & n2135 ) ;
  assign n2137 = ( n2133 & n2134 ) | ( n2133 & ~n2135 ) | ( n2134 & ~n2135 ) ;
  assign n2138 = ( ~n2134 & n2136 ) | ( ~n2134 & n2137 ) | ( n2136 & n2137 ) ;
  assign n2139 = n2128 & n2138 ;
  assign n2140 = n2128 & ~n2139 ;
  assign n2141 = ~n2128 & n2138 ;
  assign n2142 = n2140 | n2141 ;
  assign n2143 = x4 & x25 ;
  assign n2144 = n91 & n1912 ;
  assign n2145 = x7 & x22 ;
  assign n2146 = n2143 & n2145 ;
  assign n2147 = n2144 | n2146 ;
  assign n2148 = x22 & x24 ;
  assign n2149 = n135 & n2148 ;
  assign n2150 = n2143 & n2149 ;
  assign n2151 = ( n2143 & ~n2147 ) | ( n2143 & n2150 ) | ( ~n2147 & n2150 ) ;
  assign n2152 = n2147 | n2149 ;
  assign n2153 = x5 & x24 ;
  assign n2154 = ( n2145 & ~n2149 ) | ( n2145 & n2153 ) | ( ~n2149 & n2153 ) ;
  assign n2155 = n2145 & n2153 ;
  assign n2156 = ( ~n2147 & n2154 ) | ( ~n2147 & n2155 ) | ( n2154 & n2155 ) ;
  assign n2157 = ~n2152 & n2156 ;
  assign n2158 = n2151 | n2157 ;
  assign n2159 = n2141 & n2158 ;
  assign n2160 = ( n2140 & n2158 ) | ( n2140 & n2159 ) | ( n2158 & n2159 ) ;
  assign n2161 = n2142 & ~n2160 ;
  assign n2162 = x28 & n668 ;
  assign n2163 = x1 & x28 ;
  assign n2164 = x15 | n2163 ;
  assign n2165 = ~n2162 & n2164 ;
  assign n2166 = n1937 | n2165 ;
  assign n2167 = n1937 & n2165 ;
  assign n2168 = n2166 & ~n2167 ;
  assign n2169 = n1917 & n2168 ;
  assign n2170 = n1917 | n2168 ;
  assign n2171 = ~n2169 & n2170 ;
  assign n2172 = n2158 & n2171 ;
  assign n2173 = ~n2142 & n2172 ;
  assign n2174 = ( n2161 & n2171 ) | ( n2161 & n2173 ) | ( n2171 & n2173 ) ;
  assign n2175 = ( n2158 & ~n2160 ) | ( n2158 & n2171 ) | ( ~n2160 & n2171 ) ;
  assign n2176 = ( n2142 & ~n2160 ) | ( n2142 & n2175 ) | ( ~n2160 & n2175 ) ;
  assign n2177 = ~n2174 & n2176 ;
  assign n2178 = n2113 & n2177 ;
  assign n2179 = n2113 | n2177 ;
  assign n2180 = ~n2178 & n2179 ;
  assign n2181 = n2093 & n2180 ;
  assign n2182 = n2093 & ~n2181 ;
  assign n2183 = ~n2093 & n2180 ;
  assign n2184 = n2182 | n2183 ;
  assign n2185 = n2092 & n2184 ;
  assign n2186 = ( ~n2092 & n2182 ) | ( ~n2092 & n2183 ) | ( n2182 & n2183 ) ;
  assign n2187 = n2092 | n2186 ;
  assign n2188 = ~n2185 & n2187 ;
  assign n2189 = n2032 | n2035 ;
  assign n2190 = ( n2049 & n2188 ) | ( n2049 & ~n2189 ) | ( n2188 & ~n2189 ) ;
  assign n2191 = ( ~n2188 & n2189 ) | ( ~n2188 & n2190 ) | ( n2189 & n2190 ) ;
  assign n2192 = ( ~n2049 & n2190 ) | ( ~n2049 & n2191 ) | ( n2190 & n2191 ) ;
  assign n2193 = n2188 & n2189 ;
  assign n2194 = n2188 | n2189 ;
  assign n2195 = n2193 | n2194 ;
  assign n2196 = ( n2049 & n2193 ) | ( n2049 & n2195 ) | ( n2193 & n2195 ) ;
  assign n2197 = n2181 | n2185 ;
  assign n2198 = x0 & x30 ;
  assign n2199 = n2162 & n2198 ;
  assign n2200 = n2162 & ~n2199 ;
  assign n2201 = ~n2162 & n2198 ;
  assign n2202 = n2200 | n2201 ;
  assign n2203 = x1 & x29 ;
  assign n2204 = n790 & n2203 ;
  assign n2205 = n2203 & ~n2204 ;
  assign n2206 = n790 & ~n2204 ;
  assign n2207 = n2205 | n2206 ;
  assign n2208 = ~n2202 & n2207 ;
  assign n2209 = n2202 & ~n2207 ;
  assign n2210 = n2208 | n2209 ;
  assign n2211 = n1917 | n2167 ;
  assign n2212 = ( n2167 & n2168 ) | ( n2167 & n2211 ) | ( n2168 & n2211 ) ;
  assign n2213 = n2210 | n2212 ;
  assign n2214 = n2210 & n2212 ;
  assign n2215 = n2213 & ~n2214 ;
  assign n2216 = n2070 | n2083 ;
  assign n2217 = n2215 | n2216 ;
  assign n2218 = n2215 & n2216 ;
  assign n2219 = n2217 & ~n2218 ;
  assign n2220 = n2113 | n2174 ;
  assign n2221 = ( n2174 & n2177 ) | ( n2174 & n2220 ) | ( n2177 & n2220 ) ;
  assign n2222 = n2219 | n2221 ;
  assign n2223 = n2219 & n2221 ;
  assign n2224 = n2222 & ~n2223 ;
  assign n2225 = n2098 | n2149 ;
  assign n2226 = n2147 | n2225 ;
  assign n2227 = n2098 & n2149 ;
  assign n2228 = ( n2098 & n2147 ) | ( n2098 & n2227 ) | ( n2147 & n2227 ) ;
  assign n2229 = n2226 & ~n2228 ;
  assign n2230 = x2 & x28 ;
  assign n2231 = x9 & x21 ;
  assign n2232 = n2230 | n2231 ;
  assign n2233 = x13 & x17 ;
  assign n2234 = ( n2230 & n2231 ) | ( n2230 & n2233 ) | ( n2231 & n2233 ) ;
  assign n2235 = n2232 & ~n2234 ;
  assign n2236 = n2230 & n2231 ;
  assign n2237 = n2233 & ~n2236 ;
  assign n2238 = ~n2232 & n2233 ;
  assign n2239 = ( n2233 & ~n2237 ) | ( n2233 & n2238 ) | ( ~n2237 & n2238 ) ;
  assign n2240 = n2235 | n2239 ;
  assign n2241 = n2229 & n2240 ;
  assign n2242 = n2229 & ~n2241 ;
  assign n2243 = n2240 & ~n2241 ;
  assign n2244 = n2242 | n2243 ;
  assign n2245 = n2139 | n2244 ;
  assign n2246 = n2160 | n2245 ;
  assign n2247 = n2139 & n2244 ;
  assign n2248 = ( n2160 & n2244 ) | ( n2160 & n2247 ) | ( n2244 & n2247 ) ;
  assign n2249 = n2246 & ~n2248 ;
  assign n2250 = ~n2133 & n2135 ;
  assign n2251 = ( n2133 & n2134 ) | ( n2133 & n2250 ) | ( n2134 & n2250 ) ;
  assign n2252 = n2121 | n2251 ;
  assign n2253 = n2121 & n2251 ;
  assign n2254 = n2252 & ~n2253 ;
  assign n2255 = n2079 | n2254 ;
  assign n2256 = n2079 & n2254 ;
  assign n2257 = n2255 & ~n2256 ;
  assign n2258 = n2249 & n2257 ;
  assign n2259 = n2249 | n2257 ;
  assign n2260 = ~n2258 & n2259 ;
  assign n2261 = n2224 & n2260 ;
  assign n2262 = n2224 | n2260 ;
  assign n2263 = ~n2261 & n2262 ;
  assign n2312 = n2105 | n2110 ;
  assign n2313 = ( n2105 & n2108 ) | ( n2105 & n2312 ) | ( n2108 & n2312 ) ;
  assign n2264 = x4 & x26 ;
  assign n2265 = x8 & x22 ;
  assign n2266 = n2264 & n2265 ;
  assign n2267 = x26 & x27 ;
  assign n2268 = n79 & n2267 ;
  assign n2269 = x8 & x27 ;
  assign n2270 = n1591 & n2269 ;
  assign n2271 = n2268 | n2270 ;
  assign n2272 = x27 & n2266 ;
  assign n2273 = ( x27 & ~n2271 ) | ( x27 & n2272 ) | ( ~n2271 & n2272 ) ;
  assign n2274 = x3 & n2273 ;
  assign n2275 = ( n2264 & n2265 ) | ( n2264 & ~n2271 ) | ( n2265 & ~n2271 ) ;
  assign n2276 = ( ~n2266 & n2274 ) | ( ~n2266 & n2275 ) | ( n2274 & n2275 ) ;
  assign n2277 = n135 & n1557 ;
  assign n2278 = n204 & n1912 ;
  assign n2279 = n2277 | n2278 ;
  assign n2280 = n200 & n1686 ;
  assign n2281 = x25 & n2280 ;
  assign n2282 = ( x25 & ~n2279 ) | ( x25 & n2281 ) | ( ~n2279 & n2281 ) ;
  assign n2283 = x5 & n2282 ;
  assign n2284 = n2279 | n2280 ;
  assign n2285 = x6 & x24 ;
  assign n2286 = x7 & x23 ;
  assign n2287 = ( ~n2280 & n2285 ) | ( ~n2280 & n2286 ) | ( n2285 & n2286 ) ;
  assign n2288 = n2285 & n2286 ;
  assign n2289 = ( ~n2279 & n2287 ) | ( ~n2279 & n2288 ) | ( n2287 & n2288 ) ;
  assign n2290 = ~n2284 & n2289 ;
  assign n2291 = n2283 | n2290 ;
  assign n2292 = n2276 & n2291 ;
  assign n2293 = n2276 & ~n2292 ;
  assign n2294 = n2291 & ~n2292 ;
  assign n2295 = n2293 | n2294 ;
  assign n2296 = n363 & n1285 ;
  assign n2297 = n618 & n1437 ;
  assign n2298 = n2296 | n2297 ;
  assign n2299 = n490 & n1077 ;
  assign n2300 = x20 & n2299 ;
  assign n2301 = ( x20 & ~n2298 ) | ( x20 & n2300 ) | ( ~n2298 & n2300 ) ;
  assign n2302 = x10 & n2301 ;
  assign n2303 = n2298 | n2299 ;
  assign n2304 = x11 & x19 ;
  assign n2305 = x12 & x18 ;
  assign n2306 = ( ~n2299 & n2304 ) | ( ~n2299 & n2305 ) | ( n2304 & n2305 ) ;
  assign n2307 = n2304 & n2305 ;
  assign n2308 = ( ~n2298 & n2306 ) | ( ~n2298 & n2307 ) | ( n2306 & n2307 ) ;
  assign n2309 = ~n2303 & n2308 ;
  assign n2310 = n2302 | n2309 ;
  assign n2311 = ~n2295 & n2310 ;
  assign n2314 = n2311 & n2313 ;
  assign n2315 = n2295 & ~n2310 ;
  assign n2316 = ( n2313 & n2314 ) | ( n2313 & n2315 ) | ( n2314 & n2315 ) ;
  assign n2317 = n2311 | n2313 ;
  assign n2318 = n2315 | n2317 ;
  assign n2319 = ~n2316 & n2318 ;
  assign n2320 = ( n2017 & n2020 ) | ( n2017 & n2060 ) | ( n2020 & n2060 ) ;
  assign n2321 = ( n2059 & n2086 ) | ( n2059 & n2320 ) | ( n2086 & n2320 ) ;
  assign n2322 = n2319 | n2321 ;
  assign n2323 = n2319 & n2321 ;
  assign n2324 = n2322 & ~n2323 ;
  assign n2325 = n2056 | n2089 ;
  assign n2326 = ( n2056 & n2057 ) | ( n2056 & n2325 ) | ( n2057 & n2325 ) ;
  assign n2327 = n2324 & n2326 ;
  assign n2328 = n2324 | n2326 ;
  assign n2329 = ~n2327 & n2328 ;
  assign n2330 = n2263 & n2329 ;
  assign n2331 = n2263 | n2329 ;
  assign n2332 = ~n2330 & n2331 ;
  assign n2333 = ( n2196 & n2197 ) | ( n2196 & ~n2332 ) | ( n2197 & ~n2332 ) ;
  assign n2334 = ( ~n2197 & n2332 ) | ( ~n2197 & n2333 ) | ( n2332 & n2333 ) ;
  assign n2335 = ( ~n2196 & n2333 ) | ( ~n2196 & n2334 ) | ( n2333 & n2334 ) ;
  assign n2490 = n2197 & n2332 ;
  assign n2491 = n2197 | n2332 ;
  assign n2492 = n2193 & n2491 ;
  assign n2493 = n2490 | n2492 ;
  assign n2494 = n2490 | n2491 ;
  assign n2495 = ( n2195 & n2490 ) | ( n2195 & n2494 ) | ( n2490 & n2494 ) ;
  assign n2496 = ( n2042 & n2493 ) | ( n2042 & n2495 ) | ( n2493 & n2495 ) ;
  assign n2497 = n2493 | n2495 ;
  assign n2498 = ( n2048 & n2496 ) | ( n2048 & n2497 ) | ( n2496 & n2497 ) ;
  assign n2336 = x23 & x26 ;
  assign n2337 = n222 & n2336 ;
  assign n2338 = n251 & n1686 ;
  assign n2339 = n2337 | n2338 ;
  assign n2340 = x24 & x26 ;
  assign n2341 = n135 & n2340 ;
  assign n2342 = x23 & n2341 ;
  assign n2343 = ( x23 & ~n2339 ) | ( x23 & n2342 ) | ( ~n2339 & n2342 ) ;
  assign n2344 = x8 & n2343 ;
  assign n2345 = n2339 | n2341 ;
  assign n2346 = x5 & x26 ;
  assign n2347 = x7 & x24 ;
  assign n2348 = ( ~n2341 & n2346 ) | ( ~n2341 & n2347 ) | ( n2346 & n2347 ) ;
  assign n2349 = n2346 & n2347 ;
  assign n2350 = ( ~n2339 & n2348 ) | ( ~n2339 & n2349 ) | ( n2348 & n2349 ) ;
  assign n2351 = ~n2345 & n2350 ;
  assign n2352 = n2344 | n2351 ;
  assign n2353 = x14 & x17 ;
  assign n2354 = n795 | n2353 ;
  assign n2355 = n792 & n1023 ;
  assign n2356 = x6 & x25 ;
  assign n2357 = ~n2355 & n2356 ;
  assign n2358 = n2354 | n2355 ;
  assign n2359 = ( n2355 & n2357 ) | ( n2355 & n2358 ) | ( n2357 & n2358 ) ;
  assign n2360 = n2354 & ~n2359 ;
  assign n2361 = ( ~n2354 & n2355 ) | ( ~n2354 & n2356 ) | ( n2355 & n2356 ) ;
  assign n2362 = n2356 & n2361 ;
  assign n2363 = n2360 | n2362 ;
  assign n2364 = n2352 & n2363 ;
  assign n2365 = n2352 & ~n2364 ;
  assign n2366 = n2363 & ~n2364 ;
  assign n2367 = n2365 | n2366 ;
  assign n2368 = n119 & n2075 ;
  assign n2369 = x28 & x29 ;
  assign n2370 = n77 & n2369 ;
  assign n2371 = n2368 | n2370 ;
  assign n2372 = x27 & x28 ;
  assign n2373 = n79 & n2372 ;
  assign n2374 = x29 & n2373 ;
  assign n2375 = ( x29 & ~n2371 ) | ( x29 & n2374 ) | ( ~n2371 & n2374 ) ;
  assign n2376 = x2 & n2375 ;
  assign n2377 = n2371 | n2373 ;
  assign n2378 = x3 & x28 ;
  assign n2379 = x4 & x27 ;
  assign n2380 = ( ~n2373 & n2378 ) | ( ~n2373 & n2379 ) | ( n2378 & n2379 ) ;
  assign n2381 = n2378 & n2379 ;
  assign n2382 = ( ~n2371 & n2380 ) | ( ~n2371 & n2381 ) | ( n2380 & n2381 ) ;
  assign n2383 = ~n2377 & n2382 ;
  assign n2384 = n2376 | n2383 ;
  assign n2385 = ~n2367 & n2384 ;
  assign n2386 = n2367 & ~n2384 ;
  assign n2387 = n2385 | n2386 ;
  assign n2420 = n2199 | n2207 ;
  assign n2421 = ( n2199 & n2202 ) | ( n2199 & n2420 ) | ( n2202 & n2420 ) ;
  assign n2388 = x10 & x31 ;
  assign n2389 = n1129 & n2388 ;
  assign n2390 = n360 & n1585 ;
  assign n2391 = n2389 | n2390 ;
  assign n2392 = x22 & x31 ;
  assign n2393 = n218 & n2392 ;
  assign n2394 = x21 & n2393 ;
  assign n2395 = ( x21 & ~n2391 ) | ( x21 & n2394 ) | ( ~n2391 & n2394 ) ;
  assign n2396 = x10 & n2395 ;
  assign n2397 = n2391 | n2393 ;
  assign n2398 = x0 & x31 ;
  assign n2399 = x9 & x22 ;
  assign n2400 = ( ~n2393 & n2398 ) | ( ~n2393 & n2399 ) | ( n2398 & n2399 ) ;
  assign n2401 = n2398 & n2399 ;
  assign n2402 = ( ~n2391 & n2400 ) | ( ~n2391 & n2401 ) | ( n2400 & n2401 ) ;
  assign n2403 = ~n2397 & n2402 ;
  assign n2404 = n2396 | n2403 ;
  assign n2405 = n720 & n1285 ;
  assign n2406 = n490 & n1437 ;
  assign n2407 = n2405 | n2406 ;
  assign n2408 = n647 & n1077 ;
  assign n2409 = x20 & n2408 ;
  assign n2410 = ( x20 & ~n2407 ) | ( x20 & n2409 ) | ( ~n2407 & n2409 ) ;
  assign n2411 = x11 & n2410 ;
  assign n2412 = n2407 | n2408 ;
  assign n2413 = x12 & x19 ;
  assign n2414 = x13 & x18 ;
  assign n2415 = ( ~n2408 & n2413 ) | ( ~n2408 & n2414 ) | ( n2413 & n2414 ) ;
  assign n2416 = n2413 & n2414 ;
  assign n2417 = ( ~n2407 & n2415 ) | ( ~n2407 & n2416 ) | ( n2415 & n2416 ) ;
  assign n2418 = ~n2412 & n2417 ;
  assign n2419 = n2411 | n2418 ;
  assign n2422 = ( n2404 & ~n2419 ) | ( n2404 & n2421 ) | ( ~n2419 & n2421 ) ;
  assign n2423 = ( ~n2404 & n2419 ) | ( ~n2404 & n2422 ) | ( n2419 & n2422 ) ;
  assign n2424 = ( ~n2421 & n2422 ) | ( ~n2421 & n2423 ) | ( n2422 & n2423 ) ;
  assign n2425 = n2387 & n2424 ;
  assign n2426 = n2387 | n2424 ;
  assign n2427 = ~n2425 & n2426 ;
  assign n2428 = ( n2139 & n2244 ) | ( n2139 & n2257 ) | ( n2244 & n2257 ) ;
  assign n2429 = n2244 | n2257 ;
  assign n2430 = ( n2160 & n2428 ) | ( n2160 & n2429 ) | ( n2428 & n2429 ) ;
  assign n2431 = n2427 | n2430 ;
  assign n2432 = n2427 & n2430 ;
  assign n2433 = n2431 & ~n2432 ;
  assign n2434 = n2223 | n2260 ;
  assign n2435 = ( n2223 & n2224 ) | ( n2223 & n2434 ) | ( n2224 & n2434 ) ;
  assign n2436 = n2433 & n2435 ;
  assign n2437 = n2433 | n2435 ;
  assign n2438 = ~n2436 & n2437 ;
  assign n2439 = n2228 | n2241 ;
  assign n2440 = n2079 | n2253 ;
  assign n2441 = ( n2253 & n2254 ) | ( n2253 & n2440 ) | ( n2254 & n2440 ) ;
  assign n2442 = n2439 | n2441 ;
  assign n2443 = n2439 & n2441 ;
  assign n2444 = n2442 & ~n2443 ;
  assign n2445 = x1 & x30 ;
  assign n2446 = x16 & n2445 ;
  assign n2447 = x16 | n2445 ;
  assign n2448 = ~n2446 & n2447 ;
  assign n2449 = n2204 & n2448 ;
  assign n2450 = n2204 | n2448 ;
  assign n2451 = ~n2449 & n2450 ;
  assign n2452 = n2284 & n2451 ;
  assign n2453 = n2284 | n2451 ;
  assign n2454 = ~n2452 & n2453 ;
  assign n2455 = n2444 & n2454 ;
  assign n2456 = n2444 | n2454 ;
  assign n2457 = ~n2455 & n2456 ;
  assign n2458 = n2316 & n2457 ;
  assign n2459 = ( n2323 & n2457 ) | ( n2323 & n2458 ) | ( n2457 & n2458 ) ;
  assign n2460 = n2316 | n2457 ;
  assign n2461 = n2323 | n2460 ;
  assign n2462 = ~n2459 & n2461 ;
  assign n2463 = n2234 | n2266 ;
  assign n2464 = n2271 | n2463 ;
  assign n2465 = n2234 & n2266 ;
  assign n2466 = ( n2234 & n2271 ) | ( n2234 & n2465 ) | ( n2271 & n2465 ) ;
  assign n2467 = n2464 & ~n2466 ;
  assign n2468 = n2303 | n2467 ;
  assign n2469 = n2303 & n2467 ;
  assign n2470 = n2468 & ~n2469 ;
  assign n2471 = n2292 | n2310 ;
  assign n2472 = n2470 & n2471 ;
  assign n2473 = n2292 & n2470 ;
  assign n2474 = ( n2295 & n2472 ) | ( n2295 & n2473 ) | ( n2472 & n2473 ) ;
  assign n2475 = n2470 | n2471 ;
  assign n2476 = n2292 | n2470 ;
  assign n2477 = ( n2295 & n2475 ) | ( n2295 & n2476 ) | ( n2475 & n2476 ) ;
  assign n2478 = ~n2474 & n2477 ;
  assign n2479 = n2214 | n2216 ;
  assign n2480 = ( n2214 & n2215 ) | ( n2214 & n2479 ) | ( n2215 & n2479 ) ;
  assign n2481 = n2478 | n2480 ;
  assign n2482 = n2478 & n2480 ;
  assign n2483 = n2481 & ~n2482 ;
  assign n2484 = n2462 & n2483 ;
  assign n2485 = n2462 | n2483 ;
  assign n2486 = ~n2484 & n2485 ;
  assign n2487 = n2438 & n2486 ;
  assign n2488 = n2438 | n2486 ;
  assign n2489 = ~n2487 & n2488 ;
  assign n2499 = n2263 | n2327 ;
  assign n2500 = ( n2327 & n2329 ) | ( n2327 & n2499 ) | ( n2329 & n2499 ) ;
  assign n2501 = ( n2489 & n2498 ) | ( n2489 & ~n2500 ) | ( n2498 & ~n2500 ) ;
  assign n2502 = ( ~n2489 & n2500 ) | ( ~n2489 & n2501 ) | ( n2500 & n2501 ) ;
  assign n2503 = ( ~n2498 & n2501 ) | ( ~n2498 & n2502 ) | ( n2501 & n2502 ) ;
  assign n2504 = n2489 & n2500 ;
  assign n2505 = n2489 | n2500 ;
  assign n2506 = n2504 | n2505 ;
  assign n2507 = ( n2498 & n2504 ) | ( n2498 & n2506 ) | ( n2504 & n2506 ) ;
  assign n2508 = n181 & n2340 ;
  assign n2509 = n251 & n1912 ;
  assign n2510 = n2508 | n2509 ;
  assign n2511 = x25 & x26 ;
  assign n2512 = n200 & n2511 ;
  assign n2513 = x24 & n2512 ;
  assign n2514 = ( x24 & ~n2510 ) | ( x24 & n2513 ) | ( ~n2510 & n2513 ) ;
  assign n2515 = x8 & n2514 ;
  assign n2516 = n2510 | n2512 ;
  assign n2517 = x6 & x26 ;
  assign n2518 = x7 & x25 ;
  assign n2519 = ( ~n2512 & n2517 ) | ( ~n2512 & n2518 ) | ( n2517 & n2518 ) ;
  assign n2520 = n2517 & n2518 ;
  assign n2521 = ( ~n2510 & n2519 ) | ( ~n2510 & n2520 ) | ( n2519 & n2520 ) ;
  assign n2522 = ~n2516 & n2521 ;
  assign n2523 = n2515 | n2522 ;
  assign n2524 = x5 & x27 ;
  assign n2525 = x4 & x28 ;
  assign n2526 = n2524 | n2525 ;
  assign n2527 = n91 & n2372 ;
  assign n2528 = n2526 | n2527 ;
  assign n2529 = x9 & x23 ;
  assign n2530 = ( ~n2527 & n2528 ) | ( ~n2527 & n2529 ) | ( n2528 & n2529 ) ;
  assign n2531 = ( n2527 & n2528 ) | ( n2527 & ~n2529 ) | ( n2528 & ~n2529 ) ;
  assign n2532 = ( ~n2528 & n2530 ) | ( ~n2528 & n2531 ) | ( n2530 & n2531 ) ;
  assign n2533 = n2523 & n2532 ;
  assign n2534 = n2523 & ~n2533 ;
  assign n2535 = ~n2523 & n2532 ;
  assign n2536 = n2284 | n2449 ;
  assign n2537 = ( n2449 & n2451 ) | ( n2449 & n2536 ) | ( n2451 & n2536 ) ;
  assign n2538 = n2535 | n2537 ;
  assign n2539 = n2534 | n2538 ;
  assign n2540 = n2535 & n2537 ;
  assign n2541 = ( n2534 & n2537 ) | ( n2534 & n2540 ) | ( n2537 & n2540 ) ;
  assign n2542 = n2539 & ~n2541 ;
  assign n2543 = x0 & x32 ;
  assign n2544 = x2 & x30 ;
  assign n2545 = n2543 | n2544 ;
  assign n2546 = x30 & x32 ;
  assign n2547 = n67 & n2546 ;
  assign n2548 = n2545 & ~n2547 ;
  assign n2549 = n2446 | n2547 ;
  assign n2550 = ( n2547 & n2548 ) | ( n2547 & n2549 ) | ( n2548 & n2549 ) ;
  assign n2551 = n2545 & ~n2550 ;
  assign n2552 = n2446 & ~n2548 ;
  assign n2553 = n2551 | n2552 ;
  assign n2554 = n720 & n1432 ;
  assign n2555 = n490 & n1434 ;
  assign n2556 = n2554 | n2555 ;
  assign n2557 = n647 & n1437 ;
  assign n2558 = x21 & n2557 ;
  assign n2559 = ( x21 & ~n2556 ) | ( x21 & n2558 ) | ( ~n2556 & n2558 ) ;
  assign n2560 = x11 & n2559 ;
  assign n2561 = n2556 | n2557 ;
  assign n2562 = x12 & x20 ;
  assign n2563 = x13 & x19 ;
  assign n2564 = ( ~n2557 & n2562 ) | ( ~n2557 & n2563 ) | ( n2562 & n2563 ) ;
  assign n2565 = n2562 & n2563 ;
  assign n2566 = ( ~n2556 & n2564 ) | ( ~n2556 & n2565 ) | ( n2564 & n2565 ) ;
  assign n2567 = ~n2561 & n2566 ;
  assign n2568 = n2560 | n2567 ;
  assign n2569 = n2553 & n2568 ;
  assign n2570 = n2553 & ~n2569 ;
  assign n2571 = n2568 & ~n2569 ;
  assign n2572 = n2570 | n2571 ;
  assign n2573 = x3 & x29 ;
  assign n2574 = x10 & x22 ;
  assign n2575 = n2573 | n2574 ;
  assign n2576 = x14 & x18 ;
  assign n2577 = ( n2573 & n2574 ) | ( n2573 & n2576 ) | ( n2574 & n2576 ) ;
  assign n2578 = n2575 & ~n2577 ;
  assign n2579 = n2573 & n2574 ;
  assign n2580 = n2576 & ~n2579 ;
  assign n2581 = ~n2575 & n2576 ;
  assign n2582 = ( n2576 & ~n2580 ) | ( n2576 & n2581 ) | ( ~n2580 & n2581 ) ;
  assign n2583 = n2578 | n2582 ;
  assign n2584 = ~n2572 & n2583 ;
  assign n2585 = n2572 & ~n2583 ;
  assign n2586 = n2584 | n2585 ;
  assign n2587 = n2542 | n2586 ;
  assign n2588 = n2542 & n2586 ;
  assign n2589 = n2587 & ~n2588 ;
  assign n2590 = n2474 | n2480 ;
  assign n2591 = ( n2474 & n2478 ) | ( n2474 & n2590 ) | ( n2478 & n2590 ) ;
  assign n2592 = n2589 & n2591 ;
  assign n2593 = n2589 | n2591 ;
  assign n2594 = ~n2592 & n2593 ;
  assign n2595 = n2458 | n2483 ;
  assign n2596 = n2457 | n2483 ;
  assign n2597 = ( n2323 & n2595 ) | ( n2323 & n2596 ) | ( n2595 & n2596 ) ;
  assign n2598 = n2594 & n2597 ;
  assign n2599 = n2459 & n2594 ;
  assign n2600 = ( n2462 & n2598 ) | ( n2462 & n2599 ) | ( n2598 & n2599 ) ;
  assign n2601 = n2594 | n2597 ;
  assign n2602 = n2459 | n2594 ;
  assign n2603 = ( n2462 & n2601 ) | ( n2462 & n2602 ) | ( n2601 & n2602 ) ;
  assign n2604 = ~n2600 & n2603 ;
  assign n2605 = n2397 | n2412 ;
  assign n2606 = n2397 & n2412 ;
  assign n2607 = n2605 & ~n2606 ;
  assign n2608 = n2377 | n2607 ;
  assign n2609 = n2377 & n2607 ;
  assign n2610 = n2608 & ~n2609 ;
  assign n2611 = x1 & x31 ;
  assign n2612 = n913 | n2611 ;
  assign n2613 = n913 & n2611 ;
  assign n2614 = n2612 & ~n2613 ;
  assign n2615 = n2359 | n2614 ;
  assign n2616 = n2359 & n2614 ;
  assign n2617 = n2615 & ~n2616 ;
  assign n2618 = n2345 & n2617 ;
  assign n2619 = n2345 | n2617 ;
  assign n2620 = ~n2618 & n2619 ;
  assign n2621 = n2610 & n2620 ;
  assign n2622 = n2610 | n2620 ;
  assign n2623 = ~n2621 & n2622 ;
  assign n2624 = ( n2439 & n2441 ) | ( n2439 & n2454 ) | ( n2441 & n2454 ) ;
  assign n2625 = n2623 | n2624 ;
  assign n2626 = n2623 & n2624 ;
  assign n2627 = n2625 & ~n2626 ;
  assign n2628 = n2419 & n2421 ;
  assign n2629 = n2421 & ~n2628 ;
  assign n2630 = n2419 & ~n2628 ;
  assign n2631 = n2629 | n2630 ;
  assign n2632 = n2303 | n2466 ;
  assign n2633 = ( n2466 & n2467 ) | ( n2466 & n2632 ) | ( n2467 & n2632 ) ;
  assign n2634 = n2628 & n2633 ;
  assign n2635 = n2404 & n2633 ;
  assign n2636 = ( n2628 & n2633 ) | ( n2628 & n2635 ) | ( n2633 & n2635 ) ;
  assign n2637 = ( n2631 & n2634 ) | ( n2631 & n2636 ) | ( n2634 & n2636 ) ;
  assign n2638 = n2628 | n2633 ;
  assign n2639 = n2404 | n2633 ;
  assign n2640 = n2628 | n2639 ;
  assign n2641 = ( n2631 & n2638 ) | ( n2631 & n2640 ) | ( n2638 & n2640 ) ;
  assign n2642 = ~n2637 & n2641 ;
  assign n2643 = n2364 | n2384 ;
  assign n2644 = ( n2364 & n2367 ) | ( n2364 & n2643 ) | ( n2367 & n2643 ) ;
  assign n2645 = n2642 | n2644 ;
  assign n2646 = n2642 & n2644 ;
  assign n2647 = n2645 & ~n2646 ;
  assign n2648 = n2424 | n2430 ;
  assign n2649 = ( n2387 & n2430 ) | ( n2387 & n2648 ) | ( n2430 & n2648 ) ;
  assign n2650 = ( n2425 & n2427 ) | ( n2425 & n2649 ) | ( n2427 & n2649 ) ;
  assign n2651 = n2647 | n2650 ;
  assign n2652 = n2647 & n2650 ;
  assign n2653 = n2651 & ~n2652 ;
  assign n2654 = n2627 & n2653 ;
  assign n2655 = n2627 | n2653 ;
  assign n2656 = ~n2654 & n2655 ;
  assign n2657 = n2604 & n2656 ;
  assign n2658 = n2604 | n2656 ;
  assign n2659 = ~n2657 & n2658 ;
  assign n2660 = n2436 | n2487 ;
  assign n2661 = ( n2507 & n2659 ) | ( n2507 & ~n2660 ) | ( n2659 & ~n2660 ) ;
  assign n2662 = ( ~n2659 & n2660 ) | ( ~n2659 & n2661 ) | ( n2660 & n2661 ) ;
  assign n2663 = ( ~n2507 & n2661 ) | ( ~n2507 & n2662 ) | ( n2661 & n2662 ) ;
  assign n2664 = n2659 & n2660 ;
  assign n2665 = n2659 | n2660 ;
  assign n2666 = n2504 & n2665 ;
  assign n2667 = n2664 | n2666 ;
  assign n2668 = n2664 | n2665 ;
  assign n2669 = ( n2506 & n2664 ) | ( n2506 & n2668 ) | ( n2664 & n2668 ) ;
  assign n2670 = ( n2498 & n2667 ) | ( n2498 & n2669 ) | ( n2667 & n2669 ) ;
  assign n2671 = n2550 | n2561 ;
  assign n2672 = n2550 & n2561 ;
  assign n2673 = n2671 & ~n2672 ;
  assign n2674 = n2577 | n2673 ;
  assign n2675 = n2577 & n2673 ;
  assign n2676 = n2674 & ~n2675 ;
  assign n2677 = ~n2527 & n2529 ;
  assign n2678 = ( n2527 & n2528 ) | ( n2527 & n2677 ) | ( n2528 & n2677 ) ;
  assign n2679 = n2516 | n2678 ;
  assign n2680 = n2516 & n2678 ;
  assign n2681 = n2679 & ~n2680 ;
  assign n2682 = n432 & n2392 ;
  assign n2683 = x31 & x33 ;
  assign n2684 = n67 & n2683 ;
  assign n2685 = n2682 | n2684 ;
  assign n2686 = x22 & x33 ;
  assign n2687 = n329 & n2686 ;
  assign n2688 = x31 & n2687 ;
  assign n2689 = ( x31 & ~n2685 ) | ( x31 & n2688 ) | ( ~n2685 & n2688 ) ;
  assign n2690 = x2 & n2689 ;
  assign n2691 = n2685 | n2687 ;
  assign n2692 = x0 & x33 ;
  assign n2693 = x11 & x22 ;
  assign n2694 = ( ~n2687 & n2692 ) | ( ~n2687 & n2693 ) | ( n2692 & n2693 ) ;
  assign n2695 = n2692 & n2693 ;
  assign n2696 = ( ~n2685 & n2694 ) | ( ~n2685 & n2695 ) | ( n2694 & n2695 ) ;
  assign n2697 = ~n2691 & n2696 ;
  assign n2698 = n2690 | n2697 ;
  assign n2699 = n2681 & n2698 ;
  assign n2700 = n2681 & ~n2699 ;
  assign n2701 = n2698 & ~n2699 ;
  assign n2702 = n2700 | n2701 ;
  assign n2703 = n2676 | n2702 ;
  assign n2704 = n2676 & n2702 ;
  assign n2705 = n2703 & ~n2704 ;
  assign n2706 = x4 & x29 ;
  assign n2707 = x9 & x24 ;
  assign n2708 = n2706 & n2707 ;
  assign n2709 = x29 & x30 ;
  assign n2710 = n79 & n2709 ;
  assign n2711 = x24 & x30 ;
  assign n2712 = n357 & n2711 ;
  assign n2713 = n2710 | n2712 ;
  assign n2714 = x30 & n2708 ;
  assign n2715 = ( x30 & ~n2713 ) | ( x30 & n2714 ) | ( ~n2713 & n2714 ) ;
  assign n2716 = x3 & n2715 ;
  assign n2717 = ( n2706 & n2707 ) | ( n2706 & ~n2713 ) | ( n2707 & ~n2713 ) ;
  assign n2718 = ( ~n2708 & n2716 ) | ( ~n2708 & n2717 ) | ( n2716 & n2717 ) ;
  assign n2719 = x5 & x28 ;
  assign n2720 = n204 & n2372 ;
  assign n2721 = x8 & x25 ;
  assign n2722 = n2719 & n2721 ;
  assign n2723 = n2720 | n2722 ;
  assign n2724 = x25 & x27 ;
  assign n2725 = n181 & n2724 ;
  assign n2726 = n2719 & n2725 ;
  assign n2727 = ( n2719 & ~n2723 ) | ( n2719 & n2726 ) | ( ~n2723 & n2726 ) ;
  assign n2728 = n2723 | n2725 ;
  assign n2729 = x6 & x27 ;
  assign n2730 = ( n2721 & ~n2725 ) | ( n2721 & n2729 ) | ( ~n2725 & n2729 ) ;
  assign n2731 = n2721 & n2729 ;
  assign n2732 = ( ~n2723 & n2730 ) | ( ~n2723 & n2731 ) | ( n2730 & n2731 ) ;
  assign n2733 = ~n2728 & n2732 ;
  assign n2734 = n2727 | n2733 ;
  assign n2735 = n2718 & n2734 ;
  assign n2736 = n2718 & ~n2735 ;
  assign n2737 = x15 & x18 ;
  assign n2738 = n1023 | n2737 ;
  assign n2739 = n795 & n1020 ;
  assign n2740 = x7 & x26 ;
  assign n2741 = ~n2739 & n2740 ;
  assign n2742 = n2738 | n2739 ;
  assign n2743 = ( n2739 & n2741 ) | ( n2739 & n2742 ) | ( n2741 & n2742 ) ;
  assign n2744 = n2738 & ~n2743 ;
  assign n2745 = ( ~n2738 & n2739 ) | ( ~n2738 & n2740 ) | ( n2739 & n2740 ) ;
  assign n2746 = n2740 & n2745 ;
  assign n2747 = n2744 | n2746 ;
  assign n2748 = ~n2718 & n2734 ;
  assign n2749 = n2747 & n2748 ;
  assign n2750 = ( n2736 & n2747 ) | ( n2736 & n2749 ) | ( n2747 & n2749 ) ;
  assign n2751 = n2747 | n2748 ;
  assign n2752 = n2736 | n2751 ;
  assign n2753 = ~n2750 & n2752 ;
  assign n2754 = n2705 & ~n2753 ;
  assign n2755 = ~n2705 & n2753 ;
  assign n2756 = n2754 | n2755 ;
  assign n2757 = n2569 | n2583 ;
  assign n2758 = n2377 | n2606 ;
  assign n2759 = ( n2606 & n2607 ) | ( n2606 & n2758 ) | ( n2607 & n2758 ) ;
  assign n2760 = n2757 & n2759 ;
  assign n2761 = n2569 & n2759 ;
  assign n2762 = ( n2572 & n2760 ) | ( n2572 & n2761 ) | ( n2760 & n2761 ) ;
  assign n2763 = n2757 | n2759 ;
  assign n2764 = n2569 | n2759 ;
  assign n2765 = ( n2572 & n2763 ) | ( n2572 & n2764 ) | ( n2763 & n2764 ) ;
  assign n2766 = ~n2762 & n2765 ;
  assign n2767 = n2533 | n2541 ;
  assign n2768 = n2766 | n2767 ;
  assign n2769 = n2766 & n2767 ;
  assign n2770 = n2768 & ~n2769 ;
  assign n2771 = n2588 | n2591 ;
  assign n2772 = ( n2588 & n2589 ) | ( n2588 & n2771 ) | ( n2589 & n2771 ) ;
  assign n2773 = n2770 & n2772 ;
  assign n2774 = n2770 | n2772 ;
  assign n2775 = ~n2773 & n2774 ;
  assign n2776 = n2756 & n2775 ;
  assign n2777 = n2756 | n2775 ;
  assign n2778 = ~n2776 & n2777 ;
  assign n2779 = x1 & x32 ;
  assign n2780 = x17 & n2779 ;
  assign n2781 = x17 & ~n2779 ;
  assign n2782 = ( n2779 & ~n2780 ) | ( n2779 & n2781 ) | ( ~n2780 & n2781 ) ;
  assign n2783 = x10 & x23 ;
  assign n2784 = n2613 & n2783 ;
  assign n2785 = n2782 & ~n2784 ;
  assign n2786 = n2613 | n2783 ;
  assign n2787 = n2782 & ~n2786 ;
  assign n2788 = ( n2782 & ~n2785 ) | ( n2782 & n2787 ) | ( ~n2785 & n2787 ) ;
  assign n2789 = ~n2613 & n2786 ;
  assign n2790 = n2613 & ~n2783 ;
  assign n2791 = ( ~n2785 & n2789 ) | ( ~n2785 & n2790 ) | ( n2789 & n2790 ) ;
  assign n2792 = n2788 | n2791 ;
  assign n2793 = n487 & n1432 ;
  assign n2794 = n647 & n1434 ;
  assign n2795 = n2793 | n2794 ;
  assign n2796 = n650 & n1437 ;
  assign n2797 = x21 & n2796 ;
  assign n2798 = ( x21 & ~n2795 ) | ( x21 & n2797 ) | ( ~n2795 & n2797 ) ;
  assign n2799 = x12 & n2798 ;
  assign n2800 = n2795 | n2796 ;
  assign n2801 = x13 & x20 ;
  assign n2802 = x14 & x19 ;
  assign n2803 = ( ~n2796 & n2801 ) | ( ~n2796 & n2802 ) | ( n2801 & n2802 ) ;
  assign n2804 = n2801 & n2802 ;
  assign n2805 = ( ~n2795 & n2803 ) | ( ~n2795 & n2804 ) | ( n2803 & n2804 ) ;
  assign n2806 = ~n2800 & n2805 ;
  assign n2807 = n2799 | n2806 ;
  assign n2808 = n2792 & n2807 ;
  assign n2809 = n2792 & ~n2808 ;
  assign n2811 = n2345 | n2616 ;
  assign n2812 = ( n2616 & n2617 ) | ( n2616 & n2811 ) | ( n2617 & n2811 ) ;
  assign n2810 = ~n2792 & n2807 ;
  assign n2813 = n2810 & n2812 ;
  assign n2814 = ( n2809 & n2812 ) | ( n2809 & n2813 ) | ( n2812 & n2813 ) ;
  assign n2815 = n2810 | n2812 ;
  assign n2816 = n2809 | n2815 ;
  assign n2817 = ~n2814 & n2816 ;
  assign n2818 = n2637 | n2644 ;
  assign n2819 = ( n2637 & n2642 ) | ( n2637 & n2818 ) | ( n2642 & n2818 ) ;
  assign n2820 = n2817 | n2819 ;
  assign n2821 = n2817 & n2819 ;
  assign n2822 = n2820 & ~n2821 ;
  assign n2823 = n2621 | n2624 ;
  assign n2824 = ( n2621 & n2623 ) | ( n2621 & n2823 ) | ( n2623 & n2823 ) ;
  assign n2825 = n2822 | n2824 ;
  assign n2826 = n2822 & n2824 ;
  assign n2827 = n2825 & ~n2826 ;
  assign n2828 = n2627 | n2647 ;
  assign n2829 = ( n2627 & n2650 ) | ( n2627 & n2828 ) | ( n2650 & n2828 ) ;
  assign n2830 = ( n2652 & n2653 ) | ( n2652 & n2829 ) | ( n2653 & n2829 ) ;
  assign n2831 = n2827 & n2830 ;
  assign n2832 = n2827 | n2830 ;
  assign n2833 = ~n2831 & n2832 ;
  assign n2834 = n2778 & n2833 ;
  assign n2835 = n2778 | n2833 ;
  assign n2836 = ~n2834 & n2835 ;
  assign n2837 = n2600 | n2657 ;
  assign n2838 = ( n2670 & n2836 ) | ( n2670 & ~n2837 ) | ( n2836 & ~n2837 ) ;
  assign n2839 = ( ~n2836 & n2837 ) | ( ~n2836 & n2838 ) | ( n2837 & n2838 ) ;
  assign n2840 = ( ~n2670 & n2838 ) | ( ~n2670 & n2839 ) | ( n2838 & n2839 ) ;
  assign n2841 = ( n2613 & n2783 ) | ( n2613 & n2785 ) | ( n2783 & n2785 ) ;
  assign n2842 = n2800 | n2841 ;
  assign n2843 = n2800 & n2841 ;
  assign n2844 = n2842 & ~n2843 ;
  assign n2845 = x11 & x23 ;
  assign n2846 = x12 & x22 ;
  assign n2847 = n2845 | n2846 ;
  assign n2848 = n490 & n1932 ;
  assign n2849 = x2 & x32 ;
  assign n2850 = ~n2848 & n2849 ;
  assign n2851 = n2847 | n2848 ;
  assign n2852 = ( n2848 & n2850 ) | ( n2848 & n2851 ) | ( n2850 & n2851 ) ;
  assign n2853 = n2847 & ~n2852 ;
  assign n2854 = ( ~n2847 & n2848 ) | ( ~n2847 & n2849 ) | ( n2848 & n2849 ) ;
  assign n2855 = n2849 & n2854 ;
  assign n2856 = n2853 | n2855 ;
  assign n2857 = ~n2844 & n2856 ;
  assign n2858 = n2844 & ~n2856 ;
  assign n2859 = n2857 | n2858 ;
  assign n2860 = n2808 | n2814 ;
  assign n2861 = n2859 | n2860 ;
  assign n2862 = n2859 & n2860 ;
  assign n2863 = n2861 & ~n2862 ;
  assign n2864 = x5 & x29 ;
  assign n2865 = x9 & x25 ;
  assign n2866 = n2864 & n2865 ;
  assign n2867 = n360 & n1912 ;
  assign n2868 = x24 & x29 ;
  assign n2869 = n581 & n2868 ;
  assign n2870 = n2867 | n2869 ;
  assign n2871 = x24 & n2866 ;
  assign n2872 = ( x24 & ~n2870 ) | ( x24 & n2871 ) | ( ~n2870 & n2871 ) ;
  assign n2873 = x10 & n2872 ;
  assign n2874 = ( n2864 & n2865 ) | ( n2864 & ~n2870 ) | ( n2865 & ~n2870 ) ;
  assign n2875 = ( ~n2866 & n2873 ) | ( ~n2866 & n2874 ) | ( n2873 & n2874 ) ;
  assign n2876 = n723 & n1432 ;
  assign n2877 = n650 & n1434 ;
  assign n2878 = n2876 | n2877 ;
  assign n2879 = n792 & n1437 ;
  assign n2880 = x21 & n2879 ;
  assign n2881 = ( x21 & ~n2878 ) | ( x21 & n2880 ) | ( ~n2878 & n2880 ) ;
  assign n2882 = x13 & n2881 ;
  assign n2883 = n2878 | n2879 ;
  assign n2884 = x14 & x20 ;
  assign n2885 = x15 & x19 ;
  assign n2886 = ( ~n2879 & n2884 ) | ( ~n2879 & n2885 ) | ( n2884 & n2885 ) ;
  assign n2887 = n2884 & n2885 ;
  assign n2888 = ( ~n2878 & n2886 ) | ( ~n2878 & n2887 ) | ( n2886 & n2887 ) ;
  assign n2889 = ~n2883 & n2888 ;
  assign n2890 = n2882 | n2889 ;
  assign n2891 = n2875 & n2890 ;
  assign n2892 = n2875 & ~n2891 ;
  assign n2893 = n2890 & ~n2891 ;
  assign n2894 = n2892 | n2893 ;
  assign n2895 = x26 & x28 ;
  assign n2896 = n181 & n2895 ;
  assign n2897 = n200 & n2372 ;
  assign n2898 = n2896 | n2897 ;
  assign n2899 = n251 & n2267 ;
  assign n2900 = x28 & n2899 ;
  assign n2901 = ( x28 & ~n2898 ) | ( x28 & n2900 ) | ( ~n2898 & n2900 ) ;
  assign n2902 = x6 & n2901 ;
  assign n2903 = n2898 | n2899 ;
  assign n2904 = x7 & x27 ;
  assign n2905 = x8 & x26 ;
  assign n2906 = ( ~n2899 & n2904 ) | ( ~n2899 & n2905 ) | ( n2904 & n2905 ) ;
  assign n2907 = n2904 & n2905 ;
  assign n2908 = ( ~n2898 & n2906 ) | ( ~n2898 & n2907 ) | ( n2906 & n2907 ) ;
  assign n2909 = ~n2903 & n2908 ;
  assign n2910 = n2902 | n2909 ;
  assign n2911 = ~n2894 & n2910 ;
  assign n2912 = n2894 & ~n2910 ;
  assign n2913 = n2911 | n2912 ;
  assign n2914 = n2863 & n2913 ;
  assign n2915 = n2863 | n2913 ;
  assign n2916 = n2708 | n2713 ;
  assign n2917 = n2691 | n2916 ;
  assign n2918 = n2691 & n2916 ;
  assign n2919 = n2917 & ~n2918 ;
  assign n2920 = n2728 | n2919 ;
  assign n2921 = n2728 & n2919 ;
  assign n2922 = n2920 & ~n2921 ;
  assign n2923 = x1 & x33 ;
  assign n2924 = n1018 & n2923 ;
  assign n2925 = n1018 | n2923 ;
  assign n2926 = ~n2924 & n2925 ;
  assign n2927 = n2780 & n2926 ;
  assign n2928 = n2780 | n2926 ;
  assign n2929 = ~n2927 & n2928 ;
  assign n2930 = n2743 & n2929 ;
  assign n2931 = n2743 | n2929 ;
  assign n2932 = ~n2930 & n2931 ;
  assign n2933 = n2735 & n2932 ;
  assign n2934 = ( n2750 & n2932 ) | ( n2750 & n2933 ) | ( n2932 & n2933 ) ;
  assign n2935 = n2735 | n2932 ;
  assign n2936 = n2750 | n2935 ;
  assign n2937 = ~n2934 & n2936 ;
  assign n2938 = n2922 & n2937 ;
  assign n2939 = n2922 | n2937 ;
  assign n2940 = ~n2938 & n2939 ;
  assign n2941 = n2915 & n2940 ;
  assign n2942 = n2914 & n2915 ;
  assign n2943 = ( n2915 & ~n2941 ) | ( n2915 & n2942 ) | ( ~n2941 & n2942 ) ;
  assign n2944 = ~n2914 & n2943 ;
  assign n2945 = n2817 | n2824 ;
  assign n2946 = ( n2819 & n2824 ) | ( n2819 & n2945 ) | ( n2824 & n2945 ) ;
  assign n2947 = ( n2821 & n2822 ) | ( n2821 & n2946 ) | ( n2822 & n2946 ) ;
  assign n2948 = n2914 & n2940 ;
  assign n2949 = ( n2940 & ~n2941 ) | ( n2940 & n2948 ) | ( ~n2941 & n2948 ) ;
  assign n2950 = n2947 & n2949 ;
  assign n2951 = ( n2944 & n2947 ) | ( n2944 & n2950 ) | ( n2947 & n2950 ) ;
  assign n2952 = n2947 | n2949 ;
  assign n2953 = n2944 | n2952 ;
  assign n2954 = ~n2951 & n2953 ;
  assign n2955 = ( n2676 & n2702 ) | ( n2676 & n2753 ) | ( n2702 & n2753 ) ;
  assign n2956 = n2762 | n2767 ;
  assign n2957 = ( n2762 & n2766 ) | ( n2762 & n2956 ) | ( n2766 & n2956 ) ;
  assign n2958 = n2955 | n2957 ;
  assign n2959 = n2955 & n2957 ;
  assign n2960 = n2958 & ~n2959 ;
  assign n2961 = n2680 | n2699 ;
  assign n2962 = x31 & n71 ;
  assign n2963 = x30 & n82 ;
  assign n2964 = n2962 | n2963 ;
  assign n2965 = x30 & x31 ;
  assign n2966 = n79 & n2965 ;
  assign n2967 = x34 & ~n2966 ;
  assign n2968 = n2964 & n2967 ;
  assign n2969 = x3 & x31 ;
  assign n2970 = x4 & x30 ;
  assign n2971 = n2969 | n2970 ;
  assign n2972 = ~n2966 & n2971 ;
  assign n2973 = x0 & x34 ;
  assign n2974 = n2972 | n2973 ;
  assign n2975 = ~n2968 & n2974 ;
  assign n2976 = n2577 | n2672 ;
  assign n2977 = ( n2672 & n2673 ) | ( n2672 & n2976 ) | ( n2673 & n2976 ) ;
  assign n2978 = n2975 & n2977 ;
  assign n2979 = n2975 | n2977 ;
  assign n2980 = ~n2978 & n2979 ;
  assign n2981 = n2961 & n2980 ;
  assign n2982 = n2961 | n2980 ;
  assign n2983 = ~n2981 & n2982 ;
  assign n2984 = n2960 & n2983 ;
  assign n2985 = n2960 | n2983 ;
  assign n2986 = ~n2984 & n2985 ;
  assign n2987 = ( n2756 & n2770 ) | ( n2756 & n2772 ) | ( n2770 & n2772 ) ;
  assign n2988 = n2986 | n2987 ;
  assign n2989 = n2986 & n2987 ;
  assign n2990 = n2988 & ~n2989 ;
  assign n2991 = n2954 & n2990 ;
  assign n2992 = n2954 | n2990 ;
  assign n2993 = ~n2991 & n2992 ;
  assign n2994 = n2836 & n2837 ;
  assign n2995 = n2836 | n2837 ;
  assign n2996 = n2669 & n2995 ;
  assign n2997 = n2667 & n2995 ;
  assign n2998 = ( n2498 & n2996 ) | ( n2498 & n2997 ) | ( n2996 & n2997 ) ;
  assign n2999 = n2994 | n2998 ;
  assign n3000 = n2778 | n2831 ;
  assign n3001 = ( n2831 & n2833 ) | ( n2831 & n3000 ) | ( n2833 & n3000 ) ;
  assign n3002 = ( n2993 & ~n2999 ) | ( n2993 & n3001 ) | ( ~n2999 & n3001 ) ;
  assign n3003 = ( n2999 & ~n3001 ) | ( n2999 & n3002 ) | ( ~n3001 & n3002 ) ;
  assign n3004 = ( ~n2993 & n3002 ) | ( ~n2993 & n3003 ) | ( n3002 & n3003 ) ;
  assign n3005 = n2993 & n3001 ;
  assign n3006 = n2993 | n3001 ;
  assign n3007 = n2994 & n3006 ;
  assign n3008 = ( n2998 & n3006 ) | ( n2998 & n3007 ) | ( n3006 & n3007 ) ;
  assign n3009 = n3005 | n3008 ;
  assign n3010 = n2728 | n2918 ;
  assign n3011 = ( n2918 & n2919 ) | ( n2918 & n3010 ) | ( n2919 & n3010 ) ;
  assign n3012 = n2743 | n2927 ;
  assign n3013 = ( n2927 & n2929 ) | ( n2927 & n3012 ) | ( n2929 & n3012 ) ;
  assign n3014 = n3011 | n3013 ;
  assign n3015 = n3011 & n3013 ;
  assign n3016 = n3014 & ~n3015 ;
  assign n3017 = n2843 | n2856 ;
  assign n3018 = ( n2843 & n2844 ) | ( n2843 & n3017 ) | ( n2844 & n3017 ) ;
  assign n3019 = n3016 | n3018 ;
  assign n3020 = n3016 & n3018 ;
  assign n3021 = n3019 & ~n3020 ;
  assign n3022 = n2922 | n2933 ;
  assign n3023 = n2922 | n2932 ;
  assign n3024 = ( n2750 & n3022 ) | ( n2750 & n3023 ) | ( n3022 & n3023 ) ;
  assign n3025 = ( n2934 & n2937 ) | ( n2934 & n3024 ) | ( n2937 & n3024 ) ;
  assign n3026 = n3021 | n3025 ;
  assign n3027 = n3021 & n3025 ;
  assign n3028 = n3026 & ~n3027 ;
  assign n3029 = n2862 | n2913 ;
  assign n3030 = ( n2862 & n2863 ) | ( n2862 & n3029 ) | ( n2863 & n3029 ) ;
  assign n3031 = n3028 & n3030 ;
  assign n3032 = n3028 | n3030 ;
  assign n3033 = ~n3031 & n3032 ;
  assign n3034 = ~n2914 & n2941 ;
  assign n3035 = n3033 & n3034 ;
  assign n3036 = ( n2951 & n3033 ) | ( n2951 & n3035 ) | ( n3033 & n3035 ) ;
  assign n3037 = n3033 | n3034 ;
  assign n3038 = n2951 | n3037 ;
  assign n3039 = ~n3036 & n3038 ;
  assign n3040 = n2852 | n2883 ;
  assign n3041 = n2852 & n2883 ;
  assign n3042 = n3040 & ~n3041 ;
  assign n3043 = n2966 | n2968 ;
  assign n3044 = n3042 | n3043 ;
  assign n3045 = n3042 & n3043 ;
  assign n3046 = n3044 & ~n3045 ;
  assign n3047 = x34 & n872 ;
  assign n3048 = x1 & x34 ;
  assign n3049 = x18 | n3048 ;
  assign n3050 = ~n3047 & n3049 ;
  assign n3051 = n2903 | n3050 ;
  assign n3052 = n2903 & n3050 ;
  assign n3053 = n3051 & ~n3052 ;
  assign n3054 = n2866 | n2870 ;
  assign n3055 = n3053 & n3054 ;
  assign n3056 = n3053 | n3054 ;
  assign n3057 = ~n3055 & n3056 ;
  assign n3058 = n2891 | n2910 ;
  assign n3059 = n3057 & n3058 ;
  assign n3060 = n2891 & n3057 ;
  assign n3061 = ( n2894 & n3059 ) | ( n2894 & n3060 ) | ( n3059 & n3060 ) ;
  assign n3062 = n3057 | n3058 ;
  assign n3063 = n2891 | n3057 ;
  assign n3064 = ( n2894 & n3062 ) | ( n2894 & n3063 ) | ( n3062 & n3063 ) ;
  assign n3065 = ~n3061 & n3064 ;
  assign n3066 = n3046 & n3065 ;
  assign n3067 = n3046 | n3065 ;
  assign n3068 = ~n3066 & n3067 ;
  assign n3069 = n2955 | n2983 ;
  assign n3070 = ( n2957 & n2983 ) | ( n2957 & n3069 ) | ( n2983 & n3069 ) ;
  assign n3071 = n3068 & n3070 ;
  assign n3072 = n2959 & n3068 ;
  assign n3073 = ( n2960 & n3071 ) | ( n2960 & n3072 ) | ( n3071 & n3072 ) ;
  assign n3074 = n3068 | n3070 ;
  assign n3075 = n2959 | n3068 ;
  assign n3076 = ( n2960 & n3074 ) | ( n2960 & n3075 ) | ( n3074 & n3075 ) ;
  assign n3077 = ~n3073 & n3076 ;
  assign n3078 = n2961 | n2978 ;
  assign n3079 = ( n2978 & n2980 ) | ( n2978 & n3078 ) | ( n2980 & n3078 ) ;
  assign n3080 = x27 & x30 ;
  assign n3081 = n222 & n3080 ;
  assign n3082 = n204 & n2709 ;
  assign n3083 = n3081 | n3082 ;
  assign n3084 = n181 & n2075 ;
  assign n3085 = x30 & n3084 ;
  assign n3086 = ( x30 & ~n3083 ) | ( x30 & n3085 ) | ( ~n3083 & n3085 ) ;
  assign n3087 = x5 & n3086 ;
  assign n3088 = n3083 | n3084 ;
  assign n3089 = x6 & x29 ;
  assign n3090 = ( n2269 & ~n3084 ) | ( n2269 & n3089 ) | ( ~n3084 & n3089 ) ;
  assign n3091 = n2269 & n3089 ;
  assign n3092 = ( ~n3083 & n3090 ) | ( ~n3083 & n3091 ) | ( n3090 & n3091 ) ;
  assign n3093 = ~n3088 & n3092 ;
  assign n3094 = n3087 | n3093 ;
  assign n3095 = x16 & x19 ;
  assign n3096 = n1020 | n3095 ;
  assign n3097 = x7 & x28 ;
  assign n3098 = ( n1020 & n3095 ) | ( n1020 & n3097 ) | ( n3095 & n3097 ) ;
  assign n3099 = n3096 & ~n3098 ;
  assign n3100 = n1020 & n3095 ;
  assign n3101 = n3097 & ~n3100 ;
  assign n3102 = ~n3096 & n3097 ;
  assign n3103 = ( n3097 & ~n3101 ) | ( n3097 & n3102 ) | ( ~n3101 & n3102 ) ;
  assign n3104 = n3099 | n3103 ;
  assign n3105 = n3094 & n3104 ;
  assign n3106 = n3094 & ~n3105 ;
  assign n3107 = x9 & x26 ;
  assign n3108 = x10 & x25 ;
  assign n3109 = n3107 | n3108 ;
  assign n3110 = n360 & n2511 ;
  assign n3111 = x4 & x31 ;
  assign n3112 = ~n3110 & n3111 ;
  assign n3113 = n3109 | n3110 ;
  assign n3114 = ( n3110 & n3112 ) | ( n3110 & n3113 ) | ( n3112 & n3113 ) ;
  assign n3115 = n3109 & ~n3114 ;
  assign n3116 = ( ~n3109 & n3110 ) | ( ~n3109 & n3111 ) | ( n3110 & n3111 ) ;
  assign n3117 = n3111 & n3116 ;
  assign n3118 = n3115 | n3117 ;
  assign n3119 = ~n3094 & n3104 ;
  assign n3120 = n3118 & ~n3119 ;
  assign n3121 = ~n3106 & n3120 ;
  assign n3122 = n3079 & n3121 ;
  assign n3123 = ~n3118 & n3119 ;
  assign n3124 = ( n3106 & ~n3118 ) | ( n3106 & n3123 ) | ( ~n3118 & n3123 ) ;
  assign n3125 = ( n3079 & n3122 ) | ( n3079 & n3124 ) | ( n3122 & n3124 ) ;
  assign n3126 = x0 & x35 ;
  assign n3127 = x2 & x33 ;
  assign n3128 = n3126 | n3127 ;
  assign n3129 = x33 & x35 ;
  assign n3130 = n67 & n3129 ;
  assign n3131 = n3128 & ~n3130 ;
  assign n3132 = n2924 | n3130 ;
  assign n3133 = ( n3130 & n3131 ) | ( n3130 & n3132 ) | ( n3131 & n3132 ) ;
  assign n3134 = n3128 & ~n3133 ;
  assign n3135 = n2924 & ~n3131 ;
  assign n3136 = n3134 | n3135 ;
  assign n3137 = x11 & x24 ;
  assign n3138 = x12 & x23 ;
  assign n3139 = n3137 | n3138 ;
  assign n3140 = n490 & n1686 ;
  assign n3141 = x3 & x32 ;
  assign n3142 = ~n3140 & n3141 ;
  assign n3143 = n3139 | n3140 ;
  assign n3144 = ( n3140 & n3142 ) | ( n3140 & n3143 ) | ( n3142 & n3143 ) ;
  assign n3145 = n3139 & ~n3144 ;
  assign n3146 = ~n3139 & n3141 ;
  assign n3147 = ( n3141 & ~n3142 ) | ( n3141 & n3146 ) | ( ~n3142 & n3146 ) ;
  assign n3148 = n3145 | n3147 ;
  assign n3149 = n3136 & n3148 ;
  assign n3150 = n3136 & ~n3149 ;
  assign n3151 = n3148 & ~n3149 ;
  assign n3152 = n3150 | n3151 ;
  assign n3153 = n723 & n1710 ;
  assign n3154 = n650 & n1585 ;
  assign n3155 = n3153 | n3154 ;
  assign n3156 = n792 & n1434 ;
  assign n3157 = x22 & n3156 ;
  assign n3158 = ( x22 & ~n3155 ) | ( x22 & n3157 ) | ( ~n3155 & n3157 ) ;
  assign n3159 = x13 & n3158 ;
  assign n3160 = n3155 | n3156 ;
  assign n3161 = x14 & x21 ;
  assign n3162 = x15 & x20 ;
  assign n3163 = ( ~n3156 & n3161 ) | ( ~n3156 & n3162 ) | ( n3161 & n3162 ) ;
  assign n3164 = n3161 & n3162 ;
  assign n3165 = ( ~n3155 & n3163 ) | ( ~n3155 & n3164 ) | ( n3163 & n3164 ) ;
  assign n3166 = ~n3160 & n3165 ;
  assign n3167 = n3159 | n3166 ;
  assign n3168 = ~n3152 & n3167 ;
  assign n3169 = n3152 & ~n3167 ;
  assign n3170 = n3168 | n3169 ;
  assign n3171 = n3121 | n3124 ;
  assign n3172 = n3079 | n3171 ;
  assign n3173 = n3170 & n3172 ;
  assign n3174 = ~n3125 & n3173 ;
  assign n3175 = n3170 | n3172 ;
  assign n3176 = ( ~n3125 & n3170 ) | ( ~n3125 & n3175 ) | ( n3170 & n3175 ) ;
  assign n3177 = ~n3174 & n3176 ;
  assign n3178 = ~n3077 & n3177 ;
  assign n3179 = n3077 & ~n3177 ;
  assign n3180 = n3178 | n3179 ;
  assign n3181 = n3039 | n3180 ;
  assign n3182 = n3039 & n3180 ;
  assign n3183 = n3181 & ~n3182 ;
  assign n3184 = n2989 | n2991 ;
  assign n3185 = ( n3009 & n3183 ) | ( n3009 & ~n3184 ) | ( n3183 & ~n3184 ) ;
  assign n3186 = ( ~n3183 & n3184 ) | ( ~n3183 & n3185 ) | ( n3184 & n3185 ) ;
  assign n3187 = ( ~n3009 & n3185 ) | ( ~n3009 & n3186 ) | ( n3185 & n3186 ) ;
  assign n3188 = n3183 & n3184 ;
  assign n3189 = n3005 | n3006 ;
  assign n3190 = n3183 | n3184 ;
  assign n3191 = n3188 | n3190 ;
  assign n3192 = ( n3188 & n3189 ) | ( n3188 & n3191 ) | ( n3189 & n3191 ) ;
  assign n3193 = ( n2994 & n3005 ) | ( n2994 & n3189 ) | ( n3005 & n3189 ) ;
  assign n3194 = ( n3188 & n3191 ) | ( n3188 & n3193 ) | ( n3191 & n3193 ) ;
  assign n3195 = ( n2998 & n3192 ) | ( n2998 & n3194 ) | ( n3192 & n3194 ) ;
  assign n3196 = n3041 | n3043 ;
  assign n3197 = ( n3041 & n3042 ) | ( n3041 & n3196 ) | ( n3042 & n3196 ) ;
  assign n3198 = n3052 | n3054 ;
  assign n3199 = ( n3052 & n3053 ) | ( n3052 & n3198 ) | ( n3053 & n3198 ) ;
  assign n3200 = n3197 | n3199 ;
  assign n3201 = n3197 & n3199 ;
  assign n3202 = n3200 & ~n3201 ;
  assign n3203 = n3149 | n3167 ;
  assign n3204 = ( n3149 & n3152 ) | ( n3149 & n3203 ) | ( n3152 & n3203 ) ;
  assign n3205 = n3202 | n3204 ;
  assign n3206 = n3202 & n3204 ;
  assign n3207 = n3205 & ~n3206 ;
  assign n3208 = n3046 | n3061 ;
  assign n3209 = ( n3061 & n3065 ) | ( n3061 & n3208 ) | ( n3065 & n3208 ) ;
  assign n3210 = n3207 | n3209 ;
  assign n3211 = n3207 & n3209 ;
  assign n3212 = n3210 & ~n3211 ;
  assign n3213 = n3125 | n3174 ;
  assign n3214 = n3212 & n3213 ;
  assign n3215 = n3212 | n3213 ;
  assign n3216 = ~n3214 & n3215 ;
  assign n3217 = n3073 | n3177 ;
  assign n3218 = ( n3073 & n3077 ) | ( n3073 & n3217 ) | ( n3077 & n3217 ) ;
  assign n3219 = n3216 & n3218 ;
  assign n3220 = n3216 | n3218 ;
  assign n3221 = ~n3219 & n3220 ;
  assign n3222 = n3088 | n3114 ;
  assign n3223 = n3088 & n3114 ;
  assign n3224 = n3222 & ~n3223 ;
  assign n3225 = n3098 | n3224 ;
  assign n3226 = n3098 & n3224 ;
  assign n3227 = n3225 & ~n3226 ;
  assign n3228 = n3106 | n3119 ;
  assign n3229 = n3144 | n3160 ;
  assign n3230 = n3144 & n3160 ;
  assign n3231 = n3229 & ~n3230 ;
  assign n3232 = n3133 | n3231 ;
  assign n3233 = n3133 & n3231 ;
  assign n3234 = n3232 & ~n3233 ;
  assign n3235 = n3105 | n3118 ;
  assign n3236 = n3234 & n3235 ;
  assign n3237 = n3105 & n3234 ;
  assign n3238 = ( n3228 & n3236 ) | ( n3228 & n3237 ) | ( n3236 & n3237 ) ;
  assign n3239 = n3234 | n3235 ;
  assign n3240 = n3105 | n3234 ;
  assign n3241 = ( n3228 & n3239 ) | ( n3228 & n3240 ) | ( n3239 & n3240 ) ;
  assign n3242 = ~n3238 & n3241 ;
  assign n3243 = n3227 & n3242 ;
  assign n3244 = n3227 | n3242 ;
  assign n3245 = ~n3243 & n3244 ;
  assign n3246 = n3027 & n3245 ;
  assign n3247 = ( n3031 & n3245 ) | ( n3031 & n3246 ) | ( n3245 & n3246 ) ;
  assign n3248 = n3027 | n3030 ;
  assign n3249 = ( n3027 & n3028 ) | ( n3027 & n3248 ) | ( n3028 & n3248 ) ;
  assign n3250 = ~n3247 & n3249 ;
  assign n3251 = n3245 & ~n3246 ;
  assign n3252 = ~n3031 & n3251 ;
  assign n3253 = n360 & n2267 ;
  assign n3254 = n2346 & n2388 ;
  assign n3255 = n3253 | n3254 ;
  assign n3256 = x9 & x31 ;
  assign n3257 = n2524 & n3256 ;
  assign n3258 = x26 & n3257 ;
  assign n3259 = ( x26 & ~n3255 ) | ( x26 & n3258 ) | ( ~n3255 & n3258 ) ;
  assign n3260 = x10 & n3259 ;
  assign n3261 = n3255 | n3257 ;
  assign n3262 = x5 & x31 ;
  assign n3263 = x9 & x27 ;
  assign n3264 = ( ~n3257 & n3262 ) | ( ~n3257 & n3263 ) | ( n3262 & n3263 ) ;
  assign n3265 = n3262 & n3263 ;
  assign n3266 = ( ~n3255 & n3264 ) | ( ~n3255 & n3265 ) | ( n3264 & n3265 ) ;
  assign n3267 = ~n3261 & n3266 ;
  assign n3268 = n3260 | n3267 ;
  assign n3269 = x12 & x24 ;
  assign n3270 = x13 & x23 ;
  assign n3271 = n3269 | n3270 ;
  assign n3272 = n647 & n1686 ;
  assign n3273 = n3271 | n3272 ;
  assign n3274 = x2 & x34 ;
  assign n3275 = ( ~n3272 & n3273 ) | ( ~n3272 & n3274 ) | ( n3273 & n3274 ) ;
  assign n3276 = ( n3272 & n3273 ) | ( n3272 & ~n3274 ) | ( n3273 & ~n3274 ) ;
  assign n3277 = ( ~n3273 & n3275 ) | ( ~n3273 & n3276 ) | ( n3275 & n3276 ) ;
  assign n3278 = n3268 & n3277 ;
  assign n3279 = n3268 & ~n3278 ;
  assign n3280 = x28 & x30 ;
  assign n3281 = n181 & n3280 ;
  assign n3282 = n200 & n2709 ;
  assign n3283 = n3281 | n3282 ;
  assign n3284 = n251 & n2369 ;
  assign n3285 = x30 & n3284 ;
  assign n3286 = ( x30 & ~n3283 ) | ( x30 & n3285 ) | ( ~n3283 & n3285 ) ;
  assign n3287 = x6 & n3286 ;
  assign n3288 = n3283 | n3284 ;
  assign n3289 = x7 & x29 ;
  assign n3290 = x8 & x28 ;
  assign n3291 = ( ~n3284 & n3289 ) | ( ~n3284 & n3290 ) | ( n3289 & n3290 ) ;
  assign n3292 = n3289 & n3290 ;
  assign n3293 = ( ~n3283 & n3291 ) | ( ~n3283 & n3292 ) | ( n3291 & n3292 ) ;
  assign n3294 = ~n3288 & n3293 ;
  assign n3295 = n3287 | n3294 ;
  assign n3296 = ~n3268 & n3277 ;
  assign n3297 = n3295 & ~n3296 ;
  assign n3298 = ~n3279 & n3297 ;
  assign n3299 = ~n3295 & n3296 ;
  assign n3300 = ( n3279 & ~n3295 ) | ( n3279 & n3299 ) | ( ~n3295 & n3299 ) ;
  assign n3301 = n3298 | n3300 ;
  assign n3302 = n790 & n1710 ;
  assign n3303 = n792 & n1585 ;
  assign n3304 = n3302 | n3303 ;
  assign n3305 = n795 & n1434 ;
  assign n3306 = x22 & n3305 ;
  assign n3307 = ( x22 & ~n3304 ) | ( x22 & n3306 ) | ( ~n3304 & n3306 ) ;
  assign n3308 = x14 & n3307 ;
  assign n3309 = n3304 | n3305 ;
  assign n3310 = x15 & x21 ;
  assign n3311 = x16 & x20 ;
  assign n3312 = ( ~n3305 & n3310 ) | ( ~n3305 & n3311 ) | ( n3310 & n3311 ) ;
  assign n3313 = n3310 & n3311 ;
  assign n3314 = ( ~n3304 & n3312 ) | ( ~n3304 & n3313 ) | ( n3312 & n3313 ) ;
  assign n3315 = ~n3309 & n3314 ;
  assign n3316 = n3308 | n3315 ;
  assign n3317 = x11 & x25 ;
  assign n3318 = x3 & x33 ;
  assign n3319 = x4 & x32 ;
  assign n3320 = ( ~n3317 & n3318 ) | ( ~n3317 & n3319 ) | ( n3318 & n3319 ) ;
  assign n3321 = x32 & x33 ;
  assign n3322 = n79 & n3321 ;
  assign n3323 = n3318 | n3319 ;
  assign n3324 = ( n3317 & n3322 ) | ( n3317 & n3323 ) | ( n3322 & n3323 ) ;
  assign n3325 = ( n3317 & n3320 ) | ( n3317 & ~n3324 ) | ( n3320 & ~n3324 ) ;
  assign n3326 = n3316 & n3325 ;
  assign n3327 = n3316 & ~n3326 ;
  assign n3328 = x0 & x36 ;
  assign n3329 = n3047 & n3328 ;
  assign n3330 = n3047 & ~n3329 ;
  assign n3331 = ~n3047 & n3328 ;
  assign n3332 = n3330 | n3331 ;
  assign n3333 = x1 & x35 ;
  assign n3334 = x17 & x19 ;
  assign n3335 = n3333 & n3334 ;
  assign n3336 = n3333 & ~n3335 ;
  assign n3337 = n3334 & ~n3335 ;
  assign n3338 = n3336 | n3337 ;
  assign n3339 = ~n3332 & n3338 ;
  assign n3340 = n3332 & ~n3338 ;
  assign n3341 = n3339 | n3340 ;
  assign n3342 = ~n3316 & n3325 ;
  assign n3343 = n3341 & ~n3342 ;
  assign n3344 = ~n3327 & n3343 ;
  assign n3345 = ~n3341 & n3342 ;
  assign n3346 = ( n3327 & ~n3341 ) | ( n3327 & n3345 ) | ( ~n3341 & n3345 ) ;
  assign n3347 = n3344 | n3346 ;
  assign n3348 = n3015 | n3018 ;
  assign n3349 = ( n3015 & n3016 ) | ( n3015 & n3348 ) | ( n3016 & n3348 ) ;
  assign n3350 = n3347 & n3349 ;
  assign n3351 = n3347 & ~n3350 ;
  assign n3352 = ~n3347 & n3349 ;
  assign n3353 = n3301 & n3352 ;
  assign n3354 = ( n3301 & n3351 ) | ( n3301 & n3353 ) | ( n3351 & n3353 ) ;
  assign n3355 = n3301 | n3352 ;
  assign n3356 = n3351 | n3355 ;
  assign n3357 = ~n3354 & n3356 ;
  assign n3358 = n3252 | n3357 ;
  assign n3359 = n3250 | n3358 ;
  assign n3360 = n3252 & n3357 ;
  assign n3361 = ( n3250 & n3357 ) | ( n3250 & n3360 ) | ( n3357 & n3360 ) ;
  assign n3362 = n3359 & ~n3361 ;
  assign n3363 = n3221 & n3362 ;
  assign n3364 = n3221 | n3362 ;
  assign n3365 = ~n3363 & n3364 ;
  assign n3366 = n3036 | n3180 ;
  assign n3367 = ( n3036 & n3039 ) | ( n3036 & n3366 ) | ( n3039 & n3366 ) ;
  assign n3368 = ( n3195 & n3365 ) | ( n3195 & ~n3367 ) | ( n3365 & ~n3367 ) ;
  assign n3369 = ( ~n3365 & n3367 ) | ( ~n3365 & n3368 ) | ( n3367 & n3368 ) ;
  assign n3370 = ( ~n3195 & n3368 ) | ( ~n3195 & n3369 ) | ( n3368 & n3369 ) ;
  assign n3371 = n3365 & n3367 ;
  assign n3372 = n3365 | n3367 ;
  assign n3373 = n3371 | n3372 ;
  assign n3374 = ( n3195 & n3371 ) | ( n3195 & n3373 ) | ( n3371 & n3373 ) ;
  assign n3375 = n3329 | n3338 ;
  assign n3376 = ( n3329 & n3332 ) | ( n3329 & n3375 ) | ( n3332 & n3375 ) ;
  assign n3377 = n3261 | n3376 ;
  assign n3378 = n3261 & n3376 ;
  assign n3379 = n3377 & ~n3378 ;
  assign n3380 = n723 & n2148 ;
  assign n3381 = n650 & n1686 ;
  assign n3382 = n3380 | n3381 ;
  assign n3383 = n792 & n1932 ;
  assign n3384 = x24 & n3383 ;
  assign n3385 = ( x24 & ~n3382 ) | ( x24 & n3384 ) | ( ~n3382 & n3384 ) ;
  assign n3386 = x13 & n3385 ;
  assign n3387 = n3382 | n3383 ;
  assign n3388 = x14 & x23 ;
  assign n3389 = x15 & x22 ;
  assign n3390 = ( ~n3383 & n3388 ) | ( ~n3383 & n3389 ) | ( n3388 & n3389 ) ;
  assign n3391 = n3388 & n3389 ;
  assign n3392 = ( ~n3382 & n3390 ) | ( ~n3382 & n3391 ) | ( n3390 & n3391 ) ;
  assign n3393 = ~n3387 & n3392 ;
  assign n3394 = n3386 | n3393 ;
  assign n3395 = ~n3379 & n3394 ;
  assign n3396 = n3379 & ~n3394 ;
  assign n3397 = n3395 | n3396 ;
  assign n3398 = ~n3272 & n3274 ;
  assign n3399 = ( n3272 & n3273 ) | ( n3272 & n3398 ) | ( n3273 & n3398 ) ;
  assign n3400 = n3317 & n3318 ;
  assign n3401 = n3322 | n3400 ;
  assign n3402 = n3317 & n3319 ;
  assign n3403 = n3401 | n3402 ;
  assign n3404 = n3309 | n3403 ;
  assign n3405 = n3309 & n3403 ;
  assign n3406 = n3404 & ~n3405 ;
  assign n3407 = n3399 | n3406 ;
  assign n3408 = n3399 & n3406 ;
  assign n3409 = n3407 & ~n3408 ;
  assign n3410 = ( n3316 & n3325 ) | ( n3316 & n3341 ) | ( n3325 & n3341 ) ;
  assign n3411 = n3409 | n3410 ;
  assign n3412 = n3409 & n3410 ;
  assign n3413 = n3411 & ~n3412 ;
  assign n3414 = ~n3397 & n3413 ;
  assign n3415 = n3397 & ~n3413 ;
  assign n3416 = n3414 | n3415 ;
  assign n3417 = n3211 & n3416 ;
  assign n3418 = ( n3214 & n3416 ) | ( n3214 & n3417 ) | ( n3416 & n3417 ) ;
  assign n3419 = n3211 | n3416 ;
  assign n3420 = n3214 | n3419 ;
  assign n3421 = ~n3418 & n3420 ;
  assign n3422 = x26 & x32 ;
  assign n3423 = n377 & n3422 ;
  assign n3424 = n618 & n2267 ;
  assign n3425 = n3423 | n3424 ;
  assign n3426 = x10 & x32 ;
  assign n3427 = n2524 & n3426 ;
  assign n3428 = x26 & n3427 ;
  assign n3429 = ( x26 & ~n3425 ) | ( x26 & n3428 ) | ( ~n3425 & n3428 ) ;
  assign n3430 = x11 & n3429 ;
  assign n3431 = n3425 | n3427 ;
  assign n3432 = x5 & x32 ;
  assign n3433 = x10 & x27 ;
  assign n3434 = ( ~n3427 & n3432 ) | ( ~n3427 & n3433 ) | ( n3432 & n3433 ) ;
  assign n3435 = n3432 & n3433 ;
  assign n3436 = ( ~n3425 & n3434 ) | ( ~n3425 & n3435 ) | ( n3434 & n3435 ) ;
  assign n3437 = ~n3431 & n3436 ;
  assign n3438 = n3430 | n3437 ;
  assign n3439 = n1077 | n1281 ;
  assign n3440 = n1020 & n1437 ;
  assign n3441 = x8 & x29 ;
  assign n3442 = ~n3440 & n3441 ;
  assign n3443 = n3439 | n3440 ;
  assign n3444 = ( n3440 & n3442 ) | ( n3440 & n3443 ) | ( n3442 & n3443 ) ;
  assign n3445 = n3439 & ~n3444 ;
  assign n3446 = ( ~n3439 & n3440 ) | ( ~n3439 & n3441 ) | ( n3440 & n3441 ) ;
  assign n3447 = n3441 & n3446 ;
  assign n3448 = n3445 | n3447 ;
  assign n3449 = n3438 & n3448 ;
  assign n3450 = n3438 & ~n3449 ;
  assign n3451 = n3448 & ~n3449 ;
  assign n3452 = n3450 | n3451 ;
  assign n3453 = n3133 | n3230 ;
  assign n3454 = ( n3230 & n3231 ) | ( n3230 & n3453 ) | ( n3231 & n3453 ) ;
  assign n3455 = n3452 | n3454 ;
  assign n3456 = n3452 & n3454 ;
  assign n3457 = n3455 & ~n3456 ;
  assign n3458 = n3201 | n3202 ;
  assign n3459 = ( n3201 & n3204 ) | ( n3201 & n3458 ) | ( n3204 & n3458 ) ;
  assign n3460 = n3457 | n3459 ;
  assign n3461 = n3457 & n3459 ;
  assign n3462 = n3460 & ~n3461 ;
  assign n3463 = x25 & n358 ;
  assign n3464 = x33 & n82 ;
  assign n3465 = n3463 | n3464 ;
  assign n3466 = x25 & x33 ;
  assign n3467 = n645 & n3466 ;
  assign n3468 = x37 & ~n3467 ;
  assign n3469 = n3465 & n3468 ;
  assign n3470 = x0 & x37 ;
  assign n3471 = ~n3469 & n3470 ;
  assign n3472 = n3467 | n3469 ;
  assign n3473 = x4 & x33 ;
  assign n3474 = x12 & x25 ;
  assign n3475 = ( ~n3467 & n3473 ) | ( ~n3467 & n3474 ) | ( n3473 & n3474 ) ;
  assign n3476 = n3473 & n3474 ;
  assign n3477 = ( ~n3469 & n3475 ) | ( ~n3469 & n3476 ) | ( n3475 & n3476 ) ;
  assign n3478 = ~n3472 & n3477 ;
  assign n3479 = n3471 | n3478 ;
  assign n3480 = x2 & x35 ;
  assign n3481 = x3 & x34 ;
  assign n3482 = n3480 | n3481 ;
  assign n3483 = x34 & x35 ;
  assign n3484 = n77 & n3483 ;
  assign n3485 = x16 & x21 ;
  assign n3486 = ~n3484 & n3485 ;
  assign n3487 = n3482 | n3484 ;
  assign n3488 = ( n3484 & n3486 ) | ( n3484 & n3487 ) | ( n3486 & n3487 ) ;
  assign n3489 = n3482 & ~n3488 ;
  assign n3490 = ~n3482 & n3485 ;
  assign n3491 = ( n3485 & ~n3486 ) | ( n3485 & n3490 ) | ( ~n3486 & n3490 ) ;
  assign n3492 = n3489 | n3491 ;
  assign n3493 = n3479 & n3492 ;
  assign n3494 = n3479 & ~n3493 ;
  assign n3495 = x9 & x28 ;
  assign n3496 = n667 & n3280 ;
  assign n3497 = x6 & x31 ;
  assign n3498 = n3495 & n3497 ;
  assign n3499 = n3496 | n3498 ;
  assign n3500 = n200 & n2965 ;
  assign n3501 = n3495 & n3500 ;
  assign n3502 = ( n3495 & ~n3499 ) | ( n3495 & n3501 ) | ( ~n3499 & n3501 ) ;
  assign n3503 = n3499 | n3500 ;
  assign n3504 = x7 & x30 ;
  assign n3505 = ( n3497 & ~n3500 ) | ( n3497 & n3504 ) | ( ~n3500 & n3504 ) ;
  assign n3506 = n3497 & n3504 ;
  assign n3507 = ( ~n3499 & n3505 ) | ( ~n3499 & n3506 ) | ( n3505 & n3506 ) ;
  assign n3508 = ~n3503 & n3507 ;
  assign n3509 = n3502 | n3508 ;
  assign n3510 = ~n3492 & n3509 ;
  assign n3511 = ( n3479 & n3509 ) | ( n3479 & n3510 ) | ( n3509 & n3510 ) ;
  assign n3512 = ~n3494 & n3511 ;
  assign n3513 = n3492 & ~n3509 ;
  assign n3514 = ~n3479 & n3513 ;
  assign n3515 = ( n3494 & ~n3509 ) | ( n3494 & n3514 ) | ( ~n3509 & n3514 ) ;
  assign n3516 = n3512 | n3515 ;
  assign n3517 = n3462 | n3516 ;
  assign n3518 = n3462 & n3516 ;
  assign n3519 = n3517 & ~n3518 ;
  assign n3520 = n3421 & n3519 ;
  assign n3521 = n3421 | n3519 ;
  assign n3522 = ~n3520 & n3521 ;
  assign n3523 = n3247 | n3361 ;
  assign n3524 = n3350 | n3354 ;
  assign n3525 = x36 & n970 ;
  assign n3526 = x1 & x36 ;
  assign n3527 = x19 | n3526 ;
  assign n3528 = ~n3525 & n3527 ;
  assign n3529 = n3335 & n3528 ;
  assign n3530 = n3528 & ~n3529 ;
  assign n3531 = n3335 & ~n3528 ;
  assign n3532 = n3288 & n3531 ;
  assign n3533 = ( n3288 & n3530 ) | ( n3288 & n3532 ) | ( n3530 & n3532 ) ;
  assign n3534 = n3288 | n3531 ;
  assign n3535 = n3530 | n3534 ;
  assign n3536 = ~n3533 & n3535 ;
  assign n3537 = n3098 | n3223 ;
  assign n3538 = ( n3223 & n3224 ) | ( n3223 & n3537 ) | ( n3224 & n3537 ) ;
  assign n3539 = n3536 & n3538 ;
  assign n3540 = n3536 | n3538 ;
  assign n3541 = ~n3539 & n3540 ;
  assign n3542 = n3295 & n3296 ;
  assign n3543 = ( n3279 & n3295 ) | ( n3279 & n3542 ) | ( n3295 & n3542 ) ;
  assign n3544 = n3278 | n3543 ;
  assign n3545 = n3541 & n3544 ;
  assign n3546 = n3541 | n3544 ;
  assign n3547 = ~n3545 & n3546 ;
  assign n3548 = n3227 | n3238 ;
  assign n3549 = ( n3238 & n3242 ) | ( n3238 & n3548 ) | ( n3242 & n3548 ) ;
  assign n3550 = n3547 & n3549 ;
  assign n3551 = n3547 | n3549 ;
  assign n3552 = ~n3550 & n3551 ;
  assign n3553 = n3524 & n3552 ;
  assign n3554 = n3524 | n3552 ;
  assign n3555 = ~n3553 & n3554 ;
  assign n3556 = n3247 & n3555 ;
  assign n3557 = ( n3361 & n3555 ) | ( n3361 & n3556 ) | ( n3555 & n3556 ) ;
  assign n3558 = n3523 & ~n3557 ;
  assign n3559 = n3555 & ~n3556 ;
  assign n3560 = ~n3361 & n3559 ;
  assign n3561 = n3522 & n3560 ;
  assign n3562 = ( n3522 & n3558 ) | ( n3522 & n3561 ) | ( n3558 & n3561 ) ;
  assign n3563 = n3522 | n3560 ;
  assign n3564 = n3558 | n3563 ;
  assign n3565 = ~n3562 & n3564 ;
  assign n3566 = n3219 | n3363 ;
  assign n3567 = ( n3374 & n3565 ) | ( n3374 & ~n3566 ) | ( n3565 & ~n3566 ) ;
  assign n3568 = ( ~n3565 & n3566 ) | ( ~n3565 & n3567 ) | ( n3566 & n3567 ) ;
  assign n3569 = ( ~n3374 & n3567 ) | ( ~n3374 & n3568 ) | ( n3567 & n3568 ) ;
  assign n3570 = n3565 & n3566 ;
  assign n3571 = n3565 | n3566 ;
  assign n3572 = n3373 & n3571 ;
  assign n3573 = n3371 & n3571 ;
  assign n3574 = ( n3195 & n3572 ) | ( n3195 & n3573 ) | ( n3572 & n3573 ) ;
  assign n3575 = n3570 | n3574 ;
  assign n3576 = ( n3397 & n3409 ) | ( n3397 & n3410 ) | ( n3409 & n3410 ) ;
  assign n3577 = n3461 | n3516 ;
  assign n3578 = ( n3461 & n3462 ) | ( n3461 & n3577 ) | ( n3462 & n3577 ) ;
  assign n3579 = n3576 & ~n3578 ;
  assign n3580 = n3576 & n3578 ;
  assign n3581 = n3578 & ~n3580 ;
  assign n3582 = n3579 | n3581 ;
  assign n3583 = n3472 | n3488 ;
  assign n3584 = n3472 & n3488 ;
  assign n3585 = n3583 & ~n3584 ;
  assign n3586 = n3387 | n3585 ;
  assign n3587 = n3387 & n3585 ;
  assign n3588 = n3586 & ~n3587 ;
  assign n3589 = n3449 | n3454 ;
  assign n3590 = ( n3449 & n3452 ) | ( n3449 & n3589 ) | ( n3452 & n3589 ) ;
  assign n3591 = n3588 | n3590 ;
  assign n3592 = n3588 & n3590 ;
  assign n3593 = n3591 & ~n3592 ;
  assign n3594 = x9 & x29 ;
  assign n3595 = x29 & x31 ;
  assign n3596 = n667 & n3595 ;
  assign n3597 = n313 & n2709 ;
  assign n3598 = n3596 | n3597 ;
  assign n3599 = n251 & n2965 ;
  assign n3600 = n3594 & n3599 ;
  assign n3601 = ( n3594 & ~n3598 ) | ( n3594 & n3600 ) | ( ~n3598 & n3600 ) ;
  assign n3602 = n3598 | n3599 ;
  assign n3603 = x7 & x31 ;
  assign n3604 = x8 & x30 ;
  assign n3605 = ( ~n3599 & n3603 ) | ( ~n3599 & n3604 ) | ( n3603 & n3604 ) ;
  assign n3606 = n3603 & n3604 ;
  assign n3607 = ( ~n3598 & n3605 ) | ( ~n3598 & n3606 ) | ( n3605 & n3606 ) ;
  assign n3608 = ~n3602 & n3607 ;
  assign n3609 = n3601 | n3608 ;
  assign n3610 = n795 & n1932 ;
  assign n3611 = x17 & x23 ;
  assign n3612 = n3310 & n3611 ;
  assign n3613 = n3610 | n3612 ;
  assign n3614 = n1023 & n1585 ;
  assign n3615 = x23 & n3614 ;
  assign n3616 = ( x23 & ~n3613 ) | ( x23 & n3615 ) | ( ~n3613 & n3615 ) ;
  assign n3617 = x15 & n3616 ;
  assign n3618 = n3613 | n3614 ;
  assign n3619 = x16 & x22 ;
  assign n3620 = x17 & x21 ;
  assign n3621 = ( ~n3614 & n3619 ) | ( ~n3614 & n3620 ) | ( n3619 & n3620 ) ;
  assign n3622 = n3619 & n3620 ;
  assign n3623 = ( ~n3613 & n3621 ) | ( ~n3613 & n3622 ) | ( n3621 & n3622 ) ;
  assign n3624 = ~n3618 & n3623 ;
  assign n3625 = n3617 | n3624 ;
  assign n3626 = x10 & x28 ;
  assign n3627 = x5 & x33 ;
  assign n3628 = x6 & x32 ;
  assign n3629 = ( ~n3626 & n3627 ) | ( ~n3626 & n3628 ) | ( n3627 & n3628 ) ;
  assign n3630 = n204 & n3321 ;
  assign n3631 = n3627 | n3628 ;
  assign n3632 = ( n3626 & n3630 ) | ( n3626 & n3631 ) | ( n3630 & n3631 ) ;
  assign n3633 = ( n3626 & n3629 ) | ( n3626 & ~n3632 ) | ( n3629 & ~n3632 ) ;
  assign n3634 = ( n3609 & n3625 ) | ( n3609 & ~n3633 ) | ( n3625 & ~n3633 ) ;
  assign n3635 = ( ~n3625 & n3633 ) | ( ~n3625 & n3634 ) | ( n3633 & n3634 ) ;
  assign n3636 = ( ~n3609 & n3634 ) | ( ~n3609 & n3635 ) | ( n3634 & n3635 ) ;
  assign n3637 = n3593 & n3636 ;
  assign n3638 = n3593 | n3636 ;
  assign n3639 = ~n3637 & n3638 ;
  assign n3640 = n3410 & n3636 ;
  assign n3641 = n3409 & n3636 ;
  assign n3642 = ( n3397 & n3640 ) | ( n3397 & n3641 ) | ( n3640 & n3641 ) ;
  assign n3643 = ( n3576 & n3593 ) | ( n3576 & n3642 ) | ( n3593 & n3642 ) ;
  assign n3644 = ~n3637 & n3643 ;
  assign n3645 = ~n3578 & n3644 ;
  assign n3646 = ( n3581 & n3639 ) | ( n3581 & n3645 ) | ( n3639 & n3645 ) ;
  assign n3647 = n3582 & ~n3646 ;
  assign n3653 = n3418 | n3519 ;
  assign n3654 = ( n3418 & n3421 ) | ( n3418 & n3653 ) | ( n3421 & n3653 ) ;
  assign n3649 = n3578 | n3637 ;
  assign n3650 = ( ~n3580 & n3637 ) | ( ~n3580 & n3649 ) | ( n3637 & n3649 ) ;
  assign n3648 = ~n3578 & n3643 ;
  assign n3651 = ( n3638 & ~n3648 ) | ( n3638 & n3650 ) | ( ~n3648 & n3650 ) ;
  assign n3652 = ~n3650 & n3651 ;
  assign n3655 = n3652 & n3654 ;
  assign n3656 = ( n3647 & n3654 ) | ( n3647 & n3655 ) | ( n3654 & n3655 ) ;
  assign n3657 = n3652 | n3654 ;
  assign n3658 = n3647 | n3657 ;
  assign n3659 = ~n3656 & n3658 ;
  assign n3660 = n3492 & n3509 ;
  assign n3661 = ~n3479 & n3660 ;
  assign n3662 = ( n3494 & n3509 ) | ( n3494 & n3661 ) | ( n3509 & n3661 ) ;
  assign n3663 = n3378 | n3394 ;
  assign n3664 = ( n3378 & n3379 ) | ( n3378 & n3663 ) | ( n3379 & n3663 ) ;
  assign n3665 = n3493 | n3664 ;
  assign n3666 = n3662 | n3665 ;
  assign n3667 = n3493 & n3664 ;
  assign n3668 = ( n3662 & n3664 ) | ( n3662 & n3667 ) | ( n3664 & n3667 ) ;
  assign n3669 = n3666 & ~n3668 ;
  assign n3670 = x1 & x37 ;
  assign n3671 = n1285 & n3670 ;
  assign n3672 = n1285 | n3670 ;
  assign n3673 = ~n3671 & n3672 ;
  assign n3674 = n3444 | n3673 ;
  assign n3675 = n3444 & n3673 ;
  assign n3676 = n3674 & ~n3675 ;
  assign n3677 = n3503 & n3676 ;
  assign n3678 = n3503 | n3676 ;
  assign n3679 = ~n3677 & n3678 ;
  assign n3680 = n3669 & n3679 ;
  assign n3681 = n3669 | n3679 ;
  assign n3682 = ~n3680 & n3681 ;
  assign n3683 = n3550 | n3682 ;
  assign n3684 = n3553 | n3683 ;
  assign n3685 = n3550 & n3682 ;
  assign n3686 = ( n3553 & n3682 ) | ( n3553 & n3685 ) | ( n3682 & n3685 ) ;
  assign n3687 = n3684 & ~n3686 ;
  assign n3688 = n3529 | n3533 ;
  assign n3689 = n490 & n2267 ;
  assign n3690 = x12 & x34 ;
  assign n3691 = n2264 & n3690 ;
  assign n3692 = n3689 | n3691 ;
  assign n3693 = x27 & x34 ;
  assign n3694 = n543 & n3693 ;
  assign n3695 = x26 & n3694 ;
  assign n3696 = ( x26 & ~n3692 ) | ( x26 & n3695 ) | ( ~n3692 & n3695 ) ;
  assign n3697 = x12 & n3696 ;
  assign n3698 = n3692 | n3694 ;
  assign n3699 = x4 & x34 ;
  assign n3700 = x11 & x27 ;
  assign n3701 = ( ~n3694 & n3699 ) | ( ~n3694 & n3700 ) | ( n3699 & n3700 ) ;
  assign n3702 = n3699 & n3700 ;
  assign n3703 = ( ~n3692 & n3701 ) | ( ~n3692 & n3702 ) | ( n3701 & n3702 ) ;
  assign n3704 = ~n3698 & n3703 ;
  assign n3705 = n3697 | n3704 ;
  assign n3706 = n3688 & n3705 ;
  assign n3707 = n3688 & ~n3706 ;
  assign n3709 = n3399 | n3405 ;
  assign n3710 = ( n3405 & n3406 ) | ( n3405 & n3709 ) | ( n3406 & n3709 ) ;
  assign n3708 = ~n3688 & n3705 ;
  assign n3711 = n3708 & n3710 ;
  assign n3712 = ( n3707 & n3710 ) | ( n3707 & n3711 ) | ( n3710 & n3711 ) ;
  assign n3713 = n3708 | n3710 ;
  assign n3714 = n3707 | n3713 ;
  assign n3715 = ~n3712 & n3714 ;
  assign n3716 = x13 & x25 ;
  assign n3717 = x14 & x24 ;
  assign n3718 = n3716 | n3717 ;
  assign n3719 = n650 & n1912 ;
  assign n3720 = x3 & x35 ;
  assign n3721 = ~n3719 & n3720 ;
  assign n3722 = n3718 | n3719 ;
  assign n3723 = ( n3719 & n3721 ) | ( n3719 & n3722 ) | ( n3721 & n3722 ) ;
  assign n3724 = n3718 & ~n3723 ;
  assign n3725 = ( ~n3718 & n3719 ) | ( ~n3718 & n3720 ) | ( n3719 & n3720 ) ;
  assign n3726 = n3720 & n3725 ;
  assign n3727 = n3724 | n3726 ;
  assign n3728 = x0 & x38 ;
  assign n3729 = x2 & x36 ;
  assign n3730 = n3728 | n3729 ;
  assign n3731 = x36 & x38 ;
  assign n3732 = n67 & n3731 ;
  assign n3733 = n3730 & ~n3732 ;
  assign n3734 = ( n3431 & ~n3525 ) | ( n3431 & n3733 ) | ( ~n3525 & n3733 ) ;
  assign n3735 = ( n3431 & n3525 ) | ( n3431 & ~n3733 ) | ( n3525 & ~n3733 ) ;
  assign n3736 = ( ~n3431 & n3734 ) | ( ~n3431 & n3735 ) | ( n3734 & n3735 ) ;
  assign n3737 = n3727 & n3736 ;
  assign n3738 = n3727 | n3736 ;
  assign n3739 = ~n3737 & n3738 ;
  assign n3740 = n3539 | n3541 ;
  assign n3741 = ( n3539 & n3544 ) | ( n3539 & n3740 ) | ( n3544 & n3740 ) ;
  assign n3742 = n3739 | n3741 ;
  assign n3743 = n3739 & n3741 ;
  assign n3744 = n3742 & ~n3743 ;
  assign n3745 = n3715 & n3744 ;
  assign n3746 = n3715 | n3744 ;
  assign n3747 = ~n3745 & n3746 ;
  assign n3748 = n3687 & n3747 ;
  assign n3749 = n3687 | n3747 ;
  assign n3750 = ~n3748 & n3749 ;
  assign n3751 = n3659 | n3750 ;
  assign n3752 = n3659 & n3750 ;
  assign n3753 = n3751 & ~n3752 ;
  assign n3754 = n3557 | n3562 ;
  assign n3755 = ( n3575 & n3753 ) | ( n3575 & ~n3754 ) | ( n3753 & ~n3754 ) ;
  assign n3756 = ( ~n3753 & n3754 ) | ( ~n3753 & n3755 ) | ( n3754 & n3755 ) ;
  assign n3757 = ( ~n3575 & n3755 ) | ( ~n3575 & n3756 ) | ( n3755 & n3756 ) ;
  assign n3758 = n3753 & n3754 ;
  assign n3759 = n3753 | n3754 ;
  assign n3760 = n3570 & n3759 ;
  assign n3761 = ( n3572 & n3759 ) | ( n3572 & n3760 ) | ( n3759 & n3760 ) ;
  assign n3762 = ( n3573 & n3759 ) | ( n3573 & n3760 ) | ( n3759 & n3760 ) ;
  assign n3763 = ( n3194 & n3761 ) | ( n3194 & n3762 ) | ( n3761 & n3762 ) ;
  assign n3764 = ( n3192 & n3761 ) | ( n3192 & n3762 ) | ( n3761 & n3762 ) ;
  assign n3765 = ( n2998 & n3763 ) | ( n2998 & n3764 ) | ( n3763 & n3764 ) ;
  assign n3766 = n3758 | n3765 ;
  assign n3767 = x3 & x36 ;
  assign n3768 = x13 & x26 ;
  assign n3769 = n3767 & n3768 ;
  assign n3770 = x36 & x37 ;
  assign n3771 = n77 & n3770 ;
  assign n3772 = x13 & x37 ;
  assign n3773 = n2009 & n3772 ;
  assign n3774 = n3771 | n3773 ;
  assign n3775 = x37 & n3769 ;
  assign n3776 = ( x37 & ~n3774 ) | ( x37 & n3775 ) | ( ~n3774 & n3775 ) ;
  assign n3777 = x2 & n3776 ;
  assign n3778 = ( n3767 & n3768 ) | ( n3767 & ~n3774 ) | ( n3768 & ~n3774 ) ;
  assign n3779 = ( ~n3769 & n3777 ) | ( ~n3769 & n3778 ) | ( n3777 & n3778 ) ;
  assign n3780 = n790 & n1557 ;
  assign n3781 = n792 & n1912 ;
  assign n3782 = n3780 | n3781 ;
  assign n3783 = n795 & n1686 ;
  assign n3784 = x25 & n3783 ;
  assign n3785 = ( x25 & ~n3782 ) | ( x25 & n3784 ) | ( ~n3782 & n3784 ) ;
  assign n3786 = x14 & n3785 ;
  assign n3787 = n3782 | n3783 ;
  assign n3788 = x15 & x24 ;
  assign n3789 = x16 & x23 ;
  assign n3790 = ( ~n3783 & n3788 ) | ( ~n3783 & n3789 ) | ( n3788 & n3789 ) ;
  assign n3791 = n3788 & n3789 ;
  assign n3792 = ( ~n3782 & n3790 ) | ( ~n3782 & n3791 ) | ( n3790 & n3791 ) ;
  assign n3793 = ~n3787 & n3792 ;
  assign n3794 = n3786 | n3793 ;
  assign n3795 = n3779 & n3794 ;
  assign n3796 = n3779 & ~n3795 ;
  assign n3797 = n3794 & ~n3795 ;
  assign n3798 = n3796 | n3797 ;
  assign n3799 = x6 & x33 ;
  assign n3800 = n200 & n3321 ;
  assign n3801 = x9 & x30 ;
  assign n3802 = n3799 & n3801 ;
  assign n3803 = n3800 | n3802 ;
  assign n3804 = n667 & n2546 ;
  assign n3805 = n3799 & n3804 ;
  assign n3806 = ( n3799 & ~n3803 ) | ( n3799 & n3805 ) | ( ~n3803 & n3805 ) ;
  assign n3807 = n3803 | n3804 ;
  assign n3808 = x7 & x32 ;
  assign n3809 = ( n3801 & ~n3804 ) | ( n3801 & n3808 ) | ( ~n3804 & n3808 ) ;
  assign n3810 = n3801 & n3808 ;
  assign n3811 = ( ~n3803 & n3809 ) | ( ~n3803 & n3810 ) | ( n3809 & n3810 ) ;
  assign n3812 = ~n3807 & n3811 ;
  assign n3813 = n3806 | n3812 ;
  assign n3814 = ~n3798 & n3813 ;
  assign n3815 = n3798 & ~n3813 ;
  assign n3816 = n3814 | n3815 ;
  assign n3817 = ( n3493 & n3664 ) | ( n3493 & n3679 ) | ( n3664 & n3679 ) ;
  assign n3818 = n3664 | n3679 ;
  assign n3819 = ( n3662 & n3817 ) | ( n3662 & n3818 ) | ( n3817 & n3818 ) ;
  assign n3820 = n3816 | n3819 ;
  assign n3821 = n3816 & n3819 ;
  assign n3822 = n3820 & ~n3821 ;
  assign n3823 = n3588 | n3636 ;
  assign n3824 = ( n3590 & n3636 ) | ( n3590 & n3823 ) | ( n3636 & n3823 ) ;
  assign n3825 = ( n3592 & n3593 ) | ( n3592 & n3824 ) | ( n3593 & n3824 ) ;
  assign n3826 = n3822 & n3825 ;
  assign n3827 = n3822 | n3825 ;
  assign n3828 = ~n3826 & n3827 ;
  assign n3829 = ( n3581 & n3638 ) | ( n3581 & n3648 ) | ( n3638 & n3648 ) ;
  assign n3830 = ( n3576 & n3578 ) | ( n3576 & n3638 ) | ( n3578 & n3638 ) ;
  assign n3831 = ~n3576 & n3636 ;
  assign n3832 = n3593 & n3831 ;
  assign n3833 = ( ~n3578 & n3637 ) | ( ~n3578 & n3832 ) | ( n3637 & n3832 ) ;
  assign n3834 = n3830 & ~n3833 ;
  assign n3835 = n3602 | n3698 ;
  assign n3836 = n3602 & n3698 ;
  assign n3837 = n3835 & ~n3836 ;
  assign n3838 = n3626 & n3627 ;
  assign n3839 = n3630 | n3838 ;
  assign n3840 = n3626 & n3628 ;
  assign n3841 = n3839 | n3840 ;
  assign n3842 = n3837 | n3841 ;
  assign n3843 = n3837 & n3841 ;
  assign n3844 = n3842 & ~n3843 ;
  assign n3845 = n3706 & n3844 ;
  assign n3846 = ( n3712 & n3844 ) | ( n3712 & n3845 ) | ( n3844 & n3845 ) ;
  assign n3847 = n3706 | n3844 ;
  assign n3848 = n3712 | n3847 ;
  assign n3849 = ~n3846 & n3848 ;
  assign n3850 = x18 & x21 ;
  assign n3851 = n1437 | n3850 ;
  assign n3852 = n1077 & n1434 ;
  assign n3853 = x8 & x31 ;
  assign n3854 = ~n3852 & n3853 ;
  assign n3855 = n3851 | n3852 ;
  assign n3856 = ( n3852 & n3854 ) | ( n3852 & n3855 ) | ( n3854 & n3855 ) ;
  assign n3857 = n3851 & ~n3856 ;
  assign n3858 = ( ~n3851 & n3852 ) | ( ~n3851 & n3853 ) | ( n3852 & n3853 ) ;
  assign n3859 = n3853 & n3858 ;
  assign n3860 = n3857 | n3859 ;
  assign n3861 = x4 & x35 ;
  assign n3862 = x12 & x27 ;
  assign n3863 = n3861 | n3862 ;
  assign n3864 = x17 & x22 ;
  assign n3865 = ( n3861 & n3862 ) | ( n3861 & n3864 ) | ( n3862 & n3864 ) ;
  assign n3866 = n3863 & ~n3865 ;
  assign n3867 = n3861 & n3862 ;
  assign n3868 = n3864 & ~n3867 ;
  assign n3869 = ~n3863 & n3864 ;
  assign n3870 = ( n3864 & ~n3868 ) | ( n3864 & n3869 ) | ( ~n3868 & n3869 ) ;
  assign n3871 = n3866 | n3870 ;
  assign n3872 = n3860 & n3871 ;
  assign n3873 = n3860 & ~n3872 ;
  assign n3874 = x5 & x34 ;
  assign n3875 = n1996 & n3874 ;
  assign n3876 = n618 & n2369 ;
  assign n3877 = n3875 | n3876 ;
  assign n3878 = x29 & x34 ;
  assign n3879 = n581 & n3878 ;
  assign n3880 = n1996 & n3879 ;
  assign n3881 = ( n1996 & ~n3877 ) | ( n1996 & n3880 ) | ( ~n3877 & n3880 ) ;
  assign n3882 = n3877 | n3879 ;
  assign n3883 = x10 & x29 ;
  assign n3884 = ( n3874 & ~n3879 ) | ( n3874 & n3883 ) | ( ~n3879 & n3883 ) ;
  assign n3885 = n3874 & n3883 ;
  assign n3886 = ( ~n3877 & n3884 ) | ( ~n3877 & n3885 ) | ( n3884 & n3885 ) ;
  assign n3887 = ~n3882 & n3886 ;
  assign n3888 = n3881 | n3887 ;
  assign n3889 = ~n3860 & n3871 ;
  assign n3890 = n3888 & ~n3889 ;
  assign n3891 = ~n3873 & n3890 ;
  assign n3892 = ~n3888 & n3889 ;
  assign n3893 = ( n3873 & ~n3888 ) | ( n3873 & n3892 ) | ( ~n3888 & n3892 ) ;
  assign n3894 = n3891 | n3893 ;
  assign n3895 = n3849 & n3894 ;
  assign n3896 = n3849 | n3894 ;
  assign n3897 = ~n3832 & n3896 ;
  assign n3898 = ~n3637 & n3896 ;
  assign n3899 = ( n3578 & n3897 ) | ( n3578 & n3898 ) | ( n3897 & n3898 ) ;
  assign n3900 = ~n3895 & n3899 ;
  assign n3901 = n3834 & ~n3900 ;
  assign n3902 = n3576 & n3894 ;
  assign n3903 = ( n3576 & n3849 ) | ( n3576 & n3902 ) | ( n3849 & n3902 ) ;
  assign n3904 = ~n3895 & n3903 ;
  assign n3905 = n3578 & n3904 ;
  assign n3906 = n3834 & ~n3905 ;
  assign n3907 = ( ~n3829 & n3901 ) | ( ~n3829 & n3906 ) | ( n3901 & n3906 ) ;
  assign n3908 = n3578 & n3903 ;
  assign n3909 = n3895 & n3896 ;
  assign n3910 = ~n3895 & n3909 ;
  assign n3911 = ~n3895 & n3896 ;
  assign n3912 = ( ~n3908 & n3910 ) | ( ~n3908 & n3911 ) | ( n3910 & n3911 ) ;
  assign n3913 = n3828 | n3912 ;
  assign n3914 = ( ~n3899 & n3910 ) | ( ~n3899 & n3911 ) | ( n3910 & n3911 ) ;
  assign n3915 = n3828 | n3914 ;
  assign n3916 = ( ~n3829 & n3913 ) | ( ~n3829 & n3915 ) | ( n3913 & n3915 ) ;
  assign n3917 = n3907 | n3916 ;
  assign n3918 = ~n3828 & n3917 ;
  assign n3919 = x0 & x39 ;
  assign n3920 = n3671 & n3919 ;
  assign n3921 = n3671 & ~n3920 ;
  assign n3922 = ~n3671 & n3919 ;
  assign n3923 = n3921 | n3922 ;
  assign n3924 = x1 & ~x38 ;
  assign n3925 = ( x1 & ~n1133 ) | ( x1 & n3924 ) | ( ~n1133 & n3924 ) ;
  assign n3926 = x38 & n3925 ;
  assign n3927 = x20 & ~x38 ;
  assign n3928 = ( x20 & ~n1133 ) | ( x20 & n3927 ) | ( ~n1133 & n3927 ) ;
  assign n3929 = n3926 | n3928 ;
  assign n3930 = ~n3923 & n3929 ;
  assign n3931 = n3923 & ~n3929 ;
  assign n3932 = n3930 | n3931 ;
  assign n3933 = n3503 | n3675 ;
  assign n3934 = ( n3675 & n3676 ) | ( n3675 & n3933 ) | ( n3676 & n3933 ) ;
  assign n3935 = n3932 | n3934 ;
  assign n3936 = n3932 & n3934 ;
  assign n3937 = n3935 & ~n3936 ;
  assign n3938 = n3387 | n3488 ;
  assign n3939 = ( n3387 & n3472 ) | ( n3387 & n3938 ) | ( n3472 & n3938 ) ;
  assign n3940 = ( n3584 & n3585 ) | ( n3584 & n3939 ) | ( n3585 & n3939 ) ;
  assign n3941 = n3937 | n3940 ;
  assign n3942 = n3937 & n3940 ;
  assign n3943 = n3941 & ~n3942 ;
  assign n3944 = n3525 | n3732 ;
  assign n3945 = ( n3732 & n3733 ) | ( n3732 & n3944 ) | ( n3733 & n3944 ) ;
  assign n3946 = n3723 | n3945 ;
  assign n3947 = n3723 & n3945 ;
  assign n3948 = n3946 & ~n3947 ;
  assign n3949 = n3618 | n3948 ;
  assign n3950 = n3618 & n3948 ;
  assign n3951 = n3949 & ~n3950 ;
  assign n3952 = n3625 & n3633 ;
  assign n3953 = n3625 & ~n3952 ;
  assign n3954 = n3601 & n3633 ;
  assign n3955 = ( n3608 & n3633 ) | ( n3608 & n3954 ) | ( n3633 & n3954 ) ;
  assign n3956 = ~n3625 & n3955 ;
  assign n3957 = ( n3609 & n3953 ) | ( n3609 & n3956 ) | ( n3953 & n3956 ) ;
  assign n3958 = n3730 & ~n3945 ;
  assign n3959 = n3525 & ~n3733 ;
  assign n3960 = n3431 & n3959 ;
  assign n3961 = ( n3431 & n3958 ) | ( n3431 & n3960 ) | ( n3958 & n3960 ) ;
  assign n3962 = n3737 | n3961 ;
  assign n3963 = n3952 & n3962 ;
  assign n3964 = ( n3957 & n3962 ) | ( n3957 & n3963 ) | ( n3962 & n3963 ) ;
  assign n3965 = n3952 | n3962 ;
  assign n3966 = n3957 | n3965 ;
  assign n3967 = ~n3964 & n3966 ;
  assign n3968 = n3951 & n3967 ;
  assign n3969 = n3951 | n3967 ;
  assign n3970 = ~n3968 & n3969 ;
  assign n3971 = n3943 & n3970 ;
  assign n3972 = n3943 | n3970 ;
  assign n3973 = ~n3971 & n3972 ;
  assign n3974 = n3715 | n3743 ;
  assign n3975 = ( n3743 & n3744 ) | ( n3743 & n3974 ) | ( n3744 & n3974 ) ;
  assign n3976 = n3973 & n3975 ;
  assign n3977 = n3973 | n3975 ;
  assign n3978 = ~n3976 & n3977 ;
  assign n3979 = n3686 | n3747 ;
  assign n3980 = ( n3686 & n3687 ) | ( n3686 & n3979 ) | ( n3687 & n3979 ) ;
  assign n3981 = n3978 & n3980 ;
  assign n3982 = n3978 | n3980 ;
  assign n3983 = ~n3981 & n3982 ;
  assign n3984 = n3917 & n3983 ;
  assign n3985 = ( ~n3829 & n3912 ) | ( ~n3829 & n3914 ) | ( n3912 & n3914 ) ;
  assign n3986 = n3907 | n3985 ;
  assign n3987 = n3983 & ~n3986 ;
  assign n3988 = ( n3918 & n3984 ) | ( n3918 & n3987 ) | ( n3984 & n3987 ) ;
  assign n3989 = n3917 | n3983 ;
  assign n3990 = ~n3983 & n3986 ;
  assign n3991 = ( n3918 & n3989 ) | ( n3918 & ~n3990 ) | ( n3989 & ~n3990 ) ;
  assign n3992 = ~n3988 & n3991 ;
  assign n3993 = n3656 | n3750 ;
  assign n3994 = ( n3656 & n3659 ) | ( n3656 & n3993 ) | ( n3659 & n3993 ) ;
  assign n3995 = ( n3766 & n3992 ) | ( n3766 & ~n3994 ) | ( n3992 & ~n3994 ) ;
  assign n3996 = ( ~n3992 & n3994 ) | ( ~n3992 & n3995 ) | ( n3994 & n3995 ) ;
  assign n3997 = ( ~n3766 & n3995 ) | ( ~n3766 & n3996 ) | ( n3995 & n3996 ) ;
  assign n3998 = n3828 & n3912 ;
  assign n3999 = n3828 & n3914 ;
  assign n4000 = ( ~n3829 & n3998 ) | ( ~n3829 & n3999 ) | ( n3998 & n3999 ) ;
  assign n4001 = ( n3828 & n3907 ) | ( n3828 & n4000 ) | ( n3907 & n4000 ) ;
  assign n4002 = ( n3829 & n3900 ) | ( n3829 & n3905 ) | ( n3900 & n3905 ) ;
  assign n4003 = n4001 | n4002 ;
  assign n4004 = n3769 | n3774 ;
  assign n4005 = n3882 | n4004 ;
  assign n4006 = n3882 & n4004 ;
  assign n4007 = n4005 & ~n4006 ;
  assign n4008 = n3865 | n4007 ;
  assign n4009 = n3865 & n4007 ;
  assign n4010 = n4008 & ~n4009 ;
  assign n4011 = n3888 & n3889 ;
  assign n4012 = ( n3873 & n3888 ) | ( n3873 & n4011 ) | ( n3888 & n4011 ) ;
  assign n4013 = n3872 | n4012 ;
  assign n4014 = n3795 | n3813 ;
  assign n4015 = ( n3795 & n3798 ) | ( n3795 & n4014 ) | ( n3798 & n4014 ) ;
  assign n4016 = n4013 | n4015 ;
  assign n4017 = n4013 & n4015 ;
  assign n4018 = n4016 & ~n4017 ;
  assign n4019 = n4010 & n4018 ;
  assign n4020 = n4010 | n4018 ;
  assign n4021 = ~n4019 & n4020 ;
  assign n4022 = n3846 | n3894 ;
  assign n4023 = ( n3846 & n3849 ) | ( n3846 & n4022 ) | ( n3849 & n4022 ) ;
  assign n4024 = n4021 & n4023 ;
  assign n4025 = n4021 | n4023 ;
  assign n4026 = ~n4024 & n4025 ;
  assign n4027 = n3821 | n3826 ;
  assign n4028 = n4026 & n4027 ;
  assign n4029 = n4026 | n4027 ;
  assign n4030 = ~n4028 & n4029 ;
  assign n4031 = n4002 & n4030 ;
  assign n4032 = ( n4001 & n4030 ) | ( n4001 & n4031 ) | ( n4030 & n4031 ) ;
  assign n4033 = n4003 & ~n4032 ;
  assign n4034 = n3787 | n3807 ;
  assign n4035 = n3787 & n3807 ;
  assign n4036 = n4034 & ~n4035 ;
  assign n4037 = n3920 | n3929 ;
  assign n4038 = ( n3920 & n3923 ) | ( n3920 & n4037 ) | ( n3923 & n4037 ) ;
  assign n4039 = n4036 | n4038 ;
  assign n4040 = n4036 & n4038 ;
  assign n4041 = n4039 & ~n4040 ;
  assign n4042 = n3936 | n3940 ;
  assign n4043 = ( n3936 & n3937 ) | ( n3936 & n4042 ) | ( n3937 & n4042 ) ;
  assign n4044 = n4041 | n4043 ;
  assign n4045 = n4041 & n4043 ;
  assign n4046 = n4044 & ~n4045 ;
  assign n4047 = x0 & x40 ;
  assign n4048 = x2 & x38 ;
  assign n4049 = n4047 | n4048 ;
  assign n4050 = x38 & x40 ;
  assign n4051 = n67 & n4050 ;
  assign n4052 = n4049 & ~n4051 ;
  assign n4053 = n1410 | n4051 ;
  assign n4054 = ( n4051 & n4052 ) | ( n4051 & n4053 ) | ( n4052 & n4053 ) ;
  assign n4055 = n4049 & ~n4054 ;
  assign n4056 = n1410 & ~n4052 ;
  assign n4057 = n4055 | n4056 ;
  assign n4058 = x7 & x33 ;
  assign n4059 = n667 & n2683 ;
  assign n4060 = n251 & n3321 ;
  assign n4061 = n4059 | n4060 ;
  assign n4062 = x31 & x32 ;
  assign n4063 = n313 & n4062 ;
  assign n4064 = n4058 & n4063 ;
  assign n4065 = ( n4058 & ~n4061 ) | ( n4058 & n4064 ) | ( ~n4061 & n4064 ) ;
  assign n4066 = n4061 | n4063 ;
  assign n4067 = x8 & x32 ;
  assign n4068 = ( n3256 & ~n4063 ) | ( n3256 & n4067 ) | ( ~n4063 & n4067 ) ;
  assign n4069 = n3256 & n4067 ;
  assign n4070 = ( ~n4061 & n4068 ) | ( ~n4061 & n4069 ) | ( n4068 & n4069 ) ;
  assign n4071 = ~n4066 & n4070 ;
  assign n4072 = n4065 | n4071 ;
  assign n4073 = n4057 & n4072 ;
  assign n4074 = n4057 & ~n4073 ;
  assign n4075 = x5 & x35 ;
  assign n4076 = x12 & x28 ;
  assign n4077 = n4075 & n4076 ;
  assign n4078 = x35 & x36 ;
  assign n4079 = n91 & n4078 ;
  assign n4080 = x12 & x36 ;
  assign n4081 = n2525 & n4080 ;
  assign n4082 = n4079 | n4081 ;
  assign n4083 = x36 & n4077 ;
  assign n4084 = ( x36 & ~n4082 ) | ( x36 & n4083 ) | ( ~n4082 & n4083 ) ;
  assign n4085 = x4 & n4084 ;
  assign n4086 = ( n4075 & n4076 ) | ( n4075 & ~n4082 ) | ( n4076 & ~n4082 ) ;
  assign n4087 = ( ~n4077 & n4085 ) | ( ~n4077 & n4086 ) | ( n4085 & n4086 ) ;
  assign n4088 = ~n4057 & n4072 ;
  assign n4089 = n4087 & n4088 ;
  assign n4090 = ( n4074 & n4087 ) | ( n4074 & n4089 ) | ( n4087 & n4089 ) ;
  assign n4091 = n4087 | n4088 ;
  assign n4092 = n4074 | n4091 ;
  assign n4093 = ~n4090 & n4092 ;
  assign n4094 = n4046 | n4093 ;
  assign n4095 = n4046 & n4093 ;
  assign n4096 = n4094 & ~n4095 ;
  assign n4097 = n3971 | n3975 ;
  assign n4098 = ( n3971 & n3973 ) | ( n3971 & n4097 ) | ( n3973 & n4097 ) ;
  assign n4099 = n4096 & n4098 ;
  assign n4100 = n4096 | n4098 ;
  assign n4101 = ~n4099 & n4100 ;
  assign n4102 = n913 & n1557 ;
  assign n4103 = n795 & n1912 ;
  assign n4104 = n4102 | n4103 ;
  assign n4105 = n1023 & n1686 ;
  assign n4106 = x25 & n4105 ;
  assign n4107 = ( x25 & ~n4104 ) | ( x25 & n4106 ) | ( ~n4104 & n4106 ) ;
  assign n4108 = x15 & n4107 ;
  assign n4109 = n4104 | n4105 ;
  assign n4110 = x16 & x24 ;
  assign n4111 = ( n3611 & ~n4105 ) | ( n3611 & n4110 ) | ( ~n4105 & n4110 ) ;
  assign n4112 = n3611 & n4110 ;
  assign n4113 = ( ~n4104 & n4111 ) | ( ~n4104 & n4112 ) | ( n4111 & n4112 ) ;
  assign n4114 = ~n4109 & n4113 ;
  assign n4115 = n4108 | n4114 ;
  assign n4116 = x13 & x27 ;
  assign n4117 = x14 & x26 ;
  assign n4118 = n4116 | n4117 ;
  assign n4119 = n650 & n2267 ;
  assign n4120 = n4118 | n4119 ;
  assign n4121 = x3 & x37 ;
  assign n4122 = ( ~n4119 & n4120 ) | ( ~n4119 & n4121 ) | ( n4120 & n4121 ) ;
  assign n4123 = ( n4119 & n4120 ) | ( n4119 & ~n4121 ) | ( n4120 & ~n4121 ) ;
  assign n4124 = ( ~n4120 & n4122 ) | ( ~n4120 & n4123 ) | ( n4122 & n4123 ) ;
  assign n4125 = n4115 & n4124 ;
  assign n4126 = n4115 & ~n4125 ;
  assign n4127 = x6 & x34 ;
  assign n4128 = x10 & x30 ;
  assign n4129 = n4127 & n4128 ;
  assign n4130 = n618 & n2709 ;
  assign n4131 = x11 & x34 ;
  assign n4132 = n3089 & n4131 ;
  assign n4133 = n4130 | n4132 ;
  assign n4134 = x29 & n4129 ;
  assign n4135 = ( x29 & ~n4133 ) | ( x29 & n4134 ) | ( ~n4133 & n4134 ) ;
  assign n4136 = x11 & n4135 ;
  assign n4137 = ( n4127 & n4128 ) | ( n4127 & ~n4133 ) | ( n4128 & ~n4133 ) ;
  assign n4138 = ( ~n4129 & n4136 ) | ( ~n4129 & n4137 ) | ( n4136 & n4137 ) ;
  assign n4139 = ~n4115 & n4124 ;
  assign n4140 = n4138 & ~n4139 ;
  assign n4141 = ~n4126 & n4140 ;
  assign n4142 = ~n4138 & n4139 ;
  assign n4143 = ( n4126 & ~n4138 ) | ( n4126 & n4142 ) | ( ~n4138 & n4142 ) ;
  assign n4144 = n4141 | n4143 ;
  assign n4145 = n3951 | n3964 ;
  assign n4146 = ( n3964 & n3967 ) | ( n3964 & n4145 ) | ( n3967 & n4145 ) ;
  assign n4147 = n4144 & n4146 ;
  assign n4148 = n4144 | n4146 ;
  assign n4149 = ~n4147 & n4148 ;
  assign n4150 = n3836 | n3841 ;
  assign n4151 = ( n3836 & n3837 ) | ( n3836 & n4150 ) | ( n3837 & n4150 ) ;
  assign n4152 = n3618 | n3947 ;
  assign n4153 = ( n3947 & n3948 ) | ( n3947 & n4152 ) | ( n3948 & n4152 ) ;
  assign n4154 = n4151 | n4153 ;
  assign n4155 = n4151 & n4153 ;
  assign n4156 = n4154 & ~n4155 ;
  assign n4157 = x38 & n1133 ;
  assign n4158 = x1 & x39 ;
  assign n4159 = n1432 & n4158 ;
  assign n4160 = n1432 | n4158 ;
  assign n4161 = ~n4159 & n4160 ;
  assign n4162 = n4157 & n4161 ;
  assign n4163 = n4157 | n4161 ;
  assign n4164 = ~n4162 & n4163 ;
  assign n4165 = n3856 & n4164 ;
  assign n4166 = n3856 | n4164 ;
  assign n4167 = ~n4165 & n4166 ;
  assign n4168 = n4156 & n4167 ;
  assign n4169 = n4156 | n4167 ;
  assign n4170 = ~n4168 & n4169 ;
  assign n4171 = n4149 & n4170 ;
  assign n4172 = n4149 | n4170 ;
  assign n4173 = ~n4171 & n4172 ;
  assign n4174 = n4101 & n4173 ;
  assign n4175 = n4101 | n4173 ;
  assign n4176 = ~n4174 & n4175 ;
  assign n4177 = n4030 & ~n4031 ;
  assign n4178 = ~n4001 & n4177 ;
  assign n4179 = n4176 & n4178 ;
  assign n4180 = ( n4033 & n4176 ) | ( n4033 & n4179 ) | ( n4176 & n4179 ) ;
  assign n4181 = n4176 | n4178 ;
  assign n4182 = n4033 | n4181 ;
  assign n4183 = ~n4180 & n4182 ;
  assign n4184 = n3981 | n3988 ;
  assign n4185 = n4183 & n4184 ;
  assign n4186 = n4183 | n4184 ;
  assign n4187 = ~n4185 & n4186 ;
  assign n4188 = n3992 & n3994 ;
  assign n4189 = n3992 | n3994 ;
  assign n4190 = n3758 & n4189 ;
  assign n4191 = n4188 | n4190 ;
  assign n4192 = n4188 | n4189 ;
  assign n4193 = ( n3765 & n4191 ) | ( n3765 & n4192 ) | ( n4191 & n4192 ) ;
  assign n4194 = n4187 | n4193 ;
  assign n4195 = n4186 & n4193 ;
  assign n4196 = ~n4185 & n4195 ;
  assign n4197 = n4194 & ~n4196 ;
  assign n4198 = ~n4119 & n4121 ;
  assign n4199 = ( n4119 & n4120 ) | ( n4119 & n4198 ) | ( n4120 & n4198 ) ;
  assign n4200 = n4054 | n4109 ;
  assign n4201 = n4054 & n4109 ;
  assign n4202 = n4200 & ~n4201 ;
  assign n4203 = n4199 | n4202 ;
  assign n4204 = n4199 & n4202 ;
  assign n4205 = n4203 & ~n4204 ;
  assign n4206 = n4073 & n4205 ;
  assign n4207 = ( n4090 & n4205 ) | ( n4090 & n4206 ) | ( n4205 & n4206 ) ;
  assign n4208 = n4073 | n4205 ;
  assign n4209 = n4090 | n4208 ;
  assign n4210 = ~n4207 & n4209 ;
  assign n4211 = x40 & n1232 ;
  assign n4212 = x1 & x40 ;
  assign n4213 = x21 | n4212 ;
  assign n4214 = ~n4211 & n4213 ;
  assign n4215 = n4066 | n4214 ;
  assign n4216 = n4066 & n4214 ;
  assign n4217 = n4215 & ~n4216 ;
  assign n4218 = n4129 | n4133 ;
  assign n4219 = n4217 & n4218 ;
  assign n4220 = n4217 | n4218 ;
  assign n4221 = ~n4219 & n4220 ;
  assign n4222 = n4210 & n4221 ;
  assign n4223 = n4210 | n4221 ;
  assign n4224 = ~n4222 & n4223 ;
  assign n4225 = n4045 | n4093 ;
  assign n4226 = ( n4045 & n4046 ) | ( n4045 & n4225 ) | ( n4046 & n4225 ) ;
  assign n4227 = n4224 & n4226 ;
  assign n4228 = n4224 | n4226 ;
  assign n4229 = ~n4227 & n4228 ;
  assign n4230 = n4144 | n4170 ;
  assign n4231 = ( n4146 & n4170 ) | ( n4146 & n4230 ) | ( n4170 & n4230 ) ;
  assign n4232 = ( n4147 & n4149 ) | ( n4147 & n4231 ) | ( n4149 & n4231 ) ;
  assign n4233 = n4229 | n4232 ;
  assign n4234 = n4229 & n4232 ;
  assign n4235 = n4233 & ~n4234 ;
  assign n4236 = n4099 | n4173 ;
  assign n4237 = ( n4099 & n4101 ) | ( n4099 & n4236 ) | ( n4101 & n4236 ) ;
  assign n4238 = n4235 | n4237 ;
  assign n4239 = n4235 & n4237 ;
  assign n4240 = n4238 & ~n4239 ;
  assign n4241 = n204 & n4078 ;
  assign n4242 = x30 & x36 ;
  assign n4243 = n377 & n4242 ;
  assign n4244 = n4241 | n4243 ;
  assign n4245 = x30 & x35 ;
  assign n4246 = n717 & n4245 ;
  assign n4247 = x36 & n4246 ;
  assign n4248 = ( x36 & ~n4244 ) | ( x36 & n4247 ) | ( ~n4244 & n4247 ) ;
  assign n4249 = x5 & n4248 ;
  assign n4250 = n4244 | n4246 ;
  assign n4251 = x6 & x35 ;
  assign n4252 = x11 & x30 ;
  assign n4253 = ( ~n4246 & n4251 ) | ( ~n4246 & n4252 ) | ( n4251 & n4252 ) ;
  assign n4254 = n4251 & n4252 ;
  assign n4255 = ( ~n4244 & n4253 ) | ( ~n4244 & n4254 ) | ( n4253 & n4254 ) ;
  assign n4256 = ~n4250 & n4255 ;
  assign n4257 = n4249 | n4256 ;
  assign n4258 = x19 & x22 ;
  assign n4259 = n1434 | n4258 ;
  assign n4260 = x8 & x33 ;
  assign n4261 = ( n1434 & n4258 ) | ( n1434 & n4260 ) | ( n4258 & n4260 ) ;
  assign n4262 = n4259 & ~n4261 ;
  assign n4263 = n1434 & n4258 ;
  assign n4264 = n4260 & ~n4263 ;
  assign n4265 = ~n4259 & n4260 ;
  assign n4266 = ( n4260 & ~n4264 ) | ( n4260 & n4265 ) | ( ~n4264 & n4265 ) ;
  assign n4267 = n4262 | n4266 ;
  assign n4268 = n4257 & n4267 ;
  assign n4269 = n4257 & ~n4268 ;
  assign n4270 = ~n4257 & n4267 ;
  assign n4271 = n3856 | n4162 ;
  assign n4272 = ( n4162 & n4164 ) | ( n4162 & n4271 ) | ( n4164 & n4271 ) ;
  assign n4273 = n4270 | n4272 ;
  assign n4274 = n4269 | n4273 ;
  assign n4275 = n4270 & n4272 ;
  assign n4276 = ( n4269 & n4272 ) | ( n4269 & n4275 ) | ( n4272 & n4275 ) ;
  assign n4277 = n4274 & ~n4276 ;
  assign n4278 = n4155 | n4167 ;
  assign n4279 = ( n4155 & n4156 ) | ( n4155 & n4278 ) | ( n4156 & n4278 ) ;
  assign n4280 = n4277 | n4279 ;
  assign n4281 = n4277 & n4279 ;
  assign n4282 = n4280 & ~n4281 ;
  assign n4283 = x4 & x37 ;
  assign n4284 = x12 & x29 ;
  assign n4285 = n4283 & n4284 ;
  assign n4286 = x27 & x37 ;
  assign n4287 = n789 & n4286 ;
  assign n4288 = n487 & n2075 ;
  assign n4289 = n4287 | n4288 ;
  assign n4290 = x27 & n4285 ;
  assign n4291 = ( x27 & ~n4289 ) | ( x27 & n4290 ) | ( ~n4289 & n4290 ) ;
  assign n4292 = x14 & n4291 ;
  assign n4293 = ( n4283 & n4284 ) | ( n4283 & ~n4289 ) | ( n4284 & ~n4289 ) ;
  assign n4294 = ( ~n4285 & n4292 ) | ( ~n4285 & n4293 ) | ( n4292 & n4293 ) ;
  assign n4295 = n1018 & n1557 ;
  assign n4296 = n1023 & n1912 ;
  assign n4297 = n4295 | n4296 ;
  assign n4298 = n1020 & n1686 ;
  assign n4299 = x25 & n4298 ;
  assign n4300 = ( x25 & ~n4297 ) | ( x25 & n4299 ) | ( ~n4297 & n4299 ) ;
  assign n4301 = x16 & n4300 ;
  assign n4302 = n4297 | n4298 ;
  assign n4303 = x17 & x24 ;
  assign n4304 = x18 & x23 ;
  assign n4305 = ( ~n4298 & n4303 ) | ( ~n4298 & n4304 ) | ( n4303 & n4304 ) ;
  assign n4306 = n4303 & n4304 ;
  assign n4307 = ( ~n4297 & n4305 ) | ( ~n4297 & n4306 ) | ( n4305 & n4306 ) ;
  assign n4308 = ~n4302 & n4307 ;
  assign n4309 = n4301 | n4308 ;
  assign n4310 = n4294 & n4309 ;
  assign n4311 = n4294 & ~n4310 ;
  assign n4312 = n4309 & ~n4310 ;
  assign n4313 = n4311 | n4312 ;
  assign n4314 = n360 & n4062 ;
  assign n4315 = x7 & x34 ;
  assign n4316 = n2388 & n4315 ;
  assign n4317 = n4314 | n4316 ;
  assign n4318 = x32 & x34 ;
  assign n4319 = n667 & n4318 ;
  assign n4320 = n2388 & n4319 ;
  assign n4321 = ( n2388 & ~n4317 ) | ( n2388 & n4320 ) | ( ~n4317 & n4320 ) ;
  assign n4322 = n4317 | n4319 ;
  assign n4323 = x9 & x32 ;
  assign n4324 = ( n4315 & ~n4319 ) | ( n4315 & n4323 ) | ( ~n4319 & n4323 ) ;
  assign n4325 = n4315 & n4323 ;
  assign n4326 = ( ~n4317 & n4324 ) | ( ~n4317 & n4325 ) | ( n4324 & n4325 ) ;
  assign n4327 = ~n4322 & n4326 ;
  assign n4328 = n4321 | n4327 ;
  assign n4329 = ~n4313 & n4328 ;
  assign n4330 = n4313 & ~n4328 ;
  assign n4331 = n4329 | n4330 ;
  assign n4332 = n4282 | n4331 ;
  assign n4333 = n4282 & n4331 ;
  assign n4334 = n4332 & ~n4333 ;
  assign n4335 = n4024 & n4334 ;
  assign n4336 = ( n4028 & n4334 ) | ( n4028 & n4335 ) | ( n4334 & n4335 ) ;
  assign n4337 = ( n4024 & n4028 ) | ( n4024 & ~n4336 ) | ( n4028 & ~n4336 ) ;
  assign n4378 = n4010 | n4017 ;
  assign n4379 = ( n4017 & n4018 ) | ( n4017 & n4378 ) | ( n4018 & n4378 ) ;
  assign n4338 = n4035 | n4040 ;
  assign n4339 = n3865 | n4006 ;
  assign n4340 = ( n4006 & n4007 ) | ( n4006 & n4339 ) | ( n4007 & n4339 ) ;
  assign n4341 = n4338 | n4340 ;
  assign n4342 = n4338 & n4340 ;
  assign n4343 = n4341 & ~n4342 ;
  assign n4344 = n4138 & n4139 ;
  assign n4345 = ( n4126 & n4138 ) | ( n4126 & n4344 ) | ( n4138 & n4344 ) ;
  assign n4346 = n4125 | n4345 ;
  assign n4347 = n4343 | n4346 ;
  assign n4348 = n4343 & n4346 ;
  assign n4349 = n4347 & ~n4348 ;
  assign n4350 = x39 & x41 ;
  assign n4351 = n67 & n4350 ;
  assign n4352 = x0 & x41 ;
  assign n4353 = x2 & x39 ;
  assign n4354 = n4352 | n4353 ;
  assign n4355 = ~n4351 & n4354 ;
  assign n4356 = n4159 & n4355 ;
  assign n4357 = n4159 | n4355 ;
  assign n4358 = ~n4356 & n4357 ;
  assign n4359 = n4077 | n4082 ;
  assign n4360 = n4358 & n4359 ;
  assign n4361 = n4358 | n4359 ;
  assign n4362 = ~n4360 & n4361 ;
  assign n4363 = x13 & x28 ;
  assign n4364 = x15 & x26 ;
  assign n4365 = n4363 | n4364 ;
  assign n4366 = n723 & n2895 ;
  assign n4367 = x3 & x38 ;
  assign n4368 = ~n4366 & n4367 ;
  assign n4369 = n4365 | n4366 ;
  assign n4370 = ( n4366 & n4368 ) | ( n4366 & n4369 ) | ( n4368 & n4369 ) ;
  assign n4371 = n4365 & ~n4370 ;
  assign n4372 = ( ~n4365 & n4366 ) | ( ~n4365 & n4367 ) | ( n4366 & n4367 ) ;
  assign n4373 = n4367 & n4372 ;
  assign n4374 = n4371 | n4373 ;
  assign n4375 = ~n4362 & n4374 ;
  assign n4376 = n4362 & ~n4374 ;
  assign n4377 = n4375 | n4376 ;
  assign n4380 = ( n4349 & ~n4377 ) | ( n4349 & n4379 ) | ( ~n4377 & n4379 ) ;
  assign n4381 = ( ~n4349 & n4377 ) | ( ~n4349 & n4379 ) | ( n4377 & n4379 ) ;
  assign n4382 = ( ~n4379 & n4380 ) | ( ~n4379 & n4381 ) | ( n4380 & n4381 ) ;
  assign n4383 = ~n4024 & n4334 ;
  assign n4384 = n4382 | n4383 ;
  assign n4385 = ( ~n4028 & n4382 ) | ( ~n4028 & n4384 ) | ( n4382 & n4384 ) ;
  assign n4386 = n4337 | n4385 ;
  assign n4387 = n4382 & n4383 ;
  assign n4388 = ~n4028 & n4387 ;
  assign n4389 = ( n4337 & n4382 ) | ( n4337 & n4388 ) | ( n4382 & n4388 ) ;
  assign n4390 = n4386 & ~n4389 ;
  assign n4391 = n4240 & n4390 ;
  assign n4392 = n4240 | n4390 ;
  assign n4393 = ~n4391 & n4392 ;
  assign n4394 = n4032 & n4393 ;
  assign n4395 = ( n4180 & n4393 ) | ( n4180 & n4394 ) | ( n4393 & n4394 ) ;
  assign n4396 = n4032 | n4393 ;
  assign n4397 = n4180 | n4396 ;
  assign n4398 = ~n4395 & n4397 ;
  assign n4399 = n4186 & n4192 ;
  assign n4400 = n4185 | n4399 ;
  assign n4401 = n4185 | n4186 ;
  assign n4402 = ( n4185 & n4191 ) | ( n4185 & n4401 ) | ( n4191 & n4401 ) ;
  assign n4403 = ( n3765 & n4400 ) | ( n3765 & n4402 ) | ( n4400 & n4402 ) ;
  assign n4404 = n4398 | n4403 ;
  assign n4405 = n4398 & n4403 ;
  assign n4406 = n4404 & ~n4405 ;
  assign n4407 = n4239 | n4391 ;
  assign n4408 = n4199 | n4201 ;
  assign n4409 = ( n4201 & n4202 ) | ( n4201 & n4408 ) | ( n4202 & n4408 ) ;
  assign n4410 = n4360 | n4374 ;
  assign n4411 = ( n4360 & n4362 ) | ( n4360 & n4410 ) | ( n4362 & n4410 ) ;
  assign n4412 = n4409 | n4411 ;
  assign n4413 = n4409 & n4411 ;
  assign n4414 = n4412 & ~n4413 ;
  assign n4415 = n4310 | n4328 ;
  assign n4416 = ( n4310 & n4313 ) | ( n4310 & n4415 ) | ( n4313 & n4415 ) ;
  assign n4417 = n4414 | n4416 ;
  assign n4418 = n4414 & n4416 ;
  assign n4419 = n4417 & ~n4418 ;
  assign n4420 = n4281 | n4331 ;
  assign n4421 = ( n4281 & n4282 ) | ( n4281 & n4420 ) | ( n4282 & n4420 ) ;
  assign n4422 = n4419 & n4421 ;
  assign n4423 = n4419 | n4421 ;
  assign n4424 = ~n4422 & n4423 ;
  assign n4425 = n4377 & n4379 ;
  assign n4426 = n4379 & ~n4425 ;
  assign n4427 = n4349 & n4377 ;
  assign n4428 = ~n4379 & n4427 ;
  assign n4429 = n4425 | n4428 ;
  assign n4430 = n4349 | n4377 ;
  assign n4431 = ( n4349 & n4379 ) | ( n4349 & n4430 ) | ( n4379 & n4430 ) ;
  assign n4432 = ( n4426 & n4429 ) | ( n4426 & n4431 ) | ( n4429 & n4431 ) ;
  assign n4433 = n4424 & n4432 ;
  assign n4434 = n4424 | n4432 ;
  assign n4435 = ~n4433 & n4434 ;
  assign n4436 = n4336 & n4435 ;
  assign n4437 = ( n4389 & n4435 ) | ( n4389 & n4436 ) | ( n4435 & n4436 ) ;
  assign n4438 = n4336 | n4435 ;
  assign n4439 = n4389 | n4438 ;
  assign n4440 = ~n4437 & n4439 ;
  assign n4441 = x0 & x42 ;
  assign n4442 = n4211 & n4441 ;
  assign n4443 = n4211 & ~n4442 ;
  assign n4444 = ~n4211 & n4441 ;
  assign n4445 = n4443 | n4444 ;
  assign n4446 = x1 & x41 ;
  assign n4447 = n1710 & n4446 ;
  assign n4448 = n4446 & ~n4447 ;
  assign n4449 = n1710 & ~n4447 ;
  assign n4450 = n4448 | n4449 ;
  assign n4451 = ~n4445 & n4450 ;
  assign n4452 = n4445 & ~n4450 ;
  assign n4453 = n4451 | n4452 ;
  assign n4454 = x5 & x37 ;
  assign n4455 = x12 & x30 ;
  assign n4456 = n4454 & n4455 ;
  assign n4457 = n647 & n2709 ;
  assign n4458 = n2864 & n3772 ;
  assign n4459 = n4457 | n4458 ;
  assign n4460 = x29 & n4456 ;
  assign n4461 = ( x29 & ~n4459 ) | ( x29 & n4460 ) | ( ~n4459 & n4460 ) ;
  assign n4462 = x13 & n4461 ;
  assign n4463 = ( n4454 & n4455 ) | ( n4454 & ~n4459 ) | ( n4455 & ~n4459 ) ;
  assign n4464 = ( ~n4456 & n4462 ) | ( ~n4456 & n4463 ) | ( n4462 & n4463 ) ;
  assign n4465 = n4453 & n4464 ;
  assign n4466 = n4453 | n4464 ;
  assign n4467 = ~n4465 & n4466 ;
  assign n4468 = n4216 | n4218 ;
  assign n4469 = ( n4216 & n4217 ) | ( n4216 & n4468 ) | ( n4217 & n4468 ) ;
  assign n4470 = n4467 | n4469 ;
  assign n4471 = n4467 & n4469 ;
  assign n4472 = n4470 & ~n4471 ;
  assign n4473 = n4207 | n4221 ;
  assign n4474 = ( n4207 & n4210 ) | ( n4207 & n4473 ) | ( n4210 & n4473 ) ;
  assign n4475 = n4472 | n4474 ;
  assign n4476 = n4472 & n4474 ;
  assign n4477 = n4475 & ~n4476 ;
  assign n4478 = n4269 | n4270 ;
  assign n4479 = n4261 | n4285 ;
  assign n4480 = n4289 | n4479 ;
  assign n4481 = n4261 & n4285 ;
  assign n4482 = ( n4261 & n4289 ) | ( n4261 & n4481 ) | ( n4289 & n4481 ) ;
  assign n4483 = n4480 & ~n4482 ;
  assign n4484 = n4250 | n4483 ;
  assign n4485 = n4250 & n4483 ;
  assign n4486 = n4484 & ~n4485 ;
  assign n4487 = n4268 | n4272 ;
  assign n4488 = n4486 & n4487 ;
  assign n4489 = n4268 & n4486 ;
  assign n4490 = ( n4478 & n4488 ) | ( n4478 & n4489 ) | ( n4488 & n4489 ) ;
  assign n4491 = n4486 | n4487 ;
  assign n4492 = n4268 | n4486 ;
  assign n4493 = ( n4478 & n4491 ) | ( n4478 & n4492 ) | ( n4491 & n4492 ) ;
  assign n4494 = ~n4490 & n4493 ;
  assign n4495 = n4302 | n4370 ;
  assign n4496 = n4302 & n4370 ;
  assign n4497 = n4495 & ~n4496 ;
  assign n4498 = n4159 | n4351 ;
  assign n4499 = ( n4351 & n4355 ) | ( n4351 & n4498 ) | ( n4355 & n4498 ) ;
  assign n4500 = n4497 | n4499 ;
  assign n4501 = n4497 & n4499 ;
  assign n4502 = n4500 & ~n4501 ;
  assign n4503 = n4494 & n4502 ;
  assign n4504 = n4494 | n4502 ;
  assign n4505 = ~n4503 & n4504 ;
  assign n4506 = n4477 & n4505 ;
  assign n4507 = n4477 | n4505 ;
  assign n4508 = ~n4506 & n4507 ;
  assign n4509 = x31 & x36 ;
  assign n4510 = n717 & n4509 ;
  assign n4511 = n200 & n4078 ;
  assign n4512 = n4510 | n4511 ;
  assign n4513 = x7 & x35 ;
  assign n4514 = x11 & x31 ;
  assign n4515 = n4513 & n4514 ;
  assign n4516 = x6 & n4515 ;
  assign n4517 = ( x6 & ~n4512 ) | ( x6 & n4516 ) | ( ~n4512 & n4516 ) ;
  assign n4518 = x36 & n4517 ;
  assign n4519 = n4513 | n4514 ;
  assign n4520 = ~n4515 & n4519 ;
  assign n4521 = ~n4512 & n4520 ;
  assign n4522 = ~n4322 & n4521 ;
  assign n4523 = ( ~n4322 & n4518 ) | ( ~n4322 & n4522 ) | ( n4518 & n4522 ) ;
  assign n4524 = n4322 & ~n4521 ;
  assign n4525 = ~n4518 & n4524 ;
  assign n4526 = n4523 | n4525 ;
  assign n4527 = n249 & n4318 ;
  assign n4528 = n360 & n3321 ;
  assign n4529 = n4527 | n4528 ;
  assign n4530 = x33 & x34 ;
  assign n4531 = n313 & n4530 ;
  assign n4532 = n3426 & n4531 ;
  assign n4533 = ( n3426 & ~n4529 ) | ( n3426 & n4532 ) | ( ~n4529 & n4532 ) ;
  assign n4534 = n4529 | n4531 ;
  assign n4535 = x8 & x34 ;
  assign n4536 = x9 & x33 ;
  assign n4537 = ( ~n4531 & n4535 ) | ( ~n4531 & n4536 ) | ( n4535 & n4536 ) ;
  assign n4538 = n4535 & n4536 ;
  assign n4539 = ( ~n4529 & n4537 ) | ( ~n4529 & n4538 ) | ( n4537 & n4538 ) ;
  assign n4540 = ~n4534 & n4539 ;
  assign n4541 = n4533 | n4540 ;
  assign n4542 = n4526 & n4541 ;
  assign n4543 = n4526 | n4541 ;
  assign n4544 = ~n4542 & n4543 ;
  assign n4545 = n4342 & n4544 ;
  assign n4546 = ( n4348 & n4544 ) | ( n4348 & n4545 ) | ( n4544 & n4545 ) ;
  assign n4547 = n4342 | n4544 ;
  assign n4548 = n4348 | n4547 ;
  assign n4549 = ~n4546 & n4548 ;
  assign n4550 = x3 & x39 ;
  assign n4551 = x16 & x26 ;
  assign n4552 = n4550 & n4551 ;
  assign n4553 = x16 & x40 ;
  assign n4554 = n2009 & n4553 ;
  assign n4555 = x39 & x40 ;
  assign n4556 = n77 & n4555 ;
  assign n4557 = n4554 | n4556 ;
  assign n4558 = x40 & n4552 ;
  assign n4559 = ( x40 & ~n4557 ) | ( x40 & n4558 ) | ( ~n4557 & n4558 ) ;
  assign n4560 = x2 & n4559 ;
  assign n4561 = ( n4550 & n4551 ) | ( n4550 & ~n4557 ) | ( n4551 & ~n4557 ) ;
  assign n4562 = ( ~n4552 & n4560 ) | ( ~n4552 & n4561 ) | ( n4560 & n4561 ) ;
  assign n4563 = n1557 & n3334 ;
  assign n4564 = n1020 & n1912 ;
  assign n4565 = n4563 | n4564 ;
  assign n4566 = n1077 & n1686 ;
  assign n4567 = x25 & n4566 ;
  assign n4568 = ( x25 & ~n4565 ) | ( x25 & n4567 ) | ( ~n4565 & n4567 ) ;
  assign n4569 = x17 & n4568 ;
  assign n4570 = n4565 | n4566 ;
  assign n4571 = x18 & x24 ;
  assign n4572 = x19 & x23 ;
  assign n4573 = ( ~n4566 & n4571 ) | ( ~n4566 & n4572 ) | ( n4571 & n4572 ) ;
  assign n4574 = n4571 & n4572 ;
  assign n4575 = ( ~n4565 & n4573 ) | ( ~n4565 & n4574 ) | ( n4573 & n4574 ) ;
  assign n4576 = ~n4570 & n4575 ;
  assign n4577 = n4569 | n4576 ;
  assign n4578 = n4562 & n4577 ;
  assign n4579 = n4562 & ~n4578 ;
  assign n4580 = n4577 & ~n4578 ;
  assign n4581 = n4579 | n4580 ;
  assign n4582 = n792 & n2372 ;
  assign n4583 = x15 & x38 ;
  assign n4584 = n2379 & n4583 ;
  assign n4585 = n4582 | n4584 ;
  assign n4586 = x14 & x38 ;
  assign n4587 = n2525 & n4586 ;
  assign n4588 = x27 & n4587 ;
  assign n4589 = ( x27 & ~n4585 ) | ( x27 & n4588 ) | ( ~n4585 & n4588 ) ;
  assign n4590 = x15 & n4589 ;
  assign n4591 = n4585 | n4587 ;
  assign n4592 = x4 & x38 ;
  assign n4593 = x14 & x28 ;
  assign n4594 = ( ~n4587 & n4592 ) | ( ~n4587 & n4593 ) | ( n4592 & n4593 ) ;
  assign n4595 = n4592 & n4593 ;
  assign n4596 = ( ~n4585 & n4594 ) | ( ~n4585 & n4595 ) | ( n4594 & n4595 ) ;
  assign n4597 = ~n4591 & n4596 ;
  assign n4598 = n4590 | n4597 ;
  assign n4599 = ~n4581 & n4598 ;
  assign n4600 = n4581 & ~n4598 ;
  assign n4601 = n4599 | n4600 ;
  assign n4602 = n4549 & n4601 ;
  assign n4603 = n4549 | n4601 ;
  assign n4604 = ~n4602 & n4603 ;
  assign n4605 = n4227 | n4234 ;
  assign n4606 = ( n4508 & ~n4604 ) | ( n4508 & n4605 ) | ( ~n4604 & n4605 ) ;
  assign n4607 = ( n4604 & ~n4605 ) | ( n4604 & n4606 ) | ( ~n4605 & n4606 ) ;
  assign n4608 = ( ~n4508 & n4606 ) | ( ~n4508 & n4607 ) | ( n4606 & n4607 ) ;
  assign n4609 = n4440 & n4608 ;
  assign n4610 = n4440 & ~n4609 ;
  assign n4611 = ~n4440 & n4608 ;
  assign n4612 = n4407 & n4611 ;
  assign n4613 = ( n4407 & n4610 ) | ( n4407 & n4612 ) | ( n4610 & n4612 ) ;
  assign n4614 = n4407 | n4611 ;
  assign n4615 = n4610 | n4614 ;
  assign n4616 = ~n4613 & n4615 ;
  assign n4617 = n4395 | n4397 ;
  assign n4618 = ( n4395 & n4403 ) | ( n4395 & n4617 ) | ( n4403 & n4617 ) ;
  assign n4619 = n4616 & n4618 ;
  assign n4620 = n4616 | n4618 ;
  assign n4621 = ~n4619 & n4620 ;
  assign n4622 = n4395 & n4615 ;
  assign n4623 = n4613 | n4622 ;
  assign n4624 = n4613 | n4615 ;
  assign n4625 = ( n4613 & n4617 ) | ( n4613 & n4624 ) | ( n4617 & n4624 ) ;
  assign n4626 = ( n4403 & n4623 ) | ( n4403 & n4625 ) | ( n4623 & n4625 ) ;
  assign n4627 = n4518 | n4521 ;
  assign n4628 = ( n4322 & n4541 ) | ( n4322 & n4627 ) | ( n4541 & n4627 ) ;
  assign n4629 = x42 & n1362 ;
  assign n4630 = x1 & x42 ;
  assign n4631 = x22 | n4630 ;
  assign n4632 = ~n4629 & n4631 ;
  assign n4633 = n4447 & n4632 ;
  assign n4634 = n4447 | n4632 ;
  assign n4635 = ~n4633 & n4634 ;
  assign n4636 = n4534 & n4635 ;
  assign n4637 = n4534 | n4635 ;
  assign n4638 = ~n4636 & n4637 ;
  assign n4639 = n4628 & n4638 ;
  assign n4640 = n4628 & ~n4639 ;
  assign n4641 = ~n4628 & n4638 ;
  assign n4642 = n4640 | n4641 ;
  assign n4643 = n4578 | n4598 ;
  assign n4644 = ( n4578 & n4581 ) | ( n4578 & n4643 ) | ( n4581 & n4643 ) ;
  assign n4645 = n4642 | n4644 ;
  assign n4646 = ~n4644 & n4645 ;
  assign n4647 = ( ~n4642 & n4645 ) | ( ~n4642 & n4646 ) | ( n4645 & n4646 ) ;
  assign n4648 = n4546 | n4601 ;
  assign n4649 = ( n4546 & n4549 ) | ( n4546 & n4648 ) | ( n4549 & n4648 ) ;
  assign n4650 = n4647 & n4649 ;
  assign n4651 = n4647 | n4649 ;
  assign n4652 = ~n4650 & n4651 ;
  assign n4653 = n4476 | n4505 ;
  assign n4654 = ( n4476 & n4477 ) | ( n4476 & n4653 ) | ( n4477 & n4653 ) ;
  assign n4655 = n4652 & n4654 ;
  assign n4656 = n4652 | n4654 ;
  assign n4657 = ~n4655 & n4656 ;
  assign n4658 = n4227 & n4604 ;
  assign n4659 = ( n4234 & n4604 ) | ( n4234 & n4658 ) | ( n4604 & n4658 ) ;
  assign n4660 = n4605 & ~n4659 ;
  assign n4661 = n4508 & n4604 ;
  assign n4662 = ~n4605 & n4661 ;
  assign n4663 = ( n4508 & n4660 ) | ( n4508 & n4662 ) | ( n4660 & n4662 ) ;
  assign n4664 = n4657 & n4659 ;
  assign n4665 = ( n4657 & n4663 ) | ( n4657 & n4664 ) | ( n4663 & n4664 ) ;
  assign n4666 = n4659 | n4663 ;
  assign n4667 = ~n4665 & n4666 ;
  assign n4668 = n4657 & ~n4665 ;
  assign n4669 = n4667 | n4668 ;
  assign n4670 = n4413 | n4418 ;
  assign n4671 = x0 & x43 ;
  assign n4672 = x3 & x40 ;
  assign n4673 = n4671 & n4672 ;
  assign n4674 = n79 & n4555 ;
  assign n4675 = x4 & x43 ;
  assign n4676 = n3919 & n4675 ;
  assign n4677 = n4674 | n4676 ;
  assign n4678 = x39 & n4673 ;
  assign n4679 = ( x39 & ~n4677 ) | ( x39 & n4678 ) | ( ~n4677 & n4678 ) ;
  assign n4680 = x4 & n4679 ;
  assign n4681 = ( n4671 & n4672 ) | ( n4671 & ~n4677 ) | ( n4672 & ~n4677 ) ;
  assign n4682 = ( ~n4673 & n4680 ) | ( ~n4673 & n4681 ) | ( n4680 & n4681 ) ;
  assign n4683 = n790 & n2075 ;
  assign n4684 = n792 & n2369 ;
  assign n4685 = n4683 | n4684 ;
  assign n4686 = n795 & n2372 ;
  assign n4687 = x29 & n4686 ;
  assign n4688 = ( x29 & ~n4685 ) | ( x29 & n4687 ) | ( ~n4685 & n4687 ) ;
  assign n4689 = x14 & n4688 ;
  assign n4690 = n4685 | n4686 ;
  assign n4691 = x15 & x28 ;
  assign n4692 = x16 & x27 ;
  assign n4693 = ( ~n4686 & n4691 ) | ( ~n4686 & n4692 ) | ( n4691 & n4692 ) ;
  assign n4694 = n4691 & n4692 ;
  assign n4695 = ( ~n4685 & n4693 ) | ( ~n4685 & n4694 ) | ( n4693 & n4694 ) ;
  assign n4696 = ~n4690 & n4695 ;
  assign n4697 = n4689 | n4696 ;
  assign n4698 = n4682 & n4697 ;
  assign n4699 = n4682 & ~n4698 ;
  assign n4700 = n4697 & ~n4698 ;
  assign n4701 = n4699 | n4700 ;
  assign n4702 = n2340 & n3334 ;
  assign n4703 = n1020 & n2511 ;
  assign n4704 = n4702 | n4703 ;
  assign n4705 = n1077 & n1912 ;
  assign n4706 = x26 & n4705 ;
  assign n4707 = ( x26 & ~n4704 ) | ( x26 & n4706 ) | ( ~n4704 & n4706 ) ;
  assign n4708 = x17 & n4707 ;
  assign n4709 = n4704 | n4705 ;
  assign n4710 = x18 & x25 ;
  assign n4711 = ( n1684 & ~n4705 ) | ( n1684 & n4710 ) | ( ~n4705 & n4710 ) ;
  assign n4712 = n1684 & n4710 ;
  assign n4713 = ( ~n4704 & n4711 ) | ( ~n4704 & n4712 ) | ( n4711 & n4712 ) ;
  assign n4714 = ~n4709 & n4713 ;
  assign n4715 = n4708 | n4714 ;
  assign n4716 = ~n4701 & n4715 ;
  assign n4717 = n4701 & ~n4715 ;
  assign n4718 = n4716 | n4717 ;
  assign n4719 = n251 & n4078 ;
  assign n4720 = x10 & x36 ;
  assign n4721 = n4058 & n4720 ;
  assign n4722 = n4719 | n4721 ;
  assign n4723 = n249 & n3129 ;
  assign n4724 = x36 & n4723 ;
  assign n4725 = ( x36 & ~n4722 ) | ( x36 & n4724 ) | ( ~n4722 & n4724 ) ;
  assign n4726 = x7 & n4725 ;
  assign n4727 = n4722 | n4723 ;
  assign n4728 = x8 & x35 ;
  assign n4729 = x10 & x33 ;
  assign n4730 = ( ~n4723 & n4728 ) | ( ~n4723 & n4729 ) | ( n4728 & n4729 ) ;
  assign n4731 = n4728 & n4729 ;
  assign n4732 = ( ~n4722 & n4730 ) | ( ~n4722 & n4731 ) | ( n4730 & n4731 ) ;
  assign n4733 = ~n4727 & n4732 ;
  assign n4734 = n4726 | n4733 ;
  assign n4735 = x20 & x23 ;
  assign n4736 = n1585 | n4735 ;
  assign n4737 = n1434 & n1932 ;
  assign n4738 = x9 & x34 ;
  assign n4739 = ~n4737 & n4738 ;
  assign n4740 = n4736 | n4737 ;
  assign n4741 = ( n4737 & n4739 ) | ( n4737 & n4740 ) | ( n4739 & n4740 ) ;
  assign n4742 = n4736 & ~n4741 ;
  assign n4743 = ( ~n4736 & n4737 ) | ( ~n4736 & n4738 ) | ( n4737 & n4738 ) ;
  assign n4744 = n4738 & n4743 ;
  assign n4745 = n4742 | n4744 ;
  assign n4746 = n4734 & n4745 ;
  assign n4747 = n4734 & ~n4746 ;
  assign n4748 = n4745 & ~n4746 ;
  assign n4749 = n4747 | n4748 ;
  assign n4750 = x5 & x38 ;
  assign n4751 = x13 & x30 ;
  assign n4752 = n4750 | n4751 ;
  assign n4753 = x2 & x41 ;
  assign n4754 = ( n4750 & n4751 ) | ( n4750 & n4753 ) | ( n4751 & n4753 ) ;
  assign n4755 = n4752 & ~n4754 ;
  assign n4756 = n4750 & n4751 ;
  assign n4757 = n4753 & ~n4756 ;
  assign n4758 = ~n4752 & n4753 ;
  assign n4759 = ( n4753 & ~n4757 ) | ( n4753 & n4758 ) | ( ~n4757 & n4758 ) ;
  assign n4760 = n4755 | n4759 ;
  assign n4761 = ~n4749 & n4760 ;
  assign n4762 = n4749 & ~n4760 ;
  assign n4763 = n4761 | n4762 ;
  assign n4764 = n4718 & ~n4763 ;
  assign n4765 = ~n4718 & n4763 ;
  assign n4766 = n4764 | n4765 ;
  assign n4767 = n4670 & n4766 ;
  assign n4768 = n4670 | n4766 ;
  assign n4769 = ~n4767 & n4768 ;
  assign n4770 = n4422 | n4424 ;
  assign n4771 = ( n4422 & n4432 ) | ( n4422 & n4770 ) | ( n4432 & n4770 ) ;
  assign n4772 = n4769 | n4771 ;
  assign n4773 = n4512 | n4515 ;
  assign n4774 = n4591 | n4773 ;
  assign n4775 = n4591 & n4773 ;
  assign n4776 = n4774 & ~n4775 ;
  assign n4777 = n4570 | n4776 ;
  assign n4778 = n4570 & n4776 ;
  assign n4779 = n4777 & ~n4778 ;
  assign n4780 = n4552 | n4557 ;
  assign n4781 = n4456 | n4459 ;
  assign n4782 = n4780 | n4781 ;
  assign n4783 = n4780 & n4781 ;
  assign n4784 = n4782 & ~n4783 ;
  assign n4785 = n4442 | n4450 ;
  assign n4786 = ( n4442 & n4445 ) | ( n4442 & n4785 ) | ( n4445 & n4785 ) ;
  assign n4787 = n4784 | n4786 ;
  assign n4788 = n4784 & n4786 ;
  assign n4789 = n4787 & ~n4788 ;
  assign n4790 = n4779 | n4789 ;
  assign n4791 = n4779 & n4789 ;
  assign n4792 = n4790 & ~n4791 ;
  assign n4793 = n4465 | n4469 ;
  assign n4794 = ( n4465 & n4467 ) | ( n4465 & n4793 ) | ( n4467 & n4793 ) ;
  assign n4795 = n4792 & n4794 ;
  assign n4796 = n4792 | n4794 ;
  assign n4797 = ~n4795 & n4796 ;
  assign n4810 = n4250 | n4482 ;
  assign n4811 = ( n4482 & n4483 ) | ( n4482 & n4810 ) | ( n4483 & n4810 ) ;
  assign n4798 = x6 & x37 ;
  assign n4799 = x11 & x32 ;
  assign n4800 = n4798 & n4799 ;
  assign n4801 = n490 & n4062 ;
  assign n4802 = x12 & x37 ;
  assign n4803 = n3497 & n4802 ;
  assign n4804 = n4801 | n4803 ;
  assign n4805 = x31 & n4800 ;
  assign n4806 = ( x31 & ~n4804 ) | ( x31 & n4805 ) | ( ~n4804 & n4805 ) ;
  assign n4807 = x12 & n4806 ;
  assign n4808 = ( n4798 & n4799 ) | ( n4798 & ~n4804 ) | ( n4799 & ~n4804 ) ;
  assign n4809 = ( ~n4800 & n4807 ) | ( ~n4800 & n4808 ) | ( n4807 & n4808 ) ;
  assign n4812 = n4809 & n4811 ;
  assign n4813 = n4811 & ~n4812 ;
  assign n4815 = n4496 | n4499 ;
  assign n4816 = ( n4496 & n4497 ) | ( n4496 & n4815 ) | ( n4497 & n4815 ) ;
  assign n4814 = n4809 & ~n4811 ;
  assign n4817 = n4814 & n4816 ;
  assign n4818 = ( n4813 & n4816 ) | ( n4813 & n4817 ) | ( n4816 & n4817 ) ;
  assign n4819 = n4814 | n4816 ;
  assign n4820 = n4813 | n4819 ;
  assign n4821 = ~n4818 & n4820 ;
  assign n4822 = n4490 | n4502 ;
  assign n4823 = ( n4490 & n4494 ) | ( n4490 & n4822 ) | ( n4494 & n4822 ) ;
  assign n4824 = n4821 & n4823 ;
  assign n4825 = n4821 | n4823 ;
  assign n4826 = ~n4824 & n4825 ;
  assign n4827 = n4797 & n4826 ;
  assign n4828 = n4797 | n4826 ;
  assign n4829 = ~n4827 & n4828 ;
  assign n4830 = ( n4422 & n4424 ) | ( n4422 & n4769 ) | ( n4424 & n4769 ) ;
  assign n4831 = n4422 & n4769 ;
  assign n4832 = ( n4432 & n4830 ) | ( n4432 & n4831 ) | ( n4830 & n4831 ) ;
  assign n4833 = n4829 & ~n4832 ;
  assign n4834 = n4772 & n4833 ;
  assign n4835 = ~n4829 & n4832 ;
  assign n4836 = ( n4772 & n4829 ) | ( n4772 & ~n4835 ) | ( n4829 & ~n4835 ) ;
  assign n4837 = ~n4834 & n4836 ;
  assign n4838 = n4669 | n4837 ;
  assign n4839 = n4669 & ~n4837 ;
  assign n4840 = ( ~n4669 & n4838 ) | ( ~n4669 & n4839 ) | ( n4838 & n4839 ) ;
  assign n4841 = n4437 | n4608 ;
  assign n4842 = ( n4437 & n4440 ) | ( n4437 & n4841 ) | ( n4440 & n4841 ) ;
  assign n4843 = ( n4626 & n4840 ) | ( n4626 & ~n4842 ) | ( n4840 & ~n4842 ) ;
  assign n4844 = ( ~n4840 & n4842 ) | ( ~n4840 & n4843 ) | ( n4842 & n4843 ) ;
  assign n4845 = ( ~n4626 & n4843 ) | ( ~n4626 & n4844 ) | ( n4843 & n4844 ) ;
  assign n4846 = n4840 & n4842 ;
  assign n4847 = n4840 | n4842 ;
  assign n4848 = n4613 & n4847 ;
  assign n4849 = ( n4622 & n4847 ) | ( n4622 & n4848 ) | ( n4847 & n4848 ) ;
  assign n4850 = n4846 | n4849 ;
  assign n4851 = n4846 | n4847 ;
  assign n4852 = ( n4625 & n4846 ) | ( n4625 & n4851 ) | ( n4846 & n4851 ) ;
  assign n4853 = ( n4403 & n4850 ) | ( n4403 & n4852 ) | ( n4850 & n4852 ) ;
  assign n4854 = x6 & x38 ;
  assign n4855 = x33 & x38 ;
  assign n4856 = n717 & n4855 ;
  assign n4857 = x37 & x38 ;
  assign n4858 = n200 & n4857 ;
  assign n4859 = n4856 | n4858 ;
  assign n4860 = x11 & x37 ;
  assign n4861 = n4058 & n4860 ;
  assign n4862 = n4854 & n4861 ;
  assign n4863 = ( n4854 & ~n4859 ) | ( n4854 & n4862 ) | ( ~n4859 & n4862 ) ;
  assign n4864 = n4859 | n4861 ;
  assign n4865 = x7 & x37 ;
  assign n4866 = x11 & x33 ;
  assign n4867 = ( ~n4861 & n4865 ) | ( ~n4861 & n4866 ) | ( n4865 & n4866 ) ;
  assign n4868 = n4865 & n4866 ;
  assign n4869 = ( ~n4859 & n4867 ) | ( ~n4859 & n4868 ) | ( n4867 & n4868 ) ;
  assign n4870 = ~n4864 & n4869 ;
  assign n4871 = n4863 | n4870 ;
  assign n4872 = x15 & x29 ;
  assign n4873 = x17 & x27 ;
  assign n4874 = n4872 | n4873 ;
  assign n4875 = n913 & n2075 ;
  assign n4876 = x3 & x41 ;
  assign n4877 = ~n4875 & n4876 ;
  assign n4878 = n4874 | n4875 ;
  assign n4879 = ( n4875 & n4877 ) | ( n4875 & n4878 ) | ( n4877 & n4878 ) ;
  assign n4880 = n4874 & ~n4879 ;
  assign n4881 = ( ~n4874 & n4875 ) | ( ~n4874 & n4876 ) | ( n4875 & n4876 ) ;
  assign n4882 = n4876 & n4881 ;
  assign n4883 = n4880 | n4882 ;
  assign n4884 = x18 & x26 ;
  assign n4885 = n1285 & n2340 ;
  assign n4886 = n1077 & n2511 ;
  assign n4887 = n4885 | n4886 ;
  assign n4888 = n1437 & n1912 ;
  assign n4889 = n4884 & n4888 ;
  assign n4890 = ( n4884 & ~n4887 ) | ( n4884 & n4889 ) | ( ~n4887 & n4889 ) ;
  assign n4891 = n4887 | n4888 ;
  assign n4892 = x19 & x25 ;
  assign n4893 = x20 & x24 ;
  assign n4894 = ( ~n4888 & n4892 ) | ( ~n4888 & n4893 ) | ( n4892 & n4893 ) ;
  assign n4895 = n4892 & n4893 ;
  assign n4896 = ( ~n4887 & n4894 ) | ( ~n4887 & n4895 ) | ( n4894 & n4895 ) ;
  assign n4897 = ~n4891 & n4896 ;
  assign n4898 = n4890 | n4897 ;
  assign n4899 = ( n4871 & n4883 ) | ( n4871 & ~n4898 ) | ( n4883 & ~n4898 ) ;
  assign n4900 = ( ~n4883 & n4898 ) | ( ~n4883 & n4899 ) | ( n4898 & n4899 ) ;
  assign n4901 = ( ~n4871 & n4899 ) | ( ~n4871 & n4900 ) | ( n4899 & n4900 ) ;
  assign n4902 = x4 & x40 ;
  assign n4903 = x14 & x30 ;
  assign n4904 = n4902 & n4903 ;
  assign n4905 = n2525 & n4553 ;
  assign n4906 = n790 & n3280 ;
  assign n4907 = n4905 | n4906 ;
  assign n4908 = x28 & n4904 ;
  assign n4909 = ( x28 & ~n4907 ) | ( x28 & n4908 ) | ( ~n4907 & n4908 ) ;
  assign n4910 = x16 & n4909 ;
  assign n4911 = ( n4902 & n4903 ) | ( n4902 & ~n4907 ) | ( n4903 & ~n4907 ) ;
  assign n4912 = ( ~n4904 & n4910 ) | ( ~n4904 & n4911 ) | ( n4910 & n4911 ) ;
  assign n4913 = x8 & x36 ;
  assign n4914 = x34 & x36 ;
  assign n4915 = n249 & n4914 ;
  assign n4916 = n313 & n4078 ;
  assign n4917 = n4915 | n4916 ;
  assign n4918 = n360 & n3483 ;
  assign n4919 = n4913 & n4918 ;
  assign n4920 = ( n4913 & ~n4917 ) | ( n4913 & n4919 ) | ( ~n4917 & n4919 ) ;
  assign n4921 = n4917 | n4918 ;
  assign n4922 = x9 & x35 ;
  assign n4923 = x10 & x34 ;
  assign n4924 = ( ~n4918 & n4922 ) | ( ~n4918 & n4923 ) | ( n4922 & n4923 ) ;
  assign n4925 = n4922 & n4923 ;
  assign n4926 = ( ~n4917 & n4924 ) | ( ~n4917 & n4925 ) | ( n4924 & n4925 ) ;
  assign n4927 = ~n4921 & n4926 ;
  assign n4928 = n4920 | n4927 ;
  assign n4929 = n4912 & n4928 ;
  assign n4930 = n4912 & ~n4929 ;
  assign n4931 = x12 & x32 ;
  assign n4932 = x13 & x31 ;
  assign n4933 = n4931 | n4932 ;
  assign n4934 = n647 & n4062 ;
  assign n4935 = x5 & x39 ;
  assign n4936 = ~n4934 & n4935 ;
  assign n4937 = n4933 | n4934 ;
  assign n4938 = ( n4934 & n4936 ) | ( n4934 & n4937 ) | ( n4936 & n4937 ) ;
  assign n4939 = n4933 & ~n4938 ;
  assign n4940 = ( ~n4933 & n4934 ) | ( ~n4933 & n4935 ) | ( n4934 & n4935 ) ;
  assign n4941 = n4935 & n4940 ;
  assign n4942 = n4939 | n4941 ;
  assign n4943 = ~n4912 & n4928 ;
  assign n4944 = n4942 & n4943 ;
  assign n4945 = ( n4930 & n4942 ) | ( n4930 & n4944 ) | ( n4942 & n4944 ) ;
  assign n4946 = n4942 | n4943 ;
  assign n4947 = n4930 | n4946 ;
  assign n4948 = ~n4945 & n4947 ;
  assign n4949 = n4901 | n4948 ;
  assign n4950 = n4901 & n4948 ;
  assign n4951 = n4949 & ~n4950 ;
  assign n4952 = n4642 & n4644 ;
  assign n4953 = n4639 | n4952 ;
  assign n4954 = n4951 & n4953 ;
  assign n4955 = n4951 | n4953 ;
  assign n4956 = ~n4954 & n4955 ;
  assign n4957 = n4650 | n4654 ;
  assign n4958 = ( n4650 & n4652 ) | ( n4650 & n4957 ) | ( n4652 & n4957 ) ;
  assign n4959 = n4956 | n4958 ;
  assign n4960 = n4956 & n4958 ;
  assign n4961 = n4959 & ~n4960 ;
  assign n4962 = n4800 | n4804 ;
  assign n4963 = n4690 | n4962 ;
  assign n4964 = n4690 & n4962 ;
  assign n4965 = n4963 & ~n4964 ;
  assign n4966 = x0 & x44 ;
  assign n4967 = x2 & x42 ;
  assign n4968 = n4966 | n4967 ;
  assign n4969 = x42 & x44 ;
  assign n4970 = n67 & n4969 ;
  assign n4971 = n4968 & ~n4970 ;
  assign n4972 = n4629 | n4970 ;
  assign n4973 = ( n4970 & n4971 ) | ( n4970 & n4972 ) | ( n4971 & n4972 ) ;
  assign n4974 = n4968 & ~n4973 ;
  assign n4975 = n4629 & ~n4971 ;
  assign n4976 = n4974 | n4975 ;
  assign n4977 = n4965 & n4976 ;
  assign n4978 = n4965 & ~n4977 ;
  assign n4979 = n4976 & ~n4977 ;
  assign n4980 = n4978 | n4979 ;
  assign n4981 = x1 & x43 ;
  assign n4982 = n1337 | n4981 ;
  assign n4983 = n1337 & n4981 ;
  assign n4984 = n4982 & ~n4983 ;
  assign n4985 = n4741 | n4984 ;
  assign n4986 = n4741 & n4984 ;
  assign n4987 = n4985 & ~n4986 ;
  assign n4988 = n4727 & n4987 ;
  assign n4989 = n4727 | n4987 ;
  assign n4990 = ~n4988 & n4989 ;
  assign n4991 = n4980 & n4990 ;
  assign n4992 = n4980 & ~n4991 ;
  assign n4993 = n4812 | n4818 ;
  assign n4994 = ~n4991 & n4993 ;
  assign n4995 = n4812 & n4990 ;
  assign n4996 = ( n4818 & n4990 ) | ( n4818 & n4995 ) | ( n4990 & n4995 ) ;
  assign n4997 = ( n4992 & n4994 ) | ( n4992 & n4996 ) | ( n4994 & n4996 ) ;
  assign n4998 = n4991 & ~n4993 ;
  assign n4999 = n4812 | n4990 ;
  assign n5000 = n4818 | n4999 ;
  assign n5001 = ( n4992 & ~n4998 ) | ( n4992 & n5000 ) | ( ~n4998 & n5000 ) ;
  assign n5002 = ~n4997 & n5001 ;
  assign n5003 = n4534 | n4633 ;
  assign n5004 = ( n4633 & n4635 ) | ( n4633 & n5003 ) | ( n4635 & n5003 ) ;
  assign n5005 = n4783 & n5004 ;
  assign n5006 = ( n4788 & n5004 ) | ( n4788 & n5005 ) | ( n5004 & n5005 ) ;
  assign n5007 = n4783 | n5004 ;
  assign n5008 = n4788 | n5007 ;
  assign n5009 = ~n5006 & n5008 ;
  assign n5010 = n4570 | n4775 ;
  assign n5011 = ( n4775 & n4776 ) | ( n4775 & n5010 ) | ( n4776 & n5010 ) ;
  assign n5012 = n5009 | n5011 ;
  assign n5013 = n5009 & n5011 ;
  assign n5014 = n5012 & ~n5013 ;
  assign n5015 = n4791 | n4795 ;
  assign n5016 = n5014 & n5015 ;
  assign n5017 = n5014 | n5015 ;
  assign n5018 = ~n5016 & n5017 ;
  assign n5019 = n5002 | n5018 ;
  assign n5020 = n5002 & n5018 ;
  assign n5021 = n5019 & ~n5020 ;
  assign n5022 = ~n4961 & n5021 ;
  assign n5023 = n4961 & ~n5021 ;
  assign n5024 = n5022 | n5023 ;
  assign n5025 = n4673 | n4754 ;
  assign n5026 = n4677 | n5025 ;
  assign n5027 = n4673 & n4754 ;
  assign n5028 = ( n4677 & n4754 ) | ( n4677 & n5027 ) | ( n4754 & n5027 ) ;
  assign n5029 = n5026 & ~n5028 ;
  assign n5030 = n4709 | n5029 ;
  assign n5031 = n4709 & n5029 ;
  assign n5032 = n5030 & ~n5031 ;
  assign n5033 = n4746 | n4760 ;
  assign n5034 = ( n4746 & n4749 ) | ( n4746 & n5033 ) | ( n4749 & n5033 ) ;
  assign n5035 = n4698 | n4715 ;
  assign n5036 = ( n4698 & n4701 ) | ( n4698 & n5035 ) | ( n4701 & n5035 ) ;
  assign n5037 = n5034 | n5036 ;
  assign n5038 = n5034 & n5036 ;
  assign n5039 = n5037 & ~n5038 ;
  assign n5040 = n5032 & n5039 ;
  assign n5041 = n5032 | n5039 ;
  assign n5042 = ~n5040 & n5041 ;
  assign n5043 = ( n4670 & n4718 ) | ( n4670 & n4763 ) | ( n4718 & n4763 ) ;
  assign n5044 = n5042 & n5043 ;
  assign n5045 = n5042 | n5043 ;
  assign n5046 = ~n5044 & n5045 ;
  assign n5047 = n4797 | n4824 ;
  assign n5048 = ( n4824 & n4826 ) | ( n4824 & n5047 ) | ( n4826 & n5047 ) ;
  assign n5049 = n5046 & n5048 ;
  assign n5050 = n5046 | n5048 ;
  assign n5051 = ~n5049 & n5050 ;
  assign n5052 = n4832 & n5051 ;
  assign n5053 = ( n4834 & n5051 ) | ( n4834 & n5052 ) | ( n5051 & n5052 ) ;
  assign n5054 = n4832 | n5051 ;
  assign n5055 = n4834 | n5054 ;
  assign n5056 = ~n5053 & n5055 ;
  assign n5057 = n5024 & ~n5056 ;
  assign n5058 = ~n5024 & n5056 ;
  assign n5059 = n5057 | n5058 ;
  assign n5060 = n4665 | n4837 ;
  assign n5061 = ( n4665 & n4669 ) | ( n4665 & n5060 ) | ( n4669 & n5060 ) ;
  assign n5062 = ( n4853 & n5059 ) | ( n4853 & ~n5061 ) | ( n5059 & ~n5061 ) ;
  assign n5063 = ( ~n5059 & n5061 ) | ( ~n5059 & n5062 ) | ( n5061 & n5062 ) ;
  assign n5064 = ( ~n4853 & n5062 ) | ( ~n4853 & n5063 ) | ( n5062 & n5063 ) ;
  assign n5065 = n5059 & n5061 ;
  assign n5066 = n5059 | n5061 ;
  assign n5067 = n5065 | n5066 ;
  assign n5068 = ( n4853 & n5065 ) | ( n4853 & n5067 ) | ( n5065 & n5067 ) ;
  assign n5069 = n1285 & n2724 ;
  assign n5070 = n1077 & n2267 ;
  assign n5071 = n5069 | n5070 ;
  assign n5072 = n1437 & n2511 ;
  assign n5073 = x27 & n5072 ;
  assign n5074 = ( x27 & ~n5071 ) | ( x27 & n5073 ) | ( ~n5071 & n5073 ) ;
  assign n5075 = x18 & n5074 ;
  assign n5076 = n5071 | n5072 ;
  assign n5077 = x19 & x26 ;
  assign n5078 = ( n1847 & ~n5072 ) | ( n1847 & n5077 ) | ( ~n5072 & n5077 ) ;
  assign n5079 = n1847 & n5077 ;
  assign n5080 = ( ~n5071 & n5078 ) | ( ~n5071 & n5079 ) | ( n5078 & n5079 ) ;
  assign n5081 = ~n5076 & n5080 ;
  assign n5082 = n5075 | n5081 ;
  assign n5083 = n4921 & n5082 ;
  assign n5084 = n4921 | n5082 ;
  assign n5085 = ~n5083 & n5084 ;
  assign n5086 = x5 & x40 ;
  assign n5087 = x13 & x32 ;
  assign n5088 = n5086 & n5087 ;
  assign n5089 = n650 & n4062 ;
  assign n5090 = x14 & x40 ;
  assign n5091 = n3262 & n5090 ;
  assign n5092 = n5089 | n5091 ;
  assign n5093 = x31 & n5088 ;
  assign n5094 = ( x31 & ~n5092 ) | ( x31 & n5093 ) | ( ~n5092 & n5093 ) ;
  assign n5095 = x14 & n5094 ;
  assign n5096 = ( n5086 & n5087 ) | ( n5086 & ~n5092 ) | ( n5087 & ~n5092 ) ;
  assign n5097 = ( ~n5088 & n5095 ) | ( ~n5088 & n5096 ) | ( n5095 & n5096 ) ;
  assign n5098 = n5085 & n5097 ;
  assign n5099 = n5085 & ~n5098 ;
  assign n5100 = ~n5085 & n5097 ;
  assign n5101 = n5099 | n5100 ;
  assign n5102 = x41 & x45 ;
  assign n5103 = n82 & n5102 ;
  assign n5104 = x43 & x45 ;
  assign n5105 = n67 & n5104 ;
  assign n5106 = n5103 | n5105 ;
  assign n5107 = x41 & x43 ;
  assign n5108 = n119 & n5107 ;
  assign n5109 = x45 & n5108 ;
  assign n5110 = ( x45 & ~n5106 ) | ( x45 & n5109 ) | ( ~n5106 & n5109 ) ;
  assign n5111 = x0 & n5110 ;
  assign n5112 = n5106 | n5108 ;
  assign n5113 = x2 & x43 ;
  assign n5114 = x4 & x41 ;
  assign n5115 = ( ~n5108 & n5113 ) | ( ~n5108 & n5114 ) | ( n5113 & n5114 ) ;
  assign n5116 = n5113 & n5114 ;
  assign n5117 = ( ~n5106 & n5115 ) | ( ~n5106 & n5116 ) | ( n5115 & n5116 ) ;
  assign n5118 = ~n5112 & n5117 ;
  assign n5119 = n5111 | n5118 ;
  assign n5120 = x7 & x38 ;
  assign n5121 = n667 & n3731 ;
  assign n5122 = n251 & n4857 ;
  assign n5123 = n5121 | n5122 ;
  assign n5124 = n313 & n3770 ;
  assign n5125 = n5120 & n5124 ;
  assign n5126 = ( n5120 & ~n5123 ) | ( n5120 & n5125 ) | ( ~n5123 & n5125 ) ;
  assign n5127 = n5123 | n5124 ;
  assign n5128 = x8 & x37 ;
  assign n5129 = x9 & x36 ;
  assign n5130 = ( ~n5124 & n5128 ) | ( ~n5124 & n5129 ) | ( n5128 & n5129 ) ;
  assign n5131 = n5128 & n5129 ;
  assign n5132 = ( ~n5123 & n5130 ) | ( ~n5123 & n5131 ) | ( n5130 & n5131 ) ;
  assign n5133 = ~n5127 & n5132 ;
  assign n5134 = n5126 | n5133 ;
  assign n5135 = n5119 & n5134 ;
  assign n5136 = n5119 & ~n5135 ;
  assign n5137 = n1787 | n1932 ;
  assign n5138 = n1585 & n1686 ;
  assign n5139 = x10 & x35 ;
  assign n5140 = ~n5138 & n5139 ;
  assign n5141 = n5137 | n5138 ;
  assign n5142 = ( n5138 & n5140 ) | ( n5138 & n5141 ) | ( n5140 & n5141 ) ;
  assign n5143 = n5137 & ~n5142 ;
  assign n5144 = ( ~n5137 & n5138 ) | ( ~n5137 & n5139 ) | ( n5138 & n5139 ) ;
  assign n5145 = n5139 & n5144 ;
  assign n5146 = n5143 | n5145 ;
  assign n5147 = ~n5119 & n5134 ;
  assign n5148 = n5146 & n5147 ;
  assign n5149 = ( n5136 & n5146 ) | ( n5136 & n5148 ) | ( n5146 & n5148 ) ;
  assign n5150 = n5146 | n5147 ;
  assign n5151 = n5136 | n5150 ;
  assign n5152 = ~n5149 & n5151 ;
  assign n5153 = n5101 & n5152 ;
  assign n5154 = n5101 & ~n5153 ;
  assign n5155 = ~n5101 & n5152 ;
  assign n5156 = n5154 | n5155 ;
  assign n5157 = n5032 | n5038 ;
  assign n5158 = ( n5038 & n5039 ) | ( n5038 & n5157 ) | ( n5039 & n5157 ) ;
  assign n5159 = ~n5156 & n5158 ;
  assign n5160 = n5156 & ~n5158 ;
  assign n5161 = n5159 | n5160 ;
  assign n5162 = n5044 | n5048 ;
  assign n5163 = ( n5044 & n5046 ) | ( n5044 & n5162 ) | ( n5046 & n5162 ) ;
  assign n5164 = n5161 | n5163 ;
  assign n5165 = n5161 & n5163 ;
  assign n5166 = n5164 & ~n5165 ;
  assign n5167 = n4709 | n5028 ;
  assign n5168 = ( n5028 & n5029 ) | ( n5028 & n5167 ) | ( n5029 & n5167 ) ;
  assign n5169 = n4964 | n5168 ;
  assign n5170 = n4977 | n5169 ;
  assign n5171 = n4964 & n5168 ;
  assign n5172 = ( n4977 & n5168 ) | ( n4977 & n5171 ) | ( n5168 & n5171 ) ;
  assign n5173 = n5170 & ~n5172 ;
  assign n5174 = n4727 | n4986 ;
  assign n5175 = ( n4986 & n4987 ) | ( n4986 & n5174 ) | ( n4987 & n5174 ) ;
  assign n5176 = n5173 | n5175 ;
  assign n5177 = n5173 & n5175 ;
  assign n5178 = n5176 & ~n5177 ;
  assign n5179 = n4991 | n5178 ;
  assign n5180 = n4997 | n5179 ;
  assign n5181 = n4991 & n5178 ;
  assign n5182 = ( n4997 & n5178 ) | ( n4997 & n5181 ) | ( n5178 & n5181 ) ;
  assign n5183 = n5180 & ~n5182 ;
  assign n5184 = n4904 | n4907 ;
  assign n5185 = n4864 | n5184 ;
  assign n5186 = n4864 & n5184 ;
  assign n5187 = n5185 & ~n5186 ;
  assign n5188 = n4938 | n5187 ;
  assign n5189 = n4938 & n5187 ;
  assign n5190 = n5188 & ~n5189 ;
  assign n5191 = n4929 | n4945 ;
  assign n5192 = n4883 & n4898 ;
  assign n5193 = n4883 & ~n5192 ;
  assign n5194 = n4871 & n4898 ;
  assign n5195 = ~n4883 & n5194 ;
  assign n5196 = ( n4871 & n5193 ) | ( n4871 & n5195 ) | ( n5193 & n5195 ) ;
  assign n5197 = n5192 | n5196 ;
  assign n5198 = n5191 | n5197 ;
  assign n5199 = n5191 & n5197 ;
  assign n5200 = n5198 & ~n5199 ;
  assign n5201 = n5190 & n5200 ;
  assign n5202 = n5190 | n5200 ;
  assign n5203 = ~n5201 & n5202 ;
  assign n5204 = n5183 & n5203 ;
  assign n5205 = n5183 | n5203 ;
  assign n5206 = ~n5204 & n5205 ;
  assign n5207 = n5166 & n5206 ;
  assign n5208 = n5166 | n5206 ;
  assign n5209 = ~n5207 & n5208 ;
  assign n5210 = n4879 | n4973 ;
  assign n5211 = n4879 & n4973 ;
  assign n5212 = n5210 & ~n5211 ;
  assign n5213 = n4891 | n5212 ;
  assign n5214 = n4891 & n5212 ;
  assign n5215 = n5213 & ~n5214 ;
  assign n5216 = n5006 | n5011 ;
  assign n5217 = ( n5006 & n5009 ) | ( n5006 & n5216 ) | ( n5009 & n5216 ) ;
  assign n5218 = n5215 | n5217 ;
  assign n5219 = n5215 & n5217 ;
  assign n5220 = n5218 & ~n5219 ;
  assign n5221 = x12 & x39 ;
  assign n5222 = n3799 & n5221 ;
  assign n5223 = n490 & n4530 ;
  assign n5224 = n5222 | n5223 ;
  assign n5225 = x34 & x39 ;
  assign n5226 = n717 & n5225 ;
  assign n5227 = x33 & n5226 ;
  assign n5228 = ( x33 & ~n5224 ) | ( x33 & n5227 ) | ( ~n5224 & n5227 ) ;
  assign n5229 = x12 & n5228 ;
  assign n5230 = n5224 | n5226 ;
  assign n5231 = x6 & x39 ;
  assign n5232 = ( n4131 & ~n5226 ) | ( n4131 & n5231 ) | ( ~n5226 & n5231 ) ;
  assign n5233 = n4131 & n5231 ;
  assign n5234 = ( ~n5224 & n5232 ) | ( ~n5224 & n5233 ) | ( n5232 & n5233 ) ;
  assign n5235 = ~n5230 & n5234 ;
  assign n5236 = n5229 | n5235 ;
  assign n5237 = n913 & n3280 ;
  assign n5238 = n795 & n2709 ;
  assign n5239 = n5237 | n5238 ;
  assign n5240 = n1023 & n2369 ;
  assign n5241 = n5239 | n5240 ;
  assign n5242 = x16 & x29 ;
  assign n5243 = x17 & x28 ;
  assign n5244 = ( ~n5240 & n5242 ) | ( ~n5240 & n5243 ) | ( n5242 & n5243 ) ;
  assign n5245 = n5242 & n5243 ;
  assign n5246 = ( ~n5239 & n5244 ) | ( ~n5239 & n5245 ) | ( n5244 & n5245 ) ;
  assign n5247 = ~n5241 & n5246 ;
  assign n5248 = x15 & x30 ;
  assign n5249 = n5240 & n5248 ;
  assign n5250 = ( ~n5239 & n5248 ) | ( ~n5239 & n5249 ) | ( n5248 & n5249 ) ;
  assign n5251 = n5247 | n5250 ;
  assign n5252 = n5236 & n5251 ;
  assign n5253 = n5236 & ~n5252 ;
  assign n5254 = n5251 & ~n5252 ;
  assign n5255 = n5253 | n5254 ;
  assign n5256 = x3 & x42 ;
  assign n5257 = n4983 | n5256 ;
  assign n5258 = n4983 & n5256 ;
  assign n5259 = n5257 & ~n5258 ;
  assign n5260 = x1 & ~x44 ;
  assign n5261 = ( x1 & ~n1397 ) | ( x1 & n5260 ) | ( ~n1397 & n5260 ) ;
  assign n5262 = x44 & n5261 ;
  assign n5263 = x23 & ~x44 ;
  assign n5264 = ( x23 & ~n1397 ) | ( x23 & n5263 ) | ( ~n1397 & n5263 ) ;
  assign n5265 = n5262 | n5264 ;
  assign n5266 = n5259 & n5265 ;
  assign n5267 = n5265 & ~n5266 ;
  assign n5268 = ( n5259 & ~n5266 ) | ( n5259 & n5267 ) | ( ~n5266 & n5267 ) ;
  assign n5269 = ~n5255 & n5268 ;
  assign n5270 = n5255 & ~n5268 ;
  assign n5271 = n5269 | n5270 ;
  assign n5272 = n5220 & n5271 ;
  assign n5273 = n5220 | n5271 ;
  assign n5274 = ~n5272 & n5273 ;
  assign n5276 = n5002 | n5016 ;
  assign n5277 = ( n5016 & n5018 ) | ( n5016 & n5276 ) | ( n5018 & n5276 ) ;
  assign n5275 = n4950 | n4954 ;
  assign n5278 = n5275 | n5277 ;
  assign n5279 = ~n5275 & n5277 ;
  assign n5280 = ( ~n5277 & n5278 ) | ( ~n5277 & n5279 ) | ( n5278 & n5279 ) ;
  assign n5281 = n5274 & ~n5280 ;
  assign n5282 = ~n5274 & n5280 ;
  assign n5283 = n5281 | n5282 ;
  assign n5284 = ( n4956 & n4958 ) | ( n4956 & n5021 ) | ( n4958 & n5021 ) ;
  assign n5285 = n5283 | n5284 ;
  assign n5286 = n5283 & n5284 ;
  assign n5287 = n5285 & ~n5286 ;
  assign n5288 = n5209 & n5287 ;
  assign n5289 = n5287 & ~n5288 ;
  assign n5290 = ( n5209 & ~n5288 ) | ( n5209 & n5289 ) | ( ~n5288 & n5289 ) ;
  assign n5291 = n4832 | n4834 ;
  assign n5292 = ( n5024 & n5051 ) | ( n5024 & n5291 ) | ( n5051 & n5291 ) ;
  assign n5293 = ( n5068 & n5290 ) | ( n5068 & ~n5292 ) | ( n5290 & ~n5292 ) ;
  assign n5294 = ( ~n5290 & n5292 ) | ( ~n5290 & n5293 ) | ( n5292 & n5293 ) ;
  assign n5295 = ( ~n5068 & n5293 ) | ( ~n5068 & n5294 ) | ( n5293 & n5294 ) ;
  assign n5296 = n5288 & ~n5292 ;
  assign n5297 = n5209 | n5292 ;
  assign n5298 = ( n5289 & ~n5296 ) | ( n5289 & n5297 ) | ( ~n5296 & n5297 ) ;
  assign n5299 = n5065 & n5298 ;
  assign n5300 = ~n5288 & n5292 ;
  assign n5301 = n5209 & n5292 ;
  assign n5302 = ( n5289 & n5300 ) | ( n5289 & n5301 ) | ( n5300 & n5301 ) ;
  assign n5303 = n5299 | n5302 ;
  assign n5304 = n5298 | n5302 ;
  assign n5305 = ( n5067 & n5302 ) | ( n5067 & n5304 ) | ( n5302 & n5304 ) ;
  assign n5306 = ( n4853 & n5303 ) | ( n4853 & n5305 ) | ( n5303 & n5305 ) ;
  assign n5307 = n5286 | n5288 ;
  assign n5308 = n5182 | n5204 ;
  assign n5309 = n5153 | n5158 ;
  assign n5310 = ( n5153 & n5156 ) | ( n5153 & n5309 ) | ( n5156 & n5309 ) ;
  assign n5311 = n5308 | n5310 ;
  assign n5312 = n5308 & n5310 ;
  assign n5313 = n5311 & ~n5312 ;
  assign n5314 = x6 & x40 ;
  assign n5315 = x13 & x33 ;
  assign n5316 = n5314 & n5315 ;
  assign n5317 = n650 & n3321 ;
  assign n5318 = n3628 & n5090 ;
  assign n5319 = n5317 | n5318 ;
  assign n5320 = x32 & n5316 ;
  assign n5321 = ( x32 & ~n5319 ) | ( x32 & n5320 ) | ( ~n5319 & n5320 ) ;
  assign n5322 = x14 & n5321 ;
  assign n5323 = ( n5314 & n5315 ) | ( n5314 & ~n5319 ) | ( n5315 & ~n5319 ) ;
  assign n5324 = ( ~n5316 & n5322 ) | ( ~n5316 & n5323 ) | ( n5322 & n5323 ) ;
  assign n5325 = x5 & x41 ;
  assign n5326 = x15 & x31 ;
  assign n5327 = n5325 | n5326 ;
  assign n5328 = x31 & x41 ;
  assign n5329 = n1005 & n5328 ;
  assign n5330 = n5327 | n5329 ;
  assign n5331 = x2 & x44 ;
  assign n5332 = ( ~n5329 & n5330 ) | ( ~n5329 & n5331 ) | ( n5330 & n5331 ) ;
  assign n5333 = ( n5329 & n5330 ) | ( n5329 & ~n5331 ) | ( n5330 & ~n5331 ) ;
  assign n5334 = ( ~n5330 & n5332 ) | ( ~n5330 & n5333 ) | ( n5332 & n5333 ) ;
  assign n5335 = n5324 & n5334 ;
  assign n5336 = n5324 & ~n5335 ;
  assign n5337 = ~n5324 & n5334 ;
  assign n5338 = n4938 | n5186 ;
  assign n5339 = ( n5186 & n5187 ) | ( n5186 & n5338 ) | ( n5187 & n5338 ) ;
  assign n5340 = n5337 | n5339 ;
  assign n5341 = n5336 | n5340 ;
  assign n5342 = n5337 & n5339 ;
  assign n5343 = ( n5336 & n5339 ) | ( n5336 & n5342 ) | ( n5339 & n5342 ) ;
  assign n5344 = n5341 & ~n5343 ;
  assign n5345 = n5076 | n5241 ;
  assign n5346 = n5076 & n5241 ;
  assign n5347 = n5345 & ~n5346 ;
  assign n5348 = n5230 | n5347 ;
  assign n5349 = n5230 & n5347 ;
  assign n5350 = n5348 & ~n5349 ;
  assign n5351 = n5172 | n5175 ;
  assign n5352 = ( n5172 & n5173 ) | ( n5172 & n5351 ) | ( n5173 & n5351 ) ;
  assign n5353 = n5350 | n5352 ;
  assign n5354 = n5350 & n5352 ;
  assign n5355 = n5353 & ~n5354 ;
  assign n5356 = n5344 & n5355 ;
  assign n5357 = n5344 | n5355 ;
  assign n5358 = ~n5356 & n5357 ;
  assign n5359 = n5313 & n5358 ;
  assign n5360 = n5313 | n5358 ;
  assign n5361 = ~n5359 & n5360 ;
  assign n5362 = ( n5161 & n5163 ) | ( n5161 & n5206 ) | ( n5163 & n5206 ) ;
  assign n5363 = n5361 & n5362 ;
  assign n5364 = n5361 | n5362 ;
  assign n5365 = ~n5363 & n5364 ;
  assign n5366 = n5307 | n5365 ;
  assign n5367 = n5307 & n5365 ;
  assign n5368 = n5366 & ~n5367 ;
  assign n5369 = ( n5190 & n5191 ) | ( n5190 & n5197 ) | ( n5191 & n5197 ) ;
  assign n5370 = n5258 | n5266 ;
  assign n5371 = n1018 & n3280 ;
  assign n5372 = n1023 & n2709 ;
  assign n5373 = n5371 | n5372 ;
  assign n5374 = n1020 & n2369 ;
  assign n5375 = x30 & n5374 ;
  assign n5376 = ( x30 & ~n5373 ) | ( x30 & n5375 ) | ( ~n5373 & n5375 ) ;
  assign n5377 = x16 & n5376 ;
  assign n5378 = n5373 | n5374 ;
  assign n5379 = x17 & x29 ;
  assign n5380 = x18 & x28 ;
  assign n5381 = ( ~n5374 & n5379 ) | ( ~n5374 & n5380 ) | ( n5379 & n5380 ) ;
  assign n5382 = n5379 & n5380 ;
  assign n5383 = ( ~n5373 & n5381 ) | ( ~n5373 & n5382 ) | ( n5381 & n5382 ) ;
  assign n5384 = ~n5378 & n5383 ;
  assign n5385 = n5377 | n5384 ;
  assign n5386 = ~n5370 & n5385 ;
  assign n5387 = n5370 & ~n5385 ;
  assign n5388 = n5386 | n5387 ;
  assign n5389 = x7 & x39 ;
  assign n5390 = x8 & x38 ;
  assign n5391 = n5389 | n5390 ;
  assign n5392 = x38 & x39 ;
  assign n5393 = n251 & n5392 ;
  assign n5394 = n3690 & ~n5393 ;
  assign n5395 = n5391 | n5393 ;
  assign n5396 = ( n5393 & n5394 ) | ( n5393 & n5395 ) | ( n5394 & n5395 ) ;
  assign n5397 = n5391 & ~n5396 ;
  assign n5398 = n3690 & ~n5391 ;
  assign n5399 = ( n3690 & ~n5394 ) | ( n3690 & n5398 ) | ( ~n5394 & n5398 ) ;
  assign n5400 = n5397 | n5399 ;
  assign n5401 = n5388 & n5400 ;
  assign n5402 = n5388 | n5400 ;
  assign n5403 = ~n5401 & n5402 ;
  assign n5404 = x0 & x46 ;
  assign n5405 = x4 & x42 ;
  assign n5406 = n5404 & n5405 ;
  assign n5407 = x42 & x43 ;
  assign n5408 = n79 & n5407 ;
  assign n5409 = x3 & x46 ;
  assign n5410 = n4671 & n5409 ;
  assign n5411 = n5408 | n5410 ;
  assign n5412 = x43 & n5406 ;
  assign n5413 = ( x43 & ~n5411 ) | ( x43 & n5412 ) | ( ~n5411 & n5412 ) ;
  assign n5414 = x3 & n5413 ;
  assign n5415 = ( n5404 & n5405 ) | ( n5404 & ~n5411 ) | ( n5405 & ~n5411 ) ;
  assign n5416 = ( ~n5406 & n5414 ) | ( ~n5406 & n5415 ) | ( n5414 & n5415 ) ;
  assign n5417 = x35 & x37 ;
  assign n5418 = n969 & n5417 ;
  assign n5419 = n360 & n3770 ;
  assign n5420 = n5418 | n5419 ;
  assign n5421 = n618 & n4078 ;
  assign n5422 = x37 & n5421 ;
  assign n5423 = ( x37 & ~n5420 ) | ( x37 & n5422 ) | ( ~n5420 & n5422 ) ;
  assign n5424 = x9 & n5423 ;
  assign n5425 = n5420 | n5421 ;
  assign n5426 = x11 & x35 ;
  assign n5427 = ( n4720 & ~n5421 ) | ( n4720 & n5426 ) | ( ~n5421 & n5426 ) ;
  assign n5428 = n4720 & n5426 ;
  assign n5429 = ( ~n5420 & n5427 ) | ( ~n5420 & n5428 ) | ( n5427 & n5428 ) ;
  assign n5430 = ~n5425 & n5429 ;
  assign n5431 = n5424 | n5430 ;
  assign n5432 = n5416 & n5431 ;
  assign n5433 = n5416 & ~n5432 ;
  assign n5434 = n5431 & ~n5432 ;
  assign n5435 = n5433 | n5434 ;
  assign n5436 = n1432 & n2724 ;
  assign n5437 = n1437 & n2267 ;
  assign n5438 = n5436 | n5437 ;
  assign n5439 = n1434 & n2511 ;
  assign n5440 = x27 & n5439 ;
  assign n5441 = ( x27 & ~n5438 ) | ( x27 & n5440 ) | ( ~n5438 & n5440 ) ;
  assign n5442 = x19 & n5441 ;
  assign n5443 = n5438 | n5439 ;
  assign n5444 = x20 & x26 ;
  assign n5445 = x21 & x25 ;
  assign n5446 = ( ~n5439 & n5444 ) | ( ~n5439 & n5445 ) | ( n5444 & n5445 ) ;
  assign n5447 = n5444 & n5445 ;
  assign n5448 = ( ~n5438 & n5446 ) | ( ~n5438 & n5447 ) | ( n5446 & n5447 ) ;
  assign n5449 = ~n5443 & n5448 ;
  assign n5450 = n5442 | n5449 ;
  assign n5451 = ( n5403 & n5435 ) | ( n5403 & ~n5450 ) | ( n5435 & ~n5450 ) ;
  assign n5452 = ( n5403 & ~n5435 ) | ( n5403 & n5450 ) | ( ~n5435 & n5450 ) ;
  assign n5453 = ( ~n5403 & n5451 ) | ( ~n5403 & n5452 ) | ( n5451 & n5452 ) ;
  assign n5454 = n5369 | n5453 ;
  assign n5455 = n5369 & n5453 ;
  assign n5456 = n5454 & ~n5455 ;
  assign n5457 = n5274 | n5275 ;
  assign n5458 = n5016 | n5274 ;
  assign n5459 = ( n5020 & n5457 ) | ( n5020 & n5458 ) | ( n5457 & n5458 ) ;
  assign n5460 = n5456 & n5459 ;
  assign n5461 = ( n5016 & n5020 ) | ( n5016 & n5275 ) | ( n5020 & n5275 ) ;
  assign n5462 = n5456 & n5461 ;
  assign n5463 = ( n5280 & n5460 ) | ( n5280 & n5462 ) | ( n5460 & n5462 ) ;
  assign n5464 = n5456 | n5459 ;
  assign n5465 = n5456 | n5461 ;
  assign n5466 = ( n5280 & n5464 ) | ( n5280 & n5465 ) | ( n5464 & n5465 ) ;
  assign n5467 = ~n5463 & n5466 ;
  assign n5468 = n5135 | n5149 ;
  assign n5469 = n5083 | n5097 ;
  assign n5470 = ( n5083 & n5085 ) | ( n5083 & n5469 ) | ( n5085 & n5469 ) ;
  assign n5471 = n5468 | n5470 ;
  assign n5472 = n5468 & n5470 ;
  assign n5473 = n5471 & ~n5472 ;
  assign n5474 = n5252 | n5268 ;
  assign n5475 = ( n5252 & n5255 ) | ( n5252 & n5474 ) | ( n5255 & n5474 ) ;
  assign n5476 = n5473 | n5475 ;
  assign n5477 = n5473 & n5475 ;
  assign n5478 = n5476 & ~n5477 ;
  assign n5479 = n5088 | n5092 ;
  assign n5480 = n5112 | n5479 ;
  assign n5481 = n5112 & n5479 ;
  assign n5482 = n5480 & ~n5481 ;
  assign n5483 = n5127 | n5482 ;
  assign n5484 = n5127 & n5482 ;
  assign n5485 = n5483 & ~n5484 ;
  assign n5486 = x44 & n1397 ;
  assign n5487 = x1 & x45 ;
  assign n5488 = n2148 & n5487 ;
  assign n5489 = n2148 | n5487 ;
  assign n5490 = ~n5488 & n5489 ;
  assign n5491 = ~n5486 & n5490 ;
  assign n5492 = n5486 & ~n5490 ;
  assign n5493 = n5491 | n5492 ;
  assign n5494 = n5142 & n5493 ;
  assign n5495 = n5142 | n5493 ;
  assign n5496 = ~n5494 & n5495 ;
  assign n5497 = n4891 | n5211 ;
  assign n5498 = ( n5211 & n5212 ) | ( n5211 & n5497 ) | ( n5212 & n5497 ) ;
  assign n5499 = n5496 & n5498 ;
  assign n5500 = n5496 | n5498 ;
  assign n5501 = ~n5499 & n5500 ;
  assign n5502 = n5485 & n5501 ;
  assign n5503 = n5485 | n5501 ;
  assign n5504 = ~n5502 & n5503 ;
  assign n5505 = n5219 & n5504 ;
  assign n5506 = ( n5272 & n5504 ) | ( n5272 & n5505 ) | ( n5504 & n5505 ) ;
  assign n5507 = n5219 | n5504 ;
  assign n5508 = n5272 | n5507 ;
  assign n5509 = ~n5506 & n5508 ;
  assign n5510 = n5478 & n5509 ;
  assign n5511 = n5478 | n5509 ;
  assign n5512 = ~n5510 & n5511 ;
  assign n5513 = n5467 & n5512 ;
  assign n5514 = n5467 | n5512 ;
  assign n5515 = ~n5513 & n5514 ;
  assign n5516 = ( n5306 & n5368 ) | ( n5306 & ~n5515 ) | ( n5368 & ~n5515 ) ;
  assign n5517 = ( ~n5368 & n5515 ) | ( ~n5368 & n5516 ) | ( n5515 & n5516 ) ;
  assign n5518 = ( ~n5306 & n5516 ) | ( ~n5306 & n5517 ) | ( n5516 & n5517 ) ;
  assign n5519 = n5368 & n5515 ;
  assign n5520 = n5368 | n5515 ;
  assign n5521 = n5519 | n5520 ;
  assign n5522 = ( n5305 & n5519 ) | ( n5305 & n5521 ) | ( n5519 & n5521 ) ;
  assign n5523 = ( n5303 & n5519 ) | ( n5303 & n5521 ) | ( n5519 & n5521 ) ;
  assign n5524 = ( n4853 & n5522 ) | ( n4853 & n5523 ) | ( n5522 & n5523 ) ;
  assign n5525 = n5478 | n5506 ;
  assign n5526 = ( n5506 & n5509 ) | ( n5506 & n5525 ) | ( n5509 & n5525 ) ;
  assign n5527 = n5310 | n5358 ;
  assign n5528 = ( n5308 & n5358 ) | ( n5308 & n5527 ) | ( n5358 & n5527 ) ;
  assign n5529 = n5526 & n5528 ;
  assign n5530 = n5312 & n5526 ;
  assign n5531 = ( n5313 & n5529 ) | ( n5313 & n5530 ) | ( n5529 & n5530 ) ;
  assign n5532 = n5526 | n5528 ;
  assign n5533 = n5312 | n5526 ;
  assign n5534 = ( n5313 & n5532 ) | ( n5313 & n5533 ) | ( n5532 & n5533 ) ;
  assign n5535 = ~n5531 & n5534 ;
  assign n5536 = ~n5329 & n5331 ;
  assign n5537 = ( n5329 & n5330 ) | ( n5329 & n5536 ) | ( n5330 & n5536 ) ;
  assign n5538 = n5443 | n5537 ;
  assign n5539 = n5443 & n5537 ;
  assign n5540 = n5538 & ~n5539 ;
  assign n5541 = n5406 | n5411 ;
  assign n5542 = n5540 | n5541 ;
  assign n5543 = n5540 & n5541 ;
  assign n5544 = n5542 & ~n5543 ;
  assign n5545 = n5432 | n5450 ;
  assign n5546 = n5544 & n5545 ;
  assign n5547 = n5432 & n5544 ;
  assign n5548 = ( n5435 & n5546 ) | ( n5435 & n5547 ) | ( n5546 & n5547 ) ;
  assign n5549 = n5544 | n5545 ;
  assign n5550 = n5432 | n5544 ;
  assign n5551 = ( n5435 & n5549 ) | ( n5435 & n5550 ) | ( n5549 & n5550 ) ;
  assign n5552 = ~n5548 & n5551 ;
  assign n5553 = n5335 | n5343 ;
  assign n5554 = n5552 | n5553 ;
  assign n5555 = n5552 & n5553 ;
  assign n5556 = n5554 & ~n5555 ;
  assign n5557 = n5435 & n5450 ;
  assign n5558 = n5435 & ~n5557 ;
  assign n5559 = ~n5435 & n5450 ;
  assign n5560 = n5403 & n5559 ;
  assign n5561 = ( n5403 & n5558 ) | ( n5403 & n5560 ) | ( n5558 & n5560 ) ;
  assign n5562 = n5455 | n5561 ;
  assign n5563 = n5344 | n5354 ;
  assign n5564 = ( n5354 & n5355 ) | ( n5354 & n5563 ) | ( n5355 & n5563 ) ;
  assign n5565 = n5562 & n5564 ;
  assign n5566 = n5562 & ~n5565 ;
  assign n5567 = ~n5561 & n5564 ;
  assign n5568 = ~n5455 & n5556 ;
  assign n5569 = n5567 & n5568 ;
  assign n5570 = ( n5556 & n5566 ) | ( n5556 & n5569 ) | ( n5566 & n5569 ) ;
  assign n5571 = n5455 & ~n5556 ;
  assign n5572 = ( n5556 & n5567 ) | ( n5556 & ~n5571 ) | ( n5567 & ~n5571 ) ;
  assign n5573 = n5566 | n5572 ;
  assign n5574 = ~n5570 & n5573 ;
  assign n5575 = ~n5535 & n5574 ;
  assign n5576 = n5535 & ~n5574 ;
  assign n5577 = n5575 | n5576 ;
  assign n5578 = ( n5280 & n5459 ) | ( n5280 & n5461 ) | ( n5459 & n5461 ) ;
  assign n5579 = n5456 | n5512 ;
  assign n5580 = ( n5512 & n5578 ) | ( n5512 & n5579 ) | ( n5578 & n5579 ) ;
  assign n5581 = ( n5463 & n5467 ) | ( n5463 & n5580 ) | ( n5467 & n5580 ) ;
  assign n5582 = ( n5370 & n5385 ) | ( n5370 & n5400 ) | ( n5385 & n5400 ) ;
  assign n5583 = n5127 | n5481 ;
  assign n5584 = ( n5481 & n5482 ) | ( n5481 & n5583 ) | ( n5482 & n5583 ) ;
  assign n5585 = n5582 | n5584 ;
  assign n5586 = n5582 & n5584 ;
  assign n5587 = n5585 & ~n5586 ;
  assign n5588 = x1 & x46 ;
  assign n5589 = x24 | n5588 ;
  assign n5590 = x24 & x46 ;
  assign n5591 = x1 & n5590 ;
  assign n5592 = n5421 & ~n5591 ;
  assign n5593 = ( n5420 & ~n5591 ) | ( n5420 & n5592 ) | ( ~n5591 & n5592 ) ;
  assign n5594 = n5589 & n5593 ;
  assign n5595 = n5425 & ~n5594 ;
  assign n5596 = n5589 & ~n5591 ;
  assign n5597 = ~n5593 & n5596 ;
  assign n5598 = n5396 & n5597 ;
  assign n5599 = ( n5396 & n5595 ) | ( n5396 & n5598 ) | ( n5595 & n5598 ) ;
  assign n5600 = n5396 | n5597 ;
  assign n5601 = n5595 | n5600 ;
  assign n5602 = ~n5599 & n5601 ;
  assign n5603 = ~n5587 & n5602 ;
  assign n5604 = n5586 | n5602 ;
  assign n5605 = n5585 & ~n5604 ;
  assign n5606 = n5603 | n5605 ;
  assign n5607 = x0 & x47 ;
  assign n5608 = x2 & x45 ;
  assign n5609 = n5607 | n5608 ;
  assign n5610 = x45 & x47 ;
  assign n5611 = n67 & n5610 ;
  assign n5612 = n5609 & ~n5611 ;
  assign n5613 = n5488 | n5611 ;
  assign n5614 = ( n5611 & n5612 ) | ( n5611 & n5613 ) | ( n5612 & n5613 ) ;
  assign n5615 = n5609 & ~n5614 ;
  assign n5616 = n5488 & ~n5612 ;
  assign n5617 = n5615 | n5616 ;
  assign n5618 = n1018 & n3595 ;
  assign n5619 = n1023 & n2965 ;
  assign n5620 = n5618 | n5619 ;
  assign n5621 = n1020 & n2709 ;
  assign n5622 = x31 & n5621 ;
  assign n5623 = ( x31 & ~n5620 ) | ( x31 & n5622 ) | ( ~n5620 & n5622 ) ;
  assign n5624 = x16 & n5623 ;
  assign n5625 = n5620 | n5621 ;
  assign n5626 = x17 & x30 ;
  assign n5627 = x18 & x29 ;
  assign n5628 = ( ~n5621 & n5626 ) | ( ~n5621 & n5627 ) | ( n5626 & n5627 ) ;
  assign n5629 = n5626 & n5627 ;
  assign n5630 = ( ~n5620 & n5628 ) | ( ~n5620 & n5629 ) | ( n5628 & n5629 ) ;
  assign n5631 = ~n5625 & n5630 ;
  assign n5632 = n5624 | n5631 ;
  assign n5633 = n5617 & n5632 ;
  assign n5634 = n5617 & ~n5633 ;
  assign n5635 = n5632 & ~n5633 ;
  assign n5636 = n5634 | n5635 ;
  assign n5637 = n1432 & n2895 ;
  assign n5638 = n1437 & n2372 ;
  assign n5639 = n5637 | n5638 ;
  assign n5640 = n1434 & n2267 ;
  assign n5641 = x28 & n5640 ;
  assign n5642 = ( x28 & ~n5639 ) | ( x28 & n5641 ) | ( ~n5639 & n5641 ) ;
  assign n5643 = x19 & n5642 ;
  assign n5644 = n5639 | n5640 ;
  assign n5645 = x20 & x27 ;
  assign n5646 = ( n2132 & ~n5640 ) | ( n2132 & n5645 ) | ( ~n5640 & n5645 ) ;
  assign n5647 = n2132 & n5645 ;
  assign n5648 = ( ~n5639 & n5646 ) | ( ~n5639 & n5647 ) | ( n5646 & n5647 ) ;
  assign n5649 = ~n5644 & n5648 ;
  assign n5650 = n5643 | n5649 ;
  assign n5651 = ~n5636 & n5650 ;
  assign n5652 = n5636 & ~n5650 ;
  assign n5653 = n5651 | n5652 ;
  assign n5654 = n5316 | n5319 ;
  assign n5655 = n5378 | n5654 ;
  assign n5656 = n5378 & n5654 ;
  assign n5657 = n5655 & ~n5656 ;
  assign n5658 = x43 & x44 ;
  assign n5659 = n79 & n5658 ;
  assign n5660 = x15 & x44 ;
  assign n5661 = n3141 & n5660 ;
  assign n5662 = n5659 | n5661 ;
  assign n5663 = x32 & x43 ;
  assign n5664 = n921 & n5663 ;
  assign n5665 = x44 & n5664 ;
  assign n5666 = ( x44 & ~n5662 ) | ( x44 & n5665 ) | ( ~n5662 & n5665 ) ;
  assign n5667 = x3 & n5666 ;
  assign n5668 = n5662 | n5664 ;
  assign n5669 = x15 & x32 ;
  assign n5670 = ( n4675 & ~n5664 ) | ( n4675 & n5669 ) | ( ~n5664 & n5669 ) ;
  assign n5671 = n4675 & n5669 ;
  assign n5672 = ( ~n5662 & n5670 ) | ( ~n5662 & n5671 ) | ( n5670 & n5671 ) ;
  assign n5673 = ~n5668 & n5672 ;
  assign n5674 = n5667 | n5673 ;
  assign n5675 = n5657 & n5674 ;
  assign n5676 = n5657 & ~n5675 ;
  assign n5677 = n5674 & ~n5675 ;
  assign n5678 = n5676 | n5677 ;
  assign n5679 = n313 & n5392 ;
  assign n5680 = x11 & x39 ;
  assign n5681 = n4913 & n5680 ;
  assign n5682 = n5679 | n5681 ;
  assign n5683 = n969 & n3731 ;
  assign n5684 = x39 & n5683 ;
  assign n5685 = ( x39 & ~n5682 ) | ( x39 & n5684 ) | ( ~n5682 & n5684 ) ;
  assign n5686 = x8 & n5685 ;
  assign n5687 = n5682 | n5683 ;
  assign n5688 = x9 & x38 ;
  assign n5689 = x11 & x36 ;
  assign n5690 = ( ~n5683 & n5688 ) | ( ~n5683 & n5689 ) | ( n5688 & n5689 ) ;
  assign n5691 = n5688 & n5689 ;
  assign n5692 = ( ~n5682 & n5690 ) | ( ~n5682 & n5691 ) | ( n5690 & n5691 ) ;
  assign n5693 = ~n5687 & n5692 ;
  assign n5694 = n5686 | n5693 ;
  assign n5695 = x22 & x25 ;
  assign n5696 = n1686 | n5695 ;
  assign n5697 = n1912 & n1932 ;
  assign n5698 = x10 & x37 ;
  assign n5699 = ~n5697 & n5698 ;
  assign n5700 = n5696 | n5697 ;
  assign n5701 = ( n5697 & n5699 ) | ( n5697 & n5700 ) | ( n5699 & n5700 ) ;
  assign n5702 = n5696 & ~n5701 ;
  assign n5703 = ( ~n5696 & n5697 ) | ( ~n5696 & n5698 ) | ( n5697 & n5698 ) ;
  assign n5704 = n5698 & n5703 ;
  assign n5705 = n5702 | n5704 ;
  assign n5706 = n5694 & n5705 ;
  assign n5707 = n5694 & ~n5706 ;
  assign n5708 = n5705 & ~n5706 ;
  assign n5709 = n5707 | n5708 ;
  assign n5710 = x41 & x42 ;
  assign n5711 = n204 & n5710 ;
  assign n5712 = x14 & x42 ;
  assign n5713 = n3627 & n5712 ;
  assign n5714 = n5711 | n5713 ;
  assign n5715 = x33 & x41 ;
  assign n5716 = n1006 & n5715 ;
  assign n5717 = x42 & n5716 ;
  assign n5718 = ( x42 & ~n5714 ) | ( x42 & n5717 ) | ( ~n5714 & n5717 ) ;
  assign n5719 = x5 & n5718 ;
  assign n5720 = n5714 | n5716 ;
  assign n5721 = x6 & x41 ;
  assign n5722 = x14 & x33 ;
  assign n5723 = ( ~n5716 & n5721 ) | ( ~n5716 & n5722 ) | ( n5721 & n5722 ) ;
  assign n5724 = n5721 & n5722 ;
  assign n5725 = ( ~n5714 & n5723 ) | ( ~n5714 & n5724 ) | ( n5723 & n5724 ) ;
  assign n5726 = ~n5720 & n5725 ;
  assign n5727 = n5719 | n5726 ;
  assign n5728 = ( n5678 & n5709 ) | ( n5678 & ~n5727 ) | ( n5709 & ~n5727 ) ;
  assign n5729 = ( ~n5709 & n5727 ) | ( ~n5709 & n5728 ) | ( n5727 & n5728 ) ;
  assign n5730 = ( ~n5678 & n5728 ) | ( ~n5678 & n5729 ) | ( n5728 & n5729 ) ;
  assign n5731 = n5653 & n5730 ;
  assign n5732 = n5653 | n5730 ;
  assign n5733 = ~n5731 & n5732 ;
  assign n5734 = n5606 & ~n5733 ;
  assign n5735 = n647 & n3483 ;
  assign n5736 = x34 & x40 ;
  assign n5737 = n986 & n5736 ;
  assign n5738 = n5735 | n5737 ;
  assign n5739 = x12 & x40 ;
  assign n5740 = n4513 & n5739 ;
  assign n5741 = x34 & n5740 ;
  assign n5742 = ( x34 & ~n5738 ) | ( x34 & n5741 ) | ( ~n5738 & n5741 ) ;
  assign n5743 = x13 & n5742 ;
  assign n5744 = n5738 | n5740 ;
  assign n5745 = x7 & x40 ;
  assign n5746 = x12 & x35 ;
  assign n5747 = ( ~n5740 & n5745 ) | ( ~n5740 & n5746 ) | ( n5745 & n5746 ) ;
  assign n5748 = n5745 & n5746 ;
  assign n5749 = ( ~n5738 & n5747 ) | ( ~n5738 & n5748 ) | ( n5747 & n5748 ) ;
  assign n5750 = ~n5744 & n5749 ;
  assign n5751 = n5743 | n5750 ;
  assign n5752 = ( n5142 & n5486 ) | ( n5142 & n5490 ) | ( n5486 & n5490 ) ;
  assign n5753 = n5751 & n5752 ;
  assign n5754 = n5751 & ~n5753 ;
  assign n5755 = ~n5751 & n5752 ;
  assign n5756 = n5230 | n5346 ;
  assign n5757 = ( n5346 & n5347 ) | ( n5346 & n5756 ) | ( n5347 & n5756 ) ;
  assign n5758 = n5755 | n5757 ;
  assign n5759 = n5754 | n5758 ;
  assign n5760 = n5755 & n5757 ;
  assign n5761 = ( n5754 & n5757 ) | ( n5754 & n5760 ) | ( n5757 & n5760 ) ;
  assign n5762 = n5759 & ~n5761 ;
  assign n5763 = n5485 | n5499 ;
  assign n5764 = ( n5499 & n5501 ) | ( n5499 & n5763 ) | ( n5501 & n5763 ) ;
  assign n5765 = n5762 | n5764 ;
  assign n5766 = n5762 & n5764 ;
  assign n5767 = n5765 & ~n5766 ;
  assign n5768 = n5472 | n5475 ;
  assign n5769 = ( n5472 & n5473 ) | ( n5472 & n5768 ) | ( n5473 & n5768 ) ;
  assign n5770 = n5767 | n5769 ;
  assign n5771 = n5767 & n5769 ;
  assign n5772 = n5770 & ~n5771 ;
  assign n5773 = ( n5733 & n5734 ) | ( n5733 & n5772 ) | ( n5734 & n5772 ) ;
  assign n5774 = ( ~n5606 & n5734 ) | ( ~n5606 & n5773 ) | ( n5734 & n5773 ) ;
  assign n5775 = n5606 & n5733 ;
  assign n5776 = n5733 & ~n5775 ;
  assign n5777 = n5734 | n5772 ;
  assign n5778 = n5776 | n5777 ;
  assign n5779 = ~n5774 & n5778 ;
  assign n5780 = n5580 & n5779 ;
  assign n5781 = n5463 & n5779 ;
  assign n5782 = ( n5467 & n5780 ) | ( n5467 & n5781 ) | ( n5780 & n5781 ) ;
  assign n5783 = n5581 & ~n5782 ;
  assign n5784 = ~n5580 & n5779 ;
  assign n5785 = ~n5463 & n5779 ;
  assign n5786 = ( ~n5467 & n5784 ) | ( ~n5467 & n5785 ) | ( n5784 & n5785 ) ;
  assign n5787 = n5783 | n5786 ;
  assign n5788 = n5577 & n5787 ;
  assign n5789 = ( ~n5577 & n5783 ) | ( ~n5577 & n5786 ) | ( n5783 & n5786 ) ;
  assign n5790 = n5577 | n5789 ;
  assign n5791 = ~n5788 & n5790 ;
  assign n5792 = n5363 | n5365 ;
  assign n5793 = ( n5307 & n5363 ) | ( n5307 & n5792 ) | ( n5363 & n5792 ) ;
  assign n5794 = ( n5524 & n5791 ) | ( n5524 & ~n5793 ) | ( n5791 & ~n5793 ) ;
  assign n5795 = ( ~n5791 & n5793 ) | ( ~n5791 & n5794 ) | ( n5793 & n5794 ) ;
  assign n5796 = ( ~n5524 & n5794 ) | ( ~n5524 & n5795 ) | ( n5794 & n5795 ) ;
  assign n5797 = x9 & x39 ;
  assign n5798 = x37 & x39 ;
  assign n5799 = n969 & n5798 ;
  assign n5800 = n360 & n5392 ;
  assign n5801 = n5799 | n5800 ;
  assign n5802 = n618 & n4857 ;
  assign n5803 = n5797 & n5802 ;
  assign n5804 = ( n5797 & ~n5801 ) | ( n5797 & n5803 ) | ( ~n5801 & n5803 ) ;
  assign n5805 = n5801 | n5802 ;
  assign n5806 = x10 & x38 ;
  assign n5807 = ( n4860 & ~n5802 ) | ( n4860 & n5806 ) | ( ~n5802 & n5806 ) ;
  assign n5808 = n4860 & n5806 ;
  assign n5809 = ( ~n5801 & n5807 ) | ( ~n5801 & n5808 ) | ( n5807 & n5808 ) ;
  assign n5810 = ~n5805 & n5809 ;
  assign n5811 = n5804 | n5810 ;
  assign n5812 = x7 & x41 ;
  assign n5813 = x40 & x41 ;
  assign n5814 = n251 & n5813 ;
  assign n5815 = n4080 & n5812 ;
  assign n5816 = n5814 | n5815 ;
  assign n5817 = n4913 & n5739 ;
  assign n5818 = n5812 & n5817 ;
  assign n5819 = ( n5812 & ~n5816 ) | ( n5812 & n5818 ) | ( ~n5816 & n5818 ) ;
  assign n5820 = n5816 | n5817 ;
  assign n5821 = x8 & x40 ;
  assign n5822 = ( n4080 & ~n5817 ) | ( n4080 & n5821 ) | ( ~n5817 & n5821 ) ;
  assign n5823 = n4080 & n5821 ;
  assign n5824 = ( ~n5816 & n5822 ) | ( ~n5816 & n5823 ) | ( n5822 & n5823 ) ;
  assign n5825 = ~n5820 & n5824 ;
  assign n5826 = n5819 | n5825 ;
  assign n5827 = x6 & x42 ;
  assign n5828 = x13 & x35 ;
  assign n5829 = n5827 & n5828 ;
  assign n5830 = n650 & n3483 ;
  assign n5831 = n4127 & n5712 ;
  assign n5832 = n5830 | n5831 ;
  assign n5833 = x34 & n5829 ;
  assign n5834 = ( x34 & ~n5832 ) | ( x34 & n5833 ) | ( ~n5832 & n5833 ) ;
  assign n5835 = x14 & n5834 ;
  assign n5836 = ( n5827 & n5828 ) | ( n5827 & ~n5832 ) | ( n5828 & ~n5832 ) ;
  assign n5837 = ( ~n5829 & n5835 ) | ( ~n5829 & n5836 ) | ( n5835 & n5836 ) ;
  assign n5838 = ( n5811 & ~n5826 ) | ( n5811 & n5837 ) | ( ~n5826 & n5837 ) ;
  assign n5839 = ( n5826 & ~n5837 ) | ( n5826 & n5838 ) | ( ~n5837 & n5838 ) ;
  assign n5840 = ( ~n5811 & n5838 ) | ( ~n5811 & n5839 ) | ( n5838 & n5839 ) ;
  assign n5841 = n5753 | n5761 ;
  assign n5842 = n5840 | n5841 ;
  assign n5843 = n5840 & n5841 ;
  assign n5844 = n5842 & ~n5843 ;
  assign n5845 = x33 & x44 ;
  assign n5846 = n921 & n5845 ;
  assign n5847 = n91 & n5658 ;
  assign n5848 = n5846 | n5847 ;
  assign n5849 = x33 & x43 ;
  assign n5850 = n1005 & n5849 ;
  assign n5851 = x44 & n5850 ;
  assign n5852 = ( x44 & ~n5848 ) | ( x44 & n5851 ) | ( ~n5848 & n5851 ) ;
  assign n5853 = x4 & n5852 ;
  assign n5854 = n5848 | n5850 ;
  assign n5855 = x5 & x43 ;
  assign n5856 = x15 & x33 ;
  assign n5857 = ( ~n5850 & n5855 ) | ( ~n5850 & n5856 ) | ( n5855 & n5856 ) ;
  assign n5858 = n5855 & n5856 ;
  assign n5859 = ( ~n5848 & n5857 ) | ( ~n5848 & n5858 ) | ( n5857 & n5858 ) ;
  assign n5860 = ~n5854 & n5859 ;
  assign n5861 = n5853 | n5860 ;
  assign n5862 = n1710 & n2895 ;
  assign n5863 = n1434 & n2372 ;
  assign n5864 = n5862 | n5863 ;
  assign n5865 = n1585 & n2267 ;
  assign n5866 = x28 & n5865 ;
  assign n5867 = ( x28 & ~n5864 ) | ( x28 & n5866 ) | ( ~n5864 & n5866 ) ;
  assign n5868 = x20 & n5867 ;
  assign n5869 = n5864 | n5865 ;
  assign n5870 = x21 & x27 ;
  assign n5871 = x22 & x26 ;
  assign n5872 = ( ~n5865 & n5870 ) | ( ~n5865 & n5871 ) | ( n5870 & n5871 ) ;
  assign n5873 = n5870 & n5871 ;
  assign n5874 = ( ~n5864 & n5872 ) | ( ~n5864 & n5873 ) | ( n5872 & n5873 ) ;
  assign n5875 = ~n5869 & n5874 ;
  assign n5876 = n5868 | n5875 ;
  assign n5877 = n5861 & n5876 ;
  assign n5878 = n5861 & ~n5877 ;
  assign n5879 = n5876 & ~n5877 ;
  assign n5880 = n5878 | n5879 ;
  assign n5881 = n3334 & n3595 ;
  assign n5882 = n1020 & n2965 ;
  assign n5883 = n5881 | n5882 ;
  assign n5884 = n1077 & n2709 ;
  assign n5885 = x31 & n5884 ;
  assign n5886 = ( x31 & ~n5883 ) | ( x31 & n5885 ) | ( ~n5883 & n5885 ) ;
  assign n5887 = x17 & n5886 ;
  assign n5888 = n5883 | n5884 ;
  assign n5889 = x18 & x30 ;
  assign n5890 = x19 & x29 ;
  assign n5891 = ( ~n5884 & n5889 ) | ( ~n5884 & n5890 ) | ( n5889 & n5890 ) ;
  assign n5892 = n5889 & n5890 ;
  assign n5893 = ( ~n5883 & n5891 ) | ( ~n5883 & n5892 ) | ( n5891 & n5892 ) ;
  assign n5894 = ~n5888 & n5893 ;
  assign n5895 = n5887 | n5894 ;
  assign n5896 = ~n5880 & n5895 ;
  assign n5897 = n5880 & ~n5895 ;
  assign n5898 = n5896 | n5897 ;
  assign n5899 = n5844 | n5898 ;
  assign n5900 = n5844 & n5898 ;
  assign n5901 = n5899 & ~n5900 ;
  assign n5902 = n5766 | n5767 ;
  assign n5903 = ( n5766 & n5769 ) | ( n5766 & n5902 ) | ( n5769 & n5902 ) ;
  assign n5904 = n5901 & n5903 ;
  assign n5905 = n5901 | n5903 ;
  assign n5906 = ~n5904 & n5905 ;
  assign n5907 = n5565 & n5906 ;
  assign n5908 = ( n5570 & n5906 ) | ( n5570 & n5907 ) | ( n5906 & n5907 ) ;
  assign n5909 = n5565 | n5906 ;
  assign n5910 = n5570 | n5909 ;
  assign n5911 = ~n5908 & n5910 ;
  assign n5912 = n5531 | n5574 ;
  assign n5913 = ( n5531 & n5535 ) | ( n5531 & n5912 ) | ( n5535 & n5912 ) ;
  assign n5914 = n5911 | n5913 ;
  assign n5915 = n5911 & n5913 ;
  assign n5916 = n5914 & ~n5915 ;
  assign n5917 = ( n5586 & n5587 ) | ( n5586 & n5604 ) | ( n5587 & n5604 ) ;
  assign n5918 = n5548 | n5553 ;
  assign n5919 = ( n5548 & n5552 ) | ( n5548 & n5918 ) | ( n5552 & n5918 ) ;
  assign n5920 = n5917 | n5919 ;
  assign n5921 = n5917 & n5919 ;
  assign n5922 = n5920 & ~n5921 ;
  assign n5923 = x0 & x48 ;
  assign n5924 = n5591 & n5923 ;
  assign n5925 = n5591 & ~n5924 ;
  assign n5926 = ~n5591 & n5923 ;
  assign n5927 = n5925 | n5926 ;
  assign n5928 = x1 & x47 ;
  assign n5929 = n1557 & n5928 ;
  assign n5930 = n5928 & ~n5929 ;
  assign n5931 = n1557 & ~n5929 ;
  assign n5932 = n5930 | n5931 ;
  assign n5933 = ~n5927 & n5932 ;
  assign n5934 = n5927 & ~n5932 ;
  assign n5935 = n5933 | n5934 ;
  assign n5936 = n5539 | n5541 ;
  assign n5937 = ( n5539 & n5540 ) | ( n5539 & n5936 ) | ( n5540 & n5936 ) ;
  assign n5938 = n5935 | n5937 ;
  assign n5939 = n5935 & n5937 ;
  assign n5940 = n5938 & ~n5939 ;
  assign n5941 = n5656 | n5675 ;
  assign n5942 = n5940 | n5941 ;
  assign n5943 = n5940 & n5941 ;
  assign n5944 = n5942 & ~n5943 ;
  assign n5945 = n5922 & n5944 ;
  assign n5946 = n5922 | n5944 ;
  assign n5947 = ~n5945 & n5946 ;
  assign n5948 = n5775 & n5947 ;
  assign n5949 = ( n5774 & n5947 ) | ( n5774 & n5948 ) | ( n5947 & n5948 ) ;
  assign n5950 = n5734 | n5775 ;
  assign n5951 = ( ~n5734 & n5773 ) | ( ~n5734 & n5950 ) | ( n5773 & n5950 ) ;
  assign n5952 = ~n5949 & n5951 ;
  assign n5953 = n5644 | n5687 ;
  assign n5954 = n5644 & n5687 ;
  assign n5955 = n5953 & ~n5954 ;
  assign n5956 = n5720 | n5955 ;
  assign n5957 = n5720 & n5955 ;
  assign n5958 = n5956 & ~n5957 ;
  assign n5959 = n5706 | n5727 ;
  assign n5960 = n5958 & n5959 ;
  assign n5961 = n5706 & n5958 ;
  assign n5962 = ( n5709 & n5960 ) | ( n5709 & n5961 ) | ( n5960 & n5961 ) ;
  assign n5963 = n5958 | n5959 ;
  assign n5964 = n5706 | n5958 ;
  assign n5965 = ( n5709 & n5963 ) | ( n5709 & n5964 ) | ( n5963 & n5964 ) ;
  assign n5966 = ~n5962 & n5965 ;
  assign n5967 = n5701 | n5744 ;
  assign n5968 = n5701 & n5744 ;
  assign n5969 = n5967 & ~n5968 ;
  assign n5970 = x3 & x45 ;
  assign n5971 = x16 & x32 ;
  assign n5972 = n5970 & n5971 ;
  assign n5973 = x32 & x46 ;
  assign n5974 = n801 & n5973 ;
  assign n5975 = x45 & x46 ;
  assign n5976 = n77 & n5975 ;
  assign n5977 = n5974 | n5976 ;
  assign n5978 = x46 & n5972 ;
  assign n5979 = ( x46 & ~n5977 ) | ( x46 & n5978 ) | ( ~n5977 & n5978 ) ;
  assign n5980 = x2 & n5979 ;
  assign n5981 = ( n5970 & n5971 ) | ( n5970 & ~n5977 ) | ( n5971 & ~n5977 ) ;
  assign n5982 = ( ~n5972 & n5980 ) | ( ~n5972 & n5981 ) | ( n5980 & n5981 ) ;
  assign n5983 = n5969 & n5982 ;
  assign n5984 = n5969 & ~n5983 ;
  assign n5985 = n5982 & ~n5983 ;
  assign n5986 = n5984 | n5985 ;
  assign n5987 = n5966 | n5986 ;
  assign n5988 = n5966 & n5986 ;
  assign n5989 = n5987 & ~n5988 ;
  assign n5990 = n5709 & n5727 ;
  assign n5991 = n5709 & ~n5990 ;
  assign n5992 = ~n5709 & n5727 ;
  assign n5993 = n5678 & n5992 ;
  assign n5994 = ( n5678 & n5991 ) | ( n5678 & n5993 ) | ( n5991 & n5993 ) ;
  assign n5995 = n5731 | n5994 ;
  assign n5996 = n5989 & n5995 ;
  assign n5997 = n5989 | n5995 ;
  assign n5998 = ~n5996 & n5997 ;
  assign n5999 = n5625 | n5668 ;
  assign n6000 = n5625 & n5668 ;
  assign n6001 = n5999 & ~n6000 ;
  assign n6002 = n5614 | n6001 ;
  assign n6003 = n5614 & n6001 ;
  assign n6004 = n6002 & ~n6003 ;
  assign n6005 = n5594 | n5599 ;
  assign n6006 = n5633 | n5650 ;
  assign n6007 = n6005 & n6006 ;
  assign n6008 = n5633 & n6005 ;
  assign n6009 = ( n5636 & n6007 ) | ( n5636 & n6008 ) | ( n6007 & n6008 ) ;
  assign n6010 = n6005 | n6006 ;
  assign n6011 = n5633 | n6005 ;
  assign n6012 = ( n5636 & n6010 ) | ( n5636 & n6011 ) | ( n6010 & n6011 ) ;
  assign n6013 = ~n6009 & n6012 ;
  assign n6014 = n6004 & n6013 ;
  assign n6015 = n6004 | n6013 ;
  assign n6016 = ~n6014 & n6015 ;
  assign n6017 = n5998 & n6016 ;
  assign n6018 = n5998 | n6016 ;
  assign n6019 = ~n6017 & n6018 ;
  assign n6020 = n5947 & ~n5948 ;
  assign n6021 = ~n5774 & n6020 ;
  assign n6022 = n6019 | n6021 ;
  assign n6023 = n5952 | n6022 ;
  assign n6024 = n6019 & n6021 ;
  assign n6025 = ( n5952 & n6019 ) | ( n5952 & n6024 ) | ( n6019 & n6024 ) ;
  assign n6026 = n6023 & ~n6025 ;
  assign n6027 = n5916 & n6026 ;
  assign n6028 = n5916 | n6026 ;
  assign n6029 = ~n6027 & n6028 ;
  assign n6030 = n5577 | n5782 ;
  assign n6031 = ( n5782 & n5787 ) | ( n5782 & n6030 ) | ( n5787 & n6030 ) ;
  assign n6032 = n6029 | n6031 ;
  assign n6033 = n6029 & n6031 ;
  assign n6034 = n6032 & ~n6033 ;
  assign n6035 = n5791 & n5793 ;
  assign n6036 = n5791 | n5793 ;
  assign n6037 = n6035 | n6036 ;
  assign n6038 = ( n5524 & n6035 ) | ( n5524 & n6037 ) | ( n6035 & n6037 ) ;
  assign n6039 = n6034 | n6038 ;
  assign n6040 = n6032 & n6038 ;
  assign n6041 = ~n6033 & n6040 ;
  assign n6042 = n6039 & ~n6041 ;
  assign n6043 = n6032 & n6035 ;
  assign n6044 = n6033 | n6043 ;
  assign n6045 = n6032 | n6033 ;
  assign n6046 = ( n6033 & n6037 ) | ( n6033 & n6045 ) | ( n6037 & n6045 ) ;
  assign n6047 = ( n5524 & n6044 ) | ( n5524 & n6046 ) | ( n6044 & n6046 ) ;
  assign n6048 = x7 & x42 ;
  assign n6049 = x8 & x41 ;
  assign n6050 = n6048 | n6049 ;
  assign n6051 = n251 & n5710 ;
  assign n6052 = n6050 | n6051 ;
  assign n6053 = x13 & x36 ;
  assign n6054 = ( ~n6051 & n6052 ) | ( ~n6051 & n6053 ) | ( n6052 & n6053 ) ;
  assign n6055 = ( n6051 & n6052 ) | ( n6051 & ~n6053 ) | ( n6052 & ~n6053 ) ;
  assign n6056 = ( ~n6052 & n6054 ) | ( ~n6052 & n6055 ) | ( n6054 & n6055 ) ;
  assign n6057 = n1912 | n2336 ;
  assign n6058 = x11 & x38 ;
  assign n6059 = ( n1912 & n2336 ) | ( n1912 & n6058 ) | ( n2336 & n6058 ) ;
  assign n6060 = n6057 & ~n6059 ;
  assign n6061 = n1912 & n2336 ;
  assign n6062 = n6058 & ~n6061 ;
  assign n6063 = ~n6057 & n6058 ;
  assign n6064 = ( n6058 & ~n6062 ) | ( n6058 & n6063 ) | ( ~n6062 & n6063 ) ;
  assign n6065 = n6060 | n6064 ;
  assign n6066 = n6056 & n6065 ;
  assign n6067 = n6056 & ~n6066 ;
  assign n6068 = n6065 & ~n6066 ;
  assign n6069 = n6067 | n6068 ;
  assign n6070 = x15 & x43 ;
  assign n6071 = n4127 & n6070 ;
  assign n6072 = n792 & n3483 ;
  assign n6073 = n6071 | n6072 ;
  assign n6074 = x35 & x43 ;
  assign n6075 = n1006 & n6074 ;
  assign n6076 = x34 & n6075 ;
  assign n6077 = ( x34 & ~n6073 ) | ( x34 & n6076 ) | ( ~n6073 & n6076 ) ;
  assign n6078 = x15 & n6077 ;
  assign n6079 = n6073 | n6075 ;
  assign n6080 = x6 & x43 ;
  assign n6081 = x14 & x35 ;
  assign n6082 = ( ~n6075 & n6080 ) | ( ~n6075 & n6081 ) | ( n6080 & n6081 ) ;
  assign n6083 = n6080 & n6081 ;
  assign n6084 = ( ~n6073 & n6082 ) | ( ~n6073 & n6083 ) | ( n6082 & n6083 ) ;
  assign n6085 = ~n6079 & n6084 ;
  assign n6086 = n6078 | n6085 ;
  assign n6087 = ~n6069 & n6086 ;
  assign n6088 = n6069 & ~n6086 ;
  assign n6089 = n6087 | n6088 ;
  assign n6090 = x44 & n89 ;
  assign n6091 = x45 & n82 ;
  assign n6092 = n6090 | n6091 ;
  assign n6093 = x44 & x45 ;
  assign n6094 = n91 & n6093 ;
  assign n6095 = x49 & ~n6094 ;
  assign n6096 = n6092 & n6095 ;
  assign n6097 = x0 & x49 ;
  assign n6098 = ~n6096 & n6097 ;
  assign n6099 = n6094 | n6096 ;
  assign n6100 = x4 & x45 ;
  assign n6101 = x5 & x44 ;
  assign n6102 = ( ~n6094 & n6100 ) | ( ~n6094 & n6101 ) | ( n6100 & n6101 ) ;
  assign n6103 = n6100 & n6101 ;
  assign n6104 = ( ~n6096 & n6102 ) | ( ~n6096 & n6103 ) | ( n6102 & n6103 ) ;
  assign n6105 = ~n6099 & n6104 ;
  assign n6106 = n6098 | n6105 ;
  assign n6107 = n5924 | n5932 ;
  assign n6108 = ( n5924 & n5927 ) | ( n5924 & n6107 ) | ( n5927 & n6107 ) ;
  assign n6109 = n6106 & ~n6108 ;
  assign n6110 = ~n6106 & n6108 ;
  assign n6111 = n6109 | n6110 ;
  assign n6112 = n1018 & n2683 ;
  assign n6113 = n1023 & n3321 ;
  assign n6114 = n6112 | n6113 ;
  assign n6115 = n1020 & n4062 ;
  assign n6116 = x33 & n6115 ;
  assign n6117 = ( x33 & ~n6114 ) | ( x33 & n6116 ) | ( ~n6114 & n6116 ) ;
  assign n6118 = x16 & n6117 ;
  assign n6119 = n6114 | n6115 ;
  assign n6120 = x17 & x32 ;
  assign n6121 = x18 & x31 ;
  assign n6122 = ( ~n6115 & n6120 ) | ( ~n6115 & n6121 ) | ( n6120 & n6121 ) ;
  assign n6123 = n6120 & n6121 ;
  assign n6124 = ( ~n6114 & n6122 ) | ( ~n6114 & n6123 ) | ( n6122 & n6123 ) ;
  assign n6125 = ~n6119 & n6124 ;
  assign n6126 = n6118 | n6125 ;
  assign n6127 = n6111 & n6126 ;
  assign n6128 = n6111 | n6126 ;
  assign n6129 = ~n6127 & n6128 ;
  assign n6130 = n1432 & n3280 ;
  assign n6131 = n1437 & n2709 ;
  assign n6132 = n6130 | n6131 ;
  assign n6133 = n1434 & n2369 ;
  assign n6134 = x30 & n6133 ;
  assign n6135 = ( x30 & ~n6132 ) | ( x30 & n6134 ) | ( ~n6132 & n6134 ) ;
  assign n6136 = x19 & n6135 ;
  assign n6137 = n6132 | n6133 ;
  assign n6138 = x20 & x29 ;
  assign n6139 = x21 & x28 ;
  assign n6140 = ( ~n6133 & n6138 ) | ( ~n6133 & n6139 ) | ( n6138 & n6139 ) ;
  assign n6141 = n6138 & n6139 ;
  assign n6142 = ( ~n6132 & n6140 ) | ( ~n6132 & n6141 ) | ( n6140 & n6141 ) ;
  assign n6143 = ~n6137 & n6142 ;
  assign n6144 = n6136 | n6143 ;
  assign n6145 = x2 & x47 ;
  assign n6146 = n5409 | n6145 ;
  assign n6147 = x46 & x47 ;
  assign n6148 = n77 & n6147 ;
  assign n6149 = n6146 | n6148 ;
  assign n6150 = x22 & x27 ;
  assign n6151 = ( ~n6148 & n6149 ) | ( ~n6148 & n6150 ) | ( n6149 & n6150 ) ;
  assign n6152 = ( n6148 & n6149 ) | ( n6148 & ~n6150 ) | ( n6149 & ~n6150 ) ;
  assign n6153 = ( ~n6149 & n6151 ) | ( ~n6149 & n6152 ) | ( n6151 & n6152 ) ;
  assign n6154 = n6144 & n6153 ;
  assign n6155 = n6144 & ~n6154 ;
  assign n6156 = ~n6144 & n6153 ;
  assign n6157 = n6155 | n6156 ;
  assign n6158 = n360 & n4555 ;
  assign n6159 = x37 & x40 ;
  assign n6160 = n1108 & n6159 ;
  assign n6161 = n6158 | n6160 ;
  assign n6162 = n363 & n5798 ;
  assign n6163 = x40 & n6162 ;
  assign n6164 = ( x40 & ~n6161 ) | ( x40 & n6163 ) | ( ~n6161 & n6163 ) ;
  assign n6165 = x9 & n6164 ;
  assign n6166 = n6161 | n6162 ;
  assign n6167 = x10 & x39 ;
  assign n6168 = ( n4802 & ~n6162 ) | ( n4802 & n6167 ) | ( ~n6162 & n6167 ) ;
  assign n6169 = n4802 & n6167 ;
  assign n6170 = ( ~n6161 & n6168 ) | ( ~n6161 & n6169 ) | ( n6168 & n6169 ) ;
  assign n6171 = ~n6166 & n6170 ;
  assign n6172 = n6165 | n6171 ;
  assign n6173 = ( n6129 & n6157 ) | ( n6129 & ~n6172 ) | ( n6157 & ~n6172 ) ;
  assign n6174 = ( n6129 & ~n6157 ) | ( n6129 & n6172 ) | ( ~n6157 & n6172 ) ;
  assign n6175 = ( ~n6129 & n6173 ) | ( ~n6129 & n6174 ) | ( n6173 & n6174 ) ;
  assign n6176 = n6089 & n6175 ;
  assign n6177 = n6089 | n6175 ;
  assign n6178 = ~n6176 & n6177 ;
  assign n6179 = n5917 | n5944 ;
  assign n6180 = ( n5919 & n5944 ) | ( n5919 & n6179 ) | ( n5944 & n6179 ) ;
  assign n6181 = ( n5921 & n5922 ) | ( n5921 & n6180 ) | ( n5922 & n6180 ) ;
  assign n6182 = n6178 & n6181 ;
  assign n6183 = n6178 | n6181 ;
  assign n6184 = ~n6182 & n6183 ;
  assign n6185 = ( n5989 & n5995 ) | ( n5989 & n6016 ) | ( n5995 & n6016 ) ;
  assign n6186 = n6184 | n6185 ;
  assign n6187 = n6184 & n6185 ;
  assign n6188 = n6186 & ~n6187 ;
  assign n6189 = n5949 & n6188 ;
  assign n6190 = ( n6025 & n6188 ) | ( n6025 & n6189 ) | ( n6188 & n6189 ) ;
  assign n6191 = n5949 | n6188 ;
  assign n6192 = n6025 | n6191 ;
  assign n6193 = ~n6190 & n6192 ;
  assign n6194 = n5968 | n5983 ;
  assign n6195 = n5720 | n5954 ;
  assign n6196 = ( n5954 & n5955 ) | ( n5954 & n6195 ) | ( n5955 & n6195 ) ;
  assign n6197 = n6194 | n6196 ;
  assign n6198 = n6194 & n6196 ;
  assign n6199 = n6197 & ~n6198 ;
  assign n6200 = n5614 | n6000 ;
  assign n6201 = ( n6000 & n6001 ) | ( n6000 & n6200 ) | ( n6001 & n6200 ) ;
  assign n6202 = n6199 | n6201 ;
  assign n6203 = n6199 & n6201 ;
  assign n6204 = n6202 & ~n6203 ;
  assign n6205 = n5962 | n5986 ;
  assign n6206 = ( n5962 & n5966 ) | ( n5962 & n6205 ) | ( n5966 & n6205 ) ;
  assign n6207 = n6004 | n6009 ;
  assign n6208 = ( n6009 & n6013 ) | ( n6009 & n6207 ) | ( n6013 & n6207 ) ;
  assign n6209 = n6206 & n6208 ;
  assign n6210 = n6206 & ~n6209 ;
  assign n6211 = n6208 & ~n6209 ;
  assign n6212 = n6210 | n6211 ;
  assign n6213 = n6204 | n6212 ;
  assign n6214 = n6204 & n6212 ;
  assign n6215 = n6213 & ~n6214 ;
  assign n6216 = n5904 & n6215 ;
  assign n6217 = ( n5908 & n6215 ) | ( n5908 & n6216 ) | ( n6215 & n6216 ) ;
  assign n6218 = n5904 | n5908 ;
  assign n6219 = ~n6217 & n6218 ;
  assign n6220 = n5829 | n5832 ;
  assign n6221 = n5888 | n6220 ;
  assign n6222 = n5888 & n6220 ;
  assign n6223 = n6221 & ~n6222 ;
  assign n6224 = n5820 | n6223 ;
  assign n6225 = n5820 & n6223 ;
  assign n6226 = n6224 & ~n6225 ;
  assign n6227 = n5877 | n5895 ;
  assign n6228 = n6226 & n6227 ;
  assign n6229 = n5877 & n6226 ;
  assign n6230 = ( n5880 & n6228 ) | ( n5880 & n6229 ) | ( n6228 & n6229 ) ;
  assign n6231 = n6226 | n6227 ;
  assign n6232 = n5877 | n6226 ;
  assign n6233 = ( n5880 & n6231 ) | ( n5880 & n6232 ) | ( n6231 & n6232 ) ;
  assign n6234 = ~n6230 & n6233 ;
  assign n6235 = n5939 | n5941 ;
  assign n6236 = ( n5939 & n5940 ) | ( n5939 & n6235 ) | ( n5940 & n6235 ) ;
  assign n6237 = n6234 | n6236 ;
  assign n6238 = n6234 & n6236 ;
  assign n6239 = n6237 & ~n6238 ;
  assign n6240 = n5843 | n5898 ;
  assign n6241 = ( n5843 & n5844 ) | ( n5843 & n6240 ) | ( n5844 & n6240 ) ;
  assign n6242 = n6239 & n6241 ;
  assign n6243 = n6239 | n6241 ;
  assign n6244 = ~n6242 & n6243 ;
  assign n6245 = n5972 | n5977 ;
  assign n6246 = n5854 | n6245 ;
  assign n6247 = n5854 & n6245 ;
  assign n6248 = n6246 & ~n6247 ;
  assign n6249 = n5869 | n6248 ;
  assign n6250 = n5869 & n6248 ;
  assign n6251 = n6249 & ~n6250 ;
  assign n6252 = n5826 & n5837 ;
  assign n6253 = n5837 & ~n6252 ;
  assign n6254 = n5811 & n5826 ;
  assign n6255 = ~n5837 & n6254 ;
  assign n6256 = ( n5811 & n6253 ) | ( n5811 & n6255 ) | ( n6253 & n6255 ) ;
  assign n6257 = x48 & n1658 ;
  assign n6258 = x1 & x48 ;
  assign n6259 = x25 | n6258 ;
  assign n6260 = ~n6257 & n6259 ;
  assign n6261 = n5929 & n6260 ;
  assign n6262 = n5929 | n6260 ;
  assign n6263 = ~n6261 & n6262 ;
  assign n6264 = n5805 & n6263 ;
  assign n6265 = n5805 | n6263 ;
  assign n6266 = ~n6264 & n6265 ;
  assign n6267 = n6252 & n6266 ;
  assign n6268 = ( n6256 & n6266 ) | ( n6256 & n6267 ) | ( n6266 & n6267 ) ;
  assign n6269 = n6252 | n6266 ;
  assign n6270 = n6256 | n6269 ;
  assign n6271 = ~n6268 & n6270 ;
  assign n6272 = n6251 & n6271 ;
  assign n6273 = n6251 | n6271 ;
  assign n6274 = ~n6272 & n6273 ;
  assign n6275 = n6244 & n6274 ;
  assign n6276 = n6244 | n6274 ;
  assign n6277 = ~n6275 & n6276 ;
  assign n6278 = n6215 & ~n6216 ;
  assign n6279 = n5908 & ~n6277 ;
  assign n6280 = ( n6277 & n6278 ) | ( n6277 & ~n6279 ) | ( n6278 & ~n6279 ) ;
  assign n6281 = n6219 | n6280 ;
  assign n6282 = ~n5908 & n6277 ;
  assign n6283 = n6278 & n6282 ;
  assign n6284 = ( n6219 & n6277 ) | ( n6219 & n6283 ) | ( n6277 & n6283 ) ;
  assign n6285 = n6281 & ~n6284 ;
  assign n6286 = n6193 & n6285 ;
  assign n6287 = n6193 | n6285 ;
  assign n6288 = ~n6286 & n6287 ;
  assign n6289 = n5915 | n6026 ;
  assign n6290 = ( n5915 & n5916 ) | ( n5915 & n6289 ) | ( n5916 & n6289 ) ;
  assign n6291 = ( n6047 & n6288 ) | ( n6047 & ~n6290 ) | ( n6288 & ~n6290 ) ;
  assign n6292 = ( ~n6288 & n6290 ) | ( ~n6288 & n6291 ) | ( n6290 & n6291 ) ;
  assign n6293 = ( ~n6047 & n6291 ) | ( ~n6047 & n6292 ) | ( n6291 & n6292 ) ;
  assign n6294 = n6288 & n6290 ;
  assign n6295 = n6288 | n6290 ;
  assign n6296 = n6033 & n6295 ;
  assign n6297 = ( n6043 & n6295 ) | ( n6043 & n6296 ) | ( n6295 & n6296 ) ;
  assign n6298 = n6294 | n6297 ;
  assign n6299 = n6294 | n6295 ;
  assign n6300 = ( n6046 & n6294 ) | ( n6046 & n6299 ) | ( n6294 & n6299 ) ;
  assign n6301 = ( n5523 & n6298 ) | ( n5523 & n6300 ) | ( n6298 & n6300 ) ;
  assign n6302 = ( n5522 & n6298 ) | ( n5522 & n6300 ) | ( n6298 & n6300 ) ;
  assign n6303 = ( n4853 & n6301 ) | ( n4853 & n6302 ) | ( n6301 & n6302 ) ;
  assign n6447 = n6204 | n6209 ;
  assign n6448 = ( n6209 & n6212 ) | ( n6209 & n6447 ) | ( n6212 & n6447 ) ;
  assign n6304 = x16 & x45 ;
  assign n6305 = n3874 & n6304 ;
  assign n6306 = n795 & n3483 ;
  assign n6307 = n6305 | n6306 ;
  assign n6308 = x35 & x45 ;
  assign n6309 = n1005 & n6308 ;
  assign n6310 = x34 & n6309 ;
  assign n6311 = ( x34 & ~n6307 ) | ( x34 & n6310 ) | ( ~n6307 & n6310 ) ;
  assign n6312 = x16 & n6311 ;
  assign n6313 = n6307 | n6309 ;
  assign n6314 = x5 & x45 ;
  assign n6315 = x15 & x35 ;
  assign n6316 = ( ~n6309 & n6314 ) | ( ~n6309 & n6315 ) | ( n6314 & n6315 ) ;
  assign n6317 = n6314 & n6315 ;
  assign n6318 = ( ~n6307 & n6316 ) | ( ~n6307 & n6317 ) | ( n6316 & n6317 ) ;
  assign n6319 = ~n6313 & n6318 ;
  assign n6320 = n6312 | n6319 ;
  assign n6321 = x18 & x32 ;
  assign n6322 = x23 & x27 ;
  assign n6323 = n6321 & n6322 ;
  assign n6324 = x28 & x32 ;
  assign n6325 = n1410 & n6324 ;
  assign n6326 = n1932 & n2372 ;
  assign n6327 = n6325 | n6326 ;
  assign n6328 = x28 & n6323 ;
  assign n6329 = ( x28 & ~n6327 ) | ( x28 & n6328 ) | ( ~n6327 & n6328 ) ;
  assign n6330 = x22 & n6329 ;
  assign n6331 = ( n6321 & n6322 ) | ( n6321 & ~n6327 ) | ( n6322 & ~n6327 ) ;
  assign n6332 = ( ~n6323 & n6330 ) | ( ~n6323 & n6331 ) | ( n6330 & n6331 ) ;
  assign n6333 = n6320 & n6332 ;
  assign n6334 = n6320 & ~n6333 ;
  assign n6335 = n6332 & ~n6333 ;
  assign n6336 = n6334 | n6335 ;
  assign n6337 = n5805 | n6261 ;
  assign n6338 = ( n6261 & n6263 ) | ( n6261 & n6337 ) | ( n6263 & n6337 ) ;
  assign n6339 = n6336 | n6338 ;
  assign n6340 = n6336 & n6338 ;
  assign n6341 = n6339 & ~n6340 ;
  assign n6342 = x0 & x50 ;
  assign n6343 = x2 & x48 ;
  assign n6344 = n6342 | n6343 ;
  assign n6345 = x48 & x50 ;
  assign n6346 = n67 & n6345 ;
  assign n6347 = n6344 & ~n6346 ;
  assign n6348 = n6257 | n6346 ;
  assign n6349 = ( n6346 & n6347 ) | ( n6346 & n6348 ) | ( n6347 & n6348 ) ;
  assign n6350 = n6344 & ~n6349 ;
  assign n6351 = n6257 & ~n6347 ;
  assign n6352 = n6350 | n6351 ;
  assign n6353 = n79 & n6147 ;
  assign n6354 = x17 & x47 ;
  assign n6355 = n3318 & n6354 ;
  assign n6356 = n6353 | n6355 ;
  assign n6357 = x33 & x46 ;
  assign n6358 = n1111 & n6357 ;
  assign n6359 = x47 & n6358 ;
  assign n6360 = ( x47 & ~n6356 ) | ( x47 & n6359 ) | ( ~n6356 & n6359 ) ;
  assign n6361 = x3 & n6360 ;
  assign n6362 = n6356 | n6358 ;
  assign n6363 = x4 & x46 ;
  assign n6364 = x17 & x33 ;
  assign n6365 = ( ~n6358 & n6363 ) | ( ~n6358 & n6364 ) | ( n6363 & n6364 ) ;
  assign n6366 = n6363 & n6364 ;
  assign n6367 = ( ~n6356 & n6365 ) | ( ~n6356 & n6366 ) | ( n6365 & n6366 ) ;
  assign n6368 = ~n6362 & n6367 ;
  assign n6369 = n6361 | n6368 ;
  assign n6370 = n6352 & n6369 ;
  assign n6371 = n6352 & ~n6370 ;
  assign n6372 = n6369 & ~n6370 ;
  assign n6373 = n6371 | n6372 ;
  assign n6374 = n1432 & n3595 ;
  assign n6375 = n1437 & n2965 ;
  assign n6376 = n6374 | n6375 ;
  assign n6377 = n1434 & n2709 ;
  assign n6378 = x31 & n6377 ;
  assign n6379 = ( x31 & ~n6376 ) | ( x31 & n6378 ) | ( ~n6376 & n6378 ) ;
  assign n6380 = x19 & n6379 ;
  assign n6381 = n6376 | n6377 ;
  assign n6382 = x20 & x30 ;
  assign n6383 = x21 & x29 ;
  assign n6384 = ( ~n6377 & n6382 ) | ( ~n6377 & n6383 ) | ( n6382 & n6383 ) ;
  assign n6385 = n6382 & n6383 ;
  assign n6386 = ( ~n6376 & n6384 ) | ( ~n6376 & n6385 ) | ( n6384 & n6385 ) ;
  assign n6387 = ~n6381 & n6386 ;
  assign n6388 = n6380 | n6387 ;
  assign n6389 = ~n6373 & n6388 ;
  assign n6390 = n6373 & ~n6388 ;
  assign n6391 = n6389 | n6390 ;
  assign n6392 = x7 & x43 ;
  assign n6393 = x14 & x36 ;
  assign n6394 = n6392 & n6393 ;
  assign n6395 = n200 & n5658 ;
  assign n6396 = x36 & x44 ;
  assign n6397 = n1006 & n6396 ;
  assign n6398 = n6395 | n6397 ;
  assign n6399 = x44 & n6394 ;
  assign n6400 = ( x44 & ~n6398 ) | ( x44 & n6399 ) | ( ~n6398 & n6399 ) ;
  assign n6401 = x6 & n6400 ;
  assign n6402 = ( n6392 & n6393 ) | ( n6392 & ~n6398 ) | ( n6393 & ~n6398 ) ;
  assign n6403 = ( ~n6394 & n6401 ) | ( ~n6394 & n6402 ) | ( n6401 & n6402 ) ;
  assign n6404 = n313 & n5710 ;
  assign n6405 = x13 & x42 ;
  assign n6406 = n5128 & n6405 ;
  assign n6407 = n6404 | n6406 ;
  assign n6408 = x37 & x41 ;
  assign n6409 = n415 & n6408 ;
  assign n6410 = x42 & n6409 ;
  assign n6411 = ( x42 & ~n6407 ) | ( x42 & n6410 ) | ( ~n6407 & n6410 ) ;
  assign n6412 = x8 & n6411 ;
  assign n6413 = n6407 | n6409 ;
  assign n6414 = x9 & x41 ;
  assign n6415 = ( n3772 & ~n6409 ) | ( n3772 & n6414 ) | ( ~n6409 & n6414 ) ;
  assign n6416 = n3772 & n6414 ;
  assign n6417 = ( ~n6407 & n6415 ) | ( ~n6407 & n6416 ) | ( n6415 & n6416 ) ;
  assign n6418 = ~n6413 & n6417 ;
  assign n6419 = n6412 | n6418 ;
  assign n6420 = n6403 & n6419 ;
  assign n6421 = n6403 & ~n6420 ;
  assign n6422 = n6419 & ~n6420 ;
  assign n6423 = n6421 | n6422 ;
  assign n6424 = n363 & n4050 ;
  assign n6425 = n490 & n5392 ;
  assign n6426 = n6424 | n6425 ;
  assign n6427 = n618 & n4555 ;
  assign n6428 = x38 & n6427 ;
  assign n6429 = ( x38 & ~n6426 ) | ( x38 & n6428 ) | ( ~n6426 & n6428 ) ;
  assign n6430 = x12 & n6429 ;
  assign n6431 = n6426 | n6427 ;
  assign n6432 = x10 & x40 ;
  assign n6433 = ( n5680 & ~n6427 ) | ( n5680 & n6432 ) | ( ~n6427 & n6432 ) ;
  assign n6434 = n5680 & n6432 ;
  assign n6435 = ( ~n6426 & n6433 ) | ( ~n6426 & n6434 ) | ( n6433 & n6434 ) ;
  assign n6436 = ~n6431 & n6435 ;
  assign n6437 = n6430 | n6436 ;
  assign n6438 = ~n6423 & n6437 ;
  assign n6439 = n6423 & ~n6437 ;
  assign n6440 = n6438 | n6439 ;
  assign n6441 = n6391 & ~n6440 ;
  assign n6442 = ~n6391 & n6440 ;
  assign n6443 = n6441 | n6442 ;
  assign n6444 = n6341 & n6443 ;
  assign n6445 = n6341 | n6443 ;
  assign n6446 = ~n6444 & n6445 ;
  assign n6449 = n6446 & n6448 ;
  assign n6450 = n6448 & ~n6449 ;
  assign n6451 = n6446 & ~n6448 ;
  assign n6452 = n6450 | n6451 ;
  assign n6453 = ( n6239 & n6241 ) | ( n6239 & n6274 ) | ( n6241 & n6274 ) ;
  assign n6454 = n6446 | n6453 ;
  assign n6455 = ( ~n6448 & n6453 ) | ( ~n6448 & n6454 ) | ( n6453 & n6454 ) ;
  assign n6456 = n6450 | n6455 ;
  assign n6457 = ~n6453 & n6455 ;
  assign n6458 = ( n6450 & ~n6453 ) | ( n6450 & n6457 ) | ( ~n6453 & n6457 ) ;
  assign n6459 = ( ~n6452 & n6456 ) | ( ~n6452 & n6458 ) | ( n6456 & n6458 ) ;
  assign n6460 = n6217 & n6456 ;
  assign n6461 = n6217 & ~n6452 ;
  assign n6462 = ( n6458 & n6460 ) | ( n6458 & n6461 ) | ( n6460 & n6461 ) ;
  assign n6463 = ( n6284 & n6459 ) | ( n6284 & n6462 ) | ( n6459 & n6462 ) ;
  assign n6464 = n6217 | n6456 ;
  assign n6465 = ~n6217 & n6452 ;
  assign n6466 = ( n6458 & n6464 ) | ( n6458 & ~n6465 ) | ( n6464 & ~n6465 ) ;
  assign n6467 = n6284 | n6466 ;
  assign n6468 = ~n6463 & n6467 ;
  assign n6469 = n6251 | n6267 ;
  assign n6470 = n6251 | n6266 ;
  assign n6471 = ( n6256 & n6469 ) | ( n6256 & n6470 ) | ( n6469 & n6470 ) ;
  assign n6472 = ( n6268 & n6271 ) | ( n6268 & n6471 ) | ( n6271 & n6471 ) ;
  assign n6473 = n6230 | n6236 ;
  assign n6474 = ( n6230 & n6234 ) | ( n6230 & n6473 ) | ( n6234 & n6473 ) ;
  assign n6475 = n6472 | n6474 ;
  assign n6476 = n6472 & n6474 ;
  assign n6477 = n6475 & ~n6476 ;
  assign n6478 = n5820 | n6222 ;
  assign n6479 = ( n6222 & n6223 ) | ( n6222 & n6478 ) | ( n6223 & n6478 ) ;
  assign n6480 = n5869 | n6247 ;
  assign n6481 = ( n6247 & n6248 ) | ( n6247 & n6480 ) | ( n6248 & n6480 ) ;
  assign n6482 = n6479 | n6481 ;
  assign n6483 = n6479 & n6481 ;
  assign n6484 = n6482 & ~n6483 ;
  assign n6485 = ~n6148 & n6150 ;
  assign n6486 = ( n6148 & n6149 ) | ( n6148 & n6485 ) | ( n6149 & n6485 ) ;
  assign n6487 = n6099 | n6486 ;
  assign n6488 = n6099 & n6486 ;
  assign n6489 = n6487 & ~n6488 ;
  assign n6490 = n6079 | n6489 ;
  assign n6491 = n6079 & n6489 ;
  assign n6492 = n6490 & ~n6491 ;
  assign n6493 = n6484 & n6492 ;
  assign n6494 = n6484 | n6492 ;
  assign n6495 = ~n6493 & n6494 ;
  assign n6496 = n6477 & n6495 ;
  assign n6497 = n6477 | n6495 ;
  assign n6498 = ~n6496 & n6497 ;
  assign n6499 = n6182 | n6498 ;
  assign n6500 = n6187 | n6499 ;
  assign n6501 = n6156 & n6172 ;
  assign n6502 = ( n6155 & n6172 ) | ( n6155 & n6501 ) | ( n6172 & n6501 ) ;
  assign n6503 = ( n6106 & n6108 ) | ( n6106 & n6126 ) | ( n6108 & n6126 ) ;
  assign n6504 = n6154 | n6503 ;
  assign n6505 = n6502 | n6504 ;
  assign n6506 = n6154 & n6503 ;
  assign n6507 = ( n6502 & n6503 ) | ( n6502 & n6506 ) | ( n6503 & n6506 ) ;
  assign n6508 = n6505 & ~n6507 ;
  assign n6509 = x1 & x49 ;
  assign n6510 = n2340 & n6509 ;
  assign n6511 = n2340 | n6509 ;
  assign n6512 = ~n6510 & n6511 ;
  assign n6513 = n6059 | n6512 ;
  assign n6514 = n6059 & n6512 ;
  assign n6515 = n6513 & ~n6514 ;
  assign n6516 = n6166 & n6515 ;
  assign n6517 = n6166 | n6515 ;
  assign n6518 = ~n6516 & n6517 ;
  assign n6519 = n6508 & n6518 ;
  assign n6520 = n6508 | n6518 ;
  assign n6521 = ~n6519 & n6520 ;
  assign n6522 = ~n6051 & n6053 ;
  assign n6523 = ( n6051 & n6052 ) | ( n6051 & n6522 ) | ( n6052 & n6522 ) ;
  assign n6524 = n6119 | n6137 ;
  assign n6525 = n6119 & n6137 ;
  assign n6526 = n6524 & ~n6525 ;
  assign n6527 = n6523 | n6526 ;
  assign n6528 = n6523 & n6526 ;
  assign n6529 = n6527 & ~n6528 ;
  assign n6530 = n6066 | n6086 ;
  assign n6531 = ( n6066 & n6069 ) | ( n6066 & n6530 ) | ( n6069 & n6530 ) ;
  assign n6532 = n6529 & n6531 ;
  assign n6533 = n6529 | n6531 ;
  assign n6534 = ~n6532 & n6533 ;
  assign n6535 = ( n6194 & n6196 ) | ( n6194 & n6201 ) | ( n6196 & n6201 ) ;
  assign n6536 = n6534 | n6535 ;
  assign n6537 = n6534 & n6535 ;
  assign n6538 = n6536 & ~n6537 ;
  assign n6539 = n6157 & ~n6502 ;
  assign n6540 = ~n6156 & n6172 ;
  assign n6541 = ~n6155 & n6540 ;
  assign n6542 = n6129 & n6541 ;
  assign n6543 = ( n6129 & n6539 ) | ( n6129 & n6542 ) | ( n6539 & n6542 ) ;
  assign n6544 = n6538 & n6543 ;
  assign n6545 = ( n6176 & n6538 ) | ( n6176 & n6544 ) | ( n6538 & n6544 ) ;
  assign n6546 = n6538 | n6543 ;
  assign n6547 = n6176 | n6546 ;
  assign n6548 = ~n6545 & n6547 ;
  assign n6549 = n6521 & n6548 ;
  assign n6550 = n6521 | n6548 ;
  assign n6551 = ~n6549 & n6550 ;
  assign n6552 = ( n6182 & n6185 ) | ( n6182 & n6498 ) | ( n6185 & n6498 ) ;
  assign n6553 = n6182 & n6498 ;
  assign n6554 = ( n6184 & n6552 ) | ( n6184 & n6553 ) | ( n6552 & n6553 ) ;
  assign n6555 = n6551 & ~n6554 ;
  assign n6556 = n6500 & n6555 ;
  assign n6557 = ~n6551 & n6554 ;
  assign n6558 = ( n6500 & n6551 ) | ( n6500 & ~n6557 ) | ( n6551 & ~n6557 ) ;
  assign n6559 = ~n6556 & n6558 ;
  assign n6560 = n6468 & n6559 ;
  assign n6561 = n6468 | n6559 ;
  assign n6562 = ~n6560 & n6561 ;
  assign n6563 = n6190 | n6285 ;
  assign n6564 = ( n6190 & n6193 ) | ( n6190 & n6563 ) | ( n6193 & n6563 ) ;
  assign n6565 = ( n6303 & ~n6562 ) | ( n6303 & n6564 ) | ( ~n6562 & n6564 ) ;
  assign n6566 = ( n6562 & ~n6564 ) | ( n6562 & n6565 ) | ( ~n6564 & n6565 ) ;
  assign n6567 = ( ~n6303 & n6565 ) | ( ~n6303 & n6566 ) | ( n6565 & n6566 ) ;
  assign n6568 = n6562 & n6564 ;
  assign n6569 = n6562 | n6564 ;
  assign n6570 = n6568 | n6569 ;
  assign n6571 = ( n6303 & n6568 ) | ( n6303 & n6570 ) | ( n6568 & n6570 ) ;
  assign n6572 = x0 & x51 ;
  assign n6573 = n6510 & n6572 ;
  assign n6574 = n6510 & ~n6573 ;
  assign n6575 = ~n6510 & n6572 ;
  assign n6576 = x1 & x50 ;
  assign n6577 = x26 & n6576 ;
  assign n6578 = x26 & ~n6576 ;
  assign n6579 = ( n6576 & ~n6577 ) | ( n6576 & n6578 ) | ( ~n6577 & n6578 ) ;
  assign n6580 = ~n6575 & n6579 ;
  assign n6581 = ~n6574 & n6580 ;
  assign n6582 = n6575 & ~n6579 ;
  assign n6583 = ( n6574 & ~n6579 ) | ( n6574 & n6582 ) | ( ~n6579 & n6582 ) ;
  assign n6584 = n6581 | n6583 ;
  assign n6585 = x17 & x34 ;
  assign n6586 = n1437 & n4062 ;
  assign n6587 = x20 & x31 ;
  assign n6588 = x19 & x32 ;
  assign n6589 = n6587 | n6588 ;
  assign n6590 = ( n6585 & n6586 ) | ( n6585 & ~n6589 ) | ( n6586 & ~n6589 ) ;
  assign n6591 = n6585 & ~n6590 ;
  assign n6592 = ~n6586 & n6589 ;
  assign n6593 = n6585 | n6592 ;
  assign n6594 = ~n6591 & n6593 ;
  assign n6595 = n6584 & n6594 ;
  assign n6596 = n6584 | n6594 ;
  assign n6597 = ~n6595 & n6596 ;
  assign n6598 = n6523 | n6525 ;
  assign n6599 = ( n6525 & n6526 ) | ( n6525 & n6598 ) | ( n6526 & n6598 ) ;
  assign n6600 = n6597 | n6599 ;
  assign n6601 = n6597 & n6599 ;
  assign n6602 = n6600 & ~n6601 ;
  assign n6603 = x5 & x46 ;
  assign n6604 = x16 & x35 ;
  assign n6605 = n6603 & n6604 ;
  assign n6606 = n1292 & n6357 ;
  assign n6607 = n1018 & n3129 ;
  assign n6608 = n6606 | n6607 ;
  assign n6609 = x33 & n6605 ;
  assign n6610 = ( x33 & ~n6608 ) | ( x33 & n6609 ) | ( ~n6608 & n6609 ) ;
  assign n6611 = x18 & n6610 ;
  assign n6612 = ( n6603 & n6604 ) | ( n6603 & ~n6608 ) | ( n6604 & ~n6608 ) ;
  assign n6613 = ( ~n6605 & n6611 ) | ( ~n6605 & n6612 ) | ( n6611 & n6612 ) ;
  assign n6614 = n1337 & n3280 ;
  assign n6615 = n1585 & n2709 ;
  assign n6616 = n6614 | n6615 ;
  assign n6617 = n1932 & n2369 ;
  assign n6618 = x30 & n6617 ;
  assign n6619 = ( x30 & ~n6616 ) | ( x30 & n6618 ) | ( ~n6616 & n6618 ) ;
  assign n6620 = x21 & n6619 ;
  assign n6621 = n6616 | n6617 ;
  assign n6622 = x22 & x29 ;
  assign n6623 = x23 & x28 ;
  assign n6624 = ( ~n6617 & n6622 ) | ( ~n6617 & n6623 ) | ( n6622 & n6623 ) ;
  assign n6625 = n6622 & n6623 ;
  assign n6626 = ( ~n6616 & n6624 ) | ( ~n6616 & n6625 ) | ( n6624 & n6625 ) ;
  assign n6627 = ~n6621 & n6626 ;
  assign n6628 = n6620 | n6627 ;
  assign n6629 = n6613 & n6628 ;
  assign n6630 = n6613 & ~n6629 ;
  assign n6631 = n6628 & ~n6629 ;
  assign n6632 = n6630 | n6631 ;
  assign n6633 = n792 & n3770 ;
  assign n6634 = x15 & x36 ;
  assign n6635 = x6 & x45 ;
  assign n6636 = n6634 & n6635 ;
  assign n6637 = n6633 | n6636 ;
  assign n6638 = x37 & x45 ;
  assign n6639 = n1006 & n6638 ;
  assign n6640 = n6637 | n6639 ;
  assign n6641 = x14 & x37 ;
  assign n6642 = ( n6635 & ~n6639 ) | ( n6635 & n6641 ) | ( ~n6639 & n6641 ) ;
  assign n6643 = n6635 & n6641 ;
  assign n6644 = ( ~n6637 & n6642 ) | ( ~n6637 & n6643 ) | ( n6642 & n6643 ) ;
  assign n6645 = ~n6640 & n6644 ;
  assign n6646 = n6634 & n6639 ;
  assign n6647 = ( n6634 & ~n6637 ) | ( n6634 & n6646 ) | ( ~n6637 & n6646 ) ;
  assign n6648 = n6645 | n6647 ;
  assign n6649 = ~n6632 & n6648 ;
  assign n6650 = n6632 & ~n6648 ;
  assign n6651 = n6649 | n6650 ;
  assign n6652 = n251 & n5658 ;
  assign n6653 = x13 & x44 ;
  assign n6654 = n5120 & n6653 ;
  assign n6655 = n6652 | n6654 ;
  assign n6656 = x13 & x43 ;
  assign n6657 = n5390 & n6656 ;
  assign n6658 = x44 & n6657 ;
  assign n6659 = ( x44 & ~n6655 ) | ( x44 & n6658 ) | ( ~n6655 & n6658 ) ;
  assign n6660 = x7 & n6659 ;
  assign n6661 = n6655 | n6657 ;
  assign n6662 = x8 & x43 ;
  assign n6663 = x13 & x38 ;
  assign n6664 = ( ~n6657 & n6662 ) | ( ~n6657 & n6663 ) | ( n6662 & n6663 ) ;
  assign n6665 = n6662 & n6663 ;
  assign n6666 = ( ~n6655 & n6664 ) | ( ~n6655 & n6665 ) | ( n6664 & n6665 ) ;
  assign n6667 = ~n6661 & n6666 ;
  assign n6668 = n6660 | n6667 ;
  assign n6669 = x9 & x42 ;
  assign n6670 = n5221 & n6669 ;
  assign n6671 = n360 & n5710 ;
  assign n6672 = n6670 | n6671 ;
  assign n6673 = n363 & n4350 ;
  assign n6674 = n6669 & n6673 ;
  assign n6675 = ( n6669 & ~n6672 ) | ( n6669 & n6674 ) | ( ~n6672 & n6674 ) ;
  assign n6676 = n6672 | n6673 ;
  assign n6677 = x10 & x41 ;
  assign n6678 = ( n5221 & ~n6673 ) | ( n5221 & n6677 ) | ( ~n6673 & n6677 ) ;
  assign n6679 = n5221 & n6677 ;
  assign n6680 = ( ~n6672 & n6678 ) | ( ~n6672 & n6679 ) | ( n6678 & n6679 ) ;
  assign n6681 = ~n6676 & n6680 ;
  assign n6682 = n6675 | n6681 ;
  assign n6683 = n6668 & n6682 ;
  assign n6684 = n6668 & ~n6683 ;
  assign n6685 = x24 & x27 ;
  assign n6686 = n2511 | n6685 ;
  assign n6687 = n1912 & n2267 ;
  assign n6688 = x11 & x40 ;
  assign n6689 = ~n6687 & n6688 ;
  assign n6690 = n6686 | n6687 ;
  assign n6691 = ( n6687 & n6689 ) | ( n6687 & n6690 ) | ( n6689 & n6690 ) ;
  assign n6692 = n6686 & ~n6691 ;
  assign n6693 = ( ~n6686 & n6687 ) | ( ~n6686 & n6688 ) | ( n6687 & n6688 ) ;
  assign n6694 = n6688 & n6693 ;
  assign n6695 = n6692 | n6694 ;
  assign n6696 = ~n6668 & n6682 ;
  assign n6697 = n6695 & n6696 ;
  assign n6698 = ( n6684 & n6695 ) | ( n6684 & n6697 ) | ( n6695 & n6697 ) ;
  assign n6699 = n6695 | n6696 ;
  assign n6700 = n6684 | n6699 ;
  assign n6701 = ~n6698 & n6700 ;
  assign n6702 = n6651 & ~n6701 ;
  assign n6703 = ~n6651 & n6701 ;
  assign n6704 = n6702 | n6703 ;
  assign n6705 = n6602 & n6704 ;
  assign n6706 = n6602 | n6704 ;
  assign n6707 = ~n6705 & n6706 ;
  assign n6708 = ( n6472 & n6474 ) | ( n6472 & n6495 ) | ( n6474 & n6495 ) ;
  assign n6709 = n6707 & n6708 ;
  assign n6710 = n6707 | n6708 ;
  assign n6711 = ~n6709 & n6710 ;
  assign n6712 = n6521 | n6545 ;
  assign n6713 = ( n6545 & n6548 ) | ( n6545 & n6712 ) | ( n6548 & n6712 ) ;
  assign n6714 = n6711 & n6713 ;
  assign n6715 = n6711 | n6713 ;
  assign n6716 = ~n6714 & n6715 ;
  assign n6717 = n6554 & n6716 ;
  assign n6718 = ( n6556 & n6716 ) | ( n6556 & n6717 ) | ( n6716 & n6717 ) ;
  assign n6719 = n6554 | n6716 ;
  assign n6720 = n6556 | n6719 ;
  assign n6721 = ~n6718 & n6720 ;
  assign n6722 = n6532 | n6535 ;
  assign n6723 = ( n6532 & n6534 ) | ( n6532 & n6722 ) | ( n6534 & n6722 ) ;
  assign n6724 = ( n6154 & n6503 ) | ( n6154 & n6518 ) | ( n6503 & n6518 ) ;
  assign n6725 = n6503 | n6518 ;
  assign n6726 = ( n6502 & n6724 ) | ( n6502 & n6725 ) | ( n6724 & n6725 ) ;
  assign n6727 = n6723 | n6726 ;
  assign n6728 = n6723 & n6726 ;
  assign n6729 = n6727 & ~n6728 ;
  assign n6730 = ( n6079 & n6099 ) | ( n6079 & n6486 ) | ( n6099 & n6486 ) ;
  assign n6731 = n6166 | n6514 ;
  assign n6732 = ( n6514 & n6515 ) | ( n6514 & n6731 ) | ( n6515 & n6731 ) ;
  assign n6733 = n6730 | n6732 ;
  assign n6734 = n6730 & n6732 ;
  assign n6735 = n6733 & ~n6734 ;
  assign n6736 = n6370 | n6388 ;
  assign n6737 = n6735 | n6736 ;
  assign n6738 = n6370 | n6735 ;
  assign n6739 = ( n6373 & n6737 ) | ( n6373 & n6738 ) | ( n6737 & n6738 ) ;
  assign n6740 = n6735 & n6736 ;
  assign n6741 = n6370 & n6735 ;
  assign n6742 = ( n6373 & n6740 ) | ( n6373 & n6741 ) | ( n6740 & n6741 ) ;
  assign n6743 = n6739 & ~n6742 ;
  assign n6744 = n6729 & n6743 ;
  assign n6745 = n6729 | n6743 ;
  assign n6746 = ~n6744 & n6745 ;
  assign n6747 = ( n6448 & n6453 ) | ( n6448 & n6454 ) | ( n6453 & n6454 ) ;
  assign n6748 = ( n6449 & n6451 ) | ( n6449 & n6747 ) | ( n6451 & n6747 ) ;
  assign n6749 = n6449 | n6747 ;
  assign n6750 = ( n6450 & n6748 ) | ( n6450 & n6749 ) | ( n6748 & n6749 ) ;
  assign n6751 = n6746 & n6750 ;
  assign n6752 = n6746 | n6750 ;
  assign n6753 = ~n6751 & n6752 ;
  assign n6754 = n6313 | n6431 ;
  assign n6755 = n6313 & n6431 ;
  assign n6756 = n6754 & ~n6755 ;
  assign n6757 = x47 & x49 ;
  assign n6758 = n119 & n6757 ;
  assign n6759 = x48 & x49 ;
  assign n6760 = n77 & n6759 ;
  assign n6761 = n6758 | n6760 ;
  assign n6762 = x47 & x48 ;
  assign n6763 = n79 & n6762 ;
  assign n6764 = x49 & n6763 ;
  assign n6765 = ( x49 & ~n6761 ) | ( x49 & n6764 ) | ( ~n6761 & n6764 ) ;
  assign n6766 = x2 & n6765 ;
  assign n6767 = n6761 | n6763 ;
  assign n6768 = x3 & x48 ;
  assign n6769 = x4 & x47 ;
  assign n6770 = ( ~n6763 & n6768 ) | ( ~n6763 & n6769 ) | ( n6768 & n6769 ) ;
  assign n6771 = n6768 & n6769 ;
  assign n6772 = ( ~n6761 & n6770 ) | ( ~n6761 & n6771 ) | ( n6770 & n6771 ) ;
  assign n6773 = ~n6767 & n6772 ;
  assign n6774 = n6766 | n6773 ;
  assign n6775 = n6756 & n6774 ;
  assign n6776 = n6756 & ~n6775 ;
  assign n6777 = n6774 & ~n6775 ;
  assign n6778 = n6776 | n6777 ;
  assign n6779 = n6333 | n6338 ;
  assign n6780 = ( n6333 & n6336 ) | ( n6333 & n6779 ) | ( n6336 & n6779 ) ;
  assign n6781 = n6778 | n6780 ;
  assign n6782 = n6778 & n6780 ;
  assign n6783 = n6781 & ~n6782 ;
  assign n6784 = n6483 | n6493 ;
  assign n6785 = n6783 & n6784 ;
  assign n6786 = n6783 | n6784 ;
  assign n6787 = ~n6785 & n6786 ;
  assign n6788 = ( n6341 & n6391 ) | ( n6341 & n6440 ) | ( n6391 & n6440 ) ;
  assign n6789 = n6787 | n6788 ;
  assign n6790 = n6787 & n6788 ;
  assign n6791 = n6789 & ~n6790 ;
  assign n6792 = n6394 | n6398 ;
  assign n6793 = n6413 | n6792 ;
  assign n6794 = n6413 & n6792 ;
  assign n6795 = n6793 & ~n6794 ;
  assign n6796 = n6323 | n6327 ;
  assign n6797 = n6795 | n6796 ;
  assign n6798 = n6795 & n6796 ;
  assign n6799 = n6797 & ~n6798 ;
  assign n6800 = n6420 | n6437 ;
  assign n6801 = n6799 & n6800 ;
  assign n6802 = n6420 & n6799 ;
  assign n6803 = ( n6423 & n6801 ) | ( n6423 & n6802 ) | ( n6801 & n6802 ) ;
  assign n6804 = n6799 | n6800 ;
  assign n6805 = n6420 | n6799 ;
  assign n6806 = ( n6423 & n6804 ) | ( n6423 & n6805 ) | ( n6804 & n6805 ) ;
  assign n6807 = ~n6803 & n6806 ;
  assign n6808 = n6362 | n6381 ;
  assign n6809 = n6362 & n6381 ;
  assign n6810 = n6808 & ~n6809 ;
  assign n6811 = n6349 | n6810 ;
  assign n6812 = n6349 & n6810 ;
  assign n6813 = n6811 & ~n6812 ;
  assign n6814 = n6807 & n6813 ;
  assign n6815 = n6807 | n6813 ;
  assign n6816 = ~n6814 & n6815 ;
  assign n6817 = n6791 & n6816 ;
  assign n6818 = n6791 | n6816 ;
  assign n6819 = ~n6817 & n6818 ;
  assign n6820 = n6753 & n6819 ;
  assign n6821 = n6753 | n6819 ;
  assign n6822 = ~n6820 & n6821 ;
  assign n6823 = n6721 & n6822 ;
  assign n6824 = n6721 | n6822 ;
  assign n6825 = ~n6823 & n6824 ;
  assign n6826 = n6463 | n6559 ;
  assign n6827 = ( n6463 & n6468 ) | ( n6463 & n6826 ) | ( n6468 & n6826 ) ;
  assign n6828 = ( n6571 & n6825 ) | ( n6571 & ~n6827 ) | ( n6825 & ~n6827 ) ;
  assign n6829 = ( ~n6825 & n6827 ) | ( ~n6825 & n6828 ) | ( n6827 & n6828 ) ;
  assign n6830 = ( ~n6571 & n6828 ) | ( ~n6571 & n6829 ) | ( n6828 & n6829 ) ;
  assign n6844 = n6349 | n6809 ;
  assign n6845 = ( n6809 & n6810 ) | ( n6809 & n6844 ) | ( n6810 & n6844 ) ;
  assign n6831 = x2 & x50 ;
  assign n6832 = x3 & x49 ;
  assign n6833 = n6831 | n6832 ;
  assign n6834 = x49 & x50 ;
  assign n6835 = n77 & n6834 ;
  assign n6836 = x19 & x33 ;
  assign n6837 = ~n6835 & n6836 ;
  assign n6838 = n6833 | n6835 ;
  assign n6839 = ( n6835 & n6837 ) | ( n6835 & n6838 ) | ( n6837 & n6838 ) ;
  assign n6840 = n6833 & ~n6839 ;
  assign n6841 = ( ~n6833 & n6835 ) | ( ~n6833 & n6836 ) | ( n6835 & n6836 ) ;
  assign n6842 = n6836 & n6841 ;
  assign n6843 = n6840 | n6842 ;
  assign n6846 = n6843 & n6845 ;
  assign n6847 = n6845 & ~n6846 ;
  assign n6849 = n6794 | n6796 ;
  assign n6850 = ( n6794 & n6795 ) | ( n6794 & n6849 ) | ( n6795 & n6849 ) ;
  assign n6848 = n6843 & ~n6845 ;
  assign n6851 = n6848 & n6850 ;
  assign n6852 = ( n6847 & n6850 ) | ( n6847 & n6851 ) | ( n6850 & n6851 ) ;
  assign n6853 = n6848 | n6850 ;
  assign n6854 = n6847 | n6853 ;
  assign n6855 = ~n6852 & n6854 ;
  assign n6856 = n6782 | n6784 ;
  assign n6857 = ( n6782 & n6783 ) | ( n6782 & n6856 ) | ( n6783 & n6856 ) ;
  assign n6858 = n6855 | n6857 ;
  assign n6859 = n6855 & n6857 ;
  assign n6860 = n6858 & ~n6859 ;
  assign n6861 = n6683 | n6698 ;
  assign n6862 = n6755 | n6775 ;
  assign n6863 = x1 & x51 ;
  assign n6864 = n2724 | n6863 ;
  assign n6865 = n2724 & n6863 ;
  assign n6866 = n6864 & ~n6865 ;
  assign n6867 = n6577 & n6866 ;
  assign n6868 = n6577 | n6866 ;
  assign n6869 = ~n6867 & n6868 ;
  assign n6870 = n6691 & n6869 ;
  assign n6871 = n6691 | n6869 ;
  assign n6872 = ~n6870 & n6871 ;
  assign n6873 = n6862 & n6872 ;
  assign n6874 = n6862 | n6872 ;
  assign n6875 = ~n6873 & n6874 ;
  assign n6876 = n6861 & n6875 ;
  assign n6877 = n6861 | n6875 ;
  assign n6878 = ~n6876 & n6877 ;
  assign n6879 = n6860 & n6878 ;
  assign n6880 = n6860 | n6878 ;
  assign n6881 = ~n6879 & n6880 ;
  assign n6882 = n6709 | n6881 ;
  assign n6883 = n6714 | n6882 ;
  assign n6884 = n6709 & n6881 ;
  assign n6885 = ( n6714 & n6881 ) | ( n6714 & n6884 ) | ( n6881 & n6884 ) ;
  assign n6886 = n6883 & ~n6885 ;
  assign n6887 = n6575 & n6579 ;
  assign n6888 = ( n6574 & n6579 ) | ( n6574 & n6887 ) | ( n6579 & n6887 ) ;
  assign n6889 = n6573 | n6676 ;
  assign n6890 = n6888 | n6889 ;
  assign n6891 = n6573 & n6676 ;
  assign n6892 = ( n6676 & n6888 ) | ( n6676 & n6891 ) | ( n6888 & n6891 ) ;
  assign n6893 = n6890 & ~n6892 ;
  assign n6894 = x4 & x48 ;
  assign n6895 = x17 & x35 ;
  assign n6896 = n6894 & n6895 ;
  assign n6897 = x35 & n707 ;
  assign n6898 = x48 & n82 ;
  assign n6899 = n6897 | n6898 ;
  assign n6900 = x52 & ~n6896 ;
  assign n6901 = n6899 & n6900 ;
  assign n6902 = x0 & x52 ;
  assign n6903 = ~n6901 & n6902 ;
  assign n6904 = ( n6894 & n6895 ) | ( n6894 & ~n6901 ) | ( n6895 & ~n6901 ) ;
  assign n6905 = ( ~n6896 & n6903 ) | ( ~n6896 & n6904 ) | ( n6903 & n6904 ) ;
  assign n6906 = ~n6893 & n6905 ;
  assign n6907 = n6892 | n6905 ;
  assign n6908 = n6890 & ~n6907 ;
  assign n6909 = n6906 | n6908 ;
  assign n6910 = n6595 | n6599 ;
  assign n6911 = ( n6595 & n6597 ) | ( n6595 & n6910 ) | ( n6597 & n6910 ) ;
  assign n6912 = n6909 | n6911 ;
  assign n6913 = n6909 & n6911 ;
  assign n6914 = n6912 & ~n6913 ;
  assign n6915 = n6734 | n6742 ;
  assign n6916 = n6914 | n6915 ;
  assign n6917 = n6914 & n6915 ;
  assign n6918 = n6916 & ~n6917 ;
  assign n6919 = n6605 | n6608 ;
  assign n6920 = n6661 | n6919 ;
  assign n6921 = n6661 & n6919 ;
  assign n6922 = n6920 & ~n6921 ;
  assign n6923 = n6621 | n6922 ;
  assign n6924 = n6621 & n6922 ;
  assign n6925 = n6923 & ~n6924 ;
  assign n6926 = n6585 | n6586 ;
  assign n6927 = ( n6586 & ~n6590 ) | ( n6586 & n6926 ) | ( ~n6590 & n6926 ) ;
  assign n6928 = n6767 | n6927 ;
  assign n6929 = n6767 & n6927 ;
  assign n6930 = n6928 & ~n6929 ;
  assign n6931 = n6640 | n6930 ;
  assign n6932 = n6640 & n6930 ;
  assign n6933 = n6931 & ~n6932 ;
  assign n6934 = n6629 | n6648 ;
  assign n6935 = n6933 | n6934 ;
  assign n6936 = n6629 | n6933 ;
  assign n6937 = ( n6632 & n6935 ) | ( n6632 & n6936 ) | ( n6935 & n6936 ) ;
  assign n6938 = n6933 & n6934 ;
  assign n6939 = n6629 & n6933 ;
  assign n6940 = ( n6632 & n6938 ) | ( n6632 & n6939 ) | ( n6938 & n6939 ) ;
  assign n6941 = n6937 & ~n6940 ;
  assign n6942 = n6925 & n6941 ;
  assign n6943 = n6925 | n6941 ;
  assign n6944 = ~n6942 & n6943 ;
  assign n6945 = ( n6602 & n6651 ) | ( n6602 & n6701 ) | ( n6651 & n6701 ) ;
  assign n6946 = n6944 & ~n6945 ;
  assign n6947 = ~n6944 & n6945 ;
  assign n6948 = n6946 | n6947 ;
  assign n6949 = n6918 & n6948 ;
  assign n6950 = n6918 | n6948 ;
  assign n6951 = ~n6949 & n6950 ;
  assign n6952 = ~n6886 & n6951 ;
  assign n6953 = n6885 | n6951 ;
  assign n6954 = n6883 & ~n6953 ;
  assign n6955 = n6952 | n6954 ;
  assign n6956 = x5 & x47 ;
  assign n6957 = n204 & n6147 ;
  assign n6958 = x16 & x36 ;
  assign n6959 = n6956 & n6958 ;
  assign n6960 = n6957 | n6959 ;
  assign n6961 = x36 & x46 ;
  assign n6962 = n623 & n6961 ;
  assign n6963 = n6956 & n6962 ;
  assign n6964 = ( n6956 & ~n6960 ) | ( n6956 & n6963 ) | ( ~n6960 & n6963 ) ;
  assign n6965 = n6960 | n6962 ;
  assign n6966 = x6 & x46 ;
  assign n6967 = ( n6958 & ~n6962 ) | ( n6958 & n6966 ) | ( ~n6962 & n6966 ) ;
  assign n6968 = n6958 & n6966 ;
  assign n6969 = ( ~n6960 & n6967 ) | ( ~n6960 & n6968 ) | ( n6967 & n6968 ) ;
  assign n6970 = ~n6965 & n6969 ;
  assign n6971 = n6964 | n6970 ;
  assign n6972 = x10 & x42 ;
  assign n6973 = x40 & x42 ;
  assign n6974 = n363 & n6973 ;
  assign n6975 = n618 & n5710 ;
  assign n6976 = n6974 | n6975 ;
  assign n6977 = n490 & n5813 ;
  assign n6978 = n6972 & n6977 ;
  assign n6979 = ( n6972 & ~n6976 ) | ( n6972 & n6978 ) | ( ~n6976 & n6978 ) ;
  assign n6980 = n6976 | n6977 ;
  assign n6981 = x11 & x41 ;
  assign n6982 = ( n5739 & ~n6977 ) | ( n5739 & n6981 ) | ( ~n6977 & n6981 ) ;
  assign n6983 = n5739 & n6981 ;
  assign n6984 = ( ~n6976 & n6982 ) | ( ~n6976 & n6983 ) | ( n6982 & n6983 ) ;
  assign n6985 = ~n6980 & n6984 ;
  assign n6986 = n6979 | n6985 ;
  assign n6987 = n6971 & n6986 ;
  assign n6988 = n6971 & ~n6987 ;
  assign n6989 = n6986 & ~n6987 ;
  assign n6990 = n6988 | n6989 ;
  assign n6991 = x7 & x45 ;
  assign n6992 = x8 & x44 ;
  assign n6993 = n6991 | n6992 ;
  assign n6994 = n251 & n6093 ;
  assign n6995 = x15 & x37 ;
  assign n6996 = ~n6994 & n6995 ;
  assign n6997 = n6993 | n6994 ;
  assign n6998 = ( n6994 & n6996 ) | ( n6994 & n6997 ) | ( n6996 & n6997 ) ;
  assign n6999 = n6993 & ~n6998 ;
  assign n7000 = ( ~n6993 & n6994 ) | ( ~n6993 & n6995 ) | ( n6994 & n6995 ) ;
  assign n7001 = n6995 & n7000 ;
  assign n7002 = n6999 | n7001 ;
  assign n7003 = ~n6990 & n7002 ;
  assign n7004 = n6990 & ~n7002 ;
  assign n7005 = n7003 | n7004 ;
  assign n7006 = x31 & x34 ;
  assign n7007 = n3850 & n7006 ;
  assign n7008 = n1285 & n4318 ;
  assign n7009 = n7007 | n7008 ;
  assign n7010 = n1434 & n4062 ;
  assign n7011 = x34 & n7010 ;
  assign n7012 = ( x34 & ~n7009 ) | ( x34 & n7011 ) | ( ~n7009 & n7011 ) ;
  assign n7013 = x18 & n7012 ;
  assign n7014 = n7009 | n7010 ;
  assign n7015 = x20 & x32 ;
  assign n7016 = x21 & x31 ;
  assign n7017 = ( ~n7010 & n7015 ) | ( ~n7010 & n7016 ) | ( n7015 & n7016 ) ;
  assign n7018 = n7015 & n7016 ;
  assign n7019 = ( ~n7009 & n7017 ) | ( ~n7009 & n7018 ) | ( n7017 & n7018 ) ;
  assign n7020 = ~n7014 & n7019 ;
  assign n7021 = n7013 | n7020 ;
  assign n7022 = n2148 & n3280 ;
  assign n7023 = n1932 & n2709 ;
  assign n7024 = n7022 | n7023 ;
  assign n7025 = n1686 & n2369 ;
  assign n7026 = x30 & n7025 ;
  assign n7027 = ( x30 & ~n7024 ) | ( x30 & n7026 ) | ( ~n7024 & n7026 ) ;
  assign n7028 = x22 & n7027 ;
  assign n7029 = n7024 | n7025 ;
  assign n7030 = x23 & x29 ;
  assign n7031 = x24 & x28 ;
  assign n7032 = ( ~n7025 & n7030 ) | ( ~n7025 & n7031 ) | ( n7030 & n7031 ) ;
  assign n7033 = n7030 & n7031 ;
  assign n7034 = ( ~n7024 & n7032 ) | ( ~n7024 & n7033 ) | ( n7032 & n7033 ) ;
  assign n7035 = ~n7029 & n7034 ;
  assign n7036 = n7028 | n7035 ;
  assign n7037 = n7021 & n7036 ;
  assign n7038 = n7021 & ~n7037 ;
  assign n7039 = n7036 & ~n7037 ;
  assign n7040 = n7038 | n7039 ;
  assign n7041 = x9 & x43 ;
  assign n7042 = n4586 & n7041 ;
  assign n7043 = n650 & n5392 ;
  assign n7044 = n7042 | n7043 ;
  assign n7045 = n5797 & n6656 ;
  assign n7046 = n4586 & n7045 ;
  assign n7047 = ( n4586 & ~n7044 ) | ( n4586 & n7046 ) | ( ~n7044 & n7046 ) ;
  assign n7048 = n7044 | n7045 ;
  assign n7049 = x13 & x39 ;
  assign n7050 = ( n7041 & ~n7045 ) | ( n7041 & n7049 ) | ( ~n7045 & n7049 ) ;
  assign n7051 = n7041 & n7049 ;
  assign n7052 = ( ~n7044 & n7050 ) | ( ~n7044 & n7051 ) | ( n7050 & n7051 ) ;
  assign n7053 = ~n7048 & n7052 ;
  assign n7054 = n7047 | n7053 ;
  assign n7055 = ~n7040 & n7054 ;
  assign n7056 = n7040 & ~n7054 ;
  assign n7057 = n7055 | n7056 ;
  assign n7058 = n7005 | n7057 ;
  assign n7059 = n7005 & n7057 ;
  assign n7060 = n7058 & ~n7059 ;
  assign n7061 = n6803 | n6813 ;
  assign n7062 = ( n6803 & n6807 ) | ( n6803 & n7061 ) | ( n6807 & n7061 ) ;
  assign n7063 = n7060 & n7062 ;
  assign n7064 = n7060 | n7062 ;
  assign n7065 = ~n7063 & n7064 ;
  assign n7066 = n6726 | n6743 ;
  assign n7067 = ( n6723 & n6743 ) | ( n6723 & n7066 ) | ( n6743 & n7066 ) ;
  assign n7068 = ( n6728 & n6729 ) | ( n6728 & n7067 ) | ( n6729 & n7067 ) ;
  assign n7069 = n7065 & n7068 ;
  assign n7070 = n7065 | n7068 ;
  assign n7071 = ~n7069 & n7070 ;
  assign n7072 = ( n6787 & n6788 ) | ( n6787 & n6816 ) | ( n6788 & n6816 ) ;
  assign n7073 = n7071 | n7072 ;
  assign n7074 = n7071 & n7072 ;
  assign n7075 = n7073 & ~n7074 ;
  assign n7076 = n6746 | n6819 ;
  assign n7077 = ( n6750 & n6819 ) | ( n6750 & n7076 ) | ( n6819 & n7076 ) ;
  assign n7078 = n7075 & n7077 ;
  assign n7079 = n6751 & n7075 ;
  assign n7080 = ( n6753 & n7078 ) | ( n6753 & n7079 ) | ( n7078 & n7079 ) ;
  assign n7081 = n7075 | n7077 ;
  assign n7082 = n6751 | n7075 ;
  assign n7083 = ( n6753 & n7081 ) | ( n6753 & n7082 ) | ( n7081 & n7082 ) ;
  assign n7084 = ~n7080 & n7083 ;
  assign n7085 = n6955 & n7084 ;
  assign n7086 = n6955 | n7084 ;
  assign n7087 = ~n7085 & n7086 ;
  assign n7088 = n6718 | n6721 ;
  assign n7089 = ( n6718 & n6822 ) | ( n6718 & n7088 ) | ( n6822 & n7088 ) ;
  assign n7090 = n7087 | n7089 ;
  assign n7091 = n7087 & n7089 ;
  assign n7092 = n7090 & ~n7091 ;
  assign n7093 = n6825 & n6827 ;
  assign n7094 = n6825 | n6827 ;
  assign n7095 = n7093 | n7094 ;
  assign n7096 = ( n6570 & n7093 ) | ( n6570 & n7095 ) | ( n7093 & n7095 ) ;
  assign n7097 = ( n6568 & n7093 ) | ( n6568 & n7095 ) | ( n7093 & n7095 ) ;
  assign n7098 = ( n6303 & n7096 ) | ( n6303 & n7097 ) | ( n7096 & n7097 ) ;
  assign n7099 = n7092 | n7098 ;
  assign n7100 = n7090 & n7097 ;
  assign n7101 = n7090 & n7096 ;
  assign n7102 = ( n6303 & n7100 ) | ( n6303 & n7101 ) | ( n7100 & n7101 ) ;
  assign n7103 = ~n7091 & n7102 ;
  assign n7104 = n7099 & ~n7103 ;
  assign n7105 = n7090 | n7091 ;
  assign n7106 = ( n7091 & n7097 ) | ( n7091 & n7105 ) | ( n7097 & n7105 ) ;
  assign n7107 = ( n7091 & n7096 ) | ( n7091 & n7105 ) | ( n7096 & n7105 ) ;
  assign n7108 = ( n6303 & n7106 ) | ( n6303 & n7107 ) | ( n7106 & n7107 ) ;
  assign n7109 = x2 & x51 ;
  assign n7110 = x3 & x50 ;
  assign n7111 = n7109 | n7110 ;
  assign n7112 = x50 & x51 ;
  assign n7113 = n77 & n7112 ;
  assign n7114 = n7111 & ~n7113 ;
  assign n7115 = n6865 | n7113 ;
  assign n7116 = ( n7113 & n7114 ) | ( n7113 & n7115 ) | ( n7114 & n7115 ) ;
  assign n7117 = n7111 & ~n7116 ;
  assign n7118 = n6865 & ~n7114 ;
  assign n7119 = n7117 | n7118 ;
  assign n7120 = x17 & x36 ;
  assign n7121 = x18 & x35 ;
  assign n7122 = n7120 | n7121 ;
  assign n7123 = n1020 & n4078 ;
  assign n7124 = x4 & x49 ;
  assign n7125 = ~n7123 & n7124 ;
  assign n7126 = n7122 | n7123 ;
  assign n7127 = ( n7123 & n7125 ) | ( n7123 & n7126 ) | ( n7125 & n7126 ) ;
  assign n7128 = n7122 & ~n7127 ;
  assign n7129 = ( ~n7122 & n7123 ) | ( ~n7122 & n7124 ) | ( n7123 & n7124 ) ;
  assign n7130 = n7124 & n7129 ;
  assign n7131 = n7128 | n7130 ;
  assign n7132 = n7119 & n7131 ;
  assign n7133 = n7119 & ~n7132 ;
  assign n7134 = n7131 & ~n7132 ;
  assign n7135 = n7133 | n7134 ;
  assign n7136 = n1432 & n4318 ;
  assign n7137 = n1437 & n4530 ;
  assign n7138 = n7136 | n7137 ;
  assign n7139 = n1434 & n3321 ;
  assign n7140 = x34 & n7139 ;
  assign n7141 = ( x34 & ~n7138 ) | ( x34 & n7140 ) | ( ~n7138 & n7140 ) ;
  assign n7142 = x19 & n7141 ;
  assign n7143 = n7138 | n7139 ;
  assign n7144 = x20 & x33 ;
  assign n7145 = x21 & x32 ;
  assign n7146 = ( ~n7139 & n7144 ) | ( ~n7139 & n7145 ) | ( n7144 & n7145 ) ;
  assign n7147 = n7144 & n7145 ;
  assign n7148 = ( ~n7138 & n7146 ) | ( ~n7138 & n7147 ) | ( n7146 & n7147 ) ;
  assign n7149 = ~n7143 & n7148 ;
  assign n7150 = n7142 | n7149 ;
  assign n7151 = ~n7135 & n7150 ;
  assign n7152 = n7135 & ~n7150 ;
  assign n7153 = n7151 | n7152 ;
  assign n7154 = n6846 | n6852 ;
  assign n7155 = n7153 | n7154 ;
  assign n7156 = n7153 & n7154 ;
  assign n7157 = n7155 & ~n7156 ;
  assign n7158 = n200 & n6147 ;
  assign n7159 = x6 & x47 ;
  assign n7160 = x7 & x46 ;
  assign n7161 = n7159 | n7160 ;
  assign n7162 = ( n4583 & n7158 ) | ( n4583 & n7161 ) | ( n7158 & n7161 ) ;
  assign n7163 = ( ~n4583 & n7159 ) | ( ~n4583 & n7160 ) | ( n7159 & n7160 ) ;
  assign n7164 = ( n4583 & ~n7162 ) | ( n4583 & n7163 ) | ( ~n7162 & n7163 ) ;
  assign n7165 = n313 & n6093 ;
  assign n7166 = x8 & x45 ;
  assign n7167 = x14 & x39 ;
  assign n7168 = n7166 & n7167 ;
  assign n7169 = n7165 | n7168 ;
  assign n7170 = x14 & x44 ;
  assign n7171 = n5797 & n7170 ;
  assign n7172 = n7169 | n7171 ;
  assign n7173 = x9 & x44 ;
  assign n7174 = ( n7167 & ~n7171 ) | ( n7167 & n7173 ) | ( ~n7171 & n7173 ) ;
  assign n7175 = n7167 & n7173 ;
  assign n7176 = ( ~n7169 & n7174 ) | ( ~n7169 & n7175 ) | ( n7174 & n7175 ) ;
  assign n7177 = ~n7172 & n7176 ;
  assign n7178 = n7166 & n7171 ;
  assign n7179 = ( n7166 & ~n7169 ) | ( n7166 & n7178 ) | ( ~n7169 & n7178 ) ;
  assign n7180 = n7164 & n7179 ;
  assign n7181 = ( n7164 & n7177 ) | ( n7164 & n7180 ) | ( n7177 & n7180 ) ;
  assign n7182 = n7164 & ~n7181 ;
  assign n7183 = n7177 | n7179 ;
  assign n7184 = ~n7181 & n7183 ;
  assign n7185 = n7182 | n7184 ;
  assign n7186 = x5 & x48 ;
  assign n7187 = x16 & x37 ;
  assign n7188 = n7186 | n7187 ;
  assign n7189 = x16 & x48 ;
  assign n7190 = n4454 & n7189 ;
  assign n7191 = x0 & x53 ;
  assign n7192 = ~n7190 & n7191 ;
  assign n7193 = n7188 | n7190 ;
  assign n7194 = ( n7190 & n7192 ) | ( n7190 & n7193 ) | ( n7192 & n7193 ) ;
  assign n7195 = n7188 & ~n7194 ;
  assign n7196 = ( ~n7188 & n7190 ) | ( ~n7188 & n7191 ) | ( n7190 & n7191 ) ;
  assign n7197 = n7191 & n7196 ;
  assign n7198 = n7195 | n7197 ;
  assign n7199 = ~n7185 & n7198 ;
  assign n7200 = n7185 & ~n7198 ;
  assign n7201 = n7199 | n7200 ;
  assign n7202 = n7157 | n7201 ;
  assign n7203 = n7157 & n7201 ;
  assign n7204 = n7202 & ~n7203 ;
  assign n7205 = n6432 & n6656 ;
  assign n7206 = n647 & n5813 ;
  assign n7207 = n7205 | n7206 ;
  assign n7208 = n363 & n5107 ;
  assign n7209 = x40 & n7208 ;
  assign n7210 = ( x40 & ~n7207 ) | ( x40 & n7209 ) | ( ~n7207 & n7209 ) ;
  assign n7211 = x13 & n7210 ;
  assign n7212 = n7207 | n7208 ;
  assign n7213 = x10 & x43 ;
  assign n7214 = x12 & x41 ;
  assign n7215 = ( ~n7208 & n7213 ) | ( ~n7208 & n7214 ) | ( n7213 & n7214 ) ;
  assign n7216 = n7213 & n7214 ;
  assign n7217 = ( ~n7207 & n7215 ) | ( ~n7207 & n7216 ) | ( n7215 & n7216 ) ;
  assign n7218 = ~n7212 & n7217 ;
  assign n7219 = n7211 | n7218 ;
  assign n7220 = n2148 & n3595 ;
  assign n7221 = n1932 & n2965 ;
  assign n7222 = n7220 | n7221 ;
  assign n7223 = n1686 & n2709 ;
  assign n7224 = n2392 & n7223 ;
  assign n7225 = ( n2392 & ~n7222 ) | ( n2392 & n7224 ) | ( ~n7222 & n7224 ) ;
  assign n7226 = n7222 | n7223 ;
  assign n7227 = x23 & x30 ;
  assign n7228 = ( n2868 & ~n7223 ) | ( n2868 & n7227 ) | ( ~n7223 & n7227 ) ;
  assign n7229 = n2868 & n7227 ;
  assign n7230 = ( ~n7222 & n7228 ) | ( ~n7222 & n7229 ) | ( n7228 & n7229 ) ;
  assign n7231 = ~n7226 & n7230 ;
  assign n7232 = n7225 | n7231 ;
  assign n7233 = n7219 & n7232 ;
  assign n7234 = n7219 & ~n7233 ;
  assign n7235 = x25 & x28 ;
  assign n7236 = n2267 | n7235 ;
  assign n7237 = n2372 & n2511 ;
  assign n7238 = x11 & x42 ;
  assign n7239 = ~n7237 & n7238 ;
  assign n7240 = n7236 | n7237 ;
  assign n7241 = ( n7237 & n7239 ) | ( n7237 & n7240 ) | ( n7239 & n7240 ) ;
  assign n7242 = n7236 & ~n7241 ;
  assign n7243 = ( ~n7236 & n7237 ) | ( ~n7236 & n7238 ) | ( n7237 & n7238 ) ;
  assign n7244 = n7238 & n7243 ;
  assign n7245 = n7242 | n7244 ;
  assign n7246 = ~n7219 & n7232 ;
  assign n7247 = n7245 & n7246 ;
  assign n7248 = ( n7234 & n7245 ) | ( n7234 & n7247 ) | ( n7245 & n7247 ) ;
  assign n7249 = n7245 | n7246 ;
  assign n7250 = n7234 | n7249 ;
  assign n7251 = ~n7248 & n7250 ;
  assign n7252 = n6873 | n7251 ;
  assign n7253 = n6876 | n7252 ;
  assign n7254 = n6873 & n7251 ;
  assign n7255 = ( n6876 & n7251 ) | ( n6876 & n7254 ) | ( n7251 & n7254 ) ;
  assign n7256 = n7253 & ~n7255 ;
  assign n7257 = ( n6925 & n6933 ) | ( n6925 & n6934 ) | ( n6933 & n6934 ) ;
  assign n7258 = ( n6629 & n6925 ) | ( n6629 & n6933 ) | ( n6925 & n6933 ) ;
  assign n7259 = ( n6632 & n7257 ) | ( n6632 & n7258 ) | ( n7257 & n7258 ) ;
  assign n7260 = n7256 | n7259 ;
  assign n7261 = n7256 & n7259 ;
  assign n7262 = n7260 & ~n7261 ;
  assign n7263 = n7204 & n7262 ;
  assign n7264 = n7204 | n7262 ;
  assign n7265 = ~n7263 & n7264 ;
  assign n7266 = n6944 & n6945 ;
  assign n7267 = n6918 | n7266 ;
  assign n7268 = ( n6948 & n7266 ) | ( n6948 & n7267 ) | ( n7266 & n7267 ) ;
  assign n7269 = n7265 & n7268 ;
  assign n7270 = n7265 | n7268 ;
  assign n7271 = ~n7269 & n7270 ;
  assign n7272 = ( n6885 & n6886 ) | ( n6885 & n6953 ) | ( n6886 & n6953 ) ;
  assign n7273 = n7271 & n7272 ;
  assign n7274 = n7271 | n7272 ;
  assign n7275 = ~n7273 & n7274 ;
  assign n7276 = n6621 | n6921 ;
  assign n7277 = ( n6921 & n6922 ) | ( n6921 & n7276 ) | ( n6922 & n7276 ) ;
  assign n7278 = n6691 | n6867 ;
  assign n7279 = ( n6867 & n6869 ) | ( n6867 & n7278 ) | ( n6869 & n7278 ) ;
  assign n7280 = n7277 | n7279 ;
  assign n7281 = n7277 & n7279 ;
  assign n7282 = n7280 & ~n7281 ;
  assign n7283 = ( n6640 & n6767 ) | ( n6640 & n6927 ) | ( n6767 & n6927 ) ;
  assign n7284 = n7282 | n7283 ;
  assign n7285 = n7282 & n7283 ;
  assign n7286 = n7284 & ~n7285 ;
  assign n7287 = n6913 | n7286 ;
  assign n7288 = n6917 | n7287 ;
  assign n7289 = n6913 & n7286 ;
  assign n7290 = ( n6917 & n7286 ) | ( n6917 & n7289 ) | ( n7286 & n7289 ) ;
  assign n7291 = n7288 & ~n7290 ;
  assign n7292 = n7059 | n7062 ;
  assign n7293 = ( n7059 & n7060 ) | ( n7059 & n7292 ) | ( n7060 & n7292 ) ;
  assign n7294 = n7291 & n7293 ;
  assign n7295 = n7291 | n7293 ;
  assign n7296 = ~n7294 & n7295 ;
  assign n7297 = n7069 | n7296 ;
  assign n7298 = n7074 | n7297 ;
  assign n7299 = n6896 | n6901 ;
  assign n7300 = n6839 | n7299 ;
  assign n7301 = n6839 & n7299 ;
  assign n7302 = n7300 & ~n7301 ;
  assign n7303 = n7029 | n7302 ;
  assign n7304 = n7029 & n7302 ;
  assign n7305 = n7303 & ~n7304 ;
  assign n7306 = ( n6892 & n6893 ) | ( n6892 & n6907 ) | ( n6893 & n6907 ) ;
  assign n7307 = n7037 | n7054 ;
  assign n7308 = n7306 | n7307 ;
  assign n7309 = n7037 | n7306 ;
  assign n7310 = ( n7040 & n7308 ) | ( n7040 & n7309 ) | ( n7308 & n7309 ) ;
  assign n7311 = n7306 & n7307 ;
  assign n7312 = n7037 & n7306 ;
  assign n7313 = ( n7040 & n7311 ) | ( n7040 & n7312 ) | ( n7311 & n7312 ) ;
  assign n7314 = n7310 & ~n7313 ;
  assign n7315 = n7305 & n7314 ;
  assign n7316 = n7305 | n7314 ;
  assign n7317 = ~n7315 & n7316 ;
  assign n7318 = n6965 | n7014 ;
  assign n7319 = n6965 & n7014 ;
  assign n7320 = n7318 & ~n7319 ;
  assign n7321 = n6998 | n7320 ;
  assign n7322 = n6998 & n7320 ;
  assign n7323 = n7321 & ~n7322 ;
  assign n7324 = x52 & n1954 ;
  assign n7325 = x1 & x52 ;
  assign n7326 = x27 | n7325 ;
  assign n7327 = ~n7324 & n7326 ;
  assign n7328 = n6980 | n7327 ;
  assign n7329 = n6980 & n7327 ;
  assign n7330 = n7328 & ~n7329 ;
  assign n7331 = n7048 & n7330 ;
  assign n7332 = n7048 | n7330 ;
  assign n7333 = ~n7331 & n7332 ;
  assign n7334 = n6987 | n7002 ;
  assign n7336 = ( n7323 & n7333 ) | ( n7323 & ~n7334 ) | ( n7333 & ~n7334 ) ;
  assign n7337 = ( ~n6987 & n7323 ) | ( ~n6987 & n7333 ) | ( n7323 & n7333 ) ;
  assign n7338 = ( ~n6990 & n7336 ) | ( ~n6990 & n7337 ) | ( n7336 & n7337 ) ;
  assign n7335 = ( n6987 & n6990 ) | ( n6987 & n7334 ) | ( n6990 & n7334 ) ;
  assign n7339 = ( ~n7333 & n7335 ) | ( ~n7333 & n7338 ) | ( n7335 & n7338 ) ;
  assign n7340 = ( ~n7323 & n7338 ) | ( ~n7323 & n7339 ) | ( n7338 & n7339 ) ;
  assign n7341 = n7317 & n7340 ;
  assign n7342 = n7317 & ~n7341 ;
  assign n7343 = ( n6855 & n6857 ) | ( n6855 & n6878 ) | ( n6857 & n6878 ) ;
  assign n7344 = ~n7317 & n7340 ;
  assign n7345 = n7343 | n7344 ;
  assign n7346 = n7342 | n7345 ;
  assign n7347 = n7343 & n7344 ;
  assign n7348 = ( n7342 & n7343 ) | ( n7342 & n7347 ) | ( n7343 & n7347 ) ;
  assign n7349 = n7346 & ~n7348 ;
  assign n7350 = ( n7069 & n7072 ) | ( n7069 & n7296 ) | ( n7072 & n7296 ) ;
  assign n7351 = n7069 & n7296 ;
  assign n7352 = ( n7071 & n7350 ) | ( n7071 & n7351 ) | ( n7350 & n7351 ) ;
  assign n7353 = n7349 & ~n7352 ;
  assign n7354 = n7298 & n7353 ;
  assign n7355 = ~n7349 & n7352 ;
  assign n7356 = ( n7298 & n7349 ) | ( n7298 & ~n7355 ) | ( n7349 & ~n7355 ) ;
  assign n7357 = ~n7354 & n7356 ;
  assign n7358 = n7275 & n7357 ;
  assign n7359 = n7275 | n7357 ;
  assign n7360 = ~n7358 & n7359 ;
  assign n7361 = n6955 | n7080 ;
  assign n7362 = ( n7080 & n7084 ) | ( n7080 & n7361 ) | ( n7084 & n7361 ) ;
  assign n7363 = ( n7108 & ~n7360 ) | ( n7108 & n7362 ) | ( ~n7360 & n7362 ) ;
  assign n7364 = ( n7360 & ~n7362 ) | ( n7360 & n7363 ) | ( ~n7362 & n7363 ) ;
  assign n7365 = ( ~n7108 & n7363 ) | ( ~n7108 & n7364 ) | ( n7363 & n7364 ) ;
  assign n7366 = n7341 | n7348 ;
  assign n7367 = n7290 | n7294 ;
  assign n7368 = n7366 | n7367 ;
  assign n7369 = n7366 & n7367 ;
  assign n7370 = n7368 & ~n7369 ;
  assign n7371 = n7305 | n7313 ;
  assign n7372 = ( n7313 & n7314 ) | ( n7313 & n7371 ) | ( n7314 & n7371 ) ;
  assign n7373 = x0 & x54 ;
  assign n7374 = n7324 & n7373 ;
  assign n7375 = n7324 & ~n7374 ;
  assign n7376 = ~n7324 & n7373 ;
  assign n7377 = n7375 | n7376 ;
  assign n7378 = x1 & x53 ;
  assign n7379 = n2895 & n7378 ;
  assign n7380 = n7378 & ~n7379 ;
  assign n7381 = n2895 & ~n7379 ;
  assign n7382 = n7380 | n7381 ;
  assign n7383 = ~n7377 & n7382 ;
  assign n7384 = n7377 & ~n7382 ;
  assign n7385 = n7383 | n7384 ;
  assign n7386 = x32 & x35 ;
  assign n7387 = n4258 & n7386 ;
  assign n7388 = n1432 & n3129 ;
  assign n7389 = n7387 | n7388 ;
  assign n7390 = n1585 & n3321 ;
  assign n7391 = x35 & n7390 ;
  assign n7392 = ( x35 & ~n7389 ) | ( x35 & n7391 ) | ( ~n7389 & n7391 ) ;
  assign n7393 = x19 & n7392 ;
  assign n7394 = n7389 | n7390 ;
  assign n7395 = x21 & x33 ;
  assign n7396 = x22 & x32 ;
  assign n7397 = ( ~n7390 & n7395 ) | ( ~n7390 & n7396 ) | ( n7395 & n7396 ) ;
  assign n7398 = n7395 & n7396 ;
  assign n7399 = ( ~n7389 & n7397 ) | ( ~n7389 & n7398 ) | ( n7397 & n7398 ) ;
  assign n7400 = ~n7394 & n7399 ;
  assign n7401 = n7393 | n7400 ;
  assign n7402 = n1557 & n3595 ;
  assign n7403 = n1686 & n2965 ;
  assign n7404 = n7402 | n7403 ;
  assign n7405 = n1912 & n2709 ;
  assign n7406 = x31 & n7405 ;
  assign n7407 = ( x31 & ~n7404 ) | ( x31 & n7406 ) | ( ~n7404 & n7406 ) ;
  assign n7408 = x23 & n7407 ;
  assign n7409 = n7404 | n7405 ;
  assign n7410 = x25 & x29 ;
  assign n7411 = ( n2711 & ~n7405 ) | ( n2711 & n7410 ) | ( ~n7405 & n7410 ) ;
  assign n7412 = n2711 & n7410 ;
  assign n7413 = ( ~n7404 & n7411 ) | ( ~n7404 & n7412 ) | ( n7411 & n7412 ) ;
  assign n7414 = ~n7409 & n7413 ;
  assign n7415 = n7408 | n7414 ;
  assign n7416 = n7401 & n7415 ;
  assign n7417 = n7401 & ~n7416 ;
  assign n7418 = n7415 & ~n7416 ;
  assign n7419 = n7417 | n7418 ;
  assign n7420 = n7385 & ~n7419 ;
  assign n7421 = ~n7385 & n7419 ;
  assign n7422 = n7420 | n7421 ;
  assign n7423 = n7372 & n7422 ;
  assign n7424 = n7372 & ~n7423 ;
  assign n7425 = n7333 & n7334 ;
  assign n7426 = n6987 & n7333 ;
  assign n7427 = ( n6990 & n7425 ) | ( n6990 & n7426 ) | ( n7425 & n7426 ) ;
  assign n7428 = n7335 & ~n7427 ;
  assign n7429 = n7323 & n7333 ;
  assign n7430 = ~n7335 & n7429 ;
  assign n7431 = ( n7323 & n7428 ) | ( n7323 & n7430 ) | ( n7428 & n7430 ) ;
  assign n7432 = n7427 | n7431 ;
  assign n7433 = ~n7372 & n7422 ;
  assign n7434 = n7432 & n7433 ;
  assign n7435 = ( n7424 & n7432 ) | ( n7424 & n7434 ) | ( n7432 & n7434 ) ;
  assign n7436 = n7432 | n7433 ;
  assign n7437 = n7424 | n7436 ;
  assign n7438 = ~n7435 & n7437 ;
  assign n7439 = n7370 & ~n7438 ;
  assign n7440 = n7370 | n7438 ;
  assign n7441 = ( ~n7370 & n7439 ) | ( ~n7370 & n7440 ) | ( n7439 & n7440 ) ;
  assign n7442 = n7352 | n7354 ;
  assign n7443 = n7441 & n7442 ;
  assign n7444 = n7441 & ~n7443 ;
  assign n7445 = ( n6839 & n7029 ) | ( n6839 & n7299 ) | ( n7029 & n7299 ) ;
  assign n7446 = n6998 | n7319 ;
  assign n7447 = ( n7319 & n7320 ) | ( n7319 & n7446 ) | ( n7320 & n7446 ) ;
  assign n7448 = n7445 | n7447 ;
  assign n7449 = n7445 & n7447 ;
  assign n7450 = n7448 & ~n7449 ;
  assign n7451 = n7048 | n7329 ;
  assign n7452 = ( n7329 & n7330 ) | ( n7329 & n7451 ) | ( n7330 & n7451 ) ;
  assign n7453 = n7450 | n7452 ;
  assign n7454 = n7450 & n7452 ;
  assign n7455 = n7453 & ~n7454 ;
  assign n7456 = n7156 | n7201 ;
  assign n7457 = ( n7156 & n7157 ) | ( n7156 & n7456 ) | ( n7157 & n7456 ) ;
  assign n7458 = n7455 & n7457 ;
  assign n7459 = n7455 | n7457 ;
  assign n7460 = ~n7458 & n7459 ;
  assign n7461 = n4583 & n7159 ;
  assign n7462 = n7158 | n7461 ;
  assign n7463 = n4583 & n7160 ;
  assign n7464 = n7462 | n7463 ;
  assign n7465 = n7194 | n7464 ;
  assign n7466 = n7194 & n7464 ;
  assign n7467 = n7465 & ~n7466 ;
  assign n7468 = n7241 | n7467 ;
  assign n7469 = n7241 & n7467 ;
  assign n7470 = n7468 & ~n7469 ;
  assign n7471 = n7127 | n7143 ;
  assign n7472 = n7127 & n7143 ;
  assign n7473 = n7471 & ~n7472 ;
  assign n7474 = n7226 | n7473 ;
  assign n7475 = n7226 & n7473 ;
  assign n7476 = n7474 & ~n7475 ;
  assign n7477 = n7181 | n7198 ;
  assign n7478 = ( n7181 & n7185 ) | ( n7181 & n7477 ) | ( n7185 & n7477 ) ;
  assign n7479 = n7476 | n7478 ;
  assign n7480 = n7476 & n7478 ;
  assign n7481 = n7479 & ~n7480 ;
  assign n7482 = n7470 & n7481 ;
  assign n7483 = n7470 | n7481 ;
  assign n7484 = ~n7482 & n7483 ;
  assign n7485 = n7460 & n7484 ;
  assign n7486 = n7460 | n7484 ;
  assign n7487 = ~n7485 & n7486 ;
  assign n7488 = n7263 | n7268 ;
  assign n7489 = ( n7263 & n7265 ) | ( n7263 & n7488 ) | ( n7265 & n7488 ) ;
  assign n7490 = n7487 | n7489 ;
  assign n7491 = n7487 & n7489 ;
  assign n7492 = n7490 & ~n7491 ;
  assign n7542 = n7279 | n7283 ;
  assign n7543 = ( n7277 & n7283 ) | ( n7277 & n7542 ) | ( n7283 & n7542 ) ;
  assign n7544 = ( n7281 & n7282 ) | ( n7281 & n7543 ) | ( n7282 & n7543 ) ;
  assign n7493 = x5 & x49 ;
  assign n7494 = x18 & x36 ;
  assign n7495 = n7493 & n7494 ;
  assign n7496 = x20 & x49 ;
  assign n7497 = n3874 & n7496 ;
  assign n7498 = n1285 & n4914 ;
  assign n7499 = n7497 | n7498 ;
  assign n7500 = x34 & n7495 ;
  assign n7501 = ( x34 & ~n7499 ) | ( x34 & n7500 ) | ( ~n7499 & n7500 ) ;
  assign n7502 = x20 & n7501 ;
  assign n7503 = ( n7493 & n7494 ) | ( n7493 & ~n7499 ) | ( n7494 & ~n7499 ) ;
  assign n7504 = ( ~n7495 & n7502 ) | ( ~n7495 & n7503 ) | ( n7502 & n7503 ) ;
  assign n7505 = n720 & n5107 ;
  assign n7506 = n647 & n5710 ;
  assign n7507 = n7505 | n7506 ;
  assign n7508 = n490 & n5407 ;
  assign n7509 = x41 & n7508 ;
  assign n7510 = ( x41 & ~n7507 ) | ( x41 & n7509 ) | ( ~n7507 & n7509 ) ;
  assign n7511 = x13 & n7510 ;
  assign n7512 = n7507 | n7508 ;
  assign n7513 = x11 & x43 ;
  assign n7514 = x12 & x42 ;
  assign n7515 = ( ~n7508 & n7513 ) | ( ~n7508 & n7514 ) | ( n7513 & n7514 ) ;
  assign n7516 = n7513 & n7514 ;
  assign n7517 = ( ~n7507 & n7515 ) | ( ~n7507 & n7516 ) | ( n7515 & n7516 ) ;
  assign n7518 = ~n7512 & n7517 ;
  assign n7519 = n7511 | n7518 ;
  assign n7520 = n7504 & n7519 ;
  assign n7521 = n7504 & ~n7520 ;
  assign n7522 = n7519 & ~n7520 ;
  assign n7523 = n7521 | n7522 ;
  assign n7524 = x17 & x48 ;
  assign n7525 = n4798 & n7524 ;
  assign n7526 = n1023 & n4857 ;
  assign n7527 = n7525 | n7526 ;
  assign n7528 = x38 & x48 ;
  assign n7529 = n623 & n7528 ;
  assign n7530 = x37 & n7529 ;
  assign n7531 = ( x37 & ~n7527 ) | ( x37 & n7530 ) | ( ~n7527 & n7530 ) ;
  assign n7532 = x17 & n7531 ;
  assign n7533 = n7527 | n7529 ;
  assign n7534 = x6 & x48 ;
  assign n7535 = x16 & x38 ;
  assign n7536 = ( ~n7529 & n7534 ) | ( ~n7529 & n7535 ) | ( n7534 & n7535 ) ;
  assign n7537 = n7534 & n7535 ;
  assign n7538 = ( ~n7527 & n7536 ) | ( ~n7527 & n7537 ) | ( n7536 & n7537 ) ;
  assign n7539 = ~n7533 & n7538 ;
  assign n7540 = n7532 | n7539 ;
  assign n7541 = ~n7523 & n7540 ;
  assign n7545 = n7541 & n7544 ;
  assign n7546 = n7523 & ~n7540 ;
  assign n7547 = ( n7544 & n7545 ) | ( n7544 & n7546 ) | ( n7545 & n7546 ) ;
  assign n7548 = n7541 | n7544 ;
  assign n7549 = n7546 | n7548 ;
  assign n7550 = ~n7547 & n7549 ;
  assign n7551 = x9 & x45 ;
  assign n7552 = n360 & n6093 ;
  assign n7553 = n5090 & n7551 ;
  assign n7554 = n7552 | n7553 ;
  assign n7555 = n6432 & n7170 ;
  assign n7556 = n7551 & n7555 ;
  assign n7557 = ( n7551 & ~n7554 ) | ( n7551 & n7556 ) | ( ~n7554 & n7556 ) ;
  assign n7558 = n7554 | n7555 ;
  assign n7559 = x10 & x44 ;
  assign n7560 = ( n5090 & ~n7555 ) | ( n5090 & n7559 ) | ( ~n7555 & n7559 ) ;
  assign n7561 = n5090 & n7559 ;
  assign n7562 = ( ~n7554 & n7560 ) | ( ~n7554 & n7561 ) | ( n7560 & n7561 ) ;
  assign n7563 = ~n7558 & n7562 ;
  assign n7564 = n7557 | n7563 ;
  assign n7565 = x50 & x52 ;
  assign n7566 = n119 & n7565 ;
  assign n7567 = x51 & x52 ;
  assign n7568 = n77 & n7567 ;
  assign n7569 = n7566 | n7568 ;
  assign n7570 = n79 & n7112 ;
  assign n7571 = x52 & n7570 ;
  assign n7572 = ( x52 & ~n7569 ) | ( x52 & n7571 ) | ( ~n7569 & n7571 ) ;
  assign n7573 = x2 & n7572 ;
  assign n7574 = n7569 | n7570 ;
  assign n7575 = x3 & x51 ;
  assign n7576 = x4 & x50 ;
  assign n7577 = ( ~n7570 & n7575 ) | ( ~n7570 & n7576 ) | ( n7575 & n7576 ) ;
  assign n7578 = n7575 & n7576 ;
  assign n7579 = ( ~n7569 & n7577 ) | ( ~n7569 & n7578 ) | ( n7577 & n7578 ) ;
  assign n7580 = ~n7574 & n7579 ;
  assign n7581 = n7573 | n7580 ;
  assign n7582 = x15 & x39 ;
  assign n7583 = x7 & x47 ;
  assign n7584 = x8 & x46 ;
  assign n7585 = ( ~n7582 & n7583 ) | ( ~n7582 & n7584 ) | ( n7583 & n7584 ) ;
  assign n7586 = n251 & n6147 ;
  assign n7587 = n7583 | n7584 ;
  assign n7588 = ( n7582 & n7586 ) | ( n7582 & n7587 ) | ( n7586 & n7587 ) ;
  assign n7589 = ( n7582 & n7585 ) | ( n7582 & ~n7588 ) | ( n7585 & ~n7588 ) ;
  assign n7590 = ( n7564 & n7581 ) | ( n7564 & ~n7589 ) | ( n7581 & ~n7589 ) ;
  assign n7591 = ( ~n7581 & n7589 ) | ( ~n7581 & n7590 ) | ( n7589 & n7590 ) ;
  assign n7592 = ( ~n7564 & n7590 ) | ( ~n7564 & n7591 ) | ( n7590 & n7591 ) ;
  assign n7593 = n7550 | n7592 ;
  assign n7594 = n7550 & n7592 ;
  assign n7595 = n7593 & ~n7594 ;
  assign n7611 = n7255 | n7259 ;
  assign n7612 = ( n7255 & n7256 ) | ( n7255 & n7611 ) | ( n7256 & n7611 ) ;
  assign n7596 = n7116 | n7172 ;
  assign n7597 = n7116 & n7172 ;
  assign n7598 = n7596 & ~n7597 ;
  assign n7599 = n7212 | n7598 ;
  assign n7600 = n7212 & n7598 ;
  assign n7601 = n7599 & ~n7600 ;
  assign n7602 = n7233 | n7248 ;
  assign n7603 = n7132 | n7150 ;
  assign n7604 = ( n7132 & n7135 ) | ( n7132 & n7603 ) | ( n7135 & n7603 ) ;
  assign n7605 = n7602 | n7604 ;
  assign n7606 = n7602 & n7604 ;
  assign n7607 = n7605 & ~n7606 ;
  assign n7608 = n7601 & n7607 ;
  assign n7609 = n7601 | n7607 ;
  assign n7610 = ~n7608 & n7609 ;
  assign n7613 = n7610 & n7612 ;
  assign n7614 = n7612 & ~n7613 ;
  assign n7615 = n7610 & ~n7612 ;
  assign n7616 = n7595 & n7615 ;
  assign n7617 = ( n7595 & n7614 ) | ( n7595 & n7616 ) | ( n7614 & n7616 ) ;
  assign n7618 = n7595 | n7615 ;
  assign n7619 = n7614 | n7618 ;
  assign n7620 = ~n7617 & n7619 ;
  assign n7621 = ~n7492 & n7620 ;
  assign n7622 = n7491 | n7620 ;
  assign n7623 = n7490 & ~n7622 ;
  assign n7624 = n7621 | n7623 ;
  assign n7625 = ~n7441 & n7442 ;
  assign n7626 = ~n7624 & n7625 ;
  assign n7627 = ( n7444 & ~n7624 ) | ( n7444 & n7626 ) | ( ~n7624 & n7626 ) ;
  assign n7628 = n7624 & ~n7625 ;
  assign n7629 = ~n7444 & n7628 ;
  assign n7630 = n7627 | n7629 ;
  assign n7631 = n7273 | n7357 ;
  assign n7632 = ( n7273 & n7275 ) | ( n7273 & n7631 ) | ( n7275 & n7631 ) ;
  assign n7633 = n7630 & n7632 ;
  assign n7634 = n7630 | n7632 ;
  assign n7635 = ~n7633 & n7634 ;
  assign n7636 = n7360 & n7362 ;
  assign n7637 = n7360 | n7362 ;
  assign n7638 = n7105 & n7637 ;
  assign n7639 = n7091 & n7637 ;
  assign n7640 = ( n7096 & n7638 ) | ( n7096 & n7639 ) | ( n7638 & n7639 ) ;
  assign n7641 = ( n7097 & n7638 ) | ( n7097 & n7639 ) | ( n7638 & n7639 ) ;
  assign n7642 = ( n6303 & n7640 ) | ( n6303 & n7641 ) | ( n7640 & n7641 ) ;
  assign n7643 = n7636 | n7642 ;
  assign n7644 = n7635 | n7643 ;
  assign n7645 = n7635 & n7643 ;
  assign n7646 = n7644 & ~n7645 ;
  assign n7647 = n7633 | n7634 ;
  assign n7648 = ( n7630 & n7632 ) | ( n7630 & n7636 ) | ( n7632 & n7636 ) ;
  assign n7649 = ( n7642 & n7647 ) | ( n7642 & n7648 ) | ( n7647 & n7648 ) ;
  assign n7703 = ( n7491 & n7492 ) | ( n7491 & n7622 ) | ( n7492 & n7622 ) ;
  assign n7650 = n7613 | n7617 ;
  assign n7692 = n7455 | n7484 ;
  assign n7693 = ( n7457 & n7484 ) | ( n7457 & n7692 ) | ( n7484 & n7692 ) ;
  assign n7694 = ( n7458 & n7460 ) | ( n7458 & n7693 ) | ( n7460 & n7693 ) ;
  assign n7651 = x9 & x46 ;
  assign n7652 = x14 & x41 ;
  assign n7653 = n7651 & n7652 ;
  assign n7654 = x40 & x46 ;
  assign n7655 = n1462 & n7654 ;
  assign n7656 = n792 & n5813 ;
  assign n7657 = n7655 | n7656 ;
  assign n7658 = x40 & n7653 ;
  assign n7659 = ( x40 & ~n7657 ) | ( x40 & n7658 ) | ( ~n7657 & n7658 ) ;
  assign n7660 = x15 & n7659 ;
  assign n7661 = ( n7651 & n7652 ) | ( n7651 & ~n7657 ) | ( n7652 & ~n7657 ) ;
  assign n7662 = ( ~n7653 & n7660 ) | ( ~n7653 & n7661 ) | ( n7660 & n7661 ) ;
  assign n7663 = x6 & x49 ;
  assign n7664 = x17 & x38 ;
  assign n7665 = n7663 | n7664 ;
  assign n7666 = x17 & x49 ;
  assign n7667 = n4854 & n7666 ;
  assign n7668 = n7665 | n7667 ;
  assign n7669 = x3 & x52 ;
  assign n7670 = ( ~n7667 & n7668 ) | ( ~n7667 & n7669 ) | ( n7668 & n7669 ) ;
  assign n7671 = ( n7667 & n7668 ) | ( n7667 & ~n7669 ) | ( n7668 & ~n7669 ) ;
  assign n7672 = ( ~n7668 & n7670 ) | ( ~n7668 & n7671 ) | ( n7670 & n7671 ) ;
  assign n7673 = n7662 & n7672 ;
  assign n7674 = n7662 & ~n7673 ;
  assign n7675 = ~n7662 & n7672 ;
  assign n7676 = n7226 | n7472 ;
  assign n7677 = ( n7472 & n7473 ) | ( n7472 & n7676 ) | ( n7473 & n7676 ) ;
  assign n7678 = n7675 | n7677 ;
  assign n7679 = n7674 | n7678 ;
  assign n7680 = n7675 & n7677 ;
  assign n7681 = ( n7674 & n7677 ) | ( n7674 & n7680 ) | ( n7677 & n7680 ) ;
  assign n7682 = n7679 & ~n7681 ;
  assign n7683 = n7601 | n7606 ;
  assign n7684 = ( n7606 & n7607 ) | ( n7606 & n7683 ) | ( n7607 & n7683 ) ;
  assign n7685 = n7682 & n7684 ;
  assign n7686 = n7682 | n7684 ;
  assign n7687 = ~n7685 & n7686 ;
  assign n7688 = ( n7470 & n7476 ) | ( n7470 & n7478 ) | ( n7476 & n7478 ) ;
  assign n7689 = n7687 | n7688 ;
  assign n7690 = n7687 & n7688 ;
  assign n7691 = n7689 & ~n7690 ;
  assign n7695 = n7691 & n7694 ;
  assign n7696 = n7694 & ~n7695 ;
  assign n7697 = n7691 & ~n7694 ;
  assign n7698 = n7650 & n7697 ;
  assign n7699 = ( n7650 & n7696 ) | ( n7650 & n7698 ) | ( n7696 & n7698 ) ;
  assign n7700 = ~n7650 & n7697 ;
  assign n7701 = ( ~n7650 & n7696 ) | ( ~n7650 & n7700 ) | ( n7696 & n7700 ) ;
  assign n7702 = ( n7650 & ~n7699 ) | ( n7650 & n7701 ) | ( ~n7699 & n7701 ) ;
  assign n7704 = n7702 & n7703 ;
  assign n7705 = n7703 & ~n7704 ;
  assign n7706 = n7702 & ~n7704 ;
  assign n7707 = n7705 | n7706 ;
  assign n7708 = n7544 | n7592 ;
  assign n7709 = n7546 | n7592 ;
  assign n7710 = ( n7545 & n7708 ) | ( n7545 & n7709 ) | ( n7708 & n7709 ) ;
  assign n7711 = ( n7547 & n7550 ) | ( n7547 & n7710 ) | ( n7550 & n7710 ) ;
  assign n7712 = n7241 | n7466 ;
  assign n7713 = ( n7466 & n7467 ) | ( n7466 & n7712 ) | ( n7467 & n7712 ) ;
  assign n7714 = n7212 | n7597 ;
  assign n7715 = ( n7597 & n7598 ) | ( n7597 & n7714 ) | ( n7598 & n7714 ) ;
  assign n7716 = n7713 | n7715 ;
  assign n7717 = n7713 & n7715 ;
  assign n7718 = n7716 & ~n7717 ;
  assign n7719 = x28 & x54 ;
  assign n7720 = x1 & n7719 ;
  assign n7721 = x1 & x54 ;
  assign n7722 = x28 | n7721 ;
  assign n7723 = ~n7720 & n7722 ;
  assign n7724 = n7379 & n7723 ;
  assign n7725 = n7723 & ~n7724 ;
  assign n7726 = n7379 & ~n7723 ;
  assign n7727 = n7512 & n7726 ;
  assign n7728 = ( n7512 & n7725 ) | ( n7512 & n7727 ) | ( n7725 & n7727 ) ;
  assign n7729 = n7512 | n7726 ;
  assign n7730 = n7725 | n7729 ;
  assign n7731 = ~n7728 & n7730 ;
  assign n7732 = ~n7718 & n7731 ;
  assign n7733 = n7717 | n7731 ;
  assign n7734 = n7716 & ~n7733 ;
  assign n7735 = n7732 | n7734 ;
  assign n7736 = n7710 & n7735 ;
  assign n7737 = n7547 & n7735 ;
  assign n7738 = ( n7550 & n7736 ) | ( n7550 & n7737 ) | ( n7736 & n7737 ) ;
  assign n7739 = n7711 & ~n7738 ;
  assign n7740 = n7558 | n7574 ;
  assign n7741 = n7558 & n7574 ;
  assign n7742 = n7740 & ~n7741 ;
  assign n7743 = n7495 | n7499 ;
  assign n7744 = n7742 | n7743 ;
  assign n7745 = n7742 & n7743 ;
  assign n7746 = n7744 & ~n7745 ;
  assign n7747 = ( n7385 & n7401 ) | ( n7385 & n7415 ) | ( n7401 & n7415 ) ;
  assign n7748 = n7746 | n7747 ;
  assign n7749 = n7746 & n7747 ;
  assign n7750 = n7748 & ~n7749 ;
  assign n7751 = n7582 & n7583 ;
  assign n7752 = n7586 | n7751 ;
  assign n7753 = n7582 & n7584 ;
  assign n7754 = n7752 | n7753 ;
  assign n7755 = n7374 | n7382 ;
  assign n7756 = ( n7374 & n7377 ) | ( n7374 & n7755 ) | ( n7377 & n7755 ) ;
  assign n7757 = n7754 | n7756 ;
  assign n7758 = n7754 & n7756 ;
  assign n7759 = n7757 & ~n7758 ;
  assign n7760 = x18 & x37 ;
  assign n7761 = x19 & x36 ;
  assign n7762 = n7760 | n7761 ;
  assign n7763 = n1077 & n3770 ;
  assign n7764 = x5 & x50 ;
  assign n7765 = ~n7763 & n7764 ;
  assign n7766 = n7762 | n7763 ;
  assign n7767 = ( n7763 & n7765 ) | ( n7763 & n7766 ) | ( n7765 & n7766 ) ;
  assign n7768 = n7762 & ~n7767 ;
  assign n7769 = ( ~n7762 & n7763 ) | ( ~n7762 & n7764 ) | ( n7763 & n7764 ) ;
  assign n7770 = n7764 & n7769 ;
  assign n7771 = n7768 | n7770 ;
  assign n7772 = ~n7759 & n7771 ;
  assign n7773 = n7759 & ~n7771 ;
  assign n7774 = n7772 | n7773 ;
  assign n7775 = n7750 & ~n7774 ;
  assign n7776 = n7774 | n7775 ;
  assign n7777 = ( ~n7750 & n7775 ) | ( ~n7750 & n7776 ) | ( n7775 & n7776 ) ;
  assign n7778 = ~n7710 & n7735 ;
  assign n7779 = ~n7547 & n7735 ;
  assign n7780 = ( ~n7550 & n7778 ) | ( ~n7550 & n7779 ) | ( n7778 & n7779 ) ;
  assign n7781 = n7777 & n7780 ;
  assign n7782 = ( n7739 & n7777 ) | ( n7739 & n7781 ) | ( n7777 & n7781 ) ;
  assign n7783 = n7777 | n7780 ;
  assign n7784 = n7739 | n7783 ;
  assign n7785 = ~n7782 & n7784 ;
  assign n7786 = n7367 | n7438 ;
  assign n7787 = ( n7366 & n7438 ) | ( n7366 & n7786 ) | ( n7438 & n7786 ) ;
  assign n7788 = n7785 & n7787 ;
  assign n7789 = n7369 & n7785 ;
  assign n7790 = ( n7370 & n7788 ) | ( n7370 & n7789 ) | ( n7788 & n7789 ) ;
  assign n7791 = n7785 | n7787 ;
  assign n7792 = n7369 | n7785 ;
  assign n7793 = ( n7370 & n7791 ) | ( n7370 & n7792 ) | ( n7791 & n7792 ) ;
  assign n7794 = ~n7790 & n7793 ;
  assign n7795 = n7394 | n7409 ;
  assign n7796 = n7394 & n7409 ;
  assign n7797 = n7795 & ~n7796 ;
  assign n7798 = n7533 | n7797 ;
  assign n7799 = n7533 & n7797 ;
  assign n7800 = n7798 & ~n7799 ;
  assign n7801 = n7520 | n7540 ;
  assign n7802 = ( n7520 & n7523 ) | ( n7520 & n7801 ) | ( n7523 & n7801 ) ;
  assign n7803 = n7581 & n7589 ;
  assign n7804 = n7581 & ~n7803 ;
  assign n7805 = n7557 & n7589 ;
  assign n7806 = ( n7563 & n7589 ) | ( n7563 & n7805 ) | ( n7589 & n7805 ) ;
  assign n7807 = ~n7581 & n7806 ;
  assign n7808 = n7803 | n7807 ;
  assign n7809 = n7564 | n7803 ;
  assign n7810 = ( n7804 & n7808 ) | ( n7804 & n7809 ) | ( n7808 & n7809 ) ;
  assign n7811 = n7802 | n7810 ;
  assign n7812 = n7802 & n7810 ;
  assign n7813 = n7811 & ~n7812 ;
  assign n7814 = n7800 & n7813 ;
  assign n7815 = n7800 | n7813 ;
  assign n7816 = ~n7814 & n7815 ;
  assign n7817 = n7423 & n7816 ;
  assign n7818 = ( n7435 & n7816 ) | ( n7435 & n7817 ) | ( n7816 & n7817 ) ;
  assign n7819 = n7423 | n7816 ;
  assign n7820 = n7435 | n7819 ;
  assign n7821 = ~n7818 & n7820 ;
  assign n7822 = n618 & n6093 ;
  assign n7823 = x13 & x45 ;
  assign n7824 = n6972 & n7823 ;
  assign n7825 = n7822 | n7824 ;
  assign n7826 = n720 & n4969 ;
  assign n7827 = x45 & n7826 ;
  assign n7828 = ( x45 & ~n7825 ) | ( x45 & n7827 ) | ( ~n7825 & n7827 ) ;
  assign n7829 = x10 & n7828 ;
  assign n7830 = n7825 | n7826 ;
  assign n7831 = x11 & x44 ;
  assign n7832 = ( n6405 & ~n7826 ) | ( n6405 & n7831 ) | ( ~n7826 & n7831 ) ;
  assign n7833 = n6405 & n7831 ;
  assign n7834 = ( ~n7825 & n7832 ) | ( ~n7825 & n7833 ) | ( n7832 & n7833 ) ;
  assign n7835 = ~n7830 & n7834 ;
  assign n7836 = n7829 | n7835 ;
  assign n7837 = x26 & x29 ;
  assign n7838 = n2372 | n7837 ;
  assign n7839 = x12 & x43 ;
  assign n7840 = ( n2372 & n7837 ) | ( n2372 & n7839 ) | ( n7837 & n7839 ) ;
  assign n7841 = n7838 & ~n7840 ;
  assign n7842 = n2372 & n7837 ;
  assign n7843 = n7839 & ~n7842 ;
  assign n7844 = ~n7838 & n7839 ;
  assign n7845 = ( n7839 & ~n7843 ) | ( n7839 & n7844 ) | ( ~n7843 & n7844 ) ;
  assign n7846 = n7841 | n7845 ;
  assign n7847 = n7836 & n7846 ;
  assign n7848 = n7836 & ~n7847 ;
  assign n7849 = x7 & x48 ;
  assign n7850 = x8 & x47 ;
  assign n7851 = n7849 | n7850 ;
  assign n7852 = n251 & n6762 ;
  assign n7853 = x16 & x39 ;
  assign n7854 = ~n7852 & n7853 ;
  assign n7855 = n7851 | n7852 ;
  assign n7856 = ( n7852 & n7854 ) | ( n7852 & n7855 ) | ( n7854 & n7855 ) ;
  assign n7857 = n7851 & ~n7856 ;
  assign n7858 = ( ~n7851 & n7852 ) | ( ~n7851 & n7853 ) | ( n7852 & n7853 ) ;
  assign n7859 = n7853 & n7858 ;
  assign n7860 = n7857 | n7859 ;
  assign n7861 = ~n7836 & n7846 ;
  assign n7862 = n7860 & ~n7861 ;
  assign n7863 = ~n7848 & n7862 ;
  assign n7864 = ~n7860 & n7861 ;
  assign n7865 = ( n7848 & ~n7860 ) | ( n7848 & n7864 ) | ( ~n7860 & n7864 ) ;
  assign n7866 = n7863 | n7865 ;
  assign n7867 = ( n7445 & n7447 ) | ( n7445 & n7452 ) | ( n7447 & n7452 ) ;
  assign n7868 = n7866 | n7867 ;
  assign n7869 = n7866 & n7867 ;
  assign n7870 = n7868 & ~n7869 ;
  assign n7871 = x51 & n82 ;
  assign n7872 = x53 & n67 ;
  assign n7873 = n7871 | n7872 ;
  assign n7874 = x51 & x53 ;
  assign n7875 = n119 & n7874 ;
  assign n7876 = x55 & ~n7875 ;
  assign n7877 = n7873 & n7876 ;
  assign n7878 = x0 & x55 ;
  assign n7879 = ~n7877 & n7878 ;
  assign n7880 = n7875 | n7877 ;
  assign n7881 = x2 & x53 ;
  assign n7882 = x4 & x51 ;
  assign n7883 = ( ~n7875 & n7881 ) | ( ~n7875 & n7882 ) | ( n7881 & n7882 ) ;
  assign n7884 = n7881 & n7882 ;
  assign n7885 = ( ~n7877 & n7883 ) | ( ~n7877 & n7884 ) | ( n7883 & n7884 ) ;
  assign n7886 = ~n7880 & n7885 ;
  assign n7887 = n7879 | n7886 ;
  assign n7888 = n1710 & n3129 ;
  assign n7889 = n1434 & n3483 ;
  assign n7890 = n7888 | n7889 ;
  assign n7891 = n1585 & n4530 ;
  assign n7892 = x35 & n7891 ;
  assign n7893 = ( x35 & ~n7890 ) | ( x35 & n7892 ) | ( ~n7890 & n7892 ) ;
  assign n7894 = x20 & n7893 ;
  assign n7895 = n7890 | n7891 ;
  assign n7896 = x21 & x34 ;
  assign n7897 = ( n2686 & ~n7891 ) | ( n2686 & n7896 ) | ( ~n7891 & n7896 ) ;
  assign n7898 = n2686 & n7896 ;
  assign n7899 = ( ~n7890 & n7897 ) | ( ~n7890 & n7898 ) | ( n7897 & n7898 ) ;
  assign n7900 = ~n7895 & n7899 ;
  assign n7901 = n7894 | n7900 ;
  assign n7902 = n7887 & n7901 ;
  assign n7903 = n7887 & ~n7902 ;
  assign n7904 = x23 & x32 ;
  assign n7905 = n1557 & n2546 ;
  assign n7906 = n1686 & n4062 ;
  assign n7907 = n7905 | n7906 ;
  assign n7908 = n1912 & n2965 ;
  assign n7909 = n7904 & n7908 ;
  assign n7910 = ( n7904 & ~n7907 ) | ( n7904 & n7909 ) | ( ~n7907 & n7909 ) ;
  assign n7911 = n7907 | n7908 ;
  assign n7912 = x24 & x31 ;
  assign n7913 = x25 & x30 ;
  assign n7914 = ( ~n7908 & n7912 ) | ( ~n7908 & n7913 ) | ( n7912 & n7913 ) ;
  assign n7915 = n7912 & n7913 ;
  assign n7916 = ( ~n7907 & n7914 ) | ( ~n7907 & n7915 ) | ( n7914 & n7915 ) ;
  assign n7917 = ~n7911 & n7916 ;
  assign n7918 = n7910 | n7917 ;
  assign n7919 = ~n7901 & n7918 ;
  assign n7920 = ( n7887 & n7918 ) | ( n7887 & n7919 ) | ( n7918 & n7919 ) ;
  assign n7921 = ~n7903 & n7920 ;
  assign n7922 = n7901 & ~n7918 ;
  assign n7923 = ~n7887 & n7922 ;
  assign n7924 = ( n7903 & ~n7918 ) | ( n7903 & n7923 ) | ( ~n7918 & n7923 ) ;
  assign n7925 = n7921 | n7924 ;
  assign n7926 = n7870 & n7925 ;
  assign n7927 = n7870 | n7925 ;
  assign n7928 = ~n7926 & n7927 ;
  assign n7929 = ~n7821 & n7928 ;
  assign n7930 = n7821 & ~n7928 ;
  assign n7931 = n7929 | n7930 ;
  assign n7932 = n7794 | n7931 ;
  assign n7933 = n7794 & n7931 ;
  assign n7934 = n7932 & ~n7933 ;
  assign n7935 = n7707 & n7934 ;
  assign n7936 = n7707 | n7934 ;
  assign n7937 = ~n7935 & n7936 ;
  assign n7938 = ( n7441 & n7442 ) | ( n7441 & n7624 ) | ( n7442 & n7624 ) ;
  assign n7939 = ( n7649 & n7937 ) | ( n7649 & ~n7938 ) | ( n7937 & ~n7938 ) ;
  assign n7940 = ( ~n7937 & n7938 ) | ( ~n7937 & n7939 ) | ( n7938 & n7939 ) ;
  assign n7941 = ( ~n7649 & n7939 ) | ( ~n7649 & n7940 ) | ( n7939 & n7940 ) ;
  assign n8235 = n7937 & n7938 ;
  assign n8236 = n7937 | n7938 ;
  assign n8237 = n8235 | n8236 ;
  assign n8238 = ( n7648 & n8235 ) | ( n7648 & n8237 ) | ( n8235 & n8237 ) ;
  assign n8239 = ( n7647 & n8235 ) | ( n7647 & n8237 ) | ( n8235 & n8237 ) ;
  assign n8240 = ( n7640 & n8238 ) | ( n7640 & n8239 ) | ( n8238 & n8239 ) ;
  assign n8241 = ( n7641 & n8238 ) | ( n7641 & n8239 ) | ( n8238 & n8239 ) ;
  assign n8242 = ( n6303 & n8240 ) | ( n6303 & n8241 ) | ( n8240 & n8241 ) ;
  assign n7990 = n7790 | n7931 ;
  assign n7991 = ( n7790 & n7794 ) | ( n7790 & n7990 ) | ( n7794 & n7990 ) ;
  assign n7942 = n7724 | n7728 ;
  assign n7943 = x5 & x51 ;
  assign n7944 = x18 & x38 ;
  assign n7945 = n7943 | n7944 ;
  assign n7946 = x38 & x51 ;
  assign n7947 = n1292 & n7946 ;
  assign n7948 = x21 & x35 ;
  assign n7949 = ~n7947 & n7948 ;
  assign n7950 = n7945 | n7947 ;
  assign n7951 = ( n7947 & n7949 ) | ( n7947 & n7950 ) | ( n7949 & n7950 ) ;
  assign n7952 = n7945 & ~n7951 ;
  assign n7953 = ( ~n7945 & n7947 ) | ( ~n7945 & n7948 ) | ( n7947 & n7948 ) ;
  assign n7954 = n7948 & n7953 ;
  assign n7955 = n7952 | n7954 ;
  assign n7956 = n7942 & n7955 ;
  assign n7957 = n7942 & ~n7956 ;
  assign n7959 = n7741 | n7743 ;
  assign n7960 = ( n7741 & n7742 ) | ( n7741 & n7959 ) | ( n7742 & n7959 ) ;
  assign n7958 = ~n7942 & n7955 ;
  assign n7961 = n7958 & n7960 ;
  assign n7962 = ( n7957 & n7960 ) | ( n7957 & n7961 ) | ( n7960 & n7961 ) ;
  assign n7963 = n7958 | n7960 ;
  assign n7964 = n7957 | n7963 ;
  assign n7965 = ~n7962 & n7964 ;
  assign n7966 = n7800 | n7810 ;
  assign n7967 = ( n7800 & n7802 ) | ( n7800 & n7966 ) | ( n7802 & n7966 ) ;
  assign n7968 = n7965 & n7967 ;
  assign n7969 = n7812 & n7965 ;
  assign n7970 = ( n7813 & n7968 ) | ( n7813 & n7969 ) | ( n7968 & n7969 ) ;
  assign n7971 = n7965 | n7967 ;
  assign n7972 = n7812 | n7965 ;
  assign n7973 = ( n7813 & n7971 ) | ( n7813 & n7972 ) | ( n7971 & n7972 ) ;
  assign n7974 = ~n7970 & n7973 ;
  assign n7975 = n7750 & n7774 ;
  assign n7976 = n7749 | n7975 ;
  assign n7977 = n7974 | n7976 ;
  assign n7978 = n7974 & n7976 ;
  assign n7979 = n7977 & ~n7978 ;
  assign n7980 = n7738 | n7979 ;
  assign n7981 = n7782 | n7980 ;
  assign n7982 = n7738 & n7979 ;
  assign n7983 = ( n7782 & n7979 ) | ( n7782 & n7982 ) | ( n7979 & n7982 ) ;
  assign n7984 = n7981 & ~n7983 ;
  assign n7985 = n7818 | n7928 ;
  assign n7986 = ( n7818 & n7821 ) | ( n7818 & n7985 ) | ( n7821 & n7985 ) ;
  assign n7987 = n7984 | n7986 ;
  assign n7988 = n7984 & n7986 ;
  assign n7989 = n7987 & ~n7988 ;
  assign n7992 = n7989 & n7991 ;
  assign n7993 = n7991 & ~n7992 ;
  assign n7994 = n7989 & ~n7991 ;
  assign n7995 = n7993 | n7994 ;
  assign n7996 = n7758 | n7771 ;
  assign n7997 = ( n7758 & n7759 ) | ( n7758 & n7996 ) | ( n7759 & n7996 ) ;
  assign n7998 = n7533 | n7796 ;
  assign n7999 = ( n7796 & n7797 ) | ( n7796 & n7998 ) | ( n7797 & n7998 ) ;
  assign n8000 = n7997 | n7999 ;
  assign n8001 = n7997 & n7999 ;
  assign n8002 = n8000 & ~n8001 ;
  assign n8003 = n7901 & n7918 ;
  assign n8004 = ~n7887 & n8003 ;
  assign n8005 = n7902 | n8004 ;
  assign n8006 = n7902 | n7918 ;
  assign n8007 = ( n7903 & n8005 ) | ( n7903 & n8006 ) | ( n8005 & n8006 ) ;
  assign n8008 = n8002 | n8007 ;
  assign n8009 = n8002 & n8007 ;
  assign n8010 = n8008 & ~n8009 ;
  assign n8011 = n7869 | n7925 ;
  assign n8012 = ( n7869 & n7870 ) | ( n7869 & n8011 ) | ( n7870 & n8011 ) ;
  assign n8013 = n8010 & ~n8012 ;
  assign n8014 = n7767 | n7880 ;
  assign n8015 = n7767 & n7880 ;
  assign n8016 = n8014 & ~n8015 ;
  assign n8017 = n7653 | n7657 ;
  assign n8018 = n8016 | n8017 ;
  assign n8019 = n8016 & n8017 ;
  assign n8020 = n8018 & ~n8019 ;
  assign n8021 = n7673 | n7681 ;
  assign n8022 = n8020 | n8021 ;
  assign n8023 = n8020 & n8021 ;
  assign n8024 = n8022 & ~n8023 ;
  assign n8025 = ( n7717 & n7718 ) | ( n7717 & n7733 ) | ( n7718 & n7733 ) ;
  assign n8026 = n8024 | n8025 ;
  assign n8027 = n8024 & n8025 ;
  assign n8028 = n8026 & ~n8027 ;
  assign n8029 = ( n8012 & n8013 ) | ( n8012 & n8028 ) | ( n8013 & n8028 ) ;
  assign n8030 = ( ~n8010 & n8013 ) | ( ~n8010 & n8029 ) | ( n8013 & n8029 ) ;
  assign n8031 = n8010 & n8012 ;
  assign n8032 = n8012 & ~n8031 ;
  assign n8033 = n8013 | n8028 ;
  assign n8034 = n8032 | n8033 ;
  assign n8035 = ~n8030 & n8034 ;
  assign n8036 = n7695 & n8035 ;
  assign n8037 = ( n7699 & n8035 ) | ( n7699 & n8036 ) | ( n8035 & n8036 ) ;
  assign n8038 = n7695 | n7699 ;
  assign n8039 = ~n8037 & n8038 ;
  assign n8040 = x7 & x49 ;
  assign n8041 = x17 & x39 ;
  assign n8042 = n8040 & n8041 ;
  assign n8043 = n200 & n6834 ;
  assign n8044 = x17 & x50 ;
  assign n8045 = n5231 & n8044 ;
  assign n8046 = n8043 | n8045 ;
  assign n8047 = x50 & n8042 ;
  assign n8048 = ( x50 & ~n8046 ) | ( x50 & n8047 ) | ( ~n8046 & n8047 ) ;
  assign n8049 = x6 & n8048 ;
  assign n8050 = ( n8040 & n8041 ) | ( n8040 & ~n8046 ) | ( n8041 & ~n8046 ) ;
  assign n8051 = ( ~n8042 & n8049 ) | ( ~n8042 & n8050 ) | ( n8049 & n8050 ) ;
  assign n8052 = n720 & n5104 ;
  assign n8053 = n490 & n6093 ;
  assign n8054 = n8052 | n8053 ;
  assign n8055 = n647 & n5658 ;
  assign n8056 = x45 & n8055 ;
  assign n8057 = ( x45 & ~n8054 ) | ( x45 & n8056 ) | ( ~n8054 & n8056 ) ;
  assign n8058 = x11 & n8057 ;
  assign n8059 = n8054 | n8055 ;
  assign n8060 = x12 & x44 ;
  assign n8061 = ( n6656 & ~n8055 ) | ( n6656 & n8060 ) | ( ~n8055 & n8060 ) ;
  assign n8062 = n6656 & n8060 ;
  assign n8063 = ( ~n8054 & n8061 ) | ( ~n8054 & n8062 ) | ( n8061 & n8062 ) ;
  assign n8064 = ~n8059 & n8063 ;
  assign n8065 = n8058 | n8064 ;
  assign n8066 = n8051 & n8065 ;
  assign n8067 = n8051 & ~n8066 ;
  assign n8068 = n8065 & ~n8066 ;
  assign n8069 = n8067 | n8068 ;
  assign n8070 = x40 & x48 ;
  assign n8071 = n1454 & n8070 ;
  assign n8072 = n795 & n5813 ;
  assign n8073 = n8071 | n8072 ;
  assign n8074 = x15 & x48 ;
  assign n8075 = n6049 & n8074 ;
  assign n8076 = n4553 & n8075 ;
  assign n8077 = ( n4553 & ~n8073 ) | ( n4553 & n8076 ) | ( ~n8073 & n8076 ) ;
  assign n8078 = n8073 | n8075 ;
  assign n8079 = x8 & x48 ;
  assign n8080 = x15 & x41 ;
  assign n8081 = ( ~n8075 & n8079 ) | ( ~n8075 & n8080 ) | ( n8079 & n8080 ) ;
  assign n8082 = n8079 & n8080 ;
  assign n8083 = ( ~n8073 & n8081 ) | ( ~n8073 & n8082 ) | ( n8081 & n8082 ) ;
  assign n8084 = ~n8078 & n8083 ;
  assign n8085 = n8077 | n8084 ;
  assign n8086 = ~n8069 & n8085 ;
  assign n8087 = n8069 & ~n8085 ;
  assign n8088 = n8086 | n8087 ;
  assign n8089 = n1710 & n4914 ;
  assign n8090 = x33 & x36 ;
  assign n8091 = n4735 & n8090 ;
  assign n8092 = n8089 | n8091 ;
  assign n8093 = n1932 & n4530 ;
  assign n8094 = x36 & n8093 ;
  assign n8095 = ( x36 & ~n8092 ) | ( x36 & n8094 ) | ( ~n8092 & n8094 ) ;
  assign n8096 = x20 & n8095 ;
  assign n8097 = n8092 | n8093 ;
  assign n8098 = x22 & x34 ;
  assign n8099 = x23 & x33 ;
  assign n8100 = ( ~n8093 & n8098 ) | ( ~n8093 & n8099 ) | ( n8098 & n8099 ) ;
  assign n8101 = n8098 & n8099 ;
  assign n8102 = ( ~n8092 & n8100 ) | ( ~n8092 & n8101 ) | ( n8100 & n8101 ) ;
  assign n8103 = ~n8097 & n8102 ;
  assign n8104 = n8096 | n8103 ;
  assign n8105 = n2340 & n2546 ;
  assign n8106 = n1912 & n4062 ;
  assign n8107 = n8105 | n8106 ;
  assign n8108 = n2511 & n2965 ;
  assign n8109 = x32 & n8108 ;
  assign n8110 = ( x32 & ~n8107 ) | ( x32 & n8109 ) | ( ~n8107 & n8109 ) ;
  assign n8111 = x24 & n8110 ;
  assign n8112 = n8107 | n8108 ;
  assign n8113 = x25 & x31 ;
  assign n8114 = x26 & x30 ;
  assign n8115 = ( ~n8108 & n8113 ) | ( ~n8108 & n8114 ) | ( n8113 & n8114 ) ;
  assign n8116 = n8113 & n8114 ;
  assign n8117 = ( ~n8107 & n8115 ) | ( ~n8107 & n8116 ) | ( n8115 & n8116 ) ;
  assign n8118 = ~n8112 & n8117 ;
  assign n8119 = n8111 | n8118 ;
  assign n8120 = n8104 & n8119 ;
  assign n8121 = n8104 & ~n8120 ;
  assign n8122 = n8119 & ~n8120 ;
  assign n8123 = n8121 | n8122 ;
  assign n8124 = n360 & n6147 ;
  assign n8125 = x14 & x47 ;
  assign n8126 = n6669 & n8125 ;
  assign n8127 = n8124 | n8126 ;
  assign n8128 = x14 & x46 ;
  assign n8129 = n6972 & n8128 ;
  assign n8130 = x47 & n8129 ;
  assign n8131 = ( x47 & ~n8127 ) | ( x47 & n8130 ) | ( ~n8127 & n8130 ) ;
  assign n8132 = x9 & n8131 ;
  assign n8133 = n8127 | n8129 ;
  assign n8134 = x10 & x46 ;
  assign n8135 = ( n5712 & ~n8129 ) | ( n5712 & n8134 ) | ( ~n8129 & n8134 ) ;
  assign n8136 = n5712 & n8134 ;
  assign n8137 = ( ~n8127 & n8135 ) | ( ~n8127 & n8136 ) | ( n8135 & n8136 ) ;
  assign n8138 = ~n8133 & n8137 ;
  assign n8139 = n8132 | n8138 ;
  assign n8140 = ~n8123 & n8139 ;
  assign n8141 = n8123 & ~n8139 ;
  assign n8142 = n8140 | n8141 ;
  assign n8143 = n8088 & ~n8142 ;
  assign n8144 = ~n8088 & n8142 ;
  assign n8145 = n8143 | n8144 ;
  assign n8146 = x54 & x56 ;
  assign n8147 = n67 & n8146 ;
  assign n8148 = x0 & x56 ;
  assign n8149 = x2 & x54 ;
  assign n8150 = n8148 | n8149 ;
  assign n8151 = ~n8147 & n8150 ;
  assign n8152 = n7720 & n8151 ;
  assign n8153 = n7720 | n8151 ;
  assign n8154 = ~n8152 & n8153 ;
  assign n8155 = n7856 & n8154 ;
  assign n8156 = n7856 | n8154 ;
  assign n8157 = ~n8155 & n8156 ;
  assign n8158 = x4 & x52 ;
  assign n8159 = x19 & x37 ;
  assign n8160 = n8158 & n8159 ;
  assign n8161 = x52 & x53 ;
  assign n8162 = n79 & n8161 ;
  assign n8163 = x37 & x53 ;
  assign n8164 = n1211 & n8163 ;
  assign n8165 = n8162 | n8164 ;
  assign n8166 = x53 & n8160 ;
  assign n8167 = ( x53 & ~n8165 ) | ( x53 & n8166 ) | ( ~n8165 & n8166 ) ;
  assign n8168 = x3 & n8167 ;
  assign n8169 = ( n8158 & n8159 ) | ( n8158 & ~n8165 ) | ( n8159 & ~n8165 ) ;
  assign n8170 = ( ~n8160 & n8168 ) | ( ~n8160 & n8169 ) | ( n8168 & n8169 ) ;
  assign n8171 = n8157 & ~n8170 ;
  assign n8172 = n8157 | n8170 ;
  assign n8173 = ( ~n8157 & n8171 ) | ( ~n8157 & n8172 ) | ( n8171 & n8172 ) ;
  assign n8174 = n8145 | n8173 ;
  assign n8175 = n8145 & n8173 ;
  assign n8176 = n8174 & ~n8175 ;
  assign n8177 = n7682 | n7688 ;
  assign n8178 = ( n7684 & n7688 ) | ( n7684 & n8177 ) | ( n7688 & n8177 ) ;
  assign n8179 = ( n7685 & n7687 ) | ( n7685 & n8178 ) | ( n7687 & n8178 ) ;
  assign n8180 = ~n7667 & n7669 ;
  assign n8181 = ( n7667 & n7668 ) | ( n7667 & n8180 ) | ( n7668 & n8180 ) ;
  assign n8182 = n7895 | n7911 ;
  assign n8183 = n7895 & n7911 ;
  assign n8184 = n8182 & ~n8183 ;
  assign n8185 = n8181 | n8184 ;
  assign n8186 = n8181 & n8184 ;
  assign n8187 = n8185 & ~n8186 ;
  assign n8188 = x1 & x55 ;
  assign n8189 = n2075 | n8188 ;
  assign n8190 = n2075 & n8188 ;
  assign n8191 = n8189 & ~n8190 ;
  assign n8192 = n7840 | n8190 ;
  assign n8193 = ( n8190 & n8191 ) | ( n8190 & n8192 ) | ( n8191 & n8192 ) ;
  assign n8194 = n8189 & ~n8193 ;
  assign n8195 = n7840 & ~n8191 ;
  assign n8196 = n7830 & n8195 ;
  assign n8197 = ( n7830 & n8194 ) | ( n7830 & n8196 ) | ( n8194 & n8196 ) ;
  assign n8198 = ( n7830 & n8189 ) | ( n7830 & ~n8193 ) | ( n8189 & ~n8193 ) ;
  assign n8199 = n7830 | n8195 ;
  assign n8200 = n8198 | n8199 ;
  assign n8201 = ~n8197 & n8200 ;
  assign n8202 = n7860 & n7861 ;
  assign n8203 = ( n7848 & n7860 ) | ( n7848 & n8202 ) | ( n7860 & n8202 ) ;
  assign n8204 = n7847 & n8201 ;
  assign n8205 = ( n8201 & n8203 ) | ( n8201 & n8204 ) | ( n8203 & n8204 ) ;
  assign n8206 = n7847 | n8201 ;
  assign n8207 = n8203 | n8206 ;
  assign n8208 = ~n8205 & n8207 ;
  assign n8209 = n8187 & n8208 ;
  assign n8210 = n8187 | n8208 ;
  assign n8211 = ~n8209 & n8210 ;
  assign n8212 = n8178 & n8211 ;
  assign n8213 = n7685 & n8211 ;
  assign n8214 = ( n7687 & n8212 ) | ( n7687 & n8213 ) | ( n8212 & n8213 ) ;
  assign n8215 = n8179 & ~n8214 ;
  assign n8216 = ~n8178 & n8211 ;
  assign n8217 = ~n7685 & n8211 ;
  assign n8218 = ( ~n7687 & n8216 ) | ( ~n7687 & n8217 ) | ( n8216 & n8217 ) ;
  assign n8219 = n8176 & n8218 ;
  assign n8220 = ( n8176 & n8215 ) | ( n8176 & n8219 ) | ( n8215 & n8219 ) ;
  assign n8221 = n8176 | n8218 ;
  assign n8222 = n8215 | n8221 ;
  assign n8223 = ~n8220 & n8222 ;
  assign n8224 = ~n7695 & n8035 ;
  assign n8225 = n8223 & n8224 ;
  assign n8226 = ~n7699 & n8225 ;
  assign n8227 = ( n8039 & n8223 ) | ( n8039 & n8226 ) | ( n8223 & n8226 ) ;
  assign n8228 = n8223 | n8224 ;
  assign n8229 = ( ~n7699 & n8223 ) | ( ~n7699 & n8228 ) | ( n8223 & n8228 ) ;
  assign n8230 = n8039 | n8229 ;
  assign n8231 = ~n8227 & n8230 ;
  assign n8232 = n7995 & n8231 ;
  assign n8233 = n7995 | n8231 ;
  assign n8234 = ~n8232 & n8233 ;
  assign n8243 = n7704 | n7934 ;
  assign n8244 = ( n7704 & n7707 ) | ( n7704 & n8243 ) | ( n7707 & n8243 ) ;
  assign n8245 = ( n8234 & n8242 ) | ( n8234 & ~n8244 ) | ( n8242 & ~n8244 ) ;
  assign n8246 = ( ~n8234 & n8244 ) | ( ~n8234 & n8245 ) | ( n8244 & n8245 ) ;
  assign n8247 = ( ~n8242 & n8245 ) | ( ~n8242 & n8246 ) | ( n8245 & n8246 ) ;
  assign n8248 = n8234 & n8244 ;
  assign n8249 = n8234 | n8244 ;
  assign n8250 = n8241 & n8249 ;
  assign n8251 = n8240 & n8249 ;
  assign n8252 = ( n6303 & n8250 ) | ( n6303 & n8251 ) | ( n8250 & n8251 ) ;
  assign n8253 = n8248 | n8252 ;
  assign n8254 = n8214 | n8220 ;
  assign n8255 = ( n7847 & n8187 ) | ( n7847 & n8201 ) | ( n8187 & n8201 ) ;
  assign n8256 = n8187 | n8201 ;
  assign n8257 = ( n8203 & n8255 ) | ( n8203 & n8256 ) | ( n8255 & n8256 ) ;
  assign n8258 = n8023 | n8025 ;
  assign n8259 = ( n8023 & n8024 ) | ( n8023 & n8258 ) | ( n8024 & n8258 ) ;
  assign n8260 = n8257 | n8259 ;
  assign n8261 = n8257 & n8259 ;
  assign n8262 = n8260 & ~n8261 ;
  assign n8263 = x0 & x57 ;
  assign n8264 = n8190 & n8263 ;
  assign n8265 = n8190 & ~n8264 ;
  assign n8266 = ~n8190 & n8263 ;
  assign n8267 = x1 & x56 ;
  assign n8268 = x29 & n8267 ;
  assign n8269 = x29 & ~n8267 ;
  assign n8270 = ( n8267 & ~n8268 ) | ( n8267 & n8269 ) | ( ~n8268 & n8269 ) ;
  assign n8271 = ~n8266 & n8270 ;
  assign n8272 = ~n8265 & n8271 ;
  assign n8273 = n8266 & ~n8270 ;
  assign n8274 = ( n8265 & ~n8270 ) | ( n8265 & n8273 ) | ( ~n8270 & n8273 ) ;
  assign n8275 = n8272 | n8274 ;
  assign n8276 = n8181 | n8183 ;
  assign n8277 = ( n8183 & n8184 ) | ( n8183 & n8276 ) | ( n8184 & n8276 ) ;
  assign n8278 = n8275 | n8277 ;
  assign n8279 = n8275 & n8277 ;
  assign n8280 = n8278 & ~n8279 ;
  assign n8281 = ( n7767 & n7880 ) | ( n7767 & n8017 ) | ( n7880 & n8017 ) ;
  assign n8282 = n8280 | n8281 ;
  assign n8283 = n8280 & n8281 ;
  assign n8284 = n8282 & ~n8283 ;
  assign n8285 = n8262 & n8284 ;
  assign n8286 = n8262 | n8284 ;
  assign n8287 = ~n8285 & n8286 ;
  assign n8288 = n8031 & n8287 ;
  assign n8289 = ( n8030 & n8287 ) | ( n8030 & n8288 ) | ( n8287 & n8288 ) ;
  assign n8290 = n8013 | n8031 ;
  assign n8291 = n8010 & ~n8031 ;
  assign n8292 = ( n8029 & n8290 ) | ( n8029 & ~n8291 ) | ( n8290 & ~n8291 ) ;
  assign n8293 = n8287 | n8292 ;
  assign n8294 = ~n8289 & n8293 ;
  assign n8295 = n8254 & n8294 ;
  assign n8296 = n8254 | n8294 ;
  assign n8297 = ~n8295 & n8296 ;
  assign n8298 = n8037 & n8297 ;
  assign n8299 = ( n8227 & n8297 ) | ( n8227 & n8298 ) | ( n8297 & n8298 ) ;
  assign n8300 = n8037 | n8226 ;
  assign n8301 = n8037 | n8223 ;
  assign n8302 = ( n8039 & n8300 ) | ( n8039 & n8301 ) | ( n8300 & n8301 ) ;
  assign n8303 = ~n8299 & n8302 ;
  assign n8304 = n8297 & ~n8298 ;
  assign n8305 = ~n8227 & n8304 ;
  assign n8306 = n8303 | n8305 ;
  assign n8307 = n7840 & n8191 ;
  assign n8308 = n8197 | n8307 ;
  assign n8309 = n8155 | n8170 ;
  assign n8310 = ( n8155 & n8157 ) | ( n8155 & n8309 ) | ( n8157 & n8309 ) ;
  assign n8311 = n8308 | n8310 ;
  assign n8312 = n8308 & n8310 ;
  assign n8313 = n8311 & ~n8312 ;
  assign n8314 = n8120 | n8139 ;
  assign n8315 = ( n8120 & n8123 ) | ( n8120 & n8314 ) | ( n8123 & n8314 ) ;
  assign n8316 = n8313 | n8315 ;
  assign n8317 = n8313 & n8315 ;
  assign n8318 = n8316 & ~n8317 ;
  assign n8319 = ( n8088 & n8142 ) | ( n8088 & n8173 ) | ( n8142 & n8173 ) ;
  assign n8320 = n8318 | n8319 ;
  assign n8321 = n8318 & n8319 ;
  assign n8322 = n8320 & ~n8321 ;
  assign n8323 = n8078 | n8112 ;
  assign n8324 = n8078 & n8112 ;
  assign n8325 = n8323 & ~n8324 ;
  assign n8326 = n8042 | n8046 ;
  assign n8327 = n8325 | n8326 ;
  assign n8328 = n8325 & n8326 ;
  assign n8329 = n8327 & ~n8328 ;
  assign n8330 = n8160 | n8165 ;
  assign n8331 = n8097 | n8330 ;
  assign n8332 = n8097 & n8330 ;
  assign n8333 = n8331 & ~n8332 ;
  assign n8334 = n7720 | n8147 ;
  assign n8335 = ( n8147 & n8151 ) | ( n8147 & n8334 ) | ( n8151 & n8334 ) ;
  assign n8336 = n8333 | n8335 ;
  assign n8337 = n8333 & n8335 ;
  assign n8338 = n8336 & ~n8337 ;
  assign n8339 = n8329 & n8338 ;
  assign n8340 = n8329 | n8338 ;
  assign n8341 = ~n8339 & n8340 ;
  assign n8342 = n8066 | n8085 ;
  assign n8343 = ( n8066 & n8069 ) | ( n8066 & n8342 ) | ( n8069 & n8342 ) ;
  assign n8344 = n8341 & n8343 ;
  assign n8345 = n8341 | n8343 ;
  assign n8346 = ~n8344 & n8345 ;
  assign n8347 = n8322 & n8346 ;
  assign n8348 = n8322 | n8346 ;
  assign n8349 = ~n8347 & n8348 ;
  assign n8350 = n7983 | n7986 ;
  assign n8351 = ( n7983 & n7984 ) | ( n7983 & n8350 ) | ( n7984 & n8350 ) ;
  assign n8352 = n8349 | n8351 ;
  assign n8353 = n8349 & n8351 ;
  assign n8354 = n8352 & ~n8353 ;
  assign n8355 = x53 & x54 ;
  assign n8356 = n79 & n8355 ;
  assign n8357 = x54 & x55 ;
  assign n8358 = n77 & n8357 ;
  assign n8359 = n8356 | n8358 ;
  assign n8360 = x53 & x55 ;
  assign n8361 = n119 & n8360 ;
  assign n8362 = x54 & n8361 ;
  assign n8363 = ( x54 & ~n8359 ) | ( x54 & n8362 ) | ( ~n8359 & n8362 ) ;
  assign n8364 = x3 & n8363 ;
  assign n8365 = n8359 | n8361 ;
  assign n8366 = x2 & x55 ;
  assign n8367 = x4 & x53 ;
  assign n8368 = ( ~n8361 & n8366 ) | ( ~n8361 & n8367 ) | ( n8366 & n8367 ) ;
  assign n8369 = n8366 & n8367 ;
  assign n8370 = ( ~n8359 & n8368 ) | ( ~n8359 & n8369 ) | ( n8368 & n8369 ) ;
  assign n8371 = ~n8365 & n8370 ;
  assign n8372 = n8364 | n8371 ;
  assign n8373 = x19 & x38 ;
  assign n8374 = x20 & x37 ;
  assign n8375 = n8373 | n8374 ;
  assign n8376 = n1437 & n4857 ;
  assign n8377 = x5 & x52 ;
  assign n8378 = ~n8376 & n8377 ;
  assign n8379 = n8375 | n8376 ;
  assign n8380 = ( n8376 & n8378 ) | ( n8376 & n8379 ) | ( n8378 & n8379 ) ;
  assign n8381 = n8375 & ~n8380 ;
  assign n8382 = ( ~n8375 & n8376 ) | ( ~n8375 & n8377 ) | ( n8376 & n8377 ) ;
  assign n8383 = n8377 & n8382 ;
  assign n8384 = n8381 | n8383 ;
  assign n8385 = n8372 & n8384 ;
  assign n8386 = n8372 & ~n8385 ;
  assign n8387 = n8384 & ~n8385 ;
  assign n8388 = n8386 | n8387 ;
  assign n8389 = x9 & x48 ;
  assign n8390 = x10 & x47 ;
  assign n8391 = n8389 | n8390 ;
  assign n8392 = n360 & n6762 ;
  assign n8393 = x15 & x42 ;
  assign n8394 = ~n8392 & n8393 ;
  assign n8395 = n8391 | n8392 ;
  assign n8396 = ( n8392 & n8394 ) | ( n8392 & n8395 ) | ( n8394 & n8395 ) ;
  assign n8397 = n8391 & ~n8396 ;
  assign n8398 = ( ~n8391 & n8392 ) | ( ~n8391 & n8393 ) | ( n8392 & n8393 ) ;
  assign n8399 = n8393 & n8398 ;
  assign n8400 = n8397 | n8399 ;
  assign n8401 = ~n8388 & n8400 ;
  assign n8402 = n8388 & ~n8400 ;
  assign n8403 = n8401 | n8402 ;
  assign n8404 = n650 & n5658 ;
  assign n8405 = n7513 & n8128 ;
  assign n8406 = n8404 | n8405 ;
  assign n8407 = x44 & x46 ;
  assign n8408 = n720 & n8407 ;
  assign n8409 = x43 & n8408 ;
  assign n8410 = ( x43 & ~n8406 ) | ( x43 & n8409 ) | ( ~n8406 & n8409 ) ;
  assign n8411 = x14 & n8410 ;
  assign n8412 = n8406 | n8408 ;
  assign n8413 = x11 & x46 ;
  assign n8414 = ( n6653 & ~n8408 ) | ( n6653 & n8413 ) | ( ~n8408 & n8413 ) ;
  assign n8415 = n6653 & n8413 ;
  assign n8416 = ( ~n8406 & n8414 ) | ( ~n8406 & n8415 ) | ( n8414 & n8415 ) ;
  assign n8417 = ~n8412 & n8416 ;
  assign n8418 = n8411 | n8417 ;
  assign n8419 = n2369 | n3080 ;
  assign n8420 = n2372 & n2709 ;
  assign n8421 = x12 & x45 ;
  assign n8422 = ~n8420 & n8421 ;
  assign n8423 = n8419 | n8420 ;
  assign n8424 = ( n8420 & n8422 ) | ( n8420 & n8423 ) | ( n8422 & n8423 ) ;
  assign n8425 = n8419 & ~n8424 ;
  assign n8426 = ( ~n8419 & n8420 ) | ( ~n8419 & n8421 ) | ( n8420 & n8421 ) ;
  assign n8427 = n8421 & n8426 ;
  assign n8428 = n8425 | n8427 ;
  assign n8429 = n8418 & n8428 ;
  assign n8430 = n8418 & ~n8429 ;
  assign n8431 = n8428 & ~n8429 ;
  assign n8432 = n8430 | n8431 ;
  assign n8433 = x39 & x51 ;
  assign n8434 = n1415 & n8433 ;
  assign n8435 = n1020 & n4555 ;
  assign n8436 = n8434 | n8435 ;
  assign n8437 = x17 & x51 ;
  assign n8438 = n5314 & n8437 ;
  assign n8439 = x39 & n8438 ;
  assign n8440 = ( x39 & ~n8436 ) | ( x39 & n8439 ) | ( ~n8436 & n8439 ) ;
  assign n8441 = x18 & n8440 ;
  assign n8442 = n8436 | n8438 ;
  assign n8443 = x6 & x51 ;
  assign n8444 = x17 & x40 ;
  assign n8445 = ( ~n8438 & n8443 ) | ( ~n8438 & n8444 ) | ( n8443 & n8444 ) ;
  assign n8446 = n8443 & n8444 ;
  assign n8447 = ( ~n8436 & n8445 ) | ( ~n8436 & n8446 ) | ( n8445 & n8446 ) ;
  assign n8448 = ~n8442 & n8447 ;
  assign n8449 = n8441 | n8448 ;
  assign n8450 = ~n8432 & n8449 ;
  assign n8451 = n8432 & ~n8449 ;
  assign n8452 = n8450 | n8451 ;
  assign n8453 = n8403 | n8452 ;
  assign n8454 = n8403 & n8452 ;
  assign n8455 = n8453 & ~n8454 ;
  assign n8456 = n8001 | n8007 ;
  assign n8457 = ( n8001 & n8002 ) | ( n8001 & n8456 ) | ( n8002 & n8456 ) ;
  assign n8458 = n8455 & n8457 ;
  assign n8459 = n8455 | n8457 ;
  assign n8460 = ~n8458 & n8459 ;
  assign n8461 = n7951 | n8133 ;
  assign n8462 = n7951 & n8133 ;
  assign n8463 = n8461 & ~n8462 ;
  assign n8464 = n8059 | n8463 ;
  assign n8465 = n8059 & n8463 ;
  assign n8466 = n8464 & ~n8465 ;
  assign n8467 = n7956 & n8466 ;
  assign n8468 = ( n7962 & n8466 ) | ( n7962 & n8467 ) | ( n8466 & n8467 ) ;
  assign n8469 = n7956 | n8466 ;
  assign n8470 = n7962 | n8469 ;
  assign n8471 = ~n8468 & n8470 ;
  assign n8472 = n251 & n6834 ;
  assign n8473 = x16 & x50 ;
  assign n8474 = n5812 & n8473 ;
  assign n8475 = n8472 | n8474 ;
  assign n8476 = x16 & x49 ;
  assign n8477 = n6049 & n8476 ;
  assign n8478 = x50 & n8477 ;
  assign n8479 = ( x50 & ~n8475 ) | ( x50 & n8478 ) | ( ~n8475 & n8478 ) ;
  assign n8480 = x7 & n8479 ;
  assign n8481 = n8475 | n8477 ;
  assign n8482 = x8 & x49 ;
  assign n8483 = x16 & x41 ;
  assign n8484 = ( ~n8477 & n8482 ) | ( ~n8477 & n8483 ) | ( n8482 & n8483 ) ;
  assign n8485 = n8482 & n8483 ;
  assign n8486 = ( ~n8475 & n8484 ) | ( ~n8475 & n8485 ) | ( n8484 & n8485 ) ;
  assign n8487 = ~n8481 & n8486 ;
  assign n8488 = n8480 | n8487 ;
  assign n8489 = n1337 & n4914 ;
  assign n8490 = n1585 & n4078 ;
  assign n8491 = n8489 | n8490 ;
  assign n8492 = n1932 & n3483 ;
  assign n8493 = x36 & n8492 ;
  assign n8494 = ( x36 & ~n8491 ) | ( x36 & n8493 ) | ( ~n8491 & n8493 ) ;
  assign n8495 = x21 & n8494 ;
  assign n8496 = n8491 | n8492 ;
  assign n8497 = x22 & x35 ;
  assign n8498 = x23 & x34 ;
  assign n8499 = ( ~n8492 & n8497 ) | ( ~n8492 & n8498 ) | ( n8497 & n8498 ) ;
  assign n8500 = n8497 & n8498 ;
  assign n8501 = ( ~n8491 & n8499 ) | ( ~n8491 & n8500 ) | ( n8499 & n8500 ) ;
  assign n8502 = ~n8496 & n8501 ;
  assign n8503 = n8495 | n8502 ;
  assign n8504 = n8488 & n8503 ;
  assign n8505 = n8488 & ~n8504 ;
  assign n8506 = n8503 & ~n8504 ;
  assign n8507 = n8505 | n8506 ;
  assign n8508 = n2340 & n2683 ;
  assign n8509 = n1912 & n3321 ;
  assign n8510 = n8508 | n8509 ;
  assign n8511 = n2511 & n4062 ;
  assign n8512 = x33 & n8511 ;
  assign n8513 = ( x33 & ~n8510 ) | ( x33 & n8512 ) | ( ~n8510 & n8512 ) ;
  assign n8514 = x24 & n8513 ;
  assign n8515 = n8510 | n8511 ;
  assign n8516 = x25 & x32 ;
  assign n8517 = x26 & x31 ;
  assign n8518 = ( ~n8511 & n8516 ) | ( ~n8511 & n8517 ) | ( n8516 & n8517 ) ;
  assign n8519 = n8516 & n8517 ;
  assign n8520 = ( ~n8510 & n8518 ) | ( ~n8510 & n8519 ) | ( n8518 & n8519 ) ;
  assign n8521 = ~n8515 & n8520 ;
  assign n8522 = n8514 | n8521 ;
  assign n8523 = ~n8507 & n8522 ;
  assign n8524 = n8507 & ~n8522 ;
  assign n8525 = n8523 | n8524 ;
  assign n8526 = n8471 & n8525 ;
  assign n8527 = n8471 | n8525 ;
  assign n8528 = ~n8526 & n8527 ;
  assign n8529 = n7970 | n7976 ;
  assign n8530 = ( n7970 & n7974 ) | ( n7970 & n8529 ) | ( n7974 & n8529 ) ;
  assign n8531 = ( n8460 & ~n8528 ) | ( n8460 & n8530 ) | ( ~n8528 & n8530 ) ;
  assign n8532 = ( n8528 & ~n8530 ) | ( n8528 & n8531 ) | ( ~n8530 & n8531 ) ;
  assign n8533 = ( ~n8460 & n8531 ) | ( ~n8460 & n8532 ) | ( n8531 & n8532 ) ;
  assign n8534 = n8354 & ~n8533 ;
  assign n8535 = n8354 | n8533 ;
  assign n8536 = ( ~n8354 & n8534 ) | ( ~n8354 & n8535 ) | ( n8534 & n8535 ) ;
  assign n8537 = n8306 | n8536 ;
  assign n8538 = n8306 & ~n8536 ;
  assign n8539 = ( ~n8306 & n8537 ) | ( ~n8306 & n8538 ) | ( n8537 & n8538 ) ;
  assign n8540 = n7992 | n8231 ;
  assign n8541 = ( n7992 & n7995 ) | ( n7992 & n8540 ) | ( n7995 & n8540 ) ;
  assign n8542 = ( n8253 & n8539 ) | ( n8253 & ~n8541 ) | ( n8539 & ~n8541 ) ;
  assign n8543 = ( ~n8539 & n8541 ) | ( ~n8539 & n8542 ) | ( n8541 & n8542 ) ;
  assign n8544 = ( ~n8253 & n8542 ) | ( ~n8253 & n8543 ) | ( n8542 & n8543 ) ;
  assign n8545 = n8059 | n8462 ;
  assign n8546 = ( n8462 & n8463 ) | ( n8462 & n8545 ) | ( n8463 & n8545 ) ;
  assign n8547 = n8332 | n8335 ;
  assign n8548 = ( n8332 & n8333 ) | ( n8332 & n8547 ) | ( n8333 & n8547 ) ;
  assign n8549 = n8546 | n8548 ;
  assign n8550 = n8546 & n8548 ;
  assign n8551 = n8549 & ~n8550 ;
  assign n8552 = n8324 | n8326 ;
  assign n8553 = ( n8324 & n8325 ) | ( n8324 & n8552 ) | ( n8325 & n8552 ) ;
  assign n8554 = n8551 | n8553 ;
  assign n8555 = n8551 & n8553 ;
  assign n8556 = n8554 & ~n8555 ;
  assign n8557 = n8339 | n8344 ;
  assign n8558 = n8556 & n8557 ;
  assign n8559 = n8556 | n8557 ;
  assign n8560 = ~n8558 & n8559 ;
  assign n8561 = n8468 | n8525 ;
  assign n8562 = ( n8468 & n8471 ) | ( n8468 & n8561 ) | ( n8471 & n8561 ) ;
  assign n8563 = n8560 & n8562 ;
  assign n8564 = n8560 | n8562 ;
  assign n8565 = ~n8563 & n8564 ;
  assign n8566 = n8321 | n8346 ;
  assign n8567 = ( n8321 & n8322 ) | ( n8321 & n8566 ) | ( n8322 & n8566 ) ;
  assign n8568 = n8565 | n8567 ;
  assign n8569 = n8565 & n8567 ;
  assign n8570 = n8568 & ~n8569 ;
  assign n8571 = n8528 & n8530 ;
  assign n8572 = n8530 & ~n8571 ;
  assign n8573 = n8528 & ~n8530 ;
  assign n8574 = n8460 & ~n8573 ;
  assign n8575 = ~n8572 & n8574 ;
  assign n8576 = ( n8460 & n8571 ) | ( n8460 & ~n8575 ) | ( n8571 & ~n8575 ) ;
  assign n8577 = n8570 & n8576 ;
  assign n8578 = n8570 | n8576 ;
  assign n8579 = ~n8577 & n8578 ;
  assign n8580 = n8349 | n8531 ;
  assign n8581 = ~n8349 & n8460 ;
  assign n8582 = ( n8532 & n8580 ) | ( n8532 & ~n8581 ) | ( n8580 & ~n8581 ) ;
  assign n8583 = ( n8351 & n8533 ) | ( n8351 & n8582 ) | ( n8533 & n8582 ) ;
  assign n8584 = n8579 & n8583 ;
  assign n8585 = n8353 & n8579 ;
  assign n8586 = ( n8354 & n8584 ) | ( n8354 & n8585 ) | ( n8584 & n8585 ) ;
  assign n8587 = n8579 | n8583 ;
  assign n8588 = n8353 | n8579 ;
  assign n8589 = ( n8354 & n8587 ) | ( n8354 & n8588 ) | ( n8587 & n8588 ) ;
  assign n8590 = ~n8586 & n8589 ;
  assign n8591 = n8385 | n8400 ;
  assign n8592 = ( n8385 & n8388 ) | ( n8385 & n8591 ) | ( n8388 & n8591 ) ;
  assign n8593 = x1 & x57 ;
  assign n8594 = n3280 & n8593 ;
  assign n8595 = n3280 | n8593 ;
  assign n8596 = ~n8594 & n8595 ;
  assign n8597 = n8268 | n8596 ;
  assign n8598 = n8268 & n8596 ;
  assign n8599 = n8597 & ~n8598 ;
  assign n8600 = n8424 & n8599 ;
  assign n8601 = n8424 | n8599 ;
  assign n8602 = ~n8600 & n8601 ;
  assign n8603 = n8591 & n8602 ;
  assign n8604 = n8385 & n8602 ;
  assign n8605 = ( n8388 & n8603 ) | ( n8388 & n8604 ) | ( n8603 & n8604 ) ;
  assign n8606 = n8592 & ~n8605 ;
  assign n8607 = n8602 & ~n8605 ;
  assign n8608 = n8606 | n8607 ;
  assign n8609 = n8429 | n8449 ;
  assign n8610 = ( n8429 & n8432 ) | ( n8429 & n8609 ) | ( n8432 & n8609 ) ;
  assign n8611 = n8608 | n8610 ;
  assign n8612 = n8608 & ~n8610 ;
  assign n8613 = ( ~n8608 & n8611 ) | ( ~n8608 & n8612 ) | ( n8611 & n8612 ) ;
  assign n8614 = n8454 | n8457 ;
  assign n8615 = ( n8454 & n8455 ) | ( n8454 & n8614 ) | ( n8455 & n8614 ) ;
  assign n8616 = n8613 & n8615 ;
  assign n8617 = n8613 | n8615 ;
  assign n8618 = ~n8616 & n8617 ;
  assign n8619 = n8396 | n8515 ;
  assign n8620 = n8396 & n8515 ;
  assign n8621 = n8619 & ~n8620 ;
  assign n8622 = n8496 | n8621 ;
  assign n8623 = n8496 & n8621 ;
  assign n8624 = n8622 & ~n8623 ;
  assign n8625 = n8365 | n8380 ;
  assign n8626 = n8365 & n8380 ;
  assign n8627 = n8625 & ~n8626 ;
  assign n8628 = n8412 | n8627 ;
  assign n8629 = n8412 & n8627 ;
  assign n8630 = n8628 & ~n8629 ;
  assign n8631 = n8624 & n8630 ;
  assign n8632 = n8624 | n8630 ;
  assign n8633 = ~n8631 & n8632 ;
  assign n8634 = n8504 | n8522 ;
  assign n8635 = ( n8504 & n8507 ) | ( n8504 & n8634 ) | ( n8507 & n8634 ) ;
  assign n8636 = n8633 & n8635 ;
  assign n8637 = n8633 | n8635 ;
  assign n8638 = ~n8636 & n8637 ;
  assign n8639 = n8618 & n8638 ;
  assign n8640 = n8618 | n8638 ;
  assign n8641 = ~n8639 & n8640 ;
  assign n8642 = n8289 | n8641 ;
  assign n8643 = n8295 | n8642 ;
  assign n8644 = ( n8254 & n8289 ) | ( n8254 & n8641 ) | ( n8289 & n8641 ) ;
  assign n8645 = n8289 & n8641 ;
  assign n8646 = ( n8294 & n8644 ) | ( n8294 & n8645 ) | ( n8644 & n8645 ) ;
  assign n8647 = n8643 & ~n8646 ;
  assign n8648 = n2148 & n4914 ;
  assign n8649 = n1932 & n4078 ;
  assign n8650 = n8648 | n8649 ;
  assign n8651 = n1686 & n3483 ;
  assign n8652 = x36 & n8651 ;
  assign n8653 = ( x36 & ~n8650 ) | ( x36 & n8652 ) | ( ~n8650 & n8652 ) ;
  assign n8654 = x22 & n8653 ;
  assign n8655 = n8650 | n8651 ;
  assign n8656 = x23 & x35 ;
  assign n8657 = x24 & x34 ;
  assign n8658 = ( ~n8651 & n8656 ) | ( ~n8651 & n8657 ) | ( n8656 & n8657 ) ;
  assign n8659 = n8656 & n8657 ;
  assign n8660 = ( ~n8650 & n8658 ) | ( ~n8650 & n8659 ) | ( n8658 & n8659 ) ;
  assign n8661 = ~n8655 & n8660 ;
  assign n8662 = n8654 | n8661 ;
  assign n8663 = x7 & x51 ;
  assign n8664 = x8 & x50 ;
  assign n8665 = n8663 | n8664 ;
  assign n8666 = n251 & n7112 ;
  assign n8667 = n8665 | n8666 ;
  assign n8668 = x18 & x40 ;
  assign n8669 = ( ~n8666 & n8667 ) | ( ~n8666 & n8668 ) | ( n8667 & n8668 ) ;
  assign n8670 = ( n8666 & n8667 ) | ( n8666 & ~n8668 ) | ( n8667 & ~n8668 ) ;
  assign n8671 = ( ~n8667 & n8669 ) | ( ~n8667 & n8670 ) | ( n8669 & n8670 ) ;
  assign n8672 = n8662 & n8671 ;
  assign n8673 = n8662 & ~n8672 ;
  assign n8674 = n2683 & n2724 ;
  assign n8675 = n2511 & n3321 ;
  assign n8676 = n8674 | n8675 ;
  assign n8677 = n2267 & n4062 ;
  assign n8678 = n3466 & n8677 ;
  assign n8679 = ( n3466 & ~n8676 ) | ( n3466 & n8678 ) | ( ~n8676 & n8678 ) ;
  assign n8680 = n8676 | n8677 ;
  assign n8681 = x27 & x31 ;
  assign n8682 = ( n3422 & ~n8677 ) | ( n3422 & n8681 ) | ( ~n8677 & n8681 ) ;
  assign n8683 = n3422 & n8681 ;
  assign n8684 = ( ~n8676 & n8682 ) | ( ~n8676 & n8683 ) | ( n8682 & n8683 ) ;
  assign n8685 = ~n8680 & n8684 ;
  assign n8686 = n8679 | n8685 ;
  assign n8687 = ~n8662 & n8671 ;
  assign n8688 = n8686 & ~n8687 ;
  assign n8689 = ~n8673 & n8688 ;
  assign n8690 = ~n8686 & n8687 ;
  assign n8691 = ( n8673 & ~n8686 ) | ( n8673 & n8690 ) | ( ~n8686 & n8690 ) ;
  assign n8692 = n8689 | n8691 ;
  assign n8693 = x20 & x38 ;
  assign n8694 = x21 & x37 ;
  assign n8695 = n8693 | n8694 ;
  assign n8696 = n1434 & n4857 ;
  assign n8697 = x5 & x53 ;
  assign n8698 = ~n8696 & n8697 ;
  assign n8699 = n8695 | n8696 ;
  assign n8700 = ( n8696 & n8698 ) | ( n8696 & n8699 ) | ( n8698 & n8699 ) ;
  assign n8701 = n8695 & ~n8700 ;
  assign n8702 = ( ~n8695 & n8696 ) | ( ~n8695 & n8697 ) | ( n8696 & n8697 ) ;
  assign n8703 = n8697 & n8702 ;
  assign n8704 = n8701 | n8703 ;
  assign n8705 = x0 & x58 ;
  assign n8706 = x4 & x54 ;
  assign n8707 = n8705 & n8706 ;
  assign n8708 = x56 & x58 ;
  assign n8709 = n67 & n8708 ;
  assign n8710 = n119 & n8146 ;
  assign n8711 = n8709 | n8710 ;
  assign n8712 = x2 & x56 ;
  assign n8713 = n8707 & n8712 ;
  assign n8714 = ( ~n8711 & n8712 ) | ( ~n8711 & n8713 ) | ( n8712 & n8713 ) ;
  assign n8715 = ( n8705 & n8706 ) | ( n8705 & ~n8711 ) | ( n8706 & ~n8711 ) ;
  assign n8716 = ( ~n8707 & n8714 ) | ( ~n8707 & n8715 ) | ( n8714 & n8715 ) ;
  assign n8717 = n8704 & n8716 ;
  assign n8718 = n8704 & ~n8717 ;
  assign n8719 = n1023 & n5710 ;
  assign n8720 = n6414 & n7666 ;
  assign n8721 = n8719 | n8720 ;
  assign n8722 = x42 & x49 ;
  assign n8723 = n754 & n8722 ;
  assign n8724 = x41 & n8723 ;
  assign n8725 = ( x41 & ~n8721 ) | ( x41 & n8724 ) | ( ~n8721 & n8724 ) ;
  assign n8726 = x17 & n8725 ;
  assign n8727 = n8721 | n8723 ;
  assign n8728 = x9 & x49 ;
  assign n8729 = x16 & x42 ;
  assign n8730 = ( ~n8723 & n8728 ) | ( ~n8723 & n8729 ) | ( n8728 & n8729 ) ;
  assign n8731 = n8728 & n8729 ;
  assign n8732 = ( ~n8721 & n8730 ) | ( ~n8721 & n8731 ) | ( n8730 & n8731 ) ;
  assign n8733 = ~n8727 & n8732 ;
  assign n8734 = n8726 | n8733 ;
  assign n8735 = ~n8704 & n8716 ;
  assign n8736 = n8734 & n8735 ;
  assign n8737 = ( n8718 & n8734 ) | ( n8718 & n8736 ) | ( n8734 & n8736 ) ;
  assign n8738 = n8734 | n8735 ;
  assign n8739 = n8718 | n8738 ;
  assign n8740 = ~n8737 & n8739 ;
  assign n8741 = ~n8692 & n8740 ;
  assign n8742 = n8692 & ~n8740 ;
  assign n8743 = n8741 | n8742 ;
  assign n8744 = n8312 | n8317 ;
  assign n8745 = n8743 | n8744 ;
  assign n8746 = n8743 & n8744 ;
  assign n8747 = n8745 & ~n8746 ;
  assign n8748 = n8257 | n8284 ;
  assign n8749 = ( n8259 & n8284 ) | ( n8259 & n8748 ) | ( n8284 & n8748 ) ;
  assign n8750 = ( n8261 & n8262 ) | ( n8261 & n8749 ) | ( n8262 & n8749 ) ;
  assign n8751 = n8442 | n8481 ;
  assign n8752 = n8442 & n8481 ;
  assign n8753 = n8751 & ~n8752 ;
  assign n8754 = n8266 & n8270 ;
  assign n8755 = ( n8265 & n8270 ) | ( n8265 & n8754 ) | ( n8270 & n8754 ) ;
  assign n8756 = n8264 | n8755 ;
  assign n8757 = n8753 | n8756 ;
  assign n8758 = n8753 & n8756 ;
  assign n8759 = n8757 & ~n8758 ;
  assign n8760 = n8275 | n8281 ;
  assign n8761 = ( n8277 & n8281 ) | ( n8277 & n8760 ) | ( n8281 & n8760 ) ;
  assign n8762 = n8759 & n8761 ;
  assign n8763 = n8279 & n8759 ;
  assign n8764 = ( n8280 & n8762 ) | ( n8280 & n8763 ) | ( n8762 & n8763 ) ;
  assign n8765 = n8759 | n8761 ;
  assign n8766 = n8279 | n8759 ;
  assign n8767 = ( n8280 & n8765 ) | ( n8280 & n8766 ) | ( n8765 & n8766 ) ;
  assign n8768 = ~n8764 & n8767 ;
  assign n8769 = n618 & n6762 ;
  assign n8770 = n7213 & n8074 ;
  assign n8771 = n8769 | n8770 ;
  assign n8772 = x43 & x47 ;
  assign n8773 = n718 & n8772 ;
  assign n8774 = x48 & n8773 ;
  assign n8775 = ( x48 & ~n8771 ) | ( x48 & n8774 ) | ( ~n8771 & n8774 ) ;
  assign n8776 = x10 & n8775 ;
  assign n8777 = n8771 | n8773 ;
  assign n8778 = x11 & x47 ;
  assign n8779 = ( n6070 & ~n8773 ) | ( n6070 & n8778 ) | ( ~n8773 & n8778 ) ;
  assign n8780 = n6070 & n8778 ;
  assign n8781 = ( ~n8771 & n8779 ) | ( ~n8771 & n8780 ) | ( n8779 & n8780 ) ;
  assign n8782 = ~n8777 & n8781 ;
  assign n8783 = n8776 | n8782 ;
  assign n8784 = n487 & n8407 ;
  assign n8785 = n650 & n6093 ;
  assign n8786 = n8784 | n8785 ;
  assign n8787 = n647 & n5975 ;
  assign n8788 = n7170 & n8787 ;
  assign n8789 = ( n7170 & ~n8786 ) | ( n7170 & n8788 ) | ( ~n8786 & n8788 ) ;
  assign n8790 = n8786 | n8787 ;
  assign n8791 = x12 & x46 ;
  assign n8792 = ( n7823 & ~n8787 ) | ( n7823 & n8791 ) | ( ~n8787 & n8791 ) ;
  assign n8793 = n7823 & n8791 ;
  assign n8794 = ( ~n8786 & n8792 ) | ( ~n8786 & n8793 ) | ( n8792 & n8793 ) ;
  assign n8795 = ~n8790 & n8794 ;
  assign n8796 = n8789 | n8795 ;
  assign n8797 = n8783 & n8796 ;
  assign n8798 = n8783 & ~n8797 ;
  assign n8799 = x6 & x52 ;
  assign n8800 = x19 & x39 ;
  assign n8801 = n8799 | n8800 ;
  assign n8802 = x3 & x55 ;
  assign n8803 = ( n8799 & n8800 ) | ( n8799 & n8802 ) | ( n8800 & n8802 ) ;
  assign n8804 = n8801 & ~n8803 ;
  assign n8805 = n8799 & n8800 ;
  assign n8806 = n8802 & ~n8805 ;
  assign n8807 = ~n8801 & n8802 ;
  assign n8808 = ( n8802 & ~n8806 ) | ( n8802 & n8807 ) | ( ~n8806 & n8807 ) ;
  assign n8809 = n8804 | n8808 ;
  assign n8810 = ~n8783 & n8796 ;
  assign n8811 = n8809 & n8810 ;
  assign n8812 = ( n8798 & n8809 ) | ( n8798 & n8811 ) | ( n8809 & n8811 ) ;
  assign n8813 = n8809 | n8810 ;
  assign n8814 = n8798 | n8813 ;
  assign n8815 = ~n8812 & n8814 ;
  assign n8816 = n8768 | n8815 ;
  assign n8817 = n8768 & n8815 ;
  assign n8818 = n8816 & ~n8817 ;
  assign n8819 = n8749 & n8818 ;
  assign n8820 = n8261 & n8818 ;
  assign n8821 = ( n8262 & n8819 ) | ( n8262 & n8820 ) | ( n8819 & n8820 ) ;
  assign n8822 = n8750 & ~n8821 ;
  assign n8823 = ~n8749 & n8818 ;
  assign n8824 = ~n8261 & n8818 ;
  assign n8825 = ( ~n8262 & n8823 ) | ( ~n8262 & n8824 ) | ( n8823 & n8824 ) ;
  assign n8826 = n8747 & n8825 ;
  assign n8827 = ( n8747 & n8822 ) | ( n8747 & n8826 ) | ( n8822 & n8826 ) ;
  assign n8828 = n8747 | n8825 ;
  assign n8829 = n8822 | n8828 ;
  assign n8830 = ~n8827 & n8829 ;
  assign n8831 = ~n8646 & n8830 ;
  assign n8832 = n8643 & n8831 ;
  assign n8833 = n8647 & ~n8832 ;
  assign n8834 = n8646 & n8830 ;
  assign n8835 = ( ~n8643 & n8830 ) | ( ~n8643 & n8834 ) | ( n8830 & n8834 ) ;
  assign n8836 = n8590 & n8835 ;
  assign n8837 = ( n8590 & n8833 ) | ( n8590 & n8836 ) | ( n8833 & n8836 ) ;
  assign n8838 = n8590 | n8835 ;
  assign n8839 = n8833 | n8838 ;
  assign n8840 = ~n8837 & n8839 ;
  assign n8841 = ( n8297 & n8302 ) | ( n8297 & n8536 ) | ( n8302 & n8536 ) ;
  assign n8842 = n8840 & n8841 ;
  assign n8843 = n8840 | n8841 ;
  assign n8844 = ~n8842 & n8843 ;
  assign n8845 = n8539 & n8541 ;
  assign n8846 = n8539 | n8541 ;
  assign n8847 = n8248 & n8846 ;
  assign n8848 = n8845 | n8847 ;
  assign n8849 = n8845 | n8846 ;
  assign n8850 = ( n8252 & n8848 ) | ( n8252 & n8849 ) | ( n8848 & n8849 ) ;
  assign n8851 = n8844 | n8850 ;
  assign n8852 = n8843 & n8849 ;
  assign n8853 = n8843 & n8845 ;
  assign n8854 = ( n8843 & n8847 ) | ( n8843 & n8853 ) | ( n8847 & n8853 ) ;
  assign n8855 = ( n8252 & n8852 ) | ( n8252 & n8854 ) | ( n8852 & n8854 ) ;
  assign n8856 = ~n8842 & n8855 ;
  assign n8857 = n8851 & ~n8856 ;
  assign n8858 = n8842 | n8854 ;
  assign n8859 = n8842 | n8843 ;
  assign n8860 = ( n8842 & n8849 ) | ( n8842 & n8859 ) | ( n8849 & n8859 ) ;
  assign n8861 = ( n8252 & n8858 ) | ( n8252 & n8860 ) | ( n8858 & n8860 ) ;
  assign n8862 = n8821 | n8827 ;
  assign n8863 = n8752 | n8758 ;
  assign n8864 = n8412 | n8626 ;
  assign n8865 = ( n8626 & n8627 ) | ( n8626 & n8864 ) | ( n8627 & n8864 ) ;
  assign n8866 = n8863 | n8865 ;
  assign n8867 = n8863 & n8865 ;
  assign n8868 = n8866 & ~n8867 ;
  assign n8869 = n8496 | n8620 ;
  assign n8870 = ( n8620 & n8621 ) | ( n8620 & n8869 ) | ( n8621 & n8869 ) ;
  assign n8871 = n8868 | n8870 ;
  assign n8872 = n8868 & n8870 ;
  assign n8873 = n8871 & ~n8872 ;
  assign n8874 = n8631 | n8636 ;
  assign n8875 = n8873 & n8874 ;
  assign n8876 = n8873 | n8874 ;
  assign n8877 = ~n8875 & n8876 ;
  assign n8878 = n8764 | n8815 ;
  assign n8879 = ( n8764 & n8768 ) | ( n8764 & n8878 ) | ( n8768 & n8878 ) ;
  assign n8880 = n8877 & n8879 ;
  assign n8881 = n8877 | n8879 ;
  assign n8882 = ~n8880 & n8881 ;
  assign n8883 = n8613 | n8638 ;
  assign n8884 = ( n8615 & n8638 ) | ( n8615 & n8883 ) | ( n8638 & n8883 ) ;
  assign n8885 = n8882 & n8884 ;
  assign n8886 = n8616 & n8882 ;
  assign n8887 = ( n8618 & n8885 ) | ( n8618 & n8886 ) | ( n8885 & n8886 ) ;
  assign n8888 = n8882 | n8884 ;
  assign n8889 = n8616 | n8882 ;
  assign n8890 = ( n8618 & n8888 ) | ( n8618 & n8889 ) | ( n8888 & n8889 ) ;
  assign n8891 = ~n8887 & n8890 ;
  assign n8892 = n8862 & n8891 ;
  assign n8893 = n8862 | n8891 ;
  assign n8894 = ~n8892 & n8893 ;
  assign n8895 = n8646 | n8894 ;
  assign n8896 = n8832 | n8895 ;
  assign n8897 = n8646 & n8894 ;
  assign n8898 = ( n8832 & n8894 ) | ( n8832 & n8897 ) | ( n8894 & n8897 ) ;
  assign n8899 = n8896 & ~n8898 ;
  assign n8900 = x2 & x57 ;
  assign n8901 = x3 & x56 ;
  assign n8902 = n8900 | n8901 ;
  assign n8903 = x56 & x57 ;
  assign n8904 = n77 & n8903 ;
  assign n8905 = n8902 & ~n8904 ;
  assign n8906 = ( ~n8594 & n8680 ) | ( ~n8594 & n8905 ) | ( n8680 & n8905 ) ;
  assign n8907 = ( n8594 & n8680 ) | ( n8594 & ~n8905 ) | ( n8680 & ~n8905 ) ;
  assign n8908 = ( ~n8680 & n8906 ) | ( ~n8680 & n8907 ) | ( n8906 & n8907 ) ;
  assign n8909 = x5 & x54 ;
  assign n8910 = x19 & x40 ;
  assign n8911 = n8909 & n8910 ;
  assign n8912 = n91 & n8357 ;
  assign n8913 = x19 & x55 ;
  assign n8914 = n4902 & n8913 ;
  assign n8915 = n8912 | n8914 ;
  assign n8916 = x55 & n8911 ;
  assign n8917 = ( x55 & ~n8915 ) | ( x55 & n8916 ) | ( ~n8915 & n8916 ) ;
  assign n8918 = x4 & n8917 ;
  assign n8919 = ( n8909 & n8910 ) | ( n8909 & ~n8915 ) | ( n8910 & ~n8915 ) ;
  assign n8920 = ( ~n8911 & n8918 ) | ( ~n8911 & n8919 ) | ( n8918 & n8919 ) ;
  assign n8921 = n8908 & n8920 ;
  assign n8922 = n8908 | n8920 ;
  assign n8923 = ~n8921 & n8922 ;
  assign n8924 = n490 & n6762 ;
  assign n8925 = x45 & x48 ;
  assign n8926 = n1618 & n8925 ;
  assign n8927 = n8924 | n8926 ;
  assign n8928 = n487 & n5610 ;
  assign n8929 = x48 & n8928 ;
  assign n8930 = ( x48 & ~n8927 ) | ( x48 & n8929 ) | ( ~n8927 & n8929 ) ;
  assign n8931 = x11 & n8930 ;
  assign n8932 = n8927 | n8928 ;
  assign n8933 = x12 & x47 ;
  assign n8934 = x14 & x45 ;
  assign n8935 = ( ~n8928 & n8933 ) | ( ~n8928 & n8934 ) | ( n8933 & n8934 ) ;
  assign n8936 = n8933 & n8934 ;
  assign n8937 = ( ~n8927 & n8935 ) | ( ~n8927 & n8936 ) | ( n8935 & n8936 ) ;
  assign n8938 = ~n8932 & n8937 ;
  assign n8939 = n8931 | n8938 ;
  assign n8940 = x28 & x31 ;
  assign n8941 = n2709 | n8940 ;
  assign n8942 = x13 & x46 ;
  assign n8943 = ( n2709 & n8940 ) | ( n2709 & n8942 ) | ( n8940 & n8942 ) ;
  assign n8944 = n8941 & ~n8943 ;
  assign n8945 = n2709 & n8940 ;
  assign n8946 = n8942 & ~n8945 ;
  assign n8947 = ~n8941 & n8942 ;
  assign n8948 = ( n8942 & ~n8946 ) | ( n8942 & n8947 ) | ( ~n8946 & n8947 ) ;
  assign n8949 = n8944 | n8948 ;
  assign n8950 = n8939 & n8949 ;
  assign n8951 = n8939 & ~n8950 ;
  assign n8952 = x16 & x43 ;
  assign n8953 = x17 & x42 ;
  assign n8954 = n8952 | n8953 ;
  assign n8955 = n1023 & n5407 ;
  assign n8956 = x8 & x51 ;
  assign n8957 = ~n8955 & n8956 ;
  assign n8958 = n8954 | n8955 ;
  assign n8959 = ( n8955 & n8957 ) | ( n8955 & n8958 ) | ( n8957 & n8958 ) ;
  assign n8960 = n8954 & ~n8959 ;
  assign n8961 = ( ~n8954 & n8955 ) | ( ~n8954 & n8956 ) | ( n8955 & n8956 ) ;
  assign n8962 = n8956 & n8961 ;
  assign n8963 = n8960 | n8962 ;
  assign n8964 = ~n8939 & n8949 ;
  assign n8965 = n8963 & ~n8964 ;
  assign n8966 = ~n8951 & n8965 ;
  assign n8967 = n8923 & n8966 ;
  assign n8968 = ~n8963 & n8964 ;
  assign n8969 = ( n8951 & ~n8963 ) | ( n8951 & n8968 ) | ( ~n8963 & n8968 ) ;
  assign n8970 = ( n8923 & n8967 ) | ( n8923 & n8969 ) | ( n8967 & n8969 ) ;
  assign n8971 = n8923 | n8966 ;
  assign n8972 = n8969 | n8971 ;
  assign n8973 = ~n8970 & n8972 ;
  assign n8974 = n8605 | n8610 ;
  assign n8975 = ( n8605 & n8608 ) | ( n8605 & n8974 ) | ( n8608 & n8974 ) ;
  assign n8976 = n8973 & n8975 ;
  assign n8977 = n8973 | n8975 ;
  assign n8978 = ~n8976 & n8977 ;
  assign n8979 = n8558 | n8562 ;
  assign n8980 = ( n8558 & n8560 ) | ( n8558 & n8979 ) | ( n8560 & n8979 ) ;
  assign n8981 = n8978 | n8980 ;
  assign n8982 = n8978 & n8980 ;
  assign n8983 = n8981 & ~n8982 ;
  assign n8984 = x41 & x53 ;
  assign n8985 = n1415 & n8984 ;
  assign n8986 = n200 & n8161 ;
  assign n8987 = n8985 | n8986 ;
  assign n8988 = x18 & x52 ;
  assign n8989 = n5812 & n8988 ;
  assign n8990 = x53 & n8989 ;
  assign n8991 = ( x53 & ~n8987 ) | ( x53 & n8990 ) | ( ~n8987 & n8990 ) ;
  assign n8992 = x6 & n8991 ;
  assign n8993 = n8987 | n8989 ;
  assign n8994 = x7 & x52 ;
  assign n8995 = x18 & x41 ;
  assign n8996 = ( ~n8989 & n8994 ) | ( ~n8989 & n8995 ) | ( n8994 & n8995 ) ;
  assign n8997 = n8994 & n8995 ;
  assign n8998 = ( ~n8987 & n8996 ) | ( ~n8987 & n8997 ) | ( n8996 & n8997 ) ;
  assign n8999 = ~n8993 & n8998 ;
  assign n9000 = n8992 | n8999 ;
  assign n9001 = x44 & x50 ;
  assign n9002 = n1462 & n9001 ;
  assign n9003 = n360 & n6834 ;
  assign n9004 = n9002 | n9003 ;
  assign n9005 = x44 & x49 ;
  assign n9006 = n582 & n9005 ;
  assign n9007 = x50 & n9006 ;
  assign n9008 = ( x50 & ~n9004 ) | ( x50 & n9007 ) | ( ~n9004 & n9007 ) ;
  assign n9009 = x9 & n9008 ;
  assign n9010 = n9004 | n9006 ;
  assign n9011 = x10 & x49 ;
  assign n9012 = ( n5660 & ~n9006 ) | ( n5660 & n9011 ) | ( ~n9006 & n9011 ) ;
  assign n9013 = n5660 & n9011 ;
  assign n9014 = ( ~n9004 & n9012 ) | ( ~n9004 & n9013 ) | ( n9012 & n9013 ) ;
  assign n9015 = ~n9010 & n9014 ;
  assign n9016 = n9009 | n9015 ;
  assign n9017 = n9000 & n9016 ;
  assign n9018 = n9000 & ~n9017 ;
  assign n9019 = n9016 & ~n9017 ;
  assign n9020 = n9018 | n9019 ;
  assign n9021 = n8424 | n8598 ;
  assign n9022 = ( n8598 & n8599 ) | ( n8598 & n9021 ) | ( n8599 & n9021 ) ;
  assign n9023 = n9020 | n9022 ;
  assign n9024 = n9020 & n9022 ;
  assign n9025 = n9023 & ~n9024 ;
  assign n9026 = n8550 | n8553 ;
  assign n9027 = ( n8550 & n8551 ) | ( n8550 & n9026 ) | ( n8551 & n9026 ) ;
  assign n9028 = n9025 | n9027 ;
  assign n9029 = n9025 & n9027 ;
  assign n9030 = n9028 & ~n9029 ;
  assign n9031 = n1710 & n5798 ;
  assign n9032 = n1434 & n5392 ;
  assign n9033 = n9031 | n9032 ;
  assign n9034 = n1585 & n4857 ;
  assign n9035 = x39 & n9034 ;
  assign n9036 = ( x39 & ~n9033 ) | ( x39 & n9035 ) | ( ~n9033 & n9035 ) ;
  assign n9037 = x20 & n9036 ;
  assign n9038 = n9033 | n9034 ;
  assign n9039 = x21 & x38 ;
  assign n9040 = x22 & x37 ;
  assign n9041 = ( ~n9034 & n9039 ) | ( ~n9034 & n9040 ) | ( n9039 & n9040 ) ;
  assign n9042 = n9039 & n9040 ;
  assign n9043 = ( ~n9033 & n9041 ) | ( ~n9033 & n9042 ) | ( n9041 & n9042 ) ;
  assign n9044 = ~n9038 & n9043 ;
  assign n9045 = n9037 | n9044 ;
  assign n9046 = n1557 & n4914 ;
  assign n9047 = n1686 & n4078 ;
  assign n9048 = n9046 | n9047 ;
  assign n9049 = n1912 & n3483 ;
  assign n9050 = x36 & n9049 ;
  assign n9051 = ( x36 & ~n9048 ) | ( x36 & n9050 ) | ( ~n9048 & n9050 ) ;
  assign n9052 = x23 & n9051 ;
  assign n9053 = n9048 | n9049 ;
  assign n9054 = x24 & x35 ;
  assign n9055 = x25 & x34 ;
  assign n9056 = ( ~n9049 & n9054 ) | ( ~n9049 & n9055 ) | ( n9054 & n9055 ) ;
  assign n9057 = n9054 & n9055 ;
  assign n9058 = ( ~n9048 & n9056 ) | ( ~n9048 & n9057 ) | ( n9056 & n9057 ) ;
  assign n9059 = ~n9053 & n9058 ;
  assign n9060 = n9052 | n9059 ;
  assign n9061 = n9045 & n9060 ;
  assign n9062 = n9045 & ~n9061 ;
  assign n9063 = n9060 & ~n9061 ;
  assign n9064 = n9062 | n9063 ;
  assign n9065 = n2267 & n3321 ;
  assign n9066 = x26 & x59 ;
  assign n9067 = n2692 & n9066 ;
  assign n9068 = n9065 | n9067 ;
  assign n9069 = x32 & x59 ;
  assign n9070 = n1811 & n9069 ;
  assign n9071 = x33 & n9070 ;
  assign n9072 = ( x33 & ~n9068 ) | ( x33 & n9071 ) | ( ~n9068 & n9071 ) ;
  assign n9073 = x26 & n9072 ;
  assign n9074 = n9068 | n9070 ;
  assign n9075 = x0 & x59 ;
  assign n9076 = x27 & x32 ;
  assign n9077 = ( ~n9070 & n9075 ) | ( ~n9070 & n9076 ) | ( n9075 & n9076 ) ;
  assign n9078 = n9075 & n9076 ;
  assign n9079 = ( ~n9068 & n9077 ) | ( ~n9068 & n9078 ) | ( n9077 & n9078 ) ;
  assign n9080 = ~n9074 & n9079 ;
  assign n9081 = n9073 | n9080 ;
  assign n9082 = ~n9064 & n9081 ;
  assign n9083 = n9064 & ~n9081 ;
  assign n9084 = n9082 | n9083 ;
  assign n9085 = n9030 & n9084 ;
  assign n9086 = n9030 | n9084 ;
  assign n9087 = ~n9085 & n9086 ;
  assign n9088 = ~n8983 & n9087 ;
  assign n9089 = n8983 & ~n9087 ;
  assign n9090 = n9088 | n9089 ;
  assign n9120 = ( n8312 & n8692 ) | ( n8312 & n8740 ) | ( n8692 & n8740 ) ;
  assign n9121 = n8692 | n8740 ;
  assign n9122 = ( n8317 & n9120 ) | ( n8317 & n9121 ) | ( n9120 & n9121 ) ;
  assign n9091 = x58 & n2445 ;
  assign n9092 = x1 & x58 ;
  assign n9093 = x30 | n9092 ;
  assign n9094 = ~n9091 & n9093 ;
  assign n9095 = n8790 | n9094 ;
  assign n9096 = n8790 & n9094 ;
  assign n9097 = n9095 & ~n9096 ;
  assign n9098 = n8777 & n9097 ;
  assign n9099 = n8777 | n9097 ;
  assign n9100 = ~n9098 & n9099 ;
  assign n9101 = n8707 | n8803 ;
  assign n9102 = n8711 | n9101 ;
  assign n9103 = n8707 & n8803 ;
  assign n9104 = ( n8711 & n8803 ) | ( n8711 & n9103 ) | ( n8803 & n9103 ) ;
  assign n9105 = n9102 & ~n9104 ;
  assign n9106 = n8727 | n9105 ;
  assign n9107 = n8727 & n9105 ;
  assign n9108 = n9106 & ~n9107 ;
  assign n9109 = ~n8666 & n8668 ;
  assign n9110 = ( n8666 & n8667 ) | ( n8666 & n9109 ) | ( n8667 & n9109 ) ;
  assign n9111 = n8655 | n8700 ;
  assign n9112 = n8655 & n8700 ;
  assign n9113 = n9111 & ~n9112 ;
  assign n9114 = n9110 | n9113 ;
  assign n9115 = n9110 & n9113 ;
  assign n9116 = n9114 & ~n9115 ;
  assign n9117 = ( n9100 & n9108 ) | ( n9100 & ~n9116 ) | ( n9108 & ~n9116 ) ;
  assign n9118 = ( ~n9108 & n9116 ) | ( ~n9108 & n9117 ) | ( n9116 & n9117 ) ;
  assign n9119 = ( ~n9100 & n9117 ) | ( ~n9100 & n9118 ) | ( n9117 & n9118 ) ;
  assign n9123 = n9119 & n9122 ;
  assign n9124 = n9122 & ~n9123 ;
  assign n9125 = n8797 | n8812 ;
  assign n9126 = n8686 & n8687 ;
  assign n9127 = ( n8673 & n8686 ) | ( n8673 & n9126 ) | ( n8686 & n9126 ) ;
  assign n9128 = n8672 | n9127 ;
  assign n9129 = n9125 | n9128 ;
  assign n9130 = n9125 & n9128 ;
  assign n9131 = n9129 & ~n9130 ;
  assign n9132 = n8717 | n8737 ;
  assign n9133 = n9131 | n9132 ;
  assign n9134 = n9131 & n9132 ;
  assign n9135 = n9133 & ~n9134 ;
  assign n9136 = n9119 & ~n9122 ;
  assign n9137 = n9135 & n9136 ;
  assign n9138 = ( n9124 & n9135 ) | ( n9124 & n9137 ) | ( n9135 & n9137 ) ;
  assign n9139 = ( n9119 & n9122 ) | ( n9119 & ~n9123 ) | ( n9122 & ~n9123 ) ;
  assign n9140 = ( ~n9123 & n9135 ) | ( ~n9123 & n9139 ) | ( n9135 & n9139 ) ;
  assign n9141 = ~n9138 & n9140 ;
  assign n9142 = n8569 & n9141 ;
  assign n9143 = ( n8570 & n9141 ) | ( n8570 & n9142 ) | ( n9141 & n9142 ) ;
  assign n9144 = n9141 & n9142 ;
  assign n9145 = ( n8576 & n9143 ) | ( n8576 & n9144 ) | ( n9143 & n9144 ) ;
  assign n9146 = n8569 | n9141 ;
  assign n9147 = n8570 | n9146 ;
  assign n9148 = ( n8576 & n9146 ) | ( n8576 & n9147 ) | ( n9146 & n9147 ) ;
  assign n9149 = ~n9145 & n9148 ;
  assign n9150 = n9090 & n9149 ;
  assign n9151 = n9090 | n9149 ;
  assign n9152 = ~n9150 & n9151 ;
  assign n9153 = n8899 & n9152 ;
  assign n9154 = n8899 | n9152 ;
  assign n9155 = ~n9153 & n9154 ;
  assign n9156 = n8586 | n8833 ;
  assign n9157 = n8586 | n8590 ;
  assign n9158 = ( n8836 & n9156 ) | ( n8836 & n9157 ) | ( n9156 & n9157 ) ;
  assign n9159 = ( n8861 & n9155 ) | ( n8861 & ~n9158 ) | ( n9155 & ~n9158 ) ;
  assign n9160 = ( ~n9155 & n9158 ) | ( ~n9155 & n9159 ) | ( n9158 & n9159 ) ;
  assign n9161 = ( ~n8861 & n9159 ) | ( ~n8861 & n9160 ) | ( n9159 & n9160 ) ;
  assign n9162 = n9155 & n9158 ;
  assign n9163 = n9155 | n9158 ;
  assign n9164 = n8859 & n9163 ;
  assign n9165 = n8842 & n9163 ;
  assign n9166 = ( n8849 & n9164 ) | ( n8849 & n9165 ) | ( n9164 & n9165 ) ;
  assign n9167 = ( n8854 & n9163 ) | ( n8854 & n9165 ) | ( n9163 & n9165 ) ;
  assign n9168 = ( n8252 & n9166 ) | ( n8252 & n9167 ) | ( n9166 & n9167 ) ;
  assign n9169 = n9162 | n9168 ;
  assign n9170 = n9110 | n9112 ;
  assign n9171 = ( n9112 & n9113 ) | ( n9112 & n9170 ) | ( n9113 & n9170 ) ;
  assign n9172 = n8727 | n9104 ;
  assign n9173 = ( n9104 & n9105 ) | ( n9104 & n9172 ) | ( n9105 & n9172 ) ;
  assign n9174 = n9171 | n9173 ;
  assign n9175 = n9171 & n9173 ;
  assign n9176 = n9174 & ~n9175 ;
  assign n9177 = n8594 | n8904 ;
  assign n9178 = ( n8904 & n8905 ) | ( n8904 & n9177 ) | ( n8905 & n9177 ) ;
  assign n9179 = n8902 & ~n9178 ;
  assign n9180 = n8594 & ~n8905 ;
  assign n9181 = n8680 & n9180 ;
  assign n9182 = ( n8680 & n9179 ) | ( n8680 & n9181 ) | ( n9179 & n9181 ) ;
  assign n9183 = n8921 | n9182 ;
  assign n9184 = n9176 | n9183 ;
  assign n9185 = n9176 & n9183 ;
  assign n9186 = n9184 & ~n9185 ;
  assign n9187 = n9130 | n9132 ;
  assign n9188 = ( n9130 & n9131 ) | ( n9130 & n9187 ) | ( n9131 & n9187 ) ;
  assign n9189 = n9186 | n9188 ;
  assign n9190 = n9186 & n9188 ;
  assign n9191 = n9189 & ~n9190 ;
  assign n9192 = n9029 | n9084 ;
  assign n9193 = ( n9029 & n9030 ) | ( n9029 & n9192 ) | ( n9030 & n9192 ) ;
  assign n9194 = n9191 & n9193 ;
  assign n9195 = n9191 | n9193 ;
  assign n9196 = ~n9194 & n9195 ;
  assign n9197 = n9123 & n9196 ;
  assign n9198 = ( n9138 & n9196 ) | ( n9138 & n9197 ) | ( n9196 & n9197 ) ;
  assign n9199 = ( n8978 & n8980 ) | ( n8978 & n9087 ) | ( n8980 & n9087 ) ;
  assign n9200 = n9123 | n9135 ;
  assign n9201 = n9123 | n9124 ;
  assign n9202 = ( n9137 & n9200 ) | ( n9137 & n9201 ) | ( n9200 & n9201 ) ;
  assign n9203 = n9199 & n9202 ;
  assign n9204 = ( n9196 & n9199 ) | ( n9196 & n9203 ) | ( n9199 & n9203 ) ;
  assign n9205 = ~n9198 & n9204 ;
  assign n9206 = n9199 | n9202 ;
  assign n9207 = n9196 | n9206 ;
  assign n9208 = ( ~n9198 & n9199 ) | ( ~n9198 & n9207 ) | ( n9199 & n9207 ) ;
  assign n9209 = ~n9205 & n9208 ;
  assign n9210 = n9090 | n9145 ;
  assign n9211 = ( n9145 & n9149 ) | ( n9145 & n9210 ) | ( n9149 & n9210 ) ;
  assign n9212 = n9209 | n9211 ;
  assign n9213 = n9209 & n9211 ;
  assign n9214 = n9212 & ~n9213 ;
  assign n9215 = n8959 | n8993 ;
  assign n9216 = n8959 & n8993 ;
  assign n9217 = n9215 & ~n9216 ;
  assign n9218 = n8943 | n9217 ;
  assign n9219 = n8943 & n9217 ;
  assign n9220 = n9218 & ~n9219 ;
  assign n9221 = n9061 | n9081 ;
  assign n9222 = n9220 & n9221 ;
  assign n9223 = n9061 & n9220 ;
  assign n9224 = ( n9064 & n9222 ) | ( n9064 & n9223 ) | ( n9222 & n9223 ) ;
  assign n9225 = n9220 | n9221 ;
  assign n9226 = n9061 | n9220 ;
  assign n9227 = ( n9064 & n9225 ) | ( n9064 & n9226 ) | ( n9225 & n9226 ) ;
  assign n9228 = ~n9224 & n9227 ;
  assign n9229 = n8963 & n8964 ;
  assign n9230 = ( n8951 & n8963 ) | ( n8951 & n9229 ) | ( n8963 & n9229 ) ;
  assign n9231 = n8950 | n9230 ;
  assign n9232 = n9228 | n9231 ;
  assign n9233 = n9228 & n9231 ;
  assign n9234 = n9232 & ~n9233 ;
  assign n9235 = n8911 | n8915 ;
  assign n9236 = n9038 | n9235 ;
  assign n9237 = n9038 & n9235 ;
  assign n9238 = n9236 & ~n9237 ;
  assign n9239 = n9053 | n9238 ;
  assign n9240 = n9053 & n9238 ;
  assign n9241 = n9239 & ~n9240 ;
  assign n9242 = n9074 | n9178 ;
  assign n9243 = n9074 & n9178 ;
  assign n9244 = n9242 & ~n9243 ;
  assign n9245 = n9010 | n9244 ;
  assign n9246 = n9010 & n9244 ;
  assign n9247 = n9245 & ~n9246 ;
  assign n9248 = n9241 & n9247 ;
  assign n9249 = n9241 | n9247 ;
  assign n9250 = ~n9248 & n9249 ;
  assign n9251 = n9017 | n9022 ;
  assign n9252 = ( n9017 & n9020 ) | ( n9017 & n9251 ) | ( n9020 & n9251 ) ;
  assign n9253 = n9250 & n9252 ;
  assign n9254 = n9250 | n9252 ;
  assign n9255 = ~n9253 & n9254 ;
  assign n9256 = n8970 & n9255 ;
  assign n9257 = n9255 & ~n9256 ;
  assign n9258 = ~n8976 & n9257 ;
  assign n9259 = n9234 | n9258 ;
  assign n9260 = ( n8976 & n9255 ) | ( n8976 & n9256 ) | ( n9255 & n9256 ) ;
  assign n9261 = ( n8970 & n8976 ) | ( n8970 & ~n9260 ) | ( n8976 & ~n9260 ) ;
  assign n9262 = n9259 | n9261 ;
  assign n9263 = n9234 & n9258 ;
  assign n9264 = ( n9234 & n9261 ) | ( n9234 & n9263 ) | ( n9261 & n9263 ) ;
  assign n9265 = n9262 & ~n9264 ;
  assign n9266 = n8887 & n9265 ;
  assign n9267 = ( n8891 & n9265 ) | ( n8891 & n9266 ) | ( n9265 & n9266 ) ;
  assign n9268 = n9265 & n9266 ;
  assign n9269 = ( n8862 & n9267 ) | ( n8862 & n9268 ) | ( n9267 & n9268 ) ;
  assign n9270 = ( n8887 & n8892 ) | ( n8887 & ~n9269 ) | ( n8892 & ~n9269 ) ;
  assign n9371 = n8875 | n8879 ;
  assign n9372 = ( n8875 & n8877 ) | ( n8875 & n9371 ) | ( n8877 & n9371 ) ;
  assign n9271 = n119 & n8708 ;
  assign n9272 = x57 & x58 ;
  assign n9273 = n77 & n9272 ;
  assign n9274 = n9271 | n9273 ;
  assign n9275 = n79 & n8903 ;
  assign n9276 = x58 & n9275 ;
  assign n9277 = ( x58 & ~n9274 ) | ( x58 & n9276 ) | ( ~n9274 & n9276 ) ;
  assign n9278 = x2 & n9277 ;
  assign n9279 = n9274 | n9275 ;
  assign n9280 = x3 & x57 ;
  assign n9281 = x4 & x56 ;
  assign n9282 = ( ~n9275 & n9280 ) | ( ~n9275 & n9281 ) | ( n9280 & n9281 ) ;
  assign n9283 = n9280 & n9281 ;
  assign n9284 = ( ~n9274 & n9282 ) | ( ~n9274 & n9283 ) | ( n9282 & n9283 ) ;
  assign n9285 = ~n9279 & n9284 ;
  assign n9286 = n9278 | n9285 ;
  assign n9287 = n1710 & n4050 ;
  assign n9288 = n1434 & n4555 ;
  assign n9289 = n9287 | n9288 ;
  assign n9290 = n1585 & n5392 ;
  assign n9291 = x40 & n9290 ;
  assign n9292 = ( x40 & ~n9289 ) | ( x40 & n9291 ) | ( ~n9289 & n9291 ) ;
  assign n9293 = x20 & n9292 ;
  assign n9294 = n9289 | n9290 ;
  assign n9295 = x21 & x39 ;
  assign n9296 = x22 & x38 ;
  assign n9297 = ( ~n9290 & n9295 ) | ( ~n9290 & n9296 ) | ( n9295 & n9296 ) ;
  assign n9298 = n9295 & n9296 ;
  assign n9299 = ( ~n9289 & n9297 ) | ( ~n9289 & n9298 ) | ( n9297 & n9298 ) ;
  assign n9300 = ~n9294 & n9299 ;
  assign n9301 = n9293 | n9300 ;
  assign n9302 = n9286 & n9301 ;
  assign n9303 = n9286 & ~n9302 ;
  assign n9304 = n9301 & ~n9302 ;
  assign n9305 = n9303 | n9304 ;
  assign n9306 = n2340 & n4914 ;
  assign n9307 = n1912 & n4078 ;
  assign n9308 = n9306 | n9307 ;
  assign n9309 = n2511 & n3483 ;
  assign n9310 = x36 & n9309 ;
  assign n9311 = ( x36 & ~n9308 ) | ( x36 & n9310 ) | ( ~n9308 & n9310 ) ;
  assign n9312 = x24 & n9311 ;
  assign n9313 = n9308 | n9309 ;
  assign n9314 = x25 & x35 ;
  assign n9315 = x26 & x34 ;
  assign n9316 = ( ~n9309 & n9314 ) | ( ~n9309 & n9315 ) | ( n9314 & n9315 ) ;
  assign n9317 = n9314 & n9315 ;
  assign n9318 = ( ~n9308 & n9316 ) | ( ~n9308 & n9317 ) | ( n9316 & n9317 ) ;
  assign n9319 = ~n9313 & n9318 ;
  assign n9320 = n9312 | n9319 ;
  assign n9321 = ~n9305 & n9320 ;
  assign n9322 = n9305 & ~n9320 ;
  assign n9323 = n9321 | n9322 ;
  assign n9324 = ( n8863 & n8865 ) | ( n8863 & n8870 ) | ( n8865 & n8870 ) ;
  assign n9325 = n9323 | n9324 ;
  assign n9326 = n9323 & n9324 ;
  assign n9327 = n9325 & ~n9326 ;
  assign n9328 = n1023 & n5658 ;
  assign n9329 = n7041 & n8437 ;
  assign n9330 = n9328 | n9329 ;
  assign n9331 = x44 & x51 ;
  assign n9332 = n754 & n9331 ;
  assign n9333 = x43 & n9332 ;
  assign n9334 = ( x43 & ~n9330 ) | ( x43 & n9333 ) | ( ~n9330 & n9333 ) ;
  assign n9335 = x17 & n9334 ;
  assign n9336 = n9330 | n9332 ;
  assign n9337 = x9 & x51 ;
  assign n9338 = x16 & x44 ;
  assign n9339 = ( ~n9332 & n9337 ) | ( ~n9332 & n9338 ) | ( n9337 & n9338 ) ;
  assign n9340 = n9337 & n9338 ;
  assign n9341 = ( ~n9330 & n9339 ) | ( ~n9330 & n9340 ) | ( n9339 & n9340 ) ;
  assign n9342 = ~n9336 & n9341 ;
  assign n9343 = ~n8932 & n9342 ;
  assign n9344 = ( ~n8932 & n9335 ) | ( ~n8932 & n9343 ) | ( n9335 & n9343 ) ;
  assign n9345 = n8932 & ~n9342 ;
  assign n9346 = ~n9335 & n9345 ;
  assign n9347 = n9344 | n9346 ;
  assign n9348 = n618 & n6834 ;
  assign n9349 = x45 & x50 ;
  assign n9350 = n582 & n9349 ;
  assign n9351 = n9348 | n9350 ;
  assign n9352 = x45 & x49 ;
  assign n9353 = n718 & n9352 ;
  assign n9354 = x50 & n9353 ;
  assign n9355 = ( x50 & ~n9351 ) | ( x50 & n9354 ) | ( ~n9351 & n9354 ) ;
  assign n9356 = x10 & n9355 ;
  assign n9357 = n9351 | n9353 ;
  assign n9358 = x11 & x49 ;
  assign n9359 = x15 & x45 ;
  assign n9360 = ( ~n9353 & n9358 ) | ( ~n9353 & n9359 ) | ( n9358 & n9359 ) ;
  assign n9361 = n9358 & n9359 ;
  assign n9362 = ( ~n9351 & n9360 ) | ( ~n9351 & n9361 ) | ( n9360 & n9361 ) ;
  assign n9363 = ~n9357 & n9362 ;
  assign n9364 = n9356 | n9363 ;
  assign n9365 = n9347 & n9364 ;
  assign n9366 = n9347 | n9364 ;
  assign n9367 = ~n9365 & n9366 ;
  assign n9368 = n9327 | n9367 ;
  assign n9369 = n9327 & n9367 ;
  assign n9370 = n9368 & ~n9369 ;
  assign n9373 = n9370 & n9372 ;
  assign n9374 = n9372 & ~n9373 ;
  assign n9375 = x0 & x60 ;
  assign n9376 = n9091 & n9375 ;
  assign n9377 = n9091 & ~n9376 ;
  assign n9378 = ~n9091 & n9375 ;
  assign n9379 = n9377 | n9378 ;
  assign n9380 = x1 & x59 ;
  assign n9381 = n3595 & n9380 ;
  assign n9382 = n9380 & ~n9381 ;
  assign n9383 = n3595 & ~n9381 ;
  assign n9384 = n9382 | n9383 ;
  assign n9385 = ~n9379 & n9384 ;
  assign n9386 = n9379 & ~n9384 ;
  assign n9387 = n9385 | n9386 ;
  assign n9388 = n2372 & n3321 ;
  assign n9389 = n4286 & n8099 ;
  assign n9390 = n9388 | n9389 ;
  assign n9391 = x23 & x37 ;
  assign n9392 = n6324 & n9391 ;
  assign n9393 = x33 & n9392 ;
  assign n9394 = ( x33 & ~n9390 ) | ( x33 & n9393 ) | ( ~n9390 & n9393 ) ;
  assign n9395 = x27 & n9394 ;
  assign n9396 = n9390 | n9392 ;
  assign n9397 = n6324 | n9391 ;
  assign n9398 = x27 | n9397 ;
  assign n9399 = ( n9394 & n9397 ) | ( n9394 & n9398 ) | ( n9397 & n9398 ) ;
  assign n9400 = ( n9395 & ~n9396 ) | ( n9395 & n9399 ) | ( ~n9396 & n9399 ) ;
  assign n9401 = n9387 & n9400 ;
  assign n9402 = n9387 | n9400 ;
  assign n9403 = ~n9401 & n9402 ;
  assign n9404 = n8777 | n9096 ;
  assign n9405 = ( n9096 & n9097 ) | ( n9096 & n9404 ) | ( n9097 & n9404 ) ;
  assign n9406 = n9403 | n9405 ;
  assign n9407 = n9403 & n9405 ;
  assign n9408 = n9406 & ~n9407 ;
  assign n9409 = x8 & x52 ;
  assign n9410 = x18 & x42 ;
  assign n9411 = n9409 & n9410 ;
  assign n9412 = n251 & n8161 ;
  assign n9413 = x18 & x53 ;
  assign n9414 = n6048 & n9413 ;
  assign n9415 = n9412 | n9414 ;
  assign n9416 = x53 & n9411 ;
  assign n9417 = ( x53 & ~n9415 ) | ( x53 & n9416 ) | ( ~n9415 & n9416 ) ;
  assign n9418 = x7 & n9417 ;
  assign n9419 = ( n9409 & n9410 ) | ( n9409 & ~n9415 ) | ( n9410 & ~n9415 ) ;
  assign n9420 = ( ~n9411 & n9418 ) | ( ~n9411 & n9419 ) | ( n9418 & n9419 ) ;
  assign n9421 = x46 & x48 ;
  assign n9422 = n487 & n9421 ;
  assign n9423 = n650 & n6147 ;
  assign n9424 = n9422 | n9423 ;
  assign n9425 = n647 & n6762 ;
  assign n9426 = n8128 & n9425 ;
  assign n9427 = ( n8128 & ~n9424 ) | ( n8128 & n9426 ) | ( ~n9424 & n9426 ) ;
  assign n9428 = n9424 | n9425 ;
  assign n9429 = x12 & x48 ;
  assign n9430 = x13 & x47 ;
  assign n9431 = ( ~n9425 & n9429 ) | ( ~n9425 & n9430 ) | ( n9429 & n9430 ) ;
  assign n9432 = n9429 & n9430 ;
  assign n9433 = ( ~n9424 & n9431 ) | ( ~n9424 & n9432 ) | ( n9431 & n9432 ) ;
  assign n9434 = ~n9428 & n9433 ;
  assign n9435 = n9427 | n9434 ;
  assign n9436 = n9420 & n9435 ;
  assign n9437 = n9420 & ~n9436 ;
  assign n9438 = x6 & x54 ;
  assign n9439 = x19 & x41 ;
  assign n9440 = n9438 & n9439 ;
  assign n9441 = x41 & x55 ;
  assign n9442 = n1444 & n9441 ;
  assign n9443 = n204 & n8357 ;
  assign n9444 = n9442 | n9443 ;
  assign n9445 = x55 & n9440 ;
  assign n9446 = ( x55 & ~n9444 ) | ( x55 & n9445 ) | ( ~n9444 & n9445 ) ;
  assign n9447 = x5 & n9446 ;
  assign n9448 = ( n9438 & n9439 ) | ( n9438 & ~n9444 ) | ( n9439 & ~n9444 ) ;
  assign n9449 = ( ~n9440 & n9447 ) | ( ~n9440 & n9448 ) | ( n9447 & n9448 ) ;
  assign n9450 = ~n9420 & n9435 ;
  assign n9451 = n9449 & n9450 ;
  assign n9452 = ( n9437 & n9449 ) | ( n9437 & n9451 ) | ( n9449 & n9451 ) ;
  assign n9453 = n9449 | n9450 ;
  assign n9454 = n9437 | n9453 ;
  assign n9455 = ~n9452 & n9454 ;
  assign n9456 = n9408 | n9455 ;
  assign n9457 = n9408 & n9455 ;
  assign n9458 = n9456 & ~n9457 ;
  assign n9459 = n9100 & n9116 ;
  assign n9460 = n9116 & ~n9459 ;
  assign n9461 = n9100 & ~n9459 ;
  assign n9462 = n9460 | n9461 ;
  assign n9463 = n9108 | n9459 ;
  assign n9464 = ( n9459 & n9462 ) | ( n9459 & n9463 ) | ( n9462 & n9463 ) ;
  assign n9465 = n9458 & n9464 ;
  assign n9466 = n9458 | n9464 ;
  assign n9467 = ~n9465 & n9466 ;
  assign n9468 = n9373 & n9467 ;
  assign n9469 = ~n9370 & n9467 ;
  assign n9470 = ( ~n9374 & n9468 ) | ( ~n9374 & n9469 ) | ( n9468 & n9469 ) ;
  assign n9471 = n9373 | n9467 ;
  assign n9472 = n9370 & ~n9467 ;
  assign n9473 = ( n9374 & ~n9471 ) | ( n9374 & n9472 ) | ( ~n9471 & n9472 ) ;
  assign n9474 = n9470 | n9473 ;
  assign n9475 = n9265 & ~n9266 ;
  assign n9476 = n9474 | n9475 ;
  assign n9477 = ( ~n8892 & n9474 ) | ( ~n8892 & n9476 ) | ( n9474 & n9476 ) ;
  assign n9478 = n9270 | n9477 ;
  assign n9479 = n9474 & n9475 ;
  assign n9480 = ~n8892 & n9479 ;
  assign n9481 = ( n9270 & n9474 ) | ( n9270 & n9480 ) | ( n9474 & n9480 ) ;
  assign n9482 = n9478 & ~n9481 ;
  assign n9483 = n9214 & n9482 ;
  assign n9484 = n9214 | n9482 ;
  assign n9485 = ~n9483 & n9484 ;
  assign n9486 = n8898 | n9152 ;
  assign n9487 = ( n8898 & n8899 ) | ( n8898 & n9486 ) | ( n8899 & n9486 ) ;
  assign n9488 = ( n9169 & n9485 ) | ( n9169 & ~n9487 ) | ( n9485 & ~n9487 ) ;
  assign n9489 = ( ~n9485 & n9487 ) | ( ~n9485 & n9488 ) | ( n9487 & n9488 ) ;
  assign n9490 = ( ~n9169 & n9488 ) | ( ~n9169 & n9489 ) | ( n9488 & n9489 ) ;
  assign n9491 = n9485 | n9487 ;
  assign n9492 = n9485 & n9487 ;
  assign n9493 = n9491 | n9492 ;
  assign n9494 = ( n9162 & n9492 ) | ( n9162 & n9493 ) | ( n9492 & n9493 ) ;
  assign n9495 = ( n9168 & n9493 ) | ( n9168 & n9494 ) | ( n9493 & n9494 ) ;
  assign n9496 = n7041 & n8988 ;
  assign n9497 = n1020 & n5658 ;
  assign n9498 = n9496 | n9497 ;
  assign n9499 = x44 & x52 ;
  assign n9500 = n1694 & n9499 ;
  assign n9501 = x43 & n9500 ;
  assign n9502 = ( x43 & ~n9498 ) | ( x43 & n9501 ) | ( ~n9498 & n9501 ) ;
  assign n9503 = x18 & n9502 ;
  assign n9504 = n9498 | n9500 ;
  assign n9505 = x9 & x52 ;
  assign n9506 = x17 & x44 ;
  assign n9507 = ( ~n9500 & n9505 ) | ( ~n9500 & n9506 ) | ( n9505 & n9506 ) ;
  assign n9508 = n9505 & n9506 ;
  assign n9509 = ( ~n9498 & n9507 ) | ( ~n9498 & n9508 ) | ( n9507 & n9508 ) ;
  assign n9510 = ~n9504 & n9509 ;
  assign n9511 = n9503 | n9510 ;
  assign n9512 = x7 & x54 ;
  assign n9513 = x8 & x53 ;
  assign n9514 = n9512 | n9513 ;
  assign n9515 = n251 & n8355 ;
  assign n9516 = n9514 | n9515 ;
  assign n9517 = x19 & x42 ;
  assign n9518 = ( ~n9515 & n9516 ) | ( ~n9515 & n9517 ) | ( n9516 & n9517 ) ;
  assign n9519 = ( n9515 & n9516 ) | ( n9515 & ~n9517 ) | ( n9516 & ~n9517 ) ;
  assign n9520 = ( ~n9516 & n9518 ) | ( ~n9516 & n9519 ) | ( n9518 & n9519 ) ;
  assign n9521 = n9511 & n9520 ;
  assign n9522 = n9511 & ~n9521 ;
  assign n9523 = n2895 & n3129 ;
  assign n9524 = n2267 & n3483 ;
  assign n9525 = n9523 | n9524 ;
  assign n9526 = n2372 & n4530 ;
  assign n9527 = x35 & n9526 ;
  assign n9528 = ( x35 & ~n9525 ) | ( x35 & n9527 ) | ( ~n9525 & n9527 ) ;
  assign n9529 = x26 & n9528 ;
  assign n9530 = n9525 | n9526 ;
  assign n9531 = x28 & x33 ;
  assign n9532 = ( n3693 & ~n9526 ) | ( n3693 & n9531 ) | ( ~n9526 & n9531 ) ;
  assign n9533 = n3693 & n9531 ;
  assign n9534 = ( ~n9525 & n9532 ) | ( ~n9525 & n9533 ) | ( n9532 & n9533 ) ;
  assign n9535 = ~n9530 & n9534 ;
  assign n9536 = n9529 | n9535 ;
  assign n9537 = ~n9511 & n9520 ;
  assign n9538 = n9536 & ~n9537 ;
  assign n9539 = ~n9522 & n9538 ;
  assign n9540 = ~n9536 & n9537 ;
  assign n9541 = ( n9522 & ~n9536 ) | ( n9522 & n9540 ) | ( ~n9536 & n9540 ) ;
  assign n9542 = n9539 | n9541 ;
  assign n9543 = n9248 & n9542 ;
  assign n9544 = ( n9253 & n9542 ) | ( n9253 & n9543 ) | ( n9542 & n9543 ) ;
  assign n9545 = n9542 & ~n9544 ;
  assign n9546 = n9248 | n9253 ;
  assign n9547 = ~n9544 & n9546 ;
  assign n9548 = n9545 | n9547 ;
  assign n9549 = n9224 | n9231 ;
  assign n9550 = ( n9224 & n9228 ) | ( n9224 & n9549 ) | ( n9228 & n9549 ) ;
  assign n9551 = ~n9548 & n9550 ;
  assign n9552 = n9548 & ~n9550 ;
  assign n9553 = n9551 | n9552 ;
  assign n9566 = n8943 | n9216 ;
  assign n9567 = ( n9216 & n9217 ) | ( n9216 & n9566 ) | ( n9217 & n9566 ) ;
  assign n9554 = x3 & x58 ;
  assign n9555 = x4 & x57 ;
  assign n9556 = n9554 | n9555 ;
  assign n9557 = n79 & n9272 ;
  assign n9558 = x23 & x38 ;
  assign n9559 = ~n9557 & n9558 ;
  assign n9560 = n9556 | n9557 ;
  assign n9561 = ( n9557 & n9559 ) | ( n9557 & n9560 ) | ( n9559 & n9560 ) ;
  assign n9562 = n9556 & ~n9561 ;
  assign n9563 = ~n9556 & n9558 ;
  assign n9564 = ( n9558 & ~n9559 ) | ( n9558 & n9563 ) | ( ~n9559 & n9563 ) ;
  assign n9565 = n9562 | n9564 ;
  assign n9568 = n9565 & n9567 ;
  assign n9569 = n9567 & ~n9568 ;
  assign n9570 = n9010 | n9243 ;
  assign n9571 = ( n9243 & n9244 ) | ( n9243 & n9570 ) | ( n9244 & n9570 ) ;
  assign n9572 = n9565 & ~n9567 ;
  assign n9573 = n9571 & n9572 ;
  assign n9574 = ( n9569 & n9571 ) | ( n9569 & n9573 ) | ( n9571 & n9573 ) ;
  assign n9575 = n9571 | n9572 ;
  assign n9576 = n9569 | n9575 ;
  assign n9577 = ~n9574 & n9576 ;
  assign n9578 = x1 & x60 ;
  assign n9579 = x31 & n9578 ;
  assign n9580 = x31 | n9578 ;
  assign n9581 = ~n9579 & n9580 ;
  assign n9582 = n9381 & n9581 ;
  assign n9583 = n9381 | n9581 ;
  assign n9584 = ~n9582 & n9583 ;
  assign n9585 = n9428 & n9584 ;
  assign n9586 = n9428 | n9584 ;
  assign n9587 = ~n9585 & n9586 ;
  assign n9588 = n9053 | n9237 ;
  assign n9589 = ( n9237 & n9238 ) | ( n9237 & n9588 ) | ( n9238 & n9588 ) ;
  assign n9590 = n9587 & n9589 ;
  assign n9591 = n9587 | n9589 ;
  assign n9592 = ~n9590 & n9591 ;
  assign n9593 = n9335 | n9342 ;
  assign n9594 = ( n8932 & n9364 ) | ( n8932 & n9593 ) | ( n9364 & n9593 ) ;
  assign n9595 = n9592 & n9594 ;
  assign n9596 = n9592 | n9594 ;
  assign n9597 = ~n9595 & n9596 ;
  assign n9598 = n9577 & n9597 ;
  assign n9599 = n9577 & ~n9598 ;
  assign n9600 = ( n9323 & n9324 ) | ( n9323 & n9367 ) | ( n9324 & n9367 ) ;
  assign n9601 = ~n9598 & n9600 ;
  assign n9602 = n9597 & n9600 ;
  assign n9603 = ( n9599 & n9601 ) | ( n9599 & n9602 ) | ( n9601 & n9602 ) ;
  assign n9604 = n9598 & ~n9600 ;
  assign n9605 = n9597 | n9600 ;
  assign n9606 = ( n9599 & ~n9604 ) | ( n9599 & n9605 ) | ( ~n9604 & n9605 ) ;
  assign n9607 = ~n9603 & n9606 ;
  assign n9608 = n9553 & n9607 ;
  assign n9609 = n9553 & ~n9608 ;
  assign n9610 = ~n9553 & n9607 ;
  assign n9611 = n9609 | n9610 ;
  assign n9612 = ~n9373 & n9467 ;
  assign n9613 = n9370 & n9467 ;
  assign n9614 = ( n9374 & n9612 ) | ( n9374 & n9613 ) | ( n9612 & n9613 ) ;
  assign n9615 = n9373 | n9614 ;
  assign n9616 = n9611 | n9615 ;
  assign n9617 = ~n9615 & n9616 ;
  assign n9618 = ( ~n9611 & n9616 ) | ( ~n9611 & n9617 ) | ( n9616 & n9617 ) ;
  assign n9619 = n9269 & n9618 ;
  assign n9620 = ( n9481 & n9618 ) | ( n9481 & n9619 ) | ( n9618 & n9619 ) ;
  assign n9621 = n9269 | n9481 ;
  assign n9622 = ~n9620 & n9621 ;
  assign n9623 = n9618 & ~n9620 ;
  assign n9624 = n9622 | n9623 ;
  assign n9625 = n9411 | n9415 ;
  assign n9626 = n9336 | n9625 ;
  assign n9627 = n9336 & n9625 ;
  assign n9628 = n9626 & ~n9627 ;
  assign n9629 = n9376 | n9384 ;
  assign n9630 = ( n9376 & n9379 ) | ( n9376 & n9629 ) | ( n9379 & n9629 ) ;
  assign n9631 = n9628 | n9630 ;
  assign n9632 = n9628 & n9630 ;
  assign n9633 = n9631 & ~n9632 ;
  assign n9634 = n9436 & n9633 ;
  assign n9635 = ( n9452 & n9633 ) | ( n9452 & n9634 ) | ( n9633 & n9634 ) ;
  assign n9636 = n9436 | n9633 ;
  assign n9637 = n9452 | n9636 ;
  assign n9638 = ~n9635 & n9637 ;
  assign n9639 = n9401 | n9405 ;
  assign n9640 = ( n9401 & n9403 ) | ( n9401 & n9639 ) | ( n9403 & n9639 ) ;
  assign n9641 = n9638 | n9640 ;
  assign n9642 = n9638 & n9640 ;
  assign n9643 = n9641 & ~n9642 ;
  assign n9644 = n9313 | n9396 ;
  assign n9645 = n9313 & n9396 ;
  assign n9646 = n9644 & ~n9645 ;
  assign n9647 = n9294 | n9646 ;
  assign n9648 = n9294 & n9646 ;
  assign n9649 = n9647 & ~n9648 ;
  assign n9650 = n9440 | n9444 ;
  assign n9651 = n9279 | n9650 ;
  assign n9652 = n9279 & n9650 ;
  assign n9653 = n9651 & ~n9652 ;
  assign n9654 = n9357 | n9653 ;
  assign n9655 = n9357 & n9653 ;
  assign n9656 = n9654 & ~n9655 ;
  assign n9657 = n9649 | n9656 ;
  assign n9658 = n9649 & n9656 ;
  assign n9659 = n9657 & ~n9658 ;
  assign n9660 = n9302 | n9320 ;
  assign n9661 = ( n9302 & n9305 ) | ( n9302 & n9660 ) | ( n9305 & n9660 ) ;
  assign n9662 = n9659 & n9661 ;
  assign n9663 = n9659 | n9661 ;
  assign n9664 = ~n9662 & n9663 ;
  assign n9665 = n9643 & n9664 ;
  assign n9666 = n9643 | n9664 ;
  assign n9667 = ~n9665 & n9666 ;
  assign n9668 = n9457 | n9464 ;
  assign n9669 = ( n9457 & n9458 ) | ( n9457 & n9668 ) | ( n9458 & n9668 ) ;
  assign n9670 = n9667 & n9669 ;
  assign n9671 = ~n9667 & n9669 ;
  assign n9672 = ( n9667 & ~n9670 ) | ( n9667 & n9671 ) | ( ~n9670 & n9671 ) ;
  assign n9673 = n9196 | n9672 ;
  assign n9674 = n9138 | n9672 ;
  assign n9675 = ( n9197 & n9673 ) | ( n9197 & n9674 ) | ( n9673 & n9674 ) ;
  assign n9676 = n9205 | n9675 ;
  assign n9677 = n9196 & n9672 ;
  assign n9678 = n9138 & n9672 ;
  assign n9679 = ( n9197 & n9677 ) | ( n9197 & n9678 ) | ( n9677 & n9678 ) ;
  assign n9680 = ( n9205 & n9672 ) | ( n9205 & n9679 ) | ( n9672 & n9679 ) ;
  assign n9681 = n9676 & ~n9680 ;
  assign n9682 = n9260 | n9264 ;
  assign n9683 = x14 & x50 ;
  assign n9684 = n8778 & n9683 ;
  assign n9685 = n490 & n6834 ;
  assign n9686 = n9684 | n9685 ;
  assign n9687 = n487 & n6757 ;
  assign n9688 = x50 & n9687 ;
  assign n9689 = ( x50 & ~n9686 ) | ( x50 & n9688 ) | ( ~n9686 & n9688 ) ;
  assign n9690 = x11 & n9689 ;
  assign n9691 = n9686 | n9687 ;
  assign n9692 = x12 & x49 ;
  assign n9693 = ( n8125 & ~n9687 ) | ( n8125 & n9692 ) | ( ~n9687 & n9692 ) ;
  assign n9694 = n8125 & n9692 ;
  assign n9695 = ( ~n9686 & n9693 ) | ( ~n9686 & n9694 ) | ( n9693 & n9694 ) ;
  assign n9696 = ~n9691 & n9695 ;
  assign n9697 = n9690 | n9696 ;
  assign n9698 = n795 & n5975 ;
  assign n9699 = x10 & x51 ;
  assign n9700 = n6304 & n9699 ;
  assign n9701 = n9698 | n9700 ;
  assign n9702 = x46 & x51 ;
  assign n9703 = n582 & n9702 ;
  assign n9704 = n6304 & n9703 ;
  assign n9705 = ( n6304 & ~n9701 ) | ( n6304 & n9704 ) | ( ~n9701 & n9704 ) ;
  assign n9706 = n9701 | n9703 ;
  assign n9707 = x15 & x46 ;
  assign n9708 = ( n9699 & ~n9703 ) | ( n9699 & n9707 ) | ( ~n9703 & n9707 ) ;
  assign n9709 = n9699 & n9707 ;
  assign n9710 = ( ~n9701 & n9708 ) | ( ~n9701 & n9709 ) | ( n9708 & n9709 ) ;
  assign n9711 = ~n9706 & n9710 ;
  assign n9712 = n9705 | n9711 ;
  assign n9713 = n9697 & n9712 ;
  assign n9714 = n9697 & ~n9713 ;
  assign n9715 = x29 & x32 ;
  assign n9716 = n2965 | n9715 ;
  assign n9717 = n2709 & n4062 ;
  assign n9718 = x13 & x48 ;
  assign n9719 = ~n9717 & n9718 ;
  assign n9720 = n9716 | n9717 ;
  assign n9721 = ( n9717 & n9719 ) | ( n9717 & n9720 ) | ( n9719 & n9720 ) ;
  assign n9722 = n9716 & ~n9721 ;
  assign n9723 = ~n9716 & n9718 ;
  assign n9724 = ( n9718 & ~n9719 ) | ( n9718 & n9723 ) | ( ~n9719 & n9723 ) ;
  assign n9725 = n9722 | n9724 ;
  assign n9726 = ~n9697 & n9712 ;
  assign n9727 = n9725 & n9726 ;
  assign n9728 = ( n9714 & n9725 ) | ( n9714 & n9727 ) | ( n9725 & n9727 ) ;
  assign n9729 = n9725 | n9726 ;
  assign n9730 = n9714 | n9729 ;
  assign n9731 = ~n9728 & n9730 ;
  assign n9732 = n9175 | n9183 ;
  assign n9733 = ( n9175 & n9176 ) | ( n9175 & n9732 ) | ( n9176 & n9732 ) ;
  assign n9734 = n9731 | n9733 ;
  assign n9735 = n9731 & n9733 ;
  assign n9736 = n9734 & ~n9735 ;
  assign n9737 = x59 & x61 ;
  assign n9738 = n67 & n9737 ;
  assign n9739 = x5 & x61 ;
  assign n9740 = n8148 & n9739 ;
  assign n9741 = n9738 | n9740 ;
  assign n9742 = x5 & x59 ;
  assign n9743 = n8712 & n9742 ;
  assign n9744 = x61 & n9743 ;
  assign n9745 = ( x61 & ~n9741 ) | ( x61 & n9744 ) | ( ~n9741 & n9744 ) ;
  assign n9746 = x0 & n9745 ;
  assign n9747 = n9741 | n9743 ;
  assign n9748 = x2 & x59 ;
  assign n9749 = x5 & x56 ;
  assign n9750 = ( ~n9743 & n9748 ) | ( ~n9743 & n9749 ) | ( n9748 & n9749 ) ;
  assign n9751 = n9748 & n9749 ;
  assign n9752 = ( ~n9741 & n9750 ) | ( ~n9741 & n9751 ) | ( n9750 & n9751 ) ;
  assign n9753 = ~n9747 & n9752 ;
  assign n9754 = n9746 | n9753 ;
  assign n9755 = x20 & x41 ;
  assign n9756 = x21 & x40 ;
  assign n9757 = n9755 | n9756 ;
  assign n9758 = n1434 & n5813 ;
  assign n9759 = x6 & x55 ;
  assign n9760 = ~n9758 & n9759 ;
  assign n9761 = n9757 | n9758 ;
  assign n9762 = ( n9758 & n9760 ) | ( n9758 & n9761 ) | ( n9760 & n9761 ) ;
  assign n9763 = n9757 & ~n9762 ;
  assign n9764 = ~n9757 & n9759 ;
  assign n9765 = ( n9759 & ~n9760 ) | ( n9759 & n9764 ) | ( ~n9760 & n9764 ) ;
  assign n9766 = n9763 | n9765 ;
  assign n9767 = n9754 & n9766 ;
  assign n9768 = n9754 & ~n9767 ;
  assign n9769 = n9766 & ~n9767 ;
  assign n9770 = n9768 | n9769 ;
  assign n9771 = x36 & x39 ;
  assign n9772 = n5695 & n9771 ;
  assign n9773 = n2148 & n5798 ;
  assign n9774 = n9772 | n9773 ;
  assign n9775 = n1912 & n3770 ;
  assign n9776 = x39 & n9775 ;
  assign n9777 = ( x39 & ~n9774 ) | ( x39 & n9776 ) | ( ~n9774 & n9776 ) ;
  assign n9778 = x22 & n9777 ;
  assign n9779 = n9774 | n9775 ;
  assign n9780 = x24 & x37 ;
  assign n9781 = x25 & x36 ;
  assign n9782 = ( ~n9775 & n9780 ) | ( ~n9775 & n9781 ) | ( n9780 & n9781 ) ;
  assign n9783 = n9780 & n9781 ;
  assign n9784 = ( ~n9774 & n9782 ) | ( ~n9774 & n9783 ) | ( n9782 & n9783 ) ;
  assign n9785 = ~n9779 & n9784 ;
  assign n9786 = n9778 | n9785 ;
  assign n9787 = ~n9770 & n9786 ;
  assign n9788 = n9770 & ~n9786 ;
  assign n9789 = n9787 | n9788 ;
  assign n9790 = n9736 | n9789 ;
  assign n9791 = n9736 & n9789 ;
  assign n9792 = n9790 & ~n9791 ;
  assign n9793 = n9190 | n9193 ;
  assign n9794 = ( n9190 & n9191 ) | ( n9190 & n9793 ) | ( n9191 & n9793 ) ;
  assign n9795 = n9792 & n9794 ;
  assign n9796 = n9792 | n9794 ;
  assign n9797 = ~n9795 & n9796 ;
  assign n9798 = n9682 & n9797 ;
  assign n9799 = n9682 | n9797 ;
  assign n9800 = ~n9798 & n9799 ;
  assign n9801 = n9681 & n9800 ;
  assign n9802 = n9681 | n9800 ;
  assign n9803 = ~n9801 & n9802 ;
  assign n9804 = n9624 | n9803 ;
  assign n9805 = n9624 & ~n9803 ;
  assign n9806 = ( ~n9624 & n9804 ) | ( ~n9624 & n9805 ) | ( n9804 & n9805 ) ;
  assign n9807 = n9213 | n9483 ;
  assign n9808 = ( n9495 & n9806 ) | ( n9495 & ~n9807 ) | ( n9806 & ~n9807 ) ;
  assign n9809 = ( ~n9806 & n9807 ) | ( ~n9806 & n9808 ) | ( n9807 & n9808 ) ;
  assign n9810 = ( ~n9495 & n9808 ) | ( ~n9495 & n9809 ) | ( n9808 & n9809 ) ;
  assign n9811 = n9428 | n9582 ;
  assign n9812 = ( n9582 & n9584 ) | ( n9582 & n9811 ) | ( n9584 & n9811 ) ;
  assign n9813 = n9627 & n9812 ;
  assign n9814 = ( n9632 & n9812 ) | ( n9632 & n9813 ) | ( n9812 & n9813 ) ;
  assign n9815 = n9627 | n9812 ;
  assign n9816 = n9632 | n9815 ;
  assign n9817 = ~n9814 & n9816 ;
  assign n9818 = n9294 | n9645 ;
  assign n9819 = ( n9645 & n9646 ) | ( n9645 & n9818 ) | ( n9646 & n9818 ) ;
  assign n9820 = n9817 | n9819 ;
  assign n9821 = n9817 & n9819 ;
  assign n9822 = n9820 & ~n9821 ;
  assign n9823 = n9735 | n9789 ;
  assign n9824 = ( n9735 & n9736 ) | ( n9735 & n9823 ) | ( n9736 & n9823 ) ;
  assign n9825 = n9822 & ~n9824 ;
  assign n9826 = n9504 | n9706 ;
  assign n9827 = n9504 & n9706 ;
  assign n9828 = n9826 & ~n9827 ;
  assign n9829 = x57 & x59 ;
  assign n9830 = n169 & n9829 ;
  assign n9831 = x58 & x59 ;
  assign n9832 = n79 & n9831 ;
  assign n9833 = n9830 | n9832 ;
  assign n9834 = n91 & n9272 ;
  assign n9835 = x59 & n9834 ;
  assign n9836 = ( x59 & ~n9833 ) | ( x59 & n9835 ) | ( ~n9833 & n9835 ) ;
  assign n9837 = x3 & n9836 ;
  assign n9838 = n9833 | n9834 ;
  assign n9839 = x4 & x58 ;
  assign n9840 = x5 & x57 ;
  assign n9841 = ( ~n9834 & n9839 ) | ( ~n9834 & n9840 ) | ( n9839 & n9840 ) ;
  assign n9842 = n9839 & n9840 ;
  assign n9843 = ( ~n9833 & n9841 ) | ( ~n9833 & n9842 ) | ( n9841 & n9842 ) ;
  assign n9844 = ~n9838 & n9843 ;
  assign n9845 = n9837 | n9844 ;
  assign n9846 = n9828 & n9845 ;
  assign n9847 = n9828 & ~n9846 ;
  assign n9848 = n9845 & ~n9846 ;
  assign n9849 = n9847 | n9848 ;
  assign n9850 = n9536 & n9537 ;
  assign n9851 = ( n9522 & n9536 ) | ( n9522 & n9850 ) | ( n9536 & n9850 ) ;
  assign n9852 = n9521 | n9851 ;
  assign n9853 = n9849 | n9852 ;
  assign n9854 = n9849 & n9852 ;
  assign n9855 = n9853 & ~n9854 ;
  assign n9856 = n9568 | n9574 ;
  assign n9857 = n9855 | n9856 ;
  assign n9858 = n9855 & n9856 ;
  assign n9859 = n9857 & ~n9858 ;
  assign n9860 = ( n9824 & n9825 ) | ( n9824 & n9859 ) | ( n9825 & n9859 ) ;
  assign n9861 = ( ~n9822 & n9825 ) | ( ~n9822 & n9860 ) | ( n9825 & n9860 ) ;
  assign n9862 = n9822 & n9824 ;
  assign n9863 = n9824 & ~n9862 ;
  assign n9864 = n9825 | n9859 ;
  assign n9865 = n9863 | n9864 ;
  assign n9866 = ~n9861 & n9865 ;
  assign n9867 = n9611 & n9615 ;
  assign n9868 = n9608 & n9866 ;
  assign n9869 = ( n9866 & n9867 ) | ( n9866 & n9868 ) | ( n9867 & n9868 ) ;
  assign n9870 = n9608 | n9866 ;
  assign n9871 = n9867 | n9870 ;
  assign n9872 = ~n9869 & n9871 ;
  assign n9873 = n9598 | n9603 ;
  assign n9874 = n1077 & n5658 ;
  assign n9875 = x19 & x54 ;
  assign n9876 = n6662 & n9875 ;
  assign n9877 = n9874 | n9876 ;
  assign n9878 = x18 & x54 ;
  assign n9879 = n6992 & n9878 ;
  assign n9880 = x43 & n9879 ;
  assign n9881 = ( x43 & ~n9877 ) | ( x43 & n9880 ) | ( ~n9877 & n9880 ) ;
  assign n9882 = x19 & n9881 ;
  assign n9883 = n9877 | n9879 ;
  assign n9884 = x8 & x54 ;
  assign n9885 = x18 & x44 ;
  assign n9886 = ( ~n9879 & n9884 ) | ( ~n9879 & n9885 ) | ( n9884 & n9885 ) ;
  assign n9887 = n9884 & n9885 ;
  assign n9888 = ( ~n9877 & n9886 ) | ( ~n9877 & n9887 ) | ( n9886 & n9887 ) ;
  assign n9889 = ~n9883 & n9888 ;
  assign n9890 = n9882 | n9889 ;
  assign n9891 = n2075 & n3129 ;
  assign n9892 = n2372 & n3483 ;
  assign n9893 = n9891 | n9892 ;
  assign n9894 = n2369 & n4530 ;
  assign n9895 = x35 & n9894 ;
  assign n9896 = ( x35 & ~n9893 ) | ( x35 & n9895 ) | ( ~n9893 & n9895 ) ;
  assign n9897 = x27 & n9896 ;
  assign n9898 = n9893 | n9894 ;
  assign n9899 = x28 & x34 ;
  assign n9900 = x29 & x33 ;
  assign n9901 = ( ~n9894 & n9899 ) | ( ~n9894 & n9900 ) | ( n9899 & n9900 ) ;
  assign n9902 = n9899 & n9900 ;
  assign n9903 = ( ~n9893 & n9901 ) | ( ~n9893 & n9902 ) | ( n9901 & n9902 ) ;
  assign n9904 = ~n9898 & n9903 ;
  assign n9905 = n9897 | n9904 ;
  assign n9906 = n9890 & n9905 ;
  assign n9907 = n9890 & ~n9906 ;
  assign n9908 = n9905 & ~n9906 ;
  assign n9909 = n9907 | n9908 ;
  assign n9910 = n2148 & n4050 ;
  assign n9911 = n1932 & n4555 ;
  assign n9912 = n9910 | n9911 ;
  assign n9913 = n1686 & n5392 ;
  assign n9914 = x40 & n9913 ;
  assign n9915 = ( x40 & ~n9912 ) | ( x40 & n9914 ) | ( ~n9912 & n9914 ) ;
  assign n9916 = x22 & n9915 ;
  assign n9917 = n9912 | n9913 ;
  assign n9918 = x23 & x39 ;
  assign n9919 = x24 & x38 ;
  assign n9920 = ( ~n9913 & n9918 ) | ( ~n9913 & n9919 ) | ( n9918 & n9919 ) ;
  assign n9921 = n9918 & n9919 ;
  assign n9922 = ( ~n9912 & n9920 ) | ( ~n9912 & n9921 ) | ( n9920 & n9921 ) ;
  assign n9923 = ~n9917 & n9922 ;
  assign n9924 = n9916 | n9923 ;
  assign n9925 = ~n9909 & n9924 ;
  assign n9926 = n9909 & ~n9924 ;
  assign n9927 = n9925 | n9926 ;
  assign n9928 = x0 & x62 ;
  assign n9929 = x2 & x60 ;
  assign n9930 = n9928 | n9929 ;
  assign n9931 = x60 & x62 ;
  assign n9932 = n67 & n9931 ;
  assign n9933 = n9930 & ~n9932 ;
  assign n9934 = n9579 | n9932 ;
  assign n9935 = ( n9932 & n9933 ) | ( n9932 & n9934 ) | ( n9933 & n9934 ) ;
  assign n9936 = n9930 & ~n9935 ;
  assign n9937 = n9579 & ~n9933 ;
  assign n9938 = n9936 | n9937 ;
  assign n9939 = x25 & x37 ;
  assign n9940 = x26 & x36 ;
  assign n9941 = n9939 | n9940 ;
  assign n9942 = n2511 & n3770 ;
  assign n9943 = x21 & x41 ;
  assign n9944 = ~n9942 & n9943 ;
  assign n9945 = n9941 | n9942 ;
  assign n9946 = ( n9942 & n9944 ) | ( n9942 & n9945 ) | ( n9944 & n9945 ) ;
  assign n9947 = n9941 & ~n9946 ;
  assign n9948 = ~n9941 & n9943 ;
  assign n9949 = ( n9943 & ~n9944 ) | ( n9943 & n9948 ) | ( ~n9944 & n9948 ) ;
  assign n9950 = n9947 | n9949 ;
  assign n9951 = n9938 & n9950 ;
  assign n9952 = n9938 & ~n9951 ;
  assign n9953 = n9950 & ~n9951 ;
  assign n9954 = n9952 | n9953 ;
  assign n9955 = n360 & n8161 ;
  assign n9956 = x17 & x53 ;
  assign n9957 = n7551 & n9956 ;
  assign n9958 = n9955 | n9957 ;
  assign n9959 = x45 & x52 ;
  assign n9960 = n1860 & n9959 ;
  assign n9961 = x53 & n9960 ;
  assign n9962 = ( x53 & ~n9958 ) | ( x53 & n9961 ) | ( ~n9958 & n9961 ) ;
  assign n9963 = x9 & n9962 ;
  assign n9964 = n9958 | n9960 ;
  assign n9965 = x10 & x52 ;
  assign n9966 = x17 & x45 ;
  assign n9967 = ( ~n9960 & n9965 ) | ( ~n9960 & n9966 ) | ( n9965 & n9966 ) ;
  assign n9968 = n9965 & n9966 ;
  assign n9969 = ( ~n9958 & n9967 ) | ( ~n9958 & n9968 ) | ( n9967 & n9968 ) ;
  assign n9970 = ~n9964 & n9969 ;
  assign n9971 = n9963 | n9970 ;
  assign n9972 = ~n9954 & n9971 ;
  assign n9973 = n9954 & ~n9971 ;
  assign n9974 = n9972 | n9973 ;
  assign n9975 = n1846 & n9702 ;
  assign n9976 = n795 & n6147 ;
  assign n9977 = n9975 | n9976 ;
  assign n9978 = x47 & x51 ;
  assign n9979 = n718 & n9978 ;
  assign n9980 = x46 & n9979 ;
  assign n9981 = ( x46 & ~n9977 ) | ( x46 & n9980 ) | ( ~n9977 & n9980 ) ;
  assign n9982 = x16 & n9981 ;
  assign n9983 = n9977 | n9979 ;
  assign n9984 = x11 & x51 ;
  assign n9985 = x15 & x47 ;
  assign n9986 = ( ~n9979 & n9984 ) | ( ~n9979 & n9985 ) | ( n9984 & n9985 ) ;
  assign n9987 = n9984 & n9985 ;
  assign n9988 = ( ~n9977 & n9986 ) | ( ~n9977 & n9987 ) | ( n9986 & n9987 ) ;
  assign n9989 = ~n9983 & n9988 ;
  assign n9990 = n9982 | n9989 ;
  assign n9991 = n487 & n6345 ;
  assign n9992 = n647 & n6834 ;
  assign n9993 = n9991 | n9992 ;
  assign n9994 = n650 & n6759 ;
  assign n9995 = x50 & n9994 ;
  assign n9996 = ( x50 & ~n9993 ) | ( x50 & n9995 ) | ( ~n9993 & n9995 ) ;
  assign n9997 = x12 & n9996 ;
  assign n9998 = n9993 | n9994 ;
  assign n9999 = x13 & x49 ;
  assign n10000 = x14 & x48 ;
  assign n10001 = ( ~n9994 & n9999 ) | ( ~n9994 & n10000 ) | ( n9999 & n10000 ) ;
  assign n10002 = n9999 & n10000 ;
  assign n10003 = ( ~n9993 & n10001 ) | ( ~n9993 & n10002 ) | ( n10001 & n10002 ) ;
  assign n10004 = ~n9998 & n10003 ;
  assign n10005 = n9997 | n10004 ;
  assign n10006 = n9990 & n10005 ;
  assign n10007 = n9990 & ~n10006 ;
  assign n10008 = n10005 & ~n10006 ;
  assign n10009 = n10007 | n10008 ;
  assign n10010 = x6 & x56 ;
  assign n10011 = x7 & x55 ;
  assign n10012 = n10010 | n10011 ;
  assign n10013 = x55 & x56 ;
  assign n10014 = n200 & n10013 ;
  assign n10015 = x20 & x42 ;
  assign n10016 = ~n10014 & n10015 ;
  assign n10017 = n10012 | n10014 ;
  assign n10018 = ( n10014 & n10016 ) | ( n10014 & n10017 ) | ( n10016 & n10017 ) ;
  assign n10019 = n10012 & ~n10018 ;
  assign n10020 = ( ~n10012 & n10014 ) | ( ~n10012 & n10015 ) | ( n10014 & n10015 ) ;
  assign n10021 = n10015 & n10020 ;
  assign n10022 = n10019 | n10021 ;
  assign n10023 = ~n10009 & n10022 ;
  assign n10024 = n10009 & ~n10022 ;
  assign n10025 = n10023 | n10024 ;
  assign n10026 = n9974 & ~n10025 ;
  assign n10027 = ~n9974 & n10025 ;
  assign n10028 = n10026 | n10027 ;
  assign n10029 = n9927 & n10028 ;
  assign n10030 = n9927 | n10028 ;
  assign n10031 = ~n10029 & n10030 ;
  assign n10032 = n9873 & n10031 ;
  assign n10033 = n9873 & ~n10032 ;
  assign n10034 = n9665 | n9669 ;
  assign n10035 = ( n9665 & n9667 ) | ( n9665 & n10034 ) | ( n9667 & n10034 ) ;
  assign n10036 = ~n9873 & n10031 ;
  assign n10037 = n10035 & n10036 ;
  assign n10038 = ( n10033 & n10035 ) | ( n10033 & n10037 ) | ( n10035 & n10037 ) ;
  assign n10039 = n10035 | n10036 ;
  assign n10040 = n10033 | n10039 ;
  assign n10041 = ~n10038 & n10040 ;
  assign n10042 = n9872 | n10041 ;
  assign n10043 = n9872 & n10041 ;
  assign n10044 = n10042 & ~n10043 ;
  assign n10045 = n9198 | n9205 ;
  assign n10046 = ( n9672 & n9800 ) | ( n9672 & n10045 ) | ( n9800 & n10045 ) ;
  assign n10047 = n9590 | n9594 ;
  assign n10048 = ( n9590 & n9592 ) | ( n9590 & n10047 ) | ( n9592 & n10047 ) ;
  assign n10049 = n9658 & n10048 ;
  assign n10050 = ( n9662 & n10048 ) | ( n9662 & n10049 ) | ( n10048 & n10049 ) ;
  assign n10051 = n9658 | n10048 ;
  assign n10052 = n9662 | n10051 ;
  assign n10053 = ~n10050 & n10052 ;
  assign n10054 = n9635 | n9640 ;
  assign n10055 = ( n9635 & n9638 ) | ( n9635 & n10054 ) | ( n9638 & n10054 ) ;
  assign n10056 = n10053 | n10055 ;
  assign n10057 = n10053 & n10055 ;
  assign n10058 = n10056 & ~n10057 ;
  assign n10059 = n9792 | n10058 ;
  assign n10060 = ( n9794 & n10058 ) | ( n9794 & n10059 ) | ( n10058 & n10059 ) ;
  assign n10061 = n9798 | n10060 ;
  assign n10062 = n9767 | n9786 ;
  assign n10063 = n9357 | n9652 ;
  assign n10064 = ( n9652 & n9653 ) | ( n9652 & n10063 ) | ( n9653 & n10063 ) ;
  assign n10065 = n10062 & n10064 ;
  assign n10066 = n9767 & n10064 ;
  assign n10067 = ( n9770 & n10065 ) | ( n9770 & n10066 ) | ( n10065 & n10066 ) ;
  assign n10068 = n10062 | n10064 ;
  assign n10069 = n9767 | n10064 ;
  assign n10070 = ( n9770 & n10068 ) | ( n9770 & n10069 ) | ( n10068 & n10069 ) ;
  assign n10071 = ~n10067 & n10070 ;
  assign n10072 = n9713 | n9728 ;
  assign n10073 = n10071 | n10072 ;
  assign n10074 = n10071 & n10072 ;
  assign n10075 = n10073 & ~n10074 ;
  assign n10076 = n9530 | n9561 ;
  assign n10077 = n9530 & n9561 ;
  assign n10078 = n10076 & ~n10077 ;
  assign n10079 = n9779 | n10078 ;
  assign n10080 = n9779 & n10078 ;
  assign n10081 = n10079 & ~n10080 ;
  assign n10082 = x1 & x61 ;
  assign n10083 = n2546 & n10082 ;
  assign n10084 = n2546 | n10082 ;
  assign n10085 = ~n10083 & n10084 ;
  assign n10086 = n9721 | n10085 ;
  assign n10087 = n9721 & n10085 ;
  assign n10088 = n10086 & ~n10087 ;
  assign n10089 = n9691 & n10088 ;
  assign n10090 = n9691 | n10088 ;
  assign n10091 = ~n10089 & n10090 ;
  assign n10092 = n10081 & n10091 ;
  assign n10093 = n10081 & ~n10092 ;
  assign n10094 = ~n9515 & n9517 ;
  assign n10095 = ( n9515 & n9516 ) | ( n9515 & n10094 ) | ( n9516 & n10094 ) ;
  assign n10096 = n9747 | n9762 ;
  assign n10097 = n9747 & n9762 ;
  assign n10098 = n10096 & ~n10097 ;
  assign n10099 = n10095 | n10098 ;
  assign n10100 = n10095 & n10098 ;
  assign n10101 = n10099 & ~n10100 ;
  assign n10102 = n10092 & n10101 ;
  assign n10103 = ~n10091 & n10101 ;
  assign n10104 = ( ~n10093 & n10102 ) | ( ~n10093 & n10103 ) | ( n10102 & n10103 ) ;
  assign n10105 = n10092 | n10101 ;
  assign n10106 = n10091 & ~n10101 ;
  assign n10107 = ( n10093 & ~n10105 ) | ( n10093 & n10106 ) | ( ~n10105 & n10106 ) ;
  assign n10108 = n10104 | n10107 ;
  assign n10109 = n10075 & n10108 ;
  assign n10110 = ~n10075 & n10108 ;
  assign n10111 = ( n10075 & ~n10109 ) | ( n10075 & n10110 ) | ( ~n10109 & n10110 ) ;
  assign n10112 = n9544 | n9550 ;
  assign n10113 = ( n9544 & n9548 ) | ( n9544 & n10112 ) | ( n9548 & n10112 ) ;
  assign n10114 = n10111 | n10113 ;
  assign n10115 = n10111 & n10113 ;
  assign n10116 = n10114 & ~n10115 ;
  assign n10117 = ( n9260 & n9792 ) | ( n9260 & n9794 ) | ( n9792 & n9794 ) ;
  assign n10118 = ( n9264 & n9796 ) | ( n9264 & n10117 ) | ( n9796 & n10117 ) ;
  assign n10119 = ~n10058 & n10116 ;
  assign n10120 = ( n10116 & ~n10118 ) | ( n10116 & n10119 ) | ( ~n10118 & n10119 ) ;
  assign n10121 = n10061 & n10120 ;
  assign n10122 = n10058 & ~n10116 ;
  assign n10123 = n10118 & n10122 ;
  assign n10124 = ( n10061 & n10116 ) | ( n10061 & ~n10123 ) | ( n10116 & ~n10123 ) ;
  assign n10125 = ~n10121 & n10124 ;
  assign n10126 = n10046 & n10125 ;
  assign n10127 = n10046 & ~n10126 ;
  assign n10128 = ~n10046 & n10125 ;
  assign n10129 = n10127 | n10128 ;
  assign n10130 = n10044 & n10129 ;
  assign n10131 = n10044 | n10129 ;
  assign n10132 = ~n10130 & n10131 ;
  assign n10133 = n9620 | n9803 ;
  assign n10134 = ( n9620 & n9624 ) | ( n9620 & n10133 ) | ( n9624 & n10133 ) ;
  assign n10135 = n10132 & n10134 ;
  assign n10136 = n10132 | n10134 ;
  assign n10137 = ~n10135 & n10136 ;
  assign n10138 = n9806 & n9807 ;
  assign n10139 = n9806 | n9807 ;
  assign n10140 = n9494 & n10139 ;
  assign n10141 = n9493 & n10139 ;
  assign n10142 = ( n9168 & n10140 ) | ( n9168 & n10141 ) | ( n10140 & n10141 ) ;
  assign n10143 = n10138 | n10142 ;
  assign n10144 = n10137 | n10143 ;
  assign n10145 = n10136 & n10138 ;
  assign n10146 = ( n10136 & n10140 ) | ( n10136 & n10145 ) | ( n10140 & n10145 ) ;
  assign n10147 = ( n10136 & n10141 ) | ( n10136 & n10145 ) | ( n10141 & n10145 ) ;
  assign n10148 = ( n9168 & n10146 ) | ( n9168 & n10147 ) | ( n10146 & n10147 ) ;
  assign n10149 = ~n10135 & n10148 ;
  assign n10150 = n10144 & ~n10149 ;
  assign n10151 = n10135 | n10148 ;
  assign n10152 = ~n10092 & n10101 ;
  assign n10153 = n10091 & n10101 ;
  assign n10154 = ( n10093 & n10152 ) | ( n10093 & n10153 ) | ( n10152 & n10153 ) ;
  assign n10155 = n10092 | n10154 ;
  assign n10156 = n10067 | n10072 ;
  assign n10157 = ( n10067 & n10071 ) | ( n10067 & n10156 ) | ( n10071 & n10156 ) ;
  assign n10158 = n10155 | n10157 ;
  assign n10159 = n10155 & n10157 ;
  assign n10160 = n10158 & ~n10159 ;
  assign n10161 = n9854 | n9856 ;
  assign n10162 = ( n9854 & n9855 ) | ( n9854 & n10161 ) | ( n9855 & n10161 ) ;
  assign n10163 = n10160 | n10162 ;
  assign n10164 = n10160 & n10162 ;
  assign n10165 = n10163 & ~n10164 ;
  assign n10166 = n9827 | n9846 ;
  assign n10167 = n9779 | n10077 ;
  assign n10168 = ( n10077 & n10078 ) | ( n10077 & n10167 ) | ( n10078 & n10167 ) ;
  assign n10169 = n10166 | n10168 ;
  assign n10170 = n10166 & n10168 ;
  assign n10171 = n10169 & ~n10170 ;
  assign n10172 = n9691 | n10087 ;
  assign n10173 = ( n10087 & n10088 ) | ( n10087 & n10172 ) | ( n10088 & n10172 ) ;
  assign n10174 = n10171 | n10173 ;
  assign n10175 = n10171 & n10173 ;
  assign n10176 = n10174 & ~n10175 ;
  assign n10177 = ( n9927 & n9974 ) | ( n9927 & n10025 ) | ( n9974 & n10025 ) ;
  assign n10178 = n10176 | n10177 ;
  assign n10179 = n10176 & n10177 ;
  assign n10180 = n10178 & ~n10179 ;
  assign n10181 = n9917 | n10018 ;
  assign n10182 = n9917 & n10018 ;
  assign n10183 = n10181 & ~n10182 ;
  assign n10184 = n9998 | n10183 ;
  assign n10185 = n9998 & n10183 ;
  assign n10186 = n10184 & ~n10185 ;
  assign n10187 = n9838 | n9946 ;
  assign n10188 = n9838 & n9946 ;
  assign n10189 = n10187 & ~n10188 ;
  assign n10190 = n9935 | n10189 ;
  assign n10191 = n9935 & n10189 ;
  assign n10192 = n10190 & ~n10191 ;
  assign n10193 = n10095 | n10097 ;
  assign n10194 = ( n10097 & n10098 ) | ( n10097 & n10193 ) | ( n10098 & n10193 ) ;
  assign n10195 = n10192 | n10194 ;
  assign n10196 = n10192 & n10194 ;
  assign n10197 = n10195 & ~n10196 ;
  assign n10198 = n10186 & n10197 ;
  assign n10199 = n10186 | n10197 ;
  assign n10200 = ~n10198 & n10199 ;
  assign n10201 = n10180 & n10200 ;
  assign n10202 = n10180 | n10200 ;
  assign n10203 = ~n10201 & n10202 ;
  assign n10204 = n10165 & n10203 ;
  assign n10205 = n10165 | n10203 ;
  assign n10206 = ~n10204 & n10205 ;
  assign n10207 = n10032 | n10038 ;
  assign n10208 = n10206 & n10207 ;
  assign n10209 = n10207 & ~n10208 ;
  assign n10210 = ( n10206 & ~n10208 ) | ( n10206 & n10209 ) | ( ~n10208 & n10209 ) ;
  assign n10211 = n9868 | n10041 ;
  assign n10212 = n9866 | n10041 ;
  assign n10213 = ( n9867 & n10211 ) | ( n9867 & n10212 ) | ( n10211 & n10212 ) ;
  assign n10214 = ( n9869 & n9872 ) | ( n9869 & n10213 ) | ( n9872 & n10213 ) ;
  assign n10215 = n10210 | n10214 ;
  assign n10216 = n10210 & n10214 ;
  assign n10217 = n10215 & ~n10216 ;
  assign n10218 = n9898 | n9964 ;
  assign n10219 = n9898 & n9964 ;
  assign n10220 = n10218 & ~n10219 ;
  assign n10221 = n9883 | n10220 ;
  assign n10222 = n9883 & n10220 ;
  assign n10223 = n10221 & ~n10222 ;
  assign n10224 = n9906 | n9924 ;
  assign n10225 = n10223 & n10224 ;
  assign n10226 = n9906 & n10223 ;
  assign n10227 = ( n9909 & n10225 ) | ( n9909 & n10226 ) | ( n10225 & n10226 ) ;
  assign n10228 = n10223 | n10224 ;
  assign n10229 = n9906 | n10223 ;
  assign n10230 = ( n9909 & n10228 ) | ( n9909 & n10229 ) | ( n10228 & n10229 ) ;
  assign n10231 = ~n10227 & n10230 ;
  assign n10232 = n10006 | n10022 ;
  assign n10233 = ( n10006 & n10009 ) | ( n10006 & n10232 ) | ( n10009 & n10232 ) ;
  assign n10234 = n10231 | n10233 ;
  assign n10235 = n10231 & n10233 ;
  assign n10236 = n10234 & ~n10235 ;
  assign n10237 = n9814 | n9819 ;
  assign n10238 = ( n9814 & n9817 ) | ( n9814 & n10237 ) | ( n9817 & n10237 ) ;
  assign n10239 = n9951 | n9971 ;
  assign n10240 = ( n9951 & n9954 ) | ( n9951 & n10239 ) | ( n9954 & n10239 ) ;
  assign n10241 = n10238 | n10240 ;
  assign n10242 = n10238 & n10240 ;
  assign n10243 = n10241 & ~n10242 ;
  assign n10244 = x0 & x63 ;
  assign n10245 = n10083 & n10244 ;
  assign n10246 = n10083 & ~n10245 ;
  assign n10247 = ~n10083 & n10244 ;
  assign n10248 = n10246 | n10247 ;
  assign n10249 = x1 & ~x62 ;
  assign n10250 = ( x1 & ~n2779 ) | ( x1 & n10249 ) | ( ~n2779 & n10249 ) ;
  assign n10251 = x62 & n10250 ;
  assign n10252 = x32 & ~x62 ;
  assign n10253 = ( x32 & ~n2779 ) | ( x32 & n10252 ) | ( ~n2779 & n10252 ) ;
  assign n10254 = n10251 | n10253 ;
  assign n10255 = ~n10248 & n10254 ;
  assign n10256 = n10248 & ~n10254 ;
  assign n10257 = n10255 | n10256 ;
  assign n10258 = n2340 & n5798 ;
  assign n10259 = n1912 & n5392 ;
  assign n10260 = n10258 | n10259 ;
  assign n10261 = n2511 & n4857 ;
  assign n10262 = x39 & n10261 ;
  assign n10263 = ( x39 & ~n10260 ) | ( x39 & n10262 ) | ( ~n10260 & n10262 ) ;
  assign n10264 = x24 & n10263 ;
  assign n10265 = n10260 | n10261 ;
  assign n10266 = x25 & x38 ;
  assign n10267 = x26 & x37 ;
  assign n10268 = ( ~n10261 & n10266 ) | ( ~n10261 & n10267 ) | ( n10266 & n10267 ) ;
  assign n10269 = n10266 & n10267 ;
  assign n10270 = ( ~n10260 & n10268 ) | ( ~n10260 & n10269 ) | ( n10268 & n10269 ) ;
  assign n10271 = ~n10265 & n10270 ;
  assign n10272 = n10264 | n10271 ;
  assign n10273 = n2075 & n4914 ;
  assign n10274 = n2372 & n4078 ;
  assign n10275 = n10273 | n10274 ;
  assign n10276 = n2369 & n3483 ;
  assign n10277 = x36 & n10276 ;
  assign n10278 = ( x36 & ~n10275 ) | ( x36 & n10277 ) | ( ~n10275 & n10277 ) ;
  assign n10279 = x27 & n10278 ;
  assign n10280 = n10275 | n10276 ;
  assign n10281 = x28 & x35 ;
  assign n10282 = ( n3878 & ~n10276 ) | ( n3878 & n10281 ) | ( ~n10276 & n10281 ) ;
  assign n10283 = n3878 & n10281 ;
  assign n10284 = ( ~n10275 & n10282 ) | ( ~n10275 & n10283 ) | ( n10282 & n10283 ) ;
  assign n10285 = ~n10280 & n10284 ;
  assign n10286 = n10279 | n10285 ;
  assign n10287 = n10272 & n10286 ;
  assign n10288 = n10272 & ~n10287 ;
  assign n10289 = n10286 & ~n10287 ;
  assign n10290 = n10288 | n10289 ;
  assign n10291 = n10257 & ~n10290 ;
  assign n10292 = ~n10257 & n10290 ;
  assign n10293 = n10291 | n10292 ;
  assign n10294 = ~n10243 & n10293 ;
  assign n10295 = n10236 & n10294 ;
  assign n10296 = n10243 & ~n10293 ;
  assign n10297 = ( n10236 & n10295 ) | ( n10236 & n10296 ) | ( n10295 & n10296 ) ;
  assign n10298 = n10236 | n10294 ;
  assign n10299 = n10296 | n10298 ;
  assign n10300 = ~n10297 & n10299 ;
  assign n10301 = n10050 | n10055 ;
  assign n10302 = ( n10050 & n10053 ) | ( n10050 & n10301 ) | ( n10053 & n10301 ) ;
  assign n10303 = n10300 & n10302 ;
  assign n10304 = n10300 | n10302 ;
  assign n10305 = ~n10303 & n10304 ;
  assign n10306 = n10058 & n10118 ;
  assign n10307 = n10305 & n10306 ;
  assign n10308 = ( n10121 & n10305 ) | ( n10121 & n10307 ) | ( n10305 & n10307 ) ;
  assign n10309 = n10305 | n10306 ;
  assign n10310 = n10121 | n10309 ;
  assign n10311 = ~n10308 & n10310 ;
  assign n10312 = n7551 & n9878 ;
  assign n10313 = n1020 & n5975 ;
  assign n10314 = n10312 | n10313 ;
  assign n10315 = x46 & x54 ;
  assign n10316 = n1694 & n10315 ;
  assign n10317 = x45 & n10316 ;
  assign n10318 = ( x45 & ~n10314 ) | ( x45 & n10317 ) | ( ~n10314 & n10317 ) ;
  assign n10319 = x18 & n10318 ;
  assign n10320 = n10314 | n10316 ;
  assign n10321 = x9 & x54 ;
  assign n10322 = x17 & x46 ;
  assign n10323 = ( ~n10316 & n10321 ) | ( ~n10316 & n10322 ) | ( n10321 & n10322 ) ;
  assign n10324 = n10321 & n10322 ;
  assign n10325 = ( ~n10314 & n10323 ) | ( ~n10314 & n10324 ) | ( n10323 & n10324 ) ;
  assign n10326 = ~n10320 & n10325 ;
  assign n10327 = n10319 | n10326 ;
  assign n10328 = n618 & n8161 ;
  assign n10329 = x16 & x53 ;
  assign n10330 = n8390 & n10329 ;
  assign n10331 = n10328 | n10330 ;
  assign n10332 = x47 & x52 ;
  assign n10333 = n1846 & n10332 ;
  assign n10334 = x53 & n10333 ;
  assign n10335 = ( x53 & ~n10331 ) | ( x53 & n10334 ) | ( ~n10331 & n10334 ) ;
  assign n10336 = x10 & n10335 ;
  assign n10337 = n10331 | n10333 ;
  assign n10338 = x11 & x52 ;
  assign n10339 = x16 & x47 ;
  assign n10340 = ( ~n10333 & n10338 ) | ( ~n10333 & n10339 ) | ( n10338 & n10339 ) ;
  assign n10341 = n10338 & n10339 ;
  assign n10342 = ( ~n10331 & n10340 ) | ( ~n10331 & n10341 ) | ( n10340 & n10341 ) ;
  assign n10343 = ~n10337 & n10342 ;
  assign n10344 = n10336 | n10343 ;
  assign n10345 = n10327 & n10344 ;
  assign n10346 = n10327 & ~n10345 ;
  assign n10347 = n10344 & ~n10345 ;
  assign n10348 = n10346 | n10347 ;
  assign n10349 = n723 & n6345 ;
  assign n10350 = x12 & x51 ;
  assign n10351 = n8074 & n10350 ;
  assign n10352 = n10349 | n10351 ;
  assign n10353 = n647 & n7112 ;
  assign n10354 = n8074 & n10353 ;
  assign n10355 = ( n8074 & ~n10352 ) | ( n8074 & n10354 ) | ( ~n10352 & n10354 ) ;
  assign n10356 = n10352 | n10353 ;
  assign n10357 = x13 & x50 ;
  assign n10358 = ( n10350 & ~n10353 ) | ( n10350 & n10357 ) | ( ~n10353 & n10357 ) ;
  assign n10359 = n10350 & n10357 ;
  assign n10360 = ( ~n10352 & n10358 ) | ( ~n10352 & n10359 ) | ( n10358 & n10359 ) ;
  assign n10361 = ~n10356 & n10360 ;
  assign n10362 = n10355 | n10361 ;
  assign n10363 = ~n10348 & n10362 ;
  assign n10364 = n10348 & ~n10362 ;
  assign n10365 = n10363 | n10364 ;
  assign n10366 = n119 & n9737 ;
  assign n10367 = x60 & x61 ;
  assign n10368 = n77 & n10367 ;
  assign n10369 = n10366 | n10368 ;
  assign n10370 = x59 & x60 ;
  assign n10371 = n79 & n10370 ;
  assign n10372 = x2 & n10371 ;
  assign n10373 = ( x2 & ~n10369 ) | ( x2 & n10372 ) | ( ~n10369 & n10372 ) ;
  assign n10374 = x61 & n10373 ;
  assign n10375 = n10369 | n10371 ;
  assign n10376 = x3 & x60 ;
  assign n10377 = x4 & x59 ;
  assign n10378 = ( ~n10371 & n10376 ) | ( ~n10371 & n10377 ) | ( n10376 & n10377 ) ;
  assign n10379 = n10376 & n10377 ;
  assign n10380 = ( ~n10369 & n10378 ) | ( ~n10369 & n10379 ) | ( n10378 & n10379 ) ;
  assign n10381 = ~n10375 & n10380 ;
  assign n10382 = ~n9983 & n10381 ;
  assign n10383 = ( ~n9983 & n10374 ) | ( ~n9983 & n10382 ) | ( n10374 & n10382 ) ;
  assign n10384 = n9983 & ~n10381 ;
  assign n10385 = ~n10374 & n10384 ;
  assign n10386 = n10383 | n10385 ;
  assign n10387 = x21 & x42 ;
  assign n10388 = x22 & x41 ;
  assign n10389 = n10387 | n10388 ;
  assign n10390 = n1585 & n5710 ;
  assign n10391 = x5 & x58 ;
  assign n10392 = ~n10390 & n10391 ;
  assign n10393 = n10389 | n10390 ;
  assign n10394 = ( n10390 & n10392 ) | ( n10390 & n10393 ) | ( n10392 & n10393 ) ;
  assign n10395 = n10389 & ~n10394 ;
  assign n10396 = ( ~n10389 & n10390 ) | ( ~n10389 & n10391 ) | ( n10390 & n10391 ) ;
  assign n10397 = n10391 & n10396 ;
  assign n10398 = n10395 | n10397 ;
  assign n10399 = n10386 & n10398 ;
  assign n10400 = n10386 | n10398 ;
  assign n10401 = ~n10399 & n10400 ;
  assign n10402 = x6 & x57 ;
  assign n10403 = x20 & x43 ;
  assign n10404 = n10402 | n10403 ;
  assign n10405 = x23 & x40 ;
  assign n10406 = ( n10402 & n10403 ) | ( n10402 & n10405 ) | ( n10403 & n10405 ) ;
  assign n10407 = n10404 & ~n10406 ;
  assign n10408 = n10402 & n10403 ;
  assign n10409 = n10405 & ~n10408 ;
  assign n10410 = ~n10404 & n10405 ;
  assign n10411 = ( n10405 & ~n10409 ) | ( n10405 & n10410 ) | ( ~n10409 & n10410 ) ;
  assign n10412 = n10407 | n10411 ;
  assign n10413 = x30 & x33 ;
  assign n10414 = n4062 | n10413 ;
  assign n10415 = x14 & x49 ;
  assign n10416 = ( n4062 & n10413 ) | ( n4062 & n10415 ) | ( n10413 & n10415 ) ;
  assign n10417 = n10414 & ~n10416 ;
  assign n10418 = n4062 & n10413 ;
  assign n10419 = n10415 & ~n10418 ;
  assign n10420 = ~n10414 & n10415 ;
  assign n10421 = ( n10415 & ~n10419 ) | ( n10415 & n10420 ) | ( ~n10419 & n10420 ) ;
  assign n10422 = n10417 | n10421 ;
  assign n10423 = n10412 & n10422 ;
  assign n10424 = n10412 & ~n10423 ;
  assign n10425 = n10422 & ~n10423 ;
  assign n10426 = n10424 | n10425 ;
  assign n10427 = n251 & n10013 ;
  assign n10428 = x44 & x56 ;
  assign n10429 = n1682 & n10428 ;
  assign n10430 = n10427 | n10429 ;
  assign n10431 = x44 & x55 ;
  assign n10432 = n1859 & n10431 ;
  assign n10433 = x56 & n10432 ;
  assign n10434 = ( x56 & ~n10430 ) | ( x56 & n10433 ) | ( ~n10430 & n10433 ) ;
  assign n10435 = x7 & n10434 ;
  assign n10436 = n10430 | n10432 ;
  assign n10437 = x8 & x55 ;
  assign n10438 = x19 & x44 ;
  assign n10439 = ( ~n10432 & n10437 ) | ( ~n10432 & n10438 ) | ( n10437 & n10438 ) ;
  assign n10440 = n10437 & n10438 ;
  assign n10441 = ( ~n10430 & n10439 ) | ( ~n10430 & n10440 ) | ( n10439 & n10440 ) ;
  assign n10442 = ~n10436 & n10441 ;
  assign n10443 = n10435 | n10442 ;
  assign n10444 = ( n10401 & n10426 ) | ( n10401 & ~n10443 ) | ( n10426 & ~n10443 ) ;
  assign n10445 = ( n10401 & ~n10426 ) | ( n10401 & n10443 ) | ( ~n10426 & n10443 ) ;
  assign n10446 = ( ~n10401 & n10444 ) | ( ~n10401 & n10445 ) | ( n10444 & n10445 ) ;
  assign n10447 = n10365 & n10446 ;
  assign n10448 = n10365 | n10446 ;
  assign n10449 = ~n10447 & n10448 ;
  assign n10450 = n9862 & n10449 ;
  assign n10451 = ( n9861 & n10449 ) | ( n9861 & n10450 ) | ( n10449 & n10450 ) ;
  assign n10452 = n9825 | n9862 ;
  assign n10453 = ( ~n9825 & n9860 ) | ( ~n9825 & n10452 ) | ( n9860 & n10452 ) ;
  assign n10454 = ~n10451 & n10453 ;
  assign n10455 = n10109 | n10115 ;
  assign n10456 = n10449 & ~n10450 ;
  assign n10457 = ~n9861 & n10456 ;
  assign n10458 = n10455 & n10457 ;
  assign n10459 = ( n10454 & n10455 ) | ( n10454 & n10458 ) | ( n10455 & n10458 ) ;
  assign n10460 = n10455 | n10457 ;
  assign n10461 = n10454 | n10460 ;
  assign n10462 = ~n10459 & n10461 ;
  assign n10463 = n10311 & ~n10462 ;
  assign n10464 = n10311 | n10462 ;
  assign n10465 = ( ~n10311 & n10463 ) | ( ~n10311 & n10464 ) | ( n10463 & n10464 ) ;
  assign n10466 = n10217 | n10465 ;
  assign n10467 = n10217 & n10465 ;
  assign n10468 = n10466 & ~n10467 ;
  assign n10469 = n10044 | n10126 ;
  assign n10470 = ( n10126 & n10129 ) | ( n10126 & n10469 ) | ( n10129 & n10469 ) ;
  assign n10471 = ( n10151 & n10468 ) | ( n10151 & ~n10470 ) | ( n10468 & ~n10470 ) ;
  assign n10472 = ( ~n10468 & n10470 ) | ( ~n10468 & n10471 ) | ( n10470 & n10471 ) ;
  assign n10473 = ( ~n10151 & n10471 ) | ( ~n10151 & n10472 ) | ( n10471 & n10472 ) ;
  assign n10520 = n10307 | n10462 ;
  assign n10521 = n10305 | n10462 ;
  assign n10522 = ( n10121 & n10520 ) | ( n10121 & n10521 ) | ( n10520 & n10521 ) ;
  assign n10523 = ( n10308 & n10311 ) | ( n10308 & n10522 ) | ( n10311 & n10522 ) ;
  assign n10474 = n10426 & n10443 ;
  assign n10475 = n10426 & ~n10474 ;
  assign n10476 = ~n10426 & n10443 ;
  assign n10477 = n10401 & n10476 ;
  assign n10478 = ( n10401 & n10475 ) | ( n10401 & n10477 ) | ( n10475 & n10477 ) ;
  assign n10479 = n10447 | n10478 ;
  assign n10480 = n10242 | n10293 ;
  assign n10481 = ( n10242 & n10243 ) | ( n10242 & n10480 ) | ( n10243 & n10480 ) ;
  assign n10482 = n10479 | n10481 ;
  assign n10483 = n10479 & n10481 ;
  assign n10484 = n10482 & ~n10483 ;
  assign n10485 = n10316 | n10406 ;
  assign n10486 = n10314 | n10485 ;
  assign n10487 = n10316 & n10406 ;
  assign n10488 = ( n10314 & n10406 ) | ( n10314 & n10487 ) | ( n10406 & n10487 ) ;
  assign n10489 = n10486 & ~n10488 ;
  assign n10490 = n10280 | n10489 ;
  assign n10491 = n10280 & n10489 ;
  assign n10492 = n10490 & ~n10491 ;
  assign n10493 = n10375 | n10394 ;
  assign n10494 = n10375 & n10394 ;
  assign n10495 = n10493 & ~n10494 ;
  assign n10496 = n10436 | n10495 ;
  assign n10497 = n10436 & n10495 ;
  assign n10498 = n10496 & ~n10497 ;
  assign n10499 = n10492 | n10498 ;
  assign n10500 = n10492 & n10498 ;
  assign n10501 = n10499 & ~n10500 ;
  assign n10502 = ( n10257 & n10272 ) | ( n10257 & n10286 ) | ( n10272 & n10286 ) ;
  assign n10503 = n10501 & n10502 ;
  assign n10504 = n10501 | n10502 ;
  assign n10505 = ~n10503 & n10504 ;
  assign n10506 = n10484 | n10505 ;
  assign n10507 = n10484 & n10505 ;
  assign n10508 = n10506 & ~n10507 ;
  assign n10509 = n10297 | n10302 ;
  assign n10510 = ( n10297 & n10300 ) | ( n10297 & n10509 ) | ( n10300 & n10509 ) ;
  assign n10511 = n10508 & n10510 ;
  assign n10512 = n10508 & ~n10511 ;
  assign n10513 = ~n10508 & n10510 ;
  assign n10514 = n10512 | n10513 ;
  assign n10515 = n10451 | n10459 ;
  assign n10516 = n10514 & n10515 ;
  assign n10517 = n10514 & ~n10516 ;
  assign n10518 = ~n10514 & n10515 ;
  assign n10519 = n10517 | n10518 ;
  assign n10524 = n10519 & n10523 ;
  assign n10525 = n10523 & ~n10524 ;
  assign n10526 = n10265 | n10356 ;
  assign n10527 = n10265 & n10356 ;
  assign n10528 = n10526 & ~n10527 ;
  assign n10529 = n10337 | n10528 ;
  assign n10530 = n10337 & n10528 ;
  assign n10531 = n10529 & ~n10530 ;
  assign n10532 = n10423 | n10443 ;
  assign n10533 = ( n10423 & n10426 ) | ( n10423 & n10532 ) | ( n10426 & n10532 ) ;
  assign n10534 = n10531 & n10533 ;
  assign n10535 = n10531 | n10533 ;
  assign n10536 = ~n10534 & n10535 ;
  assign n10537 = n10345 | n10362 ;
  assign n10538 = ( n10345 & n10348 ) | ( n10345 & n10537 ) | ( n10348 & n10537 ) ;
  assign n10539 = n10536 | n10538 ;
  assign n10540 = n10536 & n10538 ;
  assign n10541 = n10539 & ~n10540 ;
  assign n10542 = n10159 | n10162 ;
  assign n10543 = ( n10159 & n10160 ) | ( n10159 & n10542 ) | ( n10160 & n10542 ) ;
  assign n10544 = n10541 | n10543 ;
  assign n10545 = n10541 & n10543 ;
  assign n10546 = n10544 & ~n10545 ;
  assign n10547 = n10374 | n10381 ;
  assign n10548 = ( n9983 & n10398 ) | ( n9983 & n10547 ) | ( n10398 & n10547 ) ;
  assign n10549 = n10168 | n10173 ;
  assign n10550 = ( n10166 & n10173 ) | ( n10166 & n10549 ) | ( n10173 & n10549 ) ;
  assign n10551 = n10548 & n10550 ;
  assign n10552 = n10168 & n10548 ;
  assign n10553 = n10166 & n10552 ;
  assign n10554 = ( n10171 & n10551 ) | ( n10171 & n10553 ) | ( n10551 & n10553 ) ;
  assign n10555 = n10548 | n10550 ;
  assign n10556 = n10168 | n10548 ;
  assign n10557 = ( n10166 & n10548 ) | ( n10166 & n10556 ) | ( n10548 & n10556 ) ;
  assign n10558 = ( n10171 & n10555 ) | ( n10171 & n10557 ) | ( n10555 & n10557 ) ;
  assign n10559 = ~n10554 & n10558 ;
  assign n10560 = x62 & n2779 ;
  assign n10561 = x62 & x63 ;
  assign n10562 = n2779 & n10561 ;
  assign n10563 = n10560 & ~n10562 ;
  assign n10564 = x63 & n10250 ;
  assign n10565 = n10563 | n10564 ;
  assign n10566 = n10416 & n10565 ;
  assign n10567 = n10565 & ~n10566 ;
  assign n10568 = n10416 & ~n10565 ;
  assign n10569 = n10567 | n10568 ;
  assign n10570 = x10 & x54 ;
  assign n10571 = x15 & x49 ;
  assign n10572 = n10570 & n10571 ;
  assign n10573 = x49 & x55 ;
  assign n10574 = n1462 & n10573 ;
  assign n10575 = n360 & n8357 ;
  assign n10576 = n10574 | n10575 ;
  assign n10577 = x55 & n10572 ;
  assign n10578 = ( x55 & ~n10576 ) | ( x55 & n10577 ) | ( ~n10576 & n10577 ) ;
  assign n10579 = x9 & n10578 ;
  assign n10580 = ( n10570 & n10571 ) | ( n10570 & ~n10576 ) | ( n10571 & ~n10576 ) ;
  assign n10581 = ( ~n10572 & n10579 ) | ( ~n10572 & n10580 ) | ( n10579 & n10580 ) ;
  assign n10582 = n720 & n7874 ;
  assign n10583 = n647 & n7567 ;
  assign n10584 = n10582 | n10583 ;
  assign n10585 = n490 & n8161 ;
  assign n10586 = x51 & n10585 ;
  assign n10587 = ( x51 & ~n10584 ) | ( x51 & n10586 ) | ( ~n10584 & n10586 ) ;
  assign n10588 = x13 & n10587 ;
  assign n10589 = n10584 | n10585 ;
  assign n10590 = x11 & x53 ;
  assign n10591 = x12 & x52 ;
  assign n10592 = ( ~n10585 & n10590 ) | ( ~n10585 & n10591 ) | ( n10590 & n10591 ) ;
  assign n10593 = n10590 & n10591 ;
  assign n10594 = ( ~n10584 & n10592 ) | ( ~n10584 & n10593 ) | ( n10592 & n10593 ) ;
  assign n10595 = ~n10589 & n10594 ;
  assign n10596 = n10588 | n10595 ;
  assign n10597 = n10581 & n10596 ;
  assign n10598 = n10581 & ~n10597 ;
  assign n10599 = n10596 & ~n10597 ;
  assign n10600 = n10598 | n10599 ;
  assign n10601 = n10569 & ~n10600 ;
  assign n10602 = ~n10569 & n10600 ;
  assign n10603 = n10601 | n10602 ;
  assign n10604 = ~n10559 & n10603 ;
  assign n10605 = n10559 & ~n10603 ;
  assign n10606 = n10604 | n10605 ;
  assign n10607 = n10546 | n10606 ;
  assign n10608 = n10546 & n10606 ;
  assign n10609 = n10607 & ~n10608 ;
  assign n10610 = n10204 & n10609 ;
  assign n10611 = ( n10208 & n10609 ) | ( n10208 & n10610 ) | ( n10609 & n10610 ) ;
  assign n10612 = n10204 | n10609 ;
  assign n10613 = n10208 | n10612 ;
  assign n10614 = ~n10611 & n10613 ;
  assign n10615 = n200 & n9272 ;
  assign n10616 = x17 & x58 ;
  assign n10617 = n7159 & n10616 ;
  assign n10618 = n10615 | n10617 ;
  assign n10619 = x17 & x57 ;
  assign n10620 = n7583 & n10619 ;
  assign n10621 = x58 & n10620 ;
  assign n10622 = ( x58 & ~n10618 ) | ( x58 & n10621 ) | ( ~n10618 & n10621 ) ;
  assign n10623 = x6 & n10622 ;
  assign n10624 = n10618 | n10620 ;
  assign n10625 = x7 & x57 ;
  assign n10626 = ( n6354 & ~n10620 ) | ( n6354 & n10625 ) | ( ~n10620 & n10625 ) ;
  assign n10627 = n6354 & n10625 ;
  assign n10628 = ( ~n10618 & n10626 ) | ( ~n10618 & n10627 ) | ( n10626 & n10627 ) ;
  assign n10629 = ~n10624 & n10628 ;
  assign n10630 = n10623 | n10629 ;
  assign n10631 = n1710 & n4969 ;
  assign n10632 = n1434 & n5658 ;
  assign n10633 = n10631 | n10632 ;
  assign n10634 = n1585 & n5407 ;
  assign n10635 = x44 & n10634 ;
  assign n10636 = ( x44 & ~n10633 ) | ( x44 & n10635 ) | ( ~n10633 & n10635 ) ;
  assign n10637 = x20 & n10636 ;
  assign n10638 = n10633 | n10634 ;
  assign n10639 = x21 & x43 ;
  assign n10640 = x22 & x42 ;
  assign n10641 = ( ~n10634 & n10639 ) | ( ~n10634 & n10640 ) | ( n10639 & n10640 ) ;
  assign n10642 = n10639 & n10640 ;
  assign n10643 = ( ~n10633 & n10641 ) | ( ~n10633 & n10642 ) | ( n10641 & n10642 ) ;
  assign n10644 = ~n10638 & n10643 ;
  assign n10645 = n10637 | n10644 ;
  assign n10646 = n10630 & n10645 ;
  assign n10647 = n10630 & ~n10646 ;
  assign n10648 = n10645 & ~n10646 ;
  assign n10649 = n10647 | n10648 ;
  assign n10650 = n1557 & n4350 ;
  assign n10651 = n1686 & n5813 ;
  assign n10652 = n10650 | n10651 ;
  assign n10653 = n1912 & n4555 ;
  assign n10654 = x41 & n10653 ;
  assign n10655 = ( x41 & ~n10652 ) | ( x41 & n10654 ) | ( ~n10652 & n10654 ) ;
  assign n10656 = x23 & n10655 ;
  assign n10657 = n10652 | n10653 ;
  assign n10658 = x24 & x40 ;
  assign n10659 = x25 & x39 ;
  assign n10660 = ( ~n10653 & n10658 ) | ( ~n10653 & n10659 ) | ( n10658 & n10659 ) ;
  assign n10661 = n10658 & n10659 ;
  assign n10662 = ( ~n10652 & n10660 ) | ( ~n10652 & n10661 ) | ( n10660 & n10661 ) ;
  assign n10663 = ~n10657 & n10662 ;
  assign n10664 = n10656 | n10663 ;
  assign n10665 = ~n10649 & n10664 ;
  assign n10666 = n10649 & ~n10664 ;
  assign n10667 = n10665 | n10666 ;
  assign n10668 = x18 & x46 ;
  assign n10669 = x19 & x45 ;
  assign n10670 = n10668 | n10669 ;
  assign n10671 = n1077 & n5975 ;
  assign n10672 = n10670 & ~n10671 ;
  assign n10673 = n9742 | n10671 ;
  assign n10674 = ( n10671 & n10672 ) | ( n10671 & n10673 ) | ( n10672 & n10673 ) ;
  assign n10675 = n10670 & ~n10674 ;
  assign n10676 = n9742 & ~n10672 ;
  assign n10677 = n10675 | n10676 ;
  assign n10678 = n10245 | n10254 ;
  assign n10679 = ( n10245 & n10248 ) | ( n10245 & n10678 ) | ( n10248 & n10678 ) ;
  assign n10680 = n10677 & ~n10679 ;
  assign n10681 = ~n10677 & n10679 ;
  assign n10682 = n10680 | n10681 ;
  assign n10683 = n119 & n9931 ;
  assign n10684 = x61 & x62 ;
  assign n10685 = n77 & n10684 ;
  assign n10686 = n10683 | n10685 ;
  assign n10687 = n79 & n10367 ;
  assign n10688 = x62 & n10687 ;
  assign n10689 = ( x62 & ~n10686 ) | ( x62 & n10688 ) | ( ~n10686 & n10688 ) ;
  assign n10690 = x2 & n10689 ;
  assign n10691 = n10686 | n10687 ;
  assign n10692 = x3 & x61 ;
  assign n10693 = x4 & x60 ;
  assign n10694 = ( ~n10687 & n10692 ) | ( ~n10687 & n10693 ) | ( n10692 & n10693 ) ;
  assign n10695 = n10692 & n10693 ;
  assign n10696 = ( ~n10686 & n10694 ) | ( ~n10686 & n10695 ) | ( n10694 & n10695 ) ;
  assign n10697 = ~n10691 & n10696 ;
  assign n10698 = n10690 | n10697 ;
  assign n10699 = n10682 & n10698 ;
  assign n10700 = n10682 | n10698 ;
  assign n10701 = ~n10699 & n10700 ;
  assign n10702 = n2075 & n5417 ;
  assign n10703 = n2372 & n3770 ;
  assign n10704 = n10702 | n10703 ;
  assign n10705 = n2369 & n4078 ;
  assign n10706 = n4286 & n10705 ;
  assign n10707 = ( n4286 & ~n10704 ) | ( n4286 & n10706 ) | ( ~n10704 & n10706 ) ;
  assign n10708 = n10704 | n10705 ;
  assign n10709 = x28 & x36 ;
  assign n10710 = x29 & x35 ;
  assign n10711 = ( ~n10705 & n10709 ) | ( ~n10705 & n10710 ) | ( n10709 & n10710 ) ;
  assign n10712 = n10709 & n10710 ;
  assign n10713 = ( ~n10704 & n10711 ) | ( ~n10704 & n10712 ) | ( n10711 & n10712 ) ;
  assign n10714 = ~n10708 & n10713 ;
  assign n10715 = n10707 | n10714 ;
  assign n10716 = x8 & x56 ;
  assign n10717 = n7189 | n10716 ;
  assign n10718 = x48 & x56 ;
  assign n10719 = n1454 & n10718 ;
  assign n10720 = n10717 | n10719 ;
  assign n10721 = x26 & x38 ;
  assign n10722 = ( ~n10719 & n10720 ) | ( ~n10719 & n10721 ) | ( n10720 & n10721 ) ;
  assign n10723 = ( n10719 & n10720 ) | ( n10719 & ~n10721 ) | ( n10720 & ~n10721 ) ;
  assign n10724 = ( ~n10720 & n10722 ) | ( ~n10720 & n10723 ) | ( n10722 & n10723 ) ;
  assign n10725 = n10715 & ~n10724 ;
  assign n10726 = ~n10715 & n10724 ;
  assign n10727 = n10725 | n10726 ;
  assign n10728 = x30 & x34 ;
  assign n10729 = n2683 | n10728 ;
  assign n10730 = n2965 & n4530 ;
  assign n10731 = n9683 & ~n10730 ;
  assign n10732 = n10729 | n10730 ;
  assign n10733 = ( n10730 & n10731 ) | ( n10730 & n10732 ) | ( n10731 & n10732 ) ;
  assign n10734 = n10729 & ~n10733 ;
  assign n10735 = n9683 & ~n10729 ;
  assign n10736 = ( n9683 & ~n10731 ) | ( n9683 & n10735 ) | ( ~n10731 & n10735 ) ;
  assign n10737 = n10734 | n10736 ;
  assign n10738 = n10727 & n10737 ;
  assign n10739 = n10727 | n10737 ;
  assign n10740 = ~n10738 & n10739 ;
  assign n10741 = n10701 & ~n10740 ;
  assign n10742 = ~n10701 & n10740 ;
  assign n10743 = n10741 | n10742 ;
  assign n10744 = n10667 & n10743 ;
  assign n10745 = n10667 | n10743 ;
  assign n10746 = ~n10744 & n10745 ;
  assign n10747 = n10179 | n10200 ;
  assign n10748 = ( n10179 & n10180 ) | ( n10179 & n10747 ) | ( n10180 & n10747 ) ;
  assign n10749 = n10746 & n10748 ;
  assign n10750 = n10746 | n10748 ;
  assign n10751 = ~n10749 & n10750 ;
  assign n10764 = n10186 | n10196 ;
  assign n10765 = ( n10196 & n10197 ) | ( n10196 & n10764 ) | ( n10197 & n10764 ) ;
  assign n10752 = n9998 | n10182 ;
  assign n10753 = ( n10182 & n10183 ) | ( n10182 & n10752 ) | ( n10183 & n10752 ) ;
  assign n10754 = n9883 | n10219 ;
  assign n10755 = ( n10219 & n10220 ) | ( n10219 & n10754 ) | ( n10220 & n10754 ) ;
  assign n10756 = n10753 | n10755 ;
  assign n10757 = n10753 & n10755 ;
  assign n10758 = n10756 & ~n10757 ;
  assign n10759 = n9935 | n10188 ;
  assign n10760 = ( n10188 & n10189 ) | ( n10188 & n10759 ) | ( n10189 & n10759 ) ;
  assign n10761 = n10758 | n10760 ;
  assign n10762 = n10758 & n10760 ;
  assign n10763 = n10761 & ~n10762 ;
  assign n10766 = n10227 | n10233 ;
  assign n10767 = ( n10227 & n10231 ) | ( n10227 & n10766 ) | ( n10231 & n10766 ) ;
  assign n10768 = ( n10763 & n10765 ) | ( n10763 & ~n10767 ) | ( n10765 & ~n10767 ) ;
  assign n10769 = ( ~n10763 & n10767 ) | ( ~n10763 & n10768 ) | ( n10767 & n10768 ) ;
  assign n10770 = ( ~n10765 & n10768 ) | ( ~n10765 & n10769 ) | ( n10768 & n10769 ) ;
  assign n10771 = n10751 & ~n10770 ;
  assign n10772 = n10751 | n10770 ;
  assign n10773 = ( ~n10751 & n10771 ) | ( ~n10751 & n10772 ) | ( n10771 & n10772 ) ;
  assign n10774 = n10614 & n10773 ;
  assign n10775 = n10614 | n10773 ;
  assign n10776 = ~n10774 & n10775 ;
  assign n10777 = n10519 & ~n10523 ;
  assign n10778 = n10776 & n10777 ;
  assign n10779 = ( n10525 & n10776 ) | ( n10525 & n10778 ) | ( n10776 & n10778 ) ;
  assign n10780 = n10776 | n10777 ;
  assign n10781 = n10525 | n10780 ;
  assign n10782 = ~n10779 & n10781 ;
  assign n10783 = n10216 | n10467 ;
  assign n10784 = n10782 | n10783 ;
  assign n10785 = n10782 & n10783 ;
  assign n10786 = n10784 | n10785 ;
  assign n10787 = n10468 & n10470 ;
  assign n10788 = n10468 | n10470 ;
  assign n10789 = n10135 & n10788 ;
  assign n10790 = ( n10146 & n10788 ) | ( n10146 & n10789 ) | ( n10788 & n10789 ) ;
  assign n10791 = ( n10147 & n10788 ) | ( n10147 & n10789 ) | ( n10788 & n10789 ) ;
  assign n10792 = ( n9167 & n10790 ) | ( n9167 & n10791 ) | ( n10790 & n10791 ) ;
  assign n10793 = ( n9166 & n10790 ) | ( n9166 & n10791 ) | ( n10790 & n10791 ) ;
  assign n10794 = ( n8252 & n10792 ) | ( n8252 & n10793 ) | ( n10792 & n10793 ) ;
  assign n10795 = n10787 | n10794 ;
  assign n10796 = ( n10785 & ~n10786 ) | ( n10785 & n10795 ) | ( ~n10786 & n10795 ) ;
  assign n10797 = ( n10785 & n10786 ) | ( n10785 & n10795 ) | ( n10786 & n10795 ) ;
  assign n10798 = ( n10786 & n10796 ) | ( n10786 & ~n10797 ) | ( n10796 & ~n10797 ) ;
  assign n10799 = n10784 & n10787 ;
  assign n10800 = ( n10784 & n10794 ) | ( n10784 & n10799 ) | ( n10794 & n10799 ) ;
  assign n10801 = n10785 | n10800 ;
  assign n10802 = n10524 | n10779 ;
  assign n10803 = ( n10667 & n10701 ) | ( n10667 & n10740 ) | ( n10701 & n10740 ) ;
  assign n10804 = n10554 | n10603 ;
  assign n10805 = ( n10554 & n10559 ) | ( n10554 & n10804 ) | ( n10559 & n10804 ) ;
  assign n10806 = n10803 | n10805 ;
  assign n10807 = n10803 & n10805 ;
  assign n10808 = n10806 & ~n10807 ;
  assign n10809 = n10572 | n10576 ;
  assign n10810 = n10657 | n10809 ;
  assign n10811 = n10657 & n10809 ;
  assign n10812 = n10810 & ~n10811 ;
  assign n10813 = n10624 | n10812 ;
  assign n10814 = n10624 & n10812 ;
  assign n10815 = n10813 & ~n10814 ;
  assign n10816 = ~n10719 & n10721 ;
  assign n10817 = ( n10719 & n10720 ) | ( n10719 & n10816 ) | ( n10720 & n10816 ) ;
  assign n10818 = n10674 | n10691 ;
  assign n10819 = n10674 & n10691 ;
  assign n10820 = n10818 & ~n10819 ;
  assign n10821 = n10817 | n10820 ;
  assign n10822 = n10817 & n10820 ;
  assign n10823 = n10821 & ~n10822 ;
  assign n10824 = n10815 | n10823 ;
  assign n10825 = n10815 & n10823 ;
  assign n10826 = n10824 & ~n10825 ;
  assign n10827 = ( n10569 & n10581 ) | ( n10569 & n10596 ) | ( n10581 & n10596 ) ;
  assign n10828 = n10826 & n10827 ;
  assign n10829 = n10826 | n10827 ;
  assign n10830 = ~n10828 & n10829 ;
  assign n10831 = n10808 | n10830 ;
  assign n10832 = n10808 & n10830 ;
  assign n10833 = n10831 & ~n10832 ;
  assign n10834 = n10541 | n10606 ;
  assign n10835 = ( n10543 & n10606 ) | ( n10543 & n10834 ) | ( n10606 & n10834 ) ;
  assign n10836 = ( n10545 & n10546 ) | ( n10545 & n10835 ) | ( n10546 & n10835 ) ;
  assign n10837 = n10833 & n10836 ;
  assign n10838 = n10833 | n10836 ;
  assign n10839 = ~n10837 & n10838 ;
  assign n10840 = n10749 | n10770 ;
  assign n10841 = ( n10749 & n10751 ) | ( n10749 & n10840 ) | ( n10751 & n10840 ) ;
  assign n10842 = n10839 & n10841 ;
  assign n10843 = n10839 | n10841 ;
  assign n10844 = ~n10842 & n10843 ;
  assign n10845 = n10611 | n10773 ;
  assign n10846 = ( n10611 & n10614 ) | ( n10611 & n10845 ) | ( n10614 & n10845 ) ;
  assign n10847 = n10844 | n10846 ;
  assign n10848 = n10844 & n10846 ;
  assign n10849 = n10847 & ~n10848 ;
  assign n10850 = ( n10677 & n10679 ) | ( n10677 & n10698 ) | ( n10679 & n10698 ) ;
  assign n10851 = n10757 | n10760 ;
  assign n10852 = ( n10757 & n10758 ) | ( n10757 & n10851 ) | ( n10758 & n10851 ) ;
  assign n10853 = n10850 | n10852 ;
  assign n10854 = n10850 & n10852 ;
  assign n10855 = n10853 & ~n10854 ;
  assign n10856 = x61 & x63 ;
  assign n10857 = n119 & n10856 ;
  assign n10858 = x4 & x61 ;
  assign n10859 = x2 & x63 ;
  assign n10860 = n10858 | n10859 ;
  assign n10861 = ~n10857 & n10860 ;
  assign n10862 = n10733 & n10861 ;
  assign n10863 = n10733 & ~n10862 ;
  assign n10864 = ~n10733 & n10861 ;
  assign n10865 = n10863 | n10864 ;
  assign n10866 = x49 & x51 ;
  assign n10867 = n790 & n10866 ;
  assign n10868 = n795 & n6834 ;
  assign n10869 = n10867 | n10868 ;
  assign n10870 = n792 & n7112 ;
  assign n10871 = n8476 & n10870 ;
  assign n10872 = ( n8476 & ~n10869 ) | ( n8476 & n10871 ) | ( ~n10869 & n10871 ) ;
  assign n10873 = n10869 | n10870 ;
  assign n10874 = x14 & x51 ;
  assign n10875 = x15 & x50 ;
  assign n10876 = ( ~n10870 & n10874 ) | ( ~n10870 & n10875 ) | ( n10874 & n10875 ) ;
  assign n10877 = n10874 & n10875 ;
  assign n10878 = ( ~n10869 & n10876 ) | ( ~n10869 & n10877 ) | ( n10876 & n10877 ) ;
  assign n10879 = ~n10873 & n10878 ;
  assign n10880 = n10872 | n10879 ;
  assign n10881 = x13 & x52 ;
  assign n10882 = x18 & x47 ;
  assign n10883 = n10881 & n10882 ;
  assign n10884 = n647 & n8161 ;
  assign n10885 = n8933 & n9413 ;
  assign n10886 = n10884 | n10885 ;
  assign n10887 = x53 & n10883 ;
  assign n10888 = ( x53 & ~n10886 ) | ( x53 & n10887 ) | ( ~n10886 & n10887 ) ;
  assign n10889 = x12 & n10888 ;
  assign n10890 = ( n10881 & n10882 ) | ( n10881 & ~n10886 ) | ( n10882 & ~n10886 ) ;
  assign n10891 = ( ~n10883 & n10889 ) | ( ~n10883 & n10890 ) | ( n10889 & n10890 ) ;
  assign n10892 = ( n10865 & ~n10880 ) | ( n10865 & n10891 ) | ( ~n10880 & n10891 ) ;
  assign n10893 = ( n10865 & n10880 ) | ( n10865 & ~n10891 ) | ( n10880 & ~n10891 ) ;
  assign n10894 = ( ~n10865 & n10892 ) | ( ~n10865 & n10893 ) | ( n10892 & n10893 ) ;
  assign n10895 = ~n10855 & n10894 ;
  assign n10896 = n10850 | n10894 ;
  assign n10897 = ( n10852 & n10894 ) | ( n10852 & n10896 ) | ( n10894 & n10896 ) ;
  assign n10898 = n10853 & ~n10897 ;
  assign n10899 = n10895 | n10898 ;
  assign n10900 = n10765 & n10767 ;
  assign n10901 = n10767 & ~n10900 ;
  assign n10902 = n10763 & n10765 ;
  assign n10903 = ~n10767 & n10902 ;
  assign n10904 = ( n10763 & n10901 ) | ( n10763 & n10903 ) | ( n10901 & n10903 ) ;
  assign n10905 = n10638 | n10708 ;
  assign n10906 = n10638 & n10708 ;
  assign n10907 = n10905 & ~n10906 ;
  assign n10908 = n10589 | n10907 ;
  assign n10909 = n10589 & n10907 ;
  assign n10910 = n10908 & ~n10909 ;
  assign n10911 = n10715 & n10724 ;
  assign n10912 = n10910 & n10911 ;
  assign n10913 = ( n10738 & n10910 ) | ( n10738 & n10912 ) | ( n10910 & n10912 ) ;
  assign n10914 = n10910 | n10911 ;
  assign n10915 = n10738 | n10914 ;
  assign n10916 = ~n10913 & n10915 ;
  assign n10917 = n10646 | n10664 ;
  assign n10918 = ( n10646 & n10649 ) | ( n10646 & n10917 ) | ( n10649 & n10917 ) ;
  assign n10919 = n10916 | n10918 ;
  assign n10920 = n10916 & n10918 ;
  assign n10921 = n10919 & ~n10920 ;
  assign n10922 = n10900 & n10921 ;
  assign n10923 = ( n10904 & n10921 ) | ( n10904 & n10922 ) | ( n10921 & n10922 ) ;
  assign n10924 = n10900 | n10903 ;
  assign n10925 = n10763 | n10765 ;
  assign n10926 = ( n10763 & n10767 ) | ( n10763 & n10925 ) | ( n10767 & n10925 ) ;
  assign n10927 = ( n10901 & n10924 ) | ( n10901 & n10926 ) | ( n10924 & n10926 ) ;
  assign n10928 = ~n10923 & n10927 ;
  assign n10929 = n10921 & ~n10922 ;
  assign n10930 = ~n10904 & n10929 ;
  assign n10931 = n10899 & n10930 ;
  assign n10932 = ( n10899 & n10928 ) | ( n10899 & n10931 ) | ( n10928 & n10931 ) ;
  assign n10933 = n10899 | n10930 ;
  assign n10934 = n10928 | n10933 ;
  assign n10935 = ~n10932 & n10934 ;
  assign n10936 = n10337 | n10527 ;
  assign n10937 = ( n10527 & n10528 ) | ( n10527 & n10936 ) | ( n10528 & n10936 ) ;
  assign n10938 = n10280 | n10488 ;
  assign n10939 = ( n10488 & n10489 ) | ( n10488 & n10938 ) | ( n10489 & n10938 ) ;
  assign n10940 = n10937 | n10939 ;
  assign n10941 = n10937 & n10939 ;
  assign n10942 = n10940 & ~n10941 ;
  assign n10943 = n10436 | n10494 ;
  assign n10944 = ( n10494 & n10495 ) | ( n10494 & n10943 ) | ( n10495 & n10943 ) ;
  assign n10945 = n10942 | n10944 ;
  assign n10946 = n10942 & n10944 ;
  assign n10947 = n10945 & ~n10946 ;
  assign n10948 = n10500 | n10502 ;
  assign n10949 = ( n10500 & n10501 ) | ( n10500 & n10948 ) | ( n10501 & n10948 ) ;
  assign n10950 = n10534 | n10538 ;
  assign n10951 = ( n10534 & n10536 ) | ( n10534 & n10950 ) | ( n10536 & n10950 ) ;
  assign n10952 = n10949 & ~n10951 ;
  assign n10953 = ~n10949 & n10951 ;
  assign n10954 = n10952 | n10953 ;
  assign n10955 = n10947 & n10954 ;
  assign n10956 = n10947 | n10954 ;
  assign n10957 = ~n10955 & n10956 ;
  assign n10958 = x21 & x44 ;
  assign n10959 = x22 & x43 ;
  assign n10960 = n10958 | n10959 ;
  assign n10961 = n1585 & n5658 ;
  assign n10962 = x8 & x57 ;
  assign n10963 = ~n10961 & n10962 ;
  assign n10964 = n10960 | n10961 ;
  assign n10965 = ( n10961 & n10963 ) | ( n10961 & n10964 ) | ( n10963 & n10964 ) ;
  assign n10966 = n10960 & ~n10965 ;
  assign n10967 = ( ~n10960 & n10961 ) | ( ~n10960 & n10962 ) | ( n10961 & n10962 ) ;
  assign n10968 = n10962 & n10967 ;
  assign n10969 = n10966 | n10968 ;
  assign n10970 = n10416 | n10562 ;
  assign n10971 = ( n10562 & n10565 ) | ( n10562 & n10970 ) | ( n10565 & n10970 ) ;
  assign n10972 = n10969 & ~n10971 ;
  assign n10973 = ~n10969 & n10971 ;
  assign n10974 = n10972 | n10973 ;
  assign n10975 = x58 & x60 ;
  assign n10976 = n135 & n10975 ;
  assign n10977 = n204 & n10370 ;
  assign n10978 = n10976 | n10977 ;
  assign n10979 = n200 & n9831 ;
  assign n10980 = x60 & n10979 ;
  assign n10981 = ( x60 & ~n10978 ) | ( x60 & n10980 ) | ( ~n10978 & n10980 ) ;
  assign n10982 = x5 & n10981 ;
  assign n10983 = n10978 | n10979 ;
  assign n10984 = x6 & x59 ;
  assign n10985 = x7 & x58 ;
  assign n10986 = ( ~n10979 & n10984 ) | ( ~n10979 & n10985 ) | ( n10984 & n10985 ) ;
  assign n10987 = n10984 & n10985 ;
  assign n10988 = ( ~n10978 & n10986 ) | ( ~n10978 & n10987 ) | ( n10986 & n10987 ) ;
  assign n10989 = ~n10983 & n10988 ;
  assign n10990 = n10982 | n10989 ;
  assign n10991 = n10974 & n10990 ;
  assign n10992 = n10974 | n10990 ;
  assign n10993 = ~n10991 & n10992 ;
  assign n10994 = x11 & x54 ;
  assign n10995 = x19 & x46 ;
  assign n10996 = n10994 | n10995 ;
  assign n10997 = x29 & x36 ;
  assign n10998 = ( n10994 & n10995 ) | ( n10994 & n10997 ) | ( n10995 & n10997 ) ;
  assign n10999 = n10996 & ~n10998 ;
  assign n11000 = n10994 & n10995 ;
  assign n11001 = n10997 & ~n11000 ;
  assign n11002 = ~n10996 & n10997 ;
  assign n11003 = ( n10997 & ~n11001 ) | ( n10997 & n11002 ) | ( ~n11001 & n11002 ) ;
  assign n11004 = n10999 | n11003 ;
  assign n11005 = n3321 & n4245 ;
  assign n11006 = n2965 & n3483 ;
  assign n11007 = n11005 | n11006 ;
  assign n11008 = n4062 & n4530 ;
  assign n11009 = n4245 & n11008 ;
  assign n11010 = ( n4245 & ~n11007 ) | ( n4245 & n11009 ) | ( ~n11007 & n11009 ) ;
  assign n11011 = n11007 | n11008 ;
  assign n11012 = ( n3321 & n7006 ) | ( n3321 & ~n11008 ) | ( n7006 & ~n11008 ) ;
  assign n11013 = n3321 & n7006 ;
  assign n11014 = ( ~n11007 & n11012 ) | ( ~n11007 & n11013 ) | ( n11012 & n11013 ) ;
  assign n11015 = ~n11011 & n11014 ;
  assign n11016 = n11010 | n11015 ;
  assign n11017 = ~n11004 & n11016 ;
  assign n11018 = n11004 & ~n11016 ;
  assign n11019 = n11017 | n11018 ;
  assign n11020 = x3 & x62 ;
  assign n11021 = x33 | n11020 ;
  assign n11022 = ( x33 & n7524 ) | ( x33 & n11020 ) | ( n7524 & n11020 ) ;
  assign n11023 = n11021 & ~n11022 ;
  assign n11024 = x33 & n11020 ;
  assign n11025 = n7524 & ~n11024 ;
  assign n11026 = n7524 & ~n11021 ;
  assign n11027 = ( n7524 & ~n11025 ) | ( n7524 & n11026 ) | ( ~n11025 & n11026 ) ;
  assign n11028 = n11023 | n11027 ;
  assign n11029 = n11019 & n11028 ;
  assign n11030 = n11019 | n11028 ;
  assign n11031 = ~n11029 & n11030 ;
  assign n11032 = n10993 & ~n11031 ;
  assign n11033 = ~n10993 & n11031 ;
  assign n11034 = n11032 | n11033 ;
  assign n11035 = x10 & x55 ;
  assign n11036 = x20 & x45 ;
  assign n11037 = n11035 & n11036 ;
  assign n11038 = x20 & x56 ;
  assign n11039 = n7551 & n11038 ;
  assign n11040 = n360 & n10013 ;
  assign n11041 = n11039 | n11040 ;
  assign n11042 = x56 & n11037 ;
  assign n11043 = ( x56 & ~n11041 ) | ( x56 & n11042 ) | ( ~n11041 & n11042 ) ;
  assign n11044 = x9 & n11043 ;
  assign n11045 = ( n11035 & n11036 ) | ( n11035 & ~n11041 ) | ( n11036 & ~n11041 ) ;
  assign n11046 = ( ~n11037 & n11044 ) | ( ~n11037 & n11045 ) | ( n11044 & n11045 ) ;
  assign n11047 = n1557 & n6973 ;
  assign n11048 = n1686 & n5710 ;
  assign n11049 = n11047 | n11048 ;
  assign n11050 = n1912 & n5813 ;
  assign n11051 = x42 & n11050 ;
  assign n11052 = ( x42 & ~n11049 ) | ( x42 & n11051 ) | ( ~n11049 & n11051 ) ;
  assign n11053 = x23 & n11052 ;
  assign n11054 = n11049 | n11050 ;
  assign n11055 = x24 & x41 ;
  assign n11056 = x25 & x40 ;
  assign n11057 = ( ~n11050 & n11055 ) | ( ~n11050 & n11056 ) | ( n11055 & n11056 ) ;
  assign n11058 = n11055 & n11056 ;
  assign n11059 = ( ~n11049 & n11057 ) | ( ~n11049 & n11058 ) | ( n11057 & n11058 ) ;
  assign n11060 = ~n11054 & n11059 ;
  assign n11061 = n11053 | n11060 ;
  assign n11062 = n11046 & n11061 ;
  assign n11063 = n11046 & ~n11062 ;
  assign n11064 = n11061 & ~n11062 ;
  assign n11065 = n11063 | n11064 ;
  assign n11066 = n2895 & n5798 ;
  assign n11067 = n2267 & n5392 ;
  assign n11068 = n11066 | n11067 ;
  assign n11069 = n2372 & n4857 ;
  assign n11070 = x39 & n11069 ;
  assign n11071 = ( x39 & ~n11068 ) | ( x39 & n11070 ) | ( ~n11068 & n11070 ) ;
  assign n11072 = x26 & n11071 ;
  assign n11073 = n11068 | n11069 ;
  assign n11074 = x27 & x38 ;
  assign n11075 = x28 & x37 ;
  assign n11076 = ( ~n11069 & n11074 ) | ( ~n11069 & n11075 ) | ( n11074 & n11075 ) ;
  assign n11077 = n11074 & n11075 ;
  assign n11078 = ( ~n11068 & n11076 ) | ( ~n11068 & n11077 ) | ( n11076 & n11077 ) ;
  assign n11079 = ~n11073 & n11078 ;
  assign n11080 = n11072 | n11079 ;
  assign n11081 = ~n11065 & n11080 ;
  assign n11082 = n11065 & ~n11080 ;
  assign n11083 = n11081 | n11082 ;
  assign n11084 = ~n11034 & n11083 ;
  assign n11085 = n11034 & ~n11083 ;
  assign n11086 = n11084 | n11085 ;
  assign n11087 = ( n10479 & n10481 ) | ( n10479 & n10505 ) | ( n10481 & n10505 ) ;
  assign n11088 = ( n10957 & n11086 ) | ( n10957 & ~n11087 ) | ( n11086 & ~n11087 ) ;
  assign n11089 = ( n10957 & ~n11086 ) | ( n10957 & n11087 ) | ( ~n11086 & n11087 ) ;
  assign n11090 = ( ~n10957 & n11088 ) | ( ~n10957 & n11089 ) | ( n11088 & n11089 ) ;
  assign n11091 = n10511 | n10515 ;
  assign n11092 = ( n10511 & n10514 ) | ( n10511 & n11091 ) | ( n10514 & n11091 ) ;
  assign n11093 = ( n10935 & n11090 ) | ( n10935 & ~n11092 ) | ( n11090 & ~n11092 ) ;
  assign n11094 = ( ~n11090 & n11092 ) | ( ~n11090 & n11093 ) | ( n11092 & n11093 ) ;
  assign n11095 = ( ~n10935 & n11093 ) | ( ~n10935 & n11094 ) | ( n11093 & n11094 ) ;
  assign n11096 = n10849 & n11095 ;
  assign n11097 = n10849 | n11095 ;
  assign n11098 = ~n11096 & n11097 ;
  assign n11099 = ( n10801 & n10802 ) | ( n10801 & ~n11098 ) | ( n10802 & ~n11098 ) ;
  assign n11100 = ( ~n10802 & n11098 ) | ( ~n10802 & n11099 ) | ( n11098 & n11099 ) ;
  assign n11101 = ( ~n10801 & n11099 ) | ( ~n10801 & n11100 ) | ( n11099 & n11100 ) ;
  assign n11102 = n10848 | n11096 ;
  assign n11103 = n11086 & n11087 ;
  assign n11104 = n11087 & ~n11103 ;
  assign n11105 = n11086 & ~n11087 ;
  assign n11106 = n10957 & n11105 ;
  assign n11107 = ( n10957 & n11104 ) | ( n10957 & n11106 ) | ( n11104 & n11106 ) ;
  assign n11108 = n11103 | n11107 ;
  assign n11109 = n10837 | n10841 ;
  assign n11110 = ( n10837 & n10839 ) | ( n10837 & n11109 ) | ( n10839 & n11109 ) ;
  assign n11111 = n11108 | n11110 ;
  assign n11112 = n169 & n10856 ;
  assign n11113 = n79 & n10561 ;
  assign n11114 = n11112 | n11113 ;
  assign n11115 = n91 & n10684 ;
  assign n11116 = x63 & n11115 ;
  assign n11117 = ( x63 & ~n11114 ) | ( x63 & n11116 ) | ( ~n11114 & n11116 ) ;
  assign n11118 = x3 & n11117 ;
  assign n11119 = n11114 | n11115 ;
  assign n11120 = x4 & x62 ;
  assign n11121 = ( n9739 & ~n11115 ) | ( n9739 & n11120 ) | ( ~n11115 & n11120 ) ;
  assign n11122 = n9739 & n11120 ;
  assign n11123 = ( ~n11114 & n11121 ) | ( ~n11114 & n11122 ) | ( n11121 & n11122 ) ;
  assign n11124 = ~n11119 & n11123 ;
  assign n11125 = n11118 | n11124 ;
  assign n11126 = n2075 & n5798 ;
  assign n11127 = n2372 & n5392 ;
  assign n11128 = n11126 | n11127 ;
  assign n11129 = n2369 & n4857 ;
  assign n11130 = x39 & n11129 ;
  assign n11131 = ( x39 & ~n11128 ) | ( x39 & n11130 ) | ( ~n11128 & n11130 ) ;
  assign n11132 = x27 & n11131 ;
  assign n11133 = n11128 | n11129 ;
  assign n11134 = x28 & x38 ;
  assign n11135 = x29 & x37 ;
  assign n11136 = ( ~n11129 & n11134 ) | ( ~n11129 & n11135 ) | ( n11134 & n11135 ) ;
  assign n11137 = n11134 & n11135 ;
  assign n11138 = ( ~n11128 & n11136 ) | ( ~n11128 & n11137 ) | ( n11136 & n11137 ) ;
  assign n11139 = ~n11133 & n11138 ;
  assign n11140 = n11132 | n11139 ;
  assign n11141 = n11125 & n11140 ;
  assign n11142 = n11125 & ~n11141 ;
  assign n11143 = n11140 & ~n11141 ;
  assign n11144 = n11142 | n11143 ;
  assign n11145 = x19 & x47 ;
  assign n11146 = x12 & x54 ;
  assign n11147 = n11145 & n11146 ;
  assign n11148 = n490 & n8357 ;
  assign n11149 = n8778 & n8913 ;
  assign n11150 = n11148 | n11149 ;
  assign n11151 = x55 & n11147 ;
  assign n11152 = ( x55 & ~n11150 ) | ( x55 & n11151 ) | ( ~n11150 & n11151 ) ;
  assign n11153 = x11 & n11152 ;
  assign n11154 = ( n11145 & n11146 ) | ( n11145 & ~n11150 ) | ( n11146 & ~n11150 ) ;
  assign n11155 = ( ~n11147 & n11153 ) | ( ~n11147 & n11154 ) | ( n11153 & n11154 ) ;
  assign n11156 = ~n11144 & n11155 ;
  assign n11157 = n11144 & ~n11155 ;
  assign n11158 = n11156 | n11157 ;
  assign n11159 = n1686 & n5407 ;
  assign n11160 = x43 & x57 ;
  assign n11161 = n2529 & n11160 ;
  assign n11162 = n11159 | n11161 ;
  assign n11163 = x24 & x57 ;
  assign n11164 = n6669 & n11163 ;
  assign n11165 = x43 & n11164 ;
  assign n11166 = ( x43 & ~n11162 ) | ( x43 & n11165 ) | ( ~n11162 & n11165 ) ;
  assign n11167 = x23 & n11166 ;
  assign n11168 = n11162 | n11164 ;
  assign n11169 = x9 & x57 ;
  assign n11170 = x24 & x42 ;
  assign n11171 = ( ~n11164 & n11169 ) | ( ~n11164 & n11170 ) | ( n11169 & n11170 ) ;
  assign n11172 = n11169 & n11170 ;
  assign n11173 = ( ~n11162 & n11171 ) | ( ~n11162 & n11172 ) | ( n11171 & n11172 ) ;
  assign n11174 = ~n11168 & n11173 ;
  assign n11175 = n11167 | n11174 ;
  assign n11176 = n1710 & n8407 ;
  assign n11177 = n1434 & n5975 ;
  assign n11178 = n11176 | n11177 ;
  assign n11179 = n1585 & n6093 ;
  assign n11180 = x46 & n11179 ;
  assign n11181 = ( x46 & ~n11178 ) | ( x46 & n11180 ) | ( ~n11178 & n11180 ) ;
  assign n11182 = x20 & n11181 ;
  assign n11183 = n11178 | n11179 ;
  assign n11184 = x21 & x45 ;
  assign n11185 = x22 & x44 ;
  assign n11186 = ( ~n11179 & n11184 ) | ( ~n11179 & n11185 ) | ( n11184 & n11185 ) ;
  assign n11187 = n11184 & n11185 ;
  assign n11188 = ( ~n11178 & n11186 ) | ( ~n11178 & n11187 ) | ( n11186 & n11187 ) ;
  assign n11189 = ~n11183 & n11188 ;
  assign n11190 = n11182 | n11189 ;
  assign n11191 = n11175 & n11190 ;
  assign n11192 = n11175 & ~n11191 ;
  assign n11193 = n11190 & ~n11191 ;
  assign n11194 = n11192 | n11193 ;
  assign n11195 = x25 & x41 ;
  assign n11196 = x26 & x40 ;
  assign n11197 = n11195 | n11196 ;
  assign n11198 = n2511 & n5813 ;
  assign n11199 = x10 & x56 ;
  assign n11200 = ~n11198 & n11199 ;
  assign n11201 = n11197 | n11198 ;
  assign n11202 = ( n11198 & n11200 ) | ( n11198 & n11201 ) | ( n11200 & n11201 ) ;
  assign n11203 = n11197 & ~n11202 ;
  assign n11204 = ( ~n11197 & n11198 ) | ( ~n11197 & n11199 ) | ( n11198 & n11199 ) ;
  assign n11205 = n11199 & n11204 ;
  assign n11206 = n11203 | n11205 ;
  assign n11207 = ~n11194 & n11206 ;
  assign n11208 = n11194 & ~n11206 ;
  assign n11209 = n11207 | n11208 ;
  assign n11210 = x31 & x35 ;
  assign n11211 = n4242 | n11210 ;
  assign n11212 = n2965 & n4078 ;
  assign n11213 = x14 & x52 ;
  assign n11214 = ~n11212 & n11213 ;
  assign n11215 = n11211 | n11212 ;
  assign n11216 = ( n11212 & n11214 ) | ( n11212 & n11215 ) | ( n11214 & n11215 ) ;
  assign n11217 = n11211 & ~n11216 ;
  assign n11218 = ( ~n11211 & n11212 ) | ( ~n11211 & n11213 ) | ( n11212 & n11213 ) ;
  assign n11219 = n11213 & n11218 ;
  assign n11220 = n11217 | n11219 ;
  assign n11221 = x13 & x53 ;
  assign n11222 = x15 & x51 ;
  assign n11223 = n11221 | n11222 ;
  assign n11224 = n723 & n7874 ;
  assign n11225 = n11223 | n11224 ;
  assign n11226 = x18 & x48 ;
  assign n11227 = ( ~n11224 & n11225 ) | ( ~n11224 & n11226 ) | ( n11225 & n11226 ) ;
  assign n11228 = ( n11224 & n11225 ) | ( n11224 & ~n11226 ) | ( n11225 & ~n11226 ) ;
  assign n11229 = ( ~n11225 & n11227 ) | ( ~n11225 & n11228 ) | ( n11227 & n11228 ) ;
  assign n11230 = n11220 & n11229 ;
  assign n11231 = n11220 & ~n11230 ;
  assign n11232 = n7666 | n8473 ;
  assign n11233 = n1023 & n6834 ;
  assign n11234 = n4318 & ~n11233 ;
  assign n11235 = n11232 | n11233 ;
  assign n11236 = ( n11233 & n11234 ) | ( n11233 & n11235 ) | ( n11234 & n11235 ) ;
  assign n11237 = n11232 & ~n11236 ;
  assign n11238 = n4318 & ~n11232 ;
  assign n11239 = ( n4318 & ~n11234 ) | ( n4318 & n11238 ) | ( ~n11234 & n11238 ) ;
  assign n11240 = n11237 | n11239 ;
  assign n11241 = ~n11220 & n11229 ;
  assign n11242 = n11240 & ~n11241 ;
  assign n11243 = ~n11231 & n11242 ;
  assign n11244 = ~n11240 & n11241 ;
  assign n11245 = ( n11231 & ~n11240 ) | ( n11231 & n11244 ) | ( ~n11240 & n11244 ) ;
  assign n11246 = n11243 | n11245 ;
  assign n11247 = n11209 & ~n11246 ;
  assign n11248 = ~n11209 & n11246 ;
  assign n11249 = n11247 | n11248 ;
  assign n11250 = n11158 & n11249 ;
  assign n11251 = n11158 | n11249 ;
  assign n11252 = ~n11250 & n11251 ;
  assign n11253 = ( n10803 & n10805 ) | ( n10803 & n10830 ) | ( n10805 & n10830 ) ;
  assign n11254 = n11252 & n11253 ;
  assign n11255 = n11252 | n11253 ;
  assign n11256 = ~n11254 & n11255 ;
  assign n11257 = n10624 | n10811 ;
  assign n11258 = ( n10811 & n10812 ) | ( n10811 & n11257 ) | ( n10812 & n11257 ) ;
  assign n11259 = n10817 | n10819 ;
  assign n11260 = ( n10819 & n10820 ) | ( n10819 & n11259 ) | ( n10820 & n11259 ) ;
  assign n11261 = n11258 | n11260 ;
  assign n11262 = n11258 & n11260 ;
  assign n11263 = n11261 & ~n11262 ;
  assign n11264 = n10589 | n10906 ;
  assign n11265 = ( n10906 & n10907 ) | ( n10906 & n11264 ) | ( n10907 & n11264 ) ;
  assign n11266 = n11263 | n11265 ;
  assign n11267 = n11263 & n11265 ;
  assign n11268 = n11266 & ~n11267 ;
  assign n11269 = n10825 | n10827 ;
  assign n11270 = ( n10825 & n10826 ) | ( n10825 & n11269 ) | ( n10826 & n11269 ) ;
  assign n11271 = n10913 | n10918 ;
  assign n11272 = ( n10913 & n10916 ) | ( n10913 & n11271 ) | ( n10916 & n11271 ) ;
  assign n11273 = n11270 & ~n11272 ;
  assign n11274 = ~n11270 & n11272 ;
  assign n11275 = n11273 | n11274 ;
  assign n11276 = n11268 & n11275 ;
  assign n11277 = n11268 | n11275 ;
  assign n11278 = ~n11276 & n11277 ;
  assign n11279 = n11256 & n11278 ;
  assign n11280 = n11256 | n11278 ;
  assign n11281 = ~n11279 & n11280 ;
  assign n11282 = ( n10837 & n10841 ) | ( n10837 & n11108 ) | ( n10841 & n11108 ) ;
  assign n11283 = n10837 & n11108 ;
  assign n11284 = ( n10839 & n11282 ) | ( n10839 & n11283 ) | ( n11282 & n11283 ) ;
  assign n11285 = n11281 & ~n11284 ;
  assign n11286 = n11111 & n11285 ;
  assign n11287 = ~n11281 & n11284 ;
  assign n11288 = ( n11111 & n11281 ) | ( n11111 & ~n11287 ) | ( n11281 & ~n11287 ) ;
  assign n11289 = ~n11286 & n11288 ;
  assign n11290 = n10511 & n10935 ;
  assign n11291 = ( n10515 & n10935 ) | ( n10515 & n11290 ) | ( n10935 & n11290 ) ;
  assign n11292 = n10935 & n11290 ;
  assign n11293 = ( n10514 & n11291 ) | ( n10514 & n11292 ) | ( n11291 & n11292 ) ;
  assign n11294 = n11092 & ~n11293 ;
  assign n11295 = n10935 & n11090 ;
  assign n11296 = ~n11290 & n11295 ;
  assign n11297 = ~n10516 & n11296 ;
  assign n11298 = ( n11090 & n11294 ) | ( n11090 & n11297 ) | ( n11294 & n11297 ) ;
  assign n11299 = n10880 & n10891 ;
  assign n11300 = n10891 & ~n11299 ;
  assign n11301 = n10880 & ~n10891 ;
  assign n11302 = n10865 & ~n11301 ;
  assign n11303 = ~n11300 & n11302 ;
  assign n11304 = ( n10865 & n11299 ) | ( n10865 & ~n11303 ) | ( n11299 & ~n11303 ) ;
  assign n11305 = n10857 & n11069 ;
  assign n11306 = ( n10857 & n11068 ) | ( n10857 & n11305 ) | ( n11068 & n11305 ) ;
  assign n11307 = ( n10862 & n11073 ) | ( n10862 & n11306 ) | ( n11073 & n11306 ) ;
  assign n11308 = n10857 | n11069 ;
  assign n11309 = n11068 | n11308 ;
  assign n11310 = n10862 | n11309 ;
  assign n11311 = ~n11307 & n11310 ;
  assign n11312 = n181 & n10975 ;
  assign n11313 = n200 & n10370 ;
  assign n11314 = n11312 | n11313 ;
  assign n11315 = n251 & n9831 ;
  assign n11316 = x60 & n11315 ;
  assign n11317 = ( x60 & ~n11314 ) | ( x60 & n11316 ) | ( ~n11314 & n11316 ) ;
  assign n11318 = x6 & n11317 ;
  assign n11319 = n11314 | n11315 ;
  assign n11320 = x7 & x59 ;
  assign n11321 = x8 & x58 ;
  assign n11322 = ( ~n11315 & n11320 ) | ( ~n11315 & n11321 ) | ( n11320 & n11321 ) ;
  assign n11323 = n11320 & n11321 ;
  assign n11324 = ( ~n11314 & n11322 ) | ( ~n11314 & n11323 ) | ( n11322 & n11323 ) ;
  assign n11325 = ~n11319 & n11324 ;
  assign n11326 = n11318 | n11325 ;
  assign n11327 = n11311 & ~n11326 ;
  assign n11328 = n11311 | n11326 ;
  assign n11329 = ( ~n11311 & n11327 ) | ( ~n11311 & n11328 ) | ( n11327 & n11328 ) ;
  assign n11330 = n11304 & n11329 ;
  assign n11331 = n11304 & ~n11330 ;
  assign n11332 = ~n11304 & n11329 ;
  assign n11333 = n10941 | n10944 ;
  assign n11334 = ( n10941 & n10942 ) | ( n10941 & n11333 ) | ( n10942 & n11333 ) ;
  assign n11335 = n11332 | n11334 ;
  assign n11336 = n11331 | n11335 ;
  assign n11337 = n11332 & n11334 ;
  assign n11338 = ( n11331 & n11334 ) | ( n11331 & n11337 ) | ( n11334 & n11337 ) ;
  assign n11339 = n11336 & ~n11338 ;
  assign n11340 = n11008 | n11022 ;
  assign n11341 = n11007 | n11340 ;
  assign n11342 = n11008 & n11022 ;
  assign n11343 = ( n11007 & n11022 ) | ( n11007 & n11342 ) | ( n11022 & n11342 ) ;
  assign n11344 = n11341 & ~n11343 ;
  assign n11345 = n10873 | n11344 ;
  assign n11346 = n10873 & n11344 ;
  assign n11347 = n11345 & ~n11346 ;
  assign n11348 = n10965 | n10983 ;
  assign n11349 = n10965 & n10983 ;
  assign n11350 = n11348 & ~n11349 ;
  assign n11351 = n10998 | n11350 ;
  assign n11352 = n10998 & n11350 ;
  assign n11353 = n11351 & ~n11352 ;
  assign n11354 = n11004 & n11016 ;
  assign n11355 = n11353 & n11354 ;
  assign n11356 = ( n11029 & n11353 ) | ( n11029 & n11355 ) | ( n11353 & n11355 ) ;
  assign n11357 = n11353 | n11354 ;
  assign n11358 = n11029 | n11357 ;
  assign n11359 = ~n11356 & n11358 ;
  assign n11360 = n11347 & n11359 ;
  assign n11361 = n11347 | n11359 ;
  assign n11362 = ~n11360 & n11361 ;
  assign n11363 = n11339 & n11362 ;
  assign n11364 = n11339 | n11362 ;
  assign n11365 = ~n11363 & n11364 ;
  assign n11366 = ( n10947 & n10949 ) | ( n10947 & n10951 ) | ( n10949 & n10951 ) ;
  assign n11367 = n11365 & n11366 ;
  assign n11368 = n11365 | n11366 ;
  assign n11369 = ~n11367 & n11368 ;
  assign n11370 = n10923 | n10932 ;
  assign n11371 = n10883 | n10886 ;
  assign n11372 = n11037 | n11041 ;
  assign n11373 = n11371 | n11372 ;
  assign n11374 = n11371 & n11372 ;
  assign n11375 = n11373 & ~n11374 ;
  assign n11376 = n11054 | n11375 ;
  assign n11377 = n11054 & n11375 ;
  assign n11378 = n11376 & ~n11377 ;
  assign n11379 = ( n10969 & n10971 ) | ( n10969 & n10990 ) | ( n10971 & n10990 ) ;
  assign n11380 = n11378 | n11379 ;
  assign n11381 = n11378 & n11379 ;
  assign n11382 = n11380 & ~n11381 ;
  assign n11383 = n11062 | n11080 ;
  assign n11384 = ( n11062 & n11065 ) | ( n11062 & n11383 ) | ( n11065 & n11383 ) ;
  assign n11385 = n11382 | n11384 ;
  assign n11386 = n11382 & n11384 ;
  assign n11387 = n11385 & ~n11386 ;
  assign n11388 = ( n10993 & n11031 ) | ( n10993 & n11083 ) | ( n11031 & n11083 ) ;
  assign n11389 = ( n10854 & n10855 ) | ( n10854 & n10897 ) | ( n10855 & n10897 ) ;
  assign n11390 = n11388 | n11389 ;
  assign n11391 = n11388 & n11389 ;
  assign n11392 = n11390 & ~n11391 ;
  assign n11393 = n11387 & n11392 ;
  assign n11394 = n11387 | n11392 ;
  assign n11395 = ~n11393 & n11394 ;
  assign n11396 = n10923 & n11395 ;
  assign n11397 = ( n10932 & n11395 ) | ( n10932 & n11396 ) | ( n11395 & n11396 ) ;
  assign n11398 = n11370 & ~n11397 ;
  assign n11399 = ~n10923 & n11395 ;
  assign n11400 = ~n10932 & n11399 ;
  assign n11401 = n11369 & n11400 ;
  assign n11402 = ( n11369 & n11398 ) | ( n11369 & n11401 ) | ( n11398 & n11401 ) ;
  assign n11403 = n11369 | n11400 ;
  assign n11404 = n11398 | n11403 ;
  assign n11405 = ~n11402 & n11404 ;
  assign n11406 = n11293 & n11405 ;
  assign n11407 = ( n11298 & n11405 ) | ( n11298 & n11406 ) | ( n11405 & n11406 ) ;
  assign n11408 = n11293 | n11405 ;
  assign n11409 = n11298 | n11408 ;
  assign n11410 = ~n11407 & n11409 ;
  assign n11411 = n11289 & ~n11410 ;
  assign n11412 = n11102 & n11411 ;
  assign n11413 = ~n11289 & n11410 ;
  assign n11414 = ( n11102 & n11412 ) | ( n11102 & n11413 ) | ( n11412 & n11413 ) ;
  assign n11415 = n11102 | n11411 ;
  assign n11416 = n11413 | n11415 ;
  assign n11417 = ~n11414 & n11416 ;
  assign n11418 = n10802 & n11098 ;
  assign n11419 = n10802 | n11098 ;
  assign n11420 = n10785 & n11419 ;
  assign n11421 = ( n10799 & n11419 ) | ( n10799 & n11420 ) | ( n11419 & n11420 ) ;
  assign n11422 = n11418 | n11421 ;
  assign n11423 = n11418 | n11419 ;
  assign n11424 = ( n10786 & n11418 ) | ( n10786 & n11423 ) | ( n11418 & n11423 ) ;
  assign n11425 = ( n10794 & n11422 ) | ( n10794 & n11424 ) | ( n11422 & n11424 ) ;
  assign n11426 = n11417 & n11425 ;
  assign n11427 = n11417 | n11425 ;
  assign n11428 = ~n11426 & n11427 ;
  assign n11429 = n11414 | n11416 ;
  assign n11430 = ( n11414 & n11424 ) | ( n11414 & n11429 ) | ( n11424 & n11429 ) ;
  assign n11431 = n11416 & n11418 ;
  assign n11432 = n11414 | n11431 ;
  assign n11433 = ( n11421 & n11429 ) | ( n11421 & n11432 ) | ( n11429 & n11432 ) ;
  assign n11434 = ( n10794 & n11430 ) | ( n10794 & n11433 ) | ( n11430 & n11433 ) ;
  assign n11435 = x14 & x53 ;
  assign n11436 = n8044 & n11435 ;
  assign n11437 = x48 & x53 ;
  assign n11438 = x14 & n11437 ;
  assign n11439 = x17 & n6345 ;
  assign n11440 = n11438 | n11439 ;
  assign n11441 = x19 & ~n11436 ;
  assign n11442 = n11440 & n11441 ;
  assign n11443 = x19 & x48 ;
  assign n11444 = ~n11442 & n11443 ;
  assign n11445 = ( n8044 & n11435 ) | ( n8044 & ~n11442 ) | ( n11435 & ~n11442 ) ;
  assign n11446 = ( ~n11436 & n11444 ) | ( ~n11436 & n11445 ) | ( n11444 & n11445 ) ;
  assign n11447 = x21 & x46 ;
  assign n11448 = x26 & x41 ;
  assign n11449 = n11447 & n11448 ;
  assign n11450 = n2511 & n5710 ;
  assign n11451 = x25 & x46 ;
  assign n11452 = n10387 & n11451 ;
  assign n11453 = n11450 | n11452 ;
  assign n11454 = x42 & n11449 ;
  assign n11455 = ( x42 & ~n11453 ) | ( x42 & n11454 ) | ( ~n11453 & n11454 ) ;
  assign n11456 = x25 & n11455 ;
  assign n11457 = ( n11447 & n11448 ) | ( n11447 & ~n11453 ) | ( n11448 & ~n11453 ) ;
  assign n11458 = ( ~n11449 & n11456 ) | ( ~n11449 & n11457 ) | ( n11456 & n11457 ) ;
  assign n11459 = n11446 & n11458 ;
  assign n11460 = n11446 & ~n11459 ;
  assign n11461 = n11458 & ~n11459 ;
  assign n11462 = n11460 | n11461 ;
  assign n11463 = x27 & x40 ;
  assign n11464 = x28 & x39 ;
  assign n11465 = n11463 | n11464 ;
  assign n11466 = n2372 & n4555 ;
  assign n11467 = x4 & x63 ;
  assign n11468 = ~n11466 & n11467 ;
  assign n11469 = n11465 | n11466 ;
  assign n11470 = ( n11466 & n11468 ) | ( n11466 & n11469 ) | ( n11468 & n11469 ) ;
  assign n11471 = n11465 & ~n11470 ;
  assign n11472 = ( ~n11465 & n11466 ) | ( ~n11465 & n11467 ) | ( n11466 & n11467 ) ;
  assign n11473 = n11467 & n11472 ;
  assign n11474 = n11471 | n11473 ;
  assign n11475 = ~n11462 & n11474 ;
  assign n11476 = n11462 & ~n11474 ;
  assign n11477 = n11475 | n11476 ;
  assign n11478 = n667 & n10975 ;
  assign n11479 = n251 & n10370 ;
  assign n11480 = n11478 | n11479 ;
  assign n11481 = n313 & n9831 ;
  assign n11482 = x60 & n11481 ;
  assign n11483 = ( x60 & ~n11480 ) | ( x60 & n11482 ) | ( ~n11480 & n11482 ) ;
  assign n11484 = x7 & n11483 ;
  assign n11485 = n11480 | n11481 ;
  assign n11486 = x8 & x59 ;
  assign n11487 = x9 & x58 ;
  assign n11488 = ( ~n11481 & n11486 ) | ( ~n11481 & n11487 ) | ( n11486 & n11487 ) ;
  assign n11489 = n11486 & n11487 ;
  assign n11490 = ( ~n11480 & n11488 ) | ( ~n11480 & n11489 ) | ( n11488 & n11489 ) ;
  assign n11491 = ~n11485 & n11490 ;
  assign n11492 = n11484 | n11491 ;
  assign n11493 = n2148 & n5104 ;
  assign n11494 = n1932 & n6093 ;
  assign n11495 = n11493 | n11494 ;
  assign n11496 = n1686 & n5658 ;
  assign n11497 = x45 & n11496 ;
  assign n11498 = ( x45 & ~n11495 ) | ( x45 & n11497 ) | ( ~n11495 & n11497 ) ;
  assign n11499 = x22 & n11498 ;
  assign n11500 = n11495 | n11496 ;
  assign n11501 = x23 & x44 ;
  assign n11502 = x24 & x43 ;
  assign n11503 = ( ~n11496 & n11501 ) | ( ~n11496 & n11502 ) | ( n11501 & n11502 ) ;
  assign n11504 = n11501 & n11502 ;
  assign n11505 = ( ~n11495 & n11503 ) | ( ~n11495 & n11504 ) | ( n11503 & n11504 ) ;
  assign n11506 = ~n11500 & n11505 ;
  assign n11507 = n11499 | n11506 ;
  assign n11508 = n11492 & n11507 ;
  assign n11509 = n11492 & ~n11508 ;
  assign n11510 = n11507 & ~n11508 ;
  assign n11511 = n11509 | n11510 ;
  assign n11512 = x16 & x51 ;
  assign n11513 = x30 & x37 ;
  assign n11514 = n11512 & n11513 ;
  assign n11515 = n795 & n7567 ;
  assign n11516 = x37 & x52 ;
  assign n11517 = n5248 & n11516 ;
  assign n11518 = n11515 | n11517 ;
  assign n11519 = x52 & n11514 ;
  assign n11520 = ( x52 & ~n11518 ) | ( x52 & n11519 ) | ( ~n11518 & n11519 ) ;
  assign n11521 = x15 & n11520 ;
  assign n11522 = ( n11512 & n11513 ) | ( n11512 & ~n11518 ) | ( n11513 & ~n11518 ) ;
  assign n11523 = ( ~n11514 & n11521 ) | ( ~n11514 & n11522 ) | ( n11521 & n11522 ) ;
  assign n11524 = ~n11511 & n11523 ;
  assign n11525 = n11511 & ~n11523 ;
  assign n11526 = n11524 | n11525 ;
  assign n11527 = x5 & x62 ;
  assign n11528 = x34 | n11527 ;
  assign n11529 = x18 & x49 ;
  assign n11530 = ( x34 & n11527 ) | ( x34 & n11529 ) | ( n11527 & n11529 ) ;
  assign n11531 = n11528 & ~n11530 ;
  assign n11532 = x62 & n3874 ;
  assign n11533 = n11528 & ~n11532 ;
  assign n11534 = n11529 & ~n11533 ;
  assign n11535 = n11531 | n11534 ;
  assign n11536 = n4509 & n4530 ;
  assign n11537 = n4062 & n4078 ;
  assign n11538 = n11536 | n11537 ;
  assign n11539 = n3321 & n3483 ;
  assign n11540 = n4509 & n11539 ;
  assign n11541 = ( n4509 & ~n11538 ) | ( n4509 & n11540 ) | ( ~n11538 & n11540 ) ;
  assign n11542 = n11538 | n11539 ;
  assign n11543 = ( n4530 & n7386 ) | ( n4530 & ~n11539 ) | ( n7386 & ~n11539 ) ;
  assign n11544 = n4530 & n7386 ;
  assign n11545 = ( ~n11538 & n11543 ) | ( ~n11538 & n11544 ) | ( n11543 & n11544 ) ;
  assign n11546 = ~n11542 & n11545 ;
  assign n11547 = n11541 | n11546 ;
  assign n11548 = ~n11535 & n11547 ;
  assign n11549 = n11535 & ~n11547 ;
  assign n11550 = n11548 | n11549 ;
  assign n11551 = x12 & x55 ;
  assign n11552 = x13 & x54 ;
  assign n11553 = n11551 | n11552 ;
  assign n11554 = n647 & n8357 ;
  assign n11555 = x29 & x38 ;
  assign n11556 = ~n11554 & n11555 ;
  assign n11557 = n11553 | n11554 ;
  assign n11558 = ( n11554 & n11556 ) | ( n11554 & n11557 ) | ( n11556 & n11557 ) ;
  assign n11559 = n11553 & ~n11558 ;
  assign n11560 = ~n11553 & n11555 ;
  assign n11561 = ( n11555 & ~n11556 ) | ( n11555 & n11560 ) | ( ~n11556 & n11560 ) ;
  assign n11562 = n11559 | n11561 ;
  assign n11563 = n11550 & n11562 ;
  assign n11564 = n11550 | n11562 ;
  assign n11565 = ~n11563 & n11564 ;
  assign n11566 = ~n11526 & n11565 ;
  assign n11567 = n11526 & ~n11565 ;
  assign n11568 = n11566 | n11567 ;
  assign n11569 = n11477 & n11568 ;
  assign n11570 = n11477 | n11568 ;
  assign n11571 = ~n11569 & n11570 ;
  assign n11572 = ( n11387 & n11388 ) | ( n11387 & n11389 ) | ( n11388 & n11389 ) ;
  assign n11573 = n11571 & n11572 ;
  assign n11574 = n11571 | n11572 ;
  assign n11575 = ~n11573 & n11574 ;
  assign n11576 = n10998 | n11349 ;
  assign n11577 = ( n11349 & n11350 ) | ( n11349 & n11576 ) | ( n11350 & n11576 ) ;
  assign n11578 = n11054 | n11374 ;
  assign n11579 = ( n11374 & n11375 ) | ( n11374 & n11578 ) | ( n11375 & n11578 ) ;
  assign n11580 = n11577 | n11579 ;
  assign n11581 = n11577 & n11579 ;
  assign n11582 = n11580 & ~n11581 ;
  assign n11583 = n10873 | n11343 ;
  assign n11584 = ( n11343 & n11344 ) | ( n11343 & n11583 ) | ( n11344 & n11583 ) ;
  assign n11585 = n11582 | n11584 ;
  assign n11586 = n11582 & n11584 ;
  assign n11587 = n11585 & ~n11586 ;
  assign n11588 = n11381 | n11386 ;
  assign n11589 = n11347 | n11356 ;
  assign n11590 = ( n11356 & n11359 ) | ( n11356 & n11589 ) | ( n11359 & n11589 ) ;
  assign n11591 = n11588 | n11590 ;
  assign n11592 = n11588 & n11590 ;
  assign n11593 = n11591 & ~n11592 ;
  assign n11594 = n11587 & n11593 ;
  assign n11595 = n11587 | n11593 ;
  assign n11596 = ~n11594 & n11595 ;
  assign n11597 = n11575 & n11596 ;
  assign n11598 = n11575 | n11596 ;
  assign n11599 = ~n11597 & n11598 ;
  assign n11600 = n11191 | n11206 ;
  assign n11601 = n11307 | n11326 ;
  assign n11602 = ( n11307 & n11311 ) | ( n11307 & n11601 ) | ( n11311 & n11601 ) ;
  assign n11603 = n11600 & n11602 ;
  assign n11604 = n11191 & n11602 ;
  assign n11605 = ( n11194 & n11603 ) | ( n11194 & n11604 ) | ( n11603 & n11604 ) ;
  assign n11606 = n11600 | n11602 ;
  assign n11607 = n11191 | n11602 ;
  assign n11608 = ( n11194 & n11606 ) | ( n11194 & n11607 ) | ( n11606 & n11607 ) ;
  assign n11609 = ~n11605 & n11608 ;
  assign n11610 = n11141 | n11155 ;
  assign n11611 = ( n11141 & n11144 ) | ( n11141 & n11610 ) | ( n11144 & n11610 ) ;
  assign n11612 = n11609 | n11611 ;
  assign n11613 = n11609 & n11611 ;
  assign n11614 = n11612 & ~n11613 ;
  assign n11615 = n11119 | n11319 ;
  assign n11616 = n11119 & n11319 ;
  assign n11617 = n11615 & ~n11616 ;
  assign n11618 = n11133 | n11617 ;
  assign n11619 = n11133 & n11617 ;
  assign n11620 = n11618 & ~n11619 ;
  assign n11621 = n11168 | n11202 ;
  assign n11622 = n11168 & n11202 ;
  assign n11623 = n11621 & ~n11622 ;
  assign n11624 = n11183 | n11623 ;
  assign n11625 = n11183 & n11623 ;
  assign n11626 = n11624 & ~n11625 ;
  assign n11627 = x6 & x61 ;
  assign n11628 = n11236 & n11627 ;
  assign n11629 = n11236 | n11627 ;
  assign n11630 = ~n11628 & n11629 ;
  assign n11631 = n11216 | n11630 ;
  assign n11632 = n11216 & n11630 ;
  assign n11633 = n11631 & ~n11632 ;
  assign n11634 = n11626 & n11633 ;
  assign n11635 = n11626 | n11633 ;
  assign n11636 = ~n11634 & n11635 ;
  assign n11637 = n11620 & n11636 ;
  assign n11638 = n11620 | n11636 ;
  assign n11639 = ~n11637 & n11638 ;
  assign n11640 = n11614 & n11639 ;
  assign n11641 = n11614 | n11639 ;
  assign n11642 = ~n11640 & n11641 ;
  assign n11643 = ( n11268 & n11270 ) | ( n11268 & n11272 ) | ( n11270 & n11272 ) ;
  assign n11644 = n11642 & n11643 ;
  assign n11645 = n11642 | n11643 ;
  assign n11646 = ~n11644 & n11645 ;
  assign n11647 = n11362 | n11366 ;
  assign n11648 = ( n11339 & n11366 ) | ( n11339 & n11647 ) | ( n11366 & n11647 ) ;
  assign n11649 = ( n11363 & n11365 ) | ( n11363 & n11648 ) | ( n11365 & n11648 ) ;
  assign n11650 = n11646 | n11649 ;
  assign n11651 = n11646 & n11649 ;
  assign n11652 = n11650 & ~n11651 ;
  assign n11653 = ~n11224 & n11226 ;
  assign n11654 = ( n11224 & n11225 ) | ( n11224 & n11653 ) | ( n11225 & n11653 ) ;
  assign n11655 = n11147 | n11150 ;
  assign n11656 = n11654 | n11655 ;
  assign n11657 = n11654 & n11655 ;
  assign n11658 = n11656 & ~n11657 ;
  assign n11659 = n618 & n8903 ;
  assign n11660 = x20 & x57 ;
  assign n11661 = n8390 & n11660 ;
  assign n11662 = n11659 | n11661 ;
  assign n11663 = n8778 & n11038 ;
  assign n11664 = x57 & n11663 ;
  assign n11665 = ( x57 & ~n11662 ) | ( x57 & n11664 ) | ( ~n11662 & n11664 ) ;
  assign n11666 = x10 & n11665 ;
  assign n11667 = n11662 | n11663 ;
  assign n11668 = x11 & x56 ;
  assign n11669 = x20 & x47 ;
  assign n11670 = ( ~n11663 & n11668 ) | ( ~n11663 & n11669 ) | ( n11668 & n11669 ) ;
  assign n11671 = n11668 & n11669 ;
  assign n11672 = ( ~n11662 & n11670 ) | ( ~n11662 & n11671 ) | ( n11670 & n11671 ) ;
  assign n11673 = ~n11667 & n11672 ;
  assign n11674 = n11666 | n11673 ;
  assign n11675 = n11658 & n11674 ;
  assign n11676 = n11658 & ~n11675 ;
  assign n11677 = n11674 & ~n11675 ;
  assign n11678 = n11676 | n11677 ;
  assign n11679 = n11240 & n11241 ;
  assign n11680 = ( n11231 & n11240 ) | ( n11231 & n11679 ) | ( n11240 & n11679 ) ;
  assign n11681 = n11230 | n11680 ;
  assign n11682 = n11678 | n11681 ;
  assign n11683 = n11678 & n11681 ;
  assign n11684 = n11682 & ~n11683 ;
  assign n11685 = n11262 | n11265 ;
  assign n11686 = ( n11262 & n11263 ) | ( n11262 & n11685 ) | ( n11263 & n11685 ) ;
  assign n11687 = n11684 | n11686 ;
  assign n11688 = n11684 & n11686 ;
  assign n11689 = n11687 & ~n11688 ;
  assign n11690 = ( n11158 & n11209 ) | ( n11158 & n11246 ) | ( n11209 & n11246 ) ;
  assign n11691 = n11330 | n11690 ;
  assign n11692 = n11338 | n11691 ;
  assign n11693 = n11330 & n11690 ;
  assign n11694 = ( n11338 & n11690 ) | ( n11338 & n11693 ) | ( n11690 & n11693 ) ;
  assign n11695 = n11692 & ~n11694 ;
  assign n11696 = n11689 & n11695 ;
  assign n11697 = n11689 | n11695 ;
  assign n11698 = ~n11696 & n11697 ;
  assign n11699 = n11652 & n11698 ;
  assign n11700 = n11652 | n11698 ;
  assign n11701 = ~n11699 & n11700 ;
  assign n11702 = n11284 & n11701 ;
  assign n11703 = ( n11286 & n11701 ) | ( n11286 & n11702 ) | ( n11701 & n11702 ) ;
  assign n11704 = n11284 | n11701 ;
  assign n11705 = n11286 | n11704 ;
  assign n11706 = ~n11703 & n11705 ;
  assign n11707 = ( n11252 & n11253 ) | ( n11252 & n11278 ) | ( n11253 & n11278 ) ;
  assign n11708 = n11397 & n11707 ;
  assign n11709 = ( n11402 & n11707 ) | ( n11402 & n11708 ) | ( n11707 & n11708 ) ;
  assign n11710 = n11397 | n11707 ;
  assign n11711 = n11402 | n11710 ;
  assign n11712 = ~n11709 & n11711 ;
  assign n11713 = ( n11599 & n11706 ) | ( n11599 & ~n11712 ) | ( n11706 & ~n11712 ) ;
  assign n11714 = ( ~n11706 & n11712 ) | ( ~n11706 & n11713 ) | ( n11712 & n11713 ) ;
  assign n11715 = ( ~n11599 & n11713 ) | ( ~n11599 & n11714 ) | ( n11713 & n11714 ) ;
  assign n11716 = n11289 | n11407 ;
  assign n11717 = ( n11407 & n11410 ) | ( n11407 & n11716 ) | ( n11410 & n11716 ) ;
  assign n11718 = ( n11434 & n11715 ) | ( n11434 & ~n11717 ) | ( n11715 & ~n11717 ) ;
  assign n11719 = ( ~n11715 & n11717 ) | ( ~n11715 & n11718 ) | ( n11717 & n11718 ) ;
  assign n11720 = ( ~n11434 & n11718 ) | ( ~n11434 & n11719 ) | ( n11718 & n11719 ) ;
  assign n11721 = n11715 & n11717 ;
  assign n11722 = n11715 | n11717 ;
  assign n11723 = n11433 & n11722 ;
  assign n11724 = n11429 & n11722 ;
  assign n11725 = n11414 & n11722 ;
  assign n11726 = ( n11424 & n11724 ) | ( n11424 & n11725 ) | ( n11724 & n11725 ) ;
  assign n11727 = ( n10794 & n11723 ) | ( n10794 & n11726 ) | ( n11723 & n11726 ) ;
  assign n11728 = n11721 | n11727 ;
  assign n11729 = n11599 | n11708 ;
  assign n11730 = n11599 | n11707 ;
  assign n11731 = ( n11402 & n11729 ) | ( n11402 & n11730 ) | ( n11729 & n11730 ) ;
  assign n11732 = ( n11709 & n11712 ) | ( n11709 & n11731 ) | ( n11712 & n11731 ) ;
  assign n11733 = n11436 | n11442 ;
  assign n11734 = n11449 | n11453 ;
  assign n11735 = n11733 | n11734 ;
  assign n11736 = n11733 & n11734 ;
  assign n11737 = n11735 & ~n11736 ;
  assign n11738 = n11558 | n11737 ;
  assign n11739 = n11558 & n11737 ;
  assign n11740 = n11738 & ~n11739 ;
  assign n11741 = n11535 & n11547 ;
  assign n11742 = n11562 | n11741 ;
  assign n11743 = ( n11550 & n11741 ) | ( n11550 & n11742 ) | ( n11741 & n11742 ) ;
  assign n11744 = n11459 | n11474 ;
  assign n11745 = ( n11459 & n11462 ) | ( n11459 & n11744 ) | ( n11462 & n11744 ) ;
  assign n11746 = n11743 | n11745 ;
  assign n11747 = n11743 & n11745 ;
  assign n11748 = n11746 & ~n11747 ;
  assign n11749 = n11740 & n11748 ;
  assign n11750 = n11740 | n11748 ;
  assign n11751 = ~n11749 & n11750 ;
  assign n11752 = n11500 | n11667 ;
  assign n11753 = n11500 & n11667 ;
  assign n11754 = n11752 & ~n11753 ;
  assign n11755 = n11485 | n11754 ;
  assign n11756 = n11485 & n11754 ;
  assign n11757 = n11755 & ~n11756 ;
  assign n11758 = n11470 | n11542 ;
  assign n11759 = n11470 & n11542 ;
  assign n11760 = n11758 & ~n11759 ;
  assign n11761 = n11514 | n11518 ;
  assign n11762 = n11760 | n11761 ;
  assign n11763 = n11760 & n11761 ;
  assign n11764 = n11762 & ~n11763 ;
  assign n11765 = n11757 & n11764 ;
  assign n11766 = n11757 | n11764 ;
  assign n11767 = ~n11765 & n11766 ;
  assign n11768 = n11581 | n11584 ;
  assign n11769 = ( n11581 & n11582 ) | ( n11581 & n11768 ) | ( n11582 & n11768 ) ;
  assign n11770 = n11767 & n11769 ;
  assign n11771 = n11767 | n11769 ;
  assign n11772 = ~n11770 & n11771 ;
  assign n11773 = n11751 & n11772 ;
  assign n11774 = n11751 | n11772 ;
  assign n11775 = ~n11773 & n11774 ;
  assign n11776 = n11587 | n11592 ;
  assign n11777 = ( n11592 & n11593 ) | ( n11592 & n11776 ) | ( n11593 & n11776 ) ;
  assign n11778 = n11775 & n11777 ;
  assign n11779 = n11775 | n11777 ;
  assign n11780 = ~n11778 & n11779 ;
  assign n11781 = n11657 | n11675 ;
  assign n11782 = n11183 | n11622 ;
  assign n11783 = ( n11622 & n11623 ) | ( n11622 & n11782 ) | ( n11623 & n11782 ) ;
  assign n11784 = n11781 | n11783 ;
  assign n11785 = n11781 & n11783 ;
  assign n11786 = n11784 & ~n11785 ;
  assign n11787 = n11508 | n11523 ;
  assign n11788 = ( n11508 & n11511 ) | ( n11508 & n11787 ) | ( n11511 & n11787 ) ;
  assign n11789 = n11786 | n11788 ;
  assign n11790 = n11786 & n11788 ;
  assign n11791 = n11789 & ~n11790 ;
  assign n11792 = n251 & n10367 ;
  assign n11793 = x8 & x60 ;
  assign n11794 = x7 & x61 ;
  assign n11795 = n11793 | n11794 ;
  assign n11796 = ~n11792 & n11795 ;
  assign n11797 = n11530 & n11796 ;
  assign n11798 = n11796 & ~n11797 ;
  assign n11799 = n11530 & ~n11796 ;
  assign n11800 = n11798 | n11799 ;
  assign n11801 = n11216 | n11628 ;
  assign n11802 = ( n11628 & n11630 ) | ( n11628 & n11801 ) | ( n11630 & n11801 ) ;
  assign n11803 = n11800 | n11802 ;
  assign n11804 = n11800 & n11802 ;
  assign n11805 = n11803 & ~n11804 ;
  assign n11806 = n11133 | n11616 ;
  assign n11807 = ( n11616 & n11617 ) | ( n11616 & n11806 ) | ( n11617 & n11806 ) ;
  assign n11808 = n11805 | n11807 ;
  assign n11809 = n11805 & n11807 ;
  assign n11810 = n11808 & ~n11809 ;
  assign n11811 = n11791 & n11810 ;
  assign n11812 = n11791 | n11810 ;
  assign n11813 = ~n11811 & n11812 ;
  assign n11814 = ( n11477 & n11526 ) | ( n11477 & n11565 ) | ( n11526 & n11565 ) ;
  assign n11815 = n11813 & n11814 ;
  assign n11816 = n11813 | n11814 ;
  assign n11817 = ~n11815 & n11816 ;
  assign n11818 = n11640 | n11643 ;
  assign n11819 = ( n11640 & n11642 ) | ( n11640 & n11818 ) | ( n11642 & n11818 ) ;
  assign n11820 = n11817 & n11819 ;
  assign n11821 = n11819 & ~n11820 ;
  assign n11822 = ( n11817 & ~n11820 ) | ( n11817 & n11821 ) | ( ~n11820 & n11821 ) ;
  assign n11823 = n11780 & ~n11822 ;
  assign n11824 = ~n11780 & n11822 ;
  assign n11825 = n11823 | n11824 ;
  assign n11826 = n11731 & n11825 ;
  assign n11827 = n11709 & n11825 ;
  assign n11828 = ( n11712 & n11826 ) | ( n11712 & n11827 ) | ( n11826 & n11827 ) ;
  assign n11829 = n11732 & ~n11828 ;
  assign n11830 = ~n11731 & n11825 ;
  assign n11831 = ~n11709 & n11825 ;
  assign n11832 = ( ~n11712 & n11830 ) | ( ~n11712 & n11831 ) | ( n11830 & n11831 ) ;
  assign n11833 = n11829 | n11832 ;
  assign n11834 = n11620 | n11634 ;
  assign n11835 = ( n11634 & n11636 ) | ( n11634 & n11834 ) | ( n11636 & n11834 ) ;
  assign n11836 = n11605 | n11611 ;
  assign n11837 = ( n11605 & n11609 ) | ( n11605 & n11836 ) | ( n11609 & n11836 ) ;
  assign n11838 = n11835 | n11837 ;
  assign n11839 = n11835 & n11837 ;
  assign n11840 = n11838 & ~n11839 ;
  assign n11841 = n11683 | n11686 ;
  assign n11842 = ( n11683 & n11684 ) | ( n11683 & n11841 ) | ( n11684 & n11841 ) ;
  assign n11843 = n11840 | n11842 ;
  assign n11844 = n11840 & n11842 ;
  assign n11845 = n11843 & ~n11844 ;
  assign n11846 = n969 & n9829 ;
  assign n11847 = n360 & n9831 ;
  assign n11848 = n11846 | n11847 ;
  assign n11849 = n618 & n9272 ;
  assign n11850 = x59 & n11849 ;
  assign n11851 = ( x59 & ~n11848 ) | ( x59 & n11850 ) | ( ~n11848 & n11850 ) ;
  assign n11852 = x9 & n11851 ;
  assign n11853 = n11848 | n11849 ;
  assign n11854 = x10 & x58 ;
  assign n11855 = x11 & x57 ;
  assign n11856 = ( ~n11849 & n11854 ) | ( ~n11849 & n11855 ) | ( n11854 & n11855 ) ;
  assign n11857 = n11854 & n11855 ;
  assign n11858 = ( ~n11848 & n11856 ) | ( ~n11848 & n11857 ) | ( n11856 & n11857 ) ;
  assign n11859 = ~n11853 & n11858 ;
  assign n11860 = n11852 | n11859 ;
  assign n11861 = n2075 & n4350 ;
  assign n11862 = n2372 & n5813 ;
  assign n11863 = n11861 | n11862 ;
  assign n11864 = n2369 & n4555 ;
  assign n11865 = x41 & n11864 ;
  assign n11866 = ( x41 & ~n11863 ) | ( x41 & n11865 ) | ( ~n11863 & n11865 ) ;
  assign n11867 = x27 & n11866 ;
  assign n11868 = n11863 | n11864 ;
  assign n11869 = x28 & x40 ;
  assign n11870 = x29 & x39 ;
  assign n11871 = ( ~n11864 & n11869 ) | ( ~n11864 & n11870 ) | ( n11869 & n11870 ) ;
  assign n11872 = n11869 & n11870 ;
  assign n11873 = ( ~n11863 & n11871 ) | ( ~n11863 & n11872 ) | ( n11871 & n11872 ) ;
  assign n11874 = ~n11868 & n11873 ;
  assign n11875 = n11867 | n11874 ;
  assign n11876 = n11860 & n11875 ;
  assign n11877 = n11860 & ~n11876 ;
  assign n11878 = n11875 & ~n11876 ;
  assign n11879 = n11877 | n11878 ;
  assign n11880 = x5 & x63 ;
  assign n11881 = x6 & x62 ;
  assign n11882 = n11880 | n11881 ;
  assign n11883 = n204 & n10561 ;
  assign n11884 = x21 & x47 ;
  assign n11885 = ~n11883 & n11884 ;
  assign n11886 = n11882 | n11883 ;
  assign n11887 = ( n11883 & n11885 ) | ( n11883 & n11886 ) | ( n11885 & n11886 ) ;
  assign n11888 = n11882 & ~n11887 ;
  assign n11889 = ( ~n11882 & n11883 ) | ( ~n11882 & n11884 ) | ( n11883 & n11884 ) ;
  assign n11890 = n11884 & n11889 ;
  assign n11891 = n11888 | n11890 ;
  assign n11892 = ~n11879 & n11891 ;
  assign n11893 = n11879 & ~n11891 ;
  assign n11894 = n11892 | n11893 ;
  assign n11895 = x18 & x50 ;
  assign n11896 = x19 & x49 ;
  assign n11897 = n11895 | n11896 ;
  assign n11898 = n1077 & n6834 ;
  assign n11899 = n3129 & ~n11898 ;
  assign n11900 = n11897 | n11898 ;
  assign n11901 = ( n11898 & n11899 ) | ( n11898 & n11900 ) | ( n11899 & n11900 ) ;
  assign n11902 = n11897 & ~n11901 ;
  assign n11903 = n3129 & ~n11897 ;
  assign n11904 = ( n3129 & ~n11899 ) | ( n3129 & n11903 ) | ( ~n11899 & n11903 ) ;
  assign n11905 = n11902 | n11904 ;
  assign n11906 = n2546 & n3731 ;
  assign n11907 = n2965 & n4857 ;
  assign n11908 = n11906 | n11907 ;
  assign n11909 = n3770 & n4062 ;
  assign n11910 = x38 & n11909 ;
  assign n11911 = ( x38 & ~n11908 ) | ( x38 & n11910 ) | ( ~n11908 & n11910 ) ;
  assign n11912 = x30 & n11911 ;
  assign n11913 = n11908 | n11909 ;
  assign n11914 = x31 & x37 ;
  assign n11915 = x32 & x36 ;
  assign n11916 = ( ~n11909 & n11914 ) | ( ~n11909 & n11915 ) | ( n11914 & n11915 ) ;
  assign n11917 = n11914 & n11915 ;
  assign n11918 = ( ~n11908 & n11916 ) | ( ~n11908 & n11917 ) | ( n11916 & n11917 ) ;
  assign n11919 = ~n11913 & n11918 ;
  assign n11920 = n11912 | n11919 ;
  assign n11921 = n11905 & n11920 ;
  assign n11922 = n11905 & ~n11921 ;
  assign n11923 = n11920 & ~n11921 ;
  assign n11924 = n11922 | n11923 ;
  assign n11925 = x12 & x56 ;
  assign n11926 = x13 & x55 ;
  assign n11927 = ( ~n8437 & n11925 ) | ( ~n8437 & n11926 ) | ( n11925 & n11926 ) ;
  assign n11928 = n647 & n10013 ;
  assign n11929 = n11925 | n11926 ;
  assign n11930 = ( n8437 & n11928 ) | ( n8437 & n11929 ) | ( n11928 & n11929 ) ;
  assign n11931 = ( n8437 & n11927 ) | ( n8437 & ~n11930 ) | ( n11927 & ~n11930 ) ;
  assign n11932 = ~n11924 & n11931 ;
  assign n11933 = n11924 & ~n11931 ;
  assign n11934 = n11932 | n11933 ;
  assign n11935 = x52 & x54 ;
  assign n11936 = n790 & n11935 ;
  assign n11937 = n792 & n8355 ;
  assign n11938 = n11936 | n11937 ;
  assign n11939 = n795 & n8161 ;
  assign n11940 = x54 & n11939 ;
  assign n11941 = ( x54 & ~n11938 ) | ( x54 & n11940 ) | ( ~n11938 & n11940 ) ;
  assign n11942 = x14 & n11941 ;
  assign n11943 = n11938 | n11939 ;
  assign n11944 = x15 & x53 ;
  assign n11945 = x16 & x52 ;
  assign n11946 = ( ~n11939 & n11944 ) | ( ~n11939 & n11945 ) | ( n11944 & n11945 ) ;
  assign n11947 = n11944 & n11945 ;
  assign n11948 = ( ~n11938 & n11946 ) | ( ~n11938 & n11947 ) | ( n11946 & n11947 ) ;
  assign n11949 = ~n11943 & n11948 ;
  assign n11950 = n11942 | n11949 ;
  assign n11951 = x20 & x48 ;
  assign n11952 = n1932 & n5975 ;
  assign n11953 = x23 & x45 ;
  assign n11954 = x22 & x46 ;
  assign n11955 = n11953 | n11954 ;
  assign n11956 = ( n11951 & n11952 ) | ( n11951 & ~n11955 ) | ( n11952 & ~n11955 ) ;
  assign n11957 = n11951 & ~n11956 ;
  assign n11958 = ~n11952 & n11955 ;
  assign n11959 = n11951 | n11958 ;
  assign n11960 = ~n11957 & n11959 ;
  assign n11961 = n11950 & n11960 ;
  assign n11962 = n11950 & ~n11961 ;
  assign n11963 = n2340 & n4969 ;
  assign n11964 = n1912 & n5658 ;
  assign n11965 = n11963 | n11964 ;
  assign n11966 = n2511 & n5407 ;
  assign n11967 = x44 & n11966 ;
  assign n11968 = ( x44 & ~n11965 ) | ( x44 & n11967 ) | ( ~n11965 & n11967 ) ;
  assign n11969 = x24 & n11968 ;
  assign n11970 = n11965 | n11966 ;
  assign n11971 = x25 & x43 ;
  assign n11972 = x26 & x42 ;
  assign n11973 = ( ~n11966 & n11971 ) | ( ~n11966 & n11972 ) | ( n11971 & n11972 ) ;
  assign n11974 = n11971 & n11972 ;
  assign n11975 = ( ~n11965 & n11973 ) | ( ~n11965 & n11974 ) | ( n11973 & n11974 ) ;
  assign n11976 = ~n11970 & n11975 ;
  assign n11977 = n11969 | n11976 ;
  assign n11978 = ~n11950 & n11960 ;
  assign n11979 = n11977 & ~n11978 ;
  assign n11980 = ~n11962 & n11979 ;
  assign n11981 = ~n11977 & n11978 ;
  assign n11982 = ( n11962 & ~n11977 ) | ( n11962 & n11981 ) | ( ~n11977 & n11981 ) ;
  assign n11983 = n11980 | n11982 ;
  assign n11984 = n11934 & ~n11983 ;
  assign n11985 = ~n11934 & n11983 ;
  assign n11986 = n11984 | n11985 ;
  assign n11987 = n11894 & n11986 ;
  assign n11988 = n11894 | n11986 ;
  assign n11989 = ~n11987 & n11988 ;
  assign n11990 = n11845 & n11989 ;
  assign n11991 = n11845 | n11989 ;
  assign n11992 = ~n11990 & n11991 ;
  assign n11993 = n11330 | n11338 ;
  assign n11994 = ( n11689 & n11690 ) | ( n11689 & n11993 ) | ( n11690 & n11993 ) ;
  assign n11995 = n11992 & n11994 ;
  assign n11996 = n11992 | n11994 ;
  assign n11997 = ~n11995 & n11996 ;
  assign n11998 = ( n11571 & n11572 ) | ( n11571 & n11596 ) | ( n11572 & n11596 ) ;
  assign n11999 = n11997 | n11998 ;
  assign n12000 = n11997 & n11998 ;
  assign n12001 = n11999 & ~n12000 ;
  assign n12002 = n11651 | n11698 ;
  assign n12003 = ( n11651 & n11652 ) | ( n11651 & n12002 ) | ( n11652 & n12002 ) ;
  assign n12004 = n12001 & n12003 ;
  assign n12005 = n12001 | n12003 ;
  assign n12006 = ~n12004 & n12005 ;
  assign n12007 = n11832 | n12006 ;
  assign n12008 = n11829 | n12007 ;
  assign n12009 = ~n12006 & n12008 ;
  assign n12010 = ( ~n11833 & n12008 ) | ( ~n11833 & n12009 ) | ( n12008 & n12009 ) ;
  assign n12011 = n11599 & n11712 ;
  assign n12012 = n11599 | n11712 ;
  assign n12013 = ~n12011 & n12012 ;
  assign n12014 = n11706 & n12013 ;
  assign n12015 = n11703 | n12014 ;
  assign n12016 = ( n11728 & n12010 ) | ( n11728 & ~n12015 ) | ( n12010 & ~n12015 ) ;
  assign n12017 = ( ~n12010 & n12015 ) | ( ~n12010 & n12016 ) | ( n12015 & n12016 ) ;
  assign n12018 = ( ~n11728 & n12016 ) | ( ~n11728 & n12017 ) | ( n12016 & n12017 ) ;
  assign n12019 = n12010 | n12015 ;
  assign n12020 = n12010 & n12015 ;
  assign n12021 = n12019 | n12020 ;
  assign n12022 = ( n11721 & n12020 ) | ( n11721 & n12021 ) | ( n12020 & n12021 ) ;
  assign n12023 = ( n11727 & n12021 ) | ( n11727 & n12022 ) | ( n12021 & n12022 ) ;
  assign n12024 = n11989 | n11994 ;
  assign n12025 = ( n11845 & n11994 ) | ( n11845 & n12024 ) | ( n11994 & n12024 ) ;
  assign n12026 = ( n11990 & n11992 ) | ( n11990 & n12025 ) | ( n11992 & n12025 ) ;
  assign n12027 = n11780 | n11820 ;
  assign n12028 = ( n11820 & n11822 ) | ( n11820 & n12027 ) | ( n11822 & n12027 ) ;
  assign n12029 = n12026 | n12028 ;
  assign n12030 = n12026 & n12028 ;
  assign n12031 = n12029 & ~n12030 ;
  assign n12032 = n3334 & n7565 ;
  assign n12033 = n1077 & n7112 ;
  assign n12034 = n12032 | n12033 ;
  assign n12035 = n1020 & n7567 ;
  assign n12036 = x50 & n12035 ;
  assign n12037 = ( x50 & ~n12034 ) | ( x50 & n12036 ) | ( ~n12034 & n12036 ) ;
  assign n12038 = x19 & n12037 ;
  assign n12039 = n12034 | n12035 ;
  assign n12040 = x17 & x52 ;
  assign n12041 = x18 & x51 ;
  assign n12042 = ( ~n12035 & n12040 ) | ( ~n12035 & n12041 ) | ( n12040 & n12041 ) ;
  assign n12043 = n12040 & n12041 ;
  assign n12044 = ( ~n12034 & n12042 ) | ( ~n12034 & n12043 ) | ( n12042 & n12043 ) ;
  assign n12045 = ~n12039 & n12044 ;
  assign n12046 = n12038 | n12045 ;
  assign n12047 = n3280 & n4350 ;
  assign n12048 = n2369 & n5813 ;
  assign n12049 = n12047 | n12048 ;
  assign n12050 = n2709 & n4555 ;
  assign n12051 = x41 & n12050 ;
  assign n12052 = ( x41 & ~n12049 ) | ( x41 & n12051 ) | ( ~n12049 & n12051 ) ;
  assign n12053 = x28 & n12052 ;
  assign n12054 = n12049 | n12050 ;
  assign n12055 = x29 & x40 ;
  assign n12056 = x30 & x39 ;
  assign n12057 = ( ~n12050 & n12055 ) | ( ~n12050 & n12056 ) | ( n12055 & n12056 ) ;
  assign n12058 = n12055 & n12056 ;
  assign n12059 = ( ~n12049 & n12057 ) | ( ~n12049 & n12058 ) | ( n12057 & n12058 ) ;
  assign n12060 = ~n12054 & n12059 ;
  assign n12061 = n12053 | n12060 ;
  assign n12062 = n12046 & n12061 ;
  assign n12063 = n12046 & ~n12062 ;
  assign n12064 = n12061 & ~n12062 ;
  assign n12065 = n12063 | n12064 ;
  assign n12066 = n11485 | n11753 ;
  assign n12067 = ( n11753 & n11754 ) | ( n11753 & n12066 ) | ( n11754 & n12066 ) ;
  assign n12068 = n12065 | n12067 ;
  assign n12069 = n12065 & n12067 ;
  assign n12070 = n12068 & ~n12069 ;
  assign n12071 = n2683 & n3731 ;
  assign n12072 = n4062 & n4857 ;
  assign n12073 = n12071 | n12072 ;
  assign n12074 = n3321 & n3770 ;
  assign n12075 = x38 & n12074 ;
  assign n12076 = ( x38 & ~n12073 ) | ( x38 & n12075 ) | ( ~n12073 & n12075 ) ;
  assign n12077 = x31 & n12076 ;
  assign n12078 = n12073 | n12074 ;
  assign n12079 = x32 & x37 ;
  assign n12080 = ( n8090 & ~n12074 ) | ( n8090 & n12079 ) | ( ~n12074 & n12079 ) ;
  assign n12081 = n8090 & n12079 ;
  assign n12082 = ( ~n12073 & n12080 ) | ( ~n12073 & n12081 ) | ( n12080 & n12081 ) ;
  assign n12083 = ~n12078 & n12082 ;
  assign n12084 = n12077 | n12083 ;
  assign n12085 = ( x35 & x62 ) | ( x35 & ~n3483 ) | ( x62 & ~n3483 ) ;
  assign n12086 = x7 | x62 ;
  assign n12087 = ~x7 & x35 ;
  assign n12088 = ( n3483 & n12086 ) | ( n3483 & ~n12087 ) | ( n12086 & ~n12087 ) ;
  assign n12089 = ( ~x7 & x35 ) | ( ~x7 & x62 ) | ( x35 & x62 ) ;
  assign n12090 = ( x7 & n3483 ) | ( x7 & ~n12089 ) | ( n3483 & ~n12089 ) ;
  assign n12091 = ( n12085 & ~n12088 ) | ( n12085 & n12090 ) | ( ~n12088 & n12090 ) ;
  assign n12092 = n12084 & n12091 ;
  assign n12093 = n12084 & ~n12092 ;
  assign n12094 = n7496 & n10329 ;
  assign n12095 = n795 & n8355 ;
  assign n12096 = x20 & x54 ;
  assign n12097 = n10571 & n12096 ;
  assign n12098 = n12095 | n12097 ;
  assign n12099 = x54 & n12094 ;
  assign n12100 = ( x54 & ~n12098 ) | ( x54 & n12099 ) | ( ~n12098 & n12099 ) ;
  assign n12101 = x15 & n12100 ;
  assign n12102 = ( n7496 & n10329 ) | ( n7496 & ~n12098 ) | ( n10329 & ~n12098 ) ;
  assign n12103 = ( ~n12094 & n12101 ) | ( ~n12094 & n12102 ) | ( n12101 & n12102 ) ;
  assign n12104 = ~n12084 & n12091 ;
  assign n12105 = n12103 & n12104 ;
  assign n12106 = ( n12093 & n12103 ) | ( n12093 & n12105 ) | ( n12103 & n12105 ) ;
  assign n12107 = n12103 | n12104 ;
  assign n12108 = n12093 | n12107 ;
  assign n12109 = ~n12106 & n12108 ;
  assign n12110 = n12070 & n12109 ;
  assign n12111 = n12070 | n12109 ;
  assign n12112 = ~n12110 & n12111 ;
  assign n12113 = n11740 | n11743 ;
  assign n12114 = ( n11740 & n11745 ) | ( n11740 & n12113 ) | ( n11745 & n12113 ) ;
  assign n12115 = ( n11747 & n11748 ) | ( n11747 & n12114 ) | ( n11748 & n12114 ) ;
  assign n12116 = n12112 & n12115 ;
  assign n12117 = n12115 & ~n12116 ;
  assign n12118 = ( n12112 & ~n12116 ) | ( n12112 & n12117 ) | ( ~n12116 & n12117 ) ;
  assign n12119 = n11811 | n11814 ;
  assign n12120 = ( n11811 & n11813 ) | ( n11811 & n12119 ) | ( n11813 & n12119 ) ;
  assign n12121 = n12118 & n12120 ;
  assign n12122 = n12118 & ~n12121 ;
  assign n12123 = n249 & n9737 ;
  assign n12124 = n313 & n10367 ;
  assign n12125 = n12123 | n12124 ;
  assign n12126 = n360 & n10370 ;
  assign n12127 = x61 & n12126 ;
  assign n12128 = ( x61 & ~n12125 ) | ( x61 & n12127 ) | ( ~n12125 & n12127 ) ;
  assign n12129 = x8 & n12128 ;
  assign n12130 = n12125 | n12126 ;
  assign n12131 = x9 & x60 ;
  assign n12132 = x10 & x59 ;
  assign n12133 = ( ~n12126 & n12131 ) | ( ~n12126 & n12132 ) | ( n12131 & n12132 ) ;
  assign n12134 = n12131 & n12132 ;
  assign n12135 = ( ~n12125 & n12133 ) | ( ~n12125 & n12134 ) | ( n12133 & n12134 ) ;
  assign n12136 = ~n12130 & n12135 ;
  assign n12137 = n12129 | n12136 ;
  assign n12138 = n1557 & n8407 ;
  assign n12139 = n1686 & n5975 ;
  assign n12140 = n12138 | n12139 ;
  assign n12141 = n1912 & n6093 ;
  assign n12142 = x46 & n12141 ;
  assign n12143 = ( x46 & ~n12140 ) | ( x46 & n12142 ) | ( ~n12140 & n12142 ) ;
  assign n12144 = x23 & n12143 ;
  assign n12145 = n12140 | n12141 ;
  assign n12146 = x24 & x45 ;
  assign n12147 = x25 & x44 ;
  assign n12148 = ( ~n12141 & n12146 ) | ( ~n12141 & n12147 ) | ( n12146 & n12147 ) ;
  assign n12149 = n12146 & n12147 ;
  assign n12150 = ( ~n12140 & n12148 ) | ( ~n12140 & n12149 ) | ( n12148 & n12149 ) ;
  assign n12151 = ~n12145 & n12150 ;
  assign n12152 = n12144 | n12151 ;
  assign n12153 = n12137 & n12152 ;
  assign n12154 = n12137 & ~n12153 ;
  assign n12155 = n12152 & ~n12153 ;
  assign n12156 = n12154 | n12155 ;
  assign n12157 = x26 & x43 ;
  assign n12158 = x27 & x42 ;
  assign n12159 = n12157 | n12158 ;
  assign n12160 = n2267 & n5407 ;
  assign n12161 = x6 & x63 ;
  assign n12162 = ~n12160 & n12161 ;
  assign n12163 = n12159 | n12160 ;
  assign n12164 = ( n12160 & n12162 ) | ( n12160 & n12163 ) | ( n12162 & n12163 ) ;
  assign n12165 = n12159 & ~n12164 ;
  assign n12166 = ( ~n12159 & n12160 ) | ( ~n12159 & n12161 ) | ( n12160 & n12161 ) ;
  assign n12167 = n12161 & n12166 ;
  assign n12168 = n12165 | n12167 ;
  assign n12169 = ~n12156 & n12168 ;
  assign n12170 = n12156 & ~n12168 ;
  assign n12171 = n12169 | n12170 ;
  assign n12172 = n11785 | n11790 ;
  assign n12173 = n12171 | n12172 ;
  assign n12174 = n12171 & n12172 ;
  assign n12175 = n12173 & ~n12174 ;
  assign n12176 = n720 & n8708 ;
  assign n12177 = n490 & n9272 ;
  assign n12178 = n12176 | n12177 ;
  assign n12179 = n647 & n8903 ;
  assign n12180 = x58 & n12179 ;
  assign n12181 = ( x58 & ~n12178 ) | ( x58 & n12180 ) | ( ~n12178 & n12180 ) ;
  assign n12182 = x11 & n12181 ;
  assign n12183 = n12178 | n12179 ;
  assign n12184 = x12 & x57 ;
  assign n12185 = x13 & x56 ;
  assign n12186 = ( ~n12179 & n12184 ) | ( ~n12179 & n12185 ) | ( n12184 & n12185 ) ;
  assign n12187 = n12184 & n12185 ;
  assign n12188 = ( ~n12178 & n12186 ) | ( ~n12178 & n12187 ) | ( n12186 & n12187 ) ;
  assign n12189 = ~n12183 & n12188 ;
  assign n12190 = n12182 | n12189 ;
  assign n12191 = n11530 | n11792 ;
  assign n12192 = ( n11792 & n11796 ) | ( n11792 & n12191 ) | ( n11796 & n12191 ) ;
  assign n12193 = n12190 & ~n12192 ;
  assign n12194 = ~n12190 & n12192 ;
  assign n12195 = n12193 | n12194 ;
  assign n12196 = x21 & x48 ;
  assign n12197 = x22 & x47 ;
  assign n12198 = n12196 | n12197 ;
  assign n12199 = n1585 & n6762 ;
  assign n12200 = x14 & x55 ;
  assign n12201 = ~n12199 & n12200 ;
  assign n12202 = n12198 | n12199 ;
  assign n12203 = ( n12199 & n12201 ) | ( n12199 & n12202 ) | ( n12201 & n12202 ) ;
  assign n12204 = n12198 & ~n12203 ;
  assign n12205 = ( ~n12198 & n12199 ) | ( ~n12198 & n12200 ) | ( n12199 & n12200 ) ;
  assign n12206 = n12200 & n12205 ;
  assign n12207 = n12204 | n12206 ;
  assign n12208 = n12195 & n12207 ;
  assign n12209 = n12195 | n12207 ;
  assign n12210 = ~n12208 & n12209 ;
  assign n12211 = n12175 & n12210 ;
  assign n12212 = n12175 | n12210 ;
  assign n12213 = ~n12211 & n12212 ;
  assign n12214 = ~n12118 & n12120 ;
  assign n12215 = n12213 & ~n12214 ;
  assign n12216 = ~n12122 & n12215 ;
  assign n12217 = ~n12213 & n12214 ;
  assign n12218 = ( n12122 & ~n12213 ) | ( n12122 & n12217 ) | ( ~n12213 & n12217 ) ;
  assign n12219 = n12216 | n12218 ;
  assign n12220 = n12031 & n12219 ;
  assign n12221 = n12031 | n12219 ;
  assign n12222 = ~n12220 & n12221 ;
  assign n12223 = n11765 | n11770 ;
  assign n12224 = n8437 & n11925 ;
  assign n12225 = n11928 | n12224 ;
  assign n12226 = n8437 & n11926 ;
  assign n12227 = n12225 | n12226 ;
  assign n12228 = n11970 | n12227 ;
  assign n12229 = n11970 & n12227 ;
  assign n12230 = n12228 & ~n12229 ;
  assign n12231 = n11868 | n12230 ;
  assign n12232 = n11868 & n12230 ;
  assign n12233 = n12231 & ~n12232 ;
  assign n12234 = ( n11558 & n11733 ) | ( n11558 & n11734 ) | ( n11733 & n11734 ) ;
  assign n12235 = n11759 | n11761 ;
  assign n12236 = ( n11759 & n11760 ) | ( n11759 & n12235 ) | ( n11760 & n12235 ) ;
  assign n12237 = n12234 | n12236 ;
  assign n12238 = n12234 & n12236 ;
  assign n12239 = n12237 & ~n12238 ;
  assign n12240 = n12233 & n12239 ;
  assign n12241 = n12233 | n12239 ;
  assign n12242 = ~n12240 & n12241 ;
  assign n12243 = n12223 & n12242 ;
  assign n12244 = n12223 | n12242 ;
  assign n12245 = ~n12243 & n12244 ;
  assign n12246 = ( n11894 & n11934 ) | ( n11894 & n11983 ) | ( n11934 & n11983 ) ;
  assign n12247 = n12245 | n12246 ;
  assign n12248 = n12245 & n12246 ;
  assign n12249 = n12247 & ~n12248 ;
  assign n12250 = n11773 | n11777 ;
  assign n12251 = ( n11773 & n11775 ) | ( n11773 & n12250 ) | ( n11775 & n12250 ) ;
  assign n12252 = n12249 | n12251 ;
  assign n12253 = n12249 & n12251 ;
  assign n12254 = n12252 & ~n12253 ;
  assign n12255 = n11977 & n11978 ;
  assign n12256 = ( n11962 & n11977 ) | ( n11962 & n12255 ) | ( n11977 & n12255 ) ;
  assign n12257 = n11961 | n12256 ;
  assign n12258 = n11921 | n11931 ;
  assign n12259 = ( n11921 & n11924 ) | ( n11921 & n12258 ) | ( n11924 & n12258 ) ;
  assign n12260 = n12257 | n12259 ;
  assign n12261 = n12257 & n12259 ;
  assign n12262 = n12260 & ~n12261 ;
  assign n12263 = n11804 | n11807 ;
  assign n12264 = ( n11804 & n11805 ) | ( n11804 & n12263 ) | ( n11805 & n12263 ) ;
  assign n12265 = n12262 | n12264 ;
  assign n12266 = n12262 & n12264 ;
  assign n12267 = n12265 & ~n12266 ;
  assign n12268 = n11853 | n11887 ;
  assign n12269 = n11853 & n11887 ;
  assign n12270 = n12268 & ~n12269 ;
  assign n12271 = n11951 | n11952 ;
  assign n12272 = ( n11952 & ~n11956 ) | ( n11952 & n12271 ) | ( ~n11956 & n12271 ) ;
  assign n12273 = n12270 | n12272 ;
  assign n12274 = n12270 & n12272 ;
  assign n12275 = n12273 & ~n12274 ;
  assign n12276 = n11901 | n11913 ;
  assign n12277 = n11901 & n11913 ;
  assign n12278 = n12276 & ~n12277 ;
  assign n12279 = n11943 | n12278 ;
  assign n12280 = n11943 & n12278 ;
  assign n12281 = n12279 & ~n12280 ;
  assign n12282 = n11876 | n11891 ;
  assign n12283 = n12281 & n12282 ;
  assign n12284 = n11876 & n12281 ;
  assign n12285 = ( n11879 & n12283 ) | ( n11879 & n12284 ) | ( n12283 & n12284 ) ;
  assign n12286 = n12281 | n12282 ;
  assign n12287 = n11876 | n12281 ;
  assign n12288 = ( n11879 & n12286 ) | ( n11879 & n12287 ) | ( n12286 & n12287 ) ;
  assign n12289 = ~n12285 & n12288 ;
  assign n12290 = n12275 & n12289 ;
  assign n12291 = n12275 | n12289 ;
  assign n12292 = ~n12290 & n12291 ;
  assign n12293 = n12267 & n12292 ;
  assign n12294 = n12267 | n12292 ;
  assign n12295 = ~n12293 & n12294 ;
  assign n12296 = n11839 | n11842 ;
  assign n12297 = ( n11839 & n11840 ) | ( n11839 & n12296 ) | ( n11840 & n12296 ) ;
  assign n12298 = n12295 | n12297 ;
  assign n12299 = n12295 & n12297 ;
  assign n12300 = n12298 & ~n12299 ;
  assign n12301 = n12254 & n12300 ;
  assign n12302 = n12254 | n12300 ;
  assign n12303 = ~n12301 & n12302 ;
  assign n12304 = n12000 | n12003 ;
  assign n12305 = ( n12000 & n12001 ) | ( n12000 & n12304 ) | ( n12001 & n12304 ) ;
  assign n12306 = n12303 & n12305 ;
  assign n12307 = n12303 | n12305 ;
  assign n12308 = ~n12306 & n12307 ;
  assign n12309 = n12222 & n12308 ;
  assign n12310 = n12308 & ~n12309 ;
  assign n12311 = ( n12222 & ~n12309 ) | ( n12222 & n12310 ) | ( ~n12309 & n12310 ) ;
  assign n12312 = ~n11832 & n12006 ;
  assign n12313 = ~n11829 & n12312 ;
  assign n12314 = ( n11828 & n12006 ) | ( n11828 & ~n12313 ) | ( n12006 & ~n12313 ) ;
  assign n12315 = ( n12023 & n12311 ) | ( n12023 & ~n12314 ) | ( n12311 & ~n12314 ) ;
  assign n12316 = ( ~n12311 & n12314 ) | ( ~n12311 & n12315 ) | ( n12314 & n12315 ) ;
  assign n12317 = ( ~n12023 & n12315 ) | ( ~n12023 & n12316 ) | ( n12315 & n12316 ) ;
  assign n12368 = n12253 | n12300 ;
  assign n12369 = ( n12253 & n12254 ) | ( n12253 & n12368 ) | ( n12254 & n12368 ) ;
  assign n12318 = n12054 | n12164 ;
  assign n12319 = n12054 & n12164 ;
  assign n12320 = n12318 & ~n12319 ;
  assign n12321 = n12145 | n12320 ;
  assign n12322 = n12145 & n12320 ;
  assign n12323 = n12321 & ~n12322 ;
  assign n12324 = x62 & n4513 ;
  assign n12325 = n3483 & ~n12324 ;
  assign n12326 = x8 & x62 ;
  assign n12327 = n12324 | n12326 ;
  assign n12328 = n12325 | n12327 ;
  assign n12329 = n12324 & n12326 ;
  assign n12330 = ( n12325 & n12326 ) | ( n12325 & n12329 ) | ( n12326 & n12329 ) ;
  assign n12331 = n12078 & ~n12330 ;
  assign n12332 = n12328 | n12330 ;
  assign n12333 = ( n12330 & n12331 ) | ( n12330 & n12332 ) | ( n12331 & n12332 ) ;
  assign n12334 = n12328 & ~n12333 ;
  assign n12335 = n12078 & ~n12328 ;
  assign n12336 = ( n12078 & ~n12331 ) | ( n12078 & n12335 ) | ( ~n12331 & n12335 ) ;
  assign n12337 = n12334 | n12336 ;
  assign n12338 = n12323 & n12337 ;
  assign n12339 = n12323 & ~n12338 ;
  assign n12340 = n12337 & ~n12338 ;
  assign n12341 = n12339 | n12340 ;
  assign n12342 = n12062 | n12067 ;
  assign n12343 = ( n12062 & n12065 ) | ( n12062 & n12342 ) | ( n12065 & n12342 ) ;
  assign n12344 = n12341 | n12343 ;
  assign n12345 = n12341 & n12343 ;
  assign n12346 = n12344 & ~n12345 ;
  assign n12347 = ( n12190 & n12192 ) | ( n12190 & n12207 ) | ( n12192 & n12207 ) ;
  assign n12348 = n12153 | n12168 ;
  assign n12349 = n12347 | n12348 ;
  assign n12350 = n12153 | n12347 ;
  assign n12351 = ( n12156 & n12349 ) | ( n12156 & n12350 ) | ( n12349 & n12350 ) ;
  assign n12352 = n12347 & n12348 ;
  assign n12353 = n12153 & n12347 ;
  assign n12354 = ( n12156 & n12352 ) | ( n12156 & n12353 ) | ( n12352 & n12353 ) ;
  assign n12355 = n12351 & ~n12354 ;
  assign n12356 = n12092 | n12106 ;
  assign n12357 = n12355 | n12356 ;
  assign n12358 = n12355 & n12356 ;
  assign n12359 = n12357 & ~n12358 ;
  assign n12360 = n12110 & n12359 ;
  assign n12361 = ( n12116 & n12359 ) | ( n12116 & n12360 ) | ( n12359 & n12360 ) ;
  assign n12362 = n12110 | n12359 ;
  assign n12363 = n12116 | n12362 ;
  assign n12364 = ~n12361 & n12363 ;
  assign n12365 = n12346 | n12364 ;
  assign n12366 = n12346 & n12364 ;
  assign n12367 = n12365 & ~n12366 ;
  assign n12370 = n12367 & n12369 ;
  assign n12371 = n12369 & ~n12370 ;
  assign n12372 = n12094 | n12098 ;
  assign n12373 = n12039 | n12372 ;
  assign n12374 = n12039 & n12372 ;
  assign n12375 = n12373 & ~n12374 ;
  assign n12376 = n3321 & n4857 ;
  assign n12377 = x34 & x38 ;
  assign n12378 = n11915 & n12377 ;
  assign n12379 = n12376 | n12378 ;
  assign n12380 = n3770 & n4530 ;
  assign n12381 = x38 & n12380 ;
  assign n12382 = ( x38 & ~n12379 ) | ( x38 & n12381 ) | ( ~n12379 & n12381 ) ;
  assign n12383 = x32 & n12382 ;
  assign n12384 = n12379 | n12380 ;
  assign n12385 = x33 & x37 ;
  assign n12386 = ( n4914 & ~n12380 ) | ( n4914 & n12385 ) | ( ~n12380 & n12385 ) ;
  assign n12387 = n4914 & n12385 ;
  assign n12388 = ( ~n12379 & n12386 ) | ( ~n12379 & n12387 ) | ( n12386 & n12387 ) ;
  assign n12389 = ~n12384 & n12388 ;
  assign n12390 = n12383 | n12389 ;
  assign n12391 = n12375 & n12390 ;
  assign n12392 = n12375 & ~n12391 ;
  assign n12393 = n12390 & ~n12391 ;
  assign n12394 = n12392 | n12393 ;
  assign n12395 = n12233 | n12238 ;
  assign n12396 = ( n12238 & n12239 ) | ( n12238 & n12395 ) | ( n12239 & n12395 ) ;
  assign n12397 = n12394 & n12396 ;
  assign n12398 = n12394 | n12396 ;
  assign n12399 = ~n12397 & n12398 ;
  assign n12400 = n969 & n9737 ;
  assign n12401 = n360 & n10367 ;
  assign n12402 = n12400 | n12401 ;
  assign n12403 = n618 & n10370 ;
  assign n12404 = x61 & n12403 ;
  assign n12405 = ( x61 & ~n12402 ) | ( x61 & n12404 ) | ( ~n12402 & n12404 ) ;
  assign n12406 = x9 & n12405 ;
  assign n12407 = n12402 | n12403 ;
  assign n12408 = x10 & x60 ;
  assign n12409 = x11 & x59 ;
  assign n12410 = ( ~n12403 & n12408 ) | ( ~n12403 & n12409 ) | ( n12408 & n12409 ) ;
  assign n12411 = n12408 & n12409 ;
  assign n12412 = ( ~n12402 & n12410 ) | ( ~n12402 & n12411 ) | ( n12410 & n12411 ) ;
  assign n12413 = ~n12407 & n12412 ;
  assign n12414 = n12406 | n12413 ;
  assign n12415 = n1018 & n11935 ;
  assign n12416 = n1020 & n8161 ;
  assign n12417 = n12415 | n12416 ;
  assign n12418 = n1023 & n8355 ;
  assign n12419 = n8988 & n12418 ;
  assign n12420 = ( n8988 & ~n12417 ) | ( n8988 & n12419 ) | ( ~n12417 & n12419 ) ;
  assign n12421 = n12417 | n12418 ;
  assign n12422 = x16 & x54 ;
  assign n12423 = ( n9956 & ~n12418 ) | ( n9956 & n12422 ) | ( ~n12418 & n12422 ) ;
  assign n12424 = n9956 & n12422 ;
  assign n12425 = ( ~n12417 & n12423 ) | ( ~n12417 & n12424 ) | ( n12423 & n12424 ) ;
  assign n12426 = ~n12421 & n12425 ;
  assign n12427 = n12420 | n12426 ;
  assign n12428 = n12414 & n12427 ;
  assign n12429 = n12414 & ~n12428 ;
  assign n12430 = n647 & n9272 ;
  assign n12431 = x24 & x58 ;
  assign n12432 = n8791 & n12431 ;
  assign n12433 = n12430 | n12432 ;
  assign n12434 = n8942 & n11163 ;
  assign n12435 = x58 & n12434 ;
  assign n12436 = ( x58 & ~n12433 ) | ( x58 & n12435 ) | ( ~n12433 & n12435 ) ;
  assign n12437 = x12 & n12436 ;
  assign n12438 = n12433 | n12434 ;
  assign n12439 = x13 & x57 ;
  assign n12440 = ( n5590 & ~n12434 ) | ( n5590 & n12439 ) | ( ~n12434 & n12439 ) ;
  assign n12441 = n5590 & n12439 ;
  assign n12442 = ( ~n12433 & n12440 ) | ( ~n12433 & n12441 ) | ( n12440 & n12441 ) ;
  assign n12443 = ~n12438 & n12442 ;
  assign n12444 = n12437 | n12443 ;
  assign n12445 = ~n12414 & n12427 ;
  assign n12446 = n12444 & n12445 ;
  assign n12447 = ( n12429 & n12444 ) | ( n12429 & n12446 ) | ( n12444 & n12446 ) ;
  assign n12448 = n12444 | n12445 ;
  assign n12449 = n12429 | n12448 ;
  assign n12450 = ~n12447 & n12449 ;
  assign n12451 = n12399 & n12450 ;
  assign n12452 = n12399 | n12450 ;
  assign n12453 = ~n12451 & n12452 ;
  assign n12454 = n12243 | n12246 ;
  assign n12455 = ( n12243 & n12245 ) | ( n12243 & n12454 ) | ( n12245 & n12454 ) ;
  assign n12456 = n12453 & n12455 ;
  assign n12457 = n12453 | n12455 ;
  assign n12458 = ~n12456 & n12457 ;
  assign n12542 = n12275 | n12285 ;
  assign n12543 = ( n12285 & n12289 ) | ( n12285 & n12542 ) | ( n12289 & n12542 ) ;
  assign n12459 = n3595 & n4350 ;
  assign n12460 = n2709 & n5813 ;
  assign n12461 = n12459 | n12460 ;
  assign n12462 = n2965 & n4555 ;
  assign n12463 = x41 & n12462 ;
  assign n12464 = ( x41 & ~n12461 ) | ( x41 & n12463 ) | ( ~n12461 & n12463 ) ;
  assign n12465 = x29 & n12464 ;
  assign n12466 = n12461 | n12462 ;
  assign n12467 = x30 & x40 ;
  assign n12468 = x31 & x39 ;
  assign n12469 = ( ~n12462 & n12467 ) | ( ~n12462 & n12468 ) | ( n12467 & n12468 ) ;
  assign n12470 = n12467 & n12468 ;
  assign n12471 = ( ~n12461 & n12469 ) | ( ~n12461 & n12470 ) | ( n12469 & n12470 ) ;
  assign n12472 = ~n12466 & n12471 ;
  assign n12473 = n12465 | n12472 ;
  assign n12474 = x7 & x63 ;
  assign n12475 = x23 & x47 ;
  assign n12476 = n12474 | n12475 ;
  assign n12477 = x28 & x42 ;
  assign n12478 = ( n12474 & n12475 ) | ( n12474 & n12477 ) | ( n12475 & n12477 ) ;
  assign n12479 = n12476 & ~n12478 ;
  assign n12480 = n12474 & n12475 ;
  assign n12481 = n12477 & ~n12480 ;
  assign n12482 = ~n12476 & n12477 ;
  assign n12483 = ( n12477 & ~n12481 ) | ( n12477 & n12482 ) | ( ~n12481 & n12482 ) ;
  assign n12484 = n12479 | n12483 ;
  assign n12485 = n12473 & n12484 ;
  assign n12486 = n12473 & ~n12485 ;
  assign n12487 = ~n12473 & n12484 ;
  assign n12488 = n11943 | n12277 ;
  assign n12489 = ( n12277 & n12278 ) | ( n12277 & n12488 ) | ( n12278 & n12488 ) ;
  assign n12490 = n12487 | n12489 ;
  assign n12491 = n12486 | n12490 ;
  assign n12492 = n12487 & n12489 ;
  assign n12493 = ( n12486 & n12489 ) | ( n12486 & n12492 ) | ( n12489 & n12492 ) ;
  assign n12494 = n12491 & ~n12493 ;
  assign n12495 = n2724 & n5104 ;
  assign n12496 = n2511 & n6093 ;
  assign n12497 = n12495 | n12496 ;
  assign n12498 = n2267 & n5658 ;
  assign n12499 = x45 & n12498 ;
  assign n12500 = ( x45 & ~n12497 ) | ( x45 & n12499 ) | ( ~n12497 & n12499 ) ;
  assign n12501 = x25 & n12500 ;
  assign n12502 = n12497 | n12498 ;
  assign n12503 = x26 & x44 ;
  assign n12504 = x27 & x43 ;
  assign n12505 = ( ~n12498 & n12503 ) | ( ~n12498 & n12504 ) | ( n12503 & n12504 ) ;
  assign n12506 = n12503 & n12504 ;
  assign n12507 = ( ~n12497 & n12505 ) | ( ~n12497 & n12506 ) | ( n12505 & n12506 ) ;
  assign n12508 = ~n12502 & n12507 ;
  assign n12509 = n12501 | n12508 ;
  assign n12510 = x14 & x56 ;
  assign n12511 = x15 & x55 ;
  assign n12512 = n12510 | n12511 ;
  assign n12513 = n792 & n10013 ;
  assign n12514 = n12512 | n12513 ;
  assign n12515 = x22 & x48 ;
  assign n12516 = ( ~n12513 & n12514 ) | ( ~n12513 & n12515 ) | ( n12514 & n12515 ) ;
  assign n12517 = ( n12513 & n12514 ) | ( n12513 & ~n12515 ) | ( n12514 & ~n12515 ) ;
  assign n12518 = ( ~n12514 & n12516 ) | ( ~n12514 & n12517 ) | ( n12516 & n12517 ) ;
  assign n12519 = n12509 & n12518 ;
  assign n12520 = n12509 & ~n12519 ;
  assign n12521 = n1432 & n10866 ;
  assign n12522 = n1434 & n6834 ;
  assign n12523 = n12521 | n12522 ;
  assign n12524 = n1437 & n7112 ;
  assign n12525 = x49 & n12524 ;
  assign n12526 = ( x49 & ~n12523 ) | ( x49 & n12525 ) | ( ~n12523 & n12525 ) ;
  assign n12527 = x21 & n12526 ;
  assign n12528 = n12523 | n12524 ;
  assign n12529 = x19 & x51 ;
  assign n12530 = x20 & x50 ;
  assign n12531 = ( ~n12524 & n12529 ) | ( ~n12524 & n12530 ) | ( n12529 & n12530 ) ;
  assign n12532 = n12529 & n12530 ;
  assign n12533 = ( ~n12523 & n12531 ) | ( ~n12523 & n12532 ) | ( n12531 & n12532 ) ;
  assign n12534 = ~n12528 & n12533 ;
  assign n12535 = n12527 | n12534 ;
  assign n12536 = ~n12509 & n12518 ;
  assign n12537 = n12535 & ~n12536 ;
  assign n12538 = ~n12520 & n12537 ;
  assign n12539 = ~n12535 & n12536 ;
  assign n12540 = ( n12520 & ~n12535 ) | ( n12520 & n12539 ) | ( ~n12535 & n12539 ) ;
  assign n12541 = n12538 | n12540 ;
  assign n12544 = ( n12494 & ~n12541 ) | ( n12494 & n12543 ) | ( ~n12541 & n12543 ) ;
  assign n12545 = ( ~n12494 & n12541 ) | ( ~n12494 & n12543 ) | ( n12541 & n12543 ) ;
  assign n12546 = ( ~n12543 & n12544 ) | ( ~n12543 & n12545 ) | ( n12544 & n12545 ) ;
  assign n12547 = n12458 & n12546 ;
  assign n12548 = n12458 & ~n12547 ;
  assign n12549 = ~n12458 & n12546 ;
  assign n12550 = n12548 | n12549 ;
  assign n12551 = n12370 & n12550 ;
  assign n12552 = ~n12367 & n12549 ;
  assign n12553 = ( ~n12367 & n12548 ) | ( ~n12367 & n12552 ) | ( n12548 & n12552 ) ;
  assign n12554 = ( ~n12371 & n12551 ) | ( ~n12371 & n12553 ) | ( n12551 & n12553 ) ;
  assign n12555 = n12370 | n12550 ;
  assign n12556 = n12367 & ~n12549 ;
  assign n12557 = ~n12548 & n12556 ;
  assign n12558 = ( n12371 & ~n12555 ) | ( n12371 & n12557 ) | ( ~n12555 & n12557 ) ;
  assign n12559 = n12554 | n12558 ;
  assign n12599 = n12030 | n12219 ;
  assign n12600 = ( n12030 & n12031 ) | ( n12030 & n12599 ) | ( n12031 & n12599 ) ;
  assign n12576 = n12261 | n12264 ;
  assign n12577 = ( n12261 & n12262 ) | ( n12261 & n12576 ) | ( n12262 & n12576 ) ;
  assign n12560 = n12130 | n12183 ;
  assign n12561 = n12130 & n12183 ;
  assign n12562 = n12560 & ~n12561 ;
  assign n12563 = n12203 | n12562 ;
  assign n12564 = n12203 & n12562 ;
  assign n12565 = n12563 & ~n12564 ;
  assign n12566 = n12269 | n12272 ;
  assign n12567 = ( n12269 & n12270 ) | ( n12269 & n12566 ) | ( n12270 & n12566 ) ;
  assign n12568 = n11868 | n12229 ;
  assign n12569 = ( n12229 & n12230 ) | ( n12229 & n12568 ) | ( n12230 & n12568 ) ;
  assign n12570 = n12567 | n12569 ;
  assign n12571 = n12567 & n12569 ;
  assign n12572 = n12570 & ~n12571 ;
  assign n12573 = n12565 & n12572 ;
  assign n12574 = n12565 | n12572 ;
  assign n12575 = ~n12573 & n12574 ;
  assign n12578 = n12575 & n12577 ;
  assign n12579 = n12577 & ~n12578 ;
  assign n12580 = n12575 & ~n12577 ;
  assign n12581 = n12579 | n12580 ;
  assign n12582 = n12171 | n12210 ;
  assign n12583 = ( n12172 & n12210 ) | ( n12172 & n12582 ) | ( n12210 & n12582 ) ;
  assign n12584 = ( n12174 & n12175 ) | ( n12174 & n12583 ) | ( n12175 & n12583 ) ;
  assign n12585 = ~n12581 & n12584 ;
  assign n12586 = n12581 & ~n12584 ;
  assign n12587 = n12585 | n12586 ;
  assign n12588 = n12293 | n12297 ;
  assign n12589 = ( n12293 & n12295 ) | ( n12293 & n12588 ) | ( n12295 & n12588 ) ;
  assign n12590 = n12587 & n12589 ;
  assign n12591 = n12587 | n12589 ;
  assign n12592 = ~n12590 & n12591 ;
  assign n12593 = n12213 & n12214 ;
  assign n12594 = ( n12122 & n12213 ) | ( n12122 & n12593 ) | ( n12213 & n12593 ) ;
  assign n12595 = n12121 | n12594 ;
  assign n12596 = n12592 | n12595 ;
  assign n12597 = n12592 & n12595 ;
  assign n12598 = n12596 & ~n12597 ;
  assign n12601 = n12598 & n12600 ;
  assign n12602 = n12600 & ~n12601 ;
  assign n12603 = n12598 & ~n12600 ;
  assign n12604 = n12559 & n12603 ;
  assign n12605 = ( n12559 & n12602 ) | ( n12559 & n12604 ) | ( n12602 & n12604 ) ;
  assign n12606 = n12559 | n12603 ;
  assign n12607 = n12602 | n12606 ;
  assign n12608 = ~n12605 & n12607 ;
  assign n12609 = n12222 | n12306 ;
  assign n12610 = ( n12306 & n12308 ) | ( n12306 & n12609 ) | ( n12308 & n12609 ) ;
  assign n12611 = n12608 | n12610 ;
  assign n12612 = n12608 & n12610 ;
  assign n12613 = n12611 & ~n12612 ;
  assign n12614 = n12311 & n12314 ;
  assign n12615 = n12311 | n12314 ;
  assign n12616 = n12614 | n12615 ;
  assign n12617 = ( n12022 & n12614 ) | ( n12022 & n12616 ) | ( n12614 & n12616 ) ;
  assign n12618 = ( n12021 & n12614 ) | ( n12021 & n12616 ) | ( n12614 & n12616 ) ;
  assign n12619 = ( n11727 & n12617 ) | ( n11727 & n12618 ) | ( n12617 & n12618 ) ;
  assign n12620 = n12613 | n12619 ;
  assign n12621 = n12611 & n12618 ;
  assign n12622 = n12611 & n12616 ;
  assign n12623 = n12611 & n12614 ;
  assign n12624 = ( n12022 & n12622 ) | ( n12022 & n12623 ) | ( n12622 & n12623 ) ;
  assign n12625 = ( n11727 & n12621 ) | ( n11727 & n12624 ) | ( n12621 & n12624 ) ;
  assign n12626 = ~n12612 & n12625 ;
  assign n12627 = n12620 & ~n12626 ;
  assign n12628 = n12612 | n12624 ;
  assign n12629 = n12611 | n12612 ;
  assign n12630 = ( n12612 & n12618 ) | ( n12612 & n12629 ) | ( n12618 & n12629 ) ;
  assign n12631 = ( n11727 & n12628 ) | ( n11727 & n12630 ) | ( n12628 & n12630 ) ;
  assign n12632 = ( n12367 & ~n12370 ) | ( n12367 & n12371 ) | ( ~n12370 & n12371 ) ;
  assign n12633 = n12333 & n12374 ;
  assign n12634 = ( n12333 & n12391 ) | ( n12333 & n12633 ) | ( n12391 & n12633 ) ;
  assign n12635 = n12333 | n12374 ;
  assign n12636 = n12391 | n12635 ;
  assign n12637 = ~n12634 & n12636 ;
  assign n12638 = n12145 | n12319 ;
  assign n12639 = ( n12319 & n12320 ) | ( n12319 & n12638 ) | ( n12320 & n12638 ) ;
  assign n12640 = n12637 | n12639 ;
  assign n12641 = n12637 & n12639 ;
  assign n12642 = n12640 & ~n12641 ;
  assign n12643 = n12338 | n12343 ;
  assign n12644 = ( n12338 & n12341 ) | ( n12338 & n12643 ) | ( n12341 & n12643 ) ;
  assign n12645 = n12642 | n12644 ;
  assign n12646 = n12642 & n12644 ;
  assign n12647 = n12645 & ~n12646 ;
  assign n12648 = n12397 | n12450 ;
  assign n12649 = ( n12397 & n12399 ) | ( n12397 & n12648 ) | ( n12399 & n12648 ) ;
  assign n12650 = n12647 | n12649 ;
  assign n12651 = n12647 & n12649 ;
  assign n12652 = n12650 & ~n12651 ;
  assign n12653 = n12346 | n12361 ;
  assign n12654 = ( n12361 & n12364 ) | ( n12361 & n12653 ) | ( n12364 & n12653 ) ;
  assign n12655 = n12652 & n12654 ;
  assign n12656 = n12652 | n12654 ;
  assign n12657 = ~n12655 & n12656 ;
  assign n12658 = n12453 | n12546 ;
  assign n12659 = ( n12455 & n12546 ) | ( n12455 & n12658 ) | ( n12546 & n12658 ) ;
  assign n12660 = ( n12456 & n12458 ) | ( n12456 & n12659 ) | ( n12458 & n12659 ) ;
  assign n12661 = n12657 | n12660 ;
  assign n12662 = n12657 & n12660 ;
  assign n12663 = n12661 & ~n12662 ;
  assign n12664 = n12555 & n12663 ;
  assign n12665 = n12370 & n12663 ;
  assign n12666 = ( n12632 & n12664 ) | ( n12632 & n12665 ) | ( n12664 & n12665 ) ;
  assign n12667 = n12555 | n12663 ;
  assign n12668 = n12370 | n12663 ;
  assign n12669 = ( n12632 & n12667 ) | ( n12632 & n12668 ) | ( n12667 & n12668 ) ;
  assign n12670 = ~n12666 & n12669 ;
  assign n12671 = n12494 | n12541 ;
  assign n12672 = n12543 & n12671 ;
  assign n12673 = n12203 | n12561 ;
  assign n12674 = ( n12561 & n12562 ) | ( n12561 & n12673 ) | ( n12562 & n12673 ) ;
  assign n12675 = n12428 & n12674 ;
  assign n12676 = ( n12447 & n12674 ) | ( n12447 & n12675 ) | ( n12674 & n12675 ) ;
  assign n12677 = n12428 | n12674 ;
  assign n12678 = n12447 | n12677 ;
  assign n12679 = ~n12676 & n12678 ;
  assign n12680 = n12535 & n12536 ;
  assign n12681 = ( n12520 & n12535 ) | ( n12520 & n12680 ) | ( n12535 & n12680 ) ;
  assign n12682 = n12519 | n12681 ;
  assign n12683 = n12679 | n12682 ;
  assign n12684 = n12679 & n12682 ;
  assign n12685 = n12683 & ~n12684 ;
  assign n12686 = n12494 & n12541 ;
  assign n12687 = n12685 & n12686 ;
  assign n12688 = ( n12672 & n12685 ) | ( n12672 & n12687 ) | ( n12685 & n12687 ) ;
  assign n12689 = n12685 | n12686 ;
  assign n12690 = n12672 | n12689 ;
  assign n12691 = ~n12688 & n12690 ;
  assign n12692 = n12407 | n12438 ;
  assign n12693 = n12407 & n12438 ;
  assign n12694 = n12692 & ~n12693 ;
  assign n12695 = n12502 | n12694 ;
  assign n12696 = n12502 & n12694 ;
  assign n12697 = n12695 & ~n12696 ;
  assign n12698 = ~n12513 & n12515 ;
  assign n12699 = ( n12513 & n12514 ) | ( n12513 & n12698 ) | ( n12514 & n12698 ) ;
  assign n12700 = n12466 | n12699 ;
  assign n12701 = n12466 & n12699 ;
  assign n12702 = n12700 & ~n12701 ;
  assign n12703 = n12478 | n12702 ;
  assign n12704 = n12478 & n12702 ;
  assign n12705 = n12703 & ~n12704 ;
  assign n12706 = n12697 | n12705 ;
  assign n12707 = n12697 & n12705 ;
  assign n12708 = n12706 & ~n12707 ;
  assign n12709 = n12485 | n12493 ;
  assign n12710 = n12708 & n12709 ;
  assign n12711 = n12708 | n12709 ;
  assign n12712 = ~n12710 & n12711 ;
  assign n12713 = n12691 & n12712 ;
  assign n12714 = n12691 | n12712 ;
  assign n12715 = ~n12713 & n12714 ;
  assign n12716 = n12590 & n12715 ;
  assign n12717 = ( n12597 & n12715 ) | ( n12597 & n12716 ) | ( n12715 & n12716 ) ;
  assign n12718 = n12590 | n12715 ;
  assign n12719 = n12597 | n12718 ;
  assign n12720 = ~n12717 & n12719 ;
  assign n12721 = n1432 & n7565 ;
  assign n12722 = n1434 & n7112 ;
  assign n12723 = n12721 | n12722 ;
  assign n12724 = n1437 & n7567 ;
  assign n12725 = x50 & n12724 ;
  assign n12726 = ( x50 & ~n12723 ) | ( x50 & n12725 ) | ( ~n12723 & n12725 ) ;
  assign n12727 = x21 & n12726 ;
  assign n12728 = n12723 | n12724 ;
  assign n12729 = x19 & x52 ;
  assign n12730 = x20 & x51 ;
  assign n12731 = ( ~n12724 & n12729 ) | ( ~n12724 & n12730 ) | ( n12729 & n12730 ) ;
  assign n12732 = n12729 & n12730 ;
  assign n12733 = ( ~n12723 & n12731 ) | ( ~n12723 & n12732 ) | ( n12731 & n12732 ) ;
  assign n12734 = ~n12728 & n12733 ;
  assign n12735 = n12727 | n12734 ;
  assign n12736 = x9 & x62 ;
  assign n12737 = x36 | n12736 ;
  assign n12738 = x36 & x62 ;
  assign n12739 = ~x9 & x49 ;
  assign n12740 = ( x49 & ~n12738 ) | ( x49 & n12739 ) | ( ~n12738 & n12739 ) ;
  assign n12741 = ( x22 & x36 ) | ( x22 & n12736 ) | ( x36 & n12736 ) ;
  assign n12742 = x36 & n12736 ;
  assign n12743 = ( n12740 & n12741 ) | ( n12740 & n12742 ) | ( n12741 & n12742 ) ;
  assign n12744 = n12737 & ~n12743 ;
  assign n12745 = x22 & n12740 ;
  assign n12746 = ~x36 & x49 ;
  assign n12747 = ~n12736 & n12746 ;
  assign n12748 = x22 & n12747 ;
  assign n12749 = x22 & x49 ;
  assign n12750 = ( ~n12745 & n12748 ) | ( ~n12745 & n12749 ) | ( n12748 & n12749 ) ;
  assign n12751 = n12744 | n12750 ;
  assign n12752 = n12735 & n12751 ;
  assign n12753 = n12735 & ~n12752 ;
  assign n12754 = x34 & x37 ;
  assign n12755 = ( ~n4078 & n4855 ) | ( ~n4078 & n12754 ) | ( n4855 & n12754 ) ;
  assign n12756 = n4530 & n4857 ;
  assign n12757 = n4855 | n12754 ;
  assign n12758 = ( n4078 & n12756 ) | ( n4078 & n12757 ) | ( n12756 & n12757 ) ;
  assign n12759 = ( n4078 & n12755 ) | ( n4078 & ~n12758 ) | ( n12755 & ~n12758 ) ;
  assign n12760 = ~n12751 & n12759 ;
  assign n12761 = ( n12735 & n12759 ) | ( n12735 & n12760 ) | ( n12759 & n12760 ) ;
  assign n12762 = ~n12753 & n12761 ;
  assign n12763 = n12751 & ~n12759 ;
  assign n12764 = ~n12735 & n12763 ;
  assign n12765 = ( n12753 & ~n12759 ) | ( n12753 & n12764 ) | ( ~n12759 & n12764 ) ;
  assign n12766 = n12762 | n12765 ;
  assign n12767 = n12384 | n12421 ;
  assign n12768 = n12384 & n12421 ;
  assign n12769 = n12767 & ~n12768 ;
  assign n12770 = x60 & x63 ;
  assign n12771 = n894 & n12770 ;
  assign n12772 = n618 & n10367 ;
  assign n12773 = n12771 | n12772 ;
  assign n12774 = n249 & n10856 ;
  assign n12775 = x60 & n12774 ;
  assign n12776 = ( x60 & ~n12773 ) | ( x60 & n12775 ) | ( ~n12773 & n12775 ) ;
  assign n12777 = x11 & n12776 ;
  assign n12778 = n12773 | n12774 ;
  assign n12779 = x8 & x63 ;
  assign n12780 = x10 & x61 ;
  assign n12781 = ( ~n12774 & n12779 ) | ( ~n12774 & n12780 ) | ( n12779 & n12780 ) ;
  assign n12782 = n12779 & n12780 ;
  assign n12783 = ( ~n12773 & n12781 ) | ( ~n12773 & n12782 ) | ( n12781 & n12782 ) ;
  assign n12784 = ~n12778 & n12783 ;
  assign n12785 = n12777 | n12784 ;
  assign n12786 = n12769 & n12785 ;
  assign n12787 = n12769 & ~n12786 ;
  assign n12788 = n12785 & ~n12786 ;
  assign n12789 = n12787 | n12788 ;
  assign n12790 = n12565 | n12571 ;
  assign n12791 = ( n12571 & n12572 ) | ( n12571 & n12790 ) | ( n12572 & n12790 ) ;
  assign n12792 = n12789 & n12791 ;
  assign n12793 = n12789 | n12791 ;
  assign n12794 = ~n12792 & n12793 ;
  assign n12795 = n12766 & n12794 ;
  assign n12796 = n12766 | n12794 ;
  assign n12797 = ~n12795 & n12796 ;
  assign n12798 = n12578 | n12584 ;
  assign n12799 = ( n12578 & n12581 ) | ( n12578 & n12798 ) | ( n12581 & n12798 ) ;
  assign n12800 = n12797 & n12799 ;
  assign n12801 = n12797 | n12799 ;
  assign n12802 = ~n12800 & n12801 ;
  assign n12803 = n2075 & n4969 ;
  assign n12804 = n2372 & n5658 ;
  assign n12805 = n12803 | n12804 ;
  assign n12806 = n2369 & n5407 ;
  assign n12807 = x44 & n12806 ;
  assign n12808 = ( x44 & ~n12805 ) | ( x44 & n12807 ) | ( ~n12805 & n12807 ) ;
  assign n12809 = x27 & n12808 ;
  assign n12810 = n12805 | n12806 ;
  assign n12811 = x28 & x43 ;
  assign n12812 = x29 & x42 ;
  assign n12813 = ( ~n12806 & n12811 ) | ( ~n12806 & n12812 ) | ( n12811 & n12812 ) ;
  assign n12814 = n12811 & n12812 ;
  assign n12815 = ( ~n12805 & n12813 ) | ( ~n12805 & n12814 ) | ( n12813 & n12814 ) ;
  assign n12816 = ~n12810 & n12815 ;
  assign n12817 = n12809 | n12816 ;
  assign n12818 = n2546 & n4350 ;
  assign n12819 = n2965 & n5813 ;
  assign n12820 = n12818 | n12819 ;
  assign n12821 = n4062 & n4555 ;
  assign n12822 = x41 & n12821 ;
  assign n12823 = ( x41 & ~n12820 ) | ( x41 & n12822 ) | ( ~n12820 & n12822 ) ;
  assign n12824 = x30 & n12823 ;
  assign n12825 = n12820 | n12821 ;
  assign n12826 = x31 & x40 ;
  assign n12827 = x32 & x39 ;
  assign n12828 = ( ~n12821 & n12826 ) | ( ~n12821 & n12827 ) | ( n12826 & n12827 ) ;
  assign n12829 = n12826 & n12827 ;
  assign n12830 = ( ~n12820 & n12828 ) | ( ~n12820 & n12829 ) | ( n12828 & n12829 ) ;
  assign n12831 = ~n12825 & n12830 ;
  assign n12832 = n12824 | n12831 ;
  assign n12833 = n12817 & n12832 ;
  assign n12834 = n12817 & ~n12833 ;
  assign n12835 = n12832 & ~n12833 ;
  assign n12836 = n12834 | n12835 ;
  assign n12837 = x17 & x54 ;
  assign n12838 = n9413 | n12837 ;
  assign n12839 = n1020 & n8355 ;
  assign n12840 = x23 & x48 ;
  assign n12841 = ~n12839 & n12840 ;
  assign n12842 = n12838 | n12839 ;
  assign n12843 = ( n12839 & n12841 ) | ( n12839 & n12842 ) | ( n12841 & n12842 ) ;
  assign n12844 = n12838 & ~n12843 ;
  assign n12845 = ( ~n12838 & n12839 ) | ( ~n12838 & n12840 ) | ( n12839 & n12840 ) ;
  assign n12846 = n12840 & n12845 ;
  assign n12847 = n12844 | n12846 ;
  assign n12848 = ~n12836 & n12847 ;
  assign n12849 = n12836 & ~n12847 ;
  assign n12850 = n12848 | n12849 ;
  assign n12851 = n647 & n9831 ;
  assign n12852 = x13 & x58 ;
  assign n12853 = x12 & x59 ;
  assign n12854 = n12852 | n12853 ;
  assign n12855 = ~n12851 & n12854 ;
  assign n12856 = n12528 & n12855 ;
  assign n12857 = n12528 & ~n12856 ;
  assign n12858 = ~n12528 & n12855 ;
  assign n12859 = n12857 | n12858 ;
  assign n12860 = x55 & x57 ;
  assign n12861 = n790 & n12860 ;
  assign n12862 = n792 & n8903 ;
  assign n12863 = n12861 | n12862 ;
  assign n12864 = n795 & n10013 ;
  assign n12865 = x57 & n12864 ;
  assign n12866 = ( x57 & ~n12863 ) | ( x57 & n12865 ) | ( ~n12863 & n12865 ) ;
  assign n12867 = x14 & n12866 ;
  assign n12868 = n12863 | n12864 ;
  assign n12869 = x15 & x56 ;
  assign n12870 = x16 & x55 ;
  assign n12871 = ( ~n12864 & n12869 ) | ( ~n12864 & n12870 ) | ( n12869 & n12870 ) ;
  assign n12872 = n12869 & n12870 ;
  assign n12873 = ( ~n12863 & n12871 ) | ( ~n12863 & n12872 ) | ( n12871 & n12872 ) ;
  assign n12874 = ~n12868 & n12873 ;
  assign n12875 = n12867 | n12874 ;
  assign n12876 = n2340 & n5610 ;
  assign n12877 = n1912 & n6147 ;
  assign n12878 = n12876 | n12877 ;
  assign n12879 = n2511 & n5975 ;
  assign n12880 = x47 & n12879 ;
  assign n12881 = ( x47 & ~n12878 ) | ( x47 & n12880 ) | ( ~n12878 & n12880 ) ;
  assign n12882 = x24 & n12881 ;
  assign n12883 = n12878 | n12879 ;
  assign n12884 = x26 & x45 ;
  assign n12885 = ( n11451 & ~n12879 ) | ( n11451 & n12884 ) | ( ~n12879 & n12884 ) ;
  assign n12886 = n11451 & n12884 ;
  assign n12887 = ( ~n12878 & n12885 ) | ( ~n12878 & n12886 ) | ( n12885 & n12886 ) ;
  assign n12888 = ~n12883 & n12887 ;
  assign n12889 = n12882 | n12888 ;
  assign n12890 = n12875 & n12889 ;
  assign n12891 = n12875 & ~n12890 ;
  assign n12892 = n12889 & ~n12890 ;
  assign n12893 = n12891 | n12892 ;
  assign n12894 = n12859 & ~n12893 ;
  assign n12895 = ~n12859 & n12893 ;
  assign n12896 = n12894 | n12895 ;
  assign n12897 = n12850 & n12896 ;
  assign n12898 = n12850 | n12896 ;
  assign n12899 = ~n12897 & n12898 ;
  assign n12900 = n12354 | n12356 ;
  assign n12901 = ( n12354 & n12355 ) | ( n12354 & n12900 ) | ( n12355 & n12900 ) ;
  assign n12902 = n12899 & n12901 ;
  assign n12903 = n12899 | n12901 ;
  assign n12904 = ~n12902 & n12903 ;
  assign n12905 = n12802 & n12904 ;
  assign n12906 = n12802 | n12904 ;
  assign n12907 = ~n12905 & n12906 ;
  assign n12908 = n12720 & n12907 ;
  assign n12909 = n12720 | n12907 ;
  assign n12910 = ~n12908 & n12909 ;
  assign n12911 = n12670 | n12910 ;
  assign n12912 = n12670 & n12910 ;
  assign n12913 = n12911 & ~n12912 ;
  assign n12914 = n12601 | n12605 ;
  assign n12915 = ( n12631 & n12913 ) | ( n12631 & ~n12914 ) | ( n12913 & ~n12914 ) ;
  assign n12916 = ( ~n12913 & n12914 ) | ( ~n12913 & n12915 ) | ( n12914 & n12915 ) ;
  assign n12917 = ( ~n12631 & n12915 ) | ( ~n12631 & n12916 ) | ( n12915 & n12916 ) ;
  assign n12918 = n12707 | n12710 ;
  assign n12919 = n3595 & n5107 ;
  assign n12920 = n2709 & n5407 ;
  assign n12921 = n12919 | n12920 ;
  assign n12922 = n2965 & n5710 ;
  assign n12923 = x43 & n12922 ;
  assign n12924 = ( x43 & ~n12921 ) | ( x43 & n12923 ) | ( ~n12921 & n12923 ) ;
  assign n12925 = x29 & n12924 ;
  assign n12926 = n12921 | n12922 ;
  assign n12927 = x30 & x42 ;
  assign n12928 = ( n5328 & ~n12922 ) | ( n5328 & n12927 ) | ( ~n12922 & n12927 ) ;
  assign n12929 = n5328 & n12927 ;
  assign n12930 = ( ~n12921 & n12928 ) | ( ~n12921 & n12929 ) | ( n12928 & n12929 ) ;
  assign n12931 = ~n12926 & n12930 ;
  assign n12932 = n12925 | n12931 ;
  assign n12933 = n12768 & n12932 ;
  assign n12934 = ( n12786 & n12932 ) | ( n12786 & n12933 ) | ( n12932 & n12933 ) ;
  assign n12935 = n12768 | n12932 ;
  assign n12936 = n12786 | n12935 ;
  assign n12937 = ~n12934 & n12936 ;
  assign n12938 = n12478 | n12701 ;
  assign n12939 = ( n12701 & n12702 ) | ( n12701 & n12938 ) | ( n12702 & n12938 ) ;
  assign n12940 = n12937 | n12939 ;
  assign n12941 = n12937 & n12939 ;
  assign n12942 = n12940 & ~n12941 ;
  assign n12943 = n12918 & n12942 ;
  assign n12944 = n12918 | n12942 ;
  assign n12945 = ~n12943 & n12944 ;
  assign n12946 = n12766 | n12792 ;
  assign n12947 = ( n12792 & n12794 ) | ( n12792 & n12946 ) | ( n12794 & n12946 ) ;
  assign n12948 = n12945 | n12947 ;
  assign n12949 = n12945 & n12947 ;
  assign n12950 = n12948 & ~n12949 ;
  assign n12951 = n12685 | n12712 ;
  assign n12952 = n12672 | n12712 ;
  assign n12953 = ( n12687 & n12951 ) | ( n12687 & n12952 ) | ( n12951 & n12952 ) ;
  assign n12954 = ( n12688 & n12691 ) | ( n12688 & n12953 ) | ( n12691 & n12953 ) ;
  assign n12955 = n12950 & n12954 ;
  assign n12956 = n12950 | n12954 ;
  assign n12957 = ~n12955 & n12956 ;
  assign n12958 = ( n12797 & n12799 ) | ( n12797 & n12904 ) | ( n12799 & n12904 ) ;
  assign n12959 = n12957 | n12958 ;
  assign n12960 = n12957 & n12958 ;
  assign n12961 = n12959 & ~n12960 ;
  assign n12962 = n12717 | n12907 ;
  assign n12963 = ( n12717 & n12720 ) | ( n12717 & n12962 ) | ( n12720 & n12962 ) ;
  assign n12964 = n12961 & n12963 ;
  assign n12965 = n12961 | n12963 ;
  assign n12966 = ~n12964 & n12965 ;
  assign n12967 = n12833 | n12847 ;
  assign n12968 = n12502 | n12693 ;
  assign n12969 = ( n12693 & n12694 ) | ( n12693 & n12968 ) | ( n12694 & n12968 ) ;
  assign n12970 = n12967 & n12969 ;
  assign n12971 = n12833 & n12969 ;
  assign n12972 = ( n12836 & n12970 ) | ( n12836 & n12971 ) | ( n12970 & n12971 ) ;
  assign n12973 = n12967 | n12969 ;
  assign n12974 = n12833 | n12969 ;
  assign n12975 = ( n12836 & n12973 ) | ( n12836 & n12974 ) | ( n12973 & n12974 ) ;
  assign n12976 = ~n12972 & n12975 ;
  assign n12977 = n12751 & n12759 ;
  assign n12978 = ~n12735 & n12977 ;
  assign n12979 = n12752 | n12978 ;
  assign n12980 = n12752 | n12759 ;
  assign n12981 = ( n12753 & n12979 ) | ( n12753 & n12980 ) | ( n12979 & n12980 ) ;
  assign n12982 = n12976 | n12981 ;
  assign n12983 = n12976 & n12981 ;
  assign n12984 = n12982 & ~n12983 ;
  assign n12985 = n12897 | n12901 ;
  assign n12986 = ( n12897 & n12899 ) | ( n12897 & n12985 ) | ( n12899 & n12985 ) ;
  assign n12987 = n12984 | n12986 ;
  assign n12988 = n12984 & n12986 ;
  assign n12989 = n12987 & ~n12988 ;
  assign n12990 = n12810 | n12843 ;
  assign n12991 = n12810 & n12843 ;
  assign n12992 = n12990 & ~n12991 ;
  assign n12993 = n12825 | n12992 ;
  assign n12994 = n12825 & n12992 ;
  assign n12995 = n12993 & ~n12994 ;
  assign n12996 = n4078 & n4855 ;
  assign n12997 = n12756 | n12996 ;
  assign n12998 = n4078 & n12754 ;
  assign n12999 = n12997 | n12998 ;
  assign n13000 = n12743 | n12999 ;
  assign n13001 = n12743 & n12999 ;
  assign n13002 = n13000 & ~n13001 ;
  assign n13003 = n12728 | n13002 ;
  assign n13004 = n12728 & n13002 ;
  assign n13005 = n13003 & ~n13004 ;
  assign n13006 = n12995 & n13005 ;
  assign n13007 = n12995 | n13005 ;
  assign n13008 = ~n13006 & n13007 ;
  assign n13009 = ( n12859 & n12875 ) | ( n12859 & n12889 ) | ( n12875 & n12889 ) ;
  assign n13010 = n13008 & n13009 ;
  assign n13011 = n13008 | n13009 ;
  assign n13012 = ~n13010 & n13011 ;
  assign n13013 = n12989 & n13012 ;
  assign n13014 = n12989 | n13012 ;
  assign n13015 = ~n13013 & n13014 ;
  assign n13016 = n12655 | n12660 ;
  assign n13017 = ( n12655 & n12657 ) | ( n12655 & n13016 ) | ( n12657 & n13016 ) ;
  assign n13018 = n13015 | n13017 ;
  assign n13019 = ( n12655 & n12660 ) | ( n12655 & n13015 ) | ( n12660 & n13015 ) ;
  assign n13020 = n12655 & n13015 ;
  assign n13021 = ( n12657 & n13019 ) | ( n12657 & n13020 ) | ( n13019 & n13020 ) ;
  assign n13022 = n13018 & ~n13021 ;
  assign n13023 = x21 & x51 ;
  assign n13024 = x22 & x50 ;
  assign n13025 = n13023 | n13024 ;
  assign n13026 = n1585 & n7112 ;
  assign n13027 = n5417 & ~n13026 ;
  assign n13028 = n13025 | n13026 ;
  assign n13029 = ( n13026 & n13027 ) | ( n13026 & n13028 ) | ( n13027 & n13028 ) ;
  assign n13030 = n13025 & ~n13029 ;
  assign n13031 = n5417 & ~n13025 ;
  assign n13032 = ( n5417 & ~n13027 ) | ( n5417 & n13031 ) | ( ~n13027 & n13031 ) ;
  assign n13033 = n13030 | n13032 ;
  assign n13034 = x16 & x56 ;
  assign n13035 = x23 & x49 ;
  assign n13036 = n13034 | n13035 ;
  assign n13037 = x32 & x40 ;
  assign n13038 = ( n13034 & n13035 ) | ( n13034 & n13037 ) | ( n13035 & n13037 ) ;
  assign n13039 = n13036 & ~n13038 ;
  assign n13040 = n13034 & n13035 ;
  assign n13041 = n13037 & ~n13040 ;
  assign n13042 = ~n13036 & n13037 ;
  assign n13043 = ( n13037 & ~n13041 ) | ( n13037 & n13042 ) | ( ~n13041 & n13042 ) ;
  assign n13044 = n13039 | n13043 ;
  assign n13045 = n13033 & n13044 ;
  assign n13046 = n13033 & ~n13045 ;
  assign n13047 = x17 & x55 ;
  assign n13048 = n1020 & n8357 ;
  assign n13049 = x20 & x52 ;
  assign n13050 = n13047 & n13049 ;
  assign n13051 = n13048 | n13050 ;
  assign n13052 = n1285 & n11935 ;
  assign n13053 = n13047 & n13052 ;
  assign n13054 = ( n13047 & ~n13051 ) | ( n13047 & n13053 ) | ( ~n13051 & n13053 ) ;
  assign n13055 = n13051 | n13052 ;
  assign n13056 = ( n9878 & n13049 ) | ( n9878 & ~n13052 ) | ( n13049 & ~n13052 ) ;
  assign n13057 = n9878 & n13049 ;
  assign n13058 = ( ~n13051 & n13056 ) | ( ~n13051 & n13057 ) | ( n13056 & n13057 ) ;
  assign n13059 = ~n13055 & n13058 ;
  assign n13060 = n13054 | n13059 ;
  assign n13061 = ~n13033 & n13044 ;
  assign n13062 = n13060 & ~n13061 ;
  assign n13063 = ~n13046 & n13062 ;
  assign n13064 = ~n13060 & n13061 ;
  assign n13065 = ( n13046 & ~n13060 ) | ( n13046 & n13064 ) | ( ~n13060 & n13064 ) ;
  assign n13066 = n13063 | n13065 ;
  assign n13067 = x24 & x48 ;
  assign n13068 = x25 & x47 ;
  assign n13069 = n13067 | n13068 ;
  assign n13070 = n1912 & n6762 ;
  assign n13071 = x12 & x60 ;
  assign n13072 = ~n13070 & n13071 ;
  assign n13073 = n13069 | n13070 ;
  assign n13074 = ( n13070 & n13072 ) | ( n13070 & n13073 ) | ( n13072 & n13073 ) ;
  assign n13075 = n13069 & ~n13074 ;
  assign n13076 = ( ~n13069 & n13070 ) | ( ~n13069 & n13071 ) | ( n13070 & n13071 ) ;
  assign n13077 = n13071 & n13076 ;
  assign n13078 = n13075 | n13077 ;
  assign n13079 = n969 & n10856 ;
  assign n13080 = n360 & n10561 ;
  assign n13081 = n13079 | n13080 ;
  assign n13082 = n618 & n10684 ;
  assign n13083 = x63 & n13082 ;
  assign n13084 = ( x63 & ~n13081 ) | ( x63 & n13083 ) | ( ~n13081 & n13083 ) ;
  assign n13085 = x9 & n13084 ;
  assign n13086 = n13081 | n13082 ;
  assign n13087 = x10 & x62 ;
  assign n13088 = x11 & x61 ;
  assign n13089 = ( ~n13082 & n13087 ) | ( ~n13082 & n13088 ) | ( n13087 & n13088 ) ;
  assign n13090 = n13087 & n13088 ;
  assign n13091 = ( ~n13081 & n13089 ) | ( ~n13081 & n13090 ) | ( n13089 & n13090 ) ;
  assign n13092 = ~n13086 & n13091 ;
  assign n13093 = n13085 | n13092 ;
  assign n13094 = n12851 | n12855 ;
  assign n13095 = ( n12528 & n12851 ) | ( n12528 & n13094 ) | ( n12851 & n13094 ) ;
  assign n13096 = ( n13078 & n13093 ) | ( n13078 & ~n13095 ) | ( n13093 & ~n13095 ) ;
  assign n13097 = ( ~n13093 & n13095 ) | ( ~n13093 & n13096 ) | ( n13095 & n13096 ) ;
  assign n13098 = ( ~n13078 & n13096 ) | ( ~n13078 & n13097 ) | ( n13096 & n13097 ) ;
  assign n13099 = n13066 & n13098 ;
  assign n13100 = n13066 | n13098 ;
  assign n13101 = ~n13099 & n13100 ;
  assign n13102 = n12676 | n12682 ;
  assign n13103 = ( n12676 & n12679 ) | ( n12676 & n13102 ) | ( n12679 & n13102 ) ;
  assign n13104 = n13101 & n13103 ;
  assign n13105 = n13101 | n13103 ;
  assign n13106 = ~n13104 & n13105 ;
  assign n13107 = n12868 | n12883 ;
  assign n13108 = n12868 & n12883 ;
  assign n13109 = n13107 & ~n13108 ;
  assign n13110 = n12778 | n13109 ;
  assign n13111 = n12778 & n13109 ;
  assign n13112 = n13110 & ~n13111 ;
  assign n13113 = n12634 | n12639 ;
  assign n13114 = ( n12634 & n12637 ) | ( n12634 & n13113 ) | ( n12637 & n13113 ) ;
  assign n13115 = n13112 | n13114 ;
  assign n13116 = n13112 & n13114 ;
  assign n13117 = n13115 & ~n13116 ;
  assign n13118 = n723 & n9829 ;
  assign n13119 = n650 & n9831 ;
  assign n13120 = n13118 | n13119 ;
  assign n13121 = n792 & n9272 ;
  assign n13122 = x59 & n13121 ;
  assign n13123 = ( x59 & ~n13120 ) | ( x59 & n13122 ) | ( ~n13120 & n13122 ) ;
  assign n13124 = x13 & n13123 ;
  assign n13125 = n13120 | n13121 ;
  assign n13126 = x14 & x58 ;
  assign n13127 = x15 & x57 ;
  assign n13128 = ( ~n13121 & n13126 ) | ( ~n13121 & n13127 ) | ( n13126 & n13127 ) ;
  assign n13129 = n13126 & n13127 ;
  assign n13130 = ( ~n13120 & n13128 ) | ( ~n13120 & n13129 ) | ( n13128 & n13129 ) ;
  assign n13131 = ~n13125 & n13130 ;
  assign n13132 = n13124 | n13131 ;
  assign n13133 = n2895 & n8407 ;
  assign n13134 = n2267 & n5975 ;
  assign n13135 = n13133 | n13134 ;
  assign n13136 = n2372 & n6093 ;
  assign n13137 = x46 & n13136 ;
  assign n13138 = ( x46 & ~n13135 ) | ( x46 & n13137 ) | ( ~n13135 & n13137 ) ;
  assign n13139 = x26 & n13138 ;
  assign n13140 = n13135 | n13136 ;
  assign n13141 = x27 & x45 ;
  assign n13142 = x28 & x44 ;
  assign n13143 = ( ~n13136 & n13141 ) | ( ~n13136 & n13142 ) | ( n13141 & n13142 ) ;
  assign n13144 = n13141 & n13142 ;
  assign n13145 = ( ~n13135 & n13143 ) | ( ~n13135 & n13144 ) | ( n13143 & n13144 ) ;
  assign n13146 = ~n13140 & n13145 ;
  assign n13147 = n13139 | n13146 ;
  assign n13148 = n13132 & n13147 ;
  assign n13149 = n13132 & ~n13148 ;
  assign n13150 = n13147 & ~n13148 ;
  assign n13151 = n13149 | n13150 ;
  assign n13152 = x33 & x39 ;
  assign n13153 = n12377 | n13152 ;
  assign n13154 = n4530 & n5392 ;
  assign n13155 = x19 & x53 ;
  assign n13156 = ~n13154 & n13155 ;
  assign n13157 = n13153 | n13154 ;
  assign n13158 = ( n13154 & n13156 ) | ( n13154 & n13157 ) | ( n13156 & n13157 ) ;
  assign n13159 = n13153 & ~n13158 ;
  assign n13160 = ~n13153 & n13155 ;
  assign n13161 = ( n13155 & ~n13156 ) | ( n13155 & n13160 ) | ( ~n13156 & n13160 ) ;
  assign n13162 = n13159 | n13161 ;
  assign n13163 = ~n13151 & n13162 ;
  assign n13164 = n13151 & ~n13162 ;
  assign n13165 = n13163 | n13164 ;
  assign n13166 = n13117 | n13165 ;
  assign n13167 = n13117 & n13165 ;
  assign n13168 = n13166 & ~n13167 ;
  assign n13169 = n12646 | n12649 ;
  assign n13170 = ( n12646 & n12647 ) | ( n12646 & n13169 ) | ( n12647 & n13169 ) ;
  assign n13171 = n13168 & n13170 ;
  assign n13172 = n13168 | n13170 ;
  assign n13173 = ~n13171 & n13172 ;
  assign n13174 = n13106 & ~n13173 ;
  assign n13175 = ~n13106 & n13173 ;
  assign n13176 = n13174 | n13175 ;
  assign n13177 = n13021 | n13176 ;
  assign n13178 = n13018 & ~n13177 ;
  assign n13179 = n13176 | n13178 ;
  assign n13180 = ( ~n13022 & n13178 ) | ( ~n13022 & n13179 ) | ( n13178 & n13179 ) ;
  assign n13181 = n12966 | n13180 ;
  assign n13182 = n12966 & n13180 ;
  assign n13183 = n13181 & ~n13182 ;
  assign n13184 = n12666 | n12912 ;
  assign n13185 = n13183 | n13184 ;
  assign n13186 = n13183 & n13184 ;
  assign n13187 = n13185 | n13186 ;
  assign n13188 = n12913 & n12914 ;
  assign n13189 = n12913 | n12914 ;
  assign n13190 = n12629 & n13189 ;
  assign n13191 = n12612 & n13189 ;
  assign n13192 = ( n12618 & n13190 ) | ( n12618 & n13191 ) | ( n13190 & n13191 ) ;
  assign n13193 = ( n12624 & n13189 ) | ( n12624 & n13191 ) | ( n13189 & n13191 ) ;
  assign n13194 = ( n11723 & n13192 ) | ( n11723 & n13193 ) | ( n13192 & n13193 ) ;
  assign n13195 = ( n11726 & n13192 ) | ( n11726 & n13193 ) | ( n13192 & n13193 ) ;
  assign n13196 = ( n10794 & n13194 ) | ( n10794 & n13195 ) | ( n13194 & n13195 ) ;
  assign n13197 = n13188 | n13196 ;
  assign n13198 = ( n13186 & ~n13187 ) | ( n13186 & n13197 ) | ( ~n13187 & n13197 ) ;
  assign n13199 = ( n13186 & n13187 ) | ( n13186 & n13197 ) | ( n13187 & n13197 ) ;
  assign n13200 = ( n13187 & n13198 ) | ( n13187 & ~n13199 ) | ( n13198 & ~n13199 ) ;
  assign n13201 = n13185 & n13188 ;
  assign n13202 = ( n13185 & n13196 ) | ( n13185 & n13201 ) | ( n13196 & n13201 ) ;
  assign n13203 = n13186 | n13202 ;
  assign n13219 = n12778 | n13108 ;
  assign n13220 = ( n13108 & n13109 ) | ( n13108 & n13219 ) | ( n13109 & n13219 ) ;
  assign n13204 = n2683 & n6973 ;
  assign n13205 = n4062 & n5710 ;
  assign n13206 = n13204 | n13205 ;
  assign n13207 = n3321 & n5813 ;
  assign n13208 = x42 & n13207 ;
  assign n13209 = ( x42 & ~n13206 ) | ( x42 & n13208 ) | ( ~n13206 & n13208 ) ;
  assign n13210 = x31 & n13209 ;
  assign n13211 = n13206 | n13207 ;
  assign n13212 = x32 & x41 ;
  assign n13213 = x33 & x40 ;
  assign n13214 = ( ~n13207 & n13212 ) | ( ~n13207 & n13213 ) | ( n13212 & n13213 ) ;
  assign n13215 = n13212 & n13213 ;
  assign n13216 = ( ~n13206 & n13214 ) | ( ~n13206 & n13215 ) | ( n13214 & n13215 ) ;
  assign n13217 = ~n13211 & n13216 ;
  assign n13218 = n13210 | n13217 ;
  assign n13221 = n13218 & n13220 ;
  assign n13222 = n13220 & ~n13221 ;
  assign n13224 = n12825 | n12991 ;
  assign n13225 = ( n12991 & n12992 ) | ( n12991 & n13224 ) | ( n12992 & n13224 ) ;
  assign n13223 = n13218 & ~n13220 ;
  assign n13226 = n13223 & n13225 ;
  assign n13227 = ( n13222 & n13225 ) | ( n13222 & n13226 ) | ( n13225 & n13226 ) ;
  assign n13228 = n13223 | n13225 ;
  assign n13229 = n13222 | n13228 ;
  assign n13230 = ~n13227 & n13229 ;
  assign n13231 = n13006 | n13009 ;
  assign n13232 = ( n13006 & n13008 ) | ( n13006 & n13231 ) | ( n13008 & n13231 ) ;
  assign n13233 = n13230 & n13232 ;
  assign n13234 = n13230 | n13232 ;
  assign n13235 = ~n13233 & n13234 ;
  assign n13236 = n13116 | n13165 ;
  assign n13237 = ( n13116 & n13117 ) | ( n13116 & n13236 ) | ( n13117 & n13236 ) ;
  assign n13238 = n13235 & n13237 ;
  assign n13239 = n13235 | n13237 ;
  assign n13240 = ~n13238 & n13239 ;
  assign n13241 = n12984 | n13012 ;
  assign n13242 = ( n12986 & n13012 ) | ( n12986 & n13241 ) | ( n13012 & n13241 ) ;
  assign n13243 = n13240 & n13242 ;
  assign n13244 = n12988 & n13240 ;
  assign n13245 = ( n12989 & n13243 ) | ( n12989 & n13244 ) | ( n13243 & n13244 ) ;
  assign n13246 = n13240 | n13242 ;
  assign n13247 = n12988 | n13240 ;
  assign n13248 = ( n12989 & n13246 ) | ( n12989 & n13247 ) | ( n13246 & n13247 ) ;
  assign n13249 = ~n13245 & n13248 ;
  assign n13250 = n13106 | n13168 ;
  assign n13251 = ( n13106 & n13170 ) | ( n13106 & n13250 ) | ( n13170 & n13250 ) ;
  assign n13252 = ( n13171 & n13173 ) | ( n13171 & n13251 ) | ( n13173 & n13251 ) ;
  assign n13253 = n13249 & n13252 ;
  assign n13254 = n13249 | n13252 ;
  assign n13255 = ~n13253 & n13254 ;
  assign n13256 = ~n13021 & n13176 ;
  assign n13257 = n13018 & n13256 ;
  assign n13258 = n13021 & n13255 ;
  assign n13259 = ( n13255 & n13257 ) | ( n13255 & n13258 ) | ( n13257 & n13258 ) ;
  assign n13260 = n13021 | n13255 ;
  assign n13261 = n13257 | n13260 ;
  assign n13262 = ~n13259 & n13261 ;
  assign n13263 = n13078 & n13095 ;
  assign n13264 = n13078 & ~n13263 ;
  assign n13265 = ~n13078 & n13095 ;
  assign n13266 = n13264 | n13265 ;
  assign n13267 = n13093 | n13263 ;
  assign n13268 = n12728 | n13001 ;
  assign n13269 = ( n13001 & n13002 ) | ( n13001 & n13268 ) | ( n13002 & n13268 ) ;
  assign n13270 = n13267 & n13269 ;
  assign n13271 = n13263 & n13269 ;
  assign n13272 = ( n13266 & n13270 ) | ( n13266 & n13271 ) | ( n13270 & n13271 ) ;
  assign n13273 = n13267 | n13269 ;
  assign n13274 = n13263 | n13269 ;
  assign n13275 = ( n13266 & n13273 ) | ( n13266 & n13274 ) | ( n13273 & n13274 ) ;
  assign n13276 = ~n13272 & n13275 ;
  assign n13277 = n13148 | n13162 ;
  assign n13278 = ( n13148 & n13151 ) | ( n13148 & n13277 ) | ( n13151 & n13277 ) ;
  assign n13279 = n13276 | n13278 ;
  assign n13280 = n13276 & n13278 ;
  assign n13281 = n13279 & ~n13280 ;
  assign n13282 = n13099 | n13104 ;
  assign n13283 = n13281 | n13282 ;
  assign n13284 = n13281 & n13282 ;
  assign n13285 = n13283 & ~n13284 ;
  assign n13286 = x13 & x60 ;
  assign n13287 = n13029 & n13286 ;
  assign n13288 = n13029 | n13286 ;
  assign n13289 = ~n13287 & n13288 ;
  assign n13290 = n13158 | n13289 ;
  assign n13291 = n13158 & n13289 ;
  assign n13292 = n13290 & ~n13291 ;
  assign n13293 = n13074 | n13086 ;
  assign n13294 = n13074 & n13086 ;
  assign n13295 = n13293 & ~n13294 ;
  assign n13296 = n13055 | n13295 ;
  assign n13297 = n13055 & n13295 ;
  assign n13298 = n13296 & ~n13297 ;
  assign n13299 = n13292 & n13298 ;
  assign n13300 = n13292 | n13298 ;
  assign n13301 = ~n13299 & n13300 ;
  assign n13302 = n13060 & n13061 ;
  assign n13303 = ( n13046 & n13060 ) | ( n13046 & n13302 ) | ( n13060 & n13302 ) ;
  assign n13304 = n13045 | n13303 ;
  assign n13305 = n13301 & n13304 ;
  assign n13306 = n13301 | n13304 ;
  assign n13307 = ~n13305 & n13306 ;
  assign n13308 = n13285 & n13307 ;
  assign n13309 = n13285 | n13307 ;
  assign n13310 = ~n13308 & n13309 ;
  assign n13311 = n12955 | n12958 ;
  assign n13312 = ( n12955 & n12957 ) | ( n12955 & n13311 ) | ( n12957 & n13311 ) ;
  assign n13313 = n13310 | n13312 ;
  assign n13314 = n13310 & n13312 ;
  assign n13315 = n13313 & ~n13314 ;
  assign n13316 = n13125 | n13140 ;
  assign n13317 = n13125 & n13140 ;
  assign n13318 = n13316 & ~n13317 ;
  assign n13319 = n12926 | n13318 ;
  assign n13320 = n12926 & n13318 ;
  assign n13321 = n13319 & ~n13320 ;
  assign n13322 = n12934 | n12939 ;
  assign n13323 = ( n12934 & n12937 ) | ( n12934 & n13322 ) | ( n12937 & n13322 ) ;
  assign n13324 = n13321 & n13323 ;
  assign n13325 = n13321 | n13323 ;
  assign n13326 = ~n13324 & n13325 ;
  assign n13327 = n3280 & n5104 ;
  assign n13328 = n2369 & n6093 ;
  assign n13329 = n13327 | n13328 ;
  assign n13330 = n2709 & n5658 ;
  assign n13331 = x45 & n13330 ;
  assign n13332 = ( x45 & ~n13329 ) | ( x45 & n13331 ) | ( ~n13329 & n13331 ) ;
  assign n13333 = x28 & n13332 ;
  assign n13334 = n13329 | n13330 ;
  assign n13335 = x29 & x44 ;
  assign n13336 = x30 & x43 ;
  assign n13337 = ( ~n13330 & n13335 ) | ( ~n13330 & n13336 ) | ( n13335 & n13336 ) ;
  assign n13338 = n13335 & n13336 ;
  assign n13339 = ( ~n13329 & n13337 ) | ( ~n13329 & n13338 ) | ( n13337 & n13338 ) ;
  assign n13340 = ~n13334 & n13339 ;
  assign n13341 = n13333 | n13340 ;
  assign n13342 = x10 & x63 ;
  assign n13343 = x12 & x61 ;
  assign n13344 = n13342 | n13343 ;
  assign n13345 = n363 & n10856 ;
  assign n13346 = n13344 | n13345 ;
  assign n13347 = x25 & x48 ;
  assign n13348 = ( ~n13345 & n13346 ) | ( ~n13345 & n13347 ) | ( n13346 & n13347 ) ;
  assign n13349 = ( n13345 & n13346 ) | ( n13345 & ~n13347 ) | ( n13346 & ~n13347 ) ;
  assign n13350 = ( ~n13346 & n13348 ) | ( ~n13346 & n13349 ) | ( n13348 & n13349 ) ;
  assign n13351 = n13341 & n13350 ;
  assign n13352 = n13341 & ~n13351 ;
  assign n13353 = n3770 & n5225 ;
  assign n13354 = n3483 & n5392 ;
  assign n13355 = n13353 | n13354 ;
  assign n13356 = n4078 & n4857 ;
  assign n13357 = n5225 & n13356 ;
  assign n13358 = ( n5225 & ~n13355 ) | ( n5225 & n13357 ) | ( ~n13355 & n13357 ) ;
  assign n13359 = n13355 | n13356 ;
  assign n13360 = x35 & x38 ;
  assign n13361 = ( n3770 & ~n13356 ) | ( n3770 & n13360 ) | ( ~n13356 & n13360 ) ;
  assign n13362 = n3770 & n13360 ;
  assign n13363 = ( ~n13355 & n13361 ) | ( ~n13355 & n13362 ) | ( n13361 & n13362 ) ;
  assign n13364 = ~n13359 & n13363 ;
  assign n13365 = n13358 | n13364 ;
  assign n13366 = ~n13341 & n13350 ;
  assign n13367 = n13365 & ~n13366 ;
  assign n13368 = ~n13352 & n13367 ;
  assign n13369 = ~n13365 & n13366 ;
  assign n13370 = ( n13352 & ~n13365 ) | ( n13352 & n13369 ) | ( ~n13365 & n13369 ) ;
  assign n13371 = n13368 | n13370 ;
  assign n13372 = n13326 | n13371 ;
  assign n13373 = n13326 & n13371 ;
  assign n13374 = n13372 & ~n13373 ;
  assign n13375 = n12943 | n12947 ;
  assign n13376 = ( n12943 & n12945 ) | ( n12943 & n13375 ) | ( n12945 & n13375 ) ;
  assign n13377 = n13374 & n13376 ;
  assign n13378 = ( n12943 & n12949 ) | ( n12943 & ~n13377 ) | ( n12949 & ~n13377 ) ;
  assign n13379 = n1077 & n8357 ;
  assign n13380 = n4571 & n10573 ;
  assign n13381 = n13379 | n13380 ;
  assign n13382 = x49 & x54 ;
  assign n13383 = n1684 & n13382 ;
  assign n13384 = x55 & n13383 ;
  assign n13385 = ( x55 & ~n13381 ) | ( x55 & n13384 ) | ( ~n13381 & n13384 ) ;
  assign n13386 = x18 & n13385 ;
  assign n13387 = n13381 | n13383 ;
  assign n13388 = x24 & x49 ;
  assign n13389 = ( n9875 & ~n13383 ) | ( n9875 & n13388 ) | ( ~n13383 & n13388 ) ;
  assign n13390 = n9875 & n13388 ;
  assign n13391 = ( ~n13381 & n13389 ) | ( ~n13381 & n13390 ) | ( n13389 & n13390 ) ;
  assign n13392 = ~n13387 & n13391 ;
  assign n13393 = n13386 | n13392 ;
  assign n13394 = x11 & x62 ;
  assign n13395 = x37 | n13394 ;
  assign n13396 = x50 & ~x62 ;
  assign n13397 = ( x50 & ~n4860 ) | ( x50 & n13396 ) | ( ~n4860 & n13396 ) ;
  assign n13398 = ( x23 & x37 ) | ( x23 & n13394 ) | ( x37 & n13394 ) ;
  assign n13399 = x37 & n13394 ;
  assign n13400 = ( n13397 & n13398 ) | ( n13397 & n13399 ) | ( n13398 & n13399 ) ;
  assign n13401 = n13395 & ~n13400 ;
  assign n13402 = x23 & n13397 ;
  assign n13403 = ~x37 & x50 ;
  assign n13404 = ~n13394 & n13403 ;
  assign n13405 = x23 & n13404 ;
  assign n13406 = x23 & x50 ;
  assign n13407 = ( ~n13402 & n13405 ) | ( ~n13402 & n13406 ) | ( n13405 & n13406 ) ;
  assign n13408 = n13401 | n13407 ;
  assign n13409 = n13393 & n13408 ;
  assign n13410 = n13393 & ~n13409 ;
  assign n13411 = n1710 & n7874 ;
  assign n13412 = n1585 & n7567 ;
  assign n13413 = n13411 | n13412 ;
  assign n13414 = n1434 & n8161 ;
  assign n13415 = x51 & n13414 ;
  assign n13416 = ( x51 & ~n13413 ) | ( x51 & n13415 ) | ( ~n13413 & n13415 ) ;
  assign n13417 = x22 & n13416 ;
  assign n13418 = n13413 | n13414 ;
  assign n13419 = x20 & x53 ;
  assign n13420 = x21 & x52 ;
  assign n13421 = ( ~n13414 & n13419 ) | ( ~n13414 & n13420 ) | ( n13419 & n13420 ) ;
  assign n13422 = n13419 & n13420 ;
  assign n13423 = ( ~n13413 & n13421 ) | ( ~n13413 & n13422 ) | ( n13421 & n13422 ) ;
  assign n13424 = ~n13418 & n13423 ;
  assign n13425 = n13417 | n13424 ;
  assign n13426 = ~n13393 & n13408 ;
  assign n13427 = n13425 & ~n13426 ;
  assign n13428 = ~n13410 & n13427 ;
  assign n13429 = ~n13425 & n13426 ;
  assign n13430 = ( n13410 & ~n13425 ) | ( n13410 & n13429 ) | ( ~n13425 & n13429 ) ;
  assign n13431 = n13428 | n13430 ;
  assign n13432 = x26 & x47 ;
  assign n13433 = x27 & x46 ;
  assign n13434 = n13432 | n13433 ;
  assign n13435 = n2267 & n6147 ;
  assign n13436 = x17 & x56 ;
  assign n13437 = ~n13435 & n13436 ;
  assign n13438 = n13434 | n13435 ;
  assign n13439 = ( n13435 & n13437 ) | ( n13435 & n13438 ) | ( n13437 & n13438 ) ;
  assign n13440 = n13434 & ~n13439 ;
  assign n13441 = ( ~n13434 & n13435 ) | ( ~n13434 & n13436 ) | ( n13435 & n13436 ) ;
  assign n13442 = n13038 | n13436 ;
  assign n13443 = ( n13038 & n13441 ) | ( n13038 & n13442 ) | ( n13441 & n13442 ) ;
  assign n13444 = n13440 | n13443 ;
  assign n13445 = n13038 & n13436 ;
  assign n13446 = n13441 & n13445 ;
  assign n13447 = ( n13038 & n13440 ) | ( n13038 & n13446 ) | ( n13440 & n13446 ) ;
  assign n13448 = n13444 & ~n13447 ;
  assign n13449 = n790 & n9829 ;
  assign n13450 = n792 & n9831 ;
  assign n13451 = n13449 | n13450 ;
  assign n13452 = n795 & n9272 ;
  assign n13453 = x59 & n13452 ;
  assign n13454 = ( x59 & ~n13451 ) | ( x59 & n13453 ) | ( ~n13451 & n13453 ) ;
  assign n13455 = x14 & n13454 ;
  assign n13456 = n13451 | n13452 ;
  assign n13457 = x15 & x58 ;
  assign n13458 = x16 & x57 ;
  assign n13459 = ( ~n13452 & n13457 ) | ( ~n13452 & n13458 ) | ( n13457 & n13458 ) ;
  assign n13460 = n13457 & n13458 ;
  assign n13461 = ( ~n13451 & n13459 ) | ( ~n13451 & n13460 ) | ( n13459 & n13460 ) ;
  assign n13462 = ~n13456 & n13461 ;
  assign n13463 = n13455 | n13462 ;
  assign n13464 = ~n13448 & n13463 ;
  assign n13465 = n13448 & ~n13463 ;
  assign n13466 = n13464 | n13465 ;
  assign n13467 = n13431 & n13466 ;
  assign n13468 = n13431 & ~n13467 ;
  assign n13470 = n12972 | n12981 ;
  assign n13471 = ( n12972 & n12976 ) | ( n12972 & n13470 ) | ( n12976 & n13470 ) ;
  assign n13469 = ~n13431 & n13466 ;
  assign n13472 = n13469 & n13471 ;
  assign n13473 = ( n13468 & n13471 ) | ( n13468 & n13472 ) | ( n13471 & n13472 ) ;
  assign n13474 = n13469 | n13471 ;
  assign n13475 = n13468 | n13474 ;
  assign n13476 = ~n13473 & n13475 ;
  assign n13477 = n13374 & ~n13376 ;
  assign n13478 = n13476 & ~n13477 ;
  assign n13479 = ~n13378 & n13478 ;
  assign n13480 = ~n13476 & n13477 ;
  assign n13481 = ( n13378 & ~n13476 ) | ( n13378 & n13480 ) | ( ~n13476 & n13480 ) ;
  assign n13482 = n13479 | n13481 ;
  assign n13483 = ~n13315 & n13482 ;
  assign n13484 = n13310 | n13482 ;
  assign n13485 = ( n13312 & n13482 ) | ( n13312 & n13484 ) | ( n13482 & n13484 ) ;
  assign n13486 = n13313 & ~n13485 ;
  assign n13487 = n13483 | n13486 ;
  assign n13488 = n13262 | n13487 ;
  assign n13489 = n13262 & n13487 ;
  assign n13490 = n13488 & ~n13489 ;
  assign n13491 = n12964 | n13180 ;
  assign n13492 = ( n12964 & n12966 ) | ( n12964 & n13491 ) | ( n12966 & n13491 ) ;
  assign n13493 = ( n13203 & n13490 ) | ( n13203 & ~n13492 ) | ( n13490 & ~n13492 ) ;
  assign n13494 = ( ~n13490 & n13492 ) | ( ~n13490 & n13493 ) | ( n13492 & n13493 ) ;
  assign n13495 = ( ~n13203 & n13493 ) | ( ~n13203 & n13494 ) | ( n13493 & n13494 ) ;
  assign n13496 = n13245 | n13253 ;
  assign n13497 = n13211 | n13359 ;
  assign n13498 = n13211 & n13359 ;
  assign n13499 = n13497 & ~n13498 ;
  assign n13500 = n790 & n10975 ;
  assign n13501 = n792 & n10370 ;
  assign n13502 = n13500 | n13501 ;
  assign n13503 = n795 & n9831 ;
  assign n13504 = x60 & n13503 ;
  assign n13505 = ( x60 & ~n13502 ) | ( x60 & n13504 ) | ( ~n13502 & n13504 ) ;
  assign n13506 = x14 & n13505 ;
  assign n13507 = n13502 | n13503 ;
  assign n13508 = x15 & x59 ;
  assign n13509 = x16 & x58 ;
  assign n13510 = ( ~n13503 & n13508 ) | ( ~n13503 & n13509 ) | ( n13508 & n13509 ) ;
  assign n13511 = n13508 & n13509 ;
  assign n13512 = ( ~n13502 & n13510 ) | ( ~n13502 & n13511 ) | ( n13510 & n13511 ) ;
  assign n13513 = ~n13507 & n13512 ;
  assign n13514 = n13506 | n13513 ;
  assign n13515 = n13499 & n13514 ;
  assign n13516 = n13499 & ~n13515 ;
  assign n13517 = n13514 & ~n13515 ;
  assign n13518 = n13516 | n13517 ;
  assign n13519 = n13425 & n13426 ;
  assign n13520 = ( n13410 & n13425 ) | ( n13410 & n13519 ) | ( n13425 & n13519 ) ;
  assign n13521 = n13409 | n13520 ;
  assign n13522 = n13518 | n13521 ;
  assign n13523 = n13518 & n13521 ;
  assign n13524 = n13522 & ~n13523 ;
  assign n13525 = n13221 | n13227 ;
  assign n13526 = n13524 | n13525 ;
  assign n13527 = n13524 & n13525 ;
  assign n13528 = n13526 & ~n13527 ;
  assign n13529 = n13467 | n13471 ;
  assign n13530 = n13467 | n13468 ;
  assign n13531 = ( n13472 & n13529 ) | ( n13472 & n13530 ) | ( n13529 & n13530 ) ;
  assign n13532 = n13324 | n13371 ;
  assign n13533 = ( n13324 & n13326 ) | ( n13324 & n13532 ) | ( n13326 & n13532 ) ;
  assign n13534 = n13531 & n13533 ;
  assign n13535 = n13531 | n13533 ;
  assign n13536 = ~n13534 & n13535 ;
  assign n13537 = n13528 & n13536 ;
  assign n13538 = n13528 | n13536 ;
  assign n13539 = ~n13537 & n13538 ;
  assign n13540 = n13245 & n13539 ;
  assign n13541 = ( n13253 & n13539 ) | ( n13253 & n13540 ) | ( n13539 & n13540 ) ;
  assign n13542 = n13496 & ~n13541 ;
  assign n13543 = n13334 | n13439 ;
  assign n13544 = n13334 & n13439 ;
  assign n13545 = n13543 & ~n13544 ;
  assign n13546 = n13456 | n13545 ;
  assign n13547 = n13456 & n13545 ;
  assign n13548 = n13546 & ~n13547 ;
  assign n13549 = n13352 | n13366 ;
  assign n13550 = ~n13345 & n13347 ;
  assign n13551 = ( n13345 & n13346 ) | ( n13345 & n13550 ) | ( n13346 & n13550 ) ;
  assign n13552 = n13387 | n13418 ;
  assign n13553 = n13387 & n13418 ;
  assign n13554 = n13552 & ~n13553 ;
  assign n13555 = n13551 | n13554 ;
  assign n13556 = n13551 & n13554 ;
  assign n13557 = n13555 & ~n13556 ;
  assign n13558 = n13351 | n13365 ;
  assign n13559 = n13557 & n13558 ;
  assign n13560 = n13351 & n13557 ;
  assign n13561 = ( n13549 & n13559 ) | ( n13549 & n13560 ) | ( n13559 & n13560 ) ;
  assign n13562 = n13557 | n13558 ;
  assign n13563 = n13351 | n13557 ;
  assign n13564 = ( n13549 & n13562 ) | ( n13549 & n13563 ) | ( n13562 & n13563 ) ;
  assign n13565 = ~n13561 & n13564 ;
  assign n13566 = n13548 & n13565 ;
  assign n13567 = n13548 | n13565 ;
  assign n13568 = ~n13566 & n13567 ;
  assign n13569 = n13233 | n13568 ;
  assign n13570 = n13238 | n13569 ;
  assign n13571 = ( n13233 & n13238 ) | ( n13233 & n13568 ) | ( n13238 & n13568 ) ;
  assign n13572 = n13570 & ~n13571 ;
  assign n13573 = x18 & x56 ;
  assign n13574 = x25 & x49 ;
  assign n13575 = n13573 | n13574 ;
  assign n13576 = x25 & x56 ;
  assign n13577 = n11529 & n13576 ;
  assign n13578 = n5715 & ~n13577 ;
  assign n13579 = n13575 | n13577 ;
  assign n13580 = ( n13577 & n13578 ) | ( n13577 & n13579 ) | ( n13578 & n13579 ) ;
  assign n13581 = n13575 & ~n13580 ;
  assign n13582 = n5715 & ~n13575 ;
  assign n13583 = ( n5715 & ~n13578 ) | ( n5715 & n13582 ) | ( ~n13578 & n13582 ) ;
  assign n13584 = n13581 | n13583 ;
  assign n13585 = x11 & x63 ;
  assign n13586 = n4062 & n5407 ;
  assign n13587 = x31 & x43 ;
  assign n13588 = x32 & x42 ;
  assign n13589 = n13587 | n13588 ;
  assign n13590 = ( n13585 & n13586 ) | ( n13585 & ~n13589 ) | ( n13586 & ~n13589 ) ;
  assign n13591 = n13585 & ~n13590 ;
  assign n13592 = ~n13586 & n13589 ;
  assign n13593 = n13585 | n13592 ;
  assign n13594 = ~n13591 & n13593 ;
  assign n13595 = n13584 & n13594 ;
  assign n13596 = n13584 & ~n13595 ;
  assign n13597 = n2895 & n9421 ;
  assign n13598 = n2267 & n6762 ;
  assign n13599 = n13597 | n13598 ;
  assign n13600 = n2372 & n6147 ;
  assign n13601 = x48 & n13600 ;
  assign n13602 = ( x48 & ~n13599 ) | ( x48 & n13601 ) | ( ~n13599 & n13601 ) ;
  assign n13603 = x26 & n13602 ;
  assign n13604 = n13599 | n13600 ;
  assign n13605 = x27 & x47 ;
  assign n13606 = x28 & x46 ;
  assign n13607 = ( ~n13600 & n13605 ) | ( ~n13600 & n13606 ) | ( n13605 & n13606 ) ;
  assign n13608 = n13605 & n13606 ;
  assign n13609 = ( ~n13599 & n13607 ) | ( ~n13599 & n13608 ) | ( n13607 & n13608 ) ;
  assign n13610 = ~n13604 & n13609 ;
  assign n13611 = n13603 | n13610 ;
  assign n13612 = ~n13584 & n13594 ;
  assign n13613 = n13611 & ~n13612 ;
  assign n13614 = ~n13596 & n13613 ;
  assign n13615 = ~n13611 & n13612 ;
  assign n13616 = ( n13596 & ~n13611 ) | ( n13596 & n13615 ) | ( ~n13611 & n13615 ) ;
  assign n13617 = n13614 | n13616 ;
  assign n13618 = x52 & x55 ;
  assign n13619 = n4258 & n13618 ;
  assign n13620 = n1585 & n8161 ;
  assign n13621 = n13619 | n13620 ;
  assign n13622 = n1432 & n8360 ;
  assign n13623 = x52 & n13622 ;
  assign n13624 = ( x52 & ~n13621 ) | ( x52 & n13623 ) | ( ~n13621 & n13623 ) ;
  assign n13625 = x22 & n13624 ;
  assign n13626 = n13621 | n13622 ;
  assign n13627 = x21 & x53 ;
  assign n13628 = ( n8913 & ~n13622 ) | ( n8913 & n13627 ) | ( ~n13622 & n13627 ) ;
  assign n13629 = n8913 & n13627 ;
  assign n13630 = ( ~n13621 & n13628 ) | ( ~n13621 & n13629 ) | ( n13628 & n13629 ) ;
  assign n13631 = ~n13626 & n13630 ;
  assign n13632 = n13625 | n13631 ;
  assign n13633 = x35 & x39 ;
  assign n13634 = n5736 | n13633 ;
  assign n13635 = n3483 & n4555 ;
  assign n13636 = n12096 & ~n13635 ;
  assign n13637 = n13634 | n13635 ;
  assign n13638 = ( n13635 & n13636 ) | ( n13635 & n13637 ) | ( n13636 & n13637 ) ;
  assign n13639 = n13634 & ~n13638 ;
  assign n13640 = n12096 & ~n13634 ;
  assign n13641 = ( n12096 & ~n13636 ) | ( n12096 & n13640 ) | ( ~n13636 & n13640 ) ;
  assign n13642 = n13639 | n13641 ;
  assign n13643 = n13632 & n13642 ;
  assign n13644 = n13632 & ~n13643 ;
  assign n13645 = n13642 & ~n13643 ;
  assign n13646 = n13644 | n13645 ;
  assign n13647 = x23 & x51 ;
  assign n13648 = x24 & x50 ;
  assign n13649 = n13647 | n13648 ;
  assign n13650 = n1686 & n7112 ;
  assign n13651 = n3731 & ~n13650 ;
  assign n13652 = n13649 | n13650 ;
  assign n13653 = ( n13650 & n13651 ) | ( n13650 & n13652 ) | ( n13651 & n13652 ) ;
  assign n13654 = n13649 & ~n13653 ;
  assign n13655 = n3731 & ~n13649 ;
  assign n13656 = ( n3731 & ~n13651 ) | ( n3731 & n13655 ) | ( ~n13651 & n13655 ) ;
  assign n13657 = n13654 | n13656 ;
  assign n13658 = ~n13646 & n13657 ;
  assign n13659 = n13646 & ~n13657 ;
  assign n13660 = n13658 | n13659 ;
  assign n13661 = n13617 & ~n13660 ;
  assign n13662 = ~n13617 & n13660 ;
  assign n13663 = n13661 | n13662 ;
  assign n13664 = n647 & n10684 ;
  assign n13665 = x13 & x61 ;
  assign n13666 = x12 & x62 ;
  assign n13667 = n13665 | n13666 ;
  assign n13668 = ~n13664 & n13667 ;
  assign n13669 = n13400 & n13668 ;
  assign n13670 = n13400 & ~n13669 ;
  assign n13671 = n13668 & ~n13669 ;
  assign n13672 = n13670 | n13671 ;
  assign n13673 = n2709 & n6093 ;
  assign n13674 = x29 & x57 ;
  assign n13675 = n9966 & n13674 ;
  assign n13676 = n13673 | n13675 ;
  assign n13677 = x30 & x44 ;
  assign n13678 = n10619 & n13677 ;
  assign n13679 = x45 & n13678 ;
  assign n13680 = ( x45 & ~n13676 ) | ( x45 & n13679 ) | ( ~n13676 & n13679 ) ;
  assign n13681 = x29 & n13680 ;
  assign n13682 = n13676 | n13678 ;
  assign n13683 = n10619 | n13677 ;
  assign n13684 = x29 | n13683 ;
  assign n13685 = ( n13680 & n13683 ) | ( n13680 & n13684 ) | ( n13683 & n13684 ) ;
  assign n13686 = ( n13681 & ~n13682 ) | ( n13681 & n13685 ) | ( ~n13682 & n13685 ) ;
  assign n13687 = n13672 & n13686 ;
  assign n13688 = n13672 & ~n13687 ;
  assign n13690 = n12926 | n13317 ;
  assign n13691 = ( n13317 & n13318 ) | ( n13317 & n13690 ) | ( n13318 & n13690 ) ;
  assign n13689 = ~n13672 & n13686 ;
  assign n13692 = n13689 & n13691 ;
  assign n13693 = ( n13688 & n13691 ) | ( n13688 & n13692 ) | ( n13691 & n13692 ) ;
  assign n13694 = n13689 | n13691 ;
  assign n13695 = n13688 | n13694 ;
  assign n13696 = ~n13693 & n13695 ;
  assign n13697 = ~n13663 & n13696 ;
  assign n13698 = n13663 & ~n13696 ;
  assign n13699 = n13697 | n13698 ;
  assign n13700 = n13572 & n13699 ;
  assign n13701 = n13572 & ~n13700 ;
  assign n13702 = ~n13572 & n13699 ;
  assign n13703 = n13701 | n13702 ;
  assign n13704 = n13541 | n13703 ;
  assign n13705 = n13539 & ~n13703 ;
  assign n13706 = ( n13542 & ~n13704 ) | ( n13542 & n13705 ) | ( ~n13704 & n13705 ) ;
  assign n13707 = n13541 & n13703 ;
  assign n13708 = ~n13539 & n13703 ;
  assign n13709 = ( ~n13542 & n13707 ) | ( ~n13542 & n13708 ) | ( n13707 & n13708 ) ;
  assign n13710 = n13706 | n13709 ;
  assign n13711 = n13055 | n13294 ;
  assign n13712 = ( n13294 & n13295 ) | ( n13294 & n13711 ) | ( n13295 & n13711 ) ;
  assign n13713 = n13158 | n13287 ;
  assign n13714 = ( n13287 & n13289 ) | ( n13287 & n13713 ) | ( n13289 & n13713 ) ;
  assign n13715 = n13712 | n13714 ;
  assign n13716 = n13712 & n13714 ;
  assign n13717 = n13715 & ~n13716 ;
  assign n13718 = n13447 | n13463 ;
  assign n13719 = ( n13447 & n13448 ) | ( n13447 & n13718 ) | ( n13448 & n13718 ) ;
  assign n13720 = n13717 | n13719 ;
  assign n13721 = n13717 & n13719 ;
  assign n13722 = n13720 & ~n13721 ;
  assign n13723 = n13299 | n13305 ;
  assign n13724 = n13272 | n13278 ;
  assign n13725 = ( n13272 & n13276 ) | ( n13272 & n13724 ) | ( n13276 & n13724 ) ;
  assign n13726 = n13723 | n13725 ;
  assign n13727 = n13723 & n13725 ;
  assign n13728 = n13726 & ~n13727 ;
  assign n13729 = n13722 & n13728 ;
  assign n13730 = n13722 | n13728 ;
  assign n13731 = ~n13729 & n13730 ;
  assign n13732 = n13281 | n13307 ;
  assign n13733 = ( n13282 & n13307 ) | ( n13282 & n13732 ) | ( n13307 & n13732 ) ;
  assign n13734 = ( n13284 & n13285 ) | ( n13284 & n13733 ) | ( n13285 & n13733 ) ;
  assign n13735 = n13731 & n13734 ;
  assign n13736 = n13731 | n13734 ;
  assign n13737 = ~n13735 & n13736 ;
  assign n13738 = n13476 & n13477 ;
  assign n13739 = ( n13378 & n13476 ) | ( n13378 & n13738 ) | ( n13476 & n13738 ) ;
  assign n13740 = n13377 | n13739 ;
  assign n13741 = n13737 & n13740 ;
  assign n13742 = n13737 | n13740 ;
  assign n13743 = ~n13741 & n13742 ;
  assign n13744 = n13485 & n13743 ;
  assign n13745 = n13314 & n13743 ;
  assign n13746 = ( n13315 & n13744 ) | ( n13315 & n13745 ) | ( n13744 & n13745 ) ;
  assign n13747 = n13485 | n13743 ;
  assign n13748 = n13314 | n13743 ;
  assign n13749 = ( n13315 & n13747 ) | ( n13315 & n13748 ) | ( n13747 & n13748 ) ;
  assign n13750 = ~n13746 & n13749 ;
  assign n13751 = n13710 & n13750 ;
  assign n13752 = n13710 | n13750 ;
  assign n13753 = ~n13751 & n13752 ;
  assign n13754 = n13259 | n13489 ;
  assign n13755 = n13753 | n13754 ;
  assign n13756 = n13753 & n13754 ;
  assign n13757 = n13755 & ~n13756 ;
  assign n13758 = n13490 & n13492 ;
  assign n13759 = n13490 | n13492 ;
  assign n13760 = n13186 & n13759 ;
  assign n13761 = ( n13201 & n13759 ) | ( n13201 & n13760 ) | ( n13759 & n13760 ) ;
  assign n13762 = n13758 | n13761 ;
  assign n13763 = n13758 | n13759 ;
  assign n13764 = ( n13187 & n13758 ) | ( n13187 & n13763 ) | ( n13758 & n13763 ) ;
  assign n13765 = ( n13196 & n13762 ) | ( n13196 & n13764 ) | ( n13762 & n13764 ) ;
  assign n13766 = n13757 | n13765 ;
  assign n13767 = n13757 & n13765 ;
  assign n13768 = n13766 & ~n13767 ;
  assign n13769 = ( n13490 & n13753 ) | ( n13490 & n13754 ) | ( n13753 & n13754 ) ;
  assign n13770 = ( n13492 & n13756 ) | ( n13492 & n13769 ) | ( n13756 & n13769 ) ;
  assign n13771 = ( n13755 & n13761 ) | ( n13755 & n13770 ) | ( n13761 & n13770 ) ;
  assign n13772 = n13755 | n13756 ;
  assign n13773 = ( n13756 & n13763 ) | ( n13756 & n13772 ) | ( n13763 & n13772 ) ;
  assign n13774 = ( n13756 & n13758 ) | ( n13756 & n13772 ) | ( n13758 & n13772 ) ;
  assign n13775 = ( n13187 & n13773 ) | ( n13187 & n13774 ) | ( n13773 & n13774 ) ;
  assign n13776 = ( n13196 & n13771 ) | ( n13196 & n13775 ) | ( n13771 & n13775 ) ;
  assign n13777 = n13498 | n13515 ;
  assign n13778 = n13551 | n13553 ;
  assign n13779 = ( n13553 & n13554 ) | ( n13553 & n13778 ) | ( n13554 & n13778 ) ;
  assign n13780 = n13777 | n13779 ;
  assign n13781 = n13777 & n13779 ;
  assign n13782 = n13780 & ~n13781 ;
  assign n13783 = n13456 | n13544 ;
  assign n13784 = ( n13544 & n13545 ) | ( n13544 & n13783 ) | ( n13545 & n13783 ) ;
  assign n13785 = n13782 | n13784 ;
  assign n13786 = n13782 & n13784 ;
  assign n13787 = n13785 & ~n13786 ;
  assign n13788 = ( n13617 & n13660 ) | ( n13617 & n13696 ) | ( n13660 & n13696 ) ;
  assign n13789 = n13787 | n13788 ;
  assign n13790 = n13787 & n13788 ;
  assign n13791 = n13789 & ~n13790 ;
  assign n13792 = n13687 | n13693 ;
  assign n13793 = n13638 | n13653 ;
  assign n13794 = n13638 & n13653 ;
  assign n13795 = n13793 & ~n13794 ;
  assign n13796 = n13626 | n13795 ;
  assign n13797 = n13626 & n13795 ;
  assign n13798 = n13796 & ~n13797 ;
  assign n13799 = n13585 | n13586 ;
  assign n13800 = ( n13586 & ~n13590 ) | ( n13586 & n13799 ) | ( ~n13590 & n13799 ) ;
  assign n13801 = n13580 | n13800 ;
  assign n13802 = n13580 & n13800 ;
  assign n13803 = n13801 & ~n13802 ;
  assign n13804 = n13664 | n13669 ;
  assign n13805 = n13803 | n13804 ;
  assign n13806 = n13803 & n13804 ;
  assign n13807 = n13805 & ~n13806 ;
  assign n13808 = n13798 & n13807 ;
  assign n13809 = n13798 | n13807 ;
  assign n13810 = ~n13808 & n13809 ;
  assign n13811 = n13792 & n13810 ;
  assign n13812 = n13792 | n13810 ;
  assign n13813 = ~n13811 & n13812 ;
  assign n13814 = n13791 & n13813 ;
  assign n13815 = n13791 | n13813 ;
  assign n13816 = ~n13814 & n13815 ;
  assign n13817 = ( n13735 & n13741 ) | ( n13735 & n13816 ) | ( n13741 & n13816 ) ;
  assign n13818 = n13735 | n13740 ;
  assign n13819 = n13737 | n13816 ;
  assign n13820 = n13731 | n13816 ;
  assign n13821 = ( n13734 & n13816 ) | ( n13734 & n13820 ) | ( n13816 & n13820 ) ;
  assign n13822 = ( n13818 & n13819 ) | ( n13818 & n13821 ) | ( n13819 & n13821 ) ;
  assign n13823 = ~n13817 & n13822 ;
  assign n13824 = n790 & n9737 ;
  assign n13825 = n792 & n10367 ;
  assign n13826 = n13824 | n13825 ;
  assign n13827 = n795 & n10370 ;
  assign n13828 = x61 & n13827 ;
  assign n13829 = ( x61 & ~n13826 ) | ( x61 & n13828 ) | ( ~n13826 & n13828 ) ;
  assign n13830 = x14 & n13829 ;
  assign n13831 = n13826 | n13827 ;
  assign n13832 = x15 & x60 ;
  assign n13833 = x16 & x59 ;
  assign n13834 = ( ~n13827 & n13832 ) | ( ~n13827 & n13833 ) | ( n13832 & n13833 ) ;
  assign n13835 = n13832 & n13833 ;
  assign n13836 = ( ~n13826 & n13834 ) | ( ~n13826 & n13835 ) | ( n13834 & n13835 ) ;
  assign n13837 = ~n13831 & n13836 ;
  assign n13838 = n13830 | n13837 ;
  assign n13839 = x26 & x58 ;
  assign n13840 = n7666 & n13839 ;
  assign n13841 = n1020 & n9272 ;
  assign n13842 = n13840 | n13841 ;
  assign n13843 = x49 & x57 ;
  assign n13844 = n4884 & n13843 ;
  assign n13845 = n13842 | n13844 ;
  assign n13846 = x18 & x57 ;
  assign n13847 = x26 & x49 ;
  assign n13848 = ( ~n13844 & n13846 ) | ( ~n13844 & n13847 ) | ( n13846 & n13847 ) ;
  assign n13849 = n13846 & n13847 ;
  assign n13850 = ( ~n13842 & n13848 ) | ( ~n13842 & n13849 ) | ( n13848 & n13849 ) ;
  assign n13851 = ~n13845 & n13850 ;
  assign n13852 = n10616 & n13844 ;
  assign n13853 = ( n10616 & ~n13842 ) | ( n10616 & n13852 ) | ( ~n13842 & n13852 ) ;
  assign n13854 = n13851 | n13853 ;
  assign n13855 = n13838 & n13854 ;
  assign n13856 = n13838 & ~n13855 ;
  assign n13857 = n13854 & ~n13855 ;
  assign n13858 = n13856 | n13857 ;
  assign n13859 = n2075 & n9421 ;
  assign n13860 = n2372 & n6762 ;
  assign n13861 = n13859 | n13860 ;
  assign n13862 = n2369 & n6147 ;
  assign n13863 = x48 & n13862 ;
  assign n13864 = ( x48 & ~n13861 ) | ( x48 & n13863 ) | ( ~n13861 & n13863 ) ;
  assign n13865 = x27 & n13864 ;
  assign n13866 = n13861 | n13862 ;
  assign n13867 = x28 & x47 ;
  assign n13868 = x29 & x46 ;
  assign n13869 = ( ~n13862 & n13867 ) | ( ~n13862 & n13868 ) | ( n13867 & n13868 ) ;
  assign n13870 = n13867 & n13868 ;
  assign n13871 = ( ~n13861 & n13869 ) | ( ~n13861 & n13870 ) | ( n13869 & n13870 ) ;
  assign n13872 = ~n13866 & n13871 ;
  assign n13873 = n13865 | n13872 ;
  assign n13874 = ~n13858 & n13873 ;
  assign n13875 = n13858 & ~n13873 ;
  assign n13876 = n13874 | n13875 ;
  assign n13877 = n13604 | n13682 ;
  assign n13878 = n13604 & n13682 ;
  assign n13879 = n13877 & ~n13878 ;
  assign n13880 = n13507 | n13879 ;
  assign n13881 = n13507 & n13879 ;
  assign n13882 = n13880 & ~n13881 ;
  assign n13883 = n13611 & n13612 ;
  assign n13884 = ( n13596 & n13611 ) | ( n13596 & n13883 ) | ( n13611 & n13883 ) ;
  assign n13885 = n13595 | n13884 ;
  assign n13886 = n13643 | n13657 ;
  assign n13887 = ( n13643 & n13646 ) | ( n13643 & n13886 ) | ( n13646 & n13886 ) ;
  assign n13888 = n13885 | n13887 ;
  assign n13889 = n13885 & n13887 ;
  assign n13890 = n13888 & ~n13889 ;
  assign n13891 = n13882 & n13890 ;
  assign n13892 = n13882 | n13890 ;
  assign n13893 = ~n13891 & n13892 ;
  assign n13894 = n13722 | n13727 ;
  assign n13895 = ( n13727 & n13728 ) | ( n13727 & n13894 ) | ( n13728 & n13894 ) ;
  assign n13896 = n13893 & n13895 ;
  assign n13897 = n13893 | n13895 ;
  assign n13898 = ~n13896 & n13897 ;
  assign n13899 = x35 & x40 ;
  assign n13900 = n9771 | n13899 ;
  assign n13901 = n4078 & n4555 ;
  assign n13902 = x23 & x52 ;
  assign n13903 = ~n13901 & n13902 ;
  assign n13904 = n13900 | n13901 ;
  assign n13905 = ( n13901 & n13903 ) | ( n13901 & n13904 ) | ( n13903 & n13904 ) ;
  assign n13906 = n13900 & ~n13905 ;
  assign n13907 = ~n13900 & n13902 ;
  assign n13908 = ( n13902 & ~n13903 ) | ( n13902 & n13907 ) | ( ~n13903 & n13907 ) ;
  assign n13909 = n13906 | n13908 ;
  assign n13910 = x12 & x63 ;
  assign n13911 = x19 & x56 ;
  assign n13912 = n13910 | n13911 ;
  assign n13913 = x19 & x63 ;
  assign n13914 = n11925 & n13913 ;
  assign n13915 = n13912 | n13914 ;
  assign n13916 = x30 & x45 ;
  assign n13917 = ( ~n13914 & n13915 ) | ( ~n13914 & n13916 ) | ( n13915 & n13916 ) ;
  assign n13918 = ( n13914 & n13915 ) | ( n13914 & ~n13916 ) | ( n13915 & ~n13916 ) ;
  assign n13919 = ( ~n13915 & n13917 ) | ( ~n13915 & n13918 ) | ( n13917 & n13918 ) ;
  assign n13920 = n13909 & n13919 ;
  assign n13921 = n13909 & ~n13920 ;
  assign n13922 = ( x38 & x62 ) | ( x38 & ~n4857 ) | ( x62 & ~n4857 ) ;
  assign n13923 = x13 | x62 ;
  assign n13924 = ~x13 & x38 ;
  assign n13925 = ( n4857 & n13923 ) | ( n4857 & ~n13924 ) | ( n13923 & ~n13924 ) ;
  assign n13926 = ( ~x13 & x38 ) | ( ~x13 & x62 ) | ( x38 & x62 ) ;
  assign n13927 = ( x13 & n4857 ) | ( x13 & ~n13926 ) | ( n4857 & ~n13926 ) ;
  assign n13928 = ( n13922 & ~n13925 ) | ( n13922 & n13927 ) | ( ~n13925 & n13927 ) ;
  assign n13929 = ~n13919 & n13928 ;
  assign n13930 = ( n13909 & n13928 ) | ( n13909 & n13929 ) | ( n13928 & n13929 ) ;
  assign n13931 = ~n13921 & n13930 ;
  assign n13932 = n13919 & ~n13928 ;
  assign n13933 = ~n13909 & n13932 ;
  assign n13934 = ( n13921 & ~n13928 ) | ( n13921 & n13933 ) | ( ~n13928 & n13933 ) ;
  assign n13935 = n13931 | n13934 ;
  assign n13936 = n13716 | n13719 ;
  assign n13937 = ( n13716 & n13717 ) | ( n13716 & n13936 ) | ( n13717 & n13936 ) ;
  assign n13938 = n13935 | n13937 ;
  assign n13939 = n13935 & n13937 ;
  assign n13940 = n13938 & ~n13939 ;
  assign n13941 = ( n13876 & n13898 ) | ( n13876 & ~n13940 ) | ( n13898 & ~n13940 ) ;
  assign n13942 = ( ~n13898 & n13940 ) | ( ~n13898 & n13941 ) | ( n13940 & n13941 ) ;
  assign n13943 = ( ~n13876 & n13941 ) | ( ~n13876 & n13942 ) | ( n13941 & n13942 ) ;
  assign n13944 = n13823 | n13943 ;
  assign n13945 = n13823 & n13943 ;
  assign n13946 = n13944 & ~n13945 ;
  assign n13947 = ( n13539 & ~n13541 ) | ( n13539 & n13542 ) | ( ~n13541 & n13542 ) ;
  assign n14009 = n13528 | n13534 ;
  assign n14010 = ( n13534 & n13536 ) | ( n13534 & n14009 ) | ( n13536 & n14009 ) ;
  assign n13997 = n13548 | n13561 ;
  assign n13998 = ( n13561 & n13565 ) | ( n13561 & n13997 ) | ( n13565 & n13997 ) ;
  assign n13948 = n2683 & n4969 ;
  assign n13949 = n4062 & n5658 ;
  assign n13950 = n13948 | n13949 ;
  assign n13951 = n3321 & n5407 ;
  assign n13952 = x44 & n13951 ;
  assign n13953 = ( x44 & ~n13950 ) | ( x44 & n13952 ) | ( ~n13950 & n13952 ) ;
  assign n13954 = x31 & n13953 ;
  assign n13955 = n13950 | n13951 ;
  assign n13956 = x33 & x42 ;
  assign n13957 = ( n5663 & ~n13951 ) | ( n5663 & n13956 ) | ( ~n13951 & n13956 ) ;
  assign n13958 = n5663 & n13956 ;
  assign n13959 = ( ~n13950 & n13957 ) | ( ~n13950 & n13958 ) | ( n13957 & n13958 ) ;
  assign n13960 = ~n13955 & n13959 ;
  assign n13961 = n13954 | n13960 ;
  assign n13962 = x20 & x55 ;
  assign n13963 = x25 & x50 ;
  assign n13964 = n13962 | n13963 ;
  assign n13965 = x34 & x41 ;
  assign n13966 = ( n13962 & n13963 ) | ( n13962 & n13965 ) | ( n13963 & n13965 ) ;
  assign n13967 = n13964 & ~n13966 ;
  assign n13968 = n13962 & n13963 ;
  assign n13969 = n13965 & ~n13968 ;
  assign n13970 = ~n13964 & n13965 ;
  assign n13971 = ( n13965 & ~n13969 ) | ( n13965 & n13970 ) | ( ~n13969 & n13970 ) ;
  assign n13972 = n13967 | n13971 ;
  assign n13973 = n13961 & n13972 ;
  assign n13974 = n13961 & ~n13973 ;
  assign n13975 = n1585 & n8355 ;
  assign n13976 = x24 & x54 ;
  assign n13977 = n13023 & n13976 ;
  assign n13978 = n13975 | n13977 ;
  assign n13979 = n2148 & n7874 ;
  assign n13980 = x54 & n13979 ;
  assign n13981 = ( x54 & ~n13978 ) | ( x54 & n13980 ) | ( ~n13978 & n13980 ) ;
  assign n13982 = x21 & n13981 ;
  assign n13983 = n13978 | n13979 ;
  assign n13984 = x22 & x53 ;
  assign n13985 = x24 & x51 ;
  assign n13986 = ( ~n13979 & n13984 ) | ( ~n13979 & n13985 ) | ( n13984 & n13985 ) ;
  assign n13987 = n13984 & n13985 ;
  assign n13988 = ( ~n13978 & n13986 ) | ( ~n13978 & n13987 ) | ( n13986 & n13987 ) ;
  assign n13989 = ~n13983 & n13988 ;
  assign n13990 = n13982 | n13989 ;
  assign n13991 = ~n13961 & n13972 ;
  assign n13992 = n13990 & ~n13991 ;
  assign n13993 = ~n13974 & n13992 ;
  assign n13994 = ~n13990 & n13991 ;
  assign n13995 = ( n13974 & ~n13990 ) | ( n13974 & n13994 ) | ( ~n13990 & n13994 ) ;
  assign n13996 = n13993 | n13995 ;
  assign n13999 = n13996 & n13998 ;
  assign n14000 = n13998 & ~n13999 ;
  assign n14001 = n13996 & ~n13998 ;
  assign n14002 = n13523 | n13525 ;
  assign n14003 = ( n13523 & n13524 ) | ( n13523 & n14002 ) | ( n13524 & n14002 ) ;
  assign n14004 = ~n14001 & n14003 ;
  assign n14005 = ~n14000 & n14004 ;
  assign n14006 = n14001 & ~n14003 ;
  assign n14007 = ( n14000 & ~n14003 ) | ( n14000 & n14006 ) | ( ~n14003 & n14006 ) ;
  assign n14008 = n14005 | n14007 ;
  assign n14011 = n14008 & n14010 ;
  assign n14012 = n14010 & ~n14011 ;
  assign n14014 = n13571 | n13699 ;
  assign n14015 = ( n13571 & n13572 ) | ( n13571 & n14014 ) | ( n13572 & n14014 ) ;
  assign n14013 = n14008 & ~n14010 ;
  assign n14016 = n14013 & n14015 ;
  assign n14017 = ( n14012 & n14015 ) | ( n14012 & n14016 ) | ( n14015 & n14016 ) ;
  assign n14018 = n14013 | n14015 ;
  assign n14019 = n14012 | n14018 ;
  assign n14020 = ~n14017 & n14019 ;
  assign n14021 = n13704 & n14020 ;
  assign n14022 = n13541 & n14020 ;
  assign n14023 = ( n13947 & n14021 ) | ( n13947 & n14022 ) | ( n14021 & n14022 ) ;
  assign n14024 = n13704 | n14020 ;
  assign n14025 = n13541 | n14020 ;
  assign n14026 = ( n13947 & n14024 ) | ( n13947 & n14025 ) | ( n14024 & n14025 ) ;
  assign n14027 = ~n14023 & n14026 ;
  assign n14028 = n13946 & n14027 ;
  assign n14029 = n13946 | n14027 ;
  assign n14030 = ~n14028 & n14029 ;
  assign n14031 = n13710 | n13746 ;
  assign n14032 = ( n13746 & n13750 ) | ( n13746 & n14031 ) | ( n13750 & n14031 ) ;
  assign n14033 = ( n13776 & ~n14030 ) | ( n13776 & n14032 ) | ( ~n14030 & n14032 ) ;
  assign n14034 = ( n14030 & ~n14032 ) | ( n14030 & n14033 ) | ( ~n14032 & n14033 ) ;
  assign n14035 = ( ~n13776 & n14033 ) | ( ~n13776 & n14034 ) | ( n14033 & n14034 ) ;
  assign n14036 = n14023 | n14028 ;
  assign n14037 = n13802 | n13804 ;
  assign n14038 = ( n13802 & n13803 ) | ( n13802 & n14037 ) | ( n13803 & n14037 ) ;
  assign n14039 = n13507 | n13878 ;
  assign n14040 = ( n13878 & n13879 ) | ( n13878 & n14039 ) | ( n13879 & n14039 ) ;
  assign n14041 = n14038 | n14040 ;
  assign n14042 = n14038 & n14040 ;
  assign n14043 = n14041 & ~n14042 ;
  assign n14044 = n13626 | n13794 ;
  assign n14045 = ( n13794 & n13795 ) | ( n13794 & n14044 ) | ( n13795 & n14044 ) ;
  assign n14046 = n14043 | n14045 ;
  assign n14047 = n14043 & n14045 ;
  assign n14048 = n14046 & ~n14047 ;
  assign n14049 = n13876 | n13939 ;
  assign n14050 = ( n13939 & n13940 ) | ( n13939 & n14049 ) | ( n13940 & n14049 ) ;
  assign n14051 = n14048 & n14050 ;
  assign n14052 = n14048 | n14050 ;
  assign n14053 = ~n14051 & n14052 ;
  assign n14054 = ~n13914 & n13916 ;
  assign n14055 = ( n13914 & n13915 ) | ( n13914 & n14054 ) | ( n13915 & n14054 ) ;
  assign n14056 = n13862 | n13966 ;
  assign n14057 = n13861 | n14056 ;
  assign n14058 = n13862 & n13966 ;
  assign n14059 = ( n13861 & n13966 ) | ( n13861 & n14058 ) | ( n13966 & n14058 ) ;
  assign n14060 = n14057 & ~n14059 ;
  assign n14061 = n14055 | n14060 ;
  assign n14062 = n14055 & n14060 ;
  assign n14063 = n14061 & ~n14062 ;
  assign n14064 = n13974 | n13991 ;
  assign n14065 = n13973 | n13990 ;
  assign n14066 = x38 & x62 ;
  assign n14067 = x13 & n14066 ;
  assign n14068 = n4857 & ~n14067 ;
  assign n14069 = x14 & x62 ;
  assign n14070 = n14067 | n14069 ;
  assign n14071 = n14068 | n14070 ;
  assign n14072 = n14067 & n14069 ;
  assign n14073 = ( n14068 & n14069 ) | ( n14068 & n14072 ) | ( n14069 & n14072 ) ;
  assign n14074 = n13905 & ~n14073 ;
  assign n14075 = n14071 | n14073 ;
  assign n14076 = ( n14073 & n14074 ) | ( n14073 & n14075 ) | ( n14074 & n14075 ) ;
  assign n14077 = n14071 & ~n14076 ;
  assign n14078 = n13905 & ~n14071 ;
  assign n14079 = ( n13905 & ~n14074 ) | ( n13905 & n14078 ) | ( ~n14074 & n14078 ) ;
  assign n14080 = n14077 | n14079 ;
  assign n14081 = n14065 & n14080 ;
  assign n14082 = n13973 & n14080 ;
  assign n14083 = ( n14064 & n14081 ) | ( n14064 & n14082 ) | ( n14081 & n14082 ) ;
  assign n14084 = n14065 | n14080 ;
  assign n14085 = n13973 | n14080 ;
  assign n14086 = ( n14064 & n14084 ) | ( n14064 & n14085 ) | ( n14084 & n14085 ) ;
  assign n14087 = ~n14083 & n14086 ;
  assign n14088 = n14063 & ~n14087 ;
  assign n14089 = ~n14063 & n14087 ;
  assign n14090 = n14088 | n14089 ;
  assign n14091 = n14053 & ~n14090 ;
  assign n14092 = n14053 | n14090 ;
  assign n14093 = ( ~n14053 & n14091 ) | ( ~n14053 & n14092 ) | ( n14091 & n14092 ) ;
  assign n14094 = n14011 & n14093 ;
  assign n14095 = ( n14017 & n14093 ) | ( n14017 & n14094 ) | ( n14093 & n14094 ) ;
  assign n14096 = n14011 | n14093 ;
  assign n14097 = n14017 | n14096 ;
  assign n14098 = ~n14095 & n14097 ;
  assign n14099 = n913 & n9737 ;
  assign n14100 = n795 & n10367 ;
  assign n14101 = n14099 | n14100 ;
  assign n14102 = n1023 & n10370 ;
  assign n14103 = x61 & n14102 ;
  assign n14104 = ( x61 & ~n14101 ) | ( x61 & n14103 ) | ( ~n14101 & n14103 ) ;
  assign n14105 = x15 & n14104 ;
  assign n14106 = n14101 | n14102 ;
  assign n14107 = x16 & x60 ;
  assign n14108 = x17 & x59 ;
  assign n14109 = ( ~n14102 & n14107 ) | ( ~n14102 & n14108 ) | ( n14107 & n14108 ) ;
  assign n14110 = n14107 & n14108 ;
  assign n14111 = ( ~n14101 & n14109 ) | ( ~n14101 & n14110 ) | ( n14109 & n14110 ) ;
  assign n14112 = ~n14106 & n14111 ;
  assign n14113 = ~n13983 & n14112 ;
  assign n14114 = ( ~n13983 & n14105 ) | ( ~n13983 & n14113 ) | ( n14105 & n14113 ) ;
  assign n14115 = n13983 & ~n14112 ;
  assign n14116 = ~n14105 & n14115 ;
  assign n14117 = n14114 | n14116 ;
  assign n14118 = x26 & x50 ;
  assign n14119 = x27 & x49 ;
  assign n14120 = n14118 | n14119 ;
  assign n14121 = n2267 & n6834 ;
  assign n14122 = x18 & x58 ;
  assign n14123 = ~n14121 & n14122 ;
  assign n14124 = n14120 | n14121 ;
  assign n14125 = ( n14121 & n14123 ) | ( n14121 & n14124 ) | ( n14123 & n14124 ) ;
  assign n14126 = n14120 & ~n14125 ;
  assign n14127 = ( ~n14120 & n14121 ) | ( ~n14120 & n14122 ) | ( n14121 & n14122 ) ;
  assign n14128 = n14122 & n14127 ;
  assign n14129 = n14126 | n14128 ;
  assign n14130 = n14117 & n14129 ;
  assign n14131 = n14117 | n14129 ;
  assign n14132 = ~n14130 & n14131 ;
  assign n14133 = n14000 | n14001 ;
  assign n14134 = n13831 | n13845 ;
  assign n14135 = n13831 & n13845 ;
  assign n14136 = n14134 & ~n14135 ;
  assign n14137 = n13955 | n14136 ;
  assign n14138 = n13955 & n14136 ;
  assign n14139 = n14137 & ~n14138 ;
  assign n14140 = n13855 | n13873 ;
  assign n14141 = ( n13855 & n13858 ) | ( n13855 & n14140 ) | ( n13858 & n14140 ) ;
  assign n14142 = n13919 & n13928 ;
  assign n14143 = ~n13909 & n14142 ;
  assign n14144 = n13920 | n14143 ;
  assign n14145 = n13920 | n13928 ;
  assign n14146 = ( n13921 & n14144 ) | ( n13921 & n14145 ) | ( n14144 & n14145 ) ;
  assign n14147 = n14141 | n14146 ;
  assign n14148 = n14141 & n14146 ;
  assign n14149 = n14147 & ~n14148 ;
  assign n14150 = n14139 & n14149 ;
  assign n14151 = n14139 | n14149 ;
  assign n14152 = ~n14150 & n14151 ;
  assign n14153 = n13999 | n14003 ;
  assign n14154 = n14152 & n14153 ;
  assign n14155 = n13999 & n14152 ;
  assign n14156 = ( n14133 & n14154 ) | ( n14133 & n14155 ) | ( n14154 & n14155 ) ;
  assign n14157 = n14152 | n14153 ;
  assign n14158 = n13999 | n14152 ;
  assign n14159 = ( n14133 & n14157 ) | ( n14133 & n14158 ) | ( n14157 & n14158 ) ;
  assign n14160 = ~n14156 & n14159 ;
  assign n14161 = n3280 & n9421 ;
  assign n14162 = n2369 & n6762 ;
  assign n14163 = n14161 | n14162 ;
  assign n14164 = n2709 & n6147 ;
  assign n14165 = x48 & n14164 ;
  assign n14166 = ( x48 & ~n14163 ) | ( x48 & n14165 ) | ( ~n14163 & n14165 ) ;
  assign n14167 = x28 & n14166 ;
  assign n14168 = n14163 | n14164 ;
  assign n14169 = x29 & x47 ;
  assign n14170 = x30 & x46 ;
  assign n14171 = ( ~n14164 & n14169 ) | ( ~n14164 & n14170 ) | ( n14169 & n14170 ) ;
  assign n14172 = n14169 & n14170 ;
  assign n14173 = ( ~n14163 & n14171 ) | ( ~n14163 & n14172 ) | ( n14171 & n14172 ) ;
  assign n14174 = ~n14168 & n14173 ;
  assign n14175 = n14167 | n14174 ;
  assign n14176 = n4914 & n6973 ;
  assign n14177 = n3483 & n5710 ;
  assign n14178 = n14176 | n14177 ;
  assign n14179 = n4078 & n5813 ;
  assign n14180 = x42 & n14179 ;
  assign n14181 = ( x42 & ~n14178 ) | ( x42 & n14180 ) | ( ~n14178 & n14180 ) ;
  assign n14182 = x34 & n14181 ;
  assign n14183 = n14178 | n14179 ;
  assign n14184 = x35 & x41 ;
  assign n14185 = x36 & x40 ;
  assign n14186 = ( ~n14179 & n14184 ) | ( ~n14179 & n14185 ) | ( n14184 & n14185 ) ;
  assign n14187 = n14184 & n14185 ;
  assign n14188 = ( ~n14178 & n14186 ) | ( ~n14178 & n14187 ) | ( n14186 & n14187 ) ;
  assign n14189 = ~n14183 & n14188 ;
  assign n14190 = n14182 | n14189 ;
  assign n14191 = n14175 & n14190 ;
  assign n14192 = n14175 & ~n14191 ;
  assign n14193 = n14190 & ~n14191 ;
  assign n14194 = n14192 | n14193 ;
  assign n14195 = x24 & x52 ;
  assign n14196 = x25 & x51 ;
  assign n14197 = n14195 | n14196 ;
  assign n14198 = n1912 & n7567 ;
  assign n14199 = n5798 & ~n14198 ;
  assign n14200 = n14197 | n14198 ;
  assign n14201 = ( n14198 & n14199 ) | ( n14198 & n14200 ) | ( n14199 & n14200 ) ;
  assign n14202 = n14197 & ~n14201 ;
  assign n14203 = n5798 & ~n14197 ;
  assign n14204 = ( n5798 & ~n14199 ) | ( n5798 & n14203 ) | ( ~n14199 & n14203 ) ;
  assign n14205 = n14202 | n14204 ;
  assign n14206 = ~n14194 & n14205 ;
  assign n14207 = n14194 & ~n14205 ;
  assign n14208 = n14206 | n14207 ;
  assign n14209 = ( n13777 & n13779 ) | ( n13777 & n13784 ) | ( n13779 & n13784 ) ;
  assign n14210 = n14208 | n14209 ;
  assign n14211 = n14208 & n14209 ;
  assign n14212 = n14210 & ~n14211 ;
  assign n14213 = ( n14132 & n14160 ) | ( n14132 & ~n14212 ) | ( n14160 & ~n14212 ) ;
  assign n14214 = ( ~n14160 & n14212 ) | ( ~n14160 & n14213 ) | ( n14212 & n14213 ) ;
  assign n14215 = ( ~n14132 & n14213 ) | ( ~n14132 & n14214 ) | ( n14213 & n14214 ) ;
  assign n14216 = n14098 & n14215 ;
  assign n14217 = n14098 | n14215 ;
  assign n14218 = ~n14216 & n14217 ;
  assign n14219 = n13808 | n13811 ;
  assign n14220 = x13 & x63 ;
  assign n14221 = n4062 & n6093 ;
  assign n14222 = x31 & x45 ;
  assign n14223 = x32 & x44 ;
  assign n14224 = n14222 | n14223 ;
  assign n14225 = ( n14220 & n14221 ) | ( n14220 & ~n14224 ) | ( n14221 & ~n14224 ) ;
  assign n14226 = n14220 & ~n14225 ;
  assign n14227 = ~n14221 & n14224 ;
  assign n14228 = n14220 | n14227 ;
  assign n14229 = ~n14226 & n14228 ;
  assign n14230 = x19 & x57 ;
  assign n14231 = x23 & x53 ;
  assign n14232 = n14230 | n14231 ;
  assign n14233 = ( n5849 & n14230 ) | ( n5849 & n14231 ) | ( n14230 & n14231 ) ;
  assign n14234 = n14232 & ~n14233 ;
  assign n14235 = n14230 & n14231 ;
  assign n14236 = n5849 & ~n14235 ;
  assign n14237 = n5849 & ~n14232 ;
  assign n14238 = ( n5849 & ~n14236 ) | ( n5849 & n14237 ) | ( ~n14236 & n14237 ) ;
  assign n14239 = n14234 | n14238 ;
  assign n14240 = n14229 & n14239 ;
  assign n14241 = n14229 & ~n14240 ;
  assign n14242 = n14239 & ~n14240 ;
  assign n14243 = n14241 | n14242 ;
  assign n14244 = n1710 & n8146 ;
  assign n14245 = n1434 & n10013 ;
  assign n14246 = n14244 | n14245 ;
  assign n14247 = n1585 & n8357 ;
  assign n14248 = n11038 & n14247 ;
  assign n14249 = ( n11038 & ~n14246 ) | ( n11038 & n14248 ) | ( ~n14246 & n14248 ) ;
  assign n14250 = n14246 | n14247 ;
  assign n14251 = x21 & x55 ;
  assign n14252 = x22 & x54 ;
  assign n14253 = ( ~n14247 & n14251 ) | ( ~n14247 & n14252 ) | ( n14251 & n14252 ) ;
  assign n14254 = n14251 & n14252 ;
  assign n14255 = ( ~n14246 & n14253 ) | ( ~n14246 & n14254 ) | ( n14253 & n14254 ) ;
  assign n14256 = ~n14250 & n14255 ;
  assign n14257 = n14249 | n14256 ;
  assign n14258 = ~n14243 & n14257 ;
  assign n14259 = n14243 & ~n14257 ;
  assign n14260 = n14258 | n14259 ;
  assign n14261 = n13882 | n13889 ;
  assign n14262 = ( n13889 & n13890 ) | ( n13889 & n14261 ) | ( n13890 & n14261 ) ;
  assign n14263 = n14260 & n14262 ;
  assign n14264 = n14260 | n14262 ;
  assign n14265 = ~n14263 & n14264 ;
  assign n14266 = n14219 & n14265 ;
  assign n14267 = n14219 | n14265 ;
  assign n14268 = ~n14266 & n14267 ;
  assign n14269 = ( n13787 & n13788 ) | ( n13787 & n13813 ) | ( n13788 & n13813 ) ;
  assign n14270 = n14268 | n14269 ;
  assign n14271 = n14268 & n14269 ;
  assign n14272 = n14270 & ~n14271 ;
  assign n14273 = n13876 & n13940 ;
  assign n14274 = n13876 | n13940 ;
  assign n14275 = ~n14273 & n14274 ;
  assign n14276 = n13893 | n14275 ;
  assign n14277 = ( n13895 & n14275 ) | ( n13895 & n14276 ) | ( n14275 & n14276 ) ;
  assign n14278 = ( n13896 & n13898 ) | ( n13896 & n14277 ) | ( n13898 & n14277 ) ;
  assign n14279 = n14272 & n14278 ;
  assign n14280 = n14272 | n14278 ;
  assign n14281 = ~n14279 & n14280 ;
  assign n14282 = n13817 | n13943 ;
  assign n14283 = ( n13817 & n13823 ) | ( n13817 & n14282 ) | ( n13823 & n14282 ) ;
  assign n14284 = n14281 & n14283 ;
  assign n14285 = n14281 | n14283 ;
  assign n14286 = ~n14284 & n14285 ;
  assign n14287 = ~n14218 & n14286 ;
  assign n14288 = n14036 & n14287 ;
  assign n14289 = n14218 & ~n14286 ;
  assign n14290 = ( n14036 & n14288 ) | ( n14036 & n14289 ) | ( n14288 & n14289 ) ;
  assign n14291 = n14036 | n14287 ;
  assign n14292 = n14289 | n14291 ;
  assign n14293 = ~n14290 & n14292 ;
  assign n14294 = n14030 & n14032 ;
  assign n14295 = n14030 | n14032 ;
  assign n14296 = n13775 & n14295 ;
  assign n14297 = n14294 | n14296 ;
  assign n14298 = n14294 | n14295 ;
  assign n14299 = ( n13770 & n14294 ) | ( n13770 & n14298 ) | ( n14294 & n14298 ) ;
  assign n14300 = ( n13755 & n14294 ) | ( n13755 & n14298 ) | ( n14294 & n14298 ) ;
  assign n14301 = ( n13761 & n14299 ) | ( n13761 & n14300 ) | ( n14299 & n14300 ) ;
  assign n14302 = ( n13196 & n14297 ) | ( n13196 & n14301 ) | ( n14297 & n14301 ) ;
  assign n14303 = n14293 & n14302 ;
  assign n14304 = n14293 | n14302 ;
  assign n14305 = ~n14303 & n14304 ;
  assign n14561 = n14218 | n14284 ;
  assign n14562 = ( n14284 & n14286 ) | ( n14284 & n14561 ) | ( n14286 & n14561 ) ;
  assign n14306 = n1557 & n11935 ;
  assign n14307 = n1912 & n8161 ;
  assign n14308 = n14306 | n14307 ;
  assign n14309 = n1686 & n8355 ;
  assign n14310 = x52 & n14309 ;
  assign n14311 = ( x52 & ~n14308 ) | ( x52 & n14310 ) | ( ~n14308 & n14310 ) ;
  assign n14312 = x25 & n14311 ;
  assign n14313 = n14308 | n14309 ;
  assign n14314 = x23 & x54 ;
  assign n14315 = x24 & x53 ;
  assign n14316 = ( ~n14309 & n14314 ) | ( ~n14309 & n14315 ) | ( n14314 & n14315 ) ;
  assign n14317 = n14314 & n14315 ;
  assign n14318 = ( ~n14308 & n14316 ) | ( ~n14308 & n14317 ) | ( n14316 & n14317 ) ;
  assign n14319 = ~n14313 & n14318 ;
  assign n14320 = n14312 | n14319 ;
  assign n14321 = x22 & x55 ;
  assign n14322 = x26 & x51 ;
  assign n14323 = n14321 | n14322 ;
  assign n14324 = x34 & x43 ;
  assign n14325 = ( n14321 & n14322 ) | ( n14321 & n14324 ) | ( n14322 & n14324 ) ;
  assign n14326 = n14323 & ~n14325 ;
  assign n14327 = n14321 & n14322 ;
  assign n14328 = n14324 & ~n14327 ;
  assign n14329 = ~n14323 & n14324 ;
  assign n14330 = ( n14324 & ~n14328 ) | ( n14324 & n14329 ) | ( ~n14328 & n14329 ) ;
  assign n14331 = n14326 | n14330 ;
  assign n14332 = n14320 & n14331 ;
  assign n14333 = n14320 & ~n14332 ;
  assign n14334 = x32 & x45 ;
  assign n14335 = n5845 | n14334 ;
  assign n14336 = n3321 & n6093 ;
  assign n14337 = x16 & x61 ;
  assign n14338 = ~n14336 & n14337 ;
  assign n14339 = n14335 | n14336 ;
  assign n14340 = ( n14336 & n14338 ) | ( n14336 & n14339 ) | ( n14338 & n14339 ) ;
  assign n14341 = n14335 & ~n14340 ;
  assign n14342 = ( ~n14335 & n14336 ) | ( ~n14335 & n14337 ) | ( n14336 & n14337 ) ;
  assign n14343 = n14337 & n14342 ;
  assign n14344 = n14341 | n14343 ;
  assign n14345 = ~n14320 & n14331 ;
  assign n14346 = n14344 & ~n14345 ;
  assign n14347 = ~n14333 & n14346 ;
  assign n14348 = ~n14344 & n14345 ;
  assign n14349 = ( n14333 & ~n14344 ) | ( n14333 & n14348 ) | ( ~n14344 & n14348 ) ;
  assign n14350 = n14347 | n14349 ;
  assign n14351 = n14139 | n14146 ;
  assign n14352 = ( n14139 & n14141 ) | ( n14139 & n14351 ) | ( n14141 & n14351 ) ;
  assign n14356 = n14350 & ~n14352 ;
  assign n14357 = ~n14148 & n14350 ;
  assign n14358 = ( ~n14149 & n14356 ) | ( ~n14149 & n14357 ) | ( n14356 & n14357 ) ;
  assign n14353 = ( n14148 & n14149 ) | ( n14148 & n14352 ) | ( n14149 & n14352 ) ;
  assign n14354 = n14063 | n14083 ;
  assign n14355 = ( n14083 & n14087 ) | ( n14083 & n14354 ) | ( n14087 & n14354 ) ;
  assign n14359 = ( n14353 & n14355 ) | ( n14353 & n14358 ) | ( n14355 & n14358 ) ;
  assign n14360 = ( ~n14350 & n14358 ) | ( ~n14350 & n14359 ) | ( n14358 & n14359 ) ;
  assign n14361 = n14353 | n14355 ;
  assign n14362 = n14350 & n14352 ;
  assign n14363 = n14148 & n14350 ;
  assign n14364 = ( n14149 & n14362 ) | ( n14149 & n14363 ) | ( n14362 & n14363 ) ;
  assign n14365 = ~n14358 & n14364 ;
  assign n14366 = n14355 | n14358 ;
  assign n14367 = ( n14361 & ~n14365 ) | ( n14361 & n14366 ) | ( ~n14365 & n14366 ) ;
  assign n14368 = ~n14360 & n14367 ;
  assign n14369 = n14051 | n14090 ;
  assign n14370 = ( n14051 & n14053 ) | ( n14051 & n14369 ) | ( n14053 & n14369 ) ;
  assign n14371 = n14368 & n14370 ;
  assign n14372 = n14368 | n14370 ;
  assign n14373 = ~n14371 & n14372 ;
  assign n14374 = n14132 & n14212 ;
  assign n14375 = n14132 | n14212 ;
  assign n14376 = ~n14374 & n14375 ;
  assign n14377 = n14156 | n14376 ;
  assign n14378 = ( n14156 & n14160 ) | ( n14156 & n14377 ) | ( n14160 & n14377 ) ;
  assign n14379 = n14373 & n14378 ;
  assign n14380 = n14373 | n14378 ;
  assign n14381 = ~n14379 & n14380 ;
  assign n14382 = n14095 | n14215 ;
  assign n14383 = ( n14095 & n14098 ) | ( n14095 & n14382 ) | ( n14098 & n14382 ) ;
  assign n14384 = n14381 & n14383 ;
  assign n14385 = n14381 | n14383 ;
  assign n14386 = ~n14384 & n14385 ;
  assign n14387 = n1020 & n10370 ;
  assign n14388 = x18 & x59 ;
  assign n14389 = x17 & x60 ;
  assign n14390 = n14388 | n14389 ;
  assign n14391 = ~n14387 & n14390 ;
  assign n14392 = n14201 & n14391 ;
  assign n14393 = n14201 & ~n14392 ;
  assign n14394 = ~n14201 & n14391 ;
  assign n14395 = n14393 | n14394 ;
  assign n14396 = n13955 | n14135 ;
  assign n14397 = ( n14135 & n14136 ) | ( n14135 & n14396 ) | ( n14136 & n14396 ) ;
  assign n14398 = n14395 | n14397 ;
  assign n14399 = n14395 & n14397 ;
  assign n14400 = n14398 & ~n14399 ;
  assign n14401 = n14055 | n14059 ;
  assign n14402 = ( n14059 & n14060 ) | ( n14059 & n14401 ) | ( n14060 & n14401 ) ;
  assign n14403 = n14400 | n14402 ;
  assign n14404 = n14400 & n14402 ;
  assign n14405 = n14403 & ~n14404 ;
  assign n14406 = n14132 | n14209 ;
  assign n14407 = ( n14132 & n14208 ) | ( n14132 & n14406 ) | ( n14208 & n14406 ) ;
  assign n14408 = n14405 & n14407 ;
  assign n14409 = n14211 & n14405 ;
  assign n14410 = ( n14212 & n14408 ) | ( n14212 & n14409 ) | ( n14408 & n14409 ) ;
  assign n14411 = n14405 | n14407 ;
  assign n14412 = n14211 | n14405 ;
  assign n14413 = ( n14212 & n14411 ) | ( n14212 & n14412 ) | ( n14411 & n14412 ) ;
  assign n14414 = ~n14410 & n14413 ;
  assign n14415 = n14168 | n14250 ;
  assign n14416 = n14168 & n14250 ;
  assign n14417 = n14415 & ~n14416 ;
  assign n14418 = n14220 | n14221 ;
  assign n14419 = ( n14221 & ~n14225 ) | ( n14221 & n14418 ) | ( ~n14225 & n14418 ) ;
  assign n14420 = n14417 | n14419 ;
  assign n14421 = n14417 & n14419 ;
  assign n14422 = n14420 & ~n14421 ;
  assign n14423 = n14106 | n14125 ;
  assign n14424 = n14106 & n14125 ;
  assign n14425 = n14423 & ~n14424 ;
  assign n14426 = n14233 | n14425 ;
  assign n14427 = n14233 & n14425 ;
  assign n14428 = n14426 & ~n14427 ;
  assign n14429 = n14240 | n14257 ;
  assign n14430 = ( n14240 & n14243 ) | ( n14240 & n14429 ) | ( n14243 & n14429 ) ;
  assign n14431 = n14428 & n14430 ;
  assign n14432 = n14428 | n14430 ;
  assign n14433 = ~n14431 & n14432 ;
  assign n14434 = n14422 & n14433 ;
  assign n14435 = n14422 | n14433 ;
  assign n14436 = ~n14434 & n14435 ;
  assign n14437 = n14414 & n14436 ;
  assign n14438 = n14414 | n14436 ;
  assign n14439 = ~n14437 & n14438 ;
  assign n14440 = n14271 | n14278 ;
  assign n14441 = ( n14271 & n14272 ) | ( n14271 & n14440 ) | ( n14272 & n14440 ) ;
  assign n14442 = n14439 | n14441 ;
  assign n14443 = n14439 & n14441 ;
  assign n14444 = n14442 & ~n14443 ;
  assign n14445 = n14105 | n14112 ;
  assign n14446 = ( n13983 & n14129 ) | ( n13983 & n14445 ) | ( n14129 & n14445 ) ;
  assign n14447 = n14076 | n14446 ;
  assign n14448 = n14076 & n14446 ;
  assign n14449 = n14447 & ~n14448 ;
  assign n14450 = n14191 | n14205 ;
  assign n14451 = ( n14191 & n14194 ) | ( n14191 & n14450 ) | ( n14194 & n14450 ) ;
  assign n14452 = n14449 | n14451 ;
  assign n14453 = n14449 & n14451 ;
  assign n14454 = n14452 & ~n14453 ;
  assign n14455 = n14219 | n14260 ;
  assign n14456 = ( n14219 & n14262 ) | ( n14219 & n14455 ) | ( n14262 & n14455 ) ;
  assign n14457 = n14454 | n14456 ;
  assign n14458 = n14263 | n14454 ;
  assign n14459 = ( n14265 & n14457 ) | ( n14265 & n14458 ) | ( n14457 & n14458 ) ;
  assign n14460 = n14454 & n14456 ;
  assign n14461 = n14263 & n14454 ;
  assign n14462 = ( n14265 & n14460 ) | ( n14265 & n14461 ) | ( n14460 & n14461 ) ;
  assign n14463 = n14459 & ~n14462 ;
  assign n14464 = x30 & x47 ;
  assign n14465 = n2965 & n6147 ;
  assign n14466 = x14 & x63 ;
  assign n14467 = n14464 & n14466 ;
  assign n14468 = n14465 | n14467 ;
  assign n14469 = x31 & x63 ;
  assign n14470 = n8128 & n14469 ;
  assign n14471 = n14464 & n14470 ;
  assign n14472 = ( n14464 & ~n14468 ) | ( n14464 & n14471 ) | ( ~n14468 & n14471 ) ;
  assign n14473 = n14468 | n14470 ;
  assign n14474 = x31 & x46 ;
  assign n14475 = ( n14466 & ~n14470 ) | ( n14466 & n14474 ) | ( ~n14470 & n14474 ) ;
  assign n14476 = n14466 & n14474 ;
  assign n14477 = ( ~n14468 & n14475 ) | ( ~n14468 & n14476 ) | ( n14475 & n14476 ) ;
  assign n14478 = ~n14473 & n14477 ;
  assign n14479 = n14472 | n14478 ;
  assign n14480 = x35 & x42 ;
  assign n14481 = n5417 & n6973 ;
  assign n14482 = n4078 & n5710 ;
  assign n14483 = n14481 | n14482 ;
  assign n14484 = n3770 & n5813 ;
  assign n14485 = n14480 & n14484 ;
  assign n14486 = ( n14480 & ~n14483 ) | ( n14480 & n14485 ) | ( ~n14483 & n14485 ) ;
  assign n14487 = n14483 | n14484 ;
  assign n14488 = x36 & x41 ;
  assign n14489 = ( n6159 & ~n14484 ) | ( n6159 & n14488 ) | ( ~n14484 & n14488 ) ;
  assign n14490 = n6159 & n14488 ;
  assign n14491 = ( ~n14483 & n14489 ) | ( ~n14483 & n14490 ) | ( n14489 & n14490 ) ;
  assign n14492 = ~n14487 & n14491 ;
  assign n14493 = n14486 | n14492 ;
  assign n14494 = n14479 & n14493 ;
  assign n14495 = n14479 & ~n14494 ;
  assign n14496 = n14493 & ~n14494 ;
  assign n14497 = n14495 | n14496 ;
  assign n14498 = x62 & n7582 ;
  assign n14499 = n5392 & n14498 ;
  assign n14500 = n5392 & ~n14498 ;
  assign n14501 = n14498 | n14500 ;
  assign n14502 = x15 & x62 ;
  assign n14503 = ( x39 & ~n14498 ) | ( x39 & n14502 ) | ( ~n14498 & n14502 ) ;
  assign n14504 = x39 & n14502 ;
  assign n14505 = ( ~n14500 & n14503 ) | ( ~n14500 & n14504 ) | ( n14503 & n14504 ) ;
  assign n14506 = ~n14501 & n14505 ;
  assign n14507 = n14499 | n14506 ;
  assign n14508 = ~n14497 & n14507 ;
  assign n14509 = n14497 & ~n14507 ;
  assign n14510 = n14508 | n14509 ;
  assign n14511 = ( n14038 & n14040 ) | ( n14038 & n14045 ) | ( n14040 & n14045 ) ;
  assign n14512 = n14510 | n14511 ;
  assign n14513 = n14510 & n14511 ;
  assign n14514 = n14512 & ~n14513 ;
  assign n14515 = n1432 & n8708 ;
  assign n14516 = n1437 & n9272 ;
  assign n14517 = n14515 | n14516 ;
  assign n14518 = n1434 & n8903 ;
  assign n14519 = x58 & n14518 ;
  assign n14520 = ( x58 & ~n14517 ) | ( x58 & n14519 ) | ( ~n14517 & n14519 ) ;
  assign n14521 = x19 & n14520 ;
  assign n14522 = n14517 | n14518 ;
  assign n14523 = x21 & x56 ;
  assign n14524 = ( n11660 & ~n14518 ) | ( n11660 & n14523 ) | ( ~n14518 & n14523 ) ;
  assign n14525 = n11660 & n14523 ;
  assign n14526 = ( ~n14517 & n14524 ) | ( ~n14517 & n14525 ) | ( n14524 & n14525 ) ;
  assign n14527 = ~n14522 & n14526 ;
  assign n14528 = ~n14183 & n14527 ;
  assign n14529 = ( ~n14183 & n14521 ) | ( ~n14183 & n14528 ) | ( n14521 & n14528 ) ;
  assign n14530 = n14183 & ~n14527 ;
  assign n14531 = ~n14521 & n14530 ;
  assign n14532 = n14529 | n14531 ;
  assign n14533 = n2075 & n6345 ;
  assign n14534 = n2372 & n6834 ;
  assign n14535 = n14533 | n14534 ;
  assign n14536 = n2369 & n6759 ;
  assign n14537 = x50 & n14536 ;
  assign n14538 = ( x50 & ~n14535 ) | ( x50 & n14537 ) | ( ~n14535 & n14537 ) ;
  assign n14539 = x27 & n14538 ;
  assign n14540 = n14535 | n14536 ;
  assign n14541 = x28 & x49 ;
  assign n14542 = x29 & x48 ;
  assign n14543 = ( ~n14536 & n14541 ) | ( ~n14536 & n14542 ) | ( n14541 & n14542 ) ;
  assign n14544 = n14541 & n14542 ;
  assign n14545 = ( ~n14535 & n14543 ) | ( ~n14535 & n14544 ) | ( n14543 & n14544 ) ;
  assign n14546 = ~n14540 & n14545 ;
  assign n14547 = n14539 | n14546 ;
  assign n14548 = n14532 & n14547 ;
  assign n14549 = n14532 | n14547 ;
  assign n14550 = ~n14548 & n14549 ;
  assign n14551 = n14514 & n14550 ;
  assign n14552 = n14514 | n14550 ;
  assign n14553 = ~n14551 & n14552 ;
  assign n14554 = ~n14463 & n14553 ;
  assign n14555 = n14463 & ~n14553 ;
  assign n14556 = n14554 | n14555 ;
  assign n14557 = n14444 & n14556 ;
  assign n14558 = n14444 | n14556 ;
  assign n14559 = ~n14557 & n14558 ;
  assign n14560 = ~n14386 & n14559 ;
  assign n14563 = n14560 & n14562 ;
  assign n14564 = n14386 & ~n14559 ;
  assign n14565 = ( n14562 & n14563 ) | ( n14562 & n14564 ) | ( n14563 & n14564 ) ;
  assign n14566 = n14560 | n14562 ;
  assign n14567 = n14564 | n14566 ;
  assign n14568 = ~n14565 & n14567 ;
  assign n14569 = n14292 & n14299 ;
  assign n14570 = n14292 & n14300 ;
  assign n14571 = ( n13761 & n14569 ) | ( n13761 & n14570 ) | ( n14569 & n14570 ) ;
  assign n14572 = n14292 & n14294 ;
  assign n14573 = ( n14292 & n14295 ) | ( n14292 & n14572 ) | ( n14295 & n14572 ) ;
  assign n14574 = n14292 & n14572 ;
  assign n14575 = ( n13775 & n14573 ) | ( n13775 & n14574 ) | ( n14573 & n14574 ) ;
  assign n14576 = ( n13196 & n14571 ) | ( n13196 & n14575 ) | ( n14571 & n14575 ) ;
  assign n14577 = n14290 | n14576 ;
  assign n14578 = n14568 | n14577 ;
  assign n14579 = n14568 & n14577 ;
  assign n14580 = n14578 & ~n14579 ;
  assign n14581 = n14290 & n14567 ;
  assign n14582 = n14565 | n14581 ;
  assign n14583 = n14565 | n14567 ;
  assign n14584 = ( n14576 & n14582 ) | ( n14576 & n14583 ) | ( n14582 & n14583 ) ;
  assign n14585 = n14511 | n14550 ;
  assign n14586 = ( n14510 & n14550 ) | ( n14510 & n14585 ) | ( n14550 & n14585 ) ;
  assign n14587 = ( n14513 & n14514 ) | ( n14513 & n14586 ) | ( n14514 & n14586 ) ;
  assign n14588 = n14364 & n14587 ;
  assign n14589 = ( n14360 & n14587 ) | ( n14360 & n14588 ) | ( n14587 & n14588 ) ;
  assign n14590 = n14358 | n14364 ;
  assign n14591 = n14350 & ~n14364 ;
  assign n14592 = ( n14359 & n14590 ) | ( n14359 & ~n14591 ) | ( n14590 & ~n14591 ) ;
  assign n14593 = ~n14589 & n14592 ;
  assign n14594 = x36 & x42 ;
  assign n14595 = n6074 | n14594 ;
  assign n14596 = n4078 & n5407 ;
  assign n14597 = n14595 | n14596 ;
  assign n14598 = x23 & x55 ;
  assign n14599 = ( ~n14596 & n14597 ) | ( ~n14596 & n14598 ) | ( n14597 & n14598 ) ;
  assign n14600 = ( n14596 & n14597 ) | ( n14596 & ~n14598 ) | ( n14597 & ~n14598 ) ;
  assign n14601 = ( ~n14597 & n14599 ) | ( ~n14597 & n14600 ) | ( n14599 & n14600 ) ;
  assign n14602 = x26 & x52 ;
  assign n14603 = n4050 & n14602 ;
  assign n14604 = n6408 & n14602 ;
  assign n14605 = n4857 & n5813 ;
  assign n14606 = n14604 | n14605 ;
  assign n14607 = n6408 & n14603 ;
  assign n14608 = ( n6408 & ~n14606 ) | ( n6408 & n14607 ) | ( ~n14606 & n14607 ) ;
  assign n14609 = ( n4050 & n14602 ) | ( n4050 & ~n14606 ) | ( n14602 & ~n14606 ) ;
  assign n14610 = ( ~n14603 & n14608 ) | ( ~n14603 & n14609 ) | ( n14608 & n14609 ) ;
  assign n14611 = n14601 & n14610 ;
  assign n14612 = n14601 & ~n14611 ;
  assign n14614 = n14416 | n14419 ;
  assign n14615 = ( n14416 & n14417 ) | ( n14416 & n14614 ) | ( n14417 & n14614 ) ;
  assign n14613 = ~n14601 & n14610 ;
  assign n14616 = n14613 & n14615 ;
  assign n14617 = ( n14612 & n14615 ) | ( n14612 & n14616 ) | ( n14615 & n14616 ) ;
  assign n14618 = n14613 | n14615 ;
  assign n14619 = n14612 | n14618 ;
  assign n14620 = ~n14617 & n14619 ;
  assign n14621 = n14325 & n14518 ;
  assign n14622 = ( n14325 & n14517 ) | ( n14325 & n14621 ) | ( n14517 & n14621 ) ;
  assign n14623 = n14325 | n14518 ;
  assign n14624 = n14517 | n14623 ;
  assign n14625 = ~n14622 & n14624 ;
  assign n14626 = n14387 | n14391 ;
  assign n14627 = ( n14201 & n14387 ) | ( n14201 & n14626 ) | ( n14387 & n14626 ) ;
  assign n14628 = n14625 | n14627 ;
  assign n14629 = n14625 & n14627 ;
  assign n14630 = n14628 & ~n14629 ;
  assign n14631 = n14399 | n14402 ;
  assign n14632 = ( n14399 & n14400 ) | ( n14399 & n14631 ) | ( n14400 & n14631 ) ;
  assign n14633 = n14630 | n14632 ;
  assign n14634 = n14630 & n14632 ;
  assign n14635 = n14633 & ~n14634 ;
  assign n14636 = n14620 & n14635 ;
  assign n14637 = n14620 | n14635 ;
  assign n14638 = ~n14636 & n14637 ;
  assign n14639 = n14587 & ~n14588 ;
  assign n14640 = ~n14360 & n14638 ;
  assign n14641 = n14639 & n14640 ;
  assign n14642 = ( n14593 & n14638 ) | ( n14593 & n14641 ) | ( n14638 & n14641 ) ;
  assign n14643 = n14360 & ~n14638 ;
  assign n14644 = ( n14638 & n14639 ) | ( n14638 & ~n14643 ) | ( n14639 & ~n14643 ) ;
  assign n14645 = n14593 | n14644 ;
  assign n14646 = ~n14642 & n14645 ;
  assign n14647 = x57 & x60 ;
  assign n14648 = n3850 & n14647 ;
  assign n14649 = n1077 & n10370 ;
  assign n14650 = n14648 | n14649 ;
  assign n14651 = n1432 & n9829 ;
  assign n14652 = x60 & n14651 ;
  assign n14653 = ( x60 & ~n14650 ) | ( x60 & n14652 ) | ( ~n14650 & n14652 ) ;
  assign n14654 = x18 & n14653 ;
  assign n14655 = n14650 | n14651 ;
  assign n14656 = x19 & x59 ;
  assign n14657 = x21 & x57 ;
  assign n14658 = ( ~n14651 & n14656 ) | ( ~n14651 & n14657 ) | ( n14656 & n14657 ) ;
  assign n14659 = n14656 & n14657 ;
  assign n14660 = ( ~n14650 & n14658 ) | ( ~n14650 & n14659 ) | ( n14658 & n14659 ) ;
  assign n14661 = ~n14655 & n14660 ;
  assign n14662 = n14654 | n14661 ;
  assign n14663 = n2075 & n10866 ;
  assign n14664 = n2372 & n7112 ;
  assign n14665 = n14663 | n14664 ;
  assign n14666 = n2369 & n6834 ;
  assign n14667 = x51 & n14666 ;
  assign n14668 = ( x51 & ~n14665 ) | ( x51 & n14667 ) | ( ~n14665 & n14667 ) ;
  assign n14669 = x27 & n14668 ;
  assign n14670 = n14665 | n14666 ;
  assign n14671 = x28 & x50 ;
  assign n14672 = x29 & x49 ;
  assign n14673 = ( ~n14666 & n14671 ) | ( ~n14666 & n14672 ) | ( n14671 & n14672 ) ;
  assign n14674 = n14671 & n14672 ;
  assign n14675 = ( ~n14665 & n14673 ) | ( ~n14665 & n14674 ) | ( n14673 & n14674 ) ;
  assign n14676 = ~n14670 & n14675 ;
  assign n14677 = n14669 | n14676 ;
  assign n14678 = n14662 & n14677 ;
  assign n14679 = n14662 & ~n14678 ;
  assign n14680 = n14677 & ~n14678 ;
  assign n14681 = n14679 | n14680 ;
  assign n14682 = n913 & n10856 ;
  assign n14683 = n795 & n10561 ;
  assign n14684 = n14682 | n14683 ;
  assign n14685 = n1023 & n10684 ;
  assign n14686 = x63 & n14685 ;
  assign n14687 = ( x63 & ~n14684 ) | ( x63 & n14686 ) | ( ~n14684 & n14686 ) ;
  assign n14688 = x15 & n14687 ;
  assign n14689 = n14684 | n14685 ;
  assign n14690 = x16 & x62 ;
  assign n14691 = x17 & x61 ;
  assign n14692 = ( ~n14685 & n14690 ) | ( ~n14685 & n14691 ) | ( n14690 & n14691 ) ;
  assign n14693 = n14690 & n14691 ;
  assign n14694 = ( ~n14684 & n14692 ) | ( ~n14684 & n14693 ) | ( n14692 & n14693 ) ;
  assign n14695 = ~n14689 & n14694 ;
  assign n14696 = n14688 | n14695 ;
  assign n14697 = ~n14681 & n14696 ;
  assign n14698 = n14681 & ~n14696 ;
  assign n14699 = n14697 | n14698 ;
  assign n14700 = n4318 & n8407 ;
  assign n14701 = n3321 & n5975 ;
  assign n14702 = n14700 | n14701 ;
  assign n14703 = n4530 & n6093 ;
  assign n14704 = n5973 & n14703 ;
  assign n14705 = ( n5973 & ~n14702 ) | ( n5973 & n14704 ) | ( ~n14702 & n14704 ) ;
  assign n14706 = n14702 | n14703 ;
  assign n14707 = x33 & x45 ;
  assign n14708 = x34 & x44 ;
  assign n14709 = ( ~n14703 & n14707 ) | ( ~n14703 & n14708 ) | ( n14707 & n14708 ) ;
  assign n14710 = n14707 & n14708 ;
  assign n14711 = ( ~n14702 & n14709 ) | ( ~n14702 & n14710 ) | ( n14709 & n14710 ) ;
  assign n14712 = ~n14706 & n14711 ;
  assign n14713 = n14705 | n14712 ;
  assign n14714 = x30 & x48 ;
  assign n14715 = x31 & x47 ;
  assign n14716 = n14714 | n14715 ;
  assign n14717 = n2965 & n6762 ;
  assign n14718 = n14716 | n14717 ;
  assign n14719 = x20 & x58 ;
  assign n14720 = ( ~n14717 & n14718 ) | ( ~n14717 & n14719 ) | ( n14718 & n14719 ) ;
  assign n14721 = ( n14717 & n14718 ) | ( n14717 & ~n14719 ) | ( n14718 & ~n14719 ) ;
  assign n14722 = ( ~n14718 & n14720 ) | ( ~n14718 & n14721 ) | ( n14720 & n14721 ) ;
  assign n14723 = n14713 & ~n14722 ;
  assign n14724 = ~n14713 & n14722 ;
  assign n14725 = n14723 | n14724 ;
  assign n14726 = x53 & x56 ;
  assign n14727 = n5695 & n14726 ;
  assign n14728 = n1912 & n8355 ;
  assign n14729 = n14727 | n14728 ;
  assign n14730 = n2148 & n8146 ;
  assign n14731 = x53 & n14730 ;
  assign n14732 = ( x53 & ~n14729 ) | ( x53 & n14731 ) | ( ~n14729 & n14731 ) ;
  assign n14733 = x25 & n14732 ;
  assign n14734 = n14729 | n14730 ;
  assign n14735 = x22 & x56 ;
  assign n14736 = ( n13976 & ~n14730 ) | ( n13976 & n14735 ) | ( ~n14730 & n14735 ) ;
  assign n14737 = n13976 & n14735 ;
  assign n14738 = ( ~n14729 & n14736 ) | ( ~n14729 & n14737 ) | ( n14736 & n14737 ) ;
  assign n14739 = ~n14734 & n14738 ;
  assign n14740 = n14733 | n14739 ;
  assign n14741 = n14725 & n14740 ;
  assign n14742 = n14725 | n14740 ;
  assign n14743 = ~n14741 & n14742 ;
  assign n14744 = n14699 & ~n14743 ;
  assign n14745 = ~n14699 & n14743 ;
  assign n14746 = n14744 | n14745 ;
  assign n14747 = n14448 | n14449 ;
  assign n14748 = ( n14448 & n14451 ) | ( n14448 & n14747 ) | ( n14451 & n14747 ) ;
  assign n14749 = n14746 & n14748 ;
  assign n14750 = n14746 | n14748 ;
  assign n14751 = ~n14749 & n14750 ;
  assign n14752 = n14410 | n14436 ;
  assign n14753 = ( n14410 & n14414 ) | ( n14410 & n14752 ) | ( n14414 & n14752 ) ;
  assign n14754 = n14751 & n14753 ;
  assign n14755 = n14751 | n14753 ;
  assign n14756 = ~n14754 & n14755 ;
  assign n14757 = ( n14263 & n14265 ) | ( n14263 & n14456 ) | ( n14265 & n14456 ) ;
  assign n14758 = ( n14454 & n14553 ) | ( n14454 & n14757 ) | ( n14553 & n14757 ) ;
  assign n14759 = n14756 | n14758 ;
  assign n14760 = n14756 & n14758 ;
  assign n14761 = n14759 & ~n14760 ;
  assign n14762 = n14439 | n14556 ;
  assign n14763 = ( n14441 & n14556 ) | ( n14441 & n14762 ) | ( n14556 & n14762 ) ;
  assign n14764 = n14761 & n14763 ;
  assign n14765 = n14443 & n14761 ;
  assign n14766 = ( n14444 & n14764 ) | ( n14444 & n14765 ) | ( n14764 & n14765 ) ;
  assign n14767 = n14761 | n14763 ;
  assign n14768 = n14443 | n14761 ;
  assign n14769 = ( n14444 & n14767 ) | ( n14444 & n14768 ) | ( n14767 & n14768 ) ;
  assign n14770 = ~n14766 & n14769 ;
  assign n14771 = n14371 | n14378 ;
  assign n14772 = n14521 | n14527 ;
  assign n14773 = ( n14183 & n14547 ) | ( n14183 & n14772 ) | ( n14547 & n14772 ) ;
  assign n14774 = n14494 | n14507 ;
  assign n14775 = n14773 | n14774 ;
  assign n14776 = n14494 | n14773 ;
  assign n14777 = ( n14497 & n14775 ) | ( n14497 & n14776 ) | ( n14775 & n14776 ) ;
  assign n14778 = n14773 & n14774 ;
  assign n14779 = n14494 & n14773 ;
  assign n14780 = ( n14497 & n14778 ) | ( n14497 & n14779 ) | ( n14778 & n14779 ) ;
  assign n14781 = n14777 & ~n14780 ;
  assign n14782 = n14344 & n14345 ;
  assign n14783 = ( n14333 & n14344 ) | ( n14333 & n14782 ) | ( n14344 & n14782 ) ;
  assign n14784 = n14332 | n14783 ;
  assign n14785 = n14781 | n14784 ;
  assign n14786 = n14781 & n14784 ;
  assign n14787 = n14785 & ~n14786 ;
  assign n14788 = n14422 | n14428 ;
  assign n14789 = ( n14422 & n14430 ) | ( n14422 & n14788 ) | ( n14430 & n14788 ) ;
  assign n14790 = ( n14431 & n14433 ) | ( n14431 & n14789 ) | ( n14433 & n14789 ) ;
  assign n14791 = n14787 & n14790 ;
  assign n14792 = n14787 | n14790 ;
  assign n14793 = ~n14791 & n14792 ;
  assign n14794 = n14487 | n14501 ;
  assign n14795 = n14487 & n14501 ;
  assign n14796 = n14794 & ~n14795 ;
  assign n14797 = n14313 | n14796 ;
  assign n14798 = n14313 & n14796 ;
  assign n14799 = n14797 & ~n14798 ;
  assign n14800 = n14473 | n14540 ;
  assign n14801 = n14473 & n14540 ;
  assign n14802 = n14800 & ~n14801 ;
  assign n14803 = n14340 | n14802 ;
  assign n14804 = n14340 & n14802 ;
  assign n14805 = n14803 & ~n14804 ;
  assign n14806 = n14233 | n14424 ;
  assign n14807 = ( n14424 & n14425 ) | ( n14424 & n14806 ) | ( n14425 & n14806 ) ;
  assign n14808 = n14805 | n14807 ;
  assign n14809 = n14805 & n14807 ;
  assign n14810 = n14808 & ~n14809 ;
  assign n14811 = n14799 & n14810 ;
  assign n14812 = n14799 | n14810 ;
  assign n14813 = ~n14811 & n14812 ;
  assign n14814 = n14793 & n14813 ;
  assign n14815 = n14793 | n14813 ;
  assign n14816 = ~n14814 & n14815 ;
  assign n14817 = n14373 | n14816 ;
  assign n14818 = n14371 | n14816 ;
  assign n14819 = ( n14771 & n14817 ) | ( n14771 & n14818 ) | ( n14817 & n14818 ) ;
  assign n14820 = n14373 & n14816 ;
  assign n14821 = n14371 & n14816 ;
  assign n14822 = ( n14771 & n14820 ) | ( n14771 & n14821 ) | ( n14820 & n14821 ) ;
  assign n14823 = n14819 & ~n14822 ;
  assign n14824 = ( n14646 & n14770 ) | ( n14646 & ~n14823 ) | ( n14770 & ~n14823 ) ;
  assign n14825 = ( ~n14770 & n14823 ) | ( ~n14770 & n14824 ) | ( n14823 & n14824 ) ;
  assign n14826 = ( ~n14646 & n14824 ) | ( ~n14646 & n14825 ) | ( n14824 & n14825 ) ;
  assign n14827 = n14384 | n14559 ;
  assign n14828 = ( n14384 & n14386 ) | ( n14384 & n14827 ) | ( n14386 & n14827 ) ;
  assign n14829 = ( n14584 & n14826 ) | ( n14584 & ~n14828 ) | ( n14826 & ~n14828 ) ;
  assign n14830 = ( ~n14826 & n14828 ) | ( ~n14826 & n14829 ) | ( n14828 & n14829 ) ;
  assign n14831 = ( ~n14584 & n14829 ) | ( ~n14584 & n14830 ) | ( n14829 & n14830 ) ;
  assign n14832 = n14824 & n14828 ;
  assign n14833 = ~n14646 & n14828 ;
  assign n14834 = ( n14825 & n14832 ) | ( n14825 & n14833 ) | ( n14832 & n14833 ) ;
  assign n14835 = n14824 | n14828 ;
  assign n14836 = n14646 & ~n14828 ;
  assign n14837 = ( n14825 & n14835 ) | ( n14825 & ~n14836 ) | ( n14835 & ~n14836 ) ;
  assign n14838 = n14834 | n14837 ;
  assign n14839 = ( n14582 & n14834 ) | ( n14582 & n14838 ) | ( n14834 & n14838 ) ;
  assign n14840 = ( n14583 & n14834 ) | ( n14583 & n14838 ) | ( n14834 & n14838 ) ;
  assign n14841 = ( n14576 & n14839 ) | ( n14576 & n14840 ) | ( n14839 & n14840 ) ;
  assign n14842 = n1432 & n10975 ;
  assign n14843 = n1437 & n10370 ;
  assign n14844 = n14842 | n14843 ;
  assign n14845 = n1434 & n9831 ;
  assign n14846 = x60 & n14845 ;
  assign n14847 = ( x60 & ~n14844 ) | ( x60 & n14846 ) | ( ~n14844 & n14846 ) ;
  assign n14848 = x19 & n14847 ;
  assign n14849 = n14844 | n14845 ;
  assign n14850 = x20 & x59 ;
  assign n14851 = x21 & x58 ;
  assign n14852 = ( ~n14845 & n14850 ) | ( ~n14845 & n14851 ) | ( n14850 & n14851 ) ;
  assign n14853 = n14850 & n14851 ;
  assign n14854 = ( ~n14844 & n14852 ) | ( ~n14844 & n14853 ) | ( n14852 & n14853 ) ;
  assign n14855 = ~n14849 & n14854 ;
  assign n14856 = n14848 | n14855 ;
  assign n14857 = x29 & x50 ;
  assign n14858 = x30 & x49 ;
  assign n14859 = n14857 | n14858 ;
  assign n14860 = n2709 & n6834 ;
  assign n14861 = x22 & x57 ;
  assign n14862 = ~n14860 & n14861 ;
  assign n14863 = n14859 | n14860 ;
  assign n14864 = ( n14860 & n14862 ) | ( n14860 & n14863 ) | ( n14862 & n14863 ) ;
  assign n14865 = n14859 & ~n14864 ;
  assign n14866 = ~n14859 & n14861 ;
  assign n14867 = ( n14861 & ~n14862 ) | ( n14861 & n14866 ) | ( ~n14862 & n14866 ) ;
  assign n14868 = n14865 | n14867 ;
  assign n14869 = n14856 & n14868 ;
  assign n14870 = n14856 & ~n14869 ;
  assign n14871 = n14868 & ~n14869 ;
  assign n14872 = n14870 | n14871 ;
  assign n14873 = n2683 & n9421 ;
  assign n14874 = n4062 & n6762 ;
  assign n14875 = n14873 | n14874 ;
  assign n14876 = n3321 & n6147 ;
  assign n14877 = x48 & n14876 ;
  assign n14878 = ( x48 & ~n14875 ) | ( x48 & n14877 ) | ( ~n14875 & n14877 ) ;
  assign n14879 = x31 & n14878 ;
  assign n14880 = n14875 | n14876 ;
  assign n14881 = x32 & x47 ;
  assign n14882 = ( n6357 & ~n14876 ) | ( n6357 & n14881 ) | ( ~n14876 & n14881 ) ;
  assign n14883 = n6357 & n14881 ;
  assign n14884 = ( ~n14875 & n14882 ) | ( ~n14875 & n14883 ) | ( n14882 & n14883 ) ;
  assign n14885 = ~n14880 & n14884 ;
  assign n14886 = n14879 | n14885 ;
  assign n14887 = ~n14872 & n14886 ;
  assign n14888 = n14872 & ~n14886 ;
  assign n14889 = n14887 | n14888 ;
  assign n14890 = n2340 & n8360 ;
  assign n14891 = n1912 & n8357 ;
  assign n14892 = n14890 | n14891 ;
  assign n14893 = n2511 & n8355 ;
  assign n14894 = x55 & n14893 ;
  assign n14895 = ( x55 & ~n14892 ) | ( x55 & n14894 ) | ( ~n14892 & n14894 ) ;
  assign n14896 = x24 & n14895 ;
  assign n14897 = n14892 | n14893 ;
  assign n14898 = x25 & x54 ;
  assign n14899 = x26 & x53 ;
  assign n14900 = ( ~n14893 & n14898 ) | ( ~n14893 & n14899 ) | ( n14898 & n14899 ) ;
  assign n14901 = n14898 & n14899 ;
  assign n14902 = ( ~n14892 & n14900 ) | ( ~n14892 & n14901 ) | ( n14900 & n14901 ) ;
  assign n14903 = ~n14897 & n14902 ;
  assign n14904 = n14896 | n14903 ;
  assign n14905 = x37 & x42 ;
  assign n14906 = n4555 & n14905 ;
  assign n14907 = n4857 & n5710 ;
  assign n14908 = n14906 | n14907 ;
  assign n14909 = n5392 & n5813 ;
  assign n14910 = n14905 & n14909 ;
  assign n14911 = ( n14905 & ~n14908 ) | ( n14905 & n14910 ) | ( ~n14908 & n14910 ) ;
  assign n14912 = n14908 | n14909 ;
  assign n14913 = x38 & x41 ;
  assign n14914 = ( n4555 & ~n14909 ) | ( n4555 & n14913 ) | ( ~n14909 & n14913 ) ;
  assign n14915 = n4555 & n14913 ;
  assign n14916 = ( ~n14908 & n14914 ) | ( ~n14908 & n14915 ) | ( n14914 & n14915 ) ;
  assign n14917 = ~n14912 & n14916 ;
  assign n14918 = n14911 | n14917 ;
  assign n14919 = n14904 & n14918 ;
  assign n14920 = n14904 & ~n14919 ;
  assign n14921 = x17 & x62 ;
  assign n14922 = x40 | n14921 ;
  assign n14923 = x40 & x62 ;
  assign n14924 = ~x17 & x51 ;
  assign n14925 = ( x51 & ~n14923 ) | ( x51 & n14924 ) | ( ~n14923 & n14924 ) ;
  assign n14926 = ( x28 & x40 ) | ( x28 & n14921 ) | ( x40 & n14921 ) ;
  assign n14927 = x40 & n14921 ;
  assign n14928 = ( n14925 & n14926 ) | ( n14925 & n14927 ) | ( n14926 & n14927 ) ;
  assign n14929 = n14922 & ~n14928 ;
  assign n14930 = x28 & n14925 ;
  assign n14931 = ~x40 & x51 ;
  assign n14932 = ~n14921 & n14931 ;
  assign n14933 = x28 & n14932 ;
  assign n14934 = x28 & x51 ;
  assign n14935 = ( ~n14930 & n14933 ) | ( ~n14930 & n14934 ) | ( n14933 & n14934 ) ;
  assign n14936 = n14929 | n14935 ;
  assign n14937 = ~n14904 & n14918 ;
  assign n14938 = n14936 & n14937 ;
  assign n14939 = ( n14920 & n14936 ) | ( n14920 & n14938 ) | ( n14936 & n14938 ) ;
  assign n14940 = n14936 | n14937 ;
  assign n14941 = n14920 | n14940 ;
  assign n14942 = ~n14939 & n14941 ;
  assign n14943 = n14889 | n14942 ;
  assign n14944 = n14889 & n14942 ;
  assign n14945 = n14943 & ~n14944 ;
  assign n14946 = n14799 | n14809 ;
  assign n14947 = ( n14809 & n14810 ) | ( n14809 & n14946 ) | ( n14810 & n14946 ) ;
  assign n14948 = n14945 & n14947 ;
  assign n14949 = n14945 | n14947 ;
  assign n14950 = ~n14948 & n14949 ;
  assign n14951 = ( n14787 & n14790 ) | ( n14787 & n14813 ) | ( n14790 & n14813 ) ;
  assign n14952 = n14950 | n14951 ;
  assign n14953 = n14950 & n14951 ;
  assign n14954 = n14952 & ~n14953 ;
  assign n14955 = n14340 | n14801 ;
  assign n14956 = ( n14801 & n14802 ) | ( n14801 & n14955 ) | ( n14802 & n14955 ) ;
  assign n14957 = n14313 | n14795 ;
  assign n14958 = ( n14795 & n14796 ) | ( n14795 & n14957 ) | ( n14796 & n14957 ) ;
  assign n14959 = n14956 | n14958 ;
  assign n14960 = n14956 & n14958 ;
  assign n14961 = n14959 & ~n14960 ;
  assign n14962 = n14678 | n14696 ;
  assign n14963 = ( n14678 & n14681 ) | ( n14678 & n14962 ) | ( n14681 & n14962 ) ;
  assign n14964 = n14961 | n14963 ;
  assign n14965 = n14961 & n14963 ;
  assign n14966 = n14964 & ~n14965 ;
  assign n14967 = n14780 | n14784 ;
  assign n14968 = ( n14780 & n14781 ) | ( n14780 & n14967 ) | ( n14781 & n14967 ) ;
  assign n14969 = n14966 | n14968 ;
  assign n14970 = n14966 & n14968 ;
  assign n14971 = n14969 & ~n14970 ;
  assign n14972 = n14620 | n14634 ;
  assign n14973 = ( n14634 & n14635 ) | ( n14634 & n14972 ) | ( n14635 & n14972 ) ;
  assign n14974 = n14971 & n14973 ;
  assign n14975 = n14971 | n14973 ;
  assign n14976 = ~n14974 & n14975 ;
  assign n14977 = n14954 & n14976 ;
  assign n14978 = n14954 | n14976 ;
  assign n14979 = ~n14977 & n14978 ;
  assign n14980 = n14646 | n14822 ;
  assign n14981 = ( n14822 & n14823 ) | ( n14822 & n14980 ) | ( n14823 & n14980 ) ;
  assign n14982 = n14979 & ~n14981 ;
  assign n14983 = n14655 | n14670 ;
  assign n14984 = n14655 & n14670 ;
  assign n14985 = n14983 & ~n14984 ;
  assign n14986 = n14734 | n14985 ;
  assign n14987 = n14734 & n14985 ;
  assign n14988 = n14986 & ~n14987 ;
  assign n14989 = n14611 & n14988 ;
  assign n14990 = ( n14617 & n14988 ) | ( n14617 & n14989 ) | ( n14988 & n14989 ) ;
  assign n14991 = n14611 | n14988 ;
  assign n14992 = n14617 | n14991 ;
  assign n14993 = ~n14990 & n14992 ;
  assign n14994 = x23 & x56 ;
  assign n14995 = x27 & x52 ;
  assign n14996 = n14994 | n14995 ;
  assign n14997 = x27 & x56 ;
  assign n14998 = n13902 & n14997 ;
  assign n14999 = x36 & x43 ;
  assign n15000 = ~n14998 & n14999 ;
  assign n15001 = n14996 | n14998 ;
  assign n15002 = ( n14998 & n15000 ) | ( n14998 & n15001 ) | ( n15000 & n15001 ) ;
  assign n15003 = n14996 & ~n15002 ;
  assign n15004 = ~n14996 & n14999 ;
  assign n15005 = ( n14999 & ~n15000 ) | ( n14999 & n15004 ) | ( ~n15000 & n15004 ) ;
  assign n15006 = n15003 | n15005 ;
  assign n15007 = x34 & x45 ;
  assign n15008 = x35 & x44 ;
  assign n15009 = n15007 | n15008 ;
  assign n15010 = n3483 & n6093 ;
  assign n15011 = n15009 | n15010 ;
  assign n15012 = x16 & x63 ;
  assign n15013 = ( ~n15010 & n15011 ) | ( ~n15010 & n15012 ) | ( n15011 & n15012 ) ;
  assign n15014 = ( n15010 & n15011 ) | ( n15010 & ~n15012 ) | ( n15011 & ~n15012 ) ;
  assign n15015 = ( ~n15011 & n15013 ) | ( ~n15011 & n15014 ) | ( n15013 & n15014 ) ;
  assign n15016 = n15006 & n15015 ;
  assign n15017 = n15006 & ~n15016 ;
  assign n15018 = n14622 | n14629 ;
  assign n15019 = ~n15006 & n15015 ;
  assign n15020 = n15018 & n15019 ;
  assign n15021 = ( n15017 & n15018 ) | ( n15017 & n15020 ) | ( n15018 & n15020 ) ;
  assign n15022 = n15018 | n15019 ;
  assign n15023 = n15017 | n15022 ;
  assign n15024 = ~n15021 & n15023 ;
  assign n15025 = n14993 & n15024 ;
  assign n15026 = n14993 | n15024 ;
  assign n15027 = ~n15025 & n15026 ;
  assign n15028 = ( n14699 & n14743 ) | ( n14699 & n14748 ) | ( n14743 & n14748 ) ;
  assign n15029 = n15027 | n15028 ;
  assign n15030 = n15027 & n15028 ;
  assign n15031 = n15029 & ~n15030 ;
  assign n15032 = ~n14596 & n14598 ;
  assign n15033 = ( n14596 & n14597 ) | ( n14596 & n15032 ) | ( n14597 & n15032 ) ;
  assign n15034 = x18 & x61 ;
  assign n15035 = n14603 & n15034 ;
  assign n15036 = ( n14606 & n15034 ) | ( n14606 & n15035 ) | ( n15034 & n15035 ) ;
  assign n15037 = n14603 | n15034 ;
  assign n15038 = n14606 | n15037 ;
  assign n15039 = ~n15036 & n15038 ;
  assign n15040 = n15033 | n15039 ;
  assign n15041 = n15033 & n15039 ;
  assign n15042 = n15040 & ~n15041 ;
  assign n15043 = ~n14717 & n14719 ;
  assign n15044 = ( n14717 & n14718 ) | ( n14717 & n15043 ) | ( n14718 & n15043 ) ;
  assign n15045 = n14689 | n15044 ;
  assign n15046 = n14689 & n15044 ;
  assign n15047 = n15045 & ~n15046 ;
  assign n15048 = n14706 | n15047 ;
  assign n15049 = n14706 & n15047 ;
  assign n15050 = n15048 & ~n15049 ;
  assign n15051 = n15042 & n15050 ;
  assign n15052 = n15042 | n15050 ;
  assign n15053 = ~n15051 & n15052 ;
  assign n15054 = n14713 & n14722 ;
  assign n15055 = n14740 | n15054 ;
  assign n15056 = ( n14725 & n15054 ) | ( n14725 & n15055 ) | ( n15054 & n15055 ) ;
  assign n15057 = n15053 & n15056 ;
  assign n15058 = n15053 | n15056 ;
  assign n15059 = ~n15057 & n15058 ;
  assign n15060 = n15031 & n15059 ;
  assign n15061 = n15031 | n15059 ;
  assign n15062 = ~n15060 & n15061 ;
  assign n15063 = n14589 & n15062 ;
  assign n15064 = ( n14642 & n15062 ) | ( n14642 & n15063 ) | ( n15062 & n15063 ) ;
  assign n15065 = n14589 | n15062 ;
  assign n15066 = n14642 | n15065 ;
  assign n15067 = ~n15064 & n15066 ;
  assign n15068 = n14754 | n14758 ;
  assign n15069 = ( n14754 & n14756 ) | ( n14754 & n15068 ) | ( n14756 & n15068 ) ;
  assign n15070 = n15067 | n15069 ;
  assign n15071 = n15067 & n15069 ;
  assign n15072 = n15070 & ~n15071 ;
  assign n15073 = n14979 & n14981 ;
  assign n15074 = n14981 | n15072 ;
  assign n15075 = ( n15072 & ~n15073 ) | ( n15072 & n15074 ) | ( ~n15073 & n15074 ) ;
  assign n15076 = n14982 | n15075 ;
  assign n15077 = ( n14981 & n14982 ) | ( n14981 & n15072 ) | ( n14982 & n15072 ) ;
  assign n15078 = ( ~n14979 & n14982 ) | ( ~n14979 & n15077 ) | ( n14982 & n15077 ) ;
  assign n15079 = n15076 & ~n15078 ;
  assign n15080 = n14646 & n14823 ;
  assign n15081 = n14646 | n14823 ;
  assign n15082 = ~n15080 & n15081 ;
  assign n15083 = n14766 | n15082 ;
  assign n15084 = ( n14766 & n14770 ) | ( n14766 & n15083 ) | ( n14770 & n15083 ) ;
  assign n15085 = ( n14841 & n15079 ) | ( n14841 & ~n15084 ) | ( n15079 & ~n15084 ) ;
  assign n15086 = ( ~n15079 & n15084 ) | ( ~n15079 & n15085 ) | ( n15084 & n15085 ) ;
  assign n15087 = ( ~n14841 & n15085 ) | ( ~n14841 & n15086 ) | ( n15085 & n15086 ) ;
  assign n15088 = x54 & x57 ;
  assign n15089 = n2336 & n15088 ;
  assign n15090 = n1686 & n8903 ;
  assign n15091 = n15089 | n15090 ;
  assign n15092 = n2340 & n8146 ;
  assign n15093 = x57 & n15092 ;
  assign n15094 = ( x57 & ~n15091 ) | ( x57 & n15093 ) | ( ~n15091 & n15093 ) ;
  assign n15095 = x23 & n15094 ;
  assign n15096 = n15091 | n15092 ;
  assign n15097 = x24 & x56 ;
  assign n15098 = x26 & x54 ;
  assign n15099 = ( ~n15092 & n15097 ) | ( ~n15092 & n15098 ) | ( n15097 & n15098 ) ;
  assign n15100 = n15097 & n15098 ;
  assign n15101 = ( ~n15091 & n15099 ) | ( ~n15091 & n15100 ) | ( n15099 & n15100 ) ;
  assign n15102 = ~n15096 & n15101 ;
  assign n15103 = n15095 | n15102 ;
  assign n15104 = x37 & x43 ;
  assign n15105 = x38 & x42 ;
  assign n15106 = n15104 | n15105 ;
  assign n15107 = n4857 & n5407 ;
  assign n15108 = x25 & x55 ;
  assign n15109 = ~n15107 & n15108 ;
  assign n15110 = n15106 | n15107 ;
  assign n15111 = ( n15107 & n15109 ) | ( n15107 & n15110 ) | ( n15109 & n15110 ) ;
  assign n15112 = n15106 & ~n15111 ;
  assign n15113 = ~n15106 & n15108 ;
  assign n15114 = ( n15108 & ~n15109 ) | ( n15108 & n15113 ) | ( ~n15109 & n15113 ) ;
  assign n15115 = n15112 | n15114 ;
  assign n15116 = n15103 & n15115 ;
  assign n15117 = n15103 & ~n15116 ;
  assign n15118 = n15115 & ~n15116 ;
  assign n15119 = n15117 | n15118 ;
  assign n15120 = x27 & x53 ;
  assign n15121 = x28 & x52 ;
  assign n15122 = n15120 | n15121 ;
  assign n15123 = n2372 & n8161 ;
  assign n15124 = n4350 & ~n15123 ;
  assign n15125 = n15122 | n15123 ;
  assign n15126 = ( n15123 & n15124 ) | ( n15123 & n15125 ) | ( n15124 & n15125 ) ;
  assign n15127 = n15122 & ~n15126 ;
  assign n15128 = n4350 & ~n15122 ;
  assign n15129 = ( n4350 & ~n15124 ) | ( n4350 & n15128 ) | ( ~n15124 & n15128 ) ;
  assign n15130 = n15127 | n15129 ;
  assign n15131 = n1585 & n9831 ;
  assign n15132 = n1710 & n10975 ;
  assign n15133 = n1434 & n10370 ;
  assign n15134 = n15132 | n15133 ;
  assign n15135 = ~n15131 & n15134 ;
  assign n15136 = x21 & x59 ;
  assign n15137 = x22 & x58 ;
  assign n15138 = n15136 | n15137 ;
  assign n15139 = ~n15131 & n15138 ;
  assign n15140 = x20 & x60 ;
  assign n15141 = n15139 | n15140 ;
  assign n15142 = ~n15135 & n15141 ;
  assign n15143 = n14912 & n15142 ;
  assign n15144 = n14912 | n15142 ;
  assign n15145 = ~n15143 & n15144 ;
  assign n15146 = n2546 & n6345 ;
  assign n15147 = n2965 & n6834 ;
  assign n15148 = n15146 | n15147 ;
  assign n15149 = n4062 & n6759 ;
  assign n15150 = x50 & n15149 ;
  assign n15151 = ( x50 & ~n15148 ) | ( x50 & n15150 ) | ( ~n15148 & n15150 ) ;
  assign n15152 = x30 & n15151 ;
  assign n15153 = n15148 | n15149 ;
  assign n15154 = x31 & x49 ;
  assign n15155 = x32 & x48 ;
  assign n15156 = ( ~n15149 & n15154 ) | ( ~n15149 & n15155 ) | ( n15154 & n15155 ) ;
  assign n15157 = n15154 & n15155 ;
  assign n15158 = ( ~n15148 & n15156 ) | ( ~n15148 & n15157 ) | ( n15156 & n15157 ) ;
  assign n15159 = ~n15153 & n15158 ;
  assign n15160 = n15152 | n15159 ;
  assign n15161 = ~n15145 & n15160 ;
  assign n15162 = n15145 & ~n15160 ;
  assign n15163 = n15161 | n15162 ;
  assign n15164 = ( n15119 & ~n15130 ) | ( n15119 & n15163 ) | ( ~n15130 & n15163 ) ;
  assign n15165 = ( ~n15119 & n15130 ) | ( ~n15119 & n15164 ) | ( n15130 & n15164 ) ;
  assign n15166 = n4914 & n8407 ;
  assign n15167 = n3483 & n5975 ;
  assign n15168 = n15166 | n15167 ;
  assign n15169 = n4078 & n6093 ;
  assign n15170 = x46 & n15169 ;
  assign n15171 = ( x46 & ~n15168 ) | ( x46 & n15170 ) | ( ~n15168 & n15170 ) ;
  assign n15172 = x34 & n15171 ;
  assign n15173 = n15168 | n15169 ;
  assign n15174 = ( n6308 & n6396 ) | ( n6308 & ~n15169 ) | ( n6396 & ~n15169 ) ;
  assign n15175 = n6308 & n6396 ;
  assign n15176 = ( ~n15168 & n15174 ) | ( ~n15168 & n15175 ) | ( n15174 & n15175 ) ;
  assign n15177 = ~n15173 & n15176 ;
  assign n15178 = n15172 | n15177 ;
  assign n15179 = x17 & x63 ;
  assign n15180 = x29 & x51 ;
  assign n15181 = n15179 | n15180 ;
  assign n15182 = x29 & x63 ;
  assign n15183 = n8437 & n15182 ;
  assign n15184 = n15181 | n15183 ;
  assign n15185 = x33 & x47 ;
  assign n15186 = ( ~n15183 & n15184 ) | ( ~n15183 & n15185 ) | ( n15184 & n15185 ) ;
  assign n15187 = ( n15183 & n15184 ) | ( n15183 & ~n15185 ) | ( n15184 & ~n15185 ) ;
  assign n15188 = ( ~n15184 & n15186 ) | ( ~n15184 & n15187 ) | ( n15186 & n15187 ) ;
  assign n15189 = n15178 & n15188 ;
  assign n15190 = n15178 & ~n15189 ;
  assign n15191 = n1077 & n10684 ;
  assign n15192 = x19 & x61 ;
  assign n15193 = x18 & x62 ;
  assign n15194 = n15192 | n15193 ;
  assign n15195 = ~n15191 & n15194 ;
  assign n15196 = n14928 & n15195 ;
  assign n15197 = n14928 & ~n15196 ;
  assign n15198 = n15195 & ~n15196 ;
  assign n15199 = n15197 | n15198 ;
  assign n15200 = ~n15178 & n15188 ;
  assign n15201 = ~n15199 & n15200 ;
  assign n15202 = ( n15190 & ~n15199 ) | ( n15190 & n15201 ) | ( ~n15199 & n15201 ) ;
  assign n15203 = n15199 & ~n15200 ;
  assign n15204 = ~n15190 & n15203 ;
  assign n15205 = n15202 | n15204 ;
  assign n15206 = n15164 & n15205 ;
  assign n15207 = ~n15163 & n15205 ;
  assign n15208 = ( n15165 & n15206 ) | ( n15165 & n15207 ) | ( n15206 & n15207 ) ;
  assign n15209 = n15164 | n15205 ;
  assign n15210 = n15163 & ~n15205 ;
  assign n15211 = ( n15165 & n15209 ) | ( n15165 & ~n15210 ) | ( n15209 & ~n15210 ) ;
  assign n15212 = ~n15208 & n15211 ;
  assign n15213 = n14970 | n14973 ;
  assign n15214 = ( n14970 & n14971 ) | ( n14970 & n15213 ) | ( n14971 & n15213 ) ;
  assign n15215 = n15212 & n15214 ;
  assign n15216 = n15212 | n15214 ;
  assign n15217 = ~n15215 & n15216 ;
  assign n15218 = ( n15027 & n15028 ) | ( n15027 & n15059 ) | ( n15028 & n15059 ) ;
  assign n15219 = n15217 | n15218 ;
  assign n15220 = n15217 & n15218 ;
  assign n15221 = n15219 & ~n15220 ;
  assign n15222 = n15064 | n15069 ;
  assign n15223 = ( n15064 & n15067 ) | ( n15064 & n15222 ) | ( n15067 & n15222 ) ;
  assign n15224 = n15221 | n15223 ;
  assign n15225 = n15221 & n15223 ;
  assign n15226 = n15224 & ~n15225 ;
  assign n15227 = ~n15010 & n15012 ;
  assign n15228 = ( n15010 & n15011 ) | ( n15010 & n15227 ) | ( n15011 & n15227 ) ;
  assign n15229 = n14897 | n15228 ;
  assign n15230 = n14897 & n15228 ;
  assign n15231 = n15229 & ~n15230 ;
  assign n15232 = n15002 | n15231 ;
  assign n15233 = n15002 & n15231 ;
  assign n15234 = n15232 & ~n15233 ;
  assign n15235 = n15016 | n15234 ;
  assign n15236 = n15021 | n15235 ;
  assign n15237 = n15016 & n15234 ;
  assign n15238 = ( n15021 & n15234 ) | ( n15021 & n15237 ) | ( n15234 & n15237 ) ;
  assign n15239 = n15236 & ~n15238 ;
  assign n15240 = n14960 | n14961 ;
  assign n15241 = ( n14960 & n14963 ) | ( n14960 & n15240 ) | ( n14963 & n15240 ) ;
  assign n15242 = n15239 | n15241 ;
  assign n15243 = n15239 & n15241 ;
  assign n15244 = n15242 & ~n15243 ;
  assign n15245 = ( n14889 & n14942 ) | ( n14889 & n14947 ) | ( n14942 & n14947 ) ;
  assign n15246 = n15244 | n15245 ;
  assign n15247 = n15244 & n15245 ;
  assign n15248 = n15246 & ~n15247 ;
  assign n15249 = n14849 | n14864 ;
  assign n15250 = n14849 & n14864 ;
  assign n15251 = n15249 & ~n15250 ;
  assign n15252 = n14880 | n15251 ;
  assign n15253 = n14880 & n15251 ;
  assign n15254 = n15252 & ~n15253 ;
  assign n15255 = n14919 | n14939 ;
  assign n15256 = n14869 | n14886 ;
  assign n15257 = ( n14869 & n14872 ) | ( n14869 & n15256 ) | ( n14872 & n15256 ) ;
  assign n15258 = n15255 | n15257 ;
  assign n15259 = n15255 & n15257 ;
  assign n15260 = n15258 & ~n15259 ;
  assign n15261 = n15254 & n15260 ;
  assign n15262 = n15254 | n15260 ;
  assign n15263 = ~n15261 & n15262 ;
  assign n15264 = n15248 & n15263 ;
  assign n15265 = n15248 | n15263 ;
  assign n15266 = ~n15264 & n15265 ;
  assign n15279 = n15051 | n15056 ;
  assign n15280 = ( n15051 & n15053 ) | ( n15051 & n15279 ) | ( n15053 & n15279 ) ;
  assign n15267 = n14734 | n14984 ;
  assign n15268 = ( n14984 & n14985 ) | ( n14984 & n15267 ) | ( n14985 & n15267 ) ;
  assign n15269 = n14706 | n15046 ;
  assign n15270 = ( n15046 & n15047 ) | ( n15046 & n15269 ) | ( n15047 & n15269 ) ;
  assign n15271 = n15268 | n15270 ;
  assign n15272 = n15268 & n15270 ;
  assign n15273 = n15271 & ~n15272 ;
  assign n15274 = n15033 | n15036 ;
  assign n15275 = ( n15036 & n15039 ) | ( n15036 & n15274 ) | ( n15039 & n15274 ) ;
  assign n15276 = n15273 | n15275 ;
  assign n15277 = n15273 & n15275 ;
  assign n15278 = n15276 & ~n15277 ;
  assign n15281 = n14990 | n15024 ;
  assign n15282 = ( n14990 & n14993 ) | ( n14990 & n15281 ) | ( n14993 & n15281 ) ;
  assign n15283 = ( n15278 & n15280 ) | ( n15278 & ~n15282 ) | ( n15280 & ~n15282 ) ;
  assign n15284 = ( ~n15278 & n15282 ) | ( ~n15278 & n15283 ) | ( n15282 & n15283 ) ;
  assign n15285 = ( ~n15280 & n15283 ) | ( ~n15280 & n15284 ) | ( n15283 & n15284 ) ;
  assign n15286 = n15266 & n15285 ;
  assign n15287 = n15266 & ~n15286 ;
  assign n15288 = ~n15266 & n15285 ;
  assign n15289 = n14953 | n14976 ;
  assign n15290 = ( n14953 & n14954 ) | ( n14953 & n15289 ) | ( n14954 & n15289 ) ;
  assign n15291 = n15288 | n15290 ;
  assign n15292 = n15287 | n15291 ;
  assign n15293 = n15288 & n15290 ;
  assign n15294 = ( n15287 & n15290 ) | ( n15287 & n15293 ) | ( n15290 & n15293 ) ;
  assign n15295 = n15292 & ~n15294 ;
  assign n15296 = n15226 & n15295 ;
  assign n15297 = n15226 | n15295 ;
  assign n15298 = ~n15296 & n15297 ;
  assign n15299 = n14982 | n15073 ;
  assign n15300 = ( ~n14982 & n15077 ) | ( ~n14982 & n15299 ) | ( n15077 & n15299 ) ;
  assign n15301 = n15298 | n15300 ;
  assign n15302 = n15298 & n15300 ;
  assign n15303 = n15301 & ~n15302 ;
  assign n15304 = n15079 & n15084 ;
  assign n15305 = n15079 | n15084 ;
  assign n15306 = n14840 & n15305 ;
  assign n15307 = n15304 | n15306 ;
  assign n15308 = n15304 | n15305 ;
  assign n15309 = ( n14839 & n15304 ) | ( n14839 & n15308 ) | ( n15304 & n15308 ) ;
  assign n15310 = ( n14576 & n15307 ) | ( n14576 & n15309 ) | ( n15307 & n15309 ) ;
  assign n15311 = n15303 | n15310 ;
  assign n15312 = n15301 & n15308 ;
  assign n15313 = n15301 & n15304 ;
  assign n15314 = ( n14839 & n15312 ) | ( n14839 & n15313 ) | ( n15312 & n15313 ) ;
  assign n15315 = ( n15301 & n15306 ) | ( n15301 & n15313 ) | ( n15306 & n15313 ) ;
  assign n15316 = ( n14576 & n15314 ) | ( n14576 & n15315 ) | ( n15314 & n15315 ) ;
  assign n15317 = ~n15302 & n15316 ;
  assign n15318 = n15311 & ~n15317 ;
  assign n15319 = n15301 | n15302 ;
  assign n15320 = ( n15302 & n15304 ) | ( n15302 & n15319 ) | ( n15304 & n15319 ) ;
  assign n15321 = ( n15305 & n15319 ) | ( n15305 & n15320 ) | ( n15319 & n15320 ) ;
  assign n15322 = n15319 & n15320 ;
  assign n15323 = ( n14840 & n15321 ) | ( n14840 & n15322 ) | ( n15321 & n15322 ) ;
  assign n15324 = ( n15302 & n15308 ) | ( n15302 & n15319 ) | ( n15308 & n15319 ) ;
  assign n15325 = ( n14838 & n15320 ) | ( n14838 & n15324 ) | ( n15320 & n15324 ) ;
  assign n15326 = ( n14834 & n15320 ) | ( n14834 & n15324 ) | ( n15320 & n15324 ) ;
  assign n15327 = ( n14582 & n15325 ) | ( n14582 & n15326 ) | ( n15325 & n15326 ) ;
  assign n15328 = ( n14576 & n15323 ) | ( n14576 & n15327 ) | ( n15323 & n15327 ) ;
  assign n15329 = n15286 | n15294 ;
  assign n15330 = ( n15244 & n15245 ) | ( n15244 & n15263 ) | ( n15245 & n15263 ) ;
  assign n15331 = n15280 & n15282 ;
  assign n15332 = n15282 & ~n15331 ;
  assign n15333 = n15278 & n15280 ;
  assign n15334 = ~n15282 & n15333 ;
  assign n15335 = ( n15278 & n15332 ) | ( n15278 & n15334 ) | ( n15332 & n15334 ) ;
  assign n15336 = x56 & x59 ;
  assign n15337 = n5695 & n15336 ;
  assign n15338 = n1932 & n9831 ;
  assign n15339 = n15337 | n15338 ;
  assign n15340 = n1557 & n8708 ;
  assign n15341 = x59 & n15340 ;
  assign n15342 = ( x59 & ~n15339 ) | ( x59 & n15341 ) | ( ~n15339 & n15341 ) ;
  assign n15343 = x22 & n15342 ;
  assign n15344 = n15339 | n15340 ;
  assign n15345 = x23 & x58 ;
  assign n15346 = ( n13576 & ~n15340 ) | ( n13576 & n15345 ) | ( ~n15340 & n15345 ) ;
  assign n15347 = n13576 & n15345 ;
  assign n15348 = ( ~n15339 & n15346 ) | ( ~n15339 & n15347 ) | ( n15346 & n15347 ) ;
  assign n15349 = ~n15344 & n15348 ;
  assign n15350 = n15343 | n15349 ;
  assign n15351 = ( x41 & x62 ) | ( x41 & ~n5813 ) | ( x62 & ~n5813 ) ;
  assign n15352 = x19 | x62 ;
  assign n15353 = ~x19 & x41 ;
  assign n15354 = ( n5813 & n15352 ) | ( n5813 & ~n15353 ) | ( n15352 & ~n15353 ) ;
  assign n15355 = ( ~x19 & x41 ) | ( ~x19 & x62 ) | ( x41 & x62 ) ;
  assign n15356 = ( x19 & n5813 ) | ( x19 & ~n15355 ) | ( n5813 & ~n15355 ) ;
  assign n15357 = ( n15351 & ~n15354 ) | ( n15351 & n15356 ) | ( ~n15354 & n15356 ) ;
  assign n15358 = n15350 & n15357 ;
  assign n15359 = n15350 & ~n15358 ;
  assign n15360 = x33 & x48 ;
  assign n15361 = x34 & x47 ;
  assign n15362 = n15360 | n15361 ;
  assign n15363 = n4530 & n6762 ;
  assign n15364 = n11163 & ~n15363 ;
  assign n15365 = n15362 | n15363 ;
  assign n15366 = ( n15363 & n15364 ) | ( n15363 & n15365 ) | ( n15364 & n15365 ) ;
  assign n15367 = n15362 & ~n15366 ;
  assign n15368 = n11163 & ~n15362 ;
  assign n15369 = ( n11163 & ~n15364 ) | ( n11163 & n15368 ) | ( ~n15364 & n15368 ) ;
  assign n15370 = n15367 | n15369 ;
  assign n15371 = ~n15350 & n15357 ;
  assign n15372 = n15370 & n15371 ;
  assign n15373 = ( n15359 & n15370 ) | ( n15359 & n15372 ) | ( n15370 & n15372 ) ;
  assign n15374 = n15370 | n15371 ;
  assign n15375 = n15359 | n15374 ;
  assign n15376 = ~n15373 & n15375 ;
  assign n15377 = n15272 | n15275 ;
  assign n15378 = ( n15272 & n15273 ) | ( n15272 & n15377 ) | ( n15273 & n15377 ) ;
  assign n15379 = n15376 | n15378 ;
  assign n15380 = n15376 & n15378 ;
  assign n15381 = n15379 & ~n15380 ;
  assign n15382 = n3850 & n12770 ;
  assign n15383 = n1285 & n10856 ;
  assign n15384 = n15382 | n15383 ;
  assign n15385 = n1434 & n10367 ;
  assign n15386 = x63 & n15385 ;
  assign n15387 = ( x63 & ~n15384 ) | ( x63 & n15386 ) | ( ~n15384 & n15386 ) ;
  assign n15388 = x18 & n15387 ;
  assign n15389 = n15384 | n15385 ;
  assign n15390 = x20 & x61 ;
  assign n15391 = x21 & x60 ;
  assign n15392 = ( ~n15385 & n15390 ) | ( ~n15385 & n15391 ) | ( n15390 & n15391 ) ;
  assign n15393 = n15390 & n15391 ;
  assign n15394 = ( ~n15384 & n15392 ) | ( ~n15384 & n15393 ) | ( n15392 & n15393 ) ;
  assign n15395 = ~n15389 & n15394 ;
  assign n15396 = n15388 | n15395 ;
  assign n15397 = x35 & x46 ;
  assign n15398 = n4078 & n5975 ;
  assign n15399 = x37 & x44 ;
  assign n15400 = n15397 & n15399 ;
  assign n15401 = n15398 | n15400 ;
  assign n15402 = n3770 & n6093 ;
  assign n15403 = n15397 & n15402 ;
  assign n15404 = ( n15397 & ~n15401 ) | ( n15397 & n15403 ) | ( ~n15401 & n15403 ) ;
  assign n15405 = n15401 | n15402 ;
  assign n15406 = x36 & x45 ;
  assign n15407 = ( n15399 & ~n15402 ) | ( n15399 & n15406 ) | ( ~n15402 & n15406 ) ;
  assign n15408 = n15399 & n15406 ;
  assign n15409 = ( ~n15401 & n15407 ) | ( ~n15401 & n15408 ) | ( n15407 & n15408 ) ;
  assign n15410 = ~n15405 & n15409 ;
  assign n15411 = n15404 | n15410 ;
  assign n15412 = n15396 & n15411 ;
  assign n15413 = n15396 & ~n15412 ;
  assign n15414 = x29 & n14602 ;
  assign n15415 = x53 & n2895 ;
  assign n15416 = n15414 | n15415 ;
  assign n15417 = n2369 & n8161 ;
  assign n15418 = x55 & ~n15417 ;
  assign n15419 = n15416 & n15418 ;
  assign n15420 = x26 & x55 ;
  assign n15421 = ~n15419 & n15420 ;
  assign n15422 = n15417 | n15419 ;
  assign n15423 = x28 & x53 ;
  assign n15424 = x29 & x52 ;
  assign n15425 = ( ~n15417 & n15423 ) | ( ~n15417 & n15424 ) | ( n15423 & n15424 ) ;
  assign n15426 = n15423 & n15424 ;
  assign n15427 = ( ~n15419 & n15425 ) | ( ~n15419 & n15426 ) | ( n15425 & n15426 ) ;
  assign n15428 = ~n15422 & n15427 ;
  assign n15429 = n15421 | n15428 ;
  assign n15430 = ~n15396 & n15411 ;
  assign n15431 = n15429 & n15430 ;
  assign n15432 = ( n15413 & n15429 ) | ( n15413 & n15431 ) | ( n15429 & n15431 ) ;
  assign n15433 = n15429 | n15430 ;
  assign n15434 = n15413 | n15433 ;
  assign n15435 = ~n15432 & n15434 ;
  assign n15436 = n15381 | n15435 ;
  assign n15437 = n15381 & n15435 ;
  assign n15438 = n15436 & ~n15437 ;
  assign n15439 = n15331 & n15438 ;
  assign n15440 = ( n15335 & n15438 ) | ( n15335 & n15439 ) | ( n15438 & n15439 ) ;
  assign n15441 = n15331 | n15334 ;
  assign n15442 = n15278 | n15280 ;
  assign n15443 = ( n15278 & n15282 ) | ( n15278 & n15442 ) | ( n15282 & n15442 ) ;
  assign n15444 = ( n15332 & n15441 ) | ( n15332 & n15443 ) | ( n15441 & n15443 ) ;
  assign n15445 = n15438 | n15444 ;
  assign n15446 = ~n15440 & n15445 ;
  assign n15447 = n15330 & ~n15446 ;
  assign n15448 = n15330 & n15446 ;
  assign n15449 = n15446 & ~n15448 ;
  assign n15450 = n15447 | n15449 ;
  assign n15451 = n15329 & n15450 ;
  assign n15452 = n15329 & ~n15451 ;
  assign n15487 = n15212 | n15218 ;
  assign n15488 = ( n15214 & n15218 ) | ( n15214 & n15487 ) | ( n15218 & n15487 ) ;
  assign n15489 = ( n15215 & n15217 ) | ( n15215 & n15488 ) | ( n15217 & n15488 ) ;
  assign n15465 = n14880 | n15250 ;
  assign n15466 = ( n15250 & n15251 ) | ( n15250 & n15465 ) | ( n15251 & n15465 ) ;
  assign n15453 = x38 & x43 ;
  assign n15454 = x39 & x42 ;
  assign n15455 = n15453 | n15454 ;
  assign n15456 = n5392 & n5407 ;
  assign n15457 = x27 & x54 ;
  assign n15458 = ~n15456 & n15457 ;
  assign n15459 = n15455 | n15456 ;
  assign n15460 = ( n15456 & n15458 ) | ( n15456 & n15459 ) | ( n15458 & n15459 ) ;
  assign n15461 = n15455 & ~n15460 ;
  assign n15462 = ~n15455 & n15457 ;
  assign n15463 = ( n15457 & ~n15458 ) | ( n15457 & n15462 ) | ( ~n15458 & n15462 ) ;
  assign n15464 = n15461 | n15463 ;
  assign n15467 = n15464 & n15466 ;
  assign n15468 = n15466 & ~n15467 ;
  assign n15470 = n15002 | n15230 ;
  assign n15471 = ( n15230 & n15231 ) | ( n15230 & n15470 ) | ( n15231 & n15470 ) ;
  assign n15469 = n15464 & ~n15466 ;
  assign n15472 = n15469 & n15471 ;
  assign n15473 = ( n15468 & n15471 ) | ( n15468 & n15472 ) | ( n15471 & n15472 ) ;
  assign n15474 = n15469 | n15471 ;
  assign n15475 = n15468 | n15474 ;
  assign n15476 = ~n15473 & n15475 ;
  assign n15477 = n15238 | n15243 ;
  assign n15478 = n15254 | n15259 ;
  assign n15479 = ( n15259 & n15260 ) | ( n15259 & n15478 ) | ( n15260 & n15478 ) ;
  assign n15480 = n15477 & n15479 ;
  assign n15481 = n15477 & ~n15480 ;
  assign n15482 = n15479 & ~n15480 ;
  assign n15483 = n15481 | n15482 ;
  assign n15484 = n15476 & n15483 ;
  assign n15485 = n15476 | n15483 ;
  assign n15486 = ~n15484 & n15485 ;
  assign n15490 = n15486 & n15489 ;
  assign n15491 = n15489 & ~n15490 ;
  assign n15492 = n15190 | n15200 ;
  assign n15493 = ~n15183 & n15185 ;
  assign n15494 = ( n15183 & n15184 ) | ( n15183 & n15493 ) | ( n15184 & n15493 ) ;
  assign n15495 = n15153 | n15494 ;
  assign n15496 = n15153 & n15494 ;
  assign n15497 = n15495 & ~n15496 ;
  assign n15498 = n15131 | n15134 ;
  assign n15499 = n15497 | n15498 ;
  assign n15500 = n15497 & n15498 ;
  assign n15501 = n15499 & ~n15500 ;
  assign n15502 = n15189 | n15199 ;
  assign n15503 = n15501 & n15502 ;
  assign n15504 = n15189 & n15501 ;
  assign n15505 = ( n15492 & n15503 ) | ( n15492 & n15504 ) | ( n15503 & n15504 ) ;
  assign n15506 = n15501 | n15502 ;
  assign n15507 = n15189 | n15501 ;
  assign n15508 = ( n15492 & n15506 ) | ( n15492 & n15507 ) | ( n15506 & n15507 ) ;
  assign n15509 = ~n15505 & n15508 ;
  assign n15510 = n15169 & n15191 ;
  assign n15511 = ( n15168 & n15191 ) | ( n15168 & n15510 ) | ( n15191 & n15510 ) ;
  assign n15512 = ( n15173 & n15196 ) | ( n15173 & n15511 ) | ( n15196 & n15511 ) ;
  assign n15513 = ( ~n15173 & n15191 ) | ( ~n15173 & n15196 ) | ( n15191 & n15196 ) ;
  assign n15514 = n15173 | n15513 ;
  assign n15515 = ~n15512 & n15514 ;
  assign n15516 = n2546 & n10866 ;
  assign n15517 = n2965 & n7112 ;
  assign n15518 = n15516 | n15517 ;
  assign n15519 = n4062 & n6834 ;
  assign n15520 = x51 & n15519 ;
  assign n15521 = ( x51 & ~n15518 ) | ( x51 & n15520 ) | ( ~n15518 & n15520 ) ;
  assign n15522 = x30 & n15521 ;
  assign n15523 = n15518 | n15519 ;
  assign n15524 = x31 & x50 ;
  assign n15525 = x32 & x49 ;
  assign n15526 = ( ~n15519 & n15524 ) | ( ~n15519 & n15525 ) | ( n15524 & n15525 ) ;
  assign n15527 = n15524 & n15525 ;
  assign n15528 = ( ~n15518 & n15526 ) | ( ~n15518 & n15527 ) | ( n15526 & n15527 ) ;
  assign n15529 = ~n15523 & n15528 ;
  assign n15530 = n15522 | n15529 ;
  assign n15531 = n15515 & ~n15530 ;
  assign n15532 = n15515 | n15530 ;
  assign n15533 = ( ~n15515 & n15531 ) | ( ~n15515 & n15532 ) | ( n15531 & n15532 ) ;
  assign n15534 = n15509 & ~n15533 ;
  assign n15535 = ~n15509 & n15533 ;
  assign n15536 = n15534 | n15535 ;
  assign n15537 = n15119 & n15130 ;
  assign n15538 = n15119 & ~n15537 ;
  assign n15539 = ~n15119 & n15130 ;
  assign n15540 = n15163 & n15539 ;
  assign n15541 = ( n15163 & n15538 ) | ( n15163 & n15540 ) | ( n15538 & n15540 ) ;
  assign n15542 = n15208 | n15541 ;
  assign n15543 = n15536 | n15542 ;
  assign n15544 = n15536 & n15542 ;
  assign n15545 = n15543 & ~n15544 ;
  assign n15546 = n15111 | n15126 ;
  assign n15547 = n15111 & n15126 ;
  assign n15548 = n15546 & ~n15547 ;
  assign n15549 = n15096 | n15548 ;
  assign n15550 = n15096 & n15548 ;
  assign n15551 = n15549 & ~n15550 ;
  assign n15552 = n15116 | n15130 ;
  assign n15553 = n15143 | n15160 ;
  assign n15554 = ( n15143 & n15145 ) | ( n15143 & n15553 ) | ( n15145 & n15553 ) ;
  assign n15555 = n15552 & n15554 ;
  assign n15556 = n15116 & n15554 ;
  assign n15557 = ( n15119 & n15555 ) | ( n15119 & n15556 ) | ( n15555 & n15556 ) ;
  assign n15558 = n15552 | n15554 ;
  assign n15559 = n15116 | n15554 ;
  assign n15560 = ( n15119 & n15558 ) | ( n15119 & n15559 ) | ( n15558 & n15559 ) ;
  assign n15561 = ~n15557 & n15560 ;
  assign n15562 = n15551 & n15561 ;
  assign n15563 = n15551 | n15561 ;
  assign n15564 = ~n15562 & n15563 ;
  assign n15565 = n15545 & n15564 ;
  assign n15566 = n15545 | n15564 ;
  assign n15567 = ~n15565 & n15566 ;
  assign n15568 = n15490 | n15567 ;
  assign n15569 = n15486 & ~n15567 ;
  assign n15570 = ( n15491 & ~n15568 ) | ( n15491 & n15569 ) | ( ~n15568 & n15569 ) ;
  assign n15571 = n15490 & n15567 ;
  assign n15572 = ~n15486 & n15567 ;
  assign n15573 = ( ~n15491 & n15571 ) | ( ~n15491 & n15572 ) | ( n15571 & n15572 ) ;
  assign n15574 = n15570 | n15573 ;
  assign n15575 = ~n15329 & n15450 ;
  assign n15576 = n15574 & n15575 ;
  assign n15577 = ( n15452 & n15574 ) | ( n15452 & n15576 ) | ( n15574 & n15576 ) ;
  assign n15578 = n15574 | n15575 ;
  assign n15579 = n15452 | n15578 ;
  assign n15580 = ~n15577 & n15579 ;
  assign n15581 = n15225 | n15295 ;
  assign n15582 = ( n15225 & n15226 ) | ( n15225 & n15581 ) | ( n15226 & n15581 ) ;
  assign n15583 = ( n15328 & n15580 ) | ( n15328 & ~n15582 ) | ( n15580 & ~n15582 ) ;
  assign n15584 = ( ~n15580 & n15582 ) | ( ~n15580 & n15583 ) | ( n15582 & n15583 ) ;
  assign n15585 = ( ~n15328 & n15583 ) | ( ~n15328 & n15584 ) | ( n15583 & n15584 ) ;
  assign n15586 = n15580 & n15582 ;
  assign n15587 = n15580 | n15582 ;
  assign n15588 = n15586 | n15587 ;
  assign n15589 = ( n15327 & n15586 ) | ( n15327 & n15588 ) | ( n15586 & n15588 ) ;
  assign n15590 = ( n15322 & n15586 ) | ( n15322 & n15588 ) | ( n15586 & n15588 ) ;
  assign n15591 = ( n15321 & n15586 ) | ( n15321 & n15588 ) | ( n15586 & n15588 ) ;
  assign n15592 = ( n14840 & n15590 ) | ( n14840 & n15591 ) | ( n15590 & n15591 ) ;
  assign n15593 = ( n14575 & n15589 ) | ( n14575 & n15592 ) | ( n15589 & n15592 ) ;
  assign n15594 = ( n14571 & n15589 ) | ( n14571 & n15592 ) | ( n15589 & n15592 ) ;
  assign n15595 = ( n13196 & n15593 ) | ( n13196 & n15594 ) | ( n15593 & n15594 ) ;
  assign n15596 = n15451 | n15577 ;
  assign n15597 = ( n15486 & ~n15490 ) | ( n15486 & n15491 ) | ( ~n15490 & n15491 ) ;
  assign n15598 = ( n15490 & n15568 ) | ( n15490 & n15597 ) | ( n15568 & n15597 ) ;
  assign n15599 = x31 & x51 ;
  assign n15600 = x21 & x61 ;
  assign n15601 = n15599 & n15600 ;
  assign n15602 = x51 & x62 ;
  assign n15603 = n6587 & n15602 ;
  assign n15604 = n1434 & n10684 ;
  assign n15605 = n15603 | n15604 ;
  assign n15606 = x62 & n15601 ;
  assign n15607 = ( x62 & ~n15605 ) | ( x62 & n15606 ) | ( ~n15605 & n15606 ) ;
  assign n15608 = x20 & n15607 ;
  assign n15609 = ( n15599 & n15600 ) | ( n15599 & ~n15605 ) | ( n15600 & ~n15605 ) ;
  assign n15610 = ( ~n15601 & n15608 ) | ( ~n15601 & n15609 ) | ( n15608 & n15609 ) ;
  assign n15611 = n4318 & n6345 ;
  assign n15612 = n3321 & n6834 ;
  assign n15613 = n15611 | n15612 ;
  assign n15614 = n4530 & n6759 ;
  assign n15615 = x50 & n15614 ;
  assign n15616 = ( x50 & ~n15613 ) | ( x50 & n15615 ) | ( ~n15613 & n15615 ) ;
  assign n15617 = x32 & n15616 ;
  assign n15618 = n15613 | n15614 ;
  assign n15619 = x33 & x49 ;
  assign n15620 = x34 & x48 ;
  assign n15621 = ( ~n15614 & n15619 ) | ( ~n15614 & n15620 ) | ( n15619 & n15620 ) ;
  assign n15622 = n15619 & n15620 ;
  assign n15623 = ( ~n15613 & n15621 ) | ( ~n15613 & n15622 ) | ( n15621 & n15622 ) ;
  assign n15624 = ~n15618 & n15623 ;
  assign n15625 = n15617 | n15624 ;
  assign n15626 = n15610 & n15625 ;
  assign n15627 = n15610 & ~n15626 ;
  assign n15628 = n15625 & ~n15626 ;
  assign n15629 = n15627 | n15628 ;
  assign n15630 = n2148 & n10975 ;
  assign n15631 = n1932 & n10370 ;
  assign n15632 = n15630 | n15631 ;
  assign n15633 = n1686 & n9831 ;
  assign n15634 = x60 & n15633 ;
  assign n15635 = ( x60 & ~n15632 ) | ( x60 & n15634 ) | ( ~n15632 & n15634 ) ;
  assign n15636 = x22 & n15635 ;
  assign n15637 = n15632 | n15633 ;
  assign n15638 = x23 & x59 ;
  assign n15639 = ( n12431 & ~n15633 ) | ( n12431 & n15638 ) | ( ~n15633 & n15638 ) ;
  assign n15640 = n12431 & n15638 ;
  assign n15641 = ( ~n15632 & n15639 ) | ( ~n15632 & n15640 ) | ( n15639 & n15640 ) ;
  assign n15642 = ~n15637 & n15641 ;
  assign n15643 = n15636 | n15642 ;
  assign n15644 = ~n15629 & n15643 ;
  assign n15645 = n15629 & ~n15643 ;
  assign n15646 = n15644 | n15645 ;
  assign n15647 = n15467 | n15473 ;
  assign n15648 = n15646 | n15647 ;
  assign n15649 = n15646 & n15647 ;
  assign n15650 = n15648 & ~n15649 ;
  assign n15651 = x29 & x53 ;
  assign n15652 = x30 & x52 ;
  assign n15653 = n15651 | n15652 ;
  assign n15654 = n2709 & n8161 ;
  assign n15655 = n6973 & ~n15654 ;
  assign n15656 = n15653 | n15654 ;
  assign n15657 = ( n15654 & n15655 ) | ( n15654 & n15656 ) | ( n15655 & n15656 ) ;
  assign n15658 = n15653 & ~n15657 ;
  assign n15659 = n6973 & ~n15653 ;
  assign n15660 = ( n6973 & ~n15655 ) | ( n6973 & n15659 ) | ( ~n15655 & n15659 ) ;
  assign n15661 = n15658 | n15660 ;
  assign n15662 = x38 & x44 ;
  assign n15663 = x39 & x43 ;
  assign n15664 = n15662 | n15663 ;
  assign n15665 = n5392 & n5658 ;
  assign n15666 = n15664 | n15665 ;
  assign n15667 = x26 & x56 ;
  assign n15668 = ( ~n15665 & n15666 ) | ( ~n15665 & n15667 ) | ( n15666 & n15667 ) ;
  assign n15669 = ( n15665 & n15666 ) | ( n15665 & ~n15667 ) | ( n15666 & ~n15667 ) ;
  assign n15670 = ( ~n15666 & n15668 ) | ( ~n15666 & n15669 ) | ( n15668 & n15669 ) ;
  assign n15671 = n15661 & n15670 ;
  assign n15672 = n15661 & ~n15671 ;
  assign n15673 = x37 & x47 ;
  assign n15674 = n6308 & n15673 ;
  assign n15675 = n4078 & n6147 ;
  assign n15676 = n15674 | n15675 ;
  assign n15677 = n3770 & n5975 ;
  assign n15678 = x47 & n15677 ;
  assign n15679 = ( x47 & ~n15676 ) | ( x47 & n15678 ) | ( ~n15676 & n15678 ) ;
  assign n15680 = x35 & n15679 ;
  assign n15681 = n15676 | n15677 ;
  assign n15682 = ( n6638 & n6961 ) | ( n6638 & ~n15677 ) | ( n6961 & ~n15677 ) ;
  assign n15683 = n6638 & n6961 ;
  assign n15684 = ( ~n15676 & n15682 ) | ( ~n15676 & n15683 ) | ( n15682 & n15683 ) ;
  assign n15685 = ~n15681 & n15684 ;
  assign n15686 = n15680 | n15685 ;
  assign n15687 = ~n15661 & n15670 ;
  assign n15688 = n15686 & ~n15687 ;
  assign n15689 = ~n15672 & n15688 ;
  assign n15690 = ~n15686 & n15687 ;
  assign n15691 = ( n15672 & ~n15686 ) | ( n15672 & n15690 ) | ( ~n15686 & n15690 ) ;
  assign n15692 = n15689 | n15691 ;
  assign n15693 = n15650 | n15692 ;
  assign n15694 = n15650 & n15692 ;
  assign n15695 = n15693 & ~n15694 ;
  assign n15696 = n15476 | n15480 ;
  assign n15697 = n15695 & ~n15696 ;
  assign n15698 = ~n15480 & n15695 ;
  assign n15699 = ( ~n15483 & n15697 ) | ( ~n15483 & n15698 ) | ( n15697 & n15698 ) ;
  assign n15700 = ~n15695 & n15696 ;
  assign n15701 = n15480 & ~n15695 ;
  assign n15702 = ( n15483 & n15700 ) | ( n15483 & n15701 ) | ( n15700 & n15701 ) ;
  assign n15703 = n15699 | n15702 ;
  assign n15704 = ( n15536 & n15542 ) | ( n15536 & n15564 ) | ( n15542 & n15564 ) ;
  assign n15705 = n15703 & n15704 ;
  assign n15706 = n15703 | n15704 ;
  assign n15707 = ~n15705 & n15706 ;
  assign n15708 = n15568 & n15707 ;
  assign n15709 = n15490 & n15707 ;
  assign n15710 = ( n15597 & n15708 ) | ( n15597 & n15709 ) | ( n15708 & n15709 ) ;
  assign n15711 = n15598 & ~n15710 ;
  assign n15712 = n15366 | n15523 ;
  assign n15713 = n15366 & n15523 ;
  assign n15714 = n15712 & ~n15713 ;
  assign n15715 = n15422 | n15714 ;
  assign n15716 = n15422 & n15714 ;
  assign n15717 = n15715 & ~n15716 ;
  assign n15718 = n15344 | n15389 ;
  assign n15719 = n15344 & n15389 ;
  assign n15720 = n15718 & ~n15719 ;
  assign n15721 = n15405 | n15720 ;
  assign n15722 = n15405 & n15720 ;
  assign n15723 = n15721 & ~n15722 ;
  assign n15724 = n15412 | n15723 ;
  assign n15725 = n15432 | n15724 ;
  assign n15726 = n15412 & n15723 ;
  assign n15727 = ( n15432 & n15723 ) | ( n15432 & n15726 ) | ( n15723 & n15726 ) ;
  assign n15728 = n15725 & ~n15727 ;
  assign n15729 = n15717 & n15728 ;
  assign n15730 = n15717 | n15728 ;
  assign n15731 = ~n15729 & n15730 ;
  assign n15732 = n15380 | n15435 ;
  assign n15733 = ( n15380 & n15381 ) | ( n15380 & n15732 ) | ( n15381 & n15732 ) ;
  assign n15734 = n15731 | n15733 ;
  assign n15735 = n15731 & n15733 ;
  assign n15736 = n15734 & ~n15735 ;
  assign n15737 = n15512 | n15530 ;
  assign n15738 = ( n15512 & n15515 ) | ( n15512 & n15737 ) | ( n15515 & n15737 ) ;
  assign n15739 = n15358 & n15738 ;
  assign n15740 = ( n15373 & n15738 ) | ( n15373 & n15739 ) | ( n15738 & n15739 ) ;
  assign n15741 = n15358 | n15738 ;
  assign n15742 = n15373 | n15741 ;
  assign n15743 = ~n15740 & n15742 ;
  assign n15744 = x41 & x62 ;
  assign n15745 = x19 & n15744 ;
  assign n15746 = n5813 & ~n15745 ;
  assign n15747 = n13913 & n15745 ;
  assign n15748 = ( n13913 & n15746 ) | ( n13913 & n15747 ) | ( n15746 & n15747 ) ;
  assign n15749 = n13913 | n15745 ;
  assign n15750 = n15746 | n15749 ;
  assign n15751 = ~n15748 & n15750 ;
  assign n15752 = n15460 | n15751 ;
  assign n15753 = n15460 & n15751 ;
  assign n15754 = n15752 & ~n15753 ;
  assign n15755 = n15743 & n15754 ;
  assign n15756 = n15743 | n15754 ;
  assign n15757 = ~n15755 & n15756 ;
  assign n15758 = n15736 & n15757 ;
  assign n15759 = n15736 | n15757 ;
  assign n15760 = ~n15758 & n15759 ;
  assign n15775 = n15496 | n15498 ;
  assign n15776 = ( n15496 & n15497 ) | ( n15496 & n15775 ) | ( n15497 & n15775 ) ;
  assign n15761 = n2372 & n8357 ;
  assign n15762 = x25 & x57 ;
  assign n15763 = n7719 & n15762 ;
  assign n15764 = n15761 | n15763 ;
  assign n15765 = n2724 & n12860 ;
  assign n15766 = n7719 & n15765 ;
  assign n15767 = ( n7719 & ~n15764 ) | ( n7719 & n15766 ) | ( ~n15764 & n15766 ) ;
  assign n15768 = n15764 | n15765 ;
  assign n15769 = x27 & x55 ;
  assign n15770 = ( n15762 & ~n15765 ) | ( n15762 & n15769 ) | ( ~n15765 & n15769 ) ;
  assign n15771 = n15762 & n15769 ;
  assign n15772 = ( ~n15764 & n15770 ) | ( ~n15764 & n15771 ) | ( n15770 & n15771 ) ;
  assign n15773 = ~n15768 & n15772 ;
  assign n15774 = n15767 | n15773 ;
  assign n15777 = n15774 & n15776 ;
  assign n15778 = n15776 & ~n15777 ;
  assign n15780 = n15096 | n15547 ;
  assign n15781 = ( n15547 & n15548 ) | ( n15547 & n15780 ) | ( n15548 & n15780 ) ;
  assign n15779 = n15774 & ~n15776 ;
  assign n15782 = n15779 & n15781 ;
  assign n15783 = ( n15778 & n15781 ) | ( n15778 & n15782 ) | ( n15781 & n15782 ) ;
  assign n15784 = n15779 | n15781 ;
  assign n15785 = n15778 | n15784 ;
  assign n15786 = ~n15783 & n15785 ;
  assign n15787 = n15505 | n15533 ;
  assign n15788 = ( n15505 & n15509 ) | ( n15505 & n15787 ) | ( n15509 & n15787 ) ;
  assign n15789 = n15551 | n15557 ;
  assign n15790 = ( n15557 & n15561 ) | ( n15557 & n15789 ) | ( n15561 & n15789 ) ;
  assign n15791 = n15788 & n15790 ;
  assign n15792 = n15788 & ~n15791 ;
  assign n15793 = n15790 & ~n15791 ;
  assign n15794 = n15792 | n15793 ;
  assign n15795 = n15786 & n15794 ;
  assign n15796 = n15786 | n15794 ;
  assign n15797 = ~n15795 & n15796 ;
  assign n15798 = n15330 | n15440 ;
  assign n15799 = ( n15440 & n15446 ) | ( n15440 & n15798 ) | ( n15446 & n15798 ) ;
  assign n15800 = ( n15760 & ~n15797 ) | ( n15760 & n15799 ) | ( ~n15797 & n15799 ) ;
  assign n15801 = ( n15797 & ~n15799 ) | ( n15797 & n15800 ) | ( ~n15799 & n15800 ) ;
  assign n15802 = ( ~n15760 & n15800 ) | ( ~n15760 & n15801 ) | ( n15800 & n15801 ) ;
  assign n15803 = ~n15568 & n15707 ;
  assign n15804 = ~n15490 & n15707 ;
  assign n15805 = ( ~n15597 & n15803 ) | ( ~n15597 & n15804 ) | ( n15803 & n15804 ) ;
  assign n15806 = n15802 & n15805 ;
  assign n15807 = ( n15711 & n15802 ) | ( n15711 & n15806 ) | ( n15802 & n15806 ) ;
  assign n15808 = n15802 | n15805 ;
  assign n15809 = n15711 | n15808 ;
  assign n15810 = ~n15807 & n15809 ;
  assign n15811 = ( n15595 & n15596 ) | ( n15595 & ~n15810 ) | ( n15596 & ~n15810 ) ;
  assign n15812 = ( ~n15596 & n15810 ) | ( ~n15596 & n15811 ) | ( n15810 & n15811 ) ;
  assign n15813 = ( ~n15595 & n15811 ) | ( ~n15595 & n15812 ) | ( n15811 & n15812 ) ;
  assign n15814 = n15596 & n15810 ;
  assign n15815 = n15596 | n15810 ;
  assign n15816 = n15814 | n15815 ;
  assign n15817 = ( n15595 & n15814 ) | ( n15595 & n15816 ) | ( n15814 & n15816 ) ;
  assign n15818 = n15710 | n15807 ;
  assign n15819 = n15777 | n15783 ;
  assign n15820 = x39 & x44 ;
  assign n15821 = x40 & x43 ;
  assign n15822 = n15820 | n15821 ;
  assign n15823 = n4555 & n5658 ;
  assign n15824 = x29 & x54 ;
  assign n15825 = ~n15823 & n15824 ;
  assign n15826 = n15822 | n15823 ;
  assign n15827 = ( n15823 & n15825 ) | ( n15823 & n15826 ) | ( n15825 & n15826 ) ;
  assign n15828 = n15822 & ~n15827 ;
  assign n15829 = ( ~n15822 & n15823 ) | ( ~n15822 & n15824 ) | ( n15823 & n15824 ) ;
  assign n15830 = n15824 & n15829 ;
  assign n15831 = n15828 | n15830 ;
  assign n15832 = x42 & x62 ;
  assign n15833 = x21 & n15832 ;
  assign n15834 = n5710 & n15833 ;
  assign n15835 = n5710 & ~n15833 ;
  assign n15836 = n15833 | n15835 ;
  assign n15837 = x21 & x62 ;
  assign n15838 = ( x42 & ~n15833 ) | ( x42 & n15837 ) | ( ~n15833 & n15837 ) ;
  assign n15839 = x42 & n15837 ;
  assign n15840 = ( ~n15835 & n15838 ) | ( ~n15835 & n15839 ) | ( n15838 & n15839 ) ;
  assign n15841 = ~n15836 & n15840 ;
  assign n15842 = n15834 | n15841 ;
  assign n15843 = n15831 & n15842 ;
  assign n15844 = n15831 & ~n15843 ;
  assign n15845 = n3129 & n6345 ;
  assign n15846 = n4530 & n6834 ;
  assign n15847 = n15845 | n15846 ;
  assign n15848 = n3483 & n6759 ;
  assign n15849 = x50 & n15848 ;
  assign n15850 = ( x50 & ~n15847 ) | ( x50 & n15849 ) | ( ~n15847 & n15849 ) ;
  assign n15851 = x33 & n15850 ;
  assign n15852 = n15847 | n15848 ;
  assign n15853 = x34 & x49 ;
  assign n15854 = x35 & x48 ;
  assign n15855 = ( ~n15848 & n15853 ) | ( ~n15848 & n15854 ) | ( n15853 & n15854 ) ;
  assign n15856 = n15853 & n15854 ;
  assign n15857 = ( ~n15847 & n15855 ) | ( ~n15847 & n15856 ) | ( n15855 & n15856 ) ;
  assign n15858 = ~n15852 & n15857 ;
  assign n15859 = n15851 | n15858 ;
  assign n15860 = ~n15831 & n15842 ;
  assign n15861 = n15859 & n15860 ;
  assign n15862 = ( n15844 & n15859 ) | ( n15844 & n15861 ) | ( n15859 & n15861 ) ;
  assign n15863 = n15859 | n15860 ;
  assign n15864 = n15844 | n15863 ;
  assign n15865 = ~n15862 & n15864 ;
  assign n15866 = n15819 | n15865 ;
  assign n15867 = n15819 & n15865 ;
  assign n15868 = n15866 & ~n15867 ;
  assign n15869 = n2511 & n9272 ;
  assign n15870 = x32 & x58 ;
  assign n15871 = n14196 & n15870 ;
  assign n15872 = n15869 | n15871 ;
  assign n15873 = x51 & x57 ;
  assign n15874 = n3422 & n15873 ;
  assign n15875 = x58 & n15874 ;
  assign n15876 = ( x58 & ~n15872 ) | ( x58 & n15875 ) | ( ~n15872 & n15875 ) ;
  assign n15877 = x25 & n15876 ;
  assign n15878 = n15872 | n15874 ;
  assign n15879 = x26 & x57 ;
  assign n15880 = x32 & x51 ;
  assign n15881 = ( ~n15874 & n15879 ) | ( ~n15874 & n15880 ) | ( n15879 & n15880 ) ;
  assign n15882 = n15879 & n15880 ;
  assign n15883 = ( ~n15872 & n15881 ) | ( ~n15872 & n15882 ) | ( n15881 & n15882 ) ;
  assign n15884 = ~n15878 & n15883 ;
  assign n15885 = n15877 | n15884 ;
  assign n15886 = n3731 & n5610 ;
  assign n15887 = n3770 & n6147 ;
  assign n15888 = n15886 | n15887 ;
  assign n15889 = n4857 & n5975 ;
  assign n15890 = x47 & n15889 ;
  assign n15891 = ( x47 & ~n15888 ) | ( x47 & n15890 ) | ( ~n15888 & n15890 ) ;
  assign n15892 = x36 & n15891 ;
  assign n15893 = n15888 | n15889 ;
  assign n15894 = x37 & x46 ;
  assign n15895 = x38 & x45 ;
  assign n15896 = ( ~n15889 & n15894 ) | ( ~n15889 & n15895 ) | ( n15894 & n15895 ) ;
  assign n15897 = n15894 & n15895 ;
  assign n15898 = ( ~n15888 & n15896 ) | ( ~n15888 & n15897 ) | ( n15896 & n15897 ) ;
  assign n15899 = ~n15893 & n15898 ;
  assign n15900 = n15892 | n15899 ;
  assign n15901 = n15885 & n15900 ;
  assign n15902 = n15885 & ~n15901 ;
  assign n15903 = n15900 & ~n15901 ;
  assign n15904 = n15902 | n15903 ;
  assign n15905 = x20 & x63 ;
  assign n15906 = x22 & x61 ;
  assign n15907 = n15905 | n15906 ;
  assign n15908 = n1710 & n10856 ;
  assign n15909 = n14997 & ~n15908 ;
  assign n15910 = n15907 | n15908 ;
  assign n15911 = ( n15908 & n15909 ) | ( n15908 & n15910 ) | ( n15909 & n15910 ) ;
  assign n15912 = n15907 & ~n15911 ;
  assign n15913 = n14997 & ~n15907 ;
  assign n15914 = ( n14997 & ~n15909 ) | ( n14997 & n15913 ) | ( ~n15909 & n15913 ) ;
  assign n15915 = n15912 | n15914 ;
  assign n15916 = ~n15904 & n15915 ;
  assign n15917 = n15904 & ~n15915 ;
  assign n15918 = n15916 | n15917 ;
  assign n15919 = n15868 | n15918 ;
  assign n15920 = n15868 & n15918 ;
  assign n15921 = n15919 & ~n15920 ;
  assign n15922 = n15786 | n15791 ;
  assign n15923 = ( n15791 & n15794 ) | ( n15791 & n15922 ) | ( n15794 & n15922 ) ;
  assign n15924 = n15921 & n15923 ;
  assign n15925 = n15921 | n15923 ;
  assign n15926 = ~n15924 & n15925 ;
  assign n15927 = ( n15731 & n15733 ) | ( n15731 & n15757 ) | ( n15733 & n15757 ) ;
  assign n15928 = n15926 | n15927 ;
  assign n15929 = n15926 & n15927 ;
  assign n15930 = n15928 & ~n15929 ;
  assign n15931 = n15797 & n15799 ;
  assign n15932 = n15799 & ~n15931 ;
  assign n15933 = n15760 & n15797 ;
  assign n15934 = ~n15799 & n15933 ;
  assign n15935 = ( n15760 & n15932 ) | ( n15760 & n15934 ) | ( n15932 & n15934 ) ;
  assign n15936 = n15930 & n15931 ;
  assign n15937 = ( n15930 & n15935 ) | ( n15930 & n15936 ) | ( n15935 & n15936 ) ;
  assign n15938 = n15930 | n15931 ;
  assign n15939 = n15935 | n15938 ;
  assign n15940 = ~n15937 & n15939 ;
  assign n15941 = n15422 | n15713 ;
  assign n15942 = ( n15713 & n15714 ) | ( n15713 & n15941 ) | ( n15714 & n15941 ) ;
  assign n15943 = n15405 | n15719 ;
  assign n15944 = ( n15719 & n15720 ) | ( n15719 & n15943 ) | ( n15720 & n15943 ) ;
  assign n15945 = n15942 | n15944 ;
  assign n15946 = n15942 & n15944 ;
  assign n15947 = n15945 & ~n15946 ;
  assign n15948 = n15626 | n15643 ;
  assign n15949 = ( n15626 & n15629 ) | ( n15626 & n15948 ) | ( n15629 & n15948 ) ;
  assign n15950 = n15947 | n15949 ;
  assign n15951 = n15947 & n15949 ;
  assign n15952 = n15950 & ~n15951 ;
  assign n15978 = n15460 | n15748 ;
  assign n15979 = ( n15748 & n15751 ) | ( n15748 & n15978 ) | ( n15751 & n15978 ) ;
  assign n15953 = n1686 & n10370 ;
  assign n15954 = x24 & x59 ;
  assign n15955 = x23 & x60 ;
  assign n15956 = n15954 | n15955 ;
  assign n15957 = ~n15953 & n15956 ;
  assign n15958 = n15657 & n15957 ;
  assign n15959 = n15657 & ~n15958 ;
  assign n15960 = ~n15657 & n15957 ;
  assign n15961 = n15959 | n15960 ;
  assign n15962 = n2965 & n8161 ;
  assign n15963 = x31 & x55 ;
  assign n15964 = n15121 & n15963 ;
  assign n15965 = n15962 | n15964 ;
  assign n15966 = n3280 & n8360 ;
  assign n15967 = x52 & n15966 ;
  assign n15968 = ( x52 & ~n15965 ) | ( x52 & n15967 ) | ( ~n15965 & n15967 ) ;
  assign n15969 = x31 & n15968 ;
  assign n15970 = n15965 | n15966 ;
  assign n15971 = x28 & x55 ;
  assign n15972 = x30 & x53 ;
  assign n15973 = ( ~n15966 & n15971 ) | ( ~n15966 & n15972 ) | ( n15971 & n15972 ) ;
  assign n15974 = n15971 & n15972 ;
  assign n15975 = ( ~n15965 & n15973 ) | ( ~n15965 & n15974 ) | ( n15973 & n15974 ) ;
  assign n15976 = ~n15970 & n15975 ;
  assign n15977 = n15969 | n15976 ;
  assign n15980 = ( n15961 & ~n15977 ) | ( n15961 & n15979 ) | ( ~n15977 & n15979 ) ;
  assign n15981 = ( ~n15961 & n15977 ) | ( ~n15961 & n15980 ) | ( n15977 & n15980 ) ;
  assign n15982 = ( ~n15979 & n15980 ) | ( ~n15979 & n15981 ) | ( n15980 & n15981 ) ;
  assign n15983 = n15740 | n15754 ;
  assign n15984 = ( n15740 & n15743 ) | ( n15740 & n15983 ) | ( n15743 & n15983 ) ;
  assign n15985 = n15982 & n15984 ;
  assign n15986 = n15982 | n15984 ;
  assign n15987 = ~n15985 & n15986 ;
  assign n15988 = n15952 & n15987 ;
  assign n15989 = n15952 | n15987 ;
  assign n15990 = ~n15988 & n15989 ;
  assign n15991 = n15695 & n15990 ;
  assign n15992 = ( n15480 & n15483 ) | ( n15480 & n15696 ) | ( n15483 & n15696 ) ;
  assign n15993 = n15991 & n15992 ;
  assign n15994 = ( n15705 & n15990 ) | ( n15705 & n15993 ) | ( n15990 & n15993 ) ;
  assign n15995 = n15695 & n15696 ;
  assign n15996 = n15480 & n15695 ;
  assign n15997 = ( n15483 & n15995 ) | ( n15483 & n15996 ) | ( n15995 & n15996 ) ;
  assign n15998 = n15990 | n15997 ;
  assign n15999 = n15705 | n15998 ;
  assign n16000 = ~n15994 & n15999 ;
  assign n16001 = ~n15665 & n15667 ;
  assign n16002 = ( n15665 & n15666 ) | ( n15665 & n16001 ) | ( n15666 & n16001 ) ;
  assign n16003 = n15637 | n15681 ;
  assign n16004 = n15637 & n15681 ;
  assign n16005 = n16003 & ~n16004 ;
  assign n16006 = n16002 | n16005 ;
  assign n16007 = n16002 & n16005 ;
  assign n16008 = n16006 & ~n16007 ;
  assign n16009 = n15672 | n15687 ;
  assign n16010 = n15601 | n15605 ;
  assign n16011 = n15618 | n16010 ;
  assign n16012 = n15618 & n16010 ;
  assign n16013 = n16011 & ~n16012 ;
  assign n16014 = n15768 | n16013 ;
  assign n16015 = n15768 & n16013 ;
  assign n16016 = n16014 & ~n16015 ;
  assign n16017 = n15671 | n15686 ;
  assign n16018 = n16016 & n16017 ;
  assign n16019 = n15671 & n16016 ;
  assign n16020 = ( n16009 & n16018 ) | ( n16009 & n16019 ) | ( n16018 & n16019 ) ;
  assign n16021 = n16016 | n16017 ;
  assign n16022 = n15671 | n16016 ;
  assign n16023 = ( n16009 & n16021 ) | ( n16009 & n16022 ) | ( n16021 & n16022 ) ;
  assign n16024 = ~n16020 & n16023 ;
  assign n16025 = n16008 & n16024 ;
  assign n16026 = n16008 | n16024 ;
  assign n16027 = ~n16025 & n16026 ;
  assign n16028 = n15649 | n15692 ;
  assign n16029 = ( n15649 & n15650 ) | ( n15649 & n16028 ) | ( n15650 & n16028 ) ;
  assign n16030 = n15717 | n15727 ;
  assign n16031 = ( n15727 & n15728 ) | ( n15727 & n16030 ) | ( n15728 & n16030 ) ;
  assign n16032 = ( n16027 & n16029 ) | ( n16027 & ~n16031 ) | ( n16029 & ~n16031 ) ;
  assign n16033 = ( ~n16029 & n16031 ) | ( ~n16029 & n16032 ) | ( n16031 & n16032 ) ;
  assign n16034 = ( ~n16027 & n16032 ) | ( ~n16027 & n16033 ) | ( n16032 & n16033 ) ;
  assign n16035 = n16000 & ~n16034 ;
  assign n16036 = ~n16000 & n16034 ;
  assign n16037 = n16035 | n16036 ;
  assign n16038 = ~n15940 & n16037 ;
  assign n16039 = n15940 & ~n16037 ;
  assign n16040 = n16038 | n16039 ;
  assign n16041 = ( n15817 & n15818 ) | ( n15817 & ~n16040 ) | ( n15818 & ~n16040 ) ;
  assign n16042 = ( ~n15818 & n16040 ) | ( ~n15818 & n16041 ) | ( n16040 & n16041 ) ;
  assign n16043 = ( ~n15817 & n16041 ) | ( ~n15817 & n16042 ) | ( n16041 & n16042 ) ;
  assign n16044 = n15940 & n16037 ;
  assign n16045 = n15937 | n16044 ;
  assign n16046 = n15993 | n16034 ;
  assign n16047 = n15990 | n16034 ;
  assign n16048 = ( n15705 & n16046 ) | ( n15705 & n16047 ) | ( n16046 & n16047 ) ;
  assign n16049 = ( n15994 & n16000 ) | ( n15994 & n16048 ) | ( n16000 & n16048 ) ;
  assign n16050 = n15911 & n15953 ;
  assign n16051 = ( n15911 & n15958 ) | ( n15911 & n16050 ) | ( n15958 & n16050 ) ;
  assign n16052 = n15911 | n15953 ;
  assign n16053 = n15958 | n16052 ;
  assign n16054 = ~n16051 & n16053 ;
  assign n16055 = x31 & x53 ;
  assign n16056 = x32 & x52 ;
  assign n16057 = n16055 | n16056 ;
  assign n16058 = n4062 & n8161 ;
  assign n16059 = n13839 & ~n16058 ;
  assign n16060 = n16057 | n16058 ;
  assign n16061 = ( n16058 & n16059 ) | ( n16058 & n16060 ) | ( n16059 & n16060 ) ;
  assign n16062 = n16057 & ~n16061 ;
  assign n16063 = n13839 & ~n16057 ;
  assign n16064 = ( n13839 & ~n16059 ) | ( n13839 & n16063 ) | ( ~n16059 & n16063 ) ;
  assign n16065 = n16062 | n16064 ;
  assign n16066 = ~n16054 & n16065 ;
  assign n16067 = n16054 & ~n16065 ;
  assign n16068 = n16066 | n16067 ;
  assign n16069 = n15961 & n15977 ;
  assign n16070 = n15961 & ~n16069 ;
  assign n16071 = n15977 & n15979 ;
  assign n16072 = ~n15961 & n16071 ;
  assign n16073 = n16069 | n16072 ;
  assign n16074 = n15977 | n15979 ;
  assign n16075 = ( n15961 & n15979 ) | ( n15961 & n16074 ) | ( n15979 & n16074 ) ;
  assign n16076 = ( n16070 & n16073 ) | ( n16070 & n16075 ) | ( n16073 & n16075 ) ;
  assign n16077 = n16068 | n16076 ;
  assign n16078 = n16068 & n16076 ;
  assign n16079 = n16077 & ~n16078 ;
  assign n16080 = n15946 | n15947 ;
  assign n16081 = ( n15946 & n15949 ) | ( n15946 & n16080 ) | ( n15949 & n16080 ) ;
  assign n16082 = n16079 | n16081 ;
  assign n16083 = n16079 & n16081 ;
  assign n16084 = n16082 & ~n16083 ;
  assign n16085 = n15952 | n15985 ;
  assign n16086 = ( n15985 & n15987 ) | ( n15985 & n16085 ) | ( n15987 & n16085 ) ;
  assign n16087 = n16084 | n16086 ;
  assign n16088 = n16084 & n16086 ;
  assign n16089 = n16087 & ~n16088 ;
  assign n16090 = n1337 & n10856 ;
  assign n16091 = n1585 & n10561 ;
  assign n16092 = n16090 | n16091 ;
  assign n16093 = n1932 & n10684 ;
  assign n16094 = x63 & n16093 ;
  assign n16095 = ( x63 & ~n16092 ) | ( x63 & n16094 ) | ( ~n16092 & n16094 ) ;
  assign n16096 = x21 & n16095 ;
  assign n16097 = n16092 | n16093 ;
  assign n16098 = x22 & x62 ;
  assign n16099 = x23 & x61 ;
  assign n16100 = ( ~n16093 & n16098 ) | ( ~n16093 & n16099 ) | ( n16098 & n16099 ) ;
  assign n16101 = n16098 & n16099 ;
  assign n16102 = ( ~n16092 & n16100 ) | ( ~n16092 & n16101 ) | ( n16100 & n16101 ) ;
  assign n16103 = ~n16097 & n16102 ;
  assign n16104 = n16096 | n16103 ;
  assign n16105 = x24 & x60 ;
  assign n16106 = x25 & x59 ;
  assign n16107 = n16105 | n16106 ;
  assign n16108 = n1912 & n10370 ;
  assign n16109 = x33 & x51 ;
  assign n16110 = ~n16108 & n16109 ;
  assign n16111 = n16107 | n16108 ;
  assign n16112 = ( n16108 & n16110 ) | ( n16108 & n16111 ) | ( n16110 & n16111 ) ;
  assign n16113 = n16107 & ~n16112 ;
  assign n16114 = ( ~n16107 & n16108 ) | ( ~n16107 & n16109 ) | ( n16108 & n16109 ) ;
  assign n16115 = n16109 & n16114 ;
  assign n16116 = n16113 | n16115 ;
  assign n16117 = n16104 & n16116 ;
  assign n16118 = n16104 & ~n16117 ;
  assign n16119 = n16116 & ~n16117 ;
  assign n16120 = n16118 | n16119 ;
  assign n16121 = n4914 & n6345 ;
  assign n16122 = n3483 & n6834 ;
  assign n16123 = n16121 | n16122 ;
  assign n16124 = n4078 & n6759 ;
  assign n16125 = x50 & n16124 ;
  assign n16126 = ( x50 & ~n16123 ) | ( x50 & n16125 ) | ( ~n16123 & n16125 ) ;
  assign n16127 = x34 & n16126 ;
  assign n16128 = n16123 | n16124 ;
  assign n16129 = x35 & x49 ;
  assign n16130 = x36 & x48 ;
  assign n16131 = ( ~n16124 & n16129 ) | ( ~n16124 & n16130 ) | ( n16129 & n16130 ) ;
  assign n16132 = n16129 & n16130 ;
  assign n16133 = ( ~n16123 & n16131 ) | ( ~n16123 & n16132 ) | ( n16131 & n16132 ) ;
  assign n16134 = ~n16128 & n16133 ;
  assign n16135 = n16127 | n16134 ;
  assign n16136 = ~n16120 & n16135 ;
  assign n16137 = n16120 & ~n16135 ;
  assign n16138 = n16136 | n16137 ;
  assign n16139 = x29 & x55 ;
  assign n16140 = x38 & x46 ;
  assign n16141 = n16139 & n16140 ;
  assign n16142 = n2369 & n10013 ;
  assign n16143 = x38 & x56 ;
  assign n16144 = n13606 & n16143 ;
  assign n16145 = n16142 | n16144 ;
  assign n16146 = x56 & n16141 ;
  assign n16147 = ( x56 & ~n16145 ) | ( x56 & n16146 ) | ( ~n16145 & n16146 ) ;
  assign n16148 = x28 & n16147 ;
  assign n16149 = ( n16139 & n16140 ) | ( n16139 & ~n16145 ) | ( n16140 & ~n16145 ) ;
  assign n16150 = ( ~n16141 & n16148 ) | ( ~n16141 & n16149 ) | ( n16148 & n16149 ) ;
  assign n16151 = n4350 & n5104 ;
  assign n16152 = n4555 & n6093 ;
  assign n16153 = n16151 | n16152 ;
  assign n16154 = n5658 & n5813 ;
  assign n16155 = x45 & n16154 ;
  assign n16156 = ( x45 & ~n16153 ) | ( x45 & n16155 ) | ( ~n16153 & n16155 ) ;
  assign n16157 = x39 & n16156 ;
  assign n16158 = x40 & x44 ;
  assign n16159 = n5107 | n16158 ;
  assign n16160 = ~n16154 & n16159 ;
  assign n16161 = ~n16153 & n16160 ;
  assign n16162 = n16157 | n16161 ;
  assign n16163 = n16150 & n16162 ;
  assign n16164 = n16150 & ~n16163 ;
  assign n16165 = n16162 & ~n16163 ;
  assign n16166 = n16164 | n16165 ;
  assign n16167 = x27 & x57 ;
  assign n16168 = x30 & x54 ;
  assign n16169 = n16167 | n16168 ;
  assign n16170 = x30 & x57 ;
  assign n16171 = n15457 & n16170 ;
  assign n16172 = n15673 & ~n16171 ;
  assign n16173 = n16169 | n16171 ;
  assign n16174 = ( n16171 & n16172 ) | ( n16171 & n16173 ) | ( n16172 & n16173 ) ;
  assign n16175 = n16169 & ~n16174 ;
  assign n16176 = n15673 & ~n16169 ;
  assign n16177 = ( n15673 & ~n16172 ) | ( n15673 & n16176 ) | ( ~n16172 & n16176 ) ;
  assign n16178 = n16175 | n16177 ;
  assign n16179 = ~n16166 & n16178 ;
  assign n16180 = n16166 & ~n16178 ;
  assign n16181 = n16179 | n16180 ;
  assign n16182 = n16138 & ~n16181 ;
  assign n16183 = ~n16138 & n16181 ;
  assign n16184 = n16182 | n16183 ;
  assign n16185 = n15852 | n15893 ;
  assign n16186 = n15852 & n15893 ;
  assign n16187 = n16185 & ~n16186 ;
  assign n16188 = n15878 | n16187 ;
  assign n16189 = n15878 & n16187 ;
  assign n16190 = n16188 & ~n16189 ;
  assign n16191 = n16002 | n16004 ;
  assign n16192 = ( n16004 & n16005 ) | ( n16004 & n16191 ) | ( n16005 & n16191 ) ;
  assign n16193 = n15768 | n16012 ;
  assign n16194 = ( n16012 & n16013 ) | ( n16012 & n16193 ) | ( n16013 & n16193 ) ;
  assign n16195 = n16192 | n16194 ;
  assign n16196 = n16192 & n16194 ;
  assign n16197 = n16195 & ~n16196 ;
  assign n16198 = n16190 & n16197 ;
  assign n16199 = n16190 | n16197 ;
  assign n16200 = ~n16198 & n16199 ;
  assign n16201 = ~n16184 & n16200 ;
  assign n16202 = n16184 & ~n16200 ;
  assign n16203 = n16201 | n16202 ;
  assign n16204 = n16089 & n16203 ;
  assign n16205 = n16089 | n16203 ;
  assign n16206 = ~n16204 & n16205 ;
  assign n16207 = n16048 & n16206 ;
  assign n16208 = n15994 & n16206 ;
  assign n16209 = ( n16000 & n16207 ) | ( n16000 & n16208 ) | ( n16207 & n16208 ) ;
  assign n16210 = n16049 & ~n16209 ;
  assign n16211 = n16029 & n16031 ;
  assign n16212 = n16029 & ~n16211 ;
  assign n16213 = n16027 & n16031 ;
  assign n16214 = ~n16029 & n16213 ;
  assign n16215 = n16211 | n16214 ;
  assign n16216 = n16027 | n16031 ;
  assign n16217 = ( n16027 & n16029 ) | ( n16027 & n16216 ) | ( n16029 & n16216 ) ;
  assign n16218 = ( n16212 & n16215 ) | ( n16212 & n16217 ) | ( n16215 & n16217 ) ;
  assign n16219 = n15921 | n15927 ;
  assign n16220 = ( n15923 & n15927 ) | ( n15923 & n16219 ) | ( n15927 & n16219 ) ;
  assign n16221 = n16218 | n16220 ;
  assign n16222 = n15924 | n16218 ;
  assign n16223 = ( n15926 & n16221 ) | ( n15926 & n16222 ) | ( n16221 & n16222 ) ;
  assign n16224 = n16218 & n16220 ;
  assign n16225 = n15924 & n16218 ;
  assign n16226 = ( n15926 & n16224 ) | ( n15926 & n16225 ) | ( n16224 & n16225 ) ;
  assign n16227 = n16223 & ~n16226 ;
  assign n16228 = n15867 | n15918 ;
  assign n16229 = ( n15867 & n15868 ) | ( n15867 & n16228 ) | ( n15868 & n16228 ) ;
  assign n16230 = n16008 | n16020 ;
  assign n16231 = ( n16020 & n16024 ) | ( n16020 & n16230 ) | ( n16024 & n16230 ) ;
  assign n16232 = n16229 & n16231 ;
  assign n16233 = n16229 & ~n16232 ;
  assign n16234 = n15827 | n15836 ;
  assign n16235 = n15827 & n15836 ;
  assign n16236 = n16234 & ~n16235 ;
  assign n16237 = n15970 | n16236 ;
  assign n16238 = n15970 & n16236 ;
  assign n16239 = n16237 & ~n16238 ;
  assign n16240 = n15843 | n15862 ;
  assign n16241 = n15901 | n15915 ;
  assign n16242 = ( n15901 & n15904 ) | ( n15901 & n16241 ) | ( n15904 & n16241 ) ;
  assign n16243 = n16240 | n16242 ;
  assign n16244 = n16240 & n16242 ;
  assign n16245 = n16243 & ~n16244 ;
  assign n16246 = n16239 & n16245 ;
  assign n16247 = n16239 | n16245 ;
  assign n16248 = ~n16246 & n16247 ;
  assign n16249 = ~n16229 & n16231 ;
  assign n16250 = n16248 & n16249 ;
  assign n16251 = ( n16233 & n16248 ) | ( n16233 & n16250 ) | ( n16248 & n16250 ) ;
  assign n16252 = n16248 | n16249 ;
  assign n16253 = n16233 | n16252 ;
  assign n16254 = ~n16251 & n16253 ;
  assign n16255 = n16227 & n16254 ;
  assign n16256 = n16210 | n16255 ;
  assign n16257 = n16227 | n16254 ;
  assign n16258 = n16206 & n16254 ;
  assign n16259 = ( n16206 & n16227 ) | ( n16206 & n16258 ) | ( n16227 & n16258 ) ;
  assign n16260 = ~n16049 & n16259 ;
  assign n16261 = ( n16256 & n16257 ) | ( n16256 & ~n16260 ) | ( n16257 & ~n16260 ) ;
  assign n16262 = ~n16256 & n16261 ;
  assign n16263 = ~n16048 & n16206 ;
  assign n16264 = ~n15994 & n16206 ;
  assign n16265 = ( ~n16000 & n16263 ) | ( ~n16000 & n16264 ) | ( n16263 & n16264 ) ;
  assign n16266 = n16210 | n16265 ;
  assign n16267 = ~n16255 & n16257 ;
  assign n16268 = ~n16255 & n16259 ;
  assign n16269 = ~n16049 & n16268 ;
  assign n16270 = ( n16210 & n16267 ) | ( n16210 & n16269 ) | ( n16267 & n16269 ) ;
  assign n16271 = n16266 & ~n16270 ;
  assign n16272 = n16045 & n16271 ;
  assign n16273 = ( n16045 & n16262 ) | ( n16045 & n16272 ) | ( n16262 & n16272 ) ;
  assign n16274 = n16045 | n16271 ;
  assign n16275 = n16262 | n16274 ;
  assign n16276 = ~n16273 & n16275 ;
  assign n16277 = n15818 & n16040 ;
  assign n16278 = n15818 | n16040 ;
  assign n16279 = n15814 & n16278 ;
  assign n16280 = n16277 | n16279 ;
  assign n16281 = n16277 | n16278 ;
  assign n16282 = ( n15816 & n16277 ) | ( n15816 & n16281 ) | ( n16277 & n16281 ) ;
  assign n16283 = ( n15595 & n16280 ) | ( n15595 & n16282 ) | ( n16280 & n16282 ) ;
  assign n16284 = n16276 & n16283 ;
  assign n16285 = n16276 | n16283 ;
  assign n16286 = ~n16284 & n16285 ;
  assign n16287 = n16275 & n16280 ;
  assign n16288 = n16273 | n16287 ;
  assign n16289 = n16273 | n16275 ;
  assign n16290 = ( n16273 & n16282 ) | ( n16273 & n16289 ) | ( n16282 & n16289 ) ;
  assign n16291 = ( n15595 & n16288 ) | ( n15595 & n16290 ) | ( n16288 & n16290 ) ;
  assign n16292 = ( n16049 & n16206 ) | ( n16049 & n16267 ) | ( n16206 & n16267 ) ;
  assign n16293 = n16232 | n16251 ;
  assign n16294 = n15878 | n16186 ;
  assign n16295 = ( n16186 & n16187 ) | ( n16186 & n16294 ) | ( n16187 & n16294 ) ;
  assign n16296 = n15970 | n16235 ;
  assign n16297 = ( n16235 & n16236 ) | ( n16235 & n16296 ) | ( n16236 & n16296 ) ;
  assign n16298 = n16295 | n16297 ;
  assign n16299 = n16295 & n16297 ;
  assign n16300 = n16298 & ~n16299 ;
  assign n16301 = n16051 | n16065 ;
  assign n16302 = ( n16051 & n16054 ) | ( n16051 & n16301 ) | ( n16054 & n16301 ) ;
  assign n16303 = n16300 | n16302 ;
  assign n16304 = n16300 & n16302 ;
  assign n16305 = n16303 & ~n16304 ;
  assign n16306 = n16078 | n16081 ;
  assign n16307 = ( n16078 & n16079 ) | ( n16078 & n16306 ) | ( n16079 & n16306 ) ;
  assign n16308 = n16305 | n16307 ;
  assign n16309 = n16305 & n16307 ;
  assign n16310 = n16308 & ~n16309 ;
  assign n16311 = ( n16138 & n16181 ) | ( n16138 & n16200 ) | ( n16181 & n16200 ) ;
  assign n16312 = n16310 | n16311 ;
  assign n16313 = n16310 & n16311 ;
  assign n16314 = n16312 & ~n16313 ;
  assign n16315 = n16293 | n16314 ;
  assign n16316 = n16293 & n16314 ;
  assign n16317 = n16315 & ~n16316 ;
  assign n16318 = n16088 | n16203 ;
  assign n16319 = ( n16088 & n16089 ) | ( n16088 & n16318 ) | ( n16089 & n16318 ) ;
  assign n16320 = n16317 & n16319 ;
  assign n16321 = n16317 | n16319 ;
  assign n16322 = ~n16320 & n16321 ;
  assign n16323 = n16097 | n16128 ;
  assign n16324 = n16097 & n16128 ;
  assign n16325 = n16323 & ~n16324 ;
  assign n16326 = n16112 | n16325 ;
  assign n16327 = n16112 & n16325 ;
  assign n16328 = n16326 & ~n16327 ;
  assign n16329 = n16163 | n16178 ;
  assign n16330 = ( n16163 & n16166 ) | ( n16163 & n16329 ) | ( n16166 & n16329 ) ;
  assign n16331 = n16117 | n16135 ;
  assign n16332 = ( n16117 & n16120 ) | ( n16117 & n16331 ) | ( n16120 & n16331 ) ;
  assign n16333 = n16330 | n16332 ;
  assign n16334 = n16330 & n16332 ;
  assign n16335 = n16333 & ~n16334 ;
  assign n16336 = n16328 & n16335 ;
  assign n16337 = n16328 | n16335 ;
  assign n16338 = ~n16336 & n16337 ;
  assign n16370 = n16190 | n16196 ;
  assign n16371 = ( n16196 & n16197 ) | ( n16196 & n16370 ) | ( n16197 & n16370 ) ;
  assign n16339 = x24 & x61 ;
  assign n16340 = n16154 & n16339 ;
  assign n16341 = ( n16153 & n16339 ) | ( n16153 & n16340 ) | ( n16339 & n16340 ) ;
  assign n16342 = n16154 | n16339 ;
  assign n16343 = n16153 | n16342 ;
  assign n16344 = ~n16341 & n16343 ;
  assign n16345 = n16141 | n16145 ;
  assign n16346 = n16344 | n16345 ;
  assign n16347 = n16344 & n16345 ;
  assign n16348 = n16346 & ~n16347 ;
  assign n16349 = n16061 | n16174 ;
  assign n16350 = n16061 & n16174 ;
  assign n16351 = n16349 & ~n16350 ;
  assign n16352 = n2724 & n10975 ;
  assign n16353 = n2511 & n10370 ;
  assign n16354 = n16352 | n16353 ;
  assign n16355 = n2267 & n9831 ;
  assign n16356 = x60 & n16355 ;
  assign n16357 = ( x60 & ~n16354 ) | ( x60 & n16356 ) | ( ~n16354 & n16356 ) ;
  assign n16358 = x25 & n16357 ;
  assign n16359 = n16354 | n16355 ;
  assign n16360 = x27 & x58 ;
  assign n16361 = ( n9066 & ~n16355 ) | ( n9066 & n16360 ) | ( ~n16355 & n16360 ) ;
  assign n16362 = n9066 & n16360 ;
  assign n16363 = ( ~n16354 & n16361 ) | ( ~n16354 & n16362 ) | ( n16361 & n16362 ) ;
  assign n16364 = ~n16359 & n16363 ;
  assign n16365 = n16358 | n16364 ;
  assign n16366 = n16351 & n16365 ;
  assign n16367 = n16351 & ~n16366 ;
  assign n16368 = n16365 & ~n16366 ;
  assign n16369 = n16367 | n16368 ;
  assign n16372 = ( n16348 & ~n16369 ) | ( n16348 & n16371 ) | ( ~n16369 & n16371 ) ;
  assign n16373 = ( ~n16348 & n16369 ) | ( ~n16348 & n16371 ) | ( n16369 & n16371 ) ;
  assign n16374 = ( ~n16371 & n16372 ) | ( ~n16371 & n16373 ) | ( n16372 & n16373 ) ;
  assign n16375 = n16338 & n16374 ;
  assign n16376 = n16338 & ~n16375 ;
  assign n16377 = ~n16338 & n16374 ;
  assign n16378 = n4318 & n7874 ;
  assign n16379 = n3321 & n8161 ;
  assign n16380 = n16378 | n16379 ;
  assign n16381 = n4530 & n7567 ;
  assign n16382 = x53 & n16381 ;
  assign n16383 = ( x53 & ~n16380 ) | ( x53 & n16382 ) | ( ~n16380 & n16382 ) ;
  assign n16384 = x32 & n16383 ;
  assign n16385 = n16380 | n16381 ;
  assign n16386 = x33 & x52 ;
  assign n16387 = x34 & x51 ;
  assign n16388 = ( ~n16381 & n16386 ) | ( ~n16381 & n16387 ) | ( n16386 & n16387 ) ;
  assign n16389 = n16386 & n16387 ;
  assign n16390 = ( ~n16380 & n16388 ) | ( ~n16380 & n16389 ) | ( n16388 & n16389 ) ;
  assign n16391 = ~n16385 & n16390 ;
  assign n16392 = n16384 | n16391 ;
  assign n16393 = x22 & x63 ;
  assign n16394 = x28 & x57 ;
  assign n16395 = n16393 | n16394 ;
  assign n16396 = x35 & x50 ;
  assign n16397 = ( n16393 & n16394 ) | ( n16393 & n16396 ) | ( n16394 & n16396 ) ;
  assign n16398 = n16395 & ~n16397 ;
  assign n16399 = n16393 & n16394 ;
  assign n16400 = n16396 & ~n16399 ;
  assign n16401 = ~n16395 & n16396 ;
  assign n16402 = ( n16396 & ~n16400 ) | ( n16396 & n16401 ) | ( ~n16400 & n16401 ) ;
  assign n16403 = n16398 | n16402 ;
  assign n16404 = n16392 & n16403 ;
  assign n16405 = n16392 & ~n16404 ;
  assign n16406 = n4350 & n8407 ;
  assign n16407 = n4555 & n5975 ;
  assign n16408 = n16406 | n16407 ;
  assign n16409 = n5813 & n6093 ;
  assign n16410 = x46 & n16409 ;
  assign n16411 = ( x46 & ~n16408 ) | ( x46 & n16410 ) | ( ~n16408 & n16410 ) ;
  assign n16412 = x39 & n16411 ;
  assign n16413 = n16408 | n16409 ;
  assign n16414 = x40 & x45 ;
  assign n16415 = x41 & x44 ;
  assign n16416 = ( ~n16409 & n16414 ) | ( ~n16409 & n16415 ) | ( n16414 & n16415 ) ;
  assign n16417 = n16414 & n16415 ;
  assign n16418 = ( ~n16408 & n16416 ) | ( ~n16408 & n16417 ) | ( n16416 & n16417 ) ;
  assign n16419 = ~n16413 & n16418 ;
  assign n16420 = n16412 | n16419 ;
  assign n16421 = ~n16392 & n16403 ;
  assign n16422 = n16420 & ~n16421 ;
  assign n16423 = ~n16405 & n16422 ;
  assign n16424 = ~n16420 & n16421 ;
  assign n16425 = ( n16405 & ~n16420 ) | ( n16405 & n16424 ) | ( ~n16420 & n16424 ) ;
  assign n16426 = n16423 | n16425 ;
  assign n16427 = n3731 & n6757 ;
  assign n16428 = n3770 & n6759 ;
  assign n16429 = n16427 | n16428 ;
  assign n16430 = n4857 & n6762 ;
  assign n16431 = x49 & n16430 ;
  assign n16432 = ( x49 & ~n16429 ) | ( x49 & n16431 ) | ( ~n16429 & n16431 ) ;
  assign n16433 = x36 & n16432 ;
  assign n16434 = n16429 | n16430 ;
  assign n16435 = x37 & x48 ;
  assign n16436 = x38 & x47 ;
  assign n16437 = ( ~n16430 & n16435 ) | ( ~n16430 & n16436 ) | ( n16435 & n16436 ) ;
  assign n16438 = n16435 & n16436 ;
  assign n16439 = ( ~n16429 & n16437 ) | ( ~n16429 & n16438 ) | ( n16437 & n16438 ) ;
  assign n16440 = ~n16434 & n16439 ;
  assign n16441 = n16433 | n16440 ;
  assign n16442 = x43 & x62 ;
  assign n16443 = x23 & n16442 ;
  assign n16444 = n5407 & n16443 ;
  assign n16445 = n5407 & ~n16443 ;
  assign n16446 = n16443 | n16445 ;
  assign n16447 = x23 & x62 ;
  assign n16448 = ( x43 & ~n16443 ) | ( x43 & n16447 ) | ( ~n16443 & n16447 ) ;
  assign n16449 = x43 & n16447 ;
  assign n16450 = ( ~n16445 & n16448 ) | ( ~n16445 & n16449 ) | ( n16448 & n16449 ) ;
  assign n16451 = ~n16446 & n16450 ;
  assign n16452 = n16444 | n16451 ;
  assign n16453 = n16441 & n16452 ;
  assign n16454 = n16441 & ~n16453 ;
  assign n16455 = n3595 & n8146 ;
  assign n16456 = n2709 & n10013 ;
  assign n16457 = n16455 | n16456 ;
  assign n16458 = n2965 & n8357 ;
  assign n16459 = x56 & n16458 ;
  assign n16460 = ( x56 & ~n16457 ) | ( x56 & n16459 ) | ( ~n16457 & n16459 ) ;
  assign n16461 = x29 & n16460 ;
  assign n16462 = n16457 | n16458 ;
  assign n16463 = x30 & x55 ;
  assign n16464 = x31 & x54 ;
  assign n16465 = ( ~n16458 & n16463 ) | ( ~n16458 & n16464 ) | ( n16463 & n16464 ) ;
  assign n16466 = n16463 & n16464 ;
  assign n16467 = ( ~n16457 & n16465 ) | ( ~n16457 & n16466 ) | ( n16465 & n16466 ) ;
  assign n16468 = ~n16462 & n16467 ;
  assign n16469 = n16461 | n16468 ;
  assign n16470 = ~n16441 & n16452 ;
  assign n16471 = n16469 & n16470 ;
  assign n16472 = ( n16454 & n16469 ) | ( n16454 & n16471 ) | ( n16469 & n16471 ) ;
  assign n16473 = n16469 | n16470 ;
  assign n16474 = n16454 | n16473 ;
  assign n16475 = ~n16472 & n16474 ;
  assign n16476 = n16426 & ~n16475 ;
  assign n16477 = ~n16426 & n16475 ;
  assign n16478 = n16476 | n16477 ;
  assign n16479 = n16239 | n16244 ;
  assign n16480 = ( n16244 & n16245 ) | ( n16244 & n16479 ) | ( n16245 & n16479 ) ;
  assign n16481 = n16478 | n16480 ;
  assign n16482 = n16478 & n16480 ;
  assign n16483 = n16481 & ~n16482 ;
  assign n16484 = ~n16377 & n16483 ;
  assign n16485 = ~n16376 & n16484 ;
  assign n16486 = n16377 & ~n16483 ;
  assign n16487 = ( n16376 & ~n16483 ) | ( n16376 & n16486 ) | ( ~n16483 & n16486 ) ;
  assign n16488 = n16485 | n16487 ;
  assign n16489 = n16226 | n16254 ;
  assign n16490 = ( n16226 & n16227 ) | ( n16226 & n16489 ) | ( n16227 & n16489 ) ;
  assign n16491 = ( n16322 & n16488 ) | ( n16322 & ~n16490 ) | ( n16488 & ~n16490 ) ;
  assign n16492 = ( n16322 & ~n16488 ) | ( n16322 & n16490 ) | ( ~n16488 & n16490 ) ;
  assign n16493 = ( ~n16322 & n16491 ) | ( ~n16322 & n16492 ) | ( n16491 & n16492 ) ;
  assign n16494 = ( n16291 & ~n16292 ) | ( n16291 & n16493 ) | ( ~n16292 & n16493 ) ;
  assign n16495 = ( n16292 & ~n16493 ) | ( n16292 & n16494 ) | ( ~n16493 & n16494 ) ;
  assign n16496 = ( ~n16291 & n16494 ) | ( ~n16291 & n16495 ) | ( n16494 & n16495 ) ;
  assign n16630 = n16316 | n16319 ;
  assign n16631 = ( n16316 & n16317 ) | ( n16316 & n16630 ) | ( n16317 & n16630 ) ;
  assign n16497 = n16405 | n16421 ;
  assign n16498 = n16350 | n16366 ;
  assign n16499 = n16404 | n16420 ;
  assign n16500 = n16498 & n16499 ;
  assign n16501 = n16404 & n16498 ;
  assign n16502 = ( n16497 & n16500 ) | ( n16497 & n16501 ) | ( n16500 & n16501 ) ;
  assign n16503 = n16498 | n16499 ;
  assign n16504 = n16404 | n16498 ;
  assign n16505 = ( n16497 & n16503 ) | ( n16497 & n16504 ) | ( n16503 & n16504 ) ;
  assign n16506 = ~n16502 & n16505 ;
  assign n16507 = n16453 | n16472 ;
  assign n16508 = n16506 | n16507 ;
  assign n16509 = n16506 & n16507 ;
  assign n16510 = n16508 & ~n16509 ;
  assign n16511 = n16413 | n16462 ;
  assign n16512 = n16413 & n16462 ;
  assign n16513 = n16511 & ~n16512 ;
  assign n16514 = n16434 | n16513 ;
  assign n16515 = n16434 & n16513 ;
  assign n16516 = n16514 & ~n16515 ;
  assign n16517 = n16359 | n16385 ;
  assign n16518 = n16359 & n16385 ;
  assign n16519 = n16517 & ~n16518 ;
  assign n16520 = n16397 | n16519 ;
  assign n16521 = n16397 & n16519 ;
  assign n16522 = n16520 & ~n16521 ;
  assign n16523 = n16516 & n16522 ;
  assign n16524 = n16516 | n16522 ;
  assign n16525 = ~n16523 & n16524 ;
  assign n16526 = n16299 | n16302 ;
  assign n16527 = ( n16299 & n16300 ) | ( n16299 & n16526 ) | ( n16300 & n16526 ) ;
  assign n16528 = n16525 & n16527 ;
  assign n16529 = n16525 | n16527 ;
  assign n16530 = ~n16528 & n16529 ;
  assign n16531 = n16510 & n16530 ;
  assign n16532 = n16510 | n16530 ;
  assign n16533 = ~n16531 & n16532 ;
  assign n16534 = n3129 & n7874 ;
  assign n16535 = n4530 & n8161 ;
  assign n16536 = n16534 | n16535 ;
  assign n16537 = n3483 & n7567 ;
  assign n16538 = x53 & n16537 ;
  assign n16539 = ( x53 & ~n16536 ) | ( x53 & n16538 ) | ( ~n16536 & n16538 ) ;
  assign n16540 = x33 & n16539 ;
  assign n16541 = n16536 | n16537 ;
  assign n16542 = x34 & x52 ;
  assign n16543 = x35 & x51 ;
  assign n16544 = ( ~n16537 & n16542 ) | ( ~n16537 & n16543 ) | ( n16542 & n16543 ) ;
  assign n16545 = n16542 & n16543 ;
  assign n16546 = ( ~n16536 & n16544 ) | ( ~n16536 & n16545 ) | ( n16544 & n16545 ) ;
  assign n16547 = ~n16541 & n16546 ;
  assign n16548 = n16540 | n16547 ;
  assign n16549 = x23 & x63 ;
  assign n16550 = n3770 & n6834 ;
  assign n16551 = x36 & x50 ;
  assign n16552 = x37 & x49 ;
  assign n16553 = n16551 | n16552 ;
  assign n16554 = ( n16549 & n16550 ) | ( n16549 & ~n16553 ) | ( n16550 & ~n16553 ) ;
  assign n16555 = n16549 & ~n16554 ;
  assign n16556 = ~n16550 & n16553 ;
  assign n16557 = n16549 | n16556 ;
  assign n16558 = ~n16555 & n16557 ;
  assign n16559 = n16548 & n16558 ;
  assign n16560 = n16548 & ~n16559 ;
  assign n16561 = n13674 | n15963 ;
  assign n16562 = n3595 & n12860 ;
  assign n16563 = n7528 & ~n16562 ;
  assign n16564 = n16561 | n16562 ;
  assign n16565 = ( n16562 & n16563 ) | ( n16562 & n16564 ) | ( n16563 & n16564 ) ;
  assign n16566 = n16561 & ~n16565 ;
  assign n16567 = n7528 & ~n16561 ;
  assign n16568 = ( n7528 & ~n16563 ) | ( n7528 & n16567 ) | ( ~n16563 & n16567 ) ;
  assign n16569 = n16566 | n16568 ;
  assign n16570 = ~n16548 & n16558 ;
  assign n16571 = n16569 & ~n16570 ;
  assign n16572 = ~n16560 & n16571 ;
  assign n16573 = ~n16569 & n16570 ;
  assign n16574 = ( n16560 & ~n16569 ) | ( n16560 & n16573 ) | ( ~n16569 & n16573 ) ;
  assign n16575 = n16572 | n16574 ;
  assign n16576 = n2895 & n10975 ;
  assign n16577 = n2267 & n10370 ;
  assign n16578 = n16576 | n16577 ;
  assign n16579 = n2372 & n9831 ;
  assign n16580 = x60 & n16579 ;
  assign n16581 = ( x60 & ~n16578 ) | ( x60 & n16580 ) | ( ~n16578 & n16580 ) ;
  assign n16582 = x26 & n16581 ;
  assign n16583 = n16578 | n16579 ;
  assign n16584 = x27 & x59 ;
  assign n16585 = x28 & x58 ;
  assign n16586 = ( ~n16579 & n16584 ) | ( ~n16579 & n16585 ) | ( n16584 & n16585 ) ;
  assign n16587 = n16584 & n16585 ;
  assign n16588 = ( ~n16578 & n16586 ) | ( ~n16578 & n16587 ) | ( n16586 & n16587 ) ;
  assign n16589 = ~n16583 & n16588 ;
  assign n16590 = n16582 | n16589 ;
  assign n16591 = x32 & x54 ;
  assign n16592 = n4969 & n16591 ;
  assign n16593 = n5102 & n16591 ;
  assign n16594 = n5710 & n6093 ;
  assign n16595 = n16593 | n16594 ;
  assign n16596 = n5102 & n16592 ;
  assign n16597 = ( n5102 & ~n16595 ) | ( n5102 & n16596 ) | ( ~n16595 & n16596 ) ;
  assign n16598 = ( n4969 & n16591 ) | ( n4969 & ~n16595 ) | ( n16591 & ~n16595 ) ;
  assign n16599 = ( ~n16592 & n16597 ) | ( ~n16592 & n16598 ) | ( n16597 & n16598 ) ;
  assign n16600 = n16590 & n16599 ;
  assign n16601 = n16590 & ~n16600 ;
  assign n16602 = x39 & x47 ;
  assign n16603 = n7654 | n16602 ;
  assign n16604 = n4555 & n6147 ;
  assign n16605 = x30 & x56 ;
  assign n16606 = ~n16604 & n16605 ;
  assign n16607 = n16603 | n16604 ;
  assign n16608 = ( n16604 & n16606 ) | ( n16604 & n16607 ) | ( n16606 & n16607 ) ;
  assign n16609 = n16603 & ~n16608 ;
  assign n16610 = ( ~n16603 & n16604 ) | ( ~n16603 & n16605 ) | ( n16604 & n16605 ) ;
  assign n16611 = n16605 & n16610 ;
  assign n16612 = n16609 | n16611 ;
  assign n16613 = ~n16590 & n16599 ;
  assign n16614 = n16612 & n16613 ;
  assign n16615 = ( n16601 & n16612 ) | ( n16601 & n16614 ) | ( n16612 & n16614 ) ;
  assign n16616 = n16612 | n16613 ;
  assign n16617 = n16601 | n16616 ;
  assign n16618 = ~n16615 & n16617 ;
  assign n16619 = n16575 | n16618 ;
  assign n16620 = n16575 & n16618 ;
  assign n16621 = n16619 & ~n16620 ;
  assign n16622 = n16328 | n16334 ;
  assign n16623 = ( n16334 & n16335 ) | ( n16334 & n16622 ) | ( n16335 & n16622 ) ;
  assign n16624 = n16621 & n16623 ;
  assign n16625 = n16621 | n16623 ;
  assign n16626 = ~n16624 & n16625 ;
  assign n16627 = n16533 & n16626 ;
  assign n16628 = n16533 | n16626 ;
  assign n16629 = ~n16627 & n16628 ;
  assign n16632 = n16629 & n16631 ;
  assign n16633 = n16631 & ~n16632 ;
  assign n16634 = n16377 & n16483 ;
  assign n16635 = ( n16376 & n16483 ) | ( n16376 & n16634 ) | ( n16483 & n16634 ) ;
  assign n16636 = n16305 | n16311 ;
  assign n16637 = ( n16307 & n16311 ) | ( n16307 & n16636 ) | ( n16311 & n16636 ) ;
  assign n16638 = ( n16309 & n16310 ) | ( n16309 & n16637 ) | ( n16310 & n16637 ) ;
  assign n16639 = n16375 | n16638 ;
  assign n16640 = n16635 | n16639 ;
  assign n16641 = n16375 & n16638 ;
  assign n16642 = ( n16635 & n16638 ) | ( n16635 & n16641 ) | ( n16638 & n16641 ) ;
  assign n16643 = n16640 & ~n16642 ;
  assign n16644 = n1912 & n10684 ;
  assign n16645 = x25 & x61 ;
  assign n16646 = x24 & x62 ;
  assign n16647 = n16645 | n16646 ;
  assign n16648 = ~n16644 & n16647 ;
  assign n16649 = n16446 & n16648 ;
  assign n16650 = n16446 & ~n16649 ;
  assign n16651 = ~n16446 & n16648 ;
  assign n16652 = n16650 | n16651 ;
  assign n16653 = n16341 | n16345 ;
  assign n16654 = ( n16341 & n16344 ) | ( n16341 & n16653 ) | ( n16344 & n16653 ) ;
  assign n16655 = n16652 | n16654 ;
  assign n16656 = n16652 & n16654 ;
  assign n16657 = n16655 & ~n16656 ;
  assign n16658 = n16112 | n16324 ;
  assign n16659 = ( n16324 & n16325 ) | ( n16324 & n16658 ) | ( n16325 & n16658 ) ;
  assign n16660 = n16657 | n16659 ;
  assign n16661 = n16657 & n16659 ;
  assign n16662 = n16660 & ~n16661 ;
  assign n16663 = n16348 | n16369 ;
  assign n16664 = n16371 & n16663 ;
  assign n16665 = n16348 & n16369 ;
  assign n16666 = n16664 | n16665 ;
  assign n16667 = n16662 & n16666 ;
  assign n16668 = n16662 | n16666 ;
  assign n16669 = ~n16667 & n16668 ;
  assign n16670 = ( n16426 & n16475 ) | ( n16426 & n16480 ) | ( n16475 & n16480 ) ;
  assign n16671 = n16669 | n16670 ;
  assign n16672 = n16669 & n16670 ;
  assign n16673 = n16671 & ~n16672 ;
  assign n16674 = n16643 & n16673 ;
  assign n16675 = n16643 | n16673 ;
  assign n16676 = ~n16674 & n16675 ;
  assign n16677 = n16629 & ~n16631 ;
  assign n16678 = n16676 | n16677 ;
  assign n16679 = n16633 | n16678 ;
  assign n16680 = n16676 & n16677 ;
  assign n16681 = ( n16633 & n16676 ) | ( n16633 & n16680 ) | ( n16676 & n16680 ) ;
  assign n16682 = n16679 & ~n16681 ;
  assign n16683 = n16488 & n16490 ;
  assign n16684 = n16490 & ~n16683 ;
  assign n16685 = n16488 & ~n16490 ;
  assign n16686 = n16322 & ~n16685 ;
  assign n16687 = ~n16684 & n16686 ;
  assign n16688 = ( n16322 & n16683 ) | ( n16322 & ~n16687 ) | ( n16683 & ~n16687 ) ;
  assign n16689 = n16682 | n16688 ;
  assign n16690 = n16682 & n16688 ;
  assign n16691 = n16689 & ~n16690 ;
  assign n16692 = n16292 & n16493 ;
  assign n16693 = n16292 | n16493 ;
  assign n16694 = n16692 | n16693 ;
  assign n16695 = ( n16289 & n16692 ) | ( n16289 & n16694 ) | ( n16692 & n16694 ) ;
  assign n16696 = n16045 & n16262 ;
  assign n16697 = n16045 & n16693 ;
  assign n16698 = n16692 | n16697 ;
  assign n16699 = n16271 & n16693 ;
  assign n16700 = n16692 | n16699 ;
  assign n16701 = ( n16696 & n16698 ) | ( n16696 & n16700 ) | ( n16698 & n16700 ) ;
  assign n16702 = ( n16282 & n16695 ) | ( n16282 & n16701 ) | ( n16695 & n16701 ) ;
  assign n16703 = ( n16287 & n16694 ) | ( n16287 & n16701 ) | ( n16694 & n16701 ) ;
  assign n16704 = ( n15595 & n16702 ) | ( n15595 & n16703 ) | ( n16702 & n16703 ) ;
  assign n16705 = n16691 | n16704 ;
  assign n16706 = n16689 & n16702 ;
  assign n16707 = n16689 & n16703 ;
  assign n16708 = ( n15595 & n16706 ) | ( n15595 & n16707 ) | ( n16706 & n16707 ) ;
  assign n16709 = ~n16690 & n16708 ;
  assign n16710 = n16705 & ~n16709 ;
  assign n16711 = n16690 | n16707 ;
  assign n16712 = n16689 | n16690 ;
  assign n16713 = ( n16690 & n16702 ) | ( n16690 & n16712 ) | ( n16702 & n16712 ) ;
  assign n16714 = ( n15595 & n16711 ) | ( n15595 & n16713 ) | ( n16711 & n16713 ) ;
  assign n16715 = n16632 | n16681 ;
  assign n16716 = n16560 | n16570 ;
  assign n16717 = n16559 | n16569 ;
  assign n16718 = n16434 | n16512 ;
  assign n16719 = ( n16512 & n16513 ) | ( n16512 & n16718 ) | ( n16513 & n16718 ) ;
  assign n16720 = n16717 & n16719 ;
  assign n16721 = n16559 & n16719 ;
  assign n16722 = ( n16716 & n16720 ) | ( n16716 & n16721 ) | ( n16720 & n16721 ) ;
  assign n16723 = n16717 | n16719 ;
  assign n16724 = n16559 | n16719 ;
  assign n16725 = ( n16716 & n16723 ) | ( n16716 & n16724 ) | ( n16723 & n16724 ) ;
  assign n16726 = ~n16722 & n16725 ;
  assign n16727 = n16600 | n16615 ;
  assign n16728 = n16726 | n16727 ;
  assign n16729 = n16726 & n16727 ;
  assign n16730 = n16728 & ~n16729 ;
  assign n16731 = n16620 | n16621 ;
  assign n16732 = ( n16620 & n16623 ) | ( n16620 & n16731 ) | ( n16623 & n16731 ) ;
  assign n16733 = n16730 & n16732 ;
  assign n16734 = n16730 | n16732 ;
  assign n16735 = ~n16733 & n16734 ;
  assign n16736 = n16667 | n16672 ;
  assign n16737 = n16735 | n16736 ;
  assign n16738 = n16735 & n16736 ;
  assign n16739 = n16737 & ~n16738 ;
  assign n16740 = n16642 | n16673 ;
  assign n16741 = ( n16642 & n16643 ) | ( n16642 & n16740 ) | ( n16643 & n16740 ) ;
  assign n16742 = n16739 & n16741 ;
  assign n16743 = n16739 | n16741 ;
  assign n16744 = ~n16742 & n16743 ;
  assign n16745 = x31 & x56 ;
  assign n16746 = x33 & x54 ;
  assign n16747 = n16745 | n16746 ;
  assign n16748 = n2683 & n8146 ;
  assign n16749 = x40 & x47 ;
  assign n16750 = ~n16748 & n16749 ;
  assign n16751 = n16747 | n16748 ;
  assign n16752 = ( n16748 & n16750 ) | ( n16748 & n16751 ) | ( n16750 & n16751 ) ;
  assign n16753 = n16747 & ~n16752 ;
  assign n16754 = ( ~n16747 & n16748 ) | ( ~n16747 & n16749 ) | ( n16748 & n16749 ) ;
  assign n16755 = n16749 & n16754 ;
  assign n16756 = n16753 | n16755 ;
  assign n16757 = ( x44 & x62 ) | ( x44 & ~n5658 ) | ( x62 & ~n5658 ) ;
  assign n16758 = x25 | x62 ;
  assign n16759 = ~x25 & x44 ;
  assign n16760 = ( n5658 & n16758 ) | ( n5658 & ~n16759 ) | ( n16758 & ~n16759 ) ;
  assign n16761 = ( ~x25 & x44 ) | ( ~x25 & x62 ) | ( x44 & x62 ) ;
  assign n16762 = ( x25 & n5658 ) | ( x25 & ~n16761 ) | ( n5658 & ~n16761 ) ;
  assign n16763 = ( n16757 & ~n16760 ) | ( n16757 & n16762 ) | ( ~n16760 & n16762 ) ;
  assign n16764 = n16755 & n16763 ;
  assign n16765 = ( n16753 & n16763 ) | ( n16753 & n16764 ) | ( n16763 & n16764 ) ;
  assign n16766 = n16756 & ~n16765 ;
  assign n16767 = n16397 | n16518 ;
  assign n16768 = ( n16518 & n16519 ) | ( n16518 & n16767 ) | ( n16519 & n16767 ) ;
  assign n16769 = ~n16755 & n16763 ;
  assign n16770 = ~n16753 & n16769 ;
  assign n16771 = n16768 & n16770 ;
  assign n16772 = ( n16766 & n16768 ) | ( n16766 & n16771 ) | ( n16768 & n16771 ) ;
  assign n16773 = n16768 | n16770 ;
  assign n16774 = n16766 | n16773 ;
  assign n16775 = ~n16772 & n16774 ;
  assign n16776 = n2340 & n10856 ;
  assign n16777 = n6685 & n12770 ;
  assign n16778 = n16776 | n16777 ;
  assign n16779 = n2267 & n10367 ;
  assign n16780 = x63 & n16779 ;
  assign n16781 = ( x63 & ~n16778 ) | ( x63 & n16780 ) | ( ~n16778 & n16780 ) ;
  assign n16782 = x24 & n16781 ;
  assign n16783 = n16778 | n16779 ;
  assign n16784 = x26 & x61 ;
  assign n16785 = x27 & x60 ;
  assign n16786 = ( ~n16779 & n16784 ) | ( ~n16779 & n16785 ) | ( n16784 & n16785 ) ;
  assign n16787 = n16784 & n16785 ;
  assign n16788 = ( ~n16778 & n16786 ) | ( ~n16778 & n16787 ) | ( n16786 & n16787 ) ;
  assign n16789 = ~n16783 & n16788 ;
  assign n16790 = n16782 | n16789 ;
  assign n16791 = n5798 & n6345 ;
  assign n16792 = n4857 & n6834 ;
  assign n16793 = n16791 | n16792 ;
  assign n16794 = n5392 & n6759 ;
  assign n16795 = x50 & n16794 ;
  assign n16796 = ( x50 & ~n16793 ) | ( x50 & n16795 ) | ( ~n16793 & n16795 ) ;
  assign n16797 = x37 & n16796 ;
  assign n16798 = n16793 | n16794 ;
  assign n16799 = x38 & x49 ;
  assign n16800 = x39 & x48 ;
  assign n16801 = ( ~n16794 & n16799 ) | ( ~n16794 & n16800 ) | ( n16799 & n16800 ) ;
  assign n16802 = n16799 & n16800 ;
  assign n16803 = ( ~n16793 & n16801 ) | ( ~n16793 & n16802 ) | ( n16801 & n16802 ) ;
  assign n16804 = ~n16798 & n16803 ;
  assign n16805 = n16797 | n16804 ;
  assign n16806 = n16790 & n16805 ;
  assign n16807 = n16790 & ~n16806 ;
  assign n16808 = n16805 & ~n16806 ;
  assign n16809 = n16807 | n16808 ;
  assign n16810 = x41 & x46 ;
  assign n16811 = x42 & x45 ;
  assign n16812 = n16810 | n16811 ;
  assign n16813 = n5710 & n5975 ;
  assign n16814 = x32 & x55 ;
  assign n16815 = ~n16813 & n16814 ;
  assign n16816 = n16812 | n16813 ;
  assign n16817 = ( n16813 & n16815 ) | ( n16813 & n16816 ) | ( n16815 & n16816 ) ;
  assign n16818 = n16812 & ~n16817 ;
  assign n16819 = ( ~n16812 & n16813 ) | ( ~n16812 & n16814 ) | ( n16813 & n16814 ) ;
  assign n16820 = n16814 & n16819 ;
  assign n16821 = n16818 | n16820 ;
  assign n16822 = ~n16809 & n16821 ;
  assign n16823 = n16775 & n16822 ;
  assign n16824 = n16809 & ~n16821 ;
  assign n16825 = ( n16775 & n16823 ) | ( n16775 & n16824 ) | ( n16823 & n16824 ) ;
  assign n16826 = n16775 | n16822 ;
  assign n16827 = n16824 | n16826 ;
  assign n16828 = ~n16825 & n16827 ;
  assign n16829 = n3280 & n9829 ;
  assign n16830 = x34 & x59 ;
  assign n16831 = n15423 & n16830 ;
  assign n16832 = n16829 | n16831 ;
  assign n16833 = x34 & x53 ;
  assign n16834 = n16170 & n16833 ;
  assign n16835 = x59 & n16834 ;
  assign n16836 = ( x59 & ~n16832 ) | ( x59 & n16835 ) | ( ~n16832 & n16835 ) ;
  assign n16837 = x28 & n16836 ;
  assign n16838 = n16832 | n16834 ;
  assign n16839 = n16170 | n16833 ;
  assign n16840 = x28 | n16839 ;
  assign n16841 = ( n16836 & n16839 ) | ( n16836 & n16840 ) | ( n16839 & n16840 ) ;
  assign n16842 = ( n16837 & ~n16838 ) | ( n16837 & n16841 ) | ( ~n16838 & n16841 ) ;
  assign n16843 = n16644 | n16648 ;
  assign n16844 = ( n16446 & n16644 ) | ( n16446 & n16843 ) | ( n16644 & n16843 ) ;
  assign n16845 = n16842 & ~n16844 ;
  assign n16846 = ~n16842 & n16844 ;
  assign n16847 = n16845 | n16846 ;
  assign n16848 = x29 & x58 ;
  assign n16849 = x36 & x51 ;
  assign n16850 = n16848 & n16849 ;
  assign n16851 = n4078 & n7567 ;
  assign n16852 = x35 & x58 ;
  assign n16853 = n15424 & n16852 ;
  assign n16854 = n16851 | n16853 ;
  assign n16855 = x52 & n16850 ;
  assign n16856 = ( x52 & ~n16854 ) | ( x52 & n16855 ) | ( ~n16854 & n16855 ) ;
  assign n16857 = x35 & n16856 ;
  assign n16858 = ( n16848 & n16849 ) | ( n16848 & ~n16854 ) | ( n16849 & ~n16854 ) ;
  assign n16859 = ( ~n16850 & n16857 ) | ( ~n16850 & n16858 ) | ( n16857 & n16858 ) ;
  assign n16860 = n16847 & n16859 ;
  assign n16861 = n16847 | n16859 ;
  assign n16862 = ~n16860 & n16861 ;
  assign n16863 = n16828 & n16862 ;
  assign n16864 = n16828 | n16862 ;
  assign n16865 = ~n16863 & n16864 ;
  assign n16866 = n16531 & n16865 ;
  assign n16867 = ( n16627 & n16865 ) | ( n16627 & n16866 ) | ( n16865 & n16866 ) ;
  assign n16868 = n16531 | n16865 ;
  assign n16869 = n16627 | n16868 ;
  assign n16870 = ~n16867 & n16869 ;
  assign n16871 = n16523 | n16528 ;
  assign n16872 = n16502 | n16507 ;
  assign n16873 = ( n16502 & n16506 ) | ( n16502 & n16872 ) | ( n16506 & n16872 ) ;
  assign n16874 = n16871 | n16873 ;
  assign n16875 = n16871 & n16873 ;
  assign n16876 = n16874 & ~n16875 ;
  assign n16877 = n16592 | n16595 ;
  assign n16878 = n16608 | n16877 ;
  assign n16879 = n16608 & n16877 ;
  assign n16880 = n16878 & ~n16879 ;
  assign n16881 = n16565 | n16880 ;
  assign n16882 = n16565 & n16880 ;
  assign n16883 = n16881 & ~n16882 ;
  assign n16884 = n16541 | n16583 ;
  assign n16885 = n16541 & n16583 ;
  assign n16886 = n16884 & ~n16885 ;
  assign n16887 = n16549 | n16550 ;
  assign n16888 = ( n16550 & ~n16554 ) | ( n16550 & n16887 ) | ( ~n16554 & n16887 ) ;
  assign n16889 = n16886 | n16888 ;
  assign n16890 = n16886 & n16888 ;
  assign n16891 = n16889 & ~n16890 ;
  assign n16892 = n16883 | n16891 ;
  assign n16893 = n16883 & n16891 ;
  assign n16894 = n16892 & ~n16893 ;
  assign n16895 = n16656 | n16659 ;
  assign n16896 = ( n16656 & n16657 ) | ( n16656 & n16895 ) | ( n16657 & n16895 ) ;
  assign n16897 = n16894 & n16896 ;
  assign n16898 = n16894 | n16896 ;
  assign n16899 = ~n16897 & n16898 ;
  assign n16900 = n16876 & n16899 ;
  assign n16901 = n16876 | n16899 ;
  assign n16902 = ~n16900 & n16901 ;
  assign n16903 = ~n16870 & n16902 ;
  assign n16904 = n16870 & ~n16902 ;
  assign n16905 = n16903 | n16904 ;
  assign n16906 = n16744 | n16905 ;
  assign n16907 = n16744 & n16905 ;
  assign n16908 = n16906 & ~n16907 ;
  assign n16909 = ( n16714 & n16715 ) | ( n16714 & ~n16908 ) | ( n16715 & ~n16908 ) ;
  assign n16910 = ( ~n16715 & n16908 ) | ( ~n16715 & n16909 ) | ( n16908 & n16909 ) ;
  assign n16911 = ( ~n16714 & n16909 ) | ( ~n16714 & n16910 ) | ( n16909 & n16910 ) ;
  assign n16912 = n16715 & n16908 ;
  assign n16913 = n16715 | n16908 ;
  assign n16914 = n16912 | n16913 ;
  assign n16915 = ( n16690 & n16912 ) | ( n16690 & n16914 ) | ( n16912 & n16914 ) ;
  assign n16916 = ( n16707 & n16914 ) | ( n16707 & n16915 ) | ( n16914 & n16915 ) ;
  assign n16917 = ( n16712 & n16912 ) | ( n16712 & n16914 ) | ( n16912 & n16914 ) ;
  assign n16918 = ( n16701 & n16915 ) | ( n16701 & n16917 ) | ( n16915 & n16917 ) ;
  assign n16919 = ( n16282 & n16915 ) | ( n16282 & n16917 ) | ( n16915 & n16917 ) ;
  assign n16920 = ( n16695 & n16918 ) | ( n16695 & n16919 ) | ( n16918 & n16919 ) ;
  assign n16921 = ( n15595 & n16916 ) | ( n15595 & n16920 ) | ( n16916 & n16920 ) ;
  assign n16922 = ( n16842 & n16844 ) | ( n16842 & n16859 ) | ( n16844 & n16859 ) ;
  assign n16923 = n16885 | n16888 ;
  assign n16924 = ( n16885 & n16886 ) | ( n16885 & n16923 ) | ( n16886 & n16923 ) ;
  assign n16925 = n16922 | n16924 ;
  assign n16926 = n16922 & n16924 ;
  assign n16927 = n16925 & ~n16926 ;
  assign n16928 = n16806 | n16821 ;
  assign n16929 = ( n16806 & n16809 ) | ( n16806 & n16928 ) | ( n16809 & n16928 ) ;
  assign n16930 = n16927 | n16929 ;
  assign n16931 = n16927 & n16929 ;
  assign n16932 = n16930 & ~n16931 ;
  assign n16933 = n16824 | n16862 ;
  assign n16934 = n16775 | n16862 ;
  assign n16935 = ( n16823 & n16933 ) | ( n16823 & n16934 ) | ( n16933 & n16934 ) ;
  assign n16936 = n16932 & n16935 ;
  assign n16937 = n16825 & n16932 ;
  assign n16938 = ( n16828 & n16936 ) | ( n16828 & n16937 ) | ( n16936 & n16937 ) ;
  assign n16939 = n16932 | n16935 ;
  assign n16940 = n16825 | n16932 ;
  assign n16941 = ( n16828 & n16939 ) | ( n16828 & n16940 ) | ( n16939 & n16940 ) ;
  assign n16942 = ~n16938 & n16941 ;
  assign n16943 = n16875 | n16899 ;
  assign n16944 = ( n16875 & n16876 ) | ( n16875 & n16943 ) | ( n16876 & n16943 ) ;
  assign n16945 = n16942 & n16944 ;
  assign n16946 = n16942 | n16944 ;
  assign n16947 = ~n16945 & n16946 ;
  assign n16948 = n16867 | n16902 ;
  assign n16949 = ( n16867 & n16870 ) | ( n16867 & n16948 ) | ( n16870 & n16948 ) ;
  assign n16950 = n16947 & n16949 ;
  assign n16951 = n16947 | n16949 ;
  assign n16952 = ~n16950 & n16951 ;
  assign n16953 = n16893 | n16897 ;
  assign n16954 = n16722 | n16727 ;
  assign n16955 = ( n16722 & n16726 ) | ( n16722 & n16954 ) | ( n16726 & n16954 ) ;
  assign n16956 = n16953 | n16955 ;
  assign n16957 = n16953 & n16955 ;
  assign n16958 = n16956 & ~n16957 ;
  assign n16959 = n16783 | n16838 ;
  assign n16960 = n16783 & n16838 ;
  assign n16961 = n16959 & ~n16960 ;
  assign n16962 = n16798 | n16961 ;
  assign n16963 = n16798 & n16961 ;
  assign n16964 = n16962 & ~n16963 ;
  assign n16965 = n16850 | n16854 ;
  assign n16966 = n16752 | n16965 ;
  assign n16967 = n16752 & n16965 ;
  assign n16968 = n16966 & ~n16967 ;
  assign n16969 = x33 & x55 ;
  assign n16970 = x34 & x54 ;
  assign n16971 = n16969 | n16970 ;
  assign n16972 = n4530 & n8357 ;
  assign n16973 = n5104 & ~n16972 ;
  assign n16974 = n16971 | n16972 ;
  assign n16975 = ( n16972 & n16973 ) | ( n16972 & n16974 ) | ( n16973 & n16974 ) ;
  assign n16976 = n16971 & ~n16975 ;
  assign n16977 = n5104 & ~n16971 ;
  assign n16978 = ( n5104 & ~n16973 ) | ( n5104 & n16977 ) | ( ~n16973 & n16977 ) ;
  assign n16979 = n16976 | n16978 ;
  assign n16980 = n16968 & n16979 ;
  assign n16981 = n16968 & ~n16980 ;
  assign n16982 = n16979 & ~n16980 ;
  assign n16983 = n16981 | n16982 ;
  assign n16984 = n16765 | n16768 ;
  assign n16985 = n16765 | n16766 ;
  assign n16986 = ( n16771 & n16984 ) | ( n16771 & n16985 ) | ( n16984 & n16985 ) ;
  assign n16987 = n16983 | n16986 ;
  assign n16988 = n16983 & n16986 ;
  assign n16989 = n16987 & ~n16988 ;
  assign n16990 = n16964 & n16989 ;
  assign n16991 = n16964 | n16989 ;
  assign n16992 = ~n16990 & n16991 ;
  assign n16993 = n16958 & n16992 ;
  assign n16994 = n16958 | n16992 ;
  assign n16995 = ~n16993 & n16994 ;
  assign n16996 = x30 & x58 ;
  assign n16997 = x32 & x56 ;
  assign n16998 = n16996 | n16997 ;
  assign n16999 = n2546 & n8708 ;
  assign n17000 = n8070 & ~n16999 ;
  assign n17001 = n16998 | n16999 ;
  assign n17002 = ( n16999 & n17000 ) | ( n16999 & n17001 ) | ( n17000 & n17001 ) ;
  assign n17003 = n16998 & ~n17002 ;
  assign n17004 = n8070 & ~n16998 ;
  assign n17005 = ( n8070 & ~n17000 ) | ( n8070 & n17004 ) | ( ~n17000 & n17004 ) ;
  assign n17006 = n17003 | n17005 ;
  assign n17007 = x38 & x50 ;
  assign n17008 = x39 & x49 ;
  assign n17009 = n17007 | n17008 ;
  assign n17010 = n5392 & n6834 ;
  assign n17011 = n17009 | n17010 ;
  assign n17012 = x29 & x59 ;
  assign n17013 = ( ~n17010 & n17011 ) | ( ~n17010 & n17012 ) | ( n17011 & n17012 ) ;
  assign n17014 = ( n17010 & n17011 ) | ( n17010 & ~n17012 ) | ( n17011 & ~n17012 ) ;
  assign n17015 = ( ~n17011 & n17013 ) | ( ~n17011 & n17014 ) | ( n17013 & n17014 ) ;
  assign n17016 = n17006 & n17015 ;
  assign n17017 = n17006 & ~n17016 ;
  assign n17018 = ~n17006 & n17015 ;
  assign n17019 = n16565 | n16879 ;
  assign n17020 = ( n16879 & n16880 ) | ( n16879 & n17019 ) | ( n16880 & n17019 ) ;
  assign n17021 = n17018 | n17020 ;
  assign n17022 = n17017 | n17021 ;
  assign n17023 = n17018 & n17020 ;
  assign n17024 = ( n17017 & n17020 ) | ( n17017 & n17023 ) | ( n17020 & n17023 ) ;
  assign n17025 = n17022 & ~n17024 ;
  assign n17026 = x44 & x62 ;
  assign n17027 = x25 & n17026 ;
  assign n17028 = n5658 & ~n17027 ;
  assign n17029 = x25 & x63 ;
  assign n17030 = n17027 & n17029 ;
  assign n17031 = ( n17028 & n17029 ) | ( n17028 & n17030 ) | ( n17029 & n17030 ) ;
  assign n17032 = n17027 | n17029 ;
  assign n17033 = n17028 | n17032 ;
  assign n17034 = ~n17031 & n17033 ;
  assign n17035 = n16817 | n17034 ;
  assign n17036 = n16817 & n17034 ;
  assign n17037 = n17035 & ~n17036 ;
  assign n17038 = n17025 & n17037 ;
  assign n17039 = n17025 | n17037 ;
  assign n17040 = ~n17038 & n17039 ;
  assign n17041 = n2895 & n9931 ;
  assign n17042 = n2267 & n10684 ;
  assign n17043 = n17041 | n17042 ;
  assign n17044 = n2372 & n10367 ;
  assign n17045 = x62 & n17044 ;
  assign n17046 = ( x62 & ~n17043 ) | ( x62 & n17045 ) | ( ~n17043 & n17045 ) ;
  assign n17047 = x26 & n17046 ;
  assign n17048 = n17043 | n17044 ;
  assign n17049 = x27 & x61 ;
  assign n17050 = x28 & x60 ;
  assign n17051 = ( ~n17044 & n17049 ) | ( ~n17044 & n17050 ) | ( n17049 & n17050 ) ;
  assign n17052 = n17049 & n17050 ;
  assign n17053 = ( ~n17043 & n17051 ) | ( ~n17043 & n17052 ) | ( n17051 & n17052 ) ;
  assign n17054 = ~n17048 & n17053 ;
  assign n17055 = n17047 | n17054 ;
  assign n17056 = x42 & x46 ;
  assign n17057 = x41 & x47 ;
  assign n17058 = n17056 | n17057 ;
  assign n17059 = n5710 & n6147 ;
  assign n17060 = x31 & x57 ;
  assign n17061 = ~n17059 & n17060 ;
  assign n17062 = n17058 | n17059 ;
  assign n17063 = ( n17059 & n17061 ) | ( n17059 & n17062 ) | ( n17061 & n17062 ) ;
  assign n17064 = n17058 & ~n17063 ;
  assign n17065 = ( ~n17058 & n17059 ) | ( ~n17058 & n17060 ) | ( n17059 & n17060 ) ;
  assign n17066 = n17060 & n17065 ;
  assign n17067 = n17064 | n17066 ;
  assign n17068 = n17055 & n17067 ;
  assign n17069 = n17055 & ~n17068 ;
  assign n17070 = n17067 & ~n17068 ;
  assign n17071 = n17069 | n17070 ;
  assign n17072 = n5417 & n7874 ;
  assign n17073 = n4078 & n8161 ;
  assign n17074 = n17072 | n17073 ;
  assign n17075 = n3770 & n7567 ;
  assign n17076 = x53 & n17075 ;
  assign n17077 = ( x53 & ~n17074 ) | ( x53 & n17076 ) | ( ~n17074 & n17076 ) ;
  assign n17078 = x35 & n17077 ;
  assign n17079 = n17074 | n17075 ;
  assign n17080 = x37 & x51 ;
  assign n17081 = x36 & x52 ;
  assign n17082 = ( ~n17075 & n17080 ) | ( ~n17075 & n17081 ) | ( n17080 & n17081 ) ;
  assign n17083 = n17080 & n17081 ;
  assign n17084 = ( ~n17074 & n17082 ) | ( ~n17074 & n17083 ) | ( n17082 & n17083 ) ;
  assign n17085 = ~n17079 & n17084 ;
  assign n17086 = n17078 | n17085 ;
  assign n17087 = ~n17071 & n17086 ;
  assign n17088 = n17071 & ~n17086 ;
  assign n17089 = n17087 | n17088 ;
  assign n17090 = ~n17040 & n17089 ;
  assign n17091 = n17040 & ~n17089 ;
  assign n17092 = n17090 | n17091 ;
  assign n17094 = n16995 & n17092 ;
  assign n17095 = ( ~n16733 & n16995 ) | ( ~n16733 & n17092 ) | ( n16995 & n17092 ) ;
  assign n17096 = ( ~n16738 & n17094 ) | ( ~n16738 & n17095 ) | ( n17094 & n17095 ) ;
  assign n17093 = n16733 | n16738 ;
  assign n17097 = ( ~n17092 & n17093 ) | ( ~n17092 & n17096 ) | ( n17093 & n17096 ) ;
  assign n17098 = ( ~n16995 & n17096 ) | ( ~n16995 & n17097 ) | ( n17096 & n17097 ) ;
  assign n17099 = n16952 & ~n17098 ;
  assign n17100 = ~n16952 & n17098 ;
  assign n17101 = n17099 | n17100 ;
  assign n17102 = n16742 | n16905 ;
  assign n17103 = ( n16742 & n16744 ) | ( n16742 & n17102 ) | ( n16744 & n17102 ) ;
  assign n17104 = ( n16921 & n17101 ) | ( n16921 & ~n17103 ) | ( n17101 & ~n17103 ) ;
  assign n17105 = ( ~n17101 & n17103 ) | ( ~n17101 & n17104 ) | ( n17103 & n17104 ) ;
  assign n17106 = ( ~n16921 & n17104 ) | ( ~n16921 & n17105 ) | ( n17104 & n17105 ) ;
  assign n17107 = n17101 & n17103 ;
  assign n17108 = n17101 | n17103 ;
  assign n17109 = n16920 & n17108 ;
  assign n17110 = n16914 & n17108 ;
  assign n17111 = n16912 & n17108 ;
  assign n17112 = n16690 & n17108 ;
  assign n17113 = ( n16914 & n17111 ) | ( n16914 & n17112 ) | ( n17111 & n17112 ) ;
  assign n17114 = ( n16689 & n17110 ) | ( n16689 & n17113 ) | ( n17110 & n17113 ) ;
  assign n17115 = n17110 & n17113 ;
  assign n17116 = ( n16703 & n17114 ) | ( n16703 & n17115 ) | ( n17114 & n17115 ) ;
  assign n17117 = ( n15592 & n17109 ) | ( n15592 & n17116 ) | ( n17109 & n17116 ) ;
  assign n17118 = ( n14571 & n17109 ) | ( n14571 & n17116 ) | ( n17109 & n17116 ) ;
  assign n17119 = ( n15589 & n17117 ) | ( n15589 & n17118 ) | ( n17117 & n17118 ) ;
  assign n17120 = ( n14575 & n17109 ) | ( n14575 & n17116 ) | ( n17109 & n17116 ) ;
  assign n17121 = ( n15589 & n17117 ) | ( n15589 & n17120 ) | ( n17117 & n17120 ) ;
  assign n17122 = ( n13196 & n17119 ) | ( n13196 & n17121 ) | ( n17119 & n17121 ) ;
  assign n17123 = n17107 | n17122 ;
  assign n17124 = n17016 | n17024 ;
  assign n17125 = n17068 | n17086 ;
  assign n17126 = ( n17068 & n17071 ) | ( n17068 & n17125 ) | ( n17071 & n17125 ) ;
  assign n17127 = n17124 | n17126 ;
  assign n17128 = n17124 & n17126 ;
  assign n17129 = n17127 & ~n17128 ;
  assign n17130 = ~n17010 & n17012 ;
  assign n17131 = ( n17010 & n17011 ) | ( n17010 & n17130 ) | ( n17011 & n17130 ) ;
  assign n17132 = n17063 | n17131 ;
  assign n17133 = n17063 & n17131 ;
  assign n17134 = n17132 & ~n17133 ;
  assign n17135 = x26 & x63 ;
  assign n17136 = n4555 & n6834 ;
  assign n17137 = x39 & x50 ;
  assign n17138 = x40 & x49 ;
  assign n17139 = n17137 | n17138 ;
  assign n17140 = ( n17135 & n17136 ) | ( n17135 & ~n17139 ) | ( n17136 & ~n17139 ) ;
  assign n17141 = n17135 & ~n17140 ;
  assign n17142 = ~n17136 & n17139 ;
  assign n17143 = n17135 | n17142 ;
  assign n17144 = ~n17141 & n17143 ;
  assign n17145 = n17134 & n17144 ;
  assign n17146 = n17134 & ~n17145 ;
  assign n17147 = ~n17134 & n17144 ;
  assign n17148 = n17146 | n17147 ;
  assign n17149 = n17129 | n17148 ;
  assign n17150 = n17129 & n17148 ;
  assign n17151 = n17149 & ~n17150 ;
  assign n17152 = n17038 | n17089 ;
  assign n17153 = ( n17038 & n17040 ) | ( n17038 & n17152 ) | ( n17040 & n17152 ) ;
  assign n17154 = n17151 & n17153 ;
  assign n17155 = n17151 | n17153 ;
  assign n17156 = ~n17154 & n17155 ;
  assign n17157 = n16957 | n16992 ;
  assign n17158 = ( n16957 & n16958 ) | ( n16957 & n17157 ) | ( n16958 & n17157 ) ;
  assign n17159 = n17156 & n17158 ;
  assign n17160 = n17156 | n17158 ;
  assign n17161 = ~n17159 & n17160 ;
  assign n17162 = n16733 & n17092 ;
  assign n17163 = ( n16738 & n17092 ) | ( n16738 & n17162 ) | ( n17092 & n17162 ) ;
  assign n17164 = n17093 & ~n17163 ;
  assign n17165 = ~n17093 & n17094 ;
  assign n17166 = ( n16995 & n17164 ) | ( n16995 & n17165 ) | ( n17164 & n17165 ) ;
  assign n17167 = n17161 & n17163 ;
  assign n17168 = ( n17161 & n17166 ) | ( n17161 & n17167 ) | ( n17166 & n17167 ) ;
  assign n17169 = n17163 | n17166 ;
  assign n17170 = ~n17168 & n17169 ;
  assign n17171 = n16798 | n16960 ;
  assign n17172 = ( n16960 & n16961 ) | ( n16960 & n17171 ) | ( n16961 & n17171 ) ;
  assign n17173 = n16817 | n17031 ;
  assign n17174 = ( n17031 & n17034 ) | ( n17031 & n17173 ) | ( n17034 & n17173 ) ;
  assign n17175 = n17172 | n17174 ;
  assign n17176 = n17172 & n17174 ;
  assign n17177 = n17175 & ~n17176 ;
  assign n17178 = n16967 | n16980 ;
  assign n17179 = n17177 | n17178 ;
  assign n17180 = n17177 & n17178 ;
  assign n17181 = n17179 & ~n17180 ;
  assign n17182 = n16926 | n16927 ;
  assign n17183 = ( n16926 & n16929 ) | ( n16926 & n17182 ) | ( n16929 & n17182 ) ;
  assign n17184 = n17181 | n17183 ;
  assign n17185 = n17181 & n17183 ;
  assign n17186 = n17184 & ~n17185 ;
  assign n17187 = ( n16964 & n16983 ) | ( n16964 & n16986 ) | ( n16983 & n16986 ) ;
  assign n17188 = n17186 | n17187 ;
  assign n17189 = n17186 & n17187 ;
  assign n17190 = n17188 & ~n17189 ;
  assign n17286 = n16938 | n16944 ;
  assign n17191 = n2369 & n10367 ;
  assign n17192 = x29 & x60 ;
  assign n17193 = x28 & x61 ;
  assign n17194 = n17192 | n17193 ;
  assign n17195 = ~n17191 & n17194 ;
  assign n17196 = n16975 & n17195 ;
  assign n17197 = n16975 & ~n17196 ;
  assign n17198 = ~n16975 & n17195 ;
  assign n17199 = n17197 | n17198 ;
  assign n17200 = x42 & x47 ;
  assign n17201 = x43 & x46 ;
  assign n17202 = n17200 | n17201 ;
  assign n17203 = n5407 & n6147 ;
  assign n17204 = x34 & x55 ;
  assign n17205 = ~n17203 & n17204 ;
  assign n17206 = n17202 | n17203 ;
  assign n17207 = ( n17203 & n17205 ) | ( n17203 & n17206 ) | ( n17205 & n17206 ) ;
  assign n17208 = n17202 & ~n17207 ;
  assign n17209 = ~n17202 & n17204 ;
  assign n17210 = ( n17204 & ~n17205 ) | ( n17204 & n17209 ) | ( ~n17205 & n17209 ) ;
  assign n17211 = n17208 | n17210 ;
  assign n17212 = x45 & x62 ;
  assign n17213 = x27 & n17212 ;
  assign n17214 = n6093 & n17213 ;
  assign n17215 = n6093 & ~n17213 ;
  assign n17216 = n17213 | n17215 ;
  assign n17217 = x27 & x62 ;
  assign n17218 = ( x45 & ~n17213 ) | ( x45 & n17217 ) | ( ~n17213 & n17217 ) ;
  assign n17219 = x45 & n17217 ;
  assign n17220 = ( ~n17215 & n17218 ) | ( ~n17215 & n17219 ) | ( n17218 & n17219 ) ;
  assign n17221 = ~n17216 & n17220 ;
  assign n17222 = n17214 | n17221 ;
  assign n17223 = ( n17199 & n17211 ) | ( n17199 & ~n17222 ) | ( n17211 & ~n17222 ) ;
  assign n17224 = ( n17199 & ~n17211 ) | ( n17199 & n17222 ) | ( ~n17211 & n17222 ) ;
  assign n17225 = ( ~n17199 & n17223 ) | ( ~n17199 & n17224 ) | ( n17223 & n17224 ) ;
  assign n17226 = n17048 | n17079 ;
  assign n17227 = n17048 & n17079 ;
  assign n17228 = n17226 & ~n17227 ;
  assign n17229 = n17002 | n17228 ;
  assign n17230 = n17002 & n17228 ;
  assign n17231 = n17229 & ~n17230 ;
  assign n17232 = n17225 & n17231 ;
  assign n17233 = n17225 & ~n17232 ;
  assign n17234 = n3731 & n7874 ;
  assign n17235 = n3770 & n8161 ;
  assign n17236 = n17234 | n17235 ;
  assign n17237 = n4857 & n7567 ;
  assign n17238 = x53 & n17237 ;
  assign n17239 = ( x53 & ~n17236 ) | ( x53 & n17238 ) | ( ~n17236 & n17238 ) ;
  assign n17240 = x36 & n17239 ;
  assign n17241 = n17236 | n17237 ;
  assign n17242 = ( n7946 & n11516 ) | ( n7946 & ~n17237 ) | ( n11516 & ~n17237 ) ;
  assign n17243 = n7946 & n11516 ;
  assign n17244 = ( ~n17236 & n17242 ) | ( ~n17236 & n17243 ) | ( n17242 & n17243 ) ;
  assign n17245 = ~n17241 & n17244 ;
  assign n17246 = n17240 | n17245 ;
  assign n17247 = x33 & x56 ;
  assign n17248 = x35 & x54 ;
  assign n17249 = n17247 | n17248 ;
  assign n17250 = n3129 & n8146 ;
  assign n17251 = n17249 | n17250 ;
  assign n17252 = x41 & x48 ;
  assign n17253 = ( ~n17250 & n17251 ) | ( ~n17250 & n17252 ) | ( n17251 & n17252 ) ;
  assign n17254 = ( n17250 & n17251 ) | ( n17250 & ~n17252 ) | ( n17251 & ~n17252 ) ;
  assign n17255 = ( ~n17251 & n17253 ) | ( ~n17251 & n17254 ) | ( n17253 & n17254 ) ;
  assign n17256 = n17246 & n17255 ;
  assign n17257 = n17246 & ~n17256 ;
  assign n17258 = n2546 & n9829 ;
  assign n17259 = n2965 & n9831 ;
  assign n17260 = n17258 | n17259 ;
  assign n17261 = n4062 & n9272 ;
  assign n17262 = x59 & n17261 ;
  assign n17263 = ( x59 & ~n17260 ) | ( x59 & n17262 ) | ( ~n17260 & n17262 ) ;
  assign n17264 = x30 & n17263 ;
  assign n17265 = n17260 | n17261 ;
  assign n17266 = x31 & x58 ;
  assign n17267 = x32 & x57 ;
  assign n17268 = ( ~n17261 & n17266 ) | ( ~n17261 & n17267 ) | ( n17266 & n17267 ) ;
  assign n17269 = n17266 & n17267 ;
  assign n17270 = ( ~n17260 & n17268 ) | ( ~n17260 & n17269 ) | ( n17268 & n17269 ) ;
  assign n17271 = ~n17265 & n17270 ;
  assign n17272 = n17264 | n17271 ;
  assign n17273 = ~n17246 & n17255 ;
  assign n17274 = n17272 & ~n17273 ;
  assign n17275 = ~n17257 & n17274 ;
  assign n17276 = ~n17272 & n17273 ;
  assign n17277 = ( n17257 & ~n17272 ) | ( n17257 & n17276 ) | ( ~n17272 & n17276 ) ;
  assign n17278 = n17275 | n17277 ;
  assign n17279 = n17232 & n17278 ;
  assign n17280 = ~n17231 & n17278 ;
  assign n17281 = ( ~n17233 & n17279 ) | ( ~n17233 & n17280 ) | ( n17279 & n17280 ) ;
  assign n17282 = n17232 | n17278 ;
  assign n17283 = n17231 & ~n17278 ;
  assign n17284 = ( n17233 & ~n17282 ) | ( n17233 & n17283 ) | ( ~n17282 & n17283 ) ;
  assign n17285 = n17281 | n17284 ;
  assign n17288 = ( ~n16942 & n17190 ) | ( ~n16942 & n17285 ) | ( n17190 & n17285 ) ;
  assign n17289 = ( ~n16938 & n17190 ) | ( ~n16938 & n17285 ) | ( n17190 & n17285 ) ;
  assign n17290 = ( ~n17286 & n17288 ) | ( ~n17286 & n17289 ) | ( n17288 & n17289 ) ;
  assign n17287 = ( n16938 & n16942 ) | ( n16938 & n17286 ) | ( n16942 & n17286 ) ;
  assign n17291 = ( ~n17285 & n17287 ) | ( ~n17285 & n17290 ) | ( n17287 & n17290 ) ;
  assign n17292 = ( ~n17190 & n17290 ) | ( ~n17190 & n17291 ) | ( n17290 & n17291 ) ;
  assign n17293 = n17161 & ~n17163 ;
  assign n17294 = n17292 & n17293 ;
  assign n17295 = ~n17166 & n17294 ;
  assign n17296 = ( n17170 & n17292 ) | ( n17170 & n17295 ) | ( n17292 & n17295 ) ;
  assign n17297 = n17292 | n17293 ;
  assign n17298 = ( ~n17166 & n17292 ) | ( ~n17166 & n17297 ) | ( n17292 & n17297 ) ;
  assign n17299 = n17170 | n17298 ;
  assign n17300 = ~n17296 & n17299 ;
  assign n17301 = n16950 | n17098 ;
  assign n17302 = ( n16950 & n16952 ) | ( n16950 & n17301 ) | ( n16952 & n17301 ) ;
  assign n17303 = ( n17123 & n17300 ) | ( n17123 & ~n17302 ) | ( n17300 & ~n17302 ) ;
  assign n17304 = ( ~n17300 & n17302 ) | ( ~n17300 & n17303 ) | ( n17302 & n17303 ) ;
  assign n17305 = ( ~n17123 & n17303 ) | ( ~n17123 & n17304 ) | ( n17303 & n17304 ) ;
  assign n17306 = n16942 & n17285 ;
  assign n17307 = n16938 & n17285 ;
  assign n17308 = ( n17286 & n17306 ) | ( n17286 & n17307 ) | ( n17306 & n17307 ) ;
  assign n17309 = n17287 & ~n17308 ;
  assign n17310 = n17190 & n17285 ;
  assign n17311 = ~n17287 & n17310 ;
  assign n17312 = ( n17190 & n17309 ) | ( n17190 & n17311 ) | ( n17309 & n17311 ) ;
  assign n17313 = ~n17250 & n17252 ;
  assign n17314 = ( n17250 & n17251 ) | ( n17250 & n17313 ) | ( n17251 & n17313 ) ;
  assign n17315 = n17207 | n17216 ;
  assign n17316 = n17207 & n17216 ;
  assign n17317 = n17315 & ~n17316 ;
  assign n17318 = n17314 | n17317 ;
  assign n17319 = n17314 & n17317 ;
  assign n17320 = n17318 & ~n17319 ;
  assign n17321 = n17211 & n17222 ;
  assign n17322 = n17211 & ~n17321 ;
  assign n17323 = ~n17211 & n17222 ;
  assign n17324 = n17199 & ~n17323 ;
  assign n17325 = ~n17322 & n17324 ;
  assign n17326 = ( n17199 & n17321 ) | ( n17199 & ~n17325 ) | ( n17321 & ~n17325 ) ;
  assign n17327 = n17272 & n17273 ;
  assign n17328 = ( n17257 & n17272 ) | ( n17257 & n17327 ) | ( n17272 & n17327 ) ;
  assign n17329 = n17256 | n17328 ;
  assign n17330 = n17326 | n17329 ;
  assign n17331 = n17326 & n17329 ;
  assign n17332 = n17330 & ~n17331 ;
  assign n17333 = n17320 & n17332 ;
  assign n17334 = n17320 | n17332 ;
  assign n17335 = ~n17333 & n17334 ;
  assign n17336 = ~n17232 & n17278 ;
  assign n17337 = n17231 & n17278 ;
  assign n17338 = ( n17233 & n17336 ) | ( n17233 & n17337 ) | ( n17336 & n17337 ) ;
  assign n17339 = n17232 | n17338 ;
  assign n17340 = n17335 & n17339 ;
  assign n17341 = n17335 | n17339 ;
  assign n17342 = ~n17340 & n17341 ;
  assign n17343 = n17185 | n17187 ;
  assign n17344 = ( n17185 & n17186 ) | ( n17185 & n17343 ) | ( n17186 & n17343 ) ;
  assign n17345 = n17342 | n17344 ;
  assign n17346 = n17342 & n17344 ;
  assign n17347 = n17345 & ~n17346 ;
  assign n17348 = n17308 & n17347 ;
  assign n17349 = ( n17312 & n17347 ) | ( n17312 & n17348 ) | ( n17347 & n17348 ) ;
  assign n17350 = n17308 | n17347 ;
  assign n17351 = n17312 | n17350 ;
  assign n17352 = ~n17349 & n17351 ;
  assign n17353 = n17241 | n17265 ;
  assign n17354 = n17241 & n17265 ;
  assign n17355 = n17353 & ~n17354 ;
  assign n17356 = n17135 | n17136 ;
  assign n17357 = ( n17136 & ~n17140 ) | ( n17136 & n17356 ) | ( ~n17140 & n17356 ) ;
  assign n17358 = n17355 | n17357 ;
  assign n17359 = n17355 & n17357 ;
  assign n17360 = n17358 & ~n17359 ;
  assign n17361 = n17176 | n17178 ;
  assign n17362 = ( n17176 & n17177 ) | ( n17176 & n17361 ) | ( n17177 & n17361 ) ;
  assign n17363 = n17360 | n17362 ;
  assign n17364 = n17360 & n17362 ;
  assign n17365 = n17363 & ~n17364 ;
  assign n17366 = n3129 & n12860 ;
  assign n17367 = n3483 & n10013 ;
  assign n17368 = n17366 | n17367 ;
  assign n17369 = n4530 & n8903 ;
  assign n17370 = x55 & n17369 ;
  assign n17371 = ( x55 & ~n17368 ) | ( x55 & n17370 ) | ( ~n17368 & n17370 ) ;
  assign n17372 = x35 & n17371 ;
  assign n17373 = n17368 | n17369 ;
  assign n17374 = x33 & x57 ;
  assign n17375 = x34 & x56 ;
  assign n17376 = ( ~n17369 & n17374 ) | ( ~n17369 & n17375 ) | ( n17374 & n17375 ) ;
  assign n17377 = n17374 & n17375 ;
  assign n17378 = ( ~n17368 & n17376 ) | ( ~n17368 & n17377 ) | ( n17376 & n17377 ) ;
  assign n17379 = ~n17373 & n17378 ;
  assign n17380 = n17372 | n17379 ;
  assign n17381 = n3731 & n11935 ;
  assign n17382 = n3770 & n8355 ;
  assign n17383 = n17381 | n17382 ;
  assign n17384 = n4857 & n8161 ;
  assign n17385 = x54 & n17384 ;
  assign n17386 = ( x54 & ~n17383 ) | ( x54 & n17385 ) | ( ~n17383 & n17385 ) ;
  assign n17387 = x36 & n17386 ;
  assign n17388 = n17383 | n17384 ;
  assign n17389 = x38 & x52 ;
  assign n17390 = ( n8163 & ~n17384 ) | ( n8163 & n17389 ) | ( ~n17384 & n17389 ) ;
  assign n17391 = n8163 & n17389 ;
  assign n17392 = ( ~n17383 & n17390 ) | ( ~n17383 & n17391 ) | ( n17390 & n17391 ) ;
  assign n17393 = ~n17388 & n17392 ;
  assign n17394 = n17387 | n17393 ;
  assign n17395 = n17380 & n17394 ;
  assign n17396 = n17380 & ~n17395 ;
  assign n17397 = n17394 & ~n17395 ;
  assign n17398 = n17396 | n17397 ;
  assign n17399 = n4969 & n9421 ;
  assign n17400 = n5407 & n6762 ;
  assign n17401 = n17399 | n17400 ;
  assign n17402 = n5658 & n6147 ;
  assign n17403 = x48 & n17402 ;
  assign n17404 = ( x48 & ~n17401 ) | ( x48 & n17403 ) | ( ~n17401 & n17403 ) ;
  assign n17405 = x42 & n17404 ;
  assign n17406 = n8407 | n8772 ;
  assign n17407 = ~n17402 & n17406 ;
  assign n17408 = ~n17401 & n17407 ;
  assign n17409 = n17405 | n17408 ;
  assign n17410 = ~n17398 & n17409 ;
  assign n17411 = n17398 & ~n17409 ;
  assign n17412 = n17410 | n17411 ;
  assign n17413 = n17365 & n17412 ;
  assign n17414 = n17365 | n17412 ;
  assign n17415 = ~n17413 & n17414 ;
  assign n17416 = ~n17154 & n17415 ;
  assign n17417 = ~n17159 & n17416 ;
  assign n17418 = n17154 & n17415 ;
  assign n17419 = ( n17159 & n17415 ) | ( n17159 & n17418 ) | ( n17415 & n17418 ) ;
  assign n17420 = ( n17154 & n17159 ) | ( n17154 & ~n17419 ) | ( n17159 & ~n17419 ) ;
  assign n17421 = n17417 | n17420 ;
  assign n17433 = n17191 | n17195 ;
  assign n17434 = ( n16975 & n17191 ) | ( n16975 & n17433 ) | ( n17191 & n17433 ) ;
  assign n17422 = n4062 & n9831 ;
  assign n17423 = n2546 & n10975 ;
  assign n17424 = n2965 & n10370 ;
  assign n17425 = n17423 | n17424 ;
  assign n17426 = ~n17422 & n17425 ;
  assign n17427 = x31 & x59 ;
  assign n17428 = n15870 | n17427 ;
  assign n17429 = ~n17422 & n17428 ;
  assign n17430 = x30 & x60 ;
  assign n17431 = n17429 | n17430 ;
  assign n17432 = ~n17426 & n17431 ;
  assign n17435 = n17432 & n17434 ;
  assign n17436 = n17434 & ~n17435 ;
  assign n17437 = n2372 & n10561 ;
  assign n17438 = n2075 & n10856 ;
  assign n17439 = n17437 | n17438 ;
  assign n17440 = n2369 & n10684 ;
  assign n17441 = x63 & n17440 ;
  assign n17442 = ( x63 & ~n17439 ) | ( x63 & n17441 ) | ( ~n17439 & n17441 ) ;
  assign n17443 = x27 & n17442 ;
  assign n17444 = n17439 | n17440 ;
  assign n17445 = x28 & x62 ;
  assign n17446 = x29 & x61 ;
  assign n17447 = ( ~n17440 & n17445 ) | ( ~n17440 & n17446 ) | ( n17445 & n17446 ) ;
  assign n17448 = n17445 & n17446 ;
  assign n17449 = ( ~n17439 & n17447 ) | ( ~n17439 & n17448 ) | ( n17447 & n17448 ) ;
  assign n17450 = ~n17444 & n17449 ;
  assign n17451 = n17443 | n17450 ;
  assign n17452 = n17432 & ~n17434 ;
  assign n17453 = n17451 | n17452 ;
  assign n17454 = n17436 | n17453 ;
  assign n17455 = n17451 & n17452 ;
  assign n17456 = ( n17436 & n17451 ) | ( n17436 & n17455 ) | ( n17451 & n17455 ) ;
  assign n17457 = n17454 & ~n17456 ;
  assign n17472 = n17002 | n17227 ;
  assign n17473 = ( n17227 & n17228 ) | ( n17227 & n17472 ) | ( n17228 & n17472 ) ;
  assign n17458 = n4350 & n10866 ;
  assign n17459 = n4555 & n7112 ;
  assign n17460 = n17458 | n17459 ;
  assign n17461 = n5813 & n6834 ;
  assign n17462 = n8433 & n17461 ;
  assign n17463 = ( n8433 & ~n17460 ) | ( n8433 & n17462 ) | ( ~n17460 & n17462 ) ;
  assign n17464 = n17460 | n17461 ;
  assign n17465 = x41 & x49 ;
  assign n17466 = x40 & x50 ;
  assign n17467 = ( ~n17461 & n17465 ) | ( ~n17461 & n17466 ) | ( n17465 & n17466 ) ;
  assign n17468 = n17465 & n17466 ;
  assign n17469 = ( ~n17460 & n17467 ) | ( ~n17460 & n17468 ) | ( n17467 & n17468 ) ;
  assign n17470 = ~n17464 & n17469 ;
  assign n17471 = n17463 | n17470 ;
  assign n17474 = n17471 & n17473 ;
  assign n17475 = n17473 & ~n17474 ;
  assign n17477 = n17133 | n17144 ;
  assign n17478 = ( n17133 & n17134 ) | ( n17133 & n17477 ) | ( n17134 & n17477 ) ;
  assign n17476 = n17471 & ~n17473 ;
  assign n17479 = n17476 & n17478 ;
  assign n17480 = ( n17475 & n17478 ) | ( n17475 & n17479 ) | ( n17478 & n17479 ) ;
  assign n17481 = n17476 | n17478 ;
  assign n17482 = n17475 | n17481 ;
  assign n17483 = ~n17480 & n17482 ;
  assign n17484 = n17457 & n17483 ;
  assign n17485 = n17483 & ~n17484 ;
  assign n17486 = ( n17457 & ~n17484 ) | ( n17457 & n17485 ) | ( ~n17484 & n17485 ) ;
  assign n17487 = n17128 | n17148 ;
  assign n17488 = ( n17128 & n17129 ) | ( n17128 & n17487 ) | ( n17129 & n17487 ) ;
  assign n17489 = n17486 & n17488 ;
  assign n17490 = n17486 & ~n17489 ;
  assign n17491 = ~n17486 & n17488 ;
  assign n17492 = n17490 | n17491 ;
  assign n17493 = n17417 | n17492 ;
  assign n17494 = n17420 | n17493 ;
  assign n17495 = ~n17492 & n17494 ;
  assign n17496 = ( ~n17421 & n17494 ) | ( ~n17421 & n17495 ) | ( n17494 & n17495 ) ;
  assign n17497 = n17352 | n17496 ;
  assign n17498 = n17352 & n17496 ;
  assign n17499 = n17497 & ~n17498 ;
  assign n17500 = n17168 | n17295 ;
  assign n17501 = n17168 | n17292 ;
  assign n17502 = ( n17170 & n17500 ) | ( n17170 & n17501 ) | ( n17500 & n17501 ) ;
  assign n17503 = n17499 | n17502 ;
  assign n17504 = n17499 & n17502 ;
  assign n17505 = n17503 & ~n17504 ;
  assign n17506 = n17300 & n17302 ;
  assign n17507 = n17300 | n17302 ;
  assign n17508 = n17107 & n17507 ;
  assign n17509 = n17506 | n17508 ;
  assign n17510 = n17506 | n17507 ;
  assign n17511 = ( n17122 & n17509 ) | ( n17122 & n17510 ) | ( n17509 & n17510 ) ;
  assign n17512 = n17505 | n17511 ;
  assign n17513 = n17503 & n17510 ;
  assign n17514 = n17503 & n17506 ;
  assign n17515 = ( n17503 & n17508 ) | ( n17503 & n17514 ) | ( n17508 & n17514 ) ;
  assign n17516 = ( n17122 & n17513 ) | ( n17122 & n17515 ) | ( n17513 & n17515 ) ;
  assign n17517 = ~n17504 & n17516 ;
  assign n17518 = n17512 & ~n17517 ;
  assign n17519 = n17388 | n17444 ;
  assign n17520 = n17388 & n17444 ;
  assign n17521 = n17519 & ~n17520 ;
  assign n17522 = n17422 | n17425 ;
  assign n17523 = n17521 | n17522 ;
  assign n17524 = n17521 & n17522 ;
  assign n17525 = n17523 & ~n17524 ;
  assign n17526 = n17474 & n17525 ;
  assign n17527 = ( n17480 & n17525 ) | ( n17480 & n17526 ) | ( n17525 & n17526 ) ;
  assign n17528 = n17474 | n17525 ;
  assign n17529 = n17480 | n17528 ;
  assign n17530 = ~n17527 & n17529 ;
  assign n17531 = x43 & x48 ;
  assign n17532 = x44 & x47 ;
  assign n17533 = n17531 | n17532 ;
  assign n17534 = n5658 & n6762 ;
  assign n17535 = x35 & x56 ;
  assign n17536 = ~n17534 & n17535 ;
  assign n17537 = n17533 | n17534 ;
  assign n17538 = ( n17534 & n17536 ) | ( n17534 & n17537 ) | ( n17536 & n17537 ) ;
  assign n17539 = n17533 & ~n17538 ;
  assign n17540 = ( ~n17533 & n17534 ) | ( ~n17533 & n17535 ) | ( n17534 & n17535 ) ;
  assign n17541 = n17535 & n17540 ;
  assign n17542 = n17539 | n17541 ;
  assign n17543 = x40 & x51 ;
  assign n17544 = x41 & x50 ;
  assign n17545 = n17543 | n17544 ;
  assign n17546 = n5813 & n7112 ;
  assign n17547 = n17545 | n17546 ;
  assign n17548 = x28 & x63 ;
  assign n17549 = ( ~n17546 & n17547 ) | ( ~n17546 & n17548 ) | ( n17547 & n17548 ) ;
  assign n17550 = ( n17546 & n17547 ) | ( n17546 & ~n17548 ) | ( n17547 & ~n17548 ) ;
  assign n17551 = ( ~n17547 & n17549 ) | ( ~n17547 & n17550 ) | ( n17549 & n17550 ) ;
  assign n17552 = n17542 & n17551 ;
  assign n17553 = n17542 & ~n17552 ;
  assign n17554 = x46 & x62 ;
  assign n17555 = x29 & n17554 ;
  assign n17556 = n5975 & n17555 ;
  assign n17557 = n5975 & ~n17555 ;
  assign n17558 = n17555 | n17557 ;
  assign n17559 = x29 & x62 ;
  assign n17560 = ( x46 & ~n17555 ) | ( x46 & n17559 ) | ( ~n17555 & n17559 ) ;
  assign n17561 = x46 & n17559 ;
  assign n17562 = ( ~n17557 & n17560 ) | ( ~n17557 & n17561 ) | ( n17560 & n17561 ) ;
  assign n17563 = ~n17558 & n17562 ;
  assign n17564 = n17556 | n17563 ;
  assign n17565 = ~n17542 & n17551 ;
  assign n17566 = n17564 & ~n17565 ;
  assign n17567 = ~n17553 & n17566 ;
  assign n17568 = ~n17564 & n17565 ;
  assign n17569 = ( n17553 & ~n17564 ) | ( n17553 & n17568 ) | ( ~n17564 & n17568 ) ;
  assign n17570 = n17567 | n17569 ;
  assign n17571 = n17530 | n17570 ;
  assign n17572 = n17530 & n17570 ;
  assign n17573 = n17571 & ~n17572 ;
  assign n17574 = n17340 | n17344 ;
  assign n17575 = ( n17340 & n17342 ) | ( n17340 & n17574 ) | ( n17342 & n17574 ) ;
  assign n17576 = n17573 & n17575 ;
  assign n17577 = n17573 | n17575 ;
  assign n17578 = ~n17576 & n17577 ;
  assign n17637 = n17320 | n17331 ;
  assign n17638 = ( n17331 & n17332 ) | ( n17331 & n17637 ) | ( n17332 & n17637 ) ;
  assign n17590 = n17314 | n17316 ;
  assign n17591 = ( n17316 & n17317 ) | ( n17316 & n17590 ) | ( n17317 & n17590 ) ;
  assign n17579 = x34 & x57 ;
  assign n17580 = x36 & x55 ;
  assign n17581 = n17579 | n17580 ;
  assign n17582 = n4914 & n12860 ;
  assign n17583 = n8722 & ~n17582 ;
  assign n17584 = n17581 | n17582 ;
  assign n17585 = ( n17582 & n17583 ) | ( n17582 & n17584 ) | ( n17583 & n17584 ) ;
  assign n17586 = n17581 & ~n17585 ;
  assign n17587 = n8722 & ~n17581 ;
  assign n17588 = ( n8722 & ~n17583 ) | ( n8722 & n17587 ) | ( ~n17583 & n17587 ) ;
  assign n17589 = n17586 | n17588 ;
  assign n17592 = n17589 & n17591 ;
  assign n17593 = n17591 & ~n17592 ;
  assign n17595 = n17354 | n17357 ;
  assign n17596 = ( n17354 & n17355 ) | ( n17354 & n17595 ) | ( n17355 & n17595 ) ;
  assign n17594 = n17589 & ~n17591 ;
  assign n17597 = n17594 & n17596 ;
  assign n17598 = ( n17593 & n17596 ) | ( n17593 & n17597 ) | ( n17596 & n17597 ) ;
  assign n17599 = n17594 | n17596 ;
  assign n17600 = n17593 | n17599 ;
  assign n17601 = ~n17598 & n17600 ;
  assign n17602 = n2683 & n10975 ;
  assign n17603 = n4062 & n10370 ;
  assign n17604 = n17602 | n17603 ;
  assign n17605 = n3321 & n9831 ;
  assign n17606 = x60 & n17605 ;
  assign n17607 = ( x60 & ~n17604 ) | ( x60 & n17606 ) | ( ~n17604 & n17606 ) ;
  assign n17608 = x31 & n17607 ;
  assign n17609 = n17604 | n17605 ;
  assign n17610 = x33 & x58 ;
  assign n17611 = ( n9069 & ~n17605 ) | ( n9069 & n17610 ) | ( ~n17605 & n17610 ) ;
  assign n17612 = n9069 & n17610 ;
  assign n17613 = ( ~n17604 & n17611 ) | ( ~n17604 & n17612 ) | ( n17611 & n17612 ) ;
  assign n17614 = ~n17609 & n17613 ;
  assign n17615 = n17608 | n17614 ;
  assign n17616 = n5798 & n11935 ;
  assign n17617 = n4857 & n8355 ;
  assign n17618 = n17616 | n17617 ;
  assign n17619 = n5392 & n8161 ;
  assign n17620 = x37 & n17619 ;
  assign n17621 = ( x37 & ~n17618 ) | ( x37 & n17620 ) | ( ~n17618 & n17620 ) ;
  assign n17622 = x54 & n17621 ;
  assign n17623 = n17618 | n17619 ;
  assign n17624 = x38 & x53 ;
  assign n17625 = x39 & x52 ;
  assign n17626 = ( ~n17619 & n17624 ) | ( ~n17619 & n17625 ) | ( n17624 & n17625 ) ;
  assign n17627 = n17624 & n17625 ;
  assign n17628 = ( ~n17618 & n17626 ) | ( ~n17618 & n17627 ) | ( n17626 & n17627 ) ;
  assign n17629 = ~n17623 & n17628 ;
  assign n17630 = n17622 | n17629 ;
  assign n17631 = n17464 & n17630 ;
  assign n17632 = n17464 | n17630 ;
  assign n17633 = ~n17631 & n17632 ;
  assign n17634 = n17615 & ~n17633 ;
  assign n17635 = ~n17615 & n17633 ;
  assign n17636 = n17634 | n17635 ;
  assign n17639 = ( n17601 & ~n17636 ) | ( n17601 & n17638 ) | ( ~n17636 & n17638 ) ;
  assign n17640 = ( ~n17601 & n17636 ) | ( ~n17601 & n17638 ) | ( n17636 & n17638 ) ;
  assign n17641 = ( ~n17638 & n17639 ) | ( ~n17638 & n17640 ) | ( n17639 & n17640 ) ;
  assign n17642 = n17578 & ~n17641 ;
  assign n17643 = n17578 | n17641 ;
  assign n17644 = ( ~n17578 & n17642 ) | ( ~n17578 & n17643 ) | ( n17642 & n17643 ) ;
  assign n17645 = x30 & x61 ;
  assign n17646 = n17402 & n17645 ;
  assign n17647 = ( n17401 & n17645 ) | ( n17401 & n17646 ) | ( n17645 & n17646 ) ;
  assign n17648 = n17402 | n17645 ;
  assign n17649 = n17401 | n17648 ;
  assign n17650 = ~n17647 & n17649 ;
  assign n17651 = n17373 | n17650 ;
  assign n17652 = n17373 & n17650 ;
  assign n17653 = n17651 & ~n17652 ;
  assign n17654 = n17435 | n17456 ;
  assign n17655 = n17395 | n17409 ;
  assign n17656 = ( n17395 & n17398 ) | ( n17395 & n17655 ) | ( n17398 & n17655 ) ;
  assign n17657 = n17654 | n17656 ;
  assign n17658 = n17654 & n17656 ;
  assign n17659 = n17657 & ~n17658 ;
  assign n17660 = n17653 & n17659 ;
  assign n17661 = n17653 | n17659 ;
  assign n17662 = ~n17660 & n17661 ;
  assign n17663 = n17364 | n17412 ;
  assign n17664 = ( n17364 & n17365 ) | ( n17364 & n17663 ) | ( n17365 & n17663 ) ;
  assign n17665 = n17662 & n17664 ;
  assign n17666 = ~n17662 & n17664 ;
  assign n17667 = ( n17662 & ~n17665 ) | ( n17662 & n17666 ) | ( ~n17665 & n17666 ) ;
  assign n17668 = n17484 | n17488 ;
  assign n17669 = ( n17484 & n17486 ) | ( n17484 & n17668 ) | ( n17486 & n17668 ) ;
  assign n17670 = n17667 & n17669 ;
  assign n17671 = n17667 & ~n17670 ;
  assign n17672 = ~n17667 & n17669 ;
  assign n17673 = n17671 | n17672 ;
  assign n17674 = n17419 | n17492 ;
  assign n17675 = ( n17419 & n17421 ) | ( n17419 & n17674 ) | ( n17421 & n17674 ) ;
  assign n17676 = ( n17644 & n17673 ) | ( n17644 & ~n17675 ) | ( n17673 & ~n17675 ) ;
  assign n17677 = ( ~n17673 & n17675 ) | ( ~n17673 & n17676 ) | ( n17675 & n17676 ) ;
  assign n17678 = ( ~n17644 & n17676 ) | ( ~n17644 & n17677 ) | ( n17676 & n17677 ) ;
  assign n17679 = n17349 | n17352 ;
  assign n17680 = ( n17349 & n17496 ) | ( n17349 & n17679 ) | ( n17496 & n17679 ) ;
  assign n17681 = n17678 & n17680 ;
  assign n17682 = n17678 | n17680 ;
  assign n17683 = ~n17681 & n17682 ;
  assign n17684 = n17504 | n17515 ;
  assign n17685 = n17503 | n17504 ;
  assign n17686 = ( n17504 & n17510 ) | ( n17504 & n17685 ) | ( n17510 & n17685 ) ;
  assign n17687 = ( n17122 & n17684 ) | ( n17122 & n17686 ) | ( n17684 & n17686 ) ;
  assign n17688 = ~n17683 & n17687 ;
  assign n17689 = n17683 & ~n17687 ;
  assign n17690 = n17688 | n17689 ;
  assign n17691 = n3483 & n9272 ;
  assign n17692 = x42 & x50 ;
  assign n17693 = x34 & x58 ;
  assign n17694 = n17692 & n17693 ;
  assign n17695 = n17691 | n17694 ;
  assign n17696 = x35 & x57 ;
  assign n17697 = n17692 & n17696 ;
  assign n17698 = n17695 | n17697 ;
  assign n17700 = n17693 & n17697 ;
  assign n17701 = ( n17693 & ~n17695 ) | ( n17693 & n17700 ) | ( ~n17695 & n17700 ) ;
  assign n17699 = n17692 | n17696 ;
  assign n17702 = n17699 | n17701 ;
  assign n17703 = ( ~n17698 & n17701 ) | ( ~n17698 & n17702 ) | ( n17701 & n17702 ) ;
  assign n17704 = n5104 & n6757 ;
  assign n17705 = n5658 & n6759 ;
  assign n17706 = n17704 | n17705 ;
  assign n17707 = n6093 & n6762 ;
  assign n17708 = x49 & n17707 ;
  assign n17709 = ( x49 & ~n17706 ) | ( x49 & n17708 ) | ( ~n17706 & n17708 ) ;
  assign n17710 = x43 & n17709 ;
  assign n17711 = n17706 | n17707 ;
  assign n17712 = x44 & x48 ;
  assign n17713 = ( n5610 & ~n17707 ) | ( n5610 & n17712 ) | ( ~n17707 & n17712 ) ;
  assign n17714 = n5610 & n17712 ;
  assign n17715 = ( ~n17706 & n17713 ) | ( ~n17706 & n17714 ) | ( n17713 & n17714 ) ;
  assign n17716 = ~n17711 & n17715 ;
  assign n17717 = n17710 | n17716 ;
  assign n17718 = n17703 & n17717 ;
  assign n17719 = n17703 & ~n17718 ;
  assign n17720 = n17717 & ~n17718 ;
  assign n17721 = n17719 | n17720 ;
  assign n17722 = x33 & x59 ;
  assign n17723 = n15182 | n17722 ;
  assign n17724 = x36 & x56 ;
  assign n17725 = ( n15182 & n17722 ) | ( n15182 & n17724 ) | ( n17722 & n17724 ) ;
  assign n17726 = n17723 & ~n17725 ;
  assign n17727 = n15182 & n17722 ;
  assign n17728 = n17724 & ~n17727 ;
  assign n17729 = ~n17723 & n17724 ;
  assign n17730 = ( n17724 & ~n17728 ) | ( n17724 & n17729 ) | ( ~n17728 & n17729 ) ;
  assign n17731 = n17726 | n17730 ;
  assign n17732 = ~n17721 & n17731 ;
  assign n17733 = n17721 & ~n17731 ;
  assign n17734 = n17732 | n17733 ;
  assign n17759 = n17373 | n17647 ;
  assign n17760 = ( n17647 & n17650 ) | ( n17647 & n17759 ) | ( n17650 & n17759 ) ;
  assign n17735 = n2965 & n10684 ;
  assign n17736 = x31 & x61 ;
  assign n17737 = x30 & x62 ;
  assign n17738 = n17736 | n17737 ;
  assign n17739 = ~n17735 & n17738 ;
  assign n17740 = n17558 & n17739 ;
  assign n17741 = n17558 & ~n17740 ;
  assign n17742 = ~n17558 & n17739 ;
  assign n17743 = n17741 | n17742 ;
  assign n17744 = n4350 & n7874 ;
  assign n17745 = n4555 & n8161 ;
  assign n17746 = n17744 | n17745 ;
  assign n17747 = n5813 & n7567 ;
  assign n17748 = x53 & n17747 ;
  assign n17749 = ( x53 & ~n17746 ) | ( x53 & n17748 ) | ( ~n17746 & n17748 ) ;
  assign n17750 = x39 & n17749 ;
  assign n17751 = n17746 | n17747 ;
  assign n17752 = x40 & x52 ;
  assign n17753 = x41 & x51 ;
  assign n17754 = ( ~n17747 & n17752 ) | ( ~n17747 & n17753 ) | ( n17752 & n17753 ) ;
  assign n17755 = n17752 & n17753 ;
  assign n17756 = ( ~n17746 & n17754 ) | ( ~n17746 & n17755 ) | ( n17754 & n17755 ) ;
  assign n17757 = ~n17751 & n17756 ;
  assign n17758 = n17750 | n17757 ;
  assign n17761 = ( n17743 & ~n17758 ) | ( n17743 & n17760 ) | ( ~n17758 & n17760 ) ;
  assign n17762 = ( ~n17743 & n17758 ) | ( ~n17743 & n17761 ) | ( n17758 & n17761 ) ;
  assign n17763 = ( ~n17760 & n17761 ) | ( ~n17760 & n17762 ) | ( n17761 & n17762 ) ;
  assign n17764 = n17734 | n17763 ;
  assign n17765 = n17734 & n17763 ;
  assign n17766 = n17764 & ~n17765 ;
  assign n17767 = n17653 | n17654 ;
  assign n17768 = ( n17653 & n17656 ) | ( n17653 & n17767 ) | ( n17656 & n17767 ) ;
  assign n17769 = ( n17658 & n17659 ) | ( n17658 & n17768 ) | ( n17659 & n17768 ) ;
  assign n17770 = n17766 & n17769 ;
  assign n17771 = n17766 | n17769 ;
  assign n17772 = ~n17770 & n17771 ;
  assign n17773 = n17636 & n17638 ;
  assign n17774 = n17638 & ~n17773 ;
  assign n17775 = n17601 & n17636 ;
  assign n17776 = ~n17638 & n17775 ;
  assign n17777 = n17773 | n17776 ;
  assign n17778 = n17601 | n17636 ;
  assign n17779 = ( n17601 & n17638 ) | ( n17601 & n17778 ) | ( n17638 & n17778 ) ;
  assign n17780 = ( n17774 & n17777 ) | ( n17774 & n17779 ) | ( n17777 & n17779 ) ;
  assign n17781 = n17772 & n17780 ;
  assign n17782 = n17772 | n17780 ;
  assign n17783 = ~n17781 & n17782 ;
  assign n17784 = n17665 | n17669 ;
  assign n17785 = ( n17665 & n17667 ) | ( n17665 & n17784 ) | ( n17667 & n17784 ) ;
  assign n17786 = n17783 & n17785 ;
  assign n17787 = n17783 | n17785 ;
  assign n17788 = ~n17786 & n17787 ;
  assign n17789 = n17615 | n17631 ;
  assign n17790 = ( n17631 & n17633 ) | ( n17631 & n17789 ) | ( n17633 & n17789 ) ;
  assign n17791 = n17520 | n17522 ;
  assign n17792 = ( n17520 & n17521 ) | ( n17520 & n17791 ) | ( n17521 & n17791 ) ;
  assign n17793 = n17790 & n17792 ;
  assign n17794 = n17790 | n17792 ;
  assign n17795 = ~n17793 & n17794 ;
  assign n17796 = n17564 & n17565 ;
  assign n17797 = ( n17553 & n17564 ) | ( n17553 & n17796 ) | ( n17564 & n17796 ) ;
  assign n17798 = n17552 | n17797 ;
  assign n17799 = n17795 | n17798 ;
  assign n17800 = n17795 & n17798 ;
  assign n17801 = n17799 & ~n17800 ;
  assign n17802 = n17592 | n17598 ;
  assign n17803 = ~n17546 & n17548 ;
  assign n17804 = ( n17546 & n17547 ) | ( n17546 & n17803 ) | ( n17547 & n17803 ) ;
  assign n17805 = n17609 | n17623 ;
  assign n17806 = n17609 & n17623 ;
  assign n17807 = n17805 & ~n17806 ;
  assign n17808 = n17804 | n17807 ;
  assign n17809 = n17804 & n17807 ;
  assign n17810 = n17808 & ~n17809 ;
  assign n17811 = n17538 | n17585 ;
  assign n17812 = n17538 & n17585 ;
  assign n17813 = n17811 & ~n17812 ;
  assign n17814 = x37 & x55 ;
  assign n17815 = x38 & x54 ;
  assign n17816 = n17814 | n17815 ;
  assign n17817 = n4857 & n8357 ;
  assign n17818 = n17816 & ~n17817 ;
  assign n17819 = x32 & x60 ;
  assign n17820 = n17817 | n17819 ;
  assign n17821 = ( n17817 & n17818 ) | ( n17817 & n17820 ) | ( n17818 & n17820 ) ;
  assign n17822 = n17816 & ~n17821 ;
  assign n17823 = ~n17818 & n17819 ;
  assign n17824 = n17822 | n17823 ;
  assign n17825 = n17813 & n17824 ;
  assign n17826 = n17813 & ~n17825 ;
  assign n17827 = n17824 & ~n17825 ;
  assign n17828 = n17826 | n17827 ;
  assign n17829 = n17810 | n17828 ;
  assign n17830 = n17810 & n17828 ;
  assign n17831 = n17829 & ~n17830 ;
  assign n17832 = n17802 & n17831 ;
  assign n17833 = n17802 | n17831 ;
  assign n17834 = ~n17832 & n17833 ;
  assign n17835 = n17527 | n17570 ;
  assign n17836 = ( n17527 & n17530 ) | ( n17527 & n17835 ) | ( n17530 & n17835 ) ;
  assign n17837 = n17834 & n17836 ;
  assign n17838 = n17834 | n17836 ;
  assign n17839 = ~n17837 & n17838 ;
  assign n17840 = n17801 & n17839 ;
  assign n17841 = n17801 | n17839 ;
  assign n17842 = ~n17840 & n17841 ;
  assign n17843 = n17573 | n17641 ;
  assign n17844 = ( n17575 & n17641 ) | ( n17575 & n17843 ) | ( n17641 & n17843 ) ;
  assign n17845 = n17842 & n17844 ;
  assign n17846 = n17576 & n17842 ;
  assign n17847 = ( n17578 & n17845 ) | ( n17578 & n17846 ) | ( n17845 & n17846 ) ;
  assign n17848 = n17842 | n17844 ;
  assign n17849 = n17576 | n17842 ;
  assign n17850 = ( n17578 & n17848 ) | ( n17578 & n17849 ) | ( n17848 & n17849 ) ;
  assign n17851 = ~n17847 & n17850 ;
  assign n17852 = n17788 & n17851 ;
  assign n17853 = n17788 | n17851 ;
  assign n17854 = ~n17852 & n17853 ;
  assign n17855 = n17673 & n17674 ;
  assign n17856 = n17419 & n17673 ;
  assign n17857 = ( n17421 & n17855 ) | ( n17421 & n17856 ) | ( n17855 & n17856 ) ;
  assign n17858 = n17675 & ~n17857 ;
  assign n17859 = n17673 & ~n17674 ;
  assign n17860 = ~n17419 & n17673 ;
  assign n17861 = ( ~n17421 & n17859 ) | ( ~n17421 & n17860 ) | ( n17859 & n17860 ) ;
  assign n17862 = n17644 & ~n17861 ;
  assign n17863 = ~n17858 & n17862 ;
  assign n17864 = ( n17644 & n17857 ) | ( n17644 & ~n17863 ) | ( n17857 & ~n17863 ) ;
  assign n17865 = n17854 | n17864 ;
  assign n17866 = n17854 & n17864 ;
  assign n17867 = n17865 & ~n17866 ;
  assign n17868 = n17681 | n17682 ;
  assign n17869 = ( n17681 & n17686 ) | ( n17681 & n17868 ) | ( n17686 & n17868 ) ;
  assign n17870 = ( n17504 & n17678 ) | ( n17504 & n17680 ) | ( n17678 & n17680 ) ;
  assign n17871 = ( n17515 & n17682 ) | ( n17515 & n17870 ) | ( n17682 & n17870 ) ;
  assign n17872 = ( n17122 & n17869 ) | ( n17122 & n17871 ) | ( n17869 & n17871 ) ;
  assign n17873 = n17867 | n17872 ;
  assign n17874 = n17865 & n17871 ;
  assign n17875 = n17865 & n17868 ;
  assign n17876 = n17681 & n17865 ;
  assign n17877 = ( n17686 & n17875 ) | ( n17686 & n17876 ) | ( n17875 & n17876 ) ;
  assign n17878 = ( n17122 & n17874 ) | ( n17122 & n17877 ) | ( n17874 & n17877 ) ;
  assign n17879 = ~n17866 & n17878 ;
  assign n17880 = n17873 & ~n17879 ;
  assign n17881 = n17866 | n17877 ;
  assign n17882 = n17865 | n17866 ;
  assign n17883 = ( n17866 & n17871 ) | ( n17866 & n17882 ) | ( n17871 & n17882 ) ;
  assign n17884 = ( n17122 & n17881 ) | ( n17122 & n17883 ) | ( n17881 & n17883 ) ;
  assign n17885 = n17812 | n17825 ;
  assign n17886 = n17804 | n17806 ;
  assign n17887 = ( n17806 & n17807 ) | ( n17806 & n17886 ) | ( n17807 & n17886 ) ;
  assign n17888 = n17885 | n17887 ;
  assign n17889 = n17885 & n17887 ;
  assign n17890 = n17888 & ~n17889 ;
  assign n17891 = n17718 | n17731 ;
  assign n17892 = ( n17718 & n17721 ) | ( n17718 & n17891 ) | ( n17721 & n17891 ) ;
  assign n17893 = n17890 | n17892 ;
  assign n17894 = n17890 & n17892 ;
  assign n17895 = n17893 & ~n17894 ;
  assign n17896 = n17830 | n17832 ;
  assign n17897 = n17895 & n17896 ;
  assign n17898 = n17895 | n17896 ;
  assign n17899 = ~n17897 & n17898 ;
  assign n17900 = n17698 | n17711 ;
  assign n17901 = n17698 & n17711 ;
  assign n17902 = n17900 & ~n17901 ;
  assign n17903 = n17751 | n17902 ;
  assign n17904 = n17751 & n17902 ;
  assign n17905 = n17903 & ~n17904 ;
  assign n17906 = n17725 | n17821 ;
  assign n17907 = n17725 & n17821 ;
  assign n17908 = n17906 & ~n17907 ;
  assign n17909 = n17735 | n17739 ;
  assign n17910 = ( n17558 & n17735 ) | ( n17558 & n17909 ) | ( n17735 & n17909 ) ;
  assign n17911 = n17908 | n17910 ;
  assign n17912 = n17908 & n17910 ;
  assign n17913 = n17911 & ~n17912 ;
  assign n17914 = n17905 & n17913 ;
  assign n17915 = n17905 | n17913 ;
  assign n17916 = ~n17914 & n17915 ;
  assign n17917 = n17743 & n17758 ;
  assign n17918 = n17743 & ~n17917 ;
  assign n17919 = n17758 & n17760 ;
  assign n17920 = ~n17743 & n17919 ;
  assign n17921 = n17917 | n17920 ;
  assign n17922 = n17758 | n17760 ;
  assign n17923 = ( n17743 & n17760 ) | ( n17743 & n17922 ) | ( n17760 & n17922 ) ;
  assign n17924 = ( n17918 & n17921 ) | ( n17918 & n17923 ) | ( n17921 & n17923 ) ;
  assign n17925 = n17916 & n17924 ;
  assign n17926 = n17916 | n17924 ;
  assign n17927 = ~n17925 & n17926 ;
  assign n17928 = n17899 & n17927 ;
  assign n17929 = n17899 | n17927 ;
  assign n17930 = ~n17928 & n17929 ;
  assign n17931 = n17781 | n17785 ;
  assign n17932 = ( n17781 & n17783 ) | ( n17781 & n17931 ) | ( n17783 & n17931 ) ;
  assign n17933 = n17930 | n17932 ;
  assign n17934 = n6638 & n10718 ;
  assign n17935 = n4857 & n10013 ;
  assign n17936 = n17934 | n17935 ;
  assign n17937 = x45 & x55 ;
  assign n17938 = n7528 & n17937 ;
  assign n17939 = x56 & n17938 ;
  assign n17940 = ( x56 & ~n17936 ) | ( x56 & n17939 ) | ( ~n17936 & n17939 ) ;
  assign n17941 = x37 & n17940 ;
  assign n17942 = n17936 | n17938 ;
  assign n17943 = x38 & x55 ;
  assign n17944 = ( n8925 & ~n17938 ) | ( n8925 & n17943 ) | ( ~n17938 & n17943 ) ;
  assign n17945 = n8925 & n17943 ;
  assign n17946 = ( ~n17936 & n17944 ) | ( ~n17936 & n17945 ) | ( n17944 & n17945 ) ;
  assign n17947 = ~n17942 & n17946 ;
  assign n17948 = n17941 | n17947 ;
  assign n17949 = n4969 & n10866 ;
  assign n17950 = n5407 & n7112 ;
  assign n17951 = n17949 | n17950 ;
  assign n17952 = n5658 & n6834 ;
  assign n17953 = x51 & n17952 ;
  assign n17954 = ( x51 & ~n17951 ) | ( x51 & n17953 ) | ( ~n17951 & n17953 ) ;
  assign n17955 = x42 & n17954 ;
  assign n17956 = n17951 | n17952 ;
  assign n17957 = x43 & x50 ;
  assign n17958 = ( n9005 & ~n17952 ) | ( n9005 & n17957 ) | ( ~n17952 & n17957 ) ;
  assign n17959 = n9005 & n17957 ;
  assign n17960 = ( ~n17951 & n17958 ) | ( ~n17951 & n17959 ) | ( n17958 & n17959 ) ;
  assign n17961 = ~n17956 & n17960 ;
  assign n17962 = n17955 | n17961 ;
  assign n17963 = n17948 & n17962 ;
  assign n17964 = n17948 & ~n17963 ;
  assign n17965 = n17962 & ~n17963 ;
  assign n17966 = n17964 | n17965 ;
  assign n17967 = ( x47 & x62 ) | ( x47 & ~n6147 ) | ( x62 & ~n6147 ) ;
  assign n17968 = x31 | x62 ;
  assign n17969 = ~x31 & x47 ;
  assign n17970 = ( n6147 & n17968 ) | ( n6147 & ~n17969 ) | ( n17968 & ~n17969 ) ;
  assign n17971 = ( ~x31 & x47 ) | ( ~x31 & x62 ) | ( x47 & x62 ) ;
  assign n17972 = ( x31 & n6147 ) | ( x31 & ~n17971 ) | ( n6147 & ~n17971 ) ;
  assign n17973 = ( n17967 & ~n17970 ) | ( n17967 & n17972 ) | ( ~n17970 & n17972 ) ;
  assign n17974 = ~n17966 & n17973 ;
  assign n17975 = n17966 & ~n17973 ;
  assign n17976 = n17974 | n17975 ;
  assign n17977 = n10413 & n12770 ;
  assign n17978 = n2546 & n10856 ;
  assign n17979 = n17977 | n17978 ;
  assign n17980 = n3321 & n10367 ;
  assign n17981 = x63 & n17980 ;
  assign n17982 = ( x63 & ~n17979 ) | ( x63 & n17981 ) | ( ~n17979 & n17981 ) ;
  assign n17983 = x30 & n17982 ;
  assign n17984 = n17979 | n17980 ;
  assign n17985 = x32 & x61 ;
  assign n17986 = x33 & x60 ;
  assign n17987 = ( ~n17980 & n17985 ) | ( ~n17980 & n17986 ) | ( n17985 & n17986 ) ;
  assign n17988 = n17985 & n17986 ;
  assign n17989 = ( ~n17979 & n17987 ) | ( ~n17979 & n17988 ) | ( n17987 & n17988 ) ;
  assign n17990 = ~n17984 & n17989 ;
  assign n17991 = n17983 | n17990 ;
  assign n17992 = n4078 & n9272 ;
  assign n17993 = x39 & x54 ;
  assign n17994 = n16852 & n17993 ;
  assign n17995 = n17992 | n17994 ;
  assign n17996 = n9771 & n15088 ;
  assign n17997 = n16852 & n17996 ;
  assign n17998 = ( n16852 & ~n17995 ) | ( n16852 & n17997 ) | ( ~n17995 & n17997 ) ;
  assign n17999 = n17995 | n17996 ;
  assign n18000 = x36 & x57 ;
  assign n18001 = ( n17993 & ~n17996 ) | ( n17993 & n18000 ) | ( ~n17996 & n18000 ) ;
  assign n18002 = n17993 & n18000 ;
  assign n18003 = ( ~n17995 & n18001 ) | ( ~n17995 & n18002 ) | ( n18001 & n18002 ) ;
  assign n18004 = ~n17999 & n18003 ;
  assign n18005 = n17998 | n18004 ;
  assign n18006 = n17991 & n18005 ;
  assign n18007 = n17991 & ~n18006 ;
  assign n18008 = x40 & x53 ;
  assign n18009 = x41 & x52 ;
  assign n18010 = n18008 | n18009 ;
  assign n18011 = n5813 & n8161 ;
  assign n18012 = n16830 & ~n18011 ;
  assign n18013 = n18010 | n18011 ;
  assign n18014 = ( n18011 & n18012 ) | ( n18011 & n18013 ) | ( n18012 & n18013 ) ;
  assign n18015 = n18010 & ~n18014 ;
  assign n18016 = n16830 & ~n18010 ;
  assign n18017 = ( n16830 & ~n18012 ) | ( n16830 & n18016 ) | ( ~n18012 & n18016 ) ;
  assign n18018 = n18015 | n18017 ;
  assign n18019 = ~n17991 & n18005 ;
  assign n18020 = n18018 & n18019 ;
  assign n18021 = ( n18007 & n18018 ) | ( n18007 & n18020 ) | ( n18018 & n18020 ) ;
  assign n18022 = n18018 | n18019 ;
  assign n18023 = n18007 | n18022 ;
  assign n18024 = ~n18021 & n18023 ;
  assign n18025 = n17976 | n18024 ;
  assign n18026 = n17976 & n18024 ;
  assign n18027 = n18025 & ~n18026 ;
  assign n18028 = n17793 | n17798 ;
  assign n18029 = ( n17793 & n17795 ) | ( n17793 & n18028 ) | ( n17795 & n18028 ) ;
  assign n18030 = n18027 & n18029 ;
  assign n18031 = n18027 | n18029 ;
  assign n18032 = ~n18030 & n18031 ;
  assign n18033 = n17765 | n17770 ;
  assign n18034 = n18032 & n18033 ;
  assign n18035 = n18032 | n18033 ;
  assign n18036 = ~n18034 & n18035 ;
  assign n18037 = ( n17801 & n17834 ) | ( n17801 & n17836 ) | ( n17834 & n17836 ) ;
  assign n18038 = n18036 | n18037 ;
  assign n18039 = n18036 & n18037 ;
  assign n18040 = n18038 & ~n18039 ;
  assign n18041 = ( n17781 & n17785 ) | ( n17781 & n17930 ) | ( n17785 & n17930 ) ;
  assign n18042 = n17781 & n17930 ;
  assign n18043 = ( n17783 & n18041 ) | ( n17783 & n18042 ) | ( n18041 & n18042 ) ;
  assign n18044 = n18040 & ~n18043 ;
  assign n18045 = n17933 & n18044 ;
  assign n18046 = ~n18040 & n18043 ;
  assign n18047 = ( n17933 & n18040 ) | ( n17933 & ~n18046 ) | ( n18040 & ~n18046 ) ;
  assign n18048 = ~n18045 & n18047 ;
  assign n18049 = n17788 | n17847 ;
  assign n18050 = ( n17847 & n17851 ) | ( n17847 & n18049 ) | ( n17851 & n18049 ) ;
  assign n18051 = ( n17884 & n18048 ) | ( n17884 & ~n18050 ) | ( n18048 & ~n18050 ) ;
  assign n18052 = ( ~n18048 & n18050 ) | ( ~n18048 & n18051 ) | ( n18050 & n18051 ) ;
  assign n18053 = ( ~n17884 & n18051 ) | ( ~n17884 & n18052 ) | ( n18051 & n18052 ) ;
  assign n18054 = n18048 & n18050 ;
  assign n18055 = n18048 | n18050 ;
  assign n18056 = n18054 | n18055 ;
  assign n18057 = ( n17866 & n18054 ) | ( n17866 & n18056 ) | ( n18054 & n18056 ) ;
  assign n18058 = ( n17882 & n18054 ) | ( n17882 & n18056 ) | ( n18054 & n18056 ) ;
  assign n18059 = ( n17871 & n18057 ) | ( n17871 & n18058 ) | ( n18057 & n18058 ) ;
  assign n18060 = ( n17877 & n18056 ) | ( n17877 & n18057 ) | ( n18056 & n18057 ) ;
  assign n18061 = ( n17122 & n18059 ) | ( n17122 & n18060 ) | ( n18059 & n18060 ) ;
  assign n18062 = n17907 | n17910 ;
  assign n18063 = ( n17907 & n17908 ) | ( n17907 & n18062 ) | ( n17908 & n18062 ) ;
  assign n18064 = n17751 | n17901 ;
  assign n18065 = ( n17901 & n17902 ) | ( n17901 & n18064 ) | ( n17902 & n18064 ) ;
  assign n18066 = n18063 | n18065 ;
  assign n18067 = n18063 & n18065 ;
  assign n18068 = n18066 & ~n18067 ;
  assign n18069 = n18006 | n18021 ;
  assign n18070 = n18068 | n18069 ;
  assign n18071 = n18068 & n18069 ;
  assign n18072 = n18070 & ~n18071 ;
  assign n18073 = n17914 | n17925 ;
  assign n18074 = n18072 & n18073 ;
  assign n18075 = n18072 | n18073 ;
  assign n18076 = ~n18074 & n18075 ;
  assign n18077 = n18026 | n18029 ;
  assign n18078 = ( n18026 & n18027 ) | ( n18026 & n18077 ) | ( n18027 & n18077 ) ;
  assign n18079 = n18076 & n18078 ;
  assign n18080 = n18076 | n18078 ;
  assign n18081 = ~n18079 & n18080 ;
  assign n18082 = n18034 | n18037 ;
  assign n18083 = ( n18034 & n18036 ) | ( n18034 & n18082 ) | ( n18036 & n18082 ) ;
  assign n18084 = n18081 | n18083 ;
  assign n18085 = n18081 & n18083 ;
  assign n18086 = n18084 & ~n18085 ;
  assign n18087 = x47 & x62 ;
  assign n18088 = x31 & n18087 ;
  assign n18089 = n6147 & ~n18088 ;
  assign n18090 = n14469 & n18088 ;
  assign n18091 = ( n14469 & n18089 ) | ( n14469 & n18090 ) | ( n18089 & n18090 ) ;
  assign n18092 = n14469 | n18088 ;
  assign n18093 = n18089 | n18092 ;
  assign n18094 = ~n18091 & n18093 ;
  assign n18095 = n17942 | n18094 ;
  assign n18096 = n17942 & n18094 ;
  assign n18097 = n18095 & ~n18096 ;
  assign n18098 = n17963 | n17973 ;
  assign n18099 = n18097 & n18098 ;
  assign n18100 = n17963 & n18097 ;
  assign n18101 = ( n17966 & n18099 ) | ( n17966 & n18100 ) | ( n18099 & n18100 ) ;
  assign n18102 = n18097 | n18098 ;
  assign n18103 = n17963 | n18097 ;
  assign n18104 = ( n17966 & n18102 ) | ( n17966 & n18103 ) | ( n18102 & n18103 ) ;
  assign n18105 = ~n18101 & n18104 ;
  assign n18106 = n17984 | n17999 ;
  assign n18107 = n17984 & n17999 ;
  assign n18108 = n18106 & ~n18107 ;
  assign n18109 = n18014 | n18108 ;
  assign n18110 = n18014 & n18108 ;
  assign n18111 = n18109 & ~n18110 ;
  assign n18112 = n18105 & n18111 ;
  assign n18113 = n18105 | n18111 ;
  assign n18114 = ~n18112 & n18113 ;
  assign n18115 = n17895 | n17927 ;
  assign n18116 = ( n17896 & n17927 ) | ( n17896 & n18115 ) | ( n17927 & n18115 ) ;
  assign n18117 = n18114 & n18116 ;
  assign n18118 = n17897 & n18114 ;
  assign n18119 = ( n17899 & n18117 ) | ( n17899 & n18118 ) | ( n18117 & n18118 ) ;
  assign n18120 = n18114 | n18116 ;
  assign n18121 = n17897 | n18114 ;
  assign n18122 = ( n17899 & n18120 ) | ( n17899 & n18121 ) | ( n18120 & n18121 ) ;
  assign n18123 = ~n18119 & n18122 ;
  assign n18124 = n6973 & n11935 ;
  assign n18125 = n5813 & n8355 ;
  assign n18126 = n18124 | n18125 ;
  assign n18127 = n5710 & n8161 ;
  assign n18128 = x54 & n18127 ;
  assign n18129 = ( x54 & ~n18126 ) | ( x54 & n18128 ) | ( ~n18126 & n18128 ) ;
  assign n18130 = x40 & n18129 ;
  assign n18131 = n18126 | n18127 ;
  assign n18132 = x42 & x52 ;
  assign n18133 = ( n8984 & ~n18127 ) | ( n8984 & n18132 ) | ( ~n18127 & n18132 ) ;
  assign n18134 = n8984 & n18132 ;
  assign n18135 = ( ~n18126 & n18133 ) | ( ~n18126 & n18134 ) | ( n18133 & n18134 ) ;
  assign n18136 = ~n18131 & n18135 ;
  assign n18137 = n18130 | n18136 ;
  assign n18138 = x43 & x51 ;
  assign n18139 = n9001 | n18138 ;
  assign n18140 = n5658 & n7112 ;
  assign n18141 = n18139 | n18140 ;
  assign n18142 = x36 & x58 ;
  assign n18143 = ( ~n18140 & n18141 ) | ( ~n18140 & n18142 ) | ( n18141 & n18142 ) ;
  assign n18144 = ( n18140 & n18141 ) | ( n18140 & ~n18142 ) | ( n18141 & ~n18142 ) ;
  assign n18145 = ( ~n18141 & n18143 ) | ( ~n18141 & n18144 ) | ( n18143 & n18144 ) ;
  assign n18146 = n18137 & n18145 ;
  assign n18147 = n18137 & ~n18146 ;
  assign n18148 = n9421 & n16143 ;
  assign n18149 = n9352 & n16143 ;
  assign n18150 = n5975 & n6759 ;
  assign n18151 = n18149 | n18150 ;
  assign n18152 = n9352 & n18148 ;
  assign n18153 = ( n9352 & ~n18151 ) | ( n9352 & n18152 ) | ( ~n18151 & n18152 ) ;
  assign n18154 = ( n9421 & n16143 ) | ( n9421 & ~n18151 ) | ( n16143 & ~n18151 ) ;
  assign n18155 = ( ~n18148 & n18153 ) | ( ~n18148 & n18154 ) | ( n18153 & n18154 ) ;
  assign n18156 = ~n18145 & n18155 ;
  assign n18157 = ( n18137 & n18155 ) | ( n18137 & n18156 ) | ( n18155 & n18156 ) ;
  assign n18158 = ~n18147 & n18157 ;
  assign n18159 = n18145 & ~n18155 ;
  assign n18160 = ~n18137 & n18159 ;
  assign n18161 = ( n18147 & ~n18155 ) | ( n18147 & n18160 ) | ( ~n18155 & n18160 ) ;
  assign n18162 = n18158 | n18161 ;
  assign n18163 = n17889 | n18162 ;
  assign n18164 = n17894 | n18163 ;
  assign n18165 = n17889 & n18162 ;
  assign n18166 = ( n17894 & n18162 ) | ( n17894 & n18165 ) | ( n18162 & n18165 ) ;
  assign n18167 = n18164 & ~n18166 ;
  assign n18168 = x59 & x62 ;
  assign n18169 = n7386 & n18168 ;
  assign n18170 = n3321 & n10684 ;
  assign n18171 = n18169 | n18170 ;
  assign n18172 = n3129 & n9737 ;
  assign n18173 = x62 & n18172 ;
  assign n18174 = ( x62 & ~n18171 ) | ( x62 & n18173 ) | ( ~n18171 & n18173 ) ;
  assign n18175 = x32 & n18174 ;
  assign n18176 = n18171 | n18172 ;
  assign n18177 = x33 & x61 ;
  assign n18178 = x35 & x59 ;
  assign n18179 = ( ~n18172 & n18177 ) | ( ~n18172 & n18178 ) | ( n18177 & n18178 ) ;
  assign n18180 = n18177 & n18178 ;
  assign n18181 = ( ~n18171 & n18179 ) | ( ~n18171 & n18180 ) | ( n18179 & n18180 ) ;
  assign n18182 = ~n18176 & n18181 ;
  assign n18183 = ~n17956 & n18182 ;
  assign n18184 = ( ~n17956 & n18175 ) | ( ~n17956 & n18183 ) | ( n18175 & n18183 ) ;
  assign n18185 = n17956 & ~n18182 ;
  assign n18186 = ~n18175 & n18185 ;
  assign n18187 = n18184 | n18186 ;
  assign n18188 = x34 & x60 ;
  assign n18189 = x39 & x55 ;
  assign n18190 = n18188 & n18189 ;
  assign n18191 = n5798 & n12860 ;
  assign n18192 = n12754 & n14647 ;
  assign n18193 = n18191 | n18192 ;
  assign n18194 = x57 & n18190 ;
  assign n18195 = ( x57 & ~n18193 ) | ( x57 & n18194 ) | ( ~n18193 & n18194 ) ;
  assign n18196 = x37 & n18195 ;
  assign n18197 = ( n18188 & n18189 ) | ( n18188 & ~n18193 ) | ( n18189 & ~n18193 ) ;
  assign n18198 = ( ~n18190 & n18196 ) | ( ~n18190 & n18197 ) | ( n18196 & n18197 ) ;
  assign n18199 = n18187 & n18198 ;
  assign n18200 = n18187 | n18198 ;
  assign n18201 = ~n18199 & n18200 ;
  assign n18202 = n18167 & n18201 ;
  assign n18203 = n18167 | n18201 ;
  assign n18204 = ~n18202 & n18203 ;
  assign n18205 = ~n18123 & n18204 ;
  assign n18206 = n18123 & ~n18204 ;
  assign n18207 = n18205 | n18206 ;
  assign n18208 = n18086 | n18207 ;
  assign n18209 = n18086 & n18207 ;
  assign n18210 = n18208 & ~n18209 ;
  assign n18211 = n18043 | n18045 ;
  assign n18212 = ( n18061 & n18210 ) | ( n18061 & ~n18211 ) | ( n18210 & ~n18211 ) ;
  assign n18213 = ( ~n18210 & n18211 ) | ( ~n18210 & n18212 ) | ( n18211 & n18212 ) ;
  assign n18214 = ( ~n18061 & n18212 ) | ( ~n18061 & n18213 ) | ( n18212 & n18213 ) ;
  assign n18215 = n18210 & n18211 ;
  assign n18216 = n18210 | n18211 ;
  assign n18217 = n18056 & n18216 ;
  assign n18218 = n18054 & n18216 ;
  assign n18219 = ( n17866 & n18217 ) | ( n17866 & n18218 ) | ( n18217 & n18218 ) ;
  assign n18220 = ( n17877 & n18217 ) | ( n17877 & n18219 ) | ( n18217 & n18219 ) ;
  assign n18221 = n18215 | n18220 ;
  assign n18222 = n18215 | n18216 ;
  assign n18223 = ( n18059 & n18215 ) | ( n18059 & n18222 ) | ( n18215 & n18222 ) ;
  assign n18224 = ( n17122 & n18221 ) | ( n17122 & n18223 ) | ( n18221 & n18223 ) ;
  assign n18225 = n18148 | n18151 ;
  assign n18226 = n4078 & n10370 ;
  assign n18227 = x36 & x59 ;
  assign n18228 = x35 & x60 ;
  assign n18229 = n18227 | n18228 ;
  assign n18230 = ~n18226 & n18229 ;
  assign n18231 = n18225 & n18230 ;
  assign n18232 = n18225 & ~n18231 ;
  assign n18233 = ~n18225 & n18230 ;
  assign n18234 = n18232 | n18233 ;
  assign n18235 = n17942 | n18091 ;
  assign n18236 = ( n18091 & n18094 ) | ( n18091 & n18235 ) | ( n18094 & n18235 ) ;
  assign n18237 = n18234 | n18236 ;
  assign n18238 = n18234 & n18236 ;
  assign n18239 = n18237 & ~n18238 ;
  assign n18240 = n18014 | n18107 ;
  assign n18241 = ( n18107 & n18108 ) | ( n18107 & n18240 ) | ( n18108 & n18240 ) ;
  assign n18242 = n18239 | n18241 ;
  assign n18243 = n18239 & n18241 ;
  assign n18244 = n18242 & ~n18243 ;
  assign n18245 = n18101 | n18111 ;
  assign n18246 = ( n18101 & n18105 ) | ( n18101 & n18245 ) | ( n18105 & n18245 ) ;
  assign n18247 = n18244 & n18246 ;
  assign n18248 = n18244 | n18246 ;
  assign n18249 = ~n18247 & n18248 ;
  assign n18250 = n18166 | n18201 ;
  assign n18251 = ( n18166 & n18167 ) | ( n18166 & n18250 ) | ( n18167 & n18250 ) ;
  assign n18252 = n18249 & n18251 ;
  assign n18253 = n18249 | n18251 ;
  assign n18254 = ~n18252 & n18253 ;
  assign n18255 = n18119 | n18204 ;
  assign n18256 = ( n18119 & n18123 ) | ( n18119 & n18255 ) | ( n18123 & n18255 ) ;
  assign n18257 = n18254 | n18256 ;
  assign n18258 = n18254 & n18256 ;
  assign n18259 = n18257 & ~n18258 ;
  assign n18260 = x46 & x49 ;
  assign n18261 = n9349 | n18260 ;
  assign n18262 = n5975 & n6834 ;
  assign n18263 = n18261 & ~n18262 ;
  assign n18264 = x39 & x56 ;
  assign n18265 = n18262 | n18264 ;
  assign n18266 = ( n18262 & n18263 ) | ( n18262 & n18265 ) | ( n18263 & n18265 ) ;
  assign n18267 = n18261 & ~n18266 ;
  assign n18268 = ~n18263 & n18264 ;
  assign n18269 = n18267 | n18268 ;
  assign n18270 = x48 & x62 ;
  assign n18271 = x33 & n18270 ;
  assign n18272 = n6762 & n18271 ;
  assign n18273 = n6762 & ~n18271 ;
  assign n18274 = n18271 | n18273 ;
  assign n18275 = x33 & x62 ;
  assign n18276 = ( x48 & ~n18271 ) | ( x48 & n18275 ) | ( ~n18271 & n18275 ) ;
  assign n18277 = x48 & n18275 ;
  assign n18278 = ( ~n18273 & n18276 ) | ( ~n18273 & n18277 ) | ( n18276 & n18277 ) ;
  assign n18279 = ~n18274 & n18278 ;
  assign n18280 = n18272 | n18279 ;
  assign n18281 = n18269 & n18280 ;
  assign n18282 = n18269 & ~n18281 ;
  assign n18283 = n4969 & n7874 ;
  assign n18284 = n5407 & n8161 ;
  assign n18285 = n18283 | n18284 ;
  assign n18286 = n5658 & n7567 ;
  assign n18287 = x53 & n18286 ;
  assign n18288 = ( x53 & ~n18285 ) | ( x53 & n18287 ) | ( ~n18285 & n18287 ) ;
  assign n18289 = x42 & n18288 ;
  assign n18290 = n18285 | n18286 ;
  assign n18291 = x43 & x52 ;
  assign n18292 = ( n9331 & ~n18286 ) | ( n9331 & n18291 ) | ( ~n18286 & n18291 ) ;
  assign n18293 = n9331 & n18291 ;
  assign n18294 = ( ~n18285 & n18292 ) | ( ~n18285 & n18293 ) | ( n18292 & n18293 ) ;
  assign n18295 = ~n18290 & n18294 ;
  assign n18296 = n18289 | n18295 ;
  assign n18297 = ~n18269 & n18280 ;
  assign n18298 = n18296 & n18297 ;
  assign n18299 = ( n18282 & n18296 ) | ( n18282 & n18298 ) | ( n18296 & n18298 ) ;
  assign n18300 = n18296 | n18297 ;
  assign n18301 = n18282 | n18300 ;
  assign n18302 = ~n18299 & n18301 ;
  assign n18303 = n18067 | n18068 ;
  assign n18304 = ( n18067 & n18069 ) | ( n18067 & n18303 ) | ( n18069 & n18303 ) ;
  assign n18305 = n18302 | n18304 ;
  assign n18306 = n18302 & n18304 ;
  assign n18307 = n18305 & ~n18306 ;
  assign n18308 = ~n18140 & n18142 ;
  assign n18309 = ( n18140 & n18141 ) | ( n18140 & n18308 ) | ( n18141 & n18308 ) ;
  assign n18310 = x55 & x58 ;
  assign n18311 = n6159 & n18310 ;
  assign n18312 = n4857 & n9272 ;
  assign n18313 = n18311 | n18312 ;
  assign n18314 = n4050 & n12860 ;
  assign n18315 = x37 & n18314 ;
  assign n18316 = ( x37 & ~n18313 ) | ( x37 & n18315 ) | ( ~n18313 & n18315 ) ;
  assign n18317 = x58 & n18316 ;
  assign n18318 = n18313 | n18314 ;
  assign n18319 = x38 & x57 ;
  assign n18320 = x40 & x55 ;
  assign n18321 = ( ~n18314 & n18319 ) | ( ~n18314 & n18320 ) | ( n18319 & n18320 ) ;
  assign n18322 = n18319 & n18320 ;
  assign n18323 = ( ~n18313 & n18321 ) | ( ~n18313 & n18322 ) | ( n18321 & n18322 ) ;
  assign n18324 = ~n18318 & n18323 ;
  assign n18325 = n18317 | n18324 ;
  assign n18326 = n18309 & n18325 ;
  assign n18327 = n18309 | n18325 ;
  assign n18328 = ~n18326 & n18327 ;
  assign n18329 = x32 & x63 ;
  assign n18330 = x34 & x61 ;
  assign n18331 = n18329 | n18330 ;
  assign n18332 = n4318 & n10856 ;
  assign n18333 = n18331 | n18332 ;
  assign n18334 = x41 & x54 ;
  assign n18335 = ( ~n18332 & n18333 ) | ( ~n18332 & n18334 ) | ( n18333 & n18334 ) ;
  assign n18336 = ( n18332 & n18333 ) | ( n18332 & ~n18334 ) | ( n18333 & ~n18334 ) ;
  assign n18337 = ( ~n18333 & n18335 ) | ( ~n18333 & n18336 ) | ( n18335 & n18336 ) ;
  assign n18338 = n18328 & n18337 ;
  assign n18339 = n18328 & ~n18338 ;
  assign n18340 = ~n18328 & n18337 ;
  assign n18341 = n18339 | n18340 ;
  assign n18342 = ~n18307 & n18341 ;
  assign n18343 = n18307 & ~n18341 ;
  assign n18344 = n18342 | n18343 ;
  assign n18345 = n18190 | n18193 ;
  assign n18346 = n18176 | n18345 ;
  assign n18347 = n18176 & n18345 ;
  assign n18348 = n18346 & ~n18347 ;
  assign n18349 = n18131 | n18348 ;
  assign n18350 = n18131 & n18348 ;
  assign n18351 = n18349 & ~n18350 ;
  assign n18352 = n18175 | n18182 ;
  assign n18353 = ( n17956 & n18198 ) | ( n17956 & n18352 ) | ( n18198 & n18352 ) ;
  assign n18354 = ~n18137 & n18145 ;
  assign n18355 = n18145 | n18155 ;
  assign n18356 = ( n18137 & n18155 ) | ( n18137 & n18355 ) | ( n18155 & n18355 ) ;
  assign n18357 = ( n18146 & n18354 ) | ( n18146 & n18356 ) | ( n18354 & n18356 ) ;
  assign n18358 = n18146 | n18356 ;
  assign n18359 = ( n18147 & n18357 ) | ( n18147 & n18358 ) | ( n18357 & n18358 ) ;
  assign n18360 = n18353 & n18359 ;
  assign n18361 = n18353 | n18359 ;
  assign n18362 = ~n18360 & n18361 ;
  assign n18363 = n18351 & n18362 ;
  assign n18364 = n18351 | n18362 ;
  assign n18365 = ~n18363 & n18364 ;
  assign n18366 = n18074 & n18365 ;
  assign n18367 = ( n18079 & n18365 ) | ( n18079 & n18366 ) | ( n18365 & n18366 ) ;
  assign n18368 = n18074 | n18365 ;
  assign n18369 = n18079 | n18368 ;
  assign n18370 = ~n18367 & n18369 ;
  assign n18371 = ~n18344 & n18370 ;
  assign n18372 = n18344 & ~n18370 ;
  assign n18373 = n18371 | n18372 ;
  assign n18374 = ~n18259 & n18373 ;
  assign n18375 = n18259 & ~n18373 ;
  assign n18376 = n18374 | n18375 ;
  assign n18377 = n18085 | n18207 ;
  assign n18378 = ( n18085 & n18086 ) | ( n18085 & n18377 ) | ( n18086 & n18377 ) ;
  assign n18379 = ( n18224 & n18376 ) | ( n18224 & ~n18378 ) | ( n18376 & ~n18378 ) ;
  assign n18380 = ( ~n18376 & n18378 ) | ( ~n18376 & n18379 ) | ( n18378 & n18379 ) ;
  assign n18381 = ( ~n18224 & n18379 ) | ( ~n18224 & n18380 ) | ( n18379 & n18380 ) ;
  assign n18382 = n18074 | n18079 ;
  assign n18383 = ( n18344 & n18365 ) | ( n18344 & n18382 ) | ( n18365 & n18382 ) ;
  assign n18384 = ( n18302 & n18304 ) | ( n18302 & n18341 ) | ( n18304 & n18341 ) ;
  assign n18430 = n18351 | n18353 ;
  assign n18431 = ( n18351 & n18359 ) | ( n18351 & n18430 ) | ( n18359 & n18430 ) ;
  assign n18432 = ( n18360 & n18362 ) | ( n18360 & n18431 ) | ( n18362 & n18431 ) ;
  assign n18385 = n3770 & n10370 ;
  assign n18386 = x40 & x60 ;
  assign n18387 = n17724 & n18386 ;
  assign n18388 = n18385 | n18387 ;
  assign n18389 = n6159 & n15336 ;
  assign n18390 = x60 & n18389 ;
  assign n18391 = ( x60 & ~n18388 ) | ( x60 & n18390 ) | ( ~n18388 & n18390 ) ;
  assign n18392 = x36 & n18391 ;
  assign n18393 = n18388 | n18389 ;
  assign n18394 = x37 & x59 ;
  assign n18395 = x40 & x56 ;
  assign n18396 = ( ~n18389 & n18394 ) | ( ~n18389 & n18395 ) | ( n18394 & n18395 ) ;
  assign n18397 = n18394 & n18395 ;
  assign n18398 = ( ~n18388 & n18396 ) | ( ~n18388 & n18397 ) | ( n18396 & n18397 ) ;
  assign n18399 = ~n18393 & n18398 ;
  assign n18400 = n18392 | n18399 ;
  assign n18401 = x38 & x58 ;
  assign n18402 = x39 & x57 ;
  assign n18403 = n18401 | n18402 ;
  assign n18404 = n5392 & n9272 ;
  assign n18405 = n9499 & ~n18404 ;
  assign n18406 = n18403 | n18404 ;
  assign n18407 = ( n18404 & n18405 ) | ( n18404 & n18406 ) | ( n18405 & n18406 ) ;
  assign n18408 = n18403 & ~n18407 ;
  assign n18409 = n9499 & ~n18403 ;
  assign n18410 = ( n9499 & ~n18405 ) | ( n9499 & n18409 ) | ( ~n18405 & n18409 ) ;
  assign n18411 = n18408 | n18410 ;
  assign n18412 = n18400 & n18411 ;
  assign n18413 = n18400 & ~n18412 ;
  assign n18414 = n18411 & ~n18412 ;
  assign n18415 = n18413 | n18414 ;
  assign n18416 = x45 & x51 ;
  assign n18417 = n6757 & n18416 ;
  assign n18418 = n5975 & n7112 ;
  assign n18419 = n18417 | n18418 ;
  assign n18420 = n6147 & n6834 ;
  assign n18421 = n18416 & n18420 ;
  assign n18422 = x46 & x50 ;
  assign n18423 = n6757 | n18422 ;
  assign n18424 = n18416 | n18423 ;
  assign n18425 = ( n18419 & ~n18420 ) | ( n18419 & n18424 ) | ( ~n18420 & n18424 ) ;
  assign n18426 = ( ~n18419 & n18421 ) | ( ~n18419 & n18425 ) | ( n18421 & n18425 ) ;
  assign n18427 = ~n18415 & n18426 ;
  assign n18428 = n18415 & ~n18426 ;
  assign n18429 = n18427 | n18428 ;
  assign n18433 = n18429 & n18432 ;
  assign n18434 = n18432 & ~n18433 ;
  assign n18435 = n18429 & ~n18432 ;
  assign n18436 = n18384 & n18435 ;
  assign n18437 = ( n18384 & n18434 ) | ( n18384 & n18436 ) | ( n18434 & n18436 ) ;
  assign n18438 = n18384 & ~n18437 ;
  assign n18439 = n18434 | n18435 ;
  assign n18440 = ~n18437 & n18439 ;
  assign n18441 = n18438 | n18440 ;
  assign n18442 = n18383 & n18441 ;
  assign n18443 = n18383 & ~n18442 ;
  assign n18444 = n18266 | n18274 ;
  assign n18445 = n18266 & n18274 ;
  assign n18446 = n18444 & ~n18445 ;
  assign n18447 = n18290 | n18446 ;
  assign n18448 = n18290 & n18446 ;
  assign n18449 = n18447 & ~n18448 ;
  assign n18450 = n18281 | n18299 ;
  assign n18451 = n18309 | n18337 ;
  assign n18452 = ( n18325 & n18337 ) | ( n18325 & n18451 ) | ( n18337 & n18451 ) ;
  assign n18453 = ( n18326 & n18328 ) | ( n18326 & n18452 ) | ( n18328 & n18452 ) ;
  assign n18454 = n18450 | n18453 ;
  assign n18455 = n18450 & n18453 ;
  assign n18456 = n18454 & ~n18455 ;
  assign n18457 = n18449 & n18456 ;
  assign n18458 = n18449 | n18456 ;
  assign n18459 = ~n18457 & n18458 ;
  assign n18460 = n18247 & n18459 ;
  assign n18461 = ( n18252 & n18459 ) | ( n18252 & n18460 ) | ( n18459 & n18460 ) ;
  assign n18462 = n18247 | n18459 ;
  assign n18463 = n18252 | n18462 ;
  assign n18464 = ~n18461 & n18463 ;
  assign n18465 = n3129 & n10856 ;
  assign n18466 = n4530 & n10561 ;
  assign n18467 = n18465 | n18466 ;
  assign n18468 = n3483 & n10684 ;
  assign n18469 = x63 & n18468 ;
  assign n18470 = ( x63 & ~n18467 ) | ( x63 & n18469 ) | ( ~n18467 & n18469 ) ;
  assign n18471 = x33 & n18470 ;
  assign n18472 = n18467 | n18468 ;
  assign n18473 = x34 & x62 ;
  assign n18474 = x35 & x61 ;
  assign n18475 = ( ~n18468 & n18473 ) | ( ~n18468 & n18474 ) | ( n18473 & n18474 ) ;
  assign n18476 = n18473 & n18474 ;
  assign n18477 = ( ~n18467 & n18475 ) | ( ~n18467 & n18476 ) | ( n18475 & n18476 ) ;
  assign n18478 = ~n18472 & n18477 ;
  assign n18479 = n18471 | n18478 ;
  assign n18480 = x43 & x53 ;
  assign n18481 = n9441 & n18480 ;
  assign n18482 = n5710 & n8357 ;
  assign n18483 = n18481 | n18482 ;
  assign n18484 = n5407 & n8355 ;
  assign n18485 = n9441 & n18484 ;
  assign n18486 = ( n9441 & ~n18483 ) | ( n9441 & n18485 ) | ( ~n18483 & n18485 ) ;
  assign n18487 = n18483 | n18484 ;
  assign n18488 = x42 & x54 ;
  assign n18489 = ( n18480 & ~n18484 ) | ( n18480 & n18488 ) | ( ~n18484 & n18488 ) ;
  assign n18490 = n18480 & n18488 ;
  assign n18491 = ( ~n18483 & n18489 ) | ( ~n18483 & n18490 ) | ( n18489 & n18490 ) ;
  assign n18492 = ~n18487 & n18491 ;
  assign n18493 = n18486 | n18492 ;
  assign n18494 = n18479 & n18493 ;
  assign n18495 = n18479 & ~n18494 ;
  assign n18497 = n18131 | n18347 ;
  assign n18498 = ( n18347 & n18348 ) | ( n18347 & n18497 ) | ( n18348 & n18497 ) ;
  assign n18496 = ~n18479 & n18493 ;
  assign n18499 = n18496 & n18498 ;
  assign n18500 = ( n18495 & n18498 ) | ( n18495 & n18499 ) | ( n18498 & n18499 ) ;
  assign n18501 = n18496 | n18498 ;
  assign n18502 = n18495 | n18501 ;
  assign n18503 = ~n18500 & n18502 ;
  assign n18504 = ~n18332 & n18334 ;
  assign n18505 = ( n18332 & n18333 ) | ( n18332 & n18504 ) | ( n18333 & n18504 ) ;
  assign n18506 = n18318 | n18505 ;
  assign n18507 = n18318 & n18505 ;
  assign n18508 = n18506 & ~n18507 ;
  assign n18509 = n18226 | n18230 ;
  assign n18510 = ( n18225 & n18226 ) | ( n18225 & n18509 ) | ( n18226 & n18509 ) ;
  assign n18511 = n18508 | n18510 ;
  assign n18512 = n18508 & n18510 ;
  assign n18513 = n18511 & ~n18512 ;
  assign n18514 = n18238 | n18241 ;
  assign n18515 = ( n18238 & n18239 ) | ( n18238 & n18514 ) | ( n18239 & n18514 ) ;
  assign n18516 = n18513 | n18515 ;
  assign n18517 = n18513 & n18515 ;
  assign n18518 = n18516 & ~n18517 ;
  assign n18519 = n18503 & n18518 ;
  assign n18520 = n18503 | n18518 ;
  assign n18521 = ~n18519 & n18520 ;
  assign n18522 = n18464 & n18521 ;
  assign n18523 = n18464 | n18521 ;
  assign n18524 = ~n18522 & n18523 ;
  assign n18525 = ~n18383 & n18441 ;
  assign n18526 = n18524 & n18525 ;
  assign n18527 = ( n18443 & n18524 ) | ( n18443 & n18526 ) | ( n18524 & n18526 ) ;
  assign n18528 = n18524 | n18525 ;
  assign n18529 = n18443 | n18528 ;
  assign n18530 = ~n18527 & n18529 ;
  assign n18531 = n18258 | n18373 ;
  assign n18532 = ( n18258 & n18259 ) | ( n18258 & n18531 ) | ( n18259 & n18531 ) ;
  assign n18533 = n18530 | n18532 ;
  assign n18534 = n18530 & n18532 ;
  assign n18535 = n18533 & ~n18534 ;
  assign n18536 = n18376 & n18378 ;
  assign n18537 = n18376 | n18378 ;
  assign n18538 = n18215 & n18537 ;
  assign n18539 = n18536 | n18538 ;
  assign n18540 = n18536 | n18537 ;
  assign n18541 = ( n18222 & n18536 ) | ( n18222 & n18540 ) | ( n18536 & n18540 ) ;
  assign n18542 = ( n18059 & n18539 ) | ( n18059 & n18541 ) | ( n18539 & n18541 ) ;
  assign n18543 = ( n18220 & n18539 ) | ( n18220 & n18540 ) | ( n18539 & n18540 ) ;
  assign n18544 = ( n17122 & n18542 ) | ( n17122 & n18543 ) | ( n18542 & n18543 ) ;
  assign n18545 = n18535 | n18544 ;
  assign n18546 = n18533 & n18540 ;
  assign n18547 = n18533 & n18536 ;
  assign n18548 = ( n18533 & n18538 ) | ( n18533 & n18547 ) | ( n18538 & n18547 ) ;
  assign n18549 = ( n18220 & n18546 ) | ( n18220 & n18548 ) | ( n18546 & n18548 ) ;
  assign n18550 = n18533 & n18541 ;
  assign n18551 = ( n18058 & n18548 ) | ( n18058 & n18550 ) | ( n18548 & n18550 ) ;
  assign n18552 = ( n18057 & n18548 ) | ( n18057 & n18550 ) | ( n18548 & n18550 ) ;
  assign n18553 = ( n17871 & n18551 ) | ( n17871 & n18552 ) | ( n18551 & n18552 ) ;
  assign n18554 = ( n17122 & n18549 ) | ( n17122 & n18553 ) | ( n18549 & n18553 ) ;
  assign n18555 = ~n18534 & n18554 ;
  assign n18556 = n18545 & ~n18555 ;
  assign n18557 = n18534 | n18553 ;
  assign n18558 = n18534 | n18548 ;
  assign n18559 = n18533 | n18534 ;
  assign n18560 = ( n18534 & n18540 ) | ( n18534 & n18559 ) | ( n18540 & n18559 ) ;
  assign n18561 = ( n18219 & n18558 ) | ( n18219 & n18560 ) | ( n18558 & n18560 ) ;
  assign n18562 = ( n18217 & n18558 ) | ( n18217 & n18560 ) | ( n18558 & n18560 ) ;
  assign n18563 = ( n17877 & n18561 ) | ( n17877 & n18562 ) | ( n18561 & n18562 ) ;
  assign n18564 = ( n17122 & n18557 ) | ( n17122 & n18563 ) | ( n18557 & n18563 ) ;
  assign n18565 = x36 & x61 ;
  assign n18566 = n18420 & n18565 ;
  assign n18567 = ( n18419 & n18565 ) | ( n18419 & n18566 ) | ( n18565 & n18566 ) ;
  assign n18568 = n18420 | n18565 ;
  assign n18569 = n18419 | n18568 ;
  assign n18570 = ~n18567 & n18569 ;
  assign n18571 = n18407 | n18570 ;
  assign n18572 = n18407 & n18570 ;
  assign n18573 = n18571 & ~n18572 ;
  assign n18574 = n18412 | n18426 ;
  assign n18575 = n18507 | n18510 ;
  assign n18576 = ( n18507 & n18508 ) | ( n18507 & n18575 ) | ( n18508 & n18575 ) ;
  assign n18577 = n18574 & n18576 ;
  assign n18578 = n18412 & n18576 ;
  assign n18579 = ( n18415 & n18577 ) | ( n18415 & n18578 ) | ( n18577 & n18578 ) ;
  assign n18580 = n18574 | n18576 ;
  assign n18581 = n18412 | n18576 ;
  assign n18582 = ( n18415 & n18580 ) | ( n18415 & n18581 ) | ( n18580 & n18581 ) ;
  assign n18583 = ~n18579 & n18582 ;
  assign n18584 = n18573 & n18583 ;
  assign n18585 = n18573 | n18583 ;
  assign n18586 = ~n18584 & n18585 ;
  assign n18587 = x47 & x50 ;
  assign n18588 = n9702 | n18587 ;
  assign n18589 = n6147 & n7112 ;
  assign n18590 = x40 & x57 ;
  assign n18591 = ~n18589 & n18590 ;
  assign n18592 = n18588 | n18589 ;
  assign n18593 = ( n18589 & n18591 ) | ( n18589 & n18592 ) | ( n18591 & n18592 ) ;
  assign n18594 = n18588 & ~n18593 ;
  assign n18595 = ( ~n18588 & n18589 ) | ( ~n18588 & n18590 ) | ( n18589 & n18590 ) ;
  assign n18596 = n18590 & n18595 ;
  assign n18597 = n18594 | n18596 ;
  assign n18598 = x49 & x62 ;
  assign n18599 = x35 & n18598 ;
  assign n18600 = n6759 & n18599 ;
  assign n18601 = n6759 & ~n18599 ;
  assign n18602 = n18599 | n18601 ;
  assign n18603 = x35 & x62 ;
  assign n18604 = ( x49 & ~n18599 ) | ( x49 & n18603 ) | ( ~n18599 & n18603 ) ;
  assign n18605 = x49 & n18603 ;
  assign n18606 = ( ~n18601 & n18604 ) | ( ~n18601 & n18605 ) | ( n18604 & n18605 ) ;
  assign n18607 = ~n18602 & n18606 ;
  assign n18608 = n18600 | n18607 ;
  assign n18609 = n18597 & n18608 ;
  assign n18610 = n18597 & ~n18609 ;
  assign n18612 = n18290 | n18445 ;
  assign n18613 = ( n18445 & n18446 ) | ( n18445 & n18612 ) | ( n18446 & n18612 ) ;
  assign n18611 = ~n18597 & n18608 ;
  assign n18614 = n18611 & n18613 ;
  assign n18615 = ( n18610 & n18613 ) | ( n18610 & n18614 ) | ( n18613 & n18614 ) ;
  assign n18616 = n18611 | n18613 ;
  assign n18617 = n18610 | n18616 ;
  assign n18618 = ~n18615 & n18617 ;
  assign n18619 = n18393 | n18472 ;
  assign n18620 = n18393 & n18472 ;
  assign n18621 = n18619 & ~n18620 ;
  assign n18622 = n18487 | n18621 ;
  assign n18623 = n18487 & n18621 ;
  assign n18624 = n18622 & ~n18623 ;
  assign n18625 = n18494 & n18624 ;
  assign n18626 = ( n18500 & n18624 ) | ( n18500 & n18625 ) | ( n18624 & n18625 ) ;
  assign n18627 = n18494 | n18624 ;
  assign n18628 = n18500 | n18627 ;
  assign n18629 = ~n18626 & n18628 ;
  assign n18630 = n18618 & n18629 ;
  assign n18631 = n18618 | n18629 ;
  assign n18632 = ~n18630 & n18631 ;
  assign n18633 = n18586 & n18632 ;
  assign n18634 = n18586 | n18632 ;
  assign n18635 = ~n18633 & n18634 ;
  assign n18636 = n18433 & n18635 ;
  assign n18637 = ( n18437 & n18635 ) | ( n18437 & n18636 ) | ( n18635 & n18636 ) ;
  assign n18638 = n18433 | n18635 ;
  assign n18639 = n18437 | n18638 ;
  assign n18640 = ~n18637 & n18639 ;
  assign n18641 = n18449 | n18453 ;
  assign n18642 = ( n18449 & n18450 ) | ( n18449 & n18641 ) | ( n18450 & n18641 ) ;
  assign n18643 = ( n18455 & n18456 ) | ( n18455 & n18642 ) | ( n18456 & n18642 ) ;
  assign n18644 = n5798 & n10975 ;
  assign n18645 = n4857 & n10370 ;
  assign n18646 = n18644 | n18645 ;
  assign n18647 = n5392 & n9831 ;
  assign n18648 = x60 & n18647 ;
  assign n18649 = ( x60 & ~n18646 ) | ( x60 & n18648 ) | ( ~n18646 & n18648 ) ;
  assign n18650 = x37 & n18649 ;
  assign n18651 = n18646 | n18647 ;
  assign n18652 = x38 & x59 ;
  assign n18653 = x39 & x58 ;
  assign n18654 = ( ~n18647 & n18652 ) | ( ~n18647 & n18653 ) | ( n18652 & n18653 ) ;
  assign n18655 = n18652 & n18653 ;
  assign n18656 = ( ~n18646 & n18654 ) | ( ~n18646 & n18655 ) | ( n18654 & n18655 ) ;
  assign n18657 = ~n18651 & n18656 ;
  assign n18658 = n18650 | n18657 ;
  assign n18659 = x34 & x63 ;
  assign n18660 = x41 & x56 ;
  assign n18661 = x42 & x55 ;
  assign n18662 = ( ~n18659 & n18660 ) | ( ~n18659 & n18661 ) | ( n18660 & n18661 ) ;
  assign n18663 = n5710 & n10013 ;
  assign n18664 = n18660 | n18661 ;
  assign n18665 = ( n18659 & n18663 ) | ( n18659 & n18664 ) | ( n18663 & n18664 ) ;
  assign n18666 = ( n18659 & n18662 ) | ( n18659 & ~n18665 ) | ( n18662 & ~n18665 ) ;
  assign n18667 = n18658 & n18666 ;
  assign n18668 = n18658 & ~n18667 ;
  assign n18669 = n5104 & n11935 ;
  assign n18670 = n5658 & n8355 ;
  assign n18671 = n18669 | n18670 ;
  assign n18672 = n6093 & n8161 ;
  assign n18673 = x54 & n18672 ;
  assign n18674 = ( x54 & ~n18671 ) | ( x54 & n18673 ) | ( ~n18671 & n18673 ) ;
  assign n18675 = x43 & n18674 ;
  assign n18676 = n18671 | n18672 ;
  assign n18677 = x44 & x53 ;
  assign n18678 = ( n9959 & ~n18672 ) | ( n9959 & n18677 ) | ( ~n18672 & n18677 ) ;
  assign n18679 = n9959 & n18677 ;
  assign n18680 = ( ~n18671 & n18678 ) | ( ~n18671 & n18679 ) | ( n18678 & n18679 ) ;
  assign n18681 = ~n18676 & n18680 ;
  assign n18682 = n18675 | n18681 ;
  assign n18683 = ~n18658 & n18666 ;
  assign n18684 = n18682 & n18683 ;
  assign n18685 = ( n18668 & n18682 ) | ( n18668 & n18684 ) | ( n18682 & n18684 ) ;
  assign n18686 = n18682 | n18683 ;
  assign n18687 = n18668 | n18686 ;
  assign n18688 = ~n18685 & n18687 ;
  assign n18689 = n18642 & n18688 ;
  assign n18690 = n18455 & n18688 ;
  assign n18691 = ( n18456 & n18689 ) | ( n18456 & n18690 ) | ( n18689 & n18690 ) ;
  assign n18692 = n18643 & ~n18691 ;
  assign n18693 = n18503 | n18517 ;
  assign n18694 = ( n18517 & n18518 ) | ( n18517 & n18693 ) | ( n18518 & n18693 ) ;
  assign n18695 = ~n18642 & n18688 ;
  assign n18696 = ~n18455 & n18688 ;
  assign n18697 = ( ~n18456 & n18695 ) | ( ~n18456 & n18696 ) | ( n18695 & n18696 ) ;
  assign n18698 = n18694 & n18697 ;
  assign n18699 = ( n18692 & n18694 ) | ( n18692 & n18698 ) | ( n18694 & n18698 ) ;
  assign n18700 = n18694 | n18697 ;
  assign n18701 = n18692 | n18700 ;
  assign n18702 = ~n18699 & n18701 ;
  assign n18703 = n18461 | n18521 ;
  assign n18704 = ( n18461 & n18464 ) | ( n18461 & n18703 ) | ( n18464 & n18703 ) ;
  assign n18705 = n18702 & n18704 ;
  assign n18706 = n18702 | n18704 ;
  assign n18707 = ~n18705 & n18706 ;
  assign n18708 = n18640 & n18707 ;
  assign n18709 = n18640 | n18707 ;
  assign n18710 = ~n18708 & n18709 ;
  assign n18711 = n18442 | n18524 ;
  assign n18712 = n18442 | n18443 ;
  assign n18713 = ( n18526 & n18711 ) | ( n18526 & n18712 ) | ( n18711 & n18712 ) ;
  assign n18714 = ( n18564 & ~n18710 ) | ( n18564 & n18713 ) | ( ~n18710 & n18713 ) ;
  assign n18715 = ( n18710 & ~n18713 ) | ( n18710 & n18714 ) | ( ~n18713 & n18714 ) ;
  assign n18716 = ( ~n18564 & n18714 ) | ( ~n18564 & n18715 ) | ( n18714 & n18715 ) ;
  assign n18717 = n18710 & n18713 ;
  assign n18718 = n18710 | n18713 ;
  assign n18719 = n18717 | n18718 ;
  assign n18720 = ( n18564 & n18717 ) | ( n18564 & n18719 ) | ( n18717 & n18719 ) ;
  assign n18721 = n18659 & n18660 ;
  assign n18722 = n18663 | n18721 ;
  assign n18723 = n18659 & n18661 ;
  assign n18724 = n18722 | n18723 ;
  assign n18725 = n18651 | n18724 ;
  assign n18726 = n18651 & n18724 ;
  assign n18727 = n18725 & ~n18726 ;
  assign n18728 = n18676 | n18727 ;
  assign n18729 = n18676 & n18727 ;
  assign n18730 = n18728 & ~n18729 ;
  assign n18731 = n18609 & n18730 ;
  assign n18732 = ( n18615 & n18730 ) | ( n18615 & n18731 ) | ( n18730 & n18731 ) ;
  assign n18733 = n18609 | n18730 ;
  assign n18734 = n18615 | n18733 ;
  assign n18735 = ~n18732 & n18734 ;
  assign n18736 = n6147 & n7567 ;
  assign n18737 = x48 & x52 ;
  assign n18738 = n18422 & n18737 ;
  assign n18739 = n18736 | n18738 ;
  assign n18740 = n6762 & n7112 ;
  assign n18741 = x52 & n18740 ;
  assign n18742 = ( x52 & ~n18739 ) | ( x52 & n18741 ) | ( ~n18739 & n18741 ) ;
  assign n18743 = x46 & n18742 ;
  assign n18744 = n18739 | n18740 ;
  assign n18745 = ( n6345 & n9978 ) | ( n6345 & ~n18740 ) | ( n9978 & ~n18740 ) ;
  assign n18746 = n6345 & n9978 ;
  assign n18747 = ( ~n18739 & n18745 ) | ( ~n18739 & n18746 ) | ( n18745 & n18746 ) ;
  assign n18748 = ~n18744 & n18747 ;
  assign n18749 = n18743 | n18748 ;
  assign n18750 = x39 & x59 ;
  assign n18751 = x40 & x58 ;
  assign n18752 = n18750 | n18751 ;
  assign n18753 = n4555 & n9831 ;
  assign n18754 = n18752 | n18753 ;
  assign n18755 = x45 & x53 ;
  assign n18756 = ( ~n18753 & n18754 ) | ( ~n18753 & n18755 ) | ( n18754 & n18755 ) ;
  assign n18757 = ( n18753 & n18754 ) | ( n18753 & ~n18755 ) | ( n18754 & ~n18755 ) ;
  assign n18758 = ( ~n18754 & n18756 ) | ( ~n18754 & n18757 ) | ( n18756 & n18757 ) ;
  assign n18759 = n18749 & n18758 ;
  assign n18760 = n18749 & ~n18759 ;
  assign n18761 = n3770 & n10684 ;
  assign n18762 = x37 & x61 ;
  assign n18763 = n12738 | n18762 ;
  assign n18764 = ~n18761 & n18763 ;
  assign n18765 = n18602 & n18764 ;
  assign n18766 = n18602 | n18764 ;
  assign n18767 = ~n18765 & n18766 ;
  assign n18768 = ~n18749 & n18758 ;
  assign n18769 = n18767 & ~n18768 ;
  assign n18770 = ~n18760 & n18769 ;
  assign n18771 = ~n18767 & n18768 ;
  assign n18772 = ( n18760 & ~n18767 ) | ( n18760 & n18771 ) | ( ~n18767 & n18771 ) ;
  assign n18773 = n18770 | n18772 ;
  assign n18774 = n18735 & n18773 ;
  assign n18775 = n18735 & ~n18774 ;
  assign n18776 = n18487 | n18620 ;
  assign n18777 = ( n18620 & n18621 ) | ( n18620 & n18776 ) | ( n18621 & n18776 ) ;
  assign n18778 = n18407 | n18567 ;
  assign n18779 = ( n18567 & n18570 ) | ( n18567 & n18778 ) | ( n18570 & n18778 ) ;
  assign n18780 = n18777 | n18779 ;
  assign n18781 = n18777 & n18779 ;
  assign n18782 = n18780 & ~n18781 ;
  assign n18783 = n18667 | n18685 ;
  assign n18784 = n18782 | n18783 ;
  assign n18785 = n18782 & n18783 ;
  assign n18786 = n18784 & ~n18785 ;
  assign n18787 = ~n18735 & n18773 ;
  assign n18788 = n18786 | n18787 ;
  assign n18789 = n18775 | n18788 ;
  assign n18790 = n18691 & n18789 ;
  assign n18791 = ( n18699 & n18789 ) | ( n18699 & n18790 ) | ( n18789 & n18790 ) ;
  assign n18792 = n18786 & n18787 ;
  assign n18793 = ( n18775 & n18786 ) | ( n18775 & n18792 ) | ( n18786 & n18792 ) ;
  assign n18794 = n18691 | n18789 ;
  assign n18795 = n18699 | n18794 ;
  assign n18796 = ( n18791 & ~n18793 ) | ( n18791 & n18795 ) | ( ~n18793 & n18795 ) ;
  assign n18797 = n18691 & n18793 ;
  assign n18798 = ( n18699 & n18793 ) | ( n18699 & n18797 ) | ( n18793 & n18797 ) ;
  assign n18799 = ( ~n18791 & n18796 ) | ( ~n18791 & n18798 ) | ( n18796 & n18798 ) ;
  assign n18800 = n5658 & n8357 ;
  assign n18801 = x43 & x55 ;
  assign n18802 = x44 & x54 ;
  assign n18803 = n18801 | n18802 ;
  assign n18804 = ~n18800 & n18803 ;
  assign n18805 = x35 & x63 ;
  assign n18806 = n18804 | n18805 ;
  assign n18807 = n18804 & n18805 ;
  assign n18808 = n18806 & ~n18807 ;
  assign n18809 = n18593 & n18808 ;
  assign n18810 = n18593 | n18808 ;
  assign n18811 = ~n18809 & n18810 ;
  assign n18812 = x41 & x57 ;
  assign n18813 = x42 & x56 ;
  assign n18814 = n18812 | n18813 ;
  assign n18815 = n5710 & n8903 ;
  assign n18816 = x38 & x60 ;
  assign n18817 = ~n18815 & n18816 ;
  assign n18818 = n18814 | n18815 ;
  assign n18819 = ( n18815 & n18817 ) | ( n18815 & n18818 ) | ( n18817 & n18818 ) ;
  assign n18820 = n18814 & ~n18819 ;
  assign n18821 = ~n18814 & n18816 ;
  assign n18822 = ( n18816 & ~n18817 ) | ( n18816 & n18821 ) | ( ~n18817 & n18821 ) ;
  assign n18823 = n18820 | n18822 ;
  assign n18824 = ~n18811 & n18823 ;
  assign n18825 = n18811 & ~n18823 ;
  assign n18826 = n18824 | n18825 ;
  assign n18827 = n18573 | n18579 ;
  assign n18828 = ( n18579 & n18583 ) | ( n18579 & n18827 ) | ( n18583 & n18827 ) ;
  assign n18829 = n18826 & ~n18828 ;
  assign n18830 = n18826 & n18828 ;
  assign n18831 = n18618 | n18626 ;
  assign n18832 = ( n18626 & n18629 ) | ( n18626 & n18831 ) | ( n18629 & n18831 ) ;
  assign n18833 = n18828 | n18832 ;
  assign n18834 = ( ~n18830 & n18832 ) | ( ~n18830 & n18833 ) | ( n18832 & n18833 ) ;
  assign n18835 = n18829 | n18834 ;
  assign n18836 = ( n18828 & n18829 ) | ( n18828 & n18832 ) | ( n18829 & n18832 ) ;
  assign n18837 = ( ~n18826 & n18829 ) | ( ~n18826 & n18836 ) | ( n18829 & n18836 ) ;
  assign n18838 = n18835 & ~n18837 ;
  assign n18839 = n18437 | n18633 ;
  assign n18840 = n18633 | n18635 ;
  assign n18841 = ( n18636 & n18839 ) | ( n18636 & n18840 ) | ( n18839 & n18840 ) ;
  assign n18842 = n18838 & n18841 ;
  assign n18843 = n18838 | n18841 ;
  assign n18844 = ~n18842 & n18843 ;
  assign n18845 = n18799 & n18844 ;
  assign n18846 = n18799 | n18844 ;
  assign n18847 = ~n18845 & n18846 ;
  assign n18848 = n18640 | n18705 ;
  assign n18849 = ( n18705 & n18707 ) | ( n18705 & n18848 ) | ( n18707 & n18848 ) ;
  assign n18850 = ( n18720 & n18847 ) | ( n18720 & ~n18849 ) | ( n18847 & ~n18849 ) ;
  assign n18851 = ( ~n18847 & n18849 ) | ( ~n18847 & n18850 ) | ( n18849 & n18850 ) ;
  assign n18852 = ( ~n18720 & n18850 ) | ( ~n18720 & n18851 ) | ( n18850 & n18851 ) ;
  assign n18853 = n18847 & n18849 ;
  assign n18854 = n18847 | n18849 ;
  assign n18855 = n18853 | n18854 ;
  assign n18856 = ( n18719 & n18853 ) | ( n18719 & n18855 ) | ( n18853 & n18855 ) ;
  assign n18857 = ( n18717 & n18853 ) | ( n18717 & n18855 ) | ( n18853 & n18855 ) ;
  assign n18858 = ( n18564 & n18856 ) | ( n18564 & n18857 ) | ( n18856 & n18857 ) ;
  assign n18859 = n18791 | n18793 ;
  assign n18860 = n5813 & n9831 ;
  assign n18861 = x44 & x59 ;
  assign n18862 = n18320 & n18861 ;
  assign n18863 = n18860 | n18862 ;
  assign n18864 = x41 & x58 ;
  assign n18865 = n10431 & n18864 ;
  assign n18866 = x59 & n18865 ;
  assign n18867 = ( x59 & ~n18863 ) | ( x59 & n18866 ) | ( ~n18863 & n18866 ) ;
  assign n18868 = x40 & n18867 ;
  assign n18869 = n18863 | n18865 ;
  assign n18870 = n10431 | n18864 ;
  assign n18871 = x40 | n18870 ;
  assign n18872 = ( n18867 & n18870 ) | ( n18867 & n18871 ) | ( n18870 & n18871 ) ;
  assign n18873 = ( n18868 & ~n18869 ) | ( n18868 & n18872 ) | ( ~n18869 & n18872 ) ;
  assign n18874 = n5610 & n11935 ;
  assign n18875 = n5975 & n8355 ;
  assign n18876 = n18874 | n18875 ;
  assign n18877 = n6147 & n8161 ;
  assign n18878 = x54 & n18877 ;
  assign n18879 = ( x54 & ~n18876 ) | ( x54 & n18878 ) | ( ~n18876 & n18878 ) ;
  assign n18880 = x45 & n18879 ;
  assign n18881 = n18876 | n18877 ;
  assign n18882 = x46 & x53 ;
  assign n18883 = ( n10332 & ~n18877 ) | ( n10332 & n18882 ) | ( ~n18877 & n18882 ) ;
  assign n18884 = n10332 & n18882 ;
  assign n18885 = ( ~n18876 & n18883 ) | ( ~n18876 & n18884 ) | ( n18883 & n18884 ) ;
  assign n18886 = ~n18881 & n18885 ;
  assign n18887 = n18880 | n18886 ;
  assign n18888 = n18873 & n18887 ;
  assign n18889 = n18873 & ~n18888 ;
  assign n18890 = n18887 & ~n18888 ;
  assign n18891 = n18889 | n18890 ;
  assign n18892 = x42 & x57 ;
  assign n18893 = x43 & x56 ;
  assign n18894 = n18892 | n18893 ;
  assign n18895 = n5407 & n8903 ;
  assign n18896 = x48 & x51 ;
  assign n18897 = ~n18895 & n18896 ;
  assign n18898 = n18894 | n18895 ;
  assign n18899 = ( n18895 & n18897 ) | ( n18895 & n18898 ) | ( n18897 & n18898 ) ;
  assign n18900 = n18894 & ~n18899 ;
  assign n18901 = ~n18894 & n18896 ;
  assign n18902 = ( n18896 & ~n18897 ) | ( n18896 & n18901 ) | ( ~n18897 & n18901 ) ;
  assign n18903 = n18900 | n18902 ;
  assign n18904 = ~n18891 & n18903 ;
  assign n18905 = n18891 & ~n18903 ;
  assign n18906 = n18904 | n18905 ;
  assign n18907 = n18781 | n18782 ;
  assign n18908 = ( n18781 & n18783 ) | ( n18781 & n18907 ) | ( n18783 & n18907 ) ;
  assign n18909 = n18906 | n18908 ;
  assign n18910 = n18906 & n18908 ;
  assign n18911 = n18909 & ~n18910 ;
  assign n18912 = n18732 | n18773 ;
  assign n18913 = ( n18732 & n18735 ) | ( n18732 & n18912 ) | ( n18735 & n18912 ) ;
  assign n18914 = n18911 | n18913 ;
  assign n18915 = n18911 & n18913 ;
  assign n18916 = n18914 & ~n18915 ;
  assign n18917 = n18793 & n18916 ;
  assign n18918 = ( n18791 & n18916 ) | ( n18791 & n18917 ) | ( n18916 & n18917 ) ;
  assign n18919 = n18859 & ~n18918 ;
  assign n18920 = ~n18791 & n18916 ;
  assign n18921 = ~n18917 & n18920 ;
  assign n18922 = n18919 | n18921 ;
  assign n18929 = n18676 | n18726 ;
  assign n18930 = ( n18726 & n18727 ) | ( n18726 & n18929 ) | ( n18727 & n18929 ) ;
  assign n18923 = ( x50 & x62 ) | ( x50 & ~n6834 ) | ( x62 & ~n6834 ) ;
  assign n18924 = x37 | x62 ;
  assign n18925 = ( n6834 & ~n13403 ) | ( n6834 & n18924 ) | ( ~n13403 & n18924 ) ;
  assign n18926 = ( ~x37 & x50 ) | ( ~x37 & x62 ) | ( x50 & x62 ) ;
  assign n18927 = ( x37 & n6834 ) | ( x37 & ~n18926 ) | ( n6834 & ~n18926 ) ;
  assign n18928 = ( n18923 & ~n18925 ) | ( n18923 & n18927 ) | ( ~n18925 & n18927 ) ;
  assign n18931 = n18928 & n18930 ;
  assign n18932 = n18930 & ~n18931 ;
  assign n18934 = n18809 | n18823 ;
  assign n18935 = ( n18809 & n18811 ) | ( n18809 & n18934 ) | ( n18811 & n18934 ) ;
  assign n18933 = n18928 & ~n18930 ;
  assign n18936 = n18933 & n18935 ;
  assign n18937 = ( n18932 & n18935 ) | ( n18932 & n18936 ) | ( n18935 & n18936 ) ;
  assign n18938 = n18933 | n18935 ;
  assign n18939 = n18932 | n18938 ;
  assign n18940 = ~n18937 & n18939 ;
  assign n18941 = n18761 | n18764 ;
  assign n18942 = ( n18602 & n18761 ) | ( n18602 & n18941 ) | ( n18761 & n18941 ) ;
  assign n18943 = n18819 | n18942 ;
  assign n18944 = n18819 & n18942 ;
  assign n18945 = n18943 & ~n18944 ;
  assign n18946 = n9771 & n12770 ;
  assign n18947 = n3731 & n10856 ;
  assign n18948 = n18946 | n18947 ;
  assign n18949 = n5392 & n10367 ;
  assign n18950 = x63 & n18949 ;
  assign n18951 = ( x63 & ~n18948 ) | ( x63 & n18950 ) | ( ~n18948 & n18950 ) ;
  assign n18952 = x36 & n18951 ;
  assign n18953 = n18948 | n18949 ;
  assign n18954 = x38 & x61 ;
  assign n18955 = x39 & x60 ;
  assign n18956 = ( ~n18949 & n18954 ) | ( ~n18949 & n18955 ) | ( n18954 & n18955 ) ;
  assign n18957 = n18954 & n18955 ;
  assign n18958 = ( ~n18948 & n18956 ) | ( ~n18948 & n18957 ) | ( n18956 & n18957 ) ;
  assign n18959 = ~n18953 & n18958 ;
  assign n18960 = n18952 | n18959 ;
  assign n18961 = ~n18945 & n18960 ;
  assign n18962 = n18945 & ~n18960 ;
  assign n18963 = n18961 | n18962 ;
  assign n18964 = n18760 | n18768 ;
  assign n18965 = ~n18753 & n18755 ;
  assign n18966 = ( n18753 & n18754 ) | ( n18753 & n18965 ) | ( n18754 & n18965 ) ;
  assign n18967 = n18744 | n18966 ;
  assign n18968 = n18744 & n18966 ;
  assign n18969 = n18967 & ~n18968 ;
  assign n18970 = n18800 | n18805 ;
  assign n18971 = ( n18800 & n18804 ) | ( n18800 & n18970 ) | ( n18804 & n18970 ) ;
  assign n18972 = n18969 | n18971 ;
  assign n18973 = n18969 & n18971 ;
  assign n18974 = n18972 & ~n18973 ;
  assign n18975 = n18759 | n18767 ;
  assign n18976 = n18974 & n18975 ;
  assign n18977 = n18759 & n18974 ;
  assign n18978 = ( n18964 & n18976 ) | ( n18964 & n18977 ) | ( n18976 & n18977 ) ;
  assign n18979 = n18974 | n18975 ;
  assign n18980 = n18759 | n18974 ;
  assign n18981 = ( n18964 & n18979 ) | ( n18964 & n18980 ) | ( n18979 & n18980 ) ;
  assign n18982 = ~n18978 & n18981 ;
  assign n18983 = n18963 & ~n18982 ;
  assign n18984 = ~n18963 & n18982 ;
  assign n18985 = n18983 | n18984 ;
  assign n18986 = n18940 & n18985 ;
  assign n18987 = n18940 | n18985 ;
  assign n18988 = ~n18986 & n18987 ;
  assign n18989 = n18829 | n18830 ;
  assign n18990 = ( ~n18829 & n18836 ) | ( ~n18829 & n18989 ) | ( n18836 & n18989 ) ;
  assign n18991 = n18988 & n18990 ;
  assign n18992 = n18988 | n18990 ;
  assign n18993 = ~n18991 & n18992 ;
  assign n18994 = n18922 | n18993 ;
  assign n18995 = n18922 & ~n18993 ;
  assign n18996 = ( ~n18922 & n18994 ) | ( ~n18922 & n18995 ) | ( n18994 & n18995 ) ;
  assign n18997 = n18799 | n18842 ;
  assign n18998 = ( n18842 & n18844 ) | ( n18842 & n18997 ) | ( n18844 & n18997 ) ;
  assign n18999 = ( n18858 & n18996 ) | ( n18858 & ~n18998 ) | ( n18996 & ~n18998 ) ;
  assign n19000 = ( ~n18996 & n18998 ) | ( ~n18996 & n18999 ) | ( n18998 & n18999 ) ;
  assign n19001 = ( ~n18858 & n18999 ) | ( ~n18858 & n19000 ) | ( n18999 & n19000 ) ;
  assign n19015 = n18968 | n18971 ;
  assign n19016 = ( n18968 & n18969 ) | ( n18968 & n19015 ) | ( n18969 & n19015 ) ;
  assign n19002 = n6757 & n7874 ;
  assign n19003 = n6762 & n8161 ;
  assign n19004 = n19002 | n19003 ;
  assign n19005 = n6759 & n7567 ;
  assign n19006 = x53 & n19005 ;
  assign n19007 = ( x53 & ~n19004 ) | ( x53 & n19006 ) | ( ~n19004 & n19006 ) ;
  assign n19008 = x47 & n19007 ;
  assign n19009 = n19004 | n19005 ;
  assign n19010 = ( n10866 & n18737 ) | ( n10866 & ~n19005 ) | ( n18737 & ~n19005 ) ;
  assign n19011 = n10866 & n18737 ;
  assign n19012 = ( ~n19004 & n19010 ) | ( ~n19004 & n19011 ) | ( n19010 & n19011 ) ;
  assign n19013 = ~n19009 & n19012 ;
  assign n19014 = n19008 | n19013 ;
  assign n19017 = n19014 & n19016 ;
  assign n19018 = n19016 & ~n19017 ;
  assign n19020 = n18944 | n18960 ;
  assign n19021 = ( n18944 & n18945 ) | ( n18944 & n19020 ) | ( n18945 & n19020 ) ;
  assign n19019 = n19014 & ~n19016 ;
  assign n19022 = n19019 & n19021 ;
  assign n19023 = ( n19018 & n19021 ) | ( n19018 & n19022 ) | ( n19021 & n19022 ) ;
  assign n19024 = n19019 | n19021 ;
  assign n19025 = n19018 | n19024 ;
  assign n19026 = ~n19023 & n19025 ;
  assign n19027 = n18910 | n18913 ;
  assign n19028 = ( n18910 & n18911 ) | ( n18910 & n19027 ) | ( n18911 & n19027 ) ;
  assign n19029 = n19026 | n19028 ;
  assign n19030 = n19026 & n19028 ;
  assign n19031 = n19029 & ~n19030 ;
  assign n19032 = n18881 | n18953 ;
  assign n19033 = n18881 & n18953 ;
  assign n19034 = n19032 & ~n19033 ;
  assign n19035 = n18869 | n19034 ;
  assign n19036 = n18869 & n19034 ;
  assign n19037 = n19035 & ~n19036 ;
  assign n19038 = n18888 | n18903 ;
  assign n19039 = n19037 & n19038 ;
  assign n19040 = n18888 & n19037 ;
  assign n19041 = ( n18891 & n19039 ) | ( n18891 & n19040 ) | ( n19039 & n19040 ) ;
  assign n19042 = n19037 | n19038 ;
  assign n19043 = n18888 | n19037 ;
  assign n19044 = ( n18891 & n19042 ) | ( n18891 & n19043 ) | ( n19042 & n19043 ) ;
  assign n19045 = ~n19041 & n19044 ;
  assign n19046 = x50 & x62 ;
  assign n19047 = x37 & n19046 ;
  assign n19048 = n6834 & ~n19047 ;
  assign n19049 = x37 & x63 ;
  assign n19050 = n19047 & n19049 ;
  assign n19051 = ( n19048 & n19049 ) | ( n19048 & n19050 ) | ( n19049 & n19050 ) ;
  assign n19052 = n19047 | n19049 ;
  assign n19053 = n19048 | n19052 ;
  assign n19054 = ~n19051 & n19053 ;
  assign n19055 = n18899 | n19054 ;
  assign n19056 = n18899 & n19054 ;
  assign n19057 = n19055 & ~n19056 ;
  assign n19058 = n19045 & n19057 ;
  assign n19059 = n19045 | n19057 ;
  assign n19060 = ~n19058 & n19059 ;
  assign n19061 = n19031 & n19060 ;
  assign n19062 = n19031 | n19060 ;
  assign n19063 = ~n19061 & n19062 ;
  assign n19064 = n14923 & n18816 ;
  assign n19065 = n5392 & n10684 ;
  assign n19066 = n19064 | n19065 ;
  assign n19067 = n4555 & n10367 ;
  assign n19068 = n14066 & n19067 ;
  assign n19069 = ( n14066 & ~n19066 ) | ( n14066 & n19068 ) | ( ~n19066 & n19068 ) ;
  assign n19070 = n19066 | n19067 ;
  assign n19071 = x39 & x61 ;
  assign n19072 = ( n18386 & ~n19067 ) | ( n18386 & n19071 ) | ( ~n19067 & n19071 ) ;
  assign n19073 = n18386 & n19071 ;
  assign n19074 = ( ~n19066 & n19072 ) | ( ~n19066 & n19073 ) | ( n19072 & n19073 ) ;
  assign n19075 = ~n19070 & n19074 ;
  assign n19076 = n19069 | n19075 ;
  assign n19077 = n5104 & n12860 ;
  assign n19078 = n5658 & n8903 ;
  assign n19079 = n19077 | n19078 ;
  assign n19080 = n6093 & n10013 ;
  assign n19081 = n11160 & n19080 ;
  assign n19082 = ( n11160 & ~n19079 ) | ( n11160 & n19081 ) | ( ~n19079 & n19081 ) ;
  assign n19083 = n19079 | n19080 ;
  assign n19084 = ( n10428 & n17937 ) | ( n10428 & ~n19080 ) | ( n17937 & ~n19080 ) ;
  assign n19085 = n10428 & n17937 ;
  assign n19086 = ( ~n19079 & n19084 ) | ( ~n19079 & n19085 ) | ( n19084 & n19085 ) ;
  assign n19087 = ~n19083 & n19086 ;
  assign n19088 = n19082 | n19087 ;
  assign n19089 = n19076 & n19088 ;
  assign n19090 = n19076 & ~n19089 ;
  assign n19091 = n19088 & ~n19089 ;
  assign n19092 = n19090 | n19091 ;
  assign n19093 = x41 & x59 ;
  assign n19094 = x42 & x58 ;
  assign n19095 = n19093 | n19094 ;
  assign n19096 = n5710 & n9831 ;
  assign n19097 = n10315 & ~n19096 ;
  assign n19098 = n19095 | n19096 ;
  assign n19099 = ( n19096 & n19097 ) | ( n19096 & n19098 ) | ( n19097 & n19098 ) ;
  assign n19100 = n19095 & ~n19099 ;
  assign n19101 = n10315 & ~n19095 ;
  assign n19102 = ( n10315 & ~n19097 ) | ( n10315 & n19101 ) | ( ~n19097 & n19101 ) ;
  assign n19103 = n19100 | n19102 ;
  assign n19104 = ~n19092 & n19103 ;
  assign n19105 = n19092 & ~n19103 ;
  assign n19106 = n19104 | n19105 ;
  assign n19107 = n18931 | n18937 ;
  assign n19108 = n19106 | n19107 ;
  assign n19109 = n19106 & n19107 ;
  assign n19110 = n19108 & ~n19109 ;
  assign n19111 = n18963 | n18978 ;
  assign n19112 = ( n18978 & n18982 ) | ( n18978 & n19111 ) | ( n18982 & n19111 ) ;
  assign n19113 = n19110 & n19112 ;
  assign n19114 = n19110 | n19112 ;
  assign n19115 = ~n19113 & n19114 ;
  assign n19116 = n18986 & n19115 ;
  assign n19117 = ( n18991 & n19115 ) | ( n18991 & n19116 ) | ( n19115 & n19116 ) ;
  assign n19118 = n18986 | n19115 ;
  assign n19119 = n18991 | n19118 ;
  assign n19120 = ~n19117 & n19119 ;
  assign n19121 = n19063 & n19120 ;
  assign n19122 = n19063 | n19120 ;
  assign n19123 = ~n19121 & n19122 ;
  assign n19124 = ( n18859 & n18916 ) | ( n18859 & n18993 ) | ( n18916 & n18993 ) ;
  assign n19125 = n19123 & n19124 ;
  assign n19126 = n19123 | n19124 ;
  assign n19127 = ~n19125 & n19126 ;
  assign n19128 = n18996 & n18998 ;
  assign n19129 = n18996 | n18998 ;
  assign n19130 = n18855 & n19129 ;
  assign n19131 = n18853 & n19129 ;
  assign n19132 = ( n18719 & n19130 ) | ( n18719 & n19131 ) | ( n19130 & n19131 ) ;
  assign n19133 = n19128 | n19132 ;
  assign n19134 = n19128 | n19129 ;
  assign n19135 = ( n18857 & n19128 ) | ( n18857 & n19134 ) | ( n19128 & n19134 ) ;
  assign n19136 = ( n18564 & n19133 ) | ( n18564 & n19135 ) | ( n19133 & n19135 ) ;
  assign n19137 = n19127 | n19136 ;
  assign n19138 = n19126 & n19128 ;
  assign n19139 = ( n19126 & n19132 ) | ( n19126 & n19138 ) | ( n19132 & n19138 ) ;
  assign n19140 = n19126 & n19134 ;
  assign n19141 = ( n18857 & n19138 ) | ( n18857 & n19140 ) | ( n19138 & n19140 ) ;
  assign n19142 = ( n18564 & n19139 ) | ( n18564 & n19141 ) | ( n19139 & n19141 ) ;
  assign n19143 = ~n19125 & n19142 ;
  assign n19144 = n19137 & ~n19143 ;
  assign n19145 = n19125 | n19126 ;
  assign n19146 = ( n19125 & n19128 ) | ( n19125 & n19145 ) | ( n19128 & n19145 ) ;
  assign n19147 = ( n19132 & n19145 ) | ( n19132 & n19146 ) | ( n19145 & n19146 ) ;
  assign n19148 = n19125 | n19141 ;
  assign n19149 = ( n18564 & n19147 ) | ( n18564 & n19148 ) | ( n19147 & n19148 ) ;
  assign n19150 = n19117 | n19121 ;
  assign n19151 = n19026 | n19060 ;
  assign n19152 = ( n19028 & n19060 ) | ( n19028 & n19151 ) | ( n19060 & n19151 ) ;
  assign n19153 = ( n19030 & n19031 ) | ( n19030 & n19152 ) | ( n19031 & n19152 ) ;
  assign n19154 = n15336 & n16811 ;
  assign n19155 = n5407 & n9831 ;
  assign n19156 = n19154 | n19155 ;
  assign n19157 = n5104 & n8708 ;
  assign n19158 = x59 & n19157 ;
  assign n19159 = ( x59 & ~n19156 ) | ( x59 & n19158 ) | ( ~n19156 & n19158 ) ;
  assign n19160 = x42 & n19159 ;
  assign n19161 = n19156 | n19157 ;
  assign n19162 = x43 & x58 ;
  assign n19163 = x45 & x56 ;
  assign n19164 = ( ~n19157 & n19162 ) | ( ~n19157 & n19163 ) | ( n19162 & n19163 ) ;
  assign n19165 = n19162 & n19163 ;
  assign n19166 = ( ~n19156 & n19164 ) | ( ~n19156 & n19165 ) | ( n19164 & n19165 ) ;
  assign n19167 = ~n19161 & n19166 ;
  assign n19168 = n19160 | n19167 ;
  assign n19169 = x46 & x55 ;
  assign n19170 = x47 & x54 ;
  assign n19171 = n19169 | n19170 ;
  assign n19172 = n6147 & n8357 ;
  assign n19173 = n19171 | n19172 ;
  assign n19174 = x38 & x63 ;
  assign n19175 = ( ~n19172 & n19173 ) | ( ~n19172 & n19174 ) | ( n19173 & n19174 ) ;
  assign n19176 = ( n19172 & n19173 ) | ( n19172 & ~n19174 ) | ( n19173 & ~n19174 ) ;
  assign n19177 = ( ~n19173 & n19175 ) | ( ~n19173 & n19176 ) | ( n19175 & n19176 ) ;
  assign n19178 = n19168 & n19177 ;
  assign n19179 = n19168 & ~n19178 ;
  assign n19180 = n6759 & n8161 ;
  assign n19181 = x44 & x57 ;
  assign n19182 = n11437 & n19181 ;
  assign n19183 = n19180 | n19182 ;
  assign n19184 = n9499 & n13843 ;
  assign n19185 = n11437 & n19184 ;
  assign n19186 = ( n11437 & ~n19183 ) | ( n11437 & n19185 ) | ( ~n19183 & n19185 ) ;
  assign n19187 = n19183 | n19184 ;
  assign n19188 = x49 & x52 ;
  assign n19189 = ( n19181 & ~n19184 ) | ( n19181 & n19188 ) | ( ~n19184 & n19188 ) ;
  assign n19190 = n19181 & n19188 ;
  assign n19191 = ( ~n19183 & n19189 ) | ( ~n19183 & n19190 ) | ( n19189 & n19190 ) ;
  assign n19192 = ~n19187 & n19191 ;
  assign n19193 = n19186 | n19192 ;
  assign n19194 = ~n19168 & n19177 ;
  assign n19195 = n19193 & ~n19194 ;
  assign n19196 = ~n19179 & n19195 ;
  assign n19197 = ~n19193 & n19194 ;
  assign n19198 = ( n19179 & ~n19193 ) | ( n19179 & n19197 ) | ( ~n19193 & n19197 ) ;
  assign n19199 = n19196 | n19198 ;
  assign n19200 = n19017 | n19023 ;
  assign n19201 = n19199 | n19200 ;
  assign n19202 = n19199 & n19200 ;
  assign n19203 = n19201 & ~n19202 ;
  assign n19223 = n18899 | n19051 ;
  assign n19224 = ( n19051 & n19054 ) | ( n19051 & n19223 ) | ( n19054 & n19223 ) ;
  assign n19204 = n5813 & n10367 ;
  assign n19205 = x41 & x60 ;
  assign n19206 = x40 & x61 ;
  assign n19207 = n19205 | n19206 ;
  assign n19208 = ~n19204 & n19207 ;
  assign n19209 = n19009 & n19208 ;
  assign n19210 = n19009 & ~n19209 ;
  assign n19211 = ~n19009 & n19208 ;
  assign n19212 = n19210 | n19211 ;
  assign n19213 = x62 & n8433 ;
  assign n19214 = n7112 & n19213 ;
  assign n19215 = n7112 & ~n19213 ;
  assign n19216 = n19213 | n19215 ;
  assign n19217 = x39 & x62 ;
  assign n19218 = ( x51 & ~n19213 ) | ( x51 & n19217 ) | ( ~n19213 & n19217 ) ;
  assign n19219 = x51 & n19217 ;
  assign n19220 = ( ~n19215 & n19218 ) | ( ~n19215 & n19219 ) | ( n19218 & n19219 ) ;
  assign n19221 = ~n19216 & n19220 ;
  assign n19222 = n19214 | n19221 ;
  assign n19225 = ( n19212 & ~n19222 ) | ( n19212 & n19224 ) | ( ~n19222 & n19224 ) ;
  assign n19226 = ( ~n19212 & n19222 ) | ( ~n19212 & n19225 ) | ( n19222 & n19225 ) ;
  assign n19227 = ( ~n19224 & n19225 ) | ( ~n19224 & n19226 ) | ( n19225 & n19226 ) ;
  assign n19228 = n19203 & n19227 ;
  assign n19229 = n19203 | n19227 ;
  assign n19230 = ~n19228 & n19229 ;
  assign n19231 = n19152 & n19230 ;
  assign n19232 = n19030 & n19230 ;
  assign n19233 = ( n19031 & n19231 ) | ( n19031 & n19232 ) | ( n19231 & n19232 ) ;
  assign n19234 = n19153 & ~n19233 ;
  assign n19235 = ~n19152 & n19230 ;
  assign n19236 = ~n19030 & n19230 ;
  assign n19237 = ( ~n19031 & n19235 ) | ( ~n19031 & n19236 ) | ( n19235 & n19236 ) ;
  assign n19238 = n19234 | n19237 ;
  assign n19239 = n19070 | n19099 ;
  assign n19240 = n19070 & n19099 ;
  assign n19241 = n19239 & ~n19240 ;
  assign n19242 = n19083 | n19241 ;
  assign n19243 = n19083 & n19241 ;
  assign n19244 = n19242 & ~n19243 ;
  assign n19245 = n19089 | n19103 ;
  assign n19246 = n18869 | n19033 ;
  assign n19247 = ( n19033 & n19034 ) | ( n19033 & n19246 ) | ( n19034 & n19246 ) ;
  assign n19248 = n19245 & n19247 ;
  assign n19249 = n19089 & n19247 ;
  assign n19250 = ( n19092 & n19248 ) | ( n19092 & n19249 ) | ( n19248 & n19249 ) ;
  assign n19251 = n19245 | n19247 ;
  assign n19252 = n19089 | n19247 ;
  assign n19253 = ( n19092 & n19251 ) | ( n19092 & n19252 ) | ( n19251 & n19252 ) ;
  assign n19254 = ~n19250 & n19253 ;
  assign n19255 = n19244 & n19254 ;
  assign n19256 = n19244 | n19254 ;
  assign n19257 = ~n19255 & n19256 ;
  assign n19258 = n19109 | n19112 ;
  assign n19259 = ( n19109 & n19110 ) | ( n19109 & n19258 ) | ( n19110 & n19258 ) ;
  assign n19260 = n19041 | n19057 ;
  assign n19261 = ( n19041 & n19045 ) | ( n19041 & n19260 ) | ( n19045 & n19260 ) ;
  assign n19262 = n19259 & n19261 ;
  assign n19263 = n19259 & ~n19262 ;
  assign n19264 = n19257 & n19261 ;
  assign n19265 = ~n19259 & n19264 ;
  assign n19266 = ( n19257 & n19263 ) | ( n19257 & n19265 ) | ( n19263 & n19265 ) ;
  assign n19267 = ~n19257 & n19261 ;
  assign n19268 = ~n19259 & n19267 ;
  assign n19269 = ( ~n19257 & n19263 ) | ( ~n19257 & n19268 ) | ( n19263 & n19268 ) ;
  assign n19270 = ( n19257 & ~n19266 ) | ( n19257 & n19269 ) | ( ~n19266 & n19269 ) ;
  assign n19271 = n19238 | n19270 ;
  assign n19272 = n19238 & ~n19270 ;
  assign n19273 = ( ~n19238 & n19271 ) | ( ~n19238 & n19272 ) | ( n19271 & n19272 ) ;
  assign n19274 = ( n19149 & n19150 ) | ( n19149 & ~n19273 ) | ( n19150 & ~n19273 ) ;
  assign n19275 = ( ~n19150 & n19273 ) | ( ~n19150 & n19274 ) | ( n19273 & n19274 ) ;
  assign n19276 = ( ~n19149 & n19274 ) | ( ~n19149 & n19275 ) | ( n19274 & n19275 ) ;
  assign n19277 = n19157 & n19204 ;
  assign n19278 = ( n19156 & n19204 ) | ( n19156 & n19277 ) | ( n19204 & n19277 ) ;
  assign n19279 = ( n19161 & n19209 ) | ( n19161 & n19278 ) | ( n19209 & n19278 ) ;
  assign n19280 = n19157 | n19204 ;
  assign n19281 = n19156 | n19280 ;
  assign n19282 = n19209 | n19281 ;
  assign n19283 = ~n19279 & n19282 ;
  assign n19284 = n12770 & n15454 ;
  assign n19285 = n4350 & n10856 ;
  assign n19286 = n19284 | n19285 ;
  assign n19287 = n5710 & n10367 ;
  assign n19288 = x63 & n19287 ;
  assign n19289 = ( x63 & ~n19286 ) | ( x63 & n19288 ) | ( ~n19286 & n19288 ) ;
  assign n19290 = x39 & n19289 ;
  assign n19291 = n19286 | n19287 ;
  assign n19292 = x41 & x61 ;
  assign n19293 = x42 & x60 ;
  assign n19294 = ( ~n19287 & n19292 ) | ( ~n19287 & n19293 ) | ( n19292 & n19293 ) ;
  assign n19295 = n19292 & n19293 ;
  assign n19296 = ( ~n19286 & n19294 ) | ( ~n19286 & n19295 ) | ( n19294 & n19295 ) ;
  assign n19297 = ~n19291 & n19296 ;
  assign n19298 = n19290 | n19297 ;
  assign n19299 = n19283 & ~n19298 ;
  assign n19300 = n19283 | n19298 ;
  assign n19301 = ( ~n19283 & n19299 ) | ( ~n19283 & n19300 ) | ( n19299 & n19300 ) ;
  assign n19302 = n19212 & n19222 ;
  assign n19303 = n19212 & ~n19302 ;
  assign n19304 = n19222 & n19224 ;
  assign n19305 = ~n19212 & n19304 ;
  assign n19306 = n19302 | n19305 ;
  assign n19307 = n19222 | n19224 ;
  assign n19308 = ( n19212 & n19224 ) | ( n19212 & n19307 ) | ( n19224 & n19307 ) ;
  assign n19309 = ( n19303 & n19306 ) | ( n19303 & n19308 ) | ( n19306 & n19308 ) ;
  assign n19310 = n19301 | n19309 ;
  assign n19311 = n19301 & n19309 ;
  assign n19312 = n19310 & ~n19311 ;
  assign n19313 = x43 & x59 ;
  assign n19314 = x44 & x58 ;
  assign n19315 = n19313 | n19314 ;
  assign n19316 = n5658 & n9831 ;
  assign n19317 = n14923 & ~n19316 ;
  assign n19318 = n19315 | n19316 ;
  assign n19319 = ( n19316 & n19317 ) | ( n19316 & n19318 ) | ( n19317 & n19318 ) ;
  assign n19320 = n19315 & ~n19319 ;
  assign n19321 = n14923 & ~n19315 ;
  assign n19322 = ( n14923 & ~n19317 ) | ( n14923 & n19321 ) | ( ~n19317 & n19321 ) ;
  assign n19323 = n19320 | n19322 ;
  assign n19324 = n5610 & n12860 ;
  assign n19325 = n5975 & n8903 ;
  assign n19326 = n19324 | n19325 ;
  assign n19327 = n6147 & n10013 ;
  assign n19328 = x57 & n19327 ;
  assign n19329 = ( x57 & ~n19326 ) | ( x57 & n19328 ) | ( ~n19326 & n19328 ) ;
  assign n19330 = x45 & n19329 ;
  assign n19331 = n19326 | n19327 ;
  assign n19332 = x46 & x56 ;
  assign n19333 = x47 & x55 ;
  assign n19334 = ( ~n19327 & n19332 ) | ( ~n19327 & n19333 ) | ( n19332 & n19333 ) ;
  assign n19335 = n19332 & n19333 ;
  assign n19336 = ( ~n19326 & n19334 ) | ( ~n19326 & n19335 ) | ( n19334 & n19335 ) ;
  assign n19337 = ~n19331 & n19336 ;
  assign n19338 = n19330 | n19337 ;
  assign n19339 = n19323 & n19338 ;
  assign n19340 = n19323 & ~n19339 ;
  assign n19341 = n19338 & ~n19339 ;
  assign n19342 = n19340 | n19341 ;
  assign n19343 = n6345 & n11935 ;
  assign n19344 = n6759 & n8355 ;
  assign n19345 = n19343 | n19344 ;
  assign n19346 = n6834 & n8161 ;
  assign n19347 = x54 & n19346 ;
  assign n19348 = ( x54 & ~n19345 ) | ( x54 & n19347 ) | ( ~n19345 & n19347 ) ;
  assign n19349 = x48 & n19348 ;
  assign n19350 = x49 & x53 ;
  assign n19351 = n7565 | n19350 ;
  assign n19352 = ~n19346 & n19351 ;
  assign n19353 = ~n19345 & n19352 ;
  assign n19354 = n19349 | n19353 ;
  assign n19355 = ~n19342 & n19354 ;
  assign n19356 = n19342 & ~n19354 ;
  assign n19357 = n19355 | n19356 ;
  assign n19358 = n19312 & n19357 ;
  assign n19359 = n19312 | n19357 ;
  assign n19360 = ~n19358 & n19359 ;
  assign n19361 = ( n19261 & n19358 ) | ( n19261 & ~n19359 ) | ( n19358 & ~n19359 ) ;
  assign n19362 = n19358 & ~n19359 ;
  assign n19363 = ( n19259 & n19361 ) | ( n19259 & n19362 ) | ( n19361 & n19362 ) ;
  assign n19364 = n19262 & ~n19363 ;
  assign n19365 = ( n19266 & n19360 ) | ( n19266 & n19364 ) | ( n19360 & n19364 ) ;
  assign n19366 = n19262 | n19265 ;
  assign n19367 = n19257 | n19261 ;
  assign n19368 = ( n19257 & n19259 ) | ( n19257 & n19367 ) | ( n19259 & n19367 ) ;
  assign n19369 = ( n19263 & n19366 ) | ( n19263 & n19368 ) | ( n19366 & n19368 ) ;
  assign n19370 = ~n19360 & n19369 ;
  assign n19371 = ( n19360 & ~n19365 ) | ( n19360 & n19370 ) | ( ~n19365 & n19370 ) ;
  assign n19372 = ~n19172 & n19174 ;
  assign n19373 = ( n19172 & n19173 ) | ( n19172 & n19372 ) | ( n19173 & n19372 ) ;
  assign n19374 = n19187 | n19216 ;
  assign n19375 = n19187 & n19216 ;
  assign n19376 = n19374 & ~n19375 ;
  assign n19377 = n19373 | n19376 ;
  assign n19378 = n19373 & n19376 ;
  assign n19379 = n19377 & ~n19378 ;
  assign n19380 = n19083 | n19240 ;
  assign n19381 = ( n19240 & n19241 ) | ( n19240 & n19380 ) | ( n19241 & n19380 ) ;
  assign n19382 = n19379 | n19381 ;
  assign n19383 = n19379 & n19381 ;
  assign n19384 = n19382 & ~n19383 ;
  assign n19385 = n19193 & n19194 ;
  assign n19386 = ( n19179 & n19193 ) | ( n19179 & n19385 ) | ( n19193 & n19385 ) ;
  assign n19387 = n19178 | n19386 ;
  assign n19388 = n19384 | n19387 ;
  assign n19389 = n19384 & n19387 ;
  assign n19390 = n19388 & ~n19389 ;
  assign n19391 = n19199 | n19227 ;
  assign n19392 = ( n19200 & n19227 ) | ( n19200 & n19391 ) | ( n19227 & n19391 ) ;
  assign n19393 = ( n19202 & n19203 ) | ( n19202 & n19392 ) | ( n19203 & n19392 ) ;
  assign n19394 = n19244 | n19250 ;
  assign n19395 = ( n19250 & n19254 ) | ( n19250 & n19394 ) | ( n19254 & n19394 ) ;
  assign n19396 = n19392 & n19395 ;
  assign n19397 = n19202 & n19395 ;
  assign n19398 = ( n19203 & n19396 ) | ( n19203 & n19397 ) | ( n19396 & n19397 ) ;
  assign n19399 = n19393 & ~n19398 ;
  assign n19400 = n19390 & n19395 ;
  assign n19401 = ~n19393 & n19400 ;
  assign n19402 = ( n19390 & n19399 ) | ( n19390 & n19401 ) | ( n19399 & n19401 ) ;
  assign n19403 = n19390 | n19395 ;
  assign n19404 = ( n19390 & ~n19393 ) | ( n19390 & n19403 ) | ( ~n19393 & n19403 ) ;
  assign n19405 = n19399 | n19404 ;
  assign n19406 = ~n19402 & n19405 ;
  assign n19407 = n19371 & n19406 ;
  assign n19408 = n19371 & ~n19407 ;
  assign n19409 = ~n19237 & n19270 ;
  assign n19410 = ( n19233 & n19234 ) | ( n19233 & n19270 ) | ( n19234 & n19270 ) ;
  assign n19411 = n19233 | n19270 ;
  assign n19412 = ( ~n19409 & n19410 ) | ( ~n19409 & n19411 ) | ( n19410 & n19411 ) ;
  assign n19413 = n19407 & ~n19412 ;
  assign n19414 = n19406 | n19412 ;
  assign n19415 = ( n19408 & ~n19413 ) | ( n19408 & n19414 ) | ( ~n19413 & n19414 ) ;
  assign n19416 = ~n19407 & n19412 ;
  assign n19417 = n19406 & n19412 ;
  assign n19418 = ( n19408 & n19416 ) | ( n19408 & n19417 ) | ( n19416 & n19417 ) ;
  assign n19419 = n19415 & ~n19418 ;
  assign n19420 = n19150 & n19273 ;
  assign n19421 = n19150 | n19273 ;
  assign n19422 = n19420 | n19421 ;
  assign n19423 = ( n19148 & n19420 ) | ( n19148 & n19422 ) | ( n19420 & n19422 ) ;
  assign n19424 = n19145 & n19421 ;
  assign n19425 = n19420 | n19424 ;
  assign n19426 = ( n19146 & n19420 ) | ( n19146 & n19422 ) | ( n19420 & n19422 ) ;
  assign n19427 = ( n19132 & n19425 ) | ( n19132 & n19426 ) | ( n19425 & n19426 ) ;
  assign n19428 = ( n18564 & n19423 ) | ( n18564 & n19427 ) | ( n19423 & n19427 ) ;
  assign n19429 = n19419 | n19428 ;
  assign n19430 = n19415 & n19427 ;
  assign n19431 = n19415 & n19422 ;
  assign n19432 = n19415 & n19420 ;
  assign n19433 = ( n19125 & n19431 ) | ( n19125 & n19432 ) | ( n19431 & n19432 ) ;
  assign n19434 = n19431 | n19432 ;
  assign n19435 = ( n19141 & n19433 ) | ( n19141 & n19434 ) | ( n19433 & n19434 ) ;
  assign n19436 = ( n18564 & n19430 ) | ( n18564 & n19435 ) | ( n19430 & n19435 ) ;
  assign n19437 = ~n19418 & n19436 ;
  assign n19438 = n19429 & ~n19437 ;
  assign n19550 = n19365 | n19406 ;
  assign n19551 = ( n19365 & n19371 ) | ( n19365 & n19550 ) | ( n19371 & n19550 ) ;
  assign n19439 = n6345 & n8360 ;
  assign n19440 = n6759 & n8357 ;
  assign n19441 = n19439 | n19440 ;
  assign n19442 = n6834 & n8355 ;
  assign n19443 = x55 & n19442 ;
  assign n19444 = ( x55 & ~n19441 ) | ( x55 & n19443 ) | ( ~n19441 & n19443 ) ;
  assign n19445 = x48 & n19444 ;
  assign n19446 = n19441 | n19442 ;
  assign n19447 = x50 & x53 ;
  assign n19448 = ( n13382 & ~n19442 ) | ( n13382 & n19447 ) | ( ~n19442 & n19447 ) ;
  assign n19449 = n13382 & n19447 ;
  assign n19450 = ( ~n19441 & n19448 ) | ( ~n19441 & n19449 ) | ( n19448 & n19449 ) ;
  assign n19451 = ~n19446 & n19450 ;
  assign n19452 = n19445 | n19451 ;
  assign n19453 = x46 & x57 ;
  assign n19454 = x47 & x56 ;
  assign n19455 = n19453 | n19454 ;
  assign n19456 = n6147 & n8903 ;
  assign n19457 = n19455 | n19456 ;
  assign n19458 = x43 & x60 ;
  assign n19459 = ( ~n19456 & n19457 ) | ( ~n19456 & n19458 ) | ( n19457 & n19458 ) ;
  assign n19460 = ( n19456 & n19457 ) | ( n19456 & ~n19458 ) | ( n19457 & ~n19458 ) ;
  assign n19461 = ( ~n19457 & n19459 ) | ( ~n19457 & n19460 ) | ( n19459 & n19460 ) ;
  assign n19462 = n19452 & n19461 ;
  assign n19463 = n19452 & ~n19462 ;
  assign n19464 = x52 & n15744 ;
  assign n19465 = n7567 & n19464 ;
  assign n19466 = ( x52 & ~n7567 ) | ( x52 & n15744 ) | ( ~n7567 & n15744 ) ;
  assign n19467 = x52 | n15744 ;
  assign n19468 = ( n19464 & n19466 ) | ( n19464 & n19467 ) | ( n19466 & n19467 ) ;
  assign n19469 = ( ~n19464 & n19465 ) | ( ~n19464 & n19468 ) | ( n19465 & n19468 ) ;
  assign n19470 = ~n19461 & n19469 ;
  assign n19471 = ( n19452 & n19469 ) | ( n19452 & n19470 ) | ( n19469 & n19470 ) ;
  assign n19472 = ~n19463 & n19471 ;
  assign n19473 = n19461 & ~n19469 ;
  assign n19474 = ~n19452 & n19473 ;
  assign n19475 = ( n19463 & ~n19469 ) | ( n19463 & n19474 ) | ( ~n19469 & n19474 ) ;
  assign n19476 = n19472 | n19475 ;
  assign n19477 = x40 & x63 ;
  assign n19478 = n19346 & n19477 ;
  assign n19479 = ( n19345 & n19477 ) | ( n19345 & n19478 ) | ( n19477 & n19478 ) ;
  assign n19480 = n19346 | n19477 ;
  assign n19481 = n19345 | n19480 ;
  assign n19482 = ~n19479 & n19481 ;
  assign n19483 = n19331 | n19482 ;
  assign n19484 = n19331 & n19482 ;
  assign n19485 = n19483 & ~n19484 ;
  assign n19486 = n19291 | n19319 ;
  assign n19487 = n19291 & n19319 ;
  assign n19488 = n19486 & ~n19487 ;
  assign n19489 = n4969 & n9737 ;
  assign n19490 = x45 & x61 ;
  assign n19491 = n19094 & n19490 ;
  assign n19492 = n19489 | n19491 ;
  assign n19493 = n6093 & n9831 ;
  assign n19494 = x61 & n19493 ;
  assign n19495 = ( x61 & ~n19492 ) | ( x61 & n19494 ) | ( ~n19492 & n19494 ) ;
  assign n19496 = x42 & n19495 ;
  assign n19497 = n19492 | n19493 ;
  assign n19498 = x45 & x58 ;
  assign n19499 = ( n18861 & ~n19493 ) | ( n18861 & n19498 ) | ( ~n19493 & n19498 ) ;
  assign n19500 = n18861 & n19498 ;
  assign n19501 = ( ~n19492 & n19499 ) | ( ~n19492 & n19500 ) | ( n19499 & n19500 ) ;
  assign n19502 = ~n19497 & n19501 ;
  assign n19503 = n19496 | n19502 ;
  assign n19504 = n19488 & n19503 ;
  assign n19505 = n19488 & ~n19504 ;
  assign n19506 = n19503 & ~n19504 ;
  assign n19507 = n19505 | n19506 ;
  assign n19508 = n19485 | n19507 ;
  assign n19509 = n19485 & n19507 ;
  assign n19510 = n19508 & ~n19509 ;
  assign n19511 = ~n19476 & n19510 ;
  assign n19512 = n19476 & ~n19510 ;
  assign n19513 = n19511 | n19512 ;
  assign n19514 = n19395 & n19513 ;
  assign n19515 = n19393 & n19514 ;
  assign n19516 = ( n19401 & n19513 ) | ( n19401 & n19515 ) | ( n19513 & n19515 ) ;
  assign n19517 = ( n19390 & n19513 ) | ( n19390 & n19515 ) | ( n19513 & n19515 ) ;
  assign n19518 = ( n19399 & n19516 ) | ( n19399 & n19517 ) | ( n19516 & n19517 ) ;
  assign n19519 = ( n19390 & n19392 ) | ( n19390 & n19395 ) | ( n19392 & n19395 ) ;
  assign n19520 = ( n19202 & n19390 ) | ( n19202 & n19395 ) | ( n19390 & n19395 ) ;
  assign n19521 = ( n19203 & n19519 ) | ( n19203 & n19520 ) | ( n19519 & n19520 ) ;
  assign n19522 = ~n19518 & n19521 ;
  assign n19523 = n19279 | n19298 ;
  assign n19524 = ( n19279 & n19283 ) | ( n19279 & n19523 ) | ( n19283 & n19523 ) ;
  assign n19525 = n19373 | n19375 ;
  assign n19526 = ( n19375 & n19376 ) | ( n19375 & n19525 ) | ( n19376 & n19525 ) ;
  assign n19527 = n19524 | n19526 ;
  assign n19528 = n19524 & n19526 ;
  assign n19529 = n19527 & ~n19528 ;
  assign n19530 = n19339 | n19354 ;
  assign n19531 = ( n19339 & n19342 ) | ( n19339 & n19530 ) | ( n19342 & n19530 ) ;
  assign n19532 = n19529 | n19531 ;
  assign n19533 = n19529 & n19531 ;
  assign n19534 = n19532 & ~n19533 ;
  assign n19535 = n19383 | n19389 ;
  assign n19536 = n19311 | n19357 ;
  assign n19537 = ( n19311 & n19312 ) | ( n19311 & n19536 ) | ( n19312 & n19536 ) ;
  assign n19538 = n19535 & n19537 ;
  assign n19539 = n19535 | n19537 ;
  assign n19540 = ~n19538 & n19539 ;
  assign n19541 = n19534 & n19540 ;
  assign n19542 = n19534 | n19540 ;
  assign n19543 = ~n19541 & n19542 ;
  assign n19544 = ~n19395 & n19513 ;
  assign n19545 = ( ~n19393 & n19513 ) | ( ~n19393 & n19544 ) | ( n19513 & n19544 ) ;
  assign n19546 = n19543 & n19545 ;
  assign n19547 = n19402 & n19543 ;
  assign n19548 = ( n19543 & ~n19546 ) | ( n19543 & n19547 ) | ( ~n19546 & n19547 ) ;
  assign n19549 = ~n19522 & n19548 ;
  assign n19552 = n19549 & n19551 ;
  assign n19553 = ~n19521 & n19545 ;
  assign n19554 = ~n19402 & n19553 ;
  assign n19555 = ~n19402 & n19545 ;
  assign n19556 = ( n19518 & n19554 ) | ( n19518 & n19555 ) | ( n19554 & n19555 ) ;
  assign n19557 = ( n19522 & ~n19543 ) | ( n19522 & n19556 ) | ( ~n19543 & n19556 ) ;
  assign n19558 = ( n19551 & n19552 ) | ( n19551 & n19557 ) | ( n19552 & n19557 ) ;
  assign n19559 = n19549 | n19551 ;
  assign n19560 = n19557 | n19559 ;
  assign n19561 = ~n19558 & n19560 ;
  assign n19562 = n19415 | n19418 ;
  assign n19563 = ( n19418 & n19427 ) | ( n19418 & n19562 ) | ( n19427 & n19562 ) ;
  assign n19564 = n19418 | n19435 ;
  assign n19565 = ( n18564 & n19563 ) | ( n18564 & n19564 ) | ( n19563 & n19564 ) ;
  assign n19566 = ~n19561 & n19565 ;
  assign n19567 = n19561 & ~n19565 ;
  assign n19568 = n19566 | n19567 ;
  assign n19569 = n19558 | n19560 ;
  assign n19570 = ( n19418 & n19558 ) | ( n19418 & n19569 ) | ( n19558 & n19569 ) ;
  assign n19571 = ( n19558 & n19562 ) | ( n19558 & n19569 ) | ( n19562 & n19569 ) ;
  assign n19572 = ( n19427 & n19570 ) | ( n19427 & n19571 ) | ( n19570 & n19571 ) ;
  assign n19573 = ( n19558 & n19564 ) | ( n19558 & n19569 ) | ( n19564 & n19569 ) ;
  assign n19574 = ( n18564 & n19572 ) | ( n18564 & n19573 ) | ( n19572 & n19573 ) ;
  assign n19575 = n19534 | n19535 ;
  assign n19576 = ( n19534 & n19537 ) | ( n19534 & n19575 ) | ( n19537 & n19575 ) ;
  assign n19577 = ( n19538 & n19540 ) | ( n19538 & n19576 ) | ( n19540 & n19576 ) ;
  assign n19578 = ~n19456 & n19458 ;
  assign n19579 = ( n19456 & n19457 ) | ( n19456 & n19578 ) | ( n19457 & n19578 ) ;
  assign n19580 = n19446 | n19579 ;
  assign n19581 = n19446 & n19579 ;
  assign n19582 = n19580 & ~n19581 ;
  assign n19583 = n19497 | n19582 ;
  assign n19584 = n19497 & n19582 ;
  assign n19585 = n19583 & ~n19584 ;
  assign n19586 = ~n19452 & n19461 ;
  assign n19587 = n19461 | n19469 ;
  assign n19588 = ( n19452 & n19469 ) | ( n19452 & n19587 ) | ( n19469 & n19587 ) ;
  assign n19589 = ( n19462 & n19586 ) | ( n19462 & n19588 ) | ( n19586 & n19588 ) ;
  assign n19590 = n19462 | n19588 ;
  assign n19591 = ( n19463 & n19589 ) | ( n19463 & n19590 ) | ( n19589 & n19590 ) ;
  assign n19592 = n19585 & n19591 ;
  assign n19593 = n19585 | n19591 ;
  assign n19594 = ~n19592 & n19593 ;
  assign n19595 = n5658 & n10367 ;
  assign n19596 = n6093 & n10370 ;
  assign n19597 = n19595 | n19596 ;
  assign n19598 = n5104 & n9737 ;
  assign n19599 = x60 & n19598 ;
  assign n19600 = ( x60 & ~n19597 ) | ( x60 & n19599 ) | ( ~n19597 & n19599 ) ;
  assign n19601 = x44 & n19600 ;
  assign n19602 = n19597 | n19598 ;
  assign n19603 = x43 & x61 ;
  assign n19604 = x45 & x59 ;
  assign n19605 = ( ~n19598 & n19603 ) | ( ~n19598 & n19604 ) | ( n19603 & n19604 ) ;
  assign n19606 = n19603 & n19604 ;
  assign n19607 = ( ~n19597 & n19605 ) | ( ~n19597 & n19606 ) | ( n19605 & n19606 ) ;
  assign n19608 = ~n19602 & n19607 ;
  assign n19609 = n19601 | n19608 ;
  assign n19610 = n6147 & n9272 ;
  assign n19611 = x48 & x58 ;
  assign n19612 = n19332 & n19611 ;
  assign n19613 = n19610 | n19612 ;
  assign n19614 = n6762 & n8903 ;
  assign n19615 = x58 & n19614 ;
  assign n19616 = ( x58 & ~n19613 ) | ( x58 & n19615 ) | ( ~n19613 & n19615 ) ;
  assign n19617 = x46 & n19616 ;
  assign n19618 = n19613 | n19614 ;
  assign n19619 = x47 & x57 ;
  assign n19620 = ( n10718 & ~n19614 ) | ( n10718 & n19619 ) | ( ~n19614 & n19619 ) ;
  assign n19621 = n10718 & n19619 ;
  assign n19622 = ( ~n19613 & n19620 ) | ( ~n19613 & n19621 ) | ( n19620 & n19621 ) ;
  assign n19623 = ~n19618 & n19622 ;
  assign n19624 = n19617 | n19623 ;
  assign n19625 = n19609 & n19624 ;
  assign n19626 = n19609 & ~n19625 ;
  assign n19627 = n19624 & ~n19625 ;
  assign n19628 = n19626 | n19627 ;
  assign n19629 = n7874 & n10573 ;
  assign n19630 = n6834 & n8357 ;
  assign n19631 = n19629 | n19630 ;
  assign n19632 = n7112 & n8355 ;
  assign n19633 = n10573 & n19632 ;
  assign n19634 = ( n10573 & ~n19631 ) | ( n10573 & n19633 ) | ( ~n19631 & n19633 ) ;
  assign n19635 = n19631 | n19632 ;
  assign n19636 = x50 & x54 ;
  assign n19637 = ( n7874 & ~n19632 ) | ( n7874 & n19636 ) | ( ~n19632 & n19636 ) ;
  assign n19638 = n7874 & n19636 ;
  assign n19639 = ( ~n19631 & n19637 ) | ( ~n19631 & n19638 ) | ( n19637 & n19638 ) ;
  assign n19640 = ~n19635 & n19639 ;
  assign n19641 = n19634 | n19640 ;
  assign n19642 = ~n19628 & n19641 ;
  assign n19643 = n19628 & ~n19641 ;
  assign n19644 = n19642 | n19643 ;
  assign n19645 = n19594 & n19644 ;
  assign n19646 = n19594 | n19644 ;
  assign n19647 = ~n19645 & n19646 ;
  assign n19648 = n19576 & n19647 ;
  assign n19649 = n19538 & n19647 ;
  assign n19650 = ( n19540 & n19648 ) | ( n19540 & n19649 ) | ( n19648 & n19649 ) ;
  assign n19651 = n19577 & ~n19650 ;
  assign n19652 = n19528 | n19533 ;
  assign n19653 = n19476 | n19509 ;
  assign n19654 = ( n19509 & n19510 ) | ( n19509 & n19653 ) | ( n19510 & n19653 ) ;
  assign n19655 = n19652 | n19654 ;
  assign n19656 = n19652 & n19654 ;
  assign n19657 = n19655 & ~n19656 ;
  assign n19658 = n7567 & ~n19464 ;
  assign n19659 = n19464 | n19658 ;
  assign n19660 = n5710 & n10561 ;
  assign n19661 = x41 & x63 ;
  assign n19662 = n15832 | n19661 ;
  assign n19663 = ~n19660 & n19662 ;
  assign n19664 = n19659 & n19663 ;
  assign n19665 = n19659 | n19663 ;
  assign n19666 = ~n19664 & n19665 ;
  assign n19667 = n19331 | n19479 ;
  assign n19668 = ( n19479 & n19482 ) | ( n19479 & n19667 ) | ( n19482 & n19667 ) ;
  assign n19669 = n19666 | n19668 ;
  assign n19670 = n19666 & n19668 ;
  assign n19671 = n19669 & ~n19670 ;
  assign n19672 = n19487 | n19504 ;
  assign n19673 = n19671 | n19672 ;
  assign n19674 = n19671 & n19672 ;
  assign n19675 = n19673 & ~n19674 ;
  assign n19676 = n19657 & n19675 ;
  assign n19677 = n19657 | n19675 ;
  assign n19678 = ~n19676 & n19677 ;
  assign n19679 = ~n19576 & n19647 ;
  assign n19680 = ~n19538 & n19647 ;
  assign n19681 = ( ~n19540 & n19679 ) | ( ~n19540 & n19680 ) | ( n19679 & n19680 ) ;
  assign n19682 = n19678 & n19681 ;
  assign n19683 = ( n19651 & n19678 ) | ( n19651 & n19682 ) | ( n19678 & n19682 ) ;
  assign n19684 = n19678 | n19681 ;
  assign n19685 = n19651 | n19684 ;
  assign n19686 = ~n19683 & n19685 ;
  assign n19687 = n19518 | n19522 ;
  assign n19688 = n19518 | n19543 ;
  assign n19689 = n19543 & n19555 ;
  assign n19690 = ( n19687 & n19688 ) | ( n19687 & n19689 ) | ( n19688 & n19689 ) ;
  assign n19691 = ( n19574 & n19686 ) | ( n19574 & ~n19690 ) | ( n19686 & ~n19690 ) ;
  assign n19692 = ( ~n19686 & n19690 ) | ( ~n19686 & n19691 ) | ( n19690 & n19691 ) ;
  assign n19693 = ( ~n19574 & n19691 ) | ( ~n19574 & n19692 ) | ( n19691 & n19692 ) ;
  assign n19694 = n19686 & n19690 ;
  assign n19695 = n19686 | n19690 ;
  assign n19696 = n19694 | n19695 ;
  assign n19697 = ( n19572 & n19694 ) | ( n19572 & n19696 ) | ( n19694 & n19696 ) ;
  assign n19698 = ( n19569 & n19694 ) | ( n19569 & n19696 ) | ( n19694 & n19696 ) ;
  assign n19699 = ( n19558 & n19694 ) | ( n19558 & n19696 ) | ( n19694 & n19696 ) ;
  assign n19700 = ( n19418 & n19698 ) | ( n19418 & n19699 ) | ( n19698 & n19699 ) ;
  assign n19701 = n19698 | n19699 ;
  assign n19702 = ( n19435 & n19700 ) | ( n19435 & n19701 ) | ( n19700 & n19701 ) ;
  assign n19703 = ( n18564 & n19697 ) | ( n18564 & n19702 ) | ( n19697 & n19702 ) ;
  assign n19704 = n19618 | n19635 ;
  assign n19705 = n19618 & n19635 ;
  assign n19706 = n19704 & ~n19705 ;
  assign n19707 = n19602 | n19706 ;
  assign n19708 = n19602 & n19706 ;
  assign n19709 = n19707 & ~n19708 ;
  assign n19710 = n19625 | n19641 ;
  assign n19711 = n19709 & n19710 ;
  assign n19712 = n19625 & n19709 ;
  assign n19713 = ( n19628 & n19711 ) | ( n19628 & n19712 ) | ( n19711 & n19712 ) ;
  assign n19714 = n19709 | n19710 ;
  assign n19715 = n19625 | n19709 ;
  assign n19716 = ( n19628 & n19714 ) | ( n19628 & n19715 ) | ( n19714 & n19715 ) ;
  assign n19717 = ~n19713 & n19716 ;
  assign n19718 = n19670 | n19674 ;
  assign n19719 = n19717 | n19718 ;
  assign n19720 = n19717 & n19718 ;
  assign n19721 = n19719 & ~n19720 ;
  assign n19722 = n19656 | n19675 ;
  assign n19723 = ( n19656 & n19657 ) | ( n19656 & n19722 ) | ( n19657 & n19722 ) ;
  assign n19724 = n19721 & n19723 ;
  assign n19725 = n19721 | n19723 ;
  assign n19726 = ~n19724 & n19725 ;
  assign n19727 = n8146 & n10866 ;
  assign n19728 = n6834 & n10013 ;
  assign n19729 = n19727 | n19728 ;
  assign n19730 = n7112 & n8357 ;
  assign n19731 = x56 & n19730 ;
  assign n19732 = ( x56 & ~n19729 ) | ( x56 & n19731 ) | ( ~n19729 & n19731 ) ;
  assign n19733 = x49 & n19732 ;
  assign n19734 = n19729 | n19730 ;
  assign n19735 = x51 & x54 ;
  assign n19736 = x50 & x55 ;
  assign n19737 = ( ~n19730 & n19735 ) | ( ~n19730 & n19736 ) | ( n19735 & n19736 ) ;
  assign n19738 = n19735 & n19736 ;
  assign n19739 = ( ~n19729 & n19737 ) | ( ~n19729 & n19738 ) | ( n19737 & n19738 ) ;
  assign n19740 = ~n19734 & n19739 ;
  assign n19741 = n19733 | n19740 ;
  assign n19742 = x62 & n18480 ;
  assign n19743 = n8161 & ~n19742 ;
  assign n19744 = x53 | n16442 ;
  assign n19745 = ~n19742 & n19744 ;
  assign n19746 = ~n19743 & n19745 ;
  assign n19747 = n8161 & n19742 ;
  assign n19748 = n19746 | n19747 ;
  assign n19749 = n19741 & n19748 ;
  assign n19750 = n19741 & ~n19749 ;
  assign n19752 = n19497 | n19581 ;
  assign n19753 = ( n19581 & n19582 ) | ( n19581 & n19752 ) | ( n19582 & n19752 ) ;
  assign n19751 = ~n19741 & n19748 ;
  assign n19754 = n19751 & n19753 ;
  assign n19755 = ( n19750 & n19753 ) | ( n19750 & n19754 ) | ( n19753 & n19754 ) ;
  assign n19756 = n19751 | n19753 ;
  assign n19757 = n19750 | n19756 ;
  assign n19758 = ~n19755 & n19757 ;
  assign n19759 = n12770 & n16811 ;
  assign n19760 = n4969 & n10856 ;
  assign n19761 = n19759 | n19760 ;
  assign n19762 = n6093 & n10367 ;
  assign n19763 = x42 & n19762 ;
  assign n19764 = ( x42 & ~n19761 ) | ( x42 & n19763 ) | ( ~n19761 & n19763 ) ;
  assign n19765 = x63 & n19764 ;
  assign n19766 = n19761 | n19762 ;
  assign n19767 = x44 & x61 ;
  assign n19768 = x45 & x60 ;
  assign n19769 = ( ~n19762 & n19767 ) | ( ~n19762 & n19768 ) | ( n19767 & n19768 ) ;
  assign n19770 = n19767 & n19768 ;
  assign n19771 = ( ~n19761 & n19769 ) | ( ~n19761 & n19770 ) | ( n19769 & n19770 ) ;
  assign n19772 = ~n19766 & n19771 ;
  assign n19773 = n19765 | n19772 ;
  assign n19774 = n19660 | n19663 ;
  assign n19775 = ( n19659 & n19660 ) | ( n19659 & n19774 ) | ( n19660 & n19774 ) ;
  assign n19776 = n19773 & ~n19775 ;
  assign n19777 = ~n19773 & n19775 ;
  assign n19778 = n19776 | n19777 ;
  assign n19779 = n9421 & n9829 ;
  assign n19780 = n6147 & n9831 ;
  assign n19781 = n19779 | n19780 ;
  assign n19782 = n6762 & n9272 ;
  assign n19783 = x59 & n19782 ;
  assign n19784 = ( x59 & ~n19781 ) | ( x59 & n19783 ) | ( ~n19781 & n19783 ) ;
  assign n19785 = x46 & n19784 ;
  assign n19786 = n19781 | n19782 ;
  assign n19787 = x47 & x58 ;
  assign n19788 = x48 & x57 ;
  assign n19789 = ( ~n19782 & n19787 ) | ( ~n19782 & n19788 ) | ( n19787 & n19788 ) ;
  assign n19790 = n19787 & n19788 ;
  assign n19791 = ( ~n19781 & n19789 ) | ( ~n19781 & n19790 ) | ( n19789 & n19790 ) ;
  assign n19792 = ~n19786 & n19791 ;
  assign n19793 = n19785 | n19792 ;
  assign n19794 = n19778 & n19793 ;
  assign n19795 = n19778 | n19793 ;
  assign n19796 = ~n19794 & n19795 ;
  assign n19797 = n19758 | n19796 ;
  assign n19798 = n19758 & n19796 ;
  assign n19799 = n19797 & ~n19798 ;
  assign n19800 = n19592 | n19645 ;
  assign n19801 = n19799 & n19800 ;
  assign n19802 = n19799 | n19800 ;
  assign n19803 = ~n19801 & n19802 ;
  assign n19804 = n19726 & n19803 ;
  assign n19805 = n19726 | n19803 ;
  assign n19806 = ~n19804 & n19805 ;
  assign n19807 = n19650 | n19683 ;
  assign n19808 = ( n19703 & n19806 ) | ( n19703 & ~n19807 ) | ( n19806 & ~n19807 ) ;
  assign n19809 = ( ~n19806 & n19807 ) | ( ~n19806 & n19808 ) | ( n19807 & n19808 ) ;
  assign n19810 = ( ~n19703 & n19808 ) | ( ~n19703 & n19809 ) | ( n19808 & n19809 ) ;
  assign n19811 = x43 & x63 ;
  assign n19812 = n19742 & n19811 ;
  assign n19813 = ( n19743 & n19811 ) | ( n19743 & n19812 ) | ( n19811 & n19812 ) ;
  assign n19814 = n19742 | n19811 ;
  assign n19815 = n19743 | n19814 ;
  assign n19816 = ~n19813 & n19815 ;
  assign n19817 = n19734 | n19816 ;
  assign n19818 = n19734 & n19816 ;
  assign n19819 = n19817 & ~n19818 ;
  assign n19820 = ( n19773 & n19775 ) | ( n19773 & n19793 ) | ( n19775 & n19793 ) ;
  assign n19821 = n19819 | n19820 ;
  assign n19822 = n19819 & n19820 ;
  assign n19823 = n19821 & ~n19822 ;
  assign n19824 = n19749 | n19755 ;
  assign n19825 = n19823 | n19824 ;
  assign n19826 = n19823 & n19824 ;
  assign n19827 = n19825 & ~n19826 ;
  assign n19828 = n19798 | n19799 ;
  assign n19829 = ( n19798 & n19800 ) | ( n19798 & n19828 ) | ( n19800 & n19828 ) ;
  assign n19830 = n19827 & n19829 ;
  assign n19831 = n19827 | n19829 ;
  assign n19832 = ~n19830 & n19831 ;
  assign n19888 = n19713 | n19718 ;
  assign n19889 = ( n19713 & n19717 ) | ( n19713 & n19888 ) | ( n19717 & n19888 ) ;
  assign n19833 = n6757 & n9829 ;
  assign n19834 = n6762 & n9831 ;
  assign n19835 = n19833 | n19834 ;
  assign n19836 = n6759 & n9272 ;
  assign n19837 = x59 & n19836 ;
  assign n19838 = ( x59 & ~n19835 ) | ( x59 & n19837 ) | ( ~n19835 & n19837 ) ;
  assign n19839 = x47 & n19838 ;
  assign n19840 = n19835 | n19836 ;
  assign n19841 = ( n13843 & n19611 ) | ( n13843 & ~n19836 ) | ( n19611 & ~n19836 ) ;
  assign n19842 = n13843 & n19611 ;
  assign n19843 = ( ~n19835 & n19841 ) | ( ~n19835 & n19842 ) | ( n19841 & n19842 ) ;
  assign n19844 = ~n19840 & n19843 ;
  assign n19845 = n19839 | n19844 ;
  assign n19846 = n7565 & n8146 ;
  assign n19847 = n7112 & n10013 ;
  assign n19848 = n19846 | n19847 ;
  assign n19849 = n7567 & n8357 ;
  assign n19850 = x56 & n19849 ;
  assign n19851 = ( x56 & ~n19848 ) | ( x56 & n19850 ) | ( ~n19848 & n19850 ) ;
  assign n19852 = x50 & n19851 ;
  assign n19853 = n19848 | n19849 ;
  assign n19854 = x51 & x55 ;
  assign n19855 = ( n11935 & ~n19849 ) | ( n11935 & n19854 ) | ( ~n19849 & n19854 ) ;
  assign n19856 = n11935 & n19854 ;
  assign n19857 = ( ~n19848 & n19855 ) | ( ~n19848 & n19856 ) | ( n19855 & n19856 ) ;
  assign n19858 = ~n19853 & n19857 ;
  assign n19859 = n19852 | n19858 ;
  assign n19860 = n19845 & n19859 ;
  assign n19861 = n19845 & ~n19860 ;
  assign n19862 = n19859 & ~n19860 ;
  assign n19863 = n19861 | n19862 ;
  assign n19864 = n19602 | n19705 ;
  assign n19865 = ( n19705 & n19706 ) | ( n19705 & n19864 ) | ( n19706 & n19864 ) ;
  assign n19866 = n19863 | n19865 ;
  assign n19867 = n19863 & n19865 ;
  assign n19868 = n19866 & ~n19867 ;
  assign n19869 = n19766 | n19786 ;
  assign n19870 = n19766 & n19786 ;
  assign n19871 = n19869 & ~n19870 ;
  assign n19872 = n6093 & n10684 ;
  assign n19873 = x46 & x60 ;
  assign n19874 = n17026 & n19873 ;
  assign n19875 = n19872 | n19874 ;
  assign n19876 = n5975 & n10367 ;
  assign n19877 = n17026 & n19876 ;
  assign n19878 = ( n17026 & ~n19875 ) | ( n17026 & n19877 ) | ( ~n19875 & n19877 ) ;
  assign n19879 = n19875 | n19876 ;
  assign n19880 = ( n19490 & n19873 ) | ( n19490 & ~n19876 ) | ( n19873 & ~n19876 ) ;
  assign n19881 = n19490 & n19873 ;
  assign n19882 = ( ~n19875 & n19880 ) | ( ~n19875 & n19881 ) | ( n19880 & n19881 ) ;
  assign n19883 = ~n19879 & n19882 ;
  assign n19884 = n19878 | n19883 ;
  assign n19885 = ~n19871 & n19884 ;
  assign n19886 = n19871 & ~n19884 ;
  assign n19887 = n19885 | n19886 ;
  assign n19890 = ( n19868 & ~n19887 ) | ( n19868 & n19889 ) | ( ~n19887 & n19889 ) ;
  assign n19891 = ( ~n19868 & n19887 ) | ( ~n19868 & n19889 ) | ( n19887 & n19889 ) ;
  assign n19892 = ( ~n19889 & n19890 ) | ( ~n19889 & n19891 ) | ( n19890 & n19891 ) ;
  assign n19893 = n19832 & ~n19892 ;
  assign n19894 = ~n19832 & n19892 ;
  assign n19895 = n19893 | n19894 ;
  assign n19896 = n19724 | n19803 ;
  assign n19897 = ( n19724 & n19726 ) | ( n19724 & n19896 ) | ( n19726 & n19896 ) ;
  assign n19898 = n19895 & n19897 ;
  assign n19899 = n19895 | n19897 ;
  assign n19900 = ~n19898 & n19899 ;
  assign n19901 = n19806 & n19807 ;
  assign n19902 = n19806 | n19807 ;
  assign n19903 = n19699 & n19902 ;
  assign n19904 = ( n19698 & n19902 ) | ( n19698 & n19903 ) | ( n19902 & n19903 ) ;
  assign n19905 = n19418 & n19902 ;
  assign n19906 = ( n19698 & n19903 ) | ( n19698 & n19905 ) | ( n19903 & n19905 ) ;
  assign n19907 = ( n19435 & n19904 ) | ( n19435 & n19906 ) | ( n19904 & n19906 ) ;
  assign n19908 = n19901 | n19907 ;
  assign n19909 = n19694 & n19902 ;
  assign n19910 = n19901 | n19909 ;
  assign n19911 = n19901 | n19902 ;
  assign n19912 = ( n19696 & n19901 ) | ( n19696 & n19911 ) | ( n19901 & n19911 ) ;
  assign n19913 = ( n19572 & n19910 ) | ( n19572 & n19912 ) | ( n19910 & n19912 ) ;
  assign n19914 = ( n18564 & n19908 ) | ( n18564 & n19913 ) | ( n19908 & n19913 ) ;
  assign n19915 = n19900 | n19914 ;
  assign n19916 = n19899 & n19901 ;
  assign n19917 = ( n19899 & n19907 ) | ( n19899 & n19916 ) | ( n19907 & n19916 ) ;
  assign n19918 = ( n19899 & n19909 ) | ( n19899 & n19916 ) | ( n19909 & n19916 ) ;
  assign n19919 = n19899 & n19911 ;
  assign n19920 = ( n19696 & n19916 ) | ( n19696 & n19919 ) | ( n19916 & n19919 ) ;
  assign n19921 = ( n19571 & n19918 ) | ( n19571 & n19920 ) | ( n19918 & n19920 ) ;
  assign n19922 = ( n19570 & n19918 ) | ( n19570 & n19920 ) | ( n19918 & n19920 ) ;
  assign n19923 = ( n19427 & n19921 ) | ( n19427 & n19922 ) | ( n19921 & n19922 ) ;
  assign n19924 = ( n18564 & n19917 ) | ( n18564 & n19923 ) | ( n19917 & n19923 ) ;
  assign n19925 = ~n19898 & n19924 ;
  assign n19926 = n19915 & ~n19925 ;
  assign n20015 = n19898 | n19920 ;
  assign n20016 = n19898 | n19918 ;
  assign n20017 = ( n19570 & n20015 ) | ( n19570 & n20016 ) | ( n20015 & n20016 ) ;
  assign n20018 = ( n19571 & n20015 ) | ( n19571 & n20016 ) | ( n20015 & n20016 ) ;
  assign n20019 = ( n19427 & n20017 ) | ( n19427 & n20018 ) | ( n20017 & n20018 ) ;
  assign n20020 = ( n19895 & n19897 ) | ( n19895 & n19901 ) | ( n19897 & n19901 ) ;
  assign n20021 = ( n19899 & n19906 ) | ( n19899 & n20020 ) | ( n19906 & n20020 ) ;
  assign n20022 = ( n19899 & n19904 ) | ( n19899 & n20020 ) | ( n19904 & n20020 ) ;
  assign n20023 = ( n19435 & n20021 ) | ( n19435 & n20022 ) | ( n20021 & n20022 ) ;
  assign n20024 = ( n18534 & n20019 ) | ( n18534 & n20023 ) | ( n20019 & n20023 ) ;
  assign n20025 = n20019 | n20023 ;
  assign n20026 = ( n18553 & n20024 ) | ( n18553 & n20025 ) | ( n20024 & n20025 ) ;
  assign n20027 = ( n18562 & n20019 ) | ( n18562 & n20023 ) | ( n20019 & n20023 ) ;
  assign n20028 = ( n18561 & n20019 ) | ( n18561 & n20023 ) | ( n20019 & n20023 ) ;
  assign n20029 = ( n17877 & n20027 ) | ( n17877 & n20028 ) | ( n20027 & n20028 ) ;
  assign n20030 = ( n17121 & n20026 ) | ( n17121 & n20029 ) | ( n20026 & n20029 ) ;
  assign n20031 = ( n17119 & n20026 ) | ( n17119 & n20029 ) | ( n20026 & n20029 ) ;
  assign n20032 = ( n13196 & n20030 ) | ( n13196 & n20031 ) | ( n20030 & n20031 ) ;
  assign n19927 = n19840 | n19879 ;
  assign n19928 = n19840 & n19879 ;
  assign n19929 = n19927 & ~n19928 ;
  assign n19930 = n6759 & n9831 ;
  assign n19931 = x59 & x63 ;
  assign n19932 = n17712 & n19931 ;
  assign n19933 = n19930 | n19932 ;
  assign n19934 = x58 & x63 ;
  assign n19935 = n9005 & n19934 ;
  assign n19936 = x59 & n19935 ;
  assign n19937 = ( x59 & ~n19933 ) | ( x59 & n19936 ) | ( ~n19933 & n19936 ) ;
  assign n19938 = x48 & n19937 ;
  assign n19939 = n19933 | n19935 ;
  assign n19940 = x44 & x63 ;
  assign n19941 = x49 & x58 ;
  assign n19942 = ( ~n19935 & n19940 ) | ( ~n19935 & n19941 ) | ( n19940 & n19941 ) ;
  assign n19943 = n19940 & n19941 ;
  assign n19944 = ( ~n19933 & n19942 ) | ( ~n19933 & n19943 ) | ( n19942 & n19943 ) ;
  assign n19945 = ~n19939 & n19944 ;
  assign n19946 = n19938 | n19945 ;
  assign n19947 = n19929 & n19946 ;
  assign n19948 = n19929 & ~n19947 ;
  assign n19949 = n19946 & ~n19947 ;
  assign n19950 = n19948 | n19949 ;
  assign n19951 = n6147 & n10367 ;
  assign n19952 = x47 & x60 ;
  assign n19953 = x46 & x61 ;
  assign n19954 = n19952 | n19953 ;
  assign n19955 = ~n19951 & n19954 ;
  assign n19956 = n19853 & n19955 ;
  assign n19957 = n19853 & ~n19956 ;
  assign n19958 = ~n19853 & n19955 ;
  assign n19959 = n19957 | n19958 ;
  assign n19960 = n7565 & n12860 ;
  assign n19961 = n7112 & n8903 ;
  assign n19962 = n19960 | n19961 ;
  assign n19963 = n7567 & n10013 ;
  assign n19964 = x57 & n19963 ;
  assign n19965 = ( x57 & ~n19962 ) | ( x57 & n19964 ) | ( ~n19962 & n19964 ) ;
  assign n19966 = x50 & n19965 ;
  assign n19967 = n19962 | n19963 ;
  assign n19968 = x51 & x56 ;
  assign n19969 = ( n13618 & ~n19963 ) | ( n13618 & n19968 ) | ( ~n19963 & n19968 ) ;
  assign n19970 = n13618 & n19968 ;
  assign n19971 = ( ~n19962 & n19969 ) | ( ~n19962 & n19970 ) | ( n19969 & n19970 ) ;
  assign n19972 = ~n19967 & n19971 ;
  assign n19973 = n19966 | n19972 ;
  assign n19974 = ( x54 & ~n8355 ) | ( x54 & n17212 ) | ( ~n8355 & n17212 ) ;
  assign n19975 = ( x54 & n8355 ) | ( x54 & n17212 ) | ( n8355 & n17212 ) ;
  assign n19976 = n8355 | n17212 ;
  assign n19977 = ( ~n19974 & n19975 ) | ( ~n19974 & n19976 ) | ( n19975 & n19976 ) ;
  assign n19978 = ( n8355 & n19974 ) | ( n8355 & ~n19977 ) | ( n19974 & ~n19977 ) ;
  assign n19979 = ( n19959 & n19973 ) | ( n19959 & ~n19978 ) | ( n19973 & ~n19978 ) ;
  assign n19980 = ( n19959 & ~n19973 ) | ( n19959 & n19978 ) | ( ~n19973 & n19978 ) ;
  assign n19981 = ( ~n19959 & n19979 ) | ( ~n19959 & n19980 ) | ( n19979 & n19980 ) ;
  assign n19982 = n19950 & n19981 ;
  assign n19983 = n19950 | n19981 ;
  assign n19984 = ~n19982 & n19983 ;
  assign n19985 = n19822 | n19823 ;
  assign n19986 = ( n19822 & n19824 ) | ( n19822 & n19985 ) | ( n19824 & n19985 ) ;
  assign n19987 = n19984 | n19986 ;
  assign n19988 = n19984 & n19986 ;
  assign n19989 = n19987 & ~n19988 ;
  assign n19990 = n19868 | n19887 ;
  assign n19991 = n19889 & n19990 ;
  assign n19992 = n19871 & n19884 ;
  assign n19993 = n19734 | n19813 ;
  assign n19994 = ( n19813 & n19816 ) | ( n19813 & n19993 ) | ( n19816 & n19993 ) ;
  assign n19995 = n19870 & n19994 ;
  assign n19996 = ( n19992 & n19994 ) | ( n19992 & n19995 ) | ( n19994 & n19995 ) ;
  assign n19997 = n19870 | n19994 ;
  assign n19998 = n19992 | n19997 ;
  assign n19999 = ~n19996 & n19998 ;
  assign n20000 = n19860 | n19865 ;
  assign n20001 = ( n19860 & n19863 ) | ( n19860 & n20000 ) | ( n19863 & n20000 ) ;
  assign n20002 = n19999 | n20001 ;
  assign n20003 = n19999 & n20001 ;
  assign n20004 = n20002 & ~n20003 ;
  assign n20005 = n19868 & n19887 ;
  assign n20006 = n20004 & n20005 ;
  assign n20007 = ( n19991 & n20004 ) | ( n19991 & n20006 ) | ( n20004 & n20006 ) ;
  assign n20008 = n20004 | n20005 ;
  assign n20009 = n19991 | n20008 ;
  assign n20010 = ~n20007 & n20009 ;
  assign n20011 = n19989 & n20010 ;
  assign n20012 = n19989 | n20010 ;
  assign n20013 = ~n20011 & n20012 ;
  assign n20014 = ( n19827 & n19829 ) | ( n19827 & n19892 ) | ( n19829 & n19892 ) ;
  assign n20033 = ( n20013 & ~n20014 ) | ( n20013 & n20032 ) | ( ~n20014 & n20032 ) ;
  assign n20034 = ( ~n20013 & n20014 ) | ( ~n20013 & n20033 ) | ( n20014 & n20033 ) ;
  assign n20035 = ( ~n20032 & n20033 ) | ( ~n20032 & n20034 ) | ( n20033 & n20034 ) ;
  assign n20036 = n19973 & n19978 ;
  assign n20037 = n19973 & ~n20036 ;
  assign n20038 = ~n19973 & n19978 ;
  assign n20039 = n19959 & ~n20038 ;
  assign n20040 = ~n20037 & n20039 ;
  assign n20041 = ( n19959 & n20036 ) | ( n19959 & ~n20040 ) | ( n20036 & ~n20040 ) ;
  assign n20042 = n7874 & n12860 ;
  assign n20043 = n7567 & n8903 ;
  assign n20044 = n20042 | n20043 ;
  assign n20045 = n8161 & n10013 ;
  assign n20046 = n15873 & n20045 ;
  assign n20047 = x52 & x56 ;
  assign n20048 = n8360 | n20047 ;
  assign n20049 = n15873 | n20048 ;
  assign n20050 = ( n20044 & ~n20045 ) | ( n20044 & n20049 ) | ( ~n20045 & n20049 ) ;
  assign n20051 = ( ~n20044 & n20046 ) | ( ~n20044 & n20050 ) | ( n20046 & n20050 ) ;
  assign n20052 = n19928 & n20051 ;
  assign n20053 = ( n19947 & n20051 ) | ( n19947 & n20052 ) | ( n20051 & n20052 ) ;
  assign n20054 = n19928 & ~n20051 ;
  assign n20055 = ( n19947 & ~n20051 ) | ( n19947 & n20054 ) | ( ~n20051 & n20054 ) ;
  assign n20056 = ( n20051 & ~n20053 ) | ( n20051 & n20055 ) | ( ~n20053 & n20055 ) ;
  assign n20057 = n20041 & n20056 ;
  assign n20058 = n20041 & ~n20057 ;
  assign n20059 = ~n20041 & n20056 ;
  assign n20060 = n20058 | n20059 ;
  assign n20061 = n19982 | n19988 ;
  assign n20062 = n20060 | n20061 ;
  assign n20063 = n20060 & n20061 ;
  assign n20064 = n20062 & ~n20063 ;
  assign n20065 = x54 & n17212 ;
  assign n20066 = n8355 & ~n20065 ;
  assign n20067 = n20065 | n20066 ;
  assign n20068 = n19967 | n20067 ;
  assign n20069 = n19967 & n20067 ;
  assign n20070 = n20068 & ~n20069 ;
  assign n20071 = n19939 | n20070 ;
  assign n20072 = n19939 & n20070 ;
  assign n20073 = n20071 & ~n20072 ;
  assign n20074 = n19996 | n19999 ;
  assign n20075 = ( n19996 & n20001 ) | ( n19996 & n20074 ) | ( n20001 & n20074 ) ;
  assign n20076 = n20073 | n20075 ;
  assign n20077 = n20073 & n20075 ;
  assign n20078 = n20076 & ~n20077 ;
  assign n20079 = n5610 & n10856 ;
  assign n20080 = n5975 & n10561 ;
  assign n20081 = n20079 | n20080 ;
  assign n20082 = n6147 & n10684 ;
  assign n20083 = x45 & n20082 ;
  assign n20084 = ( x45 & ~n20081 ) | ( x45 & n20083 ) | ( ~n20081 & n20083 ) ;
  assign n20085 = x63 & n20084 ;
  assign n20086 = n20081 | n20082 ;
  assign n20087 = x47 & x61 ;
  assign n20088 = ( n17554 & ~n20082 ) | ( n17554 & n20087 ) | ( ~n20082 & n20087 ) ;
  assign n20089 = n17554 & n20087 ;
  assign n20090 = ( ~n20081 & n20088 ) | ( ~n20081 & n20089 ) | ( n20088 & n20089 ) ;
  assign n20091 = ~n20086 & n20090 ;
  assign n20092 = n20085 | n20091 ;
  assign n20093 = n19951 | n19955 ;
  assign n20094 = ( n19853 & n19951 ) | ( n19853 & n20093 ) | ( n19951 & n20093 ) ;
  assign n20095 = n20092 & ~n20094 ;
  assign n20096 = ~n20092 & n20094 ;
  assign n20097 = n20095 | n20096 ;
  assign n20098 = n6345 & n10975 ;
  assign n20099 = n6759 & n10370 ;
  assign n20100 = n20098 | n20099 ;
  assign n20101 = n6834 & n9831 ;
  assign n20102 = x60 & n20101 ;
  assign n20103 = ( x60 & ~n20100 ) | ( x60 & n20102 ) | ( ~n20100 & n20102 ) ;
  assign n20104 = x48 & n20103 ;
  assign n20105 = n20100 | n20101 ;
  assign n20106 = x49 & x59 ;
  assign n20107 = x50 & x58 ;
  assign n20108 = ( ~n20101 & n20106 ) | ( ~n20101 & n20107 ) | ( n20106 & n20107 ) ;
  assign n20109 = n20106 & n20107 ;
  assign n20110 = ( ~n20100 & n20108 ) | ( ~n20100 & n20109 ) | ( n20108 & n20109 ) ;
  assign n20111 = ~n20105 & n20110 ;
  assign n20112 = n20104 | n20111 ;
  assign n20113 = n20097 & n20112 ;
  assign n20114 = n20097 | n20112 ;
  assign n20115 = ~n20113 & n20114 ;
  assign n20116 = ( n20064 & ~n20078 ) | ( n20064 & n20115 ) | ( ~n20078 & n20115 ) ;
  assign n20117 = ( ~n20064 & n20078 ) | ( ~n20064 & n20116 ) | ( n20078 & n20116 ) ;
  assign n20118 = n19989 | n20007 ;
  assign n20119 = ( n20007 & n20010 ) | ( n20007 & n20118 ) | ( n20010 & n20118 ) ;
  assign n20120 = n20116 & n20119 ;
  assign n20121 = ~n20115 & n20119 ;
  assign n20122 = ( n20117 & n20120 ) | ( n20117 & n20121 ) | ( n20120 & n20121 ) ;
  assign n20123 = n20116 | n20119 ;
  assign n20124 = n20115 & ~n20119 ;
  assign n20125 = ( n20117 & n20123 ) | ( n20117 & ~n20124 ) | ( n20123 & ~n20124 ) ;
  assign n20126 = ~n20122 & n20125 ;
  assign n20127 = n20013 & n20014 ;
  assign n20128 = n20013 | n20014 ;
  assign n20129 = n20127 | n20128 ;
  assign n20130 = ( n20032 & n20127 ) | ( n20032 & n20129 ) | ( n20127 & n20129 ) ;
  assign n20131 = n20126 | n20130 ;
  assign n20132 = n20125 & n20129 ;
  assign n20133 = n20125 & n20127 ;
  assign n20134 = ( n20032 & n20132 ) | ( n20032 & n20133 ) | ( n20132 & n20133 ) ;
  assign n20135 = ~n20122 & n20134 ;
  assign n20136 = n20131 & ~n20135 ;
  assign n20137 = n20122 | n20133 ;
  assign n20138 = n20122 | n20125 ;
  assign n20139 = ( n20122 & n20129 ) | ( n20122 & n20138 ) | ( n20129 & n20138 ) ;
  assign n20140 = ( n20032 & n20137 ) | ( n20032 & n20139 ) | ( n20137 & n20139 ) ;
  assign n20141 = n20078 & n20115 ;
  assign n20142 = n20078 | n20115 ;
  assign n20143 = ~n20141 & n20142 ;
  assign n20144 = n20064 & n20143 ;
  assign n20145 = n20063 | n20144 ;
  assign n20146 = x51 & x58 ;
  assign n20147 = n7874 & n8708 ;
  assign n20148 = n7567 & n9272 ;
  assign n20149 = n20147 | n20148 ;
  assign n20150 = n8161 & n8903 ;
  assign n20151 = n20146 & n20150 ;
  assign n20152 = ( n20146 & ~n20149 ) | ( n20146 & n20151 ) | ( ~n20149 & n20151 ) ;
  assign n20153 = n20149 | n20150 ;
  assign n20154 = x52 & x57 ;
  assign n20155 = ( n14726 & ~n20150 ) | ( n14726 & n20154 ) | ( ~n20150 & n20154 ) ;
  assign n20156 = n14726 & n20154 ;
  assign n20157 = ( ~n20149 & n20155 ) | ( ~n20149 & n20156 ) | ( n20155 & n20156 ) ;
  assign n20158 = ~n20153 & n20157 ;
  assign n20159 = n20152 | n20158 ;
  assign n20160 = n6345 & n9737 ;
  assign n20161 = n6759 & n10367 ;
  assign n20162 = n20160 | n20161 ;
  assign n20163 = n6834 & n10370 ;
  assign n20164 = x48 & n20163 ;
  assign n20165 = ( x48 & ~n20162 ) | ( x48 & n20164 ) | ( ~n20162 & n20164 ) ;
  assign n20166 = x61 & n20165 ;
  assign n20167 = n20162 | n20163 ;
  assign n20168 = x49 & x60 ;
  assign n20169 = x50 & x59 ;
  assign n20170 = ( ~n20163 & n20168 ) | ( ~n20163 & n20169 ) | ( n20168 & n20169 ) ;
  assign n20171 = n20168 & n20169 ;
  assign n20172 = ( ~n20162 & n20170 ) | ( ~n20162 & n20171 ) | ( n20170 & n20171 ) ;
  assign n20173 = ~n20167 & n20172 ;
  assign n20174 = n20166 | n20173 ;
  assign n20175 = n20086 | n20174 ;
  assign n20176 = ~n20086 & n20174 ;
  assign n20177 = ( ~n20174 & n20175 ) | ( ~n20174 & n20176 ) | ( n20175 & n20176 ) ;
  assign n20178 = n20159 & n20177 ;
  assign n20179 = n20159 | n20177 ;
  assign n20180 = ~n20178 & n20179 ;
  assign n20187 = n19939 | n20069 ;
  assign n20188 = ( n20069 & n20070 ) | ( n20069 & n20187 ) | ( n20070 & n20187 ) ;
  assign n20181 = x55 & n18087 ;
  assign n20182 = n8357 & n20181 ;
  assign n20183 = ( x55 & ~n8357 ) | ( x55 & n18087 ) | ( ~n8357 & n18087 ) ;
  assign n20184 = x55 | n18087 ;
  assign n20185 = ( n20181 & n20183 ) | ( n20181 & n20184 ) | ( n20183 & n20184 ) ;
  assign n20186 = ( ~n20181 & n20182 ) | ( ~n20181 & n20185 ) | ( n20182 & n20185 ) ;
  assign n20189 = n20186 & n20188 ;
  assign n20190 = n20188 & ~n20189 ;
  assign n20191 = n20186 & ~n20188 ;
  assign n20192 = ( n20092 & n20094 ) | ( n20092 & n20112 ) | ( n20094 & n20112 ) ;
  assign n20193 = n20191 | n20192 ;
  assign n20194 = n20190 | n20193 ;
  assign n20195 = n20191 & n20192 ;
  assign n20196 = ( n20190 & n20192 ) | ( n20190 & n20195 ) | ( n20192 & n20195 ) ;
  assign n20197 = n20194 & ~n20196 ;
  assign n20198 = n20073 | n20115 ;
  assign n20199 = ( n20075 & n20115 ) | ( n20075 & n20198 ) | ( n20115 & n20198 ) ;
  assign n20200 = n20197 & n20199 ;
  assign n20201 = n20077 & n20197 ;
  assign n20202 = ( n20078 & n20200 ) | ( n20078 & n20201 ) | ( n20200 & n20201 ) ;
  assign n20203 = n20197 | n20199 ;
  assign n20204 = n20077 | n20197 ;
  assign n20205 = ( n20078 & n20203 ) | ( n20078 & n20204 ) | ( n20203 & n20204 ) ;
  assign n20206 = ~n20202 & n20205 ;
  assign n20207 = x46 & x63 ;
  assign n20208 = n20045 & n20207 ;
  assign n20209 = ( n20044 & n20207 ) | ( n20044 & n20208 ) | ( n20207 & n20208 ) ;
  assign n20210 = n20045 | n20207 ;
  assign n20211 = n20044 | n20210 ;
  assign n20212 = ~n20209 & n20211 ;
  assign n20213 = n20105 | n20212 ;
  assign n20214 = n20105 & n20212 ;
  assign n20215 = n20213 & ~n20214 ;
  assign n20216 = n20053 & n20215 ;
  assign n20217 = ( n20056 & n20215 ) | ( n20056 & n20216 ) | ( n20215 & n20216 ) ;
  assign n20218 = ( n20041 & n20216 ) | ( n20041 & n20217 ) | ( n20216 & n20217 ) ;
  assign n20219 = n20053 | n20215 ;
  assign n20220 = n20056 | n20219 ;
  assign n20221 = ( n20041 & n20219 ) | ( n20041 & n20220 ) | ( n20219 & n20220 ) ;
  assign n20222 = ~n20218 & n20221 ;
  assign n20223 = ( n20180 & n20206 ) | ( n20180 & ~n20222 ) | ( n20206 & ~n20222 ) ;
  assign n20224 = ( ~n20206 & n20222 ) | ( ~n20206 & n20223 ) | ( n20222 & n20223 ) ;
  assign n20225 = ( ~n20180 & n20223 ) | ( ~n20180 & n20224 ) | ( n20223 & n20224 ) ;
  assign n20226 = ( n20139 & ~n20145 ) | ( n20139 & n20225 ) | ( ~n20145 & n20225 ) ;
  assign n20227 = ( n20137 & ~n20145 ) | ( n20137 & n20225 ) | ( ~n20145 & n20225 ) ;
  assign n20228 = ( n20032 & n20226 ) | ( n20032 & n20227 ) | ( n20226 & n20227 ) ;
  assign n20229 = ( n20145 & ~n20225 ) | ( n20145 & n20226 ) | ( ~n20225 & n20226 ) ;
  assign n20230 = ( n20145 & ~n20225 ) | ( n20145 & n20227 ) | ( ~n20225 & n20227 ) ;
  assign n20231 = ( n20032 & n20229 ) | ( n20032 & n20230 ) | ( n20229 & n20230 ) ;
  assign n20232 = ( ~n20140 & n20228 ) | ( ~n20140 & n20231 ) | ( n20228 & n20231 ) ;
  assign n20233 = n20153 | n20167 ;
  assign n20234 = n20153 & n20167 ;
  assign n20235 = n20233 & ~n20234 ;
  assign n20236 = n9737 & n10866 ;
  assign n20237 = n6834 & n10367 ;
  assign n20238 = n20236 | n20237 ;
  assign n20239 = n7112 & n10370 ;
  assign n20240 = x61 & n20239 ;
  assign n20241 = ( x61 & ~n20238 ) | ( x61 & n20240 ) | ( ~n20238 & n20240 ) ;
  assign n20242 = x49 & n20241 ;
  assign n20243 = n20238 | n20239 ;
  assign n20244 = x50 & x60 ;
  assign n20245 = x51 & x59 ;
  assign n20246 = ( ~n20239 & n20244 ) | ( ~n20239 & n20245 ) | ( n20244 & n20245 ) ;
  assign n20247 = n20244 & n20245 ;
  assign n20248 = ( ~n20238 & n20246 ) | ( ~n20238 & n20247 ) | ( n20246 & n20247 ) ;
  assign n20249 = ~n20243 & n20248 ;
  assign n20250 = n20242 | n20249 ;
  assign n20251 = n20235 & n20250 ;
  assign n20252 = n20235 & ~n20251 ;
  assign n20253 = n20250 & ~n20251 ;
  assign n20254 = n20252 | n20253 ;
  assign n20255 = n20086 & n20173 ;
  assign n20256 = ( n20086 & n20166 ) | ( n20086 & n20255 ) | ( n20166 & n20255 ) ;
  assign n20257 = n20159 | n20256 ;
  assign n20258 = ( n20177 & n20256 ) | ( n20177 & n20257 ) | ( n20256 & n20257 ) ;
  assign n20259 = n20254 | n20258 ;
  assign n20260 = n20254 & n20258 ;
  assign n20261 = n20259 & ~n20260 ;
  assign n20262 = n20189 | n20196 ;
  assign n20263 = n20261 | n20262 ;
  assign n20264 = n20261 & n20262 ;
  assign n20265 = n20263 & ~n20264 ;
  assign n20266 = n20180 | n20218 ;
  assign n20267 = ( n20218 & n20222 ) | ( n20218 & n20266 ) | ( n20222 & n20266 ) ;
  assign n20268 = n8357 & ~n20181 ;
  assign n20269 = n20181 | n20268 ;
  assign n20270 = n6762 & n10561 ;
  assign n20271 = x47 & x63 ;
  assign n20272 = n18270 | n20271 ;
  assign n20273 = ~n20270 & n20272 ;
  assign n20274 = n20269 & n20273 ;
  assign n20275 = n20269 | n20273 ;
  assign n20276 = ~n20274 & n20275 ;
  assign n20277 = n8161 & n9272 ;
  assign n20278 = x54 & x58 ;
  assign n20279 = n20047 & n20278 ;
  assign n20280 = n20277 | n20279 ;
  assign n20281 = n8355 & n8903 ;
  assign n20282 = x58 & n20281 ;
  assign n20283 = ( x58 & ~n20280 ) | ( x58 & n20282 ) | ( ~n20280 & n20282 ) ;
  assign n20284 = x52 & n20283 ;
  assign n20285 = n20280 | n20281 ;
  assign n20286 = x53 & x57 ;
  assign n20287 = ( n8146 & ~n20281 ) | ( n8146 & n20286 ) | ( ~n20281 & n20286 ) ;
  assign n20288 = n8146 & n20286 ;
  assign n20289 = ( ~n20280 & n20287 ) | ( ~n20280 & n20288 ) | ( n20287 & n20288 ) ;
  assign n20290 = ~n20285 & n20289 ;
  assign n20291 = n20284 | n20290 ;
  assign n20292 = n20276 & n20291 ;
  assign n20293 = n20276 & ~n20292 ;
  assign n20294 = n20291 & ~n20292 ;
  assign n20295 = n20293 | n20294 ;
  assign n20296 = n20105 | n20209 ;
  assign n20297 = ( n20209 & n20212 ) | ( n20209 & n20296 ) | ( n20212 & n20296 ) ;
  assign n20298 = n20295 | n20297 ;
  assign n20299 = n20295 & n20297 ;
  assign n20300 = n20298 & ~n20299 ;
  assign n20301 = n20267 & n20300 ;
  assign n20302 = n20267 & ~n20301 ;
  assign n20303 = ~n20267 & n20300 ;
  assign n20304 = n20265 & n20303 ;
  assign n20305 = ( n20265 & n20302 ) | ( n20265 & n20304 ) | ( n20302 & n20304 ) ;
  assign n20306 = n20265 | n20267 ;
  assign n20307 = ( n20265 & ~n20301 ) | ( n20265 & n20306 ) | ( ~n20301 & n20306 ) ;
  assign n20308 = n20303 | n20307 ;
  assign n20309 = ~n20305 & n20308 ;
  assign n20310 = n20180 & n20222 ;
  assign n20311 = n20180 | n20222 ;
  assign n20312 = ~n20310 & n20311 ;
  assign n20313 = n20202 | n20312 ;
  assign n20314 = ( n20202 & n20206 ) | ( n20202 & n20313 ) | ( n20206 & n20313 ) ;
  assign n20315 = n20309 | n20314 ;
  assign n20316 = n20309 & n20314 ;
  assign n20317 = n20315 & ~n20316 ;
  assign n20318 = n20145 & n20225 ;
  assign n20319 = n20145 | n20225 ;
  assign n20320 = n20139 & n20319 ;
  assign n20321 = n20318 | n20320 ;
  assign n20322 = n20318 | n20319 ;
  assign n20323 = ( n20137 & n20318 ) | ( n20137 & n20322 ) | ( n20318 & n20322 ) ;
  assign n20324 = ( n20032 & n20321 ) | ( n20032 & n20323 ) | ( n20321 & n20323 ) ;
  assign n20325 = n20317 | n20324 ;
  assign n20326 = n20315 & n20318 ;
  assign n20327 = ( n20315 & n20320 ) | ( n20315 & n20326 ) | ( n20320 & n20326 ) ;
  assign n20328 = n20315 & n20323 ;
  assign n20329 = ( n20032 & n20327 ) | ( n20032 & n20328 ) | ( n20327 & n20328 ) ;
  assign n20330 = ~n20316 & n20329 ;
  assign n20331 = n20325 & ~n20330 ;
  assign n20332 = n20243 | n20285 ;
  assign n20333 = n20243 & n20285 ;
  assign n20334 = n20332 & ~n20333 ;
  assign n20335 = n20270 | n20273 ;
  assign n20336 = ( n20269 & n20270 ) | ( n20269 & n20335 ) | ( n20270 & n20335 ) ;
  assign n20337 = n20334 | n20336 ;
  assign n20338 = n20334 & n20336 ;
  assign n20339 = n20337 & ~n20338 ;
  assign n20340 = n20234 | n20251 ;
  assign n20341 = n20339 | n20340 ;
  assign n20342 = n20339 & n20340 ;
  assign n20343 = n20341 & ~n20342 ;
  assign n20344 = n20292 | n20297 ;
  assign n20345 = ( n20292 & n20295 ) | ( n20292 & n20344 ) | ( n20295 & n20344 ) ;
  assign n20346 = n20343 | n20345 ;
  assign n20347 = n20343 & n20345 ;
  assign n20348 = n20346 & ~n20347 ;
  assign n20349 = n12770 & n18896 ;
  assign n20350 = n6345 & n10856 ;
  assign n20351 = n20349 | n20350 ;
  assign n20352 = n7112 & n10367 ;
  assign n20353 = x63 & n20352 ;
  assign n20354 = ( x63 & ~n20351 ) | ( x63 & n20353 ) | ( ~n20351 & n20353 ) ;
  assign n20355 = x48 & n20354 ;
  assign n20356 = n20351 | n20352 ;
  assign n20357 = x50 & x61 ;
  assign n20358 = x51 & x60 ;
  assign n20359 = ( ~n20352 & n20357 ) | ( ~n20352 & n20358 ) | ( n20357 & n20358 ) ;
  assign n20360 = n20357 & n20358 ;
  assign n20361 = ( ~n20351 & n20359 ) | ( ~n20351 & n20360 ) | ( n20359 & n20360 ) ;
  assign n20362 = ~n20356 & n20361 ;
  assign n20363 = n20355 | n20362 ;
  assign n20364 = x56 & x62 ;
  assign n20365 = x49 & n20364 ;
  assign n20366 = n10013 & n20365 ;
  assign n20367 = n10013 & ~n20365 ;
  assign n20368 = x56 | n18598 ;
  assign n20369 = ~n20365 & n20368 ;
  assign n20370 = ~n20367 & n20369 ;
  assign n20371 = n20366 | n20370 ;
  assign n20372 = n20363 & n20371 ;
  assign n20373 = n20363 & ~n20372 ;
  assign n20374 = n9829 & n11935 ;
  assign n20375 = n8161 & n9831 ;
  assign n20376 = n20374 | n20375 ;
  assign n20377 = n8355 & n9272 ;
  assign n20378 = x59 & n20377 ;
  assign n20379 = ( x59 & ~n20376 ) | ( x59 & n20378 ) | ( ~n20376 & n20378 ) ;
  assign n20380 = x52 & n20379 ;
  assign n20381 = n20376 | n20377 ;
  assign n20382 = x53 & x58 ;
  assign n20383 = ( n15088 & ~n20377 ) | ( n15088 & n20382 ) | ( ~n20377 & n20382 ) ;
  assign n20384 = n15088 & n20382 ;
  assign n20385 = ( ~n20376 & n20383 ) | ( ~n20376 & n20384 ) | ( n20383 & n20384 ) ;
  assign n20386 = ~n20381 & n20385 ;
  assign n20387 = n20380 | n20386 ;
  assign n20388 = ~n20363 & n20371 ;
  assign n20389 = n20387 & n20388 ;
  assign n20390 = ( n20373 & n20387 ) | ( n20373 & n20389 ) | ( n20387 & n20389 ) ;
  assign n20391 = n20387 | n20388 ;
  assign n20392 = n20373 | n20391 ;
  assign n20393 = ~n20390 & n20392 ;
  assign n20394 = n20260 & n20393 ;
  assign n20395 = ( n20264 & n20393 ) | ( n20264 & n20394 ) | ( n20393 & n20394 ) ;
  assign n20396 = n20260 | n20393 ;
  assign n20397 = n20264 | n20396 ;
  assign n20398 = ~n20395 & n20397 ;
  assign n20399 = n20348 & n20398 ;
  assign n20400 = n20348 | n20398 ;
  assign n20401 = ~n20399 & n20400 ;
  assign n20402 = n20301 & n20401 ;
  assign n20403 = ( n20305 & n20401 ) | ( n20305 & n20402 ) | ( n20401 & n20402 ) ;
  assign n20404 = n20301 | n20401 ;
  assign n20405 = n20305 | n20404 ;
  assign n20406 = ~n20403 & n20405 ;
  assign n20407 = n20316 | n20328 ;
  assign n20408 = n20315 | n20316 ;
  assign n20409 = ( n20316 & n20318 ) | ( n20316 & n20408 ) | ( n20318 & n20408 ) ;
  assign n20410 = ( n20320 & n20408 ) | ( n20320 & n20409 ) | ( n20408 & n20409 ) ;
  assign n20411 = ( n20032 & n20407 ) | ( n20032 & n20410 ) | ( n20407 & n20410 ) ;
  assign n20412 = ~n20406 & n20411 ;
  assign n20413 = n20406 & ~n20411 ;
  assign n20414 = n20412 | n20413 ;
  assign n20415 = n7567 & n10367 ;
  assign n20416 = x52 & n12770 ;
  assign n20417 = x51 & n10856 ;
  assign n20418 = n20416 | n20417 ;
  assign n20419 = x49 & ~n20415 ;
  assign n20420 = n20418 & n20419 ;
  assign n20421 = n20415 | n20420 ;
  assign n20422 = x51 & x61 ;
  assign n20423 = x52 & x60 ;
  assign n20424 = ( ~n20415 & n20422 ) | ( ~n20415 & n20423 ) | ( n20422 & n20423 ) ;
  assign n20425 = n20422 & n20423 ;
  assign n20426 = ( ~n20420 & n20424 ) | ( ~n20420 & n20425 ) | ( n20424 & n20425 ) ;
  assign n20427 = ~n20421 & n20426 ;
  assign n20428 = x49 & x63 ;
  assign n20429 = ~n20420 & n20428 ;
  assign n20430 = ~n20356 & n20429 ;
  assign n20431 = ( ~n20356 & n20427 ) | ( ~n20356 & n20430 ) | ( n20427 & n20430 ) ;
  assign n20432 = n20356 & ~n20429 ;
  assign n20433 = ~n20427 & n20432 ;
  assign n20434 = n20431 | n20433 ;
  assign n20435 = n8355 & n9831 ;
  assign n20436 = x55 & x59 ;
  assign n20437 = n20286 & n20436 ;
  assign n20438 = n20435 | n20437 ;
  assign n20439 = n8357 & n9272 ;
  assign n20440 = x59 & n20439 ;
  assign n20441 = ( x59 & ~n20438 ) | ( x59 & n20440 ) | ( ~n20438 & n20440 ) ;
  assign n20442 = x53 & n20441 ;
  assign n20443 = n20438 | n20439 ;
  assign n20444 = ( n12860 & n20278 ) | ( n12860 & ~n20439 ) | ( n20278 & ~n20439 ) ;
  assign n20445 = n12860 & n20278 ;
  assign n20446 = ( ~n20438 & n20444 ) | ( ~n20438 & n20445 ) | ( n20444 & n20445 ) ;
  assign n20447 = ~n20443 & n20446 ;
  assign n20448 = n20442 | n20447 ;
  assign n20449 = n20434 & n20448 ;
  assign n20450 = n20434 | n20448 ;
  assign n20451 = ~n20449 & n20450 ;
  assign n20452 = n20342 & n20451 ;
  assign n20453 = ( n20347 & n20451 ) | ( n20347 & n20452 ) | ( n20451 & n20452 ) ;
  assign n20454 = n20342 | n20451 ;
  assign n20455 = n20347 | n20454 ;
  assign n20456 = ~n20453 & n20455 ;
  assign n20457 = n19046 & n20365 ;
  assign n20458 = ( n19046 & n20367 ) | ( n19046 & n20457 ) | ( n20367 & n20457 ) ;
  assign n20459 = n19046 | n20365 ;
  assign n20460 = n20367 | n20459 ;
  assign n20461 = ~n20458 & n20460 ;
  assign n20462 = n20381 | n20461 ;
  assign n20463 = n20381 & n20461 ;
  assign n20464 = n20462 & ~n20463 ;
  assign n20465 = n20333 | n20336 ;
  assign n20466 = ( n20333 & n20334 ) | ( n20333 & n20465 ) | ( n20334 & n20465 ) ;
  assign n20467 = n20372 & n20466 ;
  assign n20468 = ( n20390 & n20466 ) | ( n20390 & n20467 ) | ( n20466 & n20467 ) ;
  assign n20469 = n20372 | n20466 ;
  assign n20470 = n20390 | n20469 ;
  assign n20471 = ~n20468 & n20470 ;
  assign n20472 = n20464 & n20471 ;
  assign n20473 = n20464 | n20471 ;
  assign n20474 = ~n20472 & n20473 ;
  assign n20475 = n20456 & n20474 ;
  assign n20476 = n20456 | n20474 ;
  assign n20477 = ~n20475 & n20476 ;
  assign n20478 = n20348 | n20395 ;
  assign n20479 = ( n20395 & n20398 ) | ( n20395 & n20478 ) | ( n20398 & n20478 ) ;
  assign n20480 = n20477 | n20479 ;
  assign n20481 = n20477 & n20479 ;
  assign n20482 = n20480 & ~n20481 ;
  assign n20483 = n20405 & n20409 ;
  assign n20484 = n20405 & n20408 ;
  assign n20485 = ( n20320 & n20483 ) | ( n20320 & n20484 ) | ( n20483 & n20484 ) ;
  assign n20486 = n20403 | n20485 ;
  assign n20487 = n20403 | n20405 ;
  assign n20488 = ( n20316 & n20403 ) | ( n20316 & n20487 ) | ( n20403 & n20487 ) ;
  assign n20489 = ( n20328 & n20487 ) | ( n20328 & n20488 ) | ( n20487 & n20488 ) ;
  assign n20490 = ( n20032 & n20486 ) | ( n20032 & n20489 ) | ( n20486 & n20489 ) ;
  assign n20491 = n20482 | n20490 ;
  assign n20492 = n20401 & n20480 ;
  assign n20493 = n20305 & n20480 ;
  assign n20494 = ( n20402 & n20492 ) | ( n20402 & n20493 ) | ( n20492 & n20493 ) ;
  assign n20495 = ( n20480 & n20485 ) | ( n20480 & n20494 ) | ( n20485 & n20494 ) ;
  assign n20496 = n20480 & n20487 ;
  assign n20497 = n20403 & n20480 ;
  assign n20498 = n20316 & n20480 ;
  assign n20499 = ( n20487 & n20497 ) | ( n20487 & n20498 ) | ( n20497 & n20498 ) ;
  assign n20500 = ( n20315 & n20496 ) | ( n20315 & n20499 ) | ( n20496 & n20499 ) ;
  assign n20501 = n20496 & n20499 ;
  assign n20502 = ( n20323 & n20500 ) | ( n20323 & n20501 ) | ( n20500 & n20501 ) ;
  assign n20503 = ( n20032 & n20495 ) | ( n20032 & n20502 ) | ( n20495 & n20502 ) ;
  assign n20504 = ~n20481 & n20503 ;
  assign n20505 = n20491 & ~n20504 ;
  assign n20506 = n20481 | n20494 ;
  assign n20507 = n20480 | n20481 ;
  assign n20508 = ( n20485 & n20506 ) | ( n20485 & n20507 ) | ( n20506 & n20507 ) ;
  assign n20509 = n20481 | n20502 ;
  assign n20510 = ( n20032 & n20508 ) | ( n20032 & n20509 ) | ( n20508 & n20509 ) ;
  assign n20511 = n20453 | n20475 ;
  assign n20512 = n8161 & n10367 ;
  assign n20513 = x53 & x60 ;
  assign n20514 = x52 & x61 ;
  assign n20515 = n20513 | n20514 ;
  assign n20516 = ~n20512 & n20515 ;
  assign n20517 = n20443 & n20516 ;
  assign n20518 = n20443 & ~n20517 ;
  assign n20519 = ~n20443 & n20516 ;
  assign n20520 = n20518 | n20519 ;
  assign n20521 = n20381 | n20458 ;
  assign n20522 = ( n20458 & n20461 ) | ( n20458 & n20521 ) | ( n20461 & n20521 ) ;
  assign n20523 = n20520 | n20522 ;
  assign n20524 = n20520 & n20522 ;
  assign n20525 = n20523 & ~n20524 ;
  assign n20526 = n20427 | n20429 ;
  assign n20527 = ( n20356 & n20448 ) | ( n20356 & n20526 ) | ( n20448 & n20526 ) ;
  assign n20528 = n20525 | n20527 ;
  assign n20529 = n20525 & n20527 ;
  assign n20530 = n20528 & ~n20529 ;
  assign n20531 = x54 & x59 ;
  assign n20532 = n18310 | n20531 ;
  assign n20533 = n8357 & n9831 ;
  assign n20534 = x50 & x63 ;
  assign n20535 = ~n20533 & n20534 ;
  assign n20536 = n20532 | n20533 ;
  assign n20537 = ( n20533 & n20535 ) | ( n20533 & n20536 ) | ( n20535 & n20536 ) ;
  assign n20538 = n20532 & ~n20537 ;
  assign n20539 = ( ~n20532 & n20533 ) | ( ~n20532 & n20534 ) | ( n20533 & n20534 ) ;
  assign n20540 = n20534 & n20539 ;
  assign n20541 = n20538 | n20540 ;
  assign n20542 = ~n20421 & n20541 ;
  assign n20543 = n20421 & ~n20541 ;
  assign n20544 = n20542 | n20543 ;
  assign n20545 = x62 & n15873 ;
  assign n20546 = n8903 & n20545 ;
  assign n20547 = n8903 & ~n20545 ;
  assign n20548 = n20545 | n20547 ;
  assign n20549 = ( x57 & n15602 ) | ( x57 & ~n20545 ) | ( n15602 & ~n20545 ) ;
  assign n20550 = x57 & n15602 ;
  assign n20551 = ( ~n20547 & n20549 ) | ( ~n20547 & n20550 ) | ( n20549 & n20550 ) ;
  assign n20552 = ~n20548 & n20551 ;
  assign n20553 = n20546 | n20552 ;
  assign n20554 = n20544 & n20553 ;
  assign n20555 = n20544 | n20553 ;
  assign n20556 = ~n20554 & n20555 ;
  assign n20557 = n20464 | n20467 ;
  assign n20558 = n20464 | n20466 ;
  assign n20559 = ( n20390 & n20557 ) | ( n20390 & n20558 ) | ( n20557 & n20558 ) ;
  assign n20560 = n20556 & n20559 ;
  assign n20561 = n20468 & n20556 ;
  assign n20562 = ( n20471 & n20560 ) | ( n20471 & n20561 ) | ( n20560 & n20561 ) ;
  assign n20563 = n20556 | n20559 ;
  assign n20564 = n20468 | n20556 ;
  assign n20565 = ( n20471 & n20563 ) | ( n20471 & n20564 ) | ( n20563 & n20564 ) ;
  assign n20566 = ~n20562 & n20565 ;
  assign n20567 = n20530 | n20566 ;
  assign n20568 = n20530 & n20566 ;
  assign n20569 = n20567 & ~n20568 ;
  assign n20570 = ( n20510 & n20511 ) | ( n20510 & ~n20569 ) | ( n20511 & ~n20569 ) ;
  assign n20571 = ( ~n20511 & n20569 ) | ( ~n20511 & n20570 ) | ( n20569 & n20570 ) ;
  assign n20572 = ( ~n20510 & n20570 ) | ( ~n20510 & n20571 ) | ( n20570 & n20571 ) ;
  assign n20573 = n20537 | n20548 ;
  assign n20574 = n20537 & n20548 ;
  assign n20575 = n20573 & ~n20574 ;
  assign n20576 = n20512 | n20516 ;
  assign n20577 = ( n20443 & n20512 ) | ( n20443 & n20576 ) | ( n20512 & n20576 ) ;
  assign n20578 = n20575 | n20577 ;
  assign n20579 = n20575 & n20577 ;
  assign n20580 = n20578 & ~n20579 ;
  assign n20581 = n20524 & n20580 ;
  assign n20582 = ( n20529 & n20580 ) | ( n20529 & n20581 ) | ( n20580 & n20581 ) ;
  assign n20583 = n20524 | n20580 ;
  assign n20584 = n20529 | n20583 ;
  assign n20585 = ~n20582 & n20584 ;
  assign n20586 = n7567 & n10561 ;
  assign n20587 = n7874 & n10856 ;
  assign n20588 = n20586 | n20587 ;
  assign n20589 = n8161 & n10684 ;
  assign n20590 = x63 & n20589 ;
  assign n20591 = ( x63 & ~n20588 ) | ( x63 & n20590 ) | ( ~n20588 & n20590 ) ;
  assign n20592 = x51 & n20591 ;
  assign n20593 = n20588 | n20589 ;
  assign n20594 = x52 & x62 ;
  assign n20595 = x53 & x61 ;
  assign n20596 = ( ~n20589 & n20594 ) | ( ~n20589 & n20595 ) | ( n20594 & n20595 ) ;
  assign n20597 = n20594 & n20595 ;
  assign n20598 = ( ~n20588 & n20596 ) | ( ~n20588 & n20597 ) | ( n20596 & n20597 ) ;
  assign n20599 = ~n20593 & n20598 ;
  assign n20600 = n20592 | n20599 ;
  assign n20601 = n8146 & n10975 ;
  assign n20602 = n8357 & n10370 ;
  assign n20603 = n20601 | n20602 ;
  assign n20604 = n9831 & n10013 ;
  assign n20605 = x60 & n20604 ;
  assign n20606 = ( x60 & ~n20603 ) | ( x60 & n20605 ) | ( ~n20603 & n20605 ) ;
  assign n20607 = x54 & n20606 ;
  assign n20608 = n8708 | n20436 ;
  assign n20609 = ~n20604 & n20608 ;
  assign n20610 = ~n20603 & n20609 ;
  assign n20611 = n20607 | n20610 ;
  assign n20612 = n20600 & n20611 ;
  assign n20613 = n20600 & ~n20612 ;
  assign n20614 = n20611 & ~n20612 ;
  assign n20615 = n20613 | n20614 ;
  assign n20616 = ( n20421 & n20541 ) | ( n20421 & n20553 ) | ( n20541 & n20553 ) ;
  assign n20617 = n20615 | n20616 ;
  assign n20618 = n20615 & n20616 ;
  assign n20619 = n20617 & ~n20618 ;
  assign n20620 = n20585 & n20619 ;
  assign n20621 = n20585 | n20619 ;
  assign n20622 = ~n20620 & n20621 ;
  assign n20623 = n20530 | n20562 ;
  assign n20624 = ( n20562 & n20566 ) | ( n20562 & n20623 ) | ( n20566 & n20623 ) ;
  assign n20625 = n20622 | n20624 ;
  assign n20626 = n20622 & n20624 ;
  assign n20627 = n20625 & ~n20626 ;
  assign n20628 = n20511 & n20569 ;
  assign n20629 = n20511 | n20569 ;
  assign n20630 = n20628 | n20629 ;
  assign n20631 = ( n20509 & n20628 ) | ( n20509 & n20630 ) | ( n20628 & n20630 ) ;
  assign n20632 = n20481 & n20629 ;
  assign n20633 = n20628 | n20632 ;
  assign n20634 = ( n20494 & n20630 ) | ( n20494 & n20633 ) | ( n20630 & n20633 ) ;
  assign n20635 = ( n20507 & n20628 ) | ( n20507 & n20630 ) | ( n20628 & n20630 ) ;
  assign n20636 = ( n20485 & n20634 ) | ( n20485 & n20635 ) | ( n20634 & n20635 ) ;
  assign n20637 = ( n20032 & n20631 ) | ( n20032 & n20636 ) | ( n20631 & n20636 ) ;
  assign n20638 = n20627 | n20637 ;
  assign n20639 = n20625 & n20630 ;
  assign n20640 = n20625 & n20628 ;
  assign n20641 = ( n20509 & n20639 ) | ( n20509 & n20640 ) | ( n20639 & n20640 ) ;
  assign n20642 = n20625 & n20634 ;
  assign n20643 = n20625 & n20635 ;
  assign n20644 = ( n20485 & n20642 ) | ( n20485 & n20643 ) | ( n20642 & n20643 ) ;
  assign n20645 = ( n20032 & n20641 ) | ( n20032 & n20644 ) | ( n20641 & n20644 ) ;
  assign n20646 = ~n20626 & n20645 ;
  assign n20647 = n20638 & ~n20646 ;
  assign n20648 = n20626 | n20644 ;
  assign n20649 = n20625 | n20626 ;
  assign n20650 = ( n20626 & n20630 ) | ( n20626 & n20649 ) | ( n20630 & n20649 ) ;
  assign n20651 = ( n20626 & n20628 ) | ( n20626 & n20649 ) | ( n20628 & n20649 ) ;
  assign n20652 = ( n20509 & n20650 ) | ( n20509 & n20651 ) | ( n20650 & n20651 ) ;
  assign n20653 = ( n20032 & n20648 ) | ( n20032 & n20652 ) | ( n20648 & n20652 ) ;
  assign n20654 = n8146 & n9737 ;
  assign n20655 = n8357 & n10367 ;
  assign n20656 = n20654 | n20655 ;
  assign n20657 = n10013 & n10370 ;
  assign n20658 = x61 & n20657 ;
  assign n20659 = ( x61 & ~n20656 ) | ( x61 & n20658 ) | ( ~n20656 & n20658 ) ;
  assign n20660 = x54 & n20659 ;
  assign n20661 = n20656 | n20657 ;
  assign n20662 = x55 & x60 ;
  assign n20663 = ( n15336 & ~n20657 ) | ( n15336 & n20662 ) | ( ~n20657 & n20662 ) ;
  assign n20664 = n15336 & n20662 ;
  assign n20665 = ( ~n20656 & n20663 ) | ( ~n20656 & n20664 ) | ( n20663 & n20664 ) ;
  assign n20666 = ~n20661 & n20665 ;
  assign n20667 = n20660 | n20666 ;
  assign n20668 = x53 & x62 ;
  assign n20669 = ( x58 & ~n9272 ) | ( x58 & n20668 ) | ( ~n9272 & n20668 ) ;
  assign n20670 = ( x58 & n9272 ) | ( x58 & n20668 ) | ( n9272 & n20668 ) ;
  assign n20671 = n9272 | n20668 ;
  assign n20672 = ( ~n20669 & n20670 ) | ( ~n20669 & n20671 ) | ( n20670 & n20671 ) ;
  assign n20673 = ( n9272 & n20669 ) | ( n9272 & ~n20672 ) | ( n20669 & ~n20672 ) ;
  assign n20674 = n20667 & n20673 ;
  assign n20675 = n20667 & ~n20674 ;
  assign n20676 = n20574 | n20577 ;
  assign n20677 = ( n20574 & n20575 ) | ( n20574 & n20676 ) | ( n20575 & n20676 ) ;
  assign n20678 = ~n20667 & n20673 ;
  assign n20679 = n20677 & n20678 ;
  assign n20680 = ( n20675 & n20677 ) | ( n20675 & n20679 ) | ( n20677 & n20679 ) ;
  assign n20681 = n20677 | n20678 ;
  assign n20682 = n20675 | n20681 ;
  assign n20683 = ~n20680 & n20682 ;
  assign n20684 = x52 & x63 ;
  assign n20685 = n20604 & n20684 ;
  assign n20686 = ( n20603 & n20684 ) | ( n20603 & n20685 ) | ( n20684 & n20685 ) ;
  assign n20687 = n20604 | n20684 ;
  assign n20688 = n20603 | n20687 ;
  assign n20689 = ~n20686 & n20688 ;
  assign n20690 = n20593 | n20689 ;
  assign n20691 = n20593 & n20689 ;
  assign n20692 = n20690 & ~n20691 ;
  assign n20693 = n20612 & n20692 ;
  assign n20694 = ( n20616 & n20692 ) | ( n20616 & n20693 ) | ( n20692 & n20693 ) ;
  assign n20695 = n20692 & n20693 ;
  assign n20696 = ( n20615 & n20694 ) | ( n20615 & n20695 ) | ( n20694 & n20695 ) ;
  assign n20697 = n20612 | n20692 ;
  assign n20698 = n20616 | n20697 ;
  assign n20699 = ( n20615 & n20697 ) | ( n20615 & n20698 ) | ( n20697 & n20698 ) ;
  assign n20700 = ~n20696 & n20699 ;
  assign n20701 = n20683 & n20700 ;
  assign n20702 = n20683 | n20700 ;
  assign n20703 = ~n20701 & n20702 ;
  assign n20704 = n20582 | n20619 ;
  assign n20705 = ( n20582 & n20585 ) | ( n20582 & n20704 ) | ( n20585 & n20704 ) ;
  assign n20706 = ( n20653 & n20703 ) | ( n20653 & ~n20705 ) | ( n20703 & ~n20705 ) ;
  assign n20707 = ( ~n20703 & n20705 ) | ( ~n20703 & n20706 ) | ( n20705 & n20706 ) ;
  assign n20708 = ( ~n20653 & n20706 ) | ( ~n20653 & n20707 ) | ( n20706 & n20707 ) ;
  assign n20709 = n20593 | n20686 ;
  assign n20710 = ( n20686 & n20689 ) | ( n20686 & n20709 ) | ( n20689 & n20709 ) ;
  assign n20711 = n20674 & n20710 ;
  assign n20712 = ( n20680 & n20710 ) | ( n20680 & n20711 ) | ( n20710 & n20711 ) ;
  assign n20713 = n20674 | n20710 ;
  assign n20714 = n20680 | n20713 ;
  assign n20715 = ~n20712 & n20714 ;
  assign n20716 = x58 & n20668 ;
  assign n20717 = n9272 & ~n20716 ;
  assign n20718 = n20716 | n20717 ;
  assign n20719 = n8355 & n10561 ;
  assign n20720 = x54 & x62 ;
  assign n20721 = x53 & x63 ;
  assign n20722 = n20720 | n20721 ;
  assign n20723 = ~n20719 & n20722 ;
  assign n20724 = n20718 & n20723 ;
  assign n20725 = n20718 & ~n20724 ;
  assign n20726 = ~n20718 & n20723 ;
  assign n20727 = n20725 | n20726 ;
  assign n20728 = n9737 & n12860 ;
  assign n20729 = n10013 & n10367 ;
  assign n20730 = n20728 | n20729 ;
  assign n20731 = n8903 & n10370 ;
  assign n20732 = x55 & n20731 ;
  assign n20733 = ( x55 & ~n20730 ) | ( x55 & n20732 ) | ( ~n20730 & n20732 ) ;
  assign n20734 = x61 & n20733 ;
  assign n20735 = n20730 | n20731 ;
  assign n20736 = x56 & x60 ;
  assign n20737 = ( n9829 & ~n20731 ) | ( n9829 & n20736 ) | ( ~n20731 & n20736 ) ;
  assign n20738 = n9829 & n20736 ;
  assign n20739 = ( ~n20730 & n20737 ) | ( ~n20730 & n20738 ) | ( n20737 & n20738 ) ;
  assign n20740 = ~n20735 & n20739 ;
  assign n20741 = n20734 | n20740 ;
  assign n20742 = n20661 & n20741 ;
  assign n20743 = n20741 & ~n20742 ;
  assign n20744 = n20661 & ~n20741 ;
  assign n20745 = n20727 & n20744 ;
  assign n20746 = ( n20727 & n20743 ) | ( n20727 & n20745 ) | ( n20743 & n20745 ) ;
  assign n20747 = n20727 | n20744 ;
  assign n20748 = n20743 | n20747 ;
  assign n20749 = ~n20746 & n20748 ;
  assign n20750 = n20715 & n20749 ;
  assign n20751 = n20715 | n20749 ;
  assign n20752 = ~n20750 & n20751 ;
  assign n20753 = n20683 | n20696 ;
  assign n20754 = ( n20696 & n20700 ) | ( n20696 & n20753 ) | ( n20700 & n20753 ) ;
  assign n20755 = n20752 | n20754 ;
  assign n20756 = n20752 & n20754 ;
  assign n20757 = n20755 & ~n20756 ;
  assign n20758 = n20703 & n20705 ;
  assign n20759 = n20703 | n20705 ;
  assign n20760 = n20649 & n20759 ;
  assign n20761 = n20626 & n20759 ;
  assign n20762 = ( n20630 & n20760 ) | ( n20630 & n20761 ) | ( n20760 & n20761 ) ;
  assign n20763 = n20758 | n20762 ;
  assign n20764 = n20758 | n20759 ;
  assign n20765 = ( n20651 & n20758 ) | ( n20651 & n20764 ) | ( n20758 & n20764 ) ;
  assign n20766 = ( n20509 & n20763 ) | ( n20509 & n20765 ) | ( n20763 & n20765 ) ;
  assign n20767 = ( n20626 & n20758 ) | ( n20626 & n20764 ) | ( n20758 & n20764 ) ;
  assign n20768 = ( n20644 & n20764 ) | ( n20644 & n20767 ) | ( n20764 & n20767 ) ;
  assign n20769 = ( n20032 & n20766 ) | ( n20032 & n20768 ) | ( n20766 & n20768 ) ;
  assign n20770 = n20757 | n20769 ;
  assign n20771 = n20755 & n20767 ;
  assign n20772 = n20755 & n20764 ;
  assign n20773 = ( n20644 & n20771 ) | ( n20644 & n20772 ) | ( n20771 & n20772 ) ;
  assign n20774 = n20755 & n20758 ;
  assign n20775 = ( n20755 & n20762 ) | ( n20755 & n20774 ) | ( n20762 & n20774 ) ;
  assign n20776 = ( n20651 & n20772 ) | ( n20651 & n20774 ) | ( n20772 & n20774 ) ;
  assign n20777 = ( n20481 & n20775 ) | ( n20481 & n20776 ) | ( n20775 & n20776 ) ;
  assign n20778 = n20775 | n20776 ;
  assign n20779 = ( n20502 & n20777 ) | ( n20502 & n20778 ) | ( n20777 & n20778 ) ;
  assign n20780 = ( n20032 & n20773 ) | ( n20032 & n20779 ) | ( n20773 & n20779 ) ;
  assign n20781 = ~n20756 & n20780 ;
  assign n20782 = n20770 & ~n20781 ;
  assign n20783 = n20755 | n20756 ;
  assign n20784 = ( n20756 & n20767 ) | ( n20756 & n20783 ) | ( n20767 & n20783 ) ;
  assign n20785 = ( n20756 & n20764 ) | ( n20756 & n20783 ) | ( n20764 & n20783 ) ;
  assign n20786 = ( n20644 & n20784 ) | ( n20644 & n20785 ) | ( n20784 & n20785 ) ;
  assign n20787 = n20756 | n20778 ;
  assign n20788 = n20756 | n20777 ;
  assign n20789 = ( n20502 & n20787 ) | ( n20502 & n20788 ) | ( n20787 & n20788 ) ;
  assign n20790 = ( n20032 & n20786 ) | ( n20032 & n20789 ) | ( n20786 & n20789 ) ;
  assign n20791 = n20719 & n20731 ;
  assign n20792 = ( n20719 & n20730 ) | ( n20719 & n20791 ) | ( n20730 & n20791 ) ;
  assign n20793 = ( n20724 & n20735 ) | ( n20724 & n20792 ) | ( n20735 & n20792 ) ;
  assign n20794 = n20719 | n20731 ;
  assign n20795 = n20730 | n20794 ;
  assign n20796 = n20724 | n20795 ;
  assign n20797 = ~n20793 & n20796 ;
  assign n20798 = n12770 & n15088 ;
  assign n20799 = n8146 & n10856 ;
  assign n20800 = n20798 | n20799 ;
  assign n20801 = n8903 & n10367 ;
  assign n20802 = x63 & n20801 ;
  assign n20803 = ( x63 & ~n20800 ) | ( x63 & n20802 ) | ( ~n20800 & n20802 ) ;
  assign n20804 = x54 & n20803 ;
  assign n20805 = n20800 | n20801 ;
  assign n20806 = x56 & x61 ;
  assign n20807 = ( n14647 & ~n20801 ) | ( n14647 & n20806 ) | ( ~n20801 & n20806 ) ;
  assign n20808 = n14647 & n20806 ;
  assign n20809 = ( ~n20800 & n20807 ) | ( ~n20800 & n20808 ) | ( n20807 & n20808 ) ;
  assign n20810 = ~n20805 & n20809 ;
  assign n20811 = n20804 | n20810 ;
  assign n20812 = ~n20797 & n20811 ;
  assign n20813 = n20797 & ~n20811 ;
  assign n20814 = n20812 | n20813 ;
  assign n20815 = ( x59 & x62 ) | ( x59 & ~n9831 ) | ( x62 & ~n9831 ) ;
  assign n20816 = x55 | x62 ;
  assign n20817 = ~x55 & x59 ;
  assign n20818 = ( n9831 & n20816 ) | ( n9831 & ~n20817 ) | ( n20816 & ~n20817 ) ;
  assign n20819 = ( ~x55 & x59 ) | ( ~x55 & x62 ) | ( x59 & x62 ) ;
  assign n20820 = ( x55 & n9831 ) | ( x55 & ~n20819 ) | ( n9831 & ~n20819 ) ;
  assign n20821 = ( n20815 & ~n20818 ) | ( n20815 & n20820 ) | ( ~n20818 & n20820 ) ;
  assign n20822 = n20742 | n20746 ;
  assign n20823 = ( n20814 & n20821 ) | ( n20814 & ~n20822 ) | ( n20821 & ~n20822 ) ;
  assign n20824 = ( ~n20821 & n20822 ) | ( ~n20821 & n20823 ) | ( n20822 & n20823 ) ;
  assign n20825 = ( ~n20814 & n20823 ) | ( ~n20814 & n20824 ) | ( n20823 & n20824 ) ;
  assign n20826 = n20712 | n20749 ;
  assign n20827 = ( n20712 & n20715 ) | ( n20712 & n20826 ) | ( n20715 & n20826 ) ;
  assign n20828 = ( n20790 & n20825 ) | ( n20790 & ~n20827 ) | ( n20825 & ~n20827 ) ;
  assign n20829 = ( ~n20825 & n20827 ) | ( ~n20825 & n20828 ) | ( n20827 & n20828 ) ;
  assign n20830 = ( ~n20790 & n20828 ) | ( ~n20790 & n20829 ) | ( n20828 & n20829 ) ;
  assign n20831 = n20825 & n20827 ;
  assign n20832 = n20825 | n20827 ;
  assign n20833 = n20831 | n20832 ;
  assign n20834 = ( n20789 & n20831 ) | ( n20789 & n20833 ) | ( n20831 & n20833 ) ;
  assign n20835 = n20783 & n20832 ;
  assign n20836 = n20756 & n20832 ;
  assign n20837 = ( n20767 & n20835 ) | ( n20767 & n20836 ) | ( n20835 & n20836 ) ;
  assign n20838 = n20831 | n20837 ;
  assign n20839 = ( n20785 & n20831 ) | ( n20785 & n20833 ) | ( n20831 & n20833 ) ;
  assign n20840 = ( n20644 & n20838 ) | ( n20644 & n20839 ) | ( n20838 & n20839 ) ;
  assign n20841 = ( n20032 & n20834 ) | ( n20032 & n20840 ) | ( n20834 & n20840 ) ;
  assign n20866 = n20793 | n20811 ;
  assign n20867 = ( n20793 & n20797 ) | ( n20793 & n20866 ) | ( n20797 & n20866 ) ;
  assign n20842 = x55 & n18168 ;
  assign n20843 = n9831 & ~n20842 ;
  assign n20844 = x55 & x63 ;
  assign n20845 = n20842 & n20844 ;
  assign n20846 = ( n20843 & n20844 ) | ( n20843 & n20845 ) | ( n20844 & n20845 ) ;
  assign n20847 = n20842 | n20844 ;
  assign n20848 = n20843 | n20847 ;
  assign n20849 = ~n20846 & n20848 ;
  assign n20850 = n20805 | n20849 ;
  assign n20851 = n20805 & n20849 ;
  assign n20852 = n20850 & ~n20851 ;
  assign n20853 = n10975 & n20364 ;
  assign n20854 = n8903 & n10684 ;
  assign n20855 = n20853 | n20854 ;
  assign n20856 = n9272 & n10367 ;
  assign n20857 = n20364 & n20856 ;
  assign n20858 = ( n20364 & ~n20855 ) | ( n20364 & n20857 ) | ( ~n20855 & n20857 ) ;
  assign n20859 = n20855 | n20856 ;
  assign n20860 = x57 & x61 ;
  assign n20861 = ( n10975 & ~n20856 ) | ( n10975 & n20860 ) | ( ~n20856 & n20860 ) ;
  assign n20862 = n10975 & n20860 ;
  assign n20863 = ( ~n20855 & n20861 ) | ( ~n20855 & n20862 ) | ( n20861 & n20862 ) ;
  assign n20864 = ~n20859 & n20863 ;
  assign n20865 = n20858 | n20864 ;
  assign n20868 = ( n20852 & ~n20865 ) | ( n20852 & n20867 ) | ( ~n20865 & n20867 ) ;
  assign n20869 = ( ~n20852 & n20865 ) | ( ~n20852 & n20867 ) | ( n20865 & n20867 ) ;
  assign n20870 = ( ~n20867 & n20868 ) | ( ~n20867 & n20869 ) | ( n20868 & n20869 ) ;
  assign n20871 = n20742 & n20821 ;
  assign n20872 = ( n20746 & n20821 ) | ( n20746 & n20871 ) | ( n20821 & n20871 ) ;
  assign n20873 = n20822 & ~n20872 ;
  assign n20874 = ~n20742 & n20821 ;
  assign n20875 = ~n20746 & n20874 ;
  assign n20876 = n20814 & ~n20875 ;
  assign n20877 = ~n20873 & n20876 ;
  assign n20878 = ( n20814 & n20872 ) | ( n20814 & ~n20877 ) | ( n20872 & ~n20877 ) ;
  assign n20879 = ( n20841 & n20870 ) | ( n20841 & ~n20878 ) | ( n20870 & ~n20878 ) ;
  assign n20880 = ( ~n20870 & n20878 ) | ( ~n20870 & n20879 ) | ( n20878 & n20879 ) ;
  assign n20881 = ( ~n20841 & n20879 ) | ( ~n20841 & n20880 ) | ( n20879 & n20880 ) ;
  assign n20882 = n20870 & n20872 ;
  assign n20883 = n20814 & n20870 ;
  assign n20884 = ( ~n20877 & n20882 ) | ( ~n20877 & n20883 ) | ( n20882 & n20883 ) ;
  assign n20885 = n20870 | n20872 ;
  assign n20886 = n20814 | n20870 ;
  assign n20887 = ( ~n20877 & n20885 ) | ( ~n20877 & n20886 ) | ( n20885 & n20886 ) ;
  assign n20888 = n20884 | n20887 ;
  assign n20889 = ( n20833 & n20884 ) | ( n20833 & n20888 ) | ( n20884 & n20888 ) ;
  assign n20890 = ( n20831 & n20884 ) | ( n20831 & n20888 ) | ( n20884 & n20888 ) ;
  assign n20891 = ( n20789 & n20889 ) | ( n20789 & n20890 ) | ( n20889 & n20890 ) ;
  assign n20892 = n20833 & n20887 ;
  assign n20893 = n20831 & n20887 ;
  assign n20894 = ( n20785 & n20892 ) | ( n20785 & n20893 ) | ( n20892 & n20893 ) ;
  assign n20895 = n20884 | n20894 ;
  assign n20896 = ( n20837 & n20888 ) | ( n20837 & n20890 ) | ( n20888 & n20890 ) ;
  assign n20897 = ( n20642 & n20895 ) | ( n20642 & n20896 ) | ( n20895 & n20896 ) ;
  assign n20898 = ( n20643 & n20895 ) | ( n20643 & n20896 ) | ( n20895 & n20896 ) ;
  assign n20899 = ( n20485 & n20897 ) | ( n20485 & n20898 ) | ( n20897 & n20898 ) ;
  assign n20900 = ( n20032 & n20891 ) | ( n20032 & n20899 ) | ( n20891 & n20899 ) ;
  assign n20901 = n8708 & n10856 ;
  assign n20902 = x58 & x61 ;
  assign n20903 = x56 & x63 ;
  assign n20904 = n20902 | n20903 ;
  assign n20905 = ~n20901 & n20904 ;
  assign n20906 = n20859 & n20905 ;
  assign n20907 = n20859 & ~n20906 ;
  assign n20908 = ~n20859 & n20905 ;
  assign n20909 = n20907 | n20908 ;
  assign n20910 = x57 & n9931 ;
  assign n20911 = n10370 & n20910 ;
  assign n20912 = n10370 & ~n20910 ;
  assign n20913 = n20910 | n20912 ;
  assign n20914 = x57 & x62 ;
  assign n20915 = ( x60 & ~n20910 ) | ( x60 & n20914 ) | ( ~n20910 & n20914 ) ;
  assign n20916 = x60 & n20914 ;
  assign n20917 = ( ~n20912 & n20915 ) | ( ~n20912 & n20916 ) | ( n20915 & n20916 ) ;
  assign n20918 = ~n20913 & n20917 ;
  assign n20919 = n20911 | n20918 ;
  assign n20920 = n20909 & n20919 ;
  assign n20921 = n20909 & ~n20920 ;
  assign n20922 = n20805 | n20846 ;
  assign n20923 = ( n20846 & n20849 ) | ( n20846 & n20922 ) | ( n20849 & n20922 ) ;
  assign n20924 = n20919 | n20923 ;
  assign n20925 = ( ~n20909 & n20923 ) | ( ~n20909 & n20924 ) | ( n20923 & n20924 ) ;
  assign n20926 = n20921 | n20925 ;
  assign n20927 = ( n20909 & n20919 ) | ( n20909 & n20923 ) | ( n20919 & n20923 ) ;
  assign n20928 = ~n20920 & n20927 ;
  assign n20929 = n20926 & ~n20928 ;
  assign n20930 = n20865 & n20867 ;
  assign n20931 = n20867 & ~n20930 ;
  assign n20932 = n20852 & n20865 ;
  assign n20933 = ~n20867 & n20932 ;
  assign n20934 = n20930 | n20933 ;
  assign n20935 = n20852 | n20930 ;
  assign n20936 = ( n20931 & n20934 ) | ( n20931 & n20935 ) | ( n20934 & n20935 ) ;
  assign n20937 = ( n20900 & n20929 ) | ( n20900 & ~n20936 ) | ( n20929 & ~n20936 ) ;
  assign n20938 = ( ~n20929 & n20936 ) | ( ~n20929 & n20937 ) | ( n20936 & n20937 ) ;
  assign n20939 = ( ~n20900 & n20937 ) | ( ~n20900 & n20938 ) | ( n20937 & n20938 ) ;
  assign n20940 = n20901 & n20910 ;
  assign n20941 = ( n20901 & n20912 ) | ( n20901 & n20940 ) | ( n20912 & n20940 ) ;
  assign n20942 = ( n20906 & n20913 ) | ( n20906 & n20941 ) | ( n20913 & n20941 ) ;
  assign n20943 = n20901 | n20910 ;
  assign n20944 = n20912 | n20943 ;
  assign n20945 = n20906 | n20944 ;
  assign n20946 = ~n20942 & n20945 ;
  assign n20947 = n9829 & n10856 ;
  assign n20948 = n9272 & n10561 ;
  assign n20949 = n20947 | n20948 ;
  assign n20950 = n9831 & n10684 ;
  assign n20951 = x63 & n20950 ;
  assign n20952 = ( x63 & ~n20949 ) | ( x63 & n20951 ) | ( ~n20949 & n20951 ) ;
  assign n20953 = x57 & n20952 ;
  assign n20954 = x58 & x62 ;
  assign n20955 = n9737 | n20954 ;
  assign n20956 = ~n20950 & n20955 ;
  assign n20957 = ~n20949 & n20956 ;
  assign n20958 = n20953 | n20957 ;
  assign n20959 = n20946 & n20958 ;
  assign n20960 = n20946 | n20958 ;
  assign n20961 = ~n20959 & n20960 ;
  assign n20962 = n20920 & n20961 ;
  assign n20963 = ( n20928 & n20961 ) | ( n20928 & n20962 ) | ( n20961 & n20962 ) ;
  assign n20964 = n20920 | n20961 ;
  assign n20965 = n20928 | n20964 ;
  assign n20966 = ~n20963 & n20965 ;
  assign n20967 = n20929 & n20936 ;
  assign n20968 = n20929 | n20936 ;
  assign n20969 = n20897 & n20968 ;
  assign n20970 = n20898 & n20968 ;
  assign n20971 = ( n20485 & n20969 ) | ( n20485 & n20970 ) | ( n20969 & n20970 ) ;
  assign n20972 = n20967 | n20971 ;
  assign n20973 = n20890 & n20968 ;
  assign n20974 = n20888 & n20968 ;
  assign n20975 = n20884 & n20968 ;
  assign n20976 = ( n20833 & n20974 ) | ( n20833 & n20975 ) | ( n20974 & n20975 ) ;
  assign n20977 = ( n20788 & n20973 ) | ( n20788 & n20976 ) | ( n20973 & n20976 ) ;
  assign n20978 = ( n20787 & n20973 ) | ( n20787 & n20976 ) | ( n20973 & n20976 ) ;
  assign n20979 = ( n20502 & n20977 ) | ( n20502 & n20978 ) | ( n20977 & n20978 ) ;
  assign n20980 = n20967 | n20979 ;
  assign n20981 = ( n20029 & n20972 ) | ( n20029 & n20980 ) | ( n20972 & n20980 ) ;
  assign n20982 = ( n20025 & n20972 ) | ( n20025 & n20980 ) | ( n20972 & n20980 ) ;
  assign n20983 = ( n20024 & n20972 ) | ( n20024 & n20980 ) | ( n20972 & n20980 ) ;
  assign n20984 = ( n18553 & n20982 ) | ( n18553 & n20983 ) | ( n20982 & n20983 ) ;
  assign n20985 = ( n17121 & n20981 ) | ( n17121 & n20984 ) | ( n20981 & n20984 ) ;
  assign n20986 = ( n17119 & n20981 ) | ( n17119 & n20984 ) | ( n20981 & n20984 ) ;
  assign n20987 = ( n13196 & n20985 ) | ( n13196 & n20986 ) | ( n20985 & n20986 ) ;
  assign n20988 = n20966 & ~n20987 ;
  assign n20989 = n20987 | n20988 ;
  assign n20990 = ( ~n20966 & n20988 ) | ( ~n20966 & n20989 ) | ( n20988 & n20989 ) ;
  assign n20991 = n20963 | n20965 ;
  assign n20992 = ( n20963 & n20987 ) | ( n20963 & n20991 ) | ( n20987 & n20991 ) ;
  assign n20993 = ~x60 & x61 ;
  assign n20994 = n18168 | n20993 ;
  assign n20995 = n18168 & n20993 ;
  assign n20996 = n20994 & ~n20995 ;
  assign n20997 = n19934 & n20950 ;
  assign n20998 = ( n19934 & n20949 ) | ( n19934 & n20997 ) | ( n20949 & n20997 ) ;
  assign n20999 = n19934 | n20950 ;
  assign n21000 = n20949 | n20999 ;
  assign n21001 = ~n20998 & n21000 ;
  assign n21002 = n20996 | n21001 ;
  assign n21003 = n20996 & n21001 ;
  assign n21004 = n21002 & ~n21003 ;
  assign n21005 = n20942 | n20958 ;
  assign n21006 = ( n20942 & n20946 ) | ( n20942 & n21005 ) | ( n20946 & n21005 ) ;
  assign n21007 = ( n20991 & n21004 ) | ( n20991 & ~n21006 ) | ( n21004 & ~n21006 ) ;
  assign n21008 = ( n20963 & n21004 ) | ( n20963 & ~n21006 ) | ( n21004 & ~n21006 ) ;
  assign n21009 = ( n20987 & n21007 ) | ( n20987 & n21008 ) | ( n21007 & n21008 ) ;
  assign n21010 = ( ~n21004 & n21006 ) | ( ~n21004 & n21007 ) | ( n21006 & n21007 ) ;
  assign n21011 = ( ~n21004 & n21006 ) | ( ~n21004 & n21008 ) | ( n21006 & n21008 ) ;
  assign n21012 = ( n20987 & n21010 ) | ( n20987 & n21011 ) | ( n21010 & n21011 ) ;
  assign n21013 = ( ~n20992 & n21009 ) | ( ~n20992 & n21012 ) | ( n21009 & n21012 ) ;
  assign n21014 = n9931 | n19931 ;
  assign n21015 = n10370 & n10561 ;
  assign n21016 = n21014 & ~n21015 ;
  assign n21017 = n10367 | n20995 ;
  assign n21018 = n21016 & n21017 ;
  assign n21019 = n21017 & ~n21018 ;
  assign n21020 = ( n21016 & ~n21018 ) | ( n21016 & n21019 ) | ( ~n21018 & n21019 ) ;
  assign n21021 = n20998 | n21003 ;
  assign n21022 = n21020 | n21021 ;
  assign n21023 = n21020 & n21021 ;
  assign n21024 = n21022 & ~n21023 ;
  assign n21025 = n21004 & n21006 ;
  assign n21026 = n21004 | n21006 ;
  assign n21027 = n21025 | n21026 ;
  assign n21028 = ( n20991 & n21025 ) | ( n20991 & n21027 ) | ( n21025 & n21027 ) ;
  assign n21029 = ( n20963 & n21025 ) | ( n20963 & n21027 ) | ( n21025 & n21027 ) ;
  assign n21030 = ( n20987 & n21028 ) | ( n20987 & n21029 ) | ( n21028 & n21029 ) ;
  assign n21031 = n21024 | n21030 ;
  assign n21032 = n21022 & n21027 ;
  assign n21033 = n21022 & n21025 ;
  assign n21034 = ( n20991 & n21032 ) | ( n20991 & n21033 ) | ( n21032 & n21033 ) ;
  assign n21035 = ( n20963 & n21032 ) | ( n20963 & n21033 ) | ( n21032 & n21033 ) ;
  assign n21036 = ( n20987 & n21034 ) | ( n20987 & n21035 ) | ( n21034 & n21035 ) ;
  assign n21037 = ~n21023 & n21036 ;
  assign n21038 = n21031 & ~n21037 ;
  assign n21039 = ~x61 & x62 ;
  assign n21040 = n12770 | n21039 ;
  assign n21041 = n12770 & n21039 ;
  assign n21042 = n21040 & ~n21041 ;
  assign n21043 = n21015 & n21042 ;
  assign n21044 = ( n21018 & n21042 ) | ( n21018 & n21043 ) | ( n21042 & n21043 ) ;
  assign n21045 = n21015 | n21042 ;
  assign n21046 = n21018 | n21045 ;
  assign n21047 = ~n21044 & n21046 ;
  assign n21048 = n21023 | n21035 ;
  assign n21049 = n21023 | n21034 ;
  assign n21050 = ( n20987 & n21048 ) | ( n20987 & n21049 ) | ( n21048 & n21049 ) ;
  assign n21051 = n21047 | n21050 ;
  assign n21052 = n21047 & n21050 ;
  assign n21053 = n21051 & ~n21052 ;
  assign n21054 = x62 & n10856 ;
  assign n21055 = n10684 | n10856 ;
  assign n21056 = n21041 | n21055 ;
  assign n21057 = ~n21054 & n21056 ;
  assign n21058 = n21044 | n21046 ;
  assign n21059 = ( n21044 & n21049 ) | ( n21044 & n21058 ) | ( n21049 & n21058 ) ;
  assign n21060 = ( n21023 & n21044 ) | ( n21023 & n21058 ) | ( n21044 & n21058 ) ;
  assign n21061 = ( n21035 & n21058 ) | ( n21035 & n21060 ) | ( n21058 & n21060 ) ;
  assign n21062 = ( n20987 & n21059 ) | ( n20987 & n21061 ) | ( n21059 & n21061 ) ;
  assign n21063 = n21057 & n21062 ;
  assign n21064 = n21057 | n21062 ;
  assign n21065 = ~n21063 & n21064 ;
  assign n21066 = n21056 & n21058 ;
  assign n21067 = n21054 | n21066 ;
  assign n21068 = n21044 & n21056 ;
  assign n21069 = n21054 | n21068 ;
  assign n21070 = ( n21049 & n21067 ) | ( n21049 & n21069 ) | ( n21067 & n21069 ) ;
  assign n21071 = n21056 & n21060 ;
  assign n21072 = n21054 | n21071 ;
  assign n21073 = ( n21035 & n21067 ) | ( n21035 & n21072 ) | ( n21067 & n21072 ) ;
  assign n21074 = ( n20987 & n21070 ) | ( n20987 & n21073 ) | ( n21070 & n21073 ) ;
  assign n21075 = ~x62 & x63 ;
  assign n21076 = n21074 & n21075 ;
  assign n21077 = n21075 & ~n21076 ;
  assign n21078 = ( n21074 & ~n21076 ) | ( n21074 & n21077 ) | ( ~n21076 & n21077 ) ;
  assign n21079 = ( n20981 & n21070 ) | ( n20981 & n21073 ) | ( n21070 & n21073 ) ;
  assign n21080 = x63 & n21079 ;
  assign n21081 = ( n20984 & n21070 ) | ( n20984 & n21073 ) | ( n21070 & n21073 ) ;
  assign n21082 = x63 & n21081 ;
  assign n21083 = ( n17122 & n21080 ) | ( n17122 & n21082 ) | ( n21080 & n21082 ) ;
  assign n21084 = n10561 | n21083 ;
  assign y0 = x0 ;
  assign y1 = 1'b0 ;
  assign y2 = n66 ;
  assign y3 = n70 ;
  assign y4 = n76 ;
  assign y5 = n87 ;
  assign y6 = n111 ;
  assign y7 = n132 ;
  assign y8 = n162 ;
  assign y9 = n194 ;
  assign y10 = n242 ;
  assign y11 = n298 ;
  assign y12 = n353 ;
  assign y13 = n405 ;
  assign y14 = n465 ;
  assign y15 = n538 ;
  assign y16 = n612 ;
  assign y17 = n691 ;
  assign y18 = n776 ;
  assign y19 = n866 ;
  assign y20 = n964 ;
  assign y21 = n1059 ;
  assign y22 = n1176 ;
  assign y23 = n1280 ;
  assign y24 = n1391 ;
  assign y25 = n1529 ;
  assign y26 = n1656 ;
  assign y27 = n1779 ;
  assign y28 = n1903 ;
  assign y29 = n2041 ;
  assign y30 = n2192 ;
  assign y31 = n2335 ;
  assign y32 = n2503 ;
  assign y33 = n2663 ;
  assign y34 = n2840 ;
  assign y35 = n3004 ;
  assign y36 = n3187 ;
  assign y37 = n3370 ;
  assign y38 = n3569 ;
  assign y39 = n3757 ;
  assign y40 = n3997 ;
  assign y41 = n4197 ;
  assign y42 = n4406 ;
  assign y43 = n4621 ;
  assign y44 = n4845 ;
  assign y45 = n5064 ;
  assign y46 = n5295 ;
  assign y47 = n5518 ;
  assign y48 = n5796 ;
  assign y49 = n6042 ;
  assign y50 = n6293 ;
  assign y51 = n6567 ;
  assign y52 = n6830 ;
  assign y53 = n7104 ;
  assign y54 = n7365 ;
  assign y55 = n7646 ;
  assign y56 = n7941 ;
  assign y57 = n8247 ;
  assign y58 = n8544 ;
  assign y59 = n8857 ;
  assign y60 = n9161 ;
  assign y61 = n9490 ;
  assign y62 = n9810 ;
  assign y63 = n10150 ;
  assign y64 = n10473 ;
  assign y65 = n10798 ;
  assign y66 = n11101 ;
  assign y67 = n11428 ;
  assign y68 = n11720 ;
  assign y69 = n12018 ;
  assign y70 = n12317 ;
  assign y71 = n12627 ;
  assign y72 = n12917 ;
  assign y73 = n13200 ;
  assign y74 = n13495 ;
  assign y75 = n13768 ;
  assign y76 = n14035 ;
  assign y77 = n14305 ;
  assign y78 = n14580 ;
  assign y79 = n14831 ;
  assign y80 = n15087 ;
  assign y81 = n15318 ;
  assign y82 = n15585 ;
  assign y83 = n15813 ;
  assign y84 = n16043 ;
  assign y85 = n16286 ;
  assign y86 = n16496 ;
  assign y87 = n16710 ;
  assign y88 = n16911 ;
  assign y89 = n17106 ;
  assign y90 = n17305 ;
  assign y91 = n17518 ;
  assign y92 = n17690 ;
  assign y93 = n17880 ;
  assign y94 = n18053 ;
  assign y95 = n18214 ;
  assign y96 = n18381 ;
  assign y97 = n18556 ;
  assign y98 = n18716 ;
  assign y99 = n18852 ;
  assign y100 = n19001 ;
  assign y101 = n19144 ;
  assign y102 = n19276 ;
  assign y103 = n19438 ;
  assign y104 = n19568 ;
  assign y105 = n19693 ;
  assign y106 = n19810 ;
  assign y107 = n19926 ;
  assign y108 = n20035 ;
  assign y109 = n20136 ;
  assign y110 = n20232 ;
  assign y111 = n20331 ;
  assign y112 = n20414 ;
  assign y113 = n20505 ;
  assign y114 = n20572 ;
  assign y115 = n20647 ;
  assign y116 = n20708 ;
  assign y117 = n20782 ;
  assign y118 = n20830 ;
  assign y119 = n20881 ;
  assign y120 = n20939 ;
  assign y121 = n20990 ;
  assign y122 = n21013 ;
  assign y123 = n21038 ;
  assign y124 = n21053 ;
  assign y125 = n21065 ;
  assign y126 = n21078 ;
  assign y127 = n21084 ;
endmodule
