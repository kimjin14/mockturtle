//Written by the Majority Logic Package Fri May  1 00:06:25 2015
module top (
            pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09, pi10, pi11, pi12, pi13, pi14, pi15, pi16, pi17, pi18, pi19, pi20, pi21, pi22, pi23, pi24, pi25, pi26, pi27, pi28, pi29, pi30, pi31, pi32, pi33, pi34, pi35, pi36, pi37, pi38, pi39, pi40, pi41, pi42, pi43, pi44, pi45, pi46, pi47, pi48, pi49, pi50, pi51, pi52, pi53, pi54, pi55, pi56, pi57, pi58, pi59, pi60, pi61, pi62, pi63, 
            po000, po001, po002, po003, po004, po005, po006, po007, po008, po009, po010, po011, po012, po013, po014, po015, po016, po017, po018, po019, po020, po021, po022, po023, po024, po025, po026, po027, po028, po029, po030, po031, po032, po033, po034, po035, po036, po037, po038, po039, po040, po041, po042, po043, po044, po045, po046, po047, po048, po049, po050, po051, po052, po053, po054, po055, po056, po057, po058, po059, po060, po061, po062, po063, po064, po065, po066, po067, po068, po069, po070, po071, po072, po073, po074, po075, po076, po077, po078, po079, po080, po081, po082, po083, po084, po085, po086, po087, po088, po089, po090, po091, po092, po093, po094, po095, po096, po097, po098, po099, po100, po101, po102, po103, po104, po105, po106, po107, po108, po109, po110, po111, po112, po113, po114, po115, po116, po117, po118, po119, po120, po121, po122, po123, po124, po125, po126);
input pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09, pi10, pi11, pi12, pi13, pi14, pi15, pi16, pi17, pi18, pi19, pi20, pi21, pi22, pi23, pi24, pi25, pi26, pi27, pi28, pi29, pi30, pi31, pi32, pi33, pi34, pi35, pi36, pi37, pi38, pi39, pi40, pi41, pi42, pi43, pi44, pi45, pi46, pi47, pi48, pi49, pi50, pi51, pi52, pi53, pi54, pi55, pi56, pi57, pi58, pi59, pi60, pi61, pi62, pi63;
output po000, po001, po002, po003, po004, po005, po006, po007, po008, po009, po010, po011, po012, po013, po014, po015, po016, po017, po018, po019, po020, po021, po022, po023, po024, po025, po026, po027, po028, po029, po030, po031, po032, po033, po034, po035, po036, po037, po038, po039, po040, po041, po042, po043, po044, po045, po046, po047, po048, po049, po050, po051, po052, po053, po054, po055, po056, po057, po058, po059, po060, po061, po062, po063, po064, po065, po066, po067, po068, po069, po070, po071, po072, po073, po074, po075, po076, po077, po078, po079, po080, po081, po082, po083, po084, po085, po086, po087, po088, po089, po090, po091, po092, po093, po094, po095, po096, po097, po098, po099, po100, po101, po102, po103, po104, po105, po106, po107, po108, po109, po110, po111, po112, po113, po114, po115, po116, po117, po118, po119, po120, po121, po122, po123, po124, po125, po126;
wire one, w0, w1, w2, w3, w4, w5, w6, w7, w8, w9, w10, w11, w12, w13, w14, w15, w16, w17, w18, w19, w20, w21, w22, w23, w24, w25, w26, w27, w28, w29, w30, w31, w32, w33, w34, w35, w36, w37, w38, w39, w40, w41, w42, w43, w44, w45, w46, w47, w48, w49, w50, w51, w52, w53, w54, w55, w56, w57, w58, w59, w60, w61, w62, w63, w64, w65, w66, w67, w68, w69, w70, w71, w72, w73, w74, w75, w76, w77, w78, w79, w80, w81, w82, w83, w84, w85, w86, w87, w88, w89, w90, w91, w92, w93, w94, w95, w96, w97, w98, w99, w100, w101, w102, w103, w104, w105, w106, w107, w108, w109, w110, w111, w112, w113, w114, w115, w116, w117, w118, w119, w120, w121, w122, w123, w124, w125, w126, w127, w128, w129, w130, w131, w132, w133, w134, w135, w136, w137, w138, w139, w140, w141, w142, w143, w144, w145, w146, w147, w148, w149, w150, w151, w152, w153, w154, w155, w156, w157, w158, w159, w160, w161, w162, w163, w164, w165, w166, w167, w168, w169, w170, w171, w172, w173, w174, w175, w176, w177, w178, w179, w180, w181, w182, w183, w184, w185, w186, w187, w188, w189, w190, w191, w192, w193, w194, w195, w196, w197, w198, w199, w200, w201, w202, w203, w204, w205, w206, w207, w208, w209, w210, w211, w212, w213, w214, w215, w216, w217, w218, w219, w220, w221, w222, w223, w224, w225, w226, w227, w228, w229, w230, w231, w232, w233, w234, w235, w236, w237, w238, w239, w240, w241, w242, w243, w244, w245, w246, w247, w248, w249, w250, w251, w252, w253, w254, w255, w256, w257, w258, w259, w260, w261, w262, w263, w264, w265, w266, w267, w268, w269, w270, w271, w272, w273, w274, w275, w276, w277, w278, w279, w280, w281, w282, w283, w284, w285, w286, w287, w288, w289, w290, w291, w292, w293, w294, w295, w296, w297, w298, w299, w300, w301, w302, w303, w304, w305, w306, w307, w308, w309, w310, w311, w312, w313, w314, w315, w316, w317, w318, w319, w320, w321, w322, w323, w324, w325, w326, w327, w328, w329, w330, w331, w332, w333, w334, w335, w336, w337, w338, w339, w340, w341, w342, w343, w344, w345, w346, w347, w348, w349, w350, w351, w352, w353, w354, w355, w356, w357, w358, w359, w360, w361, w362, w363, w364, w365, w366, w367, w368, w369, w370, w371, w372, w373, w374, w375, w376, w377, w378, w379, w380, w381, w382, w383, w384, w385, w386, w387, w388, w389, w390, w391, w392, w393, w394, w395, w396, w397, w398, w399, w400, w401, w402, w403, w404, w405, w406, w407, w408, w409, w410, w411, w412, w413, w414, w415, w416, w417, w418, w419, w420, w421, w422, w423, w424, w425, w426, w427, w428, w429, w430, w431, w432, w433, w434, w435, w436, w437, w438, w439, w440, w441, w442, w443, w444, w445, w446, w447, w448, w449, w450, w451, w452, w453, w454, w455, w456, w457, w458, w459, w460, w461, w462, w463, w464, w465, w466, w467, w468, w469, w470, w471, w472, w473, w474, w475, w476, w477, w478, w479, w480, w481, w482, w483, w484, w485, w486, w487, w488, w489, w490, w491, w492, w493, w494, w495, w496, w497, w498, w499, w500, w501, w502, w503, w504, w505, w506, w507, w508, w509, w510, w511, w512, w513, w514, w515, w516, w517, w518, w519, w520, w521, w522, w523, w524, w525, w526, w527, w528, w529, w530, w531, w532, w533, w534, w535, w536, w537, w538, w539, w540, w541, w542, w543, w544, w545, w546, w547, w548, w549, w550, w551, w552, w553, w554, w555, w556, w557, w558, w559, w560, w561, w562, w563, w564, w565, w566, w567, w568, w569, w570, w571, w572, w573, w574, w575, w576, w577, w578, w579, w580, w581, w582, w583, w584, w585, w586, w587, w588, w589, w590, w591, w592, w593, w594, w595, w596, w597, w598, w599, w600, w601, w602, w603, w604, w605, w606, w607, w608, w609, w610, w611, w612, w613, w614, w615, w616, w617, w618, w619, w620, w621, w622, w623, w624, w625, w626, w627, w628, w629, w630, w631, w632, w633, w634, w635, w636, w637, w638, w639, w640, w641, w642, w643, w644, w645, w646, w647, w648, w649, w650, w651, w652, w653, w654, w655, w656, w657, w658, w659, w660, w661, w662, w663, w664, w665, w666, w667, w668, w669, w670, w671, w672, w673, w674, w675, w676, w677, w678, w679, w680, w681, w682, w683, w684, w685, w686, w687, w688, w689, w690, w691, w692, w693, w694, w695, w696, w697, w698, w699, w700, w701, w702, w703, w704, w705, w706, w707, w708, w709, w710, w711, w712, w713, w714, w715, w716, w717, w718, w719, w720, w721, w722, w723, w724, w725, w726, w727, w728, w729, w730, w731, w732, w733, w734, w735, w736, w737, w738, w739, w740, w741, w742, w743, w744, w745, w746, w747, w748, w749, w750, w751, w752, w753, w754, w755, w756, w757, w758, w759, w760, w761, w762, w763, w764, w765, w766, w767, w768, w769, w770, w771, w772, w773, w774, w775, w776, w777, w778, w779, w780, w781, w782, w783, w784, w785, w786, w787, w788, w789, w790, w791, w792, w793, w794, w795, w796, w797, w798, w799, w800, w801, w802, w803, w804, w805, w806, w807, w808, w809, w810, w811, w812, w813, w814, w815, w816, w817, w818, w819, w820, w821, w822, w823, w824, w825, w826, w827, w828, w829, w830, w831, w832, w833, w834, w835, w836, w837, w838, w839, w840, w841, w842, w843, w844, w845, w846, w847, w848, w849, w850, w851, w852, w853, w854, w855, w856, w857, w858, w859, w860, w861, w862, w863, w864, w865, w866, w867, w868, w869, w870, w871, w872, w873, w874, w875, w876, w877, w878, w879, w880, w881, w882, w883, w884, w885, w886, w887, w888, w889, w890, w891, w892, w893, w894, w895, w896, w897, w898, w899, w900, w901, w902, w903, w904, w905, w906, w907, w908, w909, w910, w911, w912, w913, w914, w915, w916, w917, w918, w919, w920, w921, w922, w923, w924, w925, w926, w927, w928, w929, w930, w931, w932, w933, w934, w935, w936, w937, w938, w939, w940, w941, w942, w943, w944, w945, w946, w947, w948, w949, w950, w951, w952, w953, w954, w955, w956, w957, w958, w959, w960, w961, w962, w963, w964, w965, w966, w967, w968, w969, w970, w971, w972, w973, w974, w975, w976, w977, w978, w979, w980, w981, w982, w983, w984, w985, w986, w987, w988, w989, w990, w991, w992, w993, w994, w995, w996, w997, w998, w999, w1000, w1001, w1002, w1003, w1004, w1005, w1006, w1007, w1008, w1009, w1010, w1011, w1012, w1013, w1014, w1015, w1016, w1017, w1018, w1019, w1020, w1021, w1022, w1023, w1024, w1025, w1026, w1027, w1028, w1029, w1030, w1031, w1032, w1033, w1034, w1035, w1036, w1037, w1038, w1039, w1040, w1041, w1042, w1043, w1044, w1045, w1046, w1047, w1048, w1049, w1050, w1051, w1052, w1053, w1054, w1055, w1056, w1057, w1058, w1059, w1060, w1061, w1062, w1063, w1064, w1065, w1066, w1067, w1068, w1069, w1070, w1071, w1072, w1073, w1074, w1075, w1076, w1077, w1078, w1079, w1080, w1081, w1082, w1083, w1084, w1085, w1086, w1087, w1088, w1089, w1090, w1091, w1092, w1093, w1094, w1095, w1096, w1097, w1098, w1099, w1100, w1101, w1102, w1103, w1104, w1105, w1106, w1107, w1108, w1109, w1110, w1111, w1112, w1113, w1114, w1115, w1116, w1117, w1118, w1119, w1120, w1121, w1122, w1123, w1124, w1125, w1126, w1127, w1128, w1129, w1130, w1131, w1132, w1133, w1134, w1135, w1136, w1137, w1138, w1139, w1140, w1141, w1142, w1143, w1144, w1145, w1146, w1147, w1148, w1149, w1150, w1151, w1152, w1153, w1154, w1155, w1156, w1157, w1158, w1159, w1160, w1161, w1162, w1163, w1164, w1165, w1166, w1167, w1168, w1169, w1170, w1171, w1172, w1173, w1174, w1175, w1176, w1177, w1178, w1179, w1180, w1181, w1182, w1183, w1184, w1185, w1186, w1187, w1188, w1189, w1190, w1191, w1192, w1193, w1194, w1195, w1196, w1197, w1198, w1199, w1200, w1201, w1202, w1203, w1204, w1205, w1206, w1207, w1208, w1209, w1210, w1211, w1212, w1213, w1214, w1215, w1216, w1217, w1218, w1219, w1220, w1221, w1222, w1223, w1224, w1225, w1226, w1227, w1228, w1229, w1230, w1231, w1232, w1233, w1234, w1235, w1236, w1237, w1238, w1239, w1240, w1241, w1242, w1243, w1244, w1245, w1246, w1247, w1248, w1249, w1250, w1251, w1252, w1253, w1254, w1255, w1256, w1257, w1258, w1259, w1260, w1261, w1262, w1263, w1264, w1265, w1266, w1267, w1268, w1269, w1270, w1271, w1272, w1273, w1274, w1275, w1276, w1277, w1278, w1279, w1280, w1281, w1282, w1283, w1284, w1285, w1286, w1287, w1288, w1289, w1290, w1291, w1292, w1293, w1294, w1295, w1296, w1297, w1298, w1299, w1300, w1301, w1302, w1303, w1304, w1305, w1306, w1307, w1308, w1309, w1310, w1311, w1312, w1313, w1314, w1315, w1316, w1317, w1318, w1319, w1320, w1321, w1322, w1323, w1324, w1325, w1326, w1327, w1328, w1329, w1330, w1331, w1332, w1333, w1334, w1335, w1336, w1337, w1338, w1339, w1340, w1341, w1342, w1343, w1344, w1345, w1346, w1347, w1348, w1349, w1350, w1351, w1352, w1353, w1354, w1355, w1356, w1357, w1358, w1359, w1360, w1361, w1362, w1363, w1364, w1365, w1366, w1367, w1368, w1369, w1370, w1371, w1372, w1373, w1374, w1375, w1376, w1377, w1378, w1379, w1380, w1381, w1382, w1383, w1384, w1385, w1386, w1387, w1388, w1389, w1390, w1391, w1392, w1393, w1394, w1395, w1396, w1397, w1398, w1399, w1400, w1401, w1402, w1403, w1404, w1405, w1406, w1407, w1408, w1409, w1410, w1411, w1412, w1413, w1414, w1415, w1416, w1417, w1418, w1419, w1420, w1421, w1422, w1423, w1424, w1425, w1426, w1427, w1428, w1429, w1430, w1431, w1432, w1433, w1434, w1435, w1436, w1437, w1438, w1439, w1440, w1441, w1442, w1443, w1444, w1445, w1446, w1447, w1448, w1449, w1450, w1451, w1452, w1453, w1454, w1455, w1456, w1457, w1458, w1459, w1460, w1461, w1462, w1463, w1464, w1465, w1466, w1467, w1468, w1469, w1470, w1471, w1472, w1473, w1474, w1475, w1476, w1477, w1478, w1479, w1480, w1481, w1482, w1483, w1484, w1485, w1486, w1487, w1488, w1489, w1490, w1491, w1492, w1493, w1494, w1495, w1496, w1497, w1498, w1499, w1500, w1501, w1502, w1503, w1504, w1505, w1506, w1507, w1508, w1509, w1510, w1511, w1512, w1513, w1514, w1515, w1516, w1517, w1518, w1519, w1520, w1521, w1522, w1523, w1524, w1525, w1526, w1527, w1528, w1529, w1530, w1531, w1532, w1533, w1534, w1535, w1536, w1537, w1538, w1539, w1540, w1541, w1542, w1543, w1544, w1545, w1546, w1547, w1548, w1549, w1550, w1551, w1552, w1553, w1554, w1555, w1556, w1557, w1558, w1559, w1560, w1561, w1562, w1563, w1564, w1565, w1566, w1567, w1568, w1569, w1570, w1571, w1572, w1573, w1574, w1575, w1576, w1577, w1578, w1579, w1580, w1581, w1582, w1583, w1584, w1585, w1586, w1587, w1588, w1589, w1590, w1591, w1592, w1593, w1594, w1595, w1596, w1597, w1598, w1599, w1600, w1601, w1602, w1603, w1604, w1605, w1606, w1607, w1608, w1609, w1610, w1611, w1612, w1613, w1614, w1615, w1616, w1617, w1618, w1619, w1620, w1621, w1622, w1623, w1624, w1625, w1626, w1627, w1628, w1629, w1630, w1631, w1632, w1633, w1634, w1635, w1636, w1637, w1638, w1639, w1640, w1641, w1642, w1643, w1644, w1645, w1646, w1647, w1648, w1649, w1650, w1651, w1652, w1653, w1654, w1655, w1656, w1657, w1658, w1659, w1660, w1661, w1662, w1663, w1664, w1665, w1666, w1667, w1668, w1669, w1670, w1671, w1672, w1673, w1674, w1675, w1676, w1677, w1678, w1679, w1680, w1681, w1682, w1683, w1684, w1685, w1686, w1687, w1688, w1689, w1690, w1691, w1692, w1693, w1694, w1695, w1696, w1697, w1698, w1699, w1700, w1701, w1702, w1703, w1704, w1705, w1706, w1707, w1708, w1709, w1710, w1711, w1712, w1713, w1714, w1715, w1716, w1717, w1718, w1719, w1720, w1721, w1722, w1723, w1724, w1725, w1726, w1727, w1728, w1729, w1730, w1731, w1732, w1733, w1734, w1735, w1736, w1737, w1738, w1739, w1740, w1741, w1742, w1743, w1744, w1745, w1746, w1747, w1748, w1749, w1750, w1751, w1752, w1753, w1754, w1755, w1756, w1757, w1758, w1759, w1760, w1761, w1762, w1763, w1764, w1765, w1766, w1767, w1768, w1769, w1770, w1771, w1772, w1773, w1774, w1775, w1776, w1777, w1778, w1779, w1780, w1781, w1782, w1783, w1784, w1785, w1786, w1787, w1788, w1789, w1790, w1791, w1792, w1793, w1794, w1795, w1796, w1797, w1798, w1799, w1800, w1801, w1802, w1803, w1804, w1805, w1806, w1807, w1808, w1809, w1810, w1811, w1812, w1813, w1814, w1815, w1816, w1817, w1818, w1819, w1820, w1821, w1822, w1823, w1824, w1825, w1826, w1827, w1828, w1829, w1830, w1831, w1832, w1833, w1834, w1835, w1836, w1837, w1838, w1839, w1840, w1841, w1842, w1843, w1844, w1845, w1846, w1847, w1848, w1849, w1850, w1851, w1852, w1853, w1854, w1855, w1856, w1857, w1858, w1859, w1860, w1861, w1862, w1863, w1864, w1865, w1866, w1867, w1868, w1869, w1870, w1871, w1872, w1873, w1874, w1875, w1876, w1877, w1878, w1879, w1880, w1881, w1882, w1883, w1884, w1885, w1886, w1887, w1888, w1889, w1890, w1891, w1892, w1893, w1894, w1895, w1896, w1897, w1898, w1899, w1900, w1901, w1902, w1903, w1904, w1905, w1906, w1907, w1908, w1909, w1910, w1911, w1912, w1913, w1914, w1915, w1916, w1917, w1918, w1919, w1920, w1921, w1922, w1923, w1924, w1925, w1926, w1927, w1928, w1929, w1930, w1931, w1932, w1933, w1934, w1935, w1936, w1937, w1938, w1939, w1940, w1941, w1942, w1943, w1944, w1945, w1946, w1947, w1948, w1949, w1950, w1951, w1952, w1953, w1954, w1955, w1956, w1957, w1958, w1959, w1960, w1961, w1962, w1963, w1964, w1965, w1966, w1967, w1968, w1969, w1970, w1971, w1972, w1973, w1974, w1975, w1976, w1977, w1978, w1979, w1980, w1981, w1982, w1983, w1984, w1985, w1986, w1987, w1988, w1989, w1990, w1991, w1992, w1993, w1994, w1995, w1996, w1997, w1998, w1999, w2000, w2001, w2002, w2003, w2004, w2005, w2006, w2007, w2008, w2009, w2010, w2011, w2012, w2013, w2014, w2015, w2016, w2017, w2018, w2019, w2020, w2021, w2022, w2023, w2024, w2025, w2026, w2027, w2028, w2029, w2030, w2031, w2032, w2033, w2034, w2035, w2036, w2037, w2038, w2039, w2040, w2041, w2042, w2043, w2044, w2045, w2046, w2047, w2048, w2049, w2050, w2051, w2052, w2053, w2054, w2055, w2056, w2057, w2058, w2059, w2060, w2061, w2062, w2063, w2064, w2065, w2066, w2067, w2068, w2069, w2070, w2071, w2072, w2073, w2074, w2075, w2076, w2077, w2078, w2079, w2080, w2081, w2082, w2083, w2084, w2085, w2086, w2087, w2088, w2089, w2090, w2091, w2092, w2093, w2094, w2095, w2096, w2097, w2098, w2099, w2100, w2101, w2102, w2103, w2104, w2105, w2106, w2107, w2108, w2109, w2110, w2111, w2112, w2113, w2114, w2115, w2116, w2117, w2118, w2119, w2120, w2121, w2122, w2123, w2124, w2125, w2126, w2127, w2128, w2129, w2130, w2131, w2132, w2133, w2134, w2135, w2136, w2137, w2138, w2139, w2140, w2141, w2142, w2143, w2144, w2145, w2146, w2147, w2148, w2149, w2150, w2151, w2152, w2153, w2154, w2155, w2156, w2157, w2158, w2159, w2160, w2161, w2162, w2163, w2164, w2165, w2166, w2167, w2168, w2169, w2170, w2171, w2172, w2173, w2174, w2175, w2176, w2177, w2178, w2179, w2180, w2181, w2182, w2183, w2184, w2185, w2186, w2187, w2188, w2189, w2190, w2191, w2192, w2193, w2194, w2195, w2196, w2197, w2198, w2199, w2200, w2201, w2202, w2203, w2204, w2205, w2206, w2207, w2208, w2209, w2210, w2211, w2212, w2213, w2214, w2215, w2216, w2217, w2218, w2219, w2220, w2221, w2222, w2223, w2224, w2225, w2226, w2227, w2228, w2229, w2230, w2231, w2232, w2233, w2234, w2235, w2236, w2237, w2238, w2239, w2240, w2241, w2242, w2243, w2244, w2245, w2246, w2247, w2248, w2249, w2250, w2251, w2252, w2253, w2254, w2255, w2256, w2257, w2258, w2259, w2260, w2261, w2262, w2263, w2264, w2265, w2266, w2267, w2268, w2269, w2270, w2271, w2272, w2273, w2274, w2275, w2276, w2277, w2278, w2279, w2280, w2281, w2282, w2283, w2284, w2285, w2286, w2287, w2288, w2289, w2290, w2291, w2292, w2293, w2294, w2295, w2296, w2297, w2298, w2299, w2300, w2301, w2302, w2303, w2304, w2305, w2306, w2307, w2308, w2309, w2310, w2311, w2312, w2313, w2314, w2315, w2316, w2317, w2318, w2319, w2320, w2321, w2322, w2323, w2324, w2325, w2326, w2327, w2328, w2329, w2330, w2331, w2332, w2333, w2334, w2335, w2336, w2337, w2338, w2339, w2340, w2341, w2342, w2343, w2344, w2345, w2346, w2347, w2348, w2349, w2350, w2351, w2352, w2353, w2354, w2355, w2356, w2357, w2358, w2359, w2360, w2361, w2362, w2363, w2364, w2365, w2366, w2367, w2368, w2369, w2370, w2371, w2372, w2373, w2374, w2375, w2376, w2377, w2378, w2379, w2380, w2381, w2382, w2383, w2384, w2385, w2386, w2387, w2388, w2389, w2390, w2391, w2392, w2393, w2394, w2395, w2396, w2397, w2398, w2399, w2400, w2401, w2402, w2403, w2404, w2405, w2406, w2407, w2408, w2409, w2410, w2411, w2412, w2413, w2414, w2415, w2416, w2417, w2418, w2419, w2420, w2421, w2422, w2423, w2424, w2425, w2426, w2427, w2428, w2429, w2430, w2431, w2432, w2433, w2434, w2435, w2436, w2437, w2438, w2439, w2440, w2441, w2442, w2443, w2444, w2445, w2446, w2447, w2448, w2449, w2450, w2451, w2452, w2453, w2454, w2455, w2456, w2457, w2458, w2459, w2460, w2461, w2462, w2463, w2464, w2465, w2466, w2467, w2468, w2469, w2470, w2471, w2472, w2473, w2474, w2475, w2476, w2477, w2478, w2479, w2480, w2481, w2482, w2483, w2484, w2485, w2486, w2487, w2488, w2489, w2490, w2491, w2492, w2493, w2494, w2495, w2496, w2497, w2498, w2499, w2500, w2501, w2502, w2503, w2504, w2505, w2506, w2507, w2508, w2509, w2510, w2511, w2512, w2513, w2514, w2515, w2516, w2517, w2518, w2519, w2520, w2521, w2522, w2523, w2524, w2525, w2526, w2527, w2528, w2529, w2530, w2531, w2532, w2533, w2534, w2535, w2536, w2537, w2538, w2539, w2540, w2541, w2542, w2543, w2544, w2545, w2546, w2547, w2548, w2549, w2550, w2551, w2552, w2553, w2554, w2555, w2556, w2557, w2558, w2559, w2560, w2561, w2562, w2563, w2564, w2565, w2566, w2567, w2568, w2569, w2570, w2571, w2572, w2573, w2574, w2575, w2576, w2577, w2578, w2579, w2580, w2581, w2582, w2583, w2584, w2585, w2586, w2587, w2588, w2589, w2590, w2591, w2592, w2593, w2594, w2595, w2596, w2597, w2598, w2599, w2600, w2601, w2602, w2603, w2604, w2605, w2606, w2607, w2608, w2609, w2610, w2611, w2612, w2613, w2614, w2615, w2616, w2617, w2618, w2619, w2620, w2621, w2622, w2623, w2624, w2625, w2626, w2627, w2628, w2629, w2630, w2631, w2632, w2633, w2634, w2635, w2636, w2637, w2638, w2639, w2640, w2641, w2642, w2643, w2644, w2645, w2646, w2647, w2648, w2649, w2650, w2651, w2652, w2653, w2654, w2655, w2656, w2657, w2658, w2659, w2660, w2661, w2662, w2663, w2664, w2665, w2666, w2667, w2668, w2669, w2670, w2671, w2672, w2673, w2674, w2675, w2676, w2677, w2678, w2679, w2680, w2681, w2682, w2683, w2684, w2685, w2686, w2687, w2688, w2689, w2690, w2691, w2692, w2693, w2694, w2695, w2696, w2697, w2698, w2699, w2700, w2701, w2702, w2703, w2704, w2705, w2706, w2707, w2708, w2709, w2710, w2711, w2712, w2713, w2714, w2715, w2716, w2717, w2718, w2719, w2720, w2721, w2722, w2723, w2724, w2725, w2726, w2727, w2728, w2729, w2730, w2731, w2732, w2733, w2734, w2735, w2736, w2737, w2738, w2739, w2740, w2741, w2742, w2743, w2744, w2745, w2746, w2747, w2748, w2749, w2750, w2751, w2752, w2753, w2754, w2755, w2756, w2757, w2758, w2759, w2760, w2761, w2762, w2763, w2764, w2765, w2766, w2767, w2768, w2769, w2770, w2771, w2772, w2773, w2774, w2775, w2776, w2777, w2778, w2779, w2780, w2781, w2782, w2783, w2784, w2785, w2786, w2787, w2788, w2789, w2790, w2791, w2792, w2793, w2794, w2795, w2796, w2797, w2798, w2799, w2800, w2801, w2802, w2803, w2804, w2805, w2806, w2807, w2808, w2809, w2810, w2811, w2812, w2813, w2814, w2815, w2816, w2817, w2818, w2819, w2820, w2821, w2822, w2823, w2824, w2825, w2826, w2827, w2828, w2829, w2830, w2831, w2832, w2833, w2834, w2835, w2836, w2837, w2838, w2839, w2840, w2841, w2842, w2843, w2844, w2845, w2846, w2847, w2848, w2849, w2850, w2851, w2852, w2853, w2854, w2855, w2856, w2857, w2858, w2859, w2860, w2861, w2862, w2863, w2864, w2865, w2866, w2867, w2868, w2869, w2870, w2871, w2872, w2873, w2874, w2875, w2876, w2877, w2878, w2879, w2880, w2881, w2882, w2883, w2884, w2885, w2886, w2887, w2888, w2889, w2890, w2891, w2892, w2893, w2894, w2895, w2896, w2897, w2898, w2899, w2900, w2901, w2902, w2903, w2904, w2905, w2906, w2907, w2908, w2909, w2910, w2911, w2912, w2913, w2914, w2915, w2916, w2917, w2918, w2919, w2920, w2921, w2922, w2923, w2924, w2925, w2926, w2927, w2928, w2929, w2930, w2931, w2932, w2933, w2934, w2935, w2936, w2937, w2938, w2939, w2940, w2941, w2942, w2943, w2944, w2945, w2946, w2947, w2948, w2949, w2950, w2951, w2952, w2953, w2954, w2955, w2956, w2957, w2958, w2959, w2960, w2961, w2962, w2963, w2964, w2965, w2966, w2967, w2968, w2969, w2970, w2971, w2972, w2973, w2974, w2975, w2976, w2977, w2978, w2979, w2980, w2981, w2982, w2983, w2984, w2985, w2986, w2987, w2988, w2989, w2990, w2991, w2992, w2993, w2994, w2995, w2996, w2997, w2998, w2999, w3000, w3001, w3002, w3003, w3004, w3005, w3006, w3007, w3008, w3009, w3010, w3011, w3012, w3013, w3014, w3015, w3016, w3017, w3018, w3019, w3020, w3021, w3022, w3023, w3024, w3025, w3026, w3027, w3028, w3029, w3030, w3031, w3032, w3033, w3034, w3035, w3036, w3037, w3038, w3039, w3040, w3041, w3042, w3043, w3044, w3045, w3046, w3047, w3048, w3049, w3050, w3051, w3052, w3053, w3054, w3055, w3056, w3057, w3058, w3059, w3060, w3061, w3062, w3063, w3064, w3065, w3066, w3067, w3068, w3069, w3070, w3071, w3072, w3073, w3074, w3075, w3076, w3077, w3078, w3079, w3080, w3081, w3082, w3083, w3084, w3085, w3086, w3087, w3088, w3089, w3090, w3091, w3092, w3093, w3094, w3095, w3096, w3097, w3098, w3099, w3100, w3101, w3102, w3103, w3104, w3105, w3106, w3107, w3108, w3109, w3110, w3111, w3112, w3113, w3114, w3115, w3116, w3117, w3118, w3119, w3120, w3121, w3122, w3123, w3124, w3125, w3126, w3127, w3128, w3129, w3130, w3131, w3132, w3133, w3134, w3135, w3136, w3137, w3138, w3139, w3140, w3141, w3142, w3143, w3144, w3145, w3146, w3147, w3148, w3149, w3150, w3151, w3152, w3153, w3154, w3155, w3156, w3157, w3158, w3159, w3160, w3161, w3162, w3163, w3164, w3165, w3166, w3167, w3168, w3169, w3170, w3171, w3172, w3173, w3174, w3175, w3176, w3177, w3178, w3179, w3180, w3181, w3182, w3183, w3184, w3185, w3186, w3187, w3188, w3189, w3190, w3191, w3192, w3193, w3194, w3195, w3196, w3197, w3198, w3199, w3200, w3201, w3202, w3203, w3204, w3205, w3206, w3207, w3208, w3209, w3210, w3211, w3212, w3213, w3214, w3215, w3216, w3217, w3218, w3219, w3220, w3221, w3222, w3223, w3224, w3225, w3226, w3227, w3228, w3229, w3230, w3231, w3232, w3233, w3234, w3235, w3236, w3237, w3238, w3239, w3240, w3241, w3242, w3243, w3244, w3245, w3246, w3247, w3248, w3249, w3250, w3251, w3252, w3253, w3254, w3255, w3256, w3257, w3258, w3259, w3260, w3261, w3262, w3263, w3264, w3265, w3266, w3267, w3268, w3269, w3270, w3271, w3272, w3273, w3274, w3275, w3276, w3277, w3278, w3279, w3280, w3281, w3282, w3283, w3284, w3285, w3286, w3287, w3288, w3289, w3290, w3291, w3292, w3293, w3294, w3295, w3296, w3297, w3298, w3299, w3300, w3301, w3302, w3303, w3304, w3305, w3306, w3307, w3308, w3309, w3310, w3311, w3312, w3313, w3314, w3315, w3316, w3317, w3318, w3319, w3320, w3321, w3322, w3323, w3324, w3325, w3326, w3327, w3328, w3329, w3330, w3331, w3332, w3333, w3334, w3335, w3336, w3337, w3338, w3339, w3340, w3341, w3342, w3343, w3344, w3345, w3346, w3347, w3348, w3349, w3350, w3351, w3352, w3353, w3354, w3355, w3356, w3357, w3358, w3359, w3360, w3361, w3362, w3363, w3364, w3365, w3366, w3367, w3368, w3369, w3370, w3371, w3372, w3373, w3374, w3375, w3376, w3377, w3378, w3379, w3380, w3381, w3382, w3383, w3384, w3385, w3386, w3387, w3388, w3389, w3390, w3391, w3392, w3393, w3394, w3395, w3396, w3397, w3398, w3399, w3400, w3401, w3402, w3403, w3404, w3405, w3406, w3407, w3408, w3409, w3410, w3411, w3412, w3413, w3414, w3415, w3416, w3417, w3418, w3419, w3420, w3421, w3422, w3423, w3424, w3425, w3426, w3427, w3428, w3429, w3430, w3431, w3432, w3433, w3434, w3435, w3436, w3437, w3438, w3439, w3440, w3441, w3442, w3443, w3444, w3445, w3446, w3447, w3448, w3449, w3450, w3451, w3452, w3453, w3454, w3455, w3456, w3457, w3458, w3459, w3460, w3461, w3462, w3463, w3464, w3465, w3466, w3467, w3468, w3469, w3470, w3471, w3472, w3473, w3474, w3475, w3476, w3477, w3478, w3479, w3480, w3481, w3482, w3483, w3484, w3485, w3486, w3487, w3488, w3489, w3490, w3491, w3492, w3493, w3494, w3495, w3496, w3497, w3498, w3499, w3500, w3501, w3502, w3503, w3504, w3505, w3506, w3507, w3508, w3509, w3510, w3511, w3512, w3513, w3514, w3515, w3516, w3517, w3518, w3519, w3520, w3521, w3522, w3523, w3524, w3525, w3526, w3527, w3528, w3529, w3530, w3531, w3532, w3533, w3534, w3535, w3536, w3537, w3538, w3539, w3540, w3541, w3542, w3543, w3544, w3545, w3546, w3547, w3548, w3549, w3550, w3551, w3552, w3553, w3554, w3555, w3556, w3557, w3558, w3559, w3560, w3561, w3562, w3563, w3564, w3565, w3566, w3567, w3568, w3569, w3570, w3571, w3572, w3573, w3574, w3575, w3576, w3577, w3578, w3579, w3580, w3581, w3582, w3583, w3584, w3585, w3586, w3587, w3588, w3589, w3590, w3591, w3592, w3593, w3594, w3595, w3596, w3597, w3598, w3599, w3600, w3601, w3602, w3603, w3604, w3605, w3606, w3607, w3608, w3609, w3610, w3611, w3612, w3613, w3614, w3615, w3616, w3617, w3618, w3619, w3620, w3621, w3622, w3623, w3624, w3625, w3626, w3627, w3628, w3629, w3630, w3631, w3632, w3633, w3634, w3635, w3636, w3637, w3638, w3639, w3640, w3641, w3642, w3643, w3644, w3645, w3646, w3647, w3648, w3649, w3650, w3651, w3652, w3653, w3654, w3655, w3656, w3657, w3658, w3659, w3660, w3661, w3662, w3663, w3664, w3665, w3666, w3667, w3668, w3669, w3670, w3671, w3672, w3673, w3674, w3675, w3676, w3677, w3678, w3679, w3680, w3681, w3682, w3683, w3684, w3685, w3686, w3687, w3688, w3689, w3690, w3691, w3692, w3693, w3694, w3695, w3696, w3697, w3698, w3699, w3700, w3701, w3702, w3703, w3704, w3705, w3706, w3707, w3708, w3709, w3710, w3711, w3712, w3713, w3714, w3715, w3716, w3717, w3718, w3719, w3720, w3721, w3722, w3723, w3724, w3725, w3726, w3727, w3728, w3729, w3730, w3731, w3732, w3733, w3734, w3735, w3736, w3737, w3738, w3739, w3740, w3741, w3742, w3743, w3744, w3745, w3746, w3747, w3748, w3749, w3750, w3751, w3752, w3753, w3754, w3755, w3756, w3757, w3758, w3759, w3760, w3761, w3762, w3763, w3764, w3765, w3766, w3767, w3768, w3769, w3770, w3771, w3772, w3773, w3774, w3775, w3776, w3777, w3778, w3779, w3780, w3781, w3782, w3783, w3784, w3785, w3786, w3787, w3788, w3789, w3790, w3791, w3792, w3793, w3794, w3795, w3796, w3797, w3798, w3799, w3800, w3801, w3802, w3803, w3804, w3805, w3806, w3807, w3808, w3809, w3810, w3811, w3812, w3813, w3814, w3815, w3816, w3817, w3818, w3819, w3820, w3821, w3822, w3823, w3824, w3825, w3826, w3827, w3828, w3829, w3830, w3831, w3832, w3833, w3834, w3835, w3836, w3837, w3838, w3839, w3840, w3841, w3842, w3843, w3844, w3845, w3846, w3847, w3848, w3849, w3850, w3851, w3852, w3853, w3854, w3855, w3856, w3857, w3858, w3859, w3860, w3861, w3862, w3863, w3864, w3865, w3866, w3867, w3868, w3869, w3870, w3871, w3872, w3873, w3874, w3875, w3876, w3877, w3878, w3879, w3880, w3881, w3882, w3883, w3884, w3885, w3886, w3887, w3888, w3889, w3890, w3891, w3892, w3893, w3894, w3895, w3896, w3897, w3898, w3899, w3900, w3901, w3902, w3903, w3904, w3905, w3906, w3907, w3908, w3909, w3910, w3911, w3912, w3913, w3914, w3915, w3916, w3917, w3918, w3919, w3920, w3921, w3922, w3923, w3924, w3925, w3926, w3927, w3928, w3929, w3930, w3931, w3932, w3933, w3934, w3935, w3936, w3937, w3938, w3939, w3940, w3941, w3942, w3943, w3944, w3945, w3946, w3947, w3948, w3949, w3950, w3951, w3952, w3953, w3954, w3955, w3956, w3957, w3958, w3959, w3960, w3961, w3962, w3963, w3964, w3965, w3966, w3967, w3968, w3969, w3970, w3971, w3972, w3973, w3974, w3975, w3976, w3977, w3978, w3979, w3980, w3981, w3982, w3983, w3984, w3985, w3986, w3987, w3988, w3989, w3990, w3991, w3992, w3993, w3994, w3995, w3996, w3997, w3998, w3999, w4000, w4001, w4002, w4003, w4004, w4005, w4006, w4007, w4008, w4009, w4010, w4011, w4012, w4013, w4014, w4015, w4016, w4017, w4018, w4019, w4020, w4021, w4022, w4023, w4024, w4025, w4026, w4027, w4028, w4029, w4030, w4031, w4032, w4033, w4034, w4035, w4036, w4037, w4038, w4039, w4040, w4041, w4042, w4043, w4044, w4045, w4046, w4047, w4048, w4049, w4050, w4051, w4052, w4053, w4054, w4055, w4056, w4057, w4058, w4059, w4060, w4061, w4062, w4063, w4064, w4065, w4066, w4067, w4068, w4069, w4070, w4071, w4072, w4073, w4074, w4075, w4076, w4077, w4078, w4079, w4080, w4081, w4082, w4083, w4084, w4085, w4086, w4087, w4088, w4089, w4090, w4091, w4092, w4093, w4094, w4095, w4096, w4097, w4098, w4099, w4100, w4101, w4102, w4103, w4104, w4105, w4106, w4107, w4108, w4109, w4110, w4111, w4112, w4113, w4114, w4115, w4116, w4117, w4118, w4119, w4120, w4121, w4122, w4123, w4124, w4125, w4126, w4127, w4128, w4129, w4130, w4131, w4132, w4133, w4134, w4135, w4136, w4137, w4138, w4139, w4140, w4141, w4142, w4143, w4144, w4145, w4146, w4147, w4148, w4149, w4150, w4151, w4152, w4153, w4154, w4155, w4156, w4157, w4158, w4159, w4160, w4161, w4162, w4163, w4164, w4165, w4166, w4167, w4168, w4169, w4170, w4171, w4172, w4173, w4174, w4175, w4176, w4177, w4178, w4179, w4180, w4181, w4182, w4183, w4184, w4185, w4186, w4187, w4188, w4189, w4190, w4191, w4192, w4193, w4194, w4195, w4196, w4197, w4198, w4199, w4200, w4201, w4202, w4203, w4204, w4205, w4206, w4207, w4208, w4209, w4210, w4211, w4212, w4213, w4214, w4215, w4216, w4217, w4218, w4219, w4220, w4221, w4222, w4223, w4224, w4225, w4226, w4227, w4228, w4229, w4230, w4231, w4232, w4233, w4234, w4235, w4236, w4237, w4238, w4239, w4240, w4241, w4242, w4243, w4244, w4245, w4246, w4247, w4248, w4249, w4250, w4251, w4252, w4253, w4254, w4255, w4256, w4257, w4258, w4259, w4260, w4261, w4262, w4263, w4264, w4265, w4266, w4267, w4268, w4269, w4270, w4271, w4272, w4273, w4274, w4275, w4276, w4277, w4278, w4279, w4280, w4281, w4282, w4283, w4284, w4285, w4286, w4287, w4288, w4289, w4290, w4291, w4292, w4293, w4294, w4295, w4296, w4297, w4298, w4299, w4300, w4301, w4302, w4303, w4304, w4305, w4306, w4307, w4308, w4309, w4310, w4311, w4312, w4313, w4314, w4315, w4316, w4317, w4318, w4319, w4320, w4321, w4322, w4323, w4324, w4325, w4326, w4327, w4328, w4329, w4330, w4331, w4332, w4333, w4334, w4335, w4336, w4337, w4338, w4339, w4340, w4341, w4342, w4343, w4344, w4345, w4346, w4347, w4348, w4349, w4350, w4351, w4352, w4353, w4354, w4355, w4356, w4357, w4358, w4359, w4360, w4361, w4362, w4363, w4364, w4365, w4366, w4367, w4368, w4369, w4370, w4371, w4372, w4373, w4374, w4375, w4376, w4377, w4378, w4379, w4380, w4381, w4382, w4383, w4384, w4385, w4386, w4387, w4388, w4389, w4390, w4391, w4392, w4393, w4394, w4395, w4396, w4397, w4398, w4399, w4400, w4401, w4402, w4403, w4404, w4405, w4406, w4407, w4408, w4409, w4410, w4411, w4412, w4413, w4414, w4415, w4416, w4417, w4418, w4419, w4420, w4421, w4422, w4423, w4424, w4425, w4426, w4427, w4428, w4429, w4430, w4431, w4432, w4433, w4434, w4435, w4436, w4437, w4438, w4439, w4440, w4441, w4442, w4443, w4444, w4445, w4446, w4447, w4448, w4449, w4450, w4451, w4452, w4453, w4454, w4455, w4456, w4457, w4458, w4459, w4460, w4461, w4462, w4463, w4464, w4465, w4466, w4467, w4468, w4469, w4470, w4471, w4472, w4473, w4474, w4475, w4476, w4477, w4478, w4479, w4480, w4481, w4482, w4483, w4484, w4485, w4486, w4487, w4488, w4489, w4490, w4491, w4492, w4493, w4494, w4495, w4496, w4497, w4498, w4499, w4500, w4501, w4502, w4503, w4504, w4505, w4506, w4507, w4508, w4509, w4510, w4511, w4512, w4513, w4514, w4515, w4516, w4517, w4518, w4519, w4520, w4521, w4522, w4523, w4524, w4525, w4526, w4527, w4528, w4529, w4530, w4531, w4532, w4533, w4534, w4535, w4536, w4537, w4538, w4539, w4540, w4541, w4542, w4543, w4544, w4545, w4546, w4547, w4548, w4549, w4550, w4551, w4552, w4553, w4554, w4555, w4556, w4557, w4558, w4559, w4560, w4561, w4562, w4563, w4564, w4565, w4566, w4567, w4568, w4569, w4570, w4571, w4572, w4573, w4574, w4575, w4576, w4577, w4578, w4579, w4580, w4581, w4582, w4583, w4584, w4585, w4586, w4587, w4588, w4589, w4590, w4591, w4592, w4593, w4594, w4595, w4596, w4597, w4598, w4599, w4600, w4601, w4602, w4603, w4604, w4605, w4606, w4607, w4608, w4609, w4610, w4611, w4612, w4613, w4614, w4615, w4616, w4617, w4618, w4619, w4620, w4621, w4622, w4623, w4624, w4625, w4626, w4627, w4628, w4629, w4630, w4631, w4632, w4633, w4634, w4635, w4636, w4637, w4638, w4639, w4640, w4641, w4642, w4643, w4644, w4645, w4646, w4647, w4648, w4649, w4650, w4651, w4652, w4653, w4654, w4655, w4656, w4657, w4658, w4659, w4660, w4661, w4662, w4663, w4664, w4665, w4666, w4667, w4668, w4669, w4670, w4671, w4672, w4673, w4674, w4675, w4676, w4677, w4678, w4679, w4680, w4681, w4682, w4683, w4684, w4685, w4686, w4687, w4688, w4689, w4690, w4691, w4692, w4693, w4694, w4695, w4696, w4697, w4698, w4699, w4700, w4701, w4702, w4703, w4704, w4705, w4706, w4707, w4708, w4709, w4710, w4711, w4712, w4713, w4714, w4715, w4716, w4717, w4718, w4719, w4720, w4721, w4722, w4723, w4724, w4725, w4726, w4727, w4728, w4729, w4730, w4731, w4732, w4733, w4734, w4735, w4736, w4737, w4738, w4739, w4740, w4741, w4742, w4743, w4744, w4745, w4746, w4747, w4748, w4749, w4750, w4751, w4752, w4753, w4754, w4755, w4756, w4757, w4758, w4759, w4760, w4761, w4762, w4763, w4764, w4765, w4766, w4767, w4768, w4769, w4770, w4771, w4772, w4773, w4774, w4775, w4776, w4777, w4778, w4779, w4780, w4781, w4782, w4783, w4784, w4785, w4786, w4787, w4788, w4789, w4790, w4791, w4792, w4793, w4794, w4795, w4796, w4797, w4798, w4799, w4800, w4801, w4802, w4803, w4804, w4805, w4806, w4807, w4808, w4809, w4810, w4811, w4812, w4813, w4814, w4815, w4816, w4817, w4818, w4819, w4820, w4821, w4822, w4823, w4824, w4825, w4826, w4827, w4828, w4829, w4830, w4831, w4832, w4833, w4834, w4835, w4836, w4837, w4838, w4839, w4840, w4841, w4842, w4843, w4844, w4845, w4846, w4847, w4848, w4849, w4850, w4851, w4852, w4853, w4854, w4855, w4856, w4857, w4858, w4859, w4860, w4861, w4862, w4863, w4864, w4865, w4866, w4867, w4868, w4869, w4870, w4871, w4872, w4873, w4874, w4875, w4876, w4877, w4878, w4879, w4880, w4881, w4882, w4883, w4884, w4885, w4886, w4887, w4888, w4889, w4890, w4891, w4892, w4893, w4894, w4895, w4896, w4897, w4898, w4899, w4900, w4901, w4902, w4903, w4904, w4905, w4906, w4907, w4908, w4909, w4910, w4911, w4912, w4913, w4914, w4915, w4916, w4917, w4918, w4919, w4920, w4921, w4922, w4923, w4924, w4925, w4926, w4927, w4928, w4929, w4930, w4931, w4932, w4933, w4934, w4935, w4936, w4937, w4938, w4939, w4940, w4941, w4942, w4943, w4944, w4945, w4946, w4947, w4948, w4949, w4950, w4951, w4952, w4953, w4954, w4955, w4956, w4957, w4958, w4959, w4960, w4961, w4962, w4963, w4964, w4965, w4966, w4967, w4968, w4969, w4970, w4971, w4972, w4973, w4974, w4975, w4976, w4977, w4978, w4979, w4980, w4981, w4982, w4983, w4984, w4985, w4986, w4987, w4988, w4989, w4990, w4991, w4992, w4993, w4994, w4995, w4996, w4997, w4998, w4999, w5000, w5001, w5002, w5003, w5004, w5005, w5006, w5007, w5008, w5009, w5010, w5011, w5012, w5013, w5014, w5015, w5016, w5017, w5018, w5019, w5020, w5021, w5022, w5023, w5024, w5025, w5026, w5027, w5028, w5029, w5030, w5031, w5032, w5033, w5034, w5035, w5036, w5037, w5038, w5039, w5040, w5041, w5042, w5043, w5044, w5045, w5046, w5047, w5048, w5049, w5050, w5051, w5052, w5053, w5054, w5055, w5056, w5057, w5058, w5059, w5060, w5061, w5062, w5063, w5064, w5065, w5066, w5067, w5068, w5069, w5070, w5071, w5072, w5073, w5074, w5075, w5076, w5077, w5078, w5079, w5080, w5081, w5082, w5083, w5084, w5085, w5086, w5087, w5088, w5089, w5090, w5091, w5092, w5093, w5094, w5095, w5096, w5097, w5098, w5099, w5100, w5101, w5102, w5103, w5104, w5105, w5106, w5107, w5108, w5109, w5110, w5111, w5112, w5113, w5114, w5115, w5116, w5117, w5118, w5119, w5120, w5121, w5122, w5123, w5124, w5125, w5126, w5127, w5128, w5129, w5130, w5131, w5132, w5133, w5134, w5135, w5136, w5137, w5138, w5139, w5140, w5141, w5142, w5143, w5144, w5145, w5146, w5147, w5148, w5149, w5150, w5151, w5152, w5153, w5154, w5155, w5156, w5157, w5158, w5159, w5160, w5161, w5162, w5163, w5164, w5165, w5166, w5167, w5168, w5169, w5170, w5171, w5172, w5173, w5174, w5175, w5176, w5177, w5178, w5179, w5180, w5181, w5182, w5183, w5184, w5185, w5186, w5187, w5188, w5189, w5190, w5191, w5192, w5193, w5194, w5195, w5196, w5197, w5198, w5199, w5200, w5201, w5202, w5203, w5204, w5205, w5206, w5207, w5208, w5209, w5210, w5211, w5212, w5213, w5214, w5215, w5216, w5217, w5218, w5219, w5220, w5221, w5222, w5223, w5224, w5225, w5226, w5227, w5228, w5229, w5230, w5231, w5232, w5233, w5234, w5235, w5236, w5237, w5238, w5239, w5240, w5241, w5242, w5243, w5244, w5245, w5246, w5247, w5248, w5249, w5250, w5251, w5252, w5253, w5254, w5255, w5256, w5257, w5258, w5259, w5260, w5261, w5262, w5263, w5264, w5265, w5266, w5267, w5268, w5269, w5270, w5271, w5272, w5273, w5274, w5275, w5276, w5277, w5278, w5279, w5280, w5281, w5282, w5283, w5284, w5285, w5286, w5287, w5288, w5289, w5290, w5291, w5292, w5293, w5294, w5295, w5296, w5297, w5298, w5299, w5300, w5301, w5302, w5303, w5304, w5305, w5306, w5307, w5308, w5309, w5310, w5311, w5312, w5313, w5314, w5315, w5316, w5317, w5318, w5319, w5320, w5321, w5322, w5323, w5324, w5325, w5326, w5327, w5328, w5329, w5330, w5331, w5332, w5333, w5334, w5335, w5336, w5337, w5338, w5339, w5340, w5341, w5342, w5343, w5344, w5345, w5346, w5347, w5348, w5349, w5350, w5351, w5352, w5353, w5354, w5355, w5356, w5357, w5358, w5359, w5360, w5361, w5362, w5363, w5364, w5365, w5366, w5367, w5368, w5369, w5370, w5371, w5372, w5373, w5374, w5375, w5376, w5377, w5378, w5379, w5380, w5381, w5382, w5383, w5384, w5385, w5386, w5387, w5388, w5389, w5390, w5391, w5392, w5393, w5394, w5395, w5396, w5397, w5398, w5399, w5400, w5401, w5402, w5403, w5404, w5405, w5406, w5407, w5408, w5409, w5410, w5411, w5412, w5413, w5414, w5415, w5416, w5417, w5418, w5419, w5420, w5421, w5422, w5423, w5424, w5425, w5426, w5427, w5428, w5429, w5430, w5431, w5432, w5433, w5434, w5435, w5436, w5437, w5438, w5439, w5440, w5441, w5442, w5443, w5444, w5445, w5446, w5447, w5448, w5449, w5450, w5451, w5452, w5453, w5454, w5455, w5456, w5457, w5458, w5459, w5460, w5461, w5462, w5463, w5464, w5465, w5466, w5467, w5468, w5469, w5470, w5471, w5472, w5473, w5474, w5475, w5476, w5477, w5478, w5479, w5480, w5481, w5482, w5483, w5484, w5485, w5486, w5487, w5488, w5489, w5490, w5491, w5492, w5493, w5494, w5495, w5496, w5497, w5498, w5499, w5500, w5501, w5502, w5503, w5504, w5505, w5506, w5507, w5508, w5509, w5510, w5511, w5512, w5513, w5514, w5515, w5516, w5517, w5518, w5519, w5520, w5521, w5522, w5523, w5524, w5525, w5526, w5527, w5528, w5529, w5530, w5531, w5532, w5533, w5534, w5535, w5536, w5537, w5538, w5539, w5540, w5541, w5542, w5543, w5544, w5545, w5546, w5547, w5548, w5549, w5550, w5551, w5552, w5553, w5554, w5555, w5556, w5557, w5558, w5559, w5560, w5561, w5562, w5563, w5564, w5565, w5566, w5567, w5568, w5569, w5570, w5571, w5572, w5573, w5574, w5575, w5576, w5577, w5578, w5579, w5580, w5581, w5582, w5583, w5584, w5585, w5586, w5587, w5588, w5589, w5590, w5591, w5592, w5593, w5594, w5595, w5596, w5597, w5598, w5599, w5600, w5601, w5602, w5603, w5604, w5605, w5606, w5607, w5608, w5609, w5610, w5611, w5612, w5613, w5614, w5615, w5616, w5617, w5618, w5619, w5620, w5621, w5622, w5623, w5624, w5625, w5626, w5627, w5628, w5629, w5630, w5631, w5632, w5633, w5634, w5635, w5636, w5637, w5638, w5639, w5640, w5641, w5642, w5643, w5644, w5645, w5646, w5647, w5648, w5649, w5650, w5651, w5652, w5653, w5654, w5655, w5656, w5657, w5658, w5659, w5660, w5661, w5662, w5663, w5664, w5665, w5666, w5667, w5668, w5669, w5670, w5671, w5672, w5673, w5674, w5675, w5676, w5677, w5678, w5679, w5680, w5681, w5682, w5683, w5684, w5685, w5686, w5687, w5688, w5689, w5690, w5691, w5692, w5693, w5694, w5695, w5696, w5697, w5698, w5699, w5700, w5701, w5702, w5703, w5704, w5705, w5706, w5707, w5708, w5709, w5710, w5711, w5712, w5713, w5714, w5715, w5716, w5717, w5718, w5719, w5720, w5721, w5722, w5723, w5724, w5725, w5726, w5727, w5728, w5729, w5730, w5731, w5732, w5733, w5734, w5735, w5736, w5737, w5738, w5739, w5740, w5741, w5742, w5743, w5744, w5745, w5746, w5747, w5748, w5749, w5750, w5751, w5752, w5753, w5754, w5755, w5756, w5757, w5758, w5759, w5760, w5761, w5762, w5763, w5764, w5765, w5766, w5767, w5768, w5769, w5770, w5771, w5772, w5773, w5774, w5775, w5776, w5777, w5778, w5779, w5780, w5781, w5782, w5783, w5784, w5785, w5786, w5787, w5788, w5789, w5790, w5791, w5792, w5793, w5794, w5795, w5796, w5797, w5798, w5799, w5800, w5801, w5802, w5803, w5804, w5805, w5806, w5807, w5808, w5809, w5810, w5811, w5812, w5813, w5814, w5815, w5816, w5817, w5818, w5819, w5820, w5821, w5822, w5823, w5824, w5825, w5826, w5827, w5828, w5829, w5830, w5831, w5832, w5833, w5834, w5835, w5836, w5837, w5838, w5839, w5840, w5841, w5842, w5843, w5844, w5845, w5846, w5847, w5848, w5849, w5850, w5851, w5852, w5853, w5854, w5855, w5856, w5857, w5858, w5859, w5860, w5861, w5862, w5863, w5864, w5865, w5866, w5867, w5868, w5869, w5870, w5871, w5872, w5873, w5874, w5875, w5876, w5877, w5878, w5879, w5880, w5881, w5882, w5883, w5884, w5885, w5886, w5887, w5888, w5889, w5890, w5891, w5892, w5893, w5894, w5895, w5896, w5897, w5898, w5899, w5900, w5901, w5902, w5903, w5904, w5905, w5906, w5907, w5908, w5909, w5910, w5911, w5912, w5913, w5914, w5915, w5916, w5917, w5918, w5919, w5920, w5921, w5922, w5923, w5924, w5925, w5926, w5927, w5928, w5929, w5930, w5931, w5932, w5933, w5934, w5935, w5936, w5937, w5938, w5939, w5940, w5941, w5942, w5943, w5944, w5945, w5946, w5947, w5948, w5949, w5950, w5951, w5952, w5953, w5954, w5955, w5956, w5957, w5958, w5959, w5960, w5961, w5962, w5963, w5964, w5965, w5966, w5967, w5968, w5969, w5970, w5971, w5972, w5973, w5974, w5975, w5976, w5977, w5978, w5979, w5980, w5981, w5982, w5983, w5984, w5985, w5986, w5987, w5988, w5989, w5990, w5991, w5992, w5993, w5994, w5995, w5996, w5997, w5998, w5999, w6000, w6001, w6002, w6003, w6004, w6005, w6006, w6007, w6008, w6009, w6010, w6011, w6012, w6013, w6014, w6015, w6016, w6017, w6018, w6019, w6020, w6021, w6022, w6023, w6024, w6025, w6026, w6027, w6028, w6029, w6030, w6031, w6032, w6033, w6034, w6035, w6036, w6037, w6038, w6039, w6040, w6041, w6042, w6043, w6044, w6045, w6046, w6047, w6048, w6049, w6050, w6051, w6052, w6053, w6054, w6055, w6056, w6057, w6058, w6059, w6060, w6061, w6062, w6063, w6064, w6065, w6066, w6067, w6068, w6069, w6070, w6071, w6072, w6073, w6074, w6075, w6076, w6077, w6078, w6079, w6080, w6081, w6082, w6083, w6084, w6085, w6086, w6087, w6088, w6089, w6090, w6091, w6092, w6093, w6094, w6095, w6096, w6097, w6098, w6099, w6100, w6101, w6102, w6103, w6104, w6105, w6106, w6107, w6108, w6109, w6110, w6111, w6112, w6113, w6114, w6115, w6116, w6117, w6118, w6119, w6120, w6121, w6122, w6123, w6124, w6125, w6126, w6127, w6128, w6129, w6130, w6131, w6132, w6133, w6134, w6135, w6136, w6137, w6138, w6139, w6140, w6141, w6142, w6143, w6144, w6145, w6146, w6147, w6148, w6149, w6150, w6151, w6152, w6153, w6154, w6155, w6156, w6157, w6158, w6159, w6160, w6161, w6162, w6163, w6164, w6165, w6166, w6167, w6168, w6169, w6170, w6171, w6172, w6173, w6174, w6175, w6176, w6177, w6178, w6179, w6180, w6181, w6182, w6183, w6184, w6185, w6186, w6187, w6188, w6189, w6190, w6191, w6192, w6193, w6194, w6195, w6196, w6197, w6198, w6199, w6200, w6201, w6202, w6203, w6204, w6205, w6206, w6207, w6208, w6209, w6210, w6211, w6212, w6213, w6214, w6215, w6216, w6217, w6218, w6219, w6220, w6221, w6222, w6223, w6224, w6225, w6226, w6227, w6228, w6229, w6230, w6231, w6232, w6233, w6234, w6235, w6236, w6237, w6238, w6239, w6240, w6241, w6242, w6243, w6244, w6245, w6246, w6247, w6248, w6249, w6250, w6251, w6252, w6253, w6254, w6255, w6256, w6257, w6258, w6259, w6260, w6261, w6262, w6263, w6264, w6265, w6266, w6267, w6268, w6269, w6270, w6271, w6272, w6273, w6274, w6275, w6276, w6277, w6278, w6279, w6280, w6281, w6282, w6283, w6284, w6285, w6286, w6287, w6288, w6289, w6290, w6291, w6292, w6293, w6294, w6295, w6296, w6297, w6298, w6299, w6300, w6301, w6302, w6303, w6304, w6305, w6306, w6307, w6308, w6309, w6310, w6311, w6312, w6313, w6314, w6315, w6316, w6317, w6318, w6319, w6320, w6321, w6322, w6323, w6324, w6325, w6326, w6327, w6328, w6329, w6330, w6331, w6332, w6333, w6334, w6335, w6336, w6337, w6338, w6339, w6340, w6341, w6342, w6343, w6344, w6345, w6346, w6347, w6348, w6349, w6350, w6351, w6352, w6353, w6354, w6355, w6356, w6357, w6358, w6359, w6360, w6361, w6362, w6363, w6364, w6365, w6366, w6367, w6368, w6369, w6370, w6371, w6372, w6373, w6374, w6375, w6376, w6377, w6378, w6379, w6380, w6381, w6382, w6383, w6384, w6385, w6386, w6387, w6388, w6389, w6390, w6391, w6392, w6393, w6394, w6395, w6396, w6397, w6398, w6399, w6400, w6401, w6402, w6403, w6404, w6405, w6406, w6407, w6408, w6409, w6410, w6411, w6412, w6413, w6414, w6415, w6416, w6417, w6418, w6419, w6420, w6421, w6422, w6423, w6424, w6425, w6426, w6427, w6428, w6429, w6430, w6431, w6432, w6433, w6434, w6435, w6436, w6437, w6438, w6439, w6440, w6441, w6442, w6443, w6444, w6445, w6446, w6447, w6448, w6449, w6450, w6451, w6452, w6453, w6454, w6455, w6456, w6457, w6458, w6459, w6460, w6461, w6462, w6463, w6464, w6465, w6466, w6467, w6468, w6469, w6470, w6471, w6472, w6473, w6474, w6475, w6476, w6477, w6478, w6479, w6480, w6481, w6482, w6483, w6484, w6485, w6486, w6487, w6488, w6489, w6490, w6491, w6492, w6493, w6494, w6495, w6496, w6497, w6498, w6499, w6500, w6501, w6502, w6503, w6504, w6505, w6506, w6507, w6508, w6509, w6510, w6511, w6512, w6513, w6514, w6515, w6516, w6517, w6518, w6519, w6520, w6521, w6522, w6523, w6524, w6525, w6526, w6527, w6528, w6529, w6530, w6531, w6532, w6533, w6534, w6535, w6536, w6537, w6538, w6539, w6540, w6541, w6542, w6543, w6544, w6545, w6546, w6547, w6548, w6549, w6550, w6551, w6552, w6553, w6554, w6555, w6556, w6557, w6558, w6559, w6560, w6561, w6562, w6563, w6564, w6565, w6566, w6567, w6568, w6569, w6570, w6571, w6572, w6573, w6574, w6575, w6576, w6577, w6578, w6579, w6580, w6581, w6582, w6583, w6584, w6585, w6586, w6587, w6588, w6589, w6590, w6591, w6592, w6593, w6594, w6595, w6596, w6597, w6598, w6599, w6600, w6601, w6602, w6603, w6604, w6605, w6606, w6607, w6608, w6609, w6610, w6611, w6612, w6613, w6614, w6615, w6616, w6617, w6618, w6619, w6620, w6621, w6622, w6623, w6624, w6625, w6626, w6627, w6628, w6629, w6630, w6631, w6632, w6633, w6634, w6635, w6636, w6637, w6638, w6639, w6640, w6641, w6642, w6643, w6644, w6645, w6646, w6647, w6648, w6649, w6650, w6651, w6652, w6653, w6654, w6655, w6656, w6657, w6658, w6659, w6660, w6661, w6662, w6663, w6664, w6665, w6666, w6667, w6668, w6669, w6670, w6671, w6672, w6673, w6674, w6675, w6676, w6677, w6678, w6679, w6680, w6681, w6682, w6683, w6684, w6685, w6686, w6687, w6688, w6689, w6690, w6691, w6692, w6693, w6694, w6695, w6696, w6697, w6698, w6699, w6700, w6701, w6702, w6703, w6704, w6705, w6706, w6707, w6708, w6709, w6710, w6711, w6712, w6713, w6714, w6715, w6716, w6717, w6718, w6719, w6720, w6721, w6722, w6723, w6724, w6725, w6726, w6727, w6728, w6729, w6730, w6731, w6732, w6733, w6734, w6735, w6736, w6737, w6738, w6739, w6740, w6741, w6742, w6743, w6744, w6745, w6746, w6747, w6748, w6749, w6750, w6751, w6752, w6753, w6754, w6755, w6756, w6757, w6758, w6759, w6760, w6761, w6762, w6763, w6764, w6765, w6766, w6767, w6768, w6769, w6770, w6771, w6772, w6773, w6774, w6775, w6776, w6777, w6778, w6779, w6780, w6781, w6782, w6783, w6784, w6785, w6786, w6787, w6788, w6789, w6790, w6791, w6792, w6793, w6794, w6795, w6796, w6797, w6798, w6799, w6800, w6801, w6802, w6803, w6804, w6805, w6806, w6807, w6808, w6809, w6810, w6811, w6812, w6813, w6814, w6815, w6816, w6817, w6818, w6819, w6820, w6821, w6822, w6823, w6824, w6825, w6826, w6827, w6828, w6829, w6830, w6831, w6832, w6833, w6834, w6835, w6836, w6837, w6838, w6839, w6840, w6841, w6842, w6843, w6844, w6845, w6846, w6847, w6848, w6849, w6850, w6851, w6852, w6853, w6854, w6855, w6856, w6857, w6858, w6859, w6860, w6861, w6862, w6863, w6864, w6865, w6866, w6867, w6868, w6869, w6870, w6871, w6872, w6873, w6874, w6875, w6876, w6877, w6878, w6879, w6880, w6881, w6882, w6883, w6884, w6885, w6886, w6887, w6888, w6889, w6890, w6891, w6892, w6893, w6894, w6895, w6896, w6897, w6898, w6899, w6900, w6901, w6902, w6903, w6904, w6905, w6906, w6907, w6908, w6909, w6910, w6911, w6912, w6913, w6914, w6915, w6916, w6917, w6918, w6919, w6920, w6921, w6922, w6923, w6924, w6925, w6926, w6927, w6928, w6929, w6930, w6931, w6932, w6933, w6934, w6935, w6936, w6937, w6938, w6939, w6940, w6941, w6942, w6943, w6944, w6945, w6946, w6947, w6948, w6949, w6950, w6951, w6952, w6953, w6954, w6955, w6956, w6957, w6958, w6959, w6960, w6961, w6962, w6963, w6964, w6965, w6966, w6967, w6968, w6969, w6970, w6971, w6972, w6973, w6974, w6975, w6976, w6977, w6978, w6979, w6980, w6981, w6982, w6983, w6984, w6985, w6986, w6987, w6988, w6989, w6990, w6991, w6992, w6993, w6994, w6995, w6996, w6997, w6998, w6999, w7000, w7001, w7002, w7003, w7004, w7005, w7006, w7007, w7008, w7009, w7010, w7011, w7012, w7013, w7014, w7015, w7016, w7017, w7018, w7019, w7020, w7021, w7022, w7023, w7024, w7025, w7026, w7027, w7028, w7029, w7030, w7031, w7032, w7033, w7034, w7035, w7036, w7037, w7038, w7039, w7040, w7041, w7042, w7043, w7044, w7045, w7046, w7047, w7048, w7049, w7050, w7051, w7052, w7053, w7054, w7055, w7056, w7057, w7058, w7059, w7060, w7061, w7062, w7063, w7064, w7065, w7066, w7067, w7068, w7069, w7070, w7071, w7072, w7073, w7074, w7075, w7076, w7077, w7078, w7079, w7080, w7081, w7082, w7083, w7084, w7085, w7086, w7087, w7088, w7089, w7090, w7091, w7092, w7093, w7094, w7095, w7096, w7097, w7098, w7099, w7100, w7101, w7102, w7103, w7104, w7105, w7106, w7107, w7108, w7109, w7110, w7111, w7112, w7113, w7114, w7115, w7116, w7117, w7118, w7119, w7120, w7121, w7122, w7123, w7124, w7125, w7126, w7127, w7128, w7129, w7130, w7131, w7132, w7133, w7134, w7135, w7136, w7137, w7138, w7139, w7140, w7141, w7142, w7143, w7144, w7145, w7146, w7147, w7148, w7149, w7150, w7151, w7152, w7153, w7154, w7155, w7156, w7157, w7158, w7159, w7160, w7161, w7162, w7163, w7164, w7165, w7166, w7167, w7168, w7169, w7170, w7171, w7172, w7173, w7174, w7175, w7176, w7177, w7178, w7179, w7180, w7181, w7182, w7183, w7184, w7185, w7186, w7187, w7188, w7189, w7190, w7191, w7192, w7193, w7194, w7195, w7196, w7197, w7198, w7199, w7200, w7201, w7202, w7203, w7204, w7205, w7206, w7207, w7208, w7209, w7210, w7211, w7212, w7213, w7214, w7215, w7216, w7217, w7218, w7219, w7220, w7221, w7222, w7223, w7224, w7225, w7226, w7227, w7228, w7229, w7230, w7231, w7232, w7233, w7234, w7235, w7236, w7237, w7238, w7239, w7240, w7241, w7242, w7243, w7244, w7245, w7246, w7247, w7248, w7249, w7250, w7251, w7252, w7253, w7254, w7255, w7256, w7257, w7258, w7259, w7260, w7261, w7262, w7263, w7264, w7265, w7266, w7267, w7268, w7269, w7270, w7271, w7272, w7273, w7274, w7275, w7276, w7277, w7278, w7279, w7280, w7281, w7282, w7283, w7284, w7285, w7286, w7287, w7288, w7289, w7290, w7291, w7292, w7293, w7294, w7295, w7296, w7297, w7298, w7299, w7300, w7301, w7302, w7303, w7304, w7305, w7306, w7307, w7308, w7309, w7310, w7311, w7312, w7313, w7314, w7315, w7316, w7317, w7318, w7319, w7320, w7321, w7322, w7323, w7324, w7325, w7326, w7327, w7328, w7329, w7330, w7331, w7332, w7333, w7334, w7335, w7336, w7337, w7338, w7339, w7340, w7341, w7342, w7343, w7344, w7345, w7346, w7347, w7348, w7349, w7350, w7351, w7352, w7353, w7354, w7355, w7356, w7357, w7358, w7359, w7360, w7361, w7362, w7363, w7364, w7365, w7366, w7367, w7368, w7369, w7370, w7371, w7372, w7373, w7374, w7375, w7376, w7377, w7378, w7379, w7380, w7381, w7382, w7383, w7384, w7385, w7386, w7387, w7388, w7389, w7390, w7391, w7392, w7393, w7394, w7395, w7396, w7397, w7398, w7399, w7400, w7401, w7402, w7403, w7404, w7405, w7406, w7407, w7408, w7409, w7410, w7411, w7412, w7413, w7414, w7415, w7416, w7417, w7418, w7419, w7420, w7421, w7422, w7423, w7424, w7425, w7426, w7427, w7428, w7429, w7430, w7431, w7432, w7433, w7434, w7435, w7436, w7437, w7438, w7439, w7440, w7441, w7442, w7443, w7444, w7445, w7446, w7447, w7448, w7449, w7450, w7451, w7452, w7453, w7454, w7455, w7456, w7457, w7458, w7459, w7460, w7461, w7462, w7463, w7464, w7465, w7466, w7467, w7468, w7469, w7470, w7471, w7472, w7473, w7474, w7475, w7476, w7477, w7478, w7479, w7480, w7481, w7482, w7483, w7484, w7485, w7486, w7487, w7488, w7489, w7490, w7491, w7492, w7493, w7494, w7495, w7496, w7497, w7498, w7499, w7500, w7501, w7502, w7503, w7504, w7505, w7506, w7507, w7508, w7509, w7510, w7511, w7512, w7513, w7514, w7515, w7516, w7517, w7518, w7519, w7520, w7521, w7522, w7523, w7524, w7525, w7526, w7527, w7528, w7529, w7530, w7531, w7532, w7533, w7534, w7535, w7536, w7537, w7538, w7539, w7540, w7541, w7542, w7543, w7544, w7545, w7546, w7547, w7548, w7549, w7550, w7551, w7552, w7553, w7554, w7555, w7556, w7557, w7558, w7559, w7560, w7561, w7562, w7563, w7564, w7565, w7566, w7567, w7568, w7569, w7570, w7571, w7572, w7573, w7574, w7575, w7576, w7577, w7578, w7579, w7580, w7581, w7582, w7583, w7584, w7585, w7586, w7587, w7588, w7589, w7590, w7591, w7592, w7593, w7594, w7595, w7596, w7597, w7598, w7599, w7600, w7601, w7602, w7603, w7604, w7605, w7606, w7607, w7608, w7609, w7610, w7611, w7612, w7613, w7614, w7615, w7616, w7617, w7618, w7619, w7620, w7621, w7622, w7623, w7624, w7625, w7626, w7627, w7628, w7629, w7630, w7631, w7632, w7633, w7634, w7635, w7636, w7637, w7638, w7639, w7640, w7641, w7642, w7643, w7644, w7645, w7646, w7647, w7648, w7649, w7650, w7651, w7652, w7653, w7654, w7655, w7656, w7657, w7658, w7659, w7660, w7661, w7662, w7663, w7664, w7665, w7666, w7667, w7668, w7669, w7670, w7671, w7672, w7673, w7674, w7675, w7676, w7677, w7678, w7679, w7680, w7681, w7682, w7683, w7684, w7685, w7686, w7687, w7688, w7689, w7690, w7691, w7692, w7693, w7694, w7695, w7696, w7697, w7698, w7699, w7700, w7701, w7702, w7703, w7704, w7705, w7706, w7707, w7708, w7709, w7710, w7711, w7712, w7713, w7714, w7715, w7716, w7717, w7718, w7719, w7720, w7721, w7722, w7723, w7724, w7725, w7726, w7727, w7728, w7729, w7730, w7731, w7732, w7733, w7734, w7735, w7736, w7737, w7738, w7739, w7740, w7741, w7742, w7743, w7744, w7745, w7746, w7747, w7748, w7749, w7750, w7751, w7752, w7753, w7754, w7755, w7756, w7757, w7758, w7759, w7760, w7761, w7762, w7763, w7764, w7765, w7766, w7767, w7768, w7769, w7770, w7771, w7772, w7773, w7774, w7775, w7776, w7777, w7778, w7779, w7780, w7781, w7782, w7783, w7784, w7785, w7786, w7787, w7788, w7789, w7790, w7791, w7792, w7793, w7794, w7795, w7796, w7797, w7798, w7799, w7800, w7801, w7802, w7803, w7804, w7805, w7806, w7807, w7808, w7809, w7810, w7811, w7812, w7813, w7814, w7815, w7816, w7817, w7818, w7819, w7820, w7821, w7822, w7823, w7824, w7825, w7826, w7827, w7828, w7829, w7830, w7831, w7832, w7833, w7834, w7835, w7836, w7837, w7838, w7839, w7840, w7841, w7842, w7843, w7844, w7845, w7846, w7847, w7848, w7849, w7850, w7851, w7852, w7853, w7854, w7855, w7856, w7857, w7858, w7859, w7860, w7861, w7862, w7863, w7864, w7865, w7866, w7867, w7868, w7869, w7870, w7871, w7872, w7873, w7874, w7875, w7876, w7877, w7878, w7879, w7880, w7881, w7882, w7883, w7884, w7885, w7886, w7887, w7888, w7889, w7890, w7891, w7892, w7893, w7894, w7895, w7896, w7897, w7898, w7899, w7900, w7901, w7902, w7903, w7904, w7905, w7906, w7907, w7908, w7909, w7910, w7911, w7912, w7913, w7914, w7915, w7916, w7917, w7918, w7919, w7920, w7921, w7922, w7923, w7924, w7925, w7926, w7927, w7928, w7929, w7930, w7931, w7932, w7933, w7934, w7935, w7936, w7937, w7938, w7939, w7940, w7941, w7942, w7943, w7944, w7945, w7946, w7947, w7948, w7949, w7950, w7951, w7952, w7953, w7954, w7955, w7956, w7957, w7958, w7959, w7960, w7961, w7962, w7963, w7964, w7965, w7966, w7967, w7968, w7969, w7970, w7971, w7972, w7973, w7974, w7975, w7976, w7977, w7978, w7979, w7980, w7981, w7982, w7983, w7984, w7985, w7986, w7987, w7988, w7989, w7990, w7991, w7992, w7993, w7994, w7995, w7996, w7997, w7998, w7999, w8000, w8001, w8002, w8003, w8004, w8005, w8006, w8007, w8008, w8009, w8010, w8011, w8012, w8013, w8014, w8015, w8016, w8017, w8018, w8019, w8020, w8021, w8022, w8023, w8024, w8025, w8026, w8027, w8028, w8029, w8030, w8031, w8032, w8033, w8034, w8035, w8036, w8037, w8038, w8039, w8040, w8041, w8042, w8043, w8044, w8045, w8046, w8047, w8048, w8049, w8050, w8051, w8052, w8053, w8054, w8055, w8056, w8057, w8058, w8059, w8060, w8061, w8062, w8063, w8064, w8065, w8066, w8067, w8068, w8069, w8070, w8071, w8072, w8073, w8074, w8075, w8076, w8077, w8078, w8079, w8080, w8081, w8082, w8083, w8084, w8085, w8086, w8087, w8088, w8089, w8090, w8091, w8092, w8093, w8094, w8095, w8096, w8097, w8098, w8099, w8100, w8101, w8102, w8103, w8104, w8105, w8106, w8107, w8108, w8109, w8110, w8111, w8112, w8113, w8114, w8115, w8116, w8117, w8118, w8119, w8120, w8121, w8122, w8123, w8124, w8125, w8126, w8127, w8128, w8129, w8130, w8131, w8132, w8133, w8134, w8135, w8136, w8137, w8138, w8139, w8140, w8141, w8142, w8143, w8144, w8145, w8146, w8147, w8148, w8149, w8150, w8151, w8152, w8153, w8154, w8155, w8156, w8157, w8158, w8159, w8160, w8161, w8162, w8163, w8164, w8165, w8166, w8167, w8168, w8169, w8170, w8171, w8172, w8173, w8174, w8175, w8176, w8177, w8178, w8179, w8180, w8181, w8182, w8183, w8184, w8185, w8186, w8187, w8188, w8189, w8190, w8191, w8192, w8193, w8194, w8195, w8196, w8197, w8198, w8199, w8200, w8201, w8202, w8203, w8204, w8205, w8206, w8207, w8208, w8209, w8210, w8211, w8212, w8213, w8214, w8215, w8216, w8217, w8218, w8219, w8220, w8221, w8222, w8223, w8224, w8225, w8226, w8227, w8228, w8229, w8230, w8231, w8232, w8233, w8234, w8235, w8236, w8237, w8238, w8239, w8240, w8241, w8242, w8243, w8244, w8245, w8246, w8247, w8248, w8249, w8250, w8251, w8252, w8253, w8254, w8255, w8256, w8257, w8258, w8259, w8260, w8261, w8262, w8263, w8264, w8265, w8266, w8267, w8268, w8269, w8270, w8271, w8272, w8273, w8274, w8275, w8276, w8277, w8278, w8279, w8280, w8281, w8282, w8283, w8284, w8285, w8286, w8287, w8288, w8289, w8290, w8291, w8292, w8293, w8294, w8295, w8296, w8297, w8298, w8299, w8300, w8301, w8302, w8303, w8304, w8305, w8306, w8307, w8308, w8309, w8310, w8311, w8312, w8313, w8314, w8315, w8316, w8317, w8318, w8319, w8320, w8321, w8322, w8323, w8324, w8325, w8326, w8327, w8328, w8329, w8330, w8331, w8332, w8333, w8334, w8335, w8336, w8337, w8338, w8339, w8340, w8341, w8342, w8343, w8344, w8345, w8346, w8347, w8348, w8349, w8350, w8351, w8352, w8353, w8354, w8355, w8356, w8357, w8358, w8359, w8360, w8361, w8362, w8363, w8364, w8365, w8366, w8367, w8368, w8369, w8370, w8371, w8372, w8373, w8374, w8375, w8376, w8377, w8378, w8379, w8380, w8381, w8382, w8383, w8384, w8385, w8386, w8387, w8388, w8389, w8390, w8391, w8392, w8393, w8394, w8395, w8396, w8397, w8398, w8399, w8400, w8401, w8402, w8403, w8404, w8405, w8406, w8407, w8408, w8409, w8410, w8411, w8412, w8413, w8414, w8415, w8416, w8417, w8418, w8419, w8420, w8421, w8422, w8423, w8424, w8425, w8426, w8427, w8428, w8429, w8430, w8431, w8432, w8433, w8434, w8435, w8436, w8437, w8438, w8439, w8440, w8441, w8442, w8443, w8444, w8445, w8446, w8447, w8448, w8449, w8450, w8451, w8452, w8453, w8454, w8455, w8456, w8457, w8458, w8459, w8460, w8461, w8462, w8463, w8464, w8465, w8466, w8467, w8468, w8469, w8470, w8471, w8472, w8473, w8474, w8475, w8476, w8477, w8478, w8479, w8480, w8481, w8482, w8483, w8484, w8485, w8486, w8487, w8488, w8489, w8490, w8491, w8492, w8493, w8494, w8495, w8496, w8497, w8498, w8499, w8500, w8501, w8502, w8503, w8504, w8505, w8506, w8507, w8508, w8509, w8510, w8511, w8512, w8513, w8514, w8515, w8516, w8517, w8518, w8519, w8520, w8521, w8522, w8523, w8524, w8525, w8526, w8527, w8528, w8529, w8530, w8531, w8532, w8533, w8534, w8535, w8536, w8537, w8538, w8539, w8540, w8541, w8542, w8543, w8544, w8545, w8546, w8547, w8548, w8549, w8550, w8551, w8552, w8553, w8554, w8555, w8556, w8557, w8558, w8559, w8560, w8561, w8562, w8563, w8564, w8565, w8566, w8567, w8568, w8569, w8570, w8571, w8572, w8573, w8574, w8575, w8576, w8577, w8578, w8579, w8580, w8581, w8582, w8583, w8584, w8585, w8586, w8587, w8588, w8589, w8590, w8591, w8592, w8593, w8594, w8595, w8596, w8597, w8598, w8599, w8600, w8601, w8602, w8603, w8604, w8605, w8606, w8607, w8608, w8609, w8610, w8611, w8612, w8613, w8614, w8615, w8616, w8617, w8618, w8619, w8620, w8621, w8622, w8623, w8624, w8625, w8626, w8627, w8628, w8629, w8630, w8631, w8632, w8633, w8634, w8635, w8636, w8637, w8638, w8639, w8640, w8641, w8642, w8643, w8644, w8645, w8646, w8647, w8648, w8649, w8650, w8651, w8652, w8653, w8654, w8655, w8656, w8657, w8658, w8659, w8660, w8661, w8662, w8663, w8664, w8665, w8666, w8667, w8668, w8669, w8670, w8671, w8672, w8673, w8674, w8675, w8676, w8677, w8678, w8679, w8680, w8681, w8682, w8683, w8684, w8685, w8686, w8687, w8688, w8689, w8690, w8691, w8692, w8693, w8694, w8695, w8696, w8697, w8698, w8699, w8700, w8701, w8702, w8703, w8704, w8705, w8706, w8707, w8708, w8709, w8710, w8711, w8712, w8713, w8714, w8715, w8716, w8717, w8718, w8719, w8720, w8721, w8722, w8723, w8724, w8725, w8726, w8727, w8728, w8729, w8730, w8731, w8732, w8733, w8734, w8735, w8736, w8737, w8738, w8739, w8740, w8741, w8742, w8743, w8744, w8745, w8746, w8747, w8748, w8749, w8750, w8751, w8752, w8753, w8754, w8755, w8756, w8757, w8758, w8759, w8760, w8761, w8762, w8763, w8764, w8765, w8766, w8767, w8768, w8769, w8770, w8771, w8772, w8773, w8774, w8775, w8776, w8777, w8778, w8779, w8780, w8781, w8782, w8783, w8784, w8785, w8786, w8787, w8788, w8789, w8790, w8791, w8792, w8793, w8794, w8795, w8796, w8797, w8798, w8799, w8800, w8801, w8802, w8803, w8804, w8805, w8806, w8807, w8808, w8809, w8810, w8811, w8812, w8813, w8814, w8815, w8816, w8817, w8818, w8819, w8820, w8821, w8822, w8823, w8824, w8825, w8826, w8827, w8828, w8829, w8830, w8831, w8832, w8833, w8834, w8835, w8836, w8837, w8838, w8839, w8840, w8841, w8842, w8843, w8844, w8845, w8846, w8847, w8848, w8849, w8850, w8851, w8852, w8853, w8854, w8855, w8856, w8857, w8858, w8859, w8860, w8861, w8862, w8863, w8864, w8865, w8866, w8867, w8868, w8869, w8870, w8871, w8872, w8873, w8874, w8875, w8876, w8877, w8878, w8879, w8880, w8881, w8882, w8883, w8884, w8885, w8886, w8887, w8888, w8889, w8890, w8891, w8892, w8893, w8894, w8895, w8896, w8897, w8898, w8899, w8900, w8901, w8902, w8903, w8904, w8905, w8906, w8907, w8908, w8909, w8910, w8911, w8912, w8913, w8914, w8915, w8916, w8917, w8918, w8919, w8920, w8921, w8922, w8923, w8924, w8925, w8926, w8927, w8928, w8929, w8930, w8931, w8932, w8933, w8934, w8935, w8936, w8937, w8938, w8939, w8940, w8941, w8942, w8943, w8944, w8945, w8946, w8947, w8948, w8949, w8950, w8951, w8952, w8953, w8954, w8955, w8956, w8957, w8958, w8959, w8960, w8961, w8962, w8963, w8964, w8965, w8966, w8967, w8968, w8969, w8970, w8971, w8972, w8973, w8974, w8975, w8976, w8977, w8978, w8979, w8980, w8981, w8982, w8983, w8984, w8985, w8986, w8987, w8988, w8989, w8990, w8991, w8992, w8993, w8994, w8995, w8996, w8997, w8998, w8999, w9000, w9001, w9002, w9003, w9004, w9005, w9006, w9007, w9008, w9009, w9010, w9011, w9012, w9013, w9014, w9015, w9016, w9017, w9018, w9019, w9020, w9021, w9022, w9023, w9024, w9025, w9026, w9027, w9028, w9029, w9030, w9031, w9032, w9033, w9034, w9035, w9036, w9037, w9038, w9039, w9040, w9041, w9042, w9043, w9044, w9045, w9046, w9047, w9048, w9049, w9050, w9051, w9052, w9053, w9054, w9055, w9056, w9057, w9058, w9059, w9060, w9061, w9062, w9063, w9064, w9065, w9066, w9067, w9068, w9069, w9070, w9071, w9072, w9073, w9074, w9075, w9076, w9077, w9078, w9079, w9080, w9081, w9082, w9083, w9084, w9085, w9086, w9087, w9088, w9089, w9090, w9091, w9092, w9093, w9094, w9095, w9096, w9097, w9098, w9099, w9100, w9101, w9102, w9103, w9104, w9105, w9106, w9107, w9108, w9109, w9110, w9111, w9112, w9113, w9114, w9115, w9116, w9117, w9118, w9119, w9120, w9121, w9122, w9123, w9124, w9125, w9126, w9127, w9128, w9129, w9130, w9131, w9132, w9133, w9134, w9135, w9136, w9137, w9138, w9139, w9140, w9141, w9142, w9143, w9144, w9145, w9146, w9147, w9148, w9149, w9150, w9151, w9152, w9153, w9154, w9155, w9156, w9157, w9158, w9159, w9160, w9161, w9162, w9163, w9164, w9165, w9166, w9167, w9168, w9169, w9170, w9171, w9172, w9173, w9174, w9175, w9176, w9177, w9178, w9179, w9180, w9181, w9182, w9183, w9184, w9185, w9186, w9187, w9188, w9189, w9190, w9191, w9192, w9193, w9194, w9195, w9196, w9197, w9198, w9199, w9200, w9201, w9202, w9203, w9204, w9205, w9206, w9207, w9208, w9209, w9210, w9211, w9212, w9213, w9214, w9215, w9216, w9217, w9218, w9219, w9220, w9221, w9222, w9223, w9224, w9225, w9226, w9227, w9228, w9229, w9230, w9231, w9232, w9233, w9234, w9235, w9236, w9237, w9238, w9239, w9240, w9241, w9242, w9243, w9244, w9245, w9246, w9247, w9248, w9249, w9250, w9251, w9252, w9253, w9254, w9255, w9256, w9257, w9258, w9259, w9260, w9261, w9262, w9263, w9264, w9265, w9266, w9267, w9268, w9269, w9270, w9271, w9272, w9273, w9274, w9275, w9276, w9277, w9278, w9279, w9280, w9281, w9282, w9283, w9284, w9285, w9286, w9287, w9288, w9289, w9290, w9291, w9292, w9293, w9294, w9295, w9296, w9297, w9298, w9299, w9300, w9301, w9302, w9303, w9304, w9305, w9306, w9307, w9308, w9309, w9310, w9311, w9312, w9313, w9314, w9315, w9316, w9317, w9318, w9319, w9320, w9321, w9322, w9323, w9324, w9325, w9326, w9327, w9328, w9329, w9330, w9331, w9332, w9333, w9334, w9335, w9336, w9337, w9338, w9339, w9340, w9341, w9342, w9343, w9344, w9345, w9346, w9347, w9348, w9349, w9350, w9351, w9352, w9353, w9354, w9355, w9356, w9357, w9358, w9359, w9360, w9361, w9362, w9363, w9364, w9365, w9366, w9367, w9368, w9369, w9370, w9371, w9372, w9373, w9374, w9375, w9376, w9377, w9378, w9379, w9380, w9381, w9382, w9383, w9384, w9385, w9386, w9387, w9388, w9389, w9390, w9391, w9392, w9393, w9394, w9395, w9396, w9397, w9398, w9399, w9400, w9401, w9402, w9403, w9404, w9405, w9406, w9407, w9408, w9409, w9410, w9411, w9412, w9413, w9414, w9415, w9416, w9417, w9418, w9419, w9420, w9421, w9422, w9423, w9424, w9425, w9426, w9427, w9428, w9429, w9430, w9431, w9432, w9433, w9434, w9435, w9436, w9437, w9438, w9439, w9440, w9441, w9442, w9443, w9444, w9445, w9446, w9447, w9448, w9449, w9450, w9451, w9452, w9453, w9454, w9455, w9456, w9457, w9458, w9459, w9460, w9461, w9462, w9463, w9464, w9465, w9466, w9467, w9468, w9469, w9470, w9471, w9472, w9473, w9474, w9475, w9476, w9477, w9478, w9479, w9480, w9481, w9482, w9483, w9484, w9485, w9486, w9487, w9488, w9489, w9490, w9491, w9492, w9493, w9494, w9495, w9496, w9497, w9498, w9499, w9500, w9501, w9502, w9503, w9504, w9505, w9506, w9507, w9508, w9509, w9510, w9511, w9512, w9513, w9514, w9515, w9516, w9517, w9518, w9519, w9520, w9521, w9522, w9523, w9524, w9525, w9526, w9527, w9528, w9529, w9530, w9531, w9532, w9533, w9534, w9535, w9536, w9537, w9538, w9539, w9540, w9541, w9542, w9543, w9544, w9545, w9546, w9547, w9548, w9549, w9550, w9551, w9552, w9553, w9554, w9555, w9556, w9557, w9558, w9559, w9560, w9561, w9562, w9563, w9564, w9565, w9566, w9567, w9568, w9569, w9570, w9571, w9572, w9573, w9574, w9575, w9576, w9577, w9578, w9579, w9580, w9581, w9582, w9583, w9584, w9585, w9586, w9587, w9588, w9589, w9590, w9591, w9592, w9593, w9594, w9595, w9596, w9597, w9598, w9599, w9600, w9601, w9602, w9603, w9604, w9605, w9606, w9607, w9608, w9609, w9610, w9611, w9612, w9613, w9614, w9615, w9616, w9617, w9618, w9619, w9620, w9621, w9622, w9623, w9624, w9625, w9626, w9627, w9628, w9629, w9630, w9631, w9632, w9633, w9634, w9635, w9636, w9637, w9638, w9639, w9640, w9641, w9642, w9643, w9644, w9645, w9646, w9647, w9648, w9649, w9650, w9651, w9652, w9653, w9654, w9655, w9656, w9657, w9658, w9659, w9660, w9661, w9662, w9663, w9664, w9665, w9666, w9667, w9668, w9669, w9670, w9671, w9672, w9673, w9674, w9675, w9676, w9677, w9678, w9679, w9680, w9681, w9682, w9683, w9684, w9685, w9686, w9687, w9688, w9689, w9690, w9691, w9692, w9693, w9694, w9695, w9696, w9697, w9698, w9699, w9700, w9701, w9702, w9703, w9704, w9705, w9706, w9707, w9708, w9709, w9710, w9711, w9712, w9713, w9714, w9715, w9716, w9717, w9718, w9719, w9720, w9721, w9722, w9723, w9724, w9725, w9726, w9727, w9728, w9729, w9730, w9731, w9732, w9733, w9734, w9735, w9736, w9737, w9738, w9739, w9740, w9741, w9742, w9743, w9744, w9745, w9746, w9747, w9748, w9749, w9750, w9751, w9752, w9753, w9754, w9755, w9756, w9757, w9758, w9759, w9760, w9761, w9762, w9763, w9764, w9765, w9766, w9767, w9768, w9769, w9770, w9771, w9772, w9773, w9774, w9775, w9776, w9777, w9778, w9779, w9780, w9781, w9782, w9783, w9784, w9785, w9786, w9787, w9788, w9789, w9790, w9791, w9792, w9793, w9794, w9795, w9796, w9797, w9798, w9799, w9800, w9801, w9802, w9803, w9804, w9805, w9806, w9807, w9808, w9809, w9810, w9811, w9812, w9813, w9814, w9815, w9816, w9817, w9818, w9819, w9820, w9821, w9822, w9823, w9824, w9825, w9826, w9827, w9828, w9829, w9830, w9831, w9832, w9833, w9834, w9835, w9836, w9837, w9838, w9839, w9840, w9841, w9842, w9843, w9844, w9845, w9846, w9847, w9848, w9849, w9850, w9851, w9852, w9853, w9854, w9855, w9856, w9857, w9858, w9859, w9860, w9861, w9862, w9863, w9864, w9865, w9866, w9867, w9868, w9869, w9870, w9871, w9872, w9873, w9874, w9875, w9876, w9877, w9878, w9879, w9880, w9881, w9882, w9883, w9884, w9885, w9886, w9887, w9888, w9889, w9890, w9891, w9892, w9893, w9894, w9895, w9896, w9897, w9898, w9899, w9900, w9901, w9902, w9903, w9904, w9905, w9906, w9907, w9908, w9909, w9910, w9911, w9912, w9913, w9914, w9915, w9916, w9917, w9918, w9919, w9920, w9921, w9922, w9923, w9924, w9925, w9926, w9927, w9928, w9929, w9930, w9931, w9932, w9933, w9934, w9935, w9936, w9937, w9938, w9939, w9940, w9941, w9942, w9943, w9944, w9945, w9946, w9947, w9948, w9949, w9950, w9951, w9952, w9953, w9954, w9955, w9956, w9957, w9958, w9959, w9960, w9961, w9962, w9963, w9964, w9965, w9966, w9967, w9968, w9969, w9970, w9971, w9972, w9973, w9974, w9975, w9976, w9977, w9978, w9979, w9980, w9981, w9982, w9983, w9984, w9985, w9986, w9987, w9988, w9989, w9990, w9991, w9992, w9993, w9994, w9995, w9996, w9997, w9998, w9999, w10000, w10001, w10002, w10003, w10004, w10005, w10006, w10007, w10008, w10009, w10010, w10011, w10012, w10013, w10014, w10015, w10016, w10017, w10018, w10019, w10020, w10021, w10022, w10023, w10024, w10025, w10026, w10027, w10028, w10029, w10030, w10031, w10032, w10033, w10034, w10035, w10036, w10037, w10038, w10039, w10040, w10041, w10042, w10043, w10044, w10045, w10046, w10047, w10048, w10049, w10050, w10051, w10052, w10053, w10054, w10055, w10056, w10057, w10058, w10059, w10060, w10061, w10062, w10063, w10064, w10065, w10066, w10067, w10068, w10069, w10070, w10071, w10072, w10073, w10074, w10075, w10076, w10077, w10078, w10079, w10080, w10081, w10082, w10083, w10084, w10085, w10086, w10087, w10088, w10089, w10090, w10091, w10092, w10093, w10094, w10095, w10096, w10097, w10098, w10099, w10100, w10101, w10102, w10103, w10104, w10105, w10106, w10107, w10108, w10109, w10110, w10111, w10112, w10113, w10114, w10115, w10116, w10117, w10118, w10119, w10120, w10121, w10122, w10123, w10124, w10125, w10126, w10127, w10128, w10129, w10130, w10131, w10132, w10133, w10134, w10135, w10136, w10137, w10138, w10139, w10140, w10141, w10142, w10143, w10144, w10145, w10146, w10147, w10148, w10149, w10150, w10151, w10152, w10153, w10154, w10155, w10156, w10157, w10158, w10159, w10160, w10161, w10162, w10163, w10164, w10165, w10166, w10167, w10168, w10169, w10170, w10171, w10172, w10173, w10174, w10175, w10176, w10177, w10178, w10179, w10180, w10181, w10182, w10183, w10184, w10185, w10186, w10187, w10188, w10189, w10190, w10191, w10192, w10193, w10194, w10195, w10196, w10197, w10198, w10199, w10200, w10201, w10202, w10203, w10204, w10205, w10206, w10207, w10208, w10209, w10210, w10211, w10212, w10213, w10214, w10215, w10216, w10217, w10218, w10219, w10220, w10221, w10222, w10223, w10224, w10225, w10226, w10227, w10228, w10229, w10230, w10231, w10232, w10233, w10234, w10235, w10236, w10237, w10238, w10239, w10240, w10241, w10242, w10243, w10244, w10245, w10246, w10247, w10248, w10249, w10250, w10251, w10252, w10253, w10254, w10255, w10256, w10257, w10258, w10259, w10260, w10261, w10262, w10263, w10264, w10265, w10266, w10267, w10268, w10269, w10270, w10271, w10272, w10273, w10274, w10275, w10276, w10277, w10278, w10279, w10280, w10281, w10282, w10283, w10284, w10285, w10286, w10287, w10288, w10289, w10290, w10291, w10292, w10293, w10294, w10295, w10296, w10297, w10298, w10299, w10300, w10301, w10302, w10303, w10304, w10305, w10306, w10307, w10308, w10309, w10310, w10311, w10312, w10313, w10314, w10315, w10316, w10317, w10318, w10319, w10320, w10321, w10322, w10323, w10324, w10325, w10326, w10327, w10328, w10329, w10330, w10331, w10332, w10333, w10334, w10335, w10336, w10337, w10338, w10339, w10340, w10341, w10342, w10343, w10344, w10345, w10346, w10347, w10348, w10349, w10350, w10351, w10352, w10353, w10354, w10355, w10356, w10357, w10358, w10359, w10360, w10361, w10362, w10363, w10364, w10365, w10366, w10367, w10368, w10369, w10370, w10371, w10372, w10373, w10374, w10375, w10376, w10377, w10378, w10379, w10380, w10381, w10382, w10383, w10384, w10385, w10386, w10387, w10388, w10389, w10390, w10391, w10392, w10393, w10394, w10395, w10396, w10397, w10398, w10399, w10400, w10401, w10402, w10403, w10404, w10405, w10406, w10407, w10408, w10409, w10410, w10411, w10412, w10413, w10414, w10415, w10416, w10417, w10418, w10419, w10420, w10421, w10422, w10423, w10424, w10425, w10426, w10427, w10428, w10429, w10430, w10431, w10432, w10433, w10434, w10435, w10436, w10437, w10438, w10439, w10440, w10441, w10442, w10443, w10444, w10445, w10446, w10447, w10448, w10449, w10450, w10451, w10452, w10453, w10454, w10455, w10456, w10457, w10458, w10459, w10460, w10461, w10462, w10463, w10464, w10465, w10466, w10467, w10468, w10469, w10470, w10471, w10472, w10473, w10474, w10475, w10476, w10477, w10478, w10479, w10480, w10481, w10482, w10483, w10484, w10485, w10486, w10487, w10488, w10489, w10490, w10491, w10492, w10493, w10494, w10495, w10496, w10497, w10498, w10499, w10500, w10501, w10502, w10503, w10504, w10505, w10506, w10507, w10508, w10509, w10510, w10511, w10512, w10513, w10514, w10515, w10516, w10517, w10518, w10519, w10520, w10521, w10522, w10523, w10524, w10525, w10526, w10527, w10528, w10529, w10530, w10531, w10532, w10533, w10534, w10535, w10536, w10537, w10538, w10539, w10540, w10541, w10542, w10543, w10544, w10545, w10546, w10547, w10548, w10549, w10550, w10551, w10552, w10553, w10554, w10555, w10556, w10557, w10558, w10559, w10560, w10561, w10562, w10563, w10564, w10565, w10566, w10567, w10568, w10569, w10570, w10571, w10572, w10573, w10574, w10575, w10576, w10577, w10578, w10579, w10580, w10581, w10582, w10583, w10584, w10585, w10586, w10587, w10588, w10589, w10590, w10591, w10592, w10593, w10594, w10595, w10596, w10597, w10598, w10599, w10600, w10601, w10602, w10603, w10604, w10605, w10606, w10607, w10608, w10609, w10610, w10611, w10612, w10613, w10614, w10615, w10616, w10617, w10618, w10619, w10620, w10621, w10622, w10623, w10624, w10625, w10626, w10627, w10628, w10629, w10630, w10631, w10632, w10633, w10634, w10635, w10636, w10637, w10638, w10639, w10640, w10641, w10642, w10643, w10644, w10645, w10646, w10647, w10648, w10649, w10650, w10651, w10652, w10653, w10654, w10655, w10656, w10657, w10658, w10659, w10660, w10661, w10662, w10663, w10664, w10665, w10666, w10667, w10668, w10669, w10670, w10671, w10672, w10673, w10674, w10675, w10676, w10677, w10678, w10679, w10680, w10681, w10682, w10683, w10684, w10685, w10686, w10687, w10688, w10689, w10690, w10691, w10692, w10693, w10694, w10695, w10696, w10697, w10698, w10699, w10700, w10701, w10702, w10703, w10704, w10705, w10706, w10707, w10708, w10709, w10710, w10711, w10712, w10713, w10714, w10715, w10716, w10717, w10718, w10719, w10720, w10721, w10722, w10723, w10724, w10725, w10726, w10727, w10728, w10729, w10730, w10731, w10732, w10733, w10734, w10735, w10736, w10737, w10738, w10739, w10740, w10741, w10742, w10743, w10744, w10745, w10746, w10747, w10748, w10749, w10750, w10751, w10752, w10753, w10754, w10755, w10756, w10757, w10758, w10759, w10760, w10761, w10762, w10763, w10764, w10765, w10766, w10767, w10768, w10769, w10770, w10771, w10772, w10773, w10774, w10775, w10776, w10777, w10778, w10779, w10780, w10781, w10782, w10783, w10784, w10785, w10786, w10787, w10788, w10789, w10790, w10791, w10792, w10793, w10794, w10795, w10796, w10797, w10798, w10799, w10800, w10801, w10802, w10803, w10804, w10805, w10806, w10807, w10808, w10809, w10810, w10811, w10812, w10813, w10814, w10815, w10816, w10817, w10818, w10819, w10820, w10821, w10822, w10823, w10824, w10825, w10826, w10827, w10828, w10829, w10830, w10831, w10832, w10833, w10834, w10835, w10836, w10837, w10838, w10839, w10840, w10841, w10842, w10843, w10844, w10845, w10846, w10847, w10848, w10849, w10850, w10851, w10852, w10853, w10854, w10855, w10856, w10857, w10858, w10859, w10860, w10861, w10862, w10863, w10864, w10865, w10866, w10867, w10868, w10869, w10870, w10871, w10872, w10873, w10874, w10875, w10876, w10877, w10878, w10879, w10880, w10881, w10882, w10883, w10884, w10885, w10886, w10887, w10888, w10889, w10890, w10891, w10892, w10893, w10894, w10895, w10896, w10897, w10898, w10899, w10900, w10901, w10902, w10903, w10904, w10905, w10906, w10907, w10908, w10909, w10910, w10911, w10912, w10913, w10914, w10915, w10916, w10917, w10918, w10919, w10920, w10921, w10922, w10923, w10924, w10925, w10926, w10927, w10928, w10929, w10930, w10931, w10932, w10933, w10934, w10935, w10936, w10937, w10938, w10939, w10940, w10941, w10942, w10943, w10944, w10945, w10946, w10947, w10948, w10949, w10950, w10951, w10952, w10953, w10954, w10955, w10956, w10957, w10958, w10959, w10960, w10961, w10962, w10963, w10964, w10965, w10966, w10967, w10968, w10969, w10970, w10971, w10972, w10973, w10974, w10975, w10976, w10977, w10978, w10979, w10980, w10981, w10982, w10983, w10984, w10985, w10986, w10987, w10988, w10989, w10990, w10991, w10992, w10993, w10994, w10995, w10996, w10997, w10998, w10999, w11000, w11001, w11002, w11003, w11004, w11005, w11006, w11007, w11008, w11009, w11010, w11011, w11012, w11013, w11014, w11015, w11016, w11017, w11018, w11019, w11020, w11021, w11022, w11023, w11024, w11025, w11026, w11027, w11028, w11029, w11030, w11031, w11032, w11033, w11034, w11035, w11036, w11037, w11038, w11039, w11040, w11041, w11042, w11043, w11044, w11045, w11046, w11047, w11048, w11049, w11050, w11051, w11052, w11053, w11054, w11055, w11056, w11057, w11058, w11059, w11060, w11061, w11062, w11063, w11064, w11065, w11066, w11067, w11068, w11069, w11070, w11071, w11072, w11073, w11074, w11075, w11076, w11077, w11078, w11079, w11080, w11081, w11082, w11083, w11084, w11085, w11086, w11087, w11088, w11089, w11090, w11091, w11092, w11093, w11094, w11095, w11096, w11097, w11098, w11099, w11100, w11101, w11102, w11103, w11104, w11105, w11106, w11107, w11108, w11109, w11110, w11111, w11112, w11113, w11114, w11115, w11116, w11117, w11118, w11119, w11120, w11121, w11122, w11123, w11124, w11125, w11126, w11127, w11128, w11129, w11130, w11131, w11132, w11133, w11134, w11135, w11136, w11137, w11138, w11139, w11140, w11141, w11142, w11143, w11144, w11145, w11146, w11147, w11148, w11149, w11150, w11151, w11152, w11153, w11154, w11155, w11156, w11157, w11158, w11159, w11160, w11161, w11162, w11163, w11164, w11165, w11166, w11167, w11168, w11169, w11170, w11171, w11172, w11173, w11174, w11175, w11176, w11177, w11178, w11179, w11180, w11181, w11182, w11183, w11184, w11185, w11186, w11187, w11188, w11189, w11190, w11191, w11192, w11193, w11194, w11195, w11196, w11197, w11198, w11199, w11200, w11201, w11202, w11203, w11204, w11205, w11206, w11207, w11208, w11209, w11210, w11211, w11212, w11213, w11214, w11215, w11216, w11217, w11218, w11219, w11220, w11221, w11222, w11223, w11224, w11225, w11226, w11227, w11228, w11229, w11230, w11231, w11232, w11233, w11234, w11235, w11236, w11237, w11238, w11239, w11240, w11241, w11242, w11243, w11244, w11245, w11246, w11247, w11248, w11249, w11250, w11251, w11252, w11253, w11254, w11255, w11256, w11257, w11258, w11259, w11260, w11261, w11262, w11263, w11264, w11265, w11266, w11267, w11268, w11269, w11270, w11271, w11272, w11273, w11274, w11275, w11276, w11277, w11278, w11279, w11280, w11281, w11282, w11283, w11284, w11285, w11286, w11287, w11288, w11289, w11290, w11291, w11292, w11293, w11294, w11295, w11296, w11297, w11298, w11299, w11300, w11301, w11302, w11303, w11304, w11305, w11306, w11307, w11308, w11309, w11310, w11311, w11312, w11313, w11314, w11315, w11316, w11317, w11318, w11319, w11320, w11321, w11322, w11323, w11324, w11325, w11326, w11327, w11328, w11329, w11330, w11331, w11332, w11333, w11334, w11335, w11336, w11337, w11338, w11339, w11340, w11341, w11342, w11343, w11344, w11345, w11346, w11347, w11348, w11349, w11350, w11351, w11352, w11353, w11354, w11355, w11356, w11357, w11358, w11359, w11360, w11361, w11362, w11363, w11364, w11365, w11366, w11367, w11368, w11369, w11370, w11371, w11372, w11373, w11374, w11375, w11376, w11377, w11378, w11379, w11380, w11381, w11382, w11383, w11384, w11385, w11386, w11387, w11388, w11389, w11390, w11391, w11392, w11393, w11394, w11395, w11396, w11397, w11398, w11399, w11400, w11401, w11402, w11403, w11404, w11405, w11406, w11407, w11408, w11409, w11410, w11411, w11412, w11413, w11414, w11415, w11416, w11417, w11418, w11419, w11420, w11421, w11422, w11423, w11424, w11425, w11426, w11427, w11428, w11429, w11430, w11431, w11432, w11433, w11434, w11435, w11436, w11437, w11438, w11439, w11440, w11441, w11442, w11443, w11444, w11445, w11446, w11447, w11448, w11449, w11450, w11451, w11452, w11453, w11454, w11455, w11456, w11457, w11458, w11459, w11460, w11461, w11462, w11463, w11464, w11465, w11466, w11467, w11468, w11469, w11470, w11471, w11472, w11473, w11474, w11475, w11476, w11477, w11478, w11479, w11480, w11481, w11482, w11483, w11484, w11485, w11486, w11487, w11488, w11489, w11490, w11491, w11492, w11493, w11494, w11495, w11496, w11497, w11498, w11499, w11500, w11501, w11502, w11503, w11504, w11505, w11506, w11507, w11508, w11509, w11510, w11511, w11512, w11513, w11514, w11515, w11516, w11517, w11518, w11519, w11520, w11521, w11522, w11523, w11524, w11525, w11526, w11527, w11528, w11529, w11530, w11531, w11532, w11533, w11534, w11535, w11536, w11537, w11538, w11539, w11540, w11541, w11542, w11543, w11544, w11545, w11546, w11547, w11548, w11549, w11550, w11551, w11552, w11553, w11554, w11555, w11556, w11557, w11558, w11559, w11560, w11561, w11562, w11563, w11564, w11565, w11566, w11567, w11568, w11569, w11570, w11571, w11572, w11573, w11574, w11575, w11576, w11577, w11578, w11579, w11580, w11581, w11582, w11583, w11584, w11585, w11586, w11587, w11588, w11589, w11590, w11591, w11592, w11593, w11594, w11595, w11596, w11597, w11598, w11599, w11600, w11601, w11602, w11603, w11604, w11605, w11606, w11607, w11608, w11609, w11610, w11611, w11612, w11613, w11614, w11615, w11616, w11617, w11618, w11619, w11620, w11621, w11622, w11623, w11624, w11625, w11626, w11627, w11628, w11629, w11630, w11631, w11632, w11633, w11634, w11635, w11636, w11637, w11638, w11639, w11640, w11641, w11642, w11643, w11644, w11645, w11646, w11647, w11648, w11649, w11650, w11651, w11652, w11653, w11654, w11655, w11656, w11657, w11658, w11659, w11660, w11661, w11662, w11663, w11664, w11665, w11666, w11667, w11668, w11669, w11670, w11671, w11672, w11673, w11674, w11675, w11676, w11677, w11678, w11679, w11680, w11681, w11682, w11683, w11684, w11685, w11686, w11687, w11688, w11689, w11690, w11691, w11692, w11693, w11694, w11695, w11696, w11697, w11698, w11699, w11700, w11701, w11702, w11703, w11704, w11705, w11706, w11707, w11708, w11709, w11710, w11711, w11712, w11713, w11714, w11715, w11716, w11717, w11718, w11719, w11720, w11721, w11722, w11723, w11724, w11725, w11726, w11727, w11728, w11729, w11730, w11731, w11732, w11733, w11734, w11735, w11736, w11737, w11738, w11739, w11740, w11741, w11742, w11743, w11744, w11745, w11746, w11747, w11748, w11749, w11750, w11751, w11752, w11753, w11754, w11755, w11756, w11757, w11758, w11759, w11760, w11761, w11762, w11763, w11764, w11765, w11766, w11767, w11768, w11769, w11770, w11771, w11772, w11773, w11774, w11775, w11776, w11777, w11778, w11779, w11780, w11781, w11782, w11783, w11784, w11785, w11786, w11787, w11788, w11789, w11790, w11791, w11792, w11793, w11794, w11795, w11796, w11797, w11798, w11799, w11800, w11801, w11802, w11803, w11804, w11805, w11806, w11807, w11808, w11809, w11810, w11811, w11812, w11813, w11814, w11815, w11816, w11817, w11818, w11819, w11820, w11821, w11822, w11823, w11824, w11825, w11826, w11827, w11828, w11829, w11830, w11831, w11832, w11833, w11834, w11835, w11836, w11837, w11838, w11839, w11840, w11841, w11842, w11843, w11844, w11845, w11846, w11847, w11848, w11849, w11850, w11851, w11852, w11853, w11854, w11855, w11856, w11857, w11858, w11859, w11860, w11861, w11862, w11863, w11864, w11865, w11866, w11867, w11868, w11869, w11870, w11871, w11872, w11873, w11874, w11875, w11876, w11877, w11878, w11879, w11880, w11881, w11882, w11883, w11884, w11885, w11886, w11887, w11888, w11889, w11890, w11891, w11892, w11893, w11894, w11895, w11896, w11897, w11898, w11899, w11900, w11901, w11902, w11903, w11904, w11905, w11906, w11907, w11908, w11909, w11910, w11911, w11912, w11913, w11914, w11915, w11916, w11917, w11918, w11919, w11920, w11921, w11922, w11923, w11924, w11925, w11926, w11927, w11928, w11929, w11930, w11931, w11932, w11933, w11934, w11935, w11936, w11937, w11938, w11939, w11940, w11941, w11942, w11943, w11944, w11945, w11946, w11947, w11948, w11949, w11950, w11951, w11952, w11953, w11954, w11955, w11956, w11957, w11958, w11959, w11960, w11961, w11962, w11963, w11964, w11965, w11966, w11967, w11968, w11969, w11970, w11971, w11972, w11973, w11974, w11975, w11976, w11977, w11978, w11979, w11980, w11981, w11982, w11983, w11984, w11985, w11986, w11987, w11988, w11989, w11990, w11991, w11992, w11993, w11994, w11995, w11996, w11997, w11998, w11999, w12000, w12001, w12002, w12003, w12004, w12005, w12006, w12007, w12008, w12009, w12010, w12011, w12012, w12013, w12014, w12015, w12016, w12017, w12018, w12019, w12020, w12021, w12022, w12023, w12024, w12025, w12026, w12027, w12028, w12029, w12030, w12031, w12032, w12033, w12034, w12035, w12036, w12037, w12038, w12039, w12040, w12041, w12042, w12043, w12044, w12045, w12046, w12047, w12048, w12049, w12050, w12051, w12052, w12053, w12054, w12055, w12056, w12057, w12058, w12059, w12060, w12061, w12062, w12063, w12064, w12065, w12066, w12067, w12068, w12069, w12070, w12071, w12072, w12073, w12074, w12075, w12076, w12077, w12078, w12079, w12080, w12081, w12082, w12083, w12084, w12085, w12086, w12087, w12088, w12089, w12090, w12091, w12092, w12093, w12094, w12095, w12096, w12097, w12098, w12099, w12100, w12101, w12102, w12103, w12104, w12105, w12106, w12107, w12108, w12109, w12110, w12111, w12112, w12113, w12114, w12115, w12116, w12117, w12118, w12119, w12120, w12121, w12122, w12123, w12124, w12125, w12126, w12127, w12128, w12129, w12130, w12131, w12132, w12133, w12134, w12135, w12136, w12137, w12138, w12139, w12140, w12141, w12142, w12143, w12144, w12145, w12146, w12147, w12148, w12149, w12150, w12151, w12152, w12153, w12154, w12155, w12156, w12157, w12158, w12159, w12160, w12161, w12162, w12163, w12164, w12165, w12166, w12167, w12168, w12169, w12170, w12171, w12172, w12173, w12174, w12175, w12176, w12177, w12178, w12179, w12180, w12181, w12182, w12183, w12184, w12185, w12186, w12187, w12188, w12189, w12190, w12191, w12192, w12193, w12194, w12195, w12196, w12197, w12198, w12199, w12200, w12201, w12202, w12203, w12204, w12205, w12206, w12207, w12208, w12209, w12210, w12211, w12212, w12213, w12214, w12215, w12216, w12217, w12218, w12219, w12220, w12221, w12222, w12223, w12224, w12225, w12226, w12227, w12228, w12229, w12230, w12231, w12232, w12233, w12234, w12235, w12236, w12237, w12238, w12239, w12240, w12241, w12242, w12243, w12244, w12245, w12246, w12247, w12248, w12249, w12250, w12251, w12252, w12253, w12254, w12255, w12256, w12257, w12258, w12259, w12260, w12261, w12262, w12263, w12264, w12265, w12266, w12267, w12268, w12269, w12270, w12271, w12272, w12273, w12274, w12275, w12276, w12277, w12278, w12279, w12280, w12281, w12282, w12283, w12284, w12285, w12286, w12287, w12288, w12289, w12290, w12291, w12292, w12293, w12294, w12295, w12296, w12297, w12298, w12299, w12300, w12301, w12302, w12303, w12304, w12305, w12306, w12307, w12308, w12309, w12310, w12311, w12312, w12313, w12314, w12315, w12316, w12317, w12318, w12319, w12320, w12321, w12322, w12323, w12324, w12325, w12326, w12327, w12328, w12329, w12330, w12331, w12332, w12333, w12334, w12335, w12336, w12337, w12338, w12339, w12340, w12341, w12342, w12343, w12344, w12345, w12346, w12347, w12348, w12349, w12350, w12351, w12352, w12353, w12354, w12355, w12356, w12357, w12358, w12359, w12360, w12361, w12362, w12363, w12364, w12365, w12366, w12367, w12368, w12369, w12370, w12371, w12372, w12373, w12374, w12375, w12376, w12377, w12378, w12379, w12380, w12381, w12382, w12383, w12384, w12385, w12386, w12387, w12388, w12389, w12390, w12391, w12392, w12393, w12394, w12395, w12396, w12397, w12398, w12399, w12400, w12401, w12402, w12403, w12404, w12405, w12406, w12407, w12408, w12409, w12410, w12411, w12412, w12413, w12414, w12415, w12416, w12417, w12418, w12419, w12420, w12421, w12422, w12423, w12424, w12425, w12426, w12427, w12428, w12429, w12430, w12431, w12432, w12433, w12434, w12435, w12436, w12437, w12438, w12439, w12440, w12441, w12442, w12443, w12444, w12445, w12446, w12447, w12448, w12449, w12450, w12451, w12452, w12453, w12454, w12455, w12456, w12457, w12458, w12459, w12460, w12461, w12462, w12463, w12464, w12465, w12466, w12467, w12468, w12469, w12470, w12471, w12472, w12473, w12474, w12475, w12476, w12477, w12478, w12479, w12480, w12481, w12482, w12483, w12484, w12485, w12486, w12487, w12488, w12489, w12490, w12491, w12492, w12493, w12494, w12495, w12496, w12497, w12498, w12499, w12500, w12501, w12502, w12503, w12504, w12505, w12506, w12507, w12508, w12509, w12510, w12511, w12512, w12513, w12514, w12515, w12516, w12517, w12518, w12519, w12520, w12521, w12522, w12523, w12524, w12525, w12526, w12527, w12528, w12529, w12530, w12531, w12532, w12533, w12534, w12535, w12536, w12537, w12538, w12539, w12540, w12541, w12542, w12543, w12544, w12545, w12546, w12547, w12548, w12549, w12550, w12551, w12552, w12553, w12554, w12555, w12556, w12557, w12558, w12559, w12560, w12561, w12562, w12563, w12564, w12565, w12566, w12567, w12568, w12569, w12570, w12571, w12572, w12573, w12574, w12575, w12576, w12577, w12578, w12579, w12580, w12581, w12582, w12583, w12584, w12585, w12586, w12587, w12588, w12589, w12590, w12591, w12592, w12593, w12594, w12595, w12596, w12597, w12598, w12599, w12600, w12601, w12602, w12603, w12604, w12605, w12606, w12607, w12608, w12609, w12610, w12611, w12612, w12613, w12614, w12615, w12616, w12617, w12618, w12619, w12620, w12621, w12622, w12623, w12624, w12625, w12626, w12627, w12628, w12629, w12630, w12631, w12632, w12633, w12634, w12635, w12636, w12637, w12638, w12639, w12640, w12641, w12642, w12643, w12644, w12645, w12646, w12647, w12648, w12649, w12650, w12651, w12652, w12653, w12654, w12655, w12656, w12657, w12658, w12659, w12660, w12661, w12662, w12663, w12664, w12665, w12666, w12667, w12668, w12669, w12670, w12671, w12672, w12673, w12674, w12675, w12676, w12677, w12678, w12679, w12680, w12681, w12682, w12683, w12684, w12685, w12686, w12687, w12688, w12689, w12690, w12691, w12692, w12693, w12694, w12695, w12696, w12697, w12698, w12699, w12700, w12701, w12702, w12703, w12704, w12705, w12706, w12707, w12708, w12709, w12710, w12711, w12712, w12713, w12714, w12715, w12716, w12717, w12718, w12719, w12720, w12721, w12722, w12723, w12724, w12725, w12726, w12727, w12728, w12729, w12730, w12731, w12732, w12733, w12734, w12735, w12736, w12737, w12738, w12739, w12740, w12741, w12742, w12743, w12744, w12745, w12746, w12747, w12748, w12749, w12750, w12751, w12752, w12753, w12754, w12755, w12756, w12757, w12758, w12759, w12760, w12761, w12762, w12763, w12764, w12765, w12766, w12767, w12768, w12769, w12770, w12771, w12772, w12773, w12774, w12775, w12776, w12777, w12778, w12779, w12780, w12781, w12782, w12783, w12784, w12785, w12786, w12787, w12788, w12789, w12790, w12791, w12792, w12793, w12794, w12795, w12796, w12797, w12798, w12799, w12800, w12801, w12802, w12803, w12804, w12805, w12806, w12807, w12808, w12809, w12810, w12811, w12812, w12813, w12814, w12815, w12816, w12817, w12818, w12819, w12820, w12821, w12822, w12823, w12824, w12825, w12826, w12827, w12828, w12829, w12830, w12831, w12832, w12833, w12834, w12835, w12836, w12837, w12838, w12839, w12840, w12841, w12842, w12843, w12844, w12845, w12846, w12847, w12848, w12849, w12850, w12851, w12852, w12853, w12854, w12855, w12856, w12857, w12858, w12859, w12860, w12861, w12862, w12863, w12864, w12865, w12866, w12867, w12868, w12869, w12870, w12871, w12872, w12873, w12874, w12875, w12876, w12877, w12878, w12879, w12880, w12881, w12882, w12883, w12884, w12885, w12886, w12887, w12888, w12889, w12890, w12891, w12892, w12893, w12894, w12895, w12896, w12897, w12898, w12899, w12900, w12901, w12902, w12903, w12904, w12905, w12906, w12907, w12908, w12909, w12910, w12911, w12912, w12913, w12914, w12915, w12916, w12917, w12918, w12919, w12920, w12921, w12922, w12923, w12924, w12925, w12926, w12927, w12928, w12929, w12930, w12931, w12932, w12933, w12934, w12935, w12936, w12937, w12938, w12939, w12940, w12941, w12942, w12943, w12944, w12945, w12946, w12947, w12948, w12949, w12950, w12951, w12952, w12953, w12954, w12955, w12956, w12957, w12958, w12959, w12960, w12961, w12962, w12963, w12964, w12965, w12966, w12967, w12968, w12969, w12970, w12971, w12972, w12973, w12974, w12975, w12976, w12977, w12978, w12979, w12980, w12981, w12982, w12983, w12984, w12985, w12986, w12987, w12988, w12989, w12990, w12991, w12992, w12993, w12994, w12995, w12996, w12997, w12998, w12999, w13000, w13001, w13002, w13003, w13004, w13005, w13006, w13007, w13008, w13009, w13010, w13011, w13012, w13013, w13014, w13015, w13016, w13017, w13018, w13019, w13020, w13021, w13022, w13023, w13024, w13025, w13026, w13027, w13028, w13029, w13030, w13031, w13032, w13033, w13034, w13035, w13036, w13037, w13038, w13039, w13040, w13041, w13042, w13043, w13044, w13045, w13046, w13047, w13048, w13049, w13050, w13051, w13052, w13053, w13054, w13055, w13056, w13057, w13058, w13059, w13060, w13061, w13062, w13063, w13064, w13065, w13066, w13067, w13068, w13069, w13070, w13071, w13072, w13073, w13074, w13075, w13076, w13077, w13078, w13079, w13080, w13081, w13082, w13083, w13084, w13085, w13086, w13087, w13088, w13089, w13090, w13091, w13092, w13093, w13094, w13095, w13096, w13097, w13098, w13099, w13100, w13101, w13102, w13103, w13104, w13105, w13106, w13107, w13108, w13109, w13110, w13111, w13112, w13113, w13114, w13115, w13116, w13117, w13118, w13119, w13120, w13121, w13122, w13123, w13124, w13125, w13126, w13127, w13128, w13129, w13130, w13131, w13132, w13133, w13134, w13135, w13136, w13137, w13138, w13139, w13140, w13141, w13142, w13143, w13144, w13145, w13146, w13147, w13148, w13149, w13150, w13151, w13152, w13153, w13154, w13155, w13156, w13157, w13158, w13159, w13160, w13161, w13162, w13163, w13164, w13165, w13166, w13167, w13168, w13169, w13170, w13171, w13172, w13173, w13174, w13175, w13176, w13177, w13178, w13179, w13180, w13181, w13182, w13183, w13184, w13185, w13186, w13187, w13188, w13189, w13190, w13191, w13192, w13193, w13194, w13195, w13196, w13197, w13198, w13199, w13200, w13201, w13202, w13203, w13204, w13205, w13206, w13207, w13208, w13209, w13210, w13211, w13212, w13213, w13214, w13215, w13216, w13217, w13218, w13219, w13220, w13221, w13222, w13223, w13224, w13225, w13226, w13227, w13228, w13229, w13230, w13231, w13232, w13233, w13234, w13235, w13236, w13237, w13238, w13239, w13240, w13241, w13242, w13243, w13244, w13245, w13246, w13247, w13248, w13249, w13250, w13251, w13252, w13253, w13254, w13255, w13256, w13257, w13258, w13259, w13260, w13261, w13262, w13263, w13264, w13265, w13266, w13267, w13268, w13269, w13270, w13271, w13272, w13273, w13274, w13275, w13276, w13277, w13278, w13279, w13280, w13281, w13282, w13283, w13284, w13285, w13286, w13287, w13288, w13289, w13290, w13291, w13292, w13293, w13294, w13295, w13296, w13297, w13298, w13299, w13300, w13301, w13302, w13303, w13304, w13305, w13306, w13307, w13308, w13309, w13310, w13311, w13312, w13313, w13314, w13315, w13316, w13317, w13318, w13319, w13320, w13321, w13322, w13323, w13324, w13325, w13326, w13327, w13328, w13329, w13330, w13331, w13332, w13333, w13334, w13335, w13336, w13337, w13338, w13339, w13340, w13341, w13342, w13343, w13344, w13345, w13346, w13347, w13348, w13349, w13350, w13351, w13352, w13353, w13354, w13355, w13356, w13357, w13358, w13359, w13360, w13361, w13362, w13363, w13364, w13365, w13366, w13367, w13368, w13369, w13370, w13371, w13372, w13373, w13374, w13375, w13376, w13377, w13378, w13379, w13380, w13381, w13382, w13383, w13384, w13385, w13386, w13387, w13388, w13389, w13390, w13391, w13392, w13393, w13394, w13395, w13396, w13397, w13398, w13399, w13400, w13401, w13402, w13403, w13404, w13405, w13406, w13407, w13408, w13409, w13410, w13411, w13412, w13413, w13414, w13415, w13416, w13417, w13418, w13419, w13420, w13421, w13422, w13423, w13424, w13425, w13426, w13427, w13428, w13429, w13430, w13431, w13432, w13433, w13434, w13435, w13436, w13437, w13438, w13439, w13440, w13441, w13442, w13443, w13444, w13445, w13446, w13447, w13448, w13449, w13450, w13451, w13452, w13453, w13454, w13455, w13456, w13457, w13458, w13459, w13460, w13461, w13462, w13463, w13464, w13465, w13466, w13467, w13468, w13469, w13470, w13471, w13472, w13473, w13474, w13475, w13476, w13477, w13478, w13479, w13480, w13481, w13482, w13483, w13484, w13485, w13486, w13487, w13488, w13489, w13490, w13491, w13492, w13493, w13494, w13495, w13496, w13497, w13498, w13499, w13500, w13501, w13502, w13503, w13504, w13505, w13506, w13507, w13508, w13509, w13510, w13511, w13512, w13513, w13514, w13515, w13516, w13517, w13518, w13519, w13520, w13521, w13522, w13523, w13524, w13525, w13526, w13527, w13528, w13529, w13530, w13531, w13532, w13533, w13534, w13535, w13536, w13537, w13538, w13539, w13540, w13541, w13542, w13543, w13544, w13545, w13546, w13547, w13548, w13549, w13550, w13551, w13552, w13553, w13554, w13555, w13556, w13557, w13558, w13559, w13560, w13561, w13562, w13563, w13564, w13565, w13566, w13567, w13568, w13569, w13570, w13571, w13572, w13573, w13574, w13575, w13576, w13577, w13578, w13579, w13580, w13581, w13582, w13583, w13584, w13585, w13586, w13587, w13588, w13589, w13590, w13591, w13592, w13593, w13594, w13595, w13596, w13597, w13598, w13599, w13600, w13601, w13602, w13603, w13604, w13605, w13606, w13607, w13608, w13609, w13610, w13611, w13612, w13613, w13614, w13615, w13616, w13617, w13618, w13619, w13620, w13621, w13622, w13623, w13624, w13625, w13626, w13627, w13628, w13629, w13630, w13631, w13632, w13633, w13634, w13635, w13636, w13637, w13638, w13639, w13640, w13641, w13642, w13643, w13644, w13645, w13646, w13647, w13648, w13649, w13650, w13651, w13652, w13653, w13654, w13655, w13656, w13657, w13658, w13659, w13660, w13661, w13662, w13663, w13664, w13665, w13666, w13667, w13668, w13669, w13670, w13671, w13672, w13673, w13674, w13675, w13676, w13677, w13678, w13679, w13680, w13681, w13682, w13683, w13684, w13685, w13686, w13687, w13688, w13689, w13690, w13691, w13692, w13693, w13694, w13695, w13696, w13697, w13698, w13699, w13700, w13701, w13702, w13703, w13704, w13705, w13706, w13707, w13708, w13709, w13710, w13711, w13712, w13713, w13714, w13715, w13716, w13717, w13718, w13719, w13720, w13721, w13722, w13723, w13724, w13725, w13726, w13727, w13728, w13729, w13730, w13731, w13732, w13733, w13734, w13735, w13736, w13737, w13738, w13739, w13740, w13741, w13742, w13743, w13744, w13745, w13746, w13747, w13748, w13749, w13750, w13751, w13752, w13753, w13754, w13755, w13756, w13757, w13758, w13759, w13760, w13761, w13762, w13763, w13764, w13765, w13766, w13767, w13768, w13769, w13770, w13771, w13772, w13773, w13774, w13775, w13776, w13777, w13778, w13779, w13780, w13781, w13782, w13783, w13784, w13785, w13786, w13787, w13788, w13789, w13790, w13791, w13792, w13793, w13794, w13795, w13796, w13797, w13798, w13799, w13800, w13801, w13802, w13803, w13804, w13805, w13806, w13807, w13808, w13809, w13810, w13811, w13812, w13813, w13814, w13815, w13816, w13817, w13818, w13819, w13820, w13821, w13822, w13823, w13824, w13825, w13826, w13827, w13828, w13829, w13830, w13831, w13832, w13833, w13834, w13835, w13836, w13837, w13838, w13839, w13840, w13841, w13842, w13843, w13844, w13845, w13846, w13847, w13848, w13849, w13850, w13851, w13852, w13853, w13854, w13855, w13856, w13857, w13858, w13859, w13860, w13861, w13862, w13863, w13864, w13865, w13866, w13867, w13868, w13869, w13870, w13871, w13872, w13873, w13874, w13875, w13876, w13877, w13878, w13879, w13880, w13881, w13882, w13883, w13884, w13885, w13886, w13887, w13888, w13889, w13890, w13891, w13892, w13893, w13894, w13895, w13896, w13897, w13898, w13899, w13900, w13901, w13902, w13903, w13904, w13905, w13906, w13907, w13908, w13909, w13910, w13911, w13912, w13913, w13914, w13915, w13916, w13917, w13918, w13919, w13920, w13921, w13922, w13923, w13924, w13925, w13926, w13927, w13928, w13929, w13930, w13931, w13932, w13933, w13934, w13935, w13936, w13937, w13938, w13939, w13940, w13941, w13942, w13943, w13944, w13945, w13946, w13947, w13948, w13949, w13950, w13951, w13952, w13953, w13954, w13955, w13956, w13957, w13958, w13959, w13960, w13961, w13962, w13963, w13964, w13965, w13966, w13967, w13968, w13969, w13970, w13971, w13972, w13973, w13974, w13975, w13976, w13977, w13978, w13979, w13980, w13981, w13982, w13983, w13984, w13985, w13986, w13987, w13988, w13989, w13990, w13991, w13992, w13993, w13994, w13995, w13996, w13997, w13998, w13999, w14000, w14001, w14002, w14003, w14004, w14005, w14006, w14007, w14008, w14009, w14010, w14011, w14012, w14013, w14014, w14015, w14016, w14017, w14018, w14019, w14020, w14021, w14022, w14023, w14024, w14025, w14026, w14027, w14028, w14029, w14030, w14031, w14032, w14033, w14034, w14035, w14036, w14037, w14038, w14039, w14040, w14041, w14042, w14043, w14044, w14045, w14046, w14047, w14048, w14049, w14050, w14051, w14052, w14053, w14054, w14055, w14056, w14057, w14058, w14059, w14060, w14061, w14062, w14063, w14064, w14065, w14066, w14067, w14068, w14069, w14070, w14071, w14072, w14073, w14074, w14075, w14076, w14077, w14078, w14079, w14080, w14081, w14082, w14083, w14084, w14085, w14086, w14087, w14088, w14089, w14090, w14091, w14092, w14093, w14094, w14095, w14096, w14097, w14098, w14099, w14100, w14101, w14102, w14103, w14104, w14105, w14106, w14107, w14108, w14109, w14110, w14111, w14112, w14113, w14114, w14115, w14116, w14117, w14118, w14119, w14120, w14121, w14122, w14123, w14124, w14125, w14126, w14127, w14128, w14129, w14130, w14131, w14132, w14133, w14134, w14135, w14136, w14137, w14138, w14139, w14140, w14141, w14142, w14143, w14144, w14145, w14146, w14147, w14148, w14149, w14150, w14151, w14152, w14153, w14154, w14155, w14156, w14157, w14158, w14159, w14160, w14161, w14162, w14163, w14164, w14165, w14166, w14167, w14168, w14169, w14170, w14171, w14172, w14173, w14174, w14175, w14176, w14177, w14178, w14179, w14180, w14181, w14182, w14183, w14184, w14185, w14186, w14187, w14188, w14189, w14190, w14191, w14192, w14193, w14194, w14195, w14196, w14197, w14198, w14199, w14200, w14201, w14202, w14203, w14204, w14205, w14206, w14207, w14208, w14209, w14210, w14211, w14212, w14213, w14214, w14215, w14216, w14217, w14218, w14219, w14220, w14221, w14222, w14223, w14224, w14225, w14226, w14227, w14228, w14229, w14230, w14231, w14232, w14233, w14234, w14235, w14236, w14237, w14238, w14239, w14240, w14241, w14242, w14243, w14244, w14245, w14246, w14247, w14248, w14249, w14250, w14251, w14252, w14253, w14254, w14255, w14256, w14257, w14258, w14259, w14260, w14261, w14262, w14263, w14264, w14265, w14266, w14267, w14268, w14269, w14270, w14271, w14272, w14273, w14274, w14275, w14276, w14277, w14278, w14279, w14280, w14281, w14282, w14283, w14284, w14285, w14286, w14287, w14288, w14289, w14290, w14291, w14292, w14293, w14294, w14295, w14296, w14297, w14298, w14299, w14300, w14301, w14302, w14303, w14304, w14305, w14306, w14307, w14308, w14309, w14310, w14311, w14312, w14313, w14314, w14315, w14316, w14317, w14318, w14319, w14320, w14321, w14322, w14323, w14324, w14325, w14326, w14327, w14328, w14329, w14330, w14331, w14332, w14333, w14334, w14335, w14336, w14337, w14338, w14339, w14340, w14341, w14342, w14343, w14344, w14345, w14346, w14347, w14348, w14349, w14350, w14351, w14352, w14353, w14354, w14355, w14356, w14357, w14358, w14359, w14360, w14361, w14362, w14363, w14364, w14365, w14366, w14367, w14368, w14369, w14370, w14371, w14372, w14373, w14374, w14375, w14376, w14377, w14378, w14379, w14380, w14381, w14382, w14383, w14384, w14385, w14386, w14387, w14388, w14389, w14390, w14391, w14392, w14393, w14394, w14395, w14396, w14397, w14398, w14399, w14400, w14401, w14402, w14403, w14404, w14405, w14406, w14407, w14408, w14409, w14410, w14411, w14412, w14413, w14414, w14415, w14416, w14417, w14418, w14419, w14420, w14421, w14422, w14423, w14424, w14425, w14426, w14427, w14428, w14429, w14430, w14431, w14432, w14433, w14434, w14435, w14436, w14437, w14438, w14439, w14440, w14441, w14442, w14443, w14444, w14445, w14446, w14447, w14448, w14449, w14450, w14451, w14452, w14453, w14454, w14455, w14456, w14457, w14458, w14459, w14460, w14461, w14462, w14463, w14464, w14465, w14466, w14467, w14468, w14469, w14470, w14471, w14472, w14473, w14474, w14475, w14476, w14477, w14478, w14479, w14480, w14481, w14482, w14483, w14484, w14485, w14486, w14487, w14488, w14489, w14490, w14491, w14492, w14493, w14494, w14495, w14496, w14497, w14498, w14499, w14500, w14501, w14502, w14503, w14504, w14505, w14506, w14507, w14508, w14509, w14510, w14511, w14512, w14513, w14514, w14515, w14516, w14517, w14518, w14519, w14520, w14521, w14522, w14523, w14524, w14525, w14526, w14527, w14528, w14529, w14530, w14531, w14532, w14533, w14534, w14535, w14536, w14537, w14538, w14539, w14540, w14541, w14542, w14543, w14544, w14545, w14546, w14547, w14548, w14549, w14550, w14551, w14552, w14553, w14554, w14555, w14556, w14557, w14558, w14559, w14560, w14561, w14562, w14563, w14564, w14565, w14566, w14567, w14568, w14569, w14570, w14571, w14572, w14573, w14574, w14575, w14576, w14577, w14578, w14579, w14580, w14581, w14582, w14583, w14584, w14585, w14586, w14587, w14588, w14589, w14590, w14591, w14592, w14593, w14594, w14595, w14596, w14597, w14598, w14599, w14600, w14601, w14602, w14603, w14604, w14605, w14606, w14607, w14608, w14609, w14610, w14611, w14612, w14613, w14614, w14615, w14616, w14617, w14618, w14619, w14620, w14621, w14622, w14623, w14624, w14625, w14626, w14627, w14628, w14629, w14630, w14631, w14632, w14633, w14634, w14635, w14636, w14637, w14638, w14639, w14640, w14641, w14642, w14643, w14644, w14645, w14646, w14647, w14648, w14649, w14650, w14651, w14652, w14653, w14654, w14655, w14656, w14657, w14658, w14659, w14660, w14661, w14662, w14663, w14664, w14665, w14666, w14667, w14668, w14669, w14670, w14671, w14672, w14673, w14674, w14675, w14676, w14677, w14678, w14679, w14680, w14681, w14682, w14683, w14684, w14685, w14686, w14687, w14688, w14689, w14690, w14691, w14692, w14693, w14694, w14695, w14696, w14697, w14698, w14699, w14700, w14701, w14702, w14703, w14704, w14705, w14706, w14707, w14708, w14709, w14710, w14711, w14712, w14713, w14714, w14715, w14716, w14717, w14718, w14719, w14720, w14721, w14722, w14723, w14724, w14725, w14726, w14727, w14728, w14729, w14730, w14731, w14732, w14733, w14734, w14735, w14736, w14737, w14738, w14739, w14740, w14741, w14742, w14743, w14744, w14745, w14746, w14747, w14748, w14749, w14750, w14751, w14752, w14753, w14754, w14755, w14756, w14757, w14758, w14759, w14760, w14761, w14762, w14763, w14764, w14765, w14766, w14767, w14768, w14769, w14770, w14771, w14772, w14773, w14774, w14775, w14776, w14777, w14778, w14779, w14780, w14781, w14782, w14783, w14784, w14785, w14786, w14787, w14788, w14789, w14790, w14791, w14792, w14793, w14794, w14795, w14796, w14797, w14798, w14799, w14800, w14801, w14802, w14803, w14804, w14805, w14806, w14807, w14808, w14809, w14810, w14811, w14812, w14813, w14814, w14815, w14816, w14817, w14818, w14819, w14820, w14821, w14822, w14823, w14824, w14825, w14826, w14827, w14828, w14829, w14830, w14831, w14832, w14833, w14834, w14835, w14836, w14837, w14838, w14839, w14840, w14841, w14842, w14843, w14844, w14845, w14846, w14847, w14848, w14849, w14850, w14851, w14852, w14853, w14854, w14855, w14856, w14857, w14858, w14859, w14860, w14861, w14862, w14863, w14864, w14865, w14866, w14867, w14868, w14869, w14870, w14871, w14872, w14873, w14874, w14875, w14876, w14877, w14878, w14879, w14880, w14881, w14882, w14883, w14884, w14885, w14886, w14887, w14888, w14889, w14890, w14891, w14892, w14893, w14894, w14895, w14896, w14897, w14898, w14899, w14900, w14901, w14902, w14903, w14904, w14905, w14906, w14907, w14908, w14909, w14910, w14911, w14912, w14913, w14914, w14915, w14916, w14917, w14918, w14919, w14920, w14921, w14922, w14923, w14924, w14925, w14926, w14927, w14928, w14929, w14930, w14931, w14932, w14933, w14934, w14935, w14936, w14937, w14938, w14939, w14940, w14941, w14942, w14943, w14944, w14945, w14946, w14947, w14948, w14949, w14950, w14951, w14952, w14953, w14954, w14955, w14956, w14957, w14958, w14959, w14960, w14961, w14962, w14963, w14964, w14965, w14966, w14967, w14968, w14969, w14970, w14971, w14972, w14973, w14974, w14975, w14976, w14977, w14978, w14979, w14980, w14981, w14982, w14983, w14984, w14985, w14986, w14987, w14988, w14989, w14990, w14991, w14992, w14993, w14994, w14995, w14996, w14997, w14998, w14999, w15000, w15001, w15002, w15003, w15004, w15005, w15006, w15007, w15008, w15009, w15010, w15011, w15012, w15013, w15014, w15015, w15016, w15017, w15018, w15019, w15020, w15021, w15022, w15023, w15024, w15025, w15026, w15027, w15028, w15029, w15030, w15031, w15032, w15033, w15034, w15035, w15036, w15037, w15038, w15039, w15040, w15041, w15042, w15043, w15044, w15045, w15046, w15047, w15048, w15049, w15050, w15051, w15052, w15053, w15054, w15055, w15056, w15057, w15058, w15059, w15060, w15061, w15062, w15063, w15064, w15065, w15066, w15067, w15068, w15069, w15070, w15071, w15072, w15073, w15074, w15075, w15076, w15077, w15078, w15079, w15080, w15081, w15082, w15083, w15084, w15085, w15086, w15087, w15088, w15089, w15090, w15091, w15092, w15093, w15094, w15095, w15096, w15097, w15098, w15099, w15100, w15101, w15102, w15103, w15104, w15105, w15106, w15107, w15108, w15109, w15110, w15111, w15112, w15113, w15114, w15115, w15116, w15117, w15118, w15119, w15120, w15121, w15122, w15123, w15124, w15125, w15126, w15127, w15128, w15129, w15130, w15131, w15132, w15133, w15134, w15135, w15136, w15137, w15138, w15139, w15140, w15141, w15142, w15143, w15144, w15145, w15146, w15147, w15148, w15149, w15150, w15151, w15152, w15153, w15154, w15155, w15156, w15157, w15158, w15159, w15160, w15161, w15162, w15163, w15164, w15165, w15166, w15167, w15168, w15169, w15170, w15171, w15172, w15173, w15174, w15175, w15176, w15177, w15178, w15179, w15180, w15181, w15182, w15183, w15184, w15185, w15186, w15187, w15188, w15189, w15190, w15191, w15192, w15193, w15194, w15195, w15196, w15197, w15198, w15199, w15200, w15201, w15202, w15203, w15204, w15205, w15206, w15207, w15208, w15209, w15210, w15211, w15212, w15213, w15214, w15215, w15216, w15217, w15218, w15219, w15220, w15221, w15222, w15223, w15224, w15225, w15226, w15227, w15228, w15229, w15230, w15231, w15232, w15233, w15234, w15235, w15236, w15237, w15238, w15239, w15240, w15241, w15242, w15243, w15244, w15245, w15246, w15247, w15248, w15249, w15250, w15251, w15252, w15253, w15254, w15255, w15256, w15257, w15258, w15259, w15260, w15261, w15262, w15263, w15264, w15265, w15266, w15267, w15268, w15269, w15270, w15271, w15272, w15273, w15274, w15275, w15276, w15277, w15278, w15279, w15280, w15281, w15282, w15283, w15284, w15285, w15286, w15287, w15288, w15289, w15290, w15291, w15292, w15293, w15294, w15295, w15296, w15297, w15298, w15299, w15300, w15301, w15302, w15303, w15304, w15305, w15306, w15307, w15308, w15309, w15310, w15311, w15312, w15313, w15314, w15315, w15316, w15317, w15318, w15319, w15320, w15321, w15322, w15323, w15324, w15325, w15326, w15327, w15328, w15329, w15330, w15331, w15332, w15333, w15334, w15335, w15336, w15337, w15338, w15339, w15340, w15341, w15342, w15343, w15344, w15345, w15346, w15347, w15348, w15349, w15350, w15351, w15352, w15353, w15354, w15355, w15356, w15357, w15358, w15359, w15360, w15361, w15362, w15363, w15364, w15365, w15366, w15367, w15368, w15369, w15370, w15371, w15372, w15373, w15374, w15375, w15376, w15377, w15378, w15379, w15380, w15381, w15382, w15383, w15384, w15385, w15386, w15387, w15388, w15389, w15390, w15391, w15392, w15393, w15394, w15395, w15396, w15397, w15398, w15399, w15400, w15401, w15402, w15403, w15404, w15405, w15406, w15407, w15408, w15409, w15410, w15411, w15412, w15413, w15414, w15415, w15416, w15417, w15418, w15419, w15420, w15421, w15422, w15423, w15424, w15425, w15426, w15427, w15428, w15429, w15430, w15431, w15432, w15433, w15434, w15435, w15436, w15437, w15438, w15439, w15440, w15441, w15442, w15443, w15444, w15445, w15446, w15447, w15448, w15449, w15450, w15451, w15452, w15453, w15454, w15455, w15456, w15457, w15458, w15459, w15460, w15461, w15462, w15463, w15464, w15465, w15466, w15467, w15468, w15469, w15470, w15471, w15472, w15473, w15474, w15475, w15476, w15477, w15478, w15479, w15480, w15481, w15482, w15483, w15484, w15485, w15486, w15487, w15488, w15489, w15490, w15491, w15492, w15493, w15494, w15495, w15496, w15497, w15498, w15499, w15500, w15501, w15502, w15503, w15504, w15505, w15506, w15507, w15508, w15509, w15510, w15511, w15512, w15513, w15514, w15515, w15516, w15517, w15518, w15519, w15520, w15521, w15522, w15523, w15524, w15525, w15526, w15527, w15528, w15529, w15530, w15531, w15532, w15533, w15534, w15535, w15536, w15537, w15538, w15539, w15540, w15541, w15542, w15543, w15544, w15545, w15546, w15547, w15548, w15549, w15550, w15551, w15552, w15553, w15554, w15555, w15556, w15557, w15558, w15559, w15560, w15561, w15562, w15563, w15564, w15565, w15566, w15567, w15568, w15569, w15570, w15571, w15572, w15573, w15574, w15575, w15576, w15577, w15578, w15579, w15580, w15581, w15582, w15583, w15584, w15585, w15586, w15587, w15588, w15589, w15590, w15591, w15592, w15593, w15594, w15595, w15596, w15597, w15598, w15599, w15600, w15601, w15602, w15603, w15604, w15605, w15606, w15607, w15608, w15609, w15610, w15611, w15612, w15613, w15614, w15615, w15616, w15617, w15618, w15619, w15620, w15621, w15622, w15623, w15624, w15625, w15626, w15627, w15628, w15629, w15630, w15631, w15632, w15633, w15634, w15635, w15636, w15637, w15638, w15639, w15640, w15641, w15642, w15643, w15644, w15645, w15646, w15647, w15648, w15649, w15650, w15651, w15652, w15653, w15654, w15655, w15656, w15657, w15658, w15659, w15660, w15661, w15662, w15663, w15664, w15665, w15666, w15667, w15668, w15669, w15670, w15671, w15672, w15673, w15674, w15675, w15676, w15677, w15678, w15679, w15680, w15681, w15682, w15683, w15684, w15685, w15686, w15687, w15688, w15689, w15690, w15691, w15692, w15693, w15694, w15695, w15696, w15697, w15698, w15699, w15700, w15701, w15702, w15703, w15704, w15705, w15706, w15707, w15708, w15709, w15710, w15711, w15712, w15713, w15714, w15715, w15716, w15717, w15718, w15719, w15720, w15721, w15722, w15723, w15724, w15725, w15726, w15727, w15728, w15729, w15730, w15731, w15732, w15733, w15734, w15735, w15736, w15737, w15738, w15739, w15740, w15741, w15742, w15743, w15744, w15745, w15746, w15747, w15748, w15749, w15750, w15751, w15752, w15753, w15754, w15755, w15756, w15757, w15758, w15759, w15760, w15761, w15762, w15763, w15764, w15765, w15766, w15767, w15768, w15769, w15770, w15771, w15772, w15773, w15774, w15775, w15776, w15777, w15778, w15779, w15780, w15781, w15782, w15783, w15784, w15785, w15786, w15787, w15788, w15789, w15790, w15791, w15792, w15793, w15794, w15795, w15796, w15797, w15798, w15799, w15800, w15801, w15802, w15803, w15804, w15805, w15806, w15807, w15808, w15809, w15810, w15811, w15812, w15813, w15814, w15815, w15816, w15817, w15818, w15819, w15820, w15821, w15822, w15823, w15824, w15825, w15826, w15827, w15828, w15829, w15830, w15831, w15832, w15833, w15834, w15835, w15836, w15837, w15838, w15839, w15840, w15841, w15842, w15843, w15844, w15845, w15846, w15847, w15848, w15849, w15850, w15851, w15852, w15853, w15854, w15855, w15856, w15857, w15858, w15859, w15860, w15861, w15862, w15863, w15864, w15865, w15866, w15867, w15868, w15869, w15870, w15871, w15872, w15873, w15874, w15875, w15876, w15877, w15878, w15879, w15880, w15881, w15882, w15883, w15884, w15885, w15886, w15887, w15888, w15889, w15890, w15891, w15892, w15893, w15894, w15895, w15896, w15897, w15898, w15899, w15900, w15901, w15902, w15903, w15904, w15905, w15906, w15907, w15908, w15909, w15910, w15911, w15912, w15913, w15914, w15915, w15916, w15917, w15918, w15919, w15920, w15921, w15922, w15923, w15924, w15925, w15926, w15927, w15928, w15929, w15930, w15931, w15932, w15933, w15934, w15935, w15936, w15937, w15938, w15939, w15940, w15941, w15942, w15943, w15944, w15945, w15946, w15947, w15948, w15949, w15950, w15951, w15952, w15953, w15954, w15955, w15956, w15957, w15958, w15959, w15960, w15961, w15962, w15963, w15964, w15965, w15966, w15967, w15968, w15969, w15970, w15971, w15972, w15973, w15974, w15975, w15976, w15977, w15978, w15979, w15980, w15981, w15982, w15983, w15984, w15985, w15986, w15987, w15988, w15989, w15990, w15991, w15992, w15993, w15994, w15995, w15996, w15997, w15998, w15999, w16000, w16001, w16002, w16003, w16004, w16005, w16006, w16007, w16008, w16009, w16010, w16011, w16012, w16013, w16014, w16015, w16016, w16017, w16018, w16019, w16020, w16021, w16022, w16023, w16024, w16025, w16026, w16027, w16028, w16029, w16030, w16031, w16032, w16033, w16034, w16035, w16036, w16037, w16038, w16039, w16040, w16041, w16042, w16043, w16044, w16045, w16046, w16047, w16048, w16049, w16050, w16051, w16052, w16053, w16054, w16055, w16056, w16057, w16058, w16059, w16060, w16061, w16062, w16063, w16064, w16065, w16066, w16067, w16068, w16069, w16070, w16071, w16072, w16073, w16074, w16075, w16076, w16077, w16078, w16079, w16080, w16081, w16082, w16083, w16084, w16085, w16086, w16087, w16088, w16089, w16090, w16091, w16092, w16093, w16094, w16095, w16096, w16097, w16098, w16099, w16100, w16101, w16102, w16103, w16104, w16105, w16106, w16107, w16108, w16109, w16110, w16111, w16112, w16113, w16114, w16115, w16116, w16117, w16118, w16119, w16120, w16121, w16122, w16123, w16124, w16125, w16126, w16127, w16128, w16129, w16130, w16131, w16132, w16133, w16134, w16135, w16136, w16137, w16138, w16139, w16140, w16141, w16142, w16143, w16144, w16145, w16146, w16147, w16148, w16149, w16150, w16151, w16152, w16153, w16154, w16155, w16156, w16157, w16158, w16159, w16160, w16161, w16162, w16163, w16164, w16165, w16166, w16167, w16168, w16169, w16170, w16171, w16172, w16173, w16174, w16175, w16176, w16177, w16178, w16179, w16180, w16181, w16182, w16183, w16184, w16185, w16186, w16187, w16188, w16189, w16190, w16191, w16192, w16193, w16194, w16195, w16196, w16197, w16198, w16199, w16200, w16201, w16202, w16203, w16204, w16205, w16206, w16207, w16208, w16209, w16210, w16211, w16212, w16213, w16214, w16215, w16216, w16217, w16218, w16219, w16220, w16221, w16222, w16223, w16224, w16225, w16226, w16227, w16228, w16229, w16230, w16231, w16232, w16233, w16234, w16235, w16236, w16237, w16238, w16239, w16240, w16241, w16242, w16243, w16244, w16245, w16246, w16247, w16248, w16249, w16250, w16251, w16252, w16253, w16254, w16255, w16256, w16257, w16258, w16259, w16260, w16261, w16262, w16263, w16264, w16265, w16266, w16267, w16268, w16269, w16270, w16271, w16272, w16273, w16274, w16275, w16276, w16277, w16278, w16279, w16280, w16281, w16282, w16283, w16284, w16285, w16286, w16287, w16288, w16289, w16290, w16291, w16292, w16293, w16294, w16295, w16296, w16297, w16298, w16299, w16300, w16301, w16302, w16303, w16304, w16305, w16306, w16307, w16308, w16309, w16310, w16311, w16312, w16313, w16314, w16315, w16316, w16317, w16318, w16319, w16320, w16321, w16322, w16323, w16324, w16325, w16326, w16327, w16328, w16329, w16330, w16331, w16332, w16333, w16334, w16335, w16336, w16337, w16338, w16339, w16340, w16341, w16342, w16343, w16344, w16345, w16346, w16347, w16348, w16349, w16350, w16351, w16352, w16353, w16354, w16355, w16356, w16357, w16358, w16359, w16360, w16361, w16362, w16363, w16364, w16365, w16366, w16367, w16368, w16369, w16370, w16371, w16372, w16373, w16374, w16375, w16376, w16377, w16378, w16379, w16380, w16381, w16382, w16383, w16384, w16385, w16386, w16387, w16388, w16389, w16390, w16391, w16392, w16393, w16394, w16395, w16396, w16397, w16398, w16399, w16400, w16401, w16402, w16403, w16404, w16405, w16406, w16407, w16408, w16409, w16410, w16411, w16412, w16413, w16414, w16415, w16416, w16417, w16418, w16419, w16420, w16421, w16422, w16423, w16424, w16425, w16426, w16427, w16428, w16429, w16430, w16431, w16432, w16433, w16434, w16435, w16436, w16437, w16438, w16439, w16440, w16441, w16442, w16443, w16444, w16445, w16446, w16447, w16448, w16449, w16450, w16451, w16452, w16453, w16454, w16455, w16456, w16457, w16458, w16459, w16460, w16461, w16462, w16463, w16464, w16465, w16466, w16467, w16468, w16469, w16470, w16471, w16472, w16473, w16474, w16475, w16476, w16477, w16478, w16479, w16480, w16481, w16482, w16483, w16484, w16485, w16486, w16487, w16488, w16489, w16490, w16491, w16492, w16493, w16494, w16495, w16496, w16497, w16498, w16499, w16500, w16501, w16502, w16503, w16504, w16505, w16506, w16507, w16508, w16509, w16510, w16511, w16512, w16513, w16514, w16515, w16516, w16517, w16518, w16519, w16520, w16521, w16522, w16523, w16524, w16525, w16526, w16527, w16528, w16529, w16530, w16531, w16532, w16533, w16534, w16535, w16536, w16537, w16538, w16539, w16540, w16541, w16542, w16543, w16544, w16545, w16546, w16547, w16548, w16549, w16550, w16551, w16552, w16553, w16554, w16555, w16556, w16557, w16558, w16559, w16560, w16561, w16562, w16563, w16564, w16565, w16566, w16567, w16568, w16569, w16570, w16571, w16572, w16573, w16574, w16575, w16576, w16577, w16578, w16579, w16580, w16581, w16582, w16583, w16584, w16585, w16586, w16587, w16588, w16589, w16590, w16591, w16592, w16593, w16594, w16595, w16596, w16597, w16598, w16599, w16600, w16601, w16602, w16603, w16604, w16605, w16606, w16607, w16608, w16609, w16610, w16611, w16612, w16613, w16614, w16615, w16616, w16617, w16618, w16619, w16620, w16621, w16622, w16623, w16624, w16625, w16626, w16627, w16628, w16629, w16630, w16631, w16632, w16633, w16634, w16635, w16636, w16637, w16638, w16639, w16640, w16641, w16642, w16643, w16644, w16645, w16646, w16647, w16648, w16649, w16650, w16651, w16652, w16653, w16654, w16655, w16656, w16657, w16658, w16659, w16660, w16661, w16662, w16663, w16664, w16665, w16666, w16667, w16668, w16669, w16670, w16671, w16672, w16673, w16674, w16675, w16676, w16677, w16678, w16679, w16680, w16681, w16682, w16683, w16684, w16685, w16686, w16687, w16688, w16689, w16690, w16691, w16692, w16693, w16694, w16695, w16696, w16697, w16698, w16699, w16700, w16701, w16702, w16703, w16704, w16705, w16706, w16707, w16708, w16709, w16710, w16711, w16712, w16713, w16714, w16715, w16716, w16717, w16718, w16719, w16720, w16721, w16722, w16723, w16724, w16725, w16726, w16727, w16728, w16729, w16730, w16731, w16732, w16733, w16734, w16735, w16736, w16737, w16738, w16739, w16740, w16741, w16742, w16743, w16744, w16745, w16746, w16747, w16748, w16749, w16750, w16751, w16752, w16753, w16754, w16755, w16756, w16757, w16758, w16759, w16760, w16761, w16762, w16763, w16764, w16765, w16766, w16767, w16768, w16769, w16770, w16771, w16772, w16773, w16774, w16775, w16776, w16777, w16778, w16779, w16780, w16781, w16782, w16783, w16784, w16785, w16786, w16787, w16788, w16789, w16790, w16791, w16792, w16793, w16794, w16795, w16796, w16797, w16798, w16799, w16800, w16801, w16802, w16803, w16804, w16805, w16806, w16807, w16808, w16809, w16810, w16811, w16812, w16813, w16814, w16815, w16816, w16817, w16818, w16819, w16820, w16821, w16822, w16823, w16824, w16825, w16826, w16827, w16828, w16829, w16830, w16831, w16832, w16833, w16834, w16835, w16836, w16837, w16838, w16839, w16840, w16841, w16842, w16843, w16844, w16845, w16846, w16847, w16848, w16849, w16850, w16851, w16852, w16853, w16854, w16855, w16856, w16857, w16858, w16859, w16860, w16861, w16862, w16863, w16864, w16865, w16866, w16867, w16868, w16869, w16870, w16871, w16872, w16873, w16874, w16875, w16876, w16877, w16878, w16879, w16880, w16881, w16882, w16883, w16884, w16885, w16886, w16887, w16888, w16889, w16890, w16891, w16892, w16893, w16894, w16895, w16896, w16897, w16898, w16899, w16900, w16901, w16902, w16903, w16904, w16905, w16906, w16907, w16908, w16909, w16910, w16911, w16912, w16913, w16914, w16915, w16916, w16917, w16918, w16919, w16920, w16921, w16922, w16923, w16924, w16925, w16926, w16927, w16928, w16929, w16930, w16931, w16932, w16933, w16934, w16935, w16936, w16937, w16938, w16939, w16940, w16941, w16942, w16943, w16944, w16945, w16946, w16947, w16948, w16949, w16950, w16951, w16952, w16953, w16954, w16955, w16956, w16957, w16958, w16959, w16960, w16961, w16962, w16963, w16964, w16965, w16966, w16967, w16968, w16969, w16970, w16971, w16972, w16973, w16974, w16975, w16976, w16977, w16978, w16979, w16980, w16981, w16982, w16983, w16984, w16985, w16986, w16987, w16988, w16989, w16990, w16991, w16992, w16993, w16994, w16995, w16996, w16997, w16998, w16999, w17000, w17001, w17002, w17003, w17004, w17005, w17006, w17007, w17008, w17009, w17010, w17011, w17012, w17013, w17014, w17015, w17016, w17017, w17018, w17019, w17020, w17021, w17022, w17023, w17024, w17025, w17026, w17027, w17028, w17029, w17030, w17031, w17032, w17033, w17034, w17035, w17036, w17037, w17038, w17039, w17040, w17041, w17042, w17043, w17044, w17045, w17046, w17047, w17048, w17049, w17050, w17051, w17052, w17053, w17054, w17055, w17056, w17057, w17058, w17059, w17060, w17061, w17062, w17063, w17064, w17065, w17066, w17067, w17068, w17069, w17070, w17071, w17072, w17073, w17074, w17075, w17076, w17077, w17078, w17079, w17080, w17081, w17082, w17083, w17084, w17085, w17086, w17087, w17088, w17089, w17090, w17091, w17092, w17093, w17094, w17095, w17096, w17097, w17098, w17099, w17100, w17101, w17102, w17103, w17104, w17105, w17106, w17107, w17108, w17109, w17110, w17111, w17112, w17113, w17114, w17115, w17116, w17117, w17118, w17119, w17120, w17121, w17122, w17123, w17124, w17125, w17126, w17127, w17128, w17129, w17130, w17131, w17132, w17133, w17134, w17135, w17136, w17137, w17138, w17139, w17140, w17141, w17142, w17143, w17144, w17145, w17146, w17147, w17148, w17149, w17150, w17151, w17152, w17153, w17154, w17155, w17156, w17157, w17158, w17159, w17160, w17161, w17162, w17163, w17164, w17165, w17166, w17167, w17168, w17169, w17170, w17171, w17172, w17173, w17174, w17175, w17176, w17177, w17178, w17179, w17180, w17181, w17182, w17183, w17184, w17185, w17186, w17187, w17188, w17189, w17190, w17191, w17192, w17193, w17194, w17195, w17196, w17197, w17198, w17199, w17200, w17201, w17202, w17203, w17204, w17205, w17206, w17207, w17208, w17209, w17210, w17211, w17212, w17213, w17214, w17215, w17216, w17217, w17218, w17219, w17220, w17221, w17222, w17223, w17224, w17225, w17226, w17227, w17228, w17229, w17230, w17231, w17232, w17233, w17234, w17235, w17236, w17237, w17238, w17239, w17240, w17241, w17242, w17243, w17244, w17245, w17246, w17247, w17248, w17249, w17250, w17251, w17252, w17253, w17254, w17255, w17256, w17257, w17258, w17259, w17260, w17261, w17262, w17263, w17264, w17265, w17266, w17267, w17268, w17269, w17270, w17271, w17272, w17273, w17274, w17275, w17276, w17277, w17278, w17279, w17280, w17281, w17282, w17283, w17284, w17285, w17286, w17287, w17288, w17289, w17290, w17291, w17292, w17293, w17294, w17295, w17296, w17297, w17298, w17299, w17300, w17301, w17302, w17303, w17304, w17305, w17306, w17307, w17308, w17309, w17310, w17311, w17312, w17313, w17314, w17315, w17316, w17317, w17318, w17319, w17320, w17321, w17322, w17323, w17324, w17325, w17326, w17327, w17328, w17329, w17330, w17331, w17332, w17333, w17334, w17335, w17336, w17337, w17338, w17339, w17340, w17341, w17342, w17343, w17344, w17345, w17346, w17347, w17348, w17349, w17350, w17351, w17352, w17353, w17354, w17355, w17356, w17357, w17358, w17359, w17360, w17361, w17362, w17363, w17364, w17365, w17366, w17367, w17368, w17369, w17370, w17371, w17372, w17373, w17374, w17375, w17376, w17377, w17378, w17379, w17380, w17381, w17382, w17383, w17384, w17385, w17386, w17387, w17388, w17389, w17390, w17391, w17392, w17393, w17394, w17395, w17396, w17397, w17398, w17399, w17400, w17401, w17402, w17403, w17404, w17405, w17406, w17407, w17408, w17409, w17410, w17411, w17412, w17413, w17414, w17415, w17416, w17417, w17418, w17419, w17420, w17421, w17422, w17423, w17424, w17425, w17426, w17427, w17428, w17429, w17430, w17431, w17432, w17433, w17434, w17435, w17436, w17437, w17438, w17439, w17440, w17441, w17442, w17443, w17444, w17445, w17446, w17447, w17448, w17449, w17450, w17451, w17452, w17453, w17454, w17455, w17456, w17457, w17458, w17459, w17460, w17461, w17462, w17463, w17464, w17465, w17466, w17467, w17468, w17469, w17470, w17471, w17472, w17473, w17474, w17475, w17476, w17477, w17478, w17479, w17480, w17481, w17482, w17483, w17484, w17485, w17486, w17487, w17488, w17489, w17490, w17491, w17492, w17493, w17494, w17495, w17496, w17497, w17498, w17499, w17500, w17501, w17502, w17503, w17504, w17505, w17506, w17507, w17508, w17509, w17510, w17511, w17512, w17513, w17514, w17515, w17516, w17517, w17518, w17519, w17520, w17521, w17522, w17523, w17524, w17525, w17526, w17527, w17528, w17529, w17530, w17531, w17532, w17533, w17534, w17535, w17536, w17537, w17538, w17539, w17540, w17541, w17542, w17543, w17544, w17545, w17546, w17547, w17548, w17549, w17550, w17551, w17552, w17553, w17554, w17555, w17556, w17557, w17558, w17559, w17560, w17561, w17562, w17563, w17564, w17565, w17566, w17567, w17568, w17569, w17570, w17571, w17572, w17573, w17574, w17575, w17576, w17577, w17578, w17579, w17580, w17581, w17582, w17583, w17584, w17585, w17586, w17587, w17588, w17589, w17590, w17591, w17592, w17593, w17594, w17595, w17596, w17597, w17598, w17599, w17600, w17601, w17602, w17603, w17604, w17605, w17606, w17607, w17608, w17609, w17610, w17611, w17612, w17613, w17614, w17615, w17616, w17617, w17618, w17619, w17620, w17621, w17622, w17623, w17624, w17625, w17626, w17627, w17628, w17629, w17630, w17631, w17632, w17633, w17634, w17635, w17636, w17637, w17638, w17639, w17640, w17641, w17642, w17643, w17644, w17645, w17646, w17647, w17648, w17649, w17650, w17651, w17652, w17653, w17654, w17655, w17656, w17657, w17658, w17659, w17660, w17661, w17662, w17663, w17664, w17665, w17666, w17667, w17668, w17669, w17670, w17671, w17672, w17673, w17674, w17675, w17676, w17677, w17678, w17679, w17680, w17681, w17682, w17683, w17684, w17685, w17686, w17687, w17688, w17689, w17690, w17691, w17692, w17693, w17694, w17695, w17696, w17697, w17698, w17699, w17700, w17701, w17702, w17703, w17704, w17705, w17706, w17707, w17708, w17709, w17710, w17711, w17712, w17713, w17714, w17715, w17716, w17717, w17718, w17719, w17720, w17721, w17722, w17723, w17724, w17725, w17726, w17727, w17728, w17729, w17730, w17731, w17732, w17733, w17734, w17735, w17736, w17737, w17738, w17739, w17740, w17741, w17742, w17743, w17744, w17745, w17746, w17747, w17748, w17749, w17750, w17751, w17752, w17753, w17754, w17755, w17756, w17757, w17758, w17759, w17760, w17761, w17762, w17763, w17764, w17765, w17766, w17767, w17768, w17769, w17770, w17771, w17772, w17773, w17774, w17775, w17776, w17777, w17778, w17779, w17780, w17781, w17782, w17783, w17784, w17785, w17786, w17787, w17788, w17789, w17790, w17791, w17792, w17793, w17794, w17795, w17796, w17797, w17798, w17799, w17800, w17801, w17802, w17803, w17804, w17805, w17806, w17807, w17808, w17809, w17810, w17811, w17812, w17813, w17814, w17815, w17816, w17817, w17818, w17819, w17820, w17821, w17822, w17823, w17824, w17825, w17826, w17827, w17828, w17829, w17830, w17831, w17832, w17833, w17834, w17835, w17836, w17837, w17838, w17839, w17840, w17841, w17842, w17843, w17844, w17845, w17846, w17847, w17848, w17849, w17850, w17851, w17852, w17853, w17854, w17855, w17856, w17857, w17858, w17859, w17860, w17861, w17862, w17863, w17864, w17865, w17866, w17867, w17868, w17869, w17870, w17871, w17872, w17873, w17874, w17875, w17876, w17877, w17878, w17879, w17880, w17881, w17882, w17883, w17884, w17885, w17886;
assign w0 = ~pi00 & pi01;
assign w1 = ~pi01 & ~pi02;
assign w2 = pi01 & pi02;
assign w3 = pi00 & ~w1;
assign w4 = ~w2 & w3;
assign w5 = pi02 & pi03;
assign w6 = pi00 & w5;
assign w7 = pi00 & pi03;
assign w8 = pi02 & ~w0;
assign w9 = ~w7 & ~w8;
assign w10 = ~w6 & ~w9;
assign w11 = pi00 & pi04;
assign w12 = pi01 & pi03;
assign w13 = ~w11 & ~w12;
assign w14 = pi01 & pi04;
assign w15 = w7 & w14;
assign w16 = ~w13 & ~w15;
assign w17 = ~w2 & ~w16;
assign w18 = w2 & w16;
assign w19 = ~w17 & ~w18;
assign w20 = w6 & ~w19;
assign w21 = ~w6 & w19;
assign w22 = ~w20 & ~w21;
assign w23 = ~pi02 & pi03;
assign w24 = pi01 & pi05;
assign w25 = w11 & w24;
assign w26 = w15 & w25;
assign w27 = pi00 & pi05;
assign w28 = ~w14 & ~w27;
assign w29 = ~w15 & ~w25;
assign w30 = ~w28 & w29;
assign w31 = ~w30 & w16482;
assign w32 = (~w6 & ~w16) | (~w6 & w16483) | (~w16 & w16483);
assign w33 = ~w17 & ~w32;
assign w34 = w31 & ~w33;
assign w35 = (w23 & w30) | (w23 & w16484) | (w30 & w16484);
assign w36 = ~w31 & w33;
assign w37 = ~w35 & ~w36;
assign w38 = ~w34 & w37;
assign w39 = pi00 & pi06;
assign w40 = ~w5 & ~w39;
assign w41 = w5 & w39;
assign w42 = ~w40 & ~w41;
assign w43 = pi02 & pi04;
assign w44 = ~w24 & ~w43;
assign w45 = w24 & w43;
assign w46 = ~w44 & ~w45;
assign w47 = w42 & w46;
assign w48 = ~w42 & ~w46;
assign w49 = ~w47 & ~w48;
assign w50 = w29 & ~w49;
assign w51 = ~w29 & w49;
assign w52 = ~w50 & ~w51;
assign w53 = w37 & w52;
assign w54 = ~w37 & ~w52;
assign w55 = ~w53 & ~w54;
assign w56 = ~w41 & ~w47;
assign w57 = ~pi06 & w45;
assign w58 = pi01 & pi06;
assign w59 = ~pi04 & ~w58;
assign w60 = pi04 & w58;
assign w61 = ~w59 & ~w60;
assign w62 = ~w45 & ~w61;
assign w63 = ~w57 & ~w62;
assign w64 = ~w56 & w63;
assign w65 = w56 & ~w63;
assign w66 = ~w64 & ~w65;
assign w67 = pi00 & pi07;
assign w68 = pi02 & pi05;
assign w69 = pi03 & pi04;
assign w70 = ~w68 & ~w69;
assign w71 = w68 & w69;
assign w72 = ~w70 & ~w71;
assign w73 = w67 & ~w72;
assign w74 = ~w67 & w72;
assign w75 = ~w73 & ~w74;
assign w76 = ~w66 & w75;
assign w77 = w66 & ~w75;
assign w78 = ~w76 & ~w77;
assign w79 = ~w35 & ~w51;
assign w80 = (~w50 & ~w79) | (~w50 & w16485) | (~w79 & w16485);
assign w81 = w78 & w80;
assign w82 = ~w78 & ~w80;
assign w83 = ~w81 & ~w82;
assign w84 = ~w57 & ~w64;
assign w85 = pi03 & pi05;
assign w86 = pi01 & pi07;
assign w87 = ~w85 & ~w86;
assign w88 = w85 & w86;
assign w89 = ~w87 & ~w88;
assign w90 = ~w67 & ~w71;
assign w91 = ~w70 & ~w90;
assign w92 = w89 & w91;
assign w93 = ~w89 & ~w91;
assign w94 = ~w92 & ~w93;
assign w95 = pi02 & pi06;
assign w96 = pi00 & pi08;
assign w97 = ~w95 & ~w96;
assign w98 = pi02 & pi08;
assign w99 = w39 & w98;
assign w100 = ~w97 & ~w99;
assign w101 = w60 & ~w100;
assign w102 = ~w60 & w100;
assign w103 = ~w101 & ~w102;
assign w104 = w94 & ~w103;
assign w105 = ~w94 & w103;
assign w106 = ~w104 & ~w105;
assign w107 = w84 & ~w106;
assign w108 = ~w84 & w106;
assign w109 = ~w107 & ~w108;
assign w110 = ~w76 & w80;
assign w111 = ~w77 & ~w110;
assign w112 = w109 & w111;
assign w113 = ~w109 & ~w111;
assign w114 = ~w112 & ~w113;
assign w115 = ~w92 & ~w104;
assign w116 = pi08 & w24;
assign w117 = pi01 & pi08;
assign w118 = ~pi05 & ~w117;
assign w119 = ~w116 & ~w118;
assign w120 = pi00 & pi09;
assign w121 = w88 & w120;
assign w122 = ~w88 & ~w120;
assign w123 = ~w121 & ~w122;
assign w124 = w119 & w123;
assign w125 = ~w119 & ~w123;
assign w126 = ~w124 & ~w125;
assign w127 = w60 & ~w97;
assign w128 = ~w99 & ~w127;
assign w129 = pi02 & pi07;
assign w130 = pi04 & pi05;
assign w131 = pi03 & pi06;
assign w132 = ~w130 & ~w131;
assign w133 = w130 & w131;
assign w134 = ~w132 & ~w133;
assign w135 = w129 & ~w134;
assign w136 = ~w129 & w134;
assign w137 = ~w135 & ~w136;
assign w138 = ~w128 & ~w137;
assign w139 = w128 & w137;
assign w140 = ~w138 & ~w139;
assign w141 = w126 & w140;
assign w142 = ~w126 & ~w140;
assign w143 = ~w141 & ~w142;
assign w144 = ~w115 & w143;
assign w145 = w115 & ~w143;
assign w146 = ~w144 & ~w145;
assign w147 = ~w77 & ~w108;
assign w148 = (~w107 & ~w147) | (~w107 & w16486) | (~w147 & w16486);
assign w149 = w146 & w148;
assign w150 = ~w146 & ~w148;
assign w151 = ~w149 & ~w150;
assign w152 = ~w138 & ~w141;
assign w153 = pi04 & pi06;
assign w154 = pi01 & pi09;
assign w155 = ~w153 & ~w154;
assign w156 = w153 & w154;
assign w157 = ~w155 & ~w156;
assign w158 = w116 & w157;
assign w159 = ~w116 & ~w157;
assign w160 = ~w158 & ~w159;
assign w161 = ~w129 & ~w133;
assign w162 = ~w132 & ~w161;
assign w163 = w160 & w162;
assign w164 = ~w160 & ~w162;
assign w165 = ~w163 & ~w164;
assign w166 = (~w121 & ~w123) | (~w121 & w16487) | (~w123 & w16487);
assign w167 = pi03 & pi07;
assign w168 = pi00 & pi10;
assign w169 = ~w167 & ~w168;
assign w170 = w167 & w168;
assign w171 = ~w169 & ~w170;
assign w172 = w98 & ~w171;
assign w173 = ~w98 & w171;
assign w174 = ~w172 & ~w173;
assign w175 = ~w166 & ~w174;
assign w176 = w166 & w174;
assign w177 = ~w175 & ~w176;
assign w178 = w165 & w177;
assign w179 = ~w165 & ~w177;
assign w180 = ~w178 & ~w179;
assign w181 = ~w152 & w180;
assign w182 = w152 & ~w180;
assign w183 = ~w181 & ~w182;
assign w184 = ~w144 & ~w148;
assign w185 = ~w145 & ~w184;
assign w186 = w183 & w185;
assign w187 = ~w183 & ~w185;
assign w188 = ~w186 & ~w187;
assign w189 = ~w175 & ~w178;
assign w190 = pi10 & w58;
assign w191 = pi01 & pi10;
assign w192 = ~pi06 & ~w191;
assign w193 = ~w190 & ~w192;
assign w194 = ~w98 & ~w170;
assign w195 = ~w169 & ~w194;
assign w196 = w193 & w195;
assign w197 = ~w193 & ~w195;
assign w198 = ~w196 & ~w197;
assign w199 = pi03 & pi08;
assign w200 = pi02 & pi09;
assign w201 = ~w199 & ~w200;
assign w202 = w199 & w200;
assign w203 = ~w201 & ~w202;
assign w204 = w156 & ~w203;
assign w205 = ~w156 & w203;
assign w206 = ~w204 & ~w205;
assign w207 = w198 & ~w206;
assign w208 = ~w198 & w206;
assign w209 = ~w207 & ~w208;
assign w210 = (~w158 & ~w160) | (~w158 & w16488) | (~w160 & w16488);
assign w211 = pi00 & pi11;
assign w212 = pi05 & pi06;
assign w213 = pi04 & pi07;
assign w214 = ~w212 & ~w213;
assign w215 = w212 & w213;
assign w216 = ~w214 & ~w215;
assign w217 = w211 & ~w216;
assign w218 = ~w211 & w216;
assign w219 = ~w217 & ~w218;
assign w220 = ~w210 & ~w219;
assign w221 = w210 & w219;
assign w222 = ~w220 & ~w221;
assign w223 = w209 & w222;
assign w224 = ~w209 & ~w222;
assign w225 = ~w223 & ~w224;
assign w226 = w189 & ~w225;
assign w227 = ~w189 & w225;
assign w228 = ~w226 & ~w227;
assign w229 = ~w145 & ~w182;
assign w230 = ~w184 & w229;
assign w231 = ~w181 & ~w230;
assign w232 = w228 & w231;
assign w233 = ~w228 & ~w231;
assign w234 = ~w232 & ~w233;
assign w235 = ~w181 & ~w227;
assign w236 = (~w226 & w230) | (~w226 & w16489) | (w230 & w16489);
assign w237 = ~w220 & ~w223;
assign w238 = ~w211 & ~w215;
assign w239 = ~w214 & ~w238;
assign w240 = ~w156 & ~w202;
assign w241 = ~w201 & ~w240;
assign w242 = w239 & w241;
assign w243 = ~w239 & ~w241;
assign w244 = ~w242 & ~w243;
assign w245 = pi03 & pi09;
assign w246 = pi00 & pi12;
assign w247 = pi02 & pi10;
assign w248 = ~w246 & ~w247;
assign w249 = pi02 & pi12;
assign w250 = w168 & w249;
assign w251 = ~w248 & ~w250;
assign w252 = w245 & ~w251;
assign w253 = ~w245 & w251;
assign w254 = ~w252 & ~w253;
assign w255 = ~w244 & w254;
assign w256 = w244 & ~w254;
assign w257 = ~w255 & ~w256;
assign w258 = (~w196 & ~w198) | (~w196 & w16490) | (~w198 & w16490);
assign w259 = pi05 & pi07;
assign w260 = pi01 & pi11;
assign w261 = ~w259 & ~w260;
assign w262 = w259 & w260;
assign w263 = ~w261 & ~w262;
assign w264 = pi04 & pi08;
assign w265 = ~w190 & ~w264;
assign w266 = w190 & w264;
assign w267 = ~w265 & ~w266;
assign w268 = w263 & ~w267;
assign w269 = ~w263 & w267;
assign w270 = ~w268 & ~w269;
assign w271 = ~w258 & ~w270;
assign w272 = w258 & w270;
assign w273 = ~w271 & ~w272;
assign w274 = w257 & w273;
assign w275 = ~w257 & ~w273;
assign w276 = ~w274 & ~w275;
assign w277 = w237 & ~w276;
assign w278 = ~w237 & w276;
assign w279 = ~w277 & ~w278;
assign w280 = w236 & ~w279;
assign w281 = ~w236 & w279;
assign w282 = ~w280 & ~w281;
assign w283 = ~w236 & ~w278;
assign w284 = ~w277 & ~w283;
assign w285 = ~w242 & ~w256;
assign w286 = ~pi12 & w262;
assign w287 = pi12 & w86;
assign w288 = pi01 & pi12;
assign w289 = ~pi07 & ~w288;
assign w290 = ~w287 & ~w289;
assign w291 = ~w262 & ~w290;
assign w292 = ~w286 & ~w291;
assign w293 = w245 & ~w248;
assign w294 = ~w250 & ~w293;
assign w295 = ~w292 & w294;
assign w296 = w292 & ~w294;
assign w297 = ~w295 & ~w296;
assign w298 = ~w285 & w297;
assign w299 = w285 & ~w297;
assign w300 = ~w298 & ~w299;
assign w301 = (~w271 & ~w273) | (~w271 & w16491) | (~w273 & w16491);
assign w302 = ~w300 & w301;
assign w303 = w300 & ~w301;
assign w304 = ~w302 & ~w303;
assign w305 = pi03 & pi10;
assign w306 = pi04 & pi09;
assign w307 = pi00 & pi13;
assign w308 = ~w306 & ~w307;
assign w309 = w306 & w307;
assign w310 = ~w308 & ~w309;
assign w311 = w305 & ~w310;
assign w312 = ~w305 & w310;
assign w313 = ~w311 & ~w312;
assign w314 = w263 & ~w265;
assign w315 = ~w266 & ~w314;
assign w316 = ~w313 & ~w315;
assign w317 = w313 & w315;
assign w318 = ~w316 & ~w317;
assign w319 = pi02 & pi11;
assign w320 = pi06 & pi07;
assign w321 = pi05 & pi08;
assign w322 = ~w320 & ~w321;
assign w323 = w320 & w321;
assign w324 = ~w322 & ~w323;
assign w325 = w319 & ~w324;
assign w326 = ~w319 & w324;
assign w327 = ~w325 & ~w326;
assign w328 = w318 & ~w327;
assign w329 = ~w318 & w327;
assign w330 = ~w328 & ~w329;
assign w331 = ~w304 & ~w330;
assign w332 = w304 & w330;
assign w333 = ~w331 & ~w332;
assign w334 = w284 & w333;
assign w335 = ~w284 & ~w333;
assign w336 = ~w334 & ~w335;
assign w337 = ~w277 & ~w331;
assign w338 = ~w283 & w337;
assign w339 = ~w332 & ~w338;
assign w340 = ~w298 & ~w303;
assign w341 = pi04 & pi10;
assign w342 = pi05 & pi09;
assign w343 = ~w341 & ~w342;
assign w344 = w341 & w342;
assign w345 = ~w343 & ~w344;
assign w346 = w287 & ~w345;
assign w347 = ~w287 & w345;
assign w348 = ~w346 & ~w347;
assign w349 = pi00 & pi14;
assign w350 = pi03 & pi11;
assign w351 = ~w249 & ~w350;
assign w352 = w249 & w350;
assign w353 = ~w351 & ~w352;
assign w354 = w349 & ~w353;
assign w355 = ~w349 & w353;
assign w356 = ~w354 & ~w355;
assign w357 = ~w348 & ~w356;
assign w358 = w348 & w356;
assign w359 = ~w357 & ~w358;
assign w360 = (~w286 & ~w292) | (~w286 & w16807) | (~w292 & w16807);
assign w361 = ~w359 & w360;
assign w362 = w359 & ~w360;
assign w363 = ~w361 & ~w362;
assign w364 = (~w316 & ~w318) | (~w316 & w16697) | (~w318 & w16697);
assign w365 = pi06 & pi08;
assign w366 = pi01 & pi13;
assign w367 = ~w365 & ~w366;
assign w368 = w365 & w366;
assign w369 = ~w367 & ~w368;
assign w370 = ~w319 & ~w323;
assign w371 = ~w322 & ~w370;
assign w372 = w369 & w371;
assign w373 = ~w369 & ~w371;
assign w374 = ~w372 & ~w373;
assign w375 = ~w305 & ~w309;
assign w376 = ~w308 & ~w375;
assign w377 = w374 & w376;
assign w378 = ~w374 & ~w376;
assign w379 = ~w377 & ~w378;
assign w380 = ~w364 & w379;
assign w381 = w364 & ~w379;
assign w382 = ~w380 & ~w381;
assign w383 = w363 & w382;
assign w384 = ~w363 & ~w382;
assign w385 = ~w383 & ~w384;
assign w386 = ~w340 & w385;
assign w387 = w340 & ~w385;
assign w388 = ~w386 & ~w387;
assign w389 = w339 & w388;
assign w390 = ~w339 & ~w388;
assign w391 = ~w389 & ~w390;
assign w392 = ~w332 & ~w386;
assign w393 = (~w387 & w338) | (~w387 & w16492) | (w338 & w16492);
assign w394 = ~w380 & ~w383;
assign w395 = (~w372 & ~w374) | (~w372 & w16698) | (~w374 & w16698);
assign w396 = pi04 & pi11;
assign w397 = ~w368 & ~w396;
assign w398 = w368 & w396;
assign w399 = ~w397 & ~w398;
assign w400 = pi01 & pi14;
assign w401 = pi08 & w400;
assign w402 = ~pi08 & ~w400;
assign w403 = ~w401 & ~w402;
assign w404 = ~w399 & w403;
assign w405 = w399 & ~w403;
assign w406 = ~w404 & ~w405;
assign w407 = pi02 & pi13;
assign w408 = pi06 & pi09;
assign w409 = pi07 & pi08;
assign w410 = ~w408 & ~w409;
assign w411 = w408 & w409;
assign w412 = ~w410 & ~w411;
assign w413 = w407 & ~w412;
assign w414 = ~w407 & w412;
assign w415 = ~w413 & ~w414;
assign w416 = ~w406 & ~w415;
assign w417 = w406 & w415;
assign w418 = ~w416 & ~w417;
assign w419 = w395 & ~w418;
assign w420 = ~w395 & w418;
assign w421 = ~w419 & ~w420;
assign w422 = ~w349 & ~w352;
assign w423 = ~w351 & ~w422;
assign w424 = ~w287 & ~w344;
assign w425 = ~w343 & ~w424;
assign w426 = w423 & w425;
assign w427 = ~w423 & ~w425;
assign w428 = ~w426 & ~w427;
assign w429 = pi05 & pi10;
assign w430 = pi03 & pi12;
assign w431 = pi00 & pi15;
assign w432 = ~w430 & ~w431;
assign w433 = w430 & w431;
assign w434 = ~w432 & ~w433;
assign w435 = w429 & ~w434;
assign w436 = ~w429 & w434;
assign w437 = ~w435 & ~w436;
assign w438 = ~w428 & w437;
assign w439 = w428 & ~w437;
assign w440 = ~w438 & ~w439;
assign w441 = (~w357 & ~w359) | (~w357 & w16808) | (~w359 & w16808);
assign w442 = w440 & ~w441;
assign w443 = ~w440 & w441;
assign w444 = ~w442 & ~w443;
assign w445 = w421 & w444;
assign w446 = ~w421 & ~w444;
assign w447 = ~w445 & ~w446;
assign w448 = ~w394 & w447;
assign w449 = w394 & ~w447;
assign w450 = ~w448 & ~w449;
assign w451 = w393 & ~w450;
assign w452 = ~w393 & w450;
assign w453 = ~w451 & ~w452;
assign w454 = ~w442 & ~w445;
assign w455 = ~w429 & ~w433;
assign w456 = ~w432 & ~w455;
assign w457 = ~w398 & ~w403;
assign w458 = ~w397 & ~w457;
assign w459 = w456 & w458;
assign w460 = ~w456 & ~w458;
assign w461 = ~w459 & ~w460;
assign w462 = pi05 & pi11;
assign w463 = pi00 & pi16;
assign w464 = pi06 & pi10;
assign w465 = ~w463 & ~w464;
assign w466 = w463 & w464;
assign w467 = ~w465 & ~w466;
assign w468 = w462 & ~w467;
assign w469 = ~w462 & w467;
assign w470 = ~w468 & ~w469;
assign w471 = ~w461 & w470;
assign w472 = w461 & ~w470;
assign w473 = ~w471 & ~w472;
assign w474 = (~w416 & ~w418) | (~w416 & w16699) | (~w418 & w16699);
assign w475 = w473 & ~w474;
assign w476 = ~w473 & w474;
assign w477 = ~w475 & ~w476;
assign w478 = pi07 & pi09;
assign w479 = pi01 & pi15;
assign w480 = ~w478 & ~w479;
assign w481 = w478 & w479;
assign w482 = ~w480 & ~w481;
assign w483 = w401 & w482;
assign w484 = ~w401 & ~w482;
assign w485 = ~w483 & ~w484;
assign w486 = ~w407 & ~w411;
assign w487 = ~w410 & ~w486;
assign w488 = w485 & w487;
assign w489 = ~w485 & ~w487;
assign w490 = ~w488 & ~w489;
assign w491 = (~w426 & ~w428) | (~w426 & w16700) | (~w428 & w16700);
assign w492 = pi04 & pi12;
assign w493 = pi03 & pi13;
assign w494 = pi02 & pi14;
assign w495 = ~w493 & ~w494;
assign w496 = w493 & w494;
assign w497 = ~w495 & ~w496;
assign w498 = w492 & ~w497;
assign w499 = ~w492 & w497;
assign w500 = ~w498 & ~w499;
assign w501 = ~w491 & ~w500;
assign w502 = w491 & w500;
assign w503 = ~w501 & ~w502;
assign w504 = w490 & w503;
assign w505 = ~w490 & ~w503;
assign w506 = ~w504 & ~w505;
assign w507 = ~w477 & ~w506;
assign w508 = w477 & w506;
assign w509 = ~w507 & ~w508;
assign w510 = ~w454 & w509;
assign w511 = w454 & ~w509;
assign w512 = ~w510 & ~w511;
assign w513 = ~w393 & ~w448;
assign w514 = ~w449 & ~w513;
assign w515 = w512 & w514;
assign w516 = ~w512 & ~w514;
assign w517 = ~w515 & ~w516;
assign w518 = ~w475 & ~w508;
assign w519 = pi01 & pi16;
assign w520 = ~pi09 & ~w519;
assign w521 = pi16 & w154;
assign w522 = ~w520 & ~w521;
assign w523 = ~w492 & ~w496;
assign w524 = ~w495 & ~w523;
assign w525 = w522 & w524;
assign w526 = ~w522 & ~w524;
assign w527 = ~w525 & ~w526;
assign w528 = ~w462 & ~w466;
assign w529 = ~w465 & ~w528;
assign w530 = w527 & w529;
assign w531 = ~w527 & ~w529;
assign w532 = ~w530 & ~w531;
assign w533 = ~w483 & ~w488;
assign w534 = (~w459 & ~w461) | (~w459 & w16701) | (~w461 & w16701);
assign w535 = ~w533 & ~w534;
assign w536 = w533 & w534;
assign w537 = ~w535 & ~w536;
assign w538 = ~w532 & ~w537;
assign w539 = w532 & w537;
assign w540 = ~w538 & ~w539;
assign w541 = (~w501 & ~w503) | (~w501 & w16809) | (~w503 & w16809);
assign w542 = pi05 & pi12;
assign w543 = pi00 & pi17;
assign w544 = ~w542 & ~w543;
assign w545 = w542 & w543;
assign w546 = ~w544 & ~w545;
assign w547 = w481 & ~w546;
assign w548 = ~w481 & w546;
assign w549 = ~w547 & ~w548;
assign w550 = pi03 & pi14;
assign w551 = pi07 & pi10;
assign w552 = pi08 & pi09;
assign w553 = ~w551 & ~w552;
assign w554 = w551 & w552;
assign w555 = ~w553 & ~w554;
assign w556 = w550 & ~w555;
assign w557 = ~w550 & w555;
assign w558 = ~w556 & ~w557;
assign w559 = ~w549 & ~w558;
assign w560 = w549 & w558;
assign w561 = ~w559 & ~w560;
assign w562 = pi06 & pi11;
assign w563 = pi04 & pi13;
assign w564 = pi02 & pi15;
assign w565 = ~w563 & ~w564;
assign w566 = w563 & w564;
assign w567 = ~w565 & ~w566;
assign w568 = w562 & ~w567;
assign w569 = ~w562 & w567;
assign w570 = ~w568 & ~w569;
assign w571 = w561 & ~w570;
assign w572 = ~w561 & w570;
assign w573 = ~w571 & ~w572;
assign w574 = ~w541 & w573;
assign w575 = w541 & ~w573;
assign w576 = ~w574 & ~w575;
assign w577 = w540 & w576;
assign w578 = ~w540 & ~w576;
assign w579 = ~w577 & ~w578;
assign w580 = ~w518 & w579;
assign w581 = w518 & ~w579;
assign w582 = ~w580 & ~w581;
assign w583 = ~w449 & ~w511;
assign w584 = (w338 & w16810) | (w338 & w16811) | (w16810 & w16811);
assign w585 = ~w510 & ~w584;
assign w586 = w582 & w585;
assign w587 = ~w582 & ~w585;
assign w588 = ~w586 & ~w587;
assign w589 = (~w510 & ~w579) | (~w510 & w16494) | (~w579 & w16494);
assign w590 = (~w581 & w584) | (~w581 & w16495) | (w584 & w16495);
assign w591 = ~w574 & ~w577;
assign w592 = ~w481 & ~w545;
assign w593 = ~w544 & ~w592;
assign w594 = ~w550 & ~w554;
assign w595 = ~w553 & ~w594;
assign w596 = ~w562 & ~w566;
assign w597 = ~w565 & ~w596;
assign w598 = w595 & w597;
assign w599 = ~w595 & ~w597;
assign w600 = ~w598 & ~w599;
assign w601 = ~w593 & ~w600;
assign w602 = w593 & w600;
assign w603 = ~w601 & ~w602;
assign w604 = (~w525 & ~w527) | (~w525 & w16812) | (~w527 & w16812);
assign w605 = (~w559 & ~w561) | (~w559 & w16702) | (~w561 & w16702);
assign w606 = ~w604 & ~w605;
assign w607 = w604 & w605;
assign w608 = ~w606 & ~w607;
assign w609 = w603 & w608;
assign w610 = ~w603 & ~w608;
assign w611 = ~w609 & ~w610;
assign w612 = (~w535 & ~w537) | (~w535 & w16813) | (~w537 & w16813);
assign w613 = pi07 & pi11;
assign w614 = pi00 & pi18;
assign w615 = pi05 & pi13;
assign w616 = ~w614 & ~w615;
assign w617 = w614 & w615;
assign w618 = ~w616 & ~w617;
assign w619 = w613 & ~w618;
assign w620 = ~w613 & w618;
assign w621 = ~w619 & ~w620;
assign w622 = pi04 & pi14;
assign w623 = pi03 & pi15;
assign w624 = pi02 & pi16;
assign w625 = ~w623 & ~w624;
assign w626 = w623 & w624;
assign w627 = ~w625 & ~w626;
assign w628 = w622 & ~w627;
assign w629 = ~w622 & w627;
assign w630 = ~w628 & ~w629;
assign w631 = ~w621 & ~w630;
assign w632 = w621 & w630;
assign w633 = ~w631 & ~w632;
assign w634 = pi06 & pi12;
assign w635 = ~w521 & ~w634;
assign w636 = w521 & w634;
assign w637 = ~w635 & ~w636;
assign w638 = pi08 & pi10;
assign w639 = pi01 & pi17;
assign w640 = ~w638 & ~w639;
assign w641 = w638 & w639;
assign w642 = ~w640 & ~w641;
assign w643 = ~w637 & w642;
assign w644 = w637 & ~w642;
assign w645 = ~w643 & ~w644;
assign w646 = w633 & ~w645;
assign w647 = ~w633 & w645;
assign w648 = ~w646 & ~w647;
assign w649 = ~w612 & w648;
assign w650 = w612 & ~w648;
assign w651 = ~w649 & ~w650;
assign w652 = w611 & w651;
assign w653 = ~w611 & ~w651;
assign w654 = ~w652 & ~w653;
assign w655 = w591 & ~w654;
assign w656 = ~w591 & w654;
assign w657 = ~w655 & ~w656;
assign w658 = w590 & ~w657;
assign w659 = ~w590 & w657;
assign w660 = ~w658 & ~w659;
assign w661 = (~w584 & w16703) | (~w584 & w16704) | (w16703 & w16704);
assign w662 = ~w655 & ~w661;
assign w663 = ~w613 & ~w617;
assign w664 = ~w616 & ~w663;
assign w665 = ~w636 & ~w642;
assign w666 = ~w635 & ~w665;
assign w667 = w664 & w666;
assign w668 = ~w664 & ~w666;
assign w669 = ~w667 & ~w668;
assign w670 = pi03 & pi16;
assign w671 = pi09 & pi10;
assign w672 = pi08 & pi11;
assign w673 = ~w671 & ~w672;
assign w674 = w671 & w672;
assign w675 = ~w673 & ~w674;
assign w676 = w670 & ~w675;
assign w677 = ~w670 & w675;
assign w678 = ~w676 & ~w677;
assign w679 = ~w669 & w678;
assign w680 = w669 & ~w678;
assign w681 = ~w679 & ~w680;
assign w682 = (~w631 & ~w633) | (~w631 & w16705) | (~w633 & w16705);
assign w683 = ~pi18 & w641;
assign w684 = pi01 & pi18;
assign w685 = ~pi10 & ~w684;
assign w686 = pi10 & w684;
assign w687 = ~w685 & ~w686;
assign w688 = ~w641 & ~w687;
assign w689 = ~w683 & ~w688;
assign w690 = ~w622 & ~w626;
assign w691 = ~w625 & ~w690;
assign w692 = w689 & w691;
assign w693 = ~w689 & ~w691;
assign w694 = ~w692 & ~w693;
assign w695 = ~w682 & w694;
assign w696 = w682 & ~w694;
assign w697 = ~w695 & ~w696;
assign w698 = w681 & w697;
assign w699 = ~w681 & ~w697;
assign w700 = ~w698 & ~w699;
assign w701 = (~w598 & ~w600) | (~w598 & w16814) | (~w600 & w16814);
assign w702 = pi00 & pi19;
assign w703 = pi04 & pi15;
assign w704 = pi02 & pi17;
assign w705 = ~w703 & ~w704;
assign w706 = w703 & w704;
assign w707 = ~w705 & ~w706;
assign w708 = w702 & ~w707;
assign w709 = ~w702 & w707;
assign w710 = ~w708 & ~w709;
assign w711 = pi05 & pi14;
assign w712 = pi06 & pi13;
assign w713 = pi07 & pi12;
assign w714 = ~w712 & ~w713;
assign w715 = w712 & w713;
assign w716 = ~w714 & ~w715;
assign w717 = w711 & ~w716;
assign w718 = ~w711 & w716;
assign w719 = ~w717 & ~w718;
assign w720 = ~w710 & ~w719;
assign w721 = w710 & w719;
assign w722 = ~w720 & ~w721;
assign w723 = w701 & ~w722;
assign w724 = ~w701 & w722;
assign w725 = ~w723 & ~w724;
assign w726 = (~w606 & ~w608) | (~w606 & w16815) | (~w608 & w16815);
assign w727 = ~w725 & w726;
assign w728 = w725 & ~w726;
assign w729 = ~w727 & ~w728;
assign w730 = w700 & w729;
assign w731 = ~w700 & ~w729;
assign w732 = ~w730 & ~w731;
assign w733 = (~w649 & ~w651) | (~w649 & w17025) | (~w651 & w17025);
assign w734 = ~w732 & w733;
assign w735 = w732 & ~w733;
assign w736 = ~w734 & ~w735;
assign w737 = w662 & w736;
assign w738 = ~w662 & ~w736;
assign w739 = ~w737 & ~w738;
assign w740 = ~w655 & ~w734;
assign w741 = ~w661 & w740;
assign w742 = ~w735 & ~w741;
assign w743 = (~w728 & ~w729) | (~w728 & w17026) | (~w729 & w17026);
assign w744 = (~w667 & ~w669) | (~w667 & w16816) | (~w669 & w16816);
assign w745 = (~w683 & ~w689) | (~w683 & w16817) | (~w689 & w16817);
assign w746 = pi02 & pi18;
assign w747 = pi03 & pi17;
assign w748 = pi04 & pi16;
assign w749 = ~w747 & ~w748;
assign w750 = w747 & w748;
assign w751 = ~w749 & ~w750;
assign w752 = w746 & ~w751;
assign w753 = ~w746 & w751;
assign w754 = ~w752 & ~w753;
assign w755 = ~w745 & ~w754;
assign w756 = w745 & w754;
assign w757 = ~w755 & ~w756;
assign w758 = w744 & ~w757;
assign w759 = ~w744 & w757;
assign w760 = ~w758 & ~w759;
assign w761 = (~w695 & ~w697) | (~w695 & w16818) | (~w697 & w16818);
assign w762 = ~w760 & w761;
assign w763 = w760 & ~w761;
assign w764 = ~w762 & ~w763;
assign w765 = ~w711 & ~w715;
assign w766 = ~w714 & ~w765;
assign w767 = pi07 & pi13;
assign w768 = pi00 & pi20;
assign w769 = ~w767 & ~w768;
assign w770 = w767 & w768;
assign w771 = ~w769 & ~w770;
assign w772 = w686 & ~w771;
assign w773 = ~w686 & w771;
assign w774 = ~w772 & ~w773;
assign w775 = w766 & ~w774;
assign w776 = ~w766 & w774;
assign w777 = ~w775 & ~w776;
assign w778 = pi08 & pi12;
assign w779 = pi05 & pi15;
assign w780 = pi06 & pi14;
assign w781 = ~w779 & ~w780;
assign w782 = w779 & w780;
assign w783 = ~w781 & ~w782;
assign w784 = w778 & ~w783;
assign w785 = ~w778 & w783;
assign w786 = ~w784 & ~w785;
assign w787 = ~w777 & w786;
assign w788 = w777 & ~w786;
assign w789 = ~w787 & ~w788;
assign w790 = ~w720 & ~w724;
assign w791 = pi09 & pi11;
assign w792 = pi01 & pi19;
assign w793 = ~w791 & ~w792;
assign w794 = w791 & w792;
assign w795 = ~w793 & ~w794;
assign w796 = ~w670 & ~w674;
assign w797 = ~w673 & ~w796;
assign w798 = w795 & w797;
assign w799 = ~w795 & ~w797;
assign w800 = ~w798 & ~w799;
assign w801 = ~w702 & ~w706;
assign w802 = ~w705 & ~w801;
assign w803 = w800 & w802;
assign w804 = ~w800 & ~w802;
assign w805 = ~w803 & ~w804;
assign w806 = ~w790 & w805;
assign w807 = w790 & ~w805;
assign w808 = ~w806 & ~w807;
assign w809 = w789 & w808;
assign w810 = ~w789 & ~w808;
assign w811 = ~w809 & ~w810;
assign w812 = w764 & w811;
assign w813 = ~w764 & ~w811;
assign w814 = ~w812 & ~w813;
assign w815 = ~w743 & w814;
assign w816 = w743 & ~w814;
assign w817 = ~w815 & ~w816;
assign w818 = w742 & w817;
assign w819 = ~w742 & ~w817;
assign w820 = ~w818 & ~w819;
assign w821 = ~w763 & ~w812;
assign w822 = ~w746 & ~w750;
assign w823 = ~w749 & ~w822;
assign w824 = ~w778 & ~w782;
assign w825 = ~w781 & ~w824;
assign w826 = w823 & w825;
assign w827 = ~w823 & ~w825;
assign w828 = ~w826 & ~w827;
assign w829 = ~w686 & ~w770;
assign w830 = ~w769 & ~w829;
assign w831 = ~w828 & ~w830;
assign w832 = w828 & w830;
assign w833 = ~w831 & ~w832;
assign w834 = ~w759 & w17027;
assign w835 = (w833 & w759) | (w833 & w17028) | (w759 & w17028);
assign w836 = ~w834 & ~w835;
assign w837 = pi06 & pi15;
assign w838 = pi08 & pi13;
assign w839 = pi07 & pi14;
assign w840 = ~w838 & ~w839;
assign w841 = w838 & w839;
assign w842 = ~w840 & ~w841;
assign w843 = w837 & ~w842;
assign w844 = ~w837 & w842;
assign w845 = ~w843 & ~w844;
assign w846 = pi05 & pi16;
assign w847 = pi02 & pi19;
assign w848 = pi03 & pi18;
assign w849 = ~w847 & ~w848;
assign w850 = w847 & w848;
assign w851 = ~w849 & ~w850;
assign w852 = w846 & ~w851;
assign w853 = ~w846 & w851;
assign w854 = ~w852 & ~w853;
assign w855 = ~w845 & ~w854;
assign w856 = w845 & w854;
assign w857 = ~w855 & ~w856;
assign w858 = pi04 & pi17;
assign w859 = pi10 & pi11;
assign w860 = pi09 & pi12;
assign w861 = ~w859 & ~w860;
assign w862 = w859 & w860;
assign w863 = ~w861 & ~w862;
assign w864 = w858 & ~w863;
assign w865 = ~w858 & w863;
assign w866 = ~w864 & ~w865;
assign w867 = w857 & ~w866;
assign w868 = ~w857 & w866;
assign w869 = ~w867 & ~w868;
assign w870 = ~w836 & ~w869;
assign w871 = w836 & w869;
assign w872 = ~w870 & ~w871;
assign w873 = (~w798 & ~w800) | (~w798 & w16706) | (~w800 & w16706);
assign w874 = pi00 & pi21;
assign w875 = w794 & w874;
assign w876 = ~w794 & ~w874;
assign w877 = ~w875 & ~w876;
assign w878 = pi01 & pi20;
assign w879 = pi11 & w878;
assign w880 = ~pi11 & ~w878;
assign w881 = ~w879 & ~w880;
assign w882 = w877 & w881;
assign w883 = ~w877 & ~w881;
assign w884 = ~w882 & ~w883;
assign w885 = ~w873 & w884;
assign w886 = w873 & ~w884;
assign w887 = ~w885 & ~w886;
assign w888 = (~w775 & ~w777) | (~w775 & w16819) | (~w777 & w16819);
assign w889 = ~w887 & w888;
assign w890 = w887 & ~w888;
assign w891 = ~w889 & ~w890;
assign w892 = (~w806 & ~w808) | (~w806 & w17029) | (~w808 & w17029);
assign w893 = ~w891 & w892;
assign w894 = w891 & ~w892;
assign w895 = ~w893 & ~w894;
assign w896 = w872 & w895;
assign w897 = ~w872 & ~w895;
assign w898 = ~w896 & ~w897;
assign w899 = ~w821 & w898;
assign w900 = w821 & ~w898;
assign w901 = ~w899 & ~w900;
assign w902 = ~w735 & ~w815;
assign w903 = (w902 & w661) | (w902 & w16496) | (w661 & w16496);
assign w904 = ~w816 & ~w903;
assign w905 = w901 & w904;
assign w906 = ~w901 & ~w904;
assign w907 = ~w905 & ~w906;
assign w908 = ~w894 & ~w896;
assign w909 = (~w875 & ~w877) | (~w875 & w17030) | (~w877 & w17030);
assign w910 = ~w837 & ~w841;
assign w911 = ~w840 & ~w910;
assign w912 = ~w846 & ~w850;
assign w913 = ~w849 & ~w912;
assign w914 = w911 & w913;
assign w915 = ~w911 & ~w913;
assign w916 = ~w914 & ~w915;
assign w917 = w909 & ~w916;
assign w918 = ~w909 & w916;
assign w919 = ~w917 & ~w918;
assign w920 = (~w885 & ~w887) | (~w885 & w16820) | (~w887 & w16820);
assign w921 = ~w919 & w920;
assign w922 = w919 & ~w920;
assign w923 = ~w921 & ~w922;
assign w924 = pi09 & pi13;
assign w925 = pi06 & pi16;
assign w926 = pi02 & pi20;
assign w927 = ~w925 & ~w926;
assign w928 = w925 & w926;
assign w929 = ~w927 & ~w928;
assign w930 = w924 & ~w929;
assign w931 = ~w924 & w929;
assign w932 = ~w930 & ~w931;
assign w933 = pi00 & pi22;
assign w934 = pi07 & pi15;
assign w935 = pi08 & pi14;
assign w936 = ~w934 & ~w935;
assign w937 = w934 & w935;
assign w938 = ~w936 & ~w937;
assign w939 = w933 & ~w938;
assign w940 = ~w933 & w938;
assign w941 = ~w939 & ~w940;
assign w942 = ~w932 & ~w941;
assign w943 = w932 & w941;
assign w944 = ~w942 & ~w943;
assign w945 = pi03 & pi19;
assign w946 = pi05 & pi17;
assign w947 = pi04 & pi18;
assign w948 = ~w946 & ~w947;
assign w949 = w946 & w947;
assign w950 = ~w948 & ~w949;
assign w951 = w945 & ~w950;
assign w952 = ~w945 & w950;
assign w953 = ~w951 & ~w952;
assign w954 = w944 & ~w953;
assign w955 = ~w944 & w953;
assign w956 = ~w954 & ~w955;
assign w957 = ~w923 & ~w956;
assign w958 = w923 & w956;
assign w959 = ~w957 & ~w958;
assign w960 = ~w835 & ~w871;
assign w961 = (~w855 & ~w857) | (~w855 & w17282) | (~w857 & w17282);
assign w962 = (~w826 & ~w828) | (~w826 & w17031) | (~w828 & w17031);
assign w963 = pi10 & pi12;
assign w964 = pi01 & pi21;
assign w965 = ~w963 & ~w964;
assign w966 = w963 & w964;
assign w967 = ~w965 & ~w966;
assign w968 = w879 & w967;
assign w969 = ~w879 & ~w967;
assign w970 = ~w968 & ~w969;
assign w971 = ~w858 & ~w862;
assign w972 = ~w861 & ~w971;
assign w973 = w970 & w972;
assign w974 = ~w970 & ~w972;
assign w975 = ~w973 & ~w974;
assign w976 = ~w962 & w975;
assign w977 = w962 & ~w975;
assign w978 = ~w976 & ~w977;
assign w979 = ~w961 & w978;
assign w980 = w961 & ~w978;
assign w981 = ~w979 & ~w980;
assign w982 = ~w960 & w981;
assign w983 = w960 & ~w981;
assign w984 = ~w982 & ~w983;
assign w985 = w959 & w984;
assign w986 = ~w959 & ~w984;
assign w987 = ~w985 & ~w986;
assign w988 = ~w908 & w987;
assign w989 = w908 & ~w987;
assign w990 = ~w988 & ~w989;
assign w991 = (w661 & w16821) | (w661 & w16822) | (w16821 & w16822);
assign w992 = ~w900 & ~w991;
assign w993 = w990 & w992;
assign w994 = ~w990 & ~w992;
assign w995 = ~w993 & ~w994;
assign w996 = ~w982 & ~w985;
assign w997 = (~w976 & ~w978) | (~w976 & w17283) | (~w978 & w17283);
assign w998 = (~w968 & ~w970) | (~w968 & w16707) | (~w970 & w16707);
assign w999 = pi04 & pi19;
assign w1000 = pi11 & pi12;
assign w1001 = pi10 & pi13;
assign w1002 = ~w1000 & ~w1001;
assign w1003 = w1000 & w1001;
assign w1004 = ~w1002 & ~w1003;
assign w1005 = w999 & ~w1004;
assign w1006 = ~w999 & w1004;
assign w1007 = ~w1005 & ~w1006;
assign w1008 = pi06 & pi17;
assign w1009 = pi05 & pi18;
assign w1010 = pi03 & pi20;
assign w1011 = ~w1009 & ~w1010;
assign w1012 = w1009 & w1010;
assign w1013 = ~w1011 & ~w1012;
assign w1014 = w1008 & ~w1013;
assign w1015 = ~w1008 & w1013;
assign w1016 = ~w1014 & ~w1015;
assign w1017 = ~w1007 & ~w1016;
assign w1018 = w1007 & w1016;
assign w1019 = ~w1017 & ~w1018;
assign w1020 = w998 & ~w1019;
assign w1021 = ~w998 & w1019;
assign w1022 = ~w1020 & ~w1021;
assign w1023 = ~w933 & ~w937;
assign w1024 = ~w936 & ~w1023;
assign w1025 = pi00 & pi23;
assign w1026 = pi02 & pi21;
assign w1027 = ~w1025 & ~w1026;
assign w1028 = pi02 & pi23;
assign w1029 = w874 & w1028;
assign w1030 = ~w1027 & ~w1029;
assign w1031 = w966 & ~w1030;
assign w1032 = ~w966 & w1030;
assign w1033 = ~w1031 & ~w1032;
assign w1034 = w1024 & ~w1033;
assign w1035 = ~w1024 & w1033;
assign w1036 = ~w1034 & ~w1035;
assign w1037 = pi07 & pi16;
assign w1038 = pi08 & pi15;
assign w1039 = pi09 & pi14;
assign w1040 = ~w1038 & ~w1039;
assign w1041 = w1038 & w1039;
assign w1042 = ~w1040 & ~w1041;
assign w1043 = w1037 & ~w1042;
assign w1044 = ~w1037 & w1042;
assign w1045 = ~w1043 & ~w1044;
assign w1046 = w1036 & ~w1045;
assign w1047 = ~w1036 & w1045;
assign w1048 = ~w1046 & ~w1047;
assign w1049 = w1022 & w1048;
assign w1050 = ~w1022 & ~w1048;
assign w1051 = ~w1049 & ~w1050;
assign w1052 = ~w997 & w1051;
assign w1053 = w997 & ~w1051;
assign w1054 = ~w1052 & ~w1053;
assign w1055 = (~w922 & ~w923) | (~w922 & w17032) | (~w923 & w17032);
assign w1056 = pi01 & pi22;
assign w1057 = pi12 & w1056;
assign w1058 = ~pi12 & ~w1056;
assign w1059 = ~w1057 & ~w1058;
assign w1060 = ~w945 & ~w949;
assign w1061 = ~w948 & ~w1060;
assign w1062 = w1059 & w1061;
assign w1063 = ~w1059 & ~w1061;
assign w1064 = ~w1062 & ~w1063;
assign w1065 = ~w924 & ~w928;
assign w1066 = ~w927 & ~w1065;
assign w1067 = w1064 & w1066;
assign w1068 = ~w1064 & ~w1066;
assign w1069 = ~w1067 & ~w1068;
assign w1070 = (~w914 & ~w916) | (~w914 & w17033) | (~w916 & w17033);
assign w1071 = (~w942 & ~w944) | (~w942 & w16823) | (~w944 & w16823);
assign w1072 = ~w1070 & ~w1071;
assign w1073 = w1070 & w1071;
assign w1074 = ~w1072 & ~w1073;
assign w1075 = w1069 & w1074;
assign w1076 = ~w1069 & ~w1074;
assign w1077 = ~w1075 & ~w1076;
assign w1078 = ~w1055 & w1077;
assign w1079 = w1055 & ~w1077;
assign w1080 = ~w1078 & ~w1079;
assign w1081 = w1054 & w1080;
assign w1082 = ~w1054 & ~w1080;
assign w1083 = ~w1081 & ~w1082;
assign w1084 = w996 & ~w1083;
assign w1085 = ~w996 & w1083;
assign w1086 = ~w1084 & ~w1085;
assign w1087 = ~w900 & ~w989;
assign w1088 = ~w991 & w1087;
assign w1089 = ~w988 & ~w1088;
assign w1090 = w1086 & w1089;
assign w1091 = ~w1086 & ~w1089;
assign w1092 = ~w1090 & ~w1091;
assign w1093 = ~w988 & ~w1085;
assign w1094 = (~w1084 & w1088) | (~w1084 & w16498) | (w1088 & w16498);
assign w1095 = (~w1078 & ~w1080) | (~w1078 & w17284) | (~w1080 & w17284);
assign w1096 = (~w1049 & ~w1051) | (~w1049 & w17285) | (~w1051 & w17285);
assign w1097 = ~w1008 & ~w1012;
assign w1098 = ~w1011 & ~w1097;
assign w1099 = ~w999 & ~w1003;
assign w1100 = ~w1002 & ~w1099;
assign w1101 = w1098 & w1100;
assign w1102 = ~w1098 & ~w1100;
assign w1103 = ~w1101 & ~w1102;
assign w1104 = ~w1037 & ~w1041;
assign w1105 = ~w1040 & ~w1104;
assign w1106 = ~w1103 & ~w1105;
assign w1107 = w1103 & w1105;
assign w1108 = ~w1106 & ~w1107;
assign w1109 = (~w1017 & ~w1019) | (~w1017 & w16708) | (~w1019 & w16708);
assign w1110 = (~w1034 & ~w1036) | (~w1034 & w16709) | (~w1036 & w16709);
assign w1111 = ~w1109 & ~w1110;
assign w1112 = w1109 & w1110;
assign w1113 = ~w1111 & ~w1112;
assign w1114 = w1108 & w1113;
assign w1115 = ~w1108 & ~w1113;
assign w1116 = ~w1114 & ~w1115;
assign w1117 = ~w1096 & w1116;
assign w1118 = w1096 & ~w1116;
assign w1119 = ~w1117 & ~w1118;
assign w1120 = (~w1072 & ~w1074) | (~w1072 & w17034) | (~w1074 & w17034);
assign w1121 = (~w1062 & ~w1064) | (~w1062 & w17035) | (~w1064 & w17035);
assign w1122 = pi00 & pi24;
assign w1123 = w1057 & w1122;
assign w1124 = ~w1057 & ~w1122;
assign w1125 = ~w1123 & ~w1124;
assign w1126 = pi11 & pi13;
assign w1127 = pi01 & pi23;
assign w1128 = ~w1126 & ~w1127;
assign w1129 = pi11 & pi23;
assign w1130 = w366 & w1129;
assign w1131 = ~w1128 & ~w1130;
assign w1132 = w1125 & w1131;
assign w1133 = ~w1125 & ~w1131;
assign w1134 = ~w1132 & ~w1133;
assign w1135 = pi07 & pi17;
assign w1136 = pi02 & pi22;
assign w1137 = pi06 & pi18;
assign w1138 = ~w1136 & ~w1137;
assign w1139 = w1136 & w1137;
assign w1140 = ~w1138 & ~w1139;
assign w1141 = w1135 & ~w1140;
assign w1142 = ~w1135 & w1140;
assign w1143 = ~w1141 & ~w1142;
assign w1144 = w1134 & ~w1143;
assign w1145 = ~w1134 & w1143;
assign w1146 = ~w1144 & ~w1145;
assign w1147 = w1121 & ~w1146;
assign w1148 = ~w1121 & w1146;
assign w1149 = ~w1147 & ~w1148;
assign w1150 = w966 & ~w1027;
assign w1151 = ~w1029 & ~w1150;
assign w1152 = pi03 & pi21;
assign w1153 = pi05 & pi19;
assign w1154 = pi04 & pi20;
assign w1155 = ~w1153 & ~w1154;
assign w1156 = w1153 & w1154;
assign w1157 = ~w1155 & ~w1156;
assign w1158 = w1152 & ~w1157;
assign w1159 = ~w1152 & w1157;
assign w1160 = ~w1158 & ~w1159;
assign w1161 = ~w1151 & ~w1160;
assign w1162 = w1151 & w1160;
assign w1163 = ~w1161 & ~w1162;
assign w1164 = pi08 & pi16;
assign w1165 = pi09 & pi15;
assign w1166 = pi10 & pi14;
assign w1167 = ~w1165 & ~w1166;
assign w1168 = w1165 & w1166;
assign w1169 = ~w1167 & ~w1168;
assign w1170 = w1164 & ~w1169;
assign w1171 = ~w1164 & w1169;
assign w1172 = ~w1170 & ~w1171;
assign w1173 = w1163 & ~w1172;
assign w1174 = ~w1163 & w1172;
assign w1175 = ~w1173 & ~w1174;
assign w1176 = w1149 & w1175;
assign w1177 = ~w1149 & ~w1175;
assign w1178 = ~w1176 & ~w1177;
assign w1179 = ~w1120 & w1178;
assign w1180 = w1120 & ~w1178;
assign w1181 = ~w1179 & ~w1180;
assign w1182 = w1119 & w1181;
assign w1183 = ~w1119 & ~w1181;
assign w1184 = ~w1182 & ~w1183;
assign w1185 = ~w1095 & w1184;
assign w1186 = w1095 & ~w1184;
assign w1187 = ~w1185 & ~w1186;
assign w1188 = w1094 & ~w1187;
assign w1189 = ~w1094 & w1187;
assign w1190 = ~w1188 & ~w1189;
assign w1191 = ~w1117 & ~w1182;
assign w1192 = (~w1123 & ~w1125) | (~w1123 & w16710) | (~w1125 & w16710);
assign w1193 = ~w1164 & ~w1168;
assign w1194 = ~w1167 & ~w1193;
assign w1195 = ~w1135 & ~w1139;
assign w1196 = ~w1138 & ~w1195;
assign w1197 = w1194 & w1196;
assign w1198 = ~w1194 & ~w1196;
assign w1199 = ~w1197 & ~w1198;
assign w1200 = w1192 & ~w1199;
assign w1201 = ~w1192 & w1199;
assign w1202 = ~w1200 & ~w1201;
assign w1203 = (~w1161 & ~w1163) | (~w1161 & w16824) | (~w1163 & w16824);
assign w1204 = ~w1202 & w1203;
assign w1205 = w1202 & ~w1203;
assign w1206 = ~w1204 & ~w1205;
assign w1207 = (~w1144 & ~w1146) | (~w1144 & w17036) | (~w1146 & w17036);
assign w1208 = ~w1206 & w1207;
assign w1209 = w1206 & ~w1207;
assign w1210 = ~w1208 & ~w1209;
assign w1211 = (~w1176 & ~w1178) | (~w1176 & w17037) | (~w1178 & w17037);
assign w1212 = ~w1210 & w1211;
assign w1213 = w1210 & ~w1211;
assign w1214 = ~w1212 & ~w1213;
assign w1215 = pi01 & pi24;
assign w1216 = (w1215 & w1130) | (w1215 & w16825) | (w1130 & w16825);
assign w1217 = ~w1130 & w16826;
assign w1218 = ~w1216 & ~w1217;
assign w1219 = ~w1152 & ~w1156;
assign w1220 = ~w1155 & ~w1219;
assign w1221 = ~w1218 & w1220;
assign w1222 = w1218 & ~w1220;
assign w1223 = ~w1221 & ~w1222;
assign w1224 = (~w1101 & ~w1103) | (~w1101 & w17038) | (~w1103 & w17038);
assign w1225 = pi05 & pi20;
assign w1226 = pi12 & pi13;
assign w1227 = pi11 & pi14;
assign w1228 = ~w1226 & ~w1227;
assign w1229 = w1226 & w1227;
assign w1230 = ~w1228 & ~w1229;
assign w1231 = w1225 & ~w1230;
assign w1232 = ~w1225 & w1230;
assign w1233 = ~w1231 & ~w1232;
assign w1234 = ~w1224 & ~w1233;
assign w1235 = w1224 & w1233;
assign w1236 = ~w1234 & ~w1235;
assign w1237 = ~w1223 & ~w1236;
assign w1238 = w1223 & w1236;
assign w1239 = ~w1237 & ~w1238;
assign w1240 = (~w1111 & ~w1113) | (~w1111 & w16827) | (~w1113 & w16827);
assign w1241 = pi10 & pi15;
assign w1242 = pi00 & pi25;
assign w1243 = ~w1028 & ~w1242;
assign w1244 = pi02 & pi25;
assign w1245 = w1025 & w1244;
assign w1246 = ~w1243 & ~w1245;
assign w1247 = w1241 & ~w1246;
assign w1248 = ~w1241 & w1246;
assign w1249 = ~w1247 & ~w1248;
assign w1250 = pi07 & pi18;
assign w1251 = pi08 & pi17;
assign w1252 = pi09 & pi16;
assign w1253 = ~w1251 & ~w1252;
assign w1254 = w1251 & w1252;
assign w1255 = ~w1253 & ~w1254;
assign w1256 = w1250 & ~w1255;
assign w1257 = ~w1250 & w1255;
assign w1258 = ~w1256 & ~w1257;
assign w1259 = ~w1249 & ~w1258;
assign w1260 = w1249 & w1258;
assign w1261 = ~w1259 & ~w1260;
assign w1262 = pi06 & pi19;
assign w1263 = pi03 & pi22;
assign w1264 = pi04 & pi21;
assign w1265 = ~w1263 & ~w1264;
assign w1266 = w1263 & w1264;
assign w1267 = ~w1265 & ~w1266;
assign w1268 = w1262 & ~w1267;
assign w1269 = ~w1262 & w1267;
assign w1270 = ~w1268 & ~w1269;
assign w1271 = w1261 & ~w1270;
assign w1272 = ~w1261 & w1270;
assign w1273 = ~w1271 & ~w1272;
assign w1274 = ~w1240 & w1273;
assign w1275 = w1240 & ~w1273;
assign w1276 = ~w1274 & ~w1275;
assign w1277 = w1239 & w1276;
assign w1278 = ~w1239 & ~w1276;
assign w1279 = ~w1277 & ~w1278;
assign w1280 = w1214 & w1279;
assign w1281 = ~w1214 & ~w1279;
assign w1282 = ~w1280 & ~w1281;
assign w1283 = w1191 & ~w1282;
assign w1284 = ~w1191 & w1282;
assign w1285 = ~w1283 & ~w1284;
assign w1286 = ~w1094 & ~w1185;
assign w1287 = ~w1186 & ~w1286;
assign w1288 = w1285 & w1287;
assign w1289 = ~w1285 & ~w1287;
assign w1290 = ~w1288 & ~w1289;
assign w1291 = ~w1213 & ~w1280;
assign w1292 = (~w1274 & ~w1276) | (~w1274 & w17039) | (~w1276 & w17039);
assign w1293 = (~w1234 & ~w1236) | (~w1234 & w17286) | (~w1236 & w17286);
assign w1294 = (~w1259 & ~w1261) | (~w1259 & w17287) | (~w1261 & w17287);
assign w1295 = pi12 & pi14;
assign w1296 = pi01 & pi25;
assign w1297 = ~w1295 & ~w1296;
assign w1298 = w1295 & w1296;
assign w1299 = ~w1297 & ~w1298;
assign w1300 = ~w1225 & ~w1229;
assign w1301 = ~w1228 & ~w1300;
assign w1302 = w1299 & w1301;
assign w1303 = ~w1299 & ~w1301;
assign w1304 = ~w1302 & ~w1303;
assign w1305 = ~w1262 & ~w1266;
assign w1306 = ~w1265 & ~w1305;
assign w1307 = w1304 & w1306;
assign w1308 = ~w1304 & ~w1306;
assign w1309 = ~w1307 & ~w1308;
assign w1310 = ~w1294 & w1309;
assign w1311 = w1294 & ~w1309;
assign w1312 = ~w1310 & ~w1311;
assign w1313 = ~w1293 & w1312;
assign w1314 = w1293 & ~w1312;
assign w1315 = ~w1313 & ~w1314;
assign w1316 = ~w1292 & w1315;
assign w1317 = w1292 & ~w1315;
assign w1318 = ~w1316 & ~w1317;
assign w1319 = ~w1250 & ~w1254;
assign w1320 = ~w1253 & ~w1319;
assign w1321 = w1241 & ~w1243;
assign w1322 = ~w1245 & ~w1321;
assign w1323 = w1320 & ~w1322;
assign w1324 = ~w1320 & w1322;
assign w1325 = ~w1323 & ~w1324;
assign w1326 = pi13 & w1215;
assign w1327 = pi00 & pi26;
assign w1328 = pi08 & pi18;
assign w1329 = ~w1327 & ~w1328;
assign w1330 = w1327 & w1328;
assign w1331 = ~w1329 & ~w1330;
assign w1332 = w1326 & ~w1331;
assign w1333 = ~w1326 & w1331;
assign w1334 = ~w1332 & ~w1333;
assign w1335 = ~w1325 & w1334;
assign w1336 = w1325 & ~w1334;
assign w1337 = ~w1335 & ~w1336;
assign w1338 = (~w1197 & ~w1199) | (~w1197 & w16711) | (~w1199 & w16711);
assign w1339 = ~pi24 & w1130;
assign w1340 = ~w1221 & ~w1339;
assign w1341 = ~w1338 & ~w1340;
assign w1342 = w1338 & w1340;
assign w1343 = ~w1341 & ~w1342;
assign w1344 = w1337 & w1343;
assign w1345 = ~w1337 & ~w1343;
assign w1346 = ~w1344 & ~w1345;
assign w1347 = (~w1205 & ~w1206) | (~w1205 & w17040) | (~w1206 & w17040);
assign w1348 = pi02 & pi24;
assign w1349 = pi03 & pi23;
assign w1350 = pi07 & pi19;
assign w1351 = ~w1349 & ~w1350;
assign w1352 = w1349 & w1350;
assign w1353 = ~w1351 & ~w1352;
assign w1354 = w1348 & ~w1353;
assign w1355 = ~w1348 & w1353;
assign w1356 = ~w1354 & ~w1355;
assign w1357 = pi09 & pi17;
assign w1358 = pi10 & pi16;
assign w1359 = pi11 & pi15;
assign w1360 = ~w1358 & ~w1359;
assign w1361 = w1358 & w1359;
assign w1362 = ~w1360 & ~w1361;
assign w1363 = w1357 & ~w1362;
assign w1364 = ~w1357 & w1362;
assign w1365 = ~w1363 & ~w1364;
assign w1366 = ~w1356 & ~w1365;
assign w1367 = w1356 & w1365;
assign w1368 = ~w1366 & ~w1367;
assign w1369 = pi04 & pi22;
assign w1370 = pi06 & pi20;
assign w1371 = pi05 & pi21;
assign w1372 = ~w1370 & ~w1371;
assign w1373 = w1370 & w1371;
assign w1374 = ~w1372 & ~w1373;
assign w1375 = w1369 & ~w1374;
assign w1376 = ~w1369 & w1374;
assign w1377 = ~w1375 & ~w1376;
assign w1378 = w1368 & ~w1377;
assign w1379 = ~w1368 & w1377;
assign w1380 = ~w1378 & ~w1379;
assign w1381 = ~w1347 & w1380;
assign w1382 = w1347 & ~w1380;
assign w1383 = ~w1381 & ~w1382;
assign w1384 = w1346 & w1383;
assign w1385 = ~w1346 & ~w1383;
assign w1386 = ~w1384 & ~w1385;
assign w1387 = w1318 & w1386;
assign w1388 = ~w1318 & ~w1386;
assign w1389 = ~w1387 & ~w1388;
assign w1390 = ~w1291 & w1389;
assign w1391 = w1291 & ~w1389;
assign w1392 = ~w1390 & ~w1391;
assign w1393 = ~w1186 & ~w1283;
assign w1394 = (w1393 & w1094) | (w1393 & w16499) | (w1094 & w16499);
assign w1395 = ~w1284 & ~w1394;
assign w1396 = w1392 & w1395;
assign w1397 = ~w1392 & ~w1395;
assign w1398 = ~w1396 & ~w1397;
assign w1399 = ~w1316 & ~w1387;
assign w1400 = (~w1381 & ~w1383) | (~w1381 & w17288) | (~w1383 & w17288);
assign w1401 = pi26 & w400;
assign w1402 = pi01 & pi26;
assign w1403 = ~pi14 & ~w1402;
assign w1404 = ~w1401 & ~w1403;
assign w1405 = pi00 & pi27;
assign w1406 = w1298 & w1405;
assign w1407 = ~w1298 & ~w1405;
assign w1408 = ~w1406 & ~w1407;
assign w1409 = w1404 & w1408;
assign w1410 = ~w1404 & ~w1408;
assign w1411 = ~w1409 & ~w1410;
assign w1412 = pi03 & pi24;
assign w1413 = pi06 & pi21;
assign w1414 = pi04 & pi23;
assign w1415 = ~w1413 & ~w1414;
assign w1416 = w1413 & w1414;
assign w1417 = ~w1415 & ~w1416;
assign w1418 = w1412 & ~w1417;
assign w1419 = ~w1412 & w1417;
assign w1420 = ~w1418 & ~w1419;
assign w1421 = pi05 & pi22;
assign w1422 = pi12 & pi15;
assign w1423 = pi13 & pi14;
assign w1424 = ~w1422 & ~w1423;
assign w1425 = w1422 & w1423;
assign w1426 = ~w1424 & ~w1425;
assign w1427 = w1421 & ~w1426;
assign w1428 = ~w1421 & w1426;
assign w1429 = ~w1427 & ~w1428;
assign w1430 = ~w1420 & ~w1429;
assign w1431 = w1420 & w1429;
assign w1432 = ~w1430 & ~w1431;
assign w1433 = w1411 & w1432;
assign w1434 = ~w1411 & ~w1432;
assign w1435 = ~w1433 & ~w1434;
assign w1436 = ~w1369 & ~w1373;
assign w1437 = ~w1372 & ~w1436;
assign w1438 = ~w1357 & ~w1361;
assign w1439 = ~w1360 & ~w1438;
assign w1440 = w1437 & w1439;
assign w1441 = ~w1437 & ~w1439;
assign w1442 = ~w1440 & ~w1441;
assign w1443 = ~w1348 & ~w1352;
assign w1444 = ~w1351 & ~w1443;
assign w1445 = ~w1442 & ~w1444;
assign w1446 = w1442 & w1444;
assign w1447 = ~w1445 & ~w1446;
assign w1448 = (~w1341 & ~w1343) | (~w1341 & w16828) | (~w1343 & w16828);
assign w1449 = ~w1447 & w1448;
assign w1450 = w1447 & ~w1448;
assign w1451 = ~w1449 & ~w1450;
assign w1452 = w1435 & w1451;
assign w1453 = ~w1435 & ~w1451;
assign w1454 = ~w1452 & ~w1453;
assign w1455 = ~w1400 & w1454;
assign w1456 = w1400 & ~w1454;
assign w1457 = ~w1455 & ~w1456;
assign w1458 = (~w1366 & ~w1368) | (~w1366 & w16829) | (~w1368 & w16829);
assign w1459 = (~w1302 & ~w1304) | (~w1302 & w16712) | (~w1304 & w16712);
assign w1460 = (~w1323 & ~w1325) | (~w1323 & w16713) | (~w1325 & w16713);
assign w1461 = ~w1459 & ~w1460;
assign w1462 = w1459 & w1460;
assign w1463 = ~w1461 & ~w1462;
assign w1464 = w1458 & ~w1463;
assign w1465 = ~w1458 & w1463;
assign w1466 = ~w1464 & ~w1465;
assign w1467 = ~w1326 & ~w1330;
assign w1468 = ~w1329 & ~w1467;
assign w1469 = pi11 & pi16;
assign w1470 = pi07 & pi20;
assign w1471 = ~w1244 & ~w1470;
assign w1472 = w1244 & w1470;
assign w1473 = ~w1471 & ~w1472;
assign w1474 = w1469 & ~w1473;
assign w1475 = ~w1469 & w1473;
assign w1476 = ~w1474 & ~w1475;
assign w1477 = w1468 & ~w1476;
assign w1478 = ~w1468 & w1476;
assign w1479 = ~w1477 & ~w1478;
assign w1480 = pi08 & pi19;
assign w1481 = pi10 & pi17;
assign w1482 = pi09 & pi18;
assign w1483 = ~w1481 & ~w1482;
assign w1484 = w1481 & w1482;
assign w1485 = ~w1483 & ~w1484;
assign w1486 = w1480 & ~w1485;
assign w1487 = ~w1480 & w1485;
assign w1488 = ~w1486 & ~w1487;
assign w1489 = ~w1479 & w1488;
assign w1490 = w1479 & ~w1488;
assign w1491 = ~w1489 & ~w1490;
assign w1492 = ~w1310 & ~w1313;
assign w1493 = w1491 & ~w1492;
assign w1494 = ~w1491 & w1492;
assign w1495 = ~w1493 & ~w1494;
assign w1496 = w1466 & w1495;
assign w1497 = ~w1466 & ~w1495;
assign w1498 = ~w1496 & ~w1497;
assign w1499 = w1457 & w1498;
assign w1500 = ~w1457 & ~w1498;
assign w1501 = ~w1499 & ~w1500;
assign w1502 = ~w1399 & w1501;
assign w1503 = w1399 & ~w1501;
assign w1504 = ~w1502 & ~w1503;
assign w1505 = ~w1284 & ~w1390;
assign w1506 = (~w1094 & w16500) | (~w1094 & w16501) | (w16500 & w16501);
assign w1507 = ~w1391 & ~w1506;
assign w1508 = w1504 & w1507;
assign w1509 = ~w1504 & ~w1507;
assign w1510 = ~w1508 & ~w1509;
assign w1511 = (~w1406 & ~w1408) | (~w1406 & w16714) | (~w1408 & w16714);
assign w1512 = pi08 & pi20;
assign w1513 = pi03 & pi25;
assign w1514 = pi04 & pi24;
assign w1515 = ~w1513 & ~w1514;
assign w1516 = w1513 & w1514;
assign w1517 = ~w1515 & ~w1516;
assign w1518 = w1512 & ~w1517;
assign w1519 = ~w1512 & w1517;
assign w1520 = ~w1518 & ~w1519;
assign w1521 = ~w1511 & ~w1520;
assign w1522 = w1511 & w1520;
assign w1523 = ~w1521 & ~w1522;
assign w1524 = pi07 & pi21;
assign w1525 = pi06 & pi22;
assign w1526 = pi05 & pi23;
assign w1527 = ~w1525 & ~w1526;
assign w1528 = w1525 & w1526;
assign w1529 = ~w1527 & ~w1528;
assign w1530 = w1524 & ~w1529;
assign w1531 = ~w1524 & w1529;
assign w1532 = ~w1530 & ~w1531;
assign w1533 = w1523 & ~w1532;
assign w1534 = ~w1523 & w1532;
assign w1535 = ~w1533 & ~w1534;
assign w1536 = (w1451 & w17289) | (w1451 & w17290) | (w17289 & w17290);
assign w1537 = (~w1451 & w17291) | (~w1451 & w17292) | (w17291 & w17292);
assign w1538 = ~w1536 & ~w1537;
assign w1539 = ~w1430 & ~w1433;
assign w1540 = (~w1477 & ~w1479) | (~w1477 & w17293) | (~w1479 & w17293);
assign w1541 = pi13 & pi15;
assign w1542 = pi01 & pi27;
assign w1543 = ~w1541 & ~w1542;
assign w1544 = w1541 & w1542;
assign w1545 = ~w1543 & ~w1544;
assign w1546 = w1401 & w1545;
assign w1547 = ~w1401 & ~w1545;
assign w1548 = ~w1546 & ~w1547;
assign w1549 = ~w1421 & ~w1425;
assign w1550 = ~w1424 & ~w1549;
assign w1551 = w1548 & w1550;
assign w1552 = ~w1548 & ~w1550;
assign w1553 = ~w1551 & ~w1552;
assign w1554 = ~w1540 & w1553;
assign w1555 = w1540 & ~w1553;
assign w1556 = ~w1554 & ~w1555;
assign w1557 = ~w1539 & w1556;
assign w1558 = w1539 & ~w1556;
assign w1559 = ~w1557 & ~w1558;
assign w1560 = w1538 & w1559;
assign w1561 = ~w1538 & ~w1559;
assign w1562 = ~w1560 & ~w1561;
assign w1563 = ~w1455 & ~w1499;
assign w1564 = ~w1493 & ~w1496;
assign w1565 = ~w1480 & ~w1484;
assign w1566 = ~w1483 & ~w1565;
assign w1567 = ~w1412 & ~w1416;
assign w1568 = ~w1415 & ~w1567;
assign w1569 = w1566 & w1568;
assign w1570 = ~w1566 & ~w1568;
assign w1571 = ~w1569 & ~w1570;
assign w1572 = ~w1469 & ~w1472;
assign w1573 = ~w1471 & ~w1572;
assign w1574 = ~w1571 & ~w1573;
assign w1575 = w1571 & w1573;
assign w1576 = ~w1574 & ~w1575;
assign w1577 = (~w1461 & ~w1463) | (~w1461 & w16830) | (~w1463 & w16830);
assign w1578 = ~w1576 & w1577;
assign w1579 = w1576 & ~w1577;
assign w1580 = ~w1578 & ~w1579;
assign w1581 = (~w1440 & ~w1442) | (~w1440 & w16715) | (~w1442 & w16715);
assign w1582 = pi11 & pi17;
assign w1583 = pi00 & pi28;
assign w1584 = pi12 & pi16;
assign w1585 = ~w1583 & ~w1584;
assign w1586 = w1583 & w1584;
assign w1587 = ~w1585 & ~w1586;
assign w1588 = w1582 & ~w1587;
assign w1589 = ~w1582 & w1587;
assign w1590 = ~w1588 & ~w1589;
assign w1591 = pi02 & pi26;
assign w1592 = pi09 & pi19;
assign w1593 = pi10 & pi18;
assign w1594 = ~w1592 & ~w1593;
assign w1595 = w1592 & w1593;
assign w1596 = ~w1594 & ~w1595;
assign w1597 = w1591 & ~w1596;
assign w1598 = ~w1591 & w1596;
assign w1599 = ~w1597 & ~w1598;
assign w1600 = ~w1590 & ~w1599;
assign w1601 = w1590 & w1599;
assign w1602 = ~w1600 & ~w1601;
assign w1603 = w1581 & ~w1602;
assign w1604 = ~w1581 & w1602;
assign w1605 = ~w1603 & ~w1604;
assign w1606 = w1580 & w1605;
assign w1607 = ~w1580 & ~w1605;
assign w1608 = ~w1606 & ~w1607;
assign w1609 = ~w1564 & w1608;
assign w1610 = w1564 & ~w1608;
assign w1611 = ~w1609 & ~w1610;
assign w1612 = ~w1563 & w1611;
assign w1613 = w1563 & ~w1611;
assign w1614 = ~w1612 & ~w1613;
assign w1615 = ~w1562 & ~w1614;
assign w1616 = w1562 & w1614;
assign w1617 = ~w1615 & ~w1616;
assign w1618 = (~w1094 & w17042) | (~w1094 & w17043) | (w17042 & w17043);
assign w1619 = ~w1503 & ~w1618;
assign w1620 = w1617 & w1619;
assign w1621 = ~w1617 & ~w1619;
assign w1622 = ~w1620 & ~w1621;
assign w1623 = ~w1609 & ~w1612;
assign w1624 = ~w1591 & ~w1595;
assign w1625 = ~w1594 & ~w1624;
assign w1626 = ~w1582 & ~w1586;
assign w1627 = ~w1585 & ~w1626;
assign w1628 = w1625 & w1627;
assign w1629 = ~w1625 & ~w1627;
assign w1630 = ~w1628 & ~w1629;
assign w1631 = pi00 & pi29;
assign w1632 = pi02 & pi27;
assign w1633 = ~w1631 & ~w1632;
assign w1634 = pi02 & pi29;
assign w1635 = w1405 & w1634;
assign w1636 = ~w1633 & ~w1635;
assign w1637 = w1544 & ~w1636;
assign w1638 = ~w1544 & w1636;
assign w1639 = ~w1637 & ~w1638;
assign w1640 = ~w1630 & w1639;
assign w1641 = w1630 & ~w1639;
assign w1642 = ~w1640 & ~w1641;
assign w1643 = ~w1600 & ~w1604;
assign w1644 = (~w1521 & ~w1523) | (~w1521 & w16831) | (~w1523 & w16831);
assign w1645 = ~w1643 & ~w1644;
assign w1646 = w1643 & w1644;
assign w1647 = ~w1645 & ~w1646;
assign w1648 = w1642 & w1647;
assign w1649 = ~w1642 & ~w1647;
assign w1650 = ~w1648 & ~w1649;
assign w1651 = (~w1579 & ~w1580) | (~w1579 & w17044) | (~w1580 & w17044);
assign w1652 = ~w1554 & ~w1557;
assign w1653 = ~w1651 & ~w1652;
assign w1654 = w1651 & w1652;
assign w1655 = ~w1653 & ~w1654;
assign w1656 = w1650 & w1655;
assign w1657 = ~w1650 & ~w1655;
assign w1658 = ~w1656 & ~w1657;
assign w1659 = ~w1536 & ~w1560;
assign w1660 = (~w1569 & ~w1571) | (~w1569 & w17045) | (~w1571 & w17045);
assign w1661 = (~w1546 & ~w1548) | (~w1546 & w16832) | (~w1548 & w16832);
assign w1662 = pi06 & pi23;
assign w1663 = pi14 & pi15;
assign w1664 = pi13 & pi16;
assign w1665 = ~w1663 & ~w1664;
assign w1666 = w1663 & w1664;
assign w1667 = ~w1665 & ~w1666;
assign w1668 = w1662 & ~w1667;
assign w1669 = ~w1662 & w1667;
assign w1670 = ~w1668 & ~w1669;
assign w1671 = ~w1661 & ~w1670;
assign w1672 = w1661 & w1670;
assign w1673 = ~w1671 & ~w1672;
assign w1674 = w1660 & ~w1673;
assign w1675 = ~w1660 & w1673;
assign w1676 = ~w1674 & ~w1675;
assign w1677 = pi28 & w479;
assign w1678 = pi01 & pi28;
assign w1679 = ~pi15 & ~w1678;
assign w1680 = ~w1677 & ~w1679;
assign w1681 = ~w1524 & ~w1528;
assign w1682 = ~w1527 & ~w1681;
assign w1683 = w1680 & w1682;
assign w1684 = ~w1680 & ~w1682;
assign w1685 = ~w1683 & ~w1684;
assign w1686 = ~w1512 & ~w1516;
assign w1687 = ~w1515 & ~w1686;
assign w1688 = w1685 & w1687;
assign w1689 = ~w1685 & ~w1687;
assign w1690 = ~w1688 & ~w1689;
assign w1691 = pi12 & pi17;
assign w1692 = pi03 & pi26;
assign w1693 = pi08 & pi21;
assign w1694 = ~w1692 & ~w1693;
assign w1695 = w1692 & w1693;
assign w1696 = ~w1694 & ~w1695;
assign w1697 = w1691 & ~w1696;
assign w1698 = ~w1691 & w1696;
assign w1699 = ~w1697 & ~w1698;
assign w1700 = pi09 & pi20;
assign w1701 = pi10 & pi19;
assign w1702 = pi11 & pi18;
assign w1703 = ~w1701 & ~w1702;
assign w1704 = w1701 & w1702;
assign w1705 = ~w1703 & ~w1704;
assign w1706 = w1700 & ~w1705;
assign w1707 = ~w1700 & w1705;
assign w1708 = ~w1706 & ~w1707;
assign w1709 = ~w1699 & ~w1708;
assign w1710 = w1699 & w1708;
assign w1711 = ~w1709 & ~w1710;
assign w1712 = pi04 & pi25;
assign w1713 = pi07 & pi22;
assign w1714 = pi05 & pi24;
assign w1715 = ~w1713 & ~w1714;
assign w1716 = w1713 & w1714;
assign w1717 = ~w1715 & ~w1716;
assign w1718 = w1712 & ~w1717;
assign w1719 = ~w1712 & w1717;
assign w1720 = ~w1718 & ~w1719;
assign w1721 = w1711 & ~w1720;
assign w1722 = ~w1711 & w1720;
assign w1723 = ~w1721 & ~w1722;
assign w1724 = w1690 & w1723;
assign w1725 = ~w1690 & ~w1723;
assign w1726 = ~w1724 & ~w1725;
assign w1727 = w1676 & w1726;
assign w1728 = ~w1676 & ~w1726;
assign w1729 = ~w1727 & ~w1728;
assign w1730 = ~w1659 & w1729;
assign w1731 = w1659 & ~w1729;
assign w1732 = ~w1730 & ~w1731;
assign w1733 = w1658 & w1732;
assign w1734 = ~w1658 & ~w1732;
assign w1735 = ~w1733 & ~w1734;
assign w1736 = ~w1623 & w1735;
assign w1737 = w1623 & ~w1735;
assign w1738 = ~w1736 & ~w1737;
assign w1739 = ~w1503 & ~w1615;
assign w1740 = ~w1618 & w1739;
assign w1741 = ~w1616 & ~w1740;
assign w1742 = w1738 & w1741;
assign w1743 = ~w1738 & ~w1741;
assign w1744 = ~w1742 & ~w1743;
assign w1745 = ~w1730 & ~w1733;
assign w1746 = (~w1628 & ~w1630) | (~w1628 & w17046) | (~w1630 & w17046);
assign w1747 = (~w1683 & ~w1685) | (~w1683 & w16716) | (~w1685 & w16716);
assign w1748 = pi00 & pi30;
assign w1749 = w1677 & w1748;
assign w1750 = ~w1677 & ~w1748;
assign w1751 = ~w1749 & ~w1750;
assign w1752 = pi14 & pi16;
assign w1753 = pi01 & pi29;
assign w1754 = ~w1752 & ~w1753;
assign w1755 = pi14 & pi29;
assign w1756 = w519 & w1755;
assign w1757 = ~w1754 & ~w1756;
assign w1758 = w1751 & w1757;
assign w1759 = ~w1751 & ~w1757;
assign w1760 = ~w1758 & ~w1759;
assign w1761 = ~w1747 & w1760;
assign w1762 = w1747 & ~w1760;
assign w1763 = ~w1761 & ~w1762;
assign w1764 = w1746 & ~w1763;
assign w1765 = ~w1746 & w1763;
assign w1766 = ~w1764 & ~w1765;
assign w1767 = (~w1724 & ~w1726) | (~w1724 & w17294) | (~w1726 & w17294);
assign w1768 = ~w1766 & w1767;
assign w1769 = w1766 & ~w1767;
assign w1770 = ~w1768 & ~w1769;
assign w1771 = ~w1691 & ~w1695;
assign w1772 = ~w1694 & ~w1771;
assign w1773 = ~w1700 & ~w1704;
assign w1774 = ~w1703 & ~w1773;
assign w1775 = w1772 & w1774;
assign w1776 = ~w1772 & ~w1774;
assign w1777 = ~w1775 & ~w1776;
assign w1778 = w1544 & ~w1633;
assign w1779 = ~w1635 & ~w1778;
assign w1780 = ~w1777 & w1779;
assign w1781 = w1777 & ~w1779;
assign w1782 = ~w1780 & ~w1781;
assign w1783 = ~w1712 & ~w1716;
assign w1784 = ~w1715 & ~w1783;
assign w1785 = ~w1662 & ~w1666;
assign w1786 = ~w1665 & ~w1785;
assign w1787 = w1784 & w1786;
assign w1788 = ~w1784 & ~w1786;
assign w1789 = ~w1787 & ~w1788;
assign w1790 = pi13 & pi17;
assign w1791 = pi02 & pi28;
assign w1792 = pi09 & pi21;
assign w1793 = ~w1791 & ~w1792;
assign w1794 = w1791 & w1792;
assign w1795 = ~w1793 & ~w1794;
assign w1796 = w1790 & ~w1795;
assign w1797 = ~w1790 & w1795;
assign w1798 = ~w1796 & ~w1797;
assign w1799 = ~w1789 & w1798;
assign w1800 = w1789 & ~w1798;
assign w1801 = ~w1799 & ~w1800;
assign w1802 = (~w1709 & ~w1711) | (~w1709 & w16833) | (~w1711 & w16833);
assign w1803 = w1801 & ~w1802;
assign w1804 = ~w1801 & w1802;
assign w1805 = ~w1803 & ~w1804;
assign w1806 = w1782 & w1805;
assign w1807 = ~w1782 & ~w1805;
assign w1808 = ~w1806 & ~w1807;
assign w1809 = w1770 & w1808;
assign w1810 = ~w1770 & ~w1808;
assign w1811 = ~w1809 & ~w1810;
assign w1812 = (~w1653 & ~w1655) | (~w1653 & w17295) | (~w1655 & w17295);
assign w1813 = (~w1645 & ~w1647) | (~w1645 & w16834) | (~w1647 & w16834);
assign w1814 = (~w1671 & ~w1673) | (~w1671 & w17047) | (~w1673 & w17047);
assign w1815 = pi03 & pi27;
assign w1816 = pi04 & pi26;
assign w1817 = pi08 & pi22;
assign w1818 = ~w1816 & ~w1817;
assign w1819 = w1816 & w1817;
assign w1820 = ~w1818 & ~w1819;
assign w1821 = w1815 & ~w1820;
assign w1822 = ~w1815 & w1820;
assign w1823 = ~w1821 & ~w1822;
assign w1824 = pi05 & pi25;
assign w1825 = pi07 & pi23;
assign w1826 = pi06 & pi24;
assign w1827 = ~w1825 & ~w1826;
assign w1828 = w1825 & w1826;
assign w1829 = ~w1827 & ~w1828;
assign w1830 = w1824 & ~w1829;
assign w1831 = ~w1824 & w1829;
assign w1832 = ~w1830 & ~w1831;
assign w1833 = ~w1823 & ~w1832;
assign w1834 = w1823 & w1832;
assign w1835 = ~w1833 & ~w1834;
assign w1836 = pi10 & pi20;
assign w1837 = pi11 & pi19;
assign w1838 = pi12 & pi18;
assign w1839 = ~w1837 & ~w1838;
assign w1840 = w1837 & w1838;
assign w1841 = ~w1839 & ~w1840;
assign w1842 = w1836 & ~w1841;
assign w1843 = ~w1836 & w1841;
assign w1844 = ~w1842 & ~w1843;
assign w1845 = w1835 & ~w1844;
assign w1846 = ~w1835 & w1844;
assign w1847 = ~w1845 & ~w1846;
assign w1848 = ~w1814 & w1847;
assign w1849 = w1814 & ~w1847;
assign w1850 = ~w1848 & ~w1849;
assign w1851 = ~w1813 & w1850;
assign w1852 = w1813 & ~w1850;
assign w1853 = ~w1851 & ~w1852;
assign w1854 = ~w1812 & w1853;
assign w1855 = w1812 & ~w1853;
assign w1856 = ~w1854 & ~w1855;
assign w1857 = w1811 & w1856;
assign w1858 = ~w1811 & ~w1856;
assign w1859 = ~w1857 & ~w1858;
assign w1860 = ~w1745 & w1859;
assign w1861 = w1745 & ~w1859;
assign w1862 = ~w1860 & ~w1861;
assign w1863 = ~w1616 & ~w1736;
assign w1864 = (~w1737 & w1740) | (~w1737 & w16503) | (w1740 & w16503);
assign w1865 = w1862 & w1864;
assign w1866 = ~w1862 & ~w1864;
assign w1867 = ~w1865 & ~w1866;
assign w1868 = ~w1854 & ~w1857;
assign w1869 = ~w1769 & ~w1809;
assign w1870 = (~w1803 & ~w1805) | (~w1803 & w17048) | (~w1805 & w17048);
assign w1871 = (~w1749 & ~w1751) | (~w1749 & w16835) | (~w1751 & w16835);
assign w1872 = pi11 & pi20;
assign w1873 = pi12 & pi19;
assign w1874 = pi13 & pi18;
assign w1875 = ~w1873 & ~w1874;
assign w1876 = w1873 & w1874;
assign w1877 = ~w1875 & ~w1876;
assign w1878 = w1872 & ~w1877;
assign w1879 = ~w1872 & w1877;
assign w1880 = ~w1878 & ~w1879;
assign w1881 = ~w1871 & ~w1880;
assign w1882 = w1871 & w1880;
assign w1883 = ~w1881 & ~w1882;
assign w1884 = pi10 & pi21;
assign w1885 = pi00 & pi31;
assign w1886 = pi09 & pi22;
assign w1887 = ~w1885 & ~w1886;
assign w1888 = w1885 & w1886;
assign w1889 = ~w1887 & ~w1888;
assign w1890 = w1884 & ~w1889;
assign w1891 = ~w1884 & w1889;
assign w1892 = ~w1890 & ~w1891;
assign w1893 = w1883 & ~w1892;
assign w1894 = ~w1883 & w1892;
assign w1895 = ~w1893 & ~w1894;
assign w1896 = pi06 & pi25;
assign w1897 = pi15 & pi16;
assign w1898 = pi14 & pi17;
assign w1899 = ~w1897 & ~w1898;
assign w1900 = w1897 & w1898;
assign w1901 = ~w1899 & ~w1900;
assign w1902 = w1896 & ~w1901;
assign w1903 = ~w1896 & w1901;
assign w1904 = ~w1902 & ~w1903;
assign w1905 = pi08 & pi23;
assign w1906 = pi07 & pi24;
assign w1907 = pi05 & pi26;
assign w1908 = ~w1906 & ~w1907;
assign w1909 = w1906 & w1907;
assign w1910 = ~w1908 & ~w1909;
assign w1911 = w1905 & ~w1910;
assign w1912 = ~w1905 & w1910;
assign w1913 = ~w1911 & ~w1912;
assign w1914 = ~w1904 & ~w1913;
assign w1915 = w1904 & w1913;
assign w1916 = ~w1914 & ~w1915;
assign w1917 = pi04 & pi27;
assign w1918 = pi03 & pi28;
assign w1919 = ~w1917 & ~w1918;
assign w1920 = w1917 & w1918;
assign w1921 = ~w1919 & ~w1920;
assign w1922 = w1634 & ~w1921;
assign w1923 = ~w1634 & w1921;
assign w1924 = ~w1922 & ~w1923;
assign w1925 = w1916 & ~w1924;
assign w1926 = ~w1916 & w1924;
assign w1927 = ~w1925 & ~w1926;
assign w1928 = w1895 & w1927;
assign w1929 = ~w1895 & ~w1927;
assign w1930 = ~w1928 & ~w1929;
assign w1931 = ~w1870 & w1930;
assign w1932 = w1870 & ~w1930;
assign w1933 = ~w1931 & ~w1932;
assign w1934 = ~w1869 & w1933;
assign w1935 = w1869 & ~w1933;
assign w1936 = ~w1934 & ~w1935;
assign w1937 = (~w1848 & w1813) | (~w1848 & w17049) | (w1813 & w17049);
assign w1938 = pi16 & ~w1756;
assign w1939 = pi01 & pi30;
assign w1940 = ~w1938 & w1939;
assign w1941 = w1938 & ~w1939;
assign w1942 = ~w1940 & ~w1941;
assign w1943 = ~w1824 & ~w1828;
assign w1944 = ~w1827 & ~w1943;
assign w1945 = ~w1942 & w1944;
assign w1946 = w1942 & ~w1944;
assign w1947 = ~w1945 & ~w1946;
assign w1948 = ~w1787 & ~w1800;
assign w1949 = ~w1775 & ~w1781;
assign w1950 = ~w1948 & ~w1949;
assign w1951 = w1948 & w1949;
assign w1952 = ~w1950 & ~w1951;
assign w1953 = w1947 & w1952;
assign w1954 = ~w1947 & ~w1952;
assign w1955 = ~w1953 & ~w1954;
assign w1956 = ~w1937 & w1955;
assign w1957 = w1937 & ~w1955;
assign w1958 = ~w1956 & ~w1957;
assign w1959 = ~w1815 & ~w1819;
assign w1960 = ~w1818 & ~w1959;
assign w1961 = ~w1790 & ~w1794;
assign w1962 = ~w1793 & ~w1961;
assign w1963 = w1960 & w1962;
assign w1964 = ~w1960 & ~w1962;
assign w1965 = ~w1963 & ~w1964;
assign w1966 = ~w1836 & ~w1840;
assign w1967 = ~w1839 & ~w1966;
assign w1968 = ~w1965 & ~w1967;
assign w1969 = w1965 & w1967;
assign w1970 = ~w1968 & ~w1969;
assign w1971 = (~w1833 & ~w1835) | (~w1833 & w16836) | (~w1835 & w16836);
assign w1972 = ~w1970 & w1971;
assign w1973 = w1970 & ~w1971;
assign w1974 = ~w1972 & ~w1973;
assign w1975 = (~w1761 & ~w1763) | (~w1761 & w16837) | (~w1763 & w16837);
assign w1976 = ~w1974 & w1975;
assign w1977 = w1974 & ~w1975;
assign w1978 = ~w1976 & ~w1977;
assign w1979 = w1958 & w1978;
assign w1980 = ~w1958 & ~w1978;
assign w1981 = ~w1979 & ~w1980;
assign w1982 = w1936 & w1981;
assign w1983 = ~w1936 & ~w1981;
assign w1984 = ~w1982 & ~w1983;
assign w1985 = ~w1868 & w1984;
assign w1986 = w1868 & ~w1984;
assign w1987 = ~w1985 & ~w1986;
assign w1988 = ~w1860 & ~w1864;
assign w1989 = ~w1861 & ~w1988;
assign w1990 = w1987 & w1989;
assign w1991 = ~w1987 & ~w1989;
assign w1992 = ~w1990 & ~w1991;
assign w1993 = ~w1861 & ~w1986;
assign w1994 = (w1993 & w1864) | (w1993 & w16504) | (w1864 & w16504);
assign w1995 = ~w1985 & ~w1994;
assign w1996 = ~w1934 & ~w1982;
assign w1997 = ~w1956 & ~w1979;
assign w1998 = ~w1973 & ~w1977;
assign w1999 = ~pi30 & w1756;
assign w2000 = ~w1945 & ~w1999;
assign w2001 = pi09 & pi23;
assign w2002 = pi04 & pi28;
assign w2003 = pi05 & pi27;
assign w2004 = ~w2002 & ~w2003;
assign w2005 = w2002 & w2003;
assign w2006 = ~w2004 & ~w2005;
assign w2007 = w2001 & ~w2006;
assign w2008 = ~w2001 & w2006;
assign w2009 = ~w2007 & ~w2008;
assign w2010 = pi08 & pi24;
assign w2011 = pi07 & pi25;
assign w2012 = pi06 & pi26;
assign w2013 = ~w2011 & ~w2012;
assign w2014 = w2011 & w2012;
assign w2015 = ~w2013 & ~w2014;
assign w2016 = w2010 & ~w2015;
assign w2017 = ~w2010 & w2015;
assign w2018 = ~w2016 & ~w2017;
assign w2019 = ~w2009 & ~w2018;
assign w2020 = w2009 & w2018;
assign w2021 = ~w2019 & ~w2020;
assign w2022 = w2000 & ~w2021;
assign w2023 = ~w2000 & w2021;
assign w2024 = ~w2022 & ~w2023;
assign w2025 = pi16 & w1939;
assign w2026 = pi00 & pi32;
assign w2027 = pi02 & pi30;
assign w2028 = ~w2026 & ~w2027;
assign w2029 = pi02 & pi32;
assign w2030 = w1748 & w2029;
assign w2031 = ~w2028 & ~w2030;
assign w2032 = w2025 & ~w2031;
assign w2033 = ~w2025 & w2031;
assign w2034 = ~w2032 & ~w2033;
assign w2035 = pi11 & pi21;
assign w2036 = pi13 & pi19;
assign w2037 = pi12 & pi20;
assign w2038 = ~w2036 & ~w2037;
assign w2039 = w2036 & w2037;
assign w2040 = ~w2038 & ~w2039;
assign w2041 = w2035 & ~w2040;
assign w2042 = ~w2035 & w2040;
assign w2043 = ~w2041 & ~w2042;
assign w2044 = ~w2034 & ~w2043;
assign w2045 = w2034 & w2043;
assign w2046 = ~w2044 & ~w2045;
assign w2047 = pi14 & pi18;
assign w2048 = pi03 & pi29;
assign w2049 = pi10 & pi22;
assign w2050 = ~w2048 & ~w2049;
assign w2051 = w2048 & w2049;
assign w2052 = ~w2050 & ~w2051;
assign w2053 = w2047 & ~w2052;
assign w2054 = ~w2047 & w2052;
assign w2055 = ~w2053 & ~w2054;
assign w2056 = w2046 & ~w2055;
assign w2057 = ~w2046 & w2055;
assign w2058 = ~w2056 & ~w2057;
assign w2059 = ~w2024 & ~w2058;
assign w2060 = w2024 & w2058;
assign w2061 = ~w2059 & ~w2060;
assign w2062 = ~w1998 & w2061;
assign w2063 = w1998 & ~w2061;
assign w2064 = ~w2062 & ~w2063;
assign w2065 = ~w1997 & w2064;
assign w2066 = w1997 & ~w2064;
assign w2067 = ~w2065 & ~w2066;
assign w2068 = ~w1950 & ~w1953;
assign w2069 = ~w1884 & ~w1888;
assign w2070 = ~w1887 & ~w2069;
assign w2071 = ~w1872 & ~w1876;
assign w2072 = ~w1875 & ~w2071;
assign w2073 = w2070 & w2072;
assign w2074 = ~w2070 & ~w2072;
assign w2075 = ~w2073 & ~w2074;
assign w2076 = ~w1634 & ~w1920;
assign w2077 = ~w1919 & ~w2076;
assign w2078 = ~w2075 & ~w2077;
assign w2079 = w2075 & w2077;
assign w2080 = ~w2078 & ~w2079;
assign w2081 = pi15 & pi17;
assign w2082 = pi01 & pi31;
assign w2083 = ~w2081 & ~w2082;
assign w2084 = w2081 & w2082;
assign w2085 = ~w2083 & ~w2084;
assign w2086 = ~w1896 & ~w1900;
assign w2087 = ~w1899 & ~w2086;
assign w2088 = w2085 & w2087;
assign w2089 = ~w2085 & ~w2087;
assign w2090 = ~w2088 & ~w2089;
assign w2091 = ~w1905 & ~w1909;
assign w2092 = ~w1908 & ~w2091;
assign w2093 = w2090 & w2092;
assign w2094 = ~w2090 & ~w2092;
assign w2095 = ~w2093 & ~w2094;
assign w2096 = w2080 & w2095;
assign w2097 = ~w2080 & ~w2095;
assign w2098 = ~w2096 & ~w2097;
assign w2099 = w2068 & ~w2098;
assign w2100 = ~w2068 & w2098;
assign w2101 = ~w2099 & ~w2100;
assign w2102 = ~w1914 & ~w1925;
assign w2103 = (~w1881 & ~w1883) | (~w1881 & w17050) | (~w1883 & w17050);
assign w2104 = ~w1963 & ~w1969;
assign w2105 = ~w2103 & ~w2104;
assign w2106 = w2103 & w2104;
assign w2107 = ~w2105 & ~w2106;
assign w2108 = w2102 & ~w2107;
assign w2109 = ~w2102 & w2107;
assign w2110 = ~w2108 & ~w2109;
assign w2111 = ~w1928 & ~w1931;
assign w2112 = ~w2110 & w2111;
assign w2113 = w2110 & ~w2111;
assign w2114 = ~w2112 & ~w2113;
assign w2115 = w2101 & w2114;
assign w2116 = ~w2101 & ~w2114;
assign w2117 = ~w2115 & ~w2116;
assign w2118 = w2067 & w2117;
assign w2119 = ~w2067 & ~w2117;
assign w2120 = ~w2118 & ~w2119;
assign w2121 = ~w1996 & w2120;
assign w2122 = w1996 & ~w2120;
assign w2123 = ~w2121 & ~w2122;
assign w2124 = w1995 & w2123;
assign w2125 = ~w1995 & ~w2123;
assign w2126 = ~w2124 & ~w2125;
assign w2127 = ~w2035 & ~w2039;
assign w2128 = ~w2038 & ~w2127;
assign w2129 = w2025 & ~w2028;
assign w2130 = ~w2030 & ~w2129;
assign w2131 = w2128 & ~w2130;
assign w2132 = ~w2128 & w2130;
assign w2133 = ~w2131 & ~w2132;
assign w2134 = ~w2047 & ~w2051;
assign w2135 = ~w2050 & ~w2134;
assign w2136 = ~w2133 & ~w2135;
assign w2137 = w2133 & w2135;
assign w2138 = ~w2136 & ~w2137;
assign w2139 = ~w2010 & ~w2014;
assign w2140 = ~w2013 & ~w2139;
assign w2141 = ~w2001 & ~w2005;
assign w2142 = ~w2004 & ~w2141;
assign w2143 = w2140 & w2142;
assign w2144 = ~w2140 & ~w2142;
assign w2145 = ~w2143 & ~w2144;
assign w2146 = pi02 & pi31;
assign w2147 = pi00 & pi33;
assign w2148 = pi11 & pi22;
assign w2149 = ~w2147 & ~w2148;
assign w2150 = w2147 & w2148;
assign w2151 = ~w2149 & ~w2150;
assign w2152 = w2146 & ~w2151;
assign w2153 = ~w2146 & w2151;
assign w2154 = ~w2152 & ~w2153;
assign w2155 = ~w2145 & w2154;
assign w2156 = w2145 & ~w2154;
assign w2157 = ~w2155 & ~w2156;
assign w2158 = ~w2138 & ~w2157;
assign w2159 = w2138 & w2157;
assign w2160 = ~w2158 & ~w2159;
assign w2161 = pi03 & pi30;
assign w2162 = pi04 & pi29;
assign w2163 = pi09 & pi24;
assign w2164 = ~w2162 & ~w2163;
assign w2165 = w2162 & w2163;
assign w2166 = ~w2164 & ~w2165;
assign w2167 = w2161 & ~w2166;
assign w2168 = ~w2161 & w2166;
assign w2169 = ~w2167 & ~w2168;
assign w2170 = pi05 & pi28;
assign w2171 = pi08 & pi25;
assign w2172 = pi06 & pi27;
assign w2173 = ~w2171 & ~w2172;
assign w2174 = w2171 & w2172;
assign w2175 = ~w2173 & ~w2174;
assign w2176 = w2170 & ~w2175;
assign w2177 = ~w2170 & w2175;
assign w2178 = ~w2176 & ~w2177;
assign w2179 = ~w2169 & ~w2178;
assign w2180 = w2169 & w2178;
assign w2181 = ~w2179 & ~w2180;
assign w2182 = pi07 & pi26;
assign w2183 = pi16 & pi17;
assign w2184 = pi15 & pi18;
assign w2185 = ~w2183 & ~w2184;
assign w2186 = w2183 & w2184;
assign w2187 = ~w2185 & ~w2186;
assign w2188 = w2182 & ~w2187;
assign w2189 = ~w2182 & w2187;
assign w2190 = ~w2188 & ~w2189;
assign w2191 = w2181 & ~w2190;
assign w2192 = ~w2181 & w2190;
assign w2193 = ~w2191 & ~w2192;
assign w2194 = ~w2160 & ~w2193;
assign w2195 = w2160 & w2193;
assign w2196 = ~w2194 & ~w2195;
assign w2197 = ~w2019 & ~w2023;
assign w2198 = (~w2073 & ~w2075) | (~w2073 & w16838) | (~w2075 & w16838);
assign w2199 = (~w2044 & ~w2046) | (~w2044 & w16717) | (~w2046 & w16717);
assign w2200 = ~w2198 & ~w2199;
assign w2201 = w2198 & w2199;
assign w2202 = ~w2200 & ~w2201;
assign w2203 = w2197 & ~w2202;
assign w2204 = ~w2197 & w2202;
assign w2205 = ~w2203 & ~w2204;
assign w2206 = (~w2060 & w1998) | (~w2060 & w17051) | (w1998 & w17051);
assign w2207 = ~w2205 & w2206;
assign w2208 = w2205 & ~w2206;
assign w2209 = ~w2207 & ~w2208;
assign w2210 = w2196 & w2209;
assign w2211 = ~w2196 & ~w2209;
assign w2212 = ~w2210 & ~w2211;
assign w2213 = (~w2088 & ~w2090) | (~w2088 & w16839) | (~w2090 & w16839);
assign w2214 = pi10 & pi23;
assign w2215 = ~w2084 & ~w2214;
assign w2216 = w2084 & w2214;
assign w2217 = ~w2215 & ~w2216;
assign w2218 = pi01 & pi32;
assign w2219 = pi17 & w2218;
assign w2220 = ~pi17 & ~w2218;
assign w2221 = ~w2219 & ~w2220;
assign w2222 = ~w2217 & w2221;
assign w2223 = w2217 & ~w2221;
assign w2224 = ~w2222 & ~w2223;
assign w2225 = pi12 & pi21;
assign w2226 = pi13 & pi20;
assign w2227 = pi14 & pi19;
assign w2228 = ~w2226 & ~w2227;
assign w2229 = w2226 & w2227;
assign w2230 = ~w2228 & ~w2229;
assign w2231 = w2225 & ~w2230;
assign w2232 = ~w2225 & w2230;
assign w2233 = ~w2231 & ~w2232;
assign w2234 = ~w2224 & ~w2233;
assign w2235 = w2224 & w2233;
assign w2236 = ~w2234 & ~w2235;
assign w2237 = w2213 & ~w2236;
assign w2238 = ~w2213 & w2236;
assign w2239 = ~w2237 & ~w2238;
assign w2240 = (~w2105 & ~w2107) | (~w2105 & w17052) | (~w2107 & w17052);
assign w2241 = ~w2239 & w2240;
assign w2242 = w2239 & ~w2240;
assign w2243 = ~w2241 & ~w2242;
assign w2244 = (~w2096 & w2068) | (~w2096 & w17053) | (w2068 & w17053);
assign w2245 = ~w2243 & w2244;
assign w2246 = w2243 & ~w2244;
assign w2247 = ~w2245 & ~w2246;
assign w2248 = (~w2113 & ~w2114) | (~w2113 & w17054) | (~w2114 & w17054);
assign w2249 = ~w2247 & w2248;
assign w2250 = w2247 & ~w2248;
assign w2251 = ~w2249 & ~w2250;
assign w2252 = w2212 & w2251;
assign w2253 = ~w2212 & ~w2251;
assign w2254 = ~w2252 & ~w2253;
assign w2255 = (~w2065 & ~w2067) | (~w2065 & w17055) | (~w2067 & w17055);
assign w2256 = ~w2254 & w2255;
assign w2257 = w2254 & ~w2255;
assign w2258 = ~w2256 & ~w2257;
assign w2259 = ~w1985 & ~w2121;
assign w2260 = (~w1864 & w16505) | (~w1864 & w16506) | (w16505 & w16506);
assign w2261 = ~w2122 & ~w2260;
assign w2262 = w2258 & w2261;
assign w2263 = ~w2258 & ~w2261;
assign w2264 = ~w2262 & ~w2263;
assign w2265 = ~w2250 & ~w2252;
assign w2266 = (~w2208 & ~w2209) | (~w2208 & w17056) | (~w2209 & w17056);
assign w2267 = (~w2143 & ~w2145) | (~w2143 & w17057) | (~w2145 & w17057);
assign w2268 = (~w2131 & ~w2133) | (~w2131 & w16718) | (~w2133 & w16718);
assign w2269 = pi00 & pi34;
assign w2270 = pi03 & pi31;
assign w2271 = pi04 & pi30;
assign w2272 = ~w2270 & ~w2271;
assign w2273 = w2270 & w2271;
assign w2274 = ~w2272 & ~w2273;
assign w2275 = w2269 & ~w2274;
assign w2276 = ~w2269 & w2274;
assign w2277 = ~w2275 & ~w2276;
assign w2278 = ~w2268 & ~w2277;
assign w2279 = w2268 & w2277;
assign w2280 = ~w2278 & ~w2279;
assign w2281 = ~w2267 & w2280;
assign w2282 = w2267 & ~w2280;
assign w2283 = ~w2281 & ~w2282;
assign w2284 = (~w2159 & ~w2160) | (~w2159 & w16840) | (~w2160 & w16840);
assign w2285 = (~w2200 & ~w2202) | (~w2200 & w16841) | (~w2202 & w16841);
assign w2286 = ~w2284 & ~w2285;
assign w2287 = w2284 & w2285;
assign w2288 = ~w2286 & ~w2287;
assign w2289 = w2283 & w2288;
assign w2290 = ~w2283 & ~w2288;
assign w2291 = ~w2289 & ~w2290;
assign w2292 = ~w2266 & w2291;
assign w2293 = w2266 & ~w2291;
assign w2294 = ~w2292 & ~w2293;
assign w2295 = ~w2146 & ~w2150;
assign w2296 = ~w2149 & ~w2295;
assign w2297 = ~w2161 & ~w2165;
assign w2298 = ~w2164 & ~w2297;
assign w2299 = w2296 & w2298;
assign w2300 = ~w2296 & ~w2298;
assign w2301 = ~w2299 & ~w2300;
assign w2302 = ~w2170 & ~w2174;
assign w2303 = ~w2173 & ~w2302;
assign w2304 = ~w2301 & ~w2303;
assign w2305 = w2301 & w2303;
assign w2306 = ~w2304 & ~w2305;
assign w2307 = (~w2179 & ~w2181) | (~w2179 & w16719) | (~w2181 & w16719);
assign w2308 = pi16 & pi18;
assign w2309 = pi01 & pi33;
assign w2310 = ~w2308 & ~w2309;
assign w2311 = w2308 & w2309;
assign w2312 = ~w2310 & ~w2311;
assign w2313 = w2219 & w2312;
assign w2314 = ~w2219 & ~w2312;
assign w2315 = ~w2313 & ~w2314;
assign w2316 = ~w2182 & ~w2186;
assign w2317 = ~w2185 & ~w2316;
assign w2318 = w2315 & w2317;
assign w2319 = ~w2315 & ~w2317;
assign w2320 = ~w2318 & ~w2319;
assign w2321 = ~w2307 & w2320;
assign w2322 = w2307 & ~w2320;
assign w2323 = ~w2321 & ~w2322;
assign w2324 = w2306 & w2323;
assign w2325 = ~w2306 & ~w2323;
assign w2326 = ~w2324 & ~w2325;
assign w2327 = ~w2225 & ~w2229;
assign w2328 = ~w2228 & ~w2327;
assign w2329 = ~w2216 & ~w2221;
assign w2330 = ~w2215 & ~w2329;
assign w2331 = w2328 & w2330;
assign w2332 = ~w2328 & ~w2330;
assign w2333 = ~w2331 & ~w2332;
assign w2334 = pi12 & pi22;
assign w2335 = ~w1129 & ~w2334;
assign w2336 = w1129 & w2334;
assign w2337 = ~w2335 & ~w2336;
assign w2338 = w2029 & ~w2337;
assign w2339 = ~w2029 & w2337;
assign w2340 = ~w2338 & ~w2339;
assign w2341 = ~w2333 & w2340;
assign w2342 = w2333 & ~w2340;
assign w2343 = ~w2341 & ~w2342;
assign w2344 = (~w2234 & ~w2236) | (~w2234 & w16842) | (~w2236 & w16842);
assign w2345 = w2343 & ~w2344;
assign w2346 = ~w2343 & w2344;
assign w2347 = ~w2345 & ~w2346;
assign w2348 = pi10 & pi24;
assign w2349 = pi05 & pi29;
assign w2350 = pi09 & pi25;
assign w2351 = ~w2349 & ~w2350;
assign w2352 = w2349 & w2350;
assign w2353 = ~w2351 & ~w2352;
assign w2354 = w2348 & ~w2353;
assign w2355 = ~w2348 & w2353;
assign w2356 = ~w2354 & ~w2355;
assign w2357 = pi13 & pi21;
assign w2358 = pi14 & pi20;
assign w2359 = pi15 & pi19;
assign w2360 = ~w2358 & ~w2359;
assign w2361 = w2358 & w2359;
assign w2362 = ~w2360 & ~w2361;
assign w2363 = w2357 & ~w2362;
assign w2364 = ~w2357 & w2362;
assign w2365 = ~w2363 & ~w2364;
assign w2366 = ~w2356 & ~w2365;
assign w2367 = w2356 & w2365;
assign w2368 = ~w2366 & ~w2367;
assign w2369 = pi06 & pi28;
assign w2370 = pi08 & pi26;
assign w2371 = pi07 & pi27;
assign w2372 = ~w2370 & ~w2371;
assign w2373 = w2370 & w2371;
assign w2374 = ~w2372 & ~w2373;
assign w2375 = w2369 & ~w2374;
assign w2376 = ~w2369 & w2374;
assign w2377 = ~w2375 & ~w2376;
assign w2378 = w2368 & ~w2377;
assign w2379 = ~w2368 & w2377;
assign w2380 = ~w2378 & ~w2379;
assign w2381 = w2347 & w2380;
assign w2382 = ~w2347 & ~w2380;
assign w2383 = ~w2381 & ~w2382;
assign w2384 = w2326 & w2383;
assign w2385 = ~w2326 & ~w2383;
assign w2386 = ~w2384 & ~w2385;
assign w2387 = ~w2242 & ~w2246;
assign w2388 = w2386 & ~w2387;
assign w2389 = ~w2386 & w2387;
assign w2390 = ~w2388 & ~w2389;
assign w2391 = w2294 & w2390;
assign w2392 = ~w2294 & ~w2390;
assign w2393 = ~w2391 & ~w2392;
assign w2394 = ~w2265 & w2393;
assign w2395 = w2265 & ~w2393;
assign w2396 = ~w2394 & ~w2395;
assign w2397 = (~w2257 & w2260) | (~w2257 & w16507) | (w2260 & w16507);
assign w2398 = ~w2256 & ~w2397;
assign w2399 = w2396 & w2398;
assign w2400 = ~w2396 & ~w2398;
assign w2401 = ~w2399 & ~w2400;
assign w2402 = ~w2256 & ~w2395;
assign w2403 = (~w2260 & w16508) | (~w2260 & w16509) | (w16508 & w16509);
assign w2404 = ~w2394 & ~w2403;
assign w2405 = ~w2292 & ~w2391;
assign w2406 = ~w2384 & ~w2388;
assign w2407 = (~w2331 & ~w2333) | (~w2331 & w17058) | (~w2333 & w17058);
assign w2408 = (~w2299 & ~w2301) | (~w2299 & w16843) | (~w2301 & w16843);
assign w2409 = (~w2313 & ~w2315) | (~w2313 & w17059) | (~w2315 & w17059);
assign w2410 = ~w2408 & ~w2409;
assign w2411 = w2408 & w2409;
assign w2412 = ~w2410 & ~w2411;
assign w2413 = w2407 & ~w2412;
assign w2414 = ~w2407 & w2412;
assign w2415 = ~w2413 & ~w2414;
assign w2416 = (~w2321 & ~w2323) | (~w2321 & w16844) | (~w2323 & w16844);
assign w2417 = ~w2415 & w2416;
assign w2418 = w2415 & ~w2416;
assign w2419 = ~w2417 & ~w2418;
assign w2420 = (~w2345 & ~w2347) | (~w2345 & w17060) | (~w2347 & w17060);
assign w2421 = w2419 & ~w2420;
assign w2422 = ~w2419 & w2420;
assign w2423 = ~w2421 & ~w2422;
assign w2424 = ~w2406 & w2423;
assign w2425 = w2406 & ~w2423;
assign w2426 = ~w2424 & ~w2425;
assign w2427 = (~w2286 & ~w2288) | (~w2286 & w17061) | (~w2288 & w17061);
assign w2428 = ~w2029 & ~w2336;
assign w2429 = ~w2335 & ~w2428;
assign w2430 = ~w2357 & ~w2361;
assign w2431 = ~w2360 & ~w2430;
assign w2432 = w2429 & w2431;
assign w2433 = ~w2429 & ~w2431;
assign w2434 = ~w2432 & ~w2433;
assign w2435 = ~w2269 & ~w2273;
assign w2436 = ~w2272 & ~w2435;
assign w2437 = ~w2434 & ~w2436;
assign w2438 = w2434 & w2436;
assign w2439 = ~w2437 & ~w2438;
assign w2440 = (~w2366 & ~w2368) | (~w2366 & w16845) | (~w2368 & w16845);
assign w2441 = pi34 & w684;
assign w2442 = pi01 & pi34;
assign w2443 = ~pi18 & ~w2442;
assign w2444 = ~w2441 & ~w2443;
assign w2445 = ~w2369 & ~w2373;
assign w2446 = ~w2372 & ~w2445;
assign w2447 = w2444 & w2446;
assign w2448 = ~w2444 & ~w2446;
assign w2449 = ~w2447 & ~w2448;
assign w2450 = ~w2348 & ~w2352;
assign w2451 = ~w2351 & ~w2450;
assign w2452 = w2449 & w2451;
assign w2453 = ~w2449 & ~w2451;
assign w2454 = ~w2452 & ~w2453;
assign w2455 = ~w2440 & w2454;
assign w2456 = w2440 & ~w2454;
assign w2457 = ~w2455 & ~w2456;
assign w2458 = w2439 & w2457;
assign w2459 = ~w2439 & ~w2457;
assign w2460 = ~w2458 & ~w2459;
assign w2461 = ~w2427 & w2460;
assign w2462 = w2427 & ~w2460;
assign w2463 = ~w2461 & ~w2462;
assign w2464 = (~w2278 & ~w2280) | (~w2278 & w16846) | (~w2280 & w16846);
assign w2465 = pi07 & pi28;
assign w2466 = pi17 & pi18;
assign w2467 = pi16 & pi19;
assign w2468 = ~w2466 & ~w2467;
assign w2469 = w2466 & w2467;
assign w2470 = ~w2468 & ~w2469;
assign w2471 = w2465 & ~w2470;
assign w2472 = ~w2465 & w2470;
assign w2473 = ~w2471 & ~w2472;
assign w2474 = pi05 & pi30;
assign w2475 = pi08 & pi27;
assign w2476 = pi06 & pi29;
assign w2477 = ~w2475 & ~w2476;
assign w2478 = w2475 & w2476;
assign w2479 = ~w2477 & ~w2478;
assign w2480 = w2474 & ~w2479;
assign w2481 = ~w2474 & w2479;
assign w2482 = ~w2480 & ~w2481;
assign w2483 = ~w2473 & ~w2482;
assign w2484 = w2473 & w2482;
assign w2485 = ~w2483 & ~w2484;
assign w2486 = pi04 & pi31;
assign w2487 = pi09 & pi26;
assign w2488 = pi10 & pi25;
assign w2489 = ~w2487 & ~w2488;
assign w2490 = w2487 & w2488;
assign w2491 = ~w2489 & ~w2490;
assign w2492 = w2486 & ~w2491;
assign w2493 = ~w2486 & w2491;
assign w2494 = ~w2492 & ~w2493;
assign w2495 = w2485 & ~w2494;
assign w2496 = ~w2485 & w2494;
assign w2497 = ~w2495 & ~w2496;
assign w2498 = ~w2464 & w2497;
assign w2499 = w2464 & ~w2497;
assign w2500 = ~w2498 & ~w2499;
assign w2501 = pi00 & pi35;
assign w2502 = pi02 & pi33;
assign w2503 = ~w2501 & ~w2502;
assign w2504 = pi02 & pi35;
assign w2505 = w2147 & w2504;
assign w2506 = ~w2503 & ~w2505;
assign w2507 = w2311 & ~w2506;
assign w2508 = ~w2311 & w2506;
assign w2509 = ~w2507 & ~w2508;
assign w2510 = pi03 & pi32;
assign w2511 = pi12 & pi23;
assign w2512 = pi11 & pi24;
assign w2513 = ~w2511 & ~w2512;
assign w2514 = w2511 & w2512;
assign w2515 = ~w2513 & ~w2514;
assign w2516 = w2510 & ~w2515;
assign w2517 = ~w2510 & w2515;
assign w2518 = ~w2516 & ~w2517;
assign w2519 = ~w2509 & ~w2518;
assign w2520 = w2509 & w2518;
assign w2521 = ~w2519 & ~w2520;
assign w2522 = pi13 & pi22;
assign w2523 = pi15 & pi20;
assign w2524 = pi14 & pi21;
assign w2525 = ~w2523 & ~w2524;
assign w2526 = w2523 & w2524;
assign w2527 = ~w2525 & ~w2526;
assign w2528 = w2522 & ~w2527;
assign w2529 = ~w2522 & w2527;
assign w2530 = ~w2528 & ~w2529;
assign w2531 = w2521 & ~w2530;
assign w2532 = ~w2521 & w2530;
assign w2533 = ~w2531 & ~w2532;
assign w2534 = w2500 & w2533;
assign w2535 = ~w2500 & ~w2533;
assign w2536 = ~w2534 & ~w2535;
assign w2537 = w2463 & w2536;
assign w2538 = ~w2463 & ~w2536;
assign w2539 = ~w2537 & ~w2538;
assign w2540 = ~w2426 & ~w2539;
assign w2541 = w2426 & w2539;
assign w2542 = ~w2540 & ~w2541;
assign w2543 = w2405 & ~w2542;
assign w2544 = ~w2405 & w2542;
assign w2545 = ~w2543 & ~w2544;
assign w2546 = w2404 & w2545;
assign w2547 = ~w2404 & ~w2545;
assign w2548 = ~w2546 & ~w2547;
assign w2549 = (~w2424 & ~w2426) | (~w2424 & w16847) | (~w2426 & w16847);
assign w2550 = (~w2461 & ~w2463) | (~w2461 & w16848) | (~w2463 & w16848);
assign w2551 = (~w2519 & ~w2521) | (~w2519 & w16849) | (~w2521 & w16849);
assign w2552 = (~w2432 & ~w2434) | (~w2432 & w16720) | (~w2434 & w16720);
assign w2553 = (~w2447 & ~w2449) | (~w2447 & w16721) | (~w2449 & w16721);
assign w2554 = ~w2552 & ~w2553;
assign w2555 = w2552 & w2553;
assign w2556 = ~w2554 & ~w2555;
assign w2557 = w2551 & ~w2556;
assign w2558 = ~w2551 & w2556;
assign w2559 = ~w2557 & ~w2558;
assign w2560 = (~w2455 & ~w2457) | (~w2455 & w16850) | (~w2457 & w16850);
assign w2561 = ~w2559 & w2560;
assign w2562 = w2559 & ~w2560;
assign w2563 = ~w2561 & ~w2562;
assign w2564 = (~w2498 & ~w2500) | (~w2498 & w16851) | (~w2500 & w16851);
assign w2565 = w2563 & ~w2564;
assign w2566 = ~w2563 & w2564;
assign w2567 = ~w2565 & ~w2566;
assign w2568 = ~w2550 & w2567;
assign w2569 = w2550 & ~w2567;
assign w2570 = ~w2568 & ~w2569;
assign w2571 = pi02 & pi34;
assign w2572 = pi12 & pi24;
assign w2573 = pi13 & pi23;
assign w2574 = ~w2572 & ~w2573;
assign w2575 = w2572 & w2573;
assign w2576 = ~w2574 & ~w2575;
assign w2577 = w2571 & ~w2576;
assign w2578 = ~w2571 & w2576;
assign w2579 = ~w2577 & ~w2578;
assign w2580 = pi10 & pi26;
assign w2581 = pi05 & pi31;
assign w2582 = pi09 & pi27;
assign w2583 = ~w2581 & ~w2582;
assign w2584 = w2581 & w2582;
assign w2585 = ~w2583 & ~w2584;
assign w2586 = w2580 & ~w2585;
assign w2587 = ~w2580 & w2585;
assign w2588 = ~w2586 & ~w2587;
assign w2589 = ~w2579 & ~w2588;
assign w2590 = w2579 & w2588;
assign w2591 = ~w2589 & ~w2590;
assign w2592 = pi06 & pi30;
assign w2593 = pi08 & pi28;
assign w2594 = pi07 & pi29;
assign w2595 = ~w2593 & ~w2594;
assign w2596 = w2593 & w2594;
assign w2597 = ~w2595 & ~w2596;
assign w2598 = w2592 & ~w2597;
assign w2599 = ~w2592 & w2597;
assign w2600 = ~w2598 & ~w2599;
assign w2601 = w2591 & ~w2600;
assign w2602 = ~w2591 & w2600;
assign w2603 = ~w2601 & ~w2602;
assign w2604 = (~w2410 & ~w2412) | (~w2410 & w17062) | (~w2412 & w17062);
assign w2605 = pi00 & pi36;
assign w2606 = w2441 & w2605;
assign w2607 = ~w2441 & ~w2605;
assign w2608 = ~w2606 & ~w2607;
assign w2609 = pi17 & pi19;
assign w2610 = pi01 & pi35;
assign w2611 = ~w2609 & ~w2610;
assign w2612 = w2609 & w2610;
assign w2613 = ~w2611 & ~w2612;
assign w2614 = w2608 & w2613;
assign w2615 = ~w2608 & ~w2613;
assign w2616 = ~w2614 & ~w2615;
assign w2617 = pi03 & pi33;
assign w2618 = pi04 & pi32;
assign w2619 = pi11 & pi25;
assign w2620 = ~w2618 & ~w2619;
assign w2621 = w2618 & w2619;
assign w2622 = ~w2620 & ~w2621;
assign w2623 = w2617 & ~w2622;
assign w2624 = ~w2617 & w2622;
assign w2625 = ~w2623 & ~w2624;
assign w2626 = pi14 & pi22;
assign w2627 = pi15 & pi21;
assign w2628 = pi16 & pi20;
assign w2629 = ~w2627 & ~w2628;
assign w2630 = w2627 & w2628;
assign w2631 = ~w2629 & ~w2630;
assign w2632 = w2626 & ~w2631;
assign w2633 = ~w2626 & w2631;
assign w2634 = ~w2632 & ~w2633;
assign w2635 = ~w2625 & ~w2634;
assign w2636 = w2625 & w2634;
assign w2637 = ~w2635 & ~w2636;
assign w2638 = w2616 & w2637;
assign w2639 = ~w2616 & ~w2637;
assign w2640 = ~w2638 & ~w2639;
assign w2641 = ~w2604 & w2640;
assign w2642 = w2604 & ~w2640;
assign w2643 = ~w2641 & ~w2642;
assign w2644 = w2603 & w2643;
assign w2645 = ~w2603 & ~w2643;
assign w2646 = ~w2644 & ~w2645;
assign w2647 = ~w2486 & ~w2490;
assign w2648 = ~w2489 & ~w2647;
assign w2649 = ~w2474 & ~w2478;
assign w2650 = ~w2477 & ~w2649;
assign w2651 = w2648 & w2650;
assign w2652 = ~w2648 & ~w2650;
assign w2653 = ~w2651 & ~w2652;
assign w2654 = ~w2465 & ~w2469;
assign w2655 = ~w2468 & ~w2654;
assign w2656 = ~w2653 & ~w2655;
assign w2657 = w2653 & w2655;
assign w2658 = ~w2656 & ~w2657;
assign w2659 = ~w2522 & ~w2526;
assign w2660 = ~w2525 & ~w2659;
assign w2661 = ~w2510 & ~w2514;
assign w2662 = ~w2513 & ~w2661;
assign w2663 = w2660 & w2662;
assign w2664 = ~w2660 & ~w2662;
assign w2665 = ~w2663 & ~w2664;
assign w2666 = w2311 & ~w2503;
assign w2667 = ~w2505 & ~w2666;
assign w2668 = ~w2665 & w2667;
assign w2669 = w2665 & ~w2667;
assign w2670 = ~w2668 & ~w2669;
assign w2671 = (~w2483 & ~w2485) | (~w2483 & w17063) | (~w2485 & w17063);
assign w2672 = ~w2670 & w2671;
assign w2673 = w2670 & ~w2671;
assign w2674 = ~w2672 & ~w2673;
assign w2675 = w2658 & w2674;
assign w2676 = ~w2658 & ~w2674;
assign w2677 = ~w2675 & ~w2676;
assign w2678 = (w2677 & w2421) | (w2677 & w16852) | (w2421 & w16852);
assign w2679 = ~w2421 & w16853;
assign w2680 = ~w2678 & ~w2679;
assign w2681 = w2646 & w2680;
assign w2682 = ~w2646 & ~w2680;
assign w2683 = ~w2681 & ~w2682;
assign w2684 = w2570 & w2683;
assign w2685 = ~w2570 & ~w2683;
assign w2686 = ~w2684 & ~w2685;
assign w2687 = w2549 & ~w2686;
assign w2688 = ~w2549 & w2686;
assign w2689 = ~w2687 & ~w2688;
assign w2690 = ~w2394 & ~w2544;
assign w2691 = (~w2260 & w16510) | (~w2260 & w16511) | (w16510 & w16511);
assign w2692 = w2689 & w2691;
assign w2693 = ~w2689 & ~w2691;
assign w2694 = ~w2692 & ~w2693;
assign w2695 = ~w2568 & ~w2684;
assign w2696 = (~w2663 & ~w2665) | (~w2663 & w17064) | (~w2665 & w17064);
assign w2697 = pi08 & pi29;
assign w2698 = pi18 & pi19;
assign w2699 = pi17 & pi20;
assign w2700 = ~w2698 & ~w2699;
assign w2701 = w2698 & w2699;
assign w2702 = ~w2700 & ~w2701;
assign w2703 = w2697 & ~w2702;
assign w2704 = ~w2697 & w2702;
assign w2705 = ~w2703 & ~w2704;
assign w2706 = pi11 & pi26;
assign w2707 = pi05 & pi32;
assign w2708 = pi10 & pi27;
assign w2709 = ~w2707 & ~w2708;
assign w2710 = w2707 & w2708;
assign w2711 = ~w2709 & ~w2710;
assign w2712 = w2706 & ~w2711;
assign w2713 = ~w2706 & w2711;
assign w2714 = ~w2712 & ~w2713;
assign w2715 = ~w2705 & ~w2714;
assign w2716 = w2705 & w2714;
assign w2717 = ~w2715 & ~w2716;
assign w2718 = w2696 & ~w2717;
assign w2719 = ~w2696 & w2717;
assign w2720 = ~w2718 & ~w2719;
assign w2721 = (~w2554 & ~w2556) | (~w2554 & w16854) | (~w2556 & w16854);
assign w2722 = ~w2720 & w2721;
assign w2723 = w2720 & ~w2721;
assign w2724 = ~w2722 & ~w2723;
assign w2725 = pi16 & pi21;
assign w2726 = pi03 & pi34;
assign w2727 = ~w2504 & ~w2726;
assign w2728 = pi03 & pi35;
assign w2729 = w2571 & w2728;
assign w2730 = ~w2727 & ~w2729;
assign w2731 = w2725 & ~w2730;
assign w2732 = ~w2725 & w2730;
assign w2733 = ~w2731 & ~w2732;
assign w2734 = pi00 & pi37;
assign w2735 = pi12 & pi25;
assign w2736 = pi04 & pi33;
assign w2737 = ~w2735 & ~w2736;
assign w2738 = w2735 & w2736;
assign w2739 = ~w2737 & ~w2738;
assign w2740 = w2734 & ~w2739;
assign w2741 = ~w2734 & w2739;
assign w2742 = ~w2740 & ~w2741;
assign w2743 = ~w2733 & ~w2742;
assign w2744 = w2733 & w2742;
assign w2745 = ~w2743 & ~w2744;
assign w2746 = pi09 & pi28;
assign w2747 = pi06 & pi31;
assign w2748 = pi07 & pi30;
assign w2749 = ~w2747 & ~w2748;
assign w2750 = w2747 & w2748;
assign w2751 = ~w2749 & ~w2750;
assign w2752 = w2746 & ~w2751;
assign w2753 = ~w2746 & w2751;
assign w2754 = ~w2752 & ~w2753;
assign w2755 = w2745 & ~w2754;
assign w2756 = ~w2745 & w2754;
assign w2757 = ~w2755 & ~w2756;
assign w2758 = ~w2724 & ~w2757;
assign w2759 = w2724 & w2757;
assign w2760 = ~w2758 & ~w2759;
assign w2761 = (~w2606 & ~w2608) | (~w2606 & w16855) | (~w2608 & w16855);
assign w2762 = ~w2580 & ~w2584;
assign w2763 = ~w2583 & ~w2762;
assign w2764 = ~w2761 & w2763;
assign w2765 = w2761 & ~w2763;
assign w2766 = ~w2764 & ~w2765;
assign w2767 = pi13 & pi24;
assign w2768 = pi14 & pi23;
assign w2769 = pi15 & pi22;
assign w2770 = ~w2768 & ~w2769;
assign w2771 = w2768 & w2769;
assign w2772 = ~w2770 & ~w2771;
assign w2773 = w2767 & ~w2772;
assign w2774 = ~w2767 & w2772;
assign w2775 = ~w2773 & ~w2774;
assign w2776 = ~w2766 & w2775;
assign w2777 = w2766 & ~w2775;
assign w2778 = ~w2776 & ~w2777;
assign w2779 = ~w2626 & ~w2630;
assign w2780 = ~w2629 & ~w2779;
assign w2781 = ~w2617 & ~w2621;
assign w2782 = ~w2620 & ~w2781;
assign w2783 = w2780 & w2782;
assign w2784 = ~w2780 & ~w2782;
assign w2785 = ~w2783 & ~w2784;
assign w2786 = ~w2571 & ~w2575;
assign w2787 = ~w2574 & ~w2786;
assign w2788 = ~w2785 & ~w2787;
assign w2789 = w2785 & w2787;
assign w2790 = ~w2788 & ~w2789;
assign w2791 = ~w2635 & ~w2638;
assign w2792 = ~w2790 & w2791;
assign w2793 = w2790 & ~w2791;
assign w2794 = ~w2792 & ~w2793;
assign w2795 = w2778 & w2794;
assign w2796 = ~w2778 & ~w2794;
assign w2797 = ~w2795 & ~w2796;
assign w2798 = (w2797 & w2565) | (w2797 & w17065) | (w2565 & w17065);
assign w2799 = ~w2565 & w17066;
assign w2800 = ~w2798 & ~w2799;
assign w2801 = w2760 & w2800;
assign w2802 = ~w2760 & ~w2800;
assign w2803 = ~w2801 & ~w2802;
assign w2804 = (~w2678 & ~w2680) | (~w2678 & w17067) | (~w2680 & w17067);
assign w2805 = ~w2641 & ~w2644;
assign w2806 = ~w2673 & ~w2675;
assign w2807 = ~w2589 & ~w2601;
assign w2808 = (~w2651 & ~w2653) | (~w2651 & w17068) | (~w2653 & w17068);
assign w2809 = ~pi36 & w2612;
assign w2810 = pi36 & w792;
assign w2811 = pi01 & pi36;
assign w2812 = ~pi19 & ~w2811;
assign w2813 = ~w2810 & ~w2812;
assign w2814 = ~w2612 & ~w2813;
assign w2815 = ~w2809 & ~w2814;
assign w2816 = ~w2592 & ~w2596;
assign w2817 = ~w2595 & ~w2816;
assign w2818 = w2815 & w2817;
assign w2819 = ~w2815 & ~w2817;
assign w2820 = ~w2818 & ~w2819;
assign w2821 = ~w2808 & w2820;
assign w2822 = w2808 & ~w2820;
assign w2823 = ~w2821 & ~w2822;
assign w2824 = ~w2807 & w2823;
assign w2825 = w2807 & ~w2823;
assign w2826 = ~w2824 & ~w2825;
assign w2827 = ~w2806 & w2826;
assign w2828 = w2806 & ~w2826;
assign w2829 = ~w2827 & ~w2828;
assign w2830 = ~w2805 & w2829;
assign w2831 = w2805 & ~w2829;
assign w2832 = ~w2830 & ~w2831;
assign w2833 = ~w2804 & w2832;
assign w2834 = w2804 & ~w2832;
assign w2835 = ~w2833 & ~w2834;
assign w2836 = w2803 & w2835;
assign w2837 = ~w2803 & ~w2835;
assign w2838 = ~w2836 & ~w2837;
assign w2839 = ~w2695 & w2838;
assign w2840 = w2695 & ~w2838;
assign w2841 = ~w2839 & ~w2840;
assign w2842 = ~w2688 & ~w2691;
assign w2843 = ~w2687 & ~w2842;
assign w2844 = w2841 & w2843;
assign w2845 = ~w2841 & ~w2843;
assign w2846 = ~w2844 & ~w2845;
assign w2847 = ~w2833 & ~w2836;
assign w2848 = ~w2827 & ~w2830;
assign w2849 = pi18 & pi20;
assign w2850 = pi01 & pi37;
assign w2851 = ~w2849 & ~w2850;
assign w2852 = w2849 & w2850;
assign w2853 = ~w2851 & ~w2852;
assign w2854 = ~w2697 & ~w2701;
assign w2855 = ~w2700 & ~w2854;
assign w2856 = w2853 & w2855;
assign w2857 = ~w2853 & ~w2855;
assign w2858 = ~w2856 & ~w2857;
assign w2859 = ~w2746 & ~w2750;
assign w2860 = ~w2749 & ~w2859;
assign w2861 = w2858 & w2860;
assign w2862 = ~w2858 & ~w2860;
assign w2863 = ~w2861 & ~w2862;
assign w2864 = (~w2764 & ~w2766) | (~w2764 & w17069) | (~w2766 & w17069);
assign w2865 = (~w2743 & ~w2745) | (~w2743 & w17070) | (~w2745 & w17070);
assign w2866 = ~w2864 & ~w2865;
assign w2867 = w2864 & w2865;
assign w2868 = ~w2866 & ~w2867;
assign w2869 = w2863 & w2868;
assign w2870 = ~w2863 & ~w2868;
assign w2871 = ~w2869 & ~w2870;
assign w2872 = ~w2848 & w2871;
assign w2873 = w2848 & ~w2871;
assign w2874 = ~w2872 & ~w2873;
assign w2875 = (~w2783 & ~w2785) | (~w2783 & w17071) | (~w2785 & w17071);
assign w2876 = (~w2809 & ~w2815) | (~w2809 & w16856) | (~w2815 & w16856);
assign w2877 = pi12 & pi26;
assign w2878 = pi04 & pi34;
assign w2879 = pi11 & pi27;
assign w2880 = ~w2878 & ~w2879;
assign w2881 = w2878 & w2879;
assign w2882 = ~w2880 & ~w2881;
assign w2883 = w2877 & ~w2882;
assign w2884 = ~w2877 & w2882;
assign w2885 = ~w2883 & ~w2884;
assign w2886 = ~w2876 & ~w2885;
assign w2887 = w2876 & w2885;
assign w2888 = ~w2886 & ~w2887;
assign w2889 = w2875 & ~w2888;
assign w2890 = ~w2875 & w2888;
assign w2891 = ~w2889 & ~w2890;
assign w2892 = ~w2821 & ~w2824;
assign w2893 = ~w2706 & ~w2710;
assign w2894 = ~w2709 & ~w2893;
assign w2895 = pi00 & pi38;
assign w2896 = pi02 & pi36;
assign w2897 = ~w2895 & ~w2896;
assign w2898 = pi02 & pi38;
assign w2899 = w2605 & w2898;
assign w2900 = ~w2897 & ~w2899;
assign w2901 = w2810 & ~w2900;
assign w2902 = ~w2810 & w2900;
assign w2903 = ~w2901 & ~w2902;
assign w2904 = w2894 & ~w2903;
assign w2905 = ~w2894 & w2903;
assign w2906 = ~w2904 & ~w2905;
assign w2907 = pi13 & pi25;
assign w2908 = pi14 & pi24;
assign w2909 = ~w2907 & ~w2908;
assign w2910 = w2907 & w2908;
assign w2911 = ~w2909 & ~w2910;
assign w2912 = w2728 & ~w2911;
assign w2913 = ~w2728 & w2911;
assign w2914 = ~w2912 & ~w2913;
assign w2915 = w2906 & ~w2914;
assign w2916 = ~w2906 & w2914;
assign w2917 = ~w2915 & ~w2916;
assign w2918 = ~w2892 & w2917;
assign w2919 = w2892 & ~w2917;
assign w2920 = ~w2918 & ~w2919;
assign w2921 = w2891 & w2920;
assign w2922 = ~w2891 & ~w2920;
assign w2923 = ~w2921 & ~w2922;
assign w2924 = w2874 & w2923;
assign w2925 = ~w2874 & ~w2923;
assign w2926 = ~w2924 & ~w2925;
assign w2927 = ~w2734 & ~w2738;
assign w2928 = ~w2737 & ~w2927;
assign w2929 = w2725 & ~w2727;
assign w2930 = ~w2729 & ~w2929;
assign w2931 = w2928 & ~w2930;
assign w2932 = ~w2928 & w2930;
assign w2933 = ~w2931 & ~w2932;
assign w2934 = ~w2767 & ~w2771;
assign w2935 = ~w2770 & ~w2934;
assign w2936 = ~w2933 & ~w2935;
assign w2937 = w2933 & w2935;
assign w2938 = ~w2936 & ~w2937;
assign w2939 = ~w2715 & ~w2719;
assign w2940 = ~w2938 & w2939;
assign w2941 = w2938 & ~w2939;
assign w2942 = ~w2940 & ~w2941;
assign w2943 = pi05 & pi33;
assign w2944 = pi06 & pi32;
assign w2945 = pi10 & pi28;
assign w2946 = ~w2944 & ~w2945;
assign w2947 = w2944 & w2945;
assign w2948 = ~w2946 & ~w2947;
assign w2949 = w2943 & ~w2948;
assign w2950 = ~w2943 & w2948;
assign w2951 = ~w2949 & ~w2950;
assign w2952 = pi15 & pi23;
assign w2953 = pi16 & pi22;
assign w2954 = pi17 & pi21;
assign w2955 = ~w2953 & ~w2954;
assign w2956 = w2953 & w2954;
assign w2957 = ~w2955 & ~w2956;
assign w2958 = w2952 & ~w2957;
assign w2959 = ~w2952 & w2957;
assign w2960 = ~w2958 & ~w2959;
assign w2961 = ~w2951 & ~w2960;
assign w2962 = w2951 & w2960;
assign w2963 = ~w2961 & ~w2962;
assign w2964 = pi09 & pi29;
assign w2965 = pi07 & pi31;
assign w2966 = pi08 & pi30;
assign w2967 = ~w2965 & ~w2966;
assign w2968 = w2965 & w2966;
assign w2969 = ~w2967 & ~w2968;
assign w2970 = w2964 & ~w2969;
assign w2971 = ~w2964 & w2969;
assign w2972 = ~w2970 & ~w2971;
assign w2973 = w2963 & ~w2972;
assign w2974 = ~w2963 & w2972;
assign w2975 = ~w2973 & ~w2974;
assign w2976 = w2942 & w2975;
assign w2977 = ~w2942 & ~w2975;
assign w2978 = ~w2976 & ~w2977;
assign w2979 = (~w2723 & ~w2724) | (~w2723 & w17072) | (~w2724 & w17072);
assign w2980 = ~w2793 & ~w2795;
assign w2981 = ~w2979 & ~w2980;
assign w2982 = w2979 & w2980;
assign w2983 = ~w2981 & ~w2982;
assign w2984 = w2978 & w2983;
assign w2985 = ~w2978 & ~w2983;
assign w2986 = ~w2984 & ~w2985;
assign w2987 = ~w2798 & ~w2801;
assign w2988 = w2986 & ~w2987;
assign w2989 = ~w2986 & w2987;
assign w2990 = ~w2988 & ~w2989;
assign w2991 = ~w2926 & ~w2990;
assign w2992 = w2926 & w2990;
assign w2993 = ~w2991 & ~w2992;
assign w2994 = ~w2847 & w2993;
assign w2995 = w2847 & ~w2993;
assign w2996 = ~w2994 & ~w2995;
assign w2997 = ~w2687 & ~w2840;
assign w2998 = (w2997 & w2691) | (w2997 & w16512) | (w2691 & w16512);
assign w2999 = ~w2839 & ~w2998;
assign w3000 = w2996 & w2999;
assign w3001 = ~w2996 & ~w2999;
assign w3002 = ~w3000 & ~w3001;
assign w3003 = ~w2988 & ~w2992;
assign w3004 = ~w2872 & ~w2924;
assign w3005 = ~w2918 & ~w2921;
assign w3006 = ~w2931 & ~w2937;
assign w3007 = (~w2856 & ~w2858) | (~w2856 & w16857) | (~w2858 & w16857);
assign w3008 = pi38 & w878;
assign w3009 = pi01 & pi38;
assign w3010 = ~pi20 & ~w3009;
assign w3011 = ~w3008 & ~w3010;
assign w3012 = pi00 & pi39;
assign w3013 = w2852 & w3012;
assign w3014 = ~w2852 & ~w3012;
assign w3015 = ~w3013 & ~w3014;
assign w3016 = w3011 & w3015;
assign w3017 = ~w3011 & ~w3015;
assign w3018 = ~w3016 & ~w3017;
assign w3019 = ~w3007 & w3018;
assign w3020 = w3007 & ~w3018;
assign w3021 = ~w3019 & ~w3020;
assign w3022 = w3006 & ~w3021;
assign w3023 = ~w3006 & w3021;
assign w3024 = ~w3022 & ~w3023;
assign w3025 = ~w2728 & ~w2910;
assign w3026 = ~w2909 & ~w3025;
assign w3027 = ~w2810 & ~w2899;
assign w3028 = ~w2897 & ~w3027;
assign w3029 = w3026 & w3028;
assign w3030 = ~w3026 & ~w3028;
assign w3031 = ~w3029 & ~w3030;
assign w3032 = ~w2952 & ~w2956;
assign w3033 = ~w2955 & ~w3032;
assign w3034 = ~w3031 & ~w3033;
assign w3035 = w3031 & w3033;
assign w3036 = ~w3034 & ~w3035;
assign w3037 = (~w2961 & ~w2963) | (~w2961 & w16858) | (~w2963 & w16858);
assign w3038 = (~w2904 & ~w2906) | (~w2904 & w16859) | (~w2906 & w16859);
assign w3039 = ~w3037 & ~w3038;
assign w3040 = w3037 & w3038;
assign w3041 = ~w3039 & ~w3040;
assign w3042 = w3036 & w3041;
assign w3043 = ~w3036 & ~w3041;
assign w3044 = ~w3042 & ~w3043;
assign w3045 = w3024 & w3044;
assign w3046 = ~w3024 & ~w3044;
assign w3047 = ~w3045 & ~w3046;
assign w3048 = ~w3005 & w3047;
assign w3049 = w3005 & ~w3047;
assign w3050 = ~w3048 & ~w3049;
assign w3051 = ~w3004 & w3050;
assign w3052 = w3004 & ~w3050;
assign w3053 = ~w3051 & ~w3052;
assign w3054 = ~w2981 & ~w2984;
assign w3055 = ~w2877 & ~w2881;
assign w3056 = ~w2880 & ~w3055;
assign w3057 = ~w2964 & ~w2968;
assign w3058 = ~w2967 & ~w3057;
assign w3059 = w3056 & w3058;
assign w3060 = ~w3056 & ~w3058;
assign w3061 = ~w3059 & ~w3060;
assign w3062 = ~w2943 & ~w2947;
assign w3063 = ~w2946 & ~w3062;
assign w3064 = ~w3061 & ~w3063;
assign w3065 = w3061 & w3063;
assign w3066 = ~w3064 & ~w3065;
assign w3067 = (~w2886 & ~w2888) | (~w2886 & w17073) | (~w2888 & w17073);
assign w3068 = ~w3066 & w3067;
assign w3069 = w3066 & ~w3067;
assign w3070 = ~w3068 & ~w3069;
assign w3071 = pi17 & pi22;
assign w3072 = pi04 & pi35;
assign w3073 = pi12 & pi27;
assign w3074 = ~w3072 & ~w3073;
assign w3075 = w3072 & w3073;
assign w3076 = ~w3074 & ~w3075;
assign w3077 = w3071 & ~w3076;
assign w3078 = ~w3071 & w3076;
assign w3079 = ~w3077 & ~w3078;
assign w3080 = pi08 & pi31;
assign w3081 = pi19 & pi20;
assign w3082 = pi18 & pi21;
assign w3083 = ~w3081 & ~w3082;
assign w3084 = w3081 & w3082;
assign w3085 = ~w3083 & ~w3084;
assign w3086 = w3080 & ~w3085;
assign w3087 = ~w3080 & w3085;
assign w3088 = ~w3086 & ~w3087;
assign w3089 = ~w3079 & ~w3088;
assign w3090 = w3079 & w3088;
assign w3091 = ~w3089 & ~w3090;
assign w3092 = pi11 & pi28;
assign w3093 = pi10 & pi29;
assign w3094 = pi05 & pi34;
assign w3095 = ~w3093 & ~w3094;
assign w3096 = w3093 & w3094;
assign w3097 = ~w3095 & ~w3096;
assign w3098 = w3092 & ~w3097;
assign w3099 = ~w3092 & w3097;
assign w3100 = ~w3098 & ~w3099;
assign w3101 = w3091 & ~w3100;
assign w3102 = ~w3091 & w3100;
assign w3103 = ~w3101 & ~w3102;
assign w3104 = w3070 & w3103;
assign w3105 = ~w3070 & ~w3103;
assign w3106 = ~w3104 & ~w3105;
assign w3107 = ~w3054 & w3106;
assign w3108 = w3054 & ~w3106;
assign w3109 = ~w3107 & ~w3108;
assign w3110 = ~w2941 & ~w2976;
assign w3111 = ~w2866 & ~w2869;
assign w3112 = pi02 & pi37;
assign w3113 = pi03 & pi36;
assign w3114 = pi13 & pi26;
assign w3115 = ~w3113 & ~w3114;
assign w3116 = w3113 & w3114;
assign w3117 = ~w3115 & ~w3116;
assign w3118 = w3112 & ~w3117;
assign w3119 = ~w3112 & w3117;
assign w3120 = ~w3118 & ~w3119;
assign w3121 = pi14 & pi25;
assign w3122 = pi15 & pi24;
assign w3123 = pi16 & pi23;
assign w3124 = ~w3122 & ~w3123;
assign w3125 = w3122 & w3123;
assign w3126 = ~w3124 & ~w3125;
assign w3127 = w3121 & ~w3126;
assign w3128 = ~w3121 & w3126;
assign w3129 = ~w3127 & ~w3128;
assign w3130 = ~w3120 & ~w3129;
assign w3131 = w3120 & w3129;
assign w3132 = ~w3130 & ~w3131;
assign w3133 = pi06 & pi33;
assign w3134 = pi09 & pi30;
assign w3135 = pi07 & pi32;
assign w3136 = ~w3134 & ~w3135;
assign w3137 = w3134 & w3135;
assign w3138 = ~w3136 & ~w3137;
assign w3139 = w3133 & ~w3138;
assign w3140 = ~w3133 & w3138;
assign w3141 = ~w3139 & ~w3140;
assign w3142 = w3132 & ~w3141;
assign w3143 = ~w3132 & w3141;
assign w3144 = ~w3142 & ~w3143;
assign w3145 = ~w3111 & w3144;
assign w3146 = w3111 & ~w3144;
assign w3147 = ~w3145 & ~w3146;
assign w3148 = ~w3110 & w3147;
assign w3149 = w3110 & ~w3147;
assign w3150 = ~w3148 & ~w3149;
assign w3151 = w3109 & w3150;
assign w3152 = ~w3109 & ~w3150;
assign w3153 = ~w3151 & ~w3152;
assign w3154 = w3053 & w3153;
assign w3155 = ~w3053 & ~w3153;
assign w3156 = ~w3154 & ~w3155;
assign w3157 = ~w3003 & w3156;
assign w3158 = w3003 & ~w3156;
assign w3159 = ~w3157 & ~w3158;
assign w3160 = ~w2839 & ~w2994;
assign w3161 = (w2691 & w16514) | (w2691 & w16515) | (w16514 & w16515);
assign w3162 = w3159 & w3161;
assign w3163 = ~w3159 & ~w3161;
assign w3164 = ~w3162 & ~w3163;
assign w3165 = ~w3051 & ~w3154;
assign w3166 = (~w3013 & ~w3015) | (~w3013 & w16722) | (~w3015 & w16722);
assign w3167 = ~w3121 & ~w3125;
assign w3168 = ~w3124 & ~w3167;
assign w3169 = ~w3133 & ~w3137;
assign w3170 = ~w3136 & ~w3169;
assign w3171 = w3168 & w3170;
assign w3172 = ~w3168 & ~w3170;
assign w3173 = ~w3171 & ~w3172;
assign w3174 = w3166 & ~w3173;
assign w3175 = ~w3166 & w3173;
assign w3176 = ~w3174 & ~w3175;
assign w3177 = (~w3019 & ~w3021) | (~w3019 & w17074) | (~w3021 & w17074);
assign w3178 = ~w3176 & w3177;
assign w3179 = w3176 & ~w3177;
assign w3180 = ~w3178 & ~w3179;
assign w3181 = pi18 & pi22;
assign w3182 = pi00 & pi40;
assign w3183 = ~w2898 & ~w3182;
assign w3184 = pi02 & pi40;
assign w3185 = w2895 & w3184;
assign w3186 = ~w3183 & ~w3185;
assign w3187 = w3181 & ~w3186;
assign w3188 = ~w3181 & w3186;
assign w3189 = ~w3187 & ~w3188;
assign w3190 = pi07 & pi33;
assign w3191 = pi09 & pi31;
assign w3192 = pi08 & pi32;
assign w3193 = ~w3191 & ~w3192;
assign w3194 = w3191 & w3192;
assign w3195 = ~w3193 & ~w3194;
assign w3196 = w3190 & ~w3195;
assign w3197 = ~w3190 & w3195;
assign w3198 = ~w3196 & ~w3197;
assign w3199 = ~w3189 & ~w3198;
assign w3200 = w3189 & w3198;
assign w3201 = ~w3199 & ~w3200;
assign w3202 = pi04 & pi36;
assign w3203 = pi12 & pi28;
assign w3204 = pi05 & pi35;
assign w3205 = ~w3203 & ~w3204;
assign w3206 = w3203 & w3204;
assign w3207 = ~w3205 & ~w3206;
assign w3208 = w3202 & ~w3207;
assign w3209 = ~w3202 & w3207;
assign w3210 = ~w3208 & ~w3209;
assign w3211 = w3201 & ~w3210;
assign w3212 = ~w3201 & w3210;
assign w3213 = ~w3211 & ~w3212;
assign w3214 = ~w3180 & ~w3213;
assign w3215 = w3180 & w3213;
assign w3216 = ~w3214 & ~w3215;
assign w3217 = ~w3045 & ~w3048;
assign w3218 = ~w3216 & w3217;
assign w3219 = w3216 & ~w3217;
assign w3220 = ~w3218 & ~w3219;
assign w3221 = pi19 & pi21;
assign w3222 = pi01 & pi39;
assign w3223 = ~w3221 & ~w3222;
assign w3224 = w3221 & w3222;
assign w3225 = ~w3223 & ~w3224;
assign w3226 = w3008 & w3225;
assign w3227 = ~w3008 & ~w3225;
assign w3228 = ~w3226 & ~w3227;
assign w3229 = ~w3080 & ~w3084;
assign w3230 = ~w3083 & ~w3229;
assign w3231 = w3228 & w3230;
assign w3232 = ~w3228 & ~w3230;
assign w3233 = ~w3231 & ~w3232;
assign w3234 = (~w3059 & ~w3061) | (~w3059 & w16860) | (~w3061 & w16860);
assign w3235 = (~w3029 & ~w3031) | (~w3029 & w16861) | (~w3031 & w16861);
assign w3236 = ~w3234 & ~w3235;
assign w3237 = w3234 & w3235;
assign w3238 = ~w3236 & ~w3237;
assign w3239 = w3233 & w3238;
assign w3240 = ~w3233 & ~w3238;
assign w3241 = ~w3239 & ~w3240;
assign w3242 = (~w3039 & ~w3041) | (~w3039 & w17075) | (~w3041 & w17075);
assign w3243 = pi03 & pi37;
assign w3244 = pi13 & pi27;
assign w3245 = pi14 & pi26;
assign w3246 = ~w3244 & ~w3245;
assign w3247 = w3244 & w3245;
assign w3248 = ~w3246 & ~w3247;
assign w3249 = w3243 & ~w3248;
assign w3250 = ~w3243 & w3248;
assign w3251 = ~w3249 & ~w3250;
assign w3252 = pi15 & pi25;
assign w3253 = pi16 & pi24;
assign w3254 = pi17 & pi23;
assign w3255 = ~w3253 & ~w3254;
assign w3256 = w3253 & w3254;
assign w3257 = ~w3255 & ~w3256;
assign w3258 = w3252 & ~w3257;
assign w3259 = ~w3252 & w3257;
assign w3260 = ~w3258 & ~w3259;
assign w3261 = ~w3251 & ~w3260;
assign w3262 = w3251 & w3260;
assign w3263 = ~w3261 & ~w3262;
assign w3264 = pi11 & pi29;
assign w3265 = pi06 & pi34;
assign w3266 = pi10 & pi30;
assign w3267 = ~w3265 & ~w3266;
assign w3268 = w3265 & w3266;
assign w3269 = ~w3267 & ~w3268;
assign w3270 = w3264 & ~w3269;
assign w3271 = ~w3264 & w3269;
assign w3272 = ~w3270 & ~w3271;
assign w3273 = w3263 & ~w3272;
assign w3274 = ~w3263 & w3272;
assign w3275 = ~w3273 & ~w3274;
assign w3276 = ~w3242 & w3275;
assign w3277 = w3242 & ~w3275;
assign w3278 = ~w3276 & ~w3277;
assign w3279 = w3241 & w3278;
assign w3280 = ~w3241 & ~w3278;
assign w3281 = ~w3279 & ~w3280;
assign w3282 = w3220 & w3281;
assign w3283 = ~w3220 & ~w3281;
assign w3284 = ~w3282 & ~w3283;
assign w3285 = ~w3145 & ~w3148;
assign w3286 = ~w3069 & ~w3104;
assign w3287 = ~w3092 & ~w3096;
assign w3288 = ~w3095 & ~w3287;
assign w3289 = ~w3112 & ~w3116;
assign w3290 = ~w3115 & ~w3289;
assign w3291 = w3288 & w3290;
assign w3292 = ~w3288 & ~w3290;
assign w3293 = ~w3291 & ~w3292;
assign w3294 = ~w3071 & ~w3075;
assign w3295 = ~w3074 & ~w3294;
assign w3296 = ~w3293 & ~w3295;
assign w3297 = w3293 & w3295;
assign w3298 = ~w3296 & ~w3297;
assign w3299 = (~w3089 & ~w3091) | (~w3089 & w16862) | (~w3091 & w16862);
assign w3300 = (~w3130 & ~w3132) | (~w3130 & w16863) | (~w3132 & w16863);
assign w3301 = ~w3299 & ~w3300;
assign w3302 = w3299 & w3300;
assign w3303 = ~w3301 & ~w3302;
assign w3304 = w3298 & w3303;
assign w3305 = ~w3298 & ~w3303;
assign w3306 = ~w3304 & ~w3305;
assign w3307 = ~w3286 & w3306;
assign w3308 = w3286 & ~w3306;
assign w3309 = ~w3307 & ~w3308;
assign w3310 = ~w3285 & w3309;
assign w3311 = w3285 & ~w3309;
assign w3312 = ~w3310 & ~w3311;
assign w3313 = ~w3107 & ~w3151;
assign w3314 = w3312 & ~w3313;
assign w3315 = ~w3312 & w3313;
assign w3316 = ~w3314 & ~w3315;
assign w3317 = w3284 & w3316;
assign w3318 = ~w3284 & ~w3316;
assign w3319 = ~w3317 & ~w3318;
assign w3320 = ~w3165 & w3319;
assign w3321 = w3165 & ~w3319;
assign w3322 = ~w3320 & ~w3321;
assign w3323 = ~w3157 & ~w3161;
assign w3324 = ~w3158 & ~w3323;
assign w3325 = w3322 & w3324;
assign w3326 = ~w3322 & ~w3324;
assign w3327 = ~w3325 & ~w3326;
assign w3328 = ~w3314 & ~w3317;
assign w3329 = ~w3276 & ~w3279;
assign w3330 = ~w3179 & ~w3215;
assign w3331 = ~w3252 & ~w3256;
assign w3332 = ~w3255 & ~w3331;
assign w3333 = w3181 & ~w3183;
assign w3334 = ~w3185 & ~w3333;
assign w3335 = w3332 & ~w3334;
assign w3336 = ~w3332 & w3334;
assign w3337 = ~w3335 & ~w3336;
assign w3338 = ~w3243 & ~w3247;
assign w3339 = ~w3246 & ~w3338;
assign w3340 = ~w3337 & ~w3339;
assign w3341 = w3337 & w3339;
assign w3342 = ~w3340 & ~w3341;
assign w3343 = (~w3199 & ~w3201) | (~w3199 & w16864) | (~w3201 & w16864);
assign w3344 = ~w3342 & w3343;
assign w3345 = w3342 & ~w3343;
assign w3346 = ~w3344 & ~w3345;
assign w3347 = pi40 & w964;
assign w3348 = pi01 & pi40;
assign w3349 = ~pi21 & ~w3348;
assign w3350 = ~w3347 & ~w3349;
assign w3351 = ~w3190 & ~w3194;
assign w3352 = ~w3193 & ~w3351;
assign w3353 = w3350 & w3352;
assign w3354 = ~w3350 & ~w3352;
assign w3355 = ~w3353 & ~w3354;
assign w3356 = ~w3264 & ~w3268;
assign w3357 = ~w3267 & ~w3356;
assign w3358 = w3355 & w3357;
assign w3359 = ~w3355 & ~w3357;
assign w3360 = ~w3358 & ~w3359;
assign w3361 = w3346 & w3360;
assign w3362 = ~w3346 & ~w3360;
assign w3363 = ~w3361 & ~w3362;
assign w3364 = ~w3330 & w3363;
assign w3365 = w3330 & ~w3363;
assign w3366 = ~w3364 & ~w3365;
assign w3367 = w3329 & ~w3366;
assign w3368 = ~w3329 & w3366;
assign w3369 = ~w3367 & ~w3368;
assign w3370 = ~w3219 & ~w3282;
assign w3371 = ~w3369 & w3370;
assign w3372 = w3369 & ~w3370;
assign w3373 = ~w3371 & ~w3372;
assign w3374 = (~w3261 & ~w3263) | (~w3261 & w16865) | (~w3263 & w16865);
assign w3375 = (~w3171 & ~w3173) | (~w3171 & w16723) | (~w3173 & w16723);
assign w3376 = (~w3291 & ~w3293) | (~w3291 & w16724) | (~w3293 & w16724);
assign w3377 = ~w3375 & ~w3376;
assign w3378 = w3375 & w3376;
assign w3379 = ~w3377 & ~w3378;
assign w3380 = w3374 & ~w3379;
assign w3381 = ~w3374 & w3379;
assign w3382 = ~w3380 & ~w3381;
assign w3383 = ~w3202 & ~w3206;
assign w3384 = ~w3205 & ~w3383;
assign w3385 = pi00 & pi41;
assign w3386 = pi02 & pi39;
assign w3387 = ~w3385 & ~w3386;
assign w3388 = pi02 & pi41;
assign w3389 = w3012 & w3388;
assign w3390 = ~w3387 & ~w3389;
assign w3391 = w3224 & ~w3390;
assign w3392 = ~w3224 & w3390;
assign w3393 = ~w3391 & ~w3392;
assign w3394 = w3384 & ~w3393;
assign w3395 = ~w3384 & w3393;
assign w3396 = ~w3394 & ~w3395;
assign w3397 = pi03 & pi38;
assign w3398 = pi13 & pi28;
assign w3399 = pi15 & pi26;
assign w3400 = ~w3398 & ~w3399;
assign w3401 = w3398 & w3399;
assign w3402 = ~w3400 & ~w3401;
assign w3403 = w3397 & ~w3402;
assign w3404 = ~w3397 & w3402;
assign w3405 = ~w3403 & ~w3404;
assign w3406 = ~w3396 & w3405;
assign w3407 = w3396 & ~w3405;
assign w3408 = ~w3406 & ~w3407;
assign w3409 = (~w3301 & ~w3303) | (~w3301 & w17076) | (~w3303 & w17076);
assign w3410 = w3408 & ~w3409;
assign w3411 = ~w3408 & w3409;
assign w3412 = ~w3410 & ~w3411;
assign w3413 = ~w3382 & ~w3412;
assign w3414 = w3382 & w3412;
assign w3415 = ~w3413 & ~w3414;
assign w3416 = (~w3307 & w3285) | (~w3307 & w16725) | (w3285 & w16725);
assign w3417 = (~w3226 & ~w3228) | (~w3226 & w17077) | (~w3228 & w17077);
assign w3418 = pi08 & pi33;
assign w3419 = pi20 & pi21;
assign w3420 = pi19 & pi22;
assign w3421 = ~w3419 & ~w3420;
assign w3422 = w3419 & w3420;
assign w3423 = ~w3421 & ~w3422;
assign w3424 = w3418 & ~w3423;
assign w3425 = ~w3418 & w3423;
assign w3426 = ~w3424 & ~w3425;
assign w3427 = pi05 & pi36;
assign w3428 = pi06 & pi35;
assign w3429 = pi11 & pi30;
assign w3430 = ~w3428 & ~w3429;
assign w3431 = w3428 & w3429;
assign w3432 = ~w3430 & ~w3431;
assign w3433 = w3427 & ~w3432;
assign w3434 = ~w3427 & w3432;
assign w3435 = ~w3433 & ~w3434;
assign w3436 = ~w3426 & ~w3435;
assign w3437 = w3426 & w3435;
assign w3438 = ~w3436 & ~w3437;
assign w3439 = w3417 & ~w3438;
assign w3440 = ~w3417 & w3438;
assign w3441 = ~w3439 & ~w3440;
assign w3442 = (~w3236 & ~w3238) | (~w3236 & w16726) | (~w3238 & w16726);
assign w3443 = ~w3441 & w3442;
assign w3444 = w3441 & ~w3442;
assign w3445 = ~w3443 & ~w3444;
assign w3446 = pi14 & pi27;
assign w3447 = pi04 & pi37;
assign w3448 = pi12 & pi29;
assign w3449 = ~w3447 & ~w3448;
assign w3450 = w3447 & w3448;
assign w3451 = ~w3449 & ~w3450;
assign w3452 = w3446 & ~w3451;
assign w3453 = ~w3446 & w3451;
assign w3454 = ~w3452 & ~w3453;
assign w3455 = pi16 & pi25;
assign w3456 = pi17 & pi24;
assign w3457 = pi18 & pi23;
assign w3458 = ~w3456 & ~w3457;
assign w3459 = w3456 & w3457;
assign w3460 = ~w3458 & ~w3459;
assign w3461 = w3455 & ~w3460;
assign w3462 = ~w3455 & w3460;
assign w3463 = ~w3461 & ~w3462;
assign w3464 = ~w3454 & ~w3463;
assign w3465 = w3454 & w3463;
assign w3466 = ~w3464 & ~w3465;
assign w3467 = pi10 & pi31;
assign w3468 = pi09 & pi32;
assign w3469 = pi07 & pi34;
assign w3470 = ~w3468 & ~w3469;
assign w3471 = w3468 & w3469;
assign w3472 = ~w3470 & ~w3471;
assign w3473 = w3467 & ~w3472;
assign w3474 = ~w3467 & w3472;
assign w3475 = ~w3473 & ~w3474;
assign w3476 = w3466 & ~w3475;
assign w3477 = ~w3466 & w3475;
assign w3478 = ~w3476 & ~w3477;
assign w3479 = ~w3445 & ~w3478;
assign w3480 = w3445 & w3478;
assign w3481 = ~w3479 & ~w3480;
assign w3482 = ~w3416 & w3481;
assign w3483 = w3416 & ~w3481;
assign w3484 = ~w3482 & ~w3483;
assign w3485 = w3415 & w3484;
assign w3486 = ~w3415 & ~w3484;
assign w3487 = ~w3485 & ~w3486;
assign w3488 = w3373 & w3487;
assign w3489 = ~w3373 & ~w3487;
assign w3490 = ~w3488 & ~w3489;
assign w3491 = w3328 & ~w3490;
assign w3492 = ~w3328 & w3490;
assign w3493 = ~w3491 & ~w3492;
assign w3494 = ~w3158 & ~w3321;
assign w3495 = (w3494 & w3161) | (w3494 & w16516) | (w3161 & w16516);
assign w3496 = ~w3320 & ~w3495;
assign w3497 = w3493 & w3496;
assign w3498 = ~w3493 & ~w3496;
assign w3499 = ~w3497 & ~w3498;
assign w3500 = ~w3320 & ~w3492;
assign w3501 = (~w3491 & w3495) | (~w3491 & w16517) | (w3495 & w16517);
assign w3502 = ~w3372 & ~w3488;
assign w3503 = ~w3482 & ~w3485;
assign w3504 = ~w3410 & ~w3414;
assign w3505 = ~w3464 & ~w3476;
assign w3506 = ~w3335 & ~w3341;
assign w3507 = (~w3394 & ~w3396) | (~w3394 & w17078) | (~w3396 & w17078);
assign w3508 = ~w3506 & ~w3507;
assign w3509 = w3506 & w3507;
assign w3510 = ~w3508 & ~w3509;
assign w3511 = w3505 & ~w3510;
assign w3512 = ~w3505 & w3510;
assign w3513 = ~w3511 & ~w3512;
assign w3514 = (~w3444 & ~w3445) | (~w3444 & w17079) | (~w3445 & w17079);
assign w3515 = ~w3513 & w3514;
assign w3516 = w3513 & ~w3514;
assign w3517 = ~w3515 & ~w3516;
assign w3518 = ~w3504 & w3517;
assign w3519 = w3504 & ~w3517;
assign w3520 = ~w3518 & ~w3519;
assign w3521 = ~w3503 & w3520;
assign w3522 = w3503 & ~w3520;
assign w3523 = ~w3521 & ~w3522;
assign w3524 = (~w3364 & ~w3366) | (~w3364 & w16727) | (~w3366 & w16727);
assign w3525 = ~w3467 & ~w3471;
assign w3526 = ~w3470 & ~w3525;
assign w3527 = pi06 & pi36;
assign w3528 = pi07 & pi35;
assign w3529 = pi11 & pi31;
assign w3530 = ~w3528 & ~w3529;
assign w3531 = w3528 & w3529;
assign w3532 = ~w3530 & ~w3531;
assign w3533 = w3527 & ~w3532;
assign w3534 = ~w3527 & w3532;
assign w3535 = ~w3533 & ~w3534;
assign w3536 = w3526 & ~w3535;
assign w3537 = ~w3526 & w3535;
assign w3538 = ~w3536 & ~w3537;
assign w3539 = pi10 & pi32;
assign w3540 = pi09 & pi33;
assign w3541 = pi08 & pi34;
assign w3542 = ~w3540 & ~w3541;
assign w3543 = w3540 & w3541;
assign w3544 = ~w3542 & ~w3543;
assign w3545 = w3539 & ~w3544;
assign w3546 = ~w3539 & w3544;
assign w3547 = ~w3545 & ~w3546;
assign w3548 = w3538 & ~w3547;
assign w3549 = ~w3538 & w3547;
assign w3550 = ~w3548 & ~w3549;
assign w3551 = (w3550 & w3381) | (w3550 & w16728) | (w3381 & w16728);
assign w3552 = ~w3381 & w16729;
assign w3553 = ~w3551 & ~w3552;
assign w3554 = pi03 & pi39;
assign w3555 = pi16 & pi26;
assign w3556 = ~w3554 & ~w3555;
assign w3557 = w3554 & w3555;
assign w3558 = ~w3556 & ~w3557;
assign w3559 = w3184 & ~w3558;
assign w3560 = ~w3184 & w3558;
assign w3561 = ~w3559 & ~w3560;
assign w3562 = pi17 & pi25;
assign w3563 = pi18 & pi24;
assign w3564 = pi19 & pi23;
assign w3565 = ~w3563 & ~w3564;
assign w3566 = w3563 & w3564;
assign w3567 = ~w3565 & ~w3566;
assign w3568 = w3562 & ~w3567;
assign w3569 = ~w3562 & w3567;
assign w3570 = ~w3568 & ~w3569;
assign w3571 = ~w3561 & ~w3570;
assign w3572 = w3561 & w3570;
assign w3573 = ~w3571 & ~w3572;
assign w3574 = pi15 & pi27;
assign w3575 = pi04 & pi38;
assign w3576 = pi14 & pi28;
assign w3577 = ~w3575 & ~w3576;
assign w3578 = w3575 & w3576;
assign w3579 = ~w3577 & ~w3578;
assign w3580 = w3574 & ~w3579;
assign w3581 = ~w3574 & w3579;
assign w3582 = ~w3580 & ~w3581;
assign w3583 = w3573 & ~w3582;
assign w3584 = ~w3573 & w3582;
assign w3585 = ~w3583 & ~w3584;
assign w3586 = w3553 & w3585;
assign w3587 = ~w3553 & ~w3585;
assign w3588 = ~w3586 & ~w3587;
assign w3589 = ~w3524 & w3588;
assign w3590 = w3524 & ~w3588;
assign w3591 = ~w3589 & ~w3590;
assign w3592 = (~w3353 & ~w3355) | (~w3353 & w16866) | (~w3355 & w16866);
assign w3593 = pi00 & pi42;
assign w3594 = w3347 & w3593;
assign w3595 = ~w3347 & ~w3593;
assign w3596 = ~w3594 & ~w3595;
assign w3597 = pi20 & pi22;
assign w3598 = pi01 & pi41;
assign w3599 = ~w3597 & ~w3598;
assign w3600 = w3597 & w3598;
assign w3601 = ~w3599 & ~w3600;
assign w3602 = w3596 & w3601;
assign w3603 = ~w3596 & ~w3601;
assign w3604 = ~w3602 & ~w3603;
assign w3605 = pi13 & pi29;
assign w3606 = pi05 & pi37;
assign w3607 = pi12 & pi30;
assign w3608 = ~w3606 & ~w3607;
assign w3609 = w3606 & w3607;
assign w3610 = ~w3608 & ~w3609;
assign w3611 = w3605 & ~w3610;
assign w3612 = ~w3605 & w3610;
assign w3613 = ~w3611 & ~w3612;
assign w3614 = w3604 & ~w3613;
assign w3615 = ~w3604 & w3613;
assign w3616 = ~w3614 & ~w3615;
assign w3617 = w3592 & ~w3616;
assign w3618 = ~w3592 & w3616;
assign w3619 = ~w3617 & ~w3618;
assign w3620 = (~w3345 & ~w3346) | (~w3345 & w16730) | (~w3346 & w16730);
assign w3621 = ~w3619 & w3620;
assign w3622 = w3619 & ~w3620;
assign w3623 = ~w3621 & ~w3622;
assign w3624 = ~w3446 & ~w3450;
assign w3625 = ~w3449 & ~w3624;
assign w3626 = ~w3418 & ~w3422;
assign w3627 = ~w3421 & ~w3626;
assign w3628 = w3625 & w3627;
assign w3629 = ~w3625 & ~w3627;
assign w3630 = ~w3628 & ~w3629;
assign w3631 = ~w3427 & ~w3431;
assign w3632 = ~w3430 & ~w3631;
assign w3633 = ~w3630 & ~w3632;
assign w3634 = w3630 & w3632;
assign w3635 = ~w3633 & ~w3634;
assign w3636 = (~w3436 & ~w3438) | (~w3436 & w17080) | (~w3438 & w17080);
assign w3637 = ~w3635 & w3636;
assign w3638 = w3635 & ~w3636;
assign w3639 = ~w3637 & ~w3638;
assign w3640 = ~w3397 & ~w3401;
assign w3641 = ~w3400 & ~w3640;
assign w3642 = ~w3455 & ~w3459;
assign w3643 = ~w3458 & ~w3642;
assign w3644 = w3641 & w3643;
assign w3645 = ~w3641 & ~w3643;
assign w3646 = ~w3644 & ~w3645;
assign w3647 = w3224 & ~w3387;
assign w3648 = ~w3389 & ~w3647;
assign w3649 = ~w3646 & w3648;
assign w3650 = w3646 & ~w3648;
assign w3651 = ~w3649 & ~w3650;
assign w3652 = w3639 & w3651;
assign w3653 = ~w3639 & ~w3651;
assign w3654 = ~w3652 & ~w3653;
assign w3655 = w3623 & w3654;
assign w3656 = ~w3623 & ~w3654;
assign w3657 = ~w3655 & ~w3656;
assign w3658 = w3591 & w3657;
assign w3659 = ~w3591 & ~w3657;
assign w3660 = ~w3658 & ~w3659;
assign w3661 = ~w3523 & ~w3660;
assign w3662 = w3523 & w3660;
assign w3663 = ~w3661 & ~w3662;
assign w3664 = w3502 & ~w3663;
assign w3665 = ~w3502 & w3663;
assign w3666 = ~w3664 & ~w3665;
assign w3667 = w3501 & ~w3666;
assign w3668 = ~w3501 & w3666;
assign w3669 = ~w3667 & ~w3668;
assign w3670 = (~w3495 & w16518) | (~w3495 & w16519) | (w16518 & w16519);
assign w3671 = ~w3664 & ~w3670;
assign w3672 = ~w3521 & ~w3662;
assign w3673 = ~w3516 & ~w3518;
assign w3674 = ~w3508 & ~w3512;
assign w3675 = pi04 & pi39;
assign w3676 = pi00 & pi43;
assign w3677 = pi03 & pi40;
assign w3678 = ~w3676 & ~w3677;
assign w3679 = w3676 & w3677;
assign w3680 = ~w3678 & ~w3679;
assign w3681 = w3675 & ~w3680;
assign w3682 = ~w3675 & w3680;
assign w3683 = ~w3681 & ~w3682;
assign w3684 = pi15 & pi28;
assign w3685 = pi16 & pi27;
assign w3686 = ~w3684 & ~w3685;
assign w3687 = w3684 & w3685;
assign w3688 = ~w3686 & ~w3687;
assign w3689 = w1755 & ~w3688;
assign w3690 = ~w1755 & w3688;
assign w3691 = ~w3689 & ~w3690;
assign w3692 = ~w3683 & ~w3691;
assign w3693 = w3683 & w3691;
assign w3694 = ~w3692 & ~w3693;
assign w3695 = pi17 & pi26;
assign w3696 = pi19 & pi24;
assign w3697 = pi18 & pi25;
assign w3698 = ~w3696 & ~w3697;
assign w3699 = w3696 & w3697;
assign w3700 = ~w3698 & ~w3699;
assign w3701 = w3695 & ~w3700;
assign w3702 = ~w3695 & w3700;
assign w3703 = ~w3701 & ~w3702;
assign w3704 = w3694 & ~w3703;
assign w3705 = ~w3694 & w3703;
assign w3706 = ~w3704 & ~w3705;
assign w3707 = pi09 & pi34;
assign w3708 = pi21 & pi22;
assign w3709 = pi20 & pi23;
assign w3710 = ~w3708 & ~w3709;
assign w3711 = w3708 & w3709;
assign w3712 = ~w3710 & ~w3711;
assign w3713 = w3707 & ~w3712;
assign w3714 = ~w3707 & w3712;
assign w3715 = ~w3713 & ~w3714;
assign w3716 = pi07 & pi36;
assign w3717 = pi10 & pi33;
assign w3718 = pi08 & pi35;
assign w3719 = ~w3717 & ~w3718;
assign w3720 = w3717 & w3718;
assign w3721 = ~w3719 & ~w3720;
assign w3722 = w3716 & ~w3721;
assign w3723 = ~w3716 & w3721;
assign w3724 = ~w3722 & ~w3723;
assign w3725 = ~w3715 & ~w3724;
assign w3726 = w3715 & w3724;
assign w3727 = ~w3725 & ~w3726;
assign w3728 = pi05 & pi38;
assign w3729 = pi13 & pi30;
assign w3730 = ~w3728 & ~w3729;
assign w3731 = w3728 & w3729;
assign w3732 = ~w3730 & ~w3731;
assign w3733 = w3388 & ~w3732;
assign w3734 = ~w3388 & w3732;
assign w3735 = ~w3733 & ~w3734;
assign w3736 = w3727 & ~w3735;
assign w3737 = ~w3727 & w3735;
assign w3738 = ~w3736 & ~w3737;
assign w3739 = w3706 & w3738;
assign w3740 = ~w3706 & ~w3738;
assign w3741 = ~w3739 & ~w3740;
assign w3742 = ~w3674 & w3741;
assign w3743 = w3674 & ~w3741;
assign w3744 = ~w3742 & ~w3743;
assign w3745 = ~w3673 & w3744;
assign w3746 = w3673 & ~w3744;
assign w3747 = ~w3745 & ~w3746;
assign w3748 = (~w3614 & ~w3616) | (~w3614 & w16867) | (~w3616 & w16867);
assign w3749 = ~w3574 & ~w3578;
assign w3750 = ~w3577 & ~w3749;
assign w3751 = ~w3527 & ~w3531;
assign w3752 = ~w3530 & ~w3751;
assign w3753 = w3750 & w3752;
assign w3754 = ~w3750 & ~w3752;
assign w3755 = ~w3753 & ~w3754;
assign w3756 = ~w3562 & ~w3566;
assign w3757 = ~w3565 & ~w3756;
assign w3758 = ~w3755 & ~w3757;
assign w3759 = w3755 & w3757;
assign w3760 = ~w3758 & ~w3759;
assign w3761 = (~w3594 & ~w3596) | (~w3594 & w16868) | (~w3596 & w16868);
assign w3762 = ~w3184 & ~w3557;
assign w3763 = ~w3556 & ~w3762;
assign w3764 = ~w3605 & ~w3609;
assign w3765 = ~w3608 & ~w3764;
assign w3766 = w3763 & w3765;
assign w3767 = ~w3763 & ~w3765;
assign w3768 = ~w3766 & ~w3767;
assign w3769 = w3761 & ~w3768;
assign w3770 = ~w3761 & w3768;
assign w3771 = ~w3769 & ~w3770;
assign w3772 = w3760 & w3771;
assign w3773 = ~w3760 & ~w3771;
assign w3774 = ~w3772 & ~w3773;
assign w3775 = ~w3748 & w3774;
assign w3776 = w3748 & ~w3774;
assign w3777 = ~w3775 & ~w3776;
assign w3778 = (~w3644 & ~w3646) | (~w3644 & w17081) | (~w3646 & w17081);
assign w3779 = (~w3628 & ~w3630) | (~w3628 & w16731) | (~w3630 & w16731);
assign w3780 = pi12 & pi31;
assign w3781 = pi11 & pi32;
assign w3782 = pi06 & pi37;
assign w3783 = ~w3781 & ~w3782;
assign w3784 = w3781 & w3782;
assign w3785 = ~w3783 & ~w3784;
assign w3786 = w3780 & ~w3785;
assign w3787 = ~w3780 & w3785;
assign w3788 = ~w3786 & ~w3787;
assign w3789 = ~w3779 & ~w3788;
assign w3790 = w3779 & w3788;
assign w3791 = ~w3789 & ~w3790;
assign w3792 = w3778 & ~w3791;
assign w3793 = ~w3778 & w3791;
assign w3794 = ~w3792 & ~w3793;
assign w3795 = ~w3638 & ~w3652;
assign w3796 = ~w3794 & w3795;
assign w3797 = w3794 & ~w3795;
assign w3798 = ~w3796 & ~w3797;
assign w3799 = w3777 & w3798;
assign w3800 = ~w3777 & ~w3798;
assign w3801 = ~w3799 & ~w3800;
assign w3802 = w3747 & w3801;
assign w3803 = ~w3747 & ~w3801;
assign w3804 = ~w3802 & ~w3803;
assign w3805 = ~w3589 & ~w3658;
assign w3806 = (~w3622 & ~w3623) | (~w3622 & w17082) | (~w3623 & w17082);
assign w3807 = (~w3551 & ~w3553) | (~w3551 & w16869) | (~w3553 & w16869);
assign w3808 = ~w3571 & ~w3583;
assign w3809 = (~w3536 & ~w3538) | (~w3536 & w17083) | (~w3538 & w17083);
assign w3810 = ~pi42 & w3600;
assign w3811 = pi42 & w1056;
assign w3812 = pi01 & pi42;
assign w3813 = ~pi22 & ~w3812;
assign w3814 = ~w3811 & ~w3813;
assign w3815 = ~w3600 & ~w3814;
assign w3816 = ~w3810 & ~w3815;
assign w3817 = ~w3539 & ~w3543;
assign w3818 = ~w3542 & ~w3817;
assign w3819 = w3816 & w3818;
assign w3820 = ~w3816 & ~w3818;
assign w3821 = ~w3819 & ~w3820;
assign w3822 = ~w3809 & w3821;
assign w3823 = w3809 & ~w3821;
assign w3824 = ~w3822 & ~w3823;
assign w3825 = ~w3808 & w3824;
assign w3826 = w3808 & ~w3824;
assign w3827 = ~w3825 & ~w3826;
assign w3828 = ~w3807 & w3827;
assign w3829 = w3807 & ~w3827;
assign w3830 = ~w3828 & ~w3829;
assign w3831 = ~w3806 & w3830;
assign w3832 = w3806 & ~w3830;
assign w3833 = ~w3831 & ~w3832;
assign w3834 = ~w3805 & w3833;
assign w3835 = w3805 & ~w3833;
assign w3836 = ~w3834 & ~w3835;
assign w3837 = w3804 & w3836;
assign w3838 = ~w3804 & ~w3836;
assign w3839 = ~w3837 & ~w3838;
assign w3840 = ~w3672 & w3839;
assign w3841 = w3672 & ~w3839;
assign w3842 = ~w3840 & ~w3841;
assign w3843 = w3671 & w3842;
assign w3844 = ~w3671 & ~w3842;
assign w3845 = ~w3843 & ~w3844;
assign w3846 = ~w3834 & ~w3837;
assign w3847 = ~w3745 & ~w3802;
assign w3848 = ~w3797 & ~w3799;
assign w3849 = ~w3739 & ~w3742;
assign w3850 = ~w3675 & ~w3679;
assign w3851 = ~w3678 & ~w3850;
assign w3852 = ~w3388 & ~w3731;
assign w3853 = ~w3730 & ~w3852;
assign w3854 = w3851 & w3853;
assign w3855 = ~w3851 & ~w3853;
assign w3856 = ~w3854 & ~w3855;
assign w3857 = ~w3695 & ~w3699;
assign w3858 = ~w3698 & ~w3857;
assign w3859 = ~w3856 & ~w3858;
assign w3860 = w3856 & w3858;
assign w3861 = ~w3859 & ~w3860;
assign w3862 = ~w3725 & ~w3736;
assign w3863 = ~w3692 & ~w3704;
assign w3864 = ~w3862 & ~w3863;
assign w3865 = w3862 & w3863;
assign w3866 = ~w3864 & ~w3865;
assign w3867 = w3861 & w3866;
assign w3868 = ~w3861 & ~w3866;
assign w3869 = ~w3867 & ~w3868;
assign w3870 = ~w3849 & w3869;
assign w3871 = w3849 & ~w3869;
assign w3872 = ~w3870 & ~w3871;
assign w3873 = ~w3848 & w3872;
assign w3874 = w3848 & ~w3872;
assign w3875 = ~w3873 & ~w3874;
assign w3876 = ~w3847 & w3875;
assign w3877 = w3847 & ~w3875;
assign w3878 = ~w3876 & ~w3877;
assign w3879 = (~w3828 & ~w3830) | (~w3828 & w17084) | (~w3830 & w17084);
assign w3880 = ~w3822 & ~w3825;
assign w3881 = pi03 & pi41;
assign w3882 = pi15 & pi29;
assign w3883 = pi17 & pi27;
assign w3884 = ~w3882 & ~w3883;
assign w3885 = w3882 & w3883;
assign w3886 = ~w3884 & ~w3885;
assign w3887 = w3881 & ~w3886;
assign w3888 = ~w3881 & w3886;
assign w3889 = ~w3887 & ~w3888;
assign w3890 = pi18 & pi26;
assign w3891 = pi19 & pi25;
assign w3892 = pi20 & pi24;
assign w3893 = ~w3891 & ~w3892;
assign w3894 = w3891 & w3892;
assign w3895 = ~w3893 & ~w3894;
assign w3896 = w3890 & ~w3895;
assign w3897 = ~w3890 & w3895;
assign w3898 = ~w3896 & ~w3897;
assign w3899 = ~w3889 & ~w3898;
assign w3900 = w3889 & w3898;
assign w3901 = ~w3899 & ~w3900;
assign w3902 = pi06 & pi38;
assign w3903 = pi11 & pi33;
assign w3904 = pi07 & pi37;
assign w3905 = ~w3903 & ~w3904;
assign w3906 = w3903 & w3904;
assign w3907 = ~w3905 & ~w3906;
assign w3908 = w3902 & ~w3907;
assign w3909 = ~w3902 & w3907;
assign w3910 = ~w3908 & ~w3909;
assign w3911 = w3901 & ~w3910;
assign w3912 = ~w3901 & w3910;
assign w3913 = ~w3911 & ~w3912;
assign w3914 = pi08 & pi36;
assign w3915 = pi10 & pi34;
assign w3916 = pi09 & pi35;
assign w3917 = ~w3915 & ~w3916;
assign w3918 = pi10 & pi35;
assign w3919 = w3707 & w3918;
assign w3920 = ~w3917 & ~w3919;
assign w3921 = w3914 & ~w3920;
assign w3922 = ~w3914 & w3920;
assign w3923 = ~w3921 & ~w3922;
assign w3924 = pi16 & pi28;
assign w3925 = pi04 & pi40;
assign w3926 = pi14 & pi30;
assign w3927 = ~w3925 & ~w3926;
assign w3928 = w3925 & w3926;
assign w3929 = ~w3927 & ~w3928;
assign w3930 = w3924 & ~w3929;
assign w3931 = ~w3924 & w3929;
assign w3932 = ~w3930 & ~w3931;
assign w3933 = ~w3923 & ~w3932;
assign w3934 = w3923 & w3932;
assign w3935 = ~w3933 & ~w3934;
assign w3936 = pi05 & pi39;
assign w3937 = pi12 & pi32;
assign w3938 = pi13 & pi31;
assign w3939 = ~w3937 & ~w3938;
assign w3940 = w3937 & w3938;
assign w3941 = ~w3939 & ~w3940;
assign w3942 = w3936 & ~w3941;
assign w3943 = ~w3936 & w3941;
assign w3944 = ~w3942 & ~w3943;
assign w3945 = w3935 & ~w3944;
assign w3946 = ~w3935 & w3944;
assign w3947 = ~w3945 & ~w3946;
assign w3948 = w3913 & w3947;
assign w3949 = ~w3913 & ~w3947;
assign w3950 = ~w3948 & ~w3949;
assign w3951 = ~w3880 & w3950;
assign w3952 = w3880 & ~w3950;
assign w3953 = ~w3951 & ~w3952;
assign w3954 = ~w3879 & w3953;
assign w3955 = w3879 & ~w3953;
assign w3956 = ~w3954 & ~w3955;
assign w3957 = ~w1755 & ~w3687;
assign w3958 = ~w3686 & ~w3957;
assign w3959 = ~w3780 & ~w3784;
assign w3960 = ~w3783 & ~w3959;
assign w3961 = w3958 & w3960;
assign w3962 = ~w3958 & ~w3960;
assign w3963 = ~w3961 & ~w3962;
assign w3964 = pi00 & pi44;
assign w3965 = pi02 & pi42;
assign w3966 = ~w3964 & ~w3965;
assign w3967 = pi02 & pi44;
assign w3968 = w3593 & w3967;
assign w3969 = ~w3966 & ~w3968;
assign w3970 = w3811 & ~w3969;
assign w3971 = ~w3811 & w3969;
assign w3972 = ~w3970 & ~w3971;
assign w3973 = ~w3963 & w3972;
assign w3974 = w3963 & ~w3972;
assign w3975 = ~w3973 & ~w3974;
assign w3976 = pi21 & pi23;
assign w3977 = pi01 & pi43;
assign w3978 = ~w3976 & ~w3977;
assign w3979 = w3976 & w3977;
assign w3980 = ~w3978 & ~w3979;
assign w3981 = ~w3707 & ~w3711;
assign w3982 = ~w3710 & ~w3981;
assign w3983 = w3980 & w3982;
assign w3984 = ~w3980 & ~w3982;
assign w3985 = ~w3983 & ~w3984;
assign w3986 = ~w3716 & ~w3720;
assign w3987 = ~w3719 & ~w3986;
assign w3988 = w3985 & w3987;
assign w3989 = ~w3985 & ~w3987;
assign w3990 = ~w3988 & ~w3989;
assign w3991 = w3975 & w3990;
assign w3992 = ~w3975 & ~w3990;
assign w3993 = ~w3991 & ~w3992;
assign w3994 = (~w3789 & ~w3791) | (~w3789 & w16870) | (~w3791 & w16870);
assign w3995 = ~w3993 & w3994;
assign w3996 = w3993 & ~w3994;
assign w3997 = ~w3995 & ~w3996;
assign w3998 = (~w3772 & ~w3774) | (~w3772 & w16871) | (~w3774 & w16871);
assign w3999 = ~w3753 & ~w3759;
assign w4000 = (~w3766 & ~w3768) | (~w3766 & w16872) | (~w3768 & w16872);
assign w4001 = (~w3810 & ~w3816) | (~w3810 & w17085) | (~w3816 & w17085);
assign w4002 = ~w4000 & ~w4001;
assign w4003 = w4000 & w4001;
assign w4004 = ~w4002 & ~w4003;
assign w4005 = w3999 & ~w4004;
assign w4006 = ~w3999 & w4004;
assign w4007 = ~w4005 & ~w4006;
assign w4008 = ~w3998 & w4007;
assign w4009 = w3998 & ~w4007;
assign w4010 = ~w4008 & ~w4009;
assign w4011 = ~w3997 & ~w4010;
assign w4012 = w3997 & w4010;
assign w4013 = ~w4011 & ~w4012;
assign w4014 = w3956 & w4013;
assign w4015 = ~w3956 & ~w4013;
assign w4016 = ~w4014 & ~w4015;
assign w4017 = w3878 & w4016;
assign w4018 = ~w3878 & ~w4016;
assign w4019 = ~w4017 & ~w4018;
assign w4020 = ~w3846 & w4019;
assign w4021 = w3846 & ~w4019;
assign w4022 = ~w4020 & ~w4021;
assign w4023 = ~w3664 & ~w3841;
assign w4024 = ~w3670 & w4023;
assign w4025 = ~w3840 & ~w4024;
assign w4026 = w4022 & w4025;
assign w4027 = ~w4022 & ~w4025;
assign w4028 = ~w4026 & ~w4027;
assign w4029 = ~w3840 & ~w4020;
assign w4030 = (~w3670 & w16521) | (~w3670 & w16522) | (w16521 & w16522);
assign w4031 = ~w3876 & ~w4017;
assign w4032 = (~w3983 & ~w3985) | (~w3983 & w17086) | (~w3985 & w17086);
assign w4033 = (~w3961 & ~w3963) | (~w3961 & w16732) | (~w3963 & w16732);
assign w4034 = (~w3854 & ~w3856) | (~w3854 & w16733) | (~w3856 & w16733);
assign w4035 = ~w4033 & ~w4034;
assign w4036 = w4033 & w4034;
assign w4037 = ~w4035 & ~w4036;
assign w4038 = w4032 & ~w4037;
assign w4039 = ~w4032 & w4037;
assign w4040 = ~w4038 & ~w4039;
assign w4041 = ~w3991 & ~w3996;
assign w4042 = ~w4040 & w4041;
assign w4043 = w4040 & ~w4041;
assign w4044 = ~w4042 & ~w4043;
assign w4045 = ~w3902 & ~w3906;
assign w4046 = ~w3905 & ~w4045;
assign w4047 = ~w3924 & ~w3928;
assign w4048 = ~w3927 & ~w4047;
assign w4049 = w4046 & w4048;
assign w4050 = ~w4046 & ~w4048;
assign w4051 = ~w4049 & ~w4050;
assign w4052 = ~w3936 & ~w3940;
assign w4053 = ~w3939 & ~w4052;
assign w4054 = ~w4051 & ~w4053;
assign w4055 = w4051 & w4053;
assign w4056 = ~w4054 & ~w4055;
assign w4057 = (~w3933 & ~w3935) | (~w3933 & w16873) | (~w3935 & w16873);
assign w4058 = (~w3899 & ~w3901) | (~w3899 & w16874) | (~w3901 & w16874);
assign w4059 = ~w4057 & ~w4058;
assign w4060 = w4057 & w4058;
assign w4061 = ~w4059 & ~w4060;
assign w4062 = w4056 & w4061;
assign w4063 = ~w4056 & ~w4061;
assign w4064 = ~w4062 & ~w4063;
assign w4065 = w4044 & w4064;
assign w4066 = ~w4044 & ~w4064;
assign w4067 = ~w4065 & ~w4066;
assign w4068 = ~w3870 & ~w3873;
assign w4069 = ~w3864 & ~w3867;
assign w4070 = pi00 & pi45;
assign w4071 = pi02 & pi43;
assign w4072 = pi04 & pi41;
assign w4073 = ~w4071 & ~w4072;
assign w4074 = w4071 & w4072;
assign w4075 = ~w4073 & ~w4074;
assign w4076 = w4070 & ~w4075;
assign w4077 = ~w4070 & w4075;
assign w4078 = ~w4076 & ~w4077;
assign w4079 = pi07 & pi38;
assign w4080 = pi08 & pi37;
assign w4081 = pi09 & pi36;
assign w4082 = ~w4080 & ~w4081;
assign w4083 = w4080 & w4081;
assign w4084 = ~w4082 & ~w4083;
assign w4085 = w4079 & ~w4084;
assign w4086 = ~w4079 & w4084;
assign w4087 = ~w4085 & ~w4086;
assign w4088 = ~w4078 & ~w4087;
assign w4089 = w4078 & w4087;
assign w4090 = ~w4088 & ~w4089;
assign w4091 = pi22 & pi23;
assign w4092 = pi21 & pi24;
assign w4093 = ~w4091 & ~w4092;
assign w4094 = w4091 & w4092;
assign w4095 = ~w4093 & ~w4094;
assign w4096 = w3918 & ~w4095;
assign w4097 = ~w3918 & w4095;
assign w4098 = ~w4096 & ~w4097;
assign w4099 = w4090 & ~w4098;
assign w4100 = ~w4090 & w4098;
assign w4101 = ~w4099 & ~w4100;
assign w4102 = w3914 & ~w3917;
assign w4103 = ~w3919 & ~w4102;
assign w4104 = pi18 & pi27;
assign w4105 = pi20 & pi25;
assign w4106 = pi19 & pi26;
assign w4107 = ~w4105 & ~w4106;
assign w4108 = w4105 & w4106;
assign w4109 = ~w4107 & ~w4108;
assign w4110 = w4104 & ~w4109;
assign w4111 = ~w4104 & w4109;
assign w4112 = ~w4110 & ~w4111;
assign w4113 = ~w4103 & ~w4112;
assign w4114 = w4103 & w4112;
assign w4115 = ~w4113 & ~w4114;
assign w4116 = pi14 & pi31;
assign w4117 = pi13 & pi32;
assign w4118 = pi05 & pi40;
assign w4119 = ~w4117 & ~w4118;
assign w4120 = w4117 & w4118;
assign w4121 = ~w4119 & ~w4120;
assign w4122 = w4116 & ~w4121;
assign w4123 = ~w4116 & w4121;
assign w4124 = ~w4122 & ~w4123;
assign w4125 = w4115 & ~w4124;
assign w4126 = ~w4115 & w4124;
assign w4127 = ~w4125 & ~w4126;
assign w4128 = w4101 & w4127;
assign w4129 = ~w4101 & ~w4127;
assign w4130 = ~w4128 & ~w4129;
assign w4131 = ~w4069 & w4130;
assign w4132 = w4069 & ~w4130;
assign w4133 = ~w4131 & ~w4132;
assign w4134 = ~w4068 & w4133;
assign w4135 = w4068 & ~w4133;
assign w4136 = ~w4134 & ~w4135;
assign w4137 = w4067 & w4136;
assign w4138 = ~w4067 & ~w4136;
assign w4139 = ~w4137 & ~w4138;
assign w4140 = ~w3811 & ~w3968;
assign w4141 = ~w3966 & ~w4140;
assign w4142 = ~w3881 & ~w3885;
assign w4143 = ~w3884 & ~w4142;
assign w4144 = w4141 & w4143;
assign w4145 = ~w4141 & ~w4143;
assign w4146 = ~w4144 & ~w4145;
assign w4147 = ~w3890 & ~w3894;
assign w4148 = ~w3893 & ~w4147;
assign w4149 = ~w4146 & ~w4148;
assign w4150 = w4146 & w4148;
assign w4151 = ~w4149 & ~w4150;
assign w4152 = ~w4002 & ~w4006;
assign w4153 = ~w4151 & w4152;
assign w4154 = w4151 & ~w4152;
assign w4155 = ~w4153 & ~w4154;
assign w4156 = pi12 & pi33;
assign w4157 = pi11 & pi34;
assign w4158 = pi06 & pi39;
assign w4159 = ~w4157 & ~w4158;
assign w4160 = w4157 & w4158;
assign w4161 = ~w4159 & ~w4160;
assign w4162 = w4156 & ~w4161;
assign w4163 = ~w4156 & w4161;
assign w4164 = ~w4162 & ~w4163;
assign w4165 = pi15 & pi30;
assign w4166 = pi16 & pi29;
assign w4167 = pi17 & pi28;
assign w4168 = ~w4166 & ~w4167;
assign w4169 = w4166 & w4167;
assign w4170 = ~w4168 & ~w4169;
assign w4171 = w4165 & ~w4170;
assign w4172 = ~w4165 & w4170;
assign w4173 = ~w4171 & ~w4172;
assign w4174 = ~w4164 & ~w4173;
assign w4175 = w4164 & w4173;
assign w4176 = ~w4174 & ~w4175;
assign w4177 = pi44 & w1127;
assign w4178 = pi01 & pi44;
assign w4179 = ~pi23 & ~w4178;
assign w4180 = ~w4177 & ~w4179;
assign w4181 = pi03 & pi42;
assign w4182 = ~w3979 & ~w4181;
assign w4183 = w3979 & w4181;
assign w4184 = ~w4182 & ~w4183;
assign w4185 = w4180 & ~w4184;
assign w4186 = ~w4180 & w4184;
assign w4187 = ~w4185 & ~w4186;
assign w4188 = w4176 & ~w4187;
assign w4189 = ~w4176 & w4187;
assign w4190 = ~w4188 & ~w4189;
assign w4191 = w4155 & w4190;
assign w4192 = ~w4155 & ~w4190;
assign w4193 = ~w4191 & ~w4192;
assign w4194 = ~w3948 & ~w3951;
assign w4195 = (~w4008 & ~w4010) | (~w4008 & w17087) | (~w4010 & w17087);
assign w4196 = ~w4194 & ~w4195;
assign w4197 = w4194 & w4195;
assign w4198 = ~w4196 & ~w4197;
assign w4199 = w4193 & w4198;
assign w4200 = ~w4193 & ~w4198;
assign w4201 = ~w4199 & ~w4200;
assign w4202 = ~w3954 & ~w4014;
assign w4203 = w4201 & ~w4202;
assign w4204 = ~w4201 & w4202;
assign w4205 = ~w4203 & ~w4204;
assign w4206 = w4139 & w4205;
assign w4207 = ~w4139 & ~w4205;
assign w4208 = ~w4206 & ~w4207;
assign w4209 = ~w4031 & w4208;
assign w4210 = w4031 & ~w4208;
assign w4211 = ~w4209 & ~w4210;
assign w4212 = w4030 & ~w4211;
assign w4213 = ~w4030 & w4211;
assign w4214 = ~w4212 & ~w4213;
assign w4215 = (w3670 & w16523) | (w3670 & w16524) | (w16523 & w16524);
assign w4216 = ~w4210 & ~w4215;
assign w4217 = ~w4203 & ~w4206;
assign w4218 = ~w4134 & ~w4137;
assign w4219 = (~w4049 & ~w4051) | (~w4049 & w17088) | (~w4051 & w17088);
assign w4220 = pi14 & pi32;
assign w4221 = pi06 & pi40;
assign w4222 = pi13 & pi33;
assign w4223 = ~w4221 & ~w4222;
assign w4224 = w4221 & w4222;
assign w4225 = ~w4223 & ~w4224;
assign w4226 = w4220 & ~w4225;
assign w4227 = ~w4220 & w4225;
assign w4228 = ~w4226 & ~w4227;
assign w4229 = pi15 & pi31;
assign w4230 = pi05 & pi41;
assign w4231 = ~w4229 & ~w4230;
assign w4232 = w4229 & w4230;
assign w4233 = ~w4231 & ~w4232;
assign w4234 = w3967 & ~w4233;
assign w4235 = ~w3967 & w4233;
assign w4236 = ~w4234 & ~w4235;
assign w4237 = ~w4228 & ~w4236;
assign w4238 = w4228 & w4236;
assign w4239 = ~w4237 & ~w4238;
assign w4240 = w4219 & ~w4239;
assign w4241 = ~w4219 & w4239;
assign w4242 = ~w4240 & ~w4241;
assign w4243 = ~w4104 & ~w4108;
assign w4244 = ~w4107 & ~w4243;
assign w4245 = ~w4165 & ~w4169;
assign w4246 = ~w4168 & ~w4245;
assign w4247 = w4244 & w4246;
assign w4248 = ~w4244 & ~w4246;
assign w4249 = ~w4247 & ~w4248;
assign w4250 = ~w4156 & ~w4160;
assign w4251 = ~w4159 & ~w4250;
assign w4252 = ~w4249 & ~w4251;
assign w4253 = w4249 & w4251;
assign w4254 = ~w4252 & ~w4253;
assign w4255 = (~w4035 & ~w4037) | (~w4035 & w16875) | (~w4037 & w16875);
assign w4256 = ~w4254 & w4255;
assign w4257 = w4254 & ~w4255;
assign w4258 = ~w4256 & ~w4257;
assign w4259 = w4242 & w4258;
assign w4260 = ~w4242 & ~w4258;
assign w4261 = ~w4259 & ~w4260;
assign w4262 = (~w4043 & ~w4044) | (~w4043 & w17089) | (~w4044 & w17089);
assign w4263 = ~w4128 & ~w4131;
assign w4264 = ~w4262 & ~w4263;
assign w4265 = w4262 & w4263;
assign w4266 = ~w4264 & ~w4265;
assign w4267 = w4261 & w4266;
assign w4268 = ~w4261 & ~w4266;
assign w4269 = ~w4267 & ~w4268;
assign w4270 = ~w4218 & w4269;
assign w4271 = w4218 & ~w4269;
assign w4272 = ~w4270 & ~w4271;
assign w4273 = w4217 & ~w4272;
assign w4274 = ~w4217 & w4272;
assign w4275 = ~w4273 & ~w4274;
assign w4276 = ~w4196 & ~w4199;
assign w4277 = (~w4059 & ~w4061) | (~w4059 & w17090) | (~w4061 & w17090);
assign w4278 = pi03 & pi43;
assign w4279 = pi00 & pi46;
assign w4280 = pi04 & pi42;
assign w4281 = ~w4279 & ~w4280;
assign w4282 = w4279 & w4280;
assign w4283 = ~w4281 & ~w4282;
assign w4284 = w4278 & ~w4283;
assign w4285 = ~w4278 & w4283;
assign w4286 = ~w4284 & ~w4285;
assign w4287 = pi09 & pi37;
assign w4288 = pi11 & pi35;
assign w4289 = pi10 & pi36;
assign w4290 = ~w4288 & ~w4289;
assign w4291 = w4288 & w4289;
assign w4292 = ~w4290 & ~w4291;
assign w4293 = w4287 & ~w4292;
assign w4294 = ~w4287 & w4292;
assign w4295 = ~w4293 & ~w4294;
assign w4296 = ~w4286 & ~w4295;
assign w4297 = w4286 & w4295;
assign w4298 = ~w4296 & ~w4297;
assign w4299 = pi19 & pi27;
assign w4300 = pi20 & pi26;
assign w4301 = pi21 & pi25;
assign w4302 = ~w4300 & ~w4301;
assign w4303 = w4300 & w4301;
assign w4304 = ~w4302 & ~w4303;
assign w4305 = w4299 & ~w4304;
assign w4306 = ~w4299 & w4304;
assign w4307 = ~w4305 & ~w4306;
assign w4308 = w4298 & ~w4307;
assign w4309 = ~w4298 & w4307;
assign w4310 = ~w4308 & ~w4309;
assign w4311 = pi16 & pi30;
assign w4312 = pi17 & pi29;
assign w4313 = pi18 & pi28;
assign w4314 = ~w4312 & ~w4313;
assign w4315 = w4312 & w4313;
assign w4316 = ~w4314 & ~w4315;
assign w4317 = w4311 & ~w4316;
assign w4318 = ~w4311 & w4316;
assign w4319 = ~w4317 & ~w4318;
assign w4320 = ~w4180 & ~w4183;
assign w4321 = ~w4182 & ~w4320;
assign w4322 = ~w4319 & w4321;
assign w4323 = w4319 & ~w4321;
assign w4324 = ~w4322 & ~w4323;
assign w4325 = pi12 & pi34;
assign w4326 = pi08 & pi38;
assign w4327 = pi07 & pi39;
assign w4328 = ~w4326 & ~w4327;
assign w4329 = pi08 & pi39;
assign w4330 = w4079 & w4329;
assign w4331 = ~w4328 & ~w4330;
assign w4332 = w4325 & ~w4331;
assign w4333 = ~w4325 & w4331;
assign w4334 = ~w4332 & ~w4333;
assign w4335 = w4324 & ~w4334;
assign w4336 = ~w4324 & w4334;
assign w4337 = ~w4335 & ~w4336;
assign w4338 = w4310 & w4337;
assign w4339 = ~w4310 & ~w4337;
assign w4340 = ~w4338 & ~w4339;
assign w4341 = ~w4277 & w4340;
assign w4342 = w4277 & ~w4340;
assign w4343 = ~w4341 & ~w4342;
assign w4344 = ~w4276 & w4343;
assign w4345 = w4276 & ~w4343;
assign w4346 = ~w4344 & ~w4345;
assign w4347 = ~w4174 & ~w4188;
assign w4348 = ~w4113 & ~w4125;
assign w4349 = ~w4088 & ~w4099;
assign w4350 = ~w4348 & ~w4349;
assign w4351 = w4348 & w4349;
assign w4352 = ~w4350 & ~w4351;
assign w4353 = w4347 & ~w4352;
assign w4354 = ~w4347 & w4352;
assign w4355 = ~w4353 & ~w4354;
assign w4356 = ~w4154 & ~w4191;
assign w4357 = ~w4116 & ~w4120;
assign w4358 = ~w4119 & ~w4357;
assign w4359 = ~w4070 & ~w4074;
assign w4360 = ~w4073 & ~w4359;
assign w4361 = w4358 & w4360;
assign w4362 = ~w4358 & ~w4360;
assign w4363 = ~w4361 & ~w4362;
assign w4364 = ~w4079 & ~w4083;
assign w4365 = ~w4082 & ~w4364;
assign w4366 = ~w4363 & ~w4365;
assign w4367 = w4363 & w4365;
assign w4368 = ~w4366 & ~w4367;
assign w4369 = (~w4144 & ~w4146) | (~w4144 & w17091) | (~w4146 & w17091);
assign w4370 = pi22 & pi24;
assign w4371 = pi01 & pi45;
assign w4372 = ~w4370 & ~w4371;
assign w4373 = w4370 & w4371;
assign w4374 = ~w4372 & ~w4373;
assign w4375 = w4177 & w4374;
assign w4376 = ~w4177 & ~w4374;
assign w4377 = ~w4375 & ~w4376;
assign w4378 = ~w3918 & ~w4094;
assign w4379 = ~w4093 & ~w4378;
assign w4380 = w4377 & w4379;
assign w4381 = ~w4377 & ~w4379;
assign w4382 = ~w4380 & ~w4381;
assign w4383 = ~w4369 & w4382;
assign w4384 = w4369 & ~w4382;
assign w4385 = ~w4383 & ~w4384;
assign w4386 = w4368 & w4385;
assign w4387 = ~w4368 & ~w4385;
assign w4388 = ~w4386 & ~w4387;
assign w4389 = ~w4356 & w4388;
assign w4390 = w4356 & ~w4388;
assign w4391 = ~w4389 & ~w4390;
assign w4392 = w4355 & w4391;
assign w4393 = ~w4355 & ~w4391;
assign w4394 = ~w4392 & ~w4393;
assign w4395 = w4346 & w4394;
assign w4396 = ~w4346 & ~w4394;
assign w4397 = ~w4395 & ~w4396;
assign w4398 = ~w4275 & ~w4397;
assign w4399 = w4275 & w4397;
assign w4400 = ~w4398 & ~w4399;
assign w4401 = w4216 & ~w4400;
assign w4402 = ~w4216 & w4400;
assign w4403 = ~w4401 & ~w4402;
assign w4404 = ~w4270 & ~w4274;
assign w4405 = ~w3967 & ~w4232;
assign w4406 = ~w4231 & ~w4405;
assign w4407 = ~w4299 & ~w4303;
assign w4408 = ~w4302 & ~w4407;
assign w4409 = w4406 & w4408;
assign w4410 = ~w4406 & ~w4408;
assign w4411 = ~w4409 & ~w4410;
assign w4412 = ~w4278 & ~w4282;
assign w4413 = ~w4281 & ~w4412;
assign w4414 = ~w4411 & ~w4413;
assign w4415 = w4411 & w4413;
assign w4416 = ~w4414 & ~w4415;
assign w4417 = (~w4296 & ~w4298) | (~w4296 & w16876) | (~w4298 & w16876);
assign w4418 = ~w4416 & w4417;
assign w4419 = w4416 & ~w4417;
assign w4420 = ~w4418 & ~w4419;
assign w4421 = ~w4237 & ~w4241;
assign w4422 = ~w4420 & w4421;
assign w4423 = w4420 & ~w4421;
assign w4424 = ~w4422 & ~w4423;
assign w4425 = ~w4338 & ~w4341;
assign w4426 = (~w4257 & ~w4258) | (~w4257 & w17092) | (~w4258 & w17092);
assign w4427 = ~w4425 & ~w4426;
assign w4428 = w4425 & w4426;
assign w4429 = ~w4427 & ~w4428;
assign w4430 = w4424 & w4429;
assign w4431 = ~w4424 & ~w4429;
assign w4432 = ~w4430 & ~w4431;
assign w4433 = ~w4264 & ~w4267;
assign w4434 = ~w4389 & ~w4392;
assign w4435 = ~w4433 & ~w4434;
assign w4436 = w4433 & w4434;
assign w4437 = ~w4435 & ~w4436;
assign w4438 = w4432 & w4437;
assign w4439 = ~w4432 & ~w4437;
assign w4440 = ~w4438 & ~w4439;
assign w4441 = ~w4344 & ~w4395;
assign w4442 = (~w4247 & ~w4249) | (~w4247 & w17093) | (~w4249 & w17093);
assign w4443 = (~w4375 & ~w4377) | (~w4375 & w16877) | (~w4377 & w16877);
assign w4444 = pi13 & pi34;
assign w4445 = pi12 & pi35;
assign w4446 = pi07 & pi40;
assign w4447 = ~w4445 & ~w4446;
assign w4448 = w4445 & w4446;
assign w4449 = ~w4447 & ~w4448;
assign w4450 = w4444 & ~w4449;
assign w4451 = ~w4444 & w4449;
assign w4452 = ~w4450 & ~w4451;
assign w4453 = ~w4443 & ~w4452;
assign w4454 = w4443 & w4452;
assign w4455 = ~w4453 & ~w4454;
assign w4456 = w4442 & ~w4455;
assign w4457 = ~w4442 & w4455;
assign w4458 = ~w4456 & ~w4457;
assign w4459 = ~w4383 & ~w4386;
assign w4460 = ~w4458 & w4459;
assign w4461 = w4458 & ~w4459;
assign w4462 = ~w4460 & ~w4461;
assign w4463 = ~w4350 & ~w4354;
assign w4464 = ~w4462 & w4463;
assign w4465 = w4462 & ~w4463;
assign w4466 = ~w4464 & ~w4465;
assign w4467 = pi01 & pi46;
assign w4468 = ~pi24 & ~w4467;
assign w4469 = pi46 & w1215;
assign w4470 = ~w4468 & ~w4469;
assign w4471 = ~w4287 & ~w4291;
assign w4472 = ~w4290 & ~w4471;
assign w4473 = w4470 & w4472;
assign w4474 = ~w4470 & ~w4472;
assign w4475 = ~w4473 & ~w4474;
assign w4476 = w4325 & ~w4328;
assign w4477 = ~w4330 & ~w4476;
assign w4478 = w4475 & ~w4477;
assign w4479 = ~w4475 & w4477;
assign w4480 = ~w4478 & ~w4479;
assign w4481 = (~w4322 & ~w4324) | (~w4322 & w16878) | (~w4324 & w16878);
assign w4482 = (~w4361 & ~w4363) | (~w4361 & w17094) | (~w4363 & w17094);
assign w4483 = ~w4481 & ~w4482;
assign w4484 = w4481 & w4482;
assign w4485 = ~w4483 & ~w4484;
assign w4486 = ~w4480 & ~w4485;
assign w4487 = w4480 & w4485;
assign w4488 = ~w4486 & ~w4487;
assign w4489 = pi00 & pi47;
assign w4490 = pi02 & pi45;
assign w4491 = ~w4489 & ~w4490;
assign w4492 = pi02 & pi47;
assign w4493 = w4070 & w4492;
assign w4494 = ~w4491 & ~w4493;
assign w4495 = w4373 & ~w4494;
assign w4496 = ~w4373 & w4494;
assign w4497 = ~w4495 & ~w4496;
assign w4498 = pi16 & pi31;
assign w4499 = pi18 & pi29;
assign w4500 = pi17 & pi30;
assign w4501 = ~w4499 & ~w4500;
assign w4502 = w4499 & w4500;
assign w4503 = ~w4501 & ~w4502;
assign w4504 = w4498 & ~w4503;
assign w4505 = ~w4498 & w4503;
assign w4506 = ~w4504 & ~w4505;
assign w4507 = ~w4497 & ~w4506;
assign w4508 = w4497 & w4506;
assign w4509 = ~w4507 & ~w4508;
assign w4510 = pi19 & pi28;
assign w4511 = pi21 & pi26;
assign w4512 = pi20 & pi27;
assign w4513 = ~w4511 & ~w4512;
assign w4514 = w4511 & w4512;
assign w4515 = ~w4513 & ~w4514;
assign w4516 = w4510 & ~w4515;
assign w4517 = ~w4510 & w4515;
assign w4518 = ~w4516 & ~w4517;
assign w4519 = w4509 & ~w4518;
assign w4520 = ~w4509 & w4518;
assign w4521 = ~w4519 & ~w4520;
assign w4522 = ~w4311 & ~w4315;
assign w4523 = ~w4314 & ~w4522;
assign w4524 = ~w4220 & ~w4224;
assign w4525 = ~w4223 & ~w4524;
assign w4526 = w4523 & w4525;
assign w4527 = ~w4523 & ~w4525;
assign w4528 = ~w4526 & ~w4527;
assign w4529 = pi03 & pi44;
assign w4530 = pi04 & pi43;
assign w4531 = pi15 & pi32;
assign w4532 = ~w4530 & ~w4531;
assign w4533 = w4530 & w4531;
assign w4534 = ~w4532 & ~w4533;
assign w4535 = w4529 & ~w4534;
assign w4536 = ~w4529 & w4534;
assign w4537 = ~w4535 & ~w4536;
assign w4538 = ~w4528 & w4537;
assign w4539 = w4528 & ~w4537;
assign w4540 = ~w4538 & ~w4539;
assign w4541 = pi10 & pi37;
assign w4542 = pi23 & pi24;
assign w4543 = pi22 & pi25;
assign w4544 = ~w4542 & ~w4543;
assign w4545 = w4542 & w4543;
assign w4546 = ~w4544 & ~w4545;
assign w4547 = w4541 & ~w4546;
assign w4548 = ~w4541 & w4546;
assign w4549 = ~w4547 & ~w4548;
assign w4550 = pi11 & pi36;
assign w4551 = pi09 & pi38;
assign w4552 = ~w4550 & ~w4551;
assign w4553 = w4550 & w4551;
assign w4554 = ~w4552 & ~w4553;
assign w4555 = w4329 & ~w4554;
assign w4556 = ~w4329 & w4554;
assign w4557 = ~w4555 & ~w4556;
assign w4558 = ~w4549 & ~w4557;
assign w4559 = w4549 & w4557;
assign w4560 = ~w4558 & ~w4559;
assign w4561 = pi05 & pi42;
assign w4562 = pi06 & pi41;
assign w4563 = pi14 & pi33;
assign w4564 = ~w4562 & ~w4563;
assign w4565 = w4562 & w4563;
assign w4566 = ~w4564 & ~w4565;
assign w4567 = w4561 & ~w4566;
assign w4568 = ~w4561 & w4566;
assign w4569 = ~w4567 & ~w4568;
assign w4570 = w4560 & ~w4569;
assign w4571 = ~w4560 & w4569;
assign w4572 = ~w4570 & ~w4571;
assign w4573 = w4540 & w4572;
assign w4574 = ~w4540 & ~w4572;
assign w4575 = ~w4573 & ~w4574;
assign w4576 = w4521 & w4575;
assign w4577 = ~w4521 & ~w4575;
assign w4578 = ~w4576 & ~w4577;
assign w4579 = w4488 & w4578;
assign w4580 = ~w4488 & ~w4578;
assign w4581 = ~w4579 & ~w4580;
assign w4582 = w4466 & w4581;
assign w4583 = ~w4466 & ~w4581;
assign w4584 = ~w4582 & ~w4583;
assign w4585 = ~w4441 & w4584;
assign w4586 = w4441 & ~w4584;
assign w4587 = ~w4585 & ~w4586;
assign w4588 = w4440 & w4587;
assign w4589 = ~w4440 & ~w4587;
assign w4590 = ~w4588 & ~w4589;
assign w4591 = ~w4404 & w4590;
assign w4592 = w4404 & ~w4590;
assign w4593 = ~w4591 & ~w4592;
assign w4594 = ~w4210 & ~w4398;
assign w4595 = ~w4215 & w4594;
assign w4596 = ~w4399 & ~w4595;
assign w4597 = w4593 & w4596;
assign w4598 = ~w4593 & ~w4596;
assign w4599 = ~w4597 & ~w4598;
assign w4600 = ~w4399 & ~w4591;
assign w4601 = (~w4215 & w16526) | (~w4215 & w16527) | (w16526 & w16527);
assign w4602 = ~w4585 & ~w4588;
assign w4603 = ~w4435 & ~w4438;
assign w4604 = ~w4427 & ~w4430;
assign w4605 = ~w4461 & ~w4465;
assign w4606 = (~w4453 & ~w4455) | (~w4453 & w17095) | (~w4455 & w17095);
assign w4607 = pi14 & pi34;
assign w4608 = pi06 & pi42;
assign w4609 = pi13 & pi35;
assign w4610 = ~w4608 & ~w4609;
assign w4611 = w4608 & w4609;
assign w4612 = ~w4610 & ~w4611;
assign w4613 = w4607 & ~w4612;
assign w4614 = ~w4607 & w4612;
assign w4615 = ~w4613 & ~w4614;
assign w4616 = pi07 & pi41;
assign w4617 = pi12 & pi36;
assign w4618 = pi08 & pi40;
assign w4619 = ~w4617 & ~w4618;
assign w4620 = w4617 & w4618;
assign w4621 = ~w4619 & ~w4620;
assign w4622 = w4616 & ~w4621;
assign w4623 = ~w4616 & w4621;
assign w4624 = ~w4622 & ~w4623;
assign w4625 = ~w4615 & ~w4624;
assign w4626 = w4615 & w4624;
assign w4627 = ~w4625 & ~w4626;
assign w4628 = pi09 & pi39;
assign w4629 = pi11 & pi37;
assign w4630 = pi10 & pi38;
assign w4631 = ~w4629 & ~w4630;
assign w4632 = pi11 & pi38;
assign w4633 = w4541 & w4632;
assign w4634 = ~w4631 & ~w4633;
assign w4635 = w4628 & ~w4634;
assign w4636 = ~w4628 & w4634;
assign w4637 = ~w4635 & ~w4636;
assign w4638 = w4627 & ~w4637;
assign w4639 = ~w4627 & w4637;
assign w4640 = ~w4638 & ~w4639;
assign w4641 = ~w4606 & w4640;
assign w4642 = w4606 & ~w4640;
assign w4643 = ~w4641 & ~w4642;
assign w4644 = pi04 & pi44;
assign w4645 = pi05 & pi43;
assign w4646 = pi15 & pi33;
assign w4647 = ~w4645 & ~w4646;
assign w4648 = w4645 & w4646;
assign w4649 = ~w4647 & ~w4648;
assign w4650 = w4644 & ~w4649;
assign w4651 = ~w4644 & w4649;
assign w4652 = ~w4650 & ~w4651;
assign w4653 = pi20 & pi28;
assign w4654 = pi21 & pi27;
assign w4655 = pi22 & pi26;
assign w4656 = ~w4654 & ~w4655;
assign w4657 = w4654 & w4655;
assign w4658 = ~w4656 & ~w4657;
assign w4659 = w4653 & ~w4658;
assign w4660 = ~w4653 & w4658;
assign w4661 = ~w4659 & ~w4660;
assign w4662 = ~w4652 & ~w4661;
assign w4663 = w4652 & w4661;
assign w4664 = ~w4662 & ~w4663;
assign w4665 = pi17 & pi31;
assign w4666 = pi18 & pi30;
assign w4667 = pi19 & pi29;
assign w4668 = ~w4666 & ~w4667;
assign w4669 = w4666 & w4667;
assign w4670 = ~w4668 & ~w4669;
assign w4671 = w4665 & ~w4670;
assign w4672 = ~w4665 & w4670;
assign w4673 = ~w4671 & ~w4672;
assign w4674 = w4664 & ~w4673;
assign w4675 = ~w4664 & w4673;
assign w4676 = ~w4674 & ~w4675;
assign w4677 = ~w4643 & ~w4676;
assign w4678 = w4643 & w4676;
assign w4679 = ~w4677 & ~w4678;
assign w4680 = ~w4605 & w4679;
assign w4681 = w4605 & ~w4679;
assign w4682 = ~w4680 & ~w4681;
assign w4683 = ~w4604 & w4682;
assign w4684 = w4604 & ~w4682;
assign w4685 = ~w4683 & ~w4684;
assign w4686 = ~w4603 & w4685;
assign w4687 = w4603 & ~w4685;
assign w4688 = ~w4686 & ~w4687;
assign w4689 = ~w4510 & ~w4514;
assign w4690 = ~w4513 & ~w4689;
assign w4691 = ~w4329 & ~w4553;
assign w4692 = ~w4552 & ~w4691;
assign w4693 = w4690 & w4692;
assign w4694 = ~w4690 & ~w4692;
assign w4695 = ~w4693 & ~w4694;
assign w4696 = ~w4561 & ~w4565;
assign w4697 = ~w4564 & ~w4696;
assign w4698 = ~w4695 & ~w4697;
assign w4699 = w4695 & w4697;
assign w4700 = ~w4698 & ~w4699;
assign w4701 = (~w4558 & ~w4560) | (~w4558 & w16879) | (~w4560 & w16879);
assign w4702 = ~w4700 & w4701;
assign w4703 = w4700 & ~w4701;
assign w4704 = ~w4702 & ~w4703;
assign w4705 = ~w4444 & ~w4448;
assign w4706 = ~w4447 & ~w4705;
assign w4707 = ~w4541 & ~w4545;
assign w4708 = ~w4544 & ~w4707;
assign w4709 = w4706 & w4708;
assign w4710 = ~w4706 & ~w4708;
assign w4711 = ~w4709 & ~w4710;
assign w4712 = pi02 & pi46;
assign w4713 = pi03 & pi45;
assign w4714 = pi16 & pi32;
assign w4715 = ~w4713 & ~w4714;
assign w4716 = w4713 & w4714;
assign w4717 = ~w4715 & ~w4716;
assign w4718 = w4712 & ~w4717;
assign w4719 = ~w4712 & w4717;
assign w4720 = ~w4718 & ~w4719;
assign w4721 = ~w4711 & w4720;
assign w4722 = w4711 & ~w4720;
assign w4723 = ~w4721 & ~w4722;
assign w4724 = ~w4704 & ~w4723;
assign w4725 = w4704 & w4723;
assign w4726 = ~w4724 & ~w4725;
assign w4727 = ~w4573 & ~w4576;
assign w4728 = ~w4726 & w4727;
assign w4729 = w4726 & ~w4727;
assign w4730 = ~w4728 & ~w4729;
assign w4731 = ~w4498 & ~w4502;
assign w4732 = ~w4501 & ~w4731;
assign w4733 = ~w4529 & ~w4533;
assign w4734 = ~w4532 & ~w4733;
assign w4735 = w4732 & w4734;
assign w4736 = ~w4732 & ~w4734;
assign w4737 = ~w4735 & ~w4736;
assign w4738 = w4373 & ~w4491;
assign w4739 = ~w4493 & ~w4738;
assign w4740 = ~w4737 & w4739;
assign w4741 = w4737 & ~w4739;
assign w4742 = ~w4740 & ~w4741;
assign w4743 = (~w4473 & ~w4475) | (~w4473 & w17096) | (~w4475 & w17096);
assign w4744 = (~w4507 & ~w4509) | (~w4507 & w16880) | (~w4509 & w16880);
assign w4745 = ~w4743 & ~w4744;
assign w4746 = w4743 & w4744;
assign w4747 = ~w4745 & ~w4746;
assign w4748 = w4742 & w4747;
assign w4749 = ~w4742 & ~w4747;
assign w4750 = ~w4748 & ~w4749;
assign w4751 = w4730 & w4750;
assign w4752 = ~w4730 & ~w4750;
assign w4753 = ~w4751 & ~w4752;
assign w4754 = ~w4579 & ~w4582;
assign w4755 = (~w4526 & ~w4528) | (~w4526 & w17097) | (~w4528 & w17097);
assign w4756 = (~w4409 & ~w4411) | (~w4409 & w16734) | (~w4411 & w16734);
assign w4757 = pi00 & pi48;
assign w4758 = w4469 & w4757;
assign w4759 = ~w4469 & ~w4757;
assign w4760 = ~w4758 & ~w4759;
assign w4761 = pi23 & pi25;
assign w4762 = pi01 & pi47;
assign w4763 = ~w4761 & ~w4762;
assign w4764 = w4761 & w4762;
assign w4765 = ~w4763 & ~w4764;
assign w4766 = w4760 & w4765;
assign w4767 = ~w4760 & ~w4765;
assign w4768 = ~w4766 & ~w4767;
assign w4769 = ~w4756 & w4768;
assign w4770 = w4756 & ~w4768;
assign w4771 = ~w4769 & ~w4770;
assign w4772 = w4755 & ~w4771;
assign w4773 = ~w4755 & w4771;
assign w4774 = ~w4772 & ~w4773;
assign w4775 = (~w4419 & ~w4420) | (~w4419 & w17098) | (~w4420 & w17098);
assign w4776 = (~w4483 & ~w4485) | (~w4483 & w17099) | (~w4485 & w17099);
assign w4777 = ~w4775 & ~w4776;
assign w4778 = w4775 & w4776;
assign w4779 = ~w4777 & ~w4778;
assign w4780 = w4774 & w4779;
assign w4781 = ~w4774 & ~w4779;
assign w4782 = ~w4780 & ~w4781;
assign w4783 = ~w4754 & w4782;
assign w4784 = w4754 & ~w4782;
assign w4785 = ~w4783 & ~w4784;
assign w4786 = w4753 & w4785;
assign w4787 = ~w4753 & ~w4785;
assign w4788 = ~w4786 & ~w4787;
assign w4789 = w4688 & w4788;
assign w4790 = ~w4688 & ~w4788;
assign w4791 = ~w4789 & ~w4790;
assign w4792 = w4602 & ~w4791;
assign w4793 = ~w4602 & w4791;
assign w4794 = ~w4792 & ~w4793;
assign w4795 = w4601 & ~w4794;
assign w4796 = ~w4601 & w4794;
assign w4797 = ~w4795 & ~w4796;
assign w4798 = ~w4601 & ~w4793;
assign w4799 = ~w4792 & ~w4798;
assign w4800 = ~w4783 & ~w4786;
assign w4801 = ~w4729 & ~w4751;
assign w4802 = ~w4777 & ~w4780;
assign w4803 = pi22 & pi27;
assign w4804 = pi03 & pi46;
assign w4805 = ~w4492 & ~w4804;
assign w4806 = pi03 & pi47;
assign w4807 = w4712 & w4806;
assign w4808 = ~w4805 & ~w4807;
assign w4809 = w4803 & ~w4808;
assign w4810 = ~w4803 & w4808;
assign w4811 = ~w4809 & ~w4810;
assign w4812 = pi19 & pi30;
assign w4813 = pi21 & pi28;
assign w4814 = pi20 & pi29;
assign w4815 = ~w4813 & ~w4814;
assign w4816 = w4813 & w4814;
assign w4817 = ~w4815 & ~w4816;
assign w4818 = w4812 & ~w4817;
assign w4819 = ~w4812 & w4817;
assign w4820 = ~w4818 & ~w4819;
assign w4821 = ~w4811 & ~w4820;
assign w4822 = w4811 & w4820;
assign w4823 = ~w4821 & ~w4822;
assign w4824 = pi09 & pi40;
assign w4825 = pi12 & pi37;
assign w4826 = pi10 & pi39;
assign w4827 = ~w4825 & ~w4826;
assign w4828 = w4825 & w4826;
assign w4829 = ~w4827 & ~w4828;
assign w4830 = w4824 & ~w4829;
assign w4831 = ~w4824 & w4829;
assign w4832 = ~w4830 & ~w4831;
assign w4833 = w4823 & ~w4832;
assign w4834 = ~w4823 & w4832;
assign w4835 = ~w4833 & ~w4834;
assign w4836 = (~w4758 & ~w4760) | (~w4758 & w16735) | (~w4760 & w16735);
assign w4837 = pi00 & pi49;
assign w4838 = pi04 & pi45;
assign w4839 = pi05 & pi44;
assign w4840 = ~w4838 & ~w4839;
assign w4841 = pi05 & pi45;
assign w4842 = w4644 & w4841;
assign w4843 = ~w4840 & ~w4842;
assign w4844 = w4837 & ~w4843;
assign w4845 = ~w4837 & w4843;
assign w4846 = ~w4844 & ~w4845;
assign w4847 = ~w4836 & ~w4846;
assign w4848 = w4836 & w4846;
assign w4849 = ~w4847 & ~w4848;
assign w4850 = pi16 & pi33;
assign w4851 = pi17 & pi32;
assign w4852 = pi18 & pi31;
assign w4853 = ~w4851 & ~w4852;
assign w4854 = w4851 & w4852;
assign w4855 = ~w4853 & ~w4854;
assign w4856 = w4850 & ~w4855;
assign w4857 = ~w4850 & w4855;
assign w4858 = ~w4856 & ~w4857;
assign w4859 = w4849 & ~w4858;
assign w4860 = ~w4849 & w4858;
assign w4861 = ~w4859 & ~w4860;
assign w4862 = w4835 & w4861;
assign w4863 = ~w4835 & ~w4861;
assign w4864 = ~w4862 & ~w4863;
assign w4865 = pi13 & pi36;
assign w4866 = pi08 & pi41;
assign w4867 = pi07 & pi42;
assign w4868 = ~w4866 & ~w4867;
assign w4869 = pi08 & pi42;
assign w4870 = w4616 & w4869;
assign w4871 = ~w4868 & ~w4870;
assign w4872 = w4865 & ~w4871;
assign w4873 = ~w4865 & w4871;
assign w4874 = ~w4872 & ~w4873;
assign w4875 = pi24 & pi25;
assign w4876 = pi23 & pi26;
assign w4877 = ~w4875 & ~w4876;
assign w4878 = w4875 & w4876;
assign w4879 = ~w4877 & ~w4878;
assign w4880 = w4632 & ~w4879;
assign w4881 = ~w4632 & w4879;
assign w4882 = ~w4880 & ~w4881;
assign w4883 = ~w4874 & ~w4882;
assign w4884 = w4874 & w4882;
assign w4885 = ~w4883 & ~w4884;
assign w4886 = pi15 & pi34;
assign w4887 = pi06 & pi43;
assign w4888 = pi14 & pi35;
assign w4889 = ~w4887 & ~w4888;
assign w4890 = w4887 & w4888;
assign w4891 = ~w4889 & ~w4890;
assign w4892 = w4886 & ~w4891;
assign w4893 = ~w4886 & w4891;
assign w4894 = ~w4892 & ~w4893;
assign w4895 = w4885 & ~w4894;
assign w4896 = ~w4885 & w4894;
assign w4897 = ~w4895 & ~w4896;
assign w4898 = w4864 & w4897;
assign w4899 = ~w4864 & ~w4897;
assign w4900 = ~w4898 & ~w4899;
assign w4901 = ~w4802 & w4900;
assign w4902 = w4802 & ~w4900;
assign w4903 = ~w4901 & ~w4902;
assign w4904 = ~w4801 & w4903;
assign w4905 = w4801 & ~w4903;
assign w4906 = ~w4904 & ~w4905;
assign w4907 = ~w4800 & w4906;
assign w4908 = w4800 & ~w4906;
assign w4909 = ~w4907 & ~w4908;
assign w4910 = ~w4665 & ~w4669;
assign w4911 = ~w4668 & ~w4910;
assign w4912 = ~w4607 & ~w4611;
assign w4913 = ~w4610 & ~w4912;
assign w4914 = w4911 & w4913;
assign w4915 = ~w4911 & ~w4913;
assign w4916 = ~w4914 & ~w4915;
assign w4917 = ~w4616 & ~w4620;
assign w4918 = ~w4619 & ~w4917;
assign w4919 = ~w4916 & ~w4918;
assign w4920 = w4916 & w4918;
assign w4921 = ~w4919 & ~w4920;
assign w4922 = (~w4662 & ~w4664) | (~w4662 & w16881) | (~w4664 & w16881);
assign w4923 = ~w4921 & w4922;
assign w4924 = w4921 & ~w4922;
assign w4925 = ~w4923 & ~w4924;
assign w4926 = (~w4769 & ~w4771) | (~w4769 & w16882) | (~w4771 & w16882);
assign w4927 = ~w4925 & w4926;
assign w4928 = w4925 & ~w4926;
assign w4929 = ~w4927 & ~w4928;
assign w4930 = ~w4641 & ~w4678;
assign w4931 = ~w4929 & w4930;
assign w4932 = w4929 & ~w4930;
assign w4933 = ~w4931 & ~w4932;
assign w4934 = ~w4644 & ~w4648;
assign w4935 = ~w4647 & ~w4934;
assign w4936 = ~w4712 & ~w4716;
assign w4937 = ~w4715 & ~w4936;
assign w4938 = w4935 & w4937;
assign w4939 = ~w4935 & ~w4937;
assign w4940 = ~w4938 & ~w4939;
assign w4941 = ~w4653 & ~w4657;
assign w4942 = ~w4656 & ~w4941;
assign w4943 = ~w4940 & ~w4942;
assign w4944 = w4940 & w4942;
assign w4945 = ~w4943 & ~w4944;
assign w4946 = (~w4625 & ~w4627) | (~w4625 & w16883) | (~w4627 & w16883);
assign w4947 = ~pi48 & w4764;
assign w4948 = pi48 & w1296;
assign w4949 = pi01 & pi48;
assign w4950 = ~pi25 & ~w4949;
assign w4951 = ~w4948 & ~w4950;
assign w4952 = ~w4764 & ~w4951;
assign w4953 = ~w4947 & ~w4952;
assign w4954 = w4628 & ~w4631;
assign w4955 = ~w4633 & ~w4954;
assign w4956 = w4953 & ~w4955;
assign w4957 = ~w4953 & w4955;
assign w4958 = ~w4956 & ~w4957;
assign w4959 = ~w4946 & w4958;
assign w4960 = w4946 & ~w4958;
assign w4961 = ~w4959 & ~w4960;
assign w4962 = w4945 & w4961;
assign w4963 = ~w4945 & ~w4961;
assign w4964 = ~w4962 & ~w4963;
assign w4965 = w4933 & w4964;
assign w4966 = ~w4933 & ~w4964;
assign w4967 = ~w4965 & ~w4966;
assign w4968 = ~w4680 & ~w4683;
assign w4969 = (~w4735 & ~w4737) | (~w4735 & w17100) | (~w4737 & w17100);
assign w4970 = (~w4693 & ~w4695) | (~w4693 & w16736) | (~w4695 & w16736);
assign w4971 = (~w4709 & ~w4711) | (~w4709 & w16737) | (~w4711 & w16737);
assign w4972 = ~w4970 & ~w4971;
assign w4973 = w4970 & w4971;
assign w4974 = ~w4972 & ~w4973;
assign w4975 = w4969 & ~w4974;
assign w4976 = ~w4969 & w4974;
assign w4977 = ~w4975 & ~w4976;
assign w4978 = (~w4703 & ~w4704) | (~w4703 & w17101) | (~w4704 & w17101);
assign w4979 = (~w4745 & ~w4747) | (~w4745 & w17102) | (~w4747 & w17102);
assign w4980 = ~w4978 & ~w4979;
assign w4981 = w4978 & w4979;
assign w4982 = ~w4980 & ~w4981;
assign w4983 = ~w4977 & ~w4982;
assign w4984 = w4977 & w4982;
assign w4985 = ~w4983 & ~w4984;
assign w4986 = ~w4968 & w4985;
assign w4987 = w4968 & ~w4985;
assign w4988 = ~w4986 & ~w4987;
assign w4989 = w4967 & w4988;
assign w4990 = ~w4967 & ~w4988;
assign w4991 = ~w4989 & ~w4990;
assign w4992 = w4909 & w4991;
assign w4993 = ~w4909 & ~w4991;
assign w4994 = ~w4992 & ~w4993;
assign w4995 = ~w4686 & ~w4789;
assign w4996 = ~w4994 & w4995;
assign w4997 = w4994 & ~w4995;
assign w4998 = ~w4996 & ~w4997;
assign w4999 = w4799 & w4998;
assign w5000 = ~w4799 & ~w4998;
assign w5001 = ~w4999 & ~w5000;
assign w5002 = ~w4792 & ~w4996;
assign w5003 = (w5002 & w4601) | (w5002 & w16528) | (w4601 & w16528);
assign w5004 = ~w4997 & ~w5003;
assign w5005 = ~w4907 & ~w4992;
assign w5006 = ~w4986 & ~w4989;
assign w5007 = ~w4932 & ~w4965;
assign w5008 = ~w4980 & ~w4984;
assign w5009 = (~w4947 & ~w4953) | (~w4947 & w16884) | (~w4953 & w16884);
assign w5010 = pi22 & pi28;
assign w5011 = pi18 & pi32;
assign w5012 = pi23 & pi27;
assign w5013 = ~w5011 & ~w5012;
assign w5014 = w5011 & w5012;
assign w5015 = ~w5013 & ~w5014;
assign w5016 = w5010 & ~w5015;
assign w5017 = ~w5010 & w5015;
assign w5018 = ~w5016 & ~w5017;
assign w5019 = pi16 & pi34;
assign w5020 = pi15 & pi35;
assign w5021 = ~w4841 & ~w5020;
assign w5022 = w4841 & w5020;
assign w5023 = ~w5021 & ~w5022;
assign w5024 = w5019 & ~w5023;
assign w5025 = ~w5019 & w5023;
assign w5026 = ~w5024 & ~w5025;
assign w5027 = ~w5018 & ~w5026;
assign w5028 = w5018 & w5026;
assign w5029 = ~w5027 & ~w5028;
assign w5030 = w5009 & ~w5029;
assign w5031 = ~w5009 & w5029;
assign w5032 = ~w5030 & ~w5031;
assign w5033 = pi04 & pi46;
assign w5034 = pi17 & pi33;
assign w5035 = ~w5033 & ~w5034;
assign w5036 = w5033 & w5034;
assign w5037 = ~w5035 & ~w5036;
assign w5038 = w4806 & ~w5037;
assign w5039 = ~w4806 & w5037;
assign w5040 = ~w5038 & ~w5039;
assign w5041 = pi00 & pi50;
assign w5042 = pi02 & pi48;
assign w5043 = ~w5041 & ~w5042;
assign w5044 = pi02 & pi50;
assign w5045 = w4757 & w5044;
assign w5046 = ~w5043 & ~w5045;
assign w5047 = w4948 & ~w5046;
assign w5048 = ~w4948 & w5046;
assign w5049 = ~w5047 & ~w5048;
assign w5050 = ~w5040 & ~w5049;
assign w5051 = w5040 & w5049;
assign w5052 = ~w5050 & ~w5051;
assign w5053 = pi19 & pi31;
assign w5054 = pi21 & pi29;
assign w5055 = pi20 & pi30;
assign w5056 = ~w5054 & ~w5055;
assign w5057 = w5054 & w5055;
assign w5058 = ~w5056 & ~w5057;
assign w5059 = w5053 & ~w5058;
assign w5060 = ~w5053 & w5058;
assign w5061 = ~w5059 & ~w5060;
assign w5062 = w5052 & ~w5061;
assign w5063 = ~w5052 & w5061;
assign w5064 = ~w5062 & ~w5063;
assign w5065 = pi06 & pi44;
assign w5066 = pi07 & pi43;
assign w5067 = pi14 & pi36;
assign w5068 = ~w5066 & ~w5067;
assign w5069 = w5066 & w5067;
assign w5070 = ~w5068 & ~w5069;
assign w5071 = w5065 & ~w5070;
assign w5072 = ~w5065 & w5070;
assign w5073 = ~w5071 & ~w5072;
assign w5074 = pi13 & pi37;
assign w5075 = pi09 & pi41;
assign w5076 = ~w5074 & ~w5075;
assign w5077 = w5074 & w5075;
assign w5078 = ~w5076 & ~w5077;
assign w5079 = w4869 & ~w5078;
assign w5080 = ~w4869 & w5078;
assign w5081 = ~w5079 & ~w5080;
assign w5082 = ~w5073 & ~w5081;
assign w5083 = w5073 & w5081;
assign w5084 = ~w5082 & ~w5083;
assign w5085 = pi12 & pi38;
assign w5086 = pi11 & pi39;
assign w5087 = pi10 & pi40;
assign w5088 = ~w5086 & ~w5087;
assign w5089 = w5086 & w5087;
assign w5090 = ~w5088 & ~w5089;
assign w5091 = w5085 & ~w5090;
assign w5092 = ~w5085 & w5090;
assign w5093 = ~w5091 & ~w5092;
assign w5094 = w5084 & ~w5093;
assign w5095 = ~w5084 & w5093;
assign w5096 = ~w5094 & ~w5095;
assign w5097 = w5064 & w5096;
assign w5098 = ~w5064 & ~w5096;
assign w5099 = ~w5097 & ~w5098;
assign w5100 = ~w5032 & ~w5099;
assign w5101 = w5032 & w5099;
assign w5102 = ~w5100 & ~w5101;
assign w5103 = ~w5008 & w5102;
assign w5104 = w5008 & ~w5102;
assign w5105 = ~w5103 & ~w5104;
assign w5106 = ~w5007 & w5105;
assign w5107 = w5007 & ~w5105;
assign w5108 = ~w5106 & ~w5107;
assign w5109 = ~w5006 & w5108;
assign w5110 = w5006 & ~w5108;
assign w5111 = ~w5109 & ~w5110;
assign w5112 = ~w4901 & ~w4904;
assign w5113 = w4837 & ~w4840;
assign w5114 = ~w4842 & ~w5113;
assign w5115 = w4803 & ~w4805;
assign w5116 = ~w4807 & ~w5115;
assign w5117 = ~w5114 & ~w5116;
assign w5118 = w5114 & w5116;
assign w5119 = ~w5117 & ~w5118;
assign w5120 = ~w4886 & ~w4890;
assign w5121 = ~w4889 & ~w5120;
assign w5122 = ~w5119 & ~w5121;
assign w5123 = w5119 & w5121;
assign w5124 = ~w5122 & ~w5123;
assign w5125 = (~w4914 & ~w4916) | (~w4914 & w16738) | (~w4916 & w16738);
assign w5126 = (~w4938 & ~w4940) | (~w4938 & w16739) | (~w4940 & w16739);
assign w5127 = ~w5125 & ~w5126;
assign w5128 = w5125 & w5126;
assign w5129 = ~w5127 & ~w5128;
assign w5130 = w5124 & w5129;
assign w5131 = ~w5124 & ~w5129;
assign w5132 = ~w5130 & ~w5131;
assign w5133 = ~w4924 & ~w4928;
assign w5134 = (~w4959 & ~w4961) | (~w4959 & w17103) | (~w4961 & w17103);
assign w5135 = ~w5133 & ~w5134;
assign w5136 = w5133 & w5134;
assign w5137 = ~w5135 & ~w5136;
assign w5138 = w5132 & w5137;
assign w5139 = ~w5132 & ~w5137;
assign w5140 = ~w5138 & ~w5139;
assign w5141 = ~w5112 & w5140;
assign w5142 = w5112 & ~w5140;
assign w5143 = ~w5141 & ~w5142;
assign w5144 = pi24 & pi26;
assign w5145 = pi01 & pi49;
assign w5146 = ~w5144 & ~w5145;
assign w5147 = w5144 & w5145;
assign w5148 = ~w5146 & ~w5147;
assign w5149 = ~w4632 & ~w4878;
assign w5150 = ~w4877 & ~w5149;
assign w5151 = w5148 & w5150;
assign w5152 = ~w5148 & ~w5150;
assign w5153 = ~w5151 & ~w5152;
assign w5154 = ~w4824 & ~w4828;
assign w5155 = ~w4827 & ~w5154;
assign w5156 = w5153 & w5155;
assign w5157 = ~w5153 & ~w5155;
assign w5158 = ~w5156 & ~w5157;
assign w5159 = (~w4821 & ~w4823) | (~w4821 & w16885) | (~w4823 & w16885);
assign w5160 = (~w4847 & ~w4849) | (~w4847 & w16886) | (~w4849 & w16886);
assign w5161 = ~w5159 & ~w5160;
assign w5162 = w5159 & w5160;
assign w5163 = ~w5161 & ~w5162;
assign w5164 = w5158 & w5163;
assign w5165 = ~w5158 & ~w5163;
assign w5166 = ~w5164 & ~w5165;
assign w5167 = ~w4812 & ~w4816;
assign w5168 = ~w4815 & ~w5167;
assign w5169 = ~w4850 & ~w4854;
assign w5170 = ~w4853 & ~w5169;
assign w5171 = w5168 & w5170;
assign w5172 = ~w5168 & ~w5170;
assign w5173 = ~w5171 & ~w5172;
assign w5174 = w4865 & ~w4868;
assign w5175 = ~w4870 & ~w5174;
assign w5176 = ~w5173 & w5175;
assign w5177 = w5173 & ~w5175;
assign w5178 = ~w5176 & ~w5177;
assign w5179 = (~w4883 & ~w4885) | (~w4883 & w16887) | (~w4885 & w16887);
assign w5180 = ~w5178 & w5179;
assign w5181 = w5178 & ~w5179;
assign w5182 = ~w5180 & ~w5181;
assign w5183 = (~w4972 & ~w4974) | (~w4972 & w16888) | (~w4974 & w16888);
assign w5184 = ~w5182 & w5183;
assign w5185 = w5182 & ~w5183;
assign w5186 = ~w5184 & ~w5185;
assign w5187 = ~w4862 & ~w4898;
assign w5188 = ~w5186 & w5187;
assign w5189 = w5186 & ~w5187;
assign w5190 = ~w5188 & ~w5189;
assign w5191 = w5166 & w5190;
assign w5192 = ~w5166 & ~w5190;
assign w5193 = ~w5191 & ~w5192;
assign w5194 = w5143 & w5193;
assign w5195 = ~w5143 & ~w5193;
assign w5196 = ~w5194 & ~w5195;
assign w5197 = w5111 & w5196;
assign w5198 = ~w5111 & ~w5196;
assign w5199 = ~w5197 & ~w5198;
assign w5200 = ~w5005 & w5199;
assign w5201 = w5005 & ~w5199;
assign w5202 = ~w5200 & ~w5201;
assign w5203 = w5004 & w5202;
assign w5204 = ~w5004 & ~w5202;
assign w5205 = ~w5203 & ~w5204;
assign w5206 = ~w4997 & ~w5200;
assign w5207 = (w4601 & w16530) | (w4601 & w16531) | (w16530 & w16531);
assign w5208 = ~w5109 & ~w5197;
assign w5209 = ~w5141 & ~w5194;
assign w5210 = ~w5189 & ~w5191;
assign w5211 = (~w5135 & ~w5137) | (~w5135 & w17104) | (~w5137 & w17104);
assign w5212 = (~w5171 & ~w5173) | (~w5171 & w17105) | (~w5173 & w17105);
assign w5213 = pi00 & pi51;
assign w5214 = w5147 & w5213;
assign w5215 = ~w5147 & ~w5213;
assign w5216 = ~w5214 & ~w5215;
assign w5217 = pi01 & pi50;
assign w5218 = pi26 & w5217;
assign w5219 = ~pi26 & ~w5217;
assign w5220 = ~w5218 & ~w5219;
assign w5221 = w5216 & w5220;
assign w5222 = ~w5216 & ~w5220;
assign w5223 = ~w5221 & ~w5222;
assign w5224 = pi17 & pi34;
assign w5225 = pi20 & pi31;
assign w5226 = pi19 & pi32;
assign w5227 = ~w5225 & ~w5226;
assign w5228 = w5225 & w5226;
assign w5229 = ~w5227 & ~w5228;
assign w5230 = w5224 & ~w5229;
assign w5231 = ~w5224 & w5229;
assign w5232 = ~w5230 & ~w5231;
assign w5233 = w5223 & ~w5232;
assign w5234 = ~w5223 & w5232;
assign w5235 = ~w5233 & ~w5234;
assign w5236 = w5212 & ~w5235;
assign w5237 = ~w5212 & w5235;
assign w5238 = ~w5236 & ~w5237;
assign w5239 = pi18 & pi33;
assign w5240 = pi05 & pi46;
assign w5241 = pi16 & pi35;
assign w5242 = ~w5240 & ~w5241;
assign w5243 = w5240 & w5241;
assign w5244 = ~w5242 & ~w5243;
assign w5245 = w5239 & ~w5244;
assign w5246 = ~w5239 & w5244;
assign w5247 = ~w5245 & ~w5246;
assign w5248 = pi21 & pi30;
assign w5249 = pi22 & pi29;
assign w5250 = pi23 & pi28;
assign w5251 = ~w5249 & ~w5250;
assign w5252 = w5249 & w5250;
assign w5253 = ~w5251 & ~w5252;
assign w5254 = w5248 & ~w5253;
assign w5255 = ~w5248 & w5253;
assign w5256 = ~w5254 & ~w5255;
assign w5257 = ~w5247 & ~w5256;
assign w5258 = w5247 & w5256;
assign w5259 = ~w5257 & ~w5258;
assign w5260 = pi15 & pi36;
assign w5261 = pi06 & pi45;
assign w5262 = pi14 & pi37;
assign w5263 = ~w5261 & ~w5262;
assign w5264 = w5261 & w5262;
assign w5265 = ~w5263 & ~w5264;
assign w5266 = w5260 & ~w5265;
assign w5267 = ~w5260 & w5265;
assign w5268 = ~w5266 & ~w5267;
assign w5269 = w5259 & ~w5268;
assign w5270 = ~w5259 & w5268;
assign w5271 = ~w5269 & ~w5270;
assign w5272 = pi07 & pi44;
assign w5273 = pi13 & pi38;
assign w5274 = pi08 & pi43;
assign w5275 = ~w5273 & ~w5274;
assign w5276 = w5273 & w5274;
assign w5277 = ~w5275 & ~w5276;
assign w5278 = w5272 & ~w5277;
assign w5279 = ~w5272 & w5277;
assign w5280 = ~w5278 & ~w5279;
assign w5281 = pi09 & pi42;
assign w5282 = pi12 & pi39;
assign w5283 = pi10 & pi41;
assign w5284 = ~w5282 & ~w5283;
assign w5285 = w5282 & w5283;
assign w5286 = ~w5284 & ~w5285;
assign w5287 = w5281 & ~w5286;
assign w5288 = ~w5281 & w5286;
assign w5289 = ~w5287 & ~w5288;
assign w5290 = ~w5280 & ~w5289;
assign w5291 = w5280 & w5289;
assign w5292 = ~w5290 & ~w5291;
assign w5293 = pi11 & pi40;
assign w5294 = pi25 & pi26;
assign w5295 = pi24 & pi27;
assign w5296 = ~w5294 & ~w5295;
assign w5297 = w5294 & w5295;
assign w5298 = ~w5296 & ~w5297;
assign w5299 = w5293 & ~w5298;
assign w5300 = ~w5293 & w5298;
assign w5301 = ~w5299 & ~w5300;
assign w5302 = w5292 & ~w5301;
assign w5303 = ~w5292 & w5301;
assign w5304 = ~w5302 & ~w5303;
assign w5305 = w5271 & w5304;
assign w5306 = ~w5271 & ~w5304;
assign w5307 = ~w5305 & ~w5306;
assign w5308 = ~w5238 & ~w5307;
assign w5309 = w5238 & w5307;
assign w5310 = ~w5308 & ~w5309;
assign w5311 = ~w5211 & w5310;
assign w5312 = w5211 & ~w5310;
assign w5313 = ~w5311 & ~w5312;
assign w5314 = ~w5210 & w5313;
assign w5315 = w5210 & ~w5313;
assign w5316 = ~w5314 & ~w5315;
assign w5317 = ~w5209 & w5316;
assign w5318 = w5209 & ~w5316;
assign w5319 = ~w5317 & ~w5318;
assign w5320 = ~w5103 & ~w5106;
assign w5321 = ~w5050 & ~w5062;
assign w5322 = (~w5117 & ~w5119) | (~w5117 & w17106) | (~w5119 & w17106);
assign w5323 = (~w5151 & ~w5153) | (~w5151 & w17107) | (~w5153 & w17107);
assign w5324 = ~w5322 & ~w5323;
assign w5325 = w5322 & w5323;
assign w5326 = ~w5324 & ~w5325;
assign w5327 = w5321 & ~w5326;
assign w5328 = ~w5321 & w5326;
assign w5329 = ~w5327 & ~w5328;
assign w5330 = ~w5181 & ~w5185;
assign w5331 = (~w5161 & ~w5163) | (~w5161 & w17108) | (~w5163 & w17108);
assign w5332 = ~w5330 & ~w5331;
assign w5333 = w5330 & w5331;
assign w5334 = ~w5332 & ~w5333;
assign w5335 = w5329 & w5334;
assign w5336 = ~w5329 & ~w5334;
assign w5337 = ~w5335 & ~w5336;
assign w5338 = ~w5320 & w5337;
assign w5339 = w5320 & ~w5337;
assign w5340 = ~w5338 & ~w5339;
assign w5341 = ~w5097 & ~w5101;
assign w5342 = (~w5127 & ~w5129) | (~w5127 & w16889) | (~w5129 & w16889);
assign w5343 = ~w5019 & ~w5022;
assign w5344 = ~w5021 & ~w5343;
assign w5345 = ~w5085 & ~w5089;
assign w5346 = ~w5088 & ~w5345;
assign w5347 = w5344 & w5346;
assign w5348 = ~w5344 & ~w5346;
assign w5349 = ~w5347 & ~w5348;
assign w5350 = pi02 & pi49;
assign w5351 = pi03 & pi48;
assign w5352 = pi04 & pi47;
assign w5353 = ~w5351 & ~w5352;
assign w5354 = pi04 & pi48;
assign w5355 = w4806 & w5354;
assign w5356 = ~w5353 & ~w5355;
assign w5357 = w5350 & ~w5356;
assign w5358 = ~w5350 & w5356;
assign w5359 = ~w5357 & ~w5358;
assign w5360 = ~w5349 & w5359;
assign w5361 = w5349 & ~w5359;
assign w5362 = ~w5360 & ~w5361;
assign w5363 = (~w5027 & ~w5029) | (~w5027 & w16890) | (~w5029 & w16890);
assign w5364 = w5362 & ~w5363;
assign w5365 = ~w5362 & w5363;
assign w5366 = ~w5364 & ~w5365;
assign w5367 = ~w5342 & w5366;
assign w5368 = w5342 & ~w5366;
assign w5369 = ~w5367 & ~w5368;
assign w5370 = ~w5341 & w5369;
assign w5371 = w5341 & ~w5369;
assign w5372 = ~w5370 & ~w5371;
assign w5373 = ~w4869 & ~w5077;
assign w5374 = ~w5076 & ~w5373;
assign w5375 = ~w5065 & ~w5069;
assign w5376 = ~w5068 & ~w5375;
assign w5377 = w5374 & w5376;
assign w5378 = ~w5374 & ~w5376;
assign w5379 = ~w5377 & ~w5378;
assign w5380 = ~w5010 & ~w5014;
assign w5381 = ~w5013 & ~w5380;
assign w5382 = ~w5379 & ~w5381;
assign w5383 = w5379 & w5381;
assign w5384 = ~w5382 & ~w5383;
assign w5385 = ~w5082 & ~w5094;
assign w5386 = ~w5384 & w5385;
assign w5387 = w5384 & ~w5385;
assign w5388 = ~w5386 & ~w5387;
assign w5389 = ~w4806 & ~w5036;
assign w5390 = ~w5035 & ~w5389;
assign w5391 = ~w5053 & ~w5057;
assign w5392 = ~w5056 & ~w5391;
assign w5393 = w5390 & w5392;
assign w5394 = ~w5390 & ~w5392;
assign w5395 = ~w5393 & ~w5394;
assign w5396 = ~w4948 & ~w5045;
assign w5397 = ~w5043 & ~w5396;
assign w5398 = ~w5395 & ~w5397;
assign w5399 = w5395 & w5397;
assign w5400 = ~w5398 & ~w5399;
assign w5401 = w5388 & w5400;
assign w5402 = ~w5388 & ~w5400;
assign w5403 = ~w5401 & ~w5402;
assign w5404 = w5372 & w5403;
assign w5405 = ~w5372 & ~w5403;
assign w5406 = ~w5404 & ~w5405;
assign w5407 = w5340 & w5406;
assign w5408 = ~w5340 & ~w5406;
assign w5409 = ~w5407 & ~w5408;
assign w5410 = w5319 & w5409;
assign w5411 = ~w5319 & ~w5409;
assign w5412 = ~w5410 & ~w5411;
assign w5413 = ~w5208 & w5412;
assign w5414 = w5208 & ~w5412;
assign w5415 = ~w5413 & ~w5414;
assign w5416 = ~w5207 & ~w5415;
assign w5417 = w5207 & w5415;
assign w5418 = ~w5416 & ~w5417;
assign w5419 = ~w5317 & ~w5410;
assign w5420 = ~w5311 & ~w5314;
assign w5421 = (~w5377 & ~w5379) | (~w5377 & w17109) | (~w5379 & w17109);
assign w5422 = (~w5393 & ~w5395) | (~w5393 & w16740) | (~w5395 & w16740);
assign w5423 = pi19 & pi33;
assign w5424 = pi03 & pi49;
assign w5425 = ~w5044 & ~w5424;
assign w5426 = pi03 & pi50;
assign w5427 = w5350 & w5426;
assign w5428 = ~w5425 & ~w5427;
assign w5429 = w5423 & ~w5428;
assign w5430 = ~w5423 & w5428;
assign w5431 = ~w5429 & ~w5430;
assign w5432 = ~w5422 & ~w5431;
assign w5433 = w5422 & w5431;
assign w5434 = ~w5432 & ~w5433;
assign w5435 = w5421 & ~w5434;
assign w5436 = ~w5421 & w5434;
assign w5437 = ~w5435 & ~w5436;
assign w5438 = ~w5364 & ~w5367;
assign w5439 = ~w5437 & w5438;
assign w5440 = w5437 & ~w5438;
assign w5441 = ~w5439 & ~w5440;
assign w5442 = ~w5290 & ~w5302;
assign w5443 = (~w5347 & ~w5349) | (~w5347 & w17110) | (~w5349 & w17110);
assign w5444 = pi25 & pi27;
assign w5445 = pi01 & pi51;
assign w5446 = ~w5444 & ~w5445;
assign w5447 = w5444 & w5445;
assign w5448 = ~w5446 & ~w5447;
assign w5449 = w5218 & w5448;
assign w5450 = ~w5218 & ~w5448;
assign w5451 = ~w5449 & ~w5450;
assign w5452 = ~w5293 & ~w5297;
assign w5453 = ~w5296 & ~w5452;
assign w5454 = w5451 & w5453;
assign w5455 = ~w5451 & ~w5453;
assign w5456 = ~w5454 & ~w5455;
assign w5457 = ~w5443 & w5456;
assign w5458 = w5443 & ~w5456;
assign w5459 = ~w5457 & ~w5458;
assign w5460 = ~w5442 & w5459;
assign w5461 = w5442 & ~w5459;
assign w5462 = ~w5460 & ~w5461;
assign w5463 = w5441 & w5462;
assign w5464 = ~w5441 & ~w5462;
assign w5465 = ~w5463 & ~w5464;
assign w5466 = ~w5420 & w5465;
assign w5467 = w5420 & ~w5465;
assign w5468 = ~w5466 & ~w5467;
assign w5469 = ~w5324 & ~w5328;
assign w5470 = (~w5214 & ~w5216) | (~w5214 & w16741) | (~w5216 & w16741);
assign w5471 = ~w5281 & ~w5285;
assign w5472 = ~w5284 & ~w5471;
assign w5473 = ~w5470 & w5472;
assign w5474 = w5470 & ~w5472;
assign w5475 = ~w5473 & ~w5474;
assign w5476 = pi00 & pi52;
assign w5477 = pi17 & pi35;
assign w5478 = ~w5354 & ~w5477;
assign w5479 = w5354 & w5477;
assign w5480 = ~w5478 & ~w5479;
assign w5481 = w5476 & ~w5480;
assign w5482 = ~w5476 & w5480;
assign w5483 = ~w5481 & ~w5482;
assign w5484 = ~w5475 & w5483;
assign w5485 = w5475 & ~w5483;
assign w5486 = ~w5484 & ~w5485;
assign w5487 = (~w5233 & ~w5235) | (~w5233 & w17111) | (~w5235 & w17111);
assign w5488 = w5486 & ~w5487;
assign w5489 = ~w5486 & w5487;
assign w5490 = ~w5488 & ~w5489;
assign w5491 = w5469 & ~w5490;
assign w5492 = ~w5469 & w5490;
assign w5493 = ~w5491 & ~w5492;
assign w5494 = ~w5305 & ~w5309;
assign w5495 = ~w5272 & ~w5276;
assign w5496 = ~w5275 & ~w5495;
assign w5497 = ~w5239 & ~w5243;
assign w5498 = ~w5242 & ~w5497;
assign w5499 = w5496 & w5498;
assign w5500 = ~w5496 & ~w5498;
assign w5501 = ~w5499 & ~w5500;
assign w5502 = ~w5248 & ~w5252;
assign w5503 = ~w5251 & ~w5502;
assign w5504 = ~w5501 & ~w5503;
assign w5505 = w5501 & w5503;
assign w5506 = ~w5504 & ~w5505;
assign w5507 = ~w5224 & ~w5228;
assign w5508 = ~w5227 & ~w5507;
assign w5509 = w5350 & ~w5353;
assign w5510 = ~w5355 & ~w5509;
assign w5511 = w5508 & ~w5510;
assign w5512 = ~w5508 & w5510;
assign w5513 = ~w5511 & ~w5512;
assign w5514 = ~w5260 & ~w5264;
assign w5515 = ~w5263 & ~w5514;
assign w5516 = ~w5513 & ~w5515;
assign w5517 = w5513 & w5515;
assign w5518 = ~w5516 & ~w5517;
assign w5519 = ~w5257 & ~w5269;
assign w5520 = ~w5518 & w5519;
assign w5521 = w5518 & ~w5519;
assign w5522 = ~w5520 & ~w5521;
assign w5523 = w5506 & w5522;
assign w5524 = ~w5506 & ~w5522;
assign w5525 = ~w5523 & ~w5524;
assign w5526 = ~w5494 & w5525;
assign w5527 = w5494 & ~w5525;
assign w5528 = ~w5526 & ~w5527;
assign w5529 = ~w5493 & ~w5528;
assign w5530 = w5493 & w5528;
assign w5531 = ~w5529 & ~w5530;
assign w5532 = ~w5468 & ~w5531;
assign w5533 = w5468 & w5531;
assign w5534 = ~w5532 & ~w5533;
assign w5535 = ~w5370 & ~w5404;
assign w5536 = (~w5332 & ~w5334) | (~w5332 & w17112) | (~w5334 & w17112);
assign w5537 = ~w5387 & ~w5401;
assign w5538 = pi10 & pi42;
assign w5539 = pi12 & pi40;
assign w5540 = pi11 & pi41;
assign w5541 = ~w5539 & ~w5540;
assign w5542 = pi12 & pi41;
assign w5543 = w5293 & w5542;
assign w5544 = ~w5541 & ~w5543;
assign w5545 = w5538 & ~w5544;
assign w5546 = ~w5538 & w5544;
assign w5547 = ~w5545 & ~w5546;
assign w5548 = pi05 & pi47;
assign w5549 = pi16 & pi36;
assign w5550 = pi06 & pi46;
assign w5551 = ~w5549 & ~w5550;
assign w5552 = w5549 & w5550;
assign w5553 = ~w5551 & ~w5552;
assign w5554 = w5548 & ~w5553;
assign w5555 = ~w5548 & w5553;
assign w5556 = ~w5554 & ~w5555;
assign w5557 = ~w5547 & ~w5556;
assign w5558 = w5547 & w5556;
assign w5559 = ~w5557 & ~w5558;
assign w5560 = pi15 & pi37;
assign w5561 = pi08 & pi44;
assign w5562 = pi07 & pi45;
assign w5563 = ~w5561 & ~w5562;
assign w5564 = pi08 & pi45;
assign w5565 = w5272 & w5564;
assign w5566 = ~w5563 & ~w5565;
assign w5567 = w5560 & ~w5566;
assign w5568 = ~w5560 & w5566;
assign w5569 = ~w5567 & ~w5568;
assign w5570 = w5559 & ~w5569;
assign w5571 = ~w5559 & w5569;
assign w5572 = ~w5570 & ~w5571;
assign w5573 = pi18 & pi34;
assign w5574 = pi20 & pi32;
assign w5575 = pi21 & pi31;
assign w5576 = ~w5574 & ~w5575;
assign w5577 = w5574 & w5575;
assign w5578 = ~w5576 & ~w5577;
assign w5579 = w5573 & ~w5578;
assign w5580 = ~w5573 & w5578;
assign w5581 = ~w5579 & ~w5580;
assign w5582 = pi22 & pi30;
assign w5583 = pi23 & pi29;
assign w5584 = pi24 & pi28;
assign w5585 = ~w5583 & ~w5584;
assign w5586 = w5583 & w5584;
assign w5587 = ~w5585 & ~w5586;
assign w5588 = w5582 & ~w5587;
assign w5589 = ~w5582 & w5587;
assign w5590 = ~w5588 & ~w5589;
assign w5591 = ~w5581 & ~w5590;
assign w5592 = w5581 & w5590;
assign w5593 = ~w5591 & ~w5592;
assign w5594 = pi14 & pi38;
assign w5595 = pi09 & pi43;
assign w5596 = pi13 & pi39;
assign w5597 = ~w5595 & ~w5596;
assign w5598 = w5595 & w5596;
assign w5599 = ~w5597 & ~w5598;
assign w5600 = w5594 & ~w5599;
assign w5601 = ~w5594 & w5599;
assign w5602 = ~w5600 & ~w5601;
assign w5603 = w5593 & ~w5602;
assign w5604 = ~w5593 & w5602;
assign w5605 = ~w5603 & ~w5604;
assign w5606 = w5572 & w5605;
assign w5607 = ~w5572 & ~w5605;
assign w5608 = ~w5606 & ~w5607;
assign w5609 = ~w5537 & w5608;
assign w5610 = w5537 & ~w5608;
assign w5611 = ~w5609 & ~w5610;
assign w5612 = ~w5536 & w5611;
assign w5613 = w5536 & ~w5611;
assign w5614 = ~w5612 & ~w5613;
assign w5615 = w5535 & ~w5614;
assign w5616 = ~w5535 & w5614;
assign w5617 = ~w5615 & ~w5616;
assign w5618 = ~w5338 & ~w5407;
assign w5619 = ~w5617 & w5618;
assign w5620 = w5617 & ~w5618;
assign w5621 = ~w5619 & ~w5620;
assign w5622 = w5534 & w5621;
assign w5623 = ~w5534 & ~w5621;
assign w5624 = ~w5622 & ~w5623;
assign w5625 = ~w5419 & w5624;
assign w5626 = w5419 & ~w5624;
assign w5627 = ~w5414 & ~w5626;
assign w5628 = (w5627 & w5207) | (w5627 & w16532) | (w5207 & w16532);
assign w5629 = ~w5625 & w5628;
assign w5630 = ~w5625 & ~w5626;
assign w5631 = w5207 & ~w5414;
assign w5632 = ~w5413 & ~w5630;
assign w5633 = ~w5631 & w5632;
assign w5634 = ~w5629 & ~w5633;
assign w5635 = ~w5625 & ~w5628;
assign w5636 = ~w5620 & ~w5622;
assign w5637 = ~w5466 & ~w5533;
assign w5638 = ~w5526 & ~w5530;
assign w5639 = (~w5432 & ~w5434) | (~w5432 & w16891) | (~w5434 & w16891);
assign w5640 = pi02 & pi51;
assign w5641 = ~w5426 & ~w5640;
assign w5642 = pi03 & pi51;
assign w5643 = w5044 & w5642;
assign w5644 = ~w5641 & ~w5643;
assign w5645 = w5447 & ~w5644;
assign w5646 = ~w5447 & w5644;
assign w5647 = ~w5645 & ~w5646;
assign w5648 = pi04 & pi49;
assign w5649 = pi17 & pi36;
assign w5650 = pi18 & pi35;
assign w5651 = ~w5649 & ~w5650;
assign w5652 = w5649 & w5650;
assign w5653 = ~w5651 & ~w5652;
assign w5654 = w5648 & ~w5653;
assign w5655 = ~w5648 & w5653;
assign w5656 = ~w5654 & ~w5655;
assign w5657 = ~w5647 & ~w5656;
assign w5658 = w5647 & w5656;
assign w5659 = ~w5657 & ~w5658;
assign w5660 = pi19 & pi34;
assign w5661 = pi21 & pi32;
assign w5662 = pi20 & pi33;
assign w5663 = ~w5661 & ~w5662;
assign w5664 = w5661 & w5662;
assign w5665 = ~w5663 & ~w5664;
assign w5666 = w5660 & ~w5665;
assign w5667 = ~w5660 & w5665;
assign w5668 = ~w5666 & ~w5667;
assign w5669 = w5659 & ~w5668;
assign w5670 = ~w5659 & w5668;
assign w5671 = ~w5669 & ~w5670;
assign w5672 = ~w5639 & w5671;
assign w5673 = w5639 & ~w5671;
assign w5674 = ~w5672 & ~w5673;
assign w5675 = pi06 & pi47;
assign w5676 = pi07 & pi46;
assign w5677 = pi15 & pi38;
assign w5678 = ~w5676 & ~w5677;
assign w5679 = w5676 & w5677;
assign w5680 = ~w5678 & ~w5679;
assign w5681 = w5675 & ~w5680;
assign w5682 = ~w5675 & w5680;
assign w5683 = ~w5681 & ~w5682;
assign w5684 = pi14 & pi39;
assign w5685 = pi09 & pi44;
assign w5686 = ~w5684 & ~w5685;
assign w5687 = w5684 & w5685;
assign w5688 = ~w5686 & ~w5687;
assign w5689 = w5564 & ~w5688;
assign w5690 = ~w5564 & w5688;
assign w5691 = ~w5689 & ~w5690;
assign w5692 = ~w5683 & ~w5691;
assign w5693 = w5683 & w5691;
assign w5694 = ~w5692 & ~w5693;
assign w5695 = pi00 & pi53;
assign w5696 = pi05 & pi48;
assign w5697 = pi16 & pi37;
assign w5698 = ~w5696 & ~w5697;
assign w5699 = w5696 & w5697;
assign w5700 = ~w5698 & ~w5699;
assign w5701 = w5695 & ~w5700;
assign w5702 = ~w5695 & w5700;
assign w5703 = ~w5701 & ~w5702;
assign w5704 = w5694 & ~w5703;
assign w5705 = ~w5694 & w5703;
assign w5706 = ~w5704 & ~w5705;
assign w5707 = ~w5674 & ~w5706;
assign w5708 = w5674 & w5706;
assign w5709 = ~w5707 & ~w5708;
assign w5710 = ~w5521 & ~w5523;
assign w5711 = ~w5457 & ~w5460;
assign w5712 = pi13 & pi40;
assign w5713 = pi10 & pi43;
assign w5714 = ~w5542 & ~w5713;
assign w5715 = w5542 & w5713;
assign w5716 = ~w5714 & ~w5715;
assign w5717 = w5712 & ~w5716;
assign w5718 = ~w5712 & w5716;
assign w5719 = ~w5717 & ~w5718;
assign w5720 = pi22 & pi31;
assign w5721 = pi24 & pi29;
assign w5722 = pi23 & pi30;
assign w5723 = ~w5721 & ~w5722;
assign w5724 = w5721 & w5722;
assign w5725 = ~w5723 & ~w5724;
assign w5726 = w5720 & ~w5725;
assign w5727 = ~w5720 & w5725;
assign w5728 = ~w5726 & ~w5727;
assign w5729 = ~w5719 & ~w5728;
assign w5730 = w5719 & w5728;
assign w5731 = ~w5729 & ~w5730;
assign w5732 = pi11 & pi42;
assign w5733 = pi26 & pi27;
assign w5734 = pi25 & pi28;
assign w5735 = ~w5733 & ~w5734;
assign w5736 = w5733 & w5734;
assign w5737 = ~w5735 & ~w5736;
assign w5738 = w5732 & ~w5737;
assign w5739 = ~w5732 & w5737;
assign w5740 = ~w5738 & ~w5739;
assign w5741 = w5731 & ~w5740;
assign w5742 = ~w5731 & w5740;
assign w5743 = ~w5741 & ~w5742;
assign w5744 = ~w5711 & w5743;
assign w5745 = w5711 & ~w5743;
assign w5746 = ~w5744 & ~w5745;
assign w5747 = ~w5710 & w5746;
assign w5748 = w5710 & ~w5746;
assign w5749 = ~w5747 & ~w5748;
assign w5750 = w5709 & w5749;
assign w5751 = ~w5709 & ~w5749;
assign w5752 = ~w5750 & ~w5751;
assign w5753 = ~w5638 & w5752;
assign w5754 = w5638 & ~w5752;
assign w5755 = ~w5753 & ~w5754;
assign w5756 = ~w5637 & w5755;
assign w5757 = w5637 & ~w5755;
assign w5758 = ~w5756 & ~w5757;
assign w5759 = ~w5476 & ~w5479;
assign w5760 = ~w5478 & ~w5759;
assign w5761 = w5423 & ~w5425;
assign w5762 = ~w5427 & ~w5761;
assign w5763 = w5760 & ~w5762;
assign w5764 = ~w5760 & w5762;
assign w5765 = ~w5763 & ~w5764;
assign w5766 = ~w5582 & ~w5586;
assign w5767 = ~w5585 & ~w5766;
assign w5768 = ~w5765 & ~w5767;
assign w5769 = w5765 & w5767;
assign w5770 = ~w5768 & ~w5769;
assign w5771 = (~w5591 & ~w5593) | (~w5591 & w16892) | (~w5593 & w16892);
assign w5772 = (~w5473 & ~w5475) | (~w5473 & w16893) | (~w5475 & w16893);
assign w5773 = ~w5771 & ~w5772;
assign w5774 = w5771 & w5772;
assign w5775 = ~w5773 & ~w5774;
assign w5776 = w5770 & w5775;
assign w5777 = ~w5770 & ~w5775;
assign w5778 = ~w5776 & ~w5777;
assign w5779 = ~w5573 & ~w5577;
assign w5780 = ~w5576 & ~w5779;
assign w5781 = ~w5548 & ~w5552;
assign w5782 = ~w5551 & ~w5781;
assign w5783 = w5780 & w5782;
assign w5784 = ~w5780 & ~w5782;
assign w5785 = ~w5783 & ~w5784;
assign w5786 = w5560 & ~w5563;
assign w5787 = ~w5565 & ~w5786;
assign w5788 = ~w5785 & w5787;
assign w5789 = w5785 & ~w5787;
assign w5790 = ~w5788 & ~w5789;
assign w5791 = ~w5557 & ~w5570;
assign w5792 = pi52 & w1542;
assign w5793 = pi01 & pi52;
assign w5794 = ~pi27 & ~w5793;
assign w5795 = ~w5792 & ~w5794;
assign w5796 = w5538 & ~w5541;
assign w5797 = ~w5543 & ~w5796;
assign w5798 = w5795 & ~w5797;
assign w5799 = ~w5795 & w5797;
assign w5800 = ~w5798 & ~w5799;
assign w5801 = ~w5594 & ~w5598;
assign w5802 = ~w5597 & ~w5801;
assign w5803 = w5800 & w5802;
assign w5804 = ~w5800 & ~w5802;
assign w5805 = ~w5803 & ~w5804;
assign w5806 = ~w5791 & w5805;
assign w5807 = w5791 & ~w5805;
assign w5808 = ~w5806 & ~w5807;
assign w5809 = ~w5790 & ~w5808;
assign w5810 = w5790 & w5808;
assign w5811 = ~w5809 & ~w5810;
assign w5812 = ~w5778 & ~w5811;
assign w5813 = w5778 & w5811;
assign w5814 = ~w5812 & ~w5813;
assign w5815 = (~w5440 & ~w5441) | (~w5440 & w17113) | (~w5441 & w17113);
assign w5816 = ~w5814 & w5815;
assign w5817 = w5814 & ~w5815;
assign w5818 = ~w5816 & ~w5817;
assign w5819 = ~w5606 & ~w5609;
assign w5820 = (~w5511 & ~w5513) | (~w5511 & w17114) | (~w5513 & w17114);
assign w5821 = (~w5499 & ~w5501) | (~w5499 & w16742) | (~w5501 & w16742);
assign w5822 = (~w5449 & ~w5451) | (~w5449 & w16894) | (~w5451 & w16894);
assign w5823 = ~w5821 & ~w5822;
assign w5824 = w5821 & w5822;
assign w5825 = ~w5823 & ~w5824;
assign w5826 = w5820 & ~w5825;
assign w5827 = ~w5820 & w5825;
assign w5828 = ~w5826 & ~w5827;
assign w5829 = ~w5488 & ~w5492;
assign w5830 = ~w5828 & w5829;
assign w5831 = w5828 & ~w5829;
assign w5832 = ~w5830 & ~w5831;
assign w5833 = ~w5819 & w5832;
assign w5834 = w5819 & ~w5832;
assign w5835 = ~w5833 & ~w5834;
assign w5836 = ~w5612 & ~w5616;
assign w5837 = ~w5835 & w5836;
assign w5838 = w5835 & ~w5836;
assign w5839 = ~w5837 & ~w5838;
assign w5840 = w5818 & w5839;
assign w5841 = ~w5818 & ~w5839;
assign w5842 = ~w5840 & ~w5841;
assign w5843 = w5758 & w5842;
assign w5844 = ~w5758 & ~w5842;
assign w5845 = ~w5843 & ~w5844;
assign w5846 = ~w5636 & w5845;
assign w5847 = w5636 & ~w5845;
assign w5848 = ~w5846 & ~w5847;
assign w5849 = w5635 & w5848;
assign w5850 = ~w5635 & ~w5848;
assign w5851 = ~w5849 & ~w5850;
assign w5852 = ~w5756 & ~w5843;
assign w5853 = ~w5750 & ~w5753;
assign w5854 = (~w5798 & ~w5800) | (~w5798 & w17115) | (~w5800 & w17115);
assign w5855 = (~w5783 & ~w5785) | (~w5783 & w16743) | (~w5785 & w16743);
assign w5856 = (~w5763 & ~w5765) | (~w5763 & w16744) | (~w5765 & w16744);
assign w5857 = ~w5855 & ~w5856;
assign w5858 = w5855 & w5856;
assign w5859 = ~w5857 & ~w5858;
assign w5860 = w5854 & ~w5859;
assign w5861 = ~w5854 & w5859;
assign w5862 = ~w5860 & ~w5861;
assign w5863 = (~w5672 & ~w5674) | (~w5672 & w17116) | (~w5674 & w17116);
assign w5864 = ~w5862 & w5863;
assign w5865 = w5862 & ~w5863;
assign w5866 = ~w5864 & ~w5865;
assign w5867 = ~w5695 & ~w5699;
assign w5868 = ~w5698 & ~w5867;
assign w5869 = ~w5675 & ~w5679;
assign w5870 = ~w5678 & ~w5869;
assign w5871 = w5868 & w5870;
assign w5872 = ~w5868 & ~w5870;
assign w5873 = ~w5871 & ~w5872;
assign w5874 = ~w5732 & ~w5736;
assign w5875 = ~w5735 & ~w5874;
assign w5876 = ~w5873 & ~w5875;
assign w5877 = w5873 & w5875;
assign w5878 = ~w5876 & ~w5877;
assign w5879 = ~w5648 & ~w5652;
assign w5880 = ~w5651 & ~w5879;
assign w5881 = ~w5660 & ~w5664;
assign w5882 = ~w5663 & ~w5881;
assign w5883 = w5880 & w5882;
assign w5884 = ~w5880 & ~w5882;
assign w5885 = ~w5883 & ~w5884;
assign w5886 = ~w5720 & ~w5724;
assign w5887 = ~w5723 & ~w5886;
assign w5888 = ~w5885 & ~w5887;
assign w5889 = w5885 & w5887;
assign w5890 = ~w5888 & ~w5889;
assign w5891 = ~w5692 & ~w5704;
assign w5892 = ~w5890 & w5891;
assign w5893 = w5890 & ~w5891;
assign w5894 = ~w5892 & ~w5893;
assign w5895 = w5878 & w5894;
assign w5896 = ~w5878 & ~w5894;
assign w5897 = ~w5895 & ~w5896;
assign w5898 = w5866 & w5897;
assign w5899 = ~w5866 & ~w5897;
assign w5900 = ~w5898 & ~w5899;
assign w5901 = ~w5853 & w5900;
assign w5902 = w5853 & ~w5900;
assign w5903 = ~w5901 & ~w5902;
assign w5904 = (~w5823 & ~w5825) | (~w5823 & w16895) | (~w5825 & w16895);
assign w5905 = pi13 & pi41;
assign w5906 = pi12 & pi42;
assign w5907 = pi11 & pi43;
assign w5908 = ~w5906 & ~w5907;
assign w5909 = pi12 & pi43;
assign w5910 = w5732 & w5909;
assign w5911 = ~w5908 & ~w5910;
assign w5912 = w5905 & ~w5911;
assign w5913 = ~w5905 & w5911;
assign w5914 = ~w5912 & ~w5913;
assign w5915 = pi20 & pi34;
assign w5916 = pi18 & pi36;
assign w5917 = pi05 & pi49;
assign w5918 = ~w5916 & ~w5917;
assign w5919 = w5916 & w5917;
assign w5920 = ~w5918 & ~w5919;
assign w5921 = w5915 & ~w5920;
assign w5922 = ~w5915 & w5920;
assign w5923 = ~w5921 & ~w5922;
assign w5924 = ~w5914 & ~w5923;
assign w5925 = w5914 & w5923;
assign w5926 = ~w5924 & ~w5925;
assign w5927 = pi17 & pi37;
assign w5928 = pi06 & pi48;
assign w5929 = pi16 & pi38;
assign w5930 = ~w5928 & ~w5929;
assign w5931 = w5928 & w5929;
assign w5932 = ~w5930 & ~w5931;
assign w5933 = w5927 & ~w5932;
assign w5934 = ~w5927 & w5932;
assign w5935 = ~w5933 & ~w5934;
assign w5936 = w5926 & ~w5935;
assign w5937 = ~w5926 & w5935;
assign w5938 = ~w5936 & ~w5937;
assign w5939 = ~w5904 & w5938;
assign w5940 = w5904 & ~w5938;
assign w5941 = ~w5939 & ~w5940;
assign w5942 = pi02 & pi52;
assign w5943 = pi04 & pi50;
assign w5944 = ~w5642 & ~w5943;
assign w5945 = pi04 & pi51;
assign w5946 = w5426 & w5945;
assign w5947 = ~w5944 & ~w5946;
assign w5948 = w5942 & ~w5947;
assign w5949 = ~w5942 & w5947;
assign w5950 = ~w5948 & ~w5949;
assign w5951 = pi07 & pi47;
assign w5952 = pi15 & pi39;
assign w5953 = pi08 & pi46;
assign w5954 = ~w5952 & ~w5953;
assign w5955 = w5952 & w5953;
assign w5956 = ~w5954 & ~w5955;
assign w5957 = w5951 & ~w5956;
assign w5958 = ~w5951 & w5956;
assign w5959 = ~w5957 & ~w5958;
assign w5960 = ~w5950 & ~w5959;
assign w5961 = w5950 & w5959;
assign w5962 = ~w5960 & ~w5961;
assign w5963 = pi09 & pi45;
assign w5964 = pi14 & pi40;
assign w5965 = pi10 & pi44;
assign w5966 = ~w5964 & ~w5965;
assign w5967 = w5964 & w5965;
assign w5968 = ~w5966 & ~w5967;
assign w5969 = w5963 & ~w5968;
assign w5970 = ~w5963 & w5968;
assign w5971 = ~w5969 & ~w5970;
assign w5972 = w5962 & ~w5971;
assign w5973 = ~w5962 & w5971;
assign w5974 = ~w5972 & ~w5973;
assign w5975 = ~w5941 & ~w5974;
assign w5976 = w5941 & w5974;
assign w5977 = ~w5975 & ~w5976;
assign w5978 = ~w5744 & ~w5747;
assign w5979 = ~w5564 & ~w5687;
assign w5980 = ~w5686 & ~w5979;
assign w5981 = w5447 & ~w5641;
assign w5982 = ~w5643 & ~w5981;
assign w5983 = w5980 & ~w5982;
assign w5984 = ~w5980 & w5982;
assign w5985 = ~w5983 & ~w5984;
assign w5986 = ~w5712 & ~w5715;
assign w5987 = ~w5714 & ~w5986;
assign w5988 = ~w5985 & ~w5987;
assign w5989 = w5985 & w5987;
assign w5990 = ~w5988 & ~w5989;
assign w5991 = (~w5729 & ~w5731) | (~w5729 & w16896) | (~w5731 & w16896);
assign w5992 = (~w5657 & ~w5659) | (~w5657 & w16897) | (~w5659 & w16897);
assign w5993 = ~w5991 & ~w5992;
assign w5994 = w5991 & w5992;
assign w5995 = ~w5993 & ~w5994;
assign w5996 = w5990 & w5995;
assign w5997 = ~w5990 & ~w5995;
assign w5998 = ~w5996 & ~w5997;
assign w5999 = ~w5978 & w5998;
assign w6000 = w5978 & ~w5998;
assign w6001 = ~w5999 & ~w6000;
assign w6002 = ~w5977 & ~w6001;
assign w6003 = w5977 & w6001;
assign w6004 = ~w6002 & ~w6003;
assign w6005 = ~w5903 & ~w6004;
assign w6006 = w5903 & w6004;
assign w6007 = ~w6005 & ~w6006;
assign w6008 = ~w5806 & ~w5810;
assign w6009 = (~w5773 & ~w5775) | (~w5773 & w17117) | (~w5775 & w17117);
assign w6010 = pi00 & pi54;
assign w6011 = w5792 & w6010;
assign w6012 = ~w5792 & ~w6010;
assign w6013 = ~w6011 & ~w6012;
assign w6014 = pi26 & pi28;
assign w6015 = pi01 & pi53;
assign w6016 = ~w6014 & ~w6015;
assign w6017 = w6014 & w6015;
assign w6018 = ~w6016 & ~w6017;
assign w6019 = w6013 & w6018;
assign w6020 = ~w6013 & ~w6018;
assign w6021 = ~w6019 & ~w6020;
assign w6022 = pi19 & pi35;
assign w6023 = pi21 & pi33;
assign w6024 = pi22 & pi32;
assign w6025 = ~w6023 & ~w6024;
assign w6026 = w6023 & w6024;
assign w6027 = ~w6025 & ~w6026;
assign w6028 = w6022 & ~w6027;
assign w6029 = ~w6022 & w6027;
assign w6030 = ~w6028 & ~w6029;
assign w6031 = pi23 & pi31;
assign w6032 = pi24 & pi30;
assign w6033 = pi25 & pi29;
assign w6034 = ~w6032 & ~w6033;
assign w6035 = w6032 & w6033;
assign w6036 = ~w6034 & ~w6035;
assign w6037 = w6031 & ~w6036;
assign w6038 = ~w6031 & w6036;
assign w6039 = ~w6037 & ~w6038;
assign w6040 = ~w6030 & ~w6039;
assign w6041 = w6030 & w6039;
assign w6042 = ~w6040 & ~w6041;
assign w6043 = w6021 & w6042;
assign w6044 = ~w6021 & ~w6042;
assign w6045 = ~w6043 & ~w6044;
assign w6046 = ~w6009 & w6045;
assign w6047 = w6009 & ~w6045;
assign w6048 = ~w6046 & ~w6047;
assign w6049 = ~w6008 & w6048;
assign w6050 = w6008 & ~w6048;
assign w6051 = ~w6049 & ~w6050;
assign w6052 = ~w5813 & ~w5817;
assign w6053 = ~w5831 & ~w5833;
assign w6054 = ~w6052 & ~w6053;
assign w6055 = w6052 & w6053;
assign w6056 = ~w6054 & ~w6055;
assign w6057 = ~w6051 & ~w6056;
assign w6058 = w6051 & w6056;
assign w6059 = ~w6057 & ~w6058;
assign w6060 = ~w5838 & ~w5840;
assign w6061 = w6059 & ~w6060;
assign w6062 = ~w6059 & w6060;
assign w6063 = ~w6061 & ~w6062;
assign w6064 = w6007 & w6063;
assign w6065 = ~w6007 & ~w6063;
assign w6066 = ~w6064 & ~w6065;
assign w6067 = ~w5852 & w6066;
assign w6068 = w5852 & ~w6066;
assign w6069 = ~w6067 & ~w6068;
assign w6070 = ~w5625 & ~w5846;
assign w6071 = (w5207 & w16534) | (w5207 & w16535) | (w16534 & w16535);
assign w6072 = w6069 & w6071;
assign w6073 = ~w6069 & ~w6071;
assign w6074 = ~w6072 & ~w6073;
assign w6075 = ~w6061 & ~w6064;
assign w6076 = ~w6054 & ~w6058;
assign w6077 = (~w6011 & ~w6013) | (~w6011 & w16745) | (~w6013 & w16745);
assign w6078 = ~w5951 & ~w5955;
assign w6079 = ~w5954 & ~w6078;
assign w6080 = ~w6077 & w6079;
assign w6081 = w6077 & ~w6079;
assign w6082 = ~w6080 & ~w6081;
assign w6083 = pi05 & pi50;
assign w6084 = pi18 & pi37;
assign w6085 = pi19 & pi36;
assign w6086 = ~w6084 & ~w6085;
assign w6087 = w6084 & w6085;
assign w6088 = ~w6086 & ~w6087;
assign w6089 = w6083 & ~w6088;
assign w6090 = ~w6083 & w6088;
assign w6091 = ~w6089 & ~w6090;
assign w6092 = ~w6082 & w6091;
assign w6093 = w6082 & ~w6091;
assign w6094 = ~w6092 & ~w6093;
assign w6095 = ~w5963 & ~w5967;
assign w6096 = ~w5966 & ~w6095;
assign w6097 = w5942 & ~w5944;
assign w6098 = ~w5946 & ~w6097;
assign w6099 = w6096 & ~w6098;
assign w6100 = ~w6096 & w6098;
assign w6101 = ~w6099 & ~w6100;
assign w6102 = ~w5915 & ~w5919;
assign w6103 = ~w5918 & ~w6102;
assign w6104 = ~w6101 & ~w6103;
assign w6105 = w6101 & w6103;
assign w6106 = ~w6104 & ~w6105;
assign w6107 = ~w6040 & ~w6043;
assign w6108 = ~w6106 & w6107;
assign w6109 = w6106 & ~w6107;
assign w6110 = ~w6108 & ~w6109;
assign w6111 = w6094 & w6110;
assign w6112 = ~w6094 & ~w6110;
assign w6113 = ~w6111 & ~w6112;
assign w6114 = pi54 & w1678;
assign w6115 = pi01 & pi54;
assign w6116 = ~pi28 & ~w6115;
assign w6117 = ~w6114 & ~w6116;
assign w6118 = ~w6017 & ~w6117;
assign w6119 = ~pi54 & w6017;
assign w6120 = ~w6118 & ~w6119;
assign w6121 = w5905 & ~w5908;
assign w6122 = ~w5910 & ~w6121;
assign w6123 = w6120 & ~w6122;
assign w6124 = ~w6120 & w6122;
assign w6125 = ~w6123 & ~w6124;
assign w6126 = (~w5871 & ~w5873) | (~w5871 & w16746) | (~w5873 & w16746);
assign w6127 = (~w5983 & ~w5985) | (~w5983 & w16747) | (~w5985 & w16747);
assign w6128 = ~w6126 & ~w6127;
assign w6129 = w6126 & w6127;
assign w6130 = ~w6128 & ~w6129;
assign w6131 = ~w6125 & ~w6130;
assign w6132 = w6125 & w6130;
assign w6133 = ~w6131 & ~w6132;
assign w6134 = (~w5939 & ~w5941) | (~w5939 & w17118) | (~w5941 & w17118);
assign w6135 = w6133 & ~w6134;
assign w6136 = ~w6133 & w6134;
assign w6137 = ~w6135 & ~w6136;
assign w6138 = w6113 & w6137;
assign w6139 = ~w6113 & ~w6137;
assign w6140 = ~w6138 & ~w6139;
assign w6141 = ~w6076 & w6140;
assign w6142 = w6076 & ~w6140;
assign w6143 = ~w6141 & ~w6142;
assign w6144 = ~w6046 & ~w6049;
assign w6145 = ~w6022 & ~w6026;
assign w6146 = ~w6025 & ~w6145;
assign w6147 = ~w6031 & ~w6035;
assign w6148 = ~w6034 & ~w6147;
assign w6149 = w6146 & w6148;
assign w6150 = ~w6146 & ~w6148;
assign w6151 = ~w6149 & ~w6150;
assign w6152 = ~w5927 & ~w5931;
assign w6153 = ~w5930 & ~w6152;
assign w6154 = ~w6151 & ~w6153;
assign w6155 = w6151 & w6153;
assign w6156 = ~w6154 & ~w6155;
assign w6157 = (~w5924 & ~w5926) | (~w5924 & w17119) | (~w5926 & w17119);
assign w6158 = (~w5960 & ~w5962) | (~w5960 & w17120) | (~w5962 & w17120);
assign w6159 = ~w6157 & ~w6158;
assign w6160 = w6157 & w6158;
assign w6161 = ~w6159 & ~w6160;
assign w6162 = w6156 & w6161;
assign w6163 = ~w6156 & ~w6161;
assign w6164 = ~w6162 & ~w6163;
assign w6165 = ~w6144 & w6164;
assign w6166 = w6144 & ~w6164;
assign w6167 = ~w6165 & ~w6166;
assign w6168 = (~w5857 & ~w5859) | (~w5857 & w16898) | (~w5859 & w16898);
assign w6169 = pi10 & pi45;
assign w6170 = pi13 & pi42;
assign w6171 = pi11 & pi44;
assign w6172 = ~w6170 & ~w6171;
assign w6173 = pi13 & pi44;
assign w6174 = w5732 & w6173;
assign w6175 = ~w6172 & ~w6174;
assign w6176 = w6169 & ~w6175;
assign w6177 = ~w6169 & w6175;
assign w6178 = ~w6176 & ~w6177;
assign w6179 = pi27 & pi28;
assign w6180 = pi26 & pi29;
assign w6181 = ~w6179 & ~w6180;
assign w6182 = w6179 & w6180;
assign w6183 = ~w6181 & ~w6182;
assign w6184 = w5909 & ~w6183;
assign w6185 = ~w5909 & w6183;
assign w6186 = ~w6184 & ~w6185;
assign w6187 = ~w6178 & ~w6186;
assign w6188 = w6178 & w6186;
assign w6189 = ~w6187 & ~w6188;
assign w6190 = pi16 & pi39;
assign w6191 = pi08 & pi47;
assign w6192 = pi07 & pi48;
assign w6193 = ~w6191 & ~w6192;
assign w6194 = pi08 & pi48;
assign w6195 = w5951 & w6194;
assign w6196 = ~w6193 & ~w6195;
assign w6197 = w6190 & ~w6196;
assign w6198 = ~w6190 & w6196;
assign w6199 = ~w6197 & ~w6198;
assign w6200 = w6189 & ~w6199;
assign w6201 = ~w6189 & w6199;
assign w6202 = ~w6200 & ~w6201;
assign w6203 = ~w6168 & w6202;
assign w6204 = w6168 & ~w6202;
assign w6205 = ~w6203 & ~w6204;
assign w6206 = pi00 & pi55;
assign w6207 = pi02 & pi53;
assign w6208 = ~w5945 & ~w6207;
assign w6209 = w5945 & w6207;
assign w6210 = ~w6208 & ~w6209;
assign w6211 = w6206 & ~w6210;
assign w6212 = ~w6206 & w6210;
assign w6213 = ~w6211 & ~w6212;
assign w6214 = pi20 & pi35;
assign w6215 = pi22 & pi33;
assign w6216 = pi21 & pi34;
assign w6217 = ~w6215 & ~w6216;
assign w6218 = w6215 & w6216;
assign w6219 = ~w6217 & ~w6218;
assign w6220 = w6214 & ~w6219;
assign w6221 = ~w6214 & w6219;
assign w6222 = ~w6220 & ~w6221;
assign w6223 = ~w6213 & ~w6222;
assign w6224 = w6213 & w6222;
assign w6225 = ~w6223 & ~w6224;
assign w6226 = pi23 & pi32;
assign w6227 = pi25 & pi30;
assign w6228 = pi24 & pi31;
assign w6229 = ~w6227 & ~w6228;
assign w6230 = w6227 & w6228;
assign w6231 = ~w6229 & ~w6230;
assign w6232 = w6226 & ~w6231;
assign w6233 = ~w6226 & w6231;
assign w6234 = ~w6232 & ~w6233;
assign w6235 = w6225 & ~w6234;
assign w6236 = ~w6225 & w6234;
assign w6237 = ~w6235 & ~w6236;
assign w6238 = w6205 & w6237;
assign w6239 = ~w6205 & ~w6237;
assign w6240 = ~w6238 & ~w6239;
assign w6241 = w6167 & w6240;
assign w6242 = ~w6167 & ~w6240;
assign w6243 = ~w6241 & ~w6242;
assign w6244 = ~w6143 & ~w6243;
assign w6245 = w6143 & w6243;
assign w6246 = ~w6244 & ~w6245;
assign w6247 = ~w5901 & ~w6006;
assign w6248 = ~w5999 & ~w6003;
assign w6249 = ~w5865 & ~w5898;
assign w6250 = ~w5893 & ~w5895;
assign w6251 = (~w5883 & ~w5885) | (~w5883 & w16748) | (~w5885 & w16748);
assign w6252 = pi15 & pi40;
assign w6253 = pi14 & pi41;
assign w6254 = pi09 & pi46;
assign w6255 = ~w6253 & ~w6254;
assign w6256 = w6253 & w6254;
assign w6257 = ~w6255 & ~w6256;
assign w6258 = w6252 & ~w6257;
assign w6259 = ~w6252 & w6257;
assign w6260 = ~w6258 & ~w6259;
assign w6261 = pi03 & pi52;
assign w6262 = pi06 & pi49;
assign w6263 = pi17 & pi38;
assign w6264 = ~w6262 & ~w6263;
assign w6265 = w6262 & w6263;
assign w6266 = ~w6264 & ~w6265;
assign w6267 = w6261 & ~w6266;
assign w6268 = ~w6261 & w6266;
assign w6269 = ~w6267 & ~w6268;
assign w6270 = ~w6260 & ~w6269;
assign w6271 = w6260 & w6269;
assign w6272 = ~w6270 & ~w6271;
assign w6273 = w6251 & ~w6272;
assign w6274 = ~w6251 & w6272;
assign w6275 = ~w6273 & ~w6274;
assign w6276 = (~w5993 & ~w5995) | (~w5993 & w17121) | (~w5995 & w17121);
assign w6277 = ~w6275 & w6276;
assign w6278 = w6275 & ~w6276;
assign w6279 = ~w6277 & ~w6278;
assign w6280 = ~w6250 & w6279;
assign w6281 = w6250 & ~w6279;
assign w6282 = ~w6280 & ~w6281;
assign w6283 = ~w6249 & w6282;
assign w6284 = w6249 & ~w6282;
assign w6285 = ~w6283 & ~w6284;
assign w6286 = ~w6248 & w6285;
assign w6287 = w6248 & ~w6285;
assign w6288 = ~w6286 & ~w6287;
assign w6289 = ~w6247 & w6288;
assign w6290 = w6247 & ~w6288;
assign w6291 = ~w6289 & ~w6290;
assign w6292 = w6246 & w6291;
assign w6293 = ~w6246 & ~w6291;
assign w6294 = ~w6292 & ~w6293;
assign w6295 = ~w6075 & w6294;
assign w6296 = w6075 & ~w6294;
assign w6297 = ~w6295 & ~w6296;
assign w6298 = (~w5207 & w16536) | (~w5207 & w16537) | (w16536 & w16537);
assign w6299 = ~w6068 & ~w6298;
assign w6300 = w6297 & w6299;
assign w6301 = ~w6297 & ~w6299;
assign w6302 = ~w6300 & ~w6301;
assign w6303 = ~w6289 & ~w6292;
assign w6304 = ~w6278 & ~w6280;
assign w6305 = ~w6214 & ~w6218;
assign w6306 = ~w6217 & ~w6305;
assign w6307 = ~w6226 & ~w6230;
assign w6308 = ~w6229 & ~w6307;
assign w6309 = w6306 & w6308;
assign w6310 = ~w6306 & ~w6308;
assign w6311 = ~w6309 & ~w6310;
assign w6312 = ~w6261 & ~w6265;
assign w6313 = ~w6264 & ~w6312;
assign w6314 = ~w6311 & ~w6313;
assign w6315 = w6311 & w6313;
assign w6316 = ~w6314 & ~w6315;
assign w6317 = (~w6187 & ~w6189) | (~w6187 & w16899) | (~w6189 & w16899);
assign w6318 = pi27 & pi29;
assign w6319 = pi01 & pi55;
assign w6320 = ~w6318 & ~w6319;
assign w6321 = w6318 & w6319;
assign w6322 = ~w6320 & ~w6321;
assign w6323 = ~w5909 & ~w6182;
assign w6324 = ~w6181 & ~w6323;
assign w6325 = w6322 & w6324;
assign w6326 = ~w6322 & ~w6324;
assign w6327 = ~w6325 & ~w6326;
assign w6328 = w6169 & ~w6172;
assign w6329 = ~w6174 & ~w6328;
assign w6330 = w6327 & ~w6329;
assign w6331 = ~w6327 & w6329;
assign w6332 = ~w6330 & ~w6331;
assign w6333 = ~w6317 & w6332;
assign w6334 = w6317 & ~w6332;
assign w6335 = ~w6333 & ~w6334;
assign w6336 = w6316 & w6335;
assign w6337 = ~w6316 & ~w6335;
assign w6338 = ~w6336 & ~w6337;
assign w6339 = ~w6304 & w6338;
assign w6340 = w6304 & ~w6338;
assign w6341 = ~w6339 & ~w6340;
assign w6342 = w6190 & ~w6193;
assign w6343 = ~w6195 & ~w6342;
assign w6344 = pi00 & pi56;
assign w6345 = pi02 & pi54;
assign w6346 = ~w6344 & ~w6345;
assign w6347 = pi02 & pi56;
assign w6348 = w6010 & w6347;
assign w6349 = ~w6346 & ~w6348;
assign w6350 = w6114 & ~w6349;
assign w6351 = ~w6114 & w6349;
assign w6352 = ~w6350 & ~w6351;
assign w6353 = ~w6343 & ~w6352;
assign w6354 = w6343 & w6352;
assign w6355 = ~w6353 & ~w6354;
assign w6356 = pi03 & pi53;
assign w6357 = pi19 & pi37;
assign w6358 = pi04 & pi52;
assign w6359 = ~w6357 & ~w6358;
assign w6360 = w6357 & w6358;
assign w6361 = ~w6359 & ~w6360;
assign w6362 = w6356 & ~w6361;
assign w6363 = ~w6356 & w6361;
assign w6364 = ~w6362 & ~w6363;
assign w6365 = ~w6355 & w6364;
assign w6366 = w6355 & ~w6364;
assign w6367 = ~w6365 & ~w6366;
assign w6368 = pi11 & pi45;
assign w6369 = pi13 & pi43;
assign w6370 = pi12 & pi44;
assign w6371 = ~w6369 & ~w6370;
assign w6372 = w5909 & w6173;
assign w6373 = ~w6371 & ~w6372;
assign w6374 = w6368 & ~w6373;
assign w6375 = ~w6368 & w6373;
assign w6376 = ~w6374 & ~w6375;
assign w6377 = pi06 & pi50;
assign w6378 = pi07 & pi49;
assign w6379 = pi17 & pi39;
assign w6380 = ~w6378 & ~w6379;
assign w6381 = w6378 & w6379;
assign w6382 = ~w6380 & ~w6381;
assign w6383 = w6377 & ~w6382;
assign w6384 = ~w6377 & w6382;
assign w6385 = ~w6383 & ~w6384;
assign w6386 = ~w6376 & ~w6385;
assign w6387 = w6376 & w6385;
assign w6388 = ~w6386 & ~w6387;
assign w6389 = pi16 & pi40;
assign w6390 = pi15 & pi41;
assign w6391 = ~w6194 & ~w6390;
assign w6392 = w6194 & w6390;
assign w6393 = ~w6391 & ~w6392;
assign w6394 = w6389 & ~w6393;
assign w6395 = ~w6389 & w6393;
assign w6396 = ~w6394 & ~w6395;
assign w6397 = w6388 & ~w6396;
assign w6398 = ~w6388 & w6396;
assign w6399 = ~w6397 & ~w6398;
assign w6400 = pi20 & pi36;
assign w6401 = pi22 & pi34;
assign w6402 = pi23 & pi33;
assign w6403 = ~w6401 & ~w6402;
assign w6404 = w6401 & w6402;
assign w6405 = ~w6403 & ~w6404;
assign w6406 = w6400 & ~w6405;
assign w6407 = ~w6400 & w6405;
assign w6408 = ~w6406 & ~w6407;
assign w6409 = pi24 & pi32;
assign w6410 = pi25 & pi31;
assign w6411 = pi26 & pi30;
assign w6412 = ~w6410 & ~w6411;
assign w6413 = w6410 & w6411;
assign w6414 = ~w6412 & ~w6413;
assign w6415 = w6409 & ~w6414;
assign w6416 = ~w6409 & w6414;
assign w6417 = ~w6415 & ~w6416;
assign w6418 = ~w6408 & ~w6417;
assign w6419 = w6408 & w6417;
assign w6420 = ~w6418 & ~w6419;
assign w6421 = pi09 & pi47;
assign w6422 = pi14 & pi42;
assign w6423 = pi10 & pi46;
assign w6424 = ~w6422 & ~w6423;
assign w6425 = w6422 & w6423;
assign w6426 = ~w6424 & ~w6425;
assign w6427 = w6421 & ~w6426;
assign w6428 = ~w6421 & w6426;
assign w6429 = ~w6427 & ~w6428;
assign w6430 = w6420 & ~w6429;
assign w6431 = ~w6420 & w6429;
assign w6432 = ~w6430 & ~w6431;
assign w6433 = w6399 & w6432;
assign w6434 = ~w6399 & ~w6432;
assign w6435 = ~w6433 & ~w6434;
assign w6436 = w6367 & w6435;
assign w6437 = ~w6367 & ~w6435;
assign w6438 = ~w6436 & ~w6437;
assign w6439 = ~w6341 & ~w6438;
assign w6440 = w6341 & w6438;
assign w6441 = ~w6439 & ~w6440;
assign w6442 = ~w6283 & ~w6286;
assign w6443 = ~w6083 & ~w6087;
assign w6444 = ~w6086 & ~w6443;
assign w6445 = ~w6206 & ~w6209;
assign w6446 = ~w6208 & ~w6445;
assign w6447 = w6444 & w6446;
assign w6448 = ~w6444 & ~w6446;
assign w6449 = ~w6447 & ~w6448;
assign w6450 = ~w6252 & ~w6256;
assign w6451 = ~w6255 & ~w6450;
assign w6452 = ~w6449 & ~w6451;
assign w6453 = w6449 & w6451;
assign w6454 = ~w6452 & ~w6453;
assign w6455 = ~w6270 & ~w6274;
assign w6456 = ~w6454 & w6455;
assign w6457 = w6454 & ~w6455;
assign w6458 = ~w6456 & ~w6457;
assign w6459 = (~w6128 & ~w6130) | (~w6128 & w16900) | (~w6130 & w16900);
assign w6460 = ~w6458 & w6459;
assign w6461 = w6458 & ~w6459;
assign w6462 = ~w6460 & ~w6461;
assign w6463 = (~w6223 & ~w6225) | (~w6223 & w17753) | (~w6225 & w17753);
assign w6464 = (~w6149 & ~w6151) | (~w6149 & w17122) | (~w6151 & w17122);
assign w6465 = (~w6080 & ~w6082) | (~w6080 & w16901) | (~w6082 & w16901);
assign w6466 = ~w6464 & ~w6465;
assign w6467 = w6464 & w6465;
assign w6468 = ~w6466 & ~w6467;
assign w6469 = w6463 & ~w6468;
assign w6470 = ~w6463 & w6468;
assign w6471 = ~w6469 & ~w6470;
assign w6472 = (~w6203 & ~w6205) | (~w6203 & w17123) | (~w6205 & w17123);
assign w6473 = w6471 & ~w6472;
assign w6474 = ~w6471 & w6472;
assign w6475 = ~w6473 & ~w6474;
assign w6476 = w6462 & w6475;
assign w6477 = ~w6462 & ~w6475;
assign w6478 = ~w6476 & ~w6477;
assign w6479 = ~w6442 & w6478;
assign w6480 = w6442 & ~w6478;
assign w6481 = ~w6479 & ~w6480;
assign w6482 = w6441 & w6481;
assign w6483 = ~w6441 & ~w6481;
assign w6484 = ~w6482 & ~w6483;
assign w6485 = ~w6109 & ~w6111;
assign w6486 = (~w6099 & ~w6101) | (~w6099 & w17124) | (~w6101 & w17124);
assign w6487 = (~w6119 & ~w6120) | (~w6119 & w16902) | (~w6120 & w16902);
assign w6488 = pi21 & pi35;
assign w6489 = pi05 & pi51;
assign w6490 = pi18 & pi38;
assign w6491 = ~w6489 & ~w6490;
assign w6492 = w6489 & w6490;
assign w6493 = ~w6491 & ~w6492;
assign w6494 = w6488 & ~w6493;
assign w6495 = ~w6488 & w6493;
assign w6496 = ~w6494 & ~w6495;
assign w6497 = ~w6487 & ~w6496;
assign w6498 = w6487 & w6496;
assign w6499 = ~w6497 & ~w6498;
assign w6500 = w6486 & ~w6499;
assign w6501 = ~w6486 & w6499;
assign w6502 = ~w6500 & ~w6501;
assign w6503 = (~w6159 & ~w6161) | (~w6159 & w17754) | (~w6161 & w17754);
assign w6504 = ~w6502 & w6503;
assign w6505 = w6502 & ~w6503;
assign w6506 = ~w6504 & ~w6505;
assign w6507 = w6485 & ~w6506;
assign w6508 = ~w6485 & w6506;
assign w6509 = ~w6507 & ~w6508;
assign w6510 = ~w6135 & ~w6138;
assign w6511 = ~w6509 & w6510;
assign w6512 = w6509 & ~w6510;
assign w6513 = ~w6511 & ~w6512;
assign w6514 = ~w6165 & ~w6241;
assign w6515 = ~w6513 & w6514;
assign w6516 = w6513 & ~w6514;
assign w6517 = ~w6515 & ~w6516;
assign w6518 = ~w6141 & ~w6245;
assign w6519 = w6517 & ~w6518;
assign w6520 = ~w6517 & w6518;
assign w6521 = ~w6519 & ~w6520;
assign w6522 = w6484 & w6521;
assign w6523 = ~w6484 & ~w6521;
assign w6524 = ~w6522 & ~w6523;
assign w6525 = ~w6303 & w6524;
assign w6526 = w6303 & ~w6524;
assign w6527 = ~w6525 & ~w6526;
assign w6528 = ~w6068 & ~w6296;
assign w6529 = ~w6298 & w6528;
assign w6530 = ~w6295 & ~w6529;
assign w6531 = w6527 & w6530;
assign w6532 = ~w6527 & ~w6530;
assign w6533 = ~w6531 & ~w6532;
assign w6534 = ~w6519 & ~w6522;
assign w6535 = ~w6512 & ~w6516;
assign w6536 = (~w6418 & ~w6420) | (~w6418 & w17755) | (~w6420 & w17755);
assign w6537 = (~w6325 & ~w6327) | (~w6325 & w17125) | (~w6327 & w17125);
assign w6538 = (~w6353 & ~w6355) | (~w6353 & w16903) | (~w6355 & w16903);
assign w6539 = ~w6537 & ~w6538;
assign w6540 = w6537 & w6538;
assign w6541 = ~w6539 & ~w6540;
assign w6542 = w6536 & ~w6541;
assign w6543 = ~w6536 & w6541;
assign w6544 = ~w6542 & ~w6543;
assign w6545 = ~w6433 & ~w6436;
assign w6546 = ~w6544 & w6545;
assign w6547 = w6544 & ~w6545;
assign w6548 = ~w6546 & ~w6547;
assign w6549 = (~w6386 & ~w6388) | (~w6386 & w17756) | (~w6388 & w17756);
assign w6550 = ~w6389 & ~w6392;
assign w6551 = ~w6391 & ~w6550;
assign w6552 = ~w6409 & ~w6413;
assign w6553 = ~w6412 & ~w6552;
assign w6554 = w6551 & w6553;
assign w6555 = ~w6551 & ~w6553;
assign w6556 = ~w6554 & ~w6555;
assign w6557 = ~w6377 & ~w6381;
assign w6558 = ~w6380 & ~w6557;
assign w6559 = ~w6556 & ~w6558;
assign w6560 = w6556 & w6558;
assign w6561 = ~w6559 & ~w6560;
assign w6562 = ~w6400 & ~w6404;
assign w6563 = ~w6403 & ~w6562;
assign w6564 = ~w6356 & ~w6360;
assign w6565 = ~w6359 & ~w6564;
assign w6566 = w6563 & w6565;
assign w6567 = ~w6563 & ~w6565;
assign w6568 = ~w6566 & ~w6567;
assign w6569 = ~w6114 & ~w6348;
assign w6570 = ~w6346 & ~w6569;
assign w6571 = ~w6568 & ~w6570;
assign w6572 = w6568 & w6570;
assign w6573 = ~w6571 & ~w6572;
assign w6574 = w6561 & w6573;
assign w6575 = ~w6561 & ~w6573;
assign w6576 = ~w6574 & ~w6575;
assign w6577 = ~w6549 & w6576;
assign w6578 = w6549 & ~w6576;
assign w6579 = ~w6577 & ~w6578;
assign w6580 = w6548 & w6579;
assign w6581 = ~w6548 & ~w6579;
assign w6582 = ~w6580 & ~w6581;
assign w6583 = ~w6535 & w6582;
assign w6584 = w6535 & ~w6582;
assign w6585 = ~w6583 & ~w6584;
assign w6586 = ~w6505 & ~w6508;
assign w6587 = ~w6421 & ~w6425;
assign w6588 = ~w6424 & ~w6587;
assign w6589 = ~w6488 & ~w6492;
assign w6590 = ~w6491 & ~w6589;
assign w6591 = w6588 & w6590;
assign w6592 = ~w6588 & ~w6590;
assign w6593 = ~w6591 & ~w6592;
assign w6594 = w6368 & ~w6371;
assign w6595 = ~w6372 & ~w6594;
assign w6596 = ~w6593 & w6595;
assign w6597 = w6593 & ~w6595;
assign w6598 = ~w6596 & ~w6597;
assign w6599 = (~w6497 & ~w6499) | (~w6497 & w17126) | (~w6499 & w17126);
assign w6600 = ~w6598 & w6599;
assign w6601 = w6598 & ~w6599;
assign w6602 = ~w6600 & ~w6601;
assign w6603 = pi21 & pi36;
assign w6604 = pi23 & pi34;
assign w6605 = pi22 & pi35;
assign w6606 = ~w6604 & ~w6605;
assign w6607 = pi23 & pi35;
assign w6608 = w6401 & w6607;
assign w6609 = ~w6606 & ~w6608;
assign w6610 = w6603 & ~w6609;
assign w6611 = ~w6603 & w6609;
assign w6612 = ~w6610 & ~w6611;
assign w6613 = pi07 & pi50;
assign w6614 = pi08 & pi49;
assign w6615 = pi16 & pi41;
assign w6616 = ~w6614 & ~w6615;
assign w6617 = w6614 & w6615;
assign w6618 = ~w6616 & ~w6617;
assign w6619 = w6613 & ~w6618;
assign w6620 = ~w6613 & w6618;
assign w6621 = ~w6619 & ~w6620;
assign w6622 = ~w6612 & ~w6621;
assign w6623 = w6612 & w6621;
assign w6624 = ~w6622 & ~w6623;
assign w6625 = pi24 & pi33;
assign w6626 = pi26 & pi31;
assign w6627 = pi25 & pi32;
assign w6628 = ~w6626 & ~w6627;
assign w6629 = w6626 & w6627;
assign w6630 = ~w6628 & ~w6629;
assign w6631 = w6625 & ~w6630;
assign w6632 = ~w6625 & w6630;
assign w6633 = ~w6631 & ~w6632;
assign w6634 = w6624 & ~w6633;
assign w6635 = ~w6624 & w6633;
assign w6636 = ~w6634 & ~w6635;
assign w6637 = w6602 & w6636;
assign w6638 = ~w6602 & ~w6636;
assign w6639 = ~w6637 & ~w6638;
assign w6640 = ~w6586 & w6639;
assign w6641 = w6586 & ~w6639;
assign w6642 = ~w6640 & ~w6641;
assign w6643 = (~w6466 & ~w6468) | (~w6466 & w17127) | (~w6468 & w17127);
assign w6644 = pi05 & pi52;
assign w6645 = pi20 & pi37;
assign w6646 = pi19 & pi38;
assign w6647 = ~w6645 & ~w6646;
assign w6648 = pi20 & pi38;
assign w6649 = w6357 & w6648;
assign w6650 = ~w6647 & ~w6649;
assign w6651 = w6644 & ~w6650;
assign w6652 = ~w6644 & w6650;
assign w6653 = ~w6651 & ~w6652;
assign w6654 = pi03 & pi54;
assign w6655 = pi04 & pi53;
assign w6656 = pi02 & pi55;
assign w6657 = ~w6655 & ~w6656;
assign w6658 = w6655 & w6656;
assign w6659 = ~w6657 & ~w6658;
assign w6660 = w6654 & ~w6659;
assign w6661 = ~w6654 & w6659;
assign w6662 = ~w6660 & ~w6661;
assign w6663 = ~w6653 & ~w6662;
assign w6664 = w6653 & w6662;
assign w6665 = ~w6663 & ~w6664;
assign w6666 = pi15 & pi42;
assign w6667 = pi10 & pi47;
assign w6668 = pi09 & pi48;
assign w6669 = ~w6667 & ~w6668;
assign w6670 = pi10 & pi48;
assign w6671 = w6421 & w6670;
assign w6672 = ~w6669 & ~w6671;
assign w6673 = w6666 & ~w6672;
assign w6674 = ~w6666 & w6672;
assign w6675 = ~w6673 & ~w6674;
assign w6676 = w6665 & ~w6675;
assign w6677 = ~w6665 & w6675;
assign w6678 = ~w6676 & ~w6677;
assign w6679 = pi14 & pi43;
assign w6680 = pi11 & pi46;
assign w6681 = ~w6173 & ~w6680;
assign w6682 = pi13 & pi46;
assign w6683 = w6171 & w6682;
assign w6684 = ~w6681 & ~w6683;
assign w6685 = w6679 & ~w6684;
assign w6686 = ~w6679 & w6684;
assign w6687 = ~w6685 & ~w6686;
assign w6688 = pi12 & pi45;
assign w6689 = pi28 & pi29;
assign w6690 = pi27 & pi30;
assign w6691 = ~w6689 & ~w6690;
assign w6692 = w6689 & w6690;
assign w6693 = ~w6691 & ~w6692;
assign w6694 = w6688 & ~w6693;
assign w6695 = ~w6688 & w6693;
assign w6696 = ~w6694 & ~w6695;
assign w6697 = ~w6687 & ~w6696;
assign w6698 = w6687 & w6696;
assign w6699 = ~w6697 & ~w6698;
assign w6700 = pi18 & pi39;
assign w6701 = pi06 & pi51;
assign w6702 = pi17 & pi40;
assign w6703 = ~w6701 & ~w6702;
assign w6704 = w6701 & w6702;
assign w6705 = ~w6703 & ~w6704;
assign w6706 = w6700 & ~w6705;
assign w6707 = ~w6700 & w6705;
assign w6708 = ~w6706 & ~w6707;
assign w6709 = w6699 & ~w6708;
assign w6710 = ~w6699 & w6708;
assign w6711 = ~w6709 & ~w6710;
assign w6712 = w6678 & w6711;
assign w6713 = ~w6678 & ~w6711;
assign w6714 = ~w6712 & ~w6713;
assign w6715 = ~w6643 & w6714;
assign w6716 = w6643 & ~w6714;
assign w6717 = ~w6715 & ~w6716;
assign w6718 = w6642 & w6717;
assign w6719 = ~w6642 & ~w6717;
assign w6720 = ~w6718 & ~w6719;
assign w6721 = ~w6585 & ~w6720;
assign w6722 = w6585 & w6720;
assign w6723 = ~w6721 & ~w6722;
assign w6724 = ~w6479 & ~w6482;
assign w6725 = ~w6339 & ~w6440;
assign w6726 = ~w6473 & ~w6476;
assign w6727 = (~w6447 & ~w6449) | (~w6447 & w17128) | (~w6449 & w17128);
assign w6728 = (~w6309 & ~w6311) | (~w6309 & w16749) | (~w6311 & w16749);
assign w6729 = pi00 & pi57;
assign w6730 = w6321 & w6729;
assign w6731 = ~w6321 & ~w6729;
assign w6732 = ~w6730 & ~w6731;
assign w6733 = pi01 & pi56;
assign w6734 = pi29 & w6733;
assign w6735 = ~pi29 & ~w6733;
assign w6736 = ~w6734 & ~w6735;
assign w6737 = w6732 & w6736;
assign w6738 = ~w6732 & ~w6736;
assign w6739 = ~w6737 & ~w6738;
assign w6740 = ~w6728 & w6739;
assign w6741 = w6728 & ~w6739;
assign w6742 = ~w6740 & ~w6741;
assign w6743 = w6727 & ~w6742;
assign w6744 = ~w6727 & w6742;
assign w6745 = ~w6743 & ~w6744;
assign w6746 = (~w6457 & ~w6458) | (~w6457 & w16904) | (~w6458 & w16904);
assign w6747 = (~w6333 & ~w6335) | (~w6333 & w17129) | (~w6335 & w17129);
assign w6748 = ~w6746 & ~w6747;
assign w6749 = w6746 & w6747;
assign w6750 = ~w6748 & ~w6749;
assign w6751 = w6745 & w6750;
assign w6752 = ~w6745 & ~w6750;
assign w6753 = ~w6751 & ~w6752;
assign w6754 = ~w6726 & w6753;
assign w6755 = w6726 & ~w6753;
assign w6756 = ~w6754 & ~w6755;
assign w6757 = ~w6725 & w6756;
assign w6758 = w6725 & ~w6756;
assign w6759 = ~w6757 & ~w6758;
assign w6760 = ~w6724 & w6759;
assign w6761 = w6724 & ~w6759;
assign w6762 = ~w6760 & ~w6761;
assign w6763 = w6723 & w6762;
assign w6764 = ~w6723 & ~w6762;
assign w6765 = ~w6763 & ~w6764;
assign w6766 = ~w6534 & w6765;
assign w6767 = w6534 & ~w6765;
assign w6768 = ~w6766 & ~w6767;
assign w6769 = ~w6295 & ~w6525;
assign w6770 = (~w6298 & w16539) | (~w6298 & w16540) | (w16539 & w16540);
assign w6771 = w6768 & w6770;
assign w6772 = ~w6768 & ~w6770;
assign w6773 = ~w6771 & ~w6772;
assign w6774 = ~w6760 & ~w6763;
assign w6775 = ~w6583 & ~w6722;
assign w6776 = ~w6547 & ~w6580;
assign w6777 = (~w6601 & ~w6602) | (~w6601 & w17757) | (~w6602 & w17757);
assign w6778 = (~w6554 & ~w6556) | (~w6554 & w17130) | (~w6556 & w17130);
assign w6779 = (~w6591 & ~w6593) | (~w6591 & w16750) | (~w6593 & w16750);
assign w6780 = (~w6566 & ~w6568) | (~w6566 & w16751) | (~w6568 & w16751);
assign w6781 = ~w6779 & ~w6780;
assign w6782 = w6779 & w6780;
assign w6783 = ~w6781 & ~w6782;
assign w6784 = w6778 & ~w6783;
assign w6785 = ~w6778 & w6783;
assign w6786 = ~w6784 & ~w6785;
assign w6787 = (~w6574 & ~w6576) | (~w6574 & w17131) | (~w6576 & w17131);
assign w6788 = ~w6786 & w6787;
assign w6789 = w6786 & ~w6787;
assign w6790 = ~w6788 & ~w6789;
assign w6791 = ~w6777 & w6790;
assign w6792 = w6777 & ~w6790;
assign w6793 = ~w6791 & ~w6792;
assign w6794 = ~w6776 & w6793;
assign w6795 = w6776 & ~w6793;
assign w6796 = ~w6794 & ~w6795;
assign w6797 = ~w6640 & ~w6718;
assign w6798 = w6796 & ~w6797;
assign w6799 = ~w6796 & w6797;
assign w6800 = ~w6798 & ~w6799;
assign w6801 = ~w6775 & w6800;
assign w6802 = w6775 & ~w6800;
assign w6803 = ~w6801 & ~w6802;
assign w6804 = ~w6754 & ~w6757;
assign w6805 = ~w6712 & ~w6715;
assign w6806 = (~w6697 & ~w6699) | (~w6697 & w17758) | (~w6699 & w17758);
assign w6807 = (~w6663 & ~w6665) | (~w6663 & w16905) | (~w6665 & w16905);
assign w6808 = pi28 & pi30;
assign w6809 = pi01 & pi57;
assign w6810 = ~w6808 & ~w6809;
assign w6811 = w6808 & w6809;
assign w6812 = ~w6810 & ~w6811;
assign w6813 = w6734 & w6812;
assign w6814 = ~w6734 & ~w6812;
assign w6815 = ~w6813 & ~w6814;
assign w6816 = ~w6688 & ~w6692;
assign w6817 = ~w6691 & ~w6816;
assign w6818 = w6815 & w6817;
assign w6819 = ~w6815 & ~w6817;
assign w6820 = ~w6818 & ~w6819;
assign w6821 = ~w6807 & w6820;
assign w6822 = w6807 & ~w6820;
assign w6823 = ~w6821 & ~w6822;
assign w6824 = ~w6806 & w6823;
assign w6825 = w6806 & ~w6823;
assign w6826 = ~w6824 & ~w6825;
assign w6827 = ~w6805 & w6826;
assign w6828 = w6805 & ~w6826;
assign w6829 = ~w6827 & ~w6828;
assign w6830 = (~w6622 & ~w6624) | (~w6622 & w17759) | (~w6624 & w17759);
assign w6831 = ~w6625 & ~w6629;
assign w6832 = ~w6628 & ~w6831;
assign w6833 = w6666 & ~w6669;
assign w6834 = ~w6671 & ~w6833;
assign w6835 = w6832 & ~w6834;
assign w6836 = ~w6832 & w6834;
assign w6837 = ~w6835 & ~w6836;
assign w6838 = w6603 & ~w6606;
assign w6839 = ~w6608 & ~w6838;
assign w6840 = ~w6837 & w6839;
assign w6841 = w6837 & ~w6839;
assign w6842 = ~w6840 & ~w6841;
assign w6843 = ~w6654 & ~w6658;
assign w6844 = ~w6657 & ~w6843;
assign w6845 = w6644 & ~w6647;
assign w6846 = ~w6649 & ~w6845;
assign w6847 = w6844 & ~w6846;
assign w6848 = ~w6844 & w6846;
assign w6849 = ~w6847 & ~w6848;
assign w6850 = w6679 & ~w6681;
assign w6851 = ~w6683 & ~w6850;
assign w6852 = ~w6849 & w6851;
assign w6853 = w6849 & ~w6851;
assign w6854 = ~w6852 & ~w6853;
assign w6855 = w6842 & w6854;
assign w6856 = ~w6842 & ~w6854;
assign w6857 = ~w6855 & ~w6856;
assign w6858 = ~w6830 & w6857;
assign w6859 = w6830 & ~w6857;
assign w6860 = ~w6858 & ~w6859;
assign w6861 = w6829 & w6860;
assign w6862 = ~w6829 & ~w6860;
assign w6863 = ~w6861 & ~w6862;
assign w6864 = ~w6804 & w6863;
assign w6865 = w6804 & ~w6863;
assign w6866 = ~w6864 & ~w6865;
assign w6867 = (~w6748 & ~w6750) | (~w6748 & w17132) | (~w6750 & w17132);
assign w6868 = (~w6730 & ~w6732) | (~w6730 & w17133) | (~w6732 & w17133);
assign w6869 = ~w6613 & ~w6617;
assign w6870 = ~w6616 & ~w6869;
assign w6871 = ~w6700 & ~w6704;
assign w6872 = ~w6703 & ~w6871;
assign w6873 = w6870 & w6872;
assign w6874 = ~w6870 & ~w6872;
assign w6875 = ~w6873 & ~w6874;
assign w6876 = w6868 & ~w6875;
assign w6877 = ~w6868 & w6875;
assign w6878 = ~w6876 & ~w6877;
assign w6879 = (~w6740 & ~w6742) | (~w6740 & w16906) | (~w6742 & w16906);
assign w6880 = ~w6878 & w6879;
assign w6881 = w6878 & ~w6879;
assign w6882 = ~w6880 & ~w6881;
assign w6883 = pi14 & pi44;
assign w6884 = pi13 & pi45;
assign w6885 = pi12 & pi46;
assign w6886 = ~w6884 & ~w6885;
assign w6887 = w6682 & w6688;
assign w6888 = ~w6886 & ~w6887;
assign w6889 = w6883 & ~w6888;
assign w6890 = ~w6883 & w6888;
assign w6891 = ~w6889 & ~w6890;
assign w6892 = pi15 & pi43;
assign w6893 = pi11 & pi47;
assign w6894 = ~w6892 & ~w6893;
assign w6895 = w6892 & w6893;
assign w6896 = ~w6894 & ~w6895;
assign w6897 = w6670 & ~w6896;
assign w6898 = ~w6670 & w6896;
assign w6899 = ~w6897 & ~w6898;
assign w6900 = ~w6891 & ~w6899;
assign w6901 = w6891 & w6899;
assign w6902 = ~w6900 & ~w6901;
assign w6903 = pi03 & pi55;
assign w6904 = pi19 & pi39;
assign w6905 = pi06 & pi52;
assign w6906 = ~w6904 & ~w6905;
assign w6907 = w6904 & w6905;
assign w6908 = ~w6906 & ~w6907;
assign w6909 = w6903 & ~w6908;
assign w6910 = ~w6903 & w6908;
assign w6911 = ~w6909 & ~w6910;
assign w6912 = w6902 & ~w6911;
assign w6913 = ~w6902 & w6911;
assign w6914 = ~w6912 & ~w6913;
assign w6915 = ~w6882 & ~w6914;
assign w6916 = w6882 & w6914;
assign w6917 = ~w6915 & ~w6916;
assign w6918 = ~w6867 & w6917;
assign w6919 = w6867 & ~w6917;
assign w6920 = ~w6918 & ~w6919;
assign w6921 = (~w6539 & ~w6541) | (~w6539 & w17134) | (~w6541 & w17134);
assign w6922 = pi05 & pi53;
assign w6923 = pi21 & pi37;
assign w6924 = ~w6648 & ~w6923;
assign w6925 = pi21 & pi38;
assign w6926 = w6645 & w6925;
assign w6927 = ~w6924 & ~w6926;
assign w6928 = w6922 & ~w6927;
assign w6929 = ~w6922 & w6927;
assign w6930 = ~w6928 & ~w6929;
assign w6931 = pi00 & pi58;
assign w6932 = pi04 & pi54;
assign w6933 = ~w6931 & ~w6932;
assign w6934 = w6931 & w6932;
assign w6935 = ~w6933 & ~w6934;
assign w6936 = w6347 & ~w6935;
assign w6937 = ~w6347 & w6935;
assign w6938 = ~w6936 & ~w6937;
assign w6939 = ~w6930 & ~w6938;
assign w6940 = w6930 & w6938;
assign w6941 = ~w6939 & ~w6940;
assign w6942 = pi17 & pi41;
assign w6943 = pi09 & pi49;
assign w6944 = pi16 & pi42;
assign w6945 = ~w6943 & ~w6944;
assign w6946 = w6943 & w6944;
assign w6947 = ~w6945 & ~w6946;
assign w6948 = w6942 & ~w6947;
assign w6949 = ~w6942 & w6947;
assign w6950 = ~w6948 & ~w6949;
assign w6951 = w6941 & ~w6950;
assign w6952 = ~w6941 & w6950;
assign w6953 = ~w6951 & ~w6952;
assign w6954 = pi18 & pi40;
assign w6955 = pi07 & pi51;
assign w6956 = pi08 & pi50;
assign w6957 = ~w6955 & ~w6956;
assign w6958 = pi08 & pi51;
assign w6959 = w6613 & w6958;
assign w6960 = ~w6957 & ~w6959;
assign w6961 = w6954 & ~w6960;
assign w6962 = ~w6954 & w6960;
assign w6963 = ~w6961 & ~w6962;
assign w6964 = pi22 & pi36;
assign w6965 = pi24 & pi34;
assign w6966 = ~w6607 & ~w6965;
assign w6967 = pi24 & pi35;
assign w6968 = w6604 & w6967;
assign w6969 = ~w6966 & ~w6968;
assign w6970 = w6964 & ~w6969;
assign w6971 = ~w6964 & w6969;
assign w6972 = ~w6970 & ~w6971;
assign w6973 = ~w6963 & ~w6972;
assign w6974 = w6963 & w6972;
assign w6975 = ~w6973 & ~w6974;
assign w6976 = pi25 & pi33;
assign w6977 = pi26 & pi32;
assign w6978 = pi27 & pi31;
assign w6979 = ~w6977 & ~w6978;
assign w6980 = w6977 & w6978;
assign w6981 = ~w6979 & ~w6980;
assign w6982 = w6976 & ~w6981;
assign w6983 = ~w6976 & w6981;
assign w6984 = ~w6982 & ~w6983;
assign w6985 = w6975 & ~w6984;
assign w6986 = ~w6975 & w6984;
assign w6987 = ~w6985 & ~w6986;
assign w6988 = w6953 & w6987;
assign w6989 = ~w6953 & ~w6987;
assign w6990 = ~w6988 & ~w6989;
assign w6991 = ~w6921 & w6990;
assign w6992 = w6921 & ~w6990;
assign w6993 = ~w6991 & ~w6992;
assign w6994 = ~w6920 & ~w6993;
assign w6995 = w6920 & w6993;
assign w6996 = ~w6994 & ~w6995;
assign w6997 = ~w6866 & ~w6996;
assign w6998 = w6866 & w6996;
assign w6999 = ~w6997 & ~w6998;
assign w7000 = ~w6803 & ~w6999;
assign w7001 = w6803 & w6999;
assign w7002 = ~w7000 & ~w7001;
assign w7003 = ~w6774 & w7002;
assign w7004 = w6774 & ~w7002;
assign w7005 = ~w7003 & ~w7004;
assign w7006 = (w6298 & w16541) | (w6298 & w16542) | (w16541 & w16542);
assign w7007 = ~w6767 & ~w7006;
assign w7008 = w7005 & w7007;
assign w7009 = ~w7005 & ~w7007;
assign w7010 = ~w7008 & ~w7009;
assign w7011 = ~w6864 & ~w6998;
assign w7012 = (~w6918 & ~w6920) | (~w6918 & w17760) | (~w6920 & w17760);
assign w7013 = (~w6827 & ~w6829) | (~w6827 & w17761) | (~w6829 & w17761);
assign w7014 = (~w6881 & ~w6882) | (~w6881 & w17135) | (~w6882 & w17135);
assign w7015 = (~w6835 & ~w6837) | (~w6835 & w17762) | (~w6837 & w17762);
assign w7016 = (~w6873 & ~w6875) | (~w6873 & w17136) | (~w6875 & w17136);
assign w7017 = (~w6847 & ~w6849) | (~w6847 & w17137) | (~w6849 & w17137);
assign w7018 = ~w7016 & ~w7017;
assign w7019 = w7016 & w7017;
assign w7020 = ~w7018 & ~w7019;
assign w7021 = w7015 & ~w7020;
assign w7022 = ~w7015 & w7020;
assign w7023 = ~w7021 & ~w7022;
assign w7024 = (~w6855 & ~w6857) | (~w6855 & w17138) | (~w6857 & w17138);
assign w7025 = ~w7023 & w7024;
assign w7026 = w7023 & ~w7024;
assign w7027 = ~w7025 & ~w7026;
assign w7028 = ~w7014 & w7027;
assign w7029 = w7014 & ~w7027;
assign w7030 = ~w7028 & ~w7029;
assign w7031 = ~w7013 & w7030;
assign w7032 = w7013 & ~w7030;
assign w7033 = ~w7031 & ~w7032;
assign w7034 = ~w7012 & w7033;
assign w7035 = w7012 & ~w7033;
assign w7036 = ~w7034 & ~w7035;
assign w7037 = ~w7011 & w7036;
assign w7038 = w7011 & ~w7036;
assign w7039 = ~w7037 & ~w7038;
assign w7040 = ~w6794 & ~w6798;
assign w7041 = (~w6939 & ~w6941) | (~w6939 & w17763) | (~w6941 & w17763);
assign w7042 = (~w6900 & ~w6902) | (~w6900 & w16907) | (~w6902 & w16907);
assign w7043 = (~w6973 & ~w6975) | (~w6973 & w16908) | (~w6975 & w16908);
assign w7044 = ~w7042 & ~w7043;
assign w7045 = w7042 & w7043;
assign w7046 = ~w7044 & ~w7045;
assign w7047 = w7041 & ~w7046;
assign w7048 = ~w7041 & w7046;
assign w7049 = ~w7047 & ~w7048;
assign w7050 = ~w6988 & ~w6991;
assign w7051 = ~w6347 & ~w6934;
assign w7052 = ~w6933 & ~w7051;
assign w7053 = ~w6903 & ~w6907;
assign w7054 = ~w6906 & ~w7053;
assign w7055 = w7052 & w7054;
assign w7056 = ~w7052 & ~w7054;
assign w7057 = ~w7055 & ~w7056;
assign w7058 = ~w6942 & ~w6946;
assign w7059 = ~w6945 & ~w7058;
assign w7060 = ~w7057 & ~w7059;
assign w7061 = w7057 & w7059;
assign w7062 = ~w7060 & ~w7061;
assign w7063 = w6922 & ~w6924;
assign w7064 = ~w6926 & ~w7063;
assign w7065 = w6964 & ~w6966;
assign w7066 = ~w6968 & ~w7065;
assign w7067 = ~w7064 & ~w7066;
assign w7068 = w7064 & w7066;
assign w7069 = ~w7067 & ~w7068;
assign w7070 = w6954 & ~w6957;
assign w7071 = ~w6959 & ~w7070;
assign w7072 = ~w7069 & w7071;
assign w7073 = w7069 & ~w7071;
assign w7074 = ~w7072 & ~w7073;
assign w7075 = pi58 & w1939;
assign w7076 = pi01 & pi58;
assign w7077 = ~pi30 & ~w7076;
assign w7078 = ~w7075 & ~w7077;
assign w7079 = w6883 & ~w6886;
assign w7080 = ~w6887 & ~w7079;
assign w7081 = w7078 & ~w7080;
assign w7082 = ~w7078 & w7080;
assign w7083 = ~w7081 & ~w7082;
assign w7084 = ~w6670 & ~w6895;
assign w7085 = ~w6894 & ~w7084;
assign w7086 = w7083 & w7085;
assign w7087 = ~w7083 & ~w7085;
assign w7088 = ~w7086 & ~w7087;
assign w7089 = w7074 & w7088;
assign w7090 = ~w7074 & ~w7088;
assign w7091 = ~w7089 & ~w7090;
assign w7092 = w7062 & w7091;
assign w7093 = ~w7062 & ~w7091;
assign w7094 = ~w7092 & ~w7093;
assign w7095 = ~w7050 & w7094;
assign w7096 = w7050 & ~w7094;
assign w7097 = ~w7095 & ~w7096;
assign w7098 = w7049 & w7097;
assign w7099 = ~w7049 & ~w7097;
assign w7100 = ~w7098 & ~w7099;
assign w7101 = ~w7040 & w7100;
assign w7102 = w7040 & ~w7100;
assign w7103 = ~w7101 & ~w7102;
assign w7104 = (~w6789 & ~w6790) | (~w6789 & w17764) | (~w6790 & w17764);
assign w7105 = (~w6821 & ~w6823) | (~w6821 & w17139) | (~w6823 & w17139);
assign w7106 = pi29 & pi30;
assign w7107 = pi28 & pi31;
assign w7108 = ~w7106 & ~w7107;
assign w7109 = w7106 & w7107;
assign w7110 = ~w7108 & ~w7109;
assign w7111 = w6682 & ~w7110;
assign w7112 = ~w6682 & w7110;
assign w7113 = ~w7111 & ~w7112;
assign w7114 = pi11 & pi48;
assign w7115 = pi14 & pi45;
assign w7116 = pi12 & pi47;
assign w7117 = ~w7115 & ~w7116;
assign w7118 = w7115 & w7116;
assign w7119 = ~w7117 & ~w7118;
assign w7120 = w7114 & ~w7119;
assign w7121 = ~w7114 & w7119;
assign w7122 = ~w7120 & ~w7121;
assign w7123 = ~w7113 & ~w7122;
assign w7124 = w7113 & w7122;
assign w7125 = ~w7123 & ~w7124;
assign w7126 = pi16 & pi43;
assign w7127 = pi17 & pi42;
assign w7128 = ~w7126 & ~w7127;
assign w7129 = pi17 & pi43;
assign w7130 = w6944 & w7129;
assign w7131 = ~w7128 & ~w7130;
assign w7132 = w6958 & ~w7131;
assign w7133 = ~w6958 & w7131;
assign w7134 = ~w7132 & ~w7133;
assign w7135 = w7125 & ~w7134;
assign w7136 = ~w7125 & w7134;
assign w7137 = ~w7135 & ~w7136;
assign w7138 = ~w6976 & ~w6980;
assign w7139 = ~w6979 & ~w7138;
assign w7140 = pi02 & pi57;
assign w7141 = pi03 & pi56;
assign w7142 = ~w7140 & ~w7141;
assign w7143 = pi03 & pi57;
assign w7144 = w6347 & w7143;
assign w7145 = ~w7142 & ~w7144;
assign w7146 = w6811 & ~w7145;
assign w7147 = ~w6811 & w7145;
assign w7148 = ~w7146 & ~w7147;
assign w7149 = w7139 & ~w7148;
assign w7150 = ~w7139 & w7148;
assign w7151 = ~w7149 & ~w7150;
assign w7152 = pi04 & pi55;
assign w7153 = pi05 & pi54;
assign w7154 = pi19 & pi40;
assign w7155 = ~w7153 & ~w7154;
assign w7156 = w7153 & w7154;
assign w7157 = ~w7155 & ~w7156;
assign w7158 = w7152 & ~w7157;
assign w7159 = ~w7152 & w7157;
assign w7160 = ~w7158 & ~w7159;
assign w7161 = w7151 & ~w7160;
assign w7162 = ~w7151 & w7160;
assign w7163 = ~w7161 & ~w7162;
assign w7164 = w7137 & w7163;
assign w7165 = ~w7137 & ~w7163;
assign w7166 = ~w7164 & ~w7165;
assign w7167 = ~w7105 & w7166;
assign w7168 = w7105 & ~w7166;
assign w7169 = ~w7167 & ~w7168;
assign w7170 = ~w7104 & w7169;
assign w7171 = w7104 & ~w7169;
assign w7172 = ~w7170 & ~w7171;
assign w7173 = ~w6813 & ~w6818;
assign w7174 = pi06 & pi53;
assign w7175 = pi07 & pi52;
assign w7176 = pi18 & pi41;
assign w7177 = ~w7175 & ~w7176;
assign w7178 = w7175 & w7176;
assign w7179 = ~w7177 & ~w7178;
assign w7180 = w7174 & ~w7179;
assign w7181 = ~w7174 & w7179;
assign w7182 = ~w7180 & ~w7181;
assign w7183 = pi09 & pi50;
assign w7184 = pi15 & pi44;
assign w7185 = pi10 & pi49;
assign w7186 = ~w7184 & ~w7185;
assign w7187 = w7184 & w7185;
assign w7188 = ~w7186 & ~w7187;
assign w7189 = w7183 & ~w7188;
assign w7190 = ~w7183 & w7188;
assign w7191 = ~w7189 & ~w7190;
assign w7192 = ~w7182 & ~w7191;
assign w7193 = w7182 & w7191;
assign w7194 = ~w7192 & ~w7193;
assign w7195 = w7173 & ~w7194;
assign w7196 = ~w7173 & w7194;
assign w7197 = ~w7195 & ~w7196;
assign w7198 = (~w6781 & ~w6783) | (~w6781 & w16909) | (~w6783 & w16909);
assign w7199 = ~w7197 & w7198;
assign w7200 = w7197 & ~w7198;
assign w7201 = ~w7199 & ~w7200;
assign w7202 = pi20 & pi39;
assign w7203 = pi22 & pi37;
assign w7204 = ~w6925 & ~w7203;
assign w7205 = pi22 & pi38;
assign w7206 = w6923 & w7205;
assign w7207 = ~w7204 & ~w7206;
assign w7208 = w7202 & ~w7207;
assign w7209 = ~w7202 & w7207;
assign w7210 = ~w7208 & ~w7209;
assign w7211 = pi23 & pi36;
assign w7212 = pi25 & pi34;
assign w7213 = ~w6967 & ~w7212;
assign w7214 = pi25 & pi35;
assign w7215 = w6965 & w7214;
assign w7216 = ~w7213 & ~w7215;
assign w7217 = w7211 & ~w7216;
assign w7218 = ~w7211 & w7216;
assign w7219 = ~w7217 & ~w7218;
assign w7220 = ~w7210 & ~w7219;
assign w7221 = w7210 & w7219;
assign w7222 = ~w7220 & ~w7221;
assign w7223 = pi26 & pi33;
assign w7224 = pi27 & pi32;
assign w7225 = pi00 & pi59;
assign w7226 = ~w7224 & ~w7225;
assign w7227 = w7224 & w7225;
assign w7228 = ~w7226 & ~w7227;
assign w7229 = w7223 & ~w7228;
assign w7230 = ~w7223 & w7228;
assign w7231 = ~w7229 & ~w7230;
assign w7232 = w7222 & ~w7231;
assign w7233 = ~w7222 & w7231;
assign w7234 = ~w7232 & ~w7233;
assign w7235 = w7201 & w7234;
assign w7236 = ~w7201 & ~w7234;
assign w7237 = ~w7235 & ~w7236;
assign w7238 = w7172 & w7237;
assign w7239 = ~w7172 & ~w7237;
assign w7240 = ~w7238 & ~w7239;
assign w7241 = w7103 & w7240;
assign w7242 = ~w7103 & ~w7240;
assign w7243 = ~w7241 & ~w7242;
assign w7244 = w7039 & w7243;
assign w7245 = ~w7039 & ~w7243;
assign w7246 = ~w7244 & ~w7245;
assign w7247 = ~w6801 & ~w7001;
assign w7248 = ~w7246 & w7247;
assign w7249 = w7246 & ~w7247;
assign w7250 = ~w7248 & ~w7249;
assign w7251 = ~w6767 & ~w7004;
assign w7252 = ~w7006 & w7251;
assign w7253 = ~w7003 & ~w7252;
assign w7254 = w7250 & w7253;
assign w7255 = ~w7250 & ~w7253;
assign w7256 = ~w7254 & ~w7255;
assign w7257 = ~w7037 & ~w7244;
assign w7258 = ~w7101 & ~w7241;
assign w7259 = ~w7170 & ~w7238;
assign w7260 = (~w7095 & ~w7097) | (~w7095 & w17765) | (~w7097 & w17765);
assign w7261 = (~w7149 & ~w7151) | (~w7149 & w16910) | (~w7151 & w16910);
assign w7262 = (~w7067 & ~w7069) | (~w7067 & w16752) | (~w7069 & w16752);
assign w7263 = (~w7055 & ~w7057) | (~w7055 & w16753) | (~w7057 & w16753);
assign w7264 = ~w7262 & ~w7263;
assign w7265 = w7262 & w7263;
assign w7266 = ~w7264 & ~w7265;
assign w7267 = w7261 & ~w7266;
assign w7268 = ~w7261 & w7266;
assign w7269 = ~w7267 & ~w7268;
assign w7270 = (~w7044 & ~w7046) | (~w7044 & w17140) | (~w7046 & w17140);
assign w7271 = ~w7269 & w7270;
assign w7272 = w7269 & ~w7270;
assign w7273 = ~w7271 & ~w7272;
assign w7274 = (~w7200 & ~w7201) | (~w7200 & w17141) | (~w7201 & w17141);
assign w7275 = w7273 & ~w7274;
assign w7276 = ~w7273 & w7274;
assign w7277 = ~w7275 & ~w7276;
assign w7278 = ~w7260 & w7277;
assign w7279 = w7260 & ~w7277;
assign w7280 = ~w7278 & ~w7279;
assign w7281 = ~w7259 & w7280;
assign w7282 = w7259 & ~w7280;
assign w7283 = ~w7281 & ~w7282;
assign w7284 = ~w7258 & w7283;
assign w7285 = w7258 & ~w7283;
assign w7286 = ~w7284 & ~w7285;
assign w7287 = ~w7089 & ~w7092;
assign w7288 = ~w7081 & ~w7086;
assign w7289 = pi00 & pi60;
assign w7290 = w7075 & w7289;
assign w7291 = ~w7075 & ~w7289;
assign w7292 = ~w7290 & ~w7291;
assign w7293 = pi01 & pi59;
assign w7294 = pi29 & pi31;
assign w7295 = ~w7293 & ~w7294;
assign w7296 = w7293 & w7294;
assign w7297 = ~w7295 & ~w7296;
assign w7298 = w7292 & w7297;
assign w7299 = ~w7292 & ~w7297;
assign w7300 = ~w7298 & ~w7299;
assign w7301 = pi27 & pi33;
assign w7302 = pi28 & pi32;
assign w7303 = pi23 & pi37;
assign w7304 = ~w7302 & ~w7303;
assign w7305 = w7302 & w7303;
assign w7306 = ~w7304 & ~w7305;
assign w7307 = w7301 & ~w7306;
assign w7308 = ~w7301 & w7306;
assign w7309 = ~w7307 & ~w7308;
assign w7310 = w7300 & ~w7309;
assign w7311 = ~w7300 & w7309;
assign w7312 = ~w7310 & ~w7311;
assign w7313 = w7288 & ~w7312;
assign w7314 = ~w7288 & w7312;
assign w7315 = ~w7313 & ~w7314;
assign w7316 = pi14 & pi46;
assign w7317 = pi12 & pi48;
assign w7318 = pi13 & pi47;
assign w7319 = ~w7317 & ~w7318;
assign w7320 = pi13 & pi48;
assign w7321 = w7116 & w7320;
assign w7322 = ~w7319 & ~w7321;
assign w7323 = w7316 & ~w7322;
assign w7324 = ~w7316 & w7322;
assign w7325 = ~w7323 & ~w7324;
assign w7326 = pi07 & pi53;
assign w7327 = pi08 & pi52;
assign w7328 = pi18 & pi42;
assign w7329 = ~w7327 & ~w7328;
assign w7330 = w7327 & w7328;
assign w7331 = ~w7329 & ~w7330;
assign w7332 = w7326 & ~w7331;
assign w7333 = ~w7326 & w7331;
assign w7334 = ~w7332 & ~w7333;
assign w7335 = ~w7325 & ~w7334;
assign w7336 = w7325 & w7334;
assign w7337 = ~w7335 & ~w7336;
assign w7338 = pi05 & pi55;
assign w7339 = pi06 & pi54;
assign w7340 = pi19 & pi41;
assign w7341 = ~w7339 & ~w7340;
assign w7342 = w7339 & w7340;
assign w7343 = ~w7341 & ~w7342;
assign w7344 = w7338 & ~w7343;
assign w7345 = ~w7338 & w7343;
assign w7346 = ~w7344 & ~w7345;
assign w7347 = w7337 & ~w7346;
assign w7348 = ~w7337 & w7346;
assign w7349 = ~w7347 & ~w7348;
assign w7350 = ~w7315 & ~w7349;
assign w7351 = w7315 & w7349;
assign w7352 = ~w7350 & ~w7351;
assign w7353 = ~w7287 & w7352;
assign w7354 = w7287 & ~w7352;
assign w7355 = ~w7353 & ~w7354;
assign w7356 = ~w7026 & ~w7028;
assign w7357 = (~w7018 & ~w7020) | (~w7018 & w17572) | (~w7020 & w17572);
assign w7358 = pi02 & pi58;
assign w7359 = pi04 & pi56;
assign w7360 = ~w7143 & ~w7359;
assign w7361 = pi04 & pi57;
assign w7362 = w7141 & w7361;
assign w7363 = ~w7360 & ~w7362;
assign w7364 = w7358 & ~w7363;
assign w7365 = ~w7358 & w7363;
assign w7366 = ~w7364 & ~w7365;
assign w7367 = pi20 & pi40;
assign w7368 = pi21 & pi39;
assign w7369 = ~w7205 & ~w7368;
assign w7370 = pi22 & pi39;
assign w7371 = w6925 & w7370;
assign w7372 = ~w7369 & ~w7371;
assign w7373 = w7367 & ~w7372;
assign w7374 = ~w7367 & w7372;
assign w7375 = ~w7373 & ~w7374;
assign w7376 = ~w7366 & ~w7375;
assign w7377 = w7366 & w7375;
assign w7378 = ~w7376 & ~w7377;
assign w7379 = pi24 & pi36;
assign w7380 = pi26 & pi34;
assign w7381 = ~w7214 & ~w7380;
assign w7382 = pi26 & pi35;
assign w7383 = w7212 & w7382;
assign w7384 = ~w7381 & ~w7383;
assign w7385 = w7379 & ~w7384;
assign w7386 = ~w7379 & w7384;
assign w7387 = ~w7385 & ~w7386;
assign w7388 = w7378 & ~w7387;
assign w7389 = ~w7378 & w7387;
assign w7390 = ~w7388 & ~w7389;
assign w7391 = ~w7357 & w7390;
assign w7392 = w7357 & ~w7390;
assign w7393 = ~w7391 & ~w7392;
assign w7394 = ~w7114 & ~w7118;
assign w7395 = ~w7117 & ~w7394;
assign w7396 = pi09 & pi51;
assign w7397 = pi16 & pi44;
assign w7398 = ~w7396 & ~w7397;
assign w7399 = w7396 & w7397;
assign w7400 = ~w7398 & ~w7399;
assign w7401 = w7129 & ~w7400;
assign w7402 = ~w7129 & w7400;
assign w7403 = ~w7401 & ~w7402;
assign w7404 = w7395 & ~w7403;
assign w7405 = ~w7395 & w7403;
assign w7406 = ~w7404 & ~w7405;
assign w7407 = pi10 & pi50;
assign w7408 = pi15 & pi45;
assign w7409 = pi11 & pi49;
assign w7410 = ~w7408 & ~w7409;
assign w7411 = w7408 & w7409;
assign w7412 = ~w7410 & ~w7411;
assign w7413 = w7407 & ~w7412;
assign w7414 = ~w7407 & w7412;
assign w7415 = ~w7413 & ~w7414;
assign w7416 = w7406 & ~w7415;
assign w7417 = ~w7406 & w7415;
assign w7418 = ~w7416 & ~w7417;
assign w7419 = ~w7393 & ~w7418;
assign w7420 = w7393 & w7418;
assign w7421 = ~w7419 & ~w7420;
assign w7422 = ~w7356 & w7421;
assign w7423 = w7356 & ~w7421;
assign w7424 = ~w7422 & ~w7423;
assign w7425 = ~w7355 & ~w7424;
assign w7426 = w7355 & w7424;
assign w7427 = ~w7425 & ~w7426;
assign w7428 = ~w7031 & ~w7034;
assign w7429 = ~w7174 & ~w7178;
assign w7430 = ~w7177 & ~w7429;
assign w7431 = w6958 & ~w7128;
assign w7432 = ~w7130 & ~w7431;
assign w7433 = w7430 & ~w7432;
assign w7434 = ~w7430 & w7432;
assign w7435 = ~w7433 & ~w7434;
assign w7436 = ~w6682 & ~w7109;
assign w7437 = ~w7108 & ~w7436;
assign w7438 = ~w7435 & ~w7437;
assign w7439 = w7435 & w7437;
assign w7440 = ~w7438 & ~w7439;
assign w7441 = ~w7220 & ~w7232;
assign w7442 = ~w7440 & w7441;
assign w7443 = w7440 & ~w7441;
assign w7444 = ~w7442 & ~w7443;
assign w7445 = ~w7123 & ~w7135;
assign w7446 = ~w7444 & w7445;
assign w7447 = w7444 & ~w7445;
assign w7448 = ~w7446 & ~w7447;
assign w7449 = ~w7164 & ~w7167;
assign w7450 = ~w7192 & ~w7196;
assign w7451 = ~w7152 & ~w7156;
assign w7452 = ~w7155 & ~w7451;
assign w7453 = w7202 & ~w7204;
assign w7454 = ~w7206 & ~w7453;
assign w7455 = w7452 & ~w7454;
assign w7456 = ~w7452 & w7454;
assign w7457 = ~w7455 & ~w7456;
assign w7458 = w7211 & ~w7213;
assign w7459 = ~w7215 & ~w7458;
assign w7460 = ~w7457 & w7459;
assign w7461 = w7457 & ~w7459;
assign w7462 = ~w7460 & ~w7461;
assign w7463 = ~w7223 & ~w7227;
assign w7464 = ~w7226 & ~w7463;
assign w7465 = w6811 & ~w7142;
assign w7466 = ~w7144 & ~w7465;
assign w7467 = w7464 & ~w7466;
assign w7468 = ~w7464 & w7466;
assign w7469 = ~w7467 & ~w7468;
assign w7470 = ~w7183 & ~w7187;
assign w7471 = ~w7186 & ~w7470;
assign w7472 = ~w7469 & ~w7471;
assign w7473 = w7469 & w7471;
assign w7474 = ~w7472 & ~w7473;
assign w7475 = w7462 & w7474;
assign w7476 = ~w7462 & ~w7474;
assign w7477 = ~w7475 & ~w7476;
assign w7478 = ~w7450 & w7477;
assign w7479 = w7450 & ~w7477;
assign w7480 = ~w7478 & ~w7479;
assign w7481 = ~w7449 & w7480;
assign w7482 = w7449 & ~w7480;
assign w7483 = ~w7481 & ~w7482;
assign w7484 = w7448 & w7483;
assign w7485 = ~w7448 & ~w7483;
assign w7486 = ~w7484 & ~w7485;
assign w7487 = ~w7428 & w7486;
assign w7488 = w7428 & ~w7486;
assign w7489 = ~w7487 & ~w7488;
assign w7490 = w7427 & w7489;
assign w7491 = ~w7427 & ~w7489;
assign w7492 = ~w7490 & ~w7491;
assign w7493 = w7286 & w7492;
assign w7494 = ~w7286 & ~w7492;
assign w7495 = ~w7493 & ~w7494;
assign w7496 = w7257 & ~w7495;
assign w7497 = ~w7257 & w7495;
assign w7498 = ~w7496 & ~w7497;
assign w7499 = ~w7003 & ~w7249;
assign w7500 = (~w7006 & w16544) | (~w7006 & w16545) | (w16544 & w16545);
assign w7501 = w7498 & w7500;
assign w7502 = ~w7498 & ~w7500;
assign w7503 = ~w7501 & ~w7502;
assign w7504 = ~w7284 & ~w7493;
assign w7505 = (~w7481 & ~w7483) | (~w7481 & w17766) | (~w7483 & w17766);
assign w7506 = ~w7272 & ~w7275;
assign w7507 = (~w7264 & ~w7266) | (~w7264 & w16911) | (~w7266 & w16911);
assign w7508 = pi11 & pi50;
assign w7509 = pi14 & pi47;
assign w7510 = pi12 & pi49;
assign w7511 = ~w7509 & ~w7510;
assign w7512 = w7509 & w7510;
assign w7513 = ~w7511 & ~w7512;
assign w7514 = w7508 & ~w7513;
assign w7515 = ~w7508 & w7513;
assign w7516 = ~w7514 & ~w7515;
assign w7517 = pi16 & pi45;
assign w7518 = pi15 & pi46;
assign w7519 = pi10 & pi51;
assign w7520 = ~w7518 & ~w7519;
assign w7521 = w7518 & w7519;
assign w7522 = ~w7520 & ~w7521;
assign w7523 = w7517 & ~w7522;
assign w7524 = ~w7517 & w7522;
assign w7525 = ~w7523 & ~w7524;
assign w7526 = ~w7516 & ~w7525;
assign w7527 = w7516 & w7525;
assign w7528 = ~w7526 & ~w7527;
assign w7529 = pi30 & pi31;
assign w7530 = pi29 & pi32;
assign w7531 = ~w7529 & ~w7530;
assign w7532 = w7529 & w7530;
assign w7533 = ~w7531 & ~w7532;
assign w7534 = w7320 & ~w7533;
assign w7535 = ~w7320 & w7533;
assign w7536 = ~w7534 & ~w7535;
assign w7537 = w7528 & ~w7536;
assign w7538 = ~w7528 & w7536;
assign w7539 = ~w7537 & ~w7538;
assign w7540 = ~w7507 & w7539;
assign w7541 = w7507 & ~w7539;
assign w7542 = ~w7540 & ~w7541;
assign w7543 = pi06 & pi55;
assign w7544 = pi20 & pi41;
assign w7545 = pi21 & pi40;
assign w7546 = ~w7544 & ~w7545;
assign w7547 = pi21 & pi41;
assign w7548 = w7367 & w7547;
assign w7549 = ~w7546 & ~w7548;
assign w7550 = w7543 & ~w7549;
assign w7551 = ~w7543 & w7549;
assign w7552 = ~w7550 & ~w7551;
assign w7553 = pi00 & pi61;
assign w7554 = pi02 & pi59;
assign w7555 = pi05 & pi56;
assign w7556 = ~w7554 & ~w7555;
assign w7557 = w7554 & w7555;
assign w7558 = ~w7556 & ~w7557;
assign w7559 = w7553 & ~w7558;
assign w7560 = ~w7553 & w7558;
assign w7561 = ~w7559 & ~w7560;
assign w7562 = ~w7552 & ~w7561;
assign w7563 = w7552 & w7561;
assign w7564 = ~w7562 & ~w7563;
assign w7565 = pi24 & pi37;
assign w7566 = pi25 & pi36;
assign w7567 = ~w7565 & ~w7566;
assign w7568 = w7565 & w7566;
assign w7569 = ~w7567 & ~w7568;
assign w7570 = w7370 & ~w7569;
assign w7571 = ~w7370 & w7569;
assign w7572 = ~w7570 & ~w7571;
assign w7573 = w7564 & ~w7572;
assign w7574 = ~w7564 & w7572;
assign w7575 = ~w7573 & ~w7574;
assign w7576 = ~w7542 & ~w7575;
assign w7577 = w7542 & w7575;
assign w7578 = ~w7576 & ~w7577;
assign w7579 = ~w7506 & w7578;
assign w7580 = w7506 & ~w7578;
assign w7581 = ~w7579 & ~w7580;
assign w7582 = ~w7505 & w7581;
assign w7583 = w7505 & ~w7581;
assign w7584 = ~w7582 & ~w7583;
assign w7585 = ~w7278 & ~w7281;
assign w7586 = ~w7351 & ~w7353;
assign w7587 = (~w7290 & ~w7292) | (~w7290 & w17142) | (~w7292 & w17142);
assign w7588 = ~w7326 & ~w7330;
assign w7589 = ~w7329 & ~w7588;
assign w7590 = ~w7129 & ~w7399;
assign w7591 = ~w7398 & ~w7590;
assign w7592 = w7589 & w7591;
assign w7593 = ~w7589 & ~w7591;
assign w7594 = ~w7592 & ~w7593;
assign w7595 = w7587 & ~w7594;
assign w7596 = ~w7587 & w7594;
assign w7597 = ~w7595 & ~w7596;
assign w7598 = ~w7335 & ~w7347;
assign w7599 = ~w7597 & w7598;
assign w7600 = w7597 & ~w7598;
assign w7601 = ~w7599 & ~w7600;
assign w7602 = ~w7310 & ~w7314;
assign w7603 = ~w7601 & w7602;
assign w7604 = w7601 & ~w7602;
assign w7605 = ~w7603 & ~w7604;
assign w7606 = ~w7376 & ~w7388;
assign w7607 = ~w7301 & ~w7305;
assign w7608 = ~w7304 & ~w7607;
assign w7609 = w7379 & ~w7381;
assign w7610 = ~w7383 & ~w7609;
assign w7611 = w7608 & ~w7610;
assign w7612 = ~w7608 & w7610;
assign w7613 = ~w7611 & ~w7612;
assign w7614 = w7367 & ~w7369;
assign w7615 = ~w7371 & ~w7614;
assign w7616 = ~w7613 & w7615;
assign w7617 = w7613 & ~w7615;
assign w7618 = ~w7616 & ~w7617;
assign w7619 = ~w7338 & ~w7342;
assign w7620 = ~w7341 & ~w7619;
assign w7621 = w7358 & ~w7360;
assign w7622 = ~w7362 & ~w7621;
assign w7623 = w7620 & ~w7622;
assign w7624 = ~w7620 & w7622;
assign w7625 = ~w7623 & ~w7624;
assign w7626 = ~w7407 & ~w7411;
assign w7627 = ~w7410 & ~w7626;
assign w7628 = ~w7625 & ~w7627;
assign w7629 = w7625 & w7627;
assign w7630 = ~w7628 & ~w7629;
assign w7631 = w7618 & w7630;
assign w7632 = ~w7618 & ~w7630;
assign w7633 = ~w7631 & ~w7632;
assign w7634 = ~w7606 & w7633;
assign w7635 = w7606 & ~w7633;
assign w7636 = ~w7634 & ~w7635;
assign w7637 = ~w7605 & ~w7636;
assign w7638 = w7605 & w7636;
assign w7639 = ~w7637 & ~w7638;
assign w7640 = w7586 & w7639;
assign w7641 = ~w7586 & ~w7639;
assign w7642 = ~w7640 & ~w7641;
assign w7643 = ~w7585 & ~w7642;
assign w7644 = w7585 & w7642;
assign w7645 = ~w7643 & ~w7644;
assign w7646 = w7584 & w7645;
assign w7647 = ~w7584 & ~w7645;
assign w7648 = ~w7646 & ~w7647;
assign w7649 = ~w7487 & ~w7490;
assign w7650 = (~w7422 & ~w7424) | (~w7422 & w17767) | (~w7424 & w17767);
assign w7651 = (~w7391 & ~w7393) | (~w7391 & w17768) | (~w7393 & w17768);
assign w7652 = ~w7404 & ~w7416;
assign w7653 = (~w7455 & ~w7457) | (~w7455 & w17769) | (~w7457 & w17769);
assign w7654 = pi01 & pi60;
assign w7655 = ~w7296 & w17573;
assign w7656 = (w7654 & w7296) | (w7654 & w17574) | (w7296 & w17574);
assign w7657 = ~w7655 & ~w7656;
assign w7658 = w7316 & ~w7319;
assign w7659 = ~w7321 & ~w7658;
assign w7660 = ~w7657 & ~w7659;
assign w7661 = w7657 & w7659;
assign w7662 = ~w7660 & ~w7661;
assign w7663 = ~w7653 & w7662;
assign w7664 = w7653 & ~w7662;
assign w7665 = ~w7663 & ~w7664;
assign w7666 = ~w7652 & w7665;
assign w7667 = w7652 & ~w7665;
assign w7668 = ~w7666 & ~w7667;
assign w7669 = (~w7467 & ~w7469) | (~w7467 & w17770) | (~w7469 & w17770);
assign w7670 = (~w7433 & ~w7435) | (~w7433 & w17143) | (~w7435 & w17143);
assign w7671 = pi23 & pi38;
assign w7672 = pi03 & pi58;
assign w7673 = ~w7361 & ~w7672;
assign w7674 = pi04 & pi58;
assign w7675 = w7143 & w7674;
assign w7676 = ~w7673 & ~w7675;
assign w7677 = w7671 & ~w7676;
assign w7678 = ~w7671 & w7676;
assign w7679 = ~w7677 & ~w7678;
assign w7680 = ~w7670 & ~w7679;
assign w7681 = w7670 & w7679;
assign w7682 = ~w7680 & ~w7681;
assign w7683 = ~w7669 & w7682;
assign w7684 = w7669 & ~w7682;
assign w7685 = ~w7683 & ~w7684;
assign w7686 = w7668 & w7685;
assign w7687 = ~w7668 & ~w7685;
assign w7688 = ~w7686 & ~w7687;
assign w7689 = ~w7651 & w7688;
assign w7690 = w7651 & ~w7688;
assign w7691 = ~w7689 & ~w7690;
assign w7692 = ~w7443 & ~w7447;
assign w7693 = (~w7475 & ~w7477) | (~w7475 & w17771) | (~w7477 & w17771);
assign w7694 = pi19 & pi42;
assign w7695 = pi07 & pi54;
assign w7696 = pi08 & pi53;
assign w7697 = ~w7695 & ~w7696;
assign w7698 = pi08 & pi54;
assign w7699 = w7326 & w7698;
assign w7700 = ~w7697 & ~w7699;
assign w7701 = w7694 & ~w7700;
assign w7702 = ~w7694 & w7700;
assign w7703 = ~w7701 & ~w7702;
assign w7704 = pi18 & pi43;
assign w7705 = pi09 & pi52;
assign w7706 = pi17 & pi44;
assign w7707 = ~w7705 & ~w7706;
assign w7708 = w7705 & w7706;
assign w7709 = ~w7707 & ~w7708;
assign w7710 = w7704 & ~w7709;
assign w7711 = ~w7704 & w7709;
assign w7712 = ~w7710 & ~w7711;
assign w7713 = ~w7703 & ~w7712;
assign w7714 = w7703 & w7712;
assign w7715 = ~w7713 & ~w7714;
assign w7716 = pi27 & pi34;
assign w7717 = pi28 & pi33;
assign w7718 = ~w7716 & ~w7717;
assign w7719 = w7716 & w7717;
assign w7720 = ~w7718 & ~w7719;
assign w7721 = w7382 & ~w7720;
assign w7722 = ~w7382 & w7720;
assign w7723 = ~w7721 & ~w7722;
assign w7724 = w7715 & ~w7723;
assign w7725 = ~w7715 & w7723;
assign w7726 = ~w7724 & ~w7725;
assign w7727 = ~w7693 & w7726;
assign w7728 = w7693 & ~w7726;
assign w7729 = ~w7727 & ~w7728;
assign w7730 = ~w7692 & w7729;
assign w7731 = w7692 & ~w7729;
assign w7732 = ~w7730 & ~w7731;
assign w7733 = w7691 & w7732;
assign w7734 = ~w7691 & ~w7732;
assign w7735 = ~w7733 & ~w7734;
assign w7736 = ~w7650 & w7735;
assign w7737 = w7650 & ~w7735;
assign w7738 = ~w7736 & ~w7737;
assign w7739 = ~w7649 & w7738;
assign w7740 = w7649 & ~w7738;
assign w7741 = ~w7739 & ~w7740;
assign w7742 = w7648 & w7741;
assign w7743 = ~w7648 & ~w7741;
assign w7744 = ~w7742 & ~w7743;
assign w7745 = ~w7504 & w7744;
assign w7746 = w7504 & ~w7744;
assign w7747 = ~w7745 & ~w7746;
assign w7748 = (w7006 & w16546) | (w7006 & w16547) | (w16546 & w16547);
assign w7749 = ~w7496 & ~w7748;
assign w7750 = w7747 & w7749;
assign w7751 = ~w7747 & ~w7749;
assign w7752 = ~w7750 & ~w7751;
assign w7753 = ~w7496 & ~w7746;
assign w7754 = (~w7006 & w16548) | (~w7006 & w16549) | (w16548 & w16549);
assign w7755 = ~w7745 & ~w7754;
assign w7756 = ~w7739 & ~w7742;
assign w7757 = ~w7733 & ~w7736;
assign w7758 = (~w7680 & ~w7682) | (~w7680 & w17575) | (~w7682 & w17575);
assign w7759 = ~w7704 & ~w7708;
assign w7760 = ~w7707 & ~w7759;
assign w7761 = ~w7517 & ~w7521;
assign w7762 = ~w7520 & ~w7761;
assign w7763 = w7760 & w7762;
assign w7764 = ~w7760 & ~w7762;
assign w7765 = ~w7763 & ~w7764;
assign w7766 = pi03 & pi59;
assign w7767 = pi05 & pi57;
assign w7768 = ~w7674 & ~w7767;
assign w7769 = pi05 & pi58;
assign w7770 = w7361 & w7769;
assign w7771 = ~w7768 & ~w7770;
assign w7772 = w7766 & ~w7771;
assign w7773 = ~w7766 & w7771;
assign w7774 = ~w7772 & ~w7773;
assign w7775 = ~w7765 & w7774;
assign w7776 = w7765 & ~w7774;
assign w7777 = ~w7775 & ~w7776;
assign w7778 = (~w7713 & ~w7715) | (~w7713 & w17576) | (~w7715 & w17576);
assign w7779 = w7777 & ~w7778;
assign w7780 = ~w7777 & w7778;
assign w7781 = ~w7779 & ~w7780;
assign w7782 = w7758 & ~w7781;
assign w7783 = ~w7758 & w7781;
assign w7784 = ~w7782 & ~w7783;
assign w7785 = (~w7611 & ~w7613) | (~w7611 & w17772) | (~w7613 & w17772);
assign w7786 = (~w7592 & ~w7594) | (~w7592 & w17144) | (~w7594 & w17144);
assign w7787 = ~pi60 & w7296;
assign w7788 = ~w7660 & ~w7787;
assign w7789 = ~w7786 & ~w7788;
assign w7790 = w7786 & w7788;
assign w7791 = ~w7789 & ~w7790;
assign w7792 = w7785 & ~w7791;
assign w7793 = ~w7785 & w7791;
assign w7794 = ~w7792 & ~w7793;
assign w7795 = (w7542 & w17577) | (w7542 & w17578) | (w17577 & w17578);
assign w7796 = (~w7542 & w17579) | (~w7542 & w17580) | (w17579 & w17580);
assign w7797 = ~w7795 & ~w7796;
assign w7798 = w7784 & w7797;
assign w7799 = ~w7784 & ~w7797;
assign w7800 = ~w7798 & ~w7799;
assign w7801 = ~w7757 & w7800;
assign w7802 = w7757 & ~w7800;
assign w7803 = ~w7801 & ~w7802;
assign w7804 = ~w7686 & ~w7689;
assign w7805 = pi19 & pi43;
assign w7806 = pi18 & pi44;
assign w7807 = ~w7698 & ~w7806;
assign w7808 = w7698 & w7806;
assign w7809 = ~w7807 & ~w7808;
assign w7810 = w7805 & ~w7809;
assign w7811 = ~w7805 & w7809;
assign w7812 = ~w7810 & ~w7811;
assign w7813 = pi27 & pi35;
assign w7814 = pi28 & pi34;
assign w7815 = pi29 & pi33;
assign w7816 = ~w7814 & ~w7815;
assign w7817 = w7814 & w7815;
assign w7818 = ~w7816 & ~w7817;
assign w7819 = w7813 & ~w7818;
assign w7820 = ~w7813 & w7818;
assign w7821 = ~w7819 & ~w7820;
assign w7822 = ~w7812 & ~w7821;
assign w7823 = w7812 & w7821;
assign w7824 = ~w7822 & ~w7823;
assign w7825 = pi22 & pi40;
assign w7826 = pi23 & pi39;
assign w7827 = pi24 & pi38;
assign w7828 = ~w7826 & ~w7827;
assign w7829 = pi24 & pi39;
assign w7830 = w7671 & w7829;
assign w7831 = ~w7828 & ~w7830;
assign w7832 = w7825 & ~w7831;
assign w7833 = ~w7825 & w7831;
assign w7834 = ~w7832 & ~w7833;
assign w7835 = w7824 & ~w7834;
assign w7836 = ~w7824 & w7834;
assign w7837 = ~w7835 & ~w7836;
assign w7838 = pi31 & w7654;
assign w7839 = pi00 & pi62;
assign w7840 = pi02 & pi60;
assign w7841 = ~w7839 & ~w7840;
assign w7842 = pi02 & pi62;
assign w7843 = w7289 & w7842;
assign w7844 = ~w7841 & ~w7843;
assign w7845 = w7838 & ~w7844;
assign w7846 = ~w7838 & w7844;
assign w7847 = ~w7845 & ~w7846;
assign w7848 = pi25 & pi37;
assign w7849 = pi26 & pi36;
assign w7850 = ~w7848 & ~w7849;
assign w7851 = w7848 & w7849;
assign w7852 = ~w7850 & ~w7851;
assign w7853 = w7547 & ~w7852;
assign w7854 = ~w7547 & w7852;
assign w7855 = ~w7853 & ~w7854;
assign w7856 = ~w7847 & ~w7855;
assign w7857 = w7847 & w7855;
assign w7858 = ~w7856 & ~w7857;
assign w7859 = pi09 & pi53;
assign w7860 = pi17 & pi45;
assign w7861 = pi10 & pi52;
assign w7862 = ~w7860 & ~w7861;
assign w7863 = w7860 & w7861;
assign w7864 = ~w7862 & ~w7863;
assign w7865 = w7859 & ~w7864;
assign w7866 = ~w7859 & w7864;
assign w7867 = ~w7865 & ~w7866;
assign w7868 = w7858 & ~w7867;
assign w7869 = ~w7858 & w7867;
assign w7870 = ~w7868 & ~w7869;
assign w7871 = pi12 & pi50;
assign w7872 = pi13 & pi49;
assign w7873 = pi14 & pi48;
assign w7874 = ~w7872 & ~w7873;
assign w7875 = pi14 & pi49;
assign w7876 = w7320 & w7875;
assign w7877 = ~w7874 & ~w7876;
assign w7878 = w7871 & ~w7877;
assign w7879 = ~w7871 & w7877;
assign w7880 = ~w7878 & ~w7879;
assign w7881 = pi16 & pi46;
assign w7882 = pi15 & pi47;
assign w7883 = pi11 & pi51;
assign w7884 = ~w7882 & ~w7883;
assign w7885 = w7882 & w7883;
assign w7886 = ~w7884 & ~w7885;
assign w7887 = w7881 & ~w7886;
assign w7888 = ~w7881 & w7886;
assign w7889 = ~w7887 & ~w7888;
assign w7890 = ~w7880 & ~w7889;
assign w7891 = w7880 & w7889;
assign w7892 = ~w7890 & ~w7891;
assign w7893 = pi20 & pi42;
assign w7894 = pi06 & pi56;
assign w7895 = pi07 & pi55;
assign w7896 = ~w7894 & ~w7895;
assign w7897 = pi07 & pi56;
assign w7898 = w7543 & w7897;
assign w7899 = ~w7896 & ~w7898;
assign w7900 = w7893 & ~w7899;
assign w7901 = ~w7893 & w7899;
assign w7902 = ~w7900 & ~w7901;
assign w7903 = w7892 & ~w7902;
assign w7904 = ~w7892 & w7902;
assign w7905 = ~w7903 & ~w7904;
assign w7906 = w7870 & w7905;
assign w7907 = ~w7870 & ~w7905;
assign w7908 = ~w7906 & ~w7907;
assign w7909 = w7837 & w7908;
assign w7910 = ~w7837 & ~w7908;
assign w7911 = ~w7909 & ~w7910;
assign w7912 = ~w7804 & w7911;
assign w7913 = w7804 & ~w7911;
assign w7914 = ~w7912 & ~w7913;
assign w7915 = ~w7637 & ~w7640;
assign w7916 = w7914 & w7915;
assign w7917 = ~w7914 & ~w7915;
assign w7918 = ~w7916 & ~w7917;
assign w7919 = ~w7803 & ~w7918;
assign w7920 = w7803 & w7918;
assign w7921 = ~w7919 & ~w7920;
assign w7922 = ~w7643 & ~w7646;
assign w7923 = (~w7526 & ~w7528) | (~w7526 & w17581) | (~w7528 & w17581);
assign w7924 = (~w7623 & ~w7625) | (~w7623 & w17146) | (~w7625 & w17146);
assign w7925 = (~w7562 & ~w7564) | (~w7562 & w16912) | (~w7564 & w16912);
assign w7926 = ~w7924 & ~w7925;
assign w7927 = w7924 & w7925;
assign w7928 = ~w7926 & ~w7927;
assign w7929 = w7923 & ~w7928;
assign w7930 = ~w7923 & w7928;
assign w7931 = ~w7929 & ~w7930;
assign w7932 = ~w7553 & ~w7557;
assign w7933 = ~w7556 & ~w7932;
assign w7934 = w7543 & ~w7546;
assign w7935 = ~w7548 & ~w7934;
assign w7936 = w7933 & ~w7935;
assign w7937 = ~w7933 & w7935;
assign w7938 = ~w7936 & ~w7937;
assign w7939 = w7694 & ~w7697;
assign w7940 = ~w7699 & ~w7939;
assign w7941 = ~w7938 & w7940;
assign w7942 = w7938 & ~w7940;
assign w7943 = ~w7941 & ~w7942;
assign w7944 = ~w7382 & ~w7719;
assign w7945 = ~w7718 & ~w7944;
assign w7946 = w7671 & ~w7673;
assign w7947 = ~w7675 & ~w7946;
assign w7948 = w7945 & ~w7947;
assign w7949 = ~w7945 & w7947;
assign w7950 = ~w7948 & ~w7949;
assign w7951 = ~w7370 & ~w7568;
assign w7952 = ~w7567 & ~w7951;
assign w7953 = ~w7950 & ~w7952;
assign w7954 = w7950 & w7952;
assign w7955 = ~w7953 & ~w7954;
assign w7956 = pi30 & pi32;
assign w7957 = pi01 & pi61;
assign w7958 = ~w7956 & ~w7957;
assign w7959 = w7956 & w7957;
assign w7960 = ~w7958 & ~w7959;
assign w7961 = ~w7320 & ~w7532;
assign w7962 = ~w7531 & ~w7961;
assign w7963 = w7960 & w7962;
assign w7964 = ~w7960 & ~w7962;
assign w7965 = ~w7963 & ~w7964;
assign w7966 = ~w7508 & ~w7512;
assign w7967 = ~w7511 & ~w7966;
assign w7968 = w7965 & w7967;
assign w7969 = ~w7965 & ~w7967;
assign w7970 = ~w7968 & ~w7969;
assign w7971 = w7955 & w7970;
assign w7972 = ~w7955 & ~w7970;
assign w7973 = ~w7971 & ~w7972;
assign w7974 = ~w7943 & ~w7973;
assign w7975 = w7943 & w7973;
assign w7976 = ~w7974 & ~w7975;
assign w7977 = ~w7931 & ~w7976;
assign w7978 = w7931 & w7976;
assign w7979 = ~w7977 & ~w7978;
assign w7980 = ~w7727 & ~w7730;
assign w7981 = ~w7979 & w7980;
assign w7982 = w7979 & ~w7980;
assign w7983 = ~w7981 & ~w7982;
assign w7984 = ~w7600 & ~w7604;
assign w7985 = (~w7631 & ~w7633) | (~w7631 & w17773) | (~w7633 & w17773);
assign w7986 = ~w7663 & ~w7666;
assign w7987 = ~w7985 & ~w7986;
assign w7988 = w7985 & w7986;
assign w7989 = ~w7987 & ~w7988;
assign w7990 = w7984 & ~w7989;
assign w7991 = ~w7984 & w7989;
assign w7992 = ~w7990 & ~w7991;
assign w7993 = (~w7579 & ~w7581) | (~w7579 & w17774) | (~w7581 & w17774);
assign w7994 = ~w7992 & w7993;
assign w7995 = w7992 & ~w7993;
assign w7996 = ~w7994 & ~w7995;
assign w7997 = w7983 & w7996;
assign w7998 = ~w7983 & ~w7996;
assign w7999 = ~w7997 & ~w7998;
assign w8000 = ~w7922 & w7999;
assign w8001 = w7922 & ~w7999;
assign w8002 = ~w8000 & ~w8001;
assign w8003 = w7921 & w8002;
assign w8004 = ~w7921 & ~w8002;
assign w8005 = ~w8003 & ~w8004;
assign w8006 = ~w7756 & w8005;
assign w8007 = w7756 & ~w8005;
assign w8008 = ~w8006 & ~w8007;
assign w8009 = w7755 & w8008;
assign w8010 = ~w7755 & ~w8008;
assign w8011 = ~w8009 & ~w8010;
assign w8012 = ~w7745 & ~w8006;
assign w8013 = (~w7006 & w17775) | (~w7006 & w17776) | (w17775 & w17776);
assign w8014 = ~w8000 & ~w8003;
assign w8015 = ~w7995 & ~w7997;
assign w8016 = ~w7987 & ~w7991;
assign w8017 = ~w7813 & ~w7817;
assign w8018 = ~w7816 & ~w8017;
assign w8019 = ~w7859 & ~w7863;
assign w8020 = ~w7862 & ~w8019;
assign w8021 = w8018 & w8020;
assign w8022 = ~w8018 & ~w8020;
assign w8023 = ~w8021 & ~w8022;
assign w8024 = ~w7805 & ~w7808;
assign w8025 = ~w7807 & ~w8024;
assign w8026 = ~w8023 & ~w8025;
assign w8027 = w8023 & w8025;
assign w8028 = ~w8026 & ~w8027;
assign w8029 = (~w7822 & ~w7824) | (~w7822 & w16754) | (~w7824 & w16754);
assign w8030 = ~w8028 & w8029;
assign w8031 = w8028 & ~w8029;
assign w8032 = ~w8030 & ~w8031;
assign w8033 = (~w7890 & ~w7892) | (~w7890 & w17147) | (~w7892 & w17147);
assign w8034 = ~w8032 & w8033;
assign w8035 = w8032 & ~w8033;
assign w8036 = ~w8034 & ~w8035;
assign w8037 = pi00 & pi63;
assign w8038 = w7959 & w8037;
assign w8039 = ~w7959 & ~w8037;
assign w8040 = ~w8038 & ~w8039;
assign w8041 = pi01 & pi62;
assign w8042 = pi32 & ~w8041;
assign w8043 = ~pi32 & w8041;
assign w8044 = ~w8042 & ~w8043;
assign w8045 = w8040 & ~w8044;
assign w8046 = ~w8040 & w8044;
assign w8047 = ~w8045 & ~w8046;
assign w8048 = pi26 & pi37;
assign w8049 = pi25 & pi38;
assign w8050 = ~w8048 & ~w8049;
assign w8051 = pi26 & pi38;
assign w8052 = w7848 & w8051;
assign w8053 = ~w8050 & ~w8052;
assign w8054 = w7829 & ~w8053;
assign w8055 = ~w7829 & w8053;
assign w8056 = ~w8054 & ~w8055;
assign w8057 = pi27 & pi36;
assign w8058 = pi29 & pi34;
assign w8059 = pi28 & pi35;
assign w8060 = ~w8058 & ~w8059;
assign w8061 = pi29 & pi35;
assign w8062 = w7814 & w8061;
assign w8063 = ~w8060 & ~w8062;
assign w8064 = w8057 & ~w8063;
assign w8065 = ~w8057 & w8063;
assign w8066 = ~w8064 & ~w8065;
assign w8067 = ~w8056 & ~w8066;
assign w8068 = w8056 & w8066;
assign w8069 = ~w8067 & ~w8068;
assign w8070 = w8047 & w8069;
assign w8071 = ~w8047 & ~w8069;
assign w8072 = ~w8070 & ~w8071;
assign w8073 = (~w7789 & ~w7791) | (~w7789 & w17582) | (~w7791 & w17582);
assign w8074 = ~w7856 & ~w7868;
assign w8075 = ~w8073 & ~w8074;
assign w8076 = w8073 & w8074;
assign w8077 = ~w8075 & ~w8076;
assign w8078 = ~w8072 & ~w8077;
assign w8079 = w8072 & w8077;
assign w8080 = ~w8078 & ~w8079;
assign w8081 = ~w8036 & ~w8080;
assign w8082 = w8036 & w8080;
assign w8083 = ~w8081 & ~w8082;
assign w8084 = ~w8016 & w8083;
assign w8085 = w8016 & ~w8083;
assign w8086 = ~w8084 & ~w8085;
assign w8087 = ~w8015 & w8086;
assign w8088 = w8015 & ~w8086;
assign w8089 = ~w8087 & ~w8088;
assign w8090 = ~w7978 & ~w7982;
assign w8091 = (~w7795 & ~w7797) | (~w7795 & w17777) | (~w7797 & w17777);
assign w8092 = pi31 & pi32;
assign w8093 = pi30 & pi33;
assign w8094 = ~w8092 & ~w8093;
assign w8095 = w8092 & w8093;
assign w8096 = ~w8094 & ~w8095;
assign w8097 = w7875 & ~w8096;
assign w8098 = ~w7875 & w8096;
assign w8099 = ~w8097 & ~w8098;
assign w8100 = pi23 & pi40;
assign w8101 = pi06 & pi57;
assign w8102 = pi20 & pi43;
assign w8103 = ~w8101 & ~w8102;
assign w8104 = w8101 & w8102;
assign w8105 = ~w8103 & ~w8104;
assign w8106 = w8100 & ~w8105;
assign w8107 = ~w8100 & w8105;
assign w8108 = ~w8106 & ~w8107;
assign w8109 = ~w8099 & ~w8108;
assign w8110 = w8099 & w8108;
assign w8111 = ~w8109 & ~w8110;
assign w8112 = pi08 & pi55;
assign w8113 = pi19 & pi44;
assign w8114 = ~w8112 & ~w8113;
assign w8115 = w8112 & w8113;
assign w8116 = ~w8114 & ~w8115;
assign w8117 = w7897 & ~w8116;
assign w8118 = ~w7897 & w8116;
assign w8119 = ~w8117 & ~w8118;
assign w8120 = w8111 & ~w8119;
assign w8121 = ~w8111 & w8119;
assign w8122 = ~w8120 & ~w8121;
assign w8123 = ~w7881 & ~w7885;
assign w8124 = ~w7884 & ~w8123;
assign w8125 = pi02 & pi61;
assign w8126 = pi03 & pi60;
assign w8127 = pi04 & pi59;
assign w8128 = ~w8126 & ~w8127;
assign w8129 = pi04 & pi60;
assign w8130 = w7766 & w8129;
assign w8131 = ~w8128 & ~w8130;
assign w8132 = w8125 & ~w8131;
assign w8133 = ~w8125 & w8131;
assign w8134 = ~w8132 & ~w8133;
assign w8135 = w8124 & ~w8134;
assign w8136 = ~w8124 & w8134;
assign w8137 = ~w8135 & ~w8136;
assign w8138 = pi22 & pi41;
assign w8139 = pi21 & pi42;
assign w8140 = ~w8138 & ~w8139;
assign w8141 = pi22 & pi42;
assign w8142 = w7547 & w8141;
assign w8143 = ~w8140 & ~w8142;
assign w8144 = w7769 & ~w8143;
assign w8145 = ~w7769 & w8143;
assign w8146 = ~w8144 & ~w8145;
assign w8147 = w8137 & ~w8146;
assign w8148 = ~w8137 & w8146;
assign w8149 = ~w8147 & ~w8148;
assign w8150 = w8122 & w8149;
assign w8151 = ~w8122 & ~w8149;
assign w8152 = ~w8150 & ~w8151;
assign w8153 = pi18 & pi45;
assign w8154 = pi17 & pi46;
assign w8155 = pi09 & pi54;
assign w8156 = ~w8154 & ~w8155;
assign w8157 = w8154 & w8155;
assign w8158 = ~w8156 & ~w8157;
assign w8159 = w8153 & ~w8158;
assign w8160 = ~w8153 & w8158;
assign w8161 = ~w8159 & ~w8160;
assign w8162 = pi10 & pi53;
assign w8163 = pi16 & pi47;
assign w8164 = pi11 & pi52;
assign w8165 = ~w8163 & ~w8164;
assign w8166 = w8163 & w8164;
assign w8167 = ~w8165 & ~w8166;
assign w8168 = w8162 & ~w8167;
assign w8169 = ~w8162 & w8167;
assign w8170 = ~w8168 & ~w8169;
assign w8171 = ~w8161 & ~w8170;
assign w8172 = w8161 & w8170;
assign w8173 = ~w8171 & ~w8172;
assign w8174 = pi15 & pi48;
assign w8175 = pi12 & pi51;
assign w8176 = pi13 & pi50;
assign w8177 = ~w8175 & ~w8176;
assign w8178 = pi13 & pi51;
assign w8179 = w7871 & w8178;
assign w8180 = ~w8177 & ~w8179;
assign w8181 = w8174 & ~w8180;
assign w8182 = ~w8174 & w8180;
assign w8183 = ~w8181 & ~w8182;
assign w8184 = w8173 & ~w8183;
assign w8185 = ~w8173 & w8183;
assign w8186 = ~w8184 & ~w8185;
assign w8187 = w8152 & w8186;
assign w8188 = ~w8152 & ~w8186;
assign w8189 = ~w8187 & ~w8188;
assign w8190 = ~w8091 & w8189;
assign w8191 = w8091 & ~w8189;
assign w8192 = ~w8190 & ~w8191;
assign w8193 = ~w8090 & w8192;
assign w8194 = w8090 & ~w8192;
assign w8195 = ~w8193 & ~w8194;
assign w8196 = ~w8089 & ~w8195;
assign w8197 = w8089 & w8195;
assign w8198 = ~w8196 & ~w8197;
assign w8199 = ~w7801 & ~w7920;
assign w8200 = ~w7912 & ~w7916;
assign w8201 = ~w7779 & ~w7783;
assign w8202 = (~w7971 & ~w7973) | (~w7971 & w17148) | (~w7973 & w17148);
assign w8203 = (~w7926 & ~w7928) | (~w7926 & w17149) | (~w7928 & w17149);
assign w8204 = ~w8202 & ~w8203;
assign w8205 = w8202 & w8203;
assign w8206 = ~w8204 & ~w8205;
assign w8207 = w8201 & ~w8206;
assign w8208 = ~w8201 & w8206;
assign w8209 = ~w8207 & ~w8208;
assign w8210 = (~w7963 & ~w7965) | (~w7963 & w17583) | (~w7965 & w17583);
assign w8211 = (~w7763 & ~w7765) | (~w7763 & w16913) | (~w7765 & w16913);
assign w8212 = (~w7948 & ~w7950) | (~w7948 & w16914) | (~w7950 & w16914);
assign w8213 = ~w8211 & ~w8212;
assign w8214 = w8211 & w8212;
assign w8215 = ~w8213 & ~w8214;
assign w8216 = w8210 & ~w8215;
assign w8217 = ~w8210 & w8215;
assign w8218 = ~w8216 & ~w8217;
assign w8219 = (~w7906 & ~w7908) | (~w7906 & w17584) | (~w7908 & w17584);
assign w8220 = ~w8218 & w8219;
assign w8221 = w8218 & ~w8219;
assign w8222 = ~w8220 & ~w8221;
assign w8223 = w7825 & ~w7828;
assign w8224 = ~w7830 & ~w8223;
assign w8225 = w7893 & ~w7896;
assign w8226 = ~w7898 & ~w8225;
assign w8227 = ~w8224 & ~w8226;
assign w8228 = w8224 & w8226;
assign w8229 = ~w8227 & ~w8228;
assign w8230 = w7871 & ~w7874;
assign w8231 = ~w7876 & ~w8230;
assign w8232 = ~w8229 & w8231;
assign w8233 = w8229 & ~w8231;
assign w8234 = ~w8232 & ~w8233;
assign w8235 = ~w7547 & ~w7851;
assign w8236 = ~w7850 & ~w8235;
assign w8237 = w7766 & ~w7768;
assign w8238 = ~w7770 & ~w8237;
assign w8239 = w8236 & ~w8238;
assign w8240 = ~w8236 & w8238;
assign w8241 = ~w8239 & ~w8240;
assign w8242 = w7838 & ~w7841;
assign w8243 = ~w7843 & ~w8242;
assign w8244 = ~w8241 & w8243;
assign w8245 = w8241 & ~w8243;
assign w8246 = ~w8244 & ~w8245;
assign w8247 = (~w7936 & ~w7938) | (~w7936 & w16915) | (~w7938 & w16915);
assign w8248 = ~w8246 & w8247;
assign w8249 = w8246 & ~w8247;
assign w8250 = ~w8248 & ~w8249;
assign w8251 = w8234 & w8250;
assign w8252 = ~w8234 & ~w8250;
assign w8253 = ~w8251 & ~w8252;
assign w8254 = w8222 & w8253;
assign w8255 = ~w8222 & ~w8253;
assign w8256 = ~w8254 & ~w8255;
assign w8257 = ~w8209 & ~w8256;
assign w8258 = w8209 & w8256;
assign w8259 = ~w8257 & ~w8258;
assign w8260 = w8200 & ~w8259;
assign w8261 = ~w8200 & w8259;
assign w8262 = ~w8260 & ~w8261;
assign w8263 = ~w8199 & w8262;
assign w8264 = w8199 & ~w8262;
assign w8265 = ~w8263 & ~w8264;
assign w8266 = ~w8198 & ~w8265;
assign w8267 = w8198 & w8265;
assign w8268 = ~w8266 & ~w8267;
assign w8269 = w8014 & ~w8268;
assign w8270 = ~w8014 & w8268;
assign w8271 = ~w8269 & ~w8270;
assign w8272 = ~w8013 & ~w8271;
assign w8273 = w8013 & w8271;
assign w8274 = ~w8272 & ~w8273;
assign w8275 = w7829 & ~w8050;
assign w8276 = ~w8052 & ~w8275;
assign w8277 = w8174 & ~w8177;
assign w8278 = ~w8179 & ~w8277;
assign w8279 = ~w8276 & ~w8278;
assign w8280 = w8276 & w8278;
assign w8281 = ~w8279 & ~w8280;
assign w8282 = ~w8162 & ~w8166;
assign w8283 = ~w8165 & ~w8282;
assign w8284 = ~w8281 & ~w8283;
assign w8285 = w8281 & w8283;
assign w8286 = ~w8284 & ~w8285;
assign w8287 = (~w8109 & ~w8111) | (~w8109 & w17585) | (~w8111 & w17585);
assign w8288 = ~w8286 & w8287;
assign w8289 = w8286 & ~w8287;
assign w8290 = ~w8288 & ~w8289;
assign w8291 = ~w8171 & ~w8184;
assign w8292 = ~w8290 & w8291;
assign w8293 = w8290 & ~w8291;
assign w8294 = ~w8292 & ~w8293;
assign w8295 = (~w8204 & ~w8206) | (~w8204 & w17586) | (~w8206 & w17586);
assign w8296 = ~w8294 & w8295;
assign w8297 = w8294 & ~w8295;
assign w8298 = ~w8296 & ~w8297;
assign w8299 = ~w7875 & ~w8095;
assign w8300 = ~w8094 & ~w8299;
assign w8301 = pi32 & pi62;
assign w8302 = pi32 & pi63;
assign w8303 = w8041 & w8302;
assign w8304 = (pi01 & w8301) | (pi01 & w16755) | (w8301 & w16755);
assign w8305 = ~w8303 & w8304;
assign w8306 = w8300 & w8305;
assign w8307 = ~w8300 & ~w8305;
assign w8308 = ~w8306 & ~w8307;
assign w8309 = pi11 & pi53;
assign w8310 = pi12 & pi52;
assign w8311 = ~w8309 & ~w8310;
assign w8312 = pi12 & pi53;
assign w8313 = w8164 & w8312;
assign w8314 = ~w8311 & ~w8313;
assign w8315 = w8178 & ~w8314;
assign w8316 = ~w8178 & w8314;
assign w8317 = ~w8315 & ~w8316;
assign w8318 = pi09 & pi55;
assign w8319 = pi15 & pi49;
assign w8320 = pi10 & pi54;
assign w8321 = ~w8319 & ~w8320;
assign w8322 = w8319 & w8320;
assign w8323 = ~w8321 & ~w8322;
assign w8324 = w8318 & ~w8323;
assign w8325 = ~w8318 & w8323;
assign w8326 = ~w8324 & ~w8325;
assign w8327 = ~w8317 & ~w8326;
assign w8328 = w8317 & w8326;
assign w8329 = ~w8327 & ~w8328;
assign w8330 = w8308 & w8329;
assign w8331 = ~w8308 & ~w8329;
assign w8332 = ~w8330 & ~w8331;
assign w8333 = (~w8213 & ~w8215) | (~w8213 & w17150) | (~w8215 & w17150);
assign w8334 = ~w8135 & ~w8147;
assign w8335 = ~w8333 & ~w8334;
assign w8336 = w8333 & w8334;
assign w8337 = ~w8335 & ~w8336;
assign w8338 = ~w8332 & ~w8337;
assign w8339 = w8332 & w8337;
assign w8340 = ~w8338 & ~w8339;
assign w8341 = ~w8298 & ~w8340;
assign w8342 = w8298 & w8340;
assign w8343 = ~w8341 & ~w8342;
assign w8344 = ~w8258 & ~w8261;
assign w8345 = w8343 & ~w8344;
assign w8346 = ~w8343 & w8344;
assign w8347 = ~w8345 & ~w8346;
assign w8348 = (~w8221 & ~w8222) | (~w8221 & w17778) | (~w8222 & w17778);
assign w8349 = pi16 & pi48;
assign w8350 = pi08 & pi56;
assign w8351 = ~w8349 & ~w8350;
assign w8352 = w8349 & w8350;
assign w8353 = ~w8351 & ~w8352;
assign w8354 = w8051 & ~w8353;
assign w8355 = ~w8051 & w8353;
assign w8356 = ~w8354 & ~w8355;
assign w8357 = pi27 & pi37;
assign w8358 = pi28 & pi36;
assign w8359 = ~w8061 & ~w8358;
assign w8360 = w8061 & w8358;
assign w8361 = ~w8359 & ~w8360;
assign w8362 = w8357 & ~w8361;
assign w8363 = ~w8357 & w8361;
assign w8364 = ~w8362 & ~w8363;
assign w8365 = ~w8356 & ~w8364;
assign w8366 = w8356 & w8364;
assign w8367 = ~w8365 & ~w8366;
assign w8368 = pi14 & pi50;
assign w8369 = pi31 & pi33;
assign w8370 = pi30 & pi34;
assign w8371 = ~w8369 & ~w8370;
assign w8372 = w8369 & w8370;
assign w8373 = ~w8371 & ~w8372;
assign w8374 = w8368 & ~w8373;
assign w8375 = ~w8368 & w8373;
assign w8376 = ~w8374 & ~w8375;
assign w8377 = w8367 & ~w8376;
assign w8378 = ~w8367 & w8376;
assign w8379 = ~w8377 & ~w8378;
assign w8380 = (~w8038 & ~w8040) | (~w8038 & w17151) | (~w8040 & w17151);
assign w8381 = pi05 & pi59;
assign w8382 = pi18 & pi46;
assign w8383 = pi19 & pi45;
assign w8384 = ~w8382 & ~w8383;
assign w8385 = pi19 & pi46;
assign w8386 = w8153 & w8385;
assign w8387 = ~w8384 & ~w8386;
assign w8388 = w8381 & ~w8387;
assign w8389 = ~w8381 & w8387;
assign w8390 = ~w8388 & ~w8389;
assign w8391 = ~w8380 & ~w8390;
assign w8392 = w8380 & w8390;
assign w8393 = ~w8391 & ~w8392;
assign w8394 = pi03 & pi61;
assign w8395 = ~w8129 & ~w8394;
assign w8396 = pi04 & pi61;
assign w8397 = w8126 & w8396;
assign w8398 = ~w8395 & ~w8397;
assign w8399 = w7842 & ~w8398;
assign w8400 = ~w7842 & w8398;
assign w8401 = ~w8399 & ~w8400;
assign w8402 = w8393 & ~w8401;
assign w8403 = ~w8393 & w8401;
assign w8404 = ~w8402 & ~w8403;
assign w8405 = w8379 & w8404;
assign w8406 = ~w8379 & ~w8404;
assign w8407 = ~w8405 & ~w8406;
assign w8408 = pi20 & pi44;
assign w8409 = pi21 & pi43;
assign w8410 = ~w8141 & ~w8409;
assign w8411 = pi22 & pi43;
assign w8412 = w8139 & w8411;
assign w8413 = ~w8410 & ~w8412;
assign w8414 = w8408 & ~w8413;
assign w8415 = ~w8408 & w8413;
assign w8416 = ~w8414 & ~w8415;
assign w8417 = pi06 & pi58;
assign w8418 = pi17 & pi47;
assign w8419 = pi07 & pi57;
assign w8420 = ~w8418 & ~w8419;
assign w8421 = w8418 & w8419;
assign w8422 = ~w8420 & ~w8421;
assign w8423 = w8417 & ~w8422;
assign w8424 = ~w8417 & w8422;
assign w8425 = ~w8423 & ~w8424;
assign w8426 = ~w8416 & ~w8425;
assign w8427 = w8416 & w8425;
assign w8428 = ~w8426 & ~w8427;
assign w8429 = pi23 & pi41;
assign w8430 = pi24 & pi40;
assign w8431 = pi25 & pi39;
assign w8432 = ~w8430 & ~w8431;
assign w8433 = w8430 & w8431;
assign w8434 = ~w8432 & ~w8433;
assign w8435 = w8429 & ~w8434;
assign w8436 = ~w8429 & w8434;
assign w8437 = ~w8435 & ~w8436;
assign w8438 = w8428 & ~w8437;
assign w8439 = ~w8428 & w8437;
assign w8440 = ~w8438 & ~w8439;
assign w8441 = w8407 & w8440;
assign w8442 = ~w8407 & ~w8440;
assign w8443 = ~w8441 & ~w8442;
assign w8444 = ~w8348 & w8443;
assign w8445 = w8348 & ~w8443;
assign w8446 = ~w8444 & ~w8445;
assign w8447 = (~w8239 & ~w8241) | (~w8239 & w17152) | (~w8241 & w17152);
assign w8448 = (~w8227 & ~w8229) | (~w8227 & w16756) | (~w8229 & w16756);
assign w8449 = (~w8021 & ~w8023) | (~w8021 & w16757) | (~w8023 & w16757);
assign w8450 = ~w8448 & ~w8449;
assign w8451 = w8448 & w8449;
assign w8452 = ~w8450 & ~w8451;
assign w8453 = w8447 & ~w8452;
assign w8454 = ~w8447 & w8452;
assign w8455 = ~w8453 & ~w8454;
assign w8456 = (~w8031 & ~w8032) | (~w8031 & w16916) | (~w8032 & w16916);
assign w8457 = (~w8249 & ~w8250) | (~w8249 & w16917) | (~w8250 & w16917);
assign w8458 = ~w8456 & ~w8457;
assign w8459 = w8456 & w8457;
assign w8460 = ~w8458 & ~w8459;
assign w8461 = w8455 & w8460;
assign w8462 = ~w8455 & ~w8460;
assign w8463 = ~w8461 & ~w8462;
assign w8464 = w8446 & w8463;
assign w8465 = ~w8446 & ~w8463;
assign w8466 = ~w8464 & ~w8465;
assign w8467 = w8347 & w8466;
assign w8468 = ~w8347 & ~w8466;
assign w8469 = ~w8467 & ~w8468;
assign w8470 = ~w8087 & ~w8197;
assign w8471 = ~w8190 & ~w8193;
assign w8472 = (~w8082 & ~w8083) | (~w8082 & w17779) | (~w8083 & w17779);
assign w8473 = ~w8067 & ~w8070;
assign w8474 = ~w8153 & ~w8157;
assign w8475 = ~w8156 & ~w8474;
assign w8476 = ~w8100 & ~w8104;
assign w8477 = ~w8103 & ~w8476;
assign w8478 = w8475 & w8477;
assign w8479 = ~w8475 & ~w8477;
assign w8480 = ~w8478 & ~w8479;
assign w8481 = w8057 & ~w8060;
assign w8482 = ~w8062 & ~w8481;
assign w8483 = ~w8480 & w8482;
assign w8484 = w8480 & ~w8482;
assign w8485 = ~w8483 & ~w8484;
assign w8486 = w8125 & ~w8128;
assign w8487 = ~w8130 & ~w8486;
assign w8488 = w7769 & ~w8140;
assign w8489 = ~w8142 & ~w8488;
assign w8490 = ~w8487 & ~w8489;
assign w8491 = w8487 & w8489;
assign w8492 = ~w8490 & ~w8491;
assign w8493 = ~w7897 & ~w8115;
assign w8494 = ~w8114 & ~w8493;
assign w8495 = ~w8492 & ~w8494;
assign w8496 = w8492 & w8494;
assign w8497 = ~w8495 & ~w8496;
assign w8498 = w8485 & w8497;
assign w8499 = ~w8485 & ~w8497;
assign w8500 = ~w8498 & ~w8499;
assign w8501 = ~w8473 & w8500;
assign w8502 = w8473 & ~w8500;
assign w8503 = ~w8501 & ~w8502;
assign w8504 = ~w8150 & ~w8187;
assign w8505 = (~w8075 & ~w8077) | (~w8075 & w17780) | (~w8077 & w17780);
assign w8506 = ~w8504 & ~w8505;
assign w8507 = w8504 & w8505;
assign w8508 = ~w8506 & ~w8507;
assign w8509 = ~w8503 & ~w8508;
assign w8510 = w8503 & w8508;
assign w8511 = ~w8509 & ~w8510;
assign w8512 = ~w8472 & w8511;
assign w8513 = w8472 & ~w8511;
assign w8514 = ~w8512 & ~w8513;
assign w8515 = ~w8471 & w8514;
assign w8516 = w8471 & ~w8514;
assign w8517 = ~w8515 & ~w8516;
assign w8518 = ~w8470 & w8517;
assign w8519 = w8470 & ~w8517;
assign w8520 = ~w8518 & ~w8519;
assign w8521 = w8469 & w8520;
assign w8522 = ~w8469 & ~w8520;
assign w8523 = ~w8521 & ~w8522;
assign w8524 = ~w8263 & ~w8267;
assign w8525 = w8523 & ~w8524;
assign w8526 = ~w8523 & w8524;
assign w8527 = ~w8269 & ~w8526;
assign w8528 = (~w7006 & w17781) | (~w7006 & w17782) | (w17781 & w17782);
assign w8529 = ~w8525 & w8528;
assign w8530 = ~w8525 & ~w8526;
assign w8531 = w8013 & ~w8269;
assign w8532 = ~w8270 & ~w8530;
assign w8533 = ~w8531 & w8532;
assign w8534 = ~w8529 & ~w8533;
assign w8535 = ~w8525 & ~w8528;
assign w8536 = ~w8518 & ~w8521;
assign w8537 = ~w8345 & ~w8467;
assign w8538 = ~w8444 & ~w8464;
assign w8539 = (~w8297 & ~w8298) | (~w8297 & w17783) | (~w8298 & w17783);
assign w8540 = (~w8327 & ~w8329) | (~w8327 & w17587) | (~w8329 & w17587);
assign w8541 = ~w8429 & ~w8433;
assign w8542 = ~w8432 & ~w8541;
assign w8543 = ~w8318 & ~w8322;
assign w8544 = ~w8321 & ~w8543;
assign w8545 = w8542 & w8544;
assign w8546 = ~w8542 & ~w8544;
assign w8547 = ~w8545 & ~w8546;
assign w8548 = ~w8417 & ~w8421;
assign w8549 = ~w8420 & ~w8548;
assign w8550 = ~w8547 & ~w8549;
assign w8551 = w8547 & w8549;
assign w8552 = ~w8550 & ~w8551;
assign w8553 = w7842 & ~w8395;
assign w8554 = ~w8397 & ~w8553;
assign w8555 = w8381 & ~w8384;
assign w8556 = ~w8386 & ~w8555;
assign w8557 = ~w8554 & ~w8556;
assign w8558 = w8554 & w8556;
assign w8559 = ~w8557 & ~w8558;
assign w8560 = ~w8051 & ~w8352;
assign w8561 = ~w8351 & ~w8560;
assign w8562 = ~w8559 & ~w8561;
assign w8563 = w8559 & w8561;
assign w8564 = ~w8562 & ~w8563;
assign w8565 = w8552 & w8564;
assign w8566 = ~w8552 & ~w8564;
assign w8567 = ~w8565 & ~w8566;
assign w8568 = ~w8540 & w8567;
assign w8569 = w8540 & ~w8567;
assign w8570 = ~w8568 & ~w8569;
assign w8571 = (~w8405 & ~w8407) | (~w8405 & w17784) | (~w8407 & w17784);
assign w8572 = (~w8335 & ~w8337) | (~w8335 & w17588) | (~w8337 & w17588);
assign w8573 = ~w8571 & ~w8572;
assign w8574 = w8571 & w8572;
assign w8575 = ~w8573 & ~w8574;
assign w8576 = ~w8570 & ~w8575;
assign w8577 = w8570 & w8575;
assign w8578 = ~w8576 & ~w8577;
assign w8579 = ~w8539 & w8578;
assign w8580 = w8539 & ~w8578;
assign w8581 = ~w8579 & ~w8580;
assign w8582 = ~w8538 & w8581;
assign w8583 = w8538 & ~w8581;
assign w8584 = ~w8582 & ~w8583;
assign w8585 = ~w8537 & w8584;
assign w8586 = w8537 & ~w8584;
assign w8587 = ~w8585 & ~w8586;
assign w8588 = ~w8490 & ~w8496;
assign w8589 = (~w8279 & ~w8281) | (~w8279 & w17785) | (~w8281 & w17785);
assign w8590 = (~w8478 & ~w8480) | (~w8478 & w17786) | (~w8480 & w17786);
assign w8591 = ~w8589 & ~w8590;
assign w8592 = w8589 & w8590;
assign w8593 = ~w8591 & ~w8592;
assign w8594 = w8588 & ~w8593;
assign w8595 = ~w8588 & w8593;
assign w8596 = ~w8594 & ~w8595;
assign w8597 = (~w8498 & ~w8500) | (~w8498 & w17787) | (~w8500 & w17787);
assign w8598 = (~w8289 & ~w8290) | (~w8289 & w17788) | (~w8290 & w17788);
assign w8599 = ~w8597 & ~w8598;
assign w8600 = w8597 & w8598;
assign w8601 = ~w8599 & ~w8600;
assign w8602 = ~w8596 & ~w8601;
assign w8603 = w8596 & w8601;
assign w8604 = ~w8602 & ~w8603;
assign w8605 = ~w8506 & ~w8510;
assign w8606 = pi29 & pi36;
assign w8607 = pi11 & pi54;
assign w8608 = ~w8385 & ~w8607;
assign w8609 = w8385 & w8607;
assign w8610 = ~w8608 & ~w8609;
assign w8611 = w8606 & ~w8610;
assign w8612 = ~w8606 & w8610;
assign w8613 = ~w8611 & ~w8612;
assign w8614 = pi30 & pi35;
assign w8615 = pi31 & pi34;
assign w8616 = pi32 & pi33;
assign w8617 = ~w8615 & ~w8616;
assign w8618 = w8615 & w8616;
assign w8619 = ~w8617 & ~w8618;
assign w8620 = w8614 & ~w8619;
assign w8621 = ~w8614 & w8619;
assign w8622 = ~w8620 & ~w8621;
assign w8623 = ~w8613 & ~w8622;
assign w8624 = w8613 & w8622;
assign w8625 = ~w8623 & ~w8624;
assign w8626 = pi17 & pi48;
assign w8627 = pi03 & pi62;
assign w8628 = ~pi33 & ~w8627;
assign w8629 = pi33 & w8627;
assign w8630 = ~w8628 & ~w8629;
assign w8631 = w8626 & ~w8630;
assign w8632 = ~w8626 & w8630;
assign w8633 = ~w8631 & ~w8632;
assign w8634 = w8625 & ~w8633;
assign w8635 = ~w8625 & w8633;
assign w8636 = ~w8634 & ~w8635;
assign w8637 = (~w8303 & ~w8300) | (~w8303 & w16758) | (~w8300 & w16758);
assign w8638 = pi08 & pi57;
assign w8639 = pi21 & pi44;
assign w8640 = ~w8411 & ~w8639;
assign w8641 = pi22 & pi44;
assign w8642 = w8409 & w8641;
assign w8643 = ~w8640 & ~w8642;
assign w8644 = w8638 & ~w8643;
assign w8645 = ~w8638 & w8643;
assign w8646 = ~w8644 & ~w8645;
assign w8647 = ~w8637 & ~w8646;
assign w8648 = w8637 & w8646;
assign w8649 = ~w8647 & ~w8648;
assign w8650 = pi05 & pi60;
assign w8651 = pi06 & pi59;
assign w8652 = pi07 & pi58;
assign w8653 = ~w8651 & ~w8652;
assign w8654 = pi07 & pi59;
assign w8655 = w8417 & w8654;
assign w8656 = ~w8653 & ~w8655;
assign w8657 = w8650 & ~w8656;
assign w8658 = ~w8650 & w8656;
assign w8659 = ~w8657 & ~w8658;
assign w8660 = w8649 & ~w8659;
assign w8661 = ~w8649 & w8659;
assign w8662 = ~w8660 & ~w8661;
assign w8663 = w8636 & w8662;
assign w8664 = ~w8636 & ~w8662;
assign w8665 = ~w8663 & ~w8664;
assign w8666 = pi23 & pi42;
assign w8667 = pi25 & pi40;
assign w8668 = pi24 & pi41;
assign w8669 = ~w8667 & ~w8668;
assign w8670 = pi25 & pi41;
assign w8671 = w8430 & w8670;
assign w8672 = ~w8669 & ~w8671;
assign w8673 = w8666 & ~w8672;
assign w8674 = ~w8666 & w8672;
assign w8675 = ~w8673 & ~w8674;
assign w8676 = pi09 & pi56;
assign w8677 = pi10 & pi55;
assign w8678 = pi20 & pi45;
assign w8679 = ~w8677 & ~w8678;
assign w8680 = w8677 & w8678;
assign w8681 = ~w8679 & ~w8680;
assign w8682 = w8676 & ~w8681;
assign w8683 = ~w8676 & w8681;
assign w8684 = ~w8682 & ~w8683;
assign w8685 = ~w8675 & ~w8684;
assign w8686 = w8675 & w8684;
assign w8687 = ~w8685 & ~w8686;
assign w8688 = pi26 & pi39;
assign w8689 = pi28 & pi37;
assign w8690 = pi27 & pi38;
assign w8691 = ~w8689 & ~w8690;
assign w8692 = pi28 & pi38;
assign w8693 = w8357 & w8692;
assign w8694 = ~w8691 & ~w8693;
assign w8695 = w8688 & ~w8694;
assign w8696 = ~w8688 & w8694;
assign w8697 = ~w8695 & ~w8696;
assign w8698 = w8687 & ~w8697;
assign w8699 = ~w8687 & w8697;
assign w8700 = ~w8698 & ~w8699;
assign w8701 = w8665 & w8700;
assign w8702 = ~w8665 & ~w8700;
assign w8703 = ~w8701 & ~w8702;
assign w8704 = ~w8605 & w8703;
assign w8705 = w8605 & ~w8703;
assign w8706 = ~w8704 & ~w8705;
assign w8707 = w8604 & w8706;
assign w8708 = ~w8604 & ~w8706;
assign w8709 = ~w8707 & ~w8708;
assign w8710 = ~w8512 & ~w8515;
assign w8711 = pi02 & pi63;
assign w8712 = ~w8396 & ~w8711;
assign w8713 = w8396 & w8711;
assign w8714 = ~w8712 & ~w8713;
assign w8715 = ~w8368 & ~w8372;
assign w8716 = ~w8371 & ~w8715;
assign w8717 = w8714 & w8716;
assign w8718 = ~w8714 & ~w8716;
assign w8719 = ~w8717 & ~w8718;
assign w8720 = pi16 & pi49;
assign w8721 = pi15 & pi50;
assign w8722 = pi14 & pi51;
assign w8723 = ~w8721 & ~w8722;
assign w8724 = pi15 & pi51;
assign w8725 = w8368 & w8724;
assign w8726 = ~w8723 & ~w8725;
assign w8727 = w8720 & ~w8726;
assign w8728 = ~w8720 & w8726;
assign w8729 = ~w8727 & ~w8728;
assign w8730 = pi13 & pi52;
assign w8731 = pi18 & pi47;
assign w8732 = ~w8730 & ~w8731;
assign w8733 = w8730 & w8731;
assign w8734 = ~w8732 & ~w8733;
assign w8735 = w8312 & ~w8734;
assign w8736 = ~w8312 & w8734;
assign w8737 = ~w8735 & ~w8736;
assign w8738 = ~w8729 & ~w8737;
assign w8739 = w8729 & w8737;
assign w8740 = ~w8738 & ~w8739;
assign w8741 = w8719 & w8740;
assign w8742 = ~w8719 & ~w8740;
assign w8743 = ~w8741 & ~w8742;
assign w8744 = (~w8450 & ~w8452) | (~w8450 & w16918) | (~w8452 & w16918);
assign w8745 = ~w8391 & ~w8402;
assign w8746 = ~w8744 & ~w8745;
assign w8747 = w8744 & w8745;
assign w8748 = ~w8746 & ~w8747;
assign w8749 = ~w8743 & ~w8748;
assign w8750 = w8743 & w8748;
assign w8751 = ~w8749 & ~w8750;
assign w8752 = ~w8357 & ~w8360;
assign w8753 = ~w8359 & ~w8752;
assign w8754 = w8408 & ~w8410;
assign w8755 = ~w8412 & ~w8754;
assign w8756 = w8753 & ~w8755;
assign w8757 = ~w8753 & w8755;
assign w8758 = ~w8756 & ~w8757;
assign w8759 = w8178 & ~w8311;
assign w8760 = ~w8313 & ~w8759;
assign w8761 = ~w8758 & w8760;
assign w8762 = w8758 & ~w8760;
assign w8763 = ~w8761 & ~w8762;
assign w8764 = (~w8365 & ~w8367) | (~w8365 & w16919) | (~w8367 & w16919);
assign w8765 = ~w8763 & w8764;
assign w8766 = w8763 & ~w8764;
assign w8767 = ~w8765 & ~w8766;
assign w8768 = (~w8426 & ~w8428) | (~w8426 & w17589) | (~w8428 & w17589);
assign w8769 = ~w8767 & w8768;
assign w8770 = w8767 & ~w8768;
assign w8771 = ~w8769 & ~w8770;
assign w8772 = (~w8458 & ~w8460) | (~w8458 & w17153) | (~w8460 & w17153);
assign w8773 = ~w8771 & w8772;
assign w8774 = w8771 & ~w8772;
assign w8775 = ~w8773 & ~w8774;
assign w8776 = w8751 & w8775;
assign w8777 = ~w8751 & ~w8775;
assign w8778 = ~w8776 & ~w8777;
assign w8779 = ~w8710 & w8778;
assign w8780 = w8710 & ~w8778;
assign w8781 = ~w8779 & ~w8780;
assign w8782 = w8709 & w8781;
assign w8783 = ~w8709 & ~w8781;
assign w8784 = ~w8782 & ~w8783;
assign w8785 = w8587 & w8784;
assign w8786 = ~w8587 & ~w8784;
assign w8787 = ~w8785 & ~w8786;
assign w8788 = ~w8536 & w8787;
assign w8789 = w8536 & ~w8787;
assign w8790 = ~w8788 & ~w8789;
assign w8791 = w8535 & w8790;
assign w8792 = ~w8535 & ~w8790;
assign w8793 = ~w8791 & ~w8792;
assign w8794 = ~w8525 & ~w8788;
assign w8795 = (~w7006 & w17789) | (~w7006 & w17790) | (w17789 & w17790);
assign w8796 = ~w8585 & ~w8785;
assign w8797 = (~w8573 & ~w8575) | (~w8573 & w17791) | (~w8575 & w17791);
assign w8798 = pi03 & pi63;
assign w8799 = pi05 & pi61;
assign w8800 = pi04 & pi62;
assign w8801 = ~w8799 & ~w8800;
assign w8802 = pi05 & pi62;
assign w8803 = w8396 & w8802;
assign w8804 = ~w8801 & ~w8803;
assign w8805 = w8798 & ~w8804;
assign w8806 = ~w8798 & w8804;
assign w8807 = ~w8805 & ~w8806;
assign w8808 = pi27 & pi39;
assign w8809 = pi29 & pi37;
assign w8810 = ~w8692 & ~w8809;
assign w8811 = pi29 & pi38;
assign w8812 = w8689 & w8811;
assign w8813 = ~w8810 & ~w8812;
assign w8814 = w8808 & ~w8813;
assign w8815 = ~w8808 & w8813;
assign w8816 = ~w8814 & ~w8815;
assign w8817 = ~w8807 & ~w8816;
assign w8818 = w8807 & w8816;
assign w8819 = ~w8817 & ~w8818;
assign w8820 = pi11 & pi55;
assign w8821 = pi19 & pi47;
assign w8822 = pi12 & pi54;
assign w8823 = ~w8821 & ~w8822;
assign w8824 = w8821 & w8822;
assign w8825 = ~w8823 & ~w8824;
assign w8826 = w8820 & ~w8825;
assign w8827 = ~w8820 & w8825;
assign w8828 = ~w8826 & ~w8827;
assign w8829 = w8819 & ~w8828;
assign w8830 = ~w8819 & w8828;
assign w8831 = ~w8829 & ~w8830;
assign w8832 = pi20 & pi46;
assign w8833 = pi21 & pi45;
assign w8834 = ~w8641 & ~w8833;
assign w8835 = pi22 & pi45;
assign w8836 = w8639 & w8835;
assign w8837 = ~w8834 & ~w8836;
assign w8838 = w8832 & ~w8837;
assign w8839 = ~w8832 & w8837;
assign w8840 = ~w8838 & ~w8839;
assign w8841 = pi23 & pi43;
assign w8842 = pi09 & pi57;
assign w8843 = pi24 & pi42;
assign w8844 = ~w8842 & ~w8843;
assign w8845 = w8842 & w8843;
assign w8846 = ~w8844 & ~w8845;
assign w8847 = w8841 & ~w8846;
assign w8848 = ~w8841 & w8846;
assign w8849 = ~w8847 & ~w8848;
assign w8850 = ~w8840 & ~w8849;
assign w8851 = w8840 & w8849;
assign w8852 = ~w8850 & ~w8851;
assign w8853 = pi10 & pi56;
assign w8854 = pi26 & pi40;
assign w8855 = ~w8670 & ~w8854;
assign w8856 = pi26 & pi41;
assign w8857 = w8667 & w8856;
assign w8858 = ~w8855 & ~w8857;
assign w8859 = w8853 & ~w8858;
assign w8860 = ~w8853 & w8858;
assign w8861 = ~w8859 & ~w8860;
assign w8862 = w8852 & ~w8861;
assign w8863 = ~w8852 & w8861;
assign w8864 = ~w8862 & ~w8863;
assign w8865 = pi14 & pi52;
assign w8866 = pi31 & pi35;
assign w8867 = pi30 & pi36;
assign w8868 = ~w8866 & ~w8867;
assign w8869 = w8866 & w8867;
assign w8870 = ~w8868 & ~w8869;
assign w8871 = w8865 & ~w8870;
assign w8872 = ~w8865 & w8870;
assign w8873 = ~w8871 & ~w8872;
assign w8874 = pi18 & pi48;
assign w8875 = pi13 & pi53;
assign w8876 = ~w8724 & ~w8875;
assign w8877 = w8724 & w8875;
assign w8878 = ~w8876 & ~w8877;
assign w8879 = w8874 & ~w8878;
assign w8880 = ~w8874 & w8878;
assign w8881 = ~w8879 & ~w8880;
assign w8882 = ~w8873 & ~w8881;
assign w8883 = w8873 & w8881;
assign w8884 = ~w8882 & ~w8883;
assign w8885 = pi32 & pi34;
assign w8886 = pi17 & pi49;
assign w8887 = pi16 & pi50;
assign w8888 = ~w8886 & ~w8887;
assign w8889 = pi17 & pi50;
assign w8890 = w8720 & w8889;
assign w8891 = ~w8888 & ~w8890;
assign w8892 = w8885 & ~w8891;
assign w8893 = ~w8885 & w8891;
assign w8894 = ~w8892 & ~w8893;
assign w8895 = w8884 & ~w8894;
assign w8896 = ~w8884 & w8894;
assign w8897 = ~w8895 & ~w8896;
assign w8898 = w8864 & w8897;
assign w8899 = ~w8864 & ~w8897;
assign w8900 = ~w8898 & ~w8899;
assign w8901 = w8831 & w8900;
assign w8902 = ~w8831 & ~w8900;
assign w8903 = ~w8901 & ~w8902;
assign w8904 = ~w8797 & w8903;
assign w8905 = w8797 & ~w8903;
assign w8906 = ~w8904 & ~w8905;
assign w8907 = ~w8756 & ~w8762;
assign w8908 = (~w8545 & ~w8547) | (~w8545 & w17792) | (~w8547 & w17792);
assign w8909 = (~w8557 & ~w8559) | (~w8557 & w17793) | (~w8559 & w17793);
assign w8910 = ~w8908 & ~w8909;
assign w8911 = w8908 & w8909;
assign w8912 = ~w8910 & ~w8911;
assign w8913 = w8907 & ~w8912;
assign w8914 = ~w8907 & w8912;
assign w8915 = ~w8913 & ~w8914;
assign w8916 = (~w8565 & ~w8567) | (~w8565 & w17154) | (~w8567 & w17154);
assign w8917 = (~w8766 & ~w8767) | (~w8766 & w17155) | (~w8767 & w17155);
assign w8918 = ~w8916 & ~w8917;
assign w8919 = w8916 & w8917;
assign w8920 = ~w8918 & ~w8919;
assign w8921 = ~w8915 & ~w8920;
assign w8922 = w8915 & w8920;
assign w8923 = ~w8921 & ~w8922;
assign w8924 = w8906 & w8923;
assign w8925 = ~w8906 & ~w8923;
assign w8926 = ~w8924 & ~w8925;
assign w8927 = ~w8579 & ~w8582;
assign w8928 = ~w8704 & ~w8707;
assign w8929 = ~w8927 & ~w8928;
assign w8930 = w8927 & w8928;
assign w8931 = ~w8929 & ~w8930;
assign w8932 = w8926 & w8931;
assign w8933 = ~w8926 & ~w8931;
assign w8934 = ~w8932 & ~w8933;
assign w8935 = ~w8779 & ~w8782;
assign w8936 = ~w8599 & ~w8603;
assign w8937 = ~w8591 & ~w8595;
assign w8938 = (~w8713 & ~w8716) | (~w8713 & w17156) | (~w8716 & w17156);
assign w8939 = w8688 & ~w8691;
assign w8940 = ~w8693 & ~w8939;
assign w8941 = ~w8938 & ~w8940;
assign w8942 = w8938 & w8940;
assign w8943 = ~w8941 & ~w8942;
assign w8944 = pi06 & pi60;
assign w8945 = pi08 & pi58;
assign w8946 = ~w8654 & ~w8945;
assign w8947 = pi08 & pi59;
assign w8948 = w8652 & w8947;
assign w8949 = ~w8946 & ~w8948;
assign w8950 = w8944 & ~w8949;
assign w8951 = ~w8944 & w8949;
assign w8952 = ~w8950 & ~w8951;
assign w8953 = ~w8943 & w8952;
assign w8954 = w8943 & ~w8952;
assign w8955 = ~w8953 & ~w8954;
assign w8956 = ~w8738 & ~w8741;
assign w8957 = w8955 & ~w8956;
assign w8958 = ~w8955 & w8956;
assign w8959 = ~w8957 & ~w8958;
assign w8960 = w8937 & ~w8959;
assign w8961 = ~w8937 & w8959;
assign w8962 = ~w8960 & ~w8961;
assign w8963 = ~w8614 & ~w8618;
assign w8964 = ~w8617 & ~w8963;
assign w8965 = ~w8626 & ~w8629;
assign w8966 = ~w8628 & ~w8965;
assign w8967 = w8964 & w8966;
assign w8968 = ~w8964 & ~w8966;
assign w8969 = ~w8967 & ~w8968;
assign w8970 = w8720 & ~w8723;
assign w8971 = ~w8725 & ~w8970;
assign w8972 = ~w8969 & w8971;
assign w8973 = w8969 & ~w8971;
assign w8974 = ~w8972 & ~w8973;
assign w8975 = w8638 & ~w8640;
assign w8976 = ~w8642 & ~w8975;
assign w8977 = w8650 & ~w8653;
assign w8978 = ~w8655 & ~w8977;
assign w8979 = ~w8976 & ~w8978;
assign w8980 = w8976 & w8978;
assign w8981 = ~w8979 & ~w8980;
assign w8982 = ~w8606 & ~w8609;
assign w8983 = ~w8608 & ~w8982;
assign w8984 = ~w8981 & ~w8983;
assign w8985 = w8981 & w8983;
assign w8986 = ~w8984 & ~w8985;
assign w8987 = (~w8623 & ~w8625) | (~w8623 & w16920) | (~w8625 & w16920);
assign w8988 = ~w8986 & w8987;
assign w8989 = w8986 & ~w8987;
assign w8990 = ~w8988 & ~w8989;
assign w8991 = w8974 & w8990;
assign w8992 = ~w8974 & ~w8990;
assign w8993 = ~w8991 & ~w8992;
assign w8994 = w8962 & w8993;
assign w8995 = ~w8962 & ~w8993;
assign w8996 = ~w8994 & ~w8995;
assign w8997 = ~w8936 & w8996;
assign w8998 = w8936 & ~w8996;
assign w8999 = ~w8997 & ~w8998;
assign w9000 = (~w8774 & ~w8775) | (~w8774 & w17590) | (~w8775 & w17590);
assign w9001 = ~w8676 & ~w8680;
assign w9002 = ~w8679 & ~w9001;
assign w9003 = ~w8312 & ~w8733;
assign w9004 = ~w8732 & ~w9003;
assign w9005 = w9002 & w9004;
assign w9006 = ~w9002 & ~w9004;
assign w9007 = ~w9005 & ~w9006;
assign w9008 = w8666 & ~w8669;
assign w9009 = ~w8671 & ~w9008;
assign w9010 = ~w9007 & w9009;
assign w9011 = w9007 & ~w9009;
assign w9012 = ~w9010 & ~w9011;
assign w9013 = (~w8647 & ~w8649) | (~w8647 & w16921) | (~w8649 & w16921);
assign w9014 = ~w9012 & w9013;
assign w9015 = w9012 & ~w9013;
assign w9016 = ~w9014 & ~w9015;
assign w9017 = (~w8685 & ~w8687) | (~w8685 & w17591) | (~w8687 & w17591);
assign w9018 = ~w9016 & w9017;
assign w9019 = w9016 & ~w9017;
assign w9020 = ~w9018 & ~w9019;
assign w9021 = (~w8663 & ~w8665) | (~w8663 & w17592) | (~w8665 & w17592);
assign w9022 = (~w8746 & ~w8748) | (~w8746 & w17157) | (~w8748 & w17157);
assign w9023 = ~w9021 & ~w9022;
assign w9024 = w9021 & w9022;
assign w9025 = ~w9023 & ~w9024;
assign w9026 = w9020 & w9025;
assign w9027 = ~w9020 & ~w9025;
assign w9028 = ~w9026 & ~w9027;
assign w9029 = ~w9000 & w9028;
assign w9030 = w9000 & ~w9028;
assign w9031 = ~w9029 & ~w9030;
assign w9032 = ~w8999 & ~w9031;
assign w9033 = w8999 & w9031;
assign w9034 = ~w9032 & ~w9033;
assign w9035 = ~w8935 & w9034;
assign w9036 = w8935 & ~w9034;
assign w9037 = ~w9035 & ~w9036;
assign w9038 = w8934 & w9037;
assign w9039 = ~w8934 & ~w9037;
assign w9040 = ~w9038 & ~w9039;
assign w9041 = ~w8796 & w9040;
assign w9042 = w8796 & ~w9040;
assign w9043 = ~w9041 & ~w9042;
assign w9044 = w8795 & ~w9043;
assign w9045 = ~w8795 & w9043;
assign w9046 = ~w9044 & ~w9045;
assign w9047 = ~w9035 & ~w9038;
assign w9048 = ~w8929 & ~w8932;
assign w9049 = ~w8994 & ~w8997;
assign w9050 = (~w8918 & ~w8920) | (~w8918 & w17593) | (~w8920 & w17593);
assign w9051 = ~w8817 & ~w8829;
assign w9052 = (~w8850 & ~w8852) | (~w8850 & w17594) | (~w8852 & w17594);
assign w9053 = (~w8941 & ~w8943) | (~w8941 & w17595) | (~w8943 & w17595);
assign w9054 = ~w9052 & ~w9053;
assign w9055 = w9052 & w9053;
assign w9056 = ~w9054 & ~w9055;
assign w9057 = w9051 & ~w9056;
assign w9058 = ~w9051 & w9056;
assign w9059 = ~w9057 & ~w9058;
assign w9060 = w8798 & ~w8801;
assign w9061 = ~w8803 & ~w9060;
assign w9062 = w8944 & ~w8946;
assign w9063 = ~w8948 & ~w9062;
assign w9064 = ~w9061 & ~w9063;
assign w9065 = w9061 & w9063;
assign w9066 = ~w9064 & ~w9065;
assign w9067 = w8808 & ~w8810;
assign w9068 = ~w8812 & ~w9067;
assign w9069 = ~w9066 & w9068;
assign w9070 = w9066 & ~w9068;
assign w9071 = ~w9069 & ~w9070;
assign w9072 = ~w8841 & ~w8845;
assign w9073 = ~w8844 & ~w9072;
assign w9074 = w8853 & ~w8855;
assign w9075 = ~w8857 & ~w9074;
assign w9076 = w9073 & ~w9075;
assign w9077 = ~w9073 & w9075;
assign w9078 = ~w9076 & ~w9077;
assign w9079 = w8832 & ~w8834;
assign w9080 = ~w8836 & ~w9079;
assign w9081 = ~w9078 & w9080;
assign w9082 = w9078 & ~w9080;
assign w9083 = ~w9081 & ~w9082;
assign w9084 = pi06 & pi61;
assign w9085 = w8885 & ~w8888;
assign w9086 = (w9084 & w9085) | (w9084 & w16759) | (w9085 & w16759);
assign w9087 = ~w9085 & w16760;
assign w9088 = ~w9086 & ~w9087;
assign w9089 = ~w8865 & ~w8869;
assign w9090 = ~w8868 & ~w9089;
assign w9091 = ~w9088 & ~w9090;
assign w9092 = w9088 & w9090;
assign w9093 = ~w9091 & ~w9092;
assign w9094 = w9083 & w9093;
assign w9095 = ~w9083 & ~w9093;
assign w9096 = ~w9094 & ~w9095;
assign w9097 = w9071 & w9096;
assign w9098 = ~w9071 & ~w9096;
assign w9099 = ~w9097 & ~w9098;
assign w9100 = w9059 & w9099;
assign w9101 = ~w9059 & ~w9099;
assign w9102 = ~w9100 & ~w9101;
assign w9103 = ~w9050 & w9102;
assign w9104 = w9050 & ~w9102;
assign w9105 = ~w9103 & ~w9104;
assign w9106 = ~w9049 & w9105;
assign w9107 = w9049 & ~w9105;
assign w9108 = ~w9106 & ~w9107;
assign w9109 = ~w8910 & ~w8914;
assign w9110 = ~w8874 & ~w8877;
assign w9111 = ~w8876 & ~w9110;
assign w9112 = ~w8820 & ~w8824;
assign w9113 = ~w8823 & ~w9112;
assign w9114 = w9111 & w9113;
assign w9115 = ~w9111 & ~w9113;
assign w9116 = ~w9114 & ~w9115;
assign w9117 = pi10 & pi57;
assign w9118 = pi11 & pi56;
assign w9119 = pi20 & pi47;
assign w9120 = ~w9118 & ~w9119;
assign w9121 = w9118 & w9119;
assign w9122 = ~w9120 & ~w9121;
assign w9123 = w9117 & ~w9122;
assign w9124 = ~w9117 & w9122;
assign w9125 = ~w9123 & ~w9124;
assign w9126 = ~w9116 & w9125;
assign w9127 = w9116 & ~w9125;
assign w9128 = ~w9126 & ~w9127;
assign w9129 = ~w8882 & ~w8895;
assign w9130 = w9128 & ~w9129;
assign w9131 = ~w9128 & w9129;
assign w9132 = ~w9130 & ~w9131;
assign w9133 = w9109 & ~w9132;
assign w9134 = ~w9109 & w9132;
assign w9135 = ~w9133 & ~w9134;
assign w9136 = ~w8898 & ~w8901;
assign w9137 = ~w8957 & ~w8961;
assign w9138 = ~w9136 & ~w9137;
assign w9139 = w9136 & w9137;
assign w9140 = ~w9138 & ~w9139;
assign w9141 = w9135 & w9140;
assign w9142 = ~w9135 & ~w9140;
assign w9143 = ~w9141 & ~w9142;
assign w9144 = w9108 & w9143;
assign w9145 = ~w9108 & ~w9143;
assign w9146 = ~w9144 & ~w9145;
assign w9147 = ~w9048 & w9146;
assign w9148 = w9048 & ~w9146;
assign w9149 = ~w9147 & ~w9148;
assign w9150 = pi19 & pi48;
assign w9151 = pi14 & pi53;
assign w9152 = ~w8889 & ~w9151;
assign w9153 = w8889 & w9151;
assign w9154 = ~w9152 & ~w9153;
assign w9155 = w9150 & ~w9154;
assign w9156 = ~w9150 & w9154;
assign w9157 = ~w9155 & ~w9156;
assign w9158 = pi25 & pi42;
assign w9159 = pi21 & pi46;
assign w9160 = ~w8856 & ~w9159;
assign w9161 = w8856 & w9159;
assign w9162 = ~w9160 & ~w9161;
assign w9163 = w9158 & ~w9162;
assign w9164 = ~w9158 & w9162;
assign w9165 = ~w9163 & ~w9164;
assign w9166 = ~w9157 & ~w9165;
assign w9167 = w9157 & w9165;
assign w9168 = ~w9166 & ~w9167;
assign w9169 = pi04 & pi63;
assign w9170 = pi27 & pi40;
assign w9171 = pi28 & pi39;
assign w9172 = ~w9170 & ~w9171;
assign w9173 = w9170 & w9171;
assign w9174 = ~w9172 & ~w9173;
assign w9175 = w9169 & ~w9174;
assign w9176 = ~w9169 & w9174;
assign w9177 = ~w9175 & ~w9176;
assign w9178 = w9168 & ~w9177;
assign w9179 = ~w9168 & w9177;
assign w9180 = ~w9178 & ~w9179;
assign w9181 = pi18 & pi49;
assign w9182 = pi62 & w3094;
assign w9183 = ~pi34 & ~w8802;
assign w9184 = ~w9182 & ~w9183;
assign w9185 = w9181 & ~w9184;
assign w9186 = ~w9181 & w9184;
assign w9187 = ~w9185 & ~w9186;
assign w9188 = pi31 & pi36;
assign w9189 = pi33 & pi34;
assign w9190 = pi32 & pi35;
assign w9191 = ~w9189 & ~w9190;
assign w9192 = pi33 & pi35;
assign w9193 = w8885 & w9192;
assign w9194 = ~w9191 & ~w9193;
assign w9195 = w9188 & ~w9194;
assign w9196 = ~w9188 & w9194;
assign w9197 = ~w9195 & ~w9196;
assign w9198 = ~w9187 & ~w9197;
assign w9199 = w9187 & w9197;
assign w9200 = ~w9198 & ~w9199;
assign w9201 = pi12 & pi55;
assign w9202 = pi13 & pi54;
assign w9203 = ~w9201 & ~w9202;
assign w9204 = pi13 & pi55;
assign w9205 = w8822 & w9204;
assign w9206 = ~w9203 & ~w9205;
assign w9207 = w8811 & ~w9206;
assign w9208 = ~w8811 & w9206;
assign w9209 = ~w9207 & ~w9208;
assign w9210 = w9200 & ~w9209;
assign w9211 = ~w9200 & w9209;
assign w9212 = ~w9210 & ~w9211;
assign w9213 = pi07 & pi60;
assign w9214 = pi09 & pi58;
assign w9215 = ~w8947 & ~w9214;
assign w9216 = pi09 & pi59;
assign w9217 = w8945 & w9216;
assign w9218 = ~w9215 & ~w9217;
assign w9219 = w9213 & ~w9218;
assign w9220 = ~w9213 & w9218;
assign w9221 = ~w9219 & ~w9220;
assign w9222 = pi23 & pi44;
assign w9223 = pi24 & pi43;
assign w9224 = ~w9222 & ~w9223;
assign w9225 = pi24 & pi44;
assign w9226 = w8841 & w9225;
assign w9227 = ~w9224 & ~w9226;
assign w9228 = w8835 & ~w9227;
assign w9229 = ~w8835 & w9227;
assign w9230 = ~w9228 & ~w9229;
assign w9231 = ~w9221 & ~w9230;
assign w9232 = w9221 & w9230;
assign w9233 = ~w9231 & ~w9232;
assign w9234 = pi15 & pi52;
assign w9235 = pi16 & pi51;
assign w9236 = pi30 & pi37;
assign w9237 = ~w9235 & ~w9236;
assign w9238 = w9235 & w9236;
assign w9239 = ~w9237 & ~w9238;
assign w9240 = w9234 & ~w9239;
assign w9241 = ~w9234 & w9239;
assign w9242 = ~w9240 & ~w9241;
assign w9243 = w9233 & ~w9242;
assign w9244 = ~w9233 & w9242;
assign w9245 = ~w9243 & ~w9244;
assign w9246 = w9212 & w9245;
assign w9247 = ~w9212 & ~w9245;
assign w9248 = ~w9246 & ~w9247;
assign w9249 = w9180 & w9248;
assign w9250 = ~w9180 & ~w9248;
assign w9251 = ~w9249 & ~w9250;
assign w9252 = (w9025 & w17794) | (w9025 & w17795) | (w17794 & w17795);
assign w9253 = (~w9025 & w17796) | (~w9025 & w17797) | (w17796 & w17797);
assign w9254 = ~w9252 & ~w9253;
assign w9255 = (~w8967 & ~w8969) | (~w8967 & w17798) | (~w8969 & w17798);
assign w9256 = (~w8979 & ~w8981) | (~w8979 & w17158) | (~w8981 & w17158);
assign w9257 = (~w9005 & ~w9007) | (~w9005 & w17159) | (~w9007 & w17159);
assign w9258 = ~w9256 & ~w9257;
assign w9259 = w9256 & w9257;
assign w9260 = ~w9258 & ~w9259;
assign w9261 = w9255 & ~w9260;
assign w9262 = ~w9255 & w9260;
assign w9263 = ~w9261 & ~w9262;
assign w9264 = (~w8989 & ~w8990) | (~w8989 & w17160) | (~w8990 & w17160);
assign w9265 = (~w9015 & ~w9016) | (~w9015 & w17161) | (~w9016 & w17161);
assign w9266 = ~w9264 & ~w9265;
assign w9267 = w9264 & w9265;
assign w9268 = ~w9266 & ~w9267;
assign w9269 = w9263 & w9268;
assign w9270 = ~w9263 & ~w9268;
assign w9271 = ~w9269 & ~w9270;
assign w9272 = w9254 & w9271;
assign w9273 = ~w9254 & ~w9271;
assign w9274 = ~w9272 & ~w9273;
assign w9275 = (~w9029 & ~w9031) | (~w9029 & w17799) | (~w9031 & w17799);
assign w9276 = ~w8904 & ~w8924;
assign w9277 = ~w9275 & ~w9276;
assign w9278 = w9275 & w9276;
assign w9279 = ~w9277 & ~w9278;
assign w9280 = ~w9274 & ~w9279;
assign w9281 = w9274 & w9279;
assign w9282 = ~w9280 & ~w9281;
assign w9283 = w9149 & w9282;
assign w9284 = ~w9149 & ~w9282;
assign w9285 = ~w9283 & ~w9284;
assign w9286 = ~w9047 & w9285;
assign w9287 = w9047 & ~w9285;
assign w9288 = ~w9286 & ~w9287;
assign w9289 = (w7754 & w17800) | (w7754 & w17801) | (w17800 & w17801);
assign w9290 = w9288 & w9289;
assign w9291 = ~w9288 & ~w9289;
assign w9292 = ~w9290 & ~w9291;
assign w9293 = ~w9106 & ~w9144;
assign w9294 = ~w9252 & ~w9272;
assign w9295 = ~w9138 & ~w9141;
assign w9296 = ~w9130 & ~w9134;
assign w9297 = (~w9094 & ~w9096) | (~w9094 & w17802) | (~w9096 & w17802);
assign w9298 = (~w9054 & ~w9056) | (~w9054 & w17803) | (~w9056 & w17803);
assign w9299 = ~w9297 & ~w9298;
assign w9300 = w9297 & w9298;
assign w9301 = ~w9299 & ~w9300;
assign w9302 = w9296 & ~w9301;
assign w9303 = ~w9296 & w9301;
assign w9304 = ~w9302 & ~w9303;
assign w9305 = pi10 & pi58;
assign w9306 = pi11 & pi57;
assign w9307 = ~w9305 & ~w9306;
assign w9308 = pi11 & pi58;
assign w9309 = w9117 & w9308;
assign w9310 = ~w9307 & ~w9309;
assign w9311 = w9216 & ~w9310;
assign w9312 = ~w9216 & w9310;
assign w9313 = ~w9311 & ~w9312;
assign w9314 = pi27 & pi41;
assign w9315 = pi28 & pi40;
assign w9316 = pi29 & pi39;
assign w9317 = ~w9315 & ~w9316;
assign w9318 = w9315 & w9316;
assign w9319 = ~w9317 & ~w9318;
assign w9320 = w9314 & ~w9319;
assign w9321 = ~w9314 & w9319;
assign w9322 = ~w9320 & ~w9321;
assign w9323 = ~w9313 & ~w9322;
assign w9324 = w9313 & w9322;
assign w9325 = ~w9323 & ~w9324;
assign w9326 = pi21 & pi47;
assign w9327 = pi05 & pi63;
assign w9328 = pi06 & pi62;
assign w9329 = ~w9327 & ~w9328;
assign w9330 = pi06 & pi63;
assign w9331 = w8802 & w9330;
assign w9332 = ~w9329 & ~w9331;
assign w9333 = w9326 & ~w9332;
assign w9334 = ~w9326 & w9332;
assign w9335 = ~w9333 & ~w9334;
assign w9336 = w9325 & ~w9335;
assign w9337 = ~w9325 & w9335;
assign w9338 = ~w9336 & ~w9337;
assign w9339 = pi18 & pi50;
assign w9340 = pi19 & pi49;
assign w9341 = ~w9339 & ~w9340;
assign w9342 = pi19 & pi50;
assign w9343 = w9181 & w9342;
assign w9344 = ~w9341 & ~w9343;
assign w9345 = w9192 & ~w9344;
assign w9346 = ~w9192 & w9344;
assign w9347 = ~w9345 & ~w9346;
assign w9348 = pi30 & pi38;
assign w9349 = pi32 & pi36;
assign w9350 = pi31 & pi37;
assign w9351 = ~w9349 & ~w9350;
assign w9352 = w9349 & w9350;
assign w9353 = ~w9351 & ~w9352;
assign w9354 = w9348 & ~w9353;
assign w9355 = ~w9348 & w9353;
assign w9356 = ~w9354 & ~w9355;
assign w9357 = ~w9347 & ~w9356;
assign w9358 = w9347 & w9356;
assign w9359 = ~w9357 & ~w9358;
assign w9360 = pi12 & pi56;
assign w9361 = pi17 & pi51;
assign w9362 = ~w9204 & ~w9361;
assign w9363 = w9204 & w9361;
assign w9364 = ~w9362 & ~w9363;
assign w9365 = w9360 & ~w9364;
assign w9366 = ~w9360 & w9364;
assign w9367 = ~w9365 & ~w9366;
assign w9368 = w9359 & ~w9367;
assign w9369 = ~w9359 & w9367;
assign w9370 = ~w9368 & ~w9369;
assign w9371 = pi14 & pi54;
assign w9372 = pi16 & pi52;
assign w9373 = pi15 & pi53;
assign w9374 = ~w9372 & ~w9373;
assign w9375 = pi16 & pi53;
assign w9376 = w9234 & w9375;
assign w9377 = ~w9374 & ~w9376;
assign w9378 = w9371 & ~w9377;
assign w9379 = ~w9371 & w9377;
assign w9380 = ~w9378 & ~w9379;
assign w9381 = pi20 & pi48;
assign w9382 = pi22 & pi46;
assign w9383 = pi23 & pi45;
assign w9384 = ~w9382 & ~w9383;
assign w9385 = pi23 & pi46;
assign w9386 = w8835 & w9385;
assign w9387 = ~w9384 & ~w9386;
assign w9388 = w9381 & ~w9387;
assign w9389 = ~w9381 & w9387;
assign w9390 = ~w9388 & ~w9389;
assign w9391 = ~w9380 & ~w9390;
assign w9392 = w9380 & w9390;
assign w9393 = ~w9391 & ~w9392;
assign w9394 = pi25 & pi43;
assign w9395 = pi26 & pi42;
assign w9396 = ~w9394 & ~w9395;
assign w9397 = pi26 & pi43;
assign w9398 = w9158 & w9397;
assign w9399 = ~w9396 & ~w9398;
assign w9400 = w9225 & ~w9399;
assign w9401 = ~w9225 & w9399;
assign w9402 = ~w9400 & ~w9401;
assign w9403 = w9393 & ~w9402;
assign w9404 = ~w9393 & w9402;
assign w9405 = ~w9403 & ~w9404;
assign w9406 = w9370 & w9405;
assign w9407 = ~w9370 & ~w9405;
assign w9408 = ~w9406 & ~w9407;
assign w9409 = w9338 & w9408;
assign w9410 = ~w9338 & ~w9408;
assign w9411 = ~w9409 & ~w9410;
assign w9412 = w9304 & w9411;
assign w9413 = ~w9304 & ~w9411;
assign w9414 = ~w9412 & ~w9413;
assign w9415 = ~w9295 & w9414;
assign w9416 = w9295 & ~w9414;
assign w9417 = ~w9415 & ~w9416;
assign w9418 = ~w9294 & w9417;
assign w9419 = w9294 & ~w9417;
assign w9420 = ~w9418 & ~w9419;
assign w9421 = ~w9293 & w9420;
assign w9422 = w9293 & ~w9420;
assign w9423 = ~w9421 & ~w9422;
assign w9424 = ~w9277 & ~w9281;
assign w9425 = (~w9266 & ~w9268) | (~w9266 & w17599) | (~w9268 & w17599);
assign w9426 = ~w9158 & ~w9161;
assign w9427 = ~w9160 & ~w9426;
assign w9428 = ~w9150 & ~w9153;
assign w9429 = ~w9152 & ~w9428;
assign w9430 = w9427 & w9429;
assign w9431 = ~w9427 & ~w9429;
assign w9432 = ~w9430 & ~w9431;
assign w9433 = w8811 & ~w9203;
assign w9434 = ~w9205 & ~w9433;
assign w9435 = ~w9432 & w9434;
assign w9436 = w9432 & ~w9434;
assign w9437 = ~w9435 & ~w9436;
assign w9438 = (~w9166 & ~w9168) | (~w9166 & w17600) | (~w9168 & w17600);
assign w9439 = (~w9198 & ~w9200) | (~w9198 & w17601) | (~w9200 & w17601);
assign w9440 = ~w9438 & ~w9439;
assign w9441 = w9438 & w9439;
assign w9442 = ~w9440 & ~w9441;
assign w9443 = w9437 & w9442;
assign w9444 = ~w9437 & ~w9442;
assign w9445 = ~w9443 & ~w9444;
assign w9446 = (~w9258 & ~w9260) | (~w9258 & w17602) | (~w9260 & w17602);
assign w9447 = ~w9117 & ~w9121;
assign w9448 = ~w9120 & ~w9447;
assign w9449 = w8835 & ~w9224;
assign w9450 = ~w9226 & ~w9449;
assign w9451 = w9448 & ~w9450;
assign w9452 = ~w9448 & w9450;
assign w9453 = ~w9451 & ~w9452;
assign w9454 = w9213 & ~w9215;
assign w9455 = ~w9217 & ~w9454;
assign w9456 = ~w9453 & w9455;
assign w9457 = w9453 & ~w9455;
assign w9458 = ~w9456 & ~w9457;
assign w9459 = ~w9169 & ~w9173;
assign w9460 = ~w9172 & ~w9459;
assign w9461 = w9188 & ~w9191;
assign w9462 = ~w9193 & ~w9461;
assign w9463 = w9460 & ~w9462;
assign w9464 = ~w9460 & w9462;
assign w9465 = ~w9463 & ~w9464;
assign w9466 = ~w9234 & ~w9238;
assign w9467 = ~w9237 & ~w9466;
assign w9468 = ~w9465 & ~w9467;
assign w9469 = w9465 & w9467;
assign w9470 = ~w9468 & ~w9469;
assign w9471 = w9458 & w9470;
assign w9472 = ~w9458 & ~w9470;
assign w9473 = ~w9471 & ~w9472;
assign w9474 = ~w9446 & w9473;
assign w9475 = w9446 & ~w9473;
assign w9476 = ~w9474 & ~w9475;
assign w9477 = w9445 & w9476;
assign w9478 = ~w9445 & ~w9476;
assign w9479 = ~w9477 & ~w9478;
assign w9480 = ~w9425 & w9479;
assign w9481 = w9425 & ~w9479;
assign w9482 = ~w9480 & ~w9481;
assign w9483 = ~w9100 & ~w9103;
assign w9484 = ~w9246 & ~w9249;
assign w9485 = (~w9231 & ~w9233) | (~w9231 & w16922) | (~w9233 & w16922);
assign w9486 = (~w9114 & ~w9116) | (~w9114 & w16761) | (~w9116 & w16761);
assign w9487 = (~w9076 & ~w9078) | (~w9076 & w16762) | (~w9078 & w16762);
assign w9488 = ~w9486 & ~w9487;
assign w9489 = w9486 & w9487;
assign w9490 = ~w9488 & ~w9489;
assign w9491 = w9485 & ~w9490;
assign w9492 = ~w9485 & w9490;
assign w9493 = ~w9491 & ~w9492;
assign w9494 = (~w9064 & ~w9066) | (~w9064 & w17162) | (~w9066 & w17162);
assign w9495 = (~w9086 & ~w9088) | (~w9086 & w16923) | (~w9088 & w16923);
assign w9496 = pi08 & pi60;
assign w9497 = pi07 & pi61;
assign w9498 = ~w9496 & ~w9497;
assign w9499 = pi08 & pi61;
assign w9500 = w9213 & w9499;
assign w9501 = ~w9498 & ~w9500;
assign w9502 = w9181 & ~w9183;
assign w9503 = ~w9182 & ~w9502;
assign w9504 = w9501 & ~w9503;
assign w9505 = ~w9501 & w9503;
assign w9506 = ~w9504 & ~w9505;
assign w9507 = ~w9495 & w9506;
assign w9508 = w9495 & ~w9506;
assign w9509 = ~w9507 & ~w9508;
assign w9510 = w9494 & ~w9509;
assign w9511 = ~w9494 & w9509;
assign w9512 = ~w9510 & ~w9511;
assign w9513 = w9493 & w9512;
assign w9514 = ~w9493 & ~w9512;
assign w9515 = ~w9513 & ~w9514;
assign w9516 = ~w9484 & w9515;
assign w9517 = w9484 & ~w9515;
assign w9518 = ~w9516 & ~w9517;
assign w9519 = ~w9483 & w9518;
assign w9520 = w9483 & ~w9518;
assign w9521 = ~w9519 & ~w9520;
assign w9522 = ~w9482 & ~w9521;
assign w9523 = w9482 & w9521;
assign w9524 = ~w9522 & ~w9523;
assign w9525 = ~w9424 & w9524;
assign w9526 = w9424 & ~w9524;
assign w9527 = ~w9525 & ~w9526;
assign w9528 = w9423 & w9527;
assign w9529 = ~w9423 & ~w9527;
assign w9530 = ~w9528 & ~w9529;
assign w9531 = ~w9147 & ~w9283;
assign w9532 = ~w9530 & w9531;
assign w9533 = w9530 & ~w9531;
assign w9534 = ~w9532 & ~w9533;
assign w9535 = ~w9042 & ~w9287;
assign w9536 = (~w7754 & w17804) | (~w7754 & w17805) | (w17804 & w17805);
assign w9537 = w9534 & w9536;
assign w9538 = ~w9534 & ~w9536;
assign w9539 = ~w9537 & ~w9538;
assign w9540 = ~w9525 & ~w9528;
assign w9541 = ~w9418 & ~w9421;
assign w9542 = ~w9477 & ~w9480;
assign w9543 = ~w9406 & ~w9409;
assign w9544 = ~w9471 & ~w9474;
assign w9545 = ~w9360 & ~w9363;
assign w9546 = ~w9362 & ~w9545;
assign w9547 = w9225 & ~w9396;
assign w9548 = ~w9398 & ~w9547;
assign w9549 = w9546 & ~w9548;
assign w9550 = ~w9546 & w9548;
assign w9551 = ~w9549 & ~w9550;
assign w9552 = ~w9314 & ~w9318;
assign w9553 = ~w9317 & ~w9552;
assign w9554 = ~w9551 & ~w9553;
assign w9555 = w9551 & w9553;
assign w9556 = ~w9554 & ~w9555;
assign w9557 = (~w9463 & ~w9465) | (~w9463 & w16763) | (~w9465 & w16763);
assign w9558 = (~w9430 & ~w9432) | (~w9430 & w16764) | (~w9432 & w16764);
assign w9559 = ~w9557 & ~w9558;
assign w9560 = w9557 & w9558;
assign w9561 = ~w9559 & ~w9560;
assign w9562 = w9556 & w9561;
assign w9563 = ~w9556 & ~w9561;
assign w9564 = ~w9562 & ~w9563;
assign w9565 = ~w9544 & w9564;
assign w9566 = w9544 & ~w9564;
assign w9567 = ~w9565 & ~w9566;
assign w9568 = ~w9543 & w9567;
assign w9569 = w9543 & ~w9567;
assign w9570 = ~w9568 & ~w9569;
assign w9571 = ~w9542 & w9570;
assign w9572 = w9542 & ~w9570;
assign w9573 = ~w9571 & ~w9572;
assign w9574 = ~w9299 & ~w9303;
assign w9575 = (~w9507 & ~w9509) | (~w9507 & w17163) | (~w9509 & w17163);
assign w9576 = (~w9357 & ~w9359) | (~w9357 & w16924) | (~w9359 & w16924);
assign w9577 = (~w9391 & ~w9393) | (~w9391 & w16925) | (~w9393 & w16925);
assign w9578 = ~w9576 & ~w9577;
assign w9579 = w9576 & w9577;
assign w9580 = ~w9578 & ~w9579;
assign w9581 = w9575 & ~w9580;
assign w9582 = ~w9575 & w9580;
assign w9583 = ~w9581 & ~w9582;
assign w9584 = w9216 & ~w9307;
assign w9585 = ~w9309 & ~w9584;
assign w9586 = w9326 & ~w9329;
assign w9587 = ~w9331 & ~w9586;
assign w9588 = ~w9585 & ~w9587;
assign w9589 = w9585 & w9587;
assign w9590 = ~w9588 & ~w9589;
assign w9591 = w9381 & ~w9384;
assign w9592 = ~w9386 & ~w9591;
assign w9593 = ~w9590 & w9592;
assign w9594 = w9590 & ~w9592;
assign w9595 = ~w9593 & ~w9594;
assign w9596 = ~w9348 & ~w9352;
assign w9597 = ~w9351 & ~w9596;
assign w9598 = w9192 & ~w9341;
assign w9599 = ~w9343 & ~w9598;
assign w9600 = w9597 & ~w9599;
assign w9601 = ~w9597 & w9599;
assign w9602 = ~w9600 & ~w9601;
assign w9603 = w9371 & ~w9374;
assign w9604 = ~w9376 & ~w9603;
assign w9605 = ~w9602 & w9604;
assign w9606 = w9602 & ~w9604;
assign w9607 = ~w9605 & ~w9606;
assign w9608 = (~w9323 & ~w9325) | (~w9323 & w16926) | (~w9325 & w16926);
assign w9609 = ~w9607 & w9608;
assign w9610 = w9607 & ~w9608;
assign w9611 = ~w9609 & ~w9610;
assign w9612 = w9595 & w9611;
assign w9613 = ~w9595 & ~w9611;
assign w9614 = ~w9612 & ~w9613;
assign w9615 = w9583 & w9614;
assign w9616 = ~w9583 & ~w9614;
assign w9617 = ~w9615 & ~w9616;
assign w9618 = w9574 & ~w9617;
assign w9619 = ~w9574 & w9617;
assign w9620 = ~w9618 & ~w9619;
assign w9621 = w9573 & w9620;
assign w9622 = ~w9573 & ~w9620;
assign w9623 = ~w9621 & ~w9622;
assign w9624 = ~w9541 & w9623;
assign w9625 = w9541 & ~w9623;
assign w9626 = ~w9624 & ~w9625;
assign w9627 = (~w9488 & ~w9490) | (~w9488 & w16927) | (~w9490 & w16927);
assign w9628 = pi09 & pi60;
assign w9629 = pi10 & pi59;
assign w9630 = ~w9628 & ~w9629;
assign w9631 = pi10 & pi60;
assign w9632 = w9216 & w9631;
assign w9633 = ~w9630 & ~w9632;
assign w9634 = w9499 & ~w9633;
assign w9635 = ~w9499 & w9633;
assign w9636 = ~w9634 & ~w9635;
assign w9637 = pi24 & pi45;
assign w9638 = pi25 & pi44;
assign w9639 = ~w9637 & ~w9638;
assign w9640 = pi25 & pi45;
assign w9641 = w9225 & w9640;
assign w9642 = ~w9639 & ~w9641;
assign w9643 = w9385 & ~w9642;
assign w9644 = ~w9385 & w9642;
assign w9645 = ~w9643 & ~w9644;
assign w9646 = ~w9636 & ~w9645;
assign w9647 = w9636 & w9645;
assign w9648 = ~w9646 & ~w9647;
assign w9649 = pi27 & pi42;
assign w9650 = ~w9397 & ~w9649;
assign w9651 = pi27 & pi43;
assign w9652 = w9395 & w9651;
assign w9653 = ~w9650 & ~w9652;
assign w9654 = w9330 & ~w9653;
assign w9655 = ~w9330 & w9653;
assign w9656 = ~w9654 & ~w9655;
assign w9657 = w9648 & ~w9656;
assign w9658 = ~w9648 & w9656;
assign w9659 = ~w9657 & ~w9658;
assign w9660 = ~w9627 & w9659;
assign w9661 = w9627 & ~w9659;
assign w9662 = ~w9660 & ~w9661;
assign w9663 = (~w9500 & w9503) | (~w9500 & w16765) | (w9503 & w16765);
assign w9664 = pi13 & pi56;
assign w9665 = pi12 & pi57;
assign w9666 = ~w9664 & ~w9665;
assign w9667 = pi13 & pi57;
assign w9668 = w9360 & w9667;
assign w9669 = ~w9666 & ~w9668;
assign w9670 = w9308 & ~w9669;
assign w9671 = ~w9308 & w9669;
assign w9672 = ~w9670 & ~w9671;
assign w9673 = ~w9663 & ~w9672;
assign w9674 = w9663 & w9672;
assign w9675 = ~w9673 & ~w9674;
assign w9676 = pi14 & pi55;
assign w9677 = pi21 & pi48;
assign w9678 = pi22 & pi47;
assign w9679 = ~w9677 & ~w9678;
assign w9680 = pi22 & pi48;
assign w9681 = w9326 & w9680;
assign w9682 = ~w9679 & ~w9681;
assign w9683 = w9676 & ~w9682;
assign w9684 = ~w9676 & w9682;
assign w9685 = ~w9683 & ~w9684;
assign w9686 = w9675 & ~w9685;
assign w9687 = ~w9675 & w9685;
assign w9688 = ~w9686 & ~w9687;
assign w9689 = w9662 & w9688;
assign w9690 = ~w9662 & ~w9688;
assign w9691 = ~w9689 & ~w9690;
assign w9692 = ~w9513 & ~w9516;
assign w9693 = (~w9440 & ~w9442) | (~w9440 & w17806) | (~w9442 & w17806);
assign w9694 = (~w9451 & ~w9453) | (~w9451 & w17164) | (~w9453 & w17164);
assign w9695 = pi18 & pi51;
assign w9696 = pi17 & pi52;
assign w9697 = ~w9695 & ~w9696;
assign w9698 = pi18 & pi52;
assign w9699 = w9361 & w9698;
assign w9700 = ~w9697 & ~w9699;
assign w9701 = w9342 & ~w9700;
assign w9702 = ~w9342 & w9700;
assign w9703 = ~w9701 & ~w9702;
assign w9704 = pi28 & pi41;
assign w9705 = pi29 & pi40;
assign w9706 = pi30 & pi39;
assign w9707 = ~w9705 & ~w9706;
assign w9708 = w9705 & w9706;
assign w9709 = ~w9707 & ~w9708;
assign w9710 = w9704 & ~w9709;
assign w9711 = ~w9704 & w9709;
assign w9712 = ~w9710 & ~w9711;
assign w9713 = ~w9703 & ~w9712;
assign w9714 = w9703 & w9712;
assign w9715 = ~w9713 & ~w9714;
assign w9716 = w9694 & ~w9715;
assign w9717 = ~w9694 & w9715;
assign w9718 = ~w9716 & ~w9717;
assign w9719 = pi07 & pi62;
assign w9720 = ~pi34 & pi35;
assign w9721 = w9719 & ~w9720;
assign w9722 = ~w9719 & w9720;
assign w9723 = ~w9721 & ~w9722;
assign w9724 = pi31 & pi38;
assign w9725 = pi32 & pi37;
assign w9726 = pi33 & pi36;
assign w9727 = ~w9725 & ~w9726;
assign w9728 = w9725 & w9726;
assign w9729 = ~w9727 & ~w9728;
assign w9730 = w9724 & ~w9729;
assign w9731 = ~w9724 & w9729;
assign w9732 = ~w9730 & ~w9731;
assign w9733 = ~w9723 & ~w9732;
assign w9734 = w9723 & w9732;
assign w9735 = ~w9733 & ~w9734;
assign w9736 = pi15 & pi54;
assign w9737 = pi20 & pi49;
assign w9738 = ~w9375 & ~w9737;
assign w9739 = w9375 & w9737;
assign w9740 = ~w9738 & ~w9739;
assign w9741 = w9736 & ~w9740;
assign w9742 = ~w9736 & w9740;
assign w9743 = ~w9741 & ~w9742;
assign w9744 = w9735 & ~w9743;
assign w9745 = ~w9735 & w9743;
assign w9746 = ~w9744 & ~w9745;
assign w9747 = ~w9718 & ~w9746;
assign w9748 = w9718 & w9746;
assign w9749 = ~w9747 & ~w9748;
assign w9750 = w9693 & w9749;
assign w9751 = ~w9693 & ~w9749;
assign w9752 = ~w9750 & ~w9751;
assign w9753 = ~w9692 & ~w9752;
assign w9754 = w9692 & w9752;
assign w9755 = ~w9753 & ~w9754;
assign w9756 = w9691 & w9755;
assign w9757 = ~w9691 & ~w9755;
assign w9758 = ~w9756 & ~w9757;
assign w9759 = (~w9519 & ~w9521) | (~w9519 & w17807) | (~w9521 & w17807);
assign w9760 = ~w9412 & ~w9415;
assign w9761 = ~w9759 & ~w9760;
assign w9762 = w9759 & w9760;
assign w9763 = ~w9761 & ~w9762;
assign w9764 = w9758 & w9763;
assign w9765 = ~w9758 & ~w9763;
assign w9766 = ~w9764 & ~w9765;
assign w9767 = w9626 & w9766;
assign w9768 = ~w9626 & ~w9766;
assign w9769 = ~w9767 & ~w9768;
assign w9770 = ~w9540 & w9769;
assign w9771 = w9540 & ~w9769;
assign w9772 = ~w9770 & ~w9771;
assign w9773 = ~w9286 & ~w9533;
assign w9774 = (w8795 & w16560) | (w8795 & w16561) | (w16560 & w16561);
assign w9775 = w9772 & w9774;
assign w9776 = ~w9772 & ~w9774;
assign w9777 = ~w9775 & ~w9776;
assign w9778 = ~w9624 & ~w9767;
assign w9779 = (~w9571 & ~w9573) | (~w9571 & w17808) | (~w9573 & w17808);
assign w9780 = ~w9704 & ~w9708;
assign w9781 = ~w9707 & ~w9780;
assign w9782 = w9330 & ~w9650;
assign w9783 = ~w9652 & ~w9782;
assign w9784 = w9781 & ~w9783;
assign w9785 = ~w9781 & w9783;
assign w9786 = ~w9784 & ~w9785;
assign w9787 = w9385 & ~w9639;
assign w9788 = ~w9641 & ~w9787;
assign w9789 = ~w9786 & w9788;
assign w9790 = w9786 & ~w9788;
assign w9791 = ~w9789 & ~w9790;
assign w9792 = pi08 & pi62;
assign w9793 = ~pi34 & ~w9719;
assign w9794 = pi35 & ~w9793;
assign w9795 = w9792 & w9794;
assign w9796 = ~w9792 & ~w9794;
assign w9797 = ~w9795 & ~w9796;
assign w9798 = ~w9724 & ~w9728;
assign w9799 = ~w9727 & ~w9798;
assign w9800 = ~w9797 & w9799;
assign w9801 = w9797 & ~w9799;
assign w9802 = ~w9800 & ~w9801;
assign w9803 = ~w9791 & w9802;
assign w9804 = w9791 & ~w9802;
assign w9805 = ~w9803 & ~w9804;
assign w9806 = ~w9713 & ~w9717;
assign w9807 = ~w9805 & w9806;
assign w9808 = w9805 & ~w9806;
assign w9809 = ~w9807 & ~w9808;
assign w9810 = (~w9733 & ~w9735) | (~w9733 & w17452) | (~w9735 & w17452);
assign w9811 = (~w9646 & ~w9648) | (~w9646 & w16928) | (~w9648 & w16928);
assign w9812 = (~w9673 & ~w9675) | (~w9673 & w16929) | (~w9675 & w16929);
assign w9813 = ~w9811 & ~w9812;
assign w9814 = w9811 & w9812;
assign w9815 = ~w9813 & ~w9814;
assign w9816 = w9810 & ~w9815;
assign w9817 = ~w9810 & w9815;
assign w9818 = ~w9816 & ~w9817;
assign w9819 = ~w9747 & ~w9750;
assign w9820 = w9818 & w9819;
assign w9821 = ~w9818 & ~w9819;
assign w9822 = ~w9820 & ~w9821;
assign w9823 = ~w9809 & ~w9822;
assign w9824 = w9809 & w9822;
assign w9825 = ~w9823 & ~w9824;
assign w9826 = ~w9779 & w9825;
assign w9827 = w9779 & ~w9825;
assign w9828 = ~w9826 & ~w9827;
assign w9829 = (~w9565 & ~w9567) | (~w9565 & w17809) | (~w9567 & w17809);
assign w9830 = pi09 & pi61;
assign w9831 = pi11 & pi59;
assign w9832 = ~w9631 & ~w9831;
assign w9833 = pi11 & pi60;
assign w9834 = w9629 & w9833;
assign w9835 = ~w9832 & ~w9834;
assign w9836 = w9830 & ~w9835;
assign w9837 = ~w9830 & w9835;
assign w9838 = ~w9836 & ~w9837;
assign w9839 = pi17 & pi53;
assign w9840 = pi16 & pi54;
assign w9841 = ~w9839 & ~w9840;
assign w9842 = pi17 & pi54;
assign w9843 = w9375 & w9842;
assign w9844 = ~w9841 & ~w9843;
assign w9845 = w9698 & ~w9844;
assign w9846 = ~w9698 & w9844;
assign w9847 = ~w9845 & ~w9846;
assign w9848 = ~w9838 & ~w9847;
assign w9849 = w9838 & w9847;
assign w9850 = ~w9848 & ~w9849;
assign w9851 = pi12 & pi58;
assign w9852 = pi24 & pi46;
assign w9853 = ~w9667 & ~w9852;
assign w9854 = w9667 & w9852;
assign w9855 = ~w9853 & ~w9854;
assign w9856 = w9851 & ~w9855;
assign w9857 = ~w9851 & w9855;
assign w9858 = ~w9856 & ~w9857;
assign w9859 = w9850 & ~w9858;
assign w9860 = ~w9850 & w9858;
assign w9861 = ~w9859 & ~w9860;
assign w9862 = ~w9736 & ~w9739;
assign w9863 = ~w9738 & ~w9862;
assign w9864 = w9342 & ~w9697;
assign w9865 = ~w9699 & ~w9864;
assign w9866 = w9863 & ~w9865;
assign w9867 = ~w9863 & w9865;
assign w9868 = ~w9866 & ~w9867;
assign w9869 = pi32 & pi38;
assign w9870 = pi33 & pi37;
assign w9871 = pi34 & pi36;
assign w9872 = ~w9870 & ~w9871;
assign w9873 = w9870 & w9871;
assign w9874 = ~w9872 & ~w9873;
assign w9875 = w9869 & ~w9874;
assign w9876 = ~w9869 & w9874;
assign w9877 = ~w9875 & ~w9876;
assign w9878 = ~w9868 & w9877;
assign w9879 = w9868 & ~w9877;
assign w9880 = ~w9878 & ~w9879;
assign w9881 = (~w9559 & ~w9561) | (~w9559 & w16930) | (~w9561 & w16930);
assign w9882 = w9880 & ~w9881;
assign w9883 = ~w9880 & w9881;
assign w9884 = ~w9882 & ~w9883;
assign w9885 = w9861 & w9884;
assign w9886 = ~w9861 & ~w9884;
assign w9887 = ~w9885 & ~w9886;
assign w9888 = ~w9829 & w9887;
assign w9889 = w9829 & ~w9887;
assign w9890 = ~w9888 & ~w9889;
assign w9891 = (~w9610 & ~w9611) | (~w9610 & w17165) | (~w9611 & w17165);
assign w9892 = (~w9600 & ~w9602) | (~w9600 & w17166) | (~w9602 & w17166);
assign w9893 = pi28 & pi42;
assign w9894 = pi23 & pi47;
assign w9895 = pi07 & pi63;
assign w9896 = ~w9894 & ~w9895;
assign w9897 = w9894 & w9895;
assign w9898 = ~w9896 & ~w9897;
assign w9899 = w9893 & ~w9898;
assign w9900 = ~w9893 & w9898;
assign w9901 = ~w9899 & ~w9900;
assign w9902 = pi29 & pi41;
assign w9903 = pi30 & pi40;
assign w9904 = pi31 & pi39;
assign w9905 = ~w9903 & ~w9904;
assign w9906 = w9903 & w9904;
assign w9907 = ~w9905 & ~w9906;
assign w9908 = w9902 & ~w9907;
assign w9909 = ~w9902 & w9907;
assign w9910 = ~w9908 & ~w9909;
assign w9911 = ~w9901 & ~w9910;
assign w9912 = w9901 & w9910;
assign w9913 = ~w9911 & ~w9912;
assign w9914 = w9892 & ~w9913;
assign w9915 = ~w9892 & w9913;
assign w9916 = ~w9914 & ~w9915;
assign w9917 = pi14 & pi56;
assign w9918 = pi15 & pi55;
assign w9919 = ~w9917 & ~w9918;
assign w9920 = pi15 & pi56;
assign w9921 = w9676 & w9920;
assign w9922 = ~w9919 & ~w9921;
assign w9923 = w9680 & ~w9922;
assign w9924 = ~w9680 & w9922;
assign w9925 = ~w9923 & ~w9924;
assign w9926 = pi26 & pi44;
assign w9927 = ~w9651 & ~w9926;
assign w9928 = pi27 & pi44;
assign w9929 = w9397 & w9928;
assign w9930 = ~w9927 & ~w9929;
assign w9931 = w9640 & ~w9930;
assign w9932 = ~w9640 & w9930;
assign w9933 = ~w9931 & ~w9932;
assign w9934 = ~w9925 & ~w9933;
assign w9935 = w9925 & w9933;
assign w9936 = ~w9934 & ~w9935;
assign w9937 = pi21 & pi49;
assign w9938 = pi19 & pi51;
assign w9939 = pi20 & pi50;
assign w9940 = ~w9938 & ~w9939;
assign w9941 = pi20 & pi51;
assign w9942 = w9342 & w9941;
assign w9943 = ~w9940 & ~w9942;
assign w9944 = w9937 & ~w9943;
assign w9945 = ~w9937 & w9943;
assign w9946 = ~w9944 & ~w9945;
assign w9947 = w9936 & ~w9946;
assign w9948 = ~w9936 & w9946;
assign w9949 = ~w9947 & ~w9948;
assign w9950 = ~w9916 & ~w9949;
assign w9951 = w9916 & w9949;
assign w9952 = ~w9950 & ~w9951;
assign w9953 = w9891 & w9952;
assign w9954 = ~w9891 & ~w9952;
assign w9955 = ~w9953 & ~w9954;
assign w9956 = w9890 & ~w9955;
assign w9957 = ~w9890 & w9955;
assign w9958 = ~w9956 & ~w9957;
assign w9959 = w9828 & w9958;
assign w9960 = ~w9828 & ~w9958;
assign w9961 = ~w9959 & ~w9960;
assign w9962 = ~w9753 & ~w9756;
assign w9963 = ~w9615 & ~w9619;
assign w9964 = (~w9660 & ~w9662) | (~w9660 & w17167) | (~w9662 & w17167);
assign w9965 = (~w9578 & ~w9580) | (~w9578 & w17168) | (~w9580 & w17168);
assign w9966 = w9499 & ~w9630;
assign w9967 = ~w9632 & ~w9966;
assign w9968 = w9308 & ~w9666;
assign w9969 = ~w9668 & ~w9968;
assign w9970 = ~w9967 & ~w9969;
assign w9971 = w9967 & w9969;
assign w9972 = ~w9970 & ~w9971;
assign w9973 = w9676 & ~w9679;
assign w9974 = ~w9681 & ~w9973;
assign w9975 = ~w9972 & w9974;
assign w9976 = w9972 & ~w9974;
assign w9977 = ~w9975 & ~w9976;
assign w9978 = (~w9588 & ~w9590) | (~w9588 & w16766) | (~w9590 & w16766);
assign w9979 = (~w9549 & ~w9551) | (~w9549 & w16767) | (~w9551 & w16767);
assign w9980 = ~w9978 & ~w9979;
assign w9981 = w9978 & w9979;
assign w9982 = ~w9980 & ~w9981;
assign w9983 = w9977 & w9982;
assign w9984 = ~w9977 & ~w9982;
assign w9985 = ~w9983 & ~w9984;
assign w9986 = ~w9965 & w9985;
assign w9987 = w9965 & ~w9985;
assign w9988 = ~w9986 & ~w9987;
assign w9989 = ~w9964 & w9988;
assign w9990 = w9964 & ~w9988;
assign w9991 = ~w9989 & ~w9990;
assign w9992 = ~w9963 & w9991;
assign w9993 = w9963 & ~w9991;
assign w9994 = ~w9992 & ~w9993;
assign w9995 = w9962 & ~w9994;
assign w9996 = ~w9962 & w9994;
assign w9997 = ~w9995 & ~w9996;
assign w9998 = ~w9761 & ~w9764;
assign w9999 = w9997 & ~w9998;
assign w10000 = ~w9997 & w9998;
assign w10001 = ~w9999 & ~w10000;
assign w10002 = w9961 & w10001;
assign w10003 = ~w9961 & ~w10001;
assign w10004 = ~w10002 & ~w10003;
assign w10005 = ~w9778 & w10004;
assign w10006 = w9778 & ~w10004;
assign w10007 = ~w10005 & ~w10006;
assign w10008 = (~w7754 & w17605) | (~w7754 & w17606) | (w17605 & w17606);
assign w10009 = (w7754 & w17810) | (w7754 & w17811) | (w17810 & w17811);
assign w10010 = w10007 & w10009;
assign w10011 = ~w10007 & ~w10009;
assign w10012 = ~w10010 & ~w10011;
assign w10013 = ~w9771 & ~w10006;
assign w10014 = (~w7754 & w17812) | (~w7754 & w17813) | (w17812 & w17813);
assign w10015 = ~w9999 & ~w10002;
assign w10016 = ~w9888 & ~w9956;
assign w10017 = (~w9784 & ~w9786) | (~w9784 & w17169) | (~w9786 & w17169);
assign w10018 = (~w9866 & ~w9868) | (~w9866 & w16768) | (~w9868 & w16768);
assign w10019 = ~w9795 & ~w9799;
assign w10020 = ~w9796 & ~w10019;
assign w10021 = ~w10018 & w10020;
assign w10022 = w10018 & ~w10020;
assign w10023 = ~w10021 & ~w10022;
assign w10024 = w10017 & ~w10023;
assign w10025 = ~w10017 & w10023;
assign w10026 = ~w10024 & ~w10025;
assign w10027 = (~w9804 & ~w9805) | (~w9804 & w17170) | (~w9805 & w17170);
assign w10028 = ~w10026 & w10027;
assign w10029 = w10026 & ~w10027;
assign w10030 = ~w10028 & ~w10029;
assign w10031 = (~w9882 & ~w9884) | (~w9882 & w17171) | (~w9884 & w17171);
assign w10032 = ~w10030 & w10031;
assign w10033 = w10030 & ~w10031;
assign w10034 = ~w10032 & ~w10033;
assign w10035 = ~w9820 & ~w9824;
assign w10036 = ~w10034 & w10035;
assign w10037 = w10034 & ~w10035;
assign w10038 = ~w10036 & ~w10037;
assign w10039 = w10016 & ~w10038;
assign w10040 = ~w10016 & w10038;
assign w10041 = ~w10039 & ~w10040;
assign w10042 = ~w9826 & ~w9959;
assign w10043 = ~w10041 & w10042;
assign w10044 = w10041 & ~w10042;
assign w10045 = ~w10043 & ~w10044;
assign w10046 = ~w9992 & ~w9996;
assign w10047 = (~w9934 & ~w9936) | (~w9934 & w17455) | (~w9936 & w17455);
assign w10048 = (~w9848 & ~w9850) | (~w9848 & w16931) | (~w9850 & w16931);
assign w10049 = (~w9970 & ~w9972) | (~w9970 & w17172) | (~w9972 & w17172);
assign w10050 = ~w10048 & ~w10049;
assign w10051 = w10048 & w10049;
assign w10052 = ~w10050 & ~w10051;
assign w10053 = w10047 & ~w10052;
assign w10054 = ~w10047 & w10052;
assign w10055 = ~w10053 & ~w10054;
assign w10056 = ~w9950 & ~w9953;
assign w10057 = w10055 & w10056;
assign w10058 = ~w10055 & ~w10056;
assign w10059 = ~w10057 & ~w10058;
assign w10060 = ~w9911 & ~w9915;
assign w10061 = ~w9851 & ~w9854;
assign w10062 = ~w9853 & ~w10061;
assign w10063 = w9830 & ~w9832;
assign w10064 = ~w9834 & ~w10063;
assign w10065 = w10062 & ~w10064;
assign w10066 = ~w10062 & w10064;
assign w10067 = ~w10065 & ~w10066;
assign w10068 = w9640 & ~w9927;
assign w10069 = ~w9929 & ~w10068;
assign w10070 = ~w10067 & w10069;
assign w10071 = w10067 & ~w10069;
assign w10072 = ~w10070 & ~w10071;
assign w10073 = ~w9902 & ~w9906;
assign w10074 = ~w9905 & ~w10073;
assign w10075 = w9680 & ~w9919;
assign w10076 = ~w9921 & ~w10075;
assign w10077 = w10074 & ~w10076;
assign w10078 = ~w10074 & w10076;
assign w10079 = ~w10077 & ~w10078;
assign w10080 = ~w9893 & ~w9897;
assign w10081 = ~w9896 & ~w10080;
assign w10082 = ~w10079 & ~w10081;
assign w10083 = w10079 & w10081;
assign w10084 = ~w10082 & ~w10083;
assign w10085 = w10072 & w10084;
assign w10086 = ~w10072 & ~w10084;
assign w10087 = ~w10085 & ~w10086;
assign w10088 = ~w10060 & w10087;
assign w10089 = w10060 & ~w10087;
assign w10090 = ~w10088 & ~w10089;
assign w10091 = w10059 & w10090;
assign w10092 = ~w10059 & ~w10090;
assign w10093 = ~w10091 & ~w10092;
assign w10094 = ~w10046 & w10093;
assign w10095 = w10046 & ~w10093;
assign w10096 = ~w10094 & ~w10095;
assign w10097 = ~w9986 & ~w9989;
assign w10098 = pi22 & pi49;
assign w10099 = pi62 & w4081;
assign w10100 = pi09 & pi62;
assign w10101 = ~pi36 & ~w10100;
assign w10102 = ~w10099 & ~w10101;
assign w10103 = w10098 & ~w10102;
assign w10104 = ~w10098 & w10102;
assign w10105 = ~w10103 & ~w10104;
assign w10106 = pi21 & pi50;
assign w10107 = pi19 & pi52;
assign w10108 = ~w9941 & ~w10107;
assign w10109 = pi20 & pi52;
assign w10110 = w9938 & w10109;
assign w10111 = ~w10108 & ~w10110;
assign w10112 = w10106 & ~w10111;
assign w10113 = ~w10106 & w10111;
assign w10114 = ~w10112 & ~w10113;
assign w10115 = ~w10105 & ~w10114;
assign w10116 = w10105 & w10114;
assign w10117 = ~w10115 & ~w10116;
assign w10118 = pi33 & pi38;
assign w10119 = pi34 & pi37;
assign w10120 = pi35 & pi36;
assign w10121 = ~w10119 & ~w10120;
assign w10122 = w10119 & w10120;
assign w10123 = ~w10121 & ~w10122;
assign w10124 = w10118 & ~w10123;
assign w10125 = ~w10118 & w10123;
assign w10126 = ~w10124 & ~w10125;
assign w10127 = w10117 & ~w10126;
assign w10128 = ~w10117 & w10126;
assign w10129 = ~w10127 & ~w10128;
assign w10130 = ~w9869 & ~w9873;
assign w10131 = ~w9872 & ~w10130;
assign w10132 = w9698 & ~w9841;
assign w10133 = ~w9843 & ~w10132;
assign w10134 = w10131 & ~w10133;
assign w10135 = ~w10131 & w10133;
assign w10136 = ~w10134 & ~w10135;
assign w10137 = pi08 & pi63;
assign w10138 = pi10 & pi61;
assign w10139 = ~w10137 & ~w10138;
assign w10140 = w10137 & w10138;
assign w10141 = ~w10139 & ~w10140;
assign w10142 = w9833 & ~w10141;
assign w10143 = ~w9833 & w10141;
assign w10144 = ~w10142 & ~w10143;
assign w10145 = ~w10136 & w10144;
assign w10146 = w10136 & ~w10144;
assign w10147 = ~w10145 & ~w10146;
assign w10148 = (~w9980 & ~w9982) | (~w9980 & w16932) | (~w9982 & w16932);
assign w10149 = w10147 & ~w10148;
assign w10150 = ~w10147 & w10148;
assign w10151 = ~w10149 & ~w10150;
assign w10152 = w10129 & w10151;
assign w10153 = ~w10129 & ~w10151;
assign w10154 = ~w10152 & ~w10153;
assign w10155 = ~w10097 & w10154;
assign w10156 = w10097 & ~w10154;
assign w10157 = ~w10155 & ~w10156;
assign w10158 = (~w9813 & ~w9815) | (~w9813 & w17173) | (~w9815 & w17173);
assign w10159 = pi28 & pi43;
assign w10160 = pi29 & pi42;
assign w10161 = ~w10159 & ~w10160;
assign w10162 = pi29 & pi43;
assign w10163 = w9893 & w10162;
assign w10164 = ~w10161 & ~w10163;
assign w10165 = w9928 & ~w10164;
assign w10166 = ~w9928 & w10164;
assign w10167 = ~w10165 & ~w10166;
assign w10168 = pi30 & pi41;
assign w10169 = pi31 & pi40;
assign w10170 = pi32 & pi39;
assign w10171 = ~w10169 & ~w10170;
assign w10172 = w10169 & w10170;
assign w10173 = ~w10171 & ~w10172;
assign w10174 = w10168 & ~w10173;
assign w10175 = ~w10168 & w10173;
assign w10176 = ~w10174 & ~w10175;
assign w10177 = ~w10167 & ~w10176;
assign w10178 = w10167 & w10176;
assign w10179 = ~w10177 & ~w10178;
assign w10180 = pi23 & pi48;
assign w10181 = pi18 & pi53;
assign w10182 = ~w9842 & ~w10181;
assign w10183 = pi18 & pi54;
assign w10184 = w9839 & w10183;
assign w10185 = ~w10182 & ~w10184;
assign w10186 = w10180 & ~w10185;
assign w10187 = ~w10180 & w10185;
assign w10188 = ~w10186 & ~w10187;
assign w10189 = w10179 & ~w10188;
assign w10190 = ~w10179 & w10188;
assign w10191 = ~w10189 & ~w10190;
assign w10192 = pi13 & pi58;
assign w10193 = pi12 & pi59;
assign w10194 = ~w10192 & ~w10193;
assign w10195 = pi13 & pi59;
assign w10196 = w9851 & w10195;
assign w10197 = ~w10194 & ~w10196;
assign w10198 = w9937 & ~w9940;
assign w10199 = ~w9942 & ~w10198;
assign w10200 = w10197 & ~w10199;
assign w10201 = ~w10197 & w10199;
assign w10202 = ~w10200 & ~w10201;
assign w10203 = pi14 & pi57;
assign w10204 = pi16 & pi55;
assign w10205 = ~w9920 & ~w10204;
assign w10206 = pi16 & pi56;
assign w10207 = w9918 & w10206;
assign w10208 = ~w10205 & ~w10207;
assign w10209 = w10203 & ~w10208;
assign w10210 = ~w10203 & w10208;
assign w10211 = ~w10209 & ~w10210;
assign w10212 = pi24 & pi47;
assign w10213 = pi25 & pi46;
assign w10214 = pi26 & pi45;
assign w10215 = ~w10213 & ~w10214;
assign w10216 = pi26 & pi46;
assign w10217 = w9640 & w10216;
assign w10218 = ~w10215 & ~w10217;
assign w10219 = w10212 & ~w10218;
assign w10220 = ~w10212 & w10218;
assign w10221 = ~w10219 & ~w10220;
assign w10222 = ~w10211 & ~w10221;
assign w10223 = w10211 & w10221;
assign w10224 = ~w10222 & ~w10223;
assign w10225 = w10202 & w10224;
assign w10226 = ~w10202 & ~w10224;
assign w10227 = ~w10225 & ~w10226;
assign w10228 = w10191 & w10227;
assign w10229 = ~w10191 & ~w10227;
assign w10230 = ~w10228 & ~w10229;
assign w10231 = ~w10158 & w10230;
assign w10232 = w10158 & ~w10230;
assign w10233 = ~w10231 & ~w10232;
assign w10234 = w10157 & w10233;
assign w10235 = ~w10157 & ~w10233;
assign w10236 = ~w10234 & ~w10235;
assign w10237 = w10096 & w10236;
assign w10238 = ~w10096 & ~w10236;
assign w10239 = ~w10237 & ~w10238;
assign w10240 = ~w10045 & ~w10239;
assign w10241 = w10045 & w10239;
assign w10242 = ~w10240 & ~w10241;
assign w10243 = w10015 & ~w10242;
assign w10244 = ~w10015 & w10242;
assign w10245 = ~w10243 & ~w10244;
assign w10246 = w10014 & w10245;
assign w10247 = ~w10014 & ~w10245;
assign w10248 = ~w10246 & ~w10247;
assign w10249 = ~w10005 & ~w10244;
assign w10250 = (w7754 & w17814) | (w7754 & w17815) | (w17814 & w17815);
assign w10251 = (~w10155 & ~w10157) | (~w10155 & w17456) | (~w10157 & w17456);
assign w10252 = (~w10085 & ~w10087) | (~w10085 & w17174) | (~w10087 & w17174);
assign w10253 = (~w10077 & ~w10079) | (~w10077 & w17175) | (~w10079 & w17175);
assign w10254 = (~w10134 & ~w10136) | (~w10134 & w16769) | (~w10136 & w16769);
assign w10255 = pi31 & pi41;
assign w10256 = pi30 & pi42;
assign w10257 = ~w10255 & ~w10256;
assign w10258 = pi31 & pi42;
assign w10259 = w10168 & w10258;
assign w10260 = ~w10257 & ~w10259;
assign w10261 = w10162 & ~w10260;
assign w10262 = ~w10162 & w10260;
assign w10263 = ~w10261 & ~w10262;
assign w10264 = ~w10254 & ~w10263;
assign w10265 = w10254 & w10263;
assign w10266 = ~w10264 & ~w10265;
assign w10267 = w10253 & ~w10266;
assign w10268 = ~w10253 & w10266;
assign w10269 = ~w10267 & ~w10268;
assign w10270 = ~w10252 & w10269;
assign w10271 = w10252 & ~w10269;
assign w10272 = ~w10270 & ~w10271;
assign w10273 = (~w10149 & ~w10151) | (~w10149 & w17176) | (~w10151 & w17176);
assign w10274 = ~w10272 & w10273;
assign w10275 = w10272 & ~w10273;
assign w10276 = ~w10274 & ~w10275;
assign w10277 = (~w10057 & ~w10059) | (~w10057 & w17457) | (~w10059 & w17457);
assign w10278 = ~w10276 & w10277;
assign w10279 = w10276 & ~w10277;
assign w10280 = ~w10278 & ~w10279;
assign w10281 = w10251 & ~w10280;
assign w10282 = ~w10251 & w10280;
assign w10283 = ~w10281 & ~w10282;
assign w10284 = ~w10094 & ~w10237;
assign w10285 = ~w10283 & w10284;
assign w10286 = w10283 & ~w10284;
assign w10287 = ~w10285 & ~w10286;
assign w10288 = ~w10037 & ~w10040;
assign w10289 = (~w10115 & ~w10117) | (~w10115 & w17458) | (~w10117 & w17458);
assign w10290 = (~w10177 & ~w10179) | (~w10177 & w16933) | (~w10179 & w16933);
assign w10291 = (~w10065 & ~w10067) | (~w10065 & w17177) | (~w10067 & w17177);
assign w10292 = ~w10290 & ~w10291;
assign w10293 = w10290 & w10291;
assign w10294 = ~w10292 & ~w10293;
assign w10295 = w10289 & ~w10294;
assign w10296 = ~w10289 & w10294;
assign w10297 = ~w10295 & ~w10296;
assign w10298 = ~w10228 & ~w10231;
assign w10299 = ~w10297 & w10298;
assign w10300 = w10297 & ~w10298;
assign w10301 = ~w10299 & ~w10300;
assign w10302 = (~w10222 & ~w10224) | (~w10222 & w17459) | (~w10224 & w17459);
assign w10303 = w9928 & ~w10161;
assign w10304 = ~w10163 & ~w10303;
assign w10305 = w10180 & ~w10182;
assign w10306 = ~w10184 & ~w10305;
assign w10307 = ~w10304 & ~w10306;
assign w10308 = w10304 & w10306;
assign w10309 = ~w10307 & ~w10308;
assign w10310 = ~w10168 & ~w10172;
assign w10311 = ~w10171 & ~w10310;
assign w10312 = ~w10309 & ~w10311;
assign w10313 = w10309 & w10311;
assign w10314 = ~w10312 & ~w10313;
assign w10315 = w10098 & ~w10101;
assign w10316 = ~w10099 & ~w10315;
assign w10317 = ~w10118 & ~w10122;
assign w10318 = ~w10121 & ~w10317;
assign w10319 = ~w10316 & w10318;
assign w10320 = w10316 & ~w10318;
assign w10321 = ~w10319 & ~w10320;
assign w10322 = w10106 & ~w10108;
assign w10323 = ~w10110 & ~w10322;
assign w10324 = ~w10321 & w10323;
assign w10325 = w10321 & ~w10323;
assign w10326 = ~w10324 & ~w10325;
assign w10327 = w10314 & w10326;
assign w10328 = ~w10314 & ~w10326;
assign w10329 = ~w10327 & ~w10328;
assign w10330 = ~w10302 & w10329;
assign w10331 = w10302 & ~w10329;
assign w10332 = ~w10330 & ~w10331;
assign w10333 = w10301 & w10332;
assign w10334 = ~w10301 & ~w10332;
assign w10335 = ~w10333 & ~w10334;
assign w10336 = ~w10288 & w10335;
assign w10337 = w10288 & ~w10335;
assign w10338 = ~w10336 & ~w10337;
assign w10339 = (~w10050 & ~w10052) | (~w10050 & w17178) | (~w10052 & w17178);
assign w10340 = (~w10196 & w10199) | (~w10196 & w17179) | (w10199 & w17179);
assign w10341 = pi12 & pi60;
assign w10342 = pi25 & pi47;
assign w10343 = pi24 & pi48;
assign w10344 = ~w10342 & ~w10343;
assign w10345 = pi25 & pi48;
assign w10346 = w10212 & w10345;
assign w10347 = ~w10344 & ~w10346;
assign w10348 = w10341 & ~w10347;
assign w10349 = ~w10341 & w10347;
assign w10350 = ~w10348 & ~w10349;
assign w10351 = ~w10340 & ~w10350;
assign w10352 = w10340 & w10350;
assign w10353 = ~w10351 & ~w10352;
assign w10354 = pi09 & pi63;
assign w10355 = pi10 & pi62;
assign w10356 = pi11 & pi61;
assign w10357 = ~w10355 & ~w10356;
assign w10358 = pi11 & pi62;
assign w10359 = w10138 & w10358;
assign w10360 = ~w10357 & ~w10359;
assign w10361 = w10354 & ~w10360;
assign w10362 = ~w10354 & w10360;
assign w10363 = ~w10361 & ~w10362;
assign w10364 = w10353 & ~w10363;
assign w10365 = ~w10353 & w10363;
assign w10366 = ~w10364 & ~w10365;
assign w10367 = pi35 & pi37;
assign w10368 = pi21 & pi51;
assign w10369 = pi22 & pi50;
assign w10370 = ~w10368 & ~w10369;
assign w10371 = pi22 & pi51;
assign w10372 = w10106 & w10371;
assign w10373 = ~w10370 & ~w10372;
assign w10374 = w10367 & ~w10373;
assign w10375 = ~w10367 & w10373;
assign w10376 = ~w10374 & ~w10375;
assign w10377 = pi32 & pi40;
assign w10378 = pi23 & pi49;
assign w10379 = ~w10206 & ~w10378;
assign w10380 = w10206 & w10378;
assign w10381 = ~w10379 & ~w10380;
assign w10382 = w10377 & ~w10381;
assign w10383 = ~w10377 & w10381;
assign w10384 = ~w10382 & ~w10383;
assign w10385 = ~w10376 & ~w10384;
assign w10386 = w10376 & w10384;
assign w10387 = ~w10385 & ~w10386;
assign w10388 = pi17 & pi55;
assign w10389 = ~w10109 & ~w10183;
assign w10390 = w10109 & w10183;
assign w10391 = ~w10389 & ~w10390;
assign w10392 = w10388 & ~w10391;
assign w10393 = ~w10388 & w10391;
assign w10394 = ~w10392 & ~w10393;
assign w10395 = w10387 & ~w10394;
assign w10396 = ~w10387 & w10394;
assign w10397 = ~w10395 & ~w10396;
assign w10398 = w10366 & w10397;
assign w10399 = ~w10366 & ~w10397;
assign w10400 = ~w10398 & ~w10399;
assign w10401 = ~w10339 & w10400;
assign w10402 = w10339 & ~w10400;
assign w10403 = ~w10401 & ~w10402;
assign w10404 = ~w10029 & ~w10033;
assign w10405 = w10203 & ~w10205;
assign w10406 = ~w10207 & ~w10405;
assign w10407 = w10212 & ~w10215;
assign w10408 = ~w10217 & ~w10407;
assign w10409 = ~w10406 & ~w10408;
assign w10410 = w10406 & w10408;
assign w10411 = ~w10409 & ~w10410;
assign w10412 = ~w9833 & ~w10140;
assign w10413 = ~w10139 & ~w10412;
assign w10414 = ~w10411 & ~w10413;
assign w10415 = w10411 & w10413;
assign w10416 = ~w10414 & ~w10415;
assign w10417 = (~w10021 & ~w10023) | (~w10021 & w16934) | (~w10023 & w16934);
assign w10418 = ~w10416 & w10417;
assign w10419 = w10416 & ~w10417;
assign w10420 = ~w10418 & ~w10419;
assign w10421 = pi14 & pi58;
assign w10422 = pi15 & pi57;
assign w10423 = ~w10421 & ~w10422;
assign w10424 = pi15 & pi58;
assign w10425 = w10203 & w10424;
assign w10426 = ~w10423 & ~w10425;
assign w10427 = w10195 & ~w10426;
assign w10428 = ~w10195 & w10426;
assign w10429 = ~w10427 & ~w10428;
assign w10430 = pi27 & pi45;
assign w10431 = pi28 & pi44;
assign w10432 = ~w10430 & ~w10431;
assign w10433 = pi28 & pi45;
assign w10434 = w9928 & w10433;
assign w10435 = ~w10432 & ~w10434;
assign w10436 = w10216 & ~w10435;
assign w10437 = ~w10216 & w10435;
assign w10438 = ~w10436 & ~w10437;
assign w10439 = ~w10429 & ~w10438;
assign w10440 = w10429 & w10438;
assign w10441 = ~w10439 & ~w10440;
assign w10442 = pi19 & pi53;
assign w10443 = pi34 & pi38;
assign w10444 = pi33 & pi39;
assign w10445 = ~w10443 & ~w10444;
assign w10446 = pi34 & pi39;
assign w10447 = w10118 & w10446;
assign w10448 = ~w10445 & ~w10447;
assign w10449 = w10442 & ~w10448;
assign w10450 = ~w10442 & w10448;
assign w10451 = ~w10449 & ~w10450;
assign w10452 = w10441 & ~w10451;
assign w10453 = ~w10441 & w10451;
assign w10454 = ~w10452 & ~w10453;
assign w10455 = ~w10420 & ~w10454;
assign w10456 = w10420 & w10454;
assign w10457 = ~w10455 & ~w10456;
assign w10458 = ~w10404 & w10457;
assign w10459 = w10404 & ~w10457;
assign w10460 = ~w10458 & ~w10459;
assign w10461 = ~w10403 & ~w10460;
assign w10462 = w10403 & w10460;
assign w10463 = ~w10461 & ~w10462;
assign w10464 = ~w10338 & ~w10463;
assign w10465 = w10338 & w10463;
assign w10466 = ~w10464 & ~w10465;
assign w10467 = ~w10287 & ~w10466;
assign w10468 = w10287 & w10466;
assign w10469 = ~w10467 & ~w10468;
assign w10470 = ~w10044 & ~w10241;
assign w10471 = ~w10469 & w10470;
assign w10472 = w10469 & ~w10470;
assign w10473 = ~w10471 & ~w10472;
assign w10474 = w10250 & ~w10473;
assign w10475 = ~w10250 & w10473;
assign w10476 = ~w10474 & ~w10475;
assign w10477 = ~w10286 & ~w10468;
assign w10478 = ~w10336 & ~w10465;
assign w10479 = (~w10458 & ~w10460) | (~w10458 & w17460) | (~w10460 & w17460);
assign w10480 = (~w10300 & ~w10301) | (~w10300 & w17461) | (~w10301 & w17461);
assign w10481 = (~w10419 & ~w10420) | (~w10419 & w17180) | (~w10420 & w17180);
assign w10482 = ~w10307 & ~w10313;
assign w10483 = (~w10409 & ~w10411) | (~w10409 & w17181) | (~w10411 & w17181);
assign w10484 = pi33 & pi40;
assign w10485 = pi32 & pi41;
assign w10486 = ~w10484 & ~w10485;
assign w10487 = pi33 & pi41;
assign w10488 = w10377 & w10487;
assign w10489 = ~w10486 & ~w10488;
assign w10490 = w10258 & ~w10489;
assign w10491 = ~w10258 & w10489;
assign w10492 = ~w10490 & ~w10491;
assign w10493 = ~w10483 & ~w10492;
assign w10494 = w10483 & w10492;
assign w10495 = ~w10493 & ~w10494;
assign w10496 = w10482 & ~w10495;
assign w10497 = ~w10482 & w10495;
assign w10498 = ~w10496 & ~w10497;
assign w10499 = (~w10327 & ~w10329) | (~w10327 & w17182) | (~w10329 & w17182);
assign w10500 = ~w10498 & w10499;
assign w10501 = w10498 & ~w10499;
assign w10502 = ~w10500 & ~w10501;
assign w10503 = ~w10481 & w10502;
assign w10504 = w10481 & ~w10502;
assign w10505 = ~w10503 & ~w10504;
assign w10506 = ~w10480 & w10505;
assign w10507 = w10480 & ~w10505;
assign w10508 = ~w10506 & ~w10507;
assign w10509 = ~w10479 & w10508;
assign w10510 = w10479 & ~w10508;
assign w10511 = ~w10509 & ~w10510;
assign w10512 = ~w10478 & w10511;
assign w10513 = w10478 & ~w10511;
assign w10514 = ~w10512 & ~w10513;
assign w10515 = (~w10439 & ~w10441) | (~w10439 & w17816) | (~w10441 & w17816);
assign w10516 = (~w10351 & ~w10353) | (~w10351 & w17462) | (~w10353 & w17462);
assign w10517 = (~w10319 & ~w10321) | (~w10319 & w17609) | (~w10321 & w17609);
assign w10518 = ~w10516 & ~w10517;
assign w10519 = w10516 & w10517;
assign w10520 = ~w10518 & ~w10519;
assign w10521 = w10515 & ~w10520;
assign w10522 = ~w10515 & w10520;
assign w10523 = ~w10521 & ~w10522;
assign w10524 = ~w10398 & ~w10401;
assign w10525 = ~w10523 & w10524;
assign w10526 = w10523 & ~w10524;
assign w10527 = ~w10525 & ~w10526;
assign w10528 = (~w10385 & ~w10387) | (~w10385 & w17817) | (~w10387 & w17817);
assign w10529 = pi13 & pi60;
assign w10530 = w10367 & ~w10370;
assign w10531 = (w10529 & w10530) | (w10529 & w17463) | (w10530 & w17463);
assign w10532 = ~w10530 & w17464;
assign w10533 = ~w10531 & ~w10532;
assign w10534 = w10442 & ~w10445;
assign w10535 = ~w10447 & ~w10534;
assign w10536 = ~w10533 & w10535;
assign w10537 = w10533 & ~w10535;
assign w10538 = ~w10536 & ~w10537;
assign w10539 = w10354 & ~w10357;
assign w10540 = ~w10359 & ~w10539;
assign w10541 = w10341 & ~w10344;
assign w10542 = ~w10346 & ~w10541;
assign w10543 = ~w10540 & ~w10542;
assign w10544 = w10540 & w10542;
assign w10545 = ~w10543 & ~w10544;
assign w10546 = ~w10388 & ~w10390;
assign w10547 = ~w10389 & ~w10546;
assign w10548 = ~w10545 & ~w10547;
assign w10549 = w10545 & w10547;
assign w10550 = ~w10548 & ~w10549;
assign w10551 = w10538 & w10550;
assign w10552 = ~w10538 & ~w10550;
assign w10553 = ~w10551 & ~w10552;
assign w10554 = ~w10528 & w10553;
assign w10555 = w10528 & ~w10553;
assign w10556 = ~w10554 & ~w10555;
assign w10557 = w10527 & w10556;
assign w10558 = ~w10527 & ~w10556;
assign w10559 = ~w10557 & ~w10558;
assign w10560 = (w10559 & w10282) | (w10559 & w17610) | (w10282 & w17610);
assign w10561 = ~w10282 & w17611;
assign w10562 = ~w10560 & ~w10561;
assign w10563 = (~w10292 & ~w10294) | (~w10292 & w17183) | (~w10294 & w17183);
assign w10564 = ~w10377 & ~w10380;
assign w10565 = ~w10379 & ~w10564;
assign w10566 = pi17 & pi56;
assign w10567 = pi26 & pi47;
assign w10568 = pi27 & pi46;
assign w10569 = ~w10567 & ~w10568;
assign w10570 = pi27 & pi47;
assign w10571 = w10216 & w10570;
assign w10572 = ~w10569 & ~w10571;
assign w10573 = w10566 & ~w10572;
assign w10574 = ~w10566 & w10572;
assign w10575 = ~w10573 & ~w10574;
assign w10576 = w10565 & ~w10575;
assign w10577 = ~w10565 & w10575;
assign w10578 = ~w10576 & ~w10577;
assign w10579 = pi14 & pi59;
assign w10580 = pi16 & pi57;
assign w10581 = ~w10424 & ~w10580;
assign w10582 = pi16 & pi58;
assign w10583 = w10422 & w10582;
assign w10584 = ~w10581 & ~w10583;
assign w10585 = w10579 & ~w10584;
assign w10586 = ~w10579 & w10584;
assign w10587 = ~w10585 & ~w10586;
assign w10588 = w10578 & ~w10587;
assign w10589 = ~w10578 & w10587;
assign w10590 = ~w10588 & ~w10589;
assign w10591 = pi23 & pi50;
assign w10592 = pi62 & w4629;
assign w10593 = ~pi37 & ~w10358;
assign w10594 = ~w10592 & ~w10593;
assign w10595 = w10591 & ~w10594;
assign w10596 = ~w10591 & w10594;
assign w10597 = ~w10595 & ~w10596;
assign w10598 = pi18 & pi55;
assign w10599 = pi24 & pi49;
assign w10600 = pi19 & pi54;
assign w10601 = ~w10599 & ~w10600;
assign w10602 = w10599 & w10600;
assign w10603 = ~w10601 & ~w10602;
assign w10604 = w10598 & ~w10603;
assign w10605 = ~w10598 & w10603;
assign w10606 = ~w10604 & ~w10605;
assign w10607 = ~w10597 & ~w10606;
assign w10608 = w10597 & w10606;
assign w10609 = ~w10607 & ~w10608;
assign w10610 = pi20 & pi53;
assign w10611 = pi21 & pi52;
assign w10612 = ~w10610 & ~w10611;
assign w10613 = pi21 & pi53;
assign w10614 = w10109 & w10613;
assign w10615 = ~w10612 & ~w10614;
assign w10616 = w10371 & ~w10615;
assign w10617 = ~w10371 & w10615;
assign w10618 = ~w10616 & ~w10617;
assign w10619 = w10609 & ~w10618;
assign w10620 = ~w10609 & w10618;
assign w10621 = ~w10619 & ~w10620;
assign w10622 = w10590 & w10621;
assign w10623 = ~w10590 & ~w10621;
assign w10624 = ~w10622 & ~w10623;
assign w10625 = w10563 & ~w10624;
assign w10626 = ~w10563 & w10624;
assign w10627 = ~w10625 & ~w10626;
assign w10628 = ~w10270 & ~w10275;
assign w10629 = w10195 & ~w10423;
assign w10630 = ~w10425 & ~w10629;
assign w10631 = w10216 & ~w10432;
assign w10632 = ~w10434 & ~w10631;
assign w10633 = ~w10630 & ~w10632;
assign w10634 = w10630 & w10632;
assign w10635 = ~w10633 & ~w10634;
assign w10636 = w10162 & ~w10257;
assign w10637 = ~w10259 & ~w10636;
assign w10638 = ~w10635 & w10637;
assign w10639 = w10635 & ~w10637;
assign w10640 = ~w10638 & ~w10639;
assign w10641 = (~w10264 & ~w10266) | (~w10264 & w16935) | (~w10266 & w16935);
assign w10642 = ~w10640 & w10641;
assign w10643 = w10640 & ~w10641;
assign w10644 = ~w10642 & ~w10643;
assign w10645 = pi29 & pi44;
assign w10646 = pi30 & pi43;
assign w10647 = ~w10645 & ~w10646;
assign w10648 = pi30 & pi44;
assign w10649 = w10162 & w10648;
assign w10650 = ~w10647 & ~w10649;
assign w10651 = w10433 & ~w10650;
assign w10652 = ~w10433 & w10650;
assign w10653 = ~w10651 & ~w10652;
assign w10654 = pi10 & pi63;
assign w10655 = pi12 & pi61;
assign w10656 = ~w10654 & ~w10655;
assign w10657 = w10654 & w10655;
assign w10658 = ~w10656 & ~w10657;
assign w10659 = w10345 & ~w10658;
assign w10660 = ~w10345 & w10658;
assign w10661 = ~w10659 & ~w10660;
assign w10662 = ~w10653 & ~w10661;
assign w10663 = w10653 & w10661;
assign w10664 = ~w10662 & ~w10663;
assign w10665 = pi36 & pi37;
assign w10666 = pi35 & pi38;
assign w10667 = ~w10665 & ~w10666;
assign w10668 = pi36 & pi38;
assign w10669 = w10367 & w10668;
assign w10670 = ~w10667 & ~w10669;
assign w10671 = w10446 & ~w10670;
assign w10672 = ~w10446 & w10670;
assign w10673 = ~w10671 & ~w10672;
assign w10674 = w10664 & ~w10673;
assign w10675 = ~w10664 & w10673;
assign w10676 = ~w10674 & ~w10675;
assign w10677 = ~w10644 & ~w10676;
assign w10678 = w10644 & w10676;
assign w10679 = ~w10677 & ~w10678;
assign w10680 = ~w10628 & w10679;
assign w10681 = w10628 & ~w10679;
assign w10682 = ~w10680 & ~w10681;
assign w10683 = ~w10627 & ~w10682;
assign w10684 = w10627 & w10682;
assign w10685 = ~w10683 & ~w10684;
assign w10686 = ~w10562 & ~w10685;
assign w10687 = w10562 & w10685;
assign w10688 = ~w10686 & ~w10687;
assign w10689 = ~w10514 & ~w10688;
assign w10690 = w10514 & w10688;
assign w10691 = ~w10689 & ~w10690;
assign w10692 = w10477 & ~w10691;
assign w10693 = ~w10477 & w10691;
assign w10694 = ~w10692 & ~w10693;
assign w10695 = (w7754 & w17818) | (w7754 & w17819) | (w17818 & w17819);
assign w10696 = w10694 & w10695;
assign w10697 = ~w10694 & ~w10695;
assign w10698 = ~w10696 & ~w10697;
assign w10699 = ~w10512 & ~w10690;
assign w10700 = (~w10560 & ~w10562) | (~w10560 & w17820) | (~w10562 & w17820);
assign w10701 = (~w10680 & ~w10682) | (~w10680 & w17467) | (~w10682 & w17467);
assign w10702 = (~w10526 & ~w10527) | (~w10526 & w17468) | (~w10527 & w17468);
assign w10703 = (~w10576 & ~w10578) | (~w10576 & w17614) | (~w10578 & w17614);
assign w10704 = (~w10543 & ~w10545) | (~w10543 & w17469) | (~w10545 & w17469);
assign w10705 = (~w10531 & ~w10533) | (~w10531 & w17615) | (~w10533 & w17615);
assign w10706 = ~w10704 & ~w10705;
assign w10707 = w10704 & w10705;
assign w10708 = ~w10706 & ~w10707;
assign w10709 = w10703 & ~w10708;
assign w10710 = ~w10703 & w10708;
assign w10711 = ~w10709 & ~w10710;
assign w10712 = (~w10551 & ~w10553) | (~w10551 & w17616) | (~w10553 & w17616);
assign w10713 = (~w10518 & ~w10520) | (~w10518 & w17617) | (~w10520 & w17617);
assign w10714 = ~w10712 & ~w10713;
assign w10715 = w10712 & w10713;
assign w10716 = ~w10714 & ~w10715;
assign w10717 = w10711 & w10716;
assign w10718 = ~w10711 & ~w10716;
assign w10719 = ~w10717 & ~w10718;
assign w10720 = ~w10702 & w10719;
assign w10721 = w10702 & ~w10719;
assign w10722 = ~w10720 & ~w10721;
assign w10723 = ~w10701 & w10722;
assign w10724 = w10701 & ~w10722;
assign w10725 = ~w10723 & ~w10724;
assign w10726 = ~w10700 & w10725;
assign w10727 = w10700 & ~w10725;
assign w10728 = ~w10726 & ~w10727;
assign w10729 = ~w10493 & ~w10497;
assign w10730 = w10258 & ~w10486;
assign w10731 = ~w10488 & ~w10730;
assign w10732 = w10446 & ~w10667;
assign w10733 = ~w10669 & ~w10732;
assign w10734 = ~w10731 & ~w10733;
assign w10735 = w10731 & w10733;
assign w10736 = ~w10734 & ~w10735;
assign w10737 = pi14 & pi60;
assign w10738 = pi15 & pi59;
assign w10739 = ~w10582 & ~w10738;
assign w10740 = pi16 & pi59;
assign w10741 = w10424 & w10740;
assign w10742 = ~w10739 & ~w10741;
assign w10743 = w10737 & ~w10742;
assign w10744 = ~w10737 & w10742;
assign w10745 = ~w10743 & ~w10744;
assign w10746 = ~w10736 & w10745;
assign w10747 = w10736 & ~w10745;
assign w10748 = ~w10746 & ~w10747;
assign w10749 = ~w10607 & ~w10619;
assign w10750 = w10748 & ~w10749;
assign w10751 = ~w10748 & w10749;
assign w10752 = ~w10750 & ~w10751;
assign w10753 = w10729 & ~w10752;
assign w10754 = ~w10729 & w10752;
assign w10755 = ~w10753 & ~w10754;
assign w10756 = ~w10622 & ~w10626;
assign w10757 = (~w10643 & ~w10644) | (~w10643 & w17184) | (~w10644 & w17184);
assign w10758 = ~w10756 & ~w10757;
assign w10759 = w10756 & w10757;
assign w10760 = ~w10758 & ~w10759;
assign w10761 = w10755 & w10760;
assign w10762 = ~w10755 & ~w10760;
assign w10763 = ~w10761 & ~w10762;
assign w10764 = (w10763 & w10509) | (w10763 & w17618) | (w10509 & w17618);
assign w10765 = ~w10509 & w17619;
assign w10766 = ~w10764 & ~w10765;
assign w10767 = w10566 & ~w10569;
assign w10768 = ~w10571 & ~w10767;
assign w10769 = w10433 & ~w10647;
assign w10770 = ~w10649 & ~w10769;
assign w10771 = ~w10768 & ~w10770;
assign w10772 = w10768 & w10770;
assign w10773 = ~w10771 & ~w10772;
assign w10774 = w10579 & ~w10581;
assign w10775 = ~w10583 & ~w10774;
assign w10776 = ~w10773 & w10775;
assign w10777 = w10773 & ~w10775;
assign w10778 = ~w10776 & ~w10777;
assign w10779 = ~w10598 & ~w10602;
assign w10780 = ~w10601 & ~w10779;
assign w10781 = w10371 & ~w10612;
assign w10782 = ~w10614 & ~w10781;
assign w10783 = w10780 & ~w10782;
assign w10784 = ~w10780 & w10782;
assign w10785 = ~w10783 & ~w10784;
assign w10786 = ~w10345 & ~w10657;
assign w10787 = ~w10656 & ~w10786;
assign w10788 = ~w10785 & ~w10787;
assign w10789 = w10785 & w10787;
assign w10790 = ~w10788 & ~w10789;
assign w10791 = (~w10662 & ~w10664) | (~w10662 & w17470) | (~w10664 & w17470);
assign w10792 = ~w10790 & w10791;
assign w10793 = w10790 & ~w10791;
assign w10794 = ~w10792 & ~w10793;
assign w10795 = w10778 & w10794;
assign w10796 = ~w10778 & ~w10794;
assign w10797 = ~w10795 & ~w10796;
assign w10798 = (w10797 & w10503) | (w10797 & w17471) | (w10503 & w17471);
assign w10799 = ~w10503 & w17472;
assign w10800 = ~w10798 & ~w10799;
assign w10801 = ~w10633 & ~w10639;
assign w10802 = pi13 & pi61;
assign w10803 = pi12 & pi62;
assign w10804 = ~w10802 & ~w10803;
assign w10805 = pi13 & pi62;
assign w10806 = w10655 & w10805;
assign w10807 = ~w10804 & ~w10806;
assign w10808 = w10591 & ~w10593;
assign w10809 = ~w10592 & ~w10808;
assign w10810 = w10807 & ~w10809;
assign w10811 = ~w10807 & w10809;
assign w10812 = ~w10810 & ~w10811;
assign w10813 = pi29 & pi45;
assign w10814 = pi17 & pi57;
assign w10815 = ~w10648 & ~w10814;
assign w10816 = w10648 & w10814;
assign w10817 = ~w10815 & ~w10816;
assign w10818 = w10813 & ~w10817;
assign w10819 = ~w10813 & w10817;
assign w10820 = ~w10818 & ~w10819;
assign w10821 = w10812 & ~w10820;
assign w10822 = ~w10812 & w10820;
assign w10823 = ~w10821 & ~w10822;
assign w10824 = w10801 & ~w10823;
assign w10825 = ~w10801 & w10823;
assign w10826 = ~w10824 & ~w10825;
assign w10827 = pi11 & pi63;
assign w10828 = pi31 & pi43;
assign w10829 = pi32 & pi42;
assign w10830 = ~w10828 & ~w10829;
assign w10831 = pi32 & pi43;
assign w10832 = w10258 & w10831;
assign w10833 = ~w10830 & ~w10832;
assign w10834 = w10827 & ~w10833;
assign w10835 = ~w10827 & w10833;
assign w10836 = ~w10834 & ~w10835;
assign w10837 = pi18 & pi56;
assign w10838 = pi25 & pi49;
assign w10839 = ~w10837 & ~w10838;
assign w10840 = w10837 & w10838;
assign w10841 = ~w10839 & ~w10840;
assign w10842 = w10487 & ~w10841;
assign w10843 = ~w10487 & w10841;
assign w10844 = ~w10842 & ~w10843;
assign w10845 = ~w10836 & ~w10844;
assign w10846 = w10836 & w10844;
assign w10847 = ~w10845 & ~w10846;
assign w10848 = pi26 & pi48;
assign w10849 = pi28 & pi46;
assign w10850 = ~w10570 & ~w10849;
assign w10851 = pi28 & pi47;
assign w10852 = w10568 & w10851;
assign w10853 = ~w10850 & ~w10852;
assign w10854 = w10848 & ~w10853;
assign w10855 = ~w10848 & w10853;
assign w10856 = ~w10854 & ~w10855;
assign w10857 = w10847 & ~w10856;
assign w10858 = ~w10847 & w10856;
assign w10859 = ~w10857 & ~w10858;
assign w10860 = pi20 & pi54;
assign w10861 = pi35 & pi39;
assign w10862 = pi34 & pi40;
assign w10863 = ~w10861 & ~w10862;
assign w10864 = pi35 & pi40;
assign w10865 = w10446 & w10864;
assign w10866 = ~w10863 & ~w10865;
assign w10867 = w10860 & ~w10866;
assign w10868 = ~w10860 & w10866;
assign w10869 = ~w10867 & ~w10868;
assign w10870 = pi22 & pi52;
assign w10871 = pi19 & pi55;
assign w10872 = ~w10613 & ~w10871;
assign w10873 = w10613 & w10871;
assign w10874 = ~w10872 & ~w10873;
assign w10875 = w10870 & ~w10874;
assign w10876 = ~w10870 & w10874;
assign w10877 = ~w10875 & ~w10876;
assign w10878 = ~w10869 & ~w10877;
assign w10879 = w10869 & w10877;
assign w10880 = ~w10878 & ~w10879;
assign w10881 = pi23 & pi51;
assign w10882 = pi24 & pi50;
assign w10883 = ~w10881 & ~w10882;
assign w10884 = pi24 & pi51;
assign w10885 = w10591 & w10884;
assign w10886 = ~w10883 & ~w10885;
assign w10887 = w10668 & ~w10886;
assign w10888 = ~w10668 & w10886;
assign w10889 = ~w10887 & ~w10888;
assign w10890 = w10880 & ~w10889;
assign w10891 = ~w10880 & w10889;
assign w10892 = ~w10890 & ~w10891;
assign w10893 = w10859 & w10892;
assign w10894 = ~w10859 & ~w10892;
assign w10895 = ~w10893 & ~w10894;
assign w10896 = ~w10826 & ~w10895;
assign w10897 = w10826 & w10895;
assign w10898 = ~w10896 & ~w10897;
assign w10899 = ~w10800 & ~w10898;
assign w10900 = w10800 & w10898;
assign w10901 = ~w10899 & ~w10900;
assign w10902 = w10766 & w10901;
assign w10903 = ~w10766 & ~w10901;
assign w10904 = ~w10902 & ~w10903;
assign w10905 = w10728 & w10904;
assign w10906 = ~w10728 & ~w10904;
assign w10907 = ~w10905 & ~w10906;
assign w10908 = w10699 & ~w10907;
assign w10909 = ~w10699 & w10907;
assign w10910 = ~w10908 & ~w10909;
assign w10911 = ~w10471 & ~w10692;
assign w10912 = (~w8795 & w17620) | (~w8795 & w17621) | (w17620 & w17621);
assign w10913 = w10910 & w10912;
assign w10914 = ~w10910 & ~w10912;
assign w10915 = ~w10913 & ~w10914;
assign w10916 = ~w10726 & ~w10905;
assign w10917 = (~w10771 & ~w10773) | (~w10771 & w17185) | (~w10773 & w17185);
assign w10918 = (~w10734 & ~w10736) | (~w10734 & w16770) | (~w10736 & w16770);
assign w10919 = (~w10783 & ~w10785) | (~w10783 & w16771) | (~w10785 & w16771);
assign w10920 = ~w10918 & ~w10919;
assign w10921 = w10918 & w10919;
assign w10922 = ~w10920 & ~w10921;
assign w10923 = w10917 & ~w10922;
assign w10924 = ~w10917 & w10922;
assign w10925 = ~w10923 & ~w10924;
assign w10926 = (~w10893 & ~w10895) | (~w10893 & w17821) | (~w10895 & w17821);
assign w10927 = ~w10925 & w10926;
assign w10928 = w10925 & ~w10926;
assign w10929 = ~w10927 & ~w10928;
assign w10930 = ~w10821 & ~w10825;
assign w10931 = w10668 & ~w10883;
assign w10932 = ~w10885 & ~w10931;
assign w10933 = w10860 & ~w10863;
assign w10934 = ~w10865 & ~w10933;
assign w10935 = ~w10932 & ~w10934;
assign w10936 = w10932 & w10934;
assign w10937 = ~w10935 & ~w10936;
assign w10938 = ~w10870 & ~w10873;
assign w10939 = ~w10872 & ~w10938;
assign w10940 = ~w10937 & ~w10939;
assign w10941 = w10937 & w10939;
assign w10942 = ~w10940 & ~w10941;
assign w10943 = (~w10806 & w10809) | (~w10806 & w17186) | (w10809 & w17186);
assign w10944 = ~w10487 & ~w10840;
assign w10945 = ~w10839 & ~w10944;
assign w10946 = w10827 & ~w10830;
assign w10947 = ~w10832 & ~w10946;
assign w10948 = w10945 & ~w10947;
assign w10949 = ~w10945 & w10947;
assign w10950 = ~w10948 & ~w10949;
assign w10951 = w10943 & ~w10950;
assign w10952 = ~w10943 & w10950;
assign w10953 = ~w10951 & ~w10952;
assign w10954 = w10942 & w10953;
assign w10955 = ~w10942 & ~w10953;
assign w10956 = ~w10954 & ~w10955;
assign w10957 = ~w10930 & w10956;
assign w10958 = w10930 & ~w10956;
assign w10959 = ~w10957 & ~w10958;
assign w10960 = w10929 & w10959;
assign w10961 = ~w10929 & ~w10959;
assign w10962 = ~w10960 & ~w10961;
assign w10963 = (w10962 & w10723) | (w10962 & w17622) | (w10723 & w17622);
assign w10964 = ~w10723 & w17623;
assign w10965 = ~w10963 & ~w10964;
assign w10966 = (~w10714 & ~w10716) | (~w10714 & w17822) | (~w10716 & w17822);
assign w10967 = ~w10813 & ~w10816;
assign w10968 = ~w10815 & ~w10967;
assign w10969 = w10848 & ~w10850;
assign w10970 = ~w10852 & ~w10969;
assign w10971 = w10968 & ~w10970;
assign w10972 = ~w10968 & w10970;
assign w10973 = ~w10971 & ~w10972;
assign w10974 = w10737 & ~w10739;
assign w10975 = ~w10741 & ~w10974;
assign w10976 = ~w10973 & w10975;
assign w10977 = w10973 & ~w10975;
assign w10978 = ~w10976 & ~w10977;
assign w10979 = (~w10878 & ~w10880) | (~w10878 & w16936) | (~w10880 & w16936);
assign w10980 = (~w10845 & ~w10847) | (~w10845 & w16937) | (~w10847 & w16937);
assign w10981 = ~w10979 & ~w10980;
assign w10982 = w10979 & w10980;
assign w10983 = ~w10981 & ~w10982;
assign w10984 = w10978 & w10983;
assign w10985 = ~w10978 & ~w10983;
assign w10986 = ~w10984 & ~w10985;
assign w10987 = ~w10966 & w10986;
assign w10988 = w10966 & ~w10986;
assign w10989 = ~w10987 & ~w10988;
assign w10990 = (~w10706 & ~w10708) | (~w10706 & w17624) | (~w10708 & w17624);
assign w10991 = pi23 & pi52;
assign w10992 = pi36 & pi39;
assign w10993 = ~w10864 & ~w10992;
assign w10994 = w10864 & w10992;
assign w10995 = ~w10993 & ~w10994;
assign w10996 = w10991 & ~w10995;
assign w10997 = ~w10991 & w10995;
assign w10998 = ~w10996 & ~w10997;
assign w10999 = pi30 & pi45;
assign w11000 = pi12 & pi63;
assign w11001 = pi19 & pi56;
assign w11002 = ~w11000 & ~w11001;
assign w11003 = w11000 & w11001;
assign w11004 = ~w11002 & ~w11003;
assign w11005 = w10999 & ~w11004;
assign w11006 = ~w10999 & w11004;
assign w11007 = ~w11005 & ~w11006;
assign w11008 = ~w10998 & ~w11007;
assign w11009 = w10998 & w11007;
assign w11010 = ~w11008 & ~w11009;
assign w11011 = ~pi37 & pi38;
assign w11012 = w10805 & ~w11011;
assign w11013 = ~w10805 & w11011;
assign w11014 = ~w11012 & ~w11013;
assign w11015 = w11010 & ~w11014;
assign w11016 = ~w11010 & w11014;
assign w11017 = ~w11015 & ~w11016;
assign w11018 = ~w10990 & w11017;
assign w11019 = w10990 & ~w11017;
assign w11020 = ~w11018 & ~w11019;
assign w11021 = pi14 & pi61;
assign w11022 = pi15 & pi60;
assign w11023 = ~w10740 & ~w11022;
assign w11024 = pi16 & pi60;
assign w11025 = w10738 & w11024;
assign w11026 = ~w11023 & ~w11025;
assign w11027 = w11021 & ~w11026;
assign w11028 = ~w11021 & w11026;
assign w11029 = ~w11027 & ~w11028;
assign w11030 = pi17 & pi58;
assign w11031 = pi26 & pi49;
assign w11032 = pi18 & pi57;
assign w11033 = ~w11031 & ~w11032;
assign w11034 = w11031 & w11032;
assign w11035 = ~w11033 & ~w11034;
assign w11036 = w11030 & ~w11035;
assign w11037 = ~w11030 & w11035;
assign w11038 = ~w11036 & ~w11037;
assign w11039 = ~w11029 & ~w11038;
assign w11040 = w11029 & w11038;
assign w11041 = ~w11039 & ~w11040;
assign w11042 = pi27 & pi48;
assign w11043 = pi29 & pi46;
assign w11044 = ~w10851 & ~w11043;
assign w11045 = pi29 & pi47;
assign w11046 = w10849 & w11045;
assign w11047 = ~w11044 & ~w11046;
assign w11048 = w11042 & ~w11047;
assign w11049 = ~w11042 & w11047;
assign w11050 = ~w11048 & ~w11049;
assign w11051 = w11041 & ~w11050;
assign w11052 = ~w11041 & w11050;
assign w11053 = ~w11051 & ~w11052;
assign w11054 = w11020 & w11053;
assign w11055 = ~w11020 & ~w11053;
assign w11056 = ~w11054 & ~w11055;
assign w11057 = w10989 & w11056;
assign w11058 = ~w10989 & ~w11056;
assign w11059 = ~w11057 & ~w11058;
assign w11060 = ~w10965 & ~w11059;
assign w11061 = w10965 & w11059;
assign w11062 = ~w11060 & ~w11061;
assign w11063 = (~w10798 & ~w10800) | (~w10798 & w17625) | (~w10800 & w17625);
assign w11064 = (~w10758 & ~w10760) | (~w10758 & w17474) | (~w10760 & w17474);
assign w11065 = ~w10750 & ~w10754;
assign w11066 = (~w10793 & ~w10794) | (~w10793 & w17626) | (~w10794 & w17626);
assign w11067 = pi31 & pi44;
assign w11068 = pi33 & pi42;
assign w11069 = ~w10831 & ~w11068;
assign w11070 = pi33 & pi43;
assign w11071 = w10829 & w11070;
assign w11072 = ~w11069 & ~w11071;
assign w11073 = w11067 & ~w11072;
assign w11074 = ~w11067 & w11072;
assign w11075 = ~w11073 & ~w11074;
assign w11076 = pi34 & pi41;
assign w11077 = pi20 & pi55;
assign w11078 = pi25 & pi50;
assign w11079 = ~w11077 & ~w11078;
assign w11080 = w11077 & w11078;
assign w11081 = ~w11079 & ~w11080;
assign w11082 = w11076 & ~w11081;
assign w11083 = ~w11076 & w11081;
assign w11084 = ~w11082 & ~w11083;
assign w11085 = ~w11075 & ~w11084;
assign w11086 = w11075 & w11084;
assign w11087 = ~w11085 & ~w11086;
assign w11088 = pi21 & pi54;
assign w11089 = pi22 & pi53;
assign w11090 = ~w10884 & ~w11089;
assign w11091 = w10884 & w11089;
assign w11092 = ~w11090 & ~w11091;
assign w11093 = w11088 & ~w11092;
assign w11094 = ~w11088 & w11092;
assign w11095 = ~w11093 & ~w11094;
assign w11096 = w11087 & ~w11095;
assign w11097 = ~w11087 & w11095;
assign w11098 = ~w11096 & ~w11097;
assign w11099 = ~w11066 & w11098;
assign w11100 = w11066 & ~w11098;
assign w11101 = ~w11099 & ~w11100;
assign w11102 = ~w11065 & w11101;
assign w11103 = w11065 & ~w11101;
assign w11104 = ~w11102 & ~w11103;
assign w11105 = ~w11064 & w11104;
assign w11106 = w11064 & ~w11104;
assign w11107 = ~w11105 & ~w11106;
assign w11108 = w11063 & ~w11107;
assign w11109 = ~w11063 & w11107;
assign w11110 = ~w11108 & ~w11109;
assign w11111 = (~w10764 & ~w10766) | (~w10764 & w17823) | (~w10766 & w17823);
assign w11112 = ~w11110 & w11111;
assign w11113 = w11110 & ~w11111;
assign w11114 = ~w11112 & ~w11113;
assign w11115 = w11062 & w11114;
assign w11116 = ~w11062 & ~w11114;
assign w11117 = ~w11115 & ~w11116;
assign w11118 = ~w10916 & w11117;
assign w11119 = w10916 & ~w11117;
assign w11120 = ~w11118 & ~w11119;
assign w11121 = ~w10693 & ~w10909;
assign w11122 = (w8795 & w17475) | (w8795 & w17476) | (w17475 & w17476);
assign w11123 = w11120 & w11122;
assign w11124 = ~w11120 & ~w11122;
assign w11125 = ~w11123 & ~w11124;
assign w11126 = ~w11113 & ~w11115;
assign w11127 = (~w10963 & ~w10965) | (~w10963 & w17824) | (~w10965 & w17824);
assign w11128 = ~w10987 & ~w11057;
assign w11129 = ~w10928 & ~w10960;
assign w11130 = ~w10954 & ~w10957;
assign w11131 = (~w10981 & ~w10983) | (~w10981 & w17187) | (~w10983 & w17187);
assign w11132 = pi13 & pi63;
assign w11133 = pi31 & pi45;
assign w11134 = pi32 & pi44;
assign w11135 = ~w11133 & ~w11134;
assign w11136 = pi32 & pi45;
assign w11137 = w11067 & w11136;
assign w11138 = ~w11135 & ~w11137;
assign w11139 = w11132 & ~w11138;
assign w11140 = ~w11132 & w11138;
assign w11141 = ~w11139 & ~w11140;
assign w11142 = pi19 & pi57;
assign w11143 = pi23 & pi53;
assign w11144 = ~w11142 & ~w11143;
assign w11145 = w11142 & w11143;
assign w11146 = ~w11144 & ~w11145;
assign w11147 = w11070 & ~w11146;
assign w11148 = ~w11070 & w11146;
assign w11149 = ~w11147 & ~w11148;
assign w11150 = ~w11141 & ~w11149;
assign w11151 = w11141 & w11149;
assign w11152 = ~w11150 & ~w11151;
assign w11153 = pi20 & pi56;
assign w11154 = pi21 & pi55;
assign w11155 = pi22 & pi54;
assign w11156 = ~w11154 & ~w11155;
assign w11157 = pi22 & pi55;
assign w11158 = w11088 & w11157;
assign w11159 = ~w11156 & ~w11158;
assign w11160 = w11153 & ~w11159;
assign w11161 = ~w11153 & w11159;
assign w11162 = ~w11160 & ~w11161;
assign w11163 = w11152 & ~w11162;
assign w11164 = ~w11152 & w11162;
assign w11165 = ~w11163 & ~w11164;
assign w11166 = ~w11131 & w11165;
assign w11167 = w11131 & ~w11165;
assign w11168 = ~w11166 & ~w11167;
assign w11169 = ~w11130 & w11168;
assign w11170 = w11130 & ~w11168;
assign w11171 = ~w11169 & ~w11170;
assign w11172 = ~w11129 & w11171;
assign w11173 = w11129 & ~w11171;
assign w11174 = ~w11172 & ~w11173;
assign w11175 = ~w11128 & w11174;
assign w11176 = w11128 & ~w11174;
assign w11177 = ~w11175 & ~w11176;
assign w11178 = ~w11127 & w11177;
assign w11179 = w11127 & ~w11177;
assign w11180 = ~w11178 & ~w11179;
assign w11181 = ~w10935 & ~w10941;
assign w11182 = (~w10948 & ~w10950) | (~w10948 & w17188) | (~w10950 & w17188);
assign w11183 = (~w10971 & ~w10973) | (~w10971 & w17189) | (~w10973 & w17189);
assign w11184 = ~w11182 & ~w11183;
assign w11185 = w11182 & w11183;
assign w11186 = ~w11184 & ~w11185;
assign w11187 = w11181 & ~w11186;
assign w11188 = ~w11181 & w11186;
assign w11189 = ~w11187 & ~w11188;
assign w11190 = (~w11018 & ~w11020) | (~w11018 & w17825) | (~w11020 & w17825);
assign w11191 = ~w11189 & w11190;
assign w11192 = w11189 & ~w11190;
assign w11193 = ~w11191 & ~w11192;
assign w11194 = ~w11076 & ~w11080;
assign w11195 = ~w11079 & ~w11194;
assign w11196 = w11042 & ~w11044;
assign w11197 = ~w11046 & ~w11196;
assign w11198 = w11195 & ~w11197;
assign w11199 = ~w11195 & w11197;
assign w11200 = ~w11198 & ~w11199;
assign w11201 = ~w10999 & ~w11003;
assign w11202 = ~w11002 & ~w11201;
assign w11203 = ~w11200 & ~w11202;
assign w11204 = w11200 & w11202;
assign w11205 = ~w11203 & ~w11204;
assign w11206 = ~w11085 & ~w11096;
assign w11207 = pi14 & pi62;
assign w11208 = ~pi37 & ~w10805;
assign w11209 = pi38 & ~w11208;
assign w11210 = ~w11207 & ~w11209;
assign w11211 = w11207 & w11209;
assign w11212 = ~w11210 & ~w11211;
assign w11213 = ~w10991 & ~w10994;
assign w11214 = ~w10993 & ~w11213;
assign w11215 = ~w11212 & w11214;
assign w11216 = w11212 & ~w11214;
assign w11217 = ~w11215 & ~w11216;
assign w11218 = ~w11206 & ~w11217;
assign w11219 = w11206 & w11217;
assign w11220 = ~w11218 & ~w11219;
assign w11221 = ~w11205 & ~w11220;
assign w11222 = w11205 & w11220;
assign w11223 = ~w11221 & ~w11222;
assign w11224 = ~w11193 & ~w11223;
assign w11225 = w11193 & w11223;
assign w11226 = ~w11224 & ~w11225;
assign w11227 = (~w11105 & ~w11107) | (~w11105 & w17627) | (~w11107 & w17627);
assign w11228 = w11226 & ~w11227;
assign w11229 = ~w11226 & w11227;
assign w11230 = ~w11228 & ~w11229;
assign w11231 = ~w11099 & ~w11102;
assign w11232 = ~w11030 & ~w11034;
assign w11233 = ~w11033 & ~w11232;
assign w11234 = w11021 & ~w11023;
assign w11235 = ~w11025 & ~w11234;
assign w11236 = w11233 & ~w11235;
assign w11237 = ~w11233 & w11235;
assign w11238 = ~w11236 & ~w11237;
assign w11239 = w11067 & ~w11069;
assign w11240 = ~w11071 & ~w11239;
assign w11241 = ~w11238 & w11240;
assign w11242 = w11238 & ~w11240;
assign w11243 = ~w11241 & ~w11242;
assign w11244 = (~w11039 & ~w11041) | (~w11039 & w16938) | (~w11041 & w16938);
assign w11245 = (~w11008 & ~w11010) | (~w11008 & w16939) | (~w11010 & w16939);
assign w11246 = ~w11244 & ~w11245;
assign w11247 = w11244 & w11245;
assign w11248 = ~w11246 & ~w11247;
assign w11249 = w11243 & w11248;
assign w11250 = ~w11243 & ~w11248;
assign w11251 = ~w11249 & ~w11250;
assign w11252 = ~w11231 & w11251;
assign w11253 = w11231 & ~w11251;
assign w11254 = ~w11252 & ~w11253;
assign w11255 = (~w10920 & ~w10922) | (~w10920 & w16940) | (~w10922 & w16940);
assign w11256 = pi28 & pi48;
assign w11257 = pi30 & pi46;
assign w11258 = ~w11045 & ~w11257;
assign w11259 = pi30 & pi47;
assign w11260 = w11043 & w11259;
assign w11261 = ~w11258 & ~w11260;
assign w11262 = w11256 & ~w11261;
assign w11263 = ~w11256 & w11261;
assign w11264 = ~w11262 & ~w11263;
assign w11265 = pi34 & pi42;
assign w11266 = pi36 & pi40;
assign w11267 = pi35 & pi41;
assign w11268 = ~w11266 & ~w11267;
assign w11269 = pi36 & pi41;
assign w11270 = w10864 & w11269;
assign w11271 = ~w11268 & ~w11270;
assign w11272 = w11265 & ~w11271;
assign w11273 = ~w11265 & w11271;
assign w11274 = ~w11272 & ~w11273;
assign w11275 = ~w11264 & ~w11274;
assign w11276 = w11264 & w11274;
assign w11277 = ~w11275 & ~w11276;
assign w11278 = pi37 & pi39;
assign w11279 = pi25 & pi51;
assign w11280 = pi24 & pi52;
assign w11281 = ~w11279 & ~w11280;
assign w11282 = pi25 & pi52;
assign w11283 = w10884 & w11282;
assign w11284 = ~w11281 & ~w11283;
assign w11285 = w11278 & ~w11284;
assign w11286 = ~w11278 & w11284;
assign w11287 = ~w11285 & ~w11286;
assign w11288 = w11277 & ~w11287;
assign w11289 = ~w11277 & w11287;
assign w11290 = ~w11288 & ~w11289;
assign w11291 = ~w11255 & w11290;
assign w11292 = w11255 & ~w11290;
assign w11293 = ~w11291 & ~w11292;
assign w11294 = ~w11088 & ~w11091;
assign w11295 = ~w11090 & ~w11294;
assign w11296 = pi15 & pi61;
assign w11297 = pi17 & pi59;
assign w11298 = ~w11024 & ~w11297;
assign w11299 = pi17 & pi60;
assign w11300 = w10740 & w11299;
assign w11301 = ~w11298 & ~w11300;
assign w11302 = w11296 & ~w11301;
assign w11303 = ~w11296 & w11301;
assign w11304 = ~w11302 & ~w11303;
assign w11305 = w11295 & ~w11304;
assign w11306 = ~w11295 & w11304;
assign w11307 = ~w11305 & ~w11306;
assign w11308 = pi18 & pi58;
assign w11309 = pi26 & pi50;
assign w11310 = pi27 & pi49;
assign w11311 = ~w11309 & ~w11310;
assign w11312 = pi27 & pi50;
assign w11313 = w11031 & w11312;
assign w11314 = ~w11311 & ~w11313;
assign w11315 = w11308 & ~w11314;
assign w11316 = ~w11308 & w11314;
assign w11317 = ~w11315 & ~w11316;
assign w11318 = w11307 & ~w11317;
assign w11319 = ~w11307 & w11317;
assign w11320 = ~w11318 & ~w11319;
assign w11321 = w11293 & w11320;
assign w11322 = ~w11293 & ~w11320;
assign w11323 = ~w11321 & ~w11322;
assign w11324 = w11254 & w11323;
assign w11325 = ~w11254 & ~w11323;
assign w11326 = ~w11324 & ~w11325;
assign w11327 = w11230 & w11326;
assign w11328 = ~w11230 & ~w11326;
assign w11329 = ~w11327 & ~w11328;
assign w11330 = w11180 & w11329;
assign w11331 = ~w11180 & ~w11329;
assign w11332 = ~w11330 & ~w11331;
assign w11333 = ~w11126 & w11332;
assign w11334 = w11126 & ~w11332;
assign w11335 = ~w11333 & ~w11334;
assign w11336 = (w7754 & w17826) | (w7754 & w17827) | (w17826 & w17827);
assign w11337 = w11335 & w11336;
assign w11338 = ~w11335 & ~w11336;
assign w11339 = ~w11337 & ~w11338;
assign w11340 = ~w11178 & ~w11330;
assign w11341 = (~w11228 & ~w11230) | (~w11228 & w17828) | (~w11230 & w17828);
assign w11342 = ~w11252 & ~w11324;
assign w11343 = ~w11192 & ~w11225;
assign w11344 = ~w11218 & ~w11222;
assign w11345 = (~w11246 & ~w11248) | (~w11246 & w17190) | (~w11248 & w17190);
assign w11346 = pi24 & pi53;
assign w11347 = pi23 & pi54;
assign w11348 = ~w11346 & ~w11347;
assign w11349 = pi24 & pi54;
assign w11350 = w11143 & w11349;
assign w11351 = ~w11348 & ~w11350;
assign w11352 = w11282 & ~w11351;
assign w11353 = ~w11282 & w11351;
assign w11354 = ~w11352 & ~w11353;
assign w11355 = pi34 & pi43;
assign w11356 = pi26 & pi51;
assign w11357 = ~w11157 & ~w11356;
assign w11358 = w11157 & w11356;
assign w11359 = ~w11357 & ~w11358;
assign w11360 = w11355 & ~w11359;
assign w11361 = ~w11355 & w11359;
assign w11362 = ~w11360 & ~w11361;
assign w11363 = ~w11354 & ~w11362;
assign w11364 = w11354 & w11362;
assign w11365 = ~w11363 & ~w11364;
assign w11366 = pi16 & pi61;
assign w11367 = pi33 & pi44;
assign w11368 = ~w11136 & ~w11367;
assign w11369 = pi33 & pi45;
assign w11370 = w11134 & w11369;
assign w11371 = ~w11368 & ~w11370;
assign w11372 = w11366 & ~w11371;
assign w11373 = ~w11366 & w11371;
assign w11374 = ~w11372 & ~w11373;
assign w11375 = w11365 & ~w11374;
assign w11376 = ~w11365 & w11374;
assign w11377 = ~w11375 & ~w11376;
assign w11378 = ~w11345 & w11377;
assign w11379 = w11345 & ~w11377;
assign w11380 = ~w11378 & ~w11379;
assign w11381 = ~w11344 & w11380;
assign w11382 = w11344 & ~w11380;
assign w11383 = ~w11381 & ~w11382;
assign w11384 = ~w11343 & w11383;
assign w11385 = w11343 & ~w11383;
assign w11386 = ~w11384 & ~w11385;
assign w11387 = ~w11342 & w11386;
assign w11388 = w11342 & ~w11386;
assign w11389 = ~w11387 & ~w11388;
assign w11390 = ~w11341 & w11389;
assign w11391 = w11341 & ~w11389;
assign w11392 = ~w11390 & ~w11391;
assign w11393 = ~w11172 & ~w11175;
assign w11394 = (~w11198 & ~w11200) | (~w11198 & w17191) | (~w11200 & w17191);
assign w11395 = (~w11236 & ~w11238) | (~w11236 & w16772) | (~w11238 & w16772);
assign w11396 = pi18 & pi59;
assign w11397 = ~w11299 & ~w11396;
assign w11398 = pi18 & pi60;
assign w11399 = w11297 & w11398;
assign w11400 = ~w11397 & ~w11399;
assign w11401 = w11278 & ~w11281;
assign w11402 = ~w11283 & ~w11401;
assign w11403 = w11400 & ~w11402;
assign w11404 = ~w11400 & w11402;
assign w11405 = ~w11403 & ~w11404;
assign w11406 = ~w11395 & w11405;
assign w11407 = w11395 & ~w11405;
assign w11408 = ~w11406 & ~w11407;
assign w11409 = w11394 & ~w11408;
assign w11410 = ~w11394 & w11408;
assign w11411 = ~w11409 & ~w11410;
assign w11412 = (~w11291 & ~w11293) | (~w11291 & w17192) | (~w11293 & w17192);
assign w11413 = ~w11411 & w11412;
assign w11414 = w11411 & ~w11412;
assign w11415 = ~w11413 & ~w11414;
assign w11416 = w11153 & ~w11156;
assign w11417 = ~w11158 & ~w11416;
assign w11418 = w11256 & ~w11258;
assign w11419 = ~w11260 & ~w11418;
assign w11420 = ~w11417 & ~w11419;
assign w11421 = w11417 & w11419;
assign w11422 = ~w11420 & ~w11421;
assign w11423 = w11132 & ~w11135;
assign w11424 = ~w11137 & ~w11423;
assign w11425 = ~w11422 & w11424;
assign w11426 = w11422 & ~w11424;
assign w11427 = ~w11425 & ~w11426;
assign w11428 = w11296 & ~w11298;
assign w11429 = ~w11300 & ~w11428;
assign w11430 = w11308 & ~w11311;
assign w11431 = ~w11313 & ~w11430;
assign w11432 = ~w11429 & ~w11431;
assign w11433 = w11429 & w11431;
assign w11434 = ~w11432 & ~w11433;
assign w11435 = ~w11070 & ~w11145;
assign w11436 = ~w11144 & ~w11435;
assign w11437 = ~w11434 & ~w11436;
assign w11438 = w11434 & w11436;
assign w11439 = ~w11437 & ~w11438;
assign w11440 = (~w11150 & ~w11152) | (~w11150 & w17829) | (~w11152 & w17829);
assign w11441 = ~w11439 & w11440;
assign w11442 = w11439 & ~w11440;
assign w11443 = ~w11441 & ~w11442;
assign w11444 = w11427 & w11443;
assign w11445 = ~w11427 & ~w11443;
assign w11446 = ~w11444 & ~w11445;
assign w11447 = w11415 & w11446;
assign w11448 = ~w11415 & ~w11446;
assign w11449 = ~w11447 & ~w11448;
assign w11450 = ~w11393 & w11449;
assign w11451 = w11393 & ~w11449;
assign w11452 = ~w11450 & ~w11451;
assign w11453 = (~w11275 & ~w11277) | (~w11275 & w17830) | (~w11277 & w17830);
assign w11454 = (~w11305 & ~w11307) | (~w11305 & w16941) | (~w11307 & w16941);
assign w11455 = ~w11211 & ~w11214;
assign w11456 = ~w11210 & ~w11455;
assign w11457 = ~w11454 & w11456;
assign w11458 = w11454 & ~w11456;
assign w11459 = ~w11457 & ~w11458;
assign w11460 = w11453 & ~w11459;
assign w11461 = ~w11453 & w11459;
assign w11462 = ~w11460 & ~w11461;
assign w11463 = ~w11166 & ~w11169;
assign w11464 = ~w11462 & w11463;
assign w11465 = w11462 & ~w11463;
assign w11466 = ~w11464 & ~w11465;
assign w11467 = ~w11184 & ~w11188;
assign w11468 = pi35 & pi42;
assign w11469 = pi37 & pi40;
assign w11470 = ~w11269 & ~w11469;
assign w11471 = pi37 & pi41;
assign w11472 = w11266 & w11471;
assign w11473 = ~w11470 & ~w11472;
assign w11474 = w11468 & ~w11473;
assign w11475 = ~w11468 & w11473;
assign w11476 = ~w11474 & ~w11475;
assign w11477 = pi14 & pi63;
assign w11478 = pi31 & pi46;
assign w11479 = ~w11477 & ~w11478;
assign w11480 = w11477 & w11478;
assign w11481 = ~w11479 & ~w11480;
assign w11482 = w11259 & ~w11481;
assign w11483 = ~w11259 & w11481;
assign w11484 = ~w11482 & ~w11483;
assign w11485 = ~w11476 & ~w11484;
assign w11486 = w11476 & w11484;
assign w11487 = ~w11485 & ~w11486;
assign w11488 = pi15 & pi62;
assign w11489 = ~pi38 & pi39;
assign w11490 = w11488 & ~w11489;
assign w11491 = ~w11488 & w11489;
assign w11492 = ~w11490 & ~w11491;
assign w11493 = w11487 & ~w11492;
assign w11494 = ~w11487 & w11492;
assign w11495 = ~w11493 & ~w11494;
assign w11496 = ~w11467 & w11495;
assign w11497 = w11467 & ~w11495;
assign w11498 = ~w11496 & ~w11497;
assign w11499 = pi19 & pi58;
assign w11500 = pi20 & pi57;
assign w11501 = pi21 & pi56;
assign w11502 = ~w11500 & ~w11501;
assign w11503 = pi21 & pi57;
assign w11504 = w11153 & w11503;
assign w11505 = ~w11502 & ~w11504;
assign w11506 = w11499 & ~w11505;
assign w11507 = ~w11499 & w11505;
assign w11508 = ~w11506 & ~w11507;
assign w11509 = w11265 & ~w11268;
assign w11510 = ~w11270 & ~w11509;
assign w11511 = ~w11508 & ~w11510;
assign w11512 = w11508 & w11510;
assign w11513 = ~w11511 & ~w11512;
assign w11514 = pi28 & pi49;
assign w11515 = pi29 & pi48;
assign w11516 = ~w11514 & ~w11515;
assign w11517 = pi29 & pi49;
assign w11518 = w11256 & w11517;
assign w11519 = ~w11516 & ~w11518;
assign w11520 = w11312 & ~w11519;
assign w11521 = ~w11312 & w11519;
assign w11522 = ~w11520 & ~w11521;
assign w11523 = w11513 & ~w11522;
assign w11524 = ~w11513 & w11522;
assign w11525 = ~w11523 & ~w11524;
assign w11526 = w11498 & w11525;
assign w11527 = ~w11498 & ~w11525;
assign w11528 = ~w11526 & ~w11527;
assign w11529 = w11466 & w11528;
assign w11530 = ~w11466 & ~w11528;
assign w11531 = ~w11529 & ~w11530;
assign w11532 = w11452 & w11531;
assign w11533 = ~w11452 & ~w11531;
assign w11534 = ~w11532 & ~w11533;
assign w11535 = w11392 & w11534;
assign w11536 = ~w11392 & ~w11534;
assign w11537 = ~w11535 & ~w11536;
assign w11538 = ~w11340 & w11537;
assign w11539 = w11340 & ~w11537;
assign w11540 = ~w11538 & ~w11539;
assign w11541 = ~w11119 & ~w11334;
assign w11542 = (~w7754 & w17831) | (~w7754 & w17832) | (w17831 & w17832);
assign w11543 = w11540 & w11542;
assign w11544 = ~w11540 & ~w11542;
assign w11545 = ~w11543 & ~w11544;
assign w11546 = ~w11333 & ~w11538;
assign w11547 = (w8795 & w17628) | (w8795 & w17629) | (w17628 & w17629);
assign w11548 = ~w11390 & ~w11535;
assign w11549 = ~w11465 & ~w11529;
assign w11550 = ~w11414 & ~w11447;
assign w11551 = (~w11457 & ~w11459) | (~w11457 & w17193) | (~w11459 & w17193);
assign w11552 = pi27 & pi51;
assign w11553 = pi28 & pi50;
assign w11554 = ~w11517 & ~w11553;
assign w11555 = pi29 & pi50;
assign w11556 = w11514 & w11555;
assign w11557 = ~w11554 & ~w11556;
assign w11558 = w11552 & ~w11557;
assign w11559 = ~w11552 & w11557;
assign w11560 = ~w11558 & ~w11559;
assign w11561 = pi19 & pi59;
assign w11562 = ~w11503 & ~w11561;
assign w11563 = w11503 & w11561;
assign w11564 = ~w11562 & ~w11563;
assign w11565 = w11398 & ~w11564;
assign w11566 = ~w11398 & w11564;
assign w11567 = ~w11565 & ~w11566;
assign w11568 = ~w11560 & ~w11567;
assign w11569 = w11560 & w11567;
assign w11570 = ~w11568 & ~w11569;
assign w11571 = pi15 & pi63;
assign w11572 = pi16 & pi62;
assign w11573 = pi17 & pi61;
assign w11574 = ~w11572 & ~w11573;
assign w11575 = pi17 & pi62;
assign w11576 = w11366 & w11575;
assign w11577 = ~w11574 & ~w11576;
assign w11578 = w11571 & ~w11577;
assign w11579 = ~w11571 & w11577;
assign w11580 = ~w11578 & ~w11579;
assign w11581 = w11570 & ~w11580;
assign w11582 = ~w11570 & w11580;
assign w11583 = ~w11581 & ~w11582;
assign w11584 = pi32 & pi46;
assign w11585 = pi34 & pi44;
assign w11586 = ~w11369 & ~w11585;
assign w11587 = pi34 & pi45;
assign w11588 = w11367 & w11587;
assign w11589 = ~w11586 & ~w11588;
assign w11590 = w11584 & ~w11589;
assign w11591 = ~w11584 & w11589;
assign w11592 = ~w11590 & ~w11591;
assign w11593 = pi20 & pi58;
assign w11594 = pi31 & pi47;
assign w11595 = pi30 & pi48;
assign w11596 = ~w11594 & ~w11595;
assign w11597 = pi31 & pi48;
assign w11598 = w11259 & w11597;
assign w11599 = ~w11596 & ~w11598;
assign w11600 = w11593 & ~w11599;
assign w11601 = ~w11593 & w11599;
assign w11602 = ~w11600 & ~w11601;
assign w11603 = ~w11592 & ~w11602;
assign w11604 = w11592 & w11602;
assign w11605 = ~w11603 & ~w11604;
assign w11606 = pi25 & pi53;
assign w11607 = pi22 & pi56;
assign w11608 = ~w11349 & ~w11607;
assign w11609 = w11349 & w11607;
assign w11610 = ~w11608 & ~w11609;
assign w11611 = w11606 & ~w11610;
assign w11612 = ~w11606 & w11610;
assign w11613 = ~w11611 & ~w11612;
assign w11614 = w11605 & ~w11613;
assign w11615 = ~w11605 & w11613;
assign w11616 = ~w11614 & ~w11615;
assign w11617 = w11583 & w11616;
assign w11618 = ~w11583 & ~w11616;
assign w11619 = ~w11617 & ~w11618;
assign w11620 = ~w11551 & w11619;
assign w11621 = w11551 & ~w11619;
assign w11622 = ~w11620 & ~w11621;
assign w11623 = ~w11550 & w11622;
assign w11624 = w11550 & ~w11622;
assign w11625 = ~w11623 & ~w11624;
assign w11626 = w11549 & ~w11625;
assign w11627 = ~w11549 & w11625;
assign w11628 = ~w11626 & ~w11627;
assign w11629 = ~w11450 & ~w11532;
assign w11630 = ~w11628 & w11629;
assign w11631 = w11628 & ~w11629;
assign w11632 = ~w11630 & ~w11631;
assign w11633 = ~w11384 & ~w11387;
assign w11634 = (~w11363 & ~w11365) | (~w11363 & w17833) | (~w11365 & w17833);
assign w11635 = (~w11511 & ~w11513) | (~w11511 & w16942) | (~w11513 & w16942);
assign w11636 = (~w11485 & ~w11487) | (~w11485 & w16943) | (~w11487 & w16943);
assign w11637 = ~w11635 & ~w11636;
assign w11638 = w11635 & w11636;
assign w11639 = ~w11637 & ~w11638;
assign w11640 = w11634 & ~w11639;
assign w11641 = ~w11634 & w11639;
assign w11642 = ~w11640 & ~w11641;
assign w11643 = ~w11442 & ~w11444;
assign w11644 = ~w11642 & w11643;
assign w11645 = w11642 & ~w11643;
assign w11646 = ~w11644 & ~w11645;
assign w11647 = ~pi38 & ~w11488;
assign w11648 = pi39 & ~w11647;
assign w11649 = w11468 & ~w11470;
assign w11650 = ~w11472 & ~w11649;
assign w11651 = w11648 & ~w11650;
assign w11652 = ~w11648 & w11650;
assign w11653 = ~w11651 & ~w11652;
assign w11654 = w11282 & ~w11348;
assign w11655 = ~w11350 & ~w11654;
assign w11656 = ~w11653 & w11655;
assign w11657 = w11653 & ~w11655;
assign w11658 = ~w11656 & ~w11657;
assign w11659 = ~w11259 & ~w11480;
assign w11660 = ~w11479 & ~w11659;
assign w11661 = w11312 & ~w11516;
assign w11662 = ~w11518 & ~w11661;
assign w11663 = w11660 & ~w11662;
assign w11664 = ~w11660 & w11662;
assign w11665 = ~w11663 & ~w11664;
assign w11666 = w11366 & ~w11368;
assign w11667 = ~w11370 & ~w11666;
assign w11668 = ~w11665 & w11667;
assign w11669 = w11665 & ~w11667;
assign w11670 = ~w11668 & ~w11669;
assign w11671 = (~w11432 & ~w11434) | (~w11432 & w17194) | (~w11434 & w17194);
assign w11672 = ~w11670 & w11671;
assign w11673 = w11670 & ~w11671;
assign w11674 = ~w11672 & ~w11673;
assign w11675 = w11658 & w11674;
assign w11676 = ~w11658 & ~w11674;
assign w11677 = ~w11675 & ~w11676;
assign w11678 = w11646 & w11677;
assign w11679 = ~w11646 & ~w11677;
assign w11680 = ~w11678 & ~w11679;
assign w11681 = ~w11633 & w11680;
assign w11682 = w11633 & ~w11680;
assign w11683 = ~w11681 & ~w11682;
assign w11684 = (~w11420 & ~w11422) | (~w11420 & w16773) | (~w11422 & w16773);
assign w11685 = pi23 & pi55;
assign w11686 = pi35 & pi43;
assign w11687 = pi36 & pi42;
assign w11688 = ~w11686 & ~w11687;
assign w11689 = pi36 & pi43;
assign w11690 = w11468 & w11689;
assign w11691 = ~w11688 & ~w11690;
assign w11692 = w11685 & ~w11691;
assign w11693 = ~w11685 & w11691;
assign w11694 = ~w11692 & ~w11693;
assign w11695 = pi38 & pi40;
assign w11696 = pi26 & pi52;
assign w11697 = ~w11695 & ~w11696;
assign w11698 = w11695 & w11696;
assign w11699 = ~w11697 & ~w11698;
assign w11700 = w11471 & ~w11699;
assign w11701 = ~w11471 & w11699;
assign w11702 = ~w11700 & ~w11701;
assign w11703 = ~w11694 & ~w11702;
assign w11704 = w11694 & w11702;
assign w11705 = ~w11703 & ~w11704;
assign w11706 = w11684 & ~w11705;
assign w11707 = ~w11684 & w11705;
assign w11708 = ~w11706 & ~w11707;
assign w11709 = (~w11399 & w11402) | (~w11399 & w16944) | (w11402 & w16944);
assign w11710 = ~w11355 & ~w11358;
assign w11711 = ~w11357 & ~w11710;
assign w11712 = w11499 & ~w11502;
assign w11713 = ~w11504 & ~w11712;
assign w11714 = w11711 & ~w11713;
assign w11715 = ~w11711 & w11713;
assign w11716 = ~w11714 & ~w11715;
assign w11717 = w11709 & ~w11716;
assign w11718 = ~w11709 & w11716;
assign w11719 = ~w11717 & ~w11718;
assign w11720 = (~w11406 & ~w11408) | (~w11406 & w16945) | (~w11408 & w16945);
assign w11721 = ~w11719 & w11720;
assign w11722 = w11719 & ~w11720;
assign w11723 = ~w11721 & ~w11722;
assign w11724 = w11708 & w11723;
assign w11725 = ~w11708 & ~w11723;
assign w11726 = ~w11724 & ~w11725;
assign w11727 = ~w11378 & ~w11381;
assign w11728 = ~w11496 & ~w11526;
assign w11729 = ~w11727 & ~w11728;
assign w11730 = w11727 & w11728;
assign w11731 = ~w11729 & ~w11730;
assign w11732 = w11726 & w11731;
assign w11733 = ~w11726 & ~w11731;
assign w11734 = ~w11732 & ~w11733;
assign w11735 = w11683 & w11734;
assign w11736 = ~w11683 & ~w11734;
assign w11737 = ~w11735 & ~w11736;
assign w11738 = w11632 & w11737;
assign w11739 = ~w11632 & ~w11737;
assign w11740 = ~w11738 & ~w11739;
assign w11741 = ~w11548 & w11740;
assign w11742 = w11548 & ~w11740;
assign w11743 = ~w11741 & ~w11742;
assign w11744 = w11547 & ~w11743;
assign w11745 = ~w11547 & w11743;
assign w11746 = ~w11744 & ~w11745;
assign w11747 = ~w11631 & ~w11738;
assign w11748 = ~w11729 & ~w11732;
assign w11749 = ~w11617 & ~w11620;
assign w11750 = ~w11398 & ~w11563;
assign w11751 = ~w11562 & ~w11750;
assign w11752 = w11552 & ~w11554;
assign w11753 = ~w11556 & ~w11752;
assign w11754 = w11751 & ~w11753;
assign w11755 = ~w11751 & w11753;
assign w11756 = ~w11754 & ~w11755;
assign w11757 = ~w11606 & ~w11609;
assign w11758 = ~w11608 & ~w11757;
assign w11759 = ~w11756 & ~w11758;
assign w11760 = w11756 & w11758;
assign w11761 = ~w11759 & ~w11760;
assign w11762 = ~w11703 & ~w11707;
assign w11763 = ~w11761 & w11762;
assign w11764 = w11761 & ~w11762;
assign w11765 = ~w11763 & ~w11764;
assign w11766 = (~w11714 & ~w11716) | (~w11714 & w16946) | (~w11716 & w16946);
assign w11767 = pi16 & pi63;
assign w11768 = pi35 & pi44;
assign w11769 = ~w11587 & ~w11768;
assign w11770 = pi35 & pi45;
assign w11771 = w11585 & w11770;
assign w11772 = ~w11769 & ~w11771;
assign w11773 = w11767 & ~w11772;
assign w11774 = ~w11767 & w11772;
assign w11775 = ~w11773 & ~w11774;
assign w11776 = pi23 & pi56;
assign w11777 = pi27 & pi52;
assign w11778 = ~w11776 & ~w11777;
assign w11779 = w11776 & w11777;
assign w11780 = ~w11778 & ~w11779;
assign w11781 = w11689 & ~w11780;
assign w11782 = ~w11689 & w11780;
assign w11783 = ~w11781 & ~w11782;
assign w11784 = ~w11775 & ~w11783;
assign w11785 = w11775 & w11783;
assign w11786 = ~w11784 & ~w11785;
assign w11787 = w11766 & ~w11786;
assign w11788 = ~w11766 & w11786;
assign w11789 = ~w11787 & ~w11788;
assign w11790 = w11765 & w11789;
assign w11791 = ~w11765 & ~w11789;
assign w11792 = ~w11790 & ~w11791;
assign w11793 = ~w11749 & w11792;
assign w11794 = w11749 & ~w11792;
assign w11795 = ~w11793 & ~w11794;
assign w11796 = ~w11603 & ~w11614;
assign w11797 = pi18 & pi61;
assign w11798 = ~w11471 & ~w11698;
assign w11799 = ~w11798 & w17195;
assign w11800 = (~w11797 & w11798) | (~w11797 & w17196) | (w11798 & w17196);
assign w11801 = ~w11799 & ~w11800;
assign w11802 = w11685 & ~w11688;
assign w11803 = ~w11690 & ~w11802;
assign w11804 = ~w11801 & w11803;
assign w11805 = w11801 & ~w11803;
assign w11806 = ~w11804 & ~w11805;
assign w11807 = w11571 & ~w11574;
assign w11808 = ~w11576 & ~w11807;
assign w11809 = w11593 & ~w11596;
assign w11810 = ~w11598 & ~w11809;
assign w11811 = ~w11808 & ~w11810;
assign w11812 = w11808 & w11810;
assign w11813 = ~w11811 & ~w11812;
assign w11814 = w11584 & ~w11586;
assign w11815 = ~w11588 & ~w11814;
assign w11816 = ~w11813 & w11815;
assign w11817 = w11813 & ~w11815;
assign w11818 = ~w11816 & ~w11817;
assign w11819 = w11806 & w11818;
assign w11820 = ~w11806 & ~w11818;
assign w11821 = ~w11819 & ~w11820;
assign w11822 = ~w11796 & w11821;
assign w11823 = w11796 & ~w11821;
assign w11824 = ~w11822 & ~w11823;
assign w11825 = w11795 & w11824;
assign w11826 = ~w11795 & ~w11824;
assign w11827 = ~w11825 & ~w11826;
assign w11828 = ~w11748 & w11827;
assign w11829 = w11748 & ~w11827;
assign w11830 = ~w11828 & ~w11829;
assign w11831 = ~w11623 & ~w11627;
assign w11832 = ~w11830 & w11831;
assign w11833 = w11830 & ~w11831;
assign w11834 = ~w11832 & ~w11833;
assign w11835 = ~w11645 & ~w11678;
assign w11836 = (~w11673 & ~w11674) | (~w11673 & w17197) | (~w11674 & w17197);
assign w11837 = pi24 & pi55;
assign w11838 = pi26 & pi53;
assign w11839 = pi25 & pi54;
assign w11840 = ~w11838 & ~w11839;
assign w11841 = pi26 & pi54;
assign w11842 = w11606 & w11841;
assign w11843 = ~w11840 & ~w11842;
assign w11844 = w11837 & ~w11843;
assign w11845 = ~w11837 & w11843;
assign w11846 = ~w11844 & ~w11845;
assign w11847 = pi37 & pi42;
assign w11848 = pi39 & pi40;
assign w11849 = pi38 & pi41;
assign w11850 = ~w11848 & ~w11849;
assign w11851 = pi39 & pi41;
assign w11852 = w11695 & w11851;
assign w11853 = ~w11850 & ~w11852;
assign w11854 = w11847 & ~w11853;
assign w11855 = ~w11847 & w11853;
assign w11856 = ~w11854 & ~w11855;
assign w11857 = ~w11846 & ~w11856;
assign w11858 = w11846 & w11856;
assign w11859 = ~w11857 & ~w11858;
assign w11860 = pi28 & pi51;
assign w11861 = ~pi40 & ~w11575;
assign w11862 = pi62 & w6702;
assign w11863 = ~w11861 & ~w11862;
assign w11864 = w11860 & ~w11863;
assign w11865 = ~w11860 & w11863;
assign w11866 = ~w11864 & ~w11865;
assign w11867 = w11859 & ~w11866;
assign w11868 = ~w11859 & w11866;
assign w11869 = ~w11867 & ~w11868;
assign w11870 = pi19 & pi60;
assign w11871 = pi20 & pi59;
assign w11872 = pi21 & pi58;
assign w11873 = ~w11871 & ~w11872;
assign w11874 = pi21 & pi59;
assign w11875 = w11593 & w11874;
assign w11876 = ~w11873 & ~w11875;
assign w11877 = w11870 & ~w11876;
assign w11878 = ~w11870 & w11876;
assign w11879 = ~w11877 & ~w11878;
assign w11880 = pi22 & pi57;
assign w11881 = pi30 & pi49;
assign w11882 = ~w11555 & ~w11881;
assign w11883 = pi30 & pi50;
assign w11884 = w11517 & w11883;
assign w11885 = ~w11882 & ~w11884;
assign w11886 = w11880 & ~w11885;
assign w11887 = ~w11880 & w11885;
assign w11888 = ~w11886 & ~w11887;
assign w11889 = ~w11879 & ~w11888;
assign w11890 = w11879 & w11888;
assign w11891 = ~w11889 & ~w11890;
assign w11892 = pi33 & pi46;
assign w11893 = pi32 & pi47;
assign w11894 = ~w11892 & ~w11893;
assign w11895 = pi33 & pi47;
assign w11896 = w11584 & w11895;
assign w11897 = ~w11894 & ~w11896;
assign w11898 = w11597 & ~w11897;
assign w11899 = ~w11597 & w11897;
assign w11900 = ~w11898 & ~w11899;
assign w11901 = w11891 & ~w11900;
assign w11902 = ~w11891 & w11900;
assign w11903 = ~w11901 & ~w11902;
assign w11904 = w11869 & w11903;
assign w11905 = ~w11869 & ~w11903;
assign w11906 = ~w11904 & ~w11905;
assign w11907 = ~w11836 & w11906;
assign w11908 = w11836 & ~w11906;
assign w11909 = ~w11907 & ~w11908;
assign w11910 = ~w11835 & w11909;
assign w11911 = w11835 & ~w11909;
assign w11912 = ~w11910 & ~w11911;
assign w11913 = (~w11568 & ~w11570) | (~w11568 & w17198) | (~w11570 & w17198);
assign w11914 = (~w11663 & ~w11665) | (~w11663 & w16947) | (~w11665 & w16947);
assign w11915 = (~w11651 & ~w11653) | (~w11651 & w16948) | (~w11653 & w16948);
assign w11916 = ~w11914 & ~w11915;
assign w11917 = w11914 & w11915;
assign w11918 = ~w11916 & ~w11917;
assign w11919 = w11913 & ~w11918;
assign w11920 = ~w11913 & w11918;
assign w11921 = ~w11919 & ~w11920;
assign w11922 = (~w11637 & ~w11639) | (~w11637 & w17199) | (~w11639 & w17199);
assign w11923 = ~w11921 & w11922;
assign w11924 = w11921 & ~w11922;
assign w11925 = ~w11923 & ~w11924;
assign w11926 = (~w11722 & ~w11723) | (~w11722 & w17200) | (~w11723 & w17200);
assign w11927 = w11925 & ~w11926;
assign w11928 = ~w11925 & w11926;
assign w11929 = ~w11927 & ~w11928;
assign w11930 = w11912 & w11929;
assign w11931 = ~w11912 & ~w11929;
assign w11932 = ~w11930 & ~w11931;
assign w11933 = ~w11681 & ~w11735;
assign w11934 = w11932 & ~w11933;
assign w11935 = ~w11932 & w11933;
assign w11936 = ~w11934 & ~w11935;
assign w11937 = w11834 & w11936;
assign w11938 = ~w11834 & ~w11936;
assign w11939 = ~w11937 & ~w11938;
assign w11940 = ~w11747 & w11939;
assign w11941 = w11747 & ~w11939;
assign w11942 = ~w11940 & ~w11941;
assign w11943 = (w7754 & w17834) | (w7754 & w17835) | (w17834 & w17835);
assign w11944 = w11942 & w11943;
assign w11945 = ~w11942 & ~w11943;
assign w11946 = ~w11944 & ~w11945;
assign w11947 = ~w11742 & ~w11941;
assign w11948 = (~w7754 & w17836) | (~w7754 & w17837) | (w17836 & w17837);
assign w11949 = ~w11934 & ~w11937;
assign w11950 = ~w11828 & ~w11833;
assign w11951 = (~w11793 & ~w11795) | (~w11793 & w17838) | (~w11795 & w17838);
assign w11952 = pi19 & pi61;
assign w11953 = pi18 & pi62;
assign w11954 = ~w11952 & ~w11953;
assign w11955 = pi19 & pi62;
assign w11956 = w11797 & w11955;
assign w11957 = ~w11954 & ~w11956;
assign w11958 = ~w11860 & ~w11862;
assign w11959 = ~w11861 & ~w11958;
assign w11960 = w11957 & w11959;
assign w11961 = ~w11957 & ~w11959;
assign w11962 = ~w11960 & ~w11961;
assign w11963 = pi34 & pi46;
assign w11964 = pi36 & pi44;
assign w11965 = ~w11770 & ~w11964;
assign w11966 = pi36 & pi45;
assign w11967 = w11768 & w11966;
assign w11968 = ~w11965 & ~w11967;
assign w11969 = w11963 & ~w11968;
assign w11970 = ~w11963 & w11968;
assign w11971 = ~w11969 & ~w11970;
assign w11972 = pi17 & pi63;
assign w11973 = pi29 & pi51;
assign w11974 = ~w11972 & ~w11973;
assign w11975 = w11972 & w11973;
assign w11976 = ~w11974 & ~w11975;
assign w11977 = w11895 & ~w11976;
assign w11978 = ~w11895 & w11976;
assign w11979 = ~w11977 & ~w11978;
assign w11980 = ~w11971 & ~w11979;
assign w11981 = w11971 & w11979;
assign w11982 = ~w11980 & ~w11981;
assign w11983 = w11962 & w11982;
assign w11984 = ~w11962 & ~w11982;
assign w11985 = ~w11983 & ~w11984;
assign w11986 = pi20 & pi60;
assign w11987 = pi22 & pi58;
assign w11988 = ~w11874 & ~w11987;
assign w11989 = pi22 & pi59;
assign w11990 = w11872 & w11989;
assign w11991 = ~w11988 & ~w11990;
assign w11992 = w11986 & ~w11991;
assign w11993 = ~w11986 & w11991;
assign w11994 = ~w11992 & ~w11993;
assign w11995 = w11847 & ~w11850;
assign w11996 = ~w11852 & ~w11995;
assign w11997 = ~w11994 & ~w11996;
assign w11998 = w11994 & w11996;
assign w11999 = ~w11997 & ~w11998;
assign w12000 = pi31 & pi49;
assign w12001 = pi32 & pi48;
assign w12002 = ~w12000 & ~w12001;
assign w12003 = pi32 & pi49;
assign w12004 = w11597 & w12003;
assign w12005 = ~w12002 & ~w12004;
assign w12006 = w11883 & ~w12005;
assign w12007 = ~w11883 & w12005;
assign w12008 = ~w12006 & ~w12007;
assign w12009 = ~w11999 & w12008;
assign w12010 = w11999 & ~w12008;
assign w12011 = ~w12009 & ~w12010;
assign w12012 = pi25 & pi55;
assign w12013 = pi38 & pi42;
assign w12014 = pi37 & pi43;
assign w12015 = ~w12013 & ~w12014;
assign w12016 = pi38 & pi43;
assign w12017 = w11847 & w12016;
assign w12018 = ~w12015 & ~w12017;
assign w12019 = w12012 & ~w12018;
assign w12020 = ~w12012 & w12018;
assign w12021 = ~w12019 & ~w12020;
assign w12022 = pi23 & pi57;
assign w12023 = pi24 & pi56;
assign w12024 = ~w11841 & ~w12023;
assign w12025 = w11841 & w12023;
assign w12026 = ~w12024 & ~w12025;
assign w12027 = w12022 & ~w12026;
assign w12028 = ~w12022 & w12026;
assign w12029 = ~w12027 & ~w12028;
assign w12030 = ~w12021 & ~w12029;
assign w12031 = w12021 & w12029;
assign w12032 = ~w12030 & ~w12031;
assign w12033 = pi28 & pi52;
assign w12034 = pi27 & pi53;
assign w12035 = ~w12033 & ~w12034;
assign w12036 = pi28 & pi53;
assign w12037 = w11777 & w12036;
assign w12038 = ~w12035 & ~w12037;
assign w12039 = w11851 & ~w12038;
assign w12040 = ~w11851 & w12038;
assign w12041 = ~w12039 & ~w12040;
assign w12042 = w12032 & ~w12041;
assign w12043 = ~w12032 & w12041;
assign w12044 = ~w12042 & ~w12043;
assign w12045 = w12011 & w12044;
assign w12046 = ~w12011 & ~w12044;
assign w12047 = ~w12045 & ~w12046;
assign w12048 = w11985 & w12047;
assign w12049 = ~w11985 & ~w12047;
assign w12050 = ~w12048 & ~w12049;
assign w12051 = (w12050 & w11927) | (w12050 & w17839) | (w11927 & w17839);
assign w12052 = ~w11927 & w17840;
assign w12053 = ~w12051 & ~w12052;
assign w12054 = ~w11951 & w12053;
assign w12055 = w11951 & ~w12053;
assign w12056 = ~w12054 & ~w12055;
assign w12057 = ~w11950 & w12056;
assign w12058 = w11950 & ~w12056;
assign w12059 = ~w12057 & ~w12058;
assign w12060 = ~w11910 & ~w11930;
assign w12061 = ~w11904 & ~w11907;
assign w12062 = w11767 & ~w11769;
assign w12063 = ~w11771 & ~w12062;
assign w12064 = w11837 & ~w11840;
assign w12065 = ~w11842 & ~w12064;
assign w12066 = ~w12063 & ~w12065;
assign w12067 = w12063 & w12065;
assign w12068 = ~w12066 & ~w12067;
assign w12069 = ~w11689 & ~w11779;
assign w12070 = ~w11778 & ~w12069;
assign w12071 = ~w12068 & ~w12070;
assign w12072 = w12068 & w12070;
assign w12073 = ~w12071 & ~w12072;
assign w12074 = ~w11784 & ~w11788;
assign w12075 = ~w12073 & w12074;
assign w12076 = w12073 & ~w12074;
assign w12077 = ~w12075 & ~w12076;
assign w12078 = (~w11916 & ~w11918) | (~w11916 & w17201) | (~w11918 & w17201);
assign w12079 = ~w12077 & w12078;
assign w12080 = w12077 & ~w12078;
assign w12081 = ~w12079 & ~w12080;
assign w12082 = ~w12061 & w12081;
assign w12083 = w12061 & ~w12081;
assign w12084 = ~w12082 & ~w12083;
assign w12085 = w11870 & ~w11873;
assign w12086 = ~w11875 & ~w12085;
assign w12087 = w11880 & ~w11882;
assign w12088 = ~w11884 & ~w12087;
assign w12089 = ~w12086 & ~w12088;
assign w12090 = w12086 & w12088;
assign w12091 = ~w12089 & ~w12090;
assign w12092 = w11597 & ~w11894;
assign w12093 = ~w11896 & ~w12092;
assign w12094 = ~w12091 & w12093;
assign w12095 = w12091 & ~w12093;
assign w12096 = ~w12094 & ~w12095;
assign w12097 = (~w11857 & ~w11859) | (~w11857 & w17202) | (~w11859 & w17202);
assign w12098 = (~w11889 & ~w11891) | (~w11889 & w17203) | (~w11891 & w17203);
assign w12099 = ~w12097 & ~w12098;
assign w12100 = w12097 & w12098;
assign w12101 = ~w12099 & ~w12100;
assign w12102 = w12096 & w12101;
assign w12103 = ~w12096 & ~w12101;
assign w12104 = ~w12102 & ~w12103;
assign w12105 = w12084 & w12104;
assign w12106 = ~w12084 & ~w12104;
assign w12107 = ~w12105 & ~w12106;
assign w12108 = ~w11799 & ~w11805;
assign w12109 = (~w11754 & ~w11756) | (~w11754 & w17204) | (~w11756 & w17204);
assign w12110 = (~w11811 & ~w11813) | (~w11811 & w17205) | (~w11813 & w17205);
assign w12111 = ~w12109 & ~w12110;
assign w12112 = w12109 & w12110;
assign w12113 = ~w12111 & ~w12112;
assign w12114 = w12108 & ~w12113;
assign w12115 = ~w12108 & w12113;
assign w12116 = ~w12114 & ~w12115;
assign w12117 = (~w11764 & ~w11765) | (~w11764 & w16949) | (~w11765 & w16949);
assign w12118 = (~w11819 & ~w11821) | (~w11819 & w17206) | (~w11821 & w17206);
assign w12119 = ~w12117 & ~w12118;
assign w12120 = w12117 & w12118;
assign w12121 = ~w12119 & ~w12120;
assign w12122 = ~w12116 & ~w12121;
assign w12123 = w12116 & w12121;
assign w12124 = ~w12122 & ~w12123;
assign w12125 = w12107 & w12124;
assign w12126 = ~w12107 & ~w12124;
assign w12127 = ~w12125 & ~w12126;
assign w12128 = ~w12060 & w12127;
assign w12129 = w12060 & ~w12127;
assign w12130 = ~w12128 & ~w12129;
assign w12131 = w12059 & w12130;
assign w12132 = ~w12059 & ~w12130;
assign w12133 = ~w12131 & ~w12132;
assign w12134 = ~w11949 & w12133;
assign w12135 = w11949 & ~w12133;
assign w12136 = ~w12134 & ~w12135;
assign w12137 = w11948 & w12136;
assign w12138 = ~w11948 & ~w12136;
assign w12139 = ~w12137 & ~w12138;
assign w12140 = ~w11940 & ~w12134;
assign w12141 = (w8795 & w17630) | (w8795 & w17631) | (w17630 & w17631);
assign w12142 = ~w12057 & ~w12131;
assign w12143 = ~w12051 & ~w12054;
assign w12144 = ~w12066 & ~w12072;
assign w12145 = ~w12089 & ~w12095;
assign w12146 = pi27 & pi54;
assign w12147 = pi39 & pi42;
assign w12148 = ~w12016 & ~w12147;
assign w12149 = pi39 & pi43;
assign w12150 = w12013 & w12149;
assign w12151 = ~w12148 & ~w12150;
assign w12152 = w12146 & ~w12151;
assign w12153 = ~w12146 & w12151;
assign w12154 = ~w12152 & ~w12153;
assign w12155 = ~w12145 & ~w12154;
assign w12156 = w12145 & w12154;
assign w12157 = ~w12155 & ~w12156;
assign w12158 = w12144 & ~w12157;
assign w12159 = ~w12144 & w12157;
assign w12160 = ~w12158 & ~w12159;
assign w12161 = (~w12076 & ~w12077) | (~w12076 & w17207) | (~w12077 & w17207);
assign w12162 = ~w12099 & ~w12102;
assign w12163 = ~w12161 & ~w12162;
assign w12164 = w12161 & w12162;
assign w12165 = ~w12163 & ~w12164;
assign w12166 = w12160 & w12165;
assign w12167 = ~w12160 & ~w12165;
assign w12168 = ~w12166 & ~w12167;
assign w12169 = ~w12143 & w12168;
assign w12170 = w12143 & ~w12168;
assign w12171 = ~w12169 & ~w12170;
assign w12172 = w12012 & ~w12015;
assign w12173 = ~w12017 & ~w12172;
assign w12174 = w11851 & ~w12035;
assign w12175 = ~w12037 & ~w12174;
assign w12176 = ~w12173 & ~w12175;
assign w12177 = w12173 & w12175;
assign w12178 = ~w12176 & ~w12177;
assign w12179 = ~w12022 & ~w12025;
assign w12180 = ~w12024 & ~w12179;
assign w12181 = ~w12178 & ~w12180;
assign w12182 = w12178 & w12180;
assign w12183 = ~w12181 & ~w12182;
assign w12184 = (~w12030 & ~w12032) | (~w12030 & w17841) | (~w12032 & w17841);
assign w12185 = (~w11997 & ~w11999) | (~w11997 & w17842) | (~w11999 & w17842);
assign w12186 = ~w12184 & ~w12185;
assign w12187 = w12184 & w12185;
assign w12188 = ~w12186 & ~w12187;
assign w12189 = w12183 & w12188;
assign w12190 = ~w12183 & ~w12188;
assign w12191 = ~w12189 & ~w12190;
assign w12192 = ~w11956 & ~w11960;
assign w12193 = w11963 & ~w11965;
assign w12194 = ~w11967 & ~w12193;
assign w12195 = ~w12192 & ~w12194;
assign w12196 = w12192 & w12194;
assign w12197 = ~w12195 & ~w12196;
assign w12198 = pi30 & pi51;
assign w12199 = pi31 & pi50;
assign w12200 = ~w12003 & ~w12199;
assign w12201 = pi32 & pi50;
assign w12202 = w12000 & w12201;
assign w12203 = ~w12200 & ~w12202;
assign w12204 = w12198 & ~w12203;
assign w12205 = ~w12198 & w12203;
assign w12206 = ~w12204 & ~w12205;
assign w12207 = ~w12197 & w12206;
assign w12208 = w12197 & ~w12206;
assign w12209 = ~w12207 & ~w12208;
assign w12210 = ~w11895 & ~w11975;
assign w12211 = ~w11974 & ~w12210;
assign w12212 = w11883 & ~w12002;
assign w12213 = ~w12004 & ~w12212;
assign w12214 = w12211 & ~w12213;
assign w12215 = ~w12211 & w12213;
assign w12216 = ~w12214 & ~w12215;
assign w12217 = w11986 & ~w11988;
assign w12218 = ~w11990 & ~w12217;
assign w12219 = ~w12216 & w12218;
assign w12220 = w12216 & ~w12218;
assign w12221 = ~w12219 & ~w12220;
assign w12222 = (~w11980 & ~w11982) | (~w11980 & w17843) | (~w11982 & w17843);
assign w12223 = ~w12221 & w12222;
assign w12224 = w12221 & ~w12222;
assign w12225 = ~w12223 & ~w12224;
assign w12226 = w12209 & w12225;
assign w12227 = ~w12209 & ~w12225;
assign w12228 = ~w12226 & ~w12227;
assign w12229 = ~w12045 & ~w12048;
assign w12230 = w12228 & ~w12229;
assign w12231 = ~w12228 & w12229;
assign w12232 = ~w12230 & ~w12231;
assign w12233 = w12191 & w12232;
assign w12234 = ~w12191 & ~w12232;
assign w12235 = ~w12233 & ~w12234;
assign w12236 = w12171 & w12235;
assign w12237 = ~w12171 & ~w12235;
assign w12238 = ~w12236 & ~w12237;
assign w12239 = ~w12125 & ~w12128;
assign w12240 = (~w12082 & ~w12084) | (~w12082 & w17844) | (~w12084 & w17844);
assign w12241 = (~w12119 & ~w12121) | (~w12119 & w17208) | (~w12121 & w17208);
assign w12242 = (~w12111 & ~w12113) | (~w12111 & w17845) | (~w12113 & w17845);
assign w12243 = ~pi40 & pi41;
assign w12244 = w11955 & ~w12243;
assign w12245 = ~w11955 & w12243;
assign w12246 = ~w12244 & ~w12245;
assign w12247 = pi25 & pi56;
assign w12248 = pi23 & pi58;
assign w12249 = ~w12247 & ~w12248;
assign w12250 = w12247 & w12248;
assign w12251 = ~w12249 & ~w12250;
assign w12252 = w11989 & ~w12251;
assign w12253 = ~w11989 & w12251;
assign w12254 = ~w12252 & ~w12253;
assign w12255 = ~w12246 & ~w12254;
assign w12256 = w12246 & w12254;
assign w12257 = ~w12255 & ~w12256;
assign w12258 = pi24 & pi57;
assign w12259 = pi33 & pi48;
assign w12260 = pi34 & pi47;
assign w12261 = ~w12259 & ~w12260;
assign w12262 = pi34 & pi48;
assign w12263 = w11895 & w12262;
assign w12264 = ~w12261 & ~w12263;
assign w12265 = w12258 & ~w12264;
assign w12266 = ~w12258 & w12264;
assign w12267 = ~w12265 & ~w12266;
assign w12268 = w12257 & ~w12267;
assign w12269 = ~w12257 & w12267;
assign w12270 = ~w12268 & ~w12269;
assign w12271 = ~w12242 & w12270;
assign w12272 = w12242 & ~w12270;
assign w12273 = ~w12271 & ~w12272;
assign w12274 = pi18 & pi63;
assign w12275 = pi20 & pi61;
assign w12276 = pi21 & pi60;
assign w12277 = ~w12275 & ~w12276;
assign w12278 = pi21 & pi61;
assign w12279 = w11986 & w12278;
assign w12280 = ~w12277 & ~w12279;
assign w12281 = w12274 & ~w12280;
assign w12282 = ~w12274 & w12280;
assign w12283 = ~w12281 & ~w12282;
assign w12284 = pi35 & pi46;
assign w12285 = pi37 & pi44;
assign w12286 = ~w11966 & ~w12285;
assign w12287 = pi37 & pi45;
assign w12288 = w11964 & w12287;
assign w12289 = ~w12286 & ~w12288;
assign w12290 = w12284 & ~w12289;
assign w12291 = ~w12284 & w12289;
assign w12292 = ~w12290 & ~w12291;
assign w12293 = ~w12283 & ~w12292;
assign w12294 = w12283 & w12292;
assign w12295 = ~w12293 & ~w12294;
assign w12296 = pi26 & pi55;
assign w12297 = pi29 & pi52;
assign w12298 = ~w12036 & ~w12297;
assign w12299 = pi29 & pi53;
assign w12300 = w12033 & w12299;
assign w12301 = ~w12298 & ~w12300;
assign w12302 = w12296 & ~w12301;
assign w12303 = ~w12296 & w12301;
assign w12304 = ~w12302 & ~w12303;
assign w12305 = w12295 & ~w12304;
assign w12306 = ~w12295 & w12304;
assign w12307 = ~w12305 & ~w12306;
assign w12308 = ~w12273 & ~w12307;
assign w12309 = w12273 & w12307;
assign w12310 = ~w12308 & ~w12309;
assign w12311 = ~w12241 & w12310;
assign w12312 = w12241 & ~w12310;
assign w12313 = ~w12311 & ~w12312;
assign w12314 = ~w12240 & w12313;
assign w12315 = w12240 & ~w12313;
assign w12316 = ~w12314 & ~w12315;
assign w12317 = ~w12239 & w12316;
assign w12318 = w12239 & ~w12316;
assign w12319 = ~w12317 & ~w12318;
assign w12320 = w12238 & w12319;
assign w12321 = ~w12238 & ~w12319;
assign w12322 = ~w12320 & ~w12321;
assign w12323 = w12142 & ~w12322;
assign w12324 = ~w12142 & w12322;
assign w12325 = ~w12323 & ~w12324;
assign w12326 = w12141 & ~w12325;
assign w12327 = ~w12141 & w12325;
assign w12328 = ~w12326 & ~w12327;
assign w12329 = (~w7754 & w17846) | (~w7754 & w17847) | (w17846 & w17847);
assign w12330 = ~w12317 & ~w12320;
assign w12331 = (~w12311 & ~w12313) | (~w12311 & w17848) | (~w12313 & w17848);
assign w12332 = ~w12176 & ~w12182;
assign w12333 = ~w12214 & ~w12220;
assign w12334 = pi28 & pi54;
assign w12335 = pi27 & pi55;
assign w12336 = pi25 & pi57;
assign w12337 = ~w12335 & ~w12336;
assign w12338 = w12335 & w12336;
assign w12339 = ~w12337 & ~w12338;
assign w12340 = w12334 & ~w12339;
assign w12341 = ~w12334 & w12339;
assign w12342 = ~w12340 & ~w12341;
assign w12343 = ~w12333 & ~w12342;
assign w12344 = w12333 & w12342;
assign w12345 = ~w12343 & ~w12344;
assign w12346 = w12332 & ~w12345;
assign w12347 = ~w12332 & w12345;
assign w12348 = ~w12346 & ~w12347;
assign w12349 = ~w12224 & ~w12226;
assign w12350 = ~w12186 & ~w12189;
assign w12351 = ~w12349 & ~w12350;
assign w12352 = w12349 & w12350;
assign w12353 = ~w12351 & ~w12352;
assign w12354 = w12348 & w12353;
assign w12355 = ~w12348 & ~w12353;
assign w12356 = ~w12354 & ~w12355;
assign w12357 = ~w12331 & w12356;
assign w12358 = w12331 & ~w12356;
assign w12359 = ~w12357 & ~w12358;
assign w12360 = ~w12271 & ~w12309;
assign w12361 = w12198 & ~w12200;
assign w12362 = ~w12202 & ~w12361;
assign w12363 = w12258 & ~w12261;
assign w12364 = ~w12263 & ~w12363;
assign w12365 = ~w12362 & ~w12364;
assign w12366 = w12362 & w12364;
assign w12367 = ~w12365 & ~w12366;
assign w12368 = w12296 & ~w12298;
assign w12369 = ~w12300 & ~w12368;
assign w12370 = ~w12367 & w12369;
assign w12371 = w12367 & ~w12369;
assign w12372 = ~w12370 & ~w12371;
assign w12373 = ~w11989 & ~w12250;
assign w12374 = ~w12249 & ~w12373;
assign w12375 = w12274 & ~w12277;
assign w12376 = ~w12279 & ~w12375;
assign w12377 = w12374 & ~w12376;
assign w12378 = ~w12374 & w12376;
assign w12379 = ~w12377 & ~w12378;
assign w12380 = w12284 & ~w12286;
assign w12381 = ~w12288 & ~w12380;
assign w12382 = ~w12379 & w12381;
assign w12383 = w12379 & ~w12381;
assign w12384 = ~w12382 & ~w12383;
assign w12385 = ~w12293 & ~w12305;
assign w12386 = ~w12384 & w12385;
assign w12387 = w12384 & ~w12385;
assign w12388 = ~w12386 & ~w12387;
assign w12389 = w12372 & w12388;
assign w12390 = ~w12372 & ~w12388;
assign w12391 = ~w12389 & ~w12390;
assign w12392 = ~w12360 & w12391;
assign w12393 = w12360 & ~w12391;
assign w12394 = ~w12392 & ~w12393;
assign w12395 = ~w12195 & ~w12208;
assign w12396 = ~w12255 & ~w12268;
assign w12397 = ~w12395 & ~w12396;
assign w12398 = w12395 & w12396;
assign w12399 = ~w12397 & ~w12398;
assign w12400 = pi19 & pi63;
assign w12401 = ~pi40 & ~w11955;
assign w12402 = pi41 & ~w12401;
assign w12403 = ~w12400 & ~w12402;
assign w12404 = w12400 & w12402;
assign w12405 = ~w12403 & ~w12404;
assign w12406 = w12146 & ~w12148;
assign w12407 = ~w12150 & ~w12406;
assign w12408 = w12405 & ~w12407;
assign w12409 = ~w12405 & w12407;
assign w12410 = ~w12408 & ~w12409;
assign w12411 = w12399 & w12410;
assign w12412 = ~w12399 & ~w12410;
assign w12413 = ~w12411 & ~w12412;
assign w12414 = w12394 & w12413;
assign w12415 = ~w12394 & ~w12413;
assign w12416 = ~w12414 & ~w12415;
assign w12417 = w12359 & w12416;
assign w12418 = ~w12359 & ~w12416;
assign w12419 = ~w12417 & ~w12418;
assign w12420 = ~w12169 & ~w12236;
assign w12421 = ~w12230 & ~w12233;
assign w12422 = ~w12163 & ~w12166;
assign w12423 = ~w12155 & ~w12159;
assign w12424 = pi33 & pi49;
assign w12425 = ~w12262 & ~w12424;
assign w12426 = pi34 & pi49;
assign w12427 = w12259 & w12426;
assign w12428 = ~w12425 & ~w12427;
assign w12429 = w12201 & ~w12428;
assign w12430 = ~w12201 & w12428;
assign w12431 = ~w12429 & ~w12430;
assign w12432 = pi20 & pi62;
assign w12433 = pi31 & pi51;
assign w12434 = ~w12278 & ~w12433;
assign w12435 = w12278 & w12433;
assign w12436 = ~w12434 & ~w12435;
assign w12437 = w12432 & ~w12436;
assign w12438 = ~w12432 & w12436;
assign w12439 = ~w12437 & ~w12438;
assign w12440 = ~w12431 & ~w12439;
assign w12441 = w12431 & w12439;
assign w12442 = ~w12440 & ~w12441;
assign w12443 = pi22 & pi60;
assign w12444 = pi24 & pi58;
assign w12445 = pi23 & pi59;
assign w12446 = ~w12444 & ~w12445;
assign w12447 = pi24 & pi59;
assign w12448 = w12248 & w12447;
assign w12449 = ~w12446 & ~w12448;
assign w12450 = w12443 & ~w12449;
assign w12451 = ~w12443 & w12449;
assign w12452 = ~w12450 & ~w12451;
assign w12453 = w12442 & ~w12452;
assign w12454 = ~w12442 & w12452;
assign w12455 = ~w12453 & ~w12454;
assign w12456 = ~w12423 & w12455;
assign w12457 = w12423 & ~w12455;
assign w12458 = ~w12456 & ~w12457;
assign w12459 = pi40 & pi42;
assign w12460 = pi30 & pi52;
assign w12461 = ~w12299 & ~w12460;
assign w12462 = pi30 & pi53;
assign w12463 = w12297 & w12462;
assign w12464 = ~w12461 & ~w12463;
assign w12465 = w12459 & ~w12464;
assign w12466 = ~w12459 & w12464;
assign w12467 = ~w12465 & ~w12466;
assign w12468 = pi26 & pi56;
assign w12469 = pi38 & pi44;
assign w12470 = ~w12149 & ~w12469;
assign w12471 = pi39 & pi44;
assign w12472 = w12016 & w12471;
assign w12473 = ~w12470 & ~w12472;
assign w12474 = w12468 & ~w12473;
assign w12475 = ~w12468 & w12473;
assign w12476 = ~w12474 & ~w12475;
assign w12477 = ~w12467 & ~w12476;
assign w12478 = w12467 & w12476;
assign w12479 = ~w12477 & ~w12478;
assign w12480 = pi35 & pi47;
assign w12481 = pi36 & pi46;
assign w12482 = ~w12287 & ~w12481;
assign w12483 = pi37 & pi46;
assign w12484 = w11966 & w12483;
assign w12485 = ~w12482 & ~w12484;
assign w12486 = w12480 & ~w12485;
assign w12487 = ~w12480 & w12485;
assign w12488 = ~w12486 & ~w12487;
assign w12489 = w12479 & ~w12488;
assign w12490 = ~w12479 & w12488;
assign w12491 = ~w12489 & ~w12490;
assign w12492 = ~w12458 & ~w12491;
assign w12493 = w12458 & w12491;
assign w12494 = ~w12492 & ~w12493;
assign w12495 = ~w12422 & w12494;
assign w12496 = w12422 & ~w12494;
assign w12497 = ~w12495 & ~w12496;
assign w12498 = ~w12421 & w12497;
assign w12499 = w12421 & ~w12497;
assign w12500 = ~w12498 & ~w12499;
assign w12501 = ~w12420 & w12500;
assign w12502 = w12420 & ~w12500;
assign w12503 = ~w12501 & ~w12502;
assign w12504 = w12419 & w12503;
assign w12505 = ~w12419 & ~w12503;
assign w12506 = ~w12504 & ~w12505;
assign w12507 = ~w12330 & w12506;
assign w12508 = w12330 & ~w12506;
assign w12509 = ~w12507 & ~w12508;
assign w12510 = (~w10008 & w17849) | (~w10008 & w17850) | (w17849 & w17850);
assign w12511 = (w10008 & w17851) | (w10008 & w17852) | (w17851 & w17852);
assign w12512 = ~w12510 & ~w12511;
assign w12513 = ~w12501 & ~w12504;
assign w12514 = ~w12357 & ~w12417;
assign w12515 = ~w12392 & ~w12414;
assign w12516 = ~w12351 & ~w12354;
assign w12517 = ~w12343 & ~w12347;
assign w12518 = pi29 & pi54;
assign w12519 = pi40 & pi43;
assign w12520 = ~w12471 & ~w12519;
assign w12521 = pi40 & pi44;
assign w12522 = w12149 & w12521;
assign w12523 = ~w12520 & ~w12522;
assign w12524 = w12518 & ~w12523;
assign w12525 = ~w12518 & w12523;
assign w12526 = ~w12524 & ~w12525;
assign w12527 = pi21 & pi62;
assign w12528 = ~pi41 & pi42;
assign w12529 = w12527 & ~w12528;
assign w12530 = ~w12527 & w12528;
assign w12531 = ~w12529 & ~w12530;
assign w12532 = ~w12526 & ~w12531;
assign w12533 = w12526 & w12531;
assign w12534 = ~w12532 & ~w12533;
assign w12535 = pi33 & pi50;
assign w12536 = pi35 & pi48;
assign w12537 = ~w12426 & ~w12536;
assign w12538 = pi35 & pi49;
assign w12539 = w12262 & w12538;
assign w12540 = ~w12537 & ~w12539;
assign w12541 = w12535 & ~w12540;
assign w12542 = ~w12535 & w12540;
assign w12543 = ~w12541 & ~w12542;
assign w12544 = w12534 & ~w12543;
assign w12545 = ~w12534 & w12543;
assign w12546 = ~w12544 & ~w12545;
assign w12547 = ~w12517 & w12546;
assign w12548 = w12517 & ~w12546;
assign w12549 = ~w12547 & ~w12548;
assign w12550 = pi36 & pi47;
assign w12551 = pi38 & pi45;
assign w12552 = ~w12483 & ~w12551;
assign w12553 = pi38 & pi46;
assign w12554 = w12287 & w12553;
assign w12555 = ~w12552 & ~w12554;
assign w12556 = w12550 & ~w12555;
assign w12557 = ~w12550 & w12555;
assign w12558 = ~w12556 & ~w12557;
assign w12559 = pi25 & pi58;
assign w12560 = pi26 & pi57;
assign w12561 = pi32 & pi51;
assign w12562 = ~w12560 & ~w12561;
assign w12563 = w12560 & w12561;
assign w12564 = ~w12562 & ~w12563;
assign w12565 = w12559 & ~w12564;
assign w12566 = ~w12559 & w12564;
assign w12567 = ~w12565 & ~w12566;
assign w12568 = ~w12558 & ~w12567;
assign w12569 = w12558 & w12567;
assign w12570 = ~w12568 & ~w12569;
assign w12571 = pi27 & pi56;
assign w12572 = pi20 & pi63;
assign w12573 = pi22 & pi61;
assign w12574 = ~w12572 & ~w12573;
assign w12575 = w12572 & w12573;
assign w12576 = ~w12574 & ~w12575;
assign w12577 = w12571 & ~w12576;
assign w12578 = ~w12571 & w12576;
assign w12579 = ~w12577 & ~w12578;
assign w12580 = w12570 & ~w12579;
assign w12581 = ~w12570 & w12579;
assign w12582 = ~w12580 & ~w12581;
assign w12583 = ~w12549 & ~w12582;
assign w12584 = w12549 & w12582;
assign w12585 = ~w12583 & ~w12584;
assign w12586 = ~w12516 & w12585;
assign w12587 = w12516 & ~w12585;
assign w12588 = ~w12586 & ~w12587;
assign w12589 = ~w12515 & w12588;
assign w12590 = w12515 & ~w12588;
assign w12591 = ~w12589 & ~w12590;
assign w12592 = ~w12514 & w12591;
assign w12593 = w12514 & ~w12591;
assign w12594 = ~w12592 & ~w12593;
assign w12595 = w12443 & ~w12446;
assign w12596 = ~w12448 & ~w12595;
assign w12597 = w12480 & ~w12482;
assign w12598 = ~w12484 & ~w12597;
assign w12599 = ~w12596 & ~w12598;
assign w12600 = w12596 & w12598;
assign w12601 = ~w12599 & ~w12600;
assign w12602 = w12468 & ~w12470;
assign w12603 = ~w12472 & ~w12602;
assign w12604 = ~w12601 & w12603;
assign w12605 = w12601 & ~w12603;
assign w12606 = ~w12604 & ~w12605;
assign w12607 = ~w12432 & ~w12435;
assign w12608 = ~w12434 & ~w12607;
assign w12609 = w12201 & ~w12425;
assign w12610 = ~w12427 & ~w12609;
assign w12611 = w12608 & ~w12610;
assign w12612 = ~w12608 & w12610;
assign w12613 = ~w12611 & ~w12612;
assign w12614 = ~w12334 & ~w12338;
assign w12615 = ~w12337 & ~w12614;
assign w12616 = ~w12613 & ~w12615;
assign w12617 = w12613 & w12615;
assign w12618 = ~w12616 & ~w12617;
assign w12619 = ~w12477 & ~w12489;
assign w12620 = ~w12618 & w12619;
assign w12621 = w12618 & ~w12619;
assign w12622 = ~w12620 & ~w12621;
assign w12623 = w12606 & w12622;
assign w12624 = ~w12606 & ~w12622;
assign w12625 = ~w12623 & ~w12624;
assign w12626 = ~w12456 & ~w12493;
assign w12627 = ~w12387 & ~w12389;
assign w12628 = ~w12626 & ~w12627;
assign w12629 = w12626 & w12627;
assign w12630 = ~w12628 & ~w12629;
assign w12631 = w12625 & w12630;
assign w12632 = ~w12625 & ~w12630;
assign w12633 = ~w12631 & ~w12632;
assign w12634 = ~w12495 & ~w12498;
assign w12635 = ~w12440 & ~w12453;
assign w12636 = ~w12365 & ~w12371;
assign w12637 = ~w12377 & ~w12383;
assign w12638 = ~w12636 & ~w12637;
assign w12639 = w12636 & w12637;
assign w12640 = ~w12638 & ~w12639;
assign w12641 = w12635 & ~w12640;
assign w12642 = ~w12635 & w12640;
assign w12643 = ~w12641 & ~w12642;
assign w12644 = pi23 & pi60;
assign w12645 = ~w12447 & ~w12644;
assign w12646 = pi24 & pi60;
assign w12647 = w12445 & w12646;
assign w12648 = ~w12645 & ~w12647;
assign w12649 = w12459 & ~w12461;
assign w12650 = ~w12463 & ~w12649;
assign w12651 = w12648 & ~w12650;
assign w12652 = ~w12648 & w12650;
assign w12653 = ~w12651 & ~w12652;
assign w12654 = pi31 & pi52;
assign w12655 = pi28 & pi55;
assign w12656 = ~w12462 & ~w12655;
assign w12657 = w12462 & w12655;
assign w12658 = ~w12656 & ~w12657;
assign w12659 = w12654 & ~w12658;
assign w12660 = ~w12654 & w12658;
assign w12661 = ~w12659 & ~w12660;
assign w12662 = w12653 & ~w12661;
assign w12663 = ~w12653 & w12661;
assign w12664 = ~w12662 & ~w12663;
assign w12665 = ~w12404 & ~w12408;
assign w12666 = ~w12664 & w12665;
assign w12667 = w12664 & ~w12665;
assign w12668 = ~w12666 & ~w12667;
assign w12669 = ~w12397 & ~w12411;
assign w12670 = ~w12668 & w12669;
assign w12671 = w12668 & ~w12669;
assign w12672 = ~w12670 & ~w12671;
assign w12673 = w12643 & w12672;
assign w12674 = ~w12643 & ~w12672;
assign w12675 = ~w12673 & ~w12674;
assign w12676 = ~w12634 & w12675;
assign w12677 = w12634 & ~w12675;
assign w12678 = ~w12676 & ~w12677;
assign w12679 = w12633 & w12678;
assign w12680 = ~w12633 & ~w12678;
assign w12681 = ~w12679 & ~w12680;
assign w12682 = ~w12594 & ~w12681;
assign w12683 = w12594 & w12681;
assign w12684 = ~w12682 & ~w12683;
assign w12685 = ~w12513 & w12684;
assign w12686 = w12513 & ~w12684;
assign w12687 = ~w12685 & ~w12686;
assign w12688 = ~w12323 & ~w12508;
assign w12689 = (~w8795 & w17632) | (~w8795 & w17633) | (w17632 & w17633);
assign w12690 = w12687 & w12689;
assign w12691 = ~w12687 & ~w12689;
assign w12692 = ~w12690 & ~w12691;
assign w12693 = ~w12507 & ~w12685;
assign w12694 = ~w12592 & ~w12683;
assign w12695 = ~w12676 & ~w12679;
assign w12696 = ~w12638 & ~w12642;
assign w12697 = (~w12647 & w12650) | (~w12647 & w16774) | (w12650 & w16774);
assign w12698 = ~w12571 & ~w12575;
assign w12699 = ~w12574 & ~w12698;
assign w12700 = ~w12697 & w12699;
assign w12701 = w12697 & ~w12699;
assign w12702 = ~w12700 & ~w12701;
assign w12703 = pi26 & pi58;
assign w12704 = pi31 & pi53;
assign w12705 = pi32 & pi52;
assign w12706 = ~w12704 & ~w12705;
assign w12707 = pi32 & pi53;
assign w12708 = w12654 & w12707;
assign w12709 = ~w12706 & ~w12708;
assign w12710 = w12703 & ~w12709;
assign w12711 = ~w12703 & w12709;
assign w12712 = ~w12710 & ~w12711;
assign w12713 = ~w12702 & w12712;
assign w12714 = w12702 & ~w12712;
assign w12715 = ~w12713 & ~w12714;
assign w12716 = ~w12662 & ~w12667;
assign w12717 = w12715 & ~w12716;
assign w12718 = ~w12715 & w12716;
assign w12719 = ~w12717 & ~w12718;
assign w12720 = w12696 & ~w12719;
assign w12721 = ~w12696 & w12719;
assign w12722 = ~w12720 & ~w12721;
assign w12723 = ~w12671 & ~w12673;
assign w12724 = ~w12722 & w12723;
assign w12725 = w12722 & ~w12723;
assign w12726 = ~w12724 & ~w12725;
assign w12727 = w12535 & ~w12537;
assign w12728 = ~w12539 & ~w12727;
assign w12729 = w12550 & ~w12552;
assign w12730 = ~w12554 & ~w12729;
assign w12731 = ~w12728 & ~w12730;
assign w12732 = w12728 & w12730;
assign w12733 = ~w12731 & ~w12732;
assign w12734 = ~w12559 & ~w12563;
assign w12735 = ~w12562 & ~w12734;
assign w12736 = ~w12733 & ~w12735;
assign w12737 = w12733 & w12735;
assign w12738 = ~w12736 & ~w12737;
assign w12739 = (~w12599 & ~w12601) | (~w12599 & w16775) | (~w12601 & w16775);
assign w12740 = (~w12611 & ~w12613) | (~w12611 & w16776) | (~w12613 & w16776);
assign w12741 = ~w12739 & ~w12740;
assign w12742 = w12739 & w12740;
assign w12743 = ~w12741 & ~w12742;
assign w12744 = w12738 & w12743;
assign w12745 = ~w12738 & ~w12743;
assign w12746 = ~w12744 & ~w12745;
assign w12747 = pi21 & pi63;
assign w12748 = pi22 & pi62;
assign w12749 = pi23 & pi61;
assign w12750 = ~w12748 & ~w12749;
assign w12751 = pi23 & pi62;
assign w12752 = w12573 & w12751;
assign w12753 = ~w12750 & ~w12752;
assign w12754 = w12747 & ~w12753;
assign w12755 = ~w12747 & w12753;
assign w12756 = ~w12754 & ~w12755;
assign w12757 = pi33 & pi51;
assign w12758 = pi25 & pi59;
assign w12759 = ~w12646 & ~w12758;
assign w12760 = pi25 & pi60;
assign w12761 = w12447 & w12760;
assign w12762 = ~w12759 & ~w12761;
assign w12763 = w12757 & ~w12762;
assign w12764 = ~w12757 & w12762;
assign w12765 = ~w12763 & ~w12764;
assign w12766 = ~w12756 & ~w12765;
assign w12767 = w12756 & w12765;
assign w12768 = ~w12766 & ~w12767;
assign w12769 = pi34 & pi50;
assign w12770 = pi36 & pi48;
assign w12771 = ~w12538 & ~w12770;
assign w12772 = pi36 & pi49;
assign w12773 = w12536 & w12772;
assign w12774 = ~w12771 & ~w12773;
assign w12775 = w12769 & ~w12774;
assign w12776 = ~w12769 & w12774;
assign w12777 = ~w12775 & ~w12776;
assign w12778 = w12768 & ~w12777;
assign w12779 = ~w12768 & w12777;
assign w12780 = ~w12778 & ~w12779;
assign w12781 = pi39 & pi45;
assign w12782 = pi41 & pi43;
assign w12783 = ~w12521 & ~w12782;
assign w12784 = pi41 & pi44;
assign w12785 = w12519 & w12784;
assign w12786 = ~w12783 & ~w12785;
assign w12787 = w12781 & ~w12786;
assign w12788 = ~w12781 & w12786;
assign w12789 = ~w12787 & ~w12788;
assign w12790 = pi28 & pi56;
assign w12791 = pi29 & pi55;
assign w12792 = ~w12553 & ~w12791;
assign w12793 = w12553 & w12791;
assign w12794 = ~w12792 & ~w12793;
assign w12795 = w12790 & ~w12794;
assign w12796 = ~w12790 & w12794;
assign w12797 = ~w12795 & ~w12796;
assign w12798 = ~w12789 & ~w12797;
assign w12799 = w12789 & w12797;
assign w12800 = ~w12798 & ~w12799;
assign w12801 = pi37 & pi47;
assign w12802 = pi27 & pi57;
assign w12803 = pi30 & pi54;
assign w12804 = ~w12802 & ~w12803;
assign w12805 = w12802 & w12803;
assign w12806 = ~w12804 & ~w12805;
assign w12807 = w12801 & ~w12806;
assign w12808 = ~w12801 & w12806;
assign w12809 = ~w12807 & ~w12808;
assign w12810 = w12800 & ~w12809;
assign w12811 = ~w12800 & w12809;
assign w12812 = ~w12810 & ~w12811;
assign w12813 = w12780 & w12812;
assign w12814 = ~w12780 & ~w12812;
assign w12815 = ~w12813 & ~w12814;
assign w12816 = w12746 & w12815;
assign w12817 = ~w12746 & ~w12815;
assign w12818 = ~w12816 & ~w12817;
assign w12819 = w12726 & w12818;
assign w12820 = ~w12726 & ~w12818;
assign w12821 = ~w12819 & ~w12820;
assign w12822 = ~w12695 & w12821;
assign w12823 = w12695 & ~w12821;
assign w12824 = ~w12822 & ~w12823;
assign w12825 = ~pi41 & ~w12527;
assign w12826 = pi42 & ~w12825;
assign w12827 = w12518 & ~w12520;
assign w12828 = ~w12522 & ~w12827;
assign w12829 = w12826 & ~w12828;
assign w12830 = ~w12826 & w12828;
assign w12831 = ~w12829 & ~w12830;
assign w12832 = ~w12654 & ~w12657;
assign w12833 = ~w12656 & ~w12832;
assign w12834 = ~w12831 & ~w12833;
assign w12835 = w12831 & w12833;
assign w12836 = ~w12834 & ~w12835;
assign w12837 = (~w12568 & ~w12570) | (~w12568 & w16950) | (~w12570 & w16950);
assign w12838 = (~w12532 & ~w12534) | (~w12532 & w16951) | (~w12534 & w16951);
assign w12839 = ~w12837 & ~w12838;
assign w12840 = w12837 & w12838;
assign w12841 = ~w12839 & ~w12840;
assign w12842 = w12836 & w12841;
assign w12843 = ~w12836 & ~w12841;
assign w12844 = ~w12842 & ~w12843;
assign w12845 = ~w12547 & ~w12584;
assign w12846 = ~w12621 & ~w12623;
assign w12847 = ~w12845 & ~w12846;
assign w12848 = w12845 & w12846;
assign w12849 = ~w12847 & ~w12848;
assign w12850 = w12844 & w12849;
assign w12851 = ~w12844 & ~w12849;
assign w12852 = ~w12850 & ~w12851;
assign w12853 = ~w12586 & ~w12589;
assign w12854 = ~w12628 & ~w12631;
assign w12855 = ~w12853 & ~w12854;
assign w12856 = w12853 & w12854;
assign w12857 = ~w12855 & ~w12856;
assign w12858 = w12852 & w12857;
assign w12859 = ~w12852 & ~w12857;
assign w12860 = ~w12858 & ~w12859;
assign w12861 = w12824 & w12860;
assign w12862 = ~w12824 & ~w12860;
assign w12863 = ~w12861 & ~w12862;
assign w12864 = w12694 & ~w12863;
assign w12865 = ~w12694 & w12863;
assign w12866 = ~w12864 & ~w12865;
assign w12867 = (~w10008 & w17853) | (~w10008 & w17854) | (w17853 & w17854);
assign w12868 = (w10008 & w17855) | (w10008 & w17856) | (w17855 & w17856);
assign w12869 = ~w12867 & ~w12868;
assign w12870 = (w8795 & w17634) | (w8795 & w17635) | (w17634 & w17635);
assign w12871 = ~w12822 & ~w12861;
assign w12872 = ~w12847 & ~w12850;
assign w12873 = (~w12700 & ~w12702) | (~w12700 & w16952) | (~w12702 & w16952);
assign w12874 = (~w12731 & ~w12733) | (~w12731 & w16777) | (~w12733 & w16777);
assign w12875 = (~w12829 & ~w12831) | (~w12829 & w16778) | (~w12831 & w16778);
assign w12876 = ~w12874 & ~w12875;
assign w12877 = w12874 & w12875;
assign w12878 = ~w12876 & ~w12877;
assign w12879 = w12873 & ~w12878;
assign w12880 = ~w12873 & w12878;
assign w12881 = ~w12879 & ~w12880;
assign w12882 = ~w12717 & ~w12721;
assign w12883 = ~w12881 & w12882;
assign w12884 = w12881 & ~w12882;
assign w12885 = ~w12883 & ~w12884;
assign w12886 = ~w12813 & ~w12816;
assign w12887 = w12885 & ~w12886;
assign w12888 = ~w12885 & w12886;
assign w12889 = ~w12887 & ~w12888;
assign w12890 = ~w12872 & w12889;
assign w12891 = w12872 & ~w12889;
assign w12892 = ~w12890 & ~w12891;
assign w12893 = ~w12725 & ~w12819;
assign w12894 = w12892 & ~w12893;
assign w12895 = ~w12892 & w12893;
assign w12896 = ~w12894 & ~w12895;
assign w12897 = ~w12855 & ~w12858;
assign w12898 = w12747 & ~w12750;
assign w12899 = ~w12752 & ~w12898;
assign w12900 = w12769 & ~w12771;
assign w12901 = ~w12773 & ~w12900;
assign w12902 = ~w12899 & ~w12901;
assign w12903 = w12899 & w12901;
assign w12904 = ~w12902 & ~w12903;
assign w12905 = w12757 & ~w12759;
assign w12906 = ~w12761 & ~w12905;
assign w12907 = ~w12904 & w12906;
assign w12908 = w12904 & ~w12906;
assign w12909 = ~w12907 & ~w12908;
assign w12910 = (~w12798 & ~w12800) | (~w12798 & w16953) | (~w12800 & w16953);
assign w12911 = (~w12766 & ~w12768) | (~w12766 & w16954) | (~w12768 & w16954);
assign w12912 = ~w12910 & ~w12911;
assign w12913 = w12910 & w12911;
assign w12914 = ~w12912 & ~w12913;
assign w12915 = w12909 & w12914;
assign w12916 = ~w12909 & ~w12914;
assign w12917 = ~w12915 & ~w12916;
assign w12918 = (~w12741 & ~w12743) | (~w12741 & w16955) | (~w12743 & w16955);
assign w12919 = pi24 & pi61;
assign w12920 = w12781 & ~w12783;
assign w12921 = (w12919 & w12920) | (w12919 & w16779) | (w12920 & w16779);
assign w12922 = ~w12920 & w16780;
assign w12923 = ~w12921 & ~w12922;
assign w12924 = ~w12790 & ~w12793;
assign w12925 = ~w12792 & ~w12924;
assign w12926 = ~w12923 & ~w12925;
assign w12927 = w12923 & w12925;
assign w12928 = ~w12926 & ~w12927;
assign w12929 = ~w12801 & ~w12805;
assign w12930 = ~w12804 & ~w12929;
assign w12931 = w12703 & ~w12706;
assign w12932 = ~w12708 & ~w12931;
assign w12933 = w12930 & ~w12932;
assign w12934 = ~w12930 & w12932;
assign w12935 = ~w12933 & ~w12934;
assign w12936 = pi26 & pi59;
assign w12937 = pi27 & pi58;
assign w12938 = ~w12936 & ~w12937;
assign w12939 = pi27 & pi59;
assign w12940 = w12703 & w12939;
assign w12941 = ~w12938 & ~w12940;
assign w12942 = w12760 & ~w12941;
assign w12943 = ~w12760 & w12941;
assign w12944 = ~w12942 & ~w12943;
assign w12945 = ~w12935 & w12944;
assign w12946 = w12935 & ~w12944;
assign w12947 = ~w12945 & ~w12946;
assign w12948 = ~w12928 & ~w12947;
assign w12949 = w12928 & w12947;
assign w12950 = ~w12948 & ~w12949;
assign w12951 = w12918 & ~w12950;
assign w12952 = ~w12918 & w12950;
assign w12953 = ~w12951 & ~w12952;
assign w12954 = w12917 & w12953;
assign w12955 = ~w12917 & ~w12953;
assign w12956 = ~w12954 & ~w12955;
assign w12957 = (~w12839 & ~w12841) | (~w12839 & w17209) | (~w12841 & w17209);
assign w12958 = pi33 & pi52;
assign w12959 = pi34 & pi51;
assign w12960 = ~w12958 & ~w12959;
assign w12961 = pi34 & pi52;
assign w12962 = w12757 & w12961;
assign w12963 = ~w12960 & ~w12962;
assign w12964 = w12707 & ~w12963;
assign w12965 = ~w12707 & w12963;
assign w12966 = ~w12964 & ~w12965;
assign w12967 = pi35 & pi50;
assign w12968 = pi28 & pi57;
assign w12969 = pi22 & pi63;
assign w12970 = ~w12968 & ~w12969;
assign w12971 = w12968 & w12969;
assign w12972 = ~w12970 & ~w12971;
assign w12973 = w12967 & ~w12972;
assign w12974 = ~w12967 & w12972;
assign w12975 = ~w12973 & ~w12974;
assign w12976 = ~w12966 & ~w12975;
assign w12977 = w12966 & w12975;
assign w12978 = ~w12976 & ~w12977;
assign w12979 = pi39 & pi46;
assign w12980 = pi40 & pi45;
assign w12981 = ~w12784 & ~w12980;
assign w12982 = pi41 & pi45;
assign w12983 = w12521 & w12982;
assign w12984 = ~w12981 & ~w12983;
assign w12985 = w12979 & ~w12984;
assign w12986 = ~w12979 & w12984;
assign w12987 = ~w12985 & ~w12986;
assign w12988 = w12978 & ~w12987;
assign w12989 = ~w12978 & w12987;
assign w12990 = ~w12988 & ~w12989;
assign w12991 = pi37 & pi48;
assign w12992 = pi38 & pi47;
assign w12993 = ~w12991 & ~w12992;
assign w12994 = pi38 & pi48;
assign w12995 = w12801 & w12994;
assign w12996 = ~w12993 & ~w12995;
assign w12997 = w12772 & ~w12996;
assign w12998 = ~w12772 & w12996;
assign w12999 = ~w12997 & ~w12998;
assign w13000 = ~pi42 & pi43;
assign w13001 = w12751 & ~w13000;
assign w13002 = ~w12751 & w13000;
assign w13003 = ~w13001 & ~w13002;
assign w13004 = ~w12999 & ~w13003;
assign w13005 = w12999 & w13003;
assign w13006 = ~w13004 & ~w13005;
assign w13007 = pi29 & pi56;
assign w13008 = pi30 & pi55;
assign w13009 = pi31 & pi54;
assign w13010 = ~w13008 & ~w13009;
assign w13011 = pi31 & pi55;
assign w13012 = w12803 & w13011;
assign w13013 = ~w13010 & ~w13012;
assign w13014 = w13007 & ~w13013;
assign w13015 = ~w13007 & w13013;
assign w13016 = ~w13014 & ~w13015;
assign w13017 = w13006 & ~w13016;
assign w13018 = ~w13006 & w13016;
assign w13019 = ~w13017 & ~w13018;
assign w13020 = w12990 & w13019;
assign w13021 = ~w12990 & ~w13019;
assign w13022 = ~w13020 & ~w13021;
assign w13023 = ~w12957 & w13022;
assign w13024 = w12957 & ~w13022;
assign w13025 = ~w13023 & ~w13024;
assign w13026 = ~w12956 & ~w13025;
assign w13027 = w12956 & w13025;
assign w13028 = ~w13026 & ~w13027;
assign w13029 = ~w12897 & w13028;
assign w13030 = w12897 & ~w13028;
assign w13031 = ~w13029 & ~w13030;
assign w13032 = w12896 & w13031;
assign w13033 = ~w12896 & ~w13031;
assign w13034 = ~w13032 & ~w13033;
assign w13035 = ~w12871 & w13034;
assign w13036 = w12871 & ~w13034;
assign w13037 = ~w13035 & ~w13036;
assign w13038 = w12870 & w13037;
assign w13039 = ~w12870 & ~w13037;
assign w13040 = ~w13038 & ~w13039;
assign w13041 = ~w12864 & ~w13036;
assign w13042 = (~w8795 & w17636) | (~w8795 & w17637) | (w17636 & w17637);
assign w13043 = ~w13029 & ~w13032;
assign w13044 = (~w12902 & ~w12904) | (~w12902 & w17210) | (~w12904 & w17210);
assign w13045 = (~w12921 & ~w12923) | (~w12921 & w16956) | (~w12923 & w16956);
assign w13046 = pi25 & pi61;
assign w13047 = pi24 & pi62;
assign w13048 = ~w13046 & ~w13047;
assign w13049 = pi25 & pi62;
assign w13050 = w12919 & w13049;
assign w13051 = ~w13048 & ~w13050;
assign w13052 = (pi43 & w12751) | (pi43 & w16957) | (w12751 & w16957);
assign w13053 = w13051 & w13052;
assign w13054 = ~w13051 & ~w13052;
assign w13055 = ~w13053 & ~w13054;
assign w13056 = ~w13045 & w13055;
assign w13057 = w13045 & ~w13055;
assign w13058 = ~w13056 & ~w13057;
assign w13059 = w13044 & ~w13058;
assign w13060 = ~w13044 & w13058;
assign w13061 = ~w13059 & ~w13060;
assign w13062 = (w13061 & w12952) | (w13061 & w17211) | (w12952 & w17211);
assign w13063 = ~w12952 & w17212;
assign w13064 = ~w13062 & ~w13063;
assign w13065 = ~w13020 & ~w13023;
assign w13066 = w13064 & ~w13065;
assign w13067 = ~w13064 & w13065;
assign w13068 = ~w13066 & ~w13067;
assign w13069 = ~w12954 & ~w13027;
assign w13070 = ~w12884 & ~w12887;
assign w13071 = ~w13069 & ~w13070;
assign w13072 = w13069 & w13070;
assign w13073 = ~w13071 & ~w13072;
assign w13074 = w13068 & w13073;
assign w13075 = ~w13068 & ~w13073;
assign w13076 = ~w13074 & ~w13075;
assign w13077 = ~w12890 & ~w12894;
assign w13078 = (~w12912 & ~w12914) | (~w12912 & w17213) | (~w12914 & w17213);
assign w13079 = pi23 & pi63;
assign w13080 = pi36 & pi50;
assign w13081 = pi37 & pi49;
assign w13082 = ~w13080 & ~w13081;
assign w13083 = pi37 & pi50;
assign w13084 = w12772 & w13083;
assign w13085 = ~w13082 & ~w13084;
assign w13086 = w13079 & ~w13085;
assign w13087 = ~w13079 & w13085;
assign w13088 = ~w13086 & ~w13087;
assign w13089 = pi33 & pi53;
assign w13090 = pi35 & pi51;
assign w13091 = ~w12961 & ~w13090;
assign w13092 = pi35 & pi52;
assign w13093 = w12959 & w13092;
assign w13094 = ~w13091 & ~w13093;
assign w13095 = w13089 & ~w13094;
assign w13096 = ~w13089 & w13094;
assign w13097 = ~w13095 & ~w13096;
assign w13098 = ~w13088 & ~w13097;
assign w13099 = w13088 & w13097;
assign w13100 = ~w13098 & ~w13099;
assign w13101 = pi29 & pi57;
assign w13102 = ~w13011 & ~w13101;
assign w13103 = w13011 & w13101;
assign w13104 = ~w13102 & ~w13103;
assign w13105 = w12994 & ~w13104;
assign w13106 = ~w12994 & w13104;
assign w13107 = ~w13105 & ~w13106;
assign w13108 = w13100 & ~w13107;
assign w13109 = ~w13100 & w13107;
assign w13110 = ~w13108 & ~w13109;
assign w13111 = pi26 & pi60;
assign w13112 = pi28 & pi58;
assign w13113 = ~w12939 & ~w13112;
assign w13114 = pi28 & pi59;
assign w13115 = w12937 & w13114;
assign w13116 = ~w13113 & ~w13115;
assign w13117 = w13111 & ~w13116;
assign w13118 = ~w13111 & w13116;
assign w13119 = ~w13117 & ~w13118;
assign w13120 = pi42 & pi44;
assign w13121 = pi32 & pi54;
assign w13122 = ~w13120 & ~w13121;
assign w13123 = w13120 & w13121;
assign w13124 = ~w13122 & ~w13123;
assign w13125 = w12982 & ~w13124;
assign w13126 = ~w12982 & w13124;
assign w13127 = ~w13125 & ~w13126;
assign w13128 = ~w13119 & ~w13127;
assign w13129 = w13119 & w13127;
assign w13130 = ~w13128 & ~w13129;
assign w13131 = pi30 & pi56;
assign w13132 = pi40 & pi46;
assign w13133 = pi39 & pi47;
assign w13134 = ~w13132 & ~w13133;
assign w13135 = pi40 & pi47;
assign w13136 = w12979 & w13135;
assign w13137 = ~w13134 & ~w13136;
assign w13138 = w13131 & ~w13137;
assign w13139 = ~w13131 & w13137;
assign w13140 = ~w13138 & ~w13139;
assign w13141 = w13130 & ~w13140;
assign w13142 = ~w13130 & w13140;
assign w13143 = ~w13141 & ~w13142;
assign w13144 = w13110 & w13143;
assign w13145 = ~w13110 & ~w13143;
assign w13146 = ~w13144 & ~w13145;
assign w13147 = ~w13078 & w13146;
assign w13148 = w13078 & ~w13146;
assign w13149 = ~w13147 & ~w13148;
assign w13150 = ~w13004 & ~w13017;
assign w13151 = (~w12933 & ~w12935) | (~w12933 & w17214) | (~w12935 & w17214);
assign w13152 = (~w12976 & ~w12978) | (~w12976 & w16958) | (~w12978 & w16958);
assign w13153 = ~w13151 & ~w13152;
assign w13154 = w13151 & w13152;
assign w13155 = ~w13153 & ~w13154;
assign w13156 = w13150 & ~w13155;
assign w13157 = ~w13150 & w13155;
assign w13158 = ~w13156 & ~w13157;
assign w13159 = (~w12876 & ~w12878) | (~w12876 & w16959) | (~w12878 & w16959);
assign w13160 = w12979 & ~w12981;
assign w13161 = ~w12983 & ~w13160;
assign w13162 = w13007 & ~w13010;
assign w13163 = ~w13012 & ~w13162;
assign w13164 = ~w13161 & ~w13163;
assign w13165 = w13161 & w13163;
assign w13166 = ~w13164 & ~w13165;
assign w13167 = w12772 & ~w12993;
assign w13168 = ~w12995 & ~w13167;
assign w13169 = ~w13166 & w13168;
assign w13170 = w13166 & ~w13168;
assign w13171 = ~w13169 & ~w13170;
assign w13172 = w12760 & ~w12938;
assign w13173 = ~w12940 & ~w13172;
assign w13174 = w12707 & ~w12960;
assign w13175 = ~w12962 & ~w13174;
assign w13176 = ~w13173 & ~w13175;
assign w13177 = w13173 & w13175;
assign w13178 = ~w13176 & ~w13177;
assign w13179 = ~w12967 & ~w12971;
assign w13180 = ~w12970 & ~w13179;
assign w13181 = ~w13178 & ~w13180;
assign w13182 = w13178 & w13180;
assign w13183 = ~w13181 & ~w13182;
assign w13184 = w13171 & w13183;
assign w13185 = ~w13171 & ~w13183;
assign w13186 = ~w13184 & ~w13185;
assign w13187 = ~w13159 & w13186;
assign w13188 = w13159 & ~w13186;
assign w13189 = ~w13187 & ~w13188;
assign w13190 = w13158 & w13189;
assign w13191 = ~w13158 & ~w13189;
assign w13192 = ~w13190 & ~w13191;
assign w13193 = w13149 & w13192;
assign w13194 = ~w13149 & ~w13192;
assign w13195 = ~w13193 & ~w13194;
assign w13196 = ~w13077 & w13195;
assign w13197 = w13077 & ~w13195;
assign w13198 = ~w13196 & ~w13197;
assign w13199 = w13076 & w13198;
assign w13200 = ~w13076 & ~w13198;
assign w13201 = ~w13199 & ~w13200;
assign w13202 = ~w13043 & w13201;
assign w13203 = w13043 & ~w13201;
assign w13204 = ~w13202 & ~w13203;
assign w13205 = w13042 & w13204;
assign w13206 = ~w13042 & ~w13204;
assign w13207 = ~w13205 & ~w13206;
assign w13208 = ~w13035 & ~w13202;
assign w13209 = ~w13196 & ~w13199;
assign w13210 = ~w13144 & ~w13147;
assign w13211 = ~w13128 & ~w13141;
assign w13212 = (~w13164 & ~w13166) | (~w13164 & w17215) | (~w13166 & w17215);
assign w13213 = (~w13098 & ~w13100) | (~w13098 & w16960) | (~w13100 & w16960);
assign w13214 = ~w13212 & ~w13213;
assign w13215 = w13212 & w13213;
assign w13216 = ~w13214 & ~w13215;
assign w13217 = w13211 & ~w13216;
assign w13218 = ~w13211 & w13216;
assign w13219 = ~w13217 & ~w13218;
assign w13220 = ~w13210 & w13219;
assign w13221 = w13210 & ~w13219;
assign w13222 = ~w13220 & ~w13221;
assign w13223 = ~w13062 & ~w13066;
assign w13224 = ~w13222 & w13223;
assign w13225 = w13222 & ~w13223;
assign w13226 = ~w13224 & ~w13225;
assign w13227 = ~w13071 & ~w13074;
assign w13228 = ~w13226 & w13227;
assign w13229 = w13226 & ~w13227;
assign w13230 = ~w13228 & ~w13229;
assign w13231 = ~w13190 & ~w13193;
assign w13232 = (~w13176 & ~w13178) | (~w13176 & w17216) | (~w13178 & w17216);
assign w13233 = ~pi43 & pi44;
assign w13234 = w13049 & ~w13233;
assign w13235 = ~w13049 & w13233;
assign w13236 = ~w13234 & ~w13235;
assign w13237 = pi31 & pi56;
assign w13238 = pi33 & pi54;
assign w13239 = ~w13237 & ~w13238;
assign w13240 = w13237 & w13238;
assign w13241 = ~w13239 & ~w13240;
assign w13242 = w13135 & ~w13241;
assign w13243 = ~w13135 & w13241;
assign w13244 = ~w13242 & ~w13243;
assign w13245 = ~w13236 & ~w13244;
assign w13246 = w13236 & w13244;
assign w13247 = ~w13245 & ~w13246;
assign w13248 = w13232 & ~w13247;
assign w13249 = ~w13232 & w13247;
assign w13250 = ~w13248 & ~w13249;
assign w13251 = pi24 & pi63;
assign w13252 = pi26 & pi61;
assign w13253 = pi27 & pi60;
assign w13254 = ~w13252 & ~w13253;
assign w13255 = pi27 & pi61;
assign w13256 = w13111 & w13255;
assign w13257 = ~w13254 & ~w13256;
assign w13258 = w13251 & ~w13257;
assign w13259 = ~w13251 & w13257;
assign w13260 = ~w13258 & ~w13259;
assign w13261 = pi38 & pi49;
assign w13262 = pi39 & pi48;
assign w13263 = ~w13261 & ~w13262;
assign w13264 = pi39 & pi49;
assign w13265 = w12994 & w13264;
assign w13266 = ~w13263 & ~w13265;
assign w13267 = w13083 & ~w13266;
assign w13268 = ~w13083 & w13266;
assign w13269 = ~w13267 & ~w13268;
assign w13270 = ~w13260 & ~w13269;
assign w13271 = w13260 & w13269;
assign w13272 = ~w13270 & ~w13271;
assign w13273 = pi32 & pi55;
assign w13274 = pi41 & pi46;
assign w13275 = pi42 & pi45;
assign w13276 = ~w13274 & ~w13275;
assign w13277 = pi42 & pi46;
assign w13278 = w12982 & w13277;
assign w13279 = ~w13276 & ~w13278;
assign w13280 = w13273 & ~w13279;
assign w13281 = ~w13273 & w13279;
assign w13282 = ~w13280 & ~w13281;
assign w13283 = w13272 & ~w13282;
assign w13284 = ~w13272 & w13282;
assign w13285 = ~w13283 & ~w13284;
assign w13286 = ~w13250 & ~w13285;
assign w13287 = w13250 & w13285;
assign w13288 = ~w13286 & ~w13287;
assign w13289 = (~w13050 & ~w13051) | (~w13050 & w16961) | (~w13051 & w16961);
assign w13290 = pi30 & pi57;
assign w13291 = pi34 & pi53;
assign w13292 = ~w13290 & ~w13291;
assign w13293 = w13290 & w13291;
assign w13294 = ~w13292 & ~w13293;
assign w13295 = w13114 & ~w13294;
assign w13296 = ~w13114 & w13294;
assign w13297 = ~w13295 & ~w13296;
assign w13298 = ~w13289 & ~w13297;
assign w13299 = w13289 & w13297;
assign w13300 = ~w13298 & ~w13299;
assign w13301 = pi29 & pi58;
assign w13302 = pi36 & pi51;
assign w13303 = ~w13301 & ~w13302;
assign w13304 = w13301 & w13302;
assign w13305 = ~w13303 & ~w13304;
assign w13306 = w13092 & ~w13305;
assign w13307 = ~w13092 & w13305;
assign w13308 = ~w13306 & ~w13307;
assign w13309 = w13300 & ~w13308;
assign w13310 = ~w13300 & w13308;
assign w13311 = ~w13309 & ~w13310;
assign w13312 = w13288 & w13311;
assign w13313 = ~w13288 & ~w13311;
assign w13314 = ~w13312 & ~w13313;
assign w13315 = ~w13231 & w13314;
assign w13316 = w13231 & ~w13314;
assign w13317 = ~w13315 & ~w13316;
assign w13318 = (~w13056 & ~w13058) | (~w13056 & w17217) | (~w13058 & w17217);
assign w13319 = ~w12982 & ~w13123;
assign w13320 = ~w13122 & ~w13319;
assign w13321 = w13131 & ~w13134;
assign w13322 = ~w13136 & ~w13321;
assign w13323 = w13320 & ~w13322;
assign w13324 = ~w13320 & w13322;
assign w13325 = ~w13323 & ~w13324;
assign w13326 = ~w12994 & ~w13103;
assign w13327 = ~w13102 & ~w13326;
assign w13328 = ~w13325 & ~w13327;
assign w13329 = w13325 & w13327;
assign w13330 = ~w13328 & ~w13329;
assign w13331 = w13089 & ~w13091;
assign w13332 = ~w13093 & ~w13331;
assign w13333 = w13111 & ~w13113;
assign w13334 = ~w13115 & ~w13333;
assign w13335 = ~w13332 & ~w13334;
assign w13336 = w13332 & w13334;
assign w13337 = ~w13335 & ~w13336;
assign w13338 = w13079 & ~w13082;
assign w13339 = ~w13084 & ~w13338;
assign w13340 = ~w13337 & w13339;
assign w13341 = w13337 & ~w13339;
assign w13342 = ~w13340 & ~w13341;
assign w13343 = w13330 & w13342;
assign w13344 = ~w13330 & ~w13342;
assign w13345 = ~w13343 & ~w13344;
assign w13346 = ~w13318 & w13345;
assign w13347 = w13318 & ~w13345;
assign w13348 = ~w13346 & ~w13347;
assign w13349 = ~w13184 & ~w13187;
assign w13350 = (~w13153 & ~w13155) | (~w13153 & w17218) | (~w13155 & w17218);
assign w13351 = ~w13349 & ~w13350;
assign w13352 = w13349 & w13350;
assign w13353 = ~w13351 & ~w13352;
assign w13354 = w13348 & w13353;
assign w13355 = ~w13348 & ~w13353;
assign w13356 = ~w13354 & ~w13355;
assign w13357 = w13317 & w13356;
assign w13358 = ~w13317 & ~w13356;
assign w13359 = ~w13357 & ~w13358;
assign w13360 = ~w13230 & ~w13359;
assign w13361 = w13230 & w13359;
assign w13362 = ~w13360 & ~w13361;
assign w13363 = w13209 & ~w13362;
assign w13364 = ~w13209 & w13362;
assign w13365 = ~w13363 & ~w13364;
assign w13366 = (~w10008 & w17857) | (~w10008 & w17858) | (w17857 & w17858);
assign w13367 = (w10008 & w17859) | (w10008 & w17860) | (w17859 & w17860);
assign w13368 = ~w13366 & ~w13367;
assign w13369 = ~w13229 & ~w13361;
assign w13370 = ~w13315 & ~w13357;
assign w13371 = (~w13351 & ~w13353) | (~w13351 & w17219) | (~w13353 & w17219);
assign w13372 = ~w13270 & ~w13283;
assign w13373 = (~w13335 & ~w13337) | (~w13335 & w17220) | (~w13337 & w17220);
assign w13374 = (~w13298 & ~w13300) | (~w13298 & w16962) | (~w13300 & w16962);
assign w13375 = ~w13373 & ~w13374;
assign w13376 = w13373 & w13374;
assign w13377 = ~w13375 & ~w13376;
assign w13378 = w13372 & ~w13377;
assign w13379 = ~w13372 & w13377;
assign w13380 = ~w13378 & ~w13379;
assign w13381 = ~w13287 & ~w13312;
assign w13382 = ~w13380 & w13381;
assign w13383 = w13380 & ~w13381;
assign w13384 = ~w13382 & ~w13383;
assign w13385 = ~w13371 & w13384;
assign w13386 = w13371 & ~w13384;
assign w13387 = ~w13385 & ~w13386;
assign w13388 = ~w13370 & w13387;
assign w13389 = w13370 & ~w13387;
assign w13390 = ~w13388 & ~w13389;
assign w13391 = ~w13114 & ~w13293;
assign w13392 = ~w13292 & ~w13391;
assign w13393 = w13251 & ~w13254;
assign w13394 = ~w13256 & ~w13393;
assign w13395 = w13392 & ~w13394;
assign w13396 = ~w13392 & w13394;
assign w13397 = ~w13395 & ~w13396;
assign w13398 = w13083 & ~w13263;
assign w13399 = ~w13265 & ~w13398;
assign w13400 = ~w13397 & w13399;
assign w13401 = w13397 & ~w13399;
assign w13402 = ~w13400 & ~w13401;
assign w13403 = ~w13135 & ~w13240;
assign w13404 = ~w13239 & ~w13403;
assign w13405 = ~w13092 & ~w13304;
assign w13406 = ~w13303 & ~w13405;
assign w13407 = w13404 & w13406;
assign w13408 = ~w13404 & ~w13406;
assign w13409 = ~w13407 & ~w13408;
assign w13410 = pi43 & pi45;
assign w13411 = pi33 & pi55;
assign w13412 = pi34 & pi54;
assign w13413 = ~w13411 & ~w13412;
assign w13414 = pi34 & pi55;
assign w13415 = w13238 & w13414;
assign w13416 = ~w13413 & ~w13415;
assign w13417 = w13410 & ~w13416;
assign w13418 = ~w13410 & w13416;
assign w13419 = ~w13417 & ~w13418;
assign w13420 = ~w13409 & w13419;
assign w13421 = w13409 & ~w13419;
assign w13422 = ~w13420 & ~w13421;
assign w13423 = ~w13245 & ~w13249;
assign w13424 = w13422 & ~w13423;
assign w13425 = ~w13422 & w13423;
assign w13426 = ~w13424 & ~w13425;
assign w13427 = w13402 & w13426;
assign w13428 = ~w13402 & ~w13426;
assign w13429 = ~w13427 & ~w13428;
assign w13430 = (~w13343 & ~w13345) | (~w13343 & w17221) | (~w13345 & w17221);
assign w13431 = (~w13214 & ~w13216) | (~w13214 & w17222) | (~w13216 & w17222);
assign w13432 = ~w13430 & ~w13431;
assign w13433 = w13430 & w13431;
assign w13434 = ~w13432 & ~w13433;
assign w13435 = w13429 & w13434;
assign w13436 = ~w13429 & ~w13434;
assign w13437 = ~w13435 & ~w13436;
assign w13438 = ~w13220 & ~w13225;
assign w13439 = pi26 & pi62;
assign w13440 = pi28 & pi60;
assign w13441 = ~w13255 & ~w13440;
assign w13442 = pi28 & pi61;
assign w13443 = w13253 & w13442;
assign w13444 = ~w13441 & ~w13443;
assign w13445 = w13439 & ~w13444;
assign w13446 = ~w13439 & w13444;
assign w13447 = ~w13445 & ~w13446;
assign w13448 = pi31 & pi57;
assign w13449 = pi41 & pi47;
assign w13450 = ~w13277 & ~w13449;
assign w13451 = pi42 & pi47;
assign w13452 = w13274 & w13451;
assign w13453 = ~w13450 & ~w13452;
assign w13454 = w13448 & ~w13453;
assign w13455 = ~w13448 & w13453;
assign w13456 = ~w13454 & ~w13455;
assign w13457 = ~w13447 & ~w13456;
assign w13458 = w13447 & w13456;
assign w13459 = ~w13457 & ~w13458;
assign w13460 = pi35 & pi53;
assign w13461 = pi37 & pi51;
assign w13462 = pi36 & pi52;
assign w13463 = ~w13461 & ~w13462;
assign w13464 = pi37 & pi52;
assign w13465 = w13302 & w13464;
assign w13466 = ~w13463 & ~w13465;
assign w13467 = w13460 & ~w13466;
assign w13468 = ~w13460 & w13466;
assign w13469 = ~w13467 & ~w13468;
assign w13470 = w13459 & ~w13469;
assign w13471 = ~w13459 & w13469;
assign w13472 = ~w13470 & ~w13471;
assign w13473 = (~w13323 & ~w13325) | (~w13323 & w17223) | (~w13325 & w17223);
assign w13474 = pi29 & pi59;
assign w13475 = pi38 & pi50;
assign w13476 = ~w13264 & ~w13475;
assign w13477 = pi39 & pi50;
assign w13478 = w13261 & w13477;
assign w13479 = ~w13476 & ~w13478;
assign w13480 = w13474 & ~w13479;
assign w13481 = ~w13474 & w13479;
assign w13482 = ~w13480 & ~w13481;
assign w13483 = pi40 & pi48;
assign w13484 = pi30 & pi58;
assign w13485 = pi32 & pi56;
assign w13486 = ~w13484 & ~w13485;
assign w13487 = w13484 & w13485;
assign w13488 = ~w13486 & ~w13487;
assign w13489 = w13483 & ~w13488;
assign w13490 = ~w13483 & w13488;
assign w13491 = ~w13489 & ~w13490;
assign w13492 = ~w13482 & ~w13491;
assign w13493 = w13482 & w13491;
assign w13494 = ~w13492 & ~w13493;
assign w13495 = w13473 & ~w13494;
assign w13496 = ~w13473 & w13494;
assign w13497 = ~w13495 & ~w13496;
assign w13498 = pi25 & pi63;
assign w13499 = ~pi43 & ~w13049;
assign w13500 = pi44 & ~w13499;
assign w13501 = w13498 & w13500;
assign w13502 = ~w13498 & ~w13500;
assign w13503 = ~w13501 & ~w13502;
assign w13504 = w13273 & ~w13276;
assign w13505 = ~w13278 & ~w13504;
assign w13506 = ~w13503 & w13505;
assign w13507 = w13503 & ~w13505;
assign w13508 = ~w13506 & ~w13507;
assign w13509 = w13497 & w13508;
assign w13510 = ~w13497 & ~w13508;
assign w13511 = ~w13509 & ~w13510;
assign w13512 = w13472 & w13511;
assign w13513 = ~w13472 & ~w13511;
assign w13514 = ~w13512 & ~w13513;
assign w13515 = ~w13438 & w13514;
assign w13516 = w13438 & ~w13514;
assign w13517 = ~w13515 & ~w13516;
assign w13518 = w13437 & w13517;
assign w13519 = ~w13437 & ~w13517;
assign w13520 = ~w13518 & ~w13519;
assign w13521 = ~w13390 & ~w13520;
assign w13522 = w13390 & w13520;
assign w13523 = ~w13521 & ~w13522;
assign w13524 = w13369 & ~w13523;
assign w13525 = ~w13369 & w13523;
assign w13526 = ~w13524 & ~w13525;
assign w13527 = (w11122 & w17638) | (w11122 & w17639) | (w17638 & w17639);
assign w13528 = (~w11122 & w17640) | (~w11122 & w17641) | (w17640 & w17641);
assign w13529 = ~w13527 & ~w13528;
assign w13530 = ~w13388 & ~w13522;
assign w13531 = ~w13407 & ~w13421;
assign w13532 = (~w13395 & ~w13397) | (~w13395 & w17224) | (~w13397 & w17224);
assign w13533 = ~w13501 & ~w13507;
assign w13534 = ~w13532 & ~w13533;
assign w13535 = w13532 & w13533;
assign w13536 = ~w13534 & ~w13535;
assign w13537 = w13531 & ~w13536;
assign w13538 = ~w13531 & w13536;
assign w13539 = ~w13537 & ~w13538;
assign w13540 = (~w13375 & ~w13377) | (~w13375 & w17225) | (~w13377 & w17225);
assign w13541 = ~w13539 & w13540;
assign w13542 = w13539 & ~w13540;
assign w13543 = ~w13541 & ~w13542;
assign w13544 = ~w13424 & ~w13427;
assign w13545 = w13543 & ~w13544;
assign w13546 = ~w13543 & w13544;
assign w13547 = ~w13545 & ~w13546;
assign w13548 = ~w13383 & ~w13385;
assign w13549 = w13439 & ~w13441;
assign w13550 = ~w13443 & ~w13549;
assign w13551 = w13460 & ~w13463;
assign w13552 = ~w13465 & ~w13551;
assign w13553 = ~w13550 & ~w13552;
assign w13554 = w13550 & w13552;
assign w13555 = ~w13553 & ~w13554;
assign w13556 = ~w13483 & ~w13487;
assign w13557 = ~w13486 & ~w13556;
assign w13558 = ~w13555 & ~w13557;
assign w13559 = w13555 & w13557;
assign w13560 = ~w13558 & ~w13559;
assign w13561 = pi29 & pi60;
assign w13562 = ~w13442 & ~w13561;
assign w13563 = pi29 & pi61;
assign w13564 = w13440 & w13563;
assign w13565 = ~w13562 & ~w13564;
assign w13566 = w13410 & ~w13413;
assign w13567 = ~w13415 & ~w13566;
assign w13568 = w13565 & ~w13567;
assign w13569 = ~w13565 & w13567;
assign w13570 = ~w13568 & ~w13569;
assign w13571 = pi43 & pi46;
assign w13572 = ~w13451 & ~w13571;
assign w13573 = pi43 & pi47;
assign w13574 = w13277 & w13573;
assign w13575 = ~w13572 & ~w13574;
assign w13576 = w13414 & ~w13575;
assign w13577 = ~w13414 & w13575;
assign w13578 = ~w13576 & ~w13577;
assign w13579 = pi27 & pi62;
assign w13580 = ~pi44 & pi45;
assign w13581 = w13579 & ~w13580;
assign w13582 = ~w13579 & w13580;
assign w13583 = ~w13581 & ~w13582;
assign w13584 = ~w13578 & ~w13583;
assign w13585 = w13578 & w13583;
assign w13586 = ~w13584 & ~w13585;
assign w13587 = w13570 & w13586;
assign w13588 = ~w13570 & ~w13586;
assign w13589 = ~w13587 & ~w13588;
assign w13590 = ~w13560 & ~w13589;
assign w13591 = w13560 & w13589;
assign w13592 = ~w13590 & ~w13591;
assign w13593 = pi36 & pi53;
assign w13594 = pi38 & pi51;
assign w13595 = ~w13464 & ~w13594;
assign w13596 = pi38 & pi52;
assign w13597 = w13461 & w13596;
assign w13598 = ~w13595 & ~w13597;
assign w13599 = w13593 & ~w13598;
assign w13600 = ~w13593 & w13598;
assign w13601 = ~w13599 & ~w13600;
assign w13602 = pi41 & pi48;
assign w13603 = pi33 & pi56;
assign w13604 = pi35 & pi54;
assign w13605 = ~w13603 & ~w13604;
assign w13606 = w13603 & w13604;
assign w13607 = ~w13605 & ~w13606;
assign w13608 = w13602 & ~w13607;
assign w13609 = ~w13602 & w13607;
assign w13610 = ~w13608 & ~w13609;
assign w13611 = ~w13601 & ~w13610;
assign w13612 = w13601 & w13610;
assign w13613 = ~w13611 & ~w13612;
assign w13614 = pi30 & pi59;
assign w13615 = pi32 & pi57;
assign w13616 = pi31 & pi58;
assign w13617 = ~w13615 & ~w13616;
assign w13618 = pi32 & pi58;
assign w13619 = w13448 & w13618;
assign w13620 = ~w13617 & ~w13619;
assign w13621 = w13614 & ~w13620;
assign w13622 = ~w13614 & w13620;
assign w13623 = ~w13621 & ~w13622;
assign w13624 = w13613 & ~w13623;
assign w13625 = ~w13613 & w13623;
assign w13626 = ~w13624 & ~w13625;
assign w13627 = w13592 & w13626;
assign w13628 = ~w13592 & ~w13626;
assign w13629 = ~w13627 & ~w13628;
assign w13630 = ~w13548 & w13629;
assign w13631 = w13548 & ~w13629;
assign w13632 = ~w13630 & ~w13631;
assign w13633 = w13547 & w13632;
assign w13634 = ~w13547 & ~w13632;
assign w13635 = ~w13633 & ~w13634;
assign w13636 = ~w13432 & ~w13435;
assign w13637 = ~w13509 & ~w13512;
assign w13638 = w13448 & ~w13450;
assign w13639 = ~w13452 & ~w13638;
assign w13640 = w13474 & ~w13476;
assign w13641 = ~w13478 & ~w13640;
assign w13642 = ~w13639 & ~w13641;
assign w13643 = w13639 & w13641;
assign w13644 = ~w13642 & ~w13643;
assign w13645 = pi26 & pi63;
assign w13646 = pi40 & pi49;
assign w13647 = ~w13477 & ~w13646;
assign w13648 = pi40 & pi50;
assign w13649 = w13264 & w13648;
assign w13650 = ~w13647 & ~w13649;
assign w13651 = w13645 & ~w13650;
assign w13652 = ~w13645 & w13650;
assign w13653 = ~w13651 & ~w13652;
assign w13654 = ~w13644 & w13653;
assign w13655 = w13644 & ~w13653;
assign w13656 = ~w13654 & ~w13655;
assign w13657 = ~w13492 & ~w13496;
assign w13658 = ~w13457 & ~w13470;
assign w13659 = ~w13657 & ~w13658;
assign w13660 = w13657 & w13658;
assign w13661 = ~w13659 & ~w13660;
assign w13662 = ~w13656 & ~w13661;
assign w13663 = w13656 & w13661;
assign w13664 = ~w13662 & ~w13663;
assign w13665 = ~w13637 & w13664;
assign w13666 = w13637 & ~w13664;
assign w13667 = ~w13665 & ~w13666;
assign w13668 = ~w13636 & w13667;
assign w13669 = w13636 & ~w13667;
assign w13670 = ~w13668 & ~w13669;
assign w13671 = ~w13515 & ~w13518;
assign w13672 = w13670 & ~w13671;
assign w13673 = ~w13670 & w13671;
assign w13674 = ~w13672 & ~w13673;
assign w13675 = w13635 & w13674;
assign w13676 = ~w13635 & ~w13674;
assign w13677 = ~w13675 & ~w13676;
assign w13678 = ~w13530 & w13677;
assign w13679 = w13530 & ~w13677;
assign w13680 = ~w13678 & ~w13679;
assign w13681 = ~w13363 & ~w13524;
assign w13682 = (~w11122 & w17642) | (~w11122 & w17643) | (w17642 & w17643);
assign w13683 = (w11122 & w17644) | (w11122 & w17645) | (w17644 & w17645);
assign w13684 = ~w13682 & ~w13683;
assign w13685 = ~w13525 & ~w13678;
assign w13686 = ~w13672 & ~w13675;
assign w13687 = ~w13542 & ~w13545;
assign w13688 = ~w13591 & ~w13627;
assign w13689 = ~pi44 & ~w13579;
assign w13690 = pi45 & ~w13689;
assign w13691 = w13414 & ~w13572;
assign w13692 = ~w13574 & ~w13691;
assign w13693 = w13690 & ~w13692;
assign w13694 = ~w13690 & w13692;
assign w13695 = ~w13693 & ~w13694;
assign w13696 = ~w13602 & ~w13606;
assign w13697 = ~w13605 & ~w13696;
assign w13698 = ~w13695 & ~w13697;
assign w13699 = w13695 & w13697;
assign w13700 = ~w13698 & ~w13699;
assign w13701 = ~w13584 & ~w13587;
assign w13702 = ~w13611 & ~w13624;
assign w13703 = ~w13701 & ~w13702;
assign w13704 = w13701 & w13702;
assign w13705 = ~w13703 & ~w13704;
assign w13706 = w13700 & w13705;
assign w13707 = ~w13700 & ~w13705;
assign w13708 = ~w13706 & ~w13707;
assign w13709 = ~w13688 & w13708;
assign w13710 = w13688 & ~w13708;
assign w13711 = ~w13709 & ~w13710;
assign w13712 = w13687 & ~w13711;
assign w13713 = ~w13687 & w13711;
assign w13714 = ~w13712 & ~w13713;
assign w13715 = ~w13630 & ~w13633;
assign w13716 = ~w13714 & w13715;
assign w13717 = w13714 & ~w13715;
assign w13718 = ~w13716 & ~w13717;
assign w13719 = ~w13665 & ~w13668;
assign w13720 = w13614 & ~w13617;
assign w13721 = ~w13619 & ~w13720;
assign w13722 = w13593 & ~w13595;
assign w13723 = ~w13597 & ~w13722;
assign w13724 = ~w13721 & ~w13723;
assign w13725 = w13721 & w13723;
assign w13726 = ~w13724 & ~w13725;
assign w13727 = w13645 & ~w13647;
assign w13728 = ~w13649 & ~w13727;
assign w13729 = ~w13726 & w13728;
assign w13730 = w13726 & ~w13728;
assign w13731 = ~w13729 & ~w13730;
assign w13732 = ~w13534 & ~w13538;
assign w13733 = ~w13731 & w13732;
assign w13734 = w13731 & ~w13732;
assign w13735 = ~w13733 & ~w13734;
assign w13736 = pi35 & pi55;
assign w13737 = pi33 & pi57;
assign w13738 = pi34 & pi56;
assign w13739 = ~w13737 & ~w13738;
assign w13740 = pi34 & pi57;
assign w13741 = w13603 & w13740;
assign w13742 = ~w13739 & ~w13741;
assign w13743 = w13736 & ~w13742;
assign w13744 = ~w13736 & w13742;
assign w13745 = ~w13743 & ~w13744;
assign w13746 = pi36 & pi54;
assign w13747 = pi37 & pi53;
assign w13748 = ~w13596 & ~w13747;
assign w13749 = pi38 & pi53;
assign w13750 = w13464 & w13749;
assign w13751 = ~w13748 & ~w13750;
assign w13752 = w13746 & ~w13751;
assign w13753 = ~w13746 & w13751;
assign w13754 = ~w13752 & ~w13753;
assign w13755 = ~w13745 & ~w13754;
assign w13756 = w13745 & w13754;
assign w13757 = ~w13755 & ~w13756;
assign w13758 = pi42 & pi48;
assign w13759 = pi44 & pi46;
assign w13760 = ~w13573 & ~w13759;
assign w13761 = pi44 & pi47;
assign w13762 = w13571 & w13761;
assign w13763 = ~w13760 & ~w13762;
assign w13764 = w13758 & ~w13763;
assign w13765 = ~w13758 & w13763;
assign w13766 = ~w13764 & ~w13765;
assign w13767 = w13757 & ~w13766;
assign w13768 = ~w13757 & w13766;
assign w13769 = ~w13767 & ~w13768;
assign w13770 = w13735 & w13769;
assign w13771 = ~w13735 & ~w13769;
assign w13772 = ~w13770 & ~w13771;
assign w13773 = ~w13719 & w13772;
assign w13774 = w13719 & ~w13772;
assign w13775 = ~w13773 & ~w13774;
assign w13776 = ~w13659 & ~w13663;
assign w13777 = ~w13642 & ~w13655;
assign w13778 = (~w13553 & ~w13555) | (~w13553 & w17226) | (~w13555 & w17226);
assign w13779 = pi39 & pi51;
assign w13780 = pi41 & pi49;
assign w13781 = ~w13648 & ~w13780;
assign w13782 = pi41 & pi50;
assign w13783 = w13646 & w13782;
assign w13784 = ~w13781 & ~w13783;
assign w13785 = w13779 & ~w13784;
assign w13786 = ~w13779 & w13784;
assign w13787 = ~w13785 & ~w13786;
assign w13788 = ~w13778 & ~w13787;
assign w13789 = w13778 & w13787;
assign w13790 = ~w13788 & ~w13789;
assign w13791 = w13777 & ~w13790;
assign w13792 = ~w13777 & w13790;
assign w13793 = ~w13791 & ~w13792;
assign w13794 = ~w13564 & ~w13568;
assign w13795 = pi30 & pi60;
assign w13796 = pi31 & pi59;
assign w13797 = ~w13618 & ~w13796;
assign w13798 = pi32 & pi59;
assign w13799 = w13616 & w13798;
assign w13800 = ~w13797 & ~w13799;
assign w13801 = w13795 & ~w13800;
assign w13802 = ~w13795 & w13800;
assign w13803 = ~w13801 & ~w13802;
assign w13804 = ~w13794 & ~w13803;
assign w13805 = w13794 & w13803;
assign w13806 = ~w13804 & ~w13805;
assign w13807 = pi27 & pi63;
assign w13808 = pi28 & pi62;
assign w13809 = ~w13563 & ~w13808;
assign w13810 = pi29 & pi62;
assign w13811 = w13442 & w13810;
assign w13812 = ~w13809 & ~w13811;
assign w13813 = w13807 & ~w13812;
assign w13814 = ~w13807 & w13812;
assign w13815 = ~w13813 & ~w13814;
assign w13816 = w13806 & ~w13815;
assign w13817 = ~w13806 & w13815;
assign w13818 = ~w13816 & ~w13817;
assign w13819 = w13793 & w13818;
assign w13820 = ~w13793 & ~w13818;
assign w13821 = ~w13819 & ~w13820;
assign w13822 = ~w13776 & w13821;
assign w13823 = w13776 & ~w13821;
assign w13824 = ~w13822 & ~w13823;
assign w13825 = w13775 & w13824;
assign w13826 = ~w13775 & ~w13824;
assign w13827 = ~w13825 & ~w13826;
assign w13828 = ~w13718 & ~w13827;
assign w13829 = w13718 & w13827;
assign w13830 = ~w13828 & ~w13829;
assign w13831 = ~w13686 & w13830;
assign w13832 = w13686 & ~w13830;
assign w13833 = ~w13831 & ~w13832;
assign w13834 = (~w10008 & w17861) | (~w10008 & w17862) | (w17861 & w17862);
assign w13835 = (w10008 & w17863) | (w10008 & w17864) | (w17863 & w17864);
assign w13836 = ~w13834 & ~w13835;
assign w13837 = ~w13717 & ~w13829;
assign w13838 = w13746 & ~w13748;
assign w13839 = ~w13750 & ~w13838;
assign w13840 = w13807 & ~w13809;
assign w13841 = ~w13811 & ~w13840;
assign w13842 = ~w13839 & ~w13841;
assign w13843 = w13839 & w13841;
assign w13844 = ~w13842 & ~w13843;
assign w13845 = w13795 & ~w13797;
assign w13846 = ~w13799 & ~w13845;
assign w13847 = ~w13844 & w13846;
assign w13848 = w13844 & ~w13846;
assign w13849 = ~w13847 & ~w13848;
assign w13850 = ~w13788 & ~w13792;
assign w13851 = ~w13849 & w13850;
assign w13852 = w13849 & ~w13850;
assign w13853 = ~w13851 & ~w13852;
assign w13854 = pi28 & pi63;
assign w13855 = pi40 & pi51;
assign w13856 = ~w13782 & ~w13855;
assign w13857 = pi41 & pi51;
assign w13858 = w13648 & w13857;
assign w13859 = ~w13856 & ~w13858;
assign w13860 = w13854 & ~w13859;
assign w13861 = ~w13854 & w13859;
assign w13862 = ~w13860 & ~w13861;
assign w13863 = pi35 & pi56;
assign w13864 = pi43 & pi48;
assign w13865 = ~w13761 & ~w13864;
assign w13866 = pi44 & pi48;
assign w13867 = w13573 & w13866;
assign w13868 = ~w13865 & ~w13867;
assign w13869 = w13863 & ~w13868;
assign w13870 = ~w13863 & w13868;
assign w13871 = ~w13869 & ~w13870;
assign w13872 = ~w13862 & ~w13871;
assign w13873 = w13862 & w13871;
assign w13874 = ~w13872 & ~w13873;
assign w13875 = ~pi45 & pi46;
assign w13876 = w13810 & ~w13875;
assign w13877 = ~w13810 & w13875;
assign w13878 = ~w13876 & ~w13877;
assign w13879 = w13874 & ~w13878;
assign w13880 = ~w13874 & w13878;
assign w13881 = ~w13879 & ~w13880;
assign w13882 = ~w13853 & ~w13881;
assign w13883 = w13853 & w13881;
assign w13884 = ~w13882 & ~w13883;
assign w13885 = ~w13709 & ~w13713;
assign w13886 = ~w13884 & w13885;
assign w13887 = w13884 & ~w13885;
assign w13888 = ~w13886 & ~w13887;
assign w13889 = ~w13724 & ~w13730;
assign w13890 = ~w13693 & ~w13699;
assign w13891 = pi42 & pi49;
assign w13892 = pi36 & pi55;
assign w13893 = ~w13740 & ~w13892;
assign w13894 = w13740 & w13892;
assign w13895 = ~w13893 & ~w13894;
assign w13896 = w13891 & ~w13895;
assign w13897 = ~w13891 & w13895;
assign w13898 = ~w13896 & ~w13897;
assign w13899 = ~w13890 & ~w13898;
assign w13900 = w13890 & w13898;
assign w13901 = ~w13899 & ~w13900;
assign w13902 = w13889 & ~w13901;
assign w13903 = ~w13889 & w13901;
assign w13904 = ~w13902 & ~w13903;
assign w13905 = ~w13703 & ~w13706;
assign w13906 = pi37 & pi54;
assign w13907 = pi39 & pi52;
assign w13908 = ~w13749 & ~w13907;
assign w13909 = pi39 & pi53;
assign w13910 = w13596 & w13909;
assign w13911 = ~w13908 & ~w13910;
assign w13912 = w13906 & ~w13911;
assign w13913 = ~w13906 & w13911;
assign w13914 = ~w13912 & ~w13913;
assign w13915 = w13779 & ~w13781;
assign w13916 = ~w13783 & ~w13915;
assign w13917 = ~w13914 & ~w13916;
assign w13918 = w13914 & w13916;
assign w13919 = ~w13917 & ~w13918;
assign w13920 = pi31 & pi60;
assign w13921 = pi33 & pi58;
assign w13922 = ~w13798 & ~w13921;
assign w13923 = pi33 & pi59;
assign w13924 = w13618 & w13923;
assign w13925 = ~w13922 & ~w13924;
assign w13926 = w13920 & ~w13925;
assign w13927 = ~w13920 & w13925;
assign w13928 = ~w13926 & ~w13927;
assign w13929 = w13919 & ~w13928;
assign w13930 = ~w13919 & w13928;
assign w13931 = ~w13929 & ~w13930;
assign w13932 = ~w13905 & w13931;
assign w13933 = w13905 & ~w13931;
assign w13934 = ~w13932 & ~w13933;
assign w13935 = w13904 & w13934;
assign w13936 = ~w13904 & ~w13934;
assign w13937 = ~w13935 & ~w13936;
assign w13938 = w13888 & w13937;
assign w13939 = ~w13888 & ~w13937;
assign w13940 = ~w13938 & ~w13939;
assign w13941 = ~w13773 & ~w13825;
assign w13942 = ~w13819 & ~w13822;
assign w13943 = ~w13734 & ~w13770;
assign w13944 = pi30 & pi61;
assign w13945 = w13758 & ~w13760;
assign w13946 = ~w13762 & ~w13945;
assign w13947 = w13944 & ~w13946;
assign w13948 = ~w13944 & w13946;
assign w13949 = ~w13947 & ~w13948;
assign w13950 = w13736 & ~w13739;
assign w13951 = ~w13741 & ~w13950;
assign w13952 = ~w13949 & w13951;
assign w13953 = w13949 & ~w13951;
assign w13954 = ~w13952 & ~w13953;
assign w13955 = ~w13804 & ~w13816;
assign w13956 = ~w13755 & ~w13767;
assign w13957 = ~w13955 & ~w13956;
assign w13958 = w13955 & w13956;
assign w13959 = ~w13957 & ~w13958;
assign w13960 = w13954 & w13959;
assign w13961 = ~w13954 & ~w13959;
assign w13962 = ~w13960 & ~w13961;
assign w13963 = ~w13943 & w13962;
assign w13964 = w13943 & ~w13962;
assign w13965 = ~w13963 & ~w13964;
assign w13966 = ~w13942 & w13965;
assign w13967 = w13942 & ~w13965;
assign w13968 = ~w13966 & ~w13967;
assign w13969 = ~w13941 & w13968;
assign w13970 = w13941 & ~w13968;
assign w13971 = ~w13969 & ~w13970;
assign w13972 = w13940 & w13971;
assign w13973 = ~w13940 & ~w13971;
assign w13974 = ~w13972 & ~w13973;
assign w13975 = ~w13837 & w13974;
assign w13976 = w13837 & ~w13974;
assign w13977 = ~w13975 & ~w13976;
assign w13978 = (~w8795 & w17646) | (~w8795 & w17647) | (w17646 & w17647);
assign w13979 = (w11122 & w17648) | (w11122 & w17649) | (w17648 & w17649);
assign w13980 = (~w11122 & w17650) | (~w11122 & w17651) | (w17650 & w17651);
assign w13981 = ~w13979 & ~w13980;
assign w13982 = ~w13832 & ~w13976;
assign w13983 = ~w13963 & ~w13966;
assign w13984 = ~w13932 & ~w13935;
assign w13985 = ~w13957 & ~w13960;
assign w13986 = ~w13947 & ~w13953;
assign w13987 = pi31 & pi61;
assign w13988 = pi30 & pi62;
assign w13989 = ~w13987 & ~w13988;
assign w13990 = pi31 & pi62;
assign w13991 = w13944 & w13990;
assign w13992 = ~w13989 & ~w13991;
assign w13993 = ~pi45 & ~w13810;
assign w13994 = pi46 & ~w13993;
assign w13995 = w13992 & w13994;
assign w13996 = ~w13992 & ~w13994;
assign w13997 = ~w13995 & ~w13996;
assign w13998 = pi40 & pi52;
assign w13999 = ~w13857 & ~w13998;
assign w14000 = pi41 & pi52;
assign w14001 = w13855 & w14000;
assign w14002 = ~w13999 & ~w14001;
assign w14003 = w13909 & ~w14002;
assign w14004 = ~w13909 & w14002;
assign w14005 = ~w14003 & ~w14004;
assign w14006 = w13997 & ~w14005;
assign w14007 = ~w13997 & w14005;
assign w14008 = ~w14006 & ~w14007;
assign w14009 = w13986 & ~w14008;
assign w14010 = ~w13986 & w14008;
assign w14011 = ~w14009 & ~w14010;
assign w14012 = pi43 & pi49;
assign w14013 = pi45 & pi47;
assign w14014 = ~w13866 & ~w14013;
assign w14015 = pi45 & pi48;
assign w14016 = w13761 & w14015;
assign w14017 = ~w14014 & ~w14016;
assign w14018 = w14012 & ~w14017;
assign w14019 = ~w14012 & w14017;
assign w14020 = ~w14018 & ~w14019;
assign w14021 = pi34 & pi58;
assign w14022 = pi35 & pi57;
assign w14023 = pi42 & pi50;
assign w14024 = ~w14022 & ~w14023;
assign w14025 = w14022 & w14023;
assign w14026 = ~w14024 & ~w14025;
assign w14027 = w14021 & ~w14026;
assign w14028 = ~w14021 & w14026;
assign w14029 = ~w14027 & ~w14028;
assign w14030 = ~w14020 & ~w14029;
assign w14031 = w14020 & w14029;
assign w14032 = ~w14030 & ~w14031;
assign w14033 = pi36 & pi56;
assign w14034 = pi29 & pi63;
assign w14035 = ~w13923 & ~w14034;
assign w14036 = w13923 & w14034;
assign w14037 = ~w14035 & ~w14036;
assign w14038 = w14033 & ~w14037;
assign w14039 = ~w14033 & w14037;
assign w14040 = ~w14038 & ~w14039;
assign w14041 = w14032 & ~w14040;
assign w14042 = ~w14032 & w14040;
assign w14043 = ~w14041 & ~w14042;
assign w14044 = ~w14011 & ~w14043;
assign w14045 = w14011 & w14043;
assign w14046 = ~w14044 & ~w14045;
assign w14047 = ~w13985 & w14046;
assign w14048 = w13985 & ~w14046;
assign w14049 = ~w14047 & ~w14048;
assign w14050 = ~w13984 & w14049;
assign w14051 = w13984 & ~w14049;
assign w14052 = ~w14050 & ~w14051;
assign w14053 = ~w13983 & w14052;
assign w14054 = w13983 & ~w14052;
assign w14055 = ~w14053 & ~w14054;
assign w14056 = ~w13887 & ~w13938;
assign w14057 = ~w13872 & ~w13879;
assign w14058 = ~w13917 & ~w13929;
assign w14059 = ~w13842 & ~w13848;
assign w14060 = ~w14058 & ~w14059;
assign w14061 = w14058 & w14059;
assign w14062 = ~w14060 & ~w14061;
assign w14063 = w14057 & ~w14062;
assign w14064 = ~w14057 & w14062;
assign w14065 = ~w14063 & ~w14064;
assign w14066 = ~w13852 & ~w13883;
assign w14067 = ~w13899 & ~w13903;
assign w14068 = w13920 & ~w13922;
assign w14069 = ~w13924 & ~w14068;
assign w14070 = w13906 & ~w13908;
assign w14071 = ~w13910 & ~w14070;
assign w14072 = ~w14069 & ~w14071;
assign w14073 = w14069 & w14071;
assign w14074 = ~w14072 & ~w14073;
assign w14075 = w13854 & ~w13856;
assign w14076 = ~w13858 & ~w14075;
assign w14077 = ~w14074 & w14076;
assign w14078 = w14074 & ~w14076;
assign w14079 = ~w14077 & ~w14078;
assign w14080 = ~w13891 & ~w13894;
assign w14081 = ~w13893 & ~w14080;
assign w14082 = w13863 & ~w13865;
assign w14083 = ~w13867 & ~w14082;
assign w14084 = w14081 & ~w14083;
assign w14085 = ~w14081 & w14083;
assign w14086 = ~w14084 & ~w14085;
assign w14087 = pi32 & pi60;
assign w14088 = pi37 & pi55;
assign w14089 = pi38 & pi54;
assign w14090 = ~w14088 & ~w14089;
assign w14091 = pi38 & pi55;
assign w14092 = w13906 & w14091;
assign w14093 = ~w14090 & ~w14092;
assign w14094 = w14087 & ~w14093;
assign w14095 = ~w14087 & w14093;
assign w14096 = ~w14094 & ~w14095;
assign w14097 = ~w14086 & w14096;
assign w14098 = w14086 & ~w14096;
assign w14099 = ~w14097 & ~w14098;
assign w14100 = ~w14079 & ~w14099;
assign w14101 = w14079 & w14099;
assign w14102 = ~w14100 & ~w14101;
assign w14103 = ~w14067 & w14102;
assign w14104 = w14067 & ~w14102;
assign w14105 = ~w14103 & ~w14104;
assign w14106 = ~w14066 & w14105;
assign w14107 = w14066 & ~w14105;
assign w14108 = ~w14106 & ~w14107;
assign w14109 = w14065 & w14108;
assign w14110 = ~w14065 & ~w14108;
assign w14111 = ~w14109 & ~w14110;
assign w14112 = ~w14056 & w14111;
assign w14113 = w14056 & ~w14111;
assign w14114 = ~w14112 & ~w14113;
assign w14115 = w14055 & w14114;
assign w14116 = ~w14055 & ~w14114;
assign w14117 = ~w14115 & ~w14116;
assign w14118 = ~w13969 & ~w13972;
assign w14119 = w14117 & ~w14118;
assign w14120 = ~w14117 & w14118;
assign w14121 = ~w14119 & ~w14120;
assign w14122 = (w12329 & w17493) | (w12329 & w17494) | (w17493 & w17494);
assign w14123 = (~w12329 & w17495) | (~w12329 & w17496) | (w17495 & w17496);
assign w14124 = ~w14122 & ~w14123;
assign w14125 = ~w13975 & ~w14119;
assign w14126 = ~w14112 & ~w14115;
assign w14127 = ~w14050 & ~w14053;
assign w14128 = ~w14030 & ~w14041;
assign w14129 = ~w14084 & ~w14098;
assign w14130 = ~w14072 & ~w14078;
assign w14131 = ~w14129 & ~w14130;
assign w14132 = w14129 & w14130;
assign w14133 = ~w14131 & ~w14132;
assign w14134 = w14128 & ~w14133;
assign w14135 = ~w14128 & w14133;
assign w14136 = ~w14134 & ~w14135;
assign w14137 = ~w14101 & ~w14103;
assign w14138 = ~w14136 & w14137;
assign w14139 = w14136 & ~w14137;
assign w14140 = ~w14138 & ~w14139;
assign w14141 = ~w14006 & ~w14010;
assign w14142 = ~w14021 & ~w14025;
assign w14143 = ~w14024 & ~w14142;
assign w14144 = w14012 & ~w14014;
assign w14145 = ~w14016 & ~w14144;
assign w14146 = w14143 & ~w14145;
assign w14147 = ~w14143 & w14145;
assign w14148 = ~w14146 & ~w14147;
assign w14149 = w13909 & ~w13999;
assign w14150 = ~w14001 & ~w14149;
assign w14151 = ~w14148 & w14150;
assign w14152 = w14148 & ~w14150;
assign w14153 = ~w14151 & ~w14152;
assign w14154 = ~w13991 & ~w13995;
assign w14155 = ~w14033 & ~w14036;
assign w14156 = ~w14035 & ~w14155;
assign w14157 = w14087 & ~w14090;
assign w14158 = ~w14092 & ~w14157;
assign w14159 = w14156 & ~w14158;
assign w14160 = ~w14156 & w14158;
assign w14161 = ~w14159 & ~w14160;
assign w14162 = w14154 & ~w14161;
assign w14163 = ~w14154 & w14161;
assign w14164 = ~w14162 & ~w14163;
assign w14165 = w14153 & w14164;
assign w14166 = ~w14153 & ~w14164;
assign w14167 = ~w14165 & ~w14166;
assign w14168 = ~w14141 & w14167;
assign w14169 = w14141 & ~w14167;
assign w14170 = ~w14168 & ~w14169;
assign w14171 = w14140 & w14170;
assign w14172 = ~w14140 & ~w14170;
assign w14173 = ~w14171 & ~w14172;
assign w14174 = ~w14127 & w14173;
assign w14175 = w14127 & ~w14173;
assign w14176 = ~w14174 & ~w14175;
assign w14177 = ~w14106 & ~w14109;
assign w14178 = ~w14045 & ~w14047;
assign w14179 = ~w14060 & ~w14064;
assign w14180 = pi30 & pi63;
assign w14181 = pi32 & pi61;
assign w14182 = pi33 & pi60;
assign w14183 = ~w14181 & ~w14182;
assign w14184 = pi33 & pi61;
assign w14185 = w14087 & w14184;
assign w14186 = ~w14183 & ~w14185;
assign w14187 = w14180 & ~w14186;
assign w14188 = ~w14180 & w14186;
assign w14189 = ~w14187 & ~w14188;
assign w14190 = pi35 & pi58;
assign w14191 = pi36 & pi57;
assign w14192 = pi39 & pi54;
assign w14193 = ~w14191 & ~w14192;
assign w14194 = w14191 & w14192;
assign w14195 = ~w14193 & ~w14194;
assign w14196 = w14190 & ~w14195;
assign w14197 = ~w14190 & w14195;
assign w14198 = ~w14196 & ~w14197;
assign w14199 = ~w14189 & ~w14198;
assign w14200 = w14189 & w14198;
assign w14201 = ~w14199 & ~w14200;
assign w14202 = pi34 & pi59;
assign w14203 = pi40 & pi53;
assign w14204 = ~w14000 & ~w14203;
assign w14205 = pi41 & pi53;
assign w14206 = w13998 & w14205;
assign w14207 = ~w14204 & ~w14206;
assign w14208 = w14202 & ~w14207;
assign w14209 = ~w14202 & w14207;
assign w14210 = ~w14208 & ~w14209;
assign w14211 = w14201 & ~w14210;
assign w14212 = ~w14201 & w14210;
assign w14213 = ~w14211 & ~w14212;
assign w14214 = pi42 & pi51;
assign w14215 = pi44 & pi49;
assign w14216 = pi43 & pi50;
assign w14217 = ~w14215 & ~w14216;
assign w14218 = pi44 & pi50;
assign w14219 = w14012 & w14218;
assign w14220 = ~w14217 & ~w14219;
assign w14221 = w14214 & ~w14220;
assign w14222 = ~w14214 & w14220;
assign w14223 = ~w14221 & ~w14222;
assign w14224 = pi37 & pi56;
assign w14225 = ~w14015 & ~w14091;
assign w14226 = w14015 & w14091;
assign w14227 = ~w14225 & ~w14226;
assign w14228 = w14224 & ~w14227;
assign w14229 = ~w14224 & w14227;
assign w14230 = ~w14228 & ~w14229;
assign w14231 = ~w14223 & ~w14230;
assign w14232 = w14223 & w14230;
assign w14233 = ~w14231 & ~w14232;
assign w14234 = ~pi46 & pi47;
assign w14235 = w13990 & ~w14234;
assign w14236 = ~w13990 & w14234;
assign w14237 = ~w14235 & ~w14236;
assign w14238 = w14233 & ~w14237;
assign w14239 = ~w14233 & w14237;
assign w14240 = ~w14238 & ~w14239;
assign w14241 = w14213 & w14240;
assign w14242 = ~w14213 & ~w14240;
assign w14243 = ~w14241 & ~w14242;
assign w14244 = ~w14179 & w14243;
assign w14245 = w14179 & ~w14243;
assign w14246 = ~w14244 & ~w14245;
assign w14247 = ~w14178 & w14246;
assign w14248 = w14178 & ~w14246;
assign w14249 = ~w14247 & ~w14248;
assign w14250 = w14177 & ~w14249;
assign w14251 = ~w14177 & w14249;
assign w14252 = ~w14250 & ~w14251;
assign w14253 = w14176 & w14252;
assign w14254 = ~w14176 & ~w14252;
assign w14255 = ~w14253 & ~w14254;
assign w14256 = ~w14126 & w14255;
assign w14257 = w14126 & ~w14255;
assign w14258 = ~w14256 & ~w14257;
assign w14259 = (w11122 & w17652) | (w11122 & w17653) | (w17652 & w17653);
assign w14260 = (~w11122 & w17654) | (~w11122 & w17655) | (w17654 & w17655);
assign w14261 = ~w14259 & ~w14260;
assign w14262 = ~w14247 & ~w14251;
assign w14263 = ~w14241 & ~w14244;
assign w14264 = ~w14199 & ~w14211;
assign w14265 = ~w14159 & ~w14163;
assign w14266 = ~w14146 & ~w14152;
assign w14267 = ~w14265 & ~w14266;
assign w14268 = w14265 & w14266;
assign w14269 = ~w14267 & ~w14268;
assign w14270 = w14264 & ~w14269;
assign w14271 = ~w14264 & w14269;
assign w14272 = ~w14270 & ~w14271;
assign w14273 = ~w14165 & ~w14168;
assign w14274 = ~w14272 & w14273;
assign w14275 = w14272 & ~w14273;
assign w14276 = ~w14274 & ~w14275;
assign w14277 = ~w14263 & w14276;
assign w14278 = w14263 & ~w14276;
assign w14279 = ~w14277 & ~w14278;
assign w14280 = ~w14262 & w14279;
assign w14281 = w14262 & ~w14279;
assign w14282 = ~w14280 & ~w14281;
assign w14283 = ~w14139 & ~w14171;
assign w14284 = ~w14231 & ~w14238;
assign w14285 = pi31 & pi63;
assign w14286 = ~pi46 & ~w13990;
assign w14287 = pi47 & ~w14286;
assign w14288 = w14285 & w14287;
assign w14289 = ~w14285 & ~w14287;
assign w14290 = ~w14288 & ~w14289;
assign w14291 = ~w14224 & ~w14226;
assign w14292 = ~w14225 & ~w14291;
assign w14293 = w14290 & w14292;
assign w14294 = ~w14290 & ~w14292;
assign w14295 = ~w14293 & ~w14294;
assign w14296 = w14284 & ~w14295;
assign w14297 = ~w14284 & w14295;
assign w14298 = ~w14296 & ~w14297;
assign w14299 = ~w14190 & ~w14194;
assign w14300 = ~w14193 & ~w14299;
assign w14301 = w14180 & ~w14183;
assign w14302 = ~w14185 & ~w14301;
assign w14303 = w14300 & ~w14302;
assign w14304 = ~w14300 & w14302;
assign w14305 = ~w14303 & ~w14304;
assign w14306 = w14202 & ~w14204;
assign w14307 = ~w14206 & ~w14306;
assign w14308 = ~w14305 & w14307;
assign w14309 = w14305 & ~w14307;
assign w14310 = ~w14308 & ~w14309;
assign w14311 = w14298 & w14310;
assign w14312 = ~w14298 & ~w14310;
assign w14313 = ~w14311 & ~w14312;
assign w14314 = ~w14283 & w14313;
assign w14315 = w14283 & ~w14313;
assign w14316 = ~w14314 & ~w14315;
assign w14317 = ~w14131 & ~w14135;
assign w14318 = pi36 & pi58;
assign w14319 = pi43 & pi51;
assign w14320 = ~w14218 & ~w14319;
assign w14321 = pi44 & pi51;
assign w14322 = w14216 & w14321;
assign w14323 = ~w14320 & ~w14322;
assign w14324 = w14318 & ~w14323;
assign w14325 = ~w14318 & w14323;
assign w14326 = ~w14324 & ~w14325;
assign w14327 = pi40 & pi54;
assign w14328 = pi42 & pi52;
assign w14329 = ~w14205 & ~w14328;
assign w14330 = pi42 & pi53;
assign w14331 = w14000 & w14330;
assign w14332 = ~w14329 & ~w14331;
assign w14333 = w14327 & ~w14332;
assign w14334 = ~w14327 & w14332;
assign w14335 = ~w14333 & ~w14334;
assign w14336 = ~w14326 & ~w14335;
assign w14337 = w14326 & w14335;
assign w14338 = ~w14336 & ~w14337;
assign w14339 = pi45 & pi49;
assign w14340 = pi38 & pi56;
assign w14341 = pi46 & pi48;
assign w14342 = ~w14340 & ~w14341;
assign w14343 = w14340 & w14341;
assign w14344 = ~w14342 & ~w14343;
assign w14345 = w14339 & ~w14344;
assign w14346 = ~w14339 & w14344;
assign w14347 = ~w14345 & ~w14346;
assign w14348 = w14338 & ~w14347;
assign w14349 = ~w14338 & w14347;
assign w14350 = ~w14348 & ~w14349;
assign w14351 = ~w14317 & w14350;
assign w14352 = w14317 & ~w14350;
assign w14353 = ~w14351 & ~w14352;
assign w14354 = w14214 & ~w14217;
assign w14355 = ~w14219 & ~w14354;
assign w14356 = pi35 & pi59;
assign w14357 = ~w14184 & ~w14356;
assign w14358 = w14184 & w14356;
assign w14359 = ~w14357 & ~w14358;
assign w14360 = w8301 & ~w14359;
assign w14361 = ~w8301 & w14359;
assign w14362 = ~w14360 & ~w14361;
assign w14363 = ~w14355 & ~w14362;
assign w14364 = w14355 & w14362;
assign w14365 = ~w14363 & ~w14364;
assign w14366 = pi37 & pi57;
assign w14367 = pi34 & pi60;
assign w14368 = pi39 & pi55;
assign w14369 = ~w14367 & ~w14368;
assign w14370 = w14367 & w14368;
assign w14371 = ~w14369 & ~w14370;
assign w14372 = w14366 & ~w14371;
assign w14373 = ~w14366 & w14371;
assign w14374 = ~w14372 & ~w14373;
assign w14375 = w14365 & ~w14374;
assign w14376 = ~w14365 & w14374;
assign w14377 = ~w14375 & ~w14376;
assign w14378 = w14353 & w14377;
assign w14379 = ~w14353 & ~w14377;
assign w14380 = ~w14378 & ~w14379;
assign w14381 = w14316 & w14380;
assign w14382 = ~w14316 & ~w14380;
assign w14383 = ~w14381 & ~w14382;
assign w14384 = ~w14282 & ~w14383;
assign w14385 = w14282 & w14383;
assign w14386 = ~w14384 & ~w14385;
assign w14387 = ~w14174 & ~w14253;
assign w14388 = ~w14386 & w14387;
assign w14389 = w14386 & ~w14387;
assign w14390 = ~w14388 & ~w14389;
assign w14391 = (~w12329 & w17497) | (~w12329 & w17498) | (w17497 & w17498);
assign w14392 = (w12329 & w17499) | (w12329 & w17500) | (w17499 & w17500);
assign w14393 = ~w14391 & ~w14392;
assign w14394 = ~w14314 & ~w14381;
assign w14395 = ~w14351 & ~w14378;
assign w14396 = ~w14303 & ~w14309;
assign w14397 = pi36 & pi59;
assign w14398 = pi35 & pi60;
assign w14399 = ~w14397 & ~w14398;
assign w14400 = pi36 & pi60;
assign w14401 = w14356 & w14400;
assign w14402 = ~w14399 & ~w14401;
assign w14403 = ~w14339 & ~w14343;
assign w14404 = ~w14342 & ~w14403;
assign w14405 = w14402 & w14404;
assign w14406 = ~w14402 & ~w14404;
assign w14407 = ~w14405 & ~w14406;
assign w14408 = ~w14288 & ~w14293;
assign w14409 = w14407 & ~w14408;
assign w14410 = ~w14407 & w14408;
assign w14411 = ~w14409 & ~w14410;
assign w14412 = w14396 & ~w14411;
assign w14413 = ~w14396 & w14411;
assign w14414 = ~w14412 & ~w14413;
assign w14415 = ~w14297 & ~w14311;
assign w14416 = ~w14414 & w14415;
assign w14417 = w14414 & ~w14415;
assign w14418 = ~w14416 & ~w14417;
assign w14419 = ~w14395 & w14418;
assign w14420 = w14395 & ~w14418;
assign w14421 = ~w14419 & ~w14420;
assign w14422 = ~w14394 & w14421;
assign w14423 = w14394 & ~w14421;
assign w14424 = ~w14422 & ~w14423;
assign w14425 = ~w14267 & ~w14271;
assign w14426 = pi39 & pi56;
assign w14427 = pi46 & pi49;
assign w14428 = pi45 & pi50;
assign w14429 = ~w14427 & ~w14428;
assign w14430 = pi46 & pi50;
assign w14431 = w14339 & w14430;
assign w14432 = ~w14429 & ~w14431;
assign w14433 = w14426 & ~w14432;
assign w14434 = ~w14426 & w14432;
assign w14435 = ~w14433 & ~w14434;
assign w14436 = pi33 & pi62;
assign w14437 = ~pi47 & pi48;
assign w14438 = w14436 & ~w14437;
assign w14439 = ~w14436 & w14437;
assign w14440 = ~w14438 & ~w14439;
assign w14441 = ~w14435 & ~w14440;
assign w14442 = w14435 & w14440;
assign w14443 = ~w14441 & ~w14442;
assign w14444 = pi43 & pi52;
assign w14445 = ~w14321 & ~w14444;
assign w14446 = pi44 & pi52;
assign w14447 = w14319 & w14446;
assign w14448 = ~w14445 & ~w14447;
assign w14449 = w14330 & ~w14448;
assign w14450 = ~w14330 & w14448;
assign w14451 = ~w14449 & ~w14450;
assign w14452 = w14443 & ~w14451;
assign w14453 = ~w14443 & w14451;
assign w14454 = ~w14452 & ~w14453;
assign w14455 = ~w14425 & w14454;
assign w14456 = w14425 & ~w14454;
assign w14457 = ~w14455 & ~w14456;
assign w14458 = w14318 & ~w14320;
assign w14459 = ~w14322 & ~w14458;
assign w14460 = pi37 & pi58;
assign w14461 = pi40 & pi55;
assign w14462 = pi38 & pi57;
assign w14463 = ~w14461 & ~w14462;
assign w14464 = w14461 & w14462;
assign w14465 = ~w14463 & ~w14464;
assign w14466 = w14460 & ~w14465;
assign w14467 = ~w14460 & w14465;
assign w14468 = ~w14466 & ~w14467;
assign w14469 = ~w14459 & ~w14468;
assign w14470 = w14459 & w14468;
assign w14471 = ~w14469 & ~w14470;
assign w14472 = pi41 & pi54;
assign w14473 = pi34 & pi61;
assign w14474 = ~w8302 & ~w14473;
assign w14475 = w8302 & w14473;
assign w14476 = ~w14474 & ~w14475;
assign w14477 = w14472 & ~w14476;
assign w14478 = ~w14472 & w14476;
assign w14479 = ~w14477 & ~w14478;
assign w14480 = w14471 & ~w14479;
assign w14481 = ~w14471 & w14479;
assign w14482 = ~w14480 & ~w14481;
assign w14483 = ~w14457 & ~w14482;
assign w14484 = w14457 & w14482;
assign w14485 = ~w14483 & ~w14484;
assign w14486 = ~w14275 & ~w14277;
assign w14487 = ~w8301 & ~w14358;
assign w14488 = ~w14357 & ~w14487;
assign w14489 = ~w14366 & ~w14370;
assign w14490 = ~w14369 & ~w14489;
assign w14491 = w14488 & w14490;
assign w14492 = ~w14488 & ~w14490;
assign w14493 = ~w14491 & ~w14492;
assign w14494 = w14327 & ~w14329;
assign w14495 = ~w14331 & ~w14494;
assign w14496 = ~w14493 & w14495;
assign w14497 = w14493 & ~w14495;
assign w14498 = ~w14496 & ~w14497;
assign w14499 = ~w14336 & ~w14348;
assign w14500 = ~w14363 & ~w14375;
assign w14501 = ~w14499 & ~w14500;
assign w14502 = w14499 & w14500;
assign w14503 = ~w14501 & ~w14502;
assign w14504 = w14498 & w14503;
assign w14505 = ~w14498 & ~w14503;
assign w14506 = ~w14504 & ~w14505;
assign w14507 = ~w14486 & w14506;
assign w14508 = w14486 & ~w14506;
assign w14509 = ~w14507 & ~w14508;
assign w14510 = w14485 & w14509;
assign w14511 = ~w14485 & ~w14509;
assign w14512 = ~w14510 & ~w14511;
assign w14513 = ~w14424 & ~w14512;
assign w14514 = w14424 & w14512;
assign w14515 = ~w14513 & ~w14514;
assign w14516 = ~w14280 & ~w14385;
assign w14517 = w14515 & ~w14516;
assign w14518 = ~w14515 & w14516;
assign w14519 = ~w14517 & ~w14518;
assign w14520 = ~w14257 & ~w14388;
assign w14521 = (w12329 & w17501) | (w12329 & w17502) | (w17501 & w17502);
assign w14522 = (~w12329 & w17503) | (~w12329 & w17504) | (w17503 & w17504);
assign w14523 = ~w14521 & ~w14522;
assign w14524 = ~w14389 & ~w14517;
assign w14525 = ~w14422 & ~w14514;
assign w14526 = ~w14417 & ~w14419;
assign w14527 = ~pi47 & ~w14436;
assign w14528 = pi48 & ~w14527;
assign w14529 = w14426 & ~w14429;
assign w14530 = ~w14431 & ~w14529;
assign w14531 = w14528 & ~w14530;
assign w14532 = ~w14528 & w14530;
assign w14533 = ~w14531 & ~w14532;
assign w14534 = w14330 & ~w14445;
assign w14535 = ~w14447 & ~w14534;
assign w14536 = ~w14533 & w14535;
assign w14537 = w14533 & ~w14535;
assign w14538 = ~w14536 & ~w14537;
assign w14539 = ~w14469 & ~w14480;
assign w14540 = ~w14441 & ~w14452;
assign w14541 = ~w14539 & ~w14540;
assign w14542 = w14539 & w14540;
assign w14543 = ~w14541 & ~w14542;
assign w14544 = w14538 & w14543;
assign w14545 = ~w14538 & ~w14543;
assign w14546 = ~w14544 & ~w14545;
assign w14547 = ~w14526 & w14546;
assign w14548 = w14526 & ~w14546;
assign w14549 = ~w14547 & ~w14548;
assign w14550 = ~w14491 & ~w14497;
assign w14551 = pi33 & pi63;
assign w14552 = pi35 & pi61;
assign w14553 = pi34 & pi62;
assign w14554 = ~w14552 & ~w14553;
assign w14555 = pi35 & pi62;
assign w14556 = w14473 & w14555;
assign w14557 = ~w14554 & ~w14556;
assign w14558 = w14551 & ~w14557;
assign w14559 = ~w14551 & w14557;
assign w14560 = ~w14558 & ~w14559;
assign w14561 = pi41 & pi55;
assign w14562 = pi42 & pi54;
assign w14563 = pi43 & pi53;
assign w14564 = ~w14562 & ~w14563;
assign w14565 = pi43 & pi54;
assign w14566 = w14330 & w14565;
assign w14567 = ~w14564 & ~w14566;
assign w14568 = w14561 & ~w14567;
assign w14569 = ~w14561 & w14567;
assign w14570 = ~w14568 & ~w14569;
assign w14571 = ~w14560 & ~w14570;
assign w14572 = w14560 & w14570;
assign w14573 = ~w14571 & ~w14572;
assign w14574 = w14550 & ~w14573;
assign w14575 = ~w14550 & w14573;
assign w14576 = ~w14574 & ~w14575;
assign w14577 = ~w14401 & ~w14405;
assign w14578 = ~w14472 & ~w14475;
assign w14579 = ~w14474 & ~w14578;
assign w14580 = ~w14460 & ~w14464;
assign w14581 = ~w14463 & ~w14580;
assign w14582 = w14579 & w14581;
assign w14583 = ~w14579 & ~w14581;
assign w14584 = ~w14582 & ~w14583;
assign w14585 = w14577 & ~w14584;
assign w14586 = ~w14577 & w14584;
assign w14587 = ~w14585 & ~w14586;
assign w14588 = ~w14409 & ~w14413;
assign w14589 = ~w14587 & w14588;
assign w14590 = w14587 & ~w14588;
assign w14591 = ~w14589 & ~w14590;
assign w14592 = w14576 & w14591;
assign w14593 = ~w14576 & ~w14591;
assign w14594 = ~w14592 & ~w14593;
assign w14595 = w14549 & w14594;
assign w14596 = ~w14549 & ~w14594;
assign w14597 = ~w14595 & ~w14596;
assign w14598 = ~w14507 & ~w14510;
assign w14599 = ~w14455 & ~w14484;
assign w14600 = ~w14501 & ~w14504;
assign w14601 = pi39 & pi57;
assign w14602 = pi38 & pi58;
assign w14603 = ~w14601 & ~w14602;
assign w14604 = pi39 & pi58;
assign w14605 = w14462 & w14604;
assign w14606 = ~w14603 & ~w14605;
assign w14607 = w14446 & ~w14606;
assign w14608 = ~w14446 & w14606;
assign w14609 = ~w14607 & ~w14608;
assign w14610 = pi37 & pi59;
assign w14611 = pi40 & pi56;
assign w14612 = ~w14610 & ~w14611;
assign w14613 = w14610 & w14611;
assign w14614 = ~w14612 & ~w14613;
assign w14615 = w14400 & ~w14614;
assign w14616 = ~w14400 & w14614;
assign w14617 = ~w14615 & ~w14616;
assign w14618 = ~w14609 & ~w14617;
assign w14619 = w14609 & w14617;
assign w14620 = ~w14618 & ~w14619;
assign w14621 = pi45 & pi51;
assign w14622 = pi47 & pi49;
assign w14623 = ~w14430 & ~w14622;
assign w14624 = pi47 & pi50;
assign w14625 = w14427 & w14624;
assign w14626 = ~w14623 & ~w14625;
assign w14627 = w14621 & ~w14626;
assign w14628 = ~w14621 & w14626;
assign w14629 = ~w14627 & ~w14628;
assign w14630 = w14620 & ~w14629;
assign w14631 = ~w14620 & w14629;
assign w14632 = ~w14630 & ~w14631;
assign w14633 = ~w14600 & w14632;
assign w14634 = w14600 & ~w14632;
assign w14635 = ~w14633 & ~w14634;
assign w14636 = ~w14599 & w14635;
assign w14637 = w14599 & ~w14635;
assign w14638 = ~w14636 & ~w14637;
assign w14639 = ~w14598 & w14638;
assign w14640 = w14598 & ~w14638;
assign w14641 = ~w14639 & ~w14640;
assign w14642 = w14597 & w14641;
assign w14643 = ~w14597 & ~w14641;
assign w14644 = ~w14642 & ~w14643;
assign w14645 = ~w14525 & w14644;
assign w14646 = w14525 & ~w14644;
assign w14647 = ~w14645 & ~w14646;
assign w14648 = (w11122 & w17656) | (w11122 & w17657) | (w17656 & w17657);
assign w14649 = (~w11122 & w17658) | (~w11122 & w17659) | (w17658 & w17659);
assign w14650 = ~w14648 & ~w14649;
assign w14651 = ~w14639 & ~w14642;
assign w14652 = ~w14633 & ~w14636;
assign w14653 = pi36 & pi61;
assign w14654 = w14621 & ~w14623;
assign w14655 = (w14653 & w14654) | (w14653 & w16781) | (w14654 & w16781);
assign w14656 = ~w14654 & w16782;
assign w14657 = ~w14655 & ~w14656;
assign w14658 = w14446 & ~w14603;
assign w14659 = ~w14605 & ~w14658;
assign w14660 = ~w14657 & w14659;
assign w14661 = w14657 & ~w14659;
assign w14662 = ~w14660 & ~w14661;
assign w14663 = ~w14618 & ~w14630;
assign w14664 = ~w14582 & ~w14586;
assign w14665 = ~w14663 & ~w14664;
assign w14666 = w14663 & w14664;
assign w14667 = ~w14665 & ~w14666;
assign w14668 = w14662 & w14667;
assign w14669 = ~w14662 & ~w14667;
assign w14670 = ~w14668 & ~w14669;
assign w14671 = (~w14531 & ~w14533) | (~w14531 & w16783) | (~w14533 & w16783);
assign w14672 = pi40 & pi57;
assign w14673 = pi46 & pi51;
assign w14674 = ~w14624 & ~w14673;
assign w14675 = pi47 & pi51;
assign w14676 = w14430 & w14675;
assign w14677 = ~w14674 & ~w14676;
assign w14678 = w14672 & ~w14677;
assign w14679 = ~w14672 & w14677;
assign w14680 = ~w14678 & ~w14679;
assign w14681 = ~pi48 & pi49;
assign w14682 = w14555 & ~w14681;
assign w14683 = ~w14555 & w14681;
assign w14684 = ~w14682 & ~w14683;
assign w14685 = ~w14680 & ~w14684;
assign w14686 = w14680 & w14684;
assign w14687 = ~w14685 & ~w14686;
assign w14688 = w14671 & ~w14687;
assign w14689 = ~w14671 & w14687;
assign w14690 = ~w14688 & ~w14689;
assign w14691 = ~w14400 & ~w14613;
assign w14692 = ~w14612 & ~w14691;
assign w14693 = w14551 & ~w14554;
assign w14694 = ~w14556 & ~w14693;
assign w14695 = w14692 & ~w14694;
assign w14696 = ~w14692 & w14694;
assign w14697 = ~w14695 & ~w14696;
assign w14698 = w14561 & ~w14564;
assign w14699 = ~w14566 & ~w14698;
assign w14700 = ~w14697 & w14699;
assign w14701 = w14697 & ~w14699;
assign w14702 = ~w14700 & ~w14701;
assign w14703 = ~w14571 & ~w14575;
assign w14704 = ~w14702 & w14703;
assign w14705 = w14702 & ~w14703;
assign w14706 = ~w14704 & ~w14705;
assign w14707 = w14690 & w14706;
assign w14708 = ~w14690 & ~w14706;
assign w14709 = ~w14707 & ~w14708;
assign w14710 = w14670 & w14709;
assign w14711 = ~w14670 & ~w14709;
assign w14712 = ~w14710 & ~w14711;
assign w14713 = w14652 & ~w14712;
assign w14714 = ~w14652 & w14712;
assign w14715 = ~w14713 & ~w14714;
assign w14716 = ~w14547 & ~w14595;
assign w14717 = ~w14590 & ~w14592;
assign w14718 = ~w14541 & ~w14544;
assign w14719 = pi37 & pi60;
assign w14720 = pi38 & pi59;
assign w14721 = ~w14604 & ~w14720;
assign w14722 = pi39 & pi59;
assign w14723 = w14602 & w14722;
assign w14724 = ~w14721 & ~w14723;
assign w14725 = w14719 & ~w14724;
assign w14726 = ~w14719 & w14724;
assign w14727 = ~w14725 & ~w14726;
assign w14728 = pi41 & pi56;
assign w14729 = pi34 & pi63;
assign w14730 = pi42 & pi55;
assign w14731 = ~w14729 & ~w14730;
assign w14732 = w14729 & w14730;
assign w14733 = ~w14731 & ~w14732;
assign w14734 = w14728 & ~w14733;
assign w14735 = ~w14728 & w14733;
assign w14736 = ~w14734 & ~w14735;
assign w14737 = ~w14727 & ~w14736;
assign w14738 = w14727 & w14736;
assign w14739 = ~w14737 & ~w14738;
assign w14740 = pi45 & pi52;
assign w14741 = pi44 & pi53;
assign w14742 = ~w14740 & ~w14741;
assign w14743 = pi45 & pi53;
assign w14744 = w14446 & w14743;
assign w14745 = ~w14742 & ~w14744;
assign w14746 = w14565 & ~w14745;
assign w14747 = ~w14565 & w14745;
assign w14748 = ~w14746 & ~w14747;
assign w14749 = w14739 & ~w14748;
assign w14750 = ~w14739 & w14748;
assign w14751 = ~w14749 & ~w14750;
assign w14752 = ~w14718 & w14751;
assign w14753 = w14718 & ~w14751;
assign w14754 = ~w14752 & ~w14753;
assign w14755 = ~w14717 & w14754;
assign w14756 = w14717 & ~w14754;
assign w14757 = ~w14755 & ~w14756;
assign w14758 = ~w14716 & w14757;
assign w14759 = w14716 & ~w14757;
assign w14760 = ~w14758 & ~w14759;
assign w14761 = w14715 & w14760;
assign w14762 = ~w14715 & ~w14760;
assign w14763 = ~w14761 & ~w14762;
assign w14764 = ~w14651 & w14763;
assign w14765 = w14651 & ~w14763;
assign w14766 = ~w14764 & ~w14765;
assign w14767 = (~w12329 & w17505) | (~w12329 & w17506) | (w17505 & w17506);
assign w14768 = (w12329 & w17507) | (w12329 & w17508) | (w17507 & w17508);
assign w14769 = ~w14767 & ~w14768;
assign w14770 = ~w14758 & ~w14761;
assign w14771 = ~w14710 & ~w14714;
assign w14772 = ~w14705 & ~w14707;
assign w14773 = pi44 & pi54;
assign w14774 = pi43 & pi55;
assign w14775 = ~w14773 & ~w14774;
assign w14776 = pi44 & pi55;
assign w14777 = w14565 & w14776;
assign w14778 = ~w14775 & ~w14777;
assign w14779 = pi35 & pi63;
assign w14780 = ~w14778 & w14779;
assign w14781 = w14778 & ~w14779;
assign w14782 = ~w14780 & ~w14781;
assign w14783 = w14672 & ~w14674;
assign w14784 = ~w14676 & ~w14783;
assign w14785 = ~w14782 & ~w14784;
assign w14786 = w14782 & w14784;
assign w14787 = ~w14785 & ~w14786;
assign w14788 = pi38 & pi60;
assign w14789 = pi42 & pi56;
assign w14790 = pi41 & pi57;
assign w14791 = ~w14789 & ~w14790;
assign w14792 = pi42 & pi57;
assign w14793 = w14728 & w14792;
assign w14794 = ~w14791 & ~w14793;
assign w14795 = w14788 & ~w14794;
assign w14796 = ~w14788 & w14794;
assign w14797 = ~w14795 & ~w14796;
assign w14798 = ~w14787 & w14797;
assign w14799 = w14787 & ~w14797;
assign w14800 = ~w14798 & ~w14799;
assign w14801 = ~w14665 & ~w14668;
assign w14802 = w14800 & ~w14801;
assign w14803 = ~w14800 & w14801;
assign w14804 = ~w14802 & ~w14803;
assign w14805 = ~w14772 & w14804;
assign w14806 = w14772 & ~w14804;
assign w14807 = ~w14805 & ~w14806;
assign w14808 = ~w14771 & w14807;
assign w14809 = w14771 & ~w14807;
assign w14810 = ~w14808 & ~w14809;
assign w14811 = ~w14752 & ~w14755;
assign w14812 = (~w14737 & ~w14739) | (~w14737 & w16963) | (~w14739 & w16963);
assign w14813 = (~w14695 & ~w14697) | (~w14695 & w16784) | (~w14697 & w16784);
assign w14814 = (~w14655 & ~w14657) | (~w14655 & w16964) | (~w14657 & w16964);
assign w14815 = ~w14813 & ~w14814;
assign w14816 = w14813 & w14814;
assign w14817 = ~w14815 & ~w14816;
assign w14818 = w14812 & ~w14817;
assign w14819 = ~w14812 & w14817;
assign w14820 = ~w14818 & ~w14819;
assign w14821 = ~w14728 & ~w14732;
assign w14822 = ~w14731 & ~w14821;
assign w14823 = w14719 & ~w14721;
assign w14824 = ~w14723 & ~w14823;
assign w14825 = w14822 & ~w14824;
assign w14826 = ~w14822 & w14824;
assign w14827 = ~w14825 & ~w14826;
assign w14828 = w14565 & ~w14742;
assign w14829 = ~w14744 & ~w14828;
assign w14830 = ~w14827 & w14829;
assign w14831 = w14827 & ~w14829;
assign w14832 = ~w14830 & ~w14831;
assign w14833 = ~w14685 & ~w14689;
assign w14834 = ~w14832 & w14833;
assign w14835 = w14832 & ~w14833;
assign w14836 = ~w14834 & ~w14835;
assign w14837 = pi36 & pi62;
assign w14838 = pi37 & pi61;
assign w14839 = ~w14837 & ~w14838;
assign w14840 = pi37 & pi62;
assign w14841 = w14653 & w14840;
assign w14842 = ~w14839 & ~w14841;
assign w14843 = (pi49 & w14555) | (pi49 & w16965) | (w14555 & w16965);
assign w14844 = w14842 & w14843;
assign w14845 = ~w14842 & ~w14843;
assign w14846 = ~w14844 & ~w14845;
assign w14847 = pi46 & pi52;
assign w14848 = pi48 & pi50;
assign w14849 = ~w14675 & ~w14848;
assign w14850 = pi48 & pi51;
assign w14851 = w14624 & w14850;
assign w14852 = ~w14849 & ~w14851;
assign w14853 = w14847 & ~w14852;
assign w14854 = ~w14847 & w14852;
assign w14855 = ~w14853 & ~w14854;
assign w14856 = pi40 & pi58;
assign w14857 = ~w14722 & ~w14856;
assign w14858 = pi40 & pi59;
assign w14859 = w14604 & w14858;
assign w14860 = ~w14857 & ~w14859;
assign w14861 = w14743 & ~w14860;
assign w14862 = ~w14743 & w14860;
assign w14863 = ~w14861 & ~w14862;
assign w14864 = ~w14855 & ~w14863;
assign w14865 = w14855 & w14863;
assign w14866 = ~w14864 & ~w14865;
assign w14867 = w14846 & w14866;
assign w14868 = ~w14846 & ~w14866;
assign w14869 = ~w14867 & ~w14868;
assign w14870 = ~w14836 & ~w14869;
assign w14871 = w14836 & w14869;
assign w14872 = ~w14870 & ~w14871;
assign w14873 = ~w14820 & ~w14872;
assign w14874 = w14820 & w14872;
assign w14875 = ~w14873 & ~w14874;
assign w14876 = w14811 & ~w14875;
assign w14877 = ~w14811 & w14875;
assign w14878 = ~w14876 & ~w14877;
assign w14879 = w14810 & w14878;
assign w14880 = ~w14810 & ~w14878;
assign w14881 = ~w14879 & ~w14880;
assign w14882 = w14770 & ~w14881;
assign w14883 = ~w14770 & w14881;
assign w14884 = ~w14882 & ~w14883;
assign w14885 = ~w14646 & ~w14765;
assign w14886 = (w12329 & w17509) | (w12329 & w17510) | (w17509 & w17510);
assign w14887 = (~w12329 & w17511) | (~w12329 & w17512) | (w17511 & w17512);
assign w14888 = ~w14886 & ~w14887;
assign w14889 = ~w14808 & ~w14879;
assign w14890 = ~w14802 & ~w14805;
assign w14891 = (~w14785 & ~w14787) | (~w14785 & w16966) | (~w14787 & w16966);
assign w14892 = (~w14825 & ~w14827) | (~w14825 & w16785) | (~w14827 & w16785);
assign w14893 = ~pi49 & pi50;
assign w14894 = w14840 & ~w14893;
assign w14895 = ~w14840 & w14893;
assign w14896 = ~w14894 & ~w14895;
assign w14897 = ~w14892 & ~w14896;
assign w14898 = w14892 & w14896;
assign w14899 = ~w14897 & ~w14898;
assign w14900 = w14891 & ~w14899;
assign w14901 = ~w14891 & w14899;
assign w14902 = ~w14900 & ~w14901;
assign w14903 = (~w14841 & ~w14842) | (~w14841 & w16967) | (~w14842 & w16967);
assign w14904 = w14788 & ~w14791;
assign w14905 = ~w14793 & ~w14904;
assign w14906 = ~w14903 & ~w14905;
assign w14907 = w14903 & w14905;
assign w14908 = ~w14906 & ~w14907;
assign w14909 = pi36 & pi63;
assign w14910 = pi39 & pi60;
assign w14911 = pi38 & pi61;
assign w14912 = ~w14910 & ~w14911;
assign w14913 = pi39 & pi61;
assign w14914 = w14788 & w14913;
assign w14915 = ~w14912 & ~w14914;
assign w14916 = w14909 & ~w14915;
assign w14917 = ~w14909 & w14915;
assign w14918 = ~w14916 & ~w14917;
assign w14919 = ~w14908 & w14918;
assign w14920 = w14908 & ~w14918;
assign w14921 = ~w14919 & ~w14920;
assign w14922 = w14743 & ~w14857;
assign w14923 = ~w14859 & ~w14922;
assign w14924 = w14847 & ~w14849;
assign w14925 = ~w14851 & ~w14924;
assign w14926 = ~w14923 & ~w14925;
assign w14927 = w14923 & w14925;
assign w14928 = ~w14926 & ~w14927;
assign w14929 = ~w14775 & w14779;
assign w14930 = ~w14777 & ~w14929;
assign w14931 = ~w14928 & w14930;
assign w14932 = w14928 & ~w14930;
assign w14933 = ~w14931 & ~w14932;
assign w14934 = (~w14864 & ~w14866) | (~w14864 & w16968) | (~w14866 & w16968);
assign w14935 = ~w14933 & w14934;
assign w14936 = w14933 & ~w14934;
assign w14937 = ~w14935 & ~w14936;
assign w14938 = w14921 & w14937;
assign w14939 = ~w14921 & ~w14937;
assign w14940 = ~w14938 & ~w14939;
assign w14941 = ~w14902 & ~w14940;
assign w14942 = w14902 & w14940;
assign w14943 = ~w14941 & ~w14942;
assign w14944 = ~w14890 & w14943;
assign w14945 = w14890 & ~w14943;
assign w14946 = ~w14944 & ~w14945;
assign w14947 = (~w14835 & ~w14836) | (~w14835 & w16969) | (~w14836 & w16969);
assign w14948 = (~w14815 & ~w14817) | (~w14815 & w16970) | (~w14817 & w16970);
assign w14949 = pi45 & pi54;
assign w14950 = pi47 & pi52;
assign w14951 = pi46 & pi53;
assign w14952 = ~w14950 & ~w14951;
assign w14953 = pi47 & pi53;
assign w14954 = w14847 & w14953;
assign w14955 = ~w14952 & ~w14954;
assign w14956 = w14949 & ~w14955;
assign w14957 = ~w14949 & w14955;
assign w14958 = ~w14956 & ~w14957;
assign w14959 = pi41 & pi58;
assign w14960 = ~w14776 & ~w14959;
assign w14961 = w14776 & w14959;
assign w14962 = ~w14960 & ~w14961;
assign w14963 = w14858 & ~w14962;
assign w14964 = ~w14858 & w14962;
assign w14965 = ~w14963 & ~w14964;
assign w14966 = ~w14958 & ~w14965;
assign w14967 = w14958 & w14965;
assign w14968 = ~w14966 & ~w14967;
assign w14969 = pi43 & pi56;
assign w14970 = ~w14792 & ~w14969;
assign w14971 = pi43 & pi57;
assign w14972 = w14789 & w14971;
assign w14973 = ~w14970 & ~w14972;
assign w14974 = w14850 & ~w14973;
assign w14975 = ~w14850 & w14973;
assign w14976 = ~w14974 & ~w14975;
assign w14977 = w14968 & ~w14976;
assign w14978 = ~w14968 & w14976;
assign w14979 = ~w14977 & ~w14978;
assign w14980 = ~w14948 & w14979;
assign w14981 = w14948 & ~w14979;
assign w14982 = ~w14980 & ~w14981;
assign w14983 = w14947 & ~w14982;
assign w14984 = ~w14947 & w14982;
assign w14985 = ~w14983 & ~w14984;
assign w14986 = ~w14874 & ~w14877;
assign w14987 = w14985 & ~w14986;
assign w14988 = ~w14985 & w14986;
assign w14989 = ~w14987 & ~w14988;
assign w14990 = w14946 & w14989;
assign w14991 = ~w14946 & ~w14989;
assign w14992 = ~w14990 & ~w14991;
assign w14993 = ~w14889 & w14992;
assign w14994 = w14889 & ~w14992;
assign w14995 = ~w14993 & ~w14994;
assign w14996 = ~w14764 & ~w14883;
assign w14997 = (w11122 & w17660) | (w11122 & w17661) | (w17660 & w17661);
assign w14998 = (~w11122 & w17662) | (~w11122 & w17663) | (w17662 & w17663);
assign w14999 = ~w14997 & ~w14998;
assign w15000 = ~w14987 & ~w14990;
assign w15001 = (~w14906 & ~w14908) | (~w14906 & w17237) | (~w14908 & w17237);
assign w15002 = (~w14926 & ~w14928) | (~w14926 & w16786) | (~w14928 & w16786);
assign w15003 = pi49 & pi51;
assign w15004 = pi48 & pi52;
assign w15005 = ~w15003 & ~w15004;
assign w15006 = pi49 & pi52;
assign w15007 = w14850 & w15006;
assign w15008 = ~w15005 & ~w15007;
assign w15009 = w14953 & ~w15008;
assign w15010 = ~w14953 & w15008;
assign w15011 = ~w15009 & ~w15010;
assign w15012 = ~w15002 & ~w15011;
assign w15013 = w15002 & w15011;
assign w15014 = ~w15012 & ~w15013;
assign w15015 = w15001 & ~w15014;
assign w15016 = ~w15001 & w15014;
assign w15017 = ~w15015 & ~w15016;
assign w15018 = ~w14984 & w17238;
assign w15019 = (w15017 & w14984) | (w15017 & w17239) | (w14984 & w17239);
assign w15020 = ~w15018 & ~w15019;
assign w15021 = w14909 & ~w14912;
assign w15022 = ~w14914 & ~w15021;
assign w15023 = w14949 & ~w14952;
assign w15024 = ~w14954 & ~w15023;
assign w15025 = ~w15022 & ~w15024;
assign w15026 = w15022 & w15024;
assign w15027 = ~w15025 & ~w15026;
assign w15028 = ~w14858 & ~w14961;
assign w15029 = ~w14960 & ~w15028;
assign w15030 = ~w15027 & ~w15029;
assign w15031 = w15027 & w15029;
assign w15032 = ~w15030 & ~w15031;
assign w15033 = ~w14966 & ~w14977;
assign w15034 = ~w15032 & w15033;
assign w15035 = w15032 & ~w15033;
assign w15036 = ~w15034 & ~w15035;
assign w15037 = pi37 & pi63;
assign w15038 = ~pi49 & ~w14840;
assign w15039 = pi50 & ~w15038;
assign w15040 = w15037 & w15039;
assign w15041 = ~w15037 & ~w15039;
assign w15042 = ~w15040 & ~w15041;
assign w15043 = w14850 & ~w14970;
assign w15044 = ~w14972 & ~w15043;
assign w15045 = ~w15042 & w15044;
assign w15046 = w15042 & ~w15044;
assign w15047 = ~w15045 & ~w15046;
assign w15048 = w15036 & w15047;
assign w15049 = ~w15036 & ~w15047;
assign w15050 = ~w15048 & ~w15049;
assign w15051 = w15020 & w15050;
assign w15052 = ~w15020 & ~w15050;
assign w15053 = ~w15051 & ~w15052;
assign w15054 = ~w14942 & ~w14944;
assign w15055 = (~w14936 & ~w14937) | (~w14936 & w17240) | (~w14937 & w17240);
assign w15056 = (~w14897 & ~w14899) | (~w14897 & w16971) | (~w14899 & w16971);
assign w15057 = pi45 & pi55;
assign w15058 = pi44 & pi56;
assign w15059 = ~w15057 & ~w15058;
assign w15060 = pi45 & pi56;
assign w15061 = w14776 & w15060;
assign w15062 = ~w15059 & ~w15061;
assign w15063 = w14971 & ~w15062;
assign w15064 = ~w14971 & w15062;
assign w15065 = ~w15063 & ~w15064;
assign w15066 = pi38 & pi62;
assign w15067 = pi40 & pi60;
assign w15068 = ~w14913 & ~w15067;
assign w15069 = pi40 & pi61;
assign w15070 = w14910 & w15069;
assign w15071 = ~w15068 & ~w15070;
assign w15072 = w15066 & ~w15071;
assign w15073 = ~w15066 & w15071;
assign w15074 = ~w15072 & ~w15073;
assign w15075 = ~w15065 & ~w15074;
assign w15076 = w15065 & w15074;
assign w15077 = ~w15075 & ~w15076;
assign w15078 = pi46 & pi54;
assign w15079 = pi42 & pi58;
assign w15080 = pi41 & pi59;
assign w15081 = ~w15079 & ~w15080;
assign w15082 = pi42 & pi59;
assign w15083 = w14959 & w15082;
assign w15084 = ~w15081 & ~w15083;
assign w15085 = w15078 & ~w15084;
assign w15086 = ~w15078 & w15084;
assign w15087 = ~w15085 & ~w15086;
assign w15088 = w15077 & ~w15087;
assign w15089 = ~w15077 & w15087;
assign w15090 = ~w15088 & ~w15089;
assign w15091 = ~w15056 & w15090;
assign w15092 = w15056 & ~w15090;
assign w15093 = ~w15091 & ~w15092;
assign w15094 = ~w15055 & w15093;
assign w15095 = w15055 & ~w15093;
assign w15096 = ~w15094 & ~w15095;
assign w15097 = ~w15054 & w15096;
assign w15098 = w15054 & ~w15096;
assign w15099 = ~w15097 & ~w15098;
assign w15100 = w15053 & w15099;
assign w15101 = ~w15053 & ~w15099;
assign w15102 = ~w15100 & ~w15101;
assign w15103 = ~w15000 & w15102;
assign w15104 = w15000 & ~w15102;
assign w15105 = ~w15103 & ~w15104;
assign w15106 = (~w12329 & w17513) | (~w12329 & w17514) | (w17513 & w17514);
assign w15107 = (w12329 & w17515) | (w12329 & w17516) | (w17515 & w17516);
assign w15108 = ~w15106 & ~w15107;
assign w15109 = ~w14994 & ~w15104;
assign w15110 = ~w15097 & ~w15100;
assign w15111 = ~w15019 & ~w15051;
assign w15112 = (~w15012 & ~w15014) | (~w15012 & w16972) | (~w15014 & w16972);
assign w15113 = pi38 & pi63;
assign w15114 = pi47 & pi54;
assign w15115 = pi46 & pi55;
assign w15116 = ~w15114 & ~w15115;
assign w15117 = pi47 & pi55;
assign w15118 = w15078 & w15117;
assign w15119 = ~w15116 & ~w15118;
assign w15120 = w15113 & ~w15119;
assign w15121 = ~w15113 & w15119;
assign w15122 = ~w15120 & ~w15121;
assign w15123 = pi43 & pi58;
assign w15124 = ~w15060 & ~w15123;
assign w15125 = w15060 & w15123;
assign w15126 = ~w15124 & ~w15125;
assign w15127 = w15082 & ~w15126;
assign w15128 = ~w15082 & w15126;
assign w15129 = ~w15127 & ~w15128;
assign w15130 = ~w15122 & ~w15129;
assign w15131 = w15122 & w15129;
assign w15132 = ~w15130 & ~w15131;
assign w15133 = pi48 & pi53;
assign w15134 = pi44 & pi57;
assign w15135 = ~w15006 & ~w15134;
assign w15136 = w15006 & w15134;
assign w15137 = ~w15135 & ~w15136;
assign w15138 = w15133 & ~w15137;
assign w15139 = ~w15133 & w15137;
assign w15140 = ~w15138 & ~w15139;
assign w15141 = w15132 & ~w15140;
assign w15142 = ~w15132 & w15140;
assign w15143 = ~w15141 & ~w15142;
assign w15144 = ~w15112 & w15143;
assign w15145 = w15112 & ~w15143;
assign w15146 = ~w15144 & ~w15145;
assign w15147 = ~w15040 & ~w15046;
assign w15148 = pi41 & pi60;
assign w15149 = ~w15069 & ~w15148;
assign w15150 = pi41 & pi61;
assign w15151 = w15067 & w15150;
assign w15152 = ~w15149 & ~w15151;
assign w15153 = w14953 & ~w15005;
assign w15154 = ~w15007 & ~w15153;
assign w15155 = w15152 & ~w15154;
assign w15156 = ~w15152 & w15154;
assign w15157 = ~w15155 & ~w15156;
assign w15158 = pi39 & pi62;
assign w15159 = ~pi50 & pi51;
assign w15160 = w15158 & ~w15159;
assign w15161 = ~w15158 & w15159;
assign w15162 = ~w15160 & ~w15161;
assign w15163 = w15157 & ~w15162;
assign w15164 = ~w15157 & w15162;
assign w15165 = ~w15163 & ~w15164;
assign w15166 = ~w15147 & w15165;
assign w15167 = w15147 & ~w15165;
assign w15168 = ~w15166 & ~w15167;
assign w15169 = w15146 & w15168;
assign w15170 = ~w15146 & ~w15168;
assign w15171 = ~w15169 & ~w15170;
assign w15172 = ~w15111 & w15171;
assign w15173 = w15111 & ~w15171;
assign w15174 = ~w15172 & ~w15173;
assign w15175 = w15066 & ~w15068;
assign w15176 = ~w15070 & ~w15175;
assign w15177 = w15078 & ~w15081;
assign w15178 = ~w15083 & ~w15177;
assign w15179 = ~w15176 & ~w15178;
assign w15180 = w15176 & w15178;
assign w15181 = ~w15179 & ~w15180;
assign w15182 = w14971 & ~w15059;
assign w15183 = ~w15061 & ~w15182;
assign w15184 = ~w15181 & w15183;
assign w15185 = w15181 & ~w15183;
assign w15186 = ~w15184 & ~w15185;
assign w15187 = ~w15075 & ~w15088;
assign w15188 = ~w15025 & ~w15031;
assign w15189 = ~w15187 & ~w15188;
assign w15190 = w15187 & w15188;
assign w15191 = ~w15189 & ~w15190;
assign w15192 = w15186 & w15191;
assign w15193 = ~w15186 & ~w15191;
assign w15194 = ~w15192 & ~w15193;
assign w15195 = (~w15091 & ~w15093) | (~w15091 & w17245) | (~w15093 & w17245);
assign w15196 = ~w15035 & ~w15048;
assign w15197 = ~w15195 & ~w15196;
assign w15198 = w15195 & w15196;
assign w15199 = ~w15197 & ~w15198;
assign w15200 = w15194 & w15199;
assign w15201 = ~w15194 & ~w15199;
assign w15202 = ~w15200 & ~w15201;
assign w15203 = w15174 & w15202;
assign w15204 = ~w15174 & ~w15202;
assign w15205 = ~w15203 & ~w15204;
assign w15206 = ~w15110 & w15205;
assign w15207 = w15110 & ~w15205;
assign w15208 = ~w15206 & ~w15207;
assign w15209 = (w12329 & w17517) | (w12329 & w17518) | (w17517 & w17518);
assign w15210 = (~w12329 & w17519) | (~w12329 & w17520) | (w17519 & w17520);
assign w15211 = ~w15209 & ~w15210;
assign w15212 = ~w15103 & ~w15206;
assign w15213 = (~w10008 & w17521) | (~w10008 & w17522) | (w17521 & w17522);
assign w15214 = ~w15172 & ~w15203;
assign w15215 = ~w15197 & ~w15200;
assign w15216 = (~w15151 & w15154) | (~w15151 & w17248) | (w15154 & w17248);
assign w15217 = ~w15082 & ~w15125;
assign w15218 = ~w15124 & ~w15217;
assign w15219 = ~w15216 & w15218;
assign w15220 = w15216 & ~w15218;
assign w15221 = ~w15219 & ~w15220;
assign w15222 = pi39 & pi63;
assign w15223 = pi42 & pi60;
assign w15224 = ~w15150 & ~w15223;
assign w15225 = pi42 & pi61;
assign w15226 = w15148 & w15225;
assign w15227 = ~w15224 & ~w15226;
assign w15228 = w15222 & ~w15227;
assign w15229 = ~w15222 & w15227;
assign w15230 = ~w15228 & ~w15229;
assign w15231 = ~w15221 & w15230;
assign w15232 = w15221 & ~w15230;
assign w15233 = ~w15231 & ~w15232;
assign w15234 = (~w15163 & ~w15165) | (~w15163 & w17249) | (~w15165 & w17249);
assign w15235 = w15233 & ~w15234;
assign w15236 = ~w15233 & w15234;
assign w15237 = ~w15235 & ~w15236;
assign w15238 = pi40 & pi62;
assign w15239 = pi44 & pi58;
assign w15240 = pi43 & pi59;
assign w15241 = ~w15239 & ~w15240;
assign w15242 = pi44 & pi59;
assign w15243 = w15123 & w15242;
assign w15244 = ~w15241 & ~w15243;
assign w15245 = w15238 & ~w15244;
assign w15246 = ~w15238 & w15244;
assign w15247 = ~w15245 & ~w15246;
assign w15248 = pi45 & pi57;
assign w15249 = pi46 & pi56;
assign w15250 = ~w15117 & ~w15249;
assign w15251 = pi47 & pi56;
assign w15252 = w15115 & w15251;
assign w15253 = ~w15250 & ~w15252;
assign w15254 = w15248 & ~w15253;
assign w15255 = ~w15248 & w15253;
assign w15256 = ~w15254 & ~w15255;
assign w15257 = ~w15247 & ~w15256;
assign w15258 = w15247 & w15256;
assign w15259 = ~w15257 & ~w15258;
assign w15260 = pi48 & pi54;
assign w15261 = pi49 & pi53;
assign w15262 = pi50 & pi52;
assign w15263 = ~w15261 & ~w15262;
assign w15264 = pi50 & pi53;
assign w15265 = w15006 & w15264;
assign w15266 = ~w15263 & ~w15265;
assign w15267 = w15260 & ~w15266;
assign w15268 = ~w15260 & w15266;
assign w15269 = ~w15267 & ~w15268;
assign w15270 = w15259 & ~w15269;
assign w15271 = ~w15259 & w15269;
assign w15272 = ~w15270 & ~w15271;
assign w15273 = w15237 & w15272;
assign w15274 = ~w15237 & ~w15272;
assign w15275 = ~w15273 & ~w15274;
assign w15276 = ~w15215 & w15275;
assign w15277 = w15215 & ~w15275;
assign w15278 = ~w15276 & ~w15277;
assign w15279 = ~pi50 & ~w15158;
assign w15280 = pi51 & ~w15279;
assign w15281 = ~w15133 & ~w15136;
assign w15282 = ~w15135 & ~w15281;
assign w15283 = w15280 & w15282;
assign w15284 = ~w15280 & ~w15282;
assign w15285 = ~w15283 & ~w15284;
assign w15286 = w15113 & ~w15116;
assign w15287 = ~w15118 & ~w15286;
assign w15288 = ~w15285 & w15287;
assign w15289 = w15285 & ~w15287;
assign w15290 = ~w15288 & ~w15289;
assign w15291 = ~w15179 & ~w15185;
assign w15292 = ~w15290 & w15291;
assign w15293 = w15290 & ~w15291;
assign w15294 = ~w15292 & ~w15293;
assign w15295 = ~w15130 & ~w15141;
assign w15296 = ~w15294 & w15295;
assign w15297 = w15294 & ~w15295;
assign w15298 = ~w15296 & ~w15297;
assign w15299 = (~w15144 & ~w15146) | (~w15144 & w17250) | (~w15146 & w17250);
assign w15300 = ~w15189 & ~w15192;
assign w15301 = ~w15299 & ~w15300;
assign w15302 = w15299 & w15300;
assign w15303 = ~w15301 & ~w15302;
assign w15304 = w15298 & w15303;
assign w15305 = ~w15298 & ~w15303;
assign w15306 = ~w15304 & ~w15305;
assign w15307 = w15278 & w15306;
assign w15308 = ~w15278 & ~w15306;
assign w15309 = ~w15307 & ~w15308;
assign w15310 = w15214 & ~w15309;
assign w15311 = ~w15214 & w15309;
assign w15312 = ~w15310 & ~w15311;
assign w15313 = (~w10008 & w17865) | (~w10008 & w17866) | (w17865 & w17866);
assign w15314 = (w10008 & w17867) | (w10008 & w17868) | (w17867 & w17868);
assign w15315 = ~w15313 & ~w15314;
assign w15316 = ~w15257 & ~w15270;
assign w15317 = ~w15219 & ~w15232;
assign w15318 = ~w15283 & ~w15289;
assign w15319 = ~w15317 & ~w15318;
assign w15320 = w15317 & w15318;
assign w15321 = ~w15319 & ~w15320;
assign w15322 = w15316 & ~w15321;
assign w15323 = ~w15316 & w15321;
assign w15324 = ~w15322 & ~w15323;
assign w15325 = ~w15235 & ~w15273;
assign w15326 = ~w15293 & ~w15297;
assign w15327 = ~w15325 & ~w15326;
assign w15328 = w15325 & w15326;
assign w15329 = ~w15327 & ~w15328;
assign w15330 = w15324 & w15329;
assign w15331 = ~w15324 & ~w15329;
assign w15332 = ~w15330 & ~w15331;
assign w15333 = ~w15301 & ~w15304;
assign w15334 = pi40 & pi63;
assign w15335 = w15260 & ~w15263;
assign w15336 = ~w15265 & ~w15335;
assign w15337 = w15334 & ~w15336;
assign w15338 = ~w15334 & w15336;
assign w15339 = ~w15337 & ~w15338;
assign w15340 = w15248 & ~w15250;
assign w15341 = ~w15252 & ~w15340;
assign w15342 = ~w15339 & w15341;
assign w15343 = w15339 & ~w15341;
assign w15344 = ~w15342 & ~w15343;
assign w15345 = w15222 & ~w15224;
assign w15346 = ~w15226 & ~w15345;
assign w15347 = w15238 & ~w15241;
assign w15348 = ~w15243 & ~w15347;
assign w15349 = ~w15346 & ~w15348;
assign w15350 = w15346 & w15348;
assign w15351 = ~w15349 & ~w15350;
assign w15352 = pi45 & pi58;
assign w15353 = ~w15242 & ~w15352;
assign w15354 = pi45 & pi59;
assign w15355 = w15239 & w15354;
assign w15356 = ~w15353 & ~w15355;
assign w15357 = w15225 & ~w15356;
assign w15358 = ~w15225 & w15356;
assign w15359 = ~w15357 & ~w15358;
assign w15360 = ~w15351 & w15359;
assign w15361 = w15351 & ~w15359;
assign w15362 = ~w15360 & ~w15361;
assign w15363 = ~w15344 & ~w15362;
assign w15364 = w15344 & w15362;
assign w15365 = ~w15363 & ~w15364;
assign w15366 = pi43 & pi60;
assign w15367 = pi46 & pi57;
assign w15368 = ~w15251 & ~w15367;
assign w15369 = pi47 & pi57;
assign w15370 = w15249 & w15369;
assign w15371 = ~w15368 & ~w15370;
assign w15372 = w15366 & ~w15371;
assign w15373 = ~w15366 & w15371;
assign w15374 = ~w15372 & ~w15373;
assign w15375 = pi48 & pi55;
assign w15376 = pi49 & pi54;
assign w15377 = ~w15264 & ~w15376;
assign w15378 = pi50 & pi54;
assign w15379 = w15261 & w15378;
assign w15380 = ~w15377 & ~w15379;
assign w15381 = w15375 & ~w15380;
assign w15382 = ~w15375 & w15380;
assign w15383 = ~w15381 & ~w15382;
assign w15384 = ~w15374 & ~w15383;
assign w15385 = w15374 & w15383;
assign w15386 = ~w15384 & ~w15385;
assign w15387 = pi41 & pi62;
assign w15388 = ~pi51 & pi52;
assign w15389 = w15387 & ~w15388;
assign w15390 = ~w15387 & w15388;
assign w15391 = ~w15389 & ~w15390;
assign w15392 = w15386 & ~w15391;
assign w15393 = ~w15386 & w15391;
assign w15394 = ~w15392 & ~w15393;
assign w15395 = w15365 & w15394;
assign w15396 = ~w15365 & ~w15394;
assign w15397 = ~w15395 & ~w15396;
assign w15398 = ~w15333 & w15397;
assign w15399 = w15333 & ~w15397;
assign w15400 = ~w15398 & ~w15399;
assign w15401 = w15332 & w15400;
assign w15402 = ~w15332 & ~w15400;
assign w15403 = ~w15401 & ~w15402;
assign w15404 = ~w15276 & ~w15307;
assign w15405 = w15403 & ~w15404;
assign w15406 = ~w15403 & w15404;
assign w15407 = ~w15405 & ~w15406;
assign w15408 = (~w13978 & w17375) | (~w13978 & w17376) | (w17375 & w17376);
assign w15409 = (w13978 & w17377) | (w13978 & w17378) | (w17377 & w17378);
assign w15410 = ~w15408 & ~w15409;
assign w15411 = ~w15310 & ~w15406;
assign w15412 = ~w15398 & ~w15401;
assign w15413 = ~w15327 & ~w15330;
assign w15414 = w15366 & ~w15368;
assign w15415 = ~w15370 & ~w15414;
assign w15416 = w15375 & ~w15377;
assign w15417 = ~w15379 & ~w15416;
assign w15418 = ~w15415 & ~w15417;
assign w15419 = w15415 & w15417;
assign w15420 = ~w15418 & ~w15419;
assign w15421 = w15225 & ~w15353;
assign w15422 = ~w15355 & ~w15421;
assign w15423 = ~w15420 & w15422;
assign w15424 = w15420 & ~w15422;
assign w15425 = ~w15423 & ~w15424;
assign w15426 = ~w15384 & ~w15392;
assign w15427 = ~w15425 & w15426;
assign w15428 = w15425 & ~w15426;
assign w15429 = ~w15427 & ~w15428;
assign w15430 = pi46 & pi58;
assign w15431 = pi48 & pi56;
assign w15432 = ~w15369 & ~w15431;
assign w15433 = pi48 & pi57;
assign w15434 = w15251 & w15433;
assign w15435 = ~w15432 & ~w15434;
assign w15436 = w15430 & ~w15435;
assign w15437 = ~w15430 & w15435;
assign w15438 = ~w15436 & ~w15437;
assign w15439 = pi44 & pi60;
assign w15440 = pi43 & pi61;
assign w15441 = ~w15354 & ~w15440;
assign w15442 = w15354 & w15440;
assign w15443 = ~w15441 & ~w15442;
assign w15444 = w15439 & ~w15443;
assign w15445 = ~w15439 & w15443;
assign w15446 = ~w15444 & ~w15445;
assign w15447 = ~w15438 & ~w15446;
assign w15448 = w15438 & w15446;
assign w15449 = ~w15447 & ~w15448;
assign w15450 = pi49 & pi55;
assign w15451 = pi51 & pi53;
assign w15452 = ~w15378 & ~w15451;
assign w15453 = pi51 & pi54;
assign w15454 = w15264 & w15453;
assign w15455 = ~w15452 & ~w15454;
assign w15456 = w15450 & ~w15455;
assign w15457 = ~w15450 & w15455;
assign w15458 = ~w15456 & ~w15457;
assign w15459 = w15449 & ~w15458;
assign w15460 = ~w15449 & w15458;
assign w15461 = ~w15459 & ~w15460;
assign w15462 = w15429 & w15461;
assign w15463 = ~w15429 & ~w15461;
assign w15464 = ~w15462 & ~w15463;
assign w15465 = ~w15413 & w15464;
assign w15466 = w15413 & ~w15464;
assign w15467 = ~w15465 & ~w15466;
assign w15468 = ~w15337 & ~w15343;
assign w15469 = pi41 & pi63;
assign w15470 = pi42 & pi62;
assign w15471 = ~w15469 & ~w15470;
assign w15472 = pi42 & pi63;
assign w15473 = w15387 & w15472;
assign w15474 = ~w15471 & ~w15473;
assign w15475 = ~pi51 & ~w15387;
assign w15476 = pi52 & ~w15475;
assign w15477 = w15474 & w15476;
assign w15478 = ~w15474 & ~w15476;
assign w15479 = ~w15477 & ~w15478;
assign w15480 = ~w15468 & w15479;
assign w15481 = w15468 & ~w15479;
assign w15482 = ~w15480 & ~w15481;
assign w15483 = ~w15349 & ~w15361;
assign w15484 = ~w15482 & w15483;
assign w15485 = w15482 & ~w15483;
assign w15486 = ~w15484 & ~w15485;
assign w15487 = ~w15364 & ~w15395;
assign w15488 = ~w15319 & ~w15323;
assign w15489 = ~w15487 & ~w15488;
assign w15490 = w15487 & w15488;
assign w15491 = ~w15489 & ~w15490;
assign w15492 = w15486 & w15491;
assign w15493 = ~w15486 & ~w15491;
assign w15494 = ~w15492 & ~w15493;
assign w15495 = w15467 & w15494;
assign w15496 = ~w15467 & ~w15494;
assign w15497 = ~w15495 & ~w15496;
assign w15498 = ~w15412 & w15497;
assign w15499 = w15412 & ~w15497;
assign w15500 = ~w15498 & ~w15499;
assign w15501 = (w13978 & w17379) | (w13978 & w17380) | (w17379 & w17380);
assign w15502 = (~w13978 & w17381) | (~w13978 & w17382) | (w17381 & w17382);
assign w15503 = ~w15501 & ~w15502;
assign w15504 = w15430 & ~w15432;
assign w15505 = ~w15434 & ~w15504;
assign w15506 = w15450 & ~w15452;
assign w15507 = ~w15454 & ~w15506;
assign w15508 = ~w15505 & ~w15507;
assign w15509 = w15505 & w15507;
assign w15510 = ~w15508 & ~w15509;
assign w15511 = ~w15439 & ~w15442;
assign w15512 = ~w15441 & ~w15511;
assign w15513 = ~w15510 & ~w15512;
assign w15514 = w15510 & w15512;
assign w15515 = ~w15513 & ~w15514;
assign w15516 = ~w15447 & ~w15459;
assign w15517 = ~w15515 & w15516;
assign w15518 = w15515 & ~w15516;
assign w15519 = ~w15517 & ~w15518;
assign w15520 = ~w15480 & ~w15485;
assign w15521 = ~w15519 & w15520;
assign w15522 = w15519 & ~w15520;
assign w15523 = ~w15521 & ~w15522;
assign w15524 = ~w15489 & ~w15492;
assign w15525 = ~w15523 & w15524;
assign w15526 = w15523 & ~w15524;
assign w15527 = ~w15525 & ~w15526;
assign w15528 = ~w15428 & ~w15462;
assign w15529 = ~w15418 & ~w15424;
assign w15530 = pi49 & pi56;
assign w15531 = pi50 & pi55;
assign w15532 = ~w15453 & ~w15531;
assign w15533 = pi51 & pi55;
assign w15534 = w15378 & w15533;
assign w15535 = ~w15532 & ~w15534;
assign w15536 = w15530 & ~w15535;
assign w15537 = ~w15530 & w15535;
assign w15538 = ~w15536 & ~w15537;
assign w15539 = pi43 & pi62;
assign w15540 = ~pi52 & pi53;
assign w15541 = w15539 & ~w15540;
assign w15542 = ~w15539 & w15540;
assign w15543 = ~w15541 & ~w15542;
assign w15544 = ~w15538 & ~w15543;
assign w15545 = w15538 & w15543;
assign w15546 = ~w15544 & ~w15545;
assign w15547 = w15529 & ~w15546;
assign w15548 = ~w15529 & w15546;
assign w15549 = ~w15547 & ~w15548;
assign w15550 = ~w15473 & ~w15477;
assign w15551 = pi44 & pi61;
assign w15552 = pi45 & pi60;
assign w15553 = ~w15551 & ~w15552;
assign w15554 = pi45 & pi61;
assign w15555 = w15439 & w15554;
assign w15556 = ~w15553 & ~w15555;
assign w15557 = w15472 & ~w15556;
assign w15558 = ~w15472 & w15556;
assign w15559 = ~w15557 & ~w15558;
assign w15560 = ~w15550 & ~w15559;
assign w15561 = w15550 & w15559;
assign w15562 = ~w15560 & ~w15561;
assign w15563 = pi46 & pi59;
assign w15564 = pi47 & pi58;
assign w15565 = ~w15433 & ~w15564;
assign w15566 = pi48 & pi58;
assign w15567 = w15369 & w15566;
assign w15568 = ~w15565 & ~w15567;
assign w15569 = w15563 & ~w15568;
assign w15570 = ~w15563 & w15568;
assign w15571 = ~w15569 & ~w15570;
assign w15572 = w15562 & ~w15571;
assign w15573 = ~w15562 & w15571;
assign w15574 = ~w15572 & ~w15573;
assign w15575 = w15549 & w15574;
assign w15576 = ~w15549 & ~w15574;
assign w15577 = ~w15575 & ~w15576;
assign w15578 = ~w15528 & w15577;
assign w15579 = w15528 & ~w15577;
assign w15580 = ~w15578 & ~w15579;
assign w15581 = w15527 & w15580;
assign w15582 = ~w15527 & ~w15580;
assign w15583 = ~w15581 & ~w15582;
assign w15584 = ~w15465 & ~w15495;
assign w15585 = ~w15583 & w15584;
assign w15586 = w15583 & ~w15584;
assign w15587 = ~w15585 & ~w15586;
assign w15588 = ~w15405 & ~w15498;
assign w15589 = (~w12329 & w17523) | (~w12329 & w17524) | (w17523 & w17524);
assign w15590 = (w12329 & w17525) | (w12329 & w17526) | (w17525 & w17526);
assign w15591 = ~w15589 & ~w15590;
assign w15592 = ~w15526 & ~w15581;
assign w15593 = pi43 & pi63;
assign w15594 = ~pi52 & ~w15539;
assign w15595 = pi53 & ~w15594;
assign w15596 = w15593 & w15595;
assign w15597 = ~w15593 & ~w15595;
assign w15598 = ~w15596 & ~w15597;
assign w15599 = w15530 & ~w15532;
assign w15600 = ~w15534 & ~w15599;
assign w15601 = ~w15598 & w15600;
assign w15602 = w15598 & ~w15600;
assign w15603 = ~w15601 & ~w15602;
assign w15604 = ~w15560 & ~w15572;
assign w15605 = ~w15603 & w15604;
assign w15606 = w15603 & ~w15604;
assign w15607 = ~w15605 & ~w15606;
assign w15608 = ~w15544 & ~w15548;
assign w15609 = ~w15607 & w15608;
assign w15610 = w15607 & ~w15608;
assign w15611 = ~w15609 & ~w15610;
assign w15612 = ~w15575 & ~w15578;
assign w15613 = ~w15611 & w15612;
assign w15614 = w15611 & ~w15612;
assign w15615 = ~w15613 & ~w15614;
assign w15616 = ~w15518 & ~w15522;
assign w15617 = ~w15508 & ~w15514;
assign w15618 = pi47 & pi59;
assign w15619 = pi49 & pi57;
assign w15620 = ~w15566 & ~w15619;
assign w15621 = pi49 & pi58;
assign w15622 = w15433 & w15621;
assign w15623 = ~w15620 & ~w15622;
assign w15624 = w15618 & ~w15623;
assign w15625 = ~w15618 & w15623;
assign w15626 = ~w15624 & ~w15625;
assign w15627 = pi50 & pi56;
assign w15628 = pi52 & pi54;
assign w15629 = ~w15533 & ~w15628;
assign w15630 = pi52 & pi55;
assign w15631 = w15453 & w15630;
assign w15632 = ~w15629 & ~w15631;
assign w15633 = w15627 & ~w15632;
assign w15634 = ~w15627 & w15632;
assign w15635 = ~w15633 & ~w15634;
assign w15636 = ~w15626 & ~w15635;
assign w15637 = w15626 & w15635;
assign w15638 = ~w15636 & ~w15637;
assign w15639 = w15617 & ~w15638;
assign w15640 = ~w15617 & w15638;
assign w15641 = ~w15639 & ~w15640;
assign w15642 = w15472 & ~w15553;
assign w15643 = ~w15555 & ~w15642;
assign w15644 = w15563 & ~w15565;
assign w15645 = ~w15567 & ~w15644;
assign w15646 = ~w15643 & ~w15645;
assign w15647 = w15643 & w15645;
assign w15648 = ~w15646 & ~w15647;
assign w15649 = pi44 & pi62;
assign w15650 = pi46 & pi60;
assign w15651 = ~w15554 & ~w15650;
assign w15652 = pi46 & pi61;
assign w15653 = w15552 & w15652;
assign w15654 = ~w15651 & ~w15653;
assign w15655 = w15649 & ~w15654;
assign w15656 = ~w15649 & w15654;
assign w15657 = ~w15655 & ~w15656;
assign w15658 = ~w15648 & w15657;
assign w15659 = w15648 & ~w15657;
assign w15660 = ~w15658 & ~w15659;
assign w15661 = ~w15641 & ~w15660;
assign w15662 = w15641 & w15660;
assign w15663 = ~w15661 & ~w15662;
assign w15664 = w15616 & w15663;
assign w15665 = ~w15616 & ~w15663;
assign w15666 = ~w15664 & ~w15665;
assign w15667 = w15615 & ~w15666;
assign w15668 = ~w15615 & w15666;
assign w15669 = ~w15667 & ~w15668;
assign w15670 = ~w15592 & w15669;
assign w15671 = w15592 & ~w15669;
assign w15672 = ~w15670 & ~w15671;
assign w15673 = (~w13978 & w17383) | (~w13978 & w17384) | (w17383 & w17384);
assign w15674 = (w13978 & w17385) | (w13978 & w17386) | (w17385 & w17386);
assign w15675 = ~w15673 & ~w15674;
assign w15676 = ~w15585 & ~w15671;
assign w15677 = ~w15614 & ~w15667;
assign w15678 = ~w15606 & ~w15610;
assign w15679 = w15618 & ~w15620;
assign w15680 = ~w15622 & ~w15679;
assign w15681 = w15649 & ~w15651;
assign w15682 = ~w15653 & ~w15681;
assign w15683 = ~w15680 & ~w15682;
assign w15684 = w15680 & w15682;
assign w15685 = ~w15683 & ~w15684;
assign w15686 = pi48 & pi59;
assign w15687 = pi44 & pi63;
assign w15688 = ~w15621 & ~w15687;
assign w15689 = w15621 & w15687;
assign w15690 = ~w15688 & ~w15689;
assign w15691 = w15686 & ~w15690;
assign w15692 = ~w15686 & w15690;
assign w15693 = ~w15691 & ~w15692;
assign w15694 = ~w15685 & w15693;
assign w15695 = w15685 & ~w15693;
assign w15696 = ~w15694 & ~w15695;
assign w15697 = pi47 & pi60;
assign w15698 = ~w15652 & ~w15697;
assign w15699 = pi47 & pi61;
assign w15700 = w15650 & w15699;
assign w15701 = ~w15698 & ~w15700;
assign w15702 = w15627 & ~w15629;
assign w15703 = ~w15631 & ~w15702;
assign w15704 = w15701 & ~w15703;
assign w15705 = ~w15701 & w15703;
assign w15706 = ~w15704 & ~w15705;
assign w15707 = pi50 & pi57;
assign w15708 = pi51 & pi56;
assign w15709 = ~w15630 & ~w15708;
assign w15710 = pi52 & pi56;
assign w15711 = w15533 & w15710;
assign w15712 = ~w15709 & ~w15711;
assign w15713 = w15707 & ~w15712;
assign w15714 = ~w15707 & w15712;
assign w15715 = ~w15713 & ~w15714;
assign w15716 = pi45 & pi62;
assign w15717 = ~pi53 & pi54;
assign w15718 = w15716 & ~w15717;
assign w15719 = ~w15716 & w15717;
assign w15720 = ~w15718 & ~w15719;
assign w15721 = ~w15715 & ~w15720;
assign w15722 = w15715 & w15720;
assign w15723 = ~w15721 & ~w15722;
assign w15724 = w15706 & w15723;
assign w15725 = ~w15706 & ~w15723;
assign w15726 = ~w15724 & ~w15725;
assign w15727 = w15696 & w15726;
assign w15728 = ~w15696 & ~w15726;
assign w15729 = ~w15727 & ~w15728;
assign w15730 = w15678 & ~w15729;
assign w15731 = ~w15678 & w15729;
assign w15732 = ~w15730 & ~w15731;
assign w15733 = ~w15636 & ~w15640;
assign w15734 = ~w15646 & ~w15659;
assign w15735 = ~w15596 & ~w15602;
assign w15736 = ~w15734 & ~w15735;
assign w15737 = w15734 & w15735;
assign w15738 = ~w15736 & ~w15737;
assign w15739 = w15733 & ~w15738;
assign w15740 = ~w15733 & w15738;
assign w15741 = ~w15739 & ~w15740;
assign w15742 = ~w15661 & ~w15664;
assign w15743 = w15741 & w15742;
assign w15744 = ~w15741 & ~w15742;
assign w15745 = ~w15743 & ~w15744;
assign w15746 = w15732 & w15745;
assign w15747 = ~w15732 & ~w15745;
assign w15748 = ~w15746 & ~w15747;
assign w15749 = w15677 & ~w15748;
assign w15750 = ~w15677 & w15748;
assign w15751 = ~w15749 & ~w15750;
assign w15752 = (w13978 & w17387) | (w13978 & w17388) | (w17387 & w17388);
assign w15753 = (~w13978 & w17389) | (~w13978 & w17390) | (w17389 & w17390);
assign w15754 = ~w15752 & ~w15753;
assign w15755 = ~w15670 & ~w15750;
assign w15756 = ~w15743 & ~w15746;
assign w15757 = ~pi53 & ~w15716;
assign w15758 = pi54 & ~w15757;
assign w15759 = w15707 & ~w15709;
assign w15760 = ~w15711 & ~w15759;
assign w15761 = w15758 & ~w15760;
assign w15762 = ~w15758 & w15760;
assign w15763 = ~w15761 & ~w15762;
assign w15764 = ~w15686 & ~w15689;
assign w15765 = ~w15688 & ~w15764;
assign w15766 = ~w15763 & ~w15765;
assign w15767 = w15763 & w15765;
assign w15768 = ~w15766 & ~w15767;
assign w15769 = ~w15736 & ~w15740;
assign w15770 = ~w15768 & w15769;
assign w15771 = w15768 & ~w15769;
assign w15772 = ~w15770 & ~w15771;
assign w15773 = ~w15700 & ~w15704;
assign w15774 = pi45 & pi63;
assign w15775 = pi46 & pi62;
assign w15776 = ~w15699 & ~w15775;
assign w15777 = pi47 & pi62;
assign w15778 = w15652 & w15777;
assign w15779 = ~w15776 & ~w15778;
assign w15780 = w15774 & ~w15779;
assign w15781 = ~w15774 & w15779;
assign w15782 = ~w15780 & ~w15781;
assign w15783 = ~w15773 & ~w15782;
assign w15784 = w15773 & w15782;
assign w15785 = ~w15783 & ~w15784;
assign w15786 = pi48 & pi60;
assign w15787 = pi49 & pi59;
assign w15788 = pi50 & pi58;
assign w15789 = ~w15787 & ~w15788;
assign w15790 = pi50 & pi59;
assign w15791 = w15621 & w15790;
assign w15792 = ~w15789 & ~w15791;
assign w15793 = w15786 & ~w15792;
assign w15794 = ~w15786 & w15792;
assign w15795 = ~w15793 & ~w15794;
assign w15796 = w15785 & ~w15795;
assign w15797 = ~w15785 & w15795;
assign w15798 = ~w15796 & ~w15797;
assign w15799 = w15772 & w15798;
assign w15800 = ~w15772 & ~w15798;
assign w15801 = ~w15799 & ~w15800;
assign w15802 = ~w15727 & ~w15731;
assign w15803 = ~w15721 & ~w15724;
assign w15804 = ~w15683 & ~w15695;
assign w15805 = pi51 & pi57;
assign w15806 = pi53 & pi55;
assign w15807 = ~w15710 & ~w15806;
assign w15808 = pi53 & pi56;
assign w15809 = w15630 & w15808;
assign w15810 = ~w15807 & ~w15809;
assign w15811 = w15805 & ~w15810;
assign w15812 = ~w15805 & w15810;
assign w15813 = ~w15811 & ~w15812;
assign w15814 = ~w15804 & ~w15813;
assign w15815 = w15804 & w15813;
assign w15816 = ~w15814 & ~w15815;
assign w15817 = ~w15803 & w15816;
assign w15818 = w15803 & ~w15816;
assign w15819 = ~w15817 & ~w15818;
assign w15820 = ~w15802 & w15819;
assign w15821 = w15802 & ~w15819;
assign w15822 = ~w15820 & ~w15821;
assign w15823 = w15801 & w15822;
assign w15824 = ~w15801 & ~w15822;
assign w15825 = ~w15823 & ~w15824;
assign w15826 = w15756 & ~w15825;
assign w15827 = ~w15756 & w15825;
assign w15828 = ~w15826 & ~w15827;
assign w15829 = (~w12329 & w17527) | (~w12329 & w17528) | (w17527 & w17528);
assign w15830 = (w12329 & w17529) | (w12329 & w17530) | (w17529 & w17530);
assign w15831 = ~w15829 & ~w15830;
assign w15832 = ~w15820 & ~w15823;
assign w15833 = ~w15783 & ~w15796;
assign w15834 = ~w15761 & ~w15767;
assign w15835 = ~pi54 & pi55;
assign w15836 = w15777 & ~w15835;
assign w15837 = ~w15777 & w15835;
assign w15838 = ~w15836 & ~w15837;
assign w15839 = ~w15834 & ~w15838;
assign w15840 = w15834 & w15838;
assign w15841 = ~w15839 & ~w15840;
assign w15842 = w15833 & ~w15841;
assign w15843 = ~w15833 & w15841;
assign w15844 = ~w15842 & ~w15843;
assign w15845 = ~w15771 & ~w15799;
assign w15846 = ~w15844 & w15845;
assign w15847 = w15844 & ~w15845;
assign w15848 = ~w15846 & ~w15847;
assign w15849 = pi46 & pi63;
assign w15850 = w15805 & ~w15807;
assign w15851 = ~w15809 & ~w15850;
assign w15852 = w15849 & ~w15851;
assign w15853 = ~w15849 & w15851;
assign w15854 = ~w15852 & ~w15853;
assign w15855 = w15786 & ~w15789;
assign w15856 = ~w15791 & ~w15855;
assign w15857 = ~w15854 & w15856;
assign w15858 = w15854 & ~w15856;
assign w15859 = ~w15857 & ~w15858;
assign w15860 = ~w15814 & ~w15817;
assign w15861 = ~w15859 & w15860;
assign w15862 = w15859 & ~w15860;
assign w15863 = ~w15861 & ~w15862;
assign w15864 = pi48 & pi61;
assign w15865 = pi49 & pi60;
assign w15866 = ~w15790 & ~w15865;
assign w15867 = pi50 & pi60;
assign w15868 = w15787 & w15867;
assign w15869 = ~w15866 & ~w15868;
assign w15870 = w15864 & ~w15869;
assign w15871 = ~w15864 & w15869;
assign w15872 = ~w15870 & ~w15871;
assign w15873 = w15774 & ~w15776;
assign w15874 = ~w15778 & ~w15873;
assign w15875 = ~w15872 & ~w15874;
assign w15876 = w15872 & w15874;
assign w15877 = ~w15875 & ~w15876;
assign w15878 = pi51 & pi58;
assign w15879 = pi52 & pi57;
assign w15880 = ~w15808 & ~w15879;
assign w15881 = pi53 & pi57;
assign w15882 = w15710 & w15881;
assign w15883 = ~w15880 & ~w15882;
assign w15884 = w15878 & ~w15883;
assign w15885 = ~w15878 & w15883;
assign w15886 = ~w15884 & ~w15885;
assign w15887 = w15877 & ~w15886;
assign w15888 = ~w15877 & w15886;
assign w15889 = ~w15887 & ~w15888;
assign w15890 = w15863 & w15889;
assign w15891 = ~w15863 & ~w15889;
assign w15892 = ~w15890 & ~w15891;
assign w15893 = w15848 & w15892;
assign w15894 = ~w15848 & ~w15892;
assign w15895 = ~w15893 & ~w15894;
assign w15896 = ~w15832 & w15895;
assign w15897 = w15832 & ~w15895;
assign w15898 = ~w15896 & ~w15897;
assign w15899 = (~w13978 & w17391) | (~w13978 & w17392) | (w17391 & w17392);
assign w15900 = (w13978 & w17393) | (w13978 & w17394) | (w17393 & w17394);
assign w15901 = ~w15899 & ~w15900;
assign w15902 = ~w15826 & ~w15897;
assign w15903 = ~w15847 & ~w15893;
assign w15904 = ~w15839 & ~w15843;
assign w15905 = w15864 & ~w15866;
assign w15906 = ~w15868 & ~w15905;
assign w15907 = w15878 & ~w15880;
assign w15908 = ~w15882 & ~w15907;
assign w15909 = ~w15906 & ~w15908;
assign w15910 = w15906 & w15908;
assign w15911 = ~w15909 & ~w15910;
assign w15912 = pi49 & pi61;
assign w15913 = pi51 & pi59;
assign w15914 = ~w15867 & ~w15913;
assign w15915 = pi51 & pi60;
assign w15916 = w15790 & w15915;
assign w15917 = ~w15914 & ~w15916;
assign w15918 = w15912 & ~w15917;
assign w15919 = ~w15912 & w15917;
assign w15920 = ~w15918 & ~w15919;
assign w15921 = ~w15911 & w15920;
assign w15922 = w15911 & ~w15920;
assign w15923 = ~w15921 & ~w15922;
assign w15924 = ~w15875 & ~w15887;
assign w15925 = w15923 & ~w15924;
assign w15926 = ~w15923 & w15924;
assign w15927 = ~w15925 & ~w15926;
assign w15928 = w15904 & ~w15927;
assign w15929 = ~w15904 & w15927;
assign w15930 = ~w15928 & ~w15929;
assign w15931 = pi47 & pi63;
assign w15932 = pi48 & pi62;
assign w15933 = ~w15931 & ~w15932;
assign w15934 = pi48 & pi63;
assign w15935 = w15777 & w15934;
assign w15936 = ~w15933 & ~w15935;
assign w15937 = ~pi54 & ~w15777;
assign w15938 = pi55 & ~w15937;
assign w15939 = w15936 & w15938;
assign w15940 = ~w15936 & ~w15938;
assign w15941 = ~w15939 & ~w15940;
assign w15942 = pi52 & pi58;
assign w15943 = pi54 & pi56;
assign w15944 = ~w15881 & ~w15943;
assign w15945 = pi54 & pi57;
assign w15946 = w15808 & w15945;
assign w15947 = ~w15944 & ~w15946;
assign w15948 = w15942 & ~w15947;
assign w15949 = ~w15942 & w15947;
assign w15950 = ~w15948 & ~w15949;
assign w15951 = ~w15941 & w15950;
assign w15952 = w15941 & ~w15950;
assign w15953 = ~w15951 & ~w15952;
assign w15954 = ~w15852 & ~w15858;
assign w15955 = ~w15953 & w15954;
assign w15956 = w15953 & ~w15954;
assign w15957 = ~w15955 & ~w15956;
assign w15958 = ~w15862 & ~w15890;
assign w15959 = w15957 & ~w15958;
assign w15960 = ~w15957 & w15958;
assign w15961 = ~w15959 & ~w15960;
assign w15962 = w15930 & w15961;
assign w15963 = ~w15930 & ~w15961;
assign w15964 = ~w15962 & ~w15963;
assign w15965 = ~w15903 & w15964;
assign w15966 = w15903 & ~w15964;
assign w15967 = ~w15965 & ~w15966;
assign w15968 = (w13978 & w17395) | (w13978 & w17396) | (w17395 & w17396);
assign w15969 = (~w13978 & w17397) | (~w13978 & w17398) | (w17397 & w17398);
assign w15970 = ~w15968 & ~w15969;
assign w15971 = ~w15896 & ~w15965;
assign w15972 = ~w15959 & ~w15962;
assign w15973 = ~w15935 & ~w15939;
assign w15974 = w15912 & ~w15914;
assign w15975 = ~w15916 & ~w15974;
assign w15976 = w15942 & ~w15944;
assign w15977 = ~w15946 & ~w15976;
assign w15978 = ~w15975 & ~w15977;
assign w15979 = w15975 & w15977;
assign w15980 = ~w15978 & ~w15979;
assign w15981 = w15973 & ~w15980;
assign w15982 = ~w15973 & w15980;
assign w15983 = ~w15981 & ~w15982;
assign w15984 = ~w15909 & ~w15922;
assign w15985 = ~w15983 & w15984;
assign w15986 = w15983 & ~w15984;
assign w15987 = ~w15985 & ~w15986;
assign w15988 = ~w15952 & ~w15956;
assign w15989 = ~w15987 & w15988;
assign w15990 = w15987 & ~w15988;
assign w15991 = ~w15989 & ~w15990;
assign w15992 = ~w15925 & ~w15929;
assign w15993 = pi50 & pi61;
assign w15994 = ~w15915 & ~w15993;
assign w15995 = pi51 & pi61;
assign w15996 = w15867 & w15995;
assign w15997 = ~w15994 & ~w15996;
assign w15998 = w15934 & ~w15997;
assign w15999 = ~w15934 & w15997;
assign w16000 = ~w15998 & ~w15999;
assign w16001 = pi49 & pi62;
assign w16002 = ~pi55 & pi56;
assign w16003 = w16001 & ~w16002;
assign w16004 = ~w16001 & w16002;
assign w16005 = ~w16003 & ~w16004;
assign w16006 = ~w16000 & ~w16005;
assign w16007 = w16000 & w16005;
assign w16008 = ~w16006 & ~w16007;
assign w16009 = pi52 & pi59;
assign w16010 = pi53 & pi58;
assign w16011 = ~w15945 & ~w16010;
assign w16012 = pi54 & pi58;
assign w16013 = w15881 & w16012;
assign w16014 = ~w16011 & ~w16013;
assign w16015 = w16009 & ~w16014;
assign w16016 = ~w16009 & w16014;
assign w16017 = ~w16015 & ~w16016;
assign w16018 = w16008 & ~w16017;
assign w16019 = ~w16008 & w16017;
assign w16020 = ~w16018 & ~w16019;
assign w16021 = ~w15992 & w16020;
assign w16022 = w15992 & ~w16020;
assign w16023 = ~w16021 & ~w16022;
assign w16024 = w15991 & w16023;
assign w16025 = ~w15991 & ~w16023;
assign w16026 = ~w16024 & ~w16025;
assign w16027 = ~w15972 & w16026;
assign w16028 = w15972 & ~w16026;
assign w16029 = ~w16027 & ~w16028;
assign w16030 = (~w11122 & w17664) | (~w11122 & w17665) | (w17664 & w17665);
assign w16031 = (w11122 & w17666) | (w11122 & w17667) | (w17666 & w17667);
assign w16032 = ~w16030 & ~w16031;
assign w16033 = ~w16021 & ~w16024;
assign w16034 = ~w15986 & ~w15990;
assign w16035 = pi49 & pi63;
assign w16036 = pi52 & pi60;
assign w16037 = ~w15995 & ~w16036;
assign w16038 = pi52 & pi61;
assign w16039 = w15915 & w16038;
assign w16040 = ~w16037 & ~w16039;
assign w16041 = w16035 & ~w16040;
assign w16042 = ~w16035 & w16040;
assign w16043 = ~w16041 & ~w16042;
assign w16044 = w15934 & ~w15994;
assign w16045 = ~w15996 & ~w16044;
assign w16046 = ~w16043 & ~w16045;
assign w16047 = w16043 & w16045;
assign w16048 = ~w16046 & ~w16047;
assign w16049 = pi53 & pi59;
assign w16050 = pi55 & pi57;
assign w16051 = ~w16012 & ~w16050;
assign w16052 = pi55 & pi58;
assign w16053 = w15945 & w16052;
assign w16054 = ~w16051 & ~w16053;
assign w16055 = w16049 & ~w16054;
assign w16056 = ~w16049 & w16054;
assign w16057 = ~w16055 & ~w16056;
assign w16058 = w16048 & ~w16057;
assign w16059 = ~w16048 & w16057;
assign w16060 = ~w16058 & ~w16059;
assign w16061 = ~w16034 & w16060;
assign w16062 = w16034 & ~w16060;
assign w16063 = ~w16061 & ~w16062;
assign w16064 = pi50 & pi62;
assign w16065 = ~pi55 & ~w16001;
assign w16066 = pi56 & ~w16065;
assign w16067 = w16064 & w16066;
assign w16068 = ~w16064 & ~w16066;
assign w16069 = ~w16067 & ~w16068;
assign w16070 = w16009 & ~w16011;
assign w16071 = ~w16013 & ~w16070;
assign w16072 = w16069 & ~w16071;
assign w16073 = ~w16069 & w16071;
assign w16074 = ~w16072 & ~w16073;
assign w16075 = ~w15978 & ~w15982;
assign w16076 = ~w16006 & ~w16018;
assign w16077 = ~w16075 & ~w16076;
assign w16078 = w16075 & w16076;
assign w16079 = ~w16077 & ~w16078;
assign w16080 = w16074 & w16079;
assign w16081 = ~w16074 & ~w16079;
assign w16082 = ~w16080 & ~w16081;
assign w16083 = w16063 & w16082;
assign w16084 = ~w16063 & ~w16082;
assign w16085 = ~w16083 & ~w16084;
assign w16086 = ~w16033 & w16085;
assign w16087 = w16033 & ~w16085;
assign w16088 = ~w16028 & ~w16087;
assign w16089 = (w11122 & w17668) | (w11122 & w17669) | (w17668 & w17669);
assign w16090 = ~w16086 & ~w16087;
assign w16091 = ~w16027 & ~w16090;
assign w16092 = (w13978 & w17401) | (w13978 & w17402) | (w17401 & w17402);
assign w16093 = ~w16089 & ~w16092;
assign w16094 = ~w16061 & ~w16083;
assign w16095 = ~w16046 & ~w16058;
assign w16096 = pi53 & pi60;
assign w16097 = ~w16038 & ~w16096;
assign w16098 = pi53 & pi61;
assign w16099 = w16036 & w16098;
assign w16100 = ~w16097 & ~w16099;
assign w16101 = w16049 & ~w16051;
assign w16102 = ~w16053 & ~w16101;
assign w16103 = w16100 & ~w16102;
assign w16104 = ~w16100 & w16102;
assign w16105 = ~w16103 & ~w16104;
assign w16106 = ~w16067 & ~w16072;
assign w16107 = w16105 & ~w16106;
assign w16108 = ~w16105 & w16106;
assign w16109 = ~w16107 & ~w16108;
assign w16110 = w16095 & ~w16109;
assign w16111 = ~w16095 & w16109;
assign w16112 = ~w16110 & ~w16111;
assign w16113 = ~w16077 & ~w16080;
assign w16114 = pi50 & pi63;
assign w16115 = pi54 & pi59;
assign w16116 = ~w16052 & ~w16115;
assign w16117 = pi55 & pi59;
assign w16118 = w16012 & w16117;
assign w16119 = ~w16116 & ~w16118;
assign w16120 = w16114 & ~w16119;
assign w16121 = ~w16114 & w16119;
assign w16122 = ~w16120 & ~w16121;
assign w16123 = w16035 & ~w16037;
assign w16124 = ~w16039 & ~w16123;
assign w16125 = ~w16122 & ~w16124;
assign w16126 = w16122 & w16124;
assign w16127 = ~w16125 & ~w16126;
assign w16128 = pi51 & pi62;
assign w16129 = ~pi56 & pi57;
assign w16130 = w16128 & ~w16129;
assign w16131 = ~w16128 & w16129;
assign w16132 = ~w16130 & ~w16131;
assign w16133 = w16127 & ~w16132;
assign w16134 = ~w16127 & w16132;
assign w16135 = ~w16133 & ~w16134;
assign w16136 = ~w16113 & w16135;
assign w16137 = w16113 & ~w16135;
assign w16138 = ~w16136 & ~w16137;
assign w16139 = ~w16112 & ~w16138;
assign w16140 = w16112 & w16138;
assign w16141 = ~w16139 & ~w16140;
assign w16142 = w16094 & ~w16141;
assign w16143 = ~w16094 & w16141;
assign w16144 = ~w16142 & ~w16143;
assign w16145 = (w13978 & w17403) | (w13978 & w17404) | (w17403 & w17404);
assign w16146 = (~w13978 & w17405) | (~w13978 & w17406) | (w17405 & w17406);
assign w16147 = ~w16145 & ~w16146;
assign w16148 = ~w16086 & ~w16143;
assign w16149 = ~w16136 & ~w16140;
assign w16150 = ~w16099 & ~w16103;
assign w16151 = ~pi56 & ~w16128;
assign w16152 = pi57 & ~w16151;
assign w16153 = w16114 & ~w16116;
assign w16154 = ~w16118 & ~w16153;
assign w16155 = w16152 & ~w16154;
assign w16156 = ~w16152 & w16154;
assign w16157 = ~w16155 & ~w16156;
assign w16158 = w16150 & ~w16157;
assign w16159 = ~w16150 & w16157;
assign w16160 = ~w16158 & ~w16159;
assign w16161 = ~w16107 & ~w16111;
assign w16162 = ~w16160 & w16161;
assign w16163 = w16160 & ~w16161;
assign w16164 = ~w16162 & ~w16163;
assign w16165 = ~w16125 & ~w16133;
assign w16166 = pi54 & pi60;
assign w16167 = pi56 & pi58;
assign w16168 = ~w16117 & ~w16167;
assign w16169 = pi56 & pi59;
assign w16170 = w16052 & w16169;
assign w16171 = ~w16168 & ~w16170;
assign w16172 = w16166 & ~w16171;
assign w16173 = ~w16166 & w16171;
assign w16174 = ~w16172 & ~w16173;
assign w16175 = pi51 & pi63;
assign w16176 = pi52 & pi62;
assign w16177 = ~w16098 & ~w16176;
assign w16178 = pi53 & pi62;
assign w16179 = w16038 & w16178;
assign w16180 = ~w16177 & ~w16179;
assign w16181 = w16175 & ~w16180;
assign w16182 = ~w16175 & w16180;
assign w16183 = ~w16181 & ~w16182;
assign w16184 = ~w16174 & ~w16183;
assign w16185 = w16174 & w16183;
assign w16186 = ~w16184 & ~w16185;
assign w16187 = w16165 & ~w16186;
assign w16188 = ~w16165 & w16186;
assign w16189 = ~w16187 & ~w16188;
assign w16190 = w16164 & w16189;
assign w16191 = ~w16164 & ~w16189;
assign w16192 = ~w16190 & ~w16191;
assign w16193 = w16149 & ~w16192;
assign w16194 = ~w16149 & w16192;
assign w16195 = ~w16193 & ~w16194;
assign w16196 = (~w12329 & w17531) | (~w12329 & w17532) | (w17531 & w17532);
assign w16197 = (w12329 & w17533) | (w12329 & w17534) | (w17533 & w17534);
assign w16198 = ~w16196 & ~w16197;
assign w16199 = ~w16163 & ~w16190;
assign w16200 = ~w16155 & ~w16159;
assign w16201 = pi54 & pi61;
assign w16202 = pi55 & pi60;
assign w16203 = ~w16169 & ~w16202;
assign w16204 = pi56 & pi60;
assign w16205 = w16117 & w16204;
assign w16206 = ~w16203 & ~w16205;
assign w16207 = w16201 & ~w16206;
assign w16208 = ~w16201 & w16206;
assign w16209 = ~w16207 & ~w16208;
assign w16210 = ~pi57 & pi58;
assign w16211 = w16178 & ~w16210;
assign w16212 = ~w16178 & w16210;
assign w16213 = ~w16211 & ~w16212;
assign w16214 = ~w16209 & ~w16213;
assign w16215 = w16209 & w16213;
assign w16216 = ~w16214 & ~w16215;
assign w16217 = w16200 & ~w16216;
assign w16218 = ~w16200 & w16216;
assign w16219 = ~w16217 & ~w16218;
assign w16220 = pi52 & pi63;
assign w16221 = w16166 & ~w16168;
assign w16222 = ~w16170 & ~w16221;
assign w16223 = w16220 & ~w16222;
assign w16224 = ~w16220 & w16222;
assign w16225 = ~w16223 & ~w16224;
assign w16226 = w16175 & ~w16177;
assign w16227 = ~w16179 & ~w16226;
assign w16228 = ~w16225 & w16227;
assign w16229 = w16225 & ~w16227;
assign w16230 = ~w16228 & ~w16229;
assign w16231 = ~w16184 & ~w16188;
assign w16232 = ~w16230 & w16231;
assign w16233 = w16230 & ~w16231;
assign w16234 = ~w16232 & ~w16233;
assign w16235 = w16219 & w16234;
assign w16236 = ~w16219 & ~w16234;
assign w16237 = ~w16235 & ~w16236;
assign w16238 = ~w16199 & w16237;
assign w16239 = w16199 & ~w16237;
assign w16240 = ~w16238 & ~w16239;
assign w16241 = (~w13978 & w17407) | (~w13978 & w17408) | (w17407 & w17408);
assign w16242 = (w13978 & w17409) | (w13978 & w17410) | (w17409 & w17410);
assign w16243 = ~w16241 & ~w16242;
assign w16244 = ~w16193 & ~w16239;
assign w16245 = pi54 & pi62;
assign w16246 = pi53 & pi63;
assign w16247 = ~w16245 & ~w16246;
assign w16248 = pi54 & pi63;
assign w16249 = w16178 & w16248;
assign w16250 = ~w16247 & ~w16249;
assign w16251 = ~pi57 & ~w16178;
assign w16252 = pi58 & ~w16251;
assign w16253 = w16250 & w16252;
assign w16254 = ~w16250 & ~w16252;
assign w16255 = ~w16253 & ~w16254;
assign w16256 = pi55 & pi61;
assign w16257 = pi57 & pi59;
assign w16258 = ~w16204 & ~w16257;
assign w16259 = pi57 & pi60;
assign w16260 = w16169 & w16259;
assign w16261 = ~w16258 & ~w16260;
assign w16262 = w16256 & ~w16261;
assign w16263 = ~w16256 & w16261;
assign w16264 = ~w16262 & ~w16263;
assign w16265 = w16201 & ~w16203;
assign w16266 = ~w16205 & ~w16265;
assign w16267 = ~w16264 & ~w16266;
assign w16268 = w16264 & w16266;
assign w16269 = ~w16267 & ~w16268;
assign w16270 = w16255 & w16269;
assign w16271 = ~w16255 & ~w16269;
assign w16272 = ~w16270 & ~w16271;
assign w16273 = ~w16214 & ~w16218;
assign w16274 = ~w16223 & ~w16229;
assign w16275 = ~w16273 & ~w16274;
assign w16276 = w16273 & w16274;
assign w16277 = ~w16275 & ~w16276;
assign w16278 = w16272 & w16277;
assign w16279 = ~w16272 & ~w16277;
assign w16280 = ~w16278 & ~w16279;
assign w16281 = ~w16233 & ~w16235;
assign w16282 = w16280 & ~w16281;
assign w16283 = ~w16280 & w16281;
assign w16284 = ~w16282 & ~w16283;
assign w16285 = (w13978 & w17411) | (w13978 & w17412) | (w17411 & w17412);
assign w16286 = (~w13978 & w17413) | (~w13978 & w17414) | (w17413 & w17414);
assign w16287 = ~w16285 & ~w16286;
assign w16288 = ~w16238 & ~w16282;
assign w16289 = ~w16275 & ~w16278;
assign w16290 = ~w16249 & ~w16253;
assign w16291 = w16256 & ~w16258;
assign w16292 = ~w16260 & ~w16291;
assign w16293 = ~w16290 & ~w16292;
assign w16294 = w16290 & w16292;
assign w16295 = ~w16293 & ~w16294;
assign w16296 = pi56 & pi61;
assign w16297 = ~w16259 & ~w16296;
assign w16298 = pi57 & pi61;
assign w16299 = w16204 & w16298;
assign w16300 = ~w16297 & ~w16299;
assign w16301 = w16248 & ~w16300;
assign w16302 = ~w16248 & w16300;
assign w16303 = ~w16301 & ~w16302;
assign w16304 = ~w16295 & w16303;
assign w16305 = w16295 & ~w16303;
assign w16306 = ~w16304 & ~w16305;
assign w16307 = ~w16267 & ~w16270;
assign w16308 = pi55 & pi62;
assign w16309 = ~pi58 & pi59;
assign w16310 = w16308 & ~w16309;
assign w16311 = ~w16308 & w16309;
assign w16312 = ~w16310 & ~w16311;
assign w16313 = ~w16307 & ~w16312;
assign w16314 = w16307 & w16312;
assign w16315 = ~w16313 & ~w16314;
assign w16316 = w16306 & w16315;
assign w16317 = ~w16306 & ~w16315;
assign w16318 = ~w16316 & ~w16317;
assign w16319 = w16289 & ~w16318;
assign w16320 = ~w16289 & w16318;
assign w16321 = ~w16319 & ~w16320;
assign w16322 = (w11122 & w17670) | (w11122 & w17671) | (w17670 & w17671);
assign w16323 = (~w11122 & w17672) | (~w11122 & w17673) | (w17672 & w17673);
assign w16324 = ~w16322 & ~w16323;
assign w16325 = pi55 & pi63;
assign w16326 = ~pi58 & ~w16308;
assign w16327 = pi59 & ~w16326;
assign w16328 = w16325 & w16327;
assign w16329 = ~w16325 & ~w16327;
assign w16330 = ~w16328 & ~w16329;
assign w16331 = w16248 & ~w16297;
assign w16332 = ~w16299 & ~w16331;
assign w16333 = ~w16330 & w16332;
assign w16334 = w16330 & ~w16332;
assign w16335 = ~w16333 & ~w16334;
assign w16336 = ~w16293 & ~w16305;
assign w16337 = pi56 & pi62;
assign w16338 = pi58 & pi60;
assign w16339 = ~w16298 & ~w16338;
assign w16340 = pi58 & pi61;
assign w16341 = w16259 & w16340;
assign w16342 = ~w16339 & ~w16341;
assign w16343 = w16337 & ~w16342;
assign w16344 = ~w16337 & w16342;
assign w16345 = ~w16343 & ~w16344;
assign w16346 = ~w16336 & ~w16345;
assign w16347 = w16336 & w16345;
assign w16348 = ~w16346 & ~w16347;
assign w16349 = ~w16335 & ~w16348;
assign w16350 = w16335 & w16348;
assign w16351 = ~w16349 & ~w16350;
assign w16352 = ~w16313 & ~w16316;
assign w16353 = ~w16351 & w16352;
assign w16354 = w16351 & ~w16352;
assign w16355 = ~w16353 & ~w16354;
assign w16356 = (w15213 & w17325) | (w15213 & w17326) | (w17325 & w17326);
assign w16357 = (~w15213 & w17327) | (~w15213 & w17328) | (w17327 & w17328);
assign w16358 = ~w16356 & ~w16357;
assign w16359 = ~w16328 & ~w16334;
assign w16360 = pi56 & pi63;
assign w16361 = ~w16340 & ~w16360;
assign w16362 = w16340 & w16360;
assign w16363 = ~w16361 & ~w16362;
assign w16364 = w16337 & ~w16339;
assign w16365 = ~w16341 & ~w16364;
assign w16366 = w16363 & ~w16365;
assign w16367 = ~w16363 & w16365;
assign w16368 = ~w16366 & ~w16367;
assign w16369 = pi57 & pi62;
assign w16370 = ~pi59 & pi60;
assign w16371 = w16369 & ~w16370;
assign w16372 = ~w16369 & w16370;
assign w16373 = ~w16371 & ~w16372;
assign w16374 = w16368 & ~w16373;
assign w16375 = ~w16368 & w16373;
assign w16376 = ~w16374 & ~w16375;
assign w16377 = w16359 & ~w16376;
assign w16378 = ~w16359 & w16376;
assign w16379 = ~w16377 & ~w16378;
assign w16380 = ~w16346 & ~w16350;
assign w16381 = w16379 & ~w16380;
assign w16382 = ~w16379 & w16380;
assign w16383 = ~w16381 & ~w16382;
assign w16384 = ~w16319 & ~w16353;
assign w16385 = (~w15213 & w17329) | (~w15213 & w17330) | (w17329 & w17330);
assign w16386 = (w15213 & w17331) | (w15213 & w17332) | (w17331 & w17332);
assign w16387 = ~w16385 & ~w16386;
assign w16388 = ~w16354 & ~w16381;
assign w16389 = ~w16374 & ~w16378;
assign w16390 = ~w16362 & ~w16366;
assign w16391 = ~pi59 & ~w16369;
assign w16392 = pi60 & ~w16391;
assign w16393 = ~w16390 & w16392;
assign w16394 = w16390 & ~w16392;
assign w16395 = ~w16393 & ~w16394;
assign w16396 = pi57 & pi63;
assign w16397 = pi59 & pi61;
assign w16398 = pi58 & pi62;
assign w16399 = ~w16397 & ~w16398;
assign w16400 = pi59 & pi62;
assign w16401 = w16340 & w16400;
assign w16402 = ~w16399 & ~w16401;
assign w16403 = w16396 & ~w16402;
assign w16404 = ~w16396 & w16402;
assign w16405 = ~w16403 & ~w16404;
assign w16406 = w16395 & ~w16405;
assign w16407 = ~w16395 & w16405;
assign w16408 = ~w16406 & ~w16407;
assign w16409 = ~w16389 & w16408;
assign w16410 = w16389 & ~w16408;
assign w16411 = ~w16409 & ~w16410;
assign w16412 = (~w13978 & w17416) | (~w13978 & w17417) | (w17416 & w17417);
assign w16413 = (w13978 & w17418) | (w13978 & w17419) | (w17418 & w17419);
assign w16414 = ~w16412 & ~w16413;
assign w16415 = pi58 & pi63;
assign w16416 = w16396 & ~w16399;
assign w16417 = ~w16401 & ~w16416;
assign w16418 = ~w16415 & w16417;
assign w16419 = w16415 & ~w16417;
assign w16420 = ~w16418 & ~w16419;
assign w16421 = ~pi60 & pi61;
assign w16422 = w16400 & ~w16421;
assign w16423 = ~w16400 & w16421;
assign w16424 = ~w16422 & ~w16423;
assign w16425 = ~w16420 & w16424;
assign w16426 = w16420 & ~w16424;
assign w16427 = ~w16425 & ~w16426;
assign w16428 = ~w16393 & ~w16406;
assign w16429 = ~w16427 & w16428;
assign w16430 = w16427 & ~w16428;
assign w16431 = ~w16429 & ~w16430;
assign w16432 = (w15213 & w17333) | (w15213 & w17334) | (w17333 & w17334);
assign w16433 = (~w15213 & w17335) | (~w15213 & w17336) | (w17335 & w17336);
assign w16434 = ~w16432 & ~w16433;
assign w16435 = ~w16410 & ~w16429;
assign w16436 = ~w16419 & ~w16426;
assign w16437 = pi59 & pi63;
assign w16438 = pi60 & pi62;
assign w16439 = ~w16437 & ~w16438;
assign w16440 = pi60 & pi63;
assign w16441 = w16400 & w16440;
assign w16442 = ~w16439 & ~w16441;
assign w16443 = ~pi60 & ~w16400;
assign w16444 = pi61 & ~w16443;
assign w16445 = w16442 & w16444;
assign w16446 = ~w16442 & ~w16444;
assign w16447 = ~w16445 & ~w16446;
assign w16448 = w16436 & ~w16447;
assign w16449 = ~w16436 & w16447;
assign w16450 = ~w16448 & ~w16449;
assign w16451 = (w10008 & w17869) | (w10008 & w17870) | (w17869 & w17870);
assign w16452 = (~w10008 & w17871) | (~w10008 & w17872) | (w17871 & w17872);
assign w16453 = ~w16451 & ~w16452;
assign w16454 = ~w16430 & ~w16449;
assign w16455 = ~w16441 & ~w16445;
assign w16456 = ~pi61 & pi62;
assign w16457 = ~w16440 & w16456;
assign w16458 = w16440 & ~w16456;
assign w16459 = ~w16457 & ~w16458;
assign w16460 = w16455 & w16459;
assign w16461 = ~w16455 & ~w16459;
assign w16462 = ~w16460 & ~w16461;
assign w16463 = (~w10008 & w17873) | (~w10008 & w17874) | (w17873 & w17874);
assign w16464 = (w10008 & w17875) | (w10008 & w17876) | (w17875 & w17876);
assign w16465 = ~w16463 & ~w16464;
assign w16466 = pi61 & pi63;
assign w16467 = pi62 & w16466;
assign w16468 = pi62 & w16459;
assign w16469 = ~w16466 & ~w16468;
assign w16470 = ~w16467 & ~w16469;
assign w16471 = (~w10008 & w17877) | (~w10008 & w17878) | (w17877 & w17878);
assign w16472 = (w10008 & w17879) | (w10008 & w17880) | (w17879 & w17880);
assign w16473 = ~w16471 & ~w16472;
assign w16474 = ~w16460 & ~w16469;
assign w16475 = ~pi62 & pi63;
assign w16476 = (~w10008 & w17881) | (~w10008 & w17882) | (w17881 & w17882);
assign w16477 = pi63 & ~w16456;
assign w16478 = (w10008 & w17883) | (w10008 & w17884) | (w17883 & w17884);
assign w16479 = ~w16476 & ~w16478;
assign w16480 = (w10008 & w17885) | (w10008 & w17886) | (w17885 & w17886);
assign w16481 = pi63 & ~w16480;
assign w16482 = ~w26 & ~w23;
assign w16483 = ~w2 & ~w6;
assign w16484 = w26 & w23;
assign w16485 = w36 & ~w50;
assign w16486 = w110 & ~w107;
assign w16487 = ~w119 & ~w121;
assign w16488 = ~w162 & ~w158;
assign w16489 = ~w235 & ~w226;
assign w16490 = w206 & ~w196;
assign w16491 = ~w257 & ~w271;
assign w16492 = ~w392 & ~w387;
assign w16493 = ~w511 & w16682;
assign w16494 = w518 & ~w510;
assign w16495 = ~w589 & ~w581;
assign w16496 = ~w740 & w902;
assign w16497 = (w816 & ~w898) | (w816 & w16803) | (~w898 & w16803);
assign w16498 = ~w1093 & ~w1084;
assign w16499 = ~w1283 & w17337;
assign w16500 = w1505 & ~w1393;
assign w16501 = w1505 & ~w16499;
assign w16502 = w1391 & ~w1502;
assign w16503 = ~w1863 & ~w1737;
assign w16504 = w1860 & w1993;
assign w16505 = w2259 & ~w1993;
assign w16506 = w2259 & ~w16504;
assign w16507 = w2122 & ~w2257;
assign w16508 = w2402 & w2257;
assign w16509 = w2402 & ~w16507;
assign w16510 = (~w2543 & w16508) | (~w2543 & w16683) | (w16508 & w16683);
assign w16511 = (~w2543 & w16509) | (~w2543 & w16683) | (w16509 & w16683);
assign w16512 = w2688 & w2997;
assign w16513 = w3160 & ~w16512;
assign w16514 = ~w2995 & ~w16513;
assign w16515 = (~w2995 & ~w3160) | (~w2995 & w16684) | (~w3160 & w16684);
assign w16516 = ~w3321 & w16804;
assign w16517 = ~w3500 & ~w3491;
assign w16518 = ~w3665 & w3491;
assign w16519 = (~w3665 & w3500) | (~w3665 & w16518) | (w3500 & w16518);
assign w16520 = ~w4023 & w4029;
assign w16521 = ~w4021 & ~w4029;
assign w16522 = ~w4021 & ~w16520;
assign w16523 = ~w4209 & ~w16521;
assign w16524 = (~w4209 & w16520) | (~w4209 & w16685) | (w16520 & w16685);
assign w16525 = ~w4594 & w4600;
assign w16526 = ~w4592 & ~w4600;
assign w16527 = ~w4592 & ~w16525;
assign w16528 = w4793 & w5002;
assign w16529 = w5206 & ~w5002;
assign w16530 = ~w5201 & ~w16529;
assign w16531 = (~w5201 & w16528) | (~w5201 & w16686) | (w16528 & w16686);
assign w16532 = w5413 & w5627;
assign w16533 = w6070 & ~w5627;
assign w16534 = ~w5847 & ~w16533;
assign w16535 = (~w5847 & w16532) | (~w5847 & w16687) | (w16532 & w16687);
assign w16536 = ~w6067 & ~w16534;
assign w16537 = ~w6067 & ~w16535;
assign w16538 = ~w6525 & w16688;
assign w16539 = ~w6526 & ~w6769;
assign w16540 = ~w6526 & ~w16538;
assign w16541 = ~w6766 & ~w16539;
assign w16542 = ~w6766 & ~w16540;
assign w16543 = ~w7251 & w7499;
assign w16544 = ~w7248 & ~w7499;
assign w16545 = ~w7248 & ~w16543;
assign w16546 = ~w7497 & ~w16544;
assign w16547 = (~w7497 & w16543) | (~w7497 & w16689) | (w16543 & w16689);
assign w16548 = w7753 & ~w16546;
assign w16549 = w7753 & ~w16547;
assign w16550 = ~w8012 & ~w8007;
assign w16551 = ~w8270 & w8007;
assign w16552 = (~w8270 & w8012) | (~w8270 & w16551) | (w8012 & w16551);
assign w16553 = ~w8526 & w16690;
assign w16554 = w8527 & ~w16552;
assign w16555 = w8794 & ~w16553;
assign w16556 = ~w8789 & ~w16555;
assign w16557 = (~w8789 & w16554) | (~w8789 & w16691) | (w16554 & w16691);
assign w16558 = w9041 & w9535;
assign w16559 = w9773 & ~w9535;
assign w16560 = ~w9532 & ~w16559;
assign w16561 = (~w9532 & w16558) | (~w9532 & w16692) | (w16558 & w16692);
assign w16562 = (~w9770 & w16559) | (~w9770 & w17535) | (w16559 & w17535);
assign w16563 = ~w9770 & ~w16561;
assign w16564 = ~w10243 & ~w10249;
assign w16565 = (~w10243 & w10013) | (~w10243 & w16564) | (w10013 & w16564);
assign w16566 = ~w10472 & ~w16564;
assign w16567 = ~w10472 & ~w16565;
assign w16568 = w10911 & ~w16566;
assign w16569 = w10911 & ~w16567;
assign w16570 = (w11121 & w16567) | (w11121 & w17420) | (w16567 & w17420);
assign w16571 = (~w10908 & w16568) | (~w10908 & w17536) | (w16568 & w17536);
assign w16572 = ~w10908 & ~w16570;
assign w16573 = w11118 & w11541;
assign w16574 = w11546 & ~w11541;
assign w16575 = ~w11539 & ~w16574;
assign w16576 = (~w11539 & w16573) | (~w11539 & w16693) | (w16573 & w16693);
assign w16577 = ~w11741 & ~w16575;
assign w16578 = ~w11741 & ~w16576;
assign w16579 = w11947 & ~w16577;
assign w16580 = w11947 & ~w16578;
assign w16581 = w12140 & ~w16580;
assign w16582 = (~w12135 & w16579) | (~w12135 & w17338) | (w16579 & w17338);
assign w16583 = ~w12135 & ~w16581;
assign w16584 = ~w12324 & ~w16582;
assign w16585 = (~w16580 & w17421) | (~w16580 & w17422) | (w17421 & w17422);
assign w16586 = ~w12688 & w12693;
assign w16587 = ~w12686 & ~w12693;
assign w16588 = ~w12686 & ~w16586;
assign w16589 = ~w12865 & ~w16587;
assign w16590 = (~w12865 & w16586) | (~w12865 & w16694) | (w16586 & w16694);
assign w16591 = w13041 & ~w16589;
assign w16592 = w13041 & ~w16590;
assign w16593 = w13208 & ~w16592;
assign w16594 = (~w13203 & w16591) | (~w13203 & w17273) | (w16591 & w17273);
assign w16595 = ~w13203 & ~w16593;
assign w16596 = ~w13364 & ~w16594;
assign w16597 = (~w16592 & w17340) | (~w16592 & w17341) | (w17340 & w17341);
assign w16598 = (w13681 & w16594) | (w13681 & w17342) | (w16594 & w17342);
assign w16599 = w13681 & ~w16597;
assign w16600 = (w16594 & w17537) | (w16594 & w17538) | (w17537 & w17538);
assign w16601 = (~w16597 & w17674) | (~w16597 & w17537) | (w17674 & w17537);
assign w16602 = ~w13831 & ~w16600;
assign w16603 = (w16597 & w17675) | (w16597 & w17676) | (w17675 & w17676);
assign w16604 = ~w13982 & w14125;
assign w16605 = ~w14120 & ~w14125;
assign w16606 = ~w14120 & ~w16604;
assign w16607 = (~w14256 & w14125) | (~w14256 & w16695) | (w14125 & w16695);
assign w16608 = (~w14256 & w16604) | (~w14256 & w16695) | (w16604 & w16695);
assign w16609 = w14520 & ~w16607;
assign w16610 = (~w16604 & w17019) | (~w16604 & w17020) | (w17019 & w17020);
assign w16611 = w14524 & ~w16610;
assign w16612 = (~w14518 & w16609) | (~w14518 & w17275) | (w16609 & w17275);
assign w16613 = ~w14518 & ~w16611;
assign w16614 = ~w14645 & ~w16612;
assign w16615 = (~w16610 & w17343) | (~w16610 & w17344) | (w17343 & w17344);
assign w16616 = (w14885 & w16612) | (w14885 & w17345) | (w16612 & w17345);
assign w16617 = w14885 & ~w16615;
assign w16618 = (~w16612 & w17425) | (~w16612 & w17426) | (w17425 & w17426);
assign w16619 = ~w14882 & ~w16618;
assign w16620 = (~w16615 & w17540) | (~w16615 & w17541) | (w17540 & w17541);
assign w16621 = ~w14993 & ~w16619;
assign w16622 = ~w14993 & ~w16620;
assign w16623 = (~w16618 & w17677) | (~w16618 & w17678) | (w17677 & w17678);
assign w16624 = (w15109 & w16620) | (w15109 & w17542) | (w16620 & w17542);
assign w16625 = w15212 & ~w16623;
assign w16626 = w15212 & ~w16624;
assign w16627 = ~w15207 & ~w16625;
assign w16628 = ~w15207 & ~w16626;
assign w16629 = w15311 & w15411;
assign w16630 = w15588 & ~w15411;
assign w16631 = ~w15499 & ~w16630;
assign w16632 = (~w15499 & w16629) | (~w15499 & w16696) | (w16629 & w16696);
assign w16633 = (~w15586 & w16630) | (~w15586 & w16805) | (w16630 & w16805);
assign w16634 = ~w15586 & ~w16632;
assign w16635 = (~w16630 & w16806) | (~w16630 & w17021) | (w16806 & w17021);
assign w16636 = (w15676 & w16632) | (w15676 & w16806) | (w16632 & w16806);
assign w16637 = (~w16632 & w17022) | (~w16632 & w17023) | (w17022 & w17023);
assign w16638 = (~w15749 & w16635) | (~w15749 & w17277) | (w16635 & w17277);
assign w16639 = ~w15749 & ~w16637;
assign w16640 = (~w16635 & w17278) | (~w16635 & w17346) | (w17278 & w17346);
assign w16641 = (~w15827 & w16637) | (~w15827 & w17278) | (w16637 & w17278);
assign w16642 = w15902 & ~w16640;
assign w16643 = (~w16637 & w17347) | (~w16637 & w17348) | (w17347 & w17348);
assign w16644 = (w16637 & w17428) | (w16637 & w17429) | (w17428 & w17429);
assign w16645 = (~w16640 & w17543) | (~w16640 & w17544) | (w17543 & w17544);
assign w16646 = ~w15966 & ~w16644;
assign w16647 = (w16640 & w17679) | (w16640 & w17680) | (w17679 & w17680);
assign w16648 = (w16637 & w17681) | (w16637 & w17682) | (w17681 & w17682);
assign w16649 = w16088 & ~w16647;
assign w16650 = w16088 & ~w16648;
assign w16651 = w16148 & ~w16649;
assign w16652 = w16148 & ~w16650;
assign w16653 = ~w16142 & ~w16651;
assign w16654 = ~w16142 & ~w16652;
assign w16655 = ~w16194 & ~w16653;
assign w16656 = ~w16194 & ~w16654;
assign w16657 = w16244 & ~w16655;
assign w16658 = w16244 & ~w16656;
assign w16659 = w16288 & ~w16657;
assign w16660 = w16288 & ~w16658;
assign w16661 = ~w16283 & ~w16659;
assign w16662 = ~w16283 & ~w16660;
assign w16663 = w16320 & w16384;
assign w16664 = w16388 & ~w16384;
assign w16665 = w16388 & ~w16663;
assign w16666 = ~w16382 & ~w16664;
assign w16667 = ~w16382 & ~w16665;
assign w16668 = ~w16409 & ~w16666;
assign w16669 = ~w16409 & ~w16667;
assign w16670 = w16435 & ~w16668;
assign w16671 = w16435 & ~w16669;
assign w16672 = w16454 & ~w16670;
assign w16673 = w16454 & ~w16671;
assign w16674 = ~w16448 & ~w16672;
assign w16675 = ~w16448 & ~w16673;
assign w16676 = ~w16461 & ~w16674;
assign w16677 = ~w16461 & ~w16675;
assign w16678 = ~w16460 & ~w16676;
assign w16679 = ~w16460 & ~w16677;
assign w16680 = w16474 & ~w16676;
assign w16681 = w16474 & ~w16677;
assign w16682 = ~w449 & w448;
assign w16683 = ~w2690 & ~w2543;
assign w16684 = w2997 & ~w2995;
assign w16685 = w4021 & ~w4209;
assign w16686 = ~w5206 & ~w5201;
assign w16687 = ~w6070 & ~w5847;
assign w16688 = ~w6295 & ~w6528;
assign w16689 = w7248 & ~w7497;
assign w16690 = ~w8269 & ~w16551;
assign w16691 = ~w8794 & ~w8789;
assign w16692 = ~w9773 & ~w9532;
assign w16693 = ~w11546 & ~w11539;
assign w16694 = w12686 & ~w12865;
assign w16695 = w14120 & ~w14256;
assign w16696 = ~w15588 & ~w15499;
assign w16697 = w327 & ~w316;
assign w16698 = ~w376 & ~w372;
assign w16699 = w395 & ~w416;
assign w16700 = w437 & ~w426;
assign w16701 = w470 & ~w459;
assign w16702 = w570 & ~w559;
assign w16703 = ~w656 & w581;
assign w16704 = ~w656 & ~w16495;
assign w16705 = w645 & ~w631;
assign w16706 = ~w802 & ~w798;
assign w16707 = ~w972 & ~w968;
assign w16708 = w998 & ~w1017;
assign w16709 = w1045 & ~w1034;
assign w16710 = ~w1131 & ~w1123;
assign w16711 = w1192 & ~w1197;
assign w16712 = ~w1306 & ~w1302;
assign w16713 = w1334 & ~w1323;
assign w16714 = ~w1404 & ~w1406;
assign w16715 = ~w1444 & ~w1440;
assign w16716 = ~w1687 & ~w1683;
assign w16717 = w2055 & ~w2044;
assign w16718 = ~w2135 & ~w2131;
assign w16719 = w2190 & ~w2179;
assign w16720 = ~w2436 & ~w2432;
assign w16721 = ~w2451 & ~w2447;
assign w16722 = ~w3011 & ~w3013;
assign w16723 = w3166 & ~w3171;
assign w16724 = ~w3295 & ~w3291;
assign w16725 = ~w3309 & ~w3307;
assign w16726 = ~w3233 & ~w3236;
assign w16727 = w3329 & ~w3364;
assign w16728 = w3377 & w3550;
assign w16729 = ~w3377 & ~w3550;
assign w16730 = ~w3360 & ~w3345;
assign w16731 = ~w3632 & ~w3628;
assign w16732 = w3972 & ~w3961;
assign w16733 = ~w3858 & ~w3854;
assign w16734 = ~w4413 & ~w4409;
assign w16735 = ~w4765 & ~w4758;
assign w16736 = ~w4697 & ~w4693;
assign w16737 = w4720 & ~w4709;
assign w16738 = ~w4918 & ~w4914;
assign w16739 = ~w4942 & ~w4938;
assign w16740 = ~w5397 & ~w5393;
assign w16741 = ~w5220 & ~w5214;
assign w16742 = ~w5503 & ~w5499;
assign w16743 = w5787 & ~w5783;
assign w16744 = ~w5767 & ~w5763;
assign w16745 = ~w6018 & ~w6011;
assign w16746 = ~w5875 & ~w5871;
assign w16747 = ~w5987 & ~w5983;
assign w16748 = ~w5887 & ~w5883;
assign w16749 = ~w6313 & ~w6309;
assign w16750 = w6595 & ~w6591;
assign w16751 = ~w6570 & ~w6566;
assign w16752 = w7071 & ~w7067;
assign w16753 = ~w7059 & ~w7055;
assign w16754 = w7834 & ~w7822;
assign w16755 = pi63 & pi01;
assign w16756 = w8231 & ~w8227;
assign w16757 = ~w8025 & ~w8021;
assign w16758 = ~w8305 & ~w8303;
assign w16759 = w8890 & w9084;
assign w16760 = ~w8890 & ~w9084;
assign w16761 = w9125 & ~w9114;
assign w16762 = w9080 & ~w9076;
assign w16763 = ~w9467 & ~w9463;
assign w16764 = w9434 & ~w9430;
assign w16765 = ~w9501 & ~w9500;
assign w16766 = w9592 & ~w9588;
assign w16767 = ~w9553 & ~w9549;
assign w16768 = w9877 & ~w9866;
assign w16769 = w10144 & ~w10134;
assign w16770 = w10745 & ~w10734;
assign w16771 = ~w10787 & ~w10783;
assign w16772 = w11240 & ~w11236;
assign w16773 = w11424 & ~w11420;
assign w16774 = ~w12648 & ~w12647;
assign w16775 = w12603 & ~w12599;
assign w16776 = ~w12615 & ~w12611;
assign w16777 = ~w12735 & ~w12731;
assign w16778 = ~w12833 & ~w12829;
assign w16779 = w12785 & w12919;
assign w16780 = ~w12785 & ~w12919;
assign w16781 = w14625 & w14653;
assign w16782 = ~w14625 & ~w14653;
assign w16783 = w14535 & ~w14531;
assign w16784 = w14699 & ~w14695;
assign w16785 = w14829 & ~w14825;
assign w16786 = w14930 & ~w14926;
assign w16787 = ~w16320 & ~w16662;
assign w16788 = ~w16320 & ~w16661;
assign w16789 = (w16384 & w16663) | (w16384 & w16662) | (w16663 & w16662);
assign w16790 = (w16384 & w16663) | (w16384 & w16661) | (w16663 & w16661);
assign w16791 = (w16668 & w16669) | (w16668 & ~w16662) | (w16669 & ~w16662);
assign w16792 = (w16668 & w16669) | (w16668 & ~w16661) | (w16669 & ~w16661);
assign w16793 = (w16670 & w16671) | (w16670 & w16662) | (w16671 & w16662);
assign w16794 = (w16670 & w16671) | (w16670 & w16661) | (w16671 & w16661);
assign w16795 = ~w16430 & w16450;
assign w16796 = w16430 & ~w16450;
assign w16797 = (w16674 & w16675) | (w16674 & w16662) | (w16675 & w16662);
assign w16798 = (w16674 & w16675) | (w16674 & w16661) | (w16675 & w16661);
assign w16799 = (w16678 & w16679) | (w16678 & w16662) | (w16679 & w16662);
assign w16800 = (w16678 & w16679) | (w16678 & w16661) | (w16679 & w16661);
assign w16801 = (w16680 & w16681) | (w16680 & w16662) | (w16681 & w16662);
assign w16802 = (w16680 & w16681) | (w16680 & w16661) | (w16681 & w16661);
assign w16803 = w821 & w816;
assign w16804 = ~w3158 & w3157;
assign w16805 = w15499 & ~w15586;
assign w16806 = w15586 & w15676;
assign w16807 = w294 & ~w286;
assign w16808 = w360 & ~w357;
assign w16809 = ~w490 & ~w501;
assign w16810 = (w16493 & w583) | (w16493 & ~w387) | (w583 & ~w387);
assign w16811 = (w16493 & w583) | (w16493 & w16492) | (w583 & w16492);
assign w16812 = ~w529 & ~w525;
assign w16813 = ~w532 & ~w535;
assign w16814 = ~w593 & ~w598;
assign w16815 = ~w603 & ~w606;
assign w16816 = w678 & ~w667;
assign w16817 = ~w691 & ~w683;
assign w16818 = ~w681 & ~w695;
assign w16819 = w786 & ~w775;
assign w16820 = w888 & ~w885;
assign w16821 = (w16497 & ~w899) | (w16497 & w902) | (~w899 & w902);
assign w16822 = (w16497 & ~w899) | (w16497 & w16496) | (~w899 & w16496);
assign w16823 = w953 & ~w942;
assign w16824 = w1172 & ~w1161;
assign w16825 = ~pi13 & w1215;
assign w16826 = pi13 & ~w1215;
assign w16827 = ~w1108 & ~w1111;
assign w16828 = ~w1337 & ~w1341;
assign w16829 = w1377 & ~w1366;
assign w16830 = w1458 & ~w1461;
assign w16831 = w1532 & ~w1521;
assign w16832 = ~w1550 & ~w1546;
assign w16833 = w1720 & ~w1709;
assign w16834 = (~w1642 & w1643) | (~w1642 & w17024) | (w1643 & w17024);
assign w16835 = ~w1757 & ~w1749;
assign w16836 = w1844 & ~w1833;
assign w16837 = w1746 & ~w1761;
assign w16838 = ~w2077 & ~w2073;
assign w16839 = ~w2092 & ~w2088;
assign w16840 = ~w2193 & ~w2159;
assign w16841 = w2197 & ~w2200;
assign w16842 = w2213 & ~w2234;
assign w16843 = ~w2303 & ~w2299;
assign w16844 = ~w2306 & ~w2321;
assign w16845 = w2377 & ~w2366;
assign w16846 = w2267 & ~w2278;
assign w16847 = ~w2539 & ~w2424;
assign w16848 = ~w2536 & ~w2461;
assign w16849 = w2530 & ~w2519;
assign w16850 = ~w2439 & ~w2455;
assign w16851 = ~w2533 & ~w2498;
assign w16852 = w2418 & w2677;
assign w16853 = ~w2418 & ~w2677;
assign w16854 = w2551 & ~w2554;
assign w16855 = ~w2613 & ~w2606;
assign w16856 = ~w2817 & ~w2809;
assign w16857 = ~w2860 & ~w2856;
assign w16858 = w2972 & ~w2961;
assign w16859 = w2914 & ~w2904;
assign w16860 = ~w3063 & ~w3059;
assign w16861 = ~w3033 & ~w3029;
assign w16862 = w3100 & ~w3089;
assign w16863 = w3141 & ~w3130;
assign w16864 = w3210 & ~w3199;
assign w16865 = w3272 & ~w3261;
assign w16866 = ~w3357 & ~w3353;
assign w16867 = w3592 & ~w3614;
assign w16868 = ~w3601 & ~w3594;
assign w16869 = ~w3585 & ~w3551;
assign w16870 = w3778 & ~w3789;
assign w16871 = w3748 & ~w3772;
assign w16872 = w3761 & ~w3766;
assign w16873 = w3944 & ~w3933;
assign w16874 = w3910 & ~w3899;
assign w16875 = w4032 & ~w4035;
assign w16876 = w4307 & ~w4296;
assign w16877 = ~w4379 & ~w4375;
assign w16878 = w4334 & ~w4322;
assign w16879 = w4569 & ~w4558;
assign w16880 = w4518 & ~w4507;
assign w16881 = w4673 & ~w4662;
assign w16882 = w4755 & ~w4769;
assign w16883 = w4637 & ~w4625;
assign w16884 = w4955 & ~w4947;
assign w16885 = w4832 & ~w4821;
assign w16886 = w4858 & ~w4847;
assign w16887 = w4894 & ~w4883;
assign w16888 = w4969 & ~w4972;
assign w16889 = ~w5124 & ~w5127;
assign w16890 = w5009 & ~w5027;
assign w16891 = w5421 & ~w5432;
assign w16892 = w5602 & ~w5591;
assign w16893 = w5483 & ~w5473;
assign w16894 = ~w5453 & ~w5449;
assign w16895 = w5820 & ~w5823;
assign w16896 = w5740 & ~w5729;
assign w16897 = w5668 & ~w5657;
assign w16898 = w5854 & ~w5857;
assign w16899 = w6199 & ~w6187;
assign w16900 = ~w6125 & ~w6128;
assign w16901 = w6091 & ~w6080;
assign w16902 = w6122 & ~w6119;
assign w16903 = w6364 & ~w6353;
assign w16904 = w6459 & ~w6457;
assign w16905 = w6675 & ~w6663;
assign w16906 = w6727 & ~w6740;
assign w16907 = w6911 & ~w6900;
assign w16908 = w6984 & ~w6973;
assign w16909 = w6778 & ~w6781;
assign w16910 = w7160 & ~w7149;
assign w16911 = w7261 & ~w7264;
assign w16912 = w7572 & ~w7562;
assign w16913 = w7774 & ~w7763;
assign w16914 = ~w7952 & ~w7948;
assign w16915 = w7940 & ~w7936;
assign w16916 = w8033 & ~w8031;
assign w16917 = ~w8234 & ~w8249;
assign w16918 = w8447 & ~w8450;
assign w16919 = w8376 & ~w8365;
assign w16920 = w8633 & ~w8623;
assign w16921 = w8659 & ~w8647;
assign w16922 = w9242 & ~w9231;
assign w16923 = ~w9090 & ~w9086;
assign w16924 = w9367 & ~w9357;
assign w16925 = w9402 & ~w9391;
assign w16926 = w9335 & ~w9323;
assign w16927 = w9485 & ~w9488;
assign w16928 = w9656 & ~w9646;
assign w16929 = w9685 & ~w9673;
assign w16930 = ~w9556 & ~w9559;
assign w16931 = w9858 & ~w9848;
assign w16932 = ~w9977 & ~w9980;
assign w16933 = w10188 & ~w10177;
assign w16934 = w10017 & ~w10021;
assign w16935 = w10253 & ~w10264;
assign w16936 = w10889 & ~w10878;
assign w16937 = w10856 & ~w10845;
assign w16938 = w11050 & ~w11039;
assign w16939 = w11014 & ~w11008;
assign w16940 = w10917 & ~w10920;
assign w16941 = w11317 & ~w11305;
assign w16942 = w11522 & ~w11511;
assign w16943 = w11492 & ~w11485;
assign w16944 = ~w11400 & ~w11399;
assign w16945 = w11394 & ~w11406;
assign w16946 = w11709 & ~w11714;
assign w16947 = w11667 & ~w11663;
assign w16948 = w11655 & ~w11651;
assign w16949 = ~w11789 & ~w11764;
assign w16950 = w12579 & ~w12568;
assign w16951 = w12543 & ~w12532;
assign w16952 = w12712 & ~w12700;
assign w16953 = w12809 & ~w12798;
assign w16954 = w12777 & ~w12766;
assign w16955 = ~w12738 & ~w12741;
assign w16956 = ~w12925 & ~w12921;
assign w16957 = pi42 & pi43;
assign w16958 = w12987 & ~w12976;
assign w16959 = w12873 & ~w12876;
assign w16960 = w13107 & ~w13098;
assign w16961 = ~w13052 & ~w13050;
assign w16962 = w13308 & ~w13298;
assign w16963 = w14748 & ~w14737;
assign w16964 = w14659 & ~w14655;
assign w16965 = pi48 & pi49;
assign w16966 = w14797 & ~w14785;
assign w16967 = ~w14843 & ~w14841;
assign w16968 = ~w14846 & ~w14864;
assign w16969 = ~w14869 & ~w14835;
assign w16970 = w14812 & ~w14815;
assign w16971 = w14891 & ~w14897;
assign w16972 = w15001 & ~w15012;
assign w16973 = ~w15311 & ~w16628;
assign w16974 = ~w15311 & ~w16627;
assign w16975 = (w15411 & w16629) | (w15411 & w16628) | (w16629 & w16628);
assign w16976 = (w15411 & w16629) | (w15411 & w16627) | (w16629 & w16627);
assign w16977 = (w16633 & w16634) | (w16633 & ~w16628) | (w16634 & ~w16628);
assign w16978 = (w16633 & w16634) | (w16633 & ~w16627) | (w16634 & ~w16627);
assign w16979 = (w16636 & w16635) | (w16636 & w16628) | (w16635 & w16628);
assign w16980 = (w16636 & w16635) | (w16636 & w16627) | (w16635 & w16627);
assign w16981 = (w16641 & w16640) | (w16641 & ~w16628) | (w16640 & ~w16628);
assign w16982 = (w16641 & w16640) | (w16641 & ~w16627) | (w16640 & ~w16627);
assign w16983 = (w16643 & w16642) | (w16643 & w16628) | (w16642 & w16628);
assign w16984 = (w16643 & w16642) | (w16643 & w16627) | (w16642 & w16627);
assign w16985 = (w16646 & w16645) | (w16646 & w16628) | (w16645 & w16628);
assign w16986 = (w16646 & w16645) | (w16646 & w16627) | (w16645 & w16627);
assign w16987 = (w16650 & w16649) | (w16650 & w16628) | (w16649 & w16628);
assign w16988 = (w16650 & w16649) | (w16650 & w16627) | (w16649 & w16627);
assign w16989 = (w16656 & w16655) | (w16656 & ~w16628) | (w16655 & ~w16628);
assign w16990 = (w16656 & w16655) | (w16656 & ~w16627) | (w16655 & ~w16627);
assign w16991 = (w16658 & w16657) | (w16658 & w16628) | (w16657 & w16628);
assign w16992 = (w16658 & w16657) | (w16658 & w16627) | (w16657 & w16627);
assign w16993 = (w16662 & w16661) | (w16662 & w16628) | (w16661 & w16628);
assign w16994 = (w16662 & w16661) | (w16662 & w16627) | (w16661 & w16627);
assign w16995 = ~w16319 & ~w16788;
assign w16996 = ~w16319 & ~w16787;
assign w16997 = ~w16354 & ~w16790;
assign w16998 = ~w16354 & ~w16789;
assign w16999 = ~w16410 & ~w16792;
assign w17000 = ~w16410 & ~w16791;
assign w17001 = w16795 & ~w16794;
assign w17002 = w16795 & ~w16793;
assign w17003 = (~w16450 & w16796) | (~w16450 & w16794) | (w16796 & w16794);
assign w17004 = (~w16450 & w16796) | (~w16450 & w16793) | (w16796 & w16793);
assign w17005 = ~w16462 & w16798;
assign w17006 = ~w16462 & w16797;
assign w17007 = w16462 & ~w16798;
assign w17008 = w16462 & ~w16797;
assign w17009 = ~w16470 & w16800;
assign w17010 = ~w16470 & w16799;
assign w17011 = w16470 & ~w16800;
assign w17012 = w16470 & ~w16799;
assign w17013 = ~w16475 & w16802;
assign w17014 = ~w16475 & w16801;
assign w17015 = w16477 & ~w16802;
assign w17016 = w16477 & ~w16801;
assign w17017 = ~pi62 & ~w16802;
assign w17018 = ~pi62 & ~w16801;
assign w17019 = w14520 & w14256;
assign w17020 = w14520 & ~w16695;
assign w17021 = w15676 & ~w16805;
assign w17022 = w15755 & ~w15676;
assign w17023 = w15755 & ~w16806;
assign w17024 = w1644 & ~w1642;
assign w17025 = ~w611 & ~w649;
assign w17026 = ~w700 & ~w728;
assign w17027 = ~w755 & ~w833;
assign w17028 = w755 & w833;
assign w17029 = ~w789 & ~w806;
assign w17030 = ~w881 & ~w875;
assign w17031 = ~w830 & ~w826;
assign w17032 = (~w956 & w920) | (~w956 & w17279) | (w920 & w17279);
assign w17033 = w909 & ~w914;
assign w17034 = ~w1069 & ~w1072;
assign w17035 = ~w1066 & ~w1062;
assign w17036 = w1121 & ~w1144;
assign w17037 = w1120 & ~w1176;
assign w17038 = ~w1105 & ~w1101;
assign w17039 = ~w1239 & ~w1274;
assign w17040 = w1207 & ~w1205;
assign w17041 = (~w1435 & w1448) | (~w1435 & w17280) | (w1448 & w17280);
assign w17042 = (~w1502 & w16502) | (~w1502 & w16501) | (w16502 & w16501);
assign w17043 = (~w1502 & w16502) | (~w1502 & w16500) | (w16502 & w16500);
assign w17044 = (~w1605 & w1577) | (~w1605 & w17281) | (w1577 & w17281);
assign w17045 = ~w1573 & ~w1569;
assign w17046 = w1639 & ~w1628;
assign w17047 = w1660 & ~w1671;
assign w17048 = ~w1782 & ~w1803;
assign w17049 = ~w1850 & ~w1848;
assign w17050 = w1892 & ~w1881;
assign w17051 = ~w2061 & ~w2060;
assign w17052 = w2102 & ~w2105;
assign w17053 = ~w2098 & ~w2096;
assign w17054 = ~w2101 & ~w2113;
assign w17055 = ~w2117 & ~w2065;
assign w17056 = ~w2196 & ~w2208;
assign w17057 = w2154 & ~w2143;
assign w17058 = w2340 & ~w2331;
assign w17059 = ~w2317 & ~w2313;
assign w17060 = ~w2380 & ~w2345;
assign w17061 = ~w2283 & ~w2286;
assign w17062 = w2407 & ~w2410;
assign w17063 = w2494 & ~w2483;
assign w17064 = w2667 & ~w2663;
assign w17065 = w2562 & w2797;
assign w17066 = ~w2562 & ~w2797;
assign w17067 = ~w2646 & ~w2678;
assign w17068 = ~w2655 & ~w2651;
assign w17069 = w2775 & ~w2764;
assign w17070 = w2754 & ~w2743;
assign w17071 = ~w2787 & ~w2783;
assign w17072 = ~w2757 & ~w2723;
assign w17073 = w2875 & ~w2886;
assign w17074 = w3006 & ~w3019;
assign w17075 = ~w3036 & ~w3039;
assign w17076 = ~w3298 & ~w3301;
assign w17077 = ~w3230 & ~w3226;
assign w17078 = w3405 & ~w3394;
assign w17079 = ~w3478 & ~w3444;
assign w17080 = w3417 & ~w3436;
assign w17081 = w3648 & ~w3644;
assign w17082 = ~w3654 & ~w3622;
assign w17083 = w3547 & ~w3536;
assign w17084 = w3806 & ~w3828;
assign w17085 = ~w3818 & ~w3810;
assign w17086 = ~w3987 & ~w3983;
assign w17087 = ~w3997 & ~w4008;
assign w17088 = ~w4053 & ~w4049;
assign w17089 = ~w4064 & ~w4043;
assign w17090 = ~w4056 & ~w4059;
assign w17091 = ~w4148 & ~w4144;
assign w17092 = ~w4242 & ~w4257;
assign w17093 = ~w4251 & ~w4247;
assign w17094 = ~w4365 & ~w4361;
assign w17095 = w4442 & ~w4453;
assign w17096 = w4477 & ~w4473;
assign w17097 = w4537 & ~w4526;
assign w17098 = w4421 & ~w4419;
assign w17099 = ~w4480 & ~w4483;
assign w17100 = w4739 & ~w4735;
assign w17101 = ~w4723 & ~w4703;
assign w17102 = ~w4742 & ~w4745;
assign w17103 = ~w4945 & ~w4959;
assign w17104 = ~w5132 & ~w5135;
assign w17105 = w5175 & ~w5171;
assign w17106 = ~w5121 & ~w5117;
assign w17107 = ~w5155 & ~w5151;
assign w17108 = ~w5158 & ~w5161;
assign w17109 = ~w5381 & ~w5377;
assign w17110 = w5359 & ~w5347;
assign w17111 = w5212 & ~w5233;
assign w17112 = ~w5329 & ~w5332;
assign w17113 = ~w5462 & ~w5440;
assign w17114 = ~w5515 & ~w5511;
assign w17115 = ~w5802 & ~w5798;
assign w17116 = ~w5706 & ~w5672;
assign w17117 = ~w5770 & ~w5773;
assign w17118 = ~w5974 & ~w5939;
assign w17119 = w5935 & ~w5924;
assign w17120 = w5971 & ~w5960;
assign w17121 = ~w5990 & ~w5993;
assign w17122 = ~w6153 & ~w6149;
assign w17123 = ~w6237 & ~w6203;
assign w17124 = ~w6103 & ~w6099;
assign w17125 = w6329 & ~w6325;
assign w17126 = w6486 & ~w6497;
assign w17127 = w6463 & ~w6466;
assign w17128 = ~w6451 & ~w6447;
assign w17129 = ~w6316 & ~w6333;
assign w17130 = ~w6558 & ~w6554;
assign w17131 = w6549 & ~w6574;
assign w17132 = (~w6745 & w6746) | (~w6745 & w17683) | (w6746 & w17683);
assign w17133 = ~w6736 & ~w6730;
assign w17134 = w6536 & ~w6539;
assign w17135 = (~w6914 & w6879) | (~w6914 & w17684) | (w6879 & w17684);
assign w17136 = w6868 & ~w6873;
assign w17137 = w6851 & ~w6847;
assign w17138 = w6830 & ~w6855;
assign w17139 = w6806 & ~w6821;
assign w17140 = w7041 & ~w7044;
assign w17141 = (~w7234 & w7198) | (~w7234 & w17685) | (w7198 & w17685);
assign w17142 = ~w7297 & ~w7290;
assign w17143 = ~w7437 & ~w7433;
assign w17144 = w7587 & ~w7592;
assign w17145 = (~w7575 & w7507) | (~w7575 & w17546) | (w7507 & w17546);
assign w17146 = ~w7627 & ~w7623;
assign w17147 = w7902 & ~w7890;
assign w17148 = ~w7943 & ~w7971;
assign w17149 = w7923 & ~w7926;
assign w17150 = w8210 & ~w8213;
assign w17151 = w8044 & ~w8038;
assign w17152 = w8243 & ~w8239;
assign w17153 = ~w8455 & ~w8458;
assign w17154 = w8540 & ~w8565;
assign w17155 = w8768 & ~w8766;
assign w17156 = ~w8714 & ~w8713;
assign w17157 = (~w8743 & w8744) | (~w8743 & w17547) | (w8744 & w17547);
assign w17158 = ~w8983 & ~w8979;
assign w17159 = w9009 & ~w9005;
assign w17160 = ~w8974 & ~w8989;
assign w17161 = w9017 & ~w9015;
assign w17162 = w9068 & ~w9064;
assign w17163 = w9494 & ~w9507;
assign w17164 = w9455 & ~w9451;
assign w17165 = ~w9595 & ~w9610;
assign w17166 = w9604 & ~w9600;
assign w17167 = (~w9688 & w9627) | (~w9688 & w17430) | (w9627 & w17430);
assign w17168 = w9575 & ~w9578;
assign w17169 = w9788 & ~w9784;
assign w17170 = w9806 & ~w9804;
assign w17171 = (~w9861 & w9881) | (~w9861 & w17431) | (w9881 & w17431);
assign w17172 = w9974 & ~w9970;
assign w17173 = w9810 & ~w9813;
assign w17174 = w10060 & ~w10085;
assign w17175 = ~w10081 & ~w10077;
assign w17176 = (~w10129 & w10148) | (~w10129 & w17432) | (w10148 & w17432);
assign w17177 = w10069 & ~w10065;
assign w17178 = w10047 & ~w10050;
assign w17179 = ~w10197 & ~w10196;
assign w17180 = (~w10454 & w10417) | (~w10454 & w17433) | (w10417 & w17433);
assign w17181 = ~w10413 & ~w10409;
assign w17182 = w10302 & ~w10327;
assign w17183 = w10289 & ~w10292;
assign w17184 = (~w10676 & w10641) | (~w10676 & w17434) | (w10641 & w17434);
assign w17185 = w10775 & ~w10771;
assign w17186 = ~w10807 & ~w10806;
assign w17187 = ~w10978 & ~w10981;
assign w17188 = w10943 & ~w10948;
assign w17189 = w10975 & ~w10971;
assign w17190 = ~w11243 & ~w11246;
assign w17191 = ~w11202 & ~w11198;
assign w17192 = (~w11320 & w11255) | (~w11320 & w17686) | (w11255 & w17686);
assign w17193 = w11453 & ~w11457;
assign w17194 = ~w11436 & ~w11432;
assign w17195 = ~w11697 & w11797;
assign w17196 = w11697 & ~w11797;
assign w17197 = ~w11658 & ~w11673;
assign w17198 = w11580 & ~w11568;
assign w17199 = w11634 & ~w11637;
assign w17200 = (~w11708 & w11720) | (~w11708 & w17687) | (w11720 & w17687);
assign w17201 = w11913 & ~w11916;
assign w17202 = w11866 & ~w11857;
assign w17203 = w11900 & ~w11889;
assign w17204 = ~w11758 & ~w11754;
assign w17205 = w11815 & ~w11811;
assign w17206 = w11796 & ~w11819;
assign w17207 = w12078 & ~w12076;
assign w17208 = (~w12116 & w12117) | (~w12116 & w17688) | (w12117 & w17688);
assign w17209 = ~w12836 & ~w12839;
assign w17210 = w12906 & ~w12902;
assign w17211 = w12949 & w13061;
assign w17212 = ~w12949 & ~w13061;
assign w17213 = ~w12909 & ~w12912;
assign w17214 = w12944 & ~w12933;
assign w17215 = w13168 & ~w13164;
assign w17216 = ~w13180 & ~w13176;
assign w17217 = w13044 & ~w13056;
assign w17218 = w13150 & ~w13153;
assign w17219 = ~w13348 & ~w13351;
assign w17220 = w13339 & ~w13335;
assign w17221 = w13318 & ~w13343;
assign w17222 = w13211 & ~w13214;
assign w17223 = ~w13327 & ~w13323;
assign w17224 = w13399 & ~w13395;
assign w17225 = w13372 & ~w13375;
assign w17226 = ~w13557 & ~w13553;
assign w17227 = w13982 & ~w16603;
assign w17228 = (w13982 & w16600) | (w13982 & w17689) | (w16600 & w17689);
assign w17229 = (w16607 & w16608) | (w16607 & w16603) | (w16608 & w16603);
assign w17230 = (~w16600 & w17690) | (~w16600 & w17691) | (w17690 & w17691);
assign w17231 = (w16610 & w16609) | (w16610 & ~w16603) | (w16609 & ~w16603);
assign w17232 = (w16600 & w17692) | (w16600 & w17693) | (w17692 & w17693);
assign w17233 = (w16615 & w16614) | (w16615 & w16603) | (w16614 & w16603);
assign w17234 = (~w16600 & w17694) | (~w16600 & w17695) | (w17694 & w17695);
assign w17235 = (w16617 & w16616) | (w16617 & ~w16603) | (w16616 & ~w16603);
assign w17236 = (w16600 & w17696) | (w16600 & w17697) | (w17696 & w17697);
assign w17237 = w14918 & ~w14906;
assign w17238 = ~w14980 & ~w15017;
assign w17239 = w14980 & w15017;
assign w17240 = ~w14921 & ~w14936;
assign w17241 = (w16622 & w16621) | (w16622 & w16603) | (w16621 & w16603);
assign w17242 = (~w16600 & w17698) | (~w16600 & w17699) | (w17698 & w17699);
assign w17243 = (w16624 & w16623) | (w16624 & ~w16603) | (w16623 & ~w16603);
assign w17244 = (w16600 & w17700) | (w16600 & w17701) | (w17700 & w17701);
assign w17245 = w15055 & ~w15091;
assign w17246 = (w16628 & w16627) | (w16628 & ~w16603) | (w16627 & ~w16603);
assign w17247 = (w16628 & w16627) | (w16628 & ~w16602) | (w16627 & ~w16602);
assign w17248 = ~w15152 & ~w15151;
assign w17249 = w15147 & ~w15163;
assign w17250 = ~w15168 & ~w15144;
assign w17251 = ~w15310 & ~w16974;
assign w17252 = ~w15310 & ~w16973;
assign w17253 = ~w15405 & ~w16976;
assign w17254 = ~w15405 & ~w16975;
assign w17255 = ~w15585 & ~w16978;
assign w17256 = ~w15585 & ~w16977;
assign w17257 = ~w15670 & ~w16980;
assign w17258 = ~w15670 & ~w16979;
assign w17259 = ~w15826 & ~w16982;
assign w17260 = ~w15826 & ~w16981;
assign w17261 = ~w15896 & ~w16984;
assign w17262 = ~w15896 & ~w16983;
assign w17263 = ~w16028 & w16986;
assign w17264 = ~w16028 & w16985;
assign w17265 = ~w16086 & ~w16988;
assign w17266 = ~w16086 & ~w16987;
assign w17267 = ~w16193 & ~w16990;
assign w17268 = ~w16193 & ~w16989;
assign w17269 = ~w16238 & ~w16992;
assign w17270 = ~w16238 & ~w16991;
assign w17271 = (w16666 & w16667) | (w16666 & w16994) | (w16667 & w16994);
assign w17272 = (w16666 & w16667) | (w16666 & w16993) | (w16667 & w16993);
assign w17273 = ~w13208 & ~w13203;
assign w17274 = w13203 & ~w13364;
assign w17275 = ~w14524 & ~w14518;
assign w17276 = w14518 & ~w14645;
assign w17277 = ~w15755 & ~w15749;
assign w17278 = w15749 & ~w15827;
assign w17279 = ~w919 & ~w956;
assign w17280 = ~w1447 & ~w1435;
assign w17281 = ~w1576 & ~w1605;
assign w17282 = w866 & ~w855;
assign w17283 = w961 & ~w976;
assign w17284 = ~w1054 & ~w1078;
assign w17285 = w997 & ~w1049;
assign w17286 = ~w1223 & ~w1234;
assign w17287 = w1270 & ~w1259;
assign w17288 = ~w1346 & ~w1381;
assign w17289 = w1535 & ~w17041;
assign w17290 = w1535 & w1450;
assign w17291 = ~w1535 & w17041;
assign w17292 = ~w1535 & ~w1450;
assign w17293 = w1488 & ~w1477;
assign w17294 = ~w1676 & ~w1724;
assign w17295 = ~w1650 & ~w1653;
assign w17296 = w12688 & ~w16585;
assign w17297 = (w16590 & w16589) | (w16590 & w16585) | (w16589 & w16585);
assign w17298 = (w16592 & w16591) | (w16592 & ~w16585) | (w16591 & ~w16585);
assign w17299 = (w16597 & w16596) | (w16597 & w16585) | (w16596 & w16585);
assign w17300 = (~w16582 & w17440) | (~w16582 & w17441) | (w17440 & w17441);
assign w17301 = (w16599 & w16598) | (w16599 & ~w16585) | (w16598 & ~w16585);
assign w17302 = (w16582 & w17442) | (w16582 & w17443) | (w17442 & w17443);
assign w17303 = (w16603 & w16602) | (w16603 & w16585) | (w16602 & w16585);
assign w17304 = (w16603 & w16602) | (w16603 & w16584) | (w16602 & w16584);
assign w17305 = ~w13975 & ~w17228;
assign w17306 = ~w13975 & ~w17227;
assign w17307 = ~w14257 & ~w17230;
assign w17308 = ~w14257 & ~w17229;
assign w17309 = ~w14389 & ~w17232;
assign w17310 = ~w14389 & ~w17231;
assign w17311 = ~w14646 & ~w17234;
assign w17312 = ~w14646 & ~w17233;
assign w17313 = ~w14764 & ~w17236;
assign w17314 = ~w14764 & ~w17235;
assign w17315 = ~w14994 & ~w17242;
assign w17316 = ~w14994 & ~w17241;
assign w17317 = ~w15103 & ~w17244;
assign w17318 = ~w15103 & ~w17243;
assign w17319 = (~w16602 & w17702) | (~w16602 & w17703) | (w17702 & w17703);
assign w17320 = (w16632 & w16631) | (w16632 & w17246) | (w16631 & w17246);
assign w17321 = (~w16602 & w17704) | (~w16602 & w17705) | (w17704 & w17705);
assign w17322 = (w16638 & w16639) | (w16638 & w17246) | (w16639 & w17246);
assign w17323 = (~w16602 & w17706) | (~w16602 & w17707) | (w17706 & w17707);
assign w17324 = (w16654 & w16653) | (w16654 & w17246) | (w16653 & w17246);
assign w17325 = w16355 & w16996;
assign w17326 = w16355 & w16995;
assign w17327 = ~w16355 & ~w16996;
assign w17328 = ~w16355 & ~w16995;
assign w17329 = w16383 & w16998;
assign w17330 = w16383 & w16997;
assign w17331 = ~w16383 & ~w16998;
assign w17332 = ~w16383 & ~w16997;
assign w17333 = w16431 & w17000;
assign w17334 = w16431 & w16999;
assign w17335 = ~w16431 & ~w17000;
assign w17336 = ~w16431 & ~w16999;
assign w17337 = ~w1186 & w1185;
assign w17338 = ~w12140 & ~w12135;
assign w17339 = w11949 & w17708;
assign w17340 = w13203 & ~w13364;
assign w17341 = (~w13364 & w17274) | (~w13364 & w13208) | (w17274 & w13208);
assign w17342 = w13364 & w13681;
assign w17343 = w17276 & ~w14645;
assign w17344 = (~w14645 & w17276) | (~w14645 & w14524) | (w17276 & w14524);
assign w17345 = w14645 & w14885;
assign w17346 = ~w15827 & ~w17277;
assign w17347 = w15902 & w15827;
assign w17348 = w15902 & ~w17278;
assign w17349 = ~w11118 & ~w16571;
assign w17350 = (~w11118 & w16570) | (~w11118 & w17548) | (w16570 & w17548);
assign w17351 = (w11541 & w16573) | (w11541 & w16571) | (w16573 & w16571);
assign w17352 = (~w16570 & w17549) | (~w16570 & w17550) | (w17549 & w17550);
assign w17353 = (w16578 & w16577) | (w16578 & ~w16571) | (w16577 & ~w16571);
assign w17354 = (w16570 & w17551) | (w16570 & w17552) | (w17551 & w17552);
assign w17355 = (w16580 & w16579) | (w16580 & w16571) | (w16579 & w16571);
assign w17356 = (~w16570 & w17553) | (~w16570 & w17554) | (w17553 & w17554);
assign w17357 = (w16585 & w16584) | (w16585 & ~w16571) | (w16584 & ~w16571);
assign w17358 = (w16585 & w16584) | (w16585 & ~w16572) | (w16584 & ~w16572);
assign w17359 = (~w16582 & w17709) | (~w16582 & w17710) | (w17709 & w17710);
assign w17360 = ~w12507 & ~w17296;
assign w17361 = (w16582 & w17711) | (w16582 & w17712) | (w17711 & w17712);
assign w17362 = ~w12864 & ~w17297;
assign w17363 = (~w16582 & w17713) | (~w16582 & w17714) | (w17713 & w17714);
assign w17364 = ~w13035 & ~w17298;
assign w17365 = ~w13363 & ~w17299;
assign w17366 = ~w13525 & ~w17301;
assign w17367 = (~w16584 & w17444) | (~w16584 & w17445) | (w17444 & w17445);
assign w17368 = (~w16602 & w17715) | (~w16602 & w17444) | (w17715 & w17444);
assign w17369 = (~w16584 & w17446) | (~w16584 & w17447) | (w17446 & w17447);
assign w17370 = (~w16602 & w17716) | (~w16602 & w17446) | (w17716 & w17446);
assign w17371 = (~w16584 & w17448) | (~w16584 & w17449) | (w17448 & w17449);
assign w17372 = (~w16602 & w17717) | (~w16602 & w17448) | (w17717 & w17448);
assign w17373 = (~w16584 & w17450) | (~w16584 & w17451) | (w17450 & w17451);
assign w17374 = (~w16602 & w17718) | (~w16602 & w17450) | (w17718 & w17450);
assign w17375 = w15407 & w17252;
assign w17376 = w15407 & w17251;
assign w17377 = ~w15407 & ~w17252;
assign w17378 = ~w15407 & ~w17251;
assign w17379 = w15500 & w17254;
assign w17380 = w15500 & w17253;
assign w17381 = ~w15500 & ~w17254;
assign w17382 = ~w15500 & ~w17253;
assign w17383 = w15672 & w17256;
assign w17384 = w15672 & w17255;
assign w17385 = ~w15672 & ~w17256;
assign w17386 = ~w15672 & ~w17255;
assign w17387 = w15751 & w17258;
assign w17388 = w15751 & w17257;
assign w17389 = ~w15751 & ~w17258;
assign w17390 = ~w15751 & ~w17257;
assign w17391 = w15898 & w17260;
assign w17392 = w15898 & w17259;
assign w17393 = ~w15898 & ~w17260;
assign w17394 = ~w15898 & ~w17259;
assign w17395 = w15967 & w17262;
assign w17396 = w15967 & w17261;
assign w17397 = ~w15967 & ~w17262;
assign w17398 = ~w15967 & ~w17261;
assign w17399 = (w16986 & w16985) | (w16986 & ~w17304) | (w16985 & ~w17304);
assign w17400 = (w16988 & w16987) | (w16988 & ~w17304) | (w16987 & ~w17304);
assign w17401 = w16091 & ~w17264;
assign w17402 = w16091 & ~w17263;
assign w17403 = w16144 & w17266;
assign w17404 = w16144 & w17265;
assign w17405 = ~w16144 & ~w17266;
assign w17406 = ~w16144 & ~w17265;
assign w17407 = w16240 & w17268;
assign w17408 = w16240 & w17267;
assign w17409 = ~w16240 & ~w17268;
assign w17410 = ~w16240 & ~w17267;
assign w17411 = w16284 & w17270;
assign w17412 = w16284 & w17269;
assign w17413 = ~w16284 & ~w17270;
assign w17414 = ~w16284 & ~w17269;
assign w17415 = (w16994 & w16993) | (w16994 & ~w17304) | (w16993 & ~w17304);
assign w17416 = ~w16411 & w17272;
assign w17417 = ~w16411 & w17271;
assign w17418 = w16411 & ~w17272;
assign w17419 = w16411 & ~w17271;
assign w17420 = ~w10911 & w11121;
assign w17421 = w17339 & ~w12324;
assign w17422 = (~w12324 & w17339) | (~w12324 & w12140) | (w17339 & w12140);
assign w17423 = w13685 & ~w13681;
assign w17424 = (w13685 & ~w13681) | (w13685 & w17719) | (~w13681 & w17719);
assign w17425 = w14996 & ~w14885;
assign w17426 = w14996 & ~w17345;
assign w17427 = ~w15902 & w15971;
assign w17428 = w15971 & ~w17348;
assign w17429 = w15971 & ~w17347;
assign w17430 = ~w9659 & ~w9688;
assign w17431 = ~w9880 & ~w9861;
assign w17432 = ~w10147 & ~w10129;
assign w17433 = ~w10416 & ~w10454;
assign w17434 = ~w10640 & ~w10676;
assign w17435 = w12324 & w12688;
assign w17436 = w16589 & w16590;
assign w17437 = (w16590 & w16589) | (w16590 & ~w12324) | (w16589 & ~w12324);
assign w17438 = w16591 | w16592;
assign w17439 = (w16592 & w16591) | (w16592 & w12324) | (w16591 & w12324);
assign w17440 = w16596 & w16597;
assign w17441 = (w16597 & w16596) | (w16597 & ~w12324) | (w16596 & ~w12324);
assign w17442 = w16598 | w16599;
assign w17443 = (w16599 & w16598) | (w16599 & w12324) | (w16598 & w12324);
assign w17444 = ~w13832 & ~w16603;
assign w17445 = (~w13832 & w16600) | (~w13832 & w17720) | (w16600 & w17720);
assign w17446 = (w16605 & w16606) | (w16605 & ~w16603) | (w16606 & ~w16603);
assign w17447 = (w16600 & w17721) | (w16600 & w17722) | (w17721 & w17722);
assign w17448 = (w16612 & w16613) | (w16612 & ~w16603) | (w16613 & ~w16603);
assign w17449 = (w16600 & w17723) | (w16600 & w17724) | (w17723 & w17724);
assign w17450 = (w16620 & w16619) | (w16620 & ~w16603) | (w16619 & ~w16603);
assign w17451 = (w16600 & w17725) | (w16600 & w17726) | (w17725 & w17726);
assign w17452 = w9743 & ~w9733;
assign w17453 = (w10013 & w16561) | (w10013 & w17555) | (w16561 & w17555);
assign w17454 = (~w16559 & w17555) | (~w16559 & w17727) | (w17555 & w17727);
assign w17455 = w9946 & ~w9934;
assign w17456 = (~w10233 & w10097) | (~w10233 & w17556) | (w10097 & w17556);
assign w17457 = (~w10090 & ~w10056) | (~w10090 & w17557) | (~w10056 & w17557);
assign w17458 = w10126 & ~w10115;
assign w17459 = ~w10202 & ~w10222;
assign w17460 = (~w10403 & w10404) | (~w10403 & w17558) | (w10404 & w17558);
assign w17461 = (~w10332 & w10298) | (~w10332 & w17559) | (w10298 & w17559);
assign w17462 = w10363 & ~w10351;
assign w17463 = w10372 & w10529;
assign w17464 = ~w10372 & ~w10529;
assign w17465 = (~w16561 & w17560) | (~w16561 & w17561) | (w17560 & w17561);
assign w17466 = (w16566 & w16567) | (w16566 & w16562) | (w16567 & w16562);
assign w17467 = (~w10627 & w10628) | (~w10627 & w17562) | (w10628 & w17562);
assign w17468 = (~w10556 & w10524) | (~w10556 & w17563) | (w10524 & w17563);
assign w17469 = ~w10547 & ~w10543;
assign w17470 = w10673 & ~w10662;
assign w17471 = w10501 & w10797;
assign w17472 = ~w10501 & ~w10797;
assign w17473 = (w16568 & w16569) | (w16568 & ~w16562) | (w16569 & ~w16562);
assign w17474 = ~w10755 & ~w10758;
assign w17475 = (w16572 & w16571) | (w16572 & ~w16563) | (w16571 & ~w16563);
assign w17476 = (w16572 & w16571) | (w16572 & ~w16562) | (w16571 & ~w16562);
assign w17477 = ~w11119 & ~w17350;
assign w17478 = ~w11119 & ~w17349;
assign w17479 = ~w11333 & ~w17352;
assign w17480 = ~w11333 & ~w17351;
assign w17481 = ~w11742 & ~w17354;
assign w17482 = ~w11742 & ~w17353;
assign w17483 = ~w11940 & ~w17356;
assign w17484 = ~w11940 & ~w17355;
assign w17485 = ~w12323 & ~w17358;
assign w17486 = (~w16584 & w17564) | (~w16584 & w17565) | (w17564 & w17565);
assign w17487 = (w16587 & w16588) | (w16587 & ~w17358) | (w16588 & ~w17358);
assign w17488 = (~w16584 & w17566) | (~w16584 & w17567) | (w17566 & w17567);
assign w17489 = (w16594 & w16595) | (w16594 & ~w17358) | (w16595 & ~w17358);
assign w17490 = (~w16584 & w17568) | (~w16584 & w17569) | (w17568 & w17569);
assign w17491 = (w16601 & w16600) | (w16601 & ~w17358) | (w16600 & ~w17358);
assign w17492 = (~w16584 & w17570) | (~w16584 & w17571) | (w17570 & w17571);
assign w17493 = w14121 & w17306;
assign w17494 = w14121 & w17305;
assign w17495 = ~w14121 & ~w17306;
assign w17496 = ~w14121 & ~w17305;
assign w17497 = w14390 & w17308;
assign w17498 = w14390 & w17307;
assign w17499 = ~w14390 & ~w17308;
assign w17500 = ~w14390 & ~w17307;
assign w17501 = w14519 & w17310;
assign w17502 = w14519 & w17309;
assign w17503 = ~w14519 & ~w17310;
assign w17504 = ~w14519 & ~w17309;
assign w17505 = w14766 & w17312;
assign w17506 = w14766 & w17311;
assign w17507 = ~w14766 & ~w17312;
assign w17508 = ~w14766 & ~w17311;
assign w17509 = w14884 & w17314;
assign w17510 = w14884 & w17313;
assign w17511 = ~w14884 & ~w17314;
assign w17512 = ~w14884 & ~w17313;
assign w17513 = w15105 & w17316;
assign w17514 = w15105 & w17315;
assign w17515 = ~w15105 & ~w17316;
assign w17516 = ~w15105 & ~w17315;
assign w17517 = w15208 & w17318;
assign w17518 = w15208 & w17317;
assign w17519 = ~w15208 & ~w17318;
assign w17520 = ~w15208 & ~w17317;
assign w17521 = (w17247 & w17246) | (w17247 & ~w17358) | (w17246 & ~w17358);
assign w17522 = (w17247 & w17246) | (w17247 & ~w17357) | (w17246 & ~w17357);
assign w17523 = w15587 & w17320;
assign w17524 = w15587 & w17319;
assign w17525 = ~w15587 & ~w17320;
assign w17526 = ~w15587 & ~w17319;
assign w17527 = ~w15828 & w17322;
assign w17528 = ~w15828 & w17321;
assign w17529 = w15828 & ~w17322;
assign w17530 = w15828 & ~w17321;
assign w17531 = ~w16195 & w17324;
assign w17532 = ~w16195 & w17323;
assign w17533 = w16195 & ~w17324;
assign w17534 = w16195 & ~w17323;
assign w17535 = w9532 & ~w9770;
assign w17536 = ~w11121 & ~w10908;
assign w17537 = ~w13679 & ~w17423;
assign w17538 = ~w13679 & ~w17424;
assign w17539 = w13679 & ~w13831;
assign w17540 = ~w14882 & ~w14996;
assign w17541 = ~w14882 & ~w17425;
assign w17542 = w14993 & w15109;
assign w17543 = ~w15966 & ~w15971;
assign w17544 = ~w15966 & ~w17427;
assign w17545 = w15966 & ~w16027;
assign w17546 = ~w7539 & ~w7575;
assign w17547 = w8745 & ~w8743;
assign w17548 = w10908 & ~w11118;
assign w17549 = w16573 & w11541;
assign w17550 = (w11541 & w16573) | (w11541 & ~w10908) | (w16573 & ~w10908);
assign w17551 = w16577 | w16578;
assign w17552 = (w16578 & w16577) | (w16578 & w10908) | (w16577 & w10908);
assign w17553 = w16579 & w16580;
assign w17554 = (w16580 & w16579) | (w16580 & ~w10908) | (w16579 & ~w10908);
assign w17555 = w9770 & w10013;
assign w17556 = ~w10154 & ~w10233;
assign w17557 = ~w10055 & ~w10090;
assign w17558 = ~w10457 & ~w10403;
assign w17559 = ~w10297 & ~w10332;
assign w17560 = w16567 & w16566;
assign w17561 = (w16566 & w16567) | (w16566 & ~w9770) | (w16567 & ~w9770);
assign w17562 = ~w10679 & ~w10627;
assign w17563 = ~w10523 & ~w10556;
assign w17564 = ~w12323 & w16571;
assign w17565 = ~w12323 & ~w16585;
assign w17566 = (w16587 & w16588) | (w16587 & w16571) | (w16588 & w16571);
assign w17567 = (w16587 & w16588) | (w16587 & ~w16585) | (w16588 & ~w16585);
assign w17568 = (w16594 & w16595) | (w16594 & w16571) | (w16595 & w16571);
assign w17569 = (w16594 & w16595) | (w16594 & ~w16585) | (w16595 & ~w16585);
assign w17570 = (w16600 & w16601) | (w16600 & w16571) | (w16601 & w16571);
assign w17571 = (w16600 & w16601) | (w16600 & ~w16585) | (w16601 & ~w16585);
assign w17572 = w7015 & ~w7018;
assign w17573 = pi31 & ~w7654;
assign w17574 = ~pi31 & w7654;
assign w17575 = w7669 & ~w7680;
assign w17576 = w7723 & ~w7713;
assign w17577 = w7794 & ~w17145;
assign w17578 = w7794 & w7540;
assign w17579 = ~w7794 & w17145;
assign w17580 = ~w7794 & ~w7540;
assign w17581 = w7536 & ~w7526;
assign w17582 = w7785 & ~w7789;
assign w17583 = ~w7967 & ~w7963;
assign w17584 = ~w7837 & ~w7906;
assign w17585 = w8119 & ~w8109;
assign w17586 = w8201 & ~w8204;
assign w17587 = ~w8308 & ~w8327;
assign w17588 = (~w8332 & w8333) | (~w8332 & w17728) | (w8333 & w17728);
assign w17589 = w8437 & ~w8426;
assign w17590 = ~w8751 & ~w8774;
assign w17591 = w8697 & ~w8685;
assign w17592 = ~w8700 & ~w8663;
assign w17593 = ~w8915 & ~w8918;
assign w17594 = w8861 & ~w8850;
assign w17595 = w8952 & ~w8941;
assign w17596 = (~w9020 & w9022) | (~w9020 & w17729) | (w9022 & w17729);
assign w17597 = ~w9041 & ~w16557;
assign w17598 = (~w9041 & w16555) | (~w9041 & w17730) | (w16555 & w17730);
assign w17599 = ~w9263 & ~w9266;
assign w17600 = w9177 & ~w9166;
assign w17601 = w9209 & ~w9198;
assign w17602 = w9255 & ~w9258;
assign w17603 = (w9535 & w16558) | (w9535 & w16557) | (w16558 & w16557);
assign w17604 = (~w16555 & w17731) | (~w16555 & w17732) | (w17731 & w17732);
assign w17605 = (w16562 & w16563) | (w16562 & ~w16557) | (w16563 & ~w16557);
assign w17606 = (w16562 & w16563) | (w16562 & ~w16556) | (w16563 & ~w16556);
assign w17607 = (w17454 & w17453) | (w17454 & w16557) | (w17453 & w16557);
assign w17608 = (w17454 & w17453) | (w17454 & w16556) | (w17453 & w16556);
assign w17609 = w10323 & ~w10319;
assign w17610 = w10279 & w10559;
assign w17611 = ~w10279 & ~w10559;
assign w17612 = (w17466 & w17465) | (w17466 & ~w16557) | (w17465 & ~w16557);
assign w17613 = (w17466 & w17465) | (w17466 & ~w16556) | (w17465 & ~w16556);
assign w17614 = w10587 & ~w10576;
assign w17615 = w10535 & ~w10531;
assign w17616 = w10528 & ~w10551;
assign w17617 = w10515 & ~w10518;
assign w17618 = w10506 & w10763;
assign w17619 = ~w10506 & ~w10763;
assign w17620 = ~w10693 & ~w17473;
assign w17621 = (w16563 & w17733) | (w16563 & w17734) | (w17733 & w17734);
assign w17622 = w10720 & w10962;
assign w17623 = ~w10720 & ~w10962;
assign w17624 = w10703 & ~w10706;
assign w17625 = (~w10503 & w17735) | (~w10503 & w17736) | (w17735 & w17736);
assign w17626 = ~w10778 & ~w10793;
assign w17627 = w11063 & ~w11105;
assign w17628 = (w16572 & w17737) | (w16572 & w17738) | (w17737 & w17738);
assign w17629 = (w16576 & w16575) | (w16576 & w17475) | (w16575 & w17475);
assign w17630 = (w16582 & w16583) | (w16582 & w17476) | (w16583 & w17476);
assign w17631 = (w16582 & w16583) | (w16582 & w17475) | (w16583 & w17475);
assign w17632 = (w17360 & w17359) | (w17360 & ~w17476) | (w17359 & ~w17476);
assign w17633 = (w17360 & w17359) | (w17360 & ~w17475) | (w17359 & ~w17475);
assign w17634 = (w17362 & w17361) | (w17362 & w17476) | (w17361 & w17476);
assign w17635 = (w17362 & w17361) | (w17362 & w17475) | (w17361 & w17475);
assign w17636 = (w17364 & w17363) | (w17364 & ~w17476) | (w17363 & ~w17476);
assign w17637 = (w17364 & w17363) | (w17364 & ~w17475) | (w17363 & ~w17475);
assign w17638 = w13526 & w17365;
assign w17639 = ~w17300 & w17739;
assign w17640 = ~w13526 & ~w17365;
assign w17641 = (~w13526 & w17300) | (~w13526 & w17740) | (w17300 & w17740);
assign w17642 = w13680 & w17366;
assign w17643 = ~w17302 & w17741;
assign w17644 = ~w13680 & ~w17366;
assign w17645 = (~w13680 & w17302) | (~w13680 & w17742) | (w17302 & w17742);
assign w17646 = (w17304 & w17303) | (w17304 & ~w17476) | (w17303 & ~w17476);
assign w17647 = (w17304 & w17303) | (w17304 & ~w17475) | (w17303 & ~w17475);
assign w17648 = w13977 & w17368;
assign w17649 = w13977 & w17367;
assign w17650 = ~w13977 & ~w17368;
assign w17651 = ~w13977 & ~w17367;
assign w17652 = ~w14258 & w17370;
assign w17653 = ~w14258 & w17369;
assign w17654 = w14258 & ~w17370;
assign w17655 = w14258 & ~w17369;
assign w17656 = ~w14647 & w17372;
assign w17657 = ~w14647 & w17371;
assign w17658 = w14647 & ~w17372;
assign w17659 = w14647 & ~w17371;
assign w17660 = w14995 & w17374;
assign w17661 = w14995 & w17373;
assign w17662 = ~w14995 & ~w17374;
assign w17663 = ~w14995 & ~w17373;
assign w17664 = (w17303 & w17743) | (w17303 & w17744) | (w17743 & w17744);
assign w17665 = (w17304 & w17743) | (w17304 & w17744) | (w17743 & w17744);
assign w17666 = (~w17303 & w17745) | (~w17303 & w17746) | (w17745 & w17746);
assign w17667 = w16029 & w17399;
assign w17668 = (~w17303 & w17747) | (~w17303 & w17748) | (w17747 & w17748);
assign w17669 = ~w16086 & w17400;
assign w17670 = (~w17303 & w17749) | (~w17303 & w17750) | (w17749 & w17750);
assign w17671 = (~w17304 & w17749) | (~w17304 & w17750) | (w17749 & w17750);
assign w17672 = (w17303 & w17751) | (w17303 & w17752) | (w17751 & w17752);
assign w17673 = w16321 & ~w17415;
assign w17674 = ~w13679 & ~w13685;
assign w17675 = (~w13831 & w17539) | (~w13831 & w13685) | (w17539 & w13685);
assign w17676 = (~w13831 & w17539) | (~w13831 & w17423) | (w17539 & w17423);
assign w17677 = w17542 & w15109;
assign w17678 = (w15109 & w17542) | (w15109 & ~w14882) | (w17542 & ~w14882);
assign w17679 = ~w16027 & ~w17543;
assign w17680 = ~w16027 & ~w17544;
assign w17681 = (~w16027 & w17545) | (~w16027 & w17429) | (w17545 & w17429);
assign w17682 = (~w16027 & w17545) | (~w16027 & w17428) | (w17545 & w17428);
assign w17683 = w6747 & ~w6745;
assign w17684 = ~w6878 & ~w6914;
assign w17685 = ~w7197 & ~w7234;
assign w17686 = ~w11290 & ~w11320;
assign w17687 = ~w11719 & ~w11708;
assign w17688 = w12118 & ~w12116;
assign w17689 = w13831 & w13982;
assign w17690 = w16608 & w16607;
assign w17691 = (w16607 & w16608) | (w16607 & ~w13831) | (w16608 & ~w13831);
assign w17692 = w16609 | w16610;
assign w17693 = (w16610 & w16609) | (w16610 & w13831) | (w16609 & w13831);
assign w17694 = w16614 & w16615;
assign w17695 = (w16615 & w16614) | (w16615 & ~w13831) | (w16614 & ~w13831);
assign w17696 = w16616 | w16617;
assign w17697 = (w16617 & w16616) | (w16617 & w13831) | (w16616 & w13831);
assign w17698 = w16621 & w16622;
assign w17699 = (w16622 & w16621) | (w16622 & ~w13831) | (w16621 & ~w13831);
assign w17700 = w16623 | w16624;
assign w17701 = (w16624 & w16623) | (w16624 & w13831) | (w16623 & w13831);
assign w17702 = (w16632 & w16631) | (w16632 & w16628) | (w16631 & w16628);
assign w17703 = (w16632 & w16631) | (w16632 & w16627) | (w16631 & w16627);
assign w17704 = (w16638 & w16639) | (w16638 & w16628) | (w16639 & w16628);
assign w17705 = (w16638 & w16639) | (w16638 & w16627) | (w16639 & w16627);
assign w17706 = (w16654 & w16653) | (w16654 & w16628) | (w16653 & w16628);
assign w17707 = (w16654 & w16653) | (w16654 & w16627) | (w16653 & w16627);
assign w17708 = ~w12133 & ~w12324;
assign w17709 = ~w12507 & ~w12688;
assign w17710 = ~w12507 & ~w17435;
assign w17711 = ~w12864 & ~w17437;
assign w17712 = ~w12864 & ~w17436;
assign w17713 = ~w13035 & ~w17439;
assign w17714 = ~w13035 & ~w17438;
assign w17715 = ~w13832 & ~w16585;
assign w17716 = (w16605 & w16606) | (w16605 & ~w16585) | (w16606 & ~w16585);
assign w17717 = (w16612 & w16613) | (w16612 & ~w16585) | (w16613 & ~w16585);
assign w17718 = (w16620 & w16619) | (w16620 & ~w16585) | (w16619 & ~w16585);
assign w17719 = ~w13364 & w13685;
assign w17720 = w13831 & ~w13832;
assign w17721 = w16606 | w16605;
assign w17722 = (w16605 & w16606) | (w16605 & w13831) | (w16606 & w13831);
assign w17723 = w16613 | w16612;
assign w17724 = (w16612 & w16613) | (w16612 & w13831) | (w16613 & w13831);
assign w17725 = w16619 | w16620;
assign w17726 = (w16620 & w16619) | (w16620 & w13831) | (w16619 & w13831);
assign w17727 = w10013 & ~w17535;
assign w17728 = w8334 & ~w8332;
assign w17729 = w9021 & ~w9020;
assign w17730 = w8789 & ~w9041;
assign w17731 = w16558 & w9535;
assign w17732 = (w9535 & w16558) | (w9535 & ~w8789) | (w16558 & ~w8789);
assign w17733 = ~w10693 & ~w16568;
assign w17734 = ~w10693 & ~w16569;
assign w17735 = ~w10898 & ~w10797;
assign w17736 = ~w10898 & ~w17471;
assign w17737 = (w16576 & w16575) | (w16576 & ~w16562) | (w16575 & ~w16562);
assign w17738 = (w16576 & w16575) | (w16576 & w16571) | (w16575 & w16571);
assign w17739 = ~w13363 & w13526;
assign w17740 = w13363 & ~w13526;
assign w17741 = ~w13525 & w13680;
assign w17742 = w13525 & ~w13680;
assign w17743 = ~w16029 & ~w16986;
assign w17744 = ~w16029 & ~w16985;
assign w17745 = w16029 & w16986;
assign w17746 = w16029 & w16985;
assign w17747 = ~w16086 & w16988;
assign w17748 = ~w16086 & w16987;
assign w17749 = ~w16321 & w16994;
assign w17750 = ~w16321 & w16993;
assign w17751 = w16321 & ~w16994;
assign w17752 = w16321 & ~w16993;
assign w17753 = w6234 & ~w6223;
assign w17754 = ~w6156 & ~w6159;
assign w17755 = w6429 & ~w6418;
assign w17756 = w6396 & ~w6386;
assign w17757 = ~w6636 & ~w6601;
assign w17758 = w6708 & ~w6697;
assign w17759 = w6633 & ~w6622;
assign w17760 = ~w6993 & ~w6918;
assign w17761 = ~w6860 & ~w6827;
assign w17762 = w6839 & ~w6835;
assign w17763 = w6950 & ~w6939;
assign w17764 = w6777 & ~w6789;
assign w17765 = ~w7049 & ~w7095;
assign w17766 = ~w7448 & ~w7481;
assign w17767 = ~w7355 & ~w7422;
assign w17768 = ~w7418 & ~w7391;
assign w17769 = w7459 & ~w7455;
assign w17770 = ~w7471 & ~w7467;
assign w17771 = w7450 & ~w7475;
assign w17772 = w7615 & ~w7611;
assign w17773 = w7606 & ~w7631;
assign w17774 = w7505 & ~w7579;
assign w17775 = (~w8007 & w16550) | (~w8007 & w16549) | (w16550 & w16549);
assign w17776 = (~w8007 & w16550) | (~w8007 & w16548) | (w16550 & w16548);
assign w17777 = ~w7784 & ~w7795;
assign w17778 = ~w8253 & ~w8221;
assign w17779 = w8016 & ~w8082;
assign w17780 = ~w8072 & ~w8075;
assign w17781 = (w16553 & w16554) | (w16553 & w16549) | (w16554 & w16549);
assign w17782 = (w16553 & w16554) | (w16553 & w16548) | (w16554 & w16548);
assign w17783 = ~w8340 & ~w8297;
assign w17784 = ~w8440 & ~w8405;
assign w17785 = ~w8283 & ~w8279;
assign w17786 = w8482 & ~w8478;
assign w17787 = w8473 & ~w8498;
assign w17788 = w8291 & ~w8289;
assign w17789 = (w16557 & w16556) | (w16557 & w16549) | (w16556 & w16549);
assign w17790 = (w16557 & w16556) | (w16557 & w16548) | (w16556 & w16548);
assign w17791 = ~w8570 & ~w8573;
assign w17792 = ~w8549 & ~w8545;
assign w17793 = ~w8561 & ~w8557;
assign w17794 = w9251 & ~w17596;
assign w17795 = w9251 & w9023;
assign w17796 = ~w9251 & w17596;
assign w17797 = ~w9251 & ~w9023;
assign w17798 = w8971 & ~w8967;
assign w17799 = ~w8999 & ~w9029;
assign w17800 = ~w9042 & ~w17598;
assign w17801 = ~w9042 & ~w17597;
assign w17802 = ~w9071 & ~w9094;
assign w17803 = w9051 & ~w9054;
assign w17804 = ~w9286 & ~w17604;
assign w17805 = ~w9286 & ~w17603;
assign w17806 = ~w9437 & ~w9440;
assign w17807 = ~w9482 & ~w9519;
assign w17808 = ~w9620 & ~w9571;
assign w17809 = w9543 & ~w9565;
assign w17810 = ~w9771 & ~w17606;
assign w17811 = ~w9771 & ~w17605;
assign w17812 = ~w10005 & ~w17608;
assign w17813 = ~w10005 & ~w17607;
assign w17814 = (w16564 & w16565) | (w16564 & ~w17606) | (w16565 & ~w17606);
assign w17815 = (w16564 & w16565) | (w16564 & ~w17605) | (w16565 & ~w17605);
assign w17816 = w10451 & ~w10439;
assign w17817 = w10394 & ~w10385;
assign w17818 = ~w10471 & ~w17613;
assign w17819 = ~w10471 & ~w17612;
assign w17820 = ~w10685 & ~w10560;
assign w17821 = ~w10826 & ~w10893;
assign w17822 = ~w10711 & ~w10714;
assign w17823 = ~w10901 & ~w10764;
assign w17824 = ~w11059 & ~w10963;
assign w17825 = ~w11053 & ~w11018;
assign w17826 = (w17478 & w17477) | (w17478 & ~w17606) | (w17477 & ~w17606);
assign w17827 = (w17478 & w17477) | (w17478 & ~w17605) | (w17477 & ~w17605);
assign w17828 = ~w11326 & ~w11228;
assign w17829 = w11162 & ~w11150;
assign w17830 = w11287 & ~w11275;
assign w17831 = (w17480 & w17479) | (w17480 & w17606) | (w17479 & w17606);
assign w17832 = (w17480 & w17479) | (w17480 & w17605) | (w17479 & w17605);
assign w17833 = w11374 & ~w11363;
assign w17834 = (w17482 & w17481) | (w17482 & ~w17606) | (w17481 & ~w17606);
assign w17835 = (w17482 & w17481) | (w17482 & ~w17605) | (w17481 & ~w17605);
assign w17836 = (w17484 & w17483) | (w17484 & w17606) | (w17483 & w17606);
assign w17837 = (w17484 & w17483) | (w17484 & w17605) | (w17483 & w17605);
assign w17838 = ~w11824 & ~w11793;
assign w17839 = w11924 & w12050;
assign w17840 = ~w11924 & ~w12050;
assign w17841 = w12041 & ~w12030;
assign w17842 = w12008 & ~w11997;
assign w17843 = ~w11962 & ~w11980;
assign w17844 = ~w12104 & ~w12082;
assign w17845 = w12108 & ~w12111;
assign w17846 = (w17358 & w17357) | (w17358 & w17606) | (w17357 & w17606);
assign w17847 = (w17358 & w17357) | (w17358 & w17605) | (w17357 & w17605);
assign w17848 = w12240 & ~w12311;
assign w17849 = w12509 & w17486;
assign w17850 = w12509 & w17485;
assign w17851 = ~w12509 & ~w17486;
assign w17852 = ~w12509 & ~w17485;
assign w17853 = ~w12866 & w17488;
assign w17854 = ~w12866 & w17487;
assign w17855 = w12866 & ~w17488;
assign w17856 = w12866 & ~w17487;
assign w17857 = ~w13365 & w17490;
assign w17858 = ~w13365 & w17489;
assign w17859 = w13365 & ~w17490;
assign w17860 = w13365 & ~w17489;
assign w17861 = ~w13833 & w17492;
assign w17862 = ~w13833 & w17491;
assign w17863 = w13833 & ~w17492;
assign w17864 = w13833 & ~w17491;
assign w17865 = ~w15312 & w17522;
assign w17866 = ~w15312 & w17521;
assign w17867 = w15312 & ~w17522;
assign w17868 = w15312 & ~w17521;
assign w17869 = (w17002 & w17001) | (w17002 & ~w17522) | (w17001 & ~w17522);
assign w17870 = (w17002 & w17001) | (w17002 & ~w17521) | (w17001 & ~w17521);
assign w17871 = (w17004 & w17003) | (w17004 & w17522) | (w17003 & w17522);
assign w17872 = (w17004 & w17003) | (w17004 & w17521) | (w17003 & w17521);
assign w17873 = (w17006 & w17005) | (w17006 & w17522) | (w17005 & w17522);
assign w17874 = (w17006 & w17005) | (w17006 & w17521) | (w17005 & w17521);
assign w17875 = (w17008 & w17007) | (w17008 & ~w17522) | (w17007 & ~w17522);
assign w17876 = (w17008 & w17007) | (w17008 & ~w17521) | (w17007 & ~w17521);
assign w17877 = (w17010 & w17009) | (w17010 & w17522) | (w17009 & w17522);
assign w17878 = (w17010 & w17009) | (w17010 & w17521) | (w17009 & w17521);
assign w17879 = (w17012 & w17011) | (w17012 & ~w17522) | (w17011 & ~w17522);
assign w17880 = (w17012 & w17011) | (w17012 & ~w17521) | (w17011 & ~w17521);
assign w17881 = (w17014 & w17013) | (w17014 & w17522) | (w17013 & w17522);
assign w17882 = (w17014 & w17013) | (w17014 & w17521) | (w17013 & w17521);
assign w17883 = (w17016 & w17015) | (w17016 & ~w17522) | (w17015 & ~w17522);
assign w17884 = (w17016 & w17015) | (w17016 & ~w17521) | (w17015 & ~w17521);
assign w17885 = (w17018 & w17017) | (w17018 & ~w17522) | (w17017 & ~w17522);
assign w17886 = (w17018 & w17017) | (w17018 & ~w17521) | (w17017 & ~w17521);
assign one = 1;
assign po000 = pi00;// level 0
assign po001 = w0;// level 1
assign po002 = w4;// level 3
assign po003 = w10;// level 4
assign po004 = ~w22;// level 7
assign po005 = w38;// level 8
assign po006 = ~w55;// level 9
assign po007 = w83;// level 11
assign po008 = ~w114;// level 12
assign po009 = w151;// level 13
assign po010 = w188;// level 15
assign po011 = ~w234;// level 16
assign po012 = ~w282;// level 16
assign po013 = w336;// level 18
assign po014 = ~w391;// level 19
assign po015 = ~w453;// level 19
assign po016 = w517;// level 21
assign po017 = ~w588;// level 20
assign po018 = ~w660;// level 20
assign po019 = w739;// level 22
assign po020 = ~w820;// level 23
assign po021 = w907;// level 23
assign po022 = w995;// level 23
assign po023 = ~w1092;// level 24
assign po024 = ~w1190;// level 24
assign po025 = w1290;// level 26
assign po026 = ~w1398;// level 26
assign po027 = w1510;// level 26
assign po028 = w1622;// level 26
assign po029 = ~w1744;// level 27
assign po030 = w1867;// level 27
assign po031 = w1992;// level 29
assign po032 = ~w2126;// level 29
assign po033 = w2264;// level 29
assign po034 = w2401;// level 30
assign po035 = ~w2548;// level 30
assign po036 = w2694;// level 29
assign po037 = w2846;// level 31
assign po038 = ~w3002;// level 31
assign po039 = w3164;// level 30
assign po040 = w3327;// level 32
assign po041 = ~w3499;// level 32
assign po042 = ~w3669;// level 32
assign po043 = w3845;// level 33
assign po044 = ~w4028;// level 34
assign po045 = ~w4214;// level 33
assign po046 = ~w4403;// level 34
assign po047 = ~w4599;// level 35
assign po048 = ~w4797;// level 34
assign po049 = w5001;// level 36
assign po050 = ~w5205;// level 36
assign po051 = w5418;// level 35
assign po052 = w5634;// level 36
assign po053 = ~w5851;// level 37
assign po054 = w6074;// level 36
assign po055 = w6302;// level 37
assign po056 = ~w6533;// level 38
assign po057 = w6773;// level 37
assign po058 = w7010;// level 38
assign po059 = ~w7256;// level 39
assign po060 = w7503;// level 38
assign po061 = w7752;// level 39
assign po062 = ~w8011;// level 39
assign po063 = w8274;// level 38
assign po064 = w8534;// level 39
assign po065 = ~w8793;// level 39
assign po066 = ~w9046;// level 38
assign po067 = w9292;// level 39
assign po068 = ~w9539;// level 39
assign po069 = w9777;// level 39
assign po070 = w10012;// level 39
assign po071 = ~w10248;// level 39
assign po072 = ~w10476;// level 39
assign po073 = w10698;// level 39
assign po074 = ~w10915;// level 39
assign po075 = w11125;// level 39
assign po076 = w11339;// level 39
assign po077 = ~w11545;// level 39
assign po078 = ~w11746;// level 39
assign po079 = w11946;// level 39
assign po080 = ~w12139;// level 39
assign po081 = ~w12328;// level 39
assign po082 = w12512;// level 39
assign po083 = ~w12692;// level 39
assign po084 = ~w12869;// level 39
assign po085 = w13040;// level 39
assign po086 = ~w13207;// level 39
assign po087 = ~w13368;// level 39
assign po088 = w13529;// level 39
assign po089 = ~w13684;// level 39
assign po090 = ~w13836;// level 39
assign po091 = w13981;// level 39
assign po092 = ~w14124;// level 39
assign po093 = ~w14261;// level 39
assign po094 = w14393;// level 39
assign po095 = ~w14523;// level 39
assign po096 = ~w14650;// level 39
assign po097 = w14769;// level 39
assign po098 = ~w14888;// level 39
assign po099 = w14999;// level 39
assign po100 = w15108;// level 39
assign po101 = ~w15211;// level 39
assign po102 = ~w15315;// level 39
assign po103 = w15410;// level 39
assign po104 = ~w15503;// level 39
assign po105 = w15591;// level 39
assign po106 = w15675;// level 39
assign po107 = ~w15754;// level 39
assign po108 = ~w15831;// level 39
assign po109 = w15901;// level 39
assign po110 = ~w15970;// level 39
assign po111 = w16032;// level 39
assign po112 = w16093;// level 39
assign po113 = ~w16147;// level 39
assign po114 = ~w16198;// level 39
assign po115 = w16243;// level 39
assign po116 = ~w16287;// level 39
assign po117 = ~w16324;// level 39
assign po118 = w16358;// level 40
assign po119 = ~w16387;// level 40
assign po120 = ~w16414;// level 39
assign po121 = w16434;// level 40
assign po122 = ~w16453;// level 39
assign po123 = ~w16465;// level 39
assign po124 = ~w16473;// level 39
assign po125 = ~w16479;// level 39
assign po126 = w16481;// level 39
endmodule
