module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 , x147 , x148 , x149 , x150 , x151 , x152 , x153 , x154 , x155 , x156 , x157 , x158 , x159 , x160 , x161 , x162 , x163 , x164 , x165 , x166 , x167 , x168 , x169 , x170 , x171 , x172 , x173 , x174 , x175 , x176 , x177 , x178 , x179 , x180 , x181 , x182 , x183 , x184 , x185 , x186 , x187 , x188 , x189 , x190 , x191 , x192 , x193 , x194 , x195 , x196 , x197 , x198 , x199 , x200 , x201 , x202 , x203 , x204 , x205 , x206 , x207 , x208 , x209 , x210 , x211 , x212 , x213 , x214 , x215 , x216 , x217 , x218 , x219 , x220 , x221 , x222 , x223 , x224 , x225 , x226 , x227 , x228 , x229 , x230 , x231 , x232 , x233 , x234 , x235 , x236 , x237 , x238 , x239 , x240 , x241 , x242 , x243 , x244 , x245 , x246 , x247 , x248 , x249 , x250 , x251 , x252 , x253 , x254 , x255 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 , x147 , x148 , x149 , x150 , x151 , x152 , x153 , x154 , x155 , x156 , x157 , x158 , x159 , x160 , x161 , x162 , x163 , x164 , x165 , x166 , x167 , x168 , x169 , x170 , x171 , x172 , x173 , x174 , x175 , x176 , x177 , x178 , x179 , x180 , x181 , x182 , x183 , x184 , x185 , x186 , x187 , x188 , x189 , x190 , x191 , x192 , x193 , x194 , x195 , x196 , x197 , x198 , x199 , x200 , x201 , x202 , x203 , x204 , x205 , x206 , x207 , x208 , x209 , x210 , x211 , x212 , x213 , x214 , x215 , x216 , x217 , x218 , x219 , x220 , x221 , x222 , x223 , x224 , x225 , x226 , x227 , x228 , x229 , x230 , x231 , x232 , x233 , x234 , x235 , x236 , x237 , x238 , x239 , x240 , x241 , x242 , x243 , x244 , x245 , x246 , x247 , x248 , x249 , x250 , x251 , x252 , x253 , x254 , x255 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 ;
  wire n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 ;
  assign n257 = x0 & x64 ;
  assign n258 = x0 | x64 ;
  assign n259 = ~n257 & n258 ;
  assign n260 = x128 & n259 ;
  assign n261 = x128 | n259 ;
  assign n262 = ~n260 & n261 ;
  assign n263 = x192 & n262 ;
  assign n264 = x192 | n262 ;
  assign n265 = ~n263 & n264 ;
  assign n266 = n257 | n260 ;
  assign n267 = x193 & n266 ;
  assign n268 = x193 | n266 ;
  assign n269 = ~n267 & n268 ;
  assign n270 = x1 & x65 ;
  assign n271 = x1 | x65 ;
  assign n272 = ~n270 & n271 ;
  assign n273 = x129 & n272 ;
  assign n274 = x129 | n272 ;
  assign n275 = ~n273 & n274 ;
  assign n276 = n269 & n275 ;
  assign n277 = n269 | n275 ;
  assign n278 = ~n276 & n277 ;
  assign n279 = n263 | n278 ;
  assign n280 = n263 & n278 ;
  assign n281 = n279 & ~n280 ;
  assign n282 = n267 | n276 ;
  assign n283 = n270 | n273 ;
  assign n284 = x194 & n283 ;
  assign n285 = x194 | n283 ;
  assign n286 = ~n284 & n285 ;
  assign n287 = x2 & x66 ;
  assign n288 = x2 | x66 ;
  assign n289 = ~n287 & n288 ;
  assign n290 = x130 & n289 ;
  assign n291 = x130 | n289 ;
  assign n292 = ~n290 & n291 ;
  assign n293 = n286 | n292 ;
  assign n294 = n286 & n292 ;
  assign n295 = n293 & ~n294 ;
  assign n296 = n282 & n295 ;
  assign n297 = n282 | n295 ;
  assign n298 = ~n296 & n297 ;
  assign n299 = n280 & n298 ;
  assign n300 = n280 | n298 ;
  assign n301 = ~n299 & n300 ;
  assign n302 = n296 | n299 ;
  assign n303 = n284 | n294 ;
  assign n304 = n287 | n290 ;
  assign n305 = x195 & n304 ;
  assign n306 = x195 | n304 ;
  assign n307 = ~n305 & n306 ;
  assign n308 = x3 & x67 ;
  assign n309 = x3 | x67 ;
  assign n310 = ~n308 & n309 ;
  assign n311 = x131 & n310 ;
  assign n312 = x131 | n310 ;
  assign n313 = ~n311 & n312 ;
  assign n314 = n307 | n313 ;
  assign n315 = n307 & n313 ;
  assign n316 = n314 & ~n315 ;
  assign n317 = n303 & n316 ;
  assign n318 = n303 | n316 ;
  assign n319 = ~n317 & n318 ;
  assign n320 = n302 & n319 ;
  assign n321 = n302 | n319 ;
  assign n322 = ~n320 & n321 ;
  assign n323 = n317 | n320 ;
  assign n324 = n305 | n315 ;
  assign n325 = n308 | n311 ;
  assign n326 = x196 & n325 ;
  assign n327 = x196 | n325 ;
  assign n328 = ~n326 & n327 ;
  assign n329 = x4 & x68 ;
  assign n330 = x4 | x68 ;
  assign n331 = ~n329 & n330 ;
  assign n332 = x132 & n331 ;
  assign n333 = x132 | n331 ;
  assign n334 = ~n332 & n333 ;
  assign n335 = n328 | n334 ;
  assign n336 = n328 & n334 ;
  assign n337 = n335 & ~n336 ;
  assign n338 = n324 & n337 ;
  assign n339 = n324 | n337 ;
  assign n340 = ~n338 & n339 ;
  assign n341 = n323 & n340 ;
  assign n342 = n323 | n340 ;
  assign n343 = ~n341 & n342 ;
  assign n344 = n338 | n341 ;
  assign n345 = n326 | n336 ;
  assign n346 = n329 | n332 ;
  assign n347 = x197 & n346 ;
  assign n348 = x197 | n346 ;
  assign n349 = ~n347 & n348 ;
  assign n350 = x5 & x69 ;
  assign n351 = x5 | x69 ;
  assign n352 = ~n350 & n351 ;
  assign n353 = x133 & n352 ;
  assign n354 = x133 | n352 ;
  assign n355 = ~n353 & n354 ;
  assign n356 = n349 | n355 ;
  assign n357 = n349 & n355 ;
  assign n358 = n356 & ~n357 ;
  assign n359 = n345 & n358 ;
  assign n360 = n345 | n358 ;
  assign n361 = ~n359 & n360 ;
  assign n362 = n344 & n361 ;
  assign n363 = n344 | n361 ;
  assign n364 = ~n362 & n363 ;
  assign n365 = n359 | n362 ;
  assign n366 = n347 | n357 ;
  assign n367 = n350 | n353 ;
  assign n368 = x198 & n367 ;
  assign n369 = x198 | n367 ;
  assign n370 = ~n368 & n369 ;
  assign n371 = x6 & x70 ;
  assign n372 = x6 | x70 ;
  assign n373 = ~n371 & n372 ;
  assign n374 = x134 & n373 ;
  assign n375 = x134 | n373 ;
  assign n376 = ~n374 & n375 ;
  assign n377 = n370 | n376 ;
  assign n378 = n370 & n376 ;
  assign n379 = n377 & ~n378 ;
  assign n380 = n366 & n379 ;
  assign n381 = n366 | n379 ;
  assign n382 = ~n380 & n381 ;
  assign n383 = n365 & n382 ;
  assign n384 = n365 | n382 ;
  assign n385 = ~n383 & n384 ;
  assign n386 = n380 | n383 ;
  assign n387 = n368 | n378 ;
  assign n388 = n371 | n374 ;
  assign n389 = x199 & n388 ;
  assign n390 = x199 | n388 ;
  assign n391 = ~n389 & n390 ;
  assign n392 = x7 & x71 ;
  assign n393 = x7 | x71 ;
  assign n394 = ~n392 & n393 ;
  assign n395 = x135 & n394 ;
  assign n396 = x135 | n394 ;
  assign n397 = ~n395 & n396 ;
  assign n398 = n391 | n397 ;
  assign n399 = n391 & n397 ;
  assign n400 = n398 & ~n399 ;
  assign n401 = n387 & n400 ;
  assign n402 = n387 | n400 ;
  assign n403 = ~n401 & n402 ;
  assign n404 = n386 & n403 ;
  assign n405 = n386 | n403 ;
  assign n406 = ~n404 & n405 ;
  assign n407 = n401 | n404 ;
  assign n408 = n389 | n399 ;
  assign n409 = n392 | n395 ;
  assign n410 = x200 & n409 ;
  assign n411 = x200 | n409 ;
  assign n412 = ~n410 & n411 ;
  assign n413 = x8 & x72 ;
  assign n414 = x8 | x72 ;
  assign n415 = ~n413 & n414 ;
  assign n416 = x136 & n415 ;
  assign n417 = x136 | n415 ;
  assign n418 = ~n416 & n417 ;
  assign n419 = n412 & n418 ;
  assign n420 = n412 | n418 ;
  assign n421 = ~n419 & n420 ;
  assign n422 = n408 & n421 ;
  assign n423 = n408 | n421 ;
  assign n424 = ~n422 & n423 ;
  assign n425 = n407 & n424 ;
  assign n426 = n407 | n424 ;
  assign n427 = ~n425 & n426 ;
  assign n428 = n422 | n425 ;
  assign n429 = n410 | n419 ;
  assign n430 = n413 | n416 ;
  assign n431 = x201 & n430 ;
  assign n432 = x201 | n430 ;
  assign n433 = ~n431 & n432 ;
  assign n434 = x9 & x73 ;
  assign n435 = x9 | x73 ;
  assign n436 = ~n434 & n435 ;
  assign n437 = x137 & n436 ;
  assign n438 = x137 | n436 ;
  assign n439 = ~n437 & n438 ;
  assign n440 = n433 | n439 ;
  assign n441 = n433 & n439 ;
  assign n442 = n440 & ~n441 ;
  assign n443 = n429 & n442 ;
  assign n444 = n429 | n442 ;
  assign n445 = ~n443 & n444 ;
  assign n446 = n428 & n445 ;
  assign n447 = n428 | n445 ;
  assign n448 = ~n446 & n447 ;
  assign n449 = n443 | n446 ;
  assign n450 = n431 | n441 ;
  assign n451 = n434 | n437 ;
  assign n452 = x202 & n451 ;
  assign n453 = x202 | n451 ;
  assign n454 = ~n452 & n453 ;
  assign n455 = x10 & x74 ;
  assign n456 = x10 | x74 ;
  assign n457 = ~n455 & n456 ;
  assign n458 = x138 & n457 ;
  assign n459 = x138 | n457 ;
  assign n460 = ~n458 & n459 ;
  assign n461 = n454 | n460 ;
  assign n462 = n454 & n460 ;
  assign n463 = n461 & ~n462 ;
  assign n464 = n450 & n463 ;
  assign n465 = n450 | n463 ;
  assign n466 = ~n464 & n465 ;
  assign n467 = n449 & n466 ;
  assign n468 = n449 | n466 ;
  assign n469 = ~n467 & n468 ;
  assign n470 = n464 | n467 ;
  assign n471 = n452 | n462 ;
  assign n472 = n455 | n458 ;
  assign n473 = x203 & n472 ;
  assign n474 = x203 | n472 ;
  assign n475 = ~n473 & n474 ;
  assign n476 = x11 & x75 ;
  assign n477 = x11 | x75 ;
  assign n478 = ~n476 & n477 ;
  assign n479 = x139 & n478 ;
  assign n480 = x139 | n478 ;
  assign n481 = ~n479 & n480 ;
  assign n482 = n475 | n481 ;
  assign n483 = n475 & n481 ;
  assign n484 = n482 & ~n483 ;
  assign n485 = n471 & n484 ;
  assign n486 = n471 | n484 ;
  assign n487 = ~n485 & n486 ;
  assign n488 = n470 & n487 ;
  assign n489 = n470 | n487 ;
  assign n490 = ~n488 & n489 ;
  assign n491 = n485 | n488 ;
  assign n492 = n473 | n483 ;
  assign n493 = n476 | n479 ;
  assign n494 = x204 & n493 ;
  assign n495 = x204 | n493 ;
  assign n496 = ~n494 & n495 ;
  assign n497 = x12 & x76 ;
  assign n498 = x12 | x76 ;
  assign n499 = ~n497 & n498 ;
  assign n500 = x140 & n499 ;
  assign n501 = x140 | n499 ;
  assign n502 = ~n500 & n501 ;
  assign n503 = n496 | n502 ;
  assign n504 = n496 & n502 ;
  assign n505 = n503 & ~n504 ;
  assign n506 = n492 & n505 ;
  assign n507 = n492 | n505 ;
  assign n508 = ~n506 & n507 ;
  assign n509 = n491 & n508 ;
  assign n510 = n491 | n508 ;
  assign n511 = ~n509 & n510 ;
  assign n512 = n506 | n509 ;
  assign n513 = n494 | n504 ;
  assign n514 = n497 | n500 ;
  assign n515 = x205 & n514 ;
  assign n516 = x205 | n514 ;
  assign n517 = ~n515 & n516 ;
  assign n518 = x13 & x77 ;
  assign n519 = x13 | x77 ;
  assign n520 = ~n518 & n519 ;
  assign n521 = x141 & n520 ;
  assign n522 = x141 | n520 ;
  assign n523 = ~n521 & n522 ;
  assign n524 = n517 | n523 ;
  assign n525 = n517 & n523 ;
  assign n526 = n524 & ~n525 ;
  assign n527 = n513 & n526 ;
  assign n528 = n513 | n526 ;
  assign n529 = ~n527 & n528 ;
  assign n530 = n512 & n529 ;
  assign n531 = n512 | n529 ;
  assign n532 = ~n530 & n531 ;
  assign n533 = n527 | n530 ;
  assign n534 = n515 | n525 ;
  assign n535 = n518 | n521 ;
  assign n536 = x206 & n535 ;
  assign n537 = x206 | n535 ;
  assign n538 = ~n536 & n537 ;
  assign n539 = x14 & x78 ;
  assign n540 = x14 | x78 ;
  assign n541 = ~n539 & n540 ;
  assign n542 = x142 & n541 ;
  assign n543 = x142 | n541 ;
  assign n544 = ~n542 & n543 ;
  assign n545 = n538 | n544 ;
  assign n546 = n538 & n544 ;
  assign n547 = n545 & ~n546 ;
  assign n548 = n534 & n547 ;
  assign n549 = n534 | n547 ;
  assign n550 = ~n548 & n549 ;
  assign n551 = n533 & n550 ;
  assign n552 = n533 | n550 ;
  assign n553 = ~n551 & n552 ;
  assign n554 = n548 | n551 ;
  assign n555 = n536 | n546 ;
  assign n556 = n539 | n542 ;
  assign n557 = x207 & n556 ;
  assign n558 = x207 | n556 ;
  assign n559 = ~n557 & n558 ;
  assign n560 = x15 & x79 ;
  assign n561 = x15 | x79 ;
  assign n562 = ~n560 & n561 ;
  assign n563 = x143 & n562 ;
  assign n564 = x143 | n562 ;
  assign n565 = ~n563 & n564 ;
  assign n566 = n559 | n565 ;
  assign n567 = n559 & n565 ;
  assign n568 = n566 & ~n567 ;
  assign n569 = n555 & n568 ;
  assign n570 = n555 | n568 ;
  assign n571 = ~n569 & n570 ;
  assign n572 = n554 & n571 ;
  assign n573 = n554 | n571 ;
  assign n574 = ~n572 & n573 ;
  assign n575 = n569 | n572 ;
  assign n576 = n557 | n567 ;
  assign n577 = n560 | n563 ;
  assign n578 = x208 & n577 ;
  assign n579 = x208 | n577 ;
  assign n580 = ~n578 & n579 ;
  assign n581 = x16 & x80 ;
  assign n582 = x16 | x80 ;
  assign n583 = ~n581 & n582 ;
  assign n584 = x144 & n583 ;
  assign n585 = x144 | n583 ;
  assign n586 = ~n584 & n585 ;
  assign n587 = n580 | n586 ;
  assign n588 = n580 & n586 ;
  assign n589 = n587 & ~n588 ;
  assign n590 = n576 & n589 ;
  assign n591 = n576 | n589 ;
  assign n592 = ~n590 & n591 ;
  assign n593 = n575 & n592 ;
  assign n594 = n575 | n592 ;
  assign n595 = ~n593 & n594 ;
  assign n596 = n590 | n593 ;
  assign n597 = n578 | n588 ;
  assign n598 = n581 | n584 ;
  assign n599 = x209 & n598 ;
  assign n600 = x209 | n598 ;
  assign n601 = ~n599 & n600 ;
  assign n602 = x17 & x81 ;
  assign n603 = x17 | x81 ;
  assign n604 = ~n602 & n603 ;
  assign n605 = x145 & n604 ;
  assign n606 = x145 | n604 ;
  assign n607 = ~n605 & n606 ;
  assign n608 = n601 | n607 ;
  assign n609 = n601 & n607 ;
  assign n610 = n608 & ~n609 ;
  assign n611 = n597 & n610 ;
  assign n612 = n597 | n610 ;
  assign n613 = ~n611 & n612 ;
  assign n614 = n596 & n613 ;
  assign n615 = n596 | n613 ;
  assign n616 = ~n614 & n615 ;
  assign n617 = n611 | n614 ;
  assign n618 = n599 | n609 ;
  assign n619 = n602 | n605 ;
  assign n620 = x210 & n619 ;
  assign n621 = x210 | n619 ;
  assign n622 = ~n620 & n621 ;
  assign n623 = x18 & x82 ;
  assign n624 = x18 | x82 ;
  assign n625 = ~n623 & n624 ;
  assign n626 = x146 & n625 ;
  assign n627 = x146 | n625 ;
  assign n628 = ~n626 & n627 ;
  assign n629 = n622 | n628 ;
  assign n630 = n622 & n628 ;
  assign n631 = n629 & ~n630 ;
  assign n632 = n618 & n631 ;
  assign n633 = n618 | n631 ;
  assign n634 = ~n632 & n633 ;
  assign n635 = n617 & n634 ;
  assign n636 = n617 | n634 ;
  assign n637 = ~n635 & n636 ;
  assign n638 = n632 | n635 ;
  assign n639 = n620 | n630 ;
  assign n640 = n623 | n626 ;
  assign n641 = x211 & n640 ;
  assign n642 = x211 | n640 ;
  assign n643 = ~n641 & n642 ;
  assign n644 = x19 & x83 ;
  assign n645 = x19 | x83 ;
  assign n646 = ~n644 & n645 ;
  assign n647 = x147 & n646 ;
  assign n648 = x147 | n646 ;
  assign n649 = ~n647 & n648 ;
  assign n650 = n643 | n649 ;
  assign n651 = n643 & n649 ;
  assign n652 = n650 & ~n651 ;
  assign n653 = n639 & n652 ;
  assign n654 = n639 | n652 ;
  assign n655 = ~n653 & n654 ;
  assign n656 = n638 & n655 ;
  assign n657 = n638 | n655 ;
  assign n658 = ~n656 & n657 ;
  assign n659 = n653 | n656 ;
  assign n660 = n641 | n651 ;
  assign n661 = n644 | n647 ;
  assign n662 = x212 & n661 ;
  assign n663 = x212 | n661 ;
  assign n664 = ~n662 & n663 ;
  assign n665 = x20 & x84 ;
  assign n666 = x20 | x84 ;
  assign n667 = ~n665 & n666 ;
  assign n668 = x148 & n667 ;
  assign n669 = x148 | n667 ;
  assign n670 = ~n668 & n669 ;
  assign n671 = n664 | n670 ;
  assign n672 = n664 & n670 ;
  assign n673 = n671 & ~n672 ;
  assign n674 = n660 & n673 ;
  assign n675 = n660 | n673 ;
  assign n676 = ~n674 & n675 ;
  assign n677 = n659 & n676 ;
  assign n678 = n659 | n676 ;
  assign n679 = ~n677 & n678 ;
  assign n680 = n674 | n677 ;
  assign n681 = n662 | n672 ;
  assign n682 = n665 | n668 ;
  assign n683 = x213 & n682 ;
  assign n684 = x213 | n682 ;
  assign n685 = ~n683 & n684 ;
  assign n686 = x21 & x85 ;
  assign n687 = x21 | x85 ;
  assign n688 = ~n686 & n687 ;
  assign n689 = x149 & n688 ;
  assign n690 = x149 | n688 ;
  assign n691 = ~n689 & n690 ;
  assign n692 = n685 | n691 ;
  assign n693 = n685 & n691 ;
  assign n694 = n692 & ~n693 ;
  assign n695 = n681 & n694 ;
  assign n696 = n681 | n694 ;
  assign n697 = ~n695 & n696 ;
  assign n698 = n680 & n697 ;
  assign n699 = n680 | n697 ;
  assign n700 = ~n698 & n699 ;
  assign n701 = n695 | n698 ;
  assign n702 = n683 | n693 ;
  assign n703 = n686 | n689 ;
  assign n704 = x214 & n703 ;
  assign n705 = x214 | n703 ;
  assign n706 = ~n704 & n705 ;
  assign n707 = x22 & x86 ;
  assign n708 = x22 | x86 ;
  assign n709 = ~n707 & n708 ;
  assign n710 = x150 & n709 ;
  assign n711 = x150 | n709 ;
  assign n712 = ~n710 & n711 ;
  assign n713 = n706 | n712 ;
  assign n714 = n706 & n712 ;
  assign n715 = n713 & ~n714 ;
  assign n716 = n702 & n715 ;
  assign n717 = n702 | n715 ;
  assign n718 = ~n716 & n717 ;
  assign n719 = n701 & n718 ;
  assign n720 = n701 | n718 ;
  assign n721 = ~n719 & n720 ;
  assign n722 = n716 | n719 ;
  assign n723 = n704 | n714 ;
  assign n724 = n707 | n710 ;
  assign n725 = x215 & n724 ;
  assign n726 = x215 | n724 ;
  assign n727 = ~n725 & n726 ;
  assign n728 = x23 & x87 ;
  assign n729 = x23 | x87 ;
  assign n730 = ~n728 & n729 ;
  assign n731 = x151 & n730 ;
  assign n732 = x151 | n730 ;
  assign n733 = ~n731 & n732 ;
  assign n734 = n727 | n733 ;
  assign n735 = n727 & n733 ;
  assign n736 = n734 & ~n735 ;
  assign n737 = n723 & n736 ;
  assign n738 = n723 | n736 ;
  assign n739 = ~n737 & n738 ;
  assign n740 = n722 & n739 ;
  assign n741 = n722 | n739 ;
  assign n742 = ~n740 & n741 ;
  assign n743 = n737 | n740 ;
  assign n744 = n725 | n735 ;
  assign n745 = n728 | n731 ;
  assign n746 = x216 & n745 ;
  assign n747 = x216 | n745 ;
  assign n748 = ~n746 & n747 ;
  assign n749 = x24 & x88 ;
  assign n750 = x24 | x88 ;
  assign n751 = ~n749 & n750 ;
  assign n752 = x152 & n751 ;
  assign n753 = x152 | n751 ;
  assign n754 = ~n752 & n753 ;
  assign n755 = n748 | n754 ;
  assign n756 = n748 & n754 ;
  assign n757 = n755 & ~n756 ;
  assign n758 = n744 & n757 ;
  assign n759 = n744 | n757 ;
  assign n760 = ~n758 & n759 ;
  assign n761 = n743 & n760 ;
  assign n762 = n743 | n760 ;
  assign n763 = ~n761 & n762 ;
  assign n764 = n758 | n761 ;
  assign n765 = n746 | n756 ;
  assign n766 = n749 | n752 ;
  assign n767 = x217 & n766 ;
  assign n768 = x217 | n766 ;
  assign n769 = ~n767 & n768 ;
  assign n770 = x25 & x89 ;
  assign n771 = x25 | x89 ;
  assign n772 = ~n770 & n771 ;
  assign n773 = x153 & n772 ;
  assign n774 = x153 | n772 ;
  assign n775 = ~n773 & n774 ;
  assign n776 = n769 | n775 ;
  assign n777 = n769 & n775 ;
  assign n778 = n776 & ~n777 ;
  assign n779 = n765 & n778 ;
  assign n780 = n765 | n778 ;
  assign n781 = ~n779 & n780 ;
  assign n782 = n764 & n781 ;
  assign n783 = n764 | n781 ;
  assign n784 = ~n782 & n783 ;
  assign n785 = n779 | n782 ;
  assign n786 = n767 | n777 ;
  assign n787 = n770 | n773 ;
  assign n788 = x218 & n787 ;
  assign n789 = x218 | n787 ;
  assign n790 = ~n788 & n789 ;
  assign n791 = x26 & x90 ;
  assign n792 = x26 | x90 ;
  assign n793 = ~n791 & n792 ;
  assign n794 = x154 & n793 ;
  assign n795 = x154 | n793 ;
  assign n796 = ~n794 & n795 ;
  assign n797 = n790 | n796 ;
  assign n798 = n790 & n796 ;
  assign n799 = n797 & ~n798 ;
  assign n800 = n786 & n799 ;
  assign n801 = n786 | n799 ;
  assign n802 = ~n800 & n801 ;
  assign n803 = n785 & n802 ;
  assign n804 = n785 | n802 ;
  assign n805 = ~n803 & n804 ;
  assign n806 = n800 | n803 ;
  assign n807 = n788 | n798 ;
  assign n808 = n791 | n794 ;
  assign n809 = x219 & n808 ;
  assign n810 = x219 | n808 ;
  assign n811 = ~n809 & n810 ;
  assign n812 = x27 & x91 ;
  assign n813 = x27 | x91 ;
  assign n814 = ~n812 & n813 ;
  assign n815 = x155 & n814 ;
  assign n816 = x155 | n814 ;
  assign n817 = ~n815 & n816 ;
  assign n818 = n811 | n817 ;
  assign n819 = n811 & n817 ;
  assign n820 = n818 & ~n819 ;
  assign n821 = n807 & n820 ;
  assign n822 = n807 | n820 ;
  assign n823 = ~n821 & n822 ;
  assign n824 = n806 & n823 ;
  assign n825 = n806 | n823 ;
  assign n826 = ~n824 & n825 ;
  assign n827 = n821 | n824 ;
  assign n828 = n809 | n819 ;
  assign n829 = n812 | n815 ;
  assign n830 = x220 & n829 ;
  assign n831 = x220 | n829 ;
  assign n832 = ~n830 & n831 ;
  assign n833 = x28 & x92 ;
  assign n834 = x28 | x92 ;
  assign n835 = ~n833 & n834 ;
  assign n836 = x156 & n835 ;
  assign n837 = x156 | n835 ;
  assign n838 = ~n836 & n837 ;
  assign n839 = n832 | n838 ;
  assign n840 = n832 & n838 ;
  assign n841 = n839 & ~n840 ;
  assign n842 = n828 & n841 ;
  assign n843 = n828 | n841 ;
  assign n844 = ~n842 & n843 ;
  assign n845 = n827 & n844 ;
  assign n846 = n827 | n844 ;
  assign n847 = ~n845 & n846 ;
  assign n848 = n842 | n845 ;
  assign n849 = n830 | n840 ;
  assign n850 = n833 | n836 ;
  assign n851 = x221 & n850 ;
  assign n852 = x221 | n850 ;
  assign n853 = ~n851 & n852 ;
  assign n854 = x29 & x93 ;
  assign n855 = x29 | x93 ;
  assign n856 = ~n854 & n855 ;
  assign n857 = x157 & n856 ;
  assign n858 = x157 | n856 ;
  assign n859 = ~n857 & n858 ;
  assign n860 = n853 | n859 ;
  assign n861 = n853 & n859 ;
  assign n862 = n860 & ~n861 ;
  assign n863 = n849 & n862 ;
  assign n864 = n849 | n862 ;
  assign n865 = ~n863 & n864 ;
  assign n866 = n848 & n865 ;
  assign n867 = n848 | n865 ;
  assign n868 = ~n866 & n867 ;
  assign n869 = n863 | n866 ;
  assign n870 = n851 | n861 ;
  assign n871 = n854 | n857 ;
  assign n872 = x222 & n871 ;
  assign n873 = x222 | n871 ;
  assign n874 = ~n872 & n873 ;
  assign n875 = x30 & x94 ;
  assign n876 = x30 | x94 ;
  assign n877 = ~n875 & n876 ;
  assign n878 = x158 & n877 ;
  assign n879 = x158 | n877 ;
  assign n880 = ~n878 & n879 ;
  assign n881 = n874 | n880 ;
  assign n882 = n874 & n880 ;
  assign n883 = n881 & ~n882 ;
  assign n884 = n870 & n883 ;
  assign n885 = n870 | n883 ;
  assign n886 = ~n884 & n885 ;
  assign n887 = n869 & n886 ;
  assign n888 = n869 | n886 ;
  assign n889 = ~n887 & n888 ;
  assign n890 = n884 | n887 ;
  assign n891 = n872 | n882 ;
  assign n892 = n875 | n878 ;
  assign n893 = x223 & n892 ;
  assign n894 = x223 | n892 ;
  assign n895 = ~n893 & n894 ;
  assign n896 = x31 & x95 ;
  assign n897 = x31 | x95 ;
  assign n898 = ~n896 & n897 ;
  assign n899 = x159 & n898 ;
  assign n900 = x159 | n898 ;
  assign n901 = ~n899 & n900 ;
  assign n902 = n895 | n901 ;
  assign n903 = n895 & n901 ;
  assign n904 = n902 & ~n903 ;
  assign n905 = n891 & n904 ;
  assign n906 = n891 | n904 ;
  assign n907 = ~n905 & n906 ;
  assign n908 = n890 & n907 ;
  assign n909 = n890 | n907 ;
  assign n910 = ~n908 & n909 ;
  assign n911 = n905 | n908 ;
  assign n912 = n893 | n903 ;
  assign n913 = n896 | n899 ;
  assign n914 = x224 & n913 ;
  assign n915 = x224 | n913 ;
  assign n916 = ~n914 & n915 ;
  assign n917 = x32 & x96 ;
  assign n918 = x32 | x96 ;
  assign n919 = ~n917 & n918 ;
  assign n920 = x160 & n919 ;
  assign n921 = x160 | n919 ;
  assign n922 = ~n920 & n921 ;
  assign n923 = n916 | n922 ;
  assign n924 = n916 & n922 ;
  assign n925 = n923 & ~n924 ;
  assign n926 = n912 & n925 ;
  assign n927 = n912 | n925 ;
  assign n928 = ~n926 & n927 ;
  assign n929 = n911 & n928 ;
  assign n930 = n911 | n928 ;
  assign n931 = ~n929 & n930 ;
  assign n932 = n926 | n929 ;
  assign n933 = n914 | n924 ;
  assign n934 = n917 | n920 ;
  assign n935 = x225 & n934 ;
  assign n936 = x225 | n934 ;
  assign n937 = ~n935 & n936 ;
  assign n938 = x33 & x97 ;
  assign n939 = x33 | x97 ;
  assign n940 = ~n938 & n939 ;
  assign n941 = x161 & n940 ;
  assign n942 = x161 | n940 ;
  assign n943 = ~n941 & n942 ;
  assign n944 = n937 | n943 ;
  assign n945 = n937 & n943 ;
  assign n946 = n944 & ~n945 ;
  assign n947 = n933 & n946 ;
  assign n948 = n933 | n946 ;
  assign n949 = ~n947 & n948 ;
  assign n950 = n932 & n949 ;
  assign n951 = n932 | n949 ;
  assign n952 = ~n950 & n951 ;
  assign n953 = n947 | n950 ;
  assign n954 = n935 | n945 ;
  assign n955 = n938 | n941 ;
  assign n956 = x226 & n955 ;
  assign n957 = x226 | n955 ;
  assign n958 = ~n956 & n957 ;
  assign n959 = x34 & x98 ;
  assign n960 = x34 | x98 ;
  assign n961 = ~n959 & n960 ;
  assign n962 = x162 & n961 ;
  assign n963 = x162 | n961 ;
  assign n964 = ~n962 & n963 ;
  assign n965 = n958 | n964 ;
  assign n966 = n958 & n964 ;
  assign n967 = n965 & ~n966 ;
  assign n968 = n954 & n967 ;
  assign n969 = n954 | n967 ;
  assign n970 = ~n968 & n969 ;
  assign n971 = n953 & n970 ;
  assign n972 = n953 | n970 ;
  assign n973 = ~n971 & n972 ;
  assign n974 = n968 | n971 ;
  assign n975 = n956 | n966 ;
  assign n976 = n959 | n962 ;
  assign n977 = x227 & n976 ;
  assign n978 = x227 | n976 ;
  assign n979 = ~n977 & n978 ;
  assign n980 = x35 & x99 ;
  assign n981 = x35 | x99 ;
  assign n982 = ~n980 & n981 ;
  assign n983 = x163 & n982 ;
  assign n984 = x163 | n982 ;
  assign n985 = ~n983 & n984 ;
  assign n986 = n979 | n985 ;
  assign n987 = n979 & n985 ;
  assign n988 = n986 & ~n987 ;
  assign n989 = n975 & n988 ;
  assign n990 = n975 | n988 ;
  assign n991 = ~n989 & n990 ;
  assign n992 = n974 & n991 ;
  assign n993 = n974 | n991 ;
  assign n994 = ~n992 & n993 ;
  assign n995 = n989 | n992 ;
  assign n996 = n977 | n987 ;
  assign n997 = n980 | n983 ;
  assign n998 = x228 & n997 ;
  assign n999 = x228 | n997 ;
  assign n1000 = ~n998 & n999 ;
  assign n1001 = x36 & x100 ;
  assign n1002 = x36 | x100 ;
  assign n1003 = ~n1001 & n1002 ;
  assign n1004 = x164 & n1003 ;
  assign n1005 = x164 | n1003 ;
  assign n1006 = ~n1004 & n1005 ;
  assign n1007 = n1000 | n1006 ;
  assign n1008 = n1000 & n1006 ;
  assign n1009 = n1007 & ~n1008 ;
  assign n1010 = n996 & n1009 ;
  assign n1011 = n996 | n1009 ;
  assign n1012 = ~n1010 & n1011 ;
  assign n1013 = n995 & n1012 ;
  assign n1014 = n995 | n1012 ;
  assign n1015 = ~n1013 & n1014 ;
  assign n1016 = n1010 | n1013 ;
  assign n1017 = n998 | n1008 ;
  assign n1018 = n1001 | n1004 ;
  assign n1019 = x229 & n1018 ;
  assign n1020 = x229 | n1018 ;
  assign n1021 = ~n1019 & n1020 ;
  assign n1022 = x37 & x101 ;
  assign n1023 = x37 | x101 ;
  assign n1024 = ~n1022 & n1023 ;
  assign n1025 = x165 & n1024 ;
  assign n1026 = x165 | n1024 ;
  assign n1027 = ~n1025 & n1026 ;
  assign n1028 = n1021 | n1027 ;
  assign n1029 = n1021 & n1027 ;
  assign n1030 = n1028 & ~n1029 ;
  assign n1031 = n1017 & n1030 ;
  assign n1032 = n1017 | n1030 ;
  assign n1033 = ~n1031 & n1032 ;
  assign n1034 = n1016 & n1033 ;
  assign n1035 = n1016 | n1033 ;
  assign n1036 = ~n1034 & n1035 ;
  assign n1037 = n1031 | n1034 ;
  assign n1038 = n1019 | n1029 ;
  assign n1039 = n1022 | n1025 ;
  assign n1040 = x230 & n1039 ;
  assign n1041 = x230 | n1039 ;
  assign n1042 = ~n1040 & n1041 ;
  assign n1043 = x38 & x102 ;
  assign n1044 = x38 | x102 ;
  assign n1045 = ~n1043 & n1044 ;
  assign n1046 = x166 & n1045 ;
  assign n1047 = x166 | n1045 ;
  assign n1048 = ~n1046 & n1047 ;
  assign n1049 = n1042 | n1048 ;
  assign n1050 = n1042 & n1048 ;
  assign n1051 = n1049 & ~n1050 ;
  assign n1052 = n1038 & n1051 ;
  assign n1053 = n1038 | n1051 ;
  assign n1054 = ~n1052 & n1053 ;
  assign n1055 = n1037 & n1054 ;
  assign n1056 = n1037 | n1054 ;
  assign n1057 = ~n1055 & n1056 ;
  assign n1058 = n1052 | n1055 ;
  assign n1059 = n1040 | n1050 ;
  assign n1060 = n1043 | n1046 ;
  assign n1061 = x231 & n1060 ;
  assign n1062 = x231 | n1060 ;
  assign n1063 = ~n1061 & n1062 ;
  assign n1064 = x39 & x103 ;
  assign n1065 = x39 | x103 ;
  assign n1066 = ~n1064 & n1065 ;
  assign n1067 = x167 & n1066 ;
  assign n1068 = x167 | n1066 ;
  assign n1069 = ~n1067 & n1068 ;
  assign n1070 = n1063 | n1069 ;
  assign n1071 = n1063 & n1069 ;
  assign n1072 = n1070 & ~n1071 ;
  assign n1073 = n1059 & n1072 ;
  assign n1074 = n1059 | n1072 ;
  assign n1075 = ~n1073 & n1074 ;
  assign n1076 = n1058 & n1075 ;
  assign n1077 = n1058 | n1075 ;
  assign n1078 = ~n1076 & n1077 ;
  assign n1079 = n1073 | n1076 ;
  assign n1080 = n1061 | n1071 ;
  assign n1081 = n1064 | n1067 ;
  assign n1082 = x232 & n1081 ;
  assign n1083 = x232 | n1081 ;
  assign n1084 = ~n1082 & n1083 ;
  assign n1085 = x40 & x104 ;
  assign n1086 = x40 | x104 ;
  assign n1087 = ~n1085 & n1086 ;
  assign n1088 = x168 & n1087 ;
  assign n1089 = x168 | n1087 ;
  assign n1090 = ~n1088 & n1089 ;
  assign n1091 = n1084 | n1090 ;
  assign n1092 = n1084 & n1090 ;
  assign n1093 = n1091 & ~n1092 ;
  assign n1094 = n1080 & n1093 ;
  assign n1095 = n1080 | n1093 ;
  assign n1096 = ~n1094 & n1095 ;
  assign n1097 = n1079 & n1096 ;
  assign n1098 = n1079 | n1096 ;
  assign n1099 = ~n1097 & n1098 ;
  assign n1100 = n1094 | n1097 ;
  assign n1101 = n1082 | n1092 ;
  assign n1102 = n1085 | n1088 ;
  assign n1103 = x233 & n1102 ;
  assign n1104 = x233 | n1102 ;
  assign n1105 = ~n1103 & n1104 ;
  assign n1106 = x41 & x105 ;
  assign n1107 = x41 | x105 ;
  assign n1108 = ~n1106 & n1107 ;
  assign n1109 = x169 & n1108 ;
  assign n1110 = x169 | n1108 ;
  assign n1111 = ~n1109 & n1110 ;
  assign n1112 = n1105 | n1111 ;
  assign n1113 = n1105 & n1111 ;
  assign n1114 = n1112 & ~n1113 ;
  assign n1115 = n1101 & n1114 ;
  assign n1116 = n1101 | n1114 ;
  assign n1117 = ~n1115 & n1116 ;
  assign n1118 = n1100 & n1117 ;
  assign n1119 = n1100 | n1117 ;
  assign n1120 = ~n1118 & n1119 ;
  assign n1121 = n1115 | n1118 ;
  assign n1122 = n1103 | n1113 ;
  assign n1123 = n1106 | n1109 ;
  assign n1124 = x234 & n1123 ;
  assign n1125 = x234 | n1123 ;
  assign n1126 = ~n1124 & n1125 ;
  assign n1127 = x42 & x106 ;
  assign n1128 = x42 | x106 ;
  assign n1129 = ~n1127 & n1128 ;
  assign n1130 = x170 & n1129 ;
  assign n1131 = x170 | n1129 ;
  assign n1132 = ~n1130 & n1131 ;
  assign n1133 = n1126 | n1132 ;
  assign n1134 = n1126 & n1132 ;
  assign n1135 = n1133 & ~n1134 ;
  assign n1136 = n1122 & n1135 ;
  assign n1137 = n1122 | n1135 ;
  assign n1138 = ~n1136 & n1137 ;
  assign n1139 = n1121 & n1138 ;
  assign n1140 = n1121 | n1138 ;
  assign n1141 = ~n1139 & n1140 ;
  assign n1142 = n1136 | n1139 ;
  assign n1143 = n1124 | n1134 ;
  assign n1144 = n1127 | n1130 ;
  assign n1145 = x235 & n1144 ;
  assign n1146 = x235 | n1144 ;
  assign n1147 = ~n1145 & n1146 ;
  assign n1148 = x43 & x107 ;
  assign n1149 = x43 | x107 ;
  assign n1150 = ~n1148 & n1149 ;
  assign n1151 = x171 & n1150 ;
  assign n1152 = x171 | n1150 ;
  assign n1153 = ~n1151 & n1152 ;
  assign n1154 = n1147 | n1153 ;
  assign n1155 = n1147 & n1153 ;
  assign n1156 = n1154 & ~n1155 ;
  assign n1157 = n1143 & n1156 ;
  assign n1158 = n1143 | n1156 ;
  assign n1159 = ~n1157 & n1158 ;
  assign n1160 = n1142 & n1159 ;
  assign n1161 = n1142 | n1159 ;
  assign n1162 = ~n1160 & n1161 ;
  assign n1163 = n1157 | n1160 ;
  assign n1164 = n1145 | n1155 ;
  assign n1165 = n1148 | n1151 ;
  assign n1166 = x236 & n1165 ;
  assign n1167 = x236 | n1165 ;
  assign n1168 = ~n1166 & n1167 ;
  assign n1169 = x44 & x108 ;
  assign n1170 = x44 | x108 ;
  assign n1171 = ~n1169 & n1170 ;
  assign n1172 = x172 & n1171 ;
  assign n1173 = x172 | n1171 ;
  assign n1174 = ~n1172 & n1173 ;
  assign n1175 = n1168 | n1174 ;
  assign n1176 = n1168 & n1174 ;
  assign n1177 = n1175 & ~n1176 ;
  assign n1178 = n1164 & n1177 ;
  assign n1179 = n1164 | n1177 ;
  assign n1180 = ~n1178 & n1179 ;
  assign n1181 = n1163 & n1180 ;
  assign n1182 = n1163 | n1180 ;
  assign n1183 = ~n1181 & n1182 ;
  assign n1184 = n1178 | n1181 ;
  assign n1185 = n1166 | n1176 ;
  assign n1186 = n1169 | n1172 ;
  assign n1187 = x237 & n1186 ;
  assign n1188 = x237 | n1186 ;
  assign n1189 = ~n1187 & n1188 ;
  assign n1190 = x45 & x109 ;
  assign n1191 = x45 | x109 ;
  assign n1192 = ~n1190 & n1191 ;
  assign n1193 = x173 & n1192 ;
  assign n1194 = x173 | n1192 ;
  assign n1195 = ~n1193 & n1194 ;
  assign n1196 = n1189 | n1195 ;
  assign n1197 = n1189 & n1195 ;
  assign n1198 = n1196 & ~n1197 ;
  assign n1199 = n1185 & n1198 ;
  assign n1200 = n1185 | n1198 ;
  assign n1201 = ~n1199 & n1200 ;
  assign n1202 = n1184 & n1201 ;
  assign n1203 = n1184 | n1201 ;
  assign n1204 = ~n1202 & n1203 ;
  assign n1205 = n1199 | n1202 ;
  assign n1206 = n1187 | n1197 ;
  assign n1207 = n1190 | n1193 ;
  assign n1208 = x238 & n1207 ;
  assign n1209 = x238 | n1207 ;
  assign n1210 = ~n1208 & n1209 ;
  assign n1211 = x46 & x110 ;
  assign n1212 = x46 | x110 ;
  assign n1213 = ~n1211 & n1212 ;
  assign n1214 = x174 & n1213 ;
  assign n1215 = x174 | n1213 ;
  assign n1216 = ~n1214 & n1215 ;
  assign n1217 = n1210 | n1216 ;
  assign n1218 = n1210 & n1216 ;
  assign n1219 = n1217 & ~n1218 ;
  assign n1220 = n1206 & n1219 ;
  assign n1221 = n1206 | n1219 ;
  assign n1222 = ~n1220 & n1221 ;
  assign n1223 = n1205 & n1222 ;
  assign n1224 = n1205 | n1222 ;
  assign n1225 = ~n1223 & n1224 ;
  assign n1226 = n1220 | n1223 ;
  assign n1227 = n1208 | n1218 ;
  assign n1228 = n1211 | n1214 ;
  assign n1229 = x239 & n1228 ;
  assign n1230 = x239 | n1228 ;
  assign n1231 = ~n1229 & n1230 ;
  assign n1232 = x47 & x111 ;
  assign n1233 = x47 | x111 ;
  assign n1234 = ~n1232 & n1233 ;
  assign n1235 = x175 & n1234 ;
  assign n1236 = x175 | n1234 ;
  assign n1237 = ~n1235 & n1236 ;
  assign n1238 = n1231 | n1237 ;
  assign n1239 = n1231 & n1237 ;
  assign n1240 = n1238 & ~n1239 ;
  assign n1241 = n1227 & n1240 ;
  assign n1242 = n1227 | n1240 ;
  assign n1243 = ~n1241 & n1242 ;
  assign n1244 = n1226 & n1243 ;
  assign n1245 = n1226 | n1243 ;
  assign n1246 = ~n1244 & n1245 ;
  assign n1247 = n1241 | n1244 ;
  assign n1248 = n1229 | n1239 ;
  assign n1249 = n1232 | n1235 ;
  assign n1250 = x240 & n1249 ;
  assign n1251 = x240 | n1249 ;
  assign n1252 = ~n1250 & n1251 ;
  assign n1253 = x48 & x112 ;
  assign n1254 = x48 | x112 ;
  assign n1255 = ~n1253 & n1254 ;
  assign n1256 = x176 & n1255 ;
  assign n1257 = x176 | n1255 ;
  assign n1258 = ~n1256 & n1257 ;
  assign n1259 = n1252 | n1258 ;
  assign n1260 = n1252 & n1258 ;
  assign n1261 = n1259 & ~n1260 ;
  assign n1262 = n1248 & n1261 ;
  assign n1263 = n1248 | n1261 ;
  assign n1264 = ~n1262 & n1263 ;
  assign n1265 = n1247 & n1264 ;
  assign n1266 = n1247 | n1264 ;
  assign n1267 = ~n1265 & n1266 ;
  assign n1268 = n1262 | n1265 ;
  assign n1269 = n1250 | n1260 ;
  assign n1270 = n1253 | n1256 ;
  assign n1271 = x241 & n1270 ;
  assign n1272 = x241 | n1270 ;
  assign n1273 = ~n1271 & n1272 ;
  assign n1274 = x49 & x113 ;
  assign n1275 = x49 | x113 ;
  assign n1276 = ~n1274 & n1275 ;
  assign n1277 = x177 & n1276 ;
  assign n1278 = x177 | n1276 ;
  assign n1279 = ~n1277 & n1278 ;
  assign n1280 = n1273 | n1279 ;
  assign n1281 = n1273 & n1279 ;
  assign n1282 = n1280 & ~n1281 ;
  assign n1283 = n1269 & n1282 ;
  assign n1284 = n1269 | n1282 ;
  assign n1285 = ~n1283 & n1284 ;
  assign n1286 = n1268 & n1285 ;
  assign n1287 = n1268 | n1285 ;
  assign n1288 = ~n1286 & n1287 ;
  assign n1289 = n1283 | n1286 ;
  assign n1290 = n1271 | n1281 ;
  assign n1291 = n1274 | n1277 ;
  assign n1292 = x242 & n1291 ;
  assign n1293 = x242 | n1291 ;
  assign n1294 = ~n1292 & n1293 ;
  assign n1295 = x50 & x114 ;
  assign n1296 = x50 | x114 ;
  assign n1297 = ~n1295 & n1296 ;
  assign n1298 = x178 & n1297 ;
  assign n1299 = x178 | n1297 ;
  assign n1300 = ~n1298 & n1299 ;
  assign n1301 = n1294 | n1300 ;
  assign n1302 = n1294 & n1300 ;
  assign n1303 = n1301 & ~n1302 ;
  assign n1304 = n1290 & n1303 ;
  assign n1305 = n1290 | n1303 ;
  assign n1306 = ~n1304 & n1305 ;
  assign n1307 = n1289 & n1306 ;
  assign n1308 = n1289 | n1306 ;
  assign n1309 = ~n1307 & n1308 ;
  assign n1310 = n1304 | n1307 ;
  assign n1311 = n1292 | n1302 ;
  assign n1312 = n1295 | n1298 ;
  assign n1313 = x243 & n1312 ;
  assign n1314 = x243 | n1312 ;
  assign n1315 = ~n1313 & n1314 ;
  assign n1316 = x51 & x115 ;
  assign n1317 = x51 | x115 ;
  assign n1318 = ~n1316 & n1317 ;
  assign n1319 = x179 & n1318 ;
  assign n1320 = x179 | n1318 ;
  assign n1321 = ~n1319 & n1320 ;
  assign n1322 = n1315 | n1321 ;
  assign n1323 = n1315 & n1321 ;
  assign n1324 = n1322 & ~n1323 ;
  assign n1325 = n1311 & n1324 ;
  assign n1326 = n1311 | n1324 ;
  assign n1327 = ~n1325 & n1326 ;
  assign n1328 = n1310 & n1327 ;
  assign n1329 = n1310 | n1327 ;
  assign n1330 = ~n1328 & n1329 ;
  assign n1331 = n1325 | n1328 ;
  assign n1332 = n1313 | n1323 ;
  assign n1333 = n1316 | n1319 ;
  assign n1334 = x244 & n1333 ;
  assign n1335 = x244 | n1333 ;
  assign n1336 = ~n1334 & n1335 ;
  assign n1337 = x52 & x116 ;
  assign n1338 = x52 | x116 ;
  assign n1339 = ~n1337 & n1338 ;
  assign n1340 = x180 & n1339 ;
  assign n1341 = x180 | n1339 ;
  assign n1342 = ~n1340 & n1341 ;
  assign n1343 = n1336 | n1342 ;
  assign n1344 = n1336 & n1342 ;
  assign n1345 = n1343 & ~n1344 ;
  assign n1346 = n1332 & n1345 ;
  assign n1347 = n1332 | n1345 ;
  assign n1348 = ~n1346 & n1347 ;
  assign n1349 = n1331 & n1348 ;
  assign n1350 = n1331 | n1348 ;
  assign n1351 = ~n1349 & n1350 ;
  assign n1352 = n1346 | n1349 ;
  assign n1353 = n1334 | n1344 ;
  assign n1354 = n1337 | n1340 ;
  assign n1355 = x245 & n1354 ;
  assign n1356 = x245 | n1354 ;
  assign n1357 = ~n1355 & n1356 ;
  assign n1358 = x53 & x117 ;
  assign n1359 = x53 | x117 ;
  assign n1360 = ~n1358 & n1359 ;
  assign n1361 = x181 & n1360 ;
  assign n1362 = x181 | n1360 ;
  assign n1363 = ~n1361 & n1362 ;
  assign n1364 = n1357 | n1363 ;
  assign n1365 = n1357 & n1363 ;
  assign n1366 = n1364 & ~n1365 ;
  assign n1367 = n1353 & n1366 ;
  assign n1368 = n1353 | n1366 ;
  assign n1369 = ~n1367 & n1368 ;
  assign n1370 = n1352 & n1369 ;
  assign n1371 = n1352 | n1369 ;
  assign n1372 = ~n1370 & n1371 ;
  assign n1373 = n1367 | n1370 ;
  assign n1374 = n1355 | n1365 ;
  assign n1375 = n1358 | n1361 ;
  assign n1376 = x246 & n1375 ;
  assign n1377 = x246 | n1375 ;
  assign n1378 = ~n1376 & n1377 ;
  assign n1379 = x54 & x118 ;
  assign n1380 = x54 | x118 ;
  assign n1381 = ~n1379 & n1380 ;
  assign n1382 = x182 & n1381 ;
  assign n1383 = x182 | n1381 ;
  assign n1384 = ~n1382 & n1383 ;
  assign n1385 = n1378 | n1384 ;
  assign n1386 = n1378 & n1384 ;
  assign n1387 = n1385 & ~n1386 ;
  assign n1388 = n1374 & n1387 ;
  assign n1389 = n1374 | n1387 ;
  assign n1390 = ~n1388 & n1389 ;
  assign n1391 = n1373 & n1390 ;
  assign n1392 = n1373 | n1390 ;
  assign n1393 = ~n1391 & n1392 ;
  assign n1394 = n1388 | n1391 ;
  assign n1395 = n1376 | n1386 ;
  assign n1396 = n1379 | n1382 ;
  assign n1397 = x247 & n1396 ;
  assign n1398 = x247 | n1396 ;
  assign n1399 = ~n1397 & n1398 ;
  assign n1400 = x55 & x119 ;
  assign n1401 = x55 | x119 ;
  assign n1402 = ~n1400 & n1401 ;
  assign n1403 = x183 & n1402 ;
  assign n1404 = x183 | n1402 ;
  assign n1405 = ~n1403 & n1404 ;
  assign n1406 = n1399 | n1405 ;
  assign n1407 = n1399 & n1405 ;
  assign n1408 = n1406 & ~n1407 ;
  assign n1409 = n1395 & n1408 ;
  assign n1410 = n1395 | n1408 ;
  assign n1411 = ~n1409 & n1410 ;
  assign n1412 = n1394 & n1411 ;
  assign n1413 = n1394 | n1411 ;
  assign n1414 = ~n1412 & n1413 ;
  assign n1415 = n1409 | n1412 ;
  assign n1416 = n1397 | n1407 ;
  assign n1417 = n1400 | n1403 ;
  assign n1418 = x248 & n1417 ;
  assign n1419 = x248 | n1417 ;
  assign n1420 = ~n1418 & n1419 ;
  assign n1421 = x56 & x120 ;
  assign n1422 = x56 | x120 ;
  assign n1423 = ~n1421 & n1422 ;
  assign n1424 = x184 & n1423 ;
  assign n1425 = x184 | n1423 ;
  assign n1426 = ~n1424 & n1425 ;
  assign n1427 = n1420 | n1426 ;
  assign n1428 = n1420 & n1426 ;
  assign n1429 = n1427 & ~n1428 ;
  assign n1430 = n1416 & n1429 ;
  assign n1431 = n1416 | n1429 ;
  assign n1432 = ~n1430 & n1431 ;
  assign n1433 = n1415 & n1432 ;
  assign n1434 = n1415 | n1432 ;
  assign n1435 = ~n1433 & n1434 ;
  assign n1436 = n1430 | n1433 ;
  assign n1437 = n1418 | n1428 ;
  assign n1438 = n1421 | n1424 ;
  assign n1439 = x249 & n1438 ;
  assign n1440 = x249 | n1438 ;
  assign n1441 = ~n1439 & n1440 ;
  assign n1442 = x57 & x121 ;
  assign n1443 = x57 | x121 ;
  assign n1444 = ~n1442 & n1443 ;
  assign n1445 = x185 & n1444 ;
  assign n1446 = x185 | n1444 ;
  assign n1447 = ~n1445 & n1446 ;
  assign n1448 = n1441 | n1447 ;
  assign n1449 = n1441 & n1447 ;
  assign n1450 = n1448 & ~n1449 ;
  assign n1451 = n1437 & n1450 ;
  assign n1452 = n1437 | n1450 ;
  assign n1453 = ~n1451 & n1452 ;
  assign n1454 = n1436 & n1453 ;
  assign n1455 = n1436 | n1453 ;
  assign n1456 = ~n1454 & n1455 ;
  assign n1457 = n1451 | n1454 ;
  assign n1458 = n1439 | n1449 ;
  assign n1459 = n1442 | n1445 ;
  assign n1460 = x250 & n1459 ;
  assign n1461 = x250 | n1459 ;
  assign n1462 = ~n1460 & n1461 ;
  assign n1463 = x58 & x122 ;
  assign n1464 = x58 | x122 ;
  assign n1465 = ~n1463 & n1464 ;
  assign n1466 = x186 & n1465 ;
  assign n1467 = x186 | n1465 ;
  assign n1468 = ~n1466 & n1467 ;
  assign n1469 = n1462 | n1468 ;
  assign n1470 = n1462 & n1468 ;
  assign n1471 = n1469 & ~n1470 ;
  assign n1472 = n1458 & n1471 ;
  assign n1473 = n1458 | n1471 ;
  assign n1474 = ~n1472 & n1473 ;
  assign n1475 = n1457 & n1474 ;
  assign n1476 = n1457 | n1474 ;
  assign n1477 = ~n1475 & n1476 ;
  assign n1478 = n1472 | n1475 ;
  assign n1479 = n1460 | n1470 ;
  assign n1480 = n1463 | n1466 ;
  assign n1481 = x251 & n1480 ;
  assign n1482 = x251 | n1480 ;
  assign n1483 = ~n1481 & n1482 ;
  assign n1484 = x59 & x123 ;
  assign n1485 = x59 | x123 ;
  assign n1486 = ~n1484 & n1485 ;
  assign n1487 = x187 & n1486 ;
  assign n1488 = x187 | n1486 ;
  assign n1489 = ~n1487 & n1488 ;
  assign n1490 = n1483 | n1489 ;
  assign n1491 = n1483 & n1489 ;
  assign n1492 = n1490 & ~n1491 ;
  assign n1493 = n1479 & n1492 ;
  assign n1494 = n1479 | n1492 ;
  assign n1495 = ~n1493 & n1494 ;
  assign n1496 = n1478 & n1495 ;
  assign n1497 = n1478 | n1495 ;
  assign n1498 = ~n1496 & n1497 ;
  assign n1499 = n1493 | n1496 ;
  assign n1500 = n1481 | n1491 ;
  assign n1501 = n1484 | n1487 ;
  assign n1502 = x252 & n1501 ;
  assign n1503 = x252 | n1501 ;
  assign n1504 = ~n1502 & n1503 ;
  assign n1505 = x60 & x124 ;
  assign n1506 = x60 | x124 ;
  assign n1507 = ~n1505 & n1506 ;
  assign n1508 = x188 & n1507 ;
  assign n1509 = x188 | n1507 ;
  assign n1510 = ~n1508 & n1509 ;
  assign n1511 = n1504 | n1510 ;
  assign n1512 = n1504 & n1510 ;
  assign n1513 = n1511 & ~n1512 ;
  assign n1514 = n1500 & n1513 ;
  assign n1515 = n1500 | n1513 ;
  assign n1516 = ~n1514 & n1515 ;
  assign n1517 = n1499 & n1516 ;
  assign n1518 = n1499 | n1516 ;
  assign n1519 = ~n1517 & n1518 ;
  assign n1520 = n1514 | n1517 ;
  assign n1521 = n1502 | n1512 ;
  assign n1522 = n1505 | n1508 ;
  assign n1523 = x253 & n1522 ;
  assign n1524 = x253 | n1522 ;
  assign n1525 = ~n1523 & n1524 ;
  assign n1526 = x61 & x125 ;
  assign n1527 = x61 | x125 ;
  assign n1528 = ~n1526 & n1527 ;
  assign n1529 = x189 & n1528 ;
  assign n1530 = x189 | n1528 ;
  assign n1531 = ~n1529 & n1530 ;
  assign n1532 = n1525 | n1531 ;
  assign n1533 = n1525 & n1531 ;
  assign n1534 = n1532 & ~n1533 ;
  assign n1535 = n1521 & n1534 ;
  assign n1536 = n1521 | n1534 ;
  assign n1537 = ~n1535 & n1536 ;
  assign n1538 = n1520 & n1537 ;
  assign n1539 = n1520 | n1537 ;
  assign n1540 = ~n1538 & n1539 ;
  assign n1541 = n1535 | n1538 ;
  assign n1542 = n1523 | n1533 ;
  assign n1543 = n1526 | n1529 ;
  assign n1544 = x254 & n1543 ;
  assign n1545 = x254 | n1543 ;
  assign n1546 = ~n1544 & n1545 ;
  assign n1547 = x62 & x126 ;
  assign n1548 = x62 | x126 ;
  assign n1549 = ~n1547 & n1548 ;
  assign n1550 = x190 & n1549 ;
  assign n1551 = x190 | n1549 ;
  assign n1552 = ~n1550 & n1551 ;
  assign n1553 = n1546 | n1552 ;
  assign n1554 = n1546 & n1552 ;
  assign n1555 = n1553 & ~n1554 ;
  assign n1556 = n1542 & n1555 ;
  assign n1557 = n1542 | n1555 ;
  assign n1558 = ~n1556 & n1557 ;
  assign n1559 = n1541 & n1558 ;
  assign n1560 = n1541 | n1558 ;
  assign n1561 = ~n1559 & n1560 ;
  assign n1562 = n1556 | n1559 ;
  assign n1563 = n1544 | n1554 ;
  assign n1564 = x63 | x127 ;
  assign n1565 = x63 & x127 ;
  assign n1566 = n1564 & ~n1565 ;
  assign n1567 = x191 & ~n1566 ;
  assign n1568 = ~x191 & n1566 ;
  assign n1569 = n1567 | n1568 ;
  assign n1570 = n1547 | n1550 ;
  assign n1571 = ~x255 & n1570 ;
  assign n1572 = x255 & ~n1570 ;
  assign n1573 = n1571 | n1572 ;
  assign n1574 = n1569 | n1573 ;
  assign n1575 = n1569 & n1573 ;
  assign n1576 = n1574 & ~n1575 ;
  assign n1577 = n1563 & n1576 ;
  assign n1578 = n1563 | n1576 ;
  assign n1579 = ~n1577 & n1578 ;
  assign n1580 = n1562 & n1579 ;
  assign n1581 = n1562 | n1579 ;
  assign n1582 = ~n1580 & n1581 ;
  assign n1583 = n1577 | n1580 ;
  assign n1584 = n1564 & ~n1568 ;
  assign n1585 = ~n1571 & n1574 ;
  assign n1586 = n1584 | n1585 ;
  assign n1587 = n1584 & n1585 ;
  assign n1588 = n1586 & ~n1587 ;
  assign n1589 = n1583 & n1588 ;
  assign n1590 = n1583 | n1588 ;
  assign n1591 = ~n1589 & n1590 ;
  assign n1592 = n1586 & ~n1589 ;
  assign y0 = n265 ;
  assign y1 = n281 ;
  assign y2 = n301 ;
  assign y3 = n322 ;
  assign y4 = n343 ;
  assign y5 = n364 ;
  assign y6 = n385 ;
  assign y7 = n406 ;
  assign y8 = n427 ;
  assign y9 = n448 ;
  assign y10 = n469 ;
  assign y11 = n490 ;
  assign y12 = n511 ;
  assign y13 = n532 ;
  assign y14 = n553 ;
  assign y15 = n574 ;
  assign y16 = n595 ;
  assign y17 = n616 ;
  assign y18 = n637 ;
  assign y19 = n658 ;
  assign y20 = n679 ;
  assign y21 = n700 ;
  assign y22 = n721 ;
  assign y23 = n742 ;
  assign y24 = n763 ;
  assign y25 = n784 ;
  assign y26 = n805 ;
  assign y27 = n826 ;
  assign y28 = n847 ;
  assign y29 = n868 ;
  assign y30 = n889 ;
  assign y31 = n910 ;
  assign y32 = n931 ;
  assign y33 = n952 ;
  assign y34 = n973 ;
  assign y35 = n994 ;
  assign y36 = n1015 ;
  assign y37 = n1036 ;
  assign y38 = n1057 ;
  assign y39 = n1078 ;
  assign y40 = n1099 ;
  assign y41 = n1120 ;
  assign y42 = n1141 ;
  assign y43 = n1162 ;
  assign y44 = n1183 ;
  assign y45 = n1204 ;
  assign y46 = n1225 ;
  assign y47 = n1246 ;
  assign y48 = n1267 ;
  assign y49 = n1288 ;
  assign y50 = n1309 ;
  assign y51 = n1330 ;
  assign y52 = n1351 ;
  assign y53 = n1372 ;
  assign y54 = n1393 ;
  assign y55 = n1414 ;
  assign y56 = n1435 ;
  assign y57 = n1456 ;
  assign y58 = n1477 ;
  assign y59 = n1498 ;
  assign y60 = n1519 ;
  assign y61 = n1540 ;
  assign y62 = n1561 ;
  assign y63 = n1582 ;
  assign y64 = n1591 ;
  assign y65 = n1592 ;
endmodule
