module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 ;
  wire n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 ;
  assign n129 = ~x125 & x127 ;
  assign n130 = x126 & x127 ;
  assign n131 = ( x125 & ~x126 ) | ( x125 & n130 ) | ( ~x126 & n130 ) ;
  assign n132 = ( x124 & n129 ) | ( x124 & n131 ) | ( n129 & n131 ) ;
  assign n133 = ( x124 & x126 ) | ( x124 & ~n130 ) | ( x126 & ~n130 ) ;
  assign n134 = ( x122 & ~n132 ) | ( x122 & n133 ) | ( ~n132 & n133 ) ;
  assign n135 = x121 & ~n134 ;
  assign n136 = ( x123 & n132 ) | ( x123 & ~n133 ) | ( n132 & ~n133 ) ;
  assign n137 = ( ~x123 & n129 ) | ( ~x123 & n131 ) | ( n129 & n131 ) ;
  assign n138 = ( x122 & n136 ) | ( x122 & n137 ) | ( n136 & n137 ) ;
  assign n139 = ( x121 & n135 ) | ( x121 & n138 ) | ( n135 & n138 ) ;
  assign n140 = ( ~x121 & n136 ) | ( ~x121 & n137 ) | ( n136 & n137 ) ;
  assign n141 = ~x119 & n140 ;
  assign n142 = ( ~x119 & n139 ) | ( ~x119 & n141 ) | ( n139 & n141 ) ;
  assign n143 = x118 & n142 ;
  assign n144 = x120 & n140 ;
  assign n145 = ( x120 & n139 ) | ( x120 & n144 ) | ( n139 & n144 ) ;
  assign n146 = x120 | n134 ;
  assign n147 = ( x120 & ~n138 ) | ( x120 & n146 ) | ( ~n138 & n146 ) ;
  assign n148 = ( x119 & n145 ) | ( x119 & ~n147 ) | ( n145 & ~n147 ) ;
  assign n149 = ( x118 & n143 ) | ( x118 & n148 ) | ( n143 & n148 ) ;
  assign n150 = ( x118 & ~n145 ) | ( x118 & n147 ) | ( ~n145 & n147 ) ;
  assign n151 = x116 | n150 ;
  assign n152 = ( x116 & ~n149 ) | ( x116 & n151 ) | ( ~n149 & n151 ) ;
  assign n153 = x115 & ~n152 ;
  assign n154 = x117 & ~n150 ;
  assign n155 = ( x117 & n149 ) | ( x117 & n154 ) | ( n149 & n154 ) ;
  assign n156 = ~x117 & n142 ;
  assign n157 = ( ~x117 & n148 ) | ( ~x117 & n156 ) | ( n148 & n156 ) ;
  assign n158 = ( x116 & n155 ) | ( x116 & n157 ) | ( n155 & n157 ) ;
  assign n159 = ( x115 & n153 ) | ( x115 & n158 ) | ( n153 & n158 ) ;
  assign n160 = ( ~x115 & n155 ) | ( ~x115 & n157 ) | ( n155 & n157 ) ;
  assign n161 = ~x113 & n160 ;
  assign n162 = ( ~x113 & n159 ) | ( ~x113 & n161 ) | ( n159 & n161 ) ;
  assign n163 = x112 & n162 ;
  assign n164 = x114 & n160 ;
  assign n165 = ( x114 & n159 ) | ( x114 & n164 ) | ( n159 & n164 ) ;
  assign n166 = x114 | n152 ;
  assign n167 = ( x114 & ~n158 ) | ( x114 & n166 ) | ( ~n158 & n166 ) ;
  assign n168 = ( x113 & n165 ) | ( x113 & ~n167 ) | ( n165 & ~n167 ) ;
  assign n169 = ( x112 & n163 ) | ( x112 & n168 ) | ( n163 & n168 ) ;
  assign n170 = ( x112 & ~n165 ) | ( x112 & n167 ) | ( ~n165 & n167 ) ;
  assign n171 = x110 | n170 ;
  assign n172 = ( x110 & ~n169 ) | ( x110 & n171 ) | ( ~n169 & n171 ) ;
  assign n173 = x109 & ~n172 ;
  assign n174 = x111 & ~n170 ;
  assign n175 = ( x111 & n169 ) | ( x111 & n174 ) | ( n169 & n174 ) ;
  assign n176 = ~x111 & n162 ;
  assign n177 = ( ~x111 & n168 ) | ( ~x111 & n176 ) | ( n168 & n176 ) ;
  assign n178 = ( x110 & n175 ) | ( x110 & n177 ) | ( n175 & n177 ) ;
  assign n179 = ( x109 & n173 ) | ( x109 & n178 ) | ( n173 & n178 ) ;
  assign n180 = ( ~x109 & n175 ) | ( ~x109 & n177 ) | ( n175 & n177 ) ;
  assign n181 = ~x107 & n180 ;
  assign n182 = ( ~x107 & n179 ) | ( ~x107 & n181 ) | ( n179 & n181 ) ;
  assign n183 = x106 & n182 ;
  assign n184 = x108 & n180 ;
  assign n185 = ( x108 & n179 ) | ( x108 & n184 ) | ( n179 & n184 ) ;
  assign n186 = x108 | n172 ;
  assign n187 = ( x108 & ~n178 ) | ( x108 & n186 ) | ( ~n178 & n186 ) ;
  assign n188 = ( x107 & n185 ) | ( x107 & ~n187 ) | ( n185 & ~n187 ) ;
  assign n189 = ( x106 & n183 ) | ( x106 & n188 ) | ( n183 & n188 ) ;
  assign n190 = ( x106 & ~n185 ) | ( x106 & n187 ) | ( ~n185 & n187 ) ;
  assign n191 = x104 | n190 ;
  assign n192 = ( x104 & ~n189 ) | ( x104 & n191 ) | ( ~n189 & n191 ) ;
  assign n193 = x103 & ~n192 ;
  assign n194 = x105 & ~n190 ;
  assign n195 = ( x105 & n189 ) | ( x105 & n194 ) | ( n189 & n194 ) ;
  assign n196 = ~x105 & n182 ;
  assign n197 = ( ~x105 & n188 ) | ( ~x105 & n196 ) | ( n188 & n196 ) ;
  assign n198 = ( x104 & n195 ) | ( x104 & n197 ) | ( n195 & n197 ) ;
  assign n199 = ( x103 & n193 ) | ( x103 & n198 ) | ( n193 & n198 ) ;
  assign n200 = ( ~x103 & n195 ) | ( ~x103 & n197 ) | ( n195 & n197 ) ;
  assign n201 = ~x101 & n200 ;
  assign n202 = ( ~x101 & n199 ) | ( ~x101 & n201 ) | ( n199 & n201 ) ;
  assign n203 = x100 & n202 ;
  assign n204 = x102 & n200 ;
  assign n205 = ( x102 & n199 ) | ( x102 & n204 ) | ( n199 & n204 ) ;
  assign n206 = x102 | n192 ;
  assign n207 = ( x102 & ~n198 ) | ( x102 & n206 ) | ( ~n198 & n206 ) ;
  assign n208 = ( x101 & n205 ) | ( x101 & ~n207 ) | ( n205 & ~n207 ) ;
  assign n209 = ( x100 & n203 ) | ( x100 & n208 ) | ( n203 & n208 ) ;
  assign n210 = ( x100 & ~n205 ) | ( x100 & n207 ) | ( ~n205 & n207 ) ;
  assign n211 = x98 | n210 ;
  assign n212 = ( x98 & ~n209 ) | ( x98 & n211 ) | ( ~n209 & n211 ) ;
  assign n213 = x97 & ~n212 ;
  assign n214 = x99 & ~n210 ;
  assign n215 = ( x99 & n209 ) | ( x99 & n214 ) | ( n209 & n214 ) ;
  assign n216 = ~x99 & n202 ;
  assign n217 = ( ~x99 & n208 ) | ( ~x99 & n216 ) | ( n208 & n216 ) ;
  assign n218 = ( x98 & n215 ) | ( x98 & n217 ) | ( n215 & n217 ) ;
  assign n219 = ( x97 & n213 ) | ( x97 & n218 ) | ( n213 & n218 ) ;
  assign n220 = ( ~x97 & n215 ) | ( ~x97 & n217 ) | ( n215 & n217 ) ;
  assign n221 = ~x95 & n220 ;
  assign n222 = ( ~x95 & n219 ) | ( ~x95 & n221 ) | ( n219 & n221 ) ;
  assign n223 = x94 & n222 ;
  assign n224 = x96 & n220 ;
  assign n225 = ( x96 & n219 ) | ( x96 & n224 ) | ( n219 & n224 ) ;
  assign n226 = x96 | n212 ;
  assign n227 = ( x96 & ~n218 ) | ( x96 & n226 ) | ( ~n218 & n226 ) ;
  assign n228 = ( x95 & n225 ) | ( x95 & ~n227 ) | ( n225 & ~n227 ) ;
  assign n229 = ( x94 & n223 ) | ( x94 & n228 ) | ( n223 & n228 ) ;
  assign n230 = ( x94 & ~n225 ) | ( x94 & n227 ) | ( ~n225 & n227 ) ;
  assign n231 = x92 | n230 ;
  assign n232 = ( x92 & ~n229 ) | ( x92 & n231 ) | ( ~n229 & n231 ) ;
  assign n233 = x91 & ~n232 ;
  assign n234 = x93 & ~n230 ;
  assign n235 = ( x93 & n229 ) | ( x93 & n234 ) | ( n229 & n234 ) ;
  assign n236 = ~x93 & n222 ;
  assign n237 = ( ~x93 & n228 ) | ( ~x93 & n236 ) | ( n228 & n236 ) ;
  assign n238 = ( x92 & n235 ) | ( x92 & n237 ) | ( n235 & n237 ) ;
  assign n239 = ( x91 & n233 ) | ( x91 & n238 ) | ( n233 & n238 ) ;
  assign n240 = ( ~x91 & n235 ) | ( ~x91 & n237 ) | ( n235 & n237 ) ;
  assign n241 = ~x89 & n240 ;
  assign n242 = ( ~x89 & n239 ) | ( ~x89 & n241 ) | ( n239 & n241 ) ;
  assign n243 = x88 & n242 ;
  assign n244 = x90 & n240 ;
  assign n245 = ( x90 & n239 ) | ( x90 & n244 ) | ( n239 & n244 ) ;
  assign n246 = x90 | n232 ;
  assign n247 = ( x90 & ~n238 ) | ( x90 & n246 ) | ( ~n238 & n246 ) ;
  assign n248 = ( x89 & n245 ) | ( x89 & ~n247 ) | ( n245 & ~n247 ) ;
  assign n249 = ( x88 & n243 ) | ( x88 & n248 ) | ( n243 & n248 ) ;
  assign n250 = ( x88 & ~n245 ) | ( x88 & n247 ) | ( ~n245 & n247 ) ;
  assign n251 = x86 | n250 ;
  assign n252 = ( x86 & ~n249 ) | ( x86 & n251 ) | ( ~n249 & n251 ) ;
  assign n253 = x85 & ~n252 ;
  assign n254 = x87 & ~n250 ;
  assign n255 = ( x87 & n249 ) | ( x87 & n254 ) | ( n249 & n254 ) ;
  assign n256 = ~x87 & n242 ;
  assign n257 = ( ~x87 & n248 ) | ( ~x87 & n256 ) | ( n248 & n256 ) ;
  assign n258 = ( x86 & n255 ) | ( x86 & n257 ) | ( n255 & n257 ) ;
  assign n259 = ( x85 & n253 ) | ( x85 & n258 ) | ( n253 & n258 ) ;
  assign n260 = ( ~x85 & n255 ) | ( ~x85 & n257 ) | ( n255 & n257 ) ;
  assign n261 = ~x83 & n260 ;
  assign n262 = ( ~x83 & n259 ) | ( ~x83 & n261 ) | ( n259 & n261 ) ;
  assign n263 = x82 & n262 ;
  assign n264 = x84 & n260 ;
  assign n265 = ( x84 & n259 ) | ( x84 & n264 ) | ( n259 & n264 ) ;
  assign n266 = x84 | n252 ;
  assign n267 = ( x84 & ~n258 ) | ( x84 & n266 ) | ( ~n258 & n266 ) ;
  assign n268 = ( x83 & n265 ) | ( x83 & ~n267 ) | ( n265 & ~n267 ) ;
  assign n269 = ( x82 & n263 ) | ( x82 & n268 ) | ( n263 & n268 ) ;
  assign n270 = ( x82 & ~n265 ) | ( x82 & n267 ) | ( ~n265 & n267 ) ;
  assign n271 = x80 | n270 ;
  assign n272 = ( x80 & ~n269 ) | ( x80 & n271 ) | ( ~n269 & n271 ) ;
  assign n273 = x79 & ~n272 ;
  assign n274 = x81 & ~n270 ;
  assign n275 = ( x81 & n269 ) | ( x81 & n274 ) | ( n269 & n274 ) ;
  assign n276 = ~x81 & n262 ;
  assign n277 = ( ~x81 & n268 ) | ( ~x81 & n276 ) | ( n268 & n276 ) ;
  assign n278 = ( x80 & n275 ) | ( x80 & n277 ) | ( n275 & n277 ) ;
  assign n279 = ( x79 & n273 ) | ( x79 & n278 ) | ( n273 & n278 ) ;
  assign n280 = ( ~x79 & n275 ) | ( ~x79 & n277 ) | ( n275 & n277 ) ;
  assign n281 = ~x77 & n280 ;
  assign n282 = ( ~x77 & n279 ) | ( ~x77 & n281 ) | ( n279 & n281 ) ;
  assign n283 = x76 & n282 ;
  assign n284 = x78 & n280 ;
  assign n285 = ( x78 & n279 ) | ( x78 & n284 ) | ( n279 & n284 ) ;
  assign n286 = x78 | n272 ;
  assign n287 = ( x78 & ~n278 ) | ( x78 & n286 ) | ( ~n278 & n286 ) ;
  assign n288 = ( x77 & n285 ) | ( x77 & ~n287 ) | ( n285 & ~n287 ) ;
  assign n289 = ( x76 & n283 ) | ( x76 & n288 ) | ( n283 & n288 ) ;
  assign n290 = ( x76 & ~n285 ) | ( x76 & n287 ) | ( ~n285 & n287 ) ;
  assign n291 = x74 | n290 ;
  assign n292 = ( x74 & ~n289 ) | ( x74 & n291 ) | ( ~n289 & n291 ) ;
  assign n293 = x73 & ~n292 ;
  assign n294 = x75 & ~n290 ;
  assign n295 = ( x75 & n289 ) | ( x75 & n294 ) | ( n289 & n294 ) ;
  assign n296 = ~x75 & n282 ;
  assign n297 = ( ~x75 & n288 ) | ( ~x75 & n296 ) | ( n288 & n296 ) ;
  assign n298 = ( x74 & n295 ) | ( x74 & n297 ) | ( n295 & n297 ) ;
  assign n299 = ( x73 & n293 ) | ( x73 & n298 ) | ( n293 & n298 ) ;
  assign n300 = ( ~x73 & n295 ) | ( ~x73 & n297 ) | ( n295 & n297 ) ;
  assign n301 = ~x71 & n300 ;
  assign n302 = ( ~x71 & n299 ) | ( ~x71 & n301 ) | ( n299 & n301 ) ;
  assign n303 = x70 & n302 ;
  assign n304 = x72 & n300 ;
  assign n305 = ( x72 & n299 ) | ( x72 & n304 ) | ( n299 & n304 ) ;
  assign n306 = x72 | n292 ;
  assign n307 = ( x72 & ~n298 ) | ( x72 & n306 ) | ( ~n298 & n306 ) ;
  assign n308 = ( x71 & n305 ) | ( x71 & ~n307 ) | ( n305 & ~n307 ) ;
  assign n309 = ( x70 & n303 ) | ( x70 & n308 ) | ( n303 & n308 ) ;
  assign n310 = ( x70 & ~n305 ) | ( x70 & n307 ) | ( ~n305 & n307 ) ;
  assign n311 = x68 | n310 ;
  assign n312 = ( x68 & ~n309 ) | ( x68 & n311 ) | ( ~n309 & n311 ) ;
  assign n313 = x67 & ~n312 ;
  assign n314 = x69 & ~n310 ;
  assign n315 = ( x69 & n309 ) | ( x69 & n314 ) | ( n309 & n314 ) ;
  assign n316 = ~x69 & n302 ;
  assign n317 = ( ~x69 & n308 ) | ( ~x69 & n316 ) | ( n308 & n316 ) ;
  assign n318 = ( x68 & n315 ) | ( x68 & n317 ) | ( n315 & n317 ) ;
  assign n319 = ( x67 & n313 ) | ( x67 & n318 ) | ( n313 & n318 ) ;
  assign n320 = ( ~x67 & n315 ) | ( ~x67 & n317 ) | ( n315 & n317 ) ;
  assign n321 = ~x65 & n320 ;
  assign n322 = ( ~x65 & n319 ) | ( ~x65 & n321 ) | ( n319 & n321 ) ;
  assign n323 = x64 & n322 ;
  assign n324 = x66 & n320 ;
  assign n325 = ( x66 & n319 ) | ( x66 & n324 ) | ( n319 & n324 ) ;
  assign n326 = x66 | n312 ;
  assign n327 = ( x66 & ~n318 ) | ( x66 & n326 ) | ( ~n318 & n326 ) ;
  assign n328 = ( x65 & n325 ) | ( x65 & ~n327 ) | ( n325 & ~n327 ) ;
  assign n329 = ( x64 & n323 ) | ( x64 & n328 ) | ( n323 & n328 ) ;
  assign n330 = ( x64 & ~n325 ) | ( x64 & n327 ) | ( ~n325 & n327 ) ;
  assign n331 = x62 | n330 ;
  assign n332 = ( x62 & ~n329 ) | ( x62 & n331 ) | ( ~n329 & n331 ) ;
  assign n333 = x61 & ~n332 ;
  assign n334 = x63 & ~n330 ;
  assign n335 = ( x63 & n329 ) | ( x63 & n334 ) | ( n329 & n334 ) ;
  assign n336 = ~x63 & n322 ;
  assign n337 = ( ~x63 & n328 ) | ( ~x63 & n336 ) | ( n328 & n336 ) ;
  assign n338 = ( x62 & n335 ) | ( x62 & n337 ) | ( n335 & n337 ) ;
  assign n339 = ( x61 & n333 ) | ( x61 & n338 ) | ( n333 & n338 ) ;
  assign n340 = ( ~x61 & n335 ) | ( ~x61 & n337 ) | ( n335 & n337 ) ;
  assign n341 = ~x59 & n340 ;
  assign n342 = ( ~x59 & n339 ) | ( ~x59 & n341 ) | ( n339 & n341 ) ;
  assign n343 = x58 & n342 ;
  assign n344 = x60 & n340 ;
  assign n345 = ( x60 & n339 ) | ( x60 & n344 ) | ( n339 & n344 ) ;
  assign n346 = x60 | n332 ;
  assign n347 = ( x60 & ~n338 ) | ( x60 & n346 ) | ( ~n338 & n346 ) ;
  assign n348 = ( x59 & n345 ) | ( x59 & ~n347 ) | ( n345 & ~n347 ) ;
  assign n349 = ( x58 & n343 ) | ( x58 & n348 ) | ( n343 & n348 ) ;
  assign n350 = ( x58 & ~n345 ) | ( x58 & n347 ) | ( ~n345 & n347 ) ;
  assign n351 = x56 | n350 ;
  assign n352 = ( x56 & ~n349 ) | ( x56 & n351 ) | ( ~n349 & n351 ) ;
  assign n353 = x55 & ~n352 ;
  assign n354 = x57 & ~n350 ;
  assign n355 = ( x57 & n349 ) | ( x57 & n354 ) | ( n349 & n354 ) ;
  assign n356 = ~x57 & n342 ;
  assign n357 = ( ~x57 & n348 ) | ( ~x57 & n356 ) | ( n348 & n356 ) ;
  assign n358 = ( x56 & n355 ) | ( x56 & n357 ) | ( n355 & n357 ) ;
  assign n359 = ( x55 & n353 ) | ( x55 & n358 ) | ( n353 & n358 ) ;
  assign n360 = ( ~x55 & n355 ) | ( ~x55 & n357 ) | ( n355 & n357 ) ;
  assign n361 = ~x53 & n360 ;
  assign n362 = ( ~x53 & n359 ) | ( ~x53 & n361 ) | ( n359 & n361 ) ;
  assign n363 = x52 & n362 ;
  assign n364 = x54 & n360 ;
  assign n365 = ( x54 & n359 ) | ( x54 & n364 ) | ( n359 & n364 ) ;
  assign n366 = x54 | n352 ;
  assign n367 = ( x54 & ~n358 ) | ( x54 & n366 ) | ( ~n358 & n366 ) ;
  assign n368 = ( x53 & n365 ) | ( x53 & ~n367 ) | ( n365 & ~n367 ) ;
  assign n369 = ( x52 & n363 ) | ( x52 & n368 ) | ( n363 & n368 ) ;
  assign n370 = ( x52 & ~n365 ) | ( x52 & n367 ) | ( ~n365 & n367 ) ;
  assign n371 = x50 | n370 ;
  assign n372 = ( x50 & ~n369 ) | ( x50 & n371 ) | ( ~n369 & n371 ) ;
  assign n373 = x49 & ~n372 ;
  assign n374 = x51 & ~n370 ;
  assign n375 = ( x51 & n369 ) | ( x51 & n374 ) | ( n369 & n374 ) ;
  assign n376 = ~x51 & n362 ;
  assign n377 = ( ~x51 & n368 ) | ( ~x51 & n376 ) | ( n368 & n376 ) ;
  assign n378 = ( x50 & n375 ) | ( x50 & n377 ) | ( n375 & n377 ) ;
  assign n379 = ( x49 & n373 ) | ( x49 & n378 ) | ( n373 & n378 ) ;
  assign n380 = ( ~x49 & n375 ) | ( ~x49 & n377 ) | ( n375 & n377 ) ;
  assign n381 = ~x47 & n380 ;
  assign n382 = ( ~x47 & n379 ) | ( ~x47 & n381 ) | ( n379 & n381 ) ;
  assign n383 = x46 & n382 ;
  assign n384 = x48 & n380 ;
  assign n385 = ( x48 & n379 ) | ( x48 & n384 ) | ( n379 & n384 ) ;
  assign n386 = x48 | n372 ;
  assign n387 = ( x48 & ~n378 ) | ( x48 & n386 ) | ( ~n378 & n386 ) ;
  assign n388 = ( x47 & n385 ) | ( x47 & ~n387 ) | ( n385 & ~n387 ) ;
  assign n389 = ( x46 & n383 ) | ( x46 & n388 ) | ( n383 & n388 ) ;
  assign n390 = ( x46 & ~n385 ) | ( x46 & n387 ) | ( ~n385 & n387 ) ;
  assign n391 = x44 | n390 ;
  assign n392 = ( x44 & ~n389 ) | ( x44 & n391 ) | ( ~n389 & n391 ) ;
  assign n393 = x43 & ~n392 ;
  assign n394 = x45 & ~n390 ;
  assign n395 = ( x45 & n389 ) | ( x45 & n394 ) | ( n389 & n394 ) ;
  assign n396 = ~x45 & n382 ;
  assign n397 = ( ~x45 & n388 ) | ( ~x45 & n396 ) | ( n388 & n396 ) ;
  assign n398 = ( x44 & n395 ) | ( x44 & n397 ) | ( n395 & n397 ) ;
  assign n399 = ( x43 & n393 ) | ( x43 & n398 ) | ( n393 & n398 ) ;
  assign n400 = ( ~x43 & n395 ) | ( ~x43 & n397 ) | ( n395 & n397 ) ;
  assign n401 = ~x41 & n400 ;
  assign n402 = ( ~x41 & n399 ) | ( ~x41 & n401 ) | ( n399 & n401 ) ;
  assign n403 = x40 & n402 ;
  assign n404 = x42 & n400 ;
  assign n405 = ( x42 & n399 ) | ( x42 & n404 ) | ( n399 & n404 ) ;
  assign n406 = x42 | n392 ;
  assign n407 = ( x42 & ~n398 ) | ( x42 & n406 ) | ( ~n398 & n406 ) ;
  assign n408 = ( x41 & n405 ) | ( x41 & ~n407 ) | ( n405 & ~n407 ) ;
  assign n409 = ( x40 & n403 ) | ( x40 & n408 ) | ( n403 & n408 ) ;
  assign n410 = ( x40 & ~n405 ) | ( x40 & n407 ) | ( ~n405 & n407 ) ;
  assign n411 = x38 | n410 ;
  assign n412 = ( x38 & ~n409 ) | ( x38 & n411 ) | ( ~n409 & n411 ) ;
  assign n413 = x37 & ~n412 ;
  assign n414 = x39 & ~n410 ;
  assign n415 = ( x39 & n409 ) | ( x39 & n414 ) | ( n409 & n414 ) ;
  assign n416 = ~x39 & n402 ;
  assign n417 = ( ~x39 & n408 ) | ( ~x39 & n416 ) | ( n408 & n416 ) ;
  assign n418 = ( x38 & n415 ) | ( x38 & n417 ) | ( n415 & n417 ) ;
  assign n419 = ( x37 & n413 ) | ( x37 & n418 ) | ( n413 & n418 ) ;
  assign n420 = ( ~x37 & n415 ) | ( ~x37 & n417 ) | ( n415 & n417 ) ;
  assign n421 = ~x35 & n420 ;
  assign n422 = ( ~x35 & n419 ) | ( ~x35 & n421 ) | ( n419 & n421 ) ;
  assign n423 = x34 & n422 ;
  assign n424 = x36 & n420 ;
  assign n425 = ( x36 & n419 ) | ( x36 & n424 ) | ( n419 & n424 ) ;
  assign n426 = x36 | n412 ;
  assign n427 = ( x36 & ~n418 ) | ( x36 & n426 ) | ( ~n418 & n426 ) ;
  assign n428 = ( x35 & n425 ) | ( x35 & ~n427 ) | ( n425 & ~n427 ) ;
  assign n429 = ( x34 & n423 ) | ( x34 & n428 ) | ( n423 & n428 ) ;
  assign n430 = ( x34 & ~n425 ) | ( x34 & n427 ) | ( ~n425 & n427 ) ;
  assign n431 = x32 | n430 ;
  assign n432 = ( x32 & ~n429 ) | ( x32 & n431 ) | ( ~n429 & n431 ) ;
  assign n433 = x31 & ~n432 ;
  assign n434 = x33 & ~n430 ;
  assign n435 = ( x33 & n429 ) | ( x33 & n434 ) | ( n429 & n434 ) ;
  assign n436 = ~x33 & n422 ;
  assign n437 = ( ~x33 & n428 ) | ( ~x33 & n436 ) | ( n428 & n436 ) ;
  assign n438 = ( x32 & n435 ) | ( x32 & n437 ) | ( n435 & n437 ) ;
  assign n439 = ( x31 & n433 ) | ( x31 & n438 ) | ( n433 & n438 ) ;
  assign n440 = ( ~x31 & n435 ) | ( ~x31 & n437 ) | ( n435 & n437 ) ;
  assign n441 = ~x29 & n440 ;
  assign n442 = ( ~x29 & n439 ) | ( ~x29 & n441 ) | ( n439 & n441 ) ;
  assign n443 = x28 & n442 ;
  assign n444 = x30 & n440 ;
  assign n445 = ( x30 & n439 ) | ( x30 & n444 ) | ( n439 & n444 ) ;
  assign n446 = x30 | n432 ;
  assign n447 = ( x30 & ~n438 ) | ( x30 & n446 ) | ( ~n438 & n446 ) ;
  assign n448 = ( x29 & n445 ) | ( x29 & ~n447 ) | ( n445 & ~n447 ) ;
  assign n449 = ( x28 & n443 ) | ( x28 & n448 ) | ( n443 & n448 ) ;
  assign n450 = ( x28 & ~n445 ) | ( x28 & n447 ) | ( ~n445 & n447 ) ;
  assign n451 = x26 | n450 ;
  assign n452 = ( x26 & ~n449 ) | ( x26 & n451 ) | ( ~n449 & n451 ) ;
  assign n453 = x25 & ~n452 ;
  assign n454 = x27 & ~n450 ;
  assign n455 = ( x27 & n449 ) | ( x27 & n454 ) | ( n449 & n454 ) ;
  assign n456 = ~x27 & n442 ;
  assign n457 = ( ~x27 & n448 ) | ( ~x27 & n456 ) | ( n448 & n456 ) ;
  assign n458 = ( x26 & n455 ) | ( x26 & n457 ) | ( n455 & n457 ) ;
  assign n459 = ( x25 & n453 ) | ( x25 & n458 ) | ( n453 & n458 ) ;
  assign n460 = ( ~x25 & n455 ) | ( ~x25 & n457 ) | ( n455 & n457 ) ;
  assign n461 = ~x23 & n460 ;
  assign n462 = ( ~x23 & n459 ) | ( ~x23 & n461 ) | ( n459 & n461 ) ;
  assign n463 = x22 & n462 ;
  assign n464 = x24 & n460 ;
  assign n465 = ( x24 & n459 ) | ( x24 & n464 ) | ( n459 & n464 ) ;
  assign n466 = x24 | n452 ;
  assign n467 = ( x24 & ~n458 ) | ( x24 & n466 ) | ( ~n458 & n466 ) ;
  assign n468 = ( x23 & n465 ) | ( x23 & ~n467 ) | ( n465 & ~n467 ) ;
  assign n469 = ( x22 & n463 ) | ( x22 & n468 ) | ( n463 & n468 ) ;
  assign n470 = ( x22 & ~n465 ) | ( x22 & n467 ) | ( ~n465 & n467 ) ;
  assign n471 = x20 | n470 ;
  assign n472 = ( x20 & ~n469 ) | ( x20 & n471 ) | ( ~n469 & n471 ) ;
  assign n473 = x19 & ~n472 ;
  assign n474 = x21 & ~n470 ;
  assign n475 = ( x21 & n469 ) | ( x21 & n474 ) | ( n469 & n474 ) ;
  assign n476 = ~x21 & n462 ;
  assign n477 = ( ~x21 & n468 ) | ( ~x21 & n476 ) | ( n468 & n476 ) ;
  assign n478 = ( x20 & n475 ) | ( x20 & n477 ) | ( n475 & n477 ) ;
  assign n479 = ( x19 & n473 ) | ( x19 & n478 ) | ( n473 & n478 ) ;
  assign n480 = ( ~x19 & n475 ) | ( ~x19 & n477 ) | ( n475 & n477 ) ;
  assign n481 = ~x17 & n480 ;
  assign n482 = ( ~x17 & n479 ) | ( ~x17 & n481 ) | ( n479 & n481 ) ;
  assign n483 = x16 & n482 ;
  assign n484 = x18 & n480 ;
  assign n485 = ( x18 & n479 ) | ( x18 & n484 ) | ( n479 & n484 ) ;
  assign n486 = x18 | n472 ;
  assign n487 = ( x18 & ~n478 ) | ( x18 & n486 ) | ( ~n478 & n486 ) ;
  assign n488 = ( x17 & n485 ) | ( x17 & ~n487 ) | ( n485 & ~n487 ) ;
  assign n489 = ( x16 & n483 ) | ( x16 & n488 ) | ( n483 & n488 ) ;
  assign n490 = ( x16 & ~n485 ) | ( x16 & n487 ) | ( ~n485 & n487 ) ;
  assign n491 = x14 | n490 ;
  assign n492 = ( x14 & ~n489 ) | ( x14 & n491 ) | ( ~n489 & n491 ) ;
  assign n493 = x13 & ~n492 ;
  assign n494 = x15 & ~n490 ;
  assign n495 = ( x15 & n489 ) | ( x15 & n494 ) | ( n489 & n494 ) ;
  assign n496 = ~x15 & n482 ;
  assign n497 = ( ~x15 & n488 ) | ( ~x15 & n496 ) | ( n488 & n496 ) ;
  assign n498 = ( x14 & n495 ) | ( x14 & n497 ) | ( n495 & n497 ) ;
  assign n499 = ( x13 & n493 ) | ( x13 & n498 ) | ( n493 & n498 ) ;
  assign n500 = ( ~x13 & n495 ) | ( ~x13 & n497 ) | ( n495 & n497 ) ;
  assign n501 = ~x11 & n500 ;
  assign n502 = ( ~x11 & n499 ) | ( ~x11 & n501 ) | ( n499 & n501 ) ;
  assign n503 = x10 & n502 ;
  assign n504 = x12 & n500 ;
  assign n505 = ( x12 & n499 ) | ( x12 & n504 ) | ( n499 & n504 ) ;
  assign n506 = x12 | n492 ;
  assign n507 = ( x12 & ~n498 ) | ( x12 & n506 ) | ( ~n498 & n506 ) ;
  assign n508 = ( x11 & n505 ) | ( x11 & ~n507 ) | ( n505 & ~n507 ) ;
  assign n509 = ( x10 & n503 ) | ( x10 & n508 ) | ( n503 & n508 ) ;
  assign n510 = ( x10 & ~n505 ) | ( x10 & n507 ) | ( ~n505 & n507 ) ;
  assign n511 = x8 | n510 ;
  assign n512 = ( x8 & ~n509 ) | ( x8 & n511 ) | ( ~n509 & n511 ) ;
  assign n513 = x7 & ~n512 ;
  assign n514 = x9 & ~n510 ;
  assign n515 = ( x9 & n509 ) | ( x9 & n514 ) | ( n509 & n514 ) ;
  assign n516 = ~x9 & n502 ;
  assign n517 = ( ~x9 & n508 ) | ( ~x9 & n516 ) | ( n508 & n516 ) ;
  assign n518 = ( x8 & n515 ) | ( x8 & n517 ) | ( n515 & n517 ) ;
  assign n519 = ( x7 & n513 ) | ( x7 & n518 ) | ( n513 & n518 ) ;
  assign n520 = ( ~x7 & n515 ) | ( ~x7 & n517 ) | ( n515 & n517 ) ;
  assign n521 = ~x5 & n520 ;
  assign n522 = ( ~x5 & n519 ) | ( ~x5 & n521 ) | ( n519 & n521 ) ;
  assign n523 = x4 & n522 ;
  assign n524 = x6 & n520 ;
  assign n525 = ( x6 & n519 ) | ( x6 & n524 ) | ( n519 & n524 ) ;
  assign n526 = x6 | n512 ;
  assign n527 = ( x6 & ~n518 ) | ( x6 & n526 ) | ( ~n518 & n526 ) ;
  assign n528 = ( x5 & n525 ) | ( x5 & ~n527 ) | ( n525 & ~n527 ) ;
  assign n529 = ( x4 & n523 ) | ( x4 & n528 ) | ( n523 & n528 ) ;
  assign n530 = ( x4 & ~n525 ) | ( x4 & n527 ) | ( ~n525 & n527 ) ;
  assign n531 = x3 & ~n530 ;
  assign n532 = ( x3 & n529 ) | ( x3 & n531 ) | ( n529 & n531 ) ;
  assign n533 = x1 & ~x2 ;
  assign n534 = ~x3 & n522 ;
  assign n535 = ( ~x3 & n528 ) | ( ~x3 & n534 ) | ( n528 & n534 ) ;
  assign n536 = n533 | n535 ;
  assign n537 = n532 | n536 ;
  assign n538 = n530 & n533 ;
  assign n539 = ~n529 & n538 ;
  assign n540 = n537 & ~n539 ;
  assign n541 = x8 | x9 ;
  assign n542 = x12 | x13 ;
  assign n543 = x16 | x17 ;
  assign n544 = x20 | x21 ;
  assign n545 = x24 | x25 ;
  assign n546 = x28 | x29 ;
  assign n547 = x32 | x33 ;
  assign n548 = x36 | x37 ;
  assign n549 = x40 | x41 ;
  assign n550 = x44 | x45 ;
  assign n551 = x48 | x49 ;
  assign n552 = x52 | x53 ;
  assign n553 = x56 | x57 ;
  assign n554 = x60 | x61 ;
  assign n555 = x64 | x65 ;
  assign n556 = x68 | x69 ;
  assign n557 = x72 | x73 ;
  assign n558 = x76 | x77 ;
  assign n559 = x80 | x81 ;
  assign n560 = x84 | x85 ;
  assign n561 = x88 | x89 ;
  assign n562 = x92 | x93 ;
  assign n563 = x96 | x97 ;
  assign n564 = x100 | x101 ;
  assign n565 = x104 | x105 ;
  assign n566 = x108 | x109 ;
  assign n567 = x124 | x125 ;
  assign n568 = x122 | x123 ;
  assign n569 = ~n567 & n568 ;
  assign n570 = x126 | x127 ;
  assign n571 = n569 | n570 ;
  assign n572 = n567 | n570 ;
  assign n573 = x120 | x121 ;
  assign n574 = n568 | n573 ;
  assign n575 = n572 | n574 ;
  assign n576 = ~n571 & n575 ;
  assign n577 = x118 | x119 ;
  assign n578 = n571 | n577 ;
  assign n579 = ~n576 & n578 ;
  assign n580 = x114 | x115 ;
  assign n581 = n579 | n580 ;
  assign n582 = x117 | n577 ;
  assign n583 = x116 | n582 ;
  assign n584 = ( n576 & ~n578 ) | ( n576 & n583 ) | ( ~n578 & n583 ) ;
  assign n585 = ( n576 & n583 ) | ( n576 & n584 ) | ( n583 & n584 ) ;
  assign n586 = n581 & ~n585 ;
  assign n587 = x112 | x113 ;
  assign n588 = ( n580 & n583 ) | ( n580 & ~n587 ) | ( n583 & ~n587 ) ;
  assign n589 = n587 | n588 ;
  assign n590 = n575 | n589 ;
  assign n591 = ~n586 & n590 ;
  assign n592 = n566 | n591 ;
  assign n593 = x110 | x111 ;
  assign n594 = n586 | n593 ;
  assign n595 = ~n591 & n594 ;
  assign n596 = n592 & ~n595 ;
  assign n597 = n565 | n596 ;
  assign n598 = x106 | x107 ;
  assign n599 = n595 | n598 ;
  assign n600 = ~n596 & n599 ;
  assign n601 = n597 & ~n600 ;
  assign n602 = n564 | n601 ;
  assign n603 = x102 | x103 ;
  assign n604 = n600 | n603 ;
  assign n605 = ~n601 & n604 ;
  assign n606 = n602 & ~n605 ;
  assign n607 = n563 | n606 ;
  assign n608 = x98 | x99 ;
  assign n609 = n605 | n608 ;
  assign n610 = ~n606 & n609 ;
  assign n611 = n607 & ~n610 ;
  assign n612 = n562 | n611 ;
  assign n613 = x94 | x95 ;
  assign n614 = n610 | n613 ;
  assign n615 = ~n611 & n614 ;
  assign n616 = n612 & ~n615 ;
  assign n617 = n561 | n616 ;
  assign n618 = x90 | x91 ;
  assign n619 = n615 | n618 ;
  assign n620 = ~n616 & n619 ;
  assign n621 = n617 & ~n620 ;
  assign n622 = n560 | n621 ;
  assign n623 = x86 | x87 ;
  assign n624 = n620 | n623 ;
  assign n625 = ~n621 & n624 ;
  assign n626 = n622 & ~n625 ;
  assign n627 = n559 | n626 ;
  assign n628 = x82 | x83 ;
  assign n629 = n625 | n628 ;
  assign n630 = ~n626 & n629 ;
  assign n631 = n627 & ~n630 ;
  assign n632 = n558 | n631 ;
  assign n633 = x78 | x79 ;
  assign n634 = n630 | n633 ;
  assign n635 = ~n631 & n634 ;
  assign n636 = n632 & ~n635 ;
  assign n637 = n557 | n636 ;
  assign n638 = x74 | x75 ;
  assign n639 = n635 | n638 ;
  assign n640 = ~n636 & n639 ;
  assign n641 = n637 & ~n640 ;
  assign n642 = n556 | n641 ;
  assign n643 = x70 | x71 ;
  assign n644 = n640 | n643 ;
  assign n645 = ~n641 & n644 ;
  assign n646 = n642 & ~n645 ;
  assign n647 = n555 | n646 ;
  assign n648 = x66 | x67 ;
  assign n649 = n645 | n648 ;
  assign n650 = ~n646 & n649 ;
  assign n651 = n647 & ~n650 ;
  assign n652 = n554 | n651 ;
  assign n653 = x62 | x63 ;
  assign n654 = n650 | n653 ;
  assign n655 = ~n651 & n654 ;
  assign n656 = n652 & ~n655 ;
  assign n657 = n553 | n656 ;
  assign n658 = x58 | x59 ;
  assign n659 = n655 | n658 ;
  assign n660 = ~n656 & n659 ;
  assign n661 = n657 & ~n660 ;
  assign n662 = n552 | n661 ;
  assign n663 = x54 | x55 ;
  assign n664 = n660 | n663 ;
  assign n665 = ~n661 & n664 ;
  assign n666 = n662 & ~n665 ;
  assign n667 = n551 | n666 ;
  assign n668 = x50 | x51 ;
  assign n669 = n665 | n668 ;
  assign n670 = ~n666 & n669 ;
  assign n671 = n667 & ~n670 ;
  assign n672 = n550 | n671 ;
  assign n673 = x46 | x47 ;
  assign n674 = n670 | n673 ;
  assign n675 = ~n671 & n674 ;
  assign n676 = n672 & ~n675 ;
  assign n677 = n549 | n676 ;
  assign n678 = x42 | x43 ;
  assign n679 = n675 | n678 ;
  assign n680 = ~n676 & n679 ;
  assign n681 = n677 & ~n680 ;
  assign n682 = n548 | n681 ;
  assign n683 = x38 | x39 ;
  assign n684 = n680 | n683 ;
  assign n685 = ~n681 & n684 ;
  assign n686 = n682 & ~n685 ;
  assign n687 = n547 | n686 ;
  assign n688 = x34 | x35 ;
  assign n689 = n685 | n688 ;
  assign n690 = ~n686 & n689 ;
  assign n691 = n687 & ~n690 ;
  assign n692 = n546 | n691 ;
  assign n693 = x30 | x31 ;
  assign n694 = n690 | n693 ;
  assign n695 = ~n691 & n694 ;
  assign n696 = n692 & ~n695 ;
  assign n697 = n545 | n696 ;
  assign n698 = x26 | x27 ;
  assign n699 = n695 | n698 ;
  assign n700 = ~n696 & n699 ;
  assign n701 = n697 & ~n700 ;
  assign n702 = n544 | n701 ;
  assign n703 = x22 | x23 ;
  assign n704 = n700 | n703 ;
  assign n705 = ~n701 & n704 ;
  assign n706 = n702 & ~n705 ;
  assign n707 = n543 | n706 ;
  assign n708 = x18 | x19 ;
  assign n709 = n705 | n708 ;
  assign n710 = ~n706 & n709 ;
  assign n711 = n707 & ~n710 ;
  assign n712 = n542 | n711 ;
  assign n713 = x14 | x15 ;
  assign n714 = n710 | n713 ;
  assign n715 = ~n711 & n714 ;
  assign n716 = n712 & ~n715 ;
  assign n717 = n541 | n716 ;
  assign n718 = x10 | x11 ;
  assign n719 = n715 | n718 ;
  assign n720 = ~n716 & n719 ;
  assign n721 = n717 & ~n720 ;
  assign n722 = x6 | x7 ;
  assign n723 = n720 | n722 ;
  assign n724 = x2 | x3 ;
  assign n725 = x4 | x5 ;
  assign n726 = n723 | n725 ;
  assign n727 = n724 & ~n726 ;
  assign n728 = ( ~n721 & n723 ) | ( ~n721 & n727 ) | ( n723 & n727 ) ;
  assign n729 = x5 | n722 ;
  assign n730 = x4 | n729 ;
  assign n731 = x89 | n618 ;
  assign n732 = x88 | n731 ;
  assign n733 = ~n574 & n583 ;
  assign n734 = n572 | n733 ;
  assign n735 = x109 | n593 ;
  assign n736 = x108 | n735 ;
  assign n737 = x113 | x114 ;
  assign n738 = x112 | n737 ;
  assign n739 = x115 & ~n583 ;
  assign n740 = n574 | n739 ;
  assign n741 = ( ~n572 & n738 ) | ( ~n572 & n740 ) | ( n738 & n740 ) ;
  assign n742 = ~n734 & n741 ;
  assign n743 = n736 & ~n742 ;
  assign n744 = n734 | n743 ;
  assign n745 = x101 | n603 ;
  assign n746 = x100 | n745 ;
  assign n747 = n598 & ~n744 ;
  assign n748 = ( n565 & ~n744 ) | ( n565 & n747 ) | ( ~n744 & n747 ) ;
  assign n749 = n742 | n748 ;
  assign n750 = n746 & ~n749 ;
  assign n751 = n744 | n750 ;
  assign n752 = x93 | n613 ;
  assign n753 = x92 | n752 ;
  assign n754 = n608 & ~n751 ;
  assign n755 = ( n563 & ~n751 ) | ( n563 & n754 ) | ( ~n751 & n754 ) ;
  assign n756 = n749 | n755 ;
  assign n757 = n753 & ~n756 ;
  assign n758 = n751 | n757 ;
  assign n759 = n732 & ~n758 ;
  assign n760 = ~n732 & n756 ;
  assign n761 = n759 | n760 ;
  assign n762 = x85 | n623 ;
  assign n763 = x84 | n762 ;
  assign n764 = ~n761 & n763 ;
  assign n765 = n758 & ~n763 ;
  assign n766 = n764 | n765 ;
  assign n767 = x81 | n628 ;
  assign n768 = x80 | n767 ;
  assign n769 = ~n766 & n768 ;
  assign n770 = n761 & ~n768 ;
  assign n771 = n769 | n770 ;
  assign n772 = x77 | n633 ;
  assign n773 = x76 | n772 ;
  assign n774 = ~n771 & n773 ;
  assign n775 = n766 & ~n773 ;
  assign n776 = n774 | n775 ;
  assign n777 = x73 | n638 ;
  assign n778 = x72 | n777 ;
  assign n779 = ~n776 & n778 ;
  assign n780 = n771 & ~n778 ;
  assign n781 = n779 | n780 ;
  assign n782 = x69 | n643 ;
  assign n783 = x68 | n782 ;
  assign n784 = ~n781 & n783 ;
  assign n785 = n776 & ~n783 ;
  assign n786 = n784 | n785 ;
  assign n787 = x65 | n648 ;
  assign n788 = x64 | n787 ;
  assign n789 = ~n786 & n788 ;
  assign n790 = n781 & ~n788 ;
  assign n791 = n789 | n790 ;
  assign n792 = x61 | n653 ;
  assign n793 = x60 | n792 ;
  assign n794 = ~n791 & n793 ;
  assign n795 = n786 & ~n793 ;
  assign n796 = n794 | n795 ;
  assign n797 = x57 | n658 ;
  assign n798 = x56 | n797 ;
  assign n799 = ~n796 & n798 ;
  assign n800 = n791 & ~n798 ;
  assign n801 = n799 | n800 ;
  assign n802 = x53 | n663 ;
  assign n803 = x52 | n802 ;
  assign n804 = ~n801 & n803 ;
  assign n805 = n796 & ~n803 ;
  assign n806 = n804 | n805 ;
  assign n807 = x49 | n668 ;
  assign n808 = x48 | n807 ;
  assign n809 = ~n806 & n808 ;
  assign n810 = n801 & ~n808 ;
  assign n811 = n809 | n810 ;
  assign n812 = x45 | n673 ;
  assign n813 = x44 | n812 ;
  assign n814 = ~n811 & n813 ;
  assign n815 = n806 & ~n813 ;
  assign n816 = n814 | n815 ;
  assign n817 = x41 | n678 ;
  assign n818 = x40 | n817 ;
  assign n819 = ~n816 & n818 ;
  assign n820 = n811 & ~n818 ;
  assign n821 = n819 | n820 ;
  assign n822 = x37 | n683 ;
  assign n823 = x36 | n822 ;
  assign n824 = ~n821 & n823 ;
  assign n825 = n816 & ~n823 ;
  assign n826 = n824 | n825 ;
  assign n827 = x33 | n688 ;
  assign n828 = x32 | n827 ;
  assign n829 = ~n826 & n828 ;
  assign n830 = n821 & ~n828 ;
  assign n831 = n829 | n830 ;
  assign n832 = x29 | n693 ;
  assign n833 = x28 | n832 ;
  assign n834 = ~n831 & n833 ;
  assign n835 = n826 & ~n833 ;
  assign n836 = n834 | n835 ;
  assign n837 = x25 | n698 ;
  assign n838 = x24 | n837 ;
  assign n839 = ~n836 & n838 ;
  assign n840 = n831 & ~n838 ;
  assign n841 = n839 | n840 ;
  assign n842 = x21 | n703 ;
  assign n843 = x20 | n842 ;
  assign n844 = ~n841 & n843 ;
  assign n845 = n836 & ~n843 ;
  assign n846 = n844 | n845 ;
  assign n847 = x17 | n708 ;
  assign n848 = x16 | n847 ;
  assign n849 = ~n846 & n848 ;
  assign n850 = n841 & ~n848 ;
  assign n851 = n849 | n850 ;
  assign n852 = n718 & n730 ;
  assign n853 = ( n541 & n730 ) | ( n541 & n852 ) | ( n730 & n852 ) ;
  assign n854 = ( n730 & ~n851 ) | ( n730 & n853 ) | ( ~n851 & n853 ) ;
  assign n855 = x13 | n713 ;
  assign n856 = x12 | n855 ;
  assign n857 = ~n851 & n856 ;
  assign n858 = n846 & ~n856 ;
  assign n859 = n857 | n858 ;
  assign n860 = ( n730 & ~n853 ) | ( n730 & n859 ) | ( ~n853 & n859 ) ;
  assign n861 = ( ~n730 & n854 ) | ( ~n730 & n860 ) | ( n854 & n860 ) ;
  assign n862 = ( n541 & ~n718 ) | ( n541 & n856 ) | ( ~n718 & n856 ) ;
  assign n863 = n718 | n862 ;
  assign n864 = ( n565 & ~n598 ) | ( n565 & n736 ) | ( ~n598 & n736 ) ;
  assign n865 = n598 | n864 ;
  assign n866 = ~n589 & n865 ;
  assign n867 = n575 | n866 ;
  assign n868 = ( x102 & ~n564 ) | ( x102 & n608 ) | ( ~n564 & n608 ) ;
  assign n869 = n564 | n868 ;
  assign n870 = x97 | n869 ;
  assign n871 = x96 | n870 ;
  assign n872 = x103 & ~n865 ;
  assign n873 = n589 | n872 ;
  assign n874 = ( ~n575 & n871 ) | ( ~n575 & n873 ) | ( n871 & n873 ) ;
  assign n875 = ~n867 & n874 ;
  assign n876 = ( n561 & ~n618 ) | ( n561 & n753 ) | ( ~n618 & n753 ) ;
  assign n877 = n618 | n876 ;
  assign n878 = ~n875 & n877 ;
  assign n879 = n867 | n878 ;
  assign n880 = ( n559 & ~n628 ) | ( n559 & n763 ) | ( ~n628 & n763 ) ;
  assign n881 = n628 | n880 ;
  assign n882 = ~n879 & n881 ;
  assign n883 = n875 | n882 ;
  assign n884 = ( n557 & ~n638 ) | ( n557 & n773 ) | ( ~n638 & n773 ) ;
  assign n885 = n638 | n884 ;
  assign n886 = ~n883 & n885 ;
  assign n887 = n879 | n886 ;
  assign n888 = ( n555 & ~n648 ) | ( n555 & n783 ) | ( ~n648 & n783 ) ;
  assign n889 = n648 | n888 ;
  assign n890 = ~n887 & n889 ;
  assign n891 = n883 | n890 ;
  assign n892 = ( n553 & ~n658 ) | ( n553 & n793 ) | ( ~n658 & n793 ) ;
  assign n893 = n658 | n892 ;
  assign n894 = ~n891 & n893 ;
  assign n895 = n887 | n894 ;
  assign n896 = ( n551 & ~n668 ) | ( n551 & n803 ) | ( ~n668 & n803 ) ;
  assign n897 = n668 | n896 ;
  assign n898 = ~n895 & n897 ;
  assign n899 = n891 & ~n897 ;
  assign n900 = n898 | n899 ;
  assign n901 = ( n549 & ~n678 ) | ( n549 & n813 ) | ( ~n678 & n813 ) ;
  assign n902 = n678 | n901 ;
  assign n903 = ~n900 & n902 ;
  assign n904 = n895 & ~n902 ;
  assign n905 = n903 | n904 ;
  assign n906 = ( n547 & ~n688 ) | ( n547 & n823 ) | ( ~n688 & n823 ) ;
  assign n907 = n688 | n906 ;
  assign n908 = ~n905 & n907 ;
  assign n909 = n900 & ~n907 ;
  assign n910 = n908 | n909 ;
  assign n911 = ( n543 & ~n708 ) | ( n543 & n843 ) | ( ~n708 & n843 ) ;
  assign n912 = n708 | n911 ;
  assign n913 = n863 & n912 ;
  assign n914 = ( n863 & ~n910 ) | ( n863 & n913 ) | ( ~n910 & n913 ) ;
  assign n915 = ( n545 & ~n698 ) | ( n545 & n833 ) | ( ~n698 & n833 ) ;
  assign n916 = n698 | n915 ;
  assign n917 = ~n910 & n916 ;
  assign n918 = n905 & ~n916 ;
  assign n919 = n917 | n918 ;
  assign n920 = ( n863 & ~n913 ) | ( n863 & n919 ) | ( ~n913 & n919 ) ;
  assign n921 = ( ~n863 & n914 ) | ( ~n863 & n920 ) | ( n914 & n920 ) ;
  assign n922 = ( n544 & ~n703 ) | ( n544 & n916 ) | ( ~n703 & n916 ) ;
  assign n923 = n703 | n922 ;
  assign n924 = ( n543 & ~n708 ) | ( n543 & n923 ) | ( ~n708 & n923 ) ;
  assign n925 = n708 | n924 ;
  assign n926 = ( n548 & ~n683 ) | ( n548 & n902 ) | ( ~n683 & n902 ) ;
  assign n927 = n683 | n926 ;
  assign n928 = ( n547 & ~n688 ) | ( n547 & n927 ) | ( ~n688 & n927 ) ;
  assign n929 = n688 | n928 ;
  assign n930 = n925 & n929 ;
  assign n931 = x99 | n746 ;
  assign n932 = ( x98 & ~n563 ) | ( x98 & n865 ) | ( ~n563 & n865 ) ;
  assign n933 = n563 | n932 ;
  assign n934 = n931 | n933 ;
  assign n935 = ( n560 & ~n623 ) | ( n560 & n877 ) | ( ~n623 & n877 ) ;
  assign n936 = n623 | n935 ;
  assign n937 = ( n559 & ~n628 ) | ( n559 & n936 ) | ( ~n628 & n936 ) ;
  assign n938 = n628 | n937 ;
  assign n939 = x79 & ~n938 ;
  assign n940 = n934 | n939 ;
  assign n941 = ( x78 & ~n558 ) | ( x78 & n638 ) | ( ~n558 & n638 ) ;
  assign n942 = n558 | n941 ;
  assign n943 = ( ~n557 & n643 ) | ( ~n557 & n942 ) | ( n643 & n942 ) ;
  assign n944 = n557 | n943 ;
  assign n945 = x69 | n944 ;
  assign n946 = x68 | n945 ;
  assign n947 = ( n555 & ~n648 ) | ( n555 & n946 ) | ( ~n648 & n946 ) ;
  assign n948 = n648 | n947 ;
  assign n949 = ( ~n590 & n940 ) | ( ~n590 & n948 ) | ( n940 & n948 ) ;
  assign n950 = ~n934 & n938 ;
  assign n951 = n590 | n950 ;
  assign n952 = n949 & ~n951 ;
  assign n953 = ( n925 & n930 ) | ( n925 & ~n952 ) | ( n930 & ~n952 ) ;
  assign n954 = ( n552 & ~n663 ) | ( n552 & n893 ) | ( ~n663 & n893 ) ;
  assign n955 = n663 | n954 ;
  assign n956 = ( n551 & ~n668 ) | ( n551 & n955 ) | ( ~n668 & n955 ) ;
  assign n957 = n668 | n956 ;
  assign n958 = ~n952 & n957 ;
  assign n959 = n951 | n958 ;
  assign n960 = ( n925 & ~n930 ) | ( n925 & n959 ) | ( ~n930 & n959 ) ;
  assign n961 = ( ~n925 & n953 ) | ( ~n925 & n960 ) | ( n953 & n960 ) ;
  assign n962 = n590 | n934 ;
  assign n963 = x71 | n885 ;
  assign n964 = ( x70 & ~n556 ) | ( x70 & n938 ) | ( ~n556 & n938 ) ;
  assign n965 = ( n556 & ~n648 ) | ( n556 & n964 ) | ( ~n648 & n964 ) ;
  assign n966 = n648 | n965 ;
  assign n967 = ( ~n555 & n963 ) | ( ~n555 & n966 ) | ( n963 & n966 ) ;
  assign n968 = n555 | n967 ;
  assign n969 = ( n550 & ~n673 ) | ( n550 & n957 ) | ( ~n673 & n957 ) ;
  assign n970 = n673 | n969 ;
  assign n971 = ( n549 & ~n678 ) | ( n549 & n970 ) | ( ~n678 & n970 ) ;
  assign n972 = n678 | n971 ;
  assign n973 = ( n548 & ~n683 ) | ( n548 & n972 ) | ( ~n683 & n972 ) ;
  assign n974 = n683 | n973 ;
  assign n975 = ( n547 & ~n688 ) | ( n547 & n974 ) | ( ~n688 & n974 ) ;
  assign n976 = n688 | n975 ;
  assign n977 = ~n968 & n976 ;
  assign n978 = n962 | n977 ;
  assign n979 = n962 | n968 ;
  assign n980 = n925 | n976 ;
  assign n981 = n730 | n980 ;
  assign n982 = x1 | n981 ;
  assign n983 = x0 | n979 ;
  assign n984 = ( ~n724 & n863 ) | ( ~n724 & n983 ) | ( n863 & n983 ) ;
  assign n985 = n724 | n984 ;
  assign n986 = n982 | n985 ;
  assign y0 = n540 ;
  assign y1 = n728 ;
  assign y2 = n861 ;
  assign y3 = n921 ;
  assign y4 = n961 ;
  assign y5 = n978 ;
  assign y6 = n979 ;
  assign y7 = n986 ;
endmodule
