module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 ;
  wire n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 ;
  assign n97 = ( x0 & ~x1 ) | ( x0 & x2 ) | ( ~x1 & x2 ) ;
  assign n98 = ( ~x0 & x1 ) | ( ~x0 & n97 ) | ( x1 & n97 ) ;
  assign n99 = ( ~x2 & n97 ) | ( ~x2 & n98 ) | ( n97 & n98 ) ;
  assign n100 = x1 & x2 ;
  assign n101 = x1 | x2 ;
  assign n102 = x0 & n101 ;
  assign n103 = n100 | n102 ;
  assign n104 = ~x3 & n103 ;
  assign n105 = x0 | n100 ;
  assign n106 = n101 & n105 ;
  assign n107 = x3 & ~n106 ;
  assign n108 = n104 | n107 ;
  assign n109 = ( x4 & ~x5 ) | ( x4 & n108 ) | ( ~x5 & n108 ) ;
  assign n110 = x3 & n103 ;
  assign n111 = x3 | n106 ;
  assign n112 = ~n110 & n111 ;
  assign n113 = ( x5 & n109 ) | ( x5 & ~n112 ) | ( n109 & ~n112 ) ;
  assign n114 = ( ~x4 & n109 ) | ( ~x4 & n113 ) | ( n109 & n113 ) ;
  assign n115 = x0 & x1 ;
  assign n116 = ( x3 & x4 ) | ( x3 & n115 ) | ( x4 & n115 ) ;
  assign n117 = ( ~x6 & x7 ) | ( ~x6 & n116 ) | ( x7 & n116 ) ;
  assign n118 = x3 | x4 ;
  assign n119 = x3 & x4 ;
  assign n120 = n115 | n119 ;
  assign n121 = n118 & n120 ;
  assign n122 = ( x7 & ~n117 ) | ( x7 & n121 ) | ( ~n117 & n121 ) ;
  assign n123 = ( x6 & n117 ) | ( x6 & ~n122 ) | ( n117 & ~n122 ) ;
  assign n124 = ( ~x0 & x3 ) | ( ~x0 & x4 ) | ( x3 & x4 ) ;
  assign n125 = ( x1 & x3 ) | ( x1 & x4 ) | ( x3 & x4 ) ;
  assign n126 = ~n124 & n125 ;
  assign n127 = n118 & ~n119 ;
  assign n128 = x0 | x1 ;
  assign n129 = x2 & n128 ;
  assign n130 = x5 | n129 ;
  assign n131 = ( x0 & x1 ) | ( x0 & x2 ) | ( x1 & x2 ) ;
  assign n132 = x5 & n131 ;
  assign n133 = ( n127 & n130 ) | ( n127 & n132 ) | ( n130 & n132 ) ;
  assign n134 = ~n126 & n133 ;
  assign n135 = ( x8 & n123 ) | ( x8 & ~n134 ) | ( n123 & ~n134 ) ;
  assign n136 = ( ~x8 & n134 ) | ( ~x8 & n135 ) | ( n134 & n135 ) ;
  assign n137 = ( ~n123 & n135 ) | ( ~n123 & n136 ) | ( n135 & n136 ) ;
  assign n138 = x6 & x7 ;
  assign n139 = x6 | x7 ;
  assign n140 = n116 & n139 ;
  assign n141 = n138 | n140 ;
  assign n142 = x9 & x10 ;
  assign n143 = x9 | x10 ;
  assign n144 = ~n142 & n143 ;
  assign n145 = x8 | n123 ;
  assign n146 = x8 & n123 ;
  assign n147 = n134 | n146 ;
  assign n148 = n145 & n147 ;
  assign n149 = n144 & ~n148 ;
  assign n150 = n134 & n145 ;
  assign n151 = n146 | n150 ;
  assign n152 = ~n144 & n151 ;
  assign n153 = n149 | n152 ;
  assign n154 = ( x11 & ~n141 ) | ( x11 & n153 ) | ( ~n141 & n153 ) ;
  assign n155 = n144 | n148 ;
  assign n156 = n144 & n151 ;
  assign n157 = n155 & ~n156 ;
  assign n158 = ( n141 & n154 ) | ( n141 & ~n157 ) | ( n154 & ~n157 ) ;
  assign n159 = ( ~x11 & n154 ) | ( ~x11 & n158 ) | ( n154 & n158 ) ;
  assign n160 = x12 & x13 ;
  assign n161 = n141 | n142 ;
  assign n162 = n143 & n161 ;
  assign n163 = ( x12 & x13 ) | ( x12 & ~n162 ) | ( x13 & ~n162 ) ;
  assign n164 = x12 | x13 ;
  assign n165 = ~n160 & n164 ;
  assign n166 = ( x9 & x10 ) | ( x9 & n141 ) | ( x10 & n141 ) ;
  assign n167 = ~n165 & n166 ;
  assign n168 = ( ~n160 & n163 ) | ( ~n160 & n167 ) | ( n163 & n167 ) ;
  assign n169 = n141 | n144 ;
  assign n170 = n141 & n144 ;
  assign n171 = n169 & ~n170 ;
  assign n172 = ( x8 & n123 ) | ( x8 & n134 ) | ( n123 & n134 ) ;
  assign n173 = ( x11 & n171 ) | ( x11 & n172 ) | ( n171 & n172 ) ;
  assign n174 = ( x14 & n168 ) | ( x14 & ~n173 ) | ( n168 & ~n173 ) ;
  assign n175 = ( ~x14 & n173 ) | ( ~x14 & n174 ) | ( n173 & n174 ) ;
  assign n176 = ( ~n168 & n174 ) | ( ~n168 & n175 ) | ( n174 & n175 ) ;
  assign n177 = x15 & x16 ;
  assign n178 = x15 | x16 ;
  assign n179 = ~n177 & n178 ;
  assign n180 = ( x12 & x13 ) | ( x12 & n162 ) | ( x13 & n162 ) ;
  assign n181 = n179 & ~n180 ;
  assign n182 = n165 & n166 ;
  assign n183 = ( n160 & ~n179 ) | ( n160 & n182 ) | ( ~n179 & n182 ) ;
  assign n184 = n181 | n183 ;
  assign n185 = x17 & n184 ;
  assign n186 = x14 | n168 ;
  assign n187 = x14 & n168 ;
  assign n188 = n173 | n187 ;
  assign n189 = n186 & n188 ;
  assign n190 = ( x17 & n184 ) | ( x17 & ~n189 ) | ( n184 & ~n189 ) ;
  assign n191 = x17 | n184 ;
  assign n192 = ~n185 & n191 ;
  assign n193 = n186 & ~n187 ;
  assign n194 = n173 & n193 ;
  assign n195 = ( n187 & ~n192 ) | ( n187 & n194 ) | ( ~n192 & n194 ) ;
  assign n196 = ( ~n185 & n190 ) | ( ~n185 & n195 ) | ( n190 & n195 ) ;
  assign n197 = x18 & x19 ;
  assign n198 = n177 | n180 ;
  assign n199 = n178 & n198 ;
  assign n200 = ( x18 & x19 ) | ( x18 & ~n199 ) | ( x19 & ~n199 ) ;
  assign n201 = x18 | x19 ;
  assign n202 = ~n197 & n201 ;
  assign n203 = ( x15 & x16 ) | ( x15 & n180 ) | ( x16 & n180 ) ;
  assign n204 = ~n202 & n203 ;
  assign n205 = ( ~n197 & n200 ) | ( ~n197 & n204 ) | ( n200 & n204 ) ;
  assign n206 = ( x17 & n184 ) | ( x17 & n189 ) | ( n184 & n189 ) ;
  assign n207 = ( x20 & n205 ) | ( x20 & ~n206 ) | ( n205 & ~n206 ) ;
  assign n208 = ( ~x20 & n206 ) | ( ~x20 & n207 ) | ( n206 & n207 ) ;
  assign n209 = ( ~n205 & n207 ) | ( ~n205 & n208 ) | ( n207 & n208 ) ;
  assign n210 = x21 & x22 ;
  assign n211 = x21 | x22 ;
  assign n212 = ~n210 & n211 ;
  assign n213 = ( x18 & x19 ) | ( x18 & n199 ) | ( x19 & n199 ) ;
  assign n214 = n212 & ~n213 ;
  assign n215 = n202 & n203 ;
  assign n216 = ( n197 & ~n212 ) | ( n197 & n215 ) | ( ~n212 & n215 ) ;
  assign n217 = n214 | n216 ;
  assign n218 = x23 & n217 ;
  assign n219 = x20 | n205 ;
  assign n220 = x20 & n205 ;
  assign n221 = n206 | n220 ;
  assign n222 = n219 & n221 ;
  assign n223 = ( x23 & n217 ) | ( x23 & ~n222 ) | ( n217 & ~n222 ) ;
  assign n224 = x23 | n217 ;
  assign n225 = ~n218 & n224 ;
  assign n226 = n219 & ~n220 ;
  assign n227 = n206 & n226 ;
  assign n228 = ( n220 & ~n225 ) | ( n220 & n227 ) | ( ~n225 & n227 ) ;
  assign n229 = ( ~n218 & n223 ) | ( ~n218 & n228 ) | ( n223 & n228 ) ;
  assign n230 = x24 & x25 ;
  assign n231 = n210 | n213 ;
  assign n232 = n211 & n231 ;
  assign n233 = ( x24 & x25 ) | ( x24 & ~n232 ) | ( x25 & ~n232 ) ;
  assign n234 = x24 | x25 ;
  assign n235 = ~n230 & n234 ;
  assign n236 = ( x21 & x22 ) | ( x21 & n213 ) | ( x22 & n213 ) ;
  assign n237 = ~n235 & n236 ;
  assign n238 = ( ~n230 & n233 ) | ( ~n230 & n237 ) | ( n233 & n237 ) ;
  assign n239 = ( x23 & n217 ) | ( x23 & n222 ) | ( n217 & n222 ) ;
  assign n240 = ( x26 & n238 ) | ( x26 & ~n239 ) | ( n238 & ~n239 ) ;
  assign n241 = ( ~x26 & n239 ) | ( ~x26 & n240 ) | ( n239 & n240 ) ;
  assign n242 = ( ~n238 & n240 ) | ( ~n238 & n241 ) | ( n240 & n241 ) ;
  assign n243 = x27 & x28 ;
  assign n244 = x27 | x28 ;
  assign n245 = ~n243 & n244 ;
  assign n246 = ( x24 & x25 ) | ( x24 & n232 ) | ( x25 & n232 ) ;
  assign n247 = n245 & ~n246 ;
  assign n248 = n235 & n236 ;
  assign n249 = ( n230 & ~n245 ) | ( n230 & n248 ) | ( ~n245 & n248 ) ;
  assign n250 = n247 | n249 ;
  assign n251 = x29 & n250 ;
  assign n252 = x26 | n238 ;
  assign n253 = x26 & n238 ;
  assign n254 = n239 | n253 ;
  assign n255 = n252 & n254 ;
  assign n256 = ( x29 & n250 ) | ( x29 & ~n255 ) | ( n250 & ~n255 ) ;
  assign n257 = x29 | n250 ;
  assign n258 = ~n251 & n257 ;
  assign n259 = n252 & ~n253 ;
  assign n260 = n239 & n259 ;
  assign n261 = ( n253 & ~n258 ) | ( n253 & n260 ) | ( ~n258 & n260 ) ;
  assign n262 = ( ~n251 & n256 ) | ( ~n251 & n261 ) | ( n256 & n261 ) ;
  assign n263 = x30 & x31 ;
  assign n264 = n243 | n246 ;
  assign n265 = n244 & n264 ;
  assign n266 = ( x30 & x31 ) | ( x30 & ~n265 ) | ( x31 & ~n265 ) ;
  assign n267 = x30 | x31 ;
  assign n268 = ~n263 & n267 ;
  assign n269 = ( x27 & x28 ) | ( x27 & n246 ) | ( x28 & n246 ) ;
  assign n270 = ~n268 & n269 ;
  assign n271 = ( ~n263 & n266 ) | ( ~n263 & n270 ) | ( n266 & n270 ) ;
  assign n272 = ( x29 & n250 ) | ( x29 & n255 ) | ( n250 & n255 ) ;
  assign n273 = ( x32 & n271 ) | ( x32 & ~n272 ) | ( n271 & ~n272 ) ;
  assign n274 = ( ~x32 & n272 ) | ( ~x32 & n273 ) | ( n272 & n273 ) ;
  assign n275 = ( ~n271 & n273 ) | ( ~n271 & n274 ) | ( n273 & n274 ) ;
  assign n276 = x33 & x34 ;
  assign n277 = x33 | x34 ;
  assign n278 = ~n276 & n277 ;
  assign n279 = ( x30 & x31 ) | ( x30 & n265 ) | ( x31 & n265 ) ;
  assign n280 = n278 & ~n279 ;
  assign n281 = n268 & n269 ;
  assign n282 = ( n263 & ~n278 ) | ( n263 & n281 ) | ( ~n278 & n281 ) ;
  assign n283 = n280 | n282 ;
  assign n284 = x35 & n283 ;
  assign n285 = x32 | n271 ;
  assign n286 = x32 & n271 ;
  assign n287 = n272 | n286 ;
  assign n288 = n285 & n287 ;
  assign n289 = ( x35 & n283 ) | ( x35 & ~n288 ) | ( n283 & ~n288 ) ;
  assign n290 = x35 | n283 ;
  assign n291 = ~n284 & n290 ;
  assign n292 = n285 & ~n286 ;
  assign n293 = n272 & n292 ;
  assign n294 = ( n286 & ~n291 ) | ( n286 & n293 ) | ( ~n291 & n293 ) ;
  assign n295 = ( ~n284 & n289 ) | ( ~n284 & n294 ) | ( n289 & n294 ) ;
  assign n296 = x36 & x37 ;
  assign n297 = n276 | n279 ;
  assign n298 = n277 & n297 ;
  assign n299 = ( x36 & x37 ) | ( x36 & ~n298 ) | ( x37 & ~n298 ) ;
  assign n300 = x36 | x37 ;
  assign n301 = ~n296 & n300 ;
  assign n302 = ( x33 & x34 ) | ( x33 & n279 ) | ( x34 & n279 ) ;
  assign n303 = ~n301 & n302 ;
  assign n304 = ( ~n296 & n299 ) | ( ~n296 & n303 ) | ( n299 & n303 ) ;
  assign n305 = ( x35 & n283 ) | ( x35 & n288 ) | ( n283 & n288 ) ;
  assign n306 = ( x38 & n304 ) | ( x38 & ~n305 ) | ( n304 & ~n305 ) ;
  assign n307 = ( ~x38 & n305 ) | ( ~x38 & n306 ) | ( n305 & n306 ) ;
  assign n308 = ( ~n304 & n306 ) | ( ~n304 & n307 ) | ( n306 & n307 ) ;
  assign n309 = x39 & x40 ;
  assign n310 = x39 | x40 ;
  assign n311 = ~n309 & n310 ;
  assign n312 = ( x36 & x37 ) | ( x36 & n298 ) | ( x37 & n298 ) ;
  assign n313 = n311 & ~n312 ;
  assign n314 = n301 & n302 ;
  assign n315 = ( n296 & ~n311 ) | ( n296 & n314 ) | ( ~n311 & n314 ) ;
  assign n316 = n313 | n315 ;
  assign n317 = x41 & n316 ;
  assign n318 = x38 | n304 ;
  assign n319 = x38 & n304 ;
  assign n320 = n305 | n319 ;
  assign n321 = n318 & n320 ;
  assign n322 = ( x41 & n316 ) | ( x41 & ~n321 ) | ( n316 & ~n321 ) ;
  assign n323 = x41 | n316 ;
  assign n324 = ~n317 & n323 ;
  assign n325 = n318 & ~n319 ;
  assign n326 = n305 & n325 ;
  assign n327 = ( n319 & ~n324 ) | ( n319 & n326 ) | ( ~n324 & n326 ) ;
  assign n328 = ( ~n317 & n322 ) | ( ~n317 & n327 ) | ( n322 & n327 ) ;
  assign n329 = x42 & x43 ;
  assign n330 = n309 | n312 ;
  assign n331 = n310 & n330 ;
  assign n332 = ( x42 & x43 ) | ( x42 & ~n331 ) | ( x43 & ~n331 ) ;
  assign n333 = x42 | x43 ;
  assign n334 = ~n329 & n333 ;
  assign n335 = ( x39 & x40 ) | ( x39 & n312 ) | ( x40 & n312 ) ;
  assign n336 = ~n334 & n335 ;
  assign n337 = ( ~n329 & n332 ) | ( ~n329 & n336 ) | ( n332 & n336 ) ;
  assign n338 = ( x41 & n316 ) | ( x41 & n321 ) | ( n316 & n321 ) ;
  assign n339 = ( x44 & n337 ) | ( x44 & ~n338 ) | ( n337 & ~n338 ) ;
  assign n340 = ( ~x44 & n338 ) | ( ~x44 & n339 ) | ( n338 & n339 ) ;
  assign n341 = ( ~n337 & n339 ) | ( ~n337 & n340 ) | ( n339 & n340 ) ;
  assign n342 = x45 & x46 ;
  assign n343 = x45 | x46 ;
  assign n344 = ~n342 & n343 ;
  assign n345 = ( x42 & x43 ) | ( x42 & n331 ) | ( x43 & n331 ) ;
  assign n346 = n344 & ~n345 ;
  assign n347 = n334 & n335 ;
  assign n348 = ( n329 & ~n344 ) | ( n329 & n347 ) | ( ~n344 & n347 ) ;
  assign n349 = n346 | n348 ;
  assign n350 = x47 & n349 ;
  assign n351 = x44 | n337 ;
  assign n352 = x44 & n337 ;
  assign n353 = n338 | n352 ;
  assign n354 = n351 & n353 ;
  assign n355 = ( x47 & n349 ) | ( x47 & ~n354 ) | ( n349 & ~n354 ) ;
  assign n356 = x47 | n349 ;
  assign n357 = ~n350 & n356 ;
  assign n358 = n351 & ~n352 ;
  assign n359 = n338 & n358 ;
  assign n360 = ( n352 & ~n357 ) | ( n352 & n359 ) | ( ~n357 & n359 ) ;
  assign n361 = ( ~n350 & n355 ) | ( ~n350 & n360 ) | ( n355 & n360 ) ;
  assign n362 = x48 & x49 ;
  assign n363 = n342 | n345 ;
  assign n364 = n343 & n363 ;
  assign n365 = ( x48 & x49 ) | ( x48 & ~n364 ) | ( x49 & ~n364 ) ;
  assign n366 = x48 | x49 ;
  assign n367 = ~n362 & n366 ;
  assign n368 = ( x45 & x46 ) | ( x45 & n345 ) | ( x46 & n345 ) ;
  assign n369 = ~n367 & n368 ;
  assign n370 = ( ~n362 & n365 ) | ( ~n362 & n369 ) | ( n365 & n369 ) ;
  assign n371 = ( x47 & n349 ) | ( x47 & n354 ) | ( n349 & n354 ) ;
  assign n372 = ( x50 & n370 ) | ( x50 & ~n371 ) | ( n370 & ~n371 ) ;
  assign n373 = ( ~x50 & n371 ) | ( ~x50 & n372 ) | ( n371 & n372 ) ;
  assign n374 = ( ~n370 & n372 ) | ( ~n370 & n373 ) | ( n372 & n373 ) ;
  assign n375 = x51 & x52 ;
  assign n376 = x51 | x52 ;
  assign n377 = ~n375 & n376 ;
  assign n378 = ( x48 & x49 ) | ( x48 & n364 ) | ( x49 & n364 ) ;
  assign n379 = n377 & ~n378 ;
  assign n380 = n367 & n368 ;
  assign n381 = ( n362 & ~n377 ) | ( n362 & n380 ) | ( ~n377 & n380 ) ;
  assign n382 = n379 | n381 ;
  assign n383 = x53 & n382 ;
  assign n384 = x50 | n370 ;
  assign n385 = x50 & n370 ;
  assign n386 = n371 | n385 ;
  assign n387 = n384 & n386 ;
  assign n388 = ( x53 & n382 ) | ( x53 & ~n387 ) | ( n382 & ~n387 ) ;
  assign n389 = x53 | n382 ;
  assign n390 = ~n383 & n389 ;
  assign n391 = n384 & ~n385 ;
  assign n392 = n371 & n391 ;
  assign n393 = ( n385 & ~n390 ) | ( n385 & n392 ) | ( ~n390 & n392 ) ;
  assign n394 = ( ~n383 & n388 ) | ( ~n383 & n393 ) | ( n388 & n393 ) ;
  assign n395 = x54 & x55 ;
  assign n396 = n375 | n378 ;
  assign n397 = n376 & n396 ;
  assign n398 = ( x54 & x55 ) | ( x54 & ~n397 ) | ( x55 & ~n397 ) ;
  assign n399 = x54 | x55 ;
  assign n400 = ~n395 & n399 ;
  assign n401 = ( x51 & x52 ) | ( x51 & n378 ) | ( x52 & n378 ) ;
  assign n402 = ~n400 & n401 ;
  assign n403 = ( ~n395 & n398 ) | ( ~n395 & n402 ) | ( n398 & n402 ) ;
  assign n404 = ( x53 & n382 ) | ( x53 & n387 ) | ( n382 & n387 ) ;
  assign n405 = ( x56 & n403 ) | ( x56 & ~n404 ) | ( n403 & ~n404 ) ;
  assign n406 = ( ~x56 & n404 ) | ( ~x56 & n405 ) | ( n404 & n405 ) ;
  assign n407 = ( ~n403 & n405 ) | ( ~n403 & n406 ) | ( n405 & n406 ) ;
  assign n408 = x57 & x58 ;
  assign n409 = x57 | x58 ;
  assign n410 = ~n408 & n409 ;
  assign n411 = ( x54 & x55 ) | ( x54 & n397 ) | ( x55 & n397 ) ;
  assign n412 = n410 & ~n411 ;
  assign n413 = n400 & n401 ;
  assign n414 = ( n395 & ~n410 ) | ( n395 & n413 ) | ( ~n410 & n413 ) ;
  assign n415 = n412 | n414 ;
  assign n416 = x59 & n415 ;
  assign n417 = x56 | n403 ;
  assign n418 = x56 & n403 ;
  assign n419 = n404 | n418 ;
  assign n420 = n417 & n419 ;
  assign n421 = ( x59 & n415 ) | ( x59 & ~n420 ) | ( n415 & ~n420 ) ;
  assign n422 = x59 | n415 ;
  assign n423 = ~n416 & n422 ;
  assign n424 = n417 & ~n418 ;
  assign n425 = n404 & n424 ;
  assign n426 = ( n418 & ~n423 ) | ( n418 & n425 ) | ( ~n423 & n425 ) ;
  assign n427 = ( ~n416 & n421 ) | ( ~n416 & n426 ) | ( n421 & n426 ) ;
  assign n428 = x60 & x61 ;
  assign n429 = n408 | n411 ;
  assign n430 = n409 & n429 ;
  assign n431 = ( x60 & x61 ) | ( x60 & ~n430 ) | ( x61 & ~n430 ) ;
  assign n432 = x60 | x61 ;
  assign n433 = ~n428 & n432 ;
  assign n434 = ( x57 & x58 ) | ( x57 & n411 ) | ( x58 & n411 ) ;
  assign n435 = ~n433 & n434 ;
  assign n436 = ( ~n428 & n431 ) | ( ~n428 & n435 ) | ( n431 & n435 ) ;
  assign n437 = ( x59 & n415 ) | ( x59 & n420 ) | ( n415 & n420 ) ;
  assign n438 = ( x62 & n436 ) | ( x62 & ~n437 ) | ( n436 & ~n437 ) ;
  assign n439 = ( ~x62 & n437 ) | ( ~x62 & n438 ) | ( n437 & n438 ) ;
  assign n440 = ( ~n436 & n438 ) | ( ~n436 & n439 ) | ( n438 & n439 ) ;
  assign n441 = x63 & x64 ;
  assign n442 = x63 | x64 ;
  assign n443 = ~n441 & n442 ;
  assign n444 = ( x60 & x61 ) | ( x60 & n430 ) | ( x61 & n430 ) ;
  assign n445 = n443 & ~n444 ;
  assign n446 = n433 & n434 ;
  assign n447 = ( n428 & ~n443 ) | ( n428 & n446 ) | ( ~n443 & n446 ) ;
  assign n448 = n445 | n447 ;
  assign n449 = x65 & n448 ;
  assign n450 = x62 | n436 ;
  assign n451 = x62 & n436 ;
  assign n452 = n437 | n451 ;
  assign n453 = n450 & n452 ;
  assign n454 = ( x65 & n448 ) | ( x65 & ~n453 ) | ( n448 & ~n453 ) ;
  assign n455 = x65 | n448 ;
  assign n456 = ~n449 & n455 ;
  assign n457 = n450 & ~n451 ;
  assign n458 = n437 & n457 ;
  assign n459 = ( n451 & ~n456 ) | ( n451 & n458 ) | ( ~n456 & n458 ) ;
  assign n460 = ( ~n449 & n454 ) | ( ~n449 & n459 ) | ( n454 & n459 ) ;
  assign n461 = x66 & x67 ;
  assign n462 = n441 | n444 ;
  assign n463 = n442 & n462 ;
  assign n464 = ( x66 & x67 ) | ( x66 & ~n463 ) | ( x67 & ~n463 ) ;
  assign n465 = x66 | x67 ;
  assign n466 = ~n461 & n465 ;
  assign n467 = ( x63 & x64 ) | ( x63 & n444 ) | ( x64 & n444 ) ;
  assign n468 = ~n466 & n467 ;
  assign n469 = ( ~n461 & n464 ) | ( ~n461 & n468 ) | ( n464 & n468 ) ;
  assign n470 = ( x65 & n448 ) | ( x65 & n453 ) | ( n448 & n453 ) ;
  assign n471 = ( x68 & n469 ) | ( x68 & ~n470 ) | ( n469 & ~n470 ) ;
  assign n472 = ( ~x68 & n470 ) | ( ~x68 & n471 ) | ( n470 & n471 ) ;
  assign n473 = ( ~n469 & n471 ) | ( ~n469 & n472 ) | ( n471 & n472 ) ;
  assign n474 = x69 & x70 ;
  assign n475 = x69 | x70 ;
  assign n476 = ~n474 & n475 ;
  assign n477 = ( x66 & x67 ) | ( x66 & n463 ) | ( x67 & n463 ) ;
  assign n478 = n476 & ~n477 ;
  assign n479 = n466 & n467 ;
  assign n480 = ( n461 & ~n476 ) | ( n461 & n479 ) | ( ~n476 & n479 ) ;
  assign n481 = n478 | n480 ;
  assign n482 = x71 & n481 ;
  assign n483 = x68 | n469 ;
  assign n484 = x68 & n469 ;
  assign n485 = n470 | n484 ;
  assign n486 = n483 & n485 ;
  assign n487 = ( x71 & n481 ) | ( x71 & ~n486 ) | ( n481 & ~n486 ) ;
  assign n488 = x71 | n481 ;
  assign n489 = ~n482 & n488 ;
  assign n490 = n483 & ~n484 ;
  assign n491 = n470 & n490 ;
  assign n492 = ( n484 & ~n489 ) | ( n484 & n491 ) | ( ~n489 & n491 ) ;
  assign n493 = ( ~n482 & n487 ) | ( ~n482 & n492 ) | ( n487 & n492 ) ;
  assign n494 = x72 & x73 ;
  assign n495 = n474 | n477 ;
  assign n496 = n475 & n495 ;
  assign n497 = ( x72 & x73 ) | ( x72 & ~n496 ) | ( x73 & ~n496 ) ;
  assign n498 = x72 | x73 ;
  assign n499 = ~n494 & n498 ;
  assign n500 = ( x69 & x70 ) | ( x69 & n477 ) | ( x70 & n477 ) ;
  assign n501 = ~n499 & n500 ;
  assign n502 = ( ~n494 & n497 ) | ( ~n494 & n501 ) | ( n497 & n501 ) ;
  assign n503 = ( x71 & n481 ) | ( x71 & n486 ) | ( n481 & n486 ) ;
  assign n504 = ( x74 & n502 ) | ( x74 & ~n503 ) | ( n502 & ~n503 ) ;
  assign n505 = ( ~x74 & n503 ) | ( ~x74 & n504 ) | ( n503 & n504 ) ;
  assign n506 = ( ~n502 & n504 ) | ( ~n502 & n505 ) | ( n504 & n505 ) ;
  assign n507 = x75 & x76 ;
  assign n508 = x75 | x76 ;
  assign n509 = ~n507 & n508 ;
  assign n510 = ( x72 & x73 ) | ( x72 & n496 ) | ( x73 & n496 ) ;
  assign n511 = n509 & ~n510 ;
  assign n512 = n499 & n500 ;
  assign n513 = ( n494 & ~n509 ) | ( n494 & n512 ) | ( ~n509 & n512 ) ;
  assign n514 = n511 | n513 ;
  assign n515 = x77 & n514 ;
  assign n516 = x74 | n502 ;
  assign n517 = x74 & n502 ;
  assign n518 = n503 | n517 ;
  assign n519 = n516 & n518 ;
  assign n520 = ( x77 & n514 ) | ( x77 & ~n519 ) | ( n514 & ~n519 ) ;
  assign n521 = x77 | n514 ;
  assign n522 = ~n515 & n521 ;
  assign n523 = n516 & ~n517 ;
  assign n524 = n503 & n523 ;
  assign n525 = ( n517 & ~n522 ) | ( n517 & n524 ) | ( ~n522 & n524 ) ;
  assign n526 = ( ~n515 & n520 ) | ( ~n515 & n525 ) | ( n520 & n525 ) ;
  assign n527 = x78 & x79 ;
  assign n528 = n507 | n510 ;
  assign n529 = n508 & n528 ;
  assign n530 = ( x78 & x79 ) | ( x78 & ~n529 ) | ( x79 & ~n529 ) ;
  assign n531 = x78 | x79 ;
  assign n532 = ~n527 & n531 ;
  assign n533 = ( x75 & x76 ) | ( x75 & n510 ) | ( x76 & n510 ) ;
  assign n534 = ~n532 & n533 ;
  assign n535 = ( ~n527 & n530 ) | ( ~n527 & n534 ) | ( n530 & n534 ) ;
  assign n536 = ( x77 & n514 ) | ( x77 & n519 ) | ( n514 & n519 ) ;
  assign n537 = ( x80 & n535 ) | ( x80 & ~n536 ) | ( n535 & ~n536 ) ;
  assign n538 = ( ~x80 & n536 ) | ( ~x80 & n537 ) | ( n536 & n537 ) ;
  assign n539 = ( ~n535 & n537 ) | ( ~n535 & n538 ) | ( n537 & n538 ) ;
  assign n540 = x81 & x82 ;
  assign n541 = x81 | x82 ;
  assign n542 = ~n540 & n541 ;
  assign n543 = ( x78 & x79 ) | ( x78 & n529 ) | ( x79 & n529 ) ;
  assign n544 = n542 & ~n543 ;
  assign n545 = n532 & n533 ;
  assign n546 = ( n527 & ~n542 ) | ( n527 & n545 ) | ( ~n542 & n545 ) ;
  assign n547 = n544 | n546 ;
  assign n548 = x83 & n547 ;
  assign n549 = x80 | n535 ;
  assign n550 = x80 & n535 ;
  assign n551 = n536 | n550 ;
  assign n552 = n549 & n551 ;
  assign n553 = ( x83 & n547 ) | ( x83 & ~n552 ) | ( n547 & ~n552 ) ;
  assign n554 = x83 | n547 ;
  assign n555 = ~n548 & n554 ;
  assign n556 = n549 & ~n550 ;
  assign n557 = n536 & n556 ;
  assign n558 = ( n550 & ~n555 ) | ( n550 & n557 ) | ( ~n555 & n557 ) ;
  assign n559 = ( ~n548 & n553 ) | ( ~n548 & n558 ) | ( n553 & n558 ) ;
  assign n560 = x84 & x85 ;
  assign n561 = n540 | n543 ;
  assign n562 = n541 & n561 ;
  assign n563 = ( x84 & x85 ) | ( x84 & ~n562 ) | ( x85 & ~n562 ) ;
  assign n564 = x84 | x85 ;
  assign n565 = ~n560 & n564 ;
  assign n566 = ( x81 & x82 ) | ( x81 & n543 ) | ( x82 & n543 ) ;
  assign n567 = ~n565 & n566 ;
  assign n568 = ( ~n560 & n563 ) | ( ~n560 & n567 ) | ( n563 & n567 ) ;
  assign n569 = ( x83 & n547 ) | ( x83 & n552 ) | ( n547 & n552 ) ;
  assign n570 = ( x86 & n568 ) | ( x86 & ~n569 ) | ( n568 & ~n569 ) ;
  assign n571 = ( ~x86 & n569 ) | ( ~x86 & n570 ) | ( n569 & n570 ) ;
  assign n572 = ( ~n568 & n570 ) | ( ~n568 & n571 ) | ( n570 & n571 ) ;
  assign n573 = x87 & x88 ;
  assign n574 = x87 | x88 ;
  assign n575 = ~n573 & n574 ;
  assign n576 = ( x84 & x85 ) | ( x84 & n562 ) | ( x85 & n562 ) ;
  assign n577 = n575 & ~n576 ;
  assign n578 = n565 & n566 ;
  assign n579 = ( n560 & ~n575 ) | ( n560 & n578 ) | ( ~n575 & n578 ) ;
  assign n580 = n577 | n579 ;
  assign n581 = x89 & n580 ;
  assign n582 = x86 | n568 ;
  assign n583 = x86 & n568 ;
  assign n584 = n569 | n583 ;
  assign n585 = n582 & n584 ;
  assign n586 = ( x89 & n580 ) | ( x89 & ~n585 ) | ( n580 & ~n585 ) ;
  assign n587 = x89 | n580 ;
  assign n588 = ~n581 & n587 ;
  assign n589 = n582 & ~n583 ;
  assign n590 = n569 & n589 ;
  assign n591 = ( n583 & ~n588 ) | ( n583 & n590 ) | ( ~n588 & n590 ) ;
  assign n592 = ( ~n581 & n586 ) | ( ~n581 & n591 ) | ( n586 & n591 ) ;
  assign n593 = x90 & x91 ;
  assign n594 = n573 | n576 ;
  assign n595 = n574 & n594 ;
  assign n596 = ( x90 & x91 ) | ( x90 & ~n595 ) | ( x91 & ~n595 ) ;
  assign n597 = x90 | x91 ;
  assign n598 = ~n593 & n597 ;
  assign n599 = ( x87 & x88 ) | ( x87 & n576 ) | ( x88 & n576 ) ;
  assign n600 = ~n598 & n599 ;
  assign n601 = ( ~n593 & n596 ) | ( ~n593 & n600 ) | ( n596 & n600 ) ;
  assign n602 = ( x89 & n580 ) | ( x89 & n585 ) | ( n580 & n585 ) ;
  assign n603 = ( x92 & n601 ) | ( x92 & ~n602 ) | ( n601 & ~n602 ) ;
  assign n604 = ( ~x92 & n602 ) | ( ~x92 & n603 ) | ( n602 & n603 ) ;
  assign n605 = ( ~n601 & n603 ) | ( ~n601 & n604 ) | ( n603 & n604 ) ;
  assign n606 = x92 & n601 ;
  assign n607 = x92 | n601 ;
  assign n608 = n602 & n607 ;
  assign n609 = n606 | n608 ;
  assign n610 = n597 & n599 ;
  assign n611 = n593 | n610 ;
  assign n612 = ( x93 & ~x94 ) | ( x93 & n611 ) | ( ~x94 & n611 ) ;
  assign n613 = ( x90 & x91 ) | ( x90 & n595 ) | ( x91 & n595 ) ;
  assign n614 = ( x94 & n612 ) | ( x94 & ~n613 ) | ( n612 & ~n613 ) ;
  assign n615 = ( ~x93 & n612 ) | ( ~x93 & n614 ) | ( n612 & n614 ) ;
  assign n616 = ( x95 & n609 ) | ( x95 & ~n615 ) | ( n609 & ~n615 ) ;
  assign n617 = n602 | n606 ;
  assign n618 = n607 & n617 ;
  assign n619 = ( n615 & n616 ) | ( n615 & ~n618 ) | ( n616 & ~n618 ) ;
  assign n620 = ( ~x95 & n616 ) | ( ~x95 & n619 ) | ( n616 & n619 ) ;
  assign y0 = n99 ;
  assign y1 = n114 ;
  assign y2 = n137 ;
  assign y3 = n159 ;
  assign y4 = n176 ;
  assign y5 = n196 ;
  assign y6 = n209 ;
  assign y7 = n229 ;
  assign y8 = n242 ;
  assign y9 = n262 ;
  assign y10 = n275 ;
  assign y11 = n295 ;
  assign y12 = n308 ;
  assign y13 = n328 ;
  assign y14 = n341 ;
  assign y15 = n361 ;
  assign y16 = n374 ;
  assign y17 = n394 ;
  assign y18 = n407 ;
  assign y19 = n427 ;
  assign y20 = n440 ;
  assign y21 = n460 ;
  assign y22 = n473 ;
  assign y23 = n493 ;
  assign y24 = n506 ;
  assign y25 = n526 ;
  assign y26 = n539 ;
  assign y27 = n559 ;
  assign y28 = n572 ;
  assign y29 = n592 ;
  assign y30 = n605 ;
  assign y31 = n620 ;
endmodule
