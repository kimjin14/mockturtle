//Written by the Majority Logic Package Fri Nov 14 23:11:32 2014
module top (
            cin, a0, b0, b1, a1, b2, a2, b3, a3, b4, a4, b5, a5, b6, a6, b7, a7, b8, a8, b9, a9, b10, a10, b11, a11, b12, a12, b13, a13, b14, a14, b15, a15, b16, a16, b17, a17, b18, a18, b19, a19, b20, a20, b21, a21, b22, a22, b23, a23, b24, a24, b25, a25, b26, a26, b27, a27, b28, a28, b29, a29, b30, a30, b31, a31, b32, a32, b33, a33, b34, a34, b35, a35, b36, a36, b37, a37, b38, a38, b39, a39, b40, a40, b41, a41, b42, a42, b43, a43, b44, a44, b45, a45, b46, a46, b47, a47, b48, a48, b49, a49, b50, a50, b51, a51, b52, a52, b53, a53, b54, a54, b55, a55, b56, a56, b57, a57, b58, a58, b59, a59, b60, a60, b61, a61, b62, a62, b63, a63, b64, a64, b65, a65, b66, a66, b67, a67, b68, a68, b69, a69, b70, a70, b71, a71, b72, a72, b73, a73, b74, a74, b75, a75, b76, a76, b77, a77, b78, a78, b79, a79, b80, a80, b81, a81, b82, a82, b83, a83, b84, a84, b85, a85, b86, a86, b87, a87, b88, a88, b89, a89, b90, a90, b91, a91, b92, a92, b93, a93, b94, a94, b95, a95, b96, a96, b97, a97, b98, a98, b99, a99, b100, a100, b101, a101, b102, a102, b103, a103, b104, a104, b105, a105, b106, a106, b107, a107, b108, a108, b109, a109, b110, a110, b111, a111, b112, a112, b113, a113, b114, a114, b115, a115, b116, a116, b117, a117, b118, a118, b119, a119, b120, a120, b121, a121, b122, a122, b123, a123, b124, a124, b125, a125, b126, a126, a127, b127, 
            s0, s1, s2, s3, s4, s5, s6, s7, s8, s9, s10, s11, s12, s13, s14, s15, s16, s17, s18, s19, s20, s21, s22, s23, s24, s25, s26, s27, s28, s29, s30, s31, s32, s33, s34, s35, s36, s37, s38, s39, s40, s41, s42, s43, s44, s45, s46, s47, s48, s49, s50, s51, s52, s53, s54, s55, s56, s57, s58, s59, s60, s61, s62, s63, s64, s65, s66, s67, s68, s69, s70, s71, s72, s73, s74, s75, s76, s77, s78, s79, s80, s81, s82, s83, s84, s85, s86, s87, s88, s89, s90, s91, s92, s93, s94, s95, s96, s97, s98, s99, s100, s101, s102, s103, s104, s105, s106, s107, s108, s109, s110, s111, s112, s113, s114, s115, s116, s117, s118, s119, s120, s121, s122, s123, s124, s125, s126, s127, s128);
input cin, a0, b0, b1, a1, b2, a2, b3, a3, b4, a4, b5, a5, b6, a6, b7, a7, b8, a8, b9, a9, b10, a10, b11, a11, b12, a12, b13, a13, b14, a14, b15, a15, b16, a16, b17, a17, b18, a18, b19, a19, b20, a20, b21, a21, b22, a22, b23, a23, b24, a24, b25, a25, b26, a26, b27, a27, b28, a28, b29, a29, b30, a30, b31, a31, b32, a32, b33, a33, b34, a34, b35, a35, b36, a36, b37, a37, b38, a38, b39, a39, b40, a40, b41, a41, b42, a42, b43, a43, b44, a44, b45, a45, b46, a46, b47, a47, b48, a48, b49, a49, b50, a50, b51, a51, b52, a52, b53, a53, b54, a54, b55, a55, b56, a56, b57, a57, b58, a58, b59, a59, b60, a60, b61, a61, b62, a62, b63, a63, b64, a64, b65, a65, b66, a66, b67, a67, b68, a68, b69, a69, b70, a70, b71, a71, b72, a72, b73, a73, b74, a74, b75, a75, b76, a76, b77, a77, b78, a78, b79, a79, b80, a80, b81, a81, b82, a82, b83, a83, b84, a84, b85, a85, b86, a86, b87, a87, b88, a88, b89, a89, b90, a90, b91, a91, b92, a92, b93, a93, b94, a94, b95, a95, b96, a96, b97, a97, b98, a98, b99, a99, b100, a100, b101, a101, b102, a102, b103, a103, b104, a104, b105, a105, b106, a106, b107, a107, b108, a108, b109, a109, b110, a110, b111, a111, b112, a112, b113, a113, b114, a114, b115, a115, b116, a116, b117, a117, b118, a118, b119, a119, b120, a120, b121, a121, b122, a122, b123, a123, b124, a124, b125, a125, b126, a126, a127, b127;
output s0, s1, s2, s3, s4, s5, s6, s7, s8, s9, s10, s11, s12, s13, s14, s15, s16, s17, s18, s19, s20, s21, s22, s23, s24, s25, s26, s27, s28, s29, s30, s31, s32, s33, s34, s35, s36, s37, s38, s39, s40, s41, s42, s43, s44, s45, s46, s47, s48, s49, s50, s51, s52, s53, s54, s55, s56, s57, s58, s59, s60, s61, s62, s63, s64, s65, s66, s67, s68, s69, s70, s71, s72, s73, s74, s75, s76, s77, s78, s79, s80, s81, s82, s83, s84, s85, s86, s87, s88, s89, s90, s91, s92, s93, s94, s95, s96, s97, s98, s99, s100, s101, s102, s103, s104, s105, s106, s107, s108, s109, s110, s111, s112, s113, s114, s115, s116, s117, s118, s119, s120, s121, s122, s123, s124, s125, s126, s127, s128;
wire one, w0, w1, w2, w3, w4, w5, w6, w7, w8, w9, w10, w11, w12, w13, w14, w15, w16, w17, w18, w19, w20, w21, w22, w23, w24, w25, w26, w27, w28, w29, w30, w31, w32, w33, w34, w35, w36, w37, w38, w39, w40, w41, w42, w43, w44, w45, w46, w47, w48, w49, w50, w51, w52, w53, w54, w55, w56, w57, w58, w59, w60, w61, w62, w63, w64, w65, w66, w67, w68, w69, w70, w71, w72, w73, w74, w75, w76, w77, w78, w79, w80, w81, w82, w83, w84, w85, w86, w87, w88, w89, w90, w91, w92, w93, w94, w95, w96, w97, w98, w99, w100, w101, w102, w103, w104, w105, w106, w107, w108, w109, w110, w111, w112, w113, w114, w115, w116, w117, w118, w119, w120, w121, w122, w123, w124, w125, w126, w127, w128, w129, w130, w131, w132, w133, w134, w135, w136, w137, w138, w139, w140, w141, w142, w143, w144, w145, w146, w147, w148, w149, w150, w151, w152, w153, w154, w155, w156, w157, w158, w159, w160, w161, w162, w163, w164, w165, w166, w167, w168, w169, w170, w171, w172, w173, w174, w175, w176, w177, w178, w179, w180, w181, w182, w183, w184, w185, w186, w187, w188, w189, w190, w191, w192, w193, w194, w195, w196, w197, w198, w199, w200, w201, w202, w203, w204, w205, w206, w207, w208, w209, w210, w211, w212, w213, w214, w215, w216, w217, w218, w219, w220, w221, w222, w223, w224, w225, w226, w227, w228, w229, w230, w231, w232, w233, w234, w235, w236, w237, w238, w239, w240, w241, w242, w243, w244, w245, w246, w247, w248, w249, w250, w251, w252, w253, w254, w255, w256, w257, w258, w259, w260, w261, w262, w263, w264, w265, w266, w267, w268, w269, w270, w271, w272, w273, w274, w275, w276, w277, w278, w279, w280, w281, w282, w283, w284, w285, w286, w287, w288, w289, w290, w291, w292, w293, w294, w295, w296, w297, w298, w299, w300, w301, w302, w303, w304, w305, w306, w307, w308, w309, w310, w311, w312, w313, w314, w315, w316, w317, w318, w319, w320, w321, w322, w323, w324, w325, w326, w327, w328, w329, w330, w331, w332, w333, w334, w335, w336, w337, w338, w339, w340, w341, w342, w343, w344, w345, w346, w347, w348, w349, w350, w351, w352, w353, w354, w355, w356, w357, w358, w359, w360, w361, w362, w363, w364, w365, w366, w367, w368, w369, w370, w371, w372, w373, w374, w375, w376, w377, w378, w379, w380, w381, w382, w383, w384, w385, w386, w387, w388, w389, w390, w391, w392, w393, w394, w395, w396, w397, w398, w399, w400, w401, w402, w403, w404, w405, w406, w407, w408, w409, w410, w411, w412, w413, w414, w415, w416, w417, w418, w419, w420, w421, w422, w423, w424, w425, w426, w427, w428, w429, w430, w431, w432, w433, w434, w435, w436, w437, w438, w439, w440, w441, w442, w443, w444, w445, w446, w447, w448, w449, w450, w451, w452, w453, w454, w455, w456, w457, w458, w459, w460, w461, w462, w463, w464, w465, w466, w467, w468, w469, w470, w471, w472, w473, w474, w475, w476, w477, w478, w479, w480, w481, w482, w483, w484, w485, w486, w487, w488, w489, w490, w491, w492, w493, w494, w495, w496, w497, w498, w499, w500, w501, w502, w503, w504, w505, w506, w507, w508, w509, w510, w511, w512, w513, w514, w515, w516, w517, w518, w519, w520, w521, w522, w523, w524, w525, w526, w527, w528, w529, w530, w531, w532, w533, w534, w535, w536, w537, w538, w539, w540, w541, w542, w543, w544, w545, w546, w547, w548, w549, w550, w551, w552, w553, w554, w555, w556, w557, w558, w559, w560, w561, w562, w563, w564, w565, w566, w567, w568, w569, w570, w571, w572, w573, w574, w575, w576, w577, w578, w579, w580, w581, w582, w583, w584, w585, w586, w587, w588, w589, w590, w591, w592, w593, w594, w595, w596, w597, w598, w599, w600, w601, w602, w603, w604, w605, w606, w607, w608, w609, w610, w611, w612, w613, w614, w615, w616, w617, w618, w619, w620, w621, w622, w623, w624, w625, w626, w627, w628, w629, w630, w631, w632, w633, w634, w635, w636, w637, w638, w639, w640, w641, w642, w643, w644, w645, w646, w647, w648, w649, w650, w651, w652, w653, w654, w655, w656, w657, w658, w659, w660, w661, w662, w663, w664, w665, w666, w667, w668, w669, w670, w671, w672, w673, w674, w675, w676, w677, w678, w679, w680, w681, w682, w683, w684, w685, w686, w687, w688, w689, w690, w691, w692, w693, w694, w695, w696, w697, w698, w699, w700, w701, w702, w703, w704, w705, w706, w707, w708, w709, w710, w711, w712, w713, w714, w715, w716, w717, w718, w719, w720, w721, w722, w723, w724, w725, w726, w727, w728, w729, w730, w731, w732, w733, w734, w735, w736, w737, w738, w739, w740, w741, w742, w743, w744, w745, w746, w747, w748, w749, w750, w751, w752, w753, w754, w755, w756, w757, w758, w759, w760, w761, w762, w763, w764, w765, w766, w767, w768, w769, w770, w771, w772, w773, w774, w775, w776, w777, w778, w779, w780, w781, w782, w783, w784, w785, w786, w787, w788, w789, w790, w791, w792, w793, w794, w795, w796, w797, w798, w799, w800, w801, w802, w803, w804, w805, w806, w807, w808, w809, w810, w811, w812, w813, w814, w815, w816, w817, w818, w819, w820, w821, w822, w823, w824, w825, w826, w827, w828, w829, w830, w831, w832, w833, w834, w835, w836, w837, w838, w839, w840, w841, w842, w843, w844, w845, w846, w847, w848, w849, w850, w851, w852, w853, w854, w855, w856, w857, w858, w859, w860, w861, w862, w863, w864, w865, w866, w867, w868, w869, w870, w871, w872, w873, w874, w875, w876, w877, w878, w879, w880, w881, w882, w883, w884, w885, w886, w887, w888, w889, w890, w891, w892, w893, w894, w895, w896, w897, w898, w899, w900, w901, w902, w903, w904, w905, w906, w907, w908, w909, w910, w911, w912, w913, w914, w915, w916, w917, w918, w919, w920, w921, w922, w923, w924, w925, w926, w927, w928, w929, w930, w931, w932, w933, w934, w935, w936, w937, w938, w939, w940, w941, w942, w943, w944, w945, w946, w947, w948, w949, w950, w951, w952, w953, w954, w955, w956, w957, w958, w959, w960, w961, w962, w963, w964, w965, w966, w967, w968, w969, w970, w971, w972, w973, w974, w975, w976, w977, w978, w979, w980, w981, w982, w983, w984, w985, w986, w987, w988, w989, w990, w991, w992, w993, w994, w995, w996, w997, w998, w999, w1000, w1001, w1002, w1003, w1004, w1005, w1006, w1007, w1008, w1009, w1010, w1011, w1012, w1013, w1014, w1015, w1016, w1017, w1018, w1019, w1020, w1021, w1022, w1023, w1024, w1025, w1026, w1027, w1028, w1029, w1030, w1031, w1032, w1033, w1034, w1035, w1036, w1037, w1038, w1039, w1040, w1041, w1042, w1043, w1044, w1045, w1046, w1047, w1048, w1049, w1050, w1051, w1052, w1053, w1054, w1055, w1056, w1057, w1058, w1059, w1060, w1061, w1062, w1063, w1064, w1065, w1066, w1067, w1068, w1069, w1070, w1071, w1072, w1073, w1074, w1075, w1076, w1077, w1078, w1079, w1080, w1081, w1082, w1083, w1084, w1085, w1086, w1087, w1088, w1089, w1090, w1091, w1092, w1093, w1094, w1095, w1096, w1097, w1098, w1099, w1100, w1101, w1102, w1103, w1104, w1105, w1106, w1107, w1108, w1109, w1110, w1111, w1112, w1113, w1114, w1115, w1116, w1117, w1118, w1119, w1120, w1121, w1122, w1123, w1124, w1125, w1126, w1127, w1128, w1129, w1130, w1131, w1132, w1133, w1134, w1135, w1136, w1137, w1138, w1139, w1140, w1141, w1142, w1143, w1144, w1145, w1146, w1147, w1148, w1149, w1150, w1151, w1152, w1153, w1154, w1155, w1156, w1157, w1158, w1159, w1160, w1161, w1162, w1163, w1164, w1165, w1166, w1167, w1168, w1169, w1170, w1171, w1172, w1173, w1174, w1175, w1176, w1177, w1178, w1179, w1180, w1181, w1182, w1183, w1184, w1185, w1186, w1187, w1188, w1189, w1190, w1191, w1192, w1193, w1194, w1195, w1196, w1197, w1198, w1199, w1200, w1201, w1202, w1203, w1204, w1205, w1206, w1207, w1208, w1209, w1210, w1211, w1212, w1213, w1214, w1215, w1216, w1217, w1218, w1219, w1220, w1221, w1222, w1223, w1224, w1225, w1226, w1227, w1228, w1229, w1230, w1231, w1232, w1233, w1234, w1235, w1236, w1237, w1238, w1239, w1240, w1241, w1242, w1243, w1244, w1245, w1246, w1247, w1248, w1249, w1250, w1251, w1252, w1253, w1254, w1255, w1256, w1257, w1258, w1259, w1260, w1261, w1262, w1263, w1264, w1265, w1266, w1267, w1268, w1269, w1270, w1271, w1272, w1273, w1274, w1275, w1276, w1277, w1278, w1279, w1280, w1281, w1282, w1283, w1284, w1285, w1286, w1287, w1288, w1289, w1290, w1291, w1292, w1293, w1294, w1295, w1296, w1297, w1298, w1299, w1300, w1301, w1302, w1303, w1304, w1305, w1306, w1307, w1308, w1309, w1310, w1311, w1312, w1313, w1314, w1315, w1316, w1317, w1318, w1319, w1320, w1321, w1322, w1323, w1324, w1325, w1326, w1327, w1328, w1329, w1330, w1331, w1332, w1333, w1334, w1335, w1336, w1337, w1338, w1339, w1340, w1341, w1342, w1343, w1344, w1345, w1346, w1347, w1348, w1349, w1350, w1351, w1352, w1353, w1354, w1355, w1356, w1357, w1358, w1359, w1360, w1361, w1362, w1363, w1364, w1365, w1366, w1367, w1368, w1369, w1370, w1371, w1372, w1373, w1374, w1375, w1376, w1377, w1378, w1379, w1380, w1381, w1382, w1383, w1384, w1385, w1386, w1387, w1388, w1389, w1390, w1391, w1392, w1393, w1394, w1395, w1396, w1397, w1398, w1399, w1400, w1401, w1402, w1403, w1404, w1405, w1406, w1407, w1408, w1409, w1410, w1411, w1412, w1413, w1414, w1415, w1416, w1417, w1418, w1419, w1420, w1421, w1422, w1423, w1424, w1425, w1426, w1427, w1428, w1429, w1430, w1431, w1432, w1433, w1434, w1435, w1436, w1437, w1438, w1439, w1440, w1441, w1442, w1443, w1444, w1445, w1446, w1447, w1448, w1449, w1450, w1451, w1452, w1453, w1454, w1455, w1456, w1457, w1458, w1459, w1460, w1461, w1462, w1463, w1464, w1465, w1466, w1467, w1468, w1469, w1470, w1471, w1472, w1473, w1474, w1475, w1476, w1477, w1478, w1479, w1480, w1481, w1482, w1483, w1484, w1485, w1486, w1487, w1488, w1489, w1490, w1491, w1492, w1493, w1494, w1495, w1496, w1497, w1498, w1499, w1500, w1501, w1502, w1503, w1504, w1505, w1506, w1507, w1508, w1509, w1510, w1511, w1512, w1513, w1514, w1515, w1516, w1517, w1518, w1519, w1520, w1521, w1522, w1523, w1524, w1525, w1526, w1527, w1528, w1529, w1530, w1531, w1532, w1533, w1534, w1535, w1536, w1537, w1538, w1539, w1540, w1541, w1542, w1543, w1544, w1545, w1546, w1547, w1548, w1549, w1550, w1551, w1552, w1553, w1554, w1555, w1556, w1557, w1558, w1559, w1560, w1561, w1562, w1563, w1564, w1565, w1566, w1567, w1568, w1569, w1570, w1571, w1572, w1573, w1574, w1575, w1576, w1577, w1578, w1579, w1580, w1581, w1582, w1583, w1584, w1585, w1586, w1587, w1588, w1589, w1590, w1591, w1592, w1593, w1594, w1595, w1596, w1597, w1598, w1599, w1600, w1601, w1602, w1603, w1604, w1605, w1606, w1607, w1608, w1609, w1610, w1611, w1612, w1613, w1614, w1615, w1616, w1617, w1618, w1619, w1620, w1621, w1622, w1623, w1624, w1625, w1626, w1627, w1628, w1629, w1630, w1631, w1632, w1633, w1634, w1635, w1636, w1637, w1638, w1639, w1640, w1641, w1642, w1643, w1644, w1645, w1646, w1647, w1648, w1649, w1650, w1651, w1652, w1653, w1654, w1655, w1656, w1657, w1658, w1659, w1660, w1661, w1662, w1663, w1664, w1665, w1666, w1667, w1668, w1669, w1670, w1671, w1672, w1673, w1674, w1675, w1676, w1677, w1678, w1679, w1680, w1681, w1682, w1683, w1684, w1685, w1686, w1687, w1688, w1689, w1690, w1691, w1692, w1693, w1694, w1695, w1696, w1697, w1698, w1699, w1700, w1701, w1702, w1703, w1704, w1705, w1706, w1707, w1708, w1709, w1710, w1711, w1712, w1713, w1714, w1715, w1716, w1717, w1718, w1719, w1720, w1721, w1722, w1723, w1724, w1725, w1726, w1727, w1728, w1729, w1730, w1731, w1732, w1733, w1734, w1735, w1736, w1737, w1738, w1739, w1740, w1741, w1742, w1743, w1744, w1745, w1746, w1747, w1748, w1749, w1750, w1751, w1752, w1753, w1754, w1755, w1756, w1757, w1758, w1759, w1760, w1761, w1762, w1763, w1764, w1765, w1766, w1767, w1768, w1769, w1770, w1771, w1772, w1773, w1774, w1775, w1776, w1777, w1778, w1779, w1780, w1781, w1782, w1783, w1784, w1785, w1786, w1787, w1788, w1789, w1790, w1791, w1792, w1793, w1794, w1795, w1796, w1797, w1798, w1799, w1800, w1801, w1802, w1803, w1804, w1805, w1806, w1807, w1808, w1809, w1810, w1811, w1812, w1813, w1814, w1815, w1816, w1817, w1818, w1819, w1820, w1821, w1822, w1823, w1824, w1825, w1826, w1827, w1828, w1829, w1830, w1831, w1832, w1833, w1834, w1835, w1836, w1837, w1838, w1839, w1840, w1841, w1842, w1843, w1844, w1845, w1846, w1847, w1848, w1849, w1850, w1851, w1852, w1853, w1854, w1855, w1856, w1857, w1858, w1859, w1860, w1861, w1862, w1863, w1864, w1865, w1866, w1867, w1868, w1869, w1870, w1871, w1872, w1873, w1874, w1875, w1876, w1877, w1878, w1879, w1880, w1881, w1882, w1883, w1884, w1885, w1886, w1887, w1888, w1889, w1890, w1891, w1892, w1893, w1894, w1895, w1896, w1897, w1898, w1899, w1900, w1901, w1902, w1903, w1904, w1905, w1906, w1907, w1908, w1909, w1910, w1911, w1912, w1913, w1914, w1915, w1916, w1917, w1918, w1919, w1920, w1921, w1922, w1923, w1924, w1925, w1926, w1927, w1928, w1929, w1930, w1931, w1932, w1933, w1934, w1935, w1936, w1937, w1938, w1939, w1940, w1941, w1942, w1943, w1944, w1945, w1946, w1947, w1948, w1949, w1950, w1951, w1952, w1953, w1954, w1955, w1956, w1957, w1958, w1959, w1960, w1961, w1962, w1963, w1964, w1965, w1966, w1967, w1968, w1969, w1970, w1971, w1972, w1973, w1974, w1975, w1976, w1977, w1978, w1979, w1980, w1981, w1982, w1983, w1984, w1985, w1986, w1987, w1988, w1989, w1990, w1991, w1992, w1993, w1994, w1995, w1996, w1997, w1998, w1999, w2000, w2001, w2002, w2003, w2004, w2005, w2006, w2007, w2008, w2009, w2010, w2011, w2012, w2013, w2014, w2015, w2016, w2017, w2018, w2019, w2020, w2021, w2022, w2023, w2024, w2025, w2026, w2027, w2028, w2029, w2030, w2031, w2032, w2033, w2034, w2035, w2036, w2037, w2038, w2039, w2040, w2041, w2042, w2043, w2044, w2045, w2046, w2047, w2048, w2049, w2050, w2051, w2052, w2053, w2054, w2055, w2056, w2057, w2058, w2059, w2060, w2061, w2062, w2063, w2064, w2065, w2066, w2067, w2068, w2069, w2070, w2071, w2072, w2073, w2074, w2075, w2076, w2077, w2078, w2079, w2080, w2081, w2082, w2083, w2084, w2085, w2086, w2087, w2088, w2089, w2090, w2091, w2092, w2093, w2094, w2095, w2096, w2097, w2098, w2099, w2100, w2101, w2102, w2103, w2104, w2105, w2106, w2107, w2108, w2109, w2110, w2111, w2112, w2113, w2114, w2115, w2116, w2117, w2118, w2119, w2120, w2121, w2122, w2123, w2124, w2125, w2126, w2127, w2128, w2129, w2130, w2131, w2132, w2133, w2134, w2135, w2136, w2137, w2138, w2139, w2140, w2141, w2142, w2143, w2144, w2145, w2146, w2147, w2148, w2149, w2150, w2151, w2152, w2153, w2154, w2155, w2156, w2157, w2158, w2159, w2160, w2161, w2162, w2163, w2164, w2165, w2166, w2167, w2168, w2169, w2170, w2171, w2172, w2173, w2174, w2175, w2176, w2177, w2178, w2179, w2180, w2181, w2182, w2183, w2184, w2185, w2186, w2187, w2188, w2189, w2190, w2191, w2192, w2193, w2194, w2195, w2196, w2197, w2198, w2199, w2200, w2201, w2202, w2203, w2204, w2205, w2206, w2207, w2208, w2209, w2210, w2211, w2212, w2213, w2214, w2215, w2216, w2217, w2218, w2219, w2220, w2221, w2222, w2223, w2224, w2225, w2226, w2227, w2228, w2229, w2230, w2231, w2232, w2233, w2234, w2235, w2236, w2237, w2238, w2239, w2240, w2241, w2242, w2243, w2244, w2245, w2246, w2247, w2248, w2249, w2250, w2251, w2252, w2253, w2254, w2255, w2256, w2257, w2258, w2259, w2260, w2261, w2262, w2263, w2264, w2265, w2266, w2267, w2268, w2269, w2270, w2271, w2272, w2273, w2274, w2275, w2276, w2277, w2278, w2279, w2280, w2281, w2282, w2283, w2284, w2285, w2286, w2287, w2288, w2289, w2290, w2291, w2292, w2293, w2294, w2295, w2296, w2297, w2298, w2299, w2300, w2301, w2302, w2303, w2304, w2305, w2306, w2307, w2308, w2309, w2310, w2311, w2312, w2313, w2314, w2315, w2316, w2317, w2318, w2319, w2320, w2321, w2322, w2323, w2324, w2325, w2326, w2327, w2328, w2329, w2330, w2331, w2332, w2333, w2334, w2335, w2336, w2337, w2338, w2339, w2340, w2341, w2342, w2343, w2344, w2345, w2346, w2347, w2348, w2349, w2350, w2351, w2352, w2353, w2354, w2355, w2356, w2357, w2358, w2359, w2360, w2361, w2362, w2363, w2364, w2365, w2366, w2367, w2368, w2369, w2370, w2371, w2372, w2373, w2374, w2375, w2376, w2377, w2378, w2379, w2380, w2381, w2382, w2383, w2384, w2385, w2386, w2387, w2388, w2389, w2390, w2391, w2392, w2393, w2394, w2395, w2396, w2397, w2398, w2399, w2400, w2401, w2402, w2403, w2404, w2405, w2406, w2407, w2408, w2409, w2410, w2411, w2412, w2413, w2414, w2415, w2416, w2417, w2418, w2419, w2420, w2421, w2422, w2423, w2424, w2425, w2426, w2427, w2428, w2429, w2430, w2431, w2432, w2433, w2434, w2435, w2436, w2437, w2438, w2439, w2440, w2441, w2442, w2443, w2444, w2445, w2446, w2447, w2448, w2449, w2450, w2451, w2452, w2453, w2454, w2455, w2456, w2457, w2458, w2459, w2460, w2461, w2462, w2463, w2464, w2465, w2466, w2467, w2468, w2469, w2470, w2471, w2472, w2473, w2474, w2475, w2476, w2477, w2478, w2479, w2480, w2481, w2482, w2483, w2484, w2485, w2486, w2487, w2488, w2489, w2490, w2491, w2492, w2493, w2494, w2495, w2496, w2497, w2498, w2499, w2500, w2501, w2502, w2503, w2504, w2505, w2506, w2507, w2508, w2509, w2510, w2511, w2512, w2513, w2514, w2515, w2516, w2517, w2518, w2519, w2520, w2521, w2522, w2523, w2524, w2525, w2526, w2527, w2528, w2529, w2530, w2531, w2532, w2533, w2534, w2535, w2536, w2537, w2538, w2539, w2540, w2541, w2542, w2543, w2544, w2545, w2546, w2547, w2548, w2549, w2550, w2551, w2552, w2553, w2554, w2555, w2556, w2557, w2558, w2559, w2560, w2561, w2562, w2563, w2564, w2565, w2566, w2567, w2568, w2569, w2570, w2571, w2572, w2573, w2574, w2575, w2576, w2577, w2578, w2579, w2580, w2581, w2582, w2583, w2584, w2585, w2586, w2587, w2588, w2589, w2590, w2591, w2592, w2593, w2594, w2595, w2596, w2597, w2598, w2599, w2600, w2601, w2602, w2603, w2604, w2605, w2606, w2607, w2608, w2609, w2610, w2611, w2612, w2613, w2614, w2615, w2616, w2617, w2618, w2619, w2620, w2621, w2622, w2623, w2624, w2625, w2626, w2627, w2628, w2629, w2630, w2631, w2632, w2633, w2634, w2635, w2636, w2637, w2638, w2639, w2640, w2641, w2642, w2643, w2644, w2645, w2646, w2647, w2648, w2649, w2650, w2651, w2652, w2653, w2654, w2655, w2656, w2657, w2658, w2659, w2660, w2661, w2662, w2663, w2664, w2665, w2666, w2667, w2668, w2669, w2670, w2671, w2672, w2673, w2674, w2675, w2676, w2677, w2678, w2679, w2680, w2681, w2682, w2683, w2684, w2685, w2686, w2687, w2688, w2689, w2690, w2691, w2692, w2693, w2694, w2695, w2696, w2697, w2698, w2699, w2700, w2701, w2702, w2703, w2704, w2705, w2706, w2707, w2708, w2709, w2710, w2711, w2712, w2713, w2714, w2715, w2716, w2717, w2718, w2719, w2720, w2721, w2722, w2723, w2724, w2725, w2726, w2727, w2728, w2729, w2730, w2731, w2732, w2733, w2734, w2735, w2736, w2737, w2738, w2739, w2740, w2741, w2742, w2743, w2744, w2745, w2746, w2747, w2748, w2749, w2750, w2751, w2752, w2753, w2754, w2755, w2756, w2757, w2758, w2759, w2760, w2761, w2762, w2763, w2764, w2765, w2766, w2767, w2768, w2769, w2770, w2771, w2772, w2773, w2774, w2775, w2776, w2777, w2778, w2779, w2780, w2781, w2782, w2783, w2784, w2785, w2786, w2787, w2788, w2789, w2790, w2791, w2792, w2793, w2794, w2795, w2796, w2797, w2798, w2799, w2800, w2801, w2802, w2803, w2804, w2805, w2806, w2807, w2808, w2809, w2810, w2811, w2812, w2813, w2814, w2815, w2816, w2817, w2818, w2819, w2820, w2821, w2822, w2823, w2824, w2825, w2826, w2827, w2828, w2829, w2830, w2831, w2832, w2833, w2834, w2835, w2836, w2837, w2838, w2839, w2840, w2841, w2842, w2843, w2844, w2845, w2846, w2847, w2848, w2849, w2850, w2851, w2852, w2853, w2854, w2855, w2856, w2857, w2858, w2859, w2860, w2861, w2862, w2863, w2864, w2865, w2866, w2867, w2868, w2869, w2870, w2871, w2872, w2873, w2874, w2875, w2876, w2877, w2878, w2879, w2880, w2881, w2882, w2883, w2884, w2885, w2886, w2887, w2888, w2889, w2890, w2891, w2892, w2893, w2894, w2895, w2896, w2897, w2898, w2899, w2900, w2901, w2902, w2903, w2904, w2905, w2906, w2907, w2908, w2909, w2910, w2911, w2912, w2913, w2914, w2915, w2916, w2917, w2918, w2919, w2920, w2921, w2922, w2923, w2924, w2925, w2926, w2927, w2928, w2929, w2930, w2931, w2932, w2933, w2934, w2935, w2936, w2937, w2938, w2939, w2940, w2941, w2942, w2943, w2944, w2945, w2946, w2947, w2948, w2949, w2950, w2951, w2952, w2953, w2954, w2955, w2956, w2957, w2958, w2959, w2960, w2961, w2962, w2963, w2964, w2965, w2966, w2967, w2968, w2969, w2970, w2971, w2972, w2973, w2974, w2975, w2976, w2977, w2978, w2979, w2980, w2981, w2982, w2983, w2984, w2985, w2986, w2987, w2988, w2989, w2990, w2991, w2992, w2993, w2994, w2995, w2996, w2997, w2998, w2999, w3000, w3001, w3002, w3003, w3004, w3005, w3006, w3007, w3008, w3009, w3010, w3011, w3012, w3013, w3014, w3015, w3016, w3017, w3018, w3019, w3020, w3021, w3022, w3023, w3024, w3025, w3026, w3027, w3028, w3029, w3030, w3031, w3032, w3033, w3034, w3035, w3036, w3037, w3038, w3039, w3040, w3041, w3042, w3043, w3044, w3045, w3046, w3047, w3048, w3049, w3050, w3051, w3052, w3053, w3054, w3055, w3056, w3057, w3058, w3059, w3060, w3061, w3062, w3063, w3064, w3065, w3066, w3067, w3068, w3069, w3070, w3071, w3072, w3073, w3074, w3075, w3076, w3077, w3078, w3079, w3080, w3081, w3082, w3083, w3084, w3085, w3086, w3087, w3088, w3089, w3090, w3091, w3092, w3093, w3094, w3095, w3096, w3097, w3098, w3099, w3100, w3101, w3102, w3103, w3104, w3105, w3106, w3107, w3108, w3109, w3110, w3111, w3112, w3113, w3114, w3115, w3116, w3117, w3118, w3119, w3120, w3121, w3122, w3123, w3124, w3125, w3126, w3127, w3128, w3129, w3130, w3131, w3132, w3133, w3134, w3135, w3136, w3137, w3138, w3139, w3140, w3141, w3142, w3143, w3144, w3145, w3146, w3147, w3148, w3149, w3150, w3151, w3152, w3153, w3154, w3155, w3156, w3157, w3158, w3159, w3160, w3161, w3162, w3163, w3164, w3165, w3166, w3167, w3168, w3169, w3170, w3171, w3172, w3173, w3174, w3175, w3176, w3177, w3178, w3179, w3180, w3181, w3182, w3183, w3184, w3185, w3186, w3187, w3188, w3189, w3190, w3191, w3192, w3193, w3194, w3195, w3196, w3197, w3198, w3199, w3200, w3201, w3202, w3203, w3204, w3205, w3206, w3207, w3208, w3209, w3210, w3211, w3212, w3213, w3214, w3215, w3216, w3217, w3218, w3219, w3220, w3221, w3222, w3223, w3224, w3225, w3226, w3227, w3228, w3229, w3230, w3231, w3232, w3233, w3234, w3235, w3236, w3237, w3238, w3239, w3240, w3241, w3242, w3243, w3244, w3245, w3246, w3247, w3248, w3249, w3250, w3251, w3252, w3253, w3254, w3255, w3256, w3257, w3258, w3259, w3260, w3261, w3262, w3263, w3264, w3265, w3266, w3267, w3268, w3269, w3270, w3271, w3272, w3273, w3274, w3275, w3276, w3277, w3278, w3279, w3280, w3281, w3282, w3283, w3284, w3285, w3286, w3287, w3288, w3289, w3290, w3291, w3292, w3293, w3294, w3295, w3296, w3297, w3298, w3299, w3300, w3301, w3302, w3303, w3304, w3305, w3306, w3307, w3308, w3309, w3310, w3311, w3312, w3313, w3314, w3315, w3316, w3317, w3318, w3319, w3320, w3321, w3322, w3323, w3324, w3325, w3326, w3327, w3328, w3329, w3330, w3331, w3332, w3333, w3334, w3335, w3336, w3337, w3338, w3339, w3340, w3341, w3342, w3343, w3344, w3345, w3346, w3347, w3348, w3349, w3350, w3351, w3352, w3353, w3354, w3355, w3356, w3357, w3358, w3359, w3360, w3361, w3362, w3363, w3364, w3365, w3366, w3367, w3368, w3369, w3370, w3371, w3372, w3373, w3374, w3375, w3376, w3377, w3378, w3379, w3380, w3381, w3382, w3383, w3384, w3385, w3386, w3387, w3388, w3389, w3390, w3391, w3392, w3393, w3394, w3395, w3396, w3397, w3398, w3399, w3400, w3401, w3402, w3403, w3404, w3405, w3406, w3407, w3408, w3409, w3410, w3411, w3412, w3413, w3414, w3415, w3416, w3417, w3418, w3419, w3420, w3421, w3422, w3423, w3424, w3425, w3426, w3427, w3428, w3429, w3430, w3431, w3432, w3433, w3434, w3435, w3436, w3437, w3438, w3439, w3440, w3441, w3442, w3443, w3444, w3445, w3446, w3447, w3448, w3449, w3450, w3451, w3452, w3453, w3454, w3455, w3456, w3457, w3458, w3459, w3460, w3461, w3462, w3463, w3464, w3465, w3466, w3467, w3468, w3469, w3470, w3471, w3472, w3473, w3474, w3475, w3476, w3477, w3478, w3479, w3480, w3481, w3482, w3483, w3484, w3485, w3486, w3487, w3488, w3489, w3490, w3491, w3492, w3493, w3494, w3495, w3496, w3497, w3498, w3499, w3500, w3501, w3502, w3503, w3504, w3505, w3506, w3507, w3508, w3509, w3510, w3511, w3512, w3513, w3514, w3515, w3516, w3517, w3518, w3519, w3520, w3521, w3522, w3523, w3524, w3525, w3526, w3527, w3528, w3529, w3530, w3531, w3532, w3533, w3534, w3535, w3536, w3537, w3538, w3539, w3540, w3541, w3542, w3543, w3544, w3545, w3546, w3547, w3548, w3549, w3550, w3551, w3552, w3553, w3554, w3555, w3556, w3557, w3558, w3559, w3560, w3561, w3562, w3563, w3564, w3565, w3566, w3567, w3568, w3569, w3570, w3571, w3572, w3573, w3574, w3575, w3576, w3577, w3578, w3579, w3580, w3581, w3582, w3583, w3584, w3585, w3586, w3587, w3588, w3589, w3590, w3591, w3592, w3593, w3594, w3595, w3596, w3597, w3598, w3599, w3600, w3601, w3602, w3603, w3604, w3605, w3606, w3607, w3608, w3609, w3610, w3611, w3612, w3613, w3614, w3615, w3616, w3617, w3618, w3619, w3620, w3621, w3622, w3623, w3624, w3625, w3626, w3627, w3628, w3629, w3630, w3631, w3632, w3633, w3634, w3635, w3636, w3637, w3638, w3639, w3640, w3641, w3642, w3643, w3644, w3645, w3646, w3647, w3648, w3649, w3650, w3651, w3652, w3653, w3654, w3655, w3656, w3657, w3658, w3659, w3660, w3661, w3662, w3663, w3664, w3665, w3666, w3667, w3668, w3669, w3670, w3671, w3672, w3673, w3674, w3675, w3676, w3677, w3678, w3679, w3680, w3681, w3682, w3683, w3684, w3685, w3686, w3687, w3688, w3689, w3690, w3691, w3692, w3693, w3694, w3695, w3696, w3697, w3698, w3699, w3700, w3701, w3702, w3703, w3704, w3705, w3706, w3707, w3708, w3709, w3710, w3711, w3712, w3713, w3714, w3715, w3716, w3717, w3718, w3719, w3720, w3721, w3722, w3723, w3724, w3725, w3726, w3727, w3728, w3729, w3730, w3731, w3732, w3733, w3734, w3735, w3736, w3737, w3738, w3739, w3740, w3741, w3742, w3743, w3744, w3745, w3746, w3747, w3748, w3749, w3750, w3751, w3752, w3753, w3754, w3755, w3756, w3757, w3758, w3759, w3760, w3761, w3762, w3763, w3764, w3765, w3766, w3767, w3768, w3769, w3770, w3771, w3772, w3773, w3774, w3775, w3776, w3777, w3778, w3779, w3780, w3781, w3782, w3783, w3784, w3785, w3786, w3787, w3788, w3789, w3790, w3791, w3792, w3793, w3794, w3795, w3796, w3797, w3798, w3799, w3800, w3801, w3802, w3803, w3804, w3805, w3806, w3807, w3808, w3809, w3810, w3811, w3812, w3813, w3814, w3815, w3816, w3817, w3818, w3819, w3820, w3821, w3822, w3823, w3824, w3825, w3826, w3827, w3828, w3829, w3830, w3831, w3832, w3833, w3834, w3835, w3836, w3837, w3838, w3839, w3840, w3841, w3842, w3843, w3844, w3845, w3846, w3847, w3848, w3849, w3850, w3851, w3852, w3853, w3854, w3855, w3856, w3857, w3858, w3859, w3860, w3861, w3862, w3863, w3864, w3865, w3866, w3867, w3868, w3869, w3870, w3871, w3872, w3873, w3874, w3875, w3876, w3877, w3878, w3879, w3880, w3881, w3882, w3883, w3884, w3885, w3886, w3887, w3888, w3889, w3890, w3891, w3892, w3893, w3894, w3895, w3896, w3897, w3898, w3899, w3900, w3901, w3902, w3903, w3904, w3905, w3906, w3907, w3908, w3909, w3910, w3911, w3912, w3913, w3914, w3915, w3916, w3917, w3918, w3919, w3920, w3921, w3922, w3923, w3924, w3925, w3926, w3927, w3928, w3929, w3930, w3931, w3932, w3933, w3934, w3935, w3936, w3937, w3938, w3939, w3940, w3941, w3942, w3943, w3944, w3945, w3946, w3947, w3948, w3949, w3950, w3951, w3952, w3953, w3954, w3955, w3956, w3957, w3958, w3959, w3960, w3961, w3962, w3963, w3964, w3965, w3966, w3967, w3968, w3969, w3970, w3971, w3972, w3973, w3974, w3975, w3976, w3977, w3978, w3979, w3980, w3981, w3982, w3983, w3984, w3985, w3986, w3987, w3988, w3989, w3990, w3991, w3992, w3993, w3994, w3995, w3996, w3997, w3998, w3999, w4000, w4001, w4002, w4003, w4004, w4005, w4006, w4007, w4008, w4009, w4010, w4011, w4012, w4013, w4014, w4015, w4016, w4017, w4018, w4019, w4020, w4021, w4022, w4023, w4024, w4025, w4026, w4027, w4028, w4029, w4030, w4031, w4032, w4033, w4034, w4035, w4036, w4037, w4038, w4039, w4040, w4041, w4042, w4043, w4044, w4045, w4046, w4047, w4048, w4049, w4050, w4051, w4052, w4053, w4054, w4055, w4056, w4057, w4058, w4059, w4060, w4061, w4062, w4063, w4064, w4065, w4066, w4067, w4068, w4069, w4070, w4071, w4072, w4073, w4074, w4075, w4076, w4077, w4078, w4079, w4080, w4081, w4082, w4083, w4084, w4085, w4086, w4087, w4088, w4089, w4090, w4091, w4092, w4093, w4094, w4095, w4096, w4097, w4098, w4099, w4100, w4101, w4102, w4103, w4104, w4105, w4106, w4107, w4108, w4109, w4110, w4111, w4112, w4113, w4114, w4115, w4116, w4117, w4118, w4119, w4120, w4121, w4122, w4123, w4124, w4125, w4126, w4127, w4128, w4129, w4130, w4131, w4132, w4133, w4134, w4135, w4136, w4137, w4138, w4139, w4140, w4141, w4142, w4143, w4144, w4145, w4146, w4147, w4148, w4149, w4150, w4151, w4152, w4153, w4154, w4155, w4156, w4157, w4158, w4159, w4160, w4161, w4162, w4163, w4164, w4165, w4166, w4167, w4168, w4169, w4170, w4171, w4172, w4173, w4174, w4175, w4176, w4177, w4178, w4179, w4180, w4181, w4182, w4183, w4184, w4185, w4186, w4187, w4188, w4189, w4190, w4191, w4192, w4193, w4194, w4195, w4196, w4197, w4198, w4199, w4200, w4201, w4202, w4203, w4204, w4205, w4206, w4207, w4208, w4209, w4210, w4211, w4212, w4213, w4214, w4215, w4216, w4217, w4218, w4219, w4220, w4221, w4222, w4223, w4224, w4225, w4226, w4227, w4228, w4229, w4230, w4231, w4232, w4233, w4234, w4235, w4236, w4237, w4238, w4239, w4240, w4241, w4242, w4243, w4244, w4245, w4246, w4247, w4248, w4249, w4250, w4251, w4252, w4253, w4254, w4255, w4256, w4257, w4258, w4259, w4260, w4261, w4262, w4263, w4264, w4265, w4266, w4267, w4268, w4269, w4270, w4271, w4272, w4273, w4274, w4275, w4276, w4277, w4278, w4279, w4280, w4281, w4282, w4283, w4284, w4285, w4286, w4287, w4288, w4289, w4290, w4291, w4292, w4293, w4294, w4295, w4296, w4297, w4298, w4299, w4300, w4301, w4302, w4303, w4304, w4305, w4306, w4307, w4308, w4309, w4310, w4311, w4312, w4313, w4314, w4315, w4316, w4317, w4318, w4319, w4320, w4321, w4322, w4323, w4324, w4325, w4326, w4327, w4328, w4329, w4330, w4331, w4332, w4333, w4334, w4335, w4336, w4337, w4338, w4339, w4340, w4341, w4342, w4343, w4344, w4345, w4346, w4347, w4348, w4349, w4350, w4351, w4352, w4353, w4354, w4355, w4356, w4357, w4358, w4359, w4360, w4361, w4362, w4363, w4364, w4365, w4366, w4367, w4368, w4369, w4370, w4371, w4372, w4373, w4374, w4375, w4376, w4377, w4378, w4379, w4380, w4381, w4382, w4383, w4384, w4385, w4386, w4387, w4388, w4389, w4390, w4391, w4392, w4393, w4394, w4395, w4396, w4397, w4398, w4399, w4400, w4401, w4402, w4403, w4404, w4405, w4406, w4407, w4408, w4409, w4410, w4411, w4412, w4413, w4414, w4415, w4416, w4417, w4418, w4419, w4420, w4421, w4422, w4423, w4424, w4425, w4426, w4427, w4428, w4429, w4430, w4431, w4432, w4433, w4434, w4435, w4436, w4437, w4438, w4439, w4440, w4441, w4442, w4443, w4444, w4445, w4446, w4447, w4448, w4449, w4450, w4451, w4452, w4453, w4454, w4455, w4456, w4457, w4458, w4459, w4460, w4461, w4462, w4463, w4464, w4465, w4466, w4467, w4468, w4469, w4470, w4471, w4472, w4473, w4474, w4475, w4476, w4477, w4478, w4479, w4480, w4481, w4482, w4483, w4484, w4485, w4486, w4487, w4488, w4489, w4490, w4491, w4492, w4493, w4494, w4495, w4496, w4497, w4498, w4499, w4500, w4501, w4502, w4503, w4504, w4505, w4506, w4507, w4508, w4509, w4510, w4511, w4512, w4513, w4514, w4515, w4516, w4517, w4518, w4519, w4520, w4521, w4522, w4523, w4524, w4525, w4526, w4527, w4528, w4529, w4530, w4531, w4532, w4533, w4534, w4535, w4536, w4537, w4538, w4539, w4540, w4541, w4542, w4543, w4544, w4545, w4546, w4547, w4548, w4549, w4550, w4551, w4552, w4553, w4554, w4555, w4556, w4557, w4558, w4559, w4560, w4561, w4562, w4563, w4564, w4565, w4566, w4567, w4568, w4569, w4570, w4571, w4572, w4573, w4574, w4575, w4576, w4577, w4578, w4579, w4580, w4581, w4582, w4583, w4584, w4585, w4586, w4587, w4588, w4589, w4590, w4591, w4592, w4593, w4594, w4595, w4596, w4597, w4598, w4599, w4600, w4601, w4602, w4603, w4604, w4605, w4606, w4607, w4608, w4609, w4610, w4611, w4612, w4613, w4614, w4615, w4616, w4617, w4618, w4619, w4620, w4621, w4622, w4623, w4624, w4625, w4626, w4627, w4628, w4629, w4630, w4631, w4632, w4633, w4634, w4635, w4636, w4637, w4638, w4639, w4640, w4641, w4642, w4643, w4644, w4645, w4646, w4647, w4648, w4649, w4650, w4651, w4652, w4653, w4654, w4655, w4656, w4657, w4658, w4659, w4660, w4661, w4662, w4663, w4664, w4665, w4666, w4667, w4668, w4669, w4670, w4671, w4672, w4673, w4674, w4675, w4676, w4677, w4678, w4679, w4680, w4681, w4682, w4683, w4684, w4685, w4686, w4687, w4688, w4689, w4690, w4691, w4692, w4693, w4694, w4695, w4696, w4697, w4698, w4699, w4700, w4701, w4702, w4703, w4704, w4705, w4706, w4707, w4708, w4709, w4710, w4711, w4712, w4713, w4714, w4715, w4716, w4717, w4718, w4719, w4720, w4721, w4722, w4723, w4724, w4725, w4726, w4727, w4728, w4729, w4730, w4731, w4732, w4733, w4734, w4735, w4736, w4737, w4738, w4739, w4740, w4741, w4742, w4743, w4744, w4745, w4746, w4747, w4748, w4749, w4750, w4751, w4752, w4753, w4754, w4755, w4756, w4757, w4758, w4759, w4760, w4761, w4762, w4763, w4764, w4765, w4766, w4767, w4768, w4769, w4770, w4771, w4772, w4773, w4774, w4775, w4776, w4777, w4778, w4779, w4780, w4781, w4782, w4783, w4784, w4785, w4786, w4787, w4788, w4789, w4790, w4791, w4792, w4793, w4794, w4795, w4796, w4797, w4798, w4799, w4800, w4801, w4802, w4803, w4804, w4805, w4806, w4807, w4808, w4809, w4810, w4811, w4812, w4813, w4814, w4815, w4816, w4817, w4818, w4819, w4820, w4821, w4822, w4823, w4824, w4825, w4826, w4827, w4828, w4829, w4830, w4831, w4832, w4833, w4834, w4835, w4836, w4837, w4838, w4839, w4840, w4841, w4842, w4843, w4844, w4845, w4846, w4847, w4848, w4849, w4850, w4851, w4852, w4853, w4854, w4855, w4856, w4857, w4858, w4859, w4860, w4861, w4862, w4863, w4864, w4865, w4866, w4867, w4868, w4869, w4870, w4871, w4872, w4873, w4874, w4875, w4876, w4877, w4878, w4879, w4880, w4881, w4882, w4883, w4884, w4885, w4886, w4887, w4888, w4889, w4890, w4891, w4892, w4893, w4894, w4895, w4896, w4897, w4898, w4899, w4900, w4901, w4902, w4903, w4904, w4905, w4906, w4907, w4908, w4909, w4910, w4911, w4912, w4913, w4914, w4915, w4916, w4917, w4918, w4919, w4920, w4921, w4922, w4923, w4924, w4925, w4926, w4927, w4928, w4929, w4930, w4931, w4932, w4933, w4934, w4935, w4936, w4937, w4938, w4939, w4940, w4941, w4942, w4943, w4944, w4945, w4946, w4947, w4948, w4949, w4950, w4951, w4952, w4953, w4954, w4955, w4956, w4957, w4958, w4959, w4960, w4961, w4962, w4963, w4964, w4965, w4966, w4967, w4968, w4969, w4970, w4971, w4972, w4973, w4974, w4975, w4976, w4977, w4978, w4979, w4980, w4981, w4982, w4983, w4984, w4985, w4986, w4987, w4988, w4989, w4990, w4991, w4992, w4993, w4994, w4995, w4996, w4997, w4998, w4999, w5000, w5001, w5002, w5003, w5004, w5005, w5006, w5007, w5008, w5009, w5010, w5011, w5012, w5013, w5014, w5015, w5016, w5017, w5018, w5019, w5020, w5021, w5022, w5023, w5024, w5025, w5026, w5027, w5028, w5029, w5030, w5031, w5032, w5033, w5034, w5035, w5036, w5037, w5038, w5039, w5040, w5041, w5042, w5043, w5044, w5045, w5046, w5047, w5048, w5049, w5050, w5051, w5052, w5053, w5054, w5055, w5056, w5057, w5058, w5059, w5060, w5061, w5062, w5063, w5064, w5065, w5066, w5067, w5068, w5069, w5070, w5071, w5072, w5073, w5074, w5075, w5076, w5077, w5078, w5079, w5080, w5081, w5082, w5083, w5084, w5085, w5086, w5087, w5088, w5089, w5090, w5091, w5092, w5093, w5094, w5095, w5096, w5097, w5098, w5099, w5100, w5101, w5102, w5103, w5104, w5105, w5106, w5107, w5108, w5109, w5110, w5111, w5112, w5113, w5114, w5115, w5116, w5117, w5118, w5119, w5120, w5121, w5122, w5123, w5124, w5125, w5126, w5127, w5128, w5129, w5130, w5131, w5132, w5133, w5134, w5135, w5136, w5137, w5138, w5139, w5140, w5141, w5142, w5143, w5144, w5145, w5146, w5147, w5148, w5149, w5150, w5151, w5152, w5153, w5154, w5155, w5156, w5157, w5158, w5159, w5160, w5161, w5162, w5163, w5164, w5165, w5166, w5167, w5168, w5169, w5170, w5171, w5172, w5173, w5174, w5175, w5176, w5177, w5178, w5179, w5180, w5181, w5182, w5183, w5184, w5185, w5186, w5187, w5188, w5189, w5190, w5191, w5192, w5193, w5194, w5195, w5196, w5197, w5198, w5199, w5200, w5201, w5202, w5203, w5204, w5205, w5206, w5207, w5208, w5209, w5210, w5211, w5212, w5213, w5214, w5215, w5216, w5217, w5218, w5219, w5220, w5221, w5222, w5223, w5224, w5225, w5226, w5227, w5228, w5229, w5230, w5231, w5232, w5233, w5234, w5235, w5236, w5237, w5238, w5239, w5240, w5241, w5242, w5243, w5244, w5245, w5246, w5247, w5248, w5249, w5250, w5251, w5252, w5253, w5254, w5255, w5256, w5257, w5258, w5259, w5260, w5261, w5262, w5263, w5264, w5265, w5266, w5267, w5268, w5269, w5270, w5271, w5272, w5273, w5274, w5275, w5276, w5277, w5278, w5279, w5280, w5281, w5282, w5283, w5284, w5285, w5286, w5287, w5288, w5289, w5290, w5291, w5292, w5293, w5294, w5295, w5296, w5297, w5298, w5299, w5300, w5301, w5302, w5303, w5304, w5305, w5306, w5307, w5308, w5309, w5310, w5311, w5312, w5313, w5314, w5315, w5316, w5317, w5318, w5319, w5320, w5321, w5322, w5323, w5324, w5325, w5326, w5327, w5328, w5329, w5330, w5331, w5332, w5333, w5334, w5335, w5336, w5337, w5338, w5339, w5340, w5341, w5342, w5343, w5344, w5345, w5346, w5347, w5348, w5349, w5350, w5351, w5352, w5353, w5354, w5355, w5356, w5357, w5358, w5359, w5360, w5361, w5362, w5363, w5364, w5365, w5366, w5367, w5368, w5369, w5370, w5371, w5372, w5373, w5374, w5375, w5376, w5377, w5378, w5379, w5380, w5381, w5382, w5383, w5384, w5385, w5386, w5387, w5388, w5389, w5390, w5391, w5392, w5393, w5394, w5395, w5396, w5397, w5398, w5399, w5400, w5401, w5402, w5403, w5404, w5405, w5406, w5407, w5408, w5409, w5410, w5411, w5412, w5413, w5414, w5415, w5416, w5417, w5418, w5419, w5420, w5421, w5422, w5423, w5424, w5425, w5426, w5427, w5428, w5429, w5430, w5431, w5432, w5433, w5434, w5435, w5436, w5437, w5438, w5439, w5440, w5441, w5442, w5443, w5444, w5445, w5446, w5447, w5448, w5449, w5450, w5451, w5452, w5453, w5454, w5455, w5456, w5457, w5458, w5459, w5460, w5461, w5462, w5463, w5464, w5465, w5466, w5467, w5468, w5469, w5470, w5471, w5472, w5473, w5474, w5475, w5476, w5477, w5478, w5479, w5480, w5481, w5482, w5483, w5484, w5485, w5486, w5487, w5488, w5489, w5490, w5491, w5492, w5493, w5494, w5495, w5496, w5497, w5498, w5499, w5500, w5501, w5502, w5503, w5504, w5505, w5506, w5507, w5508, w5509, w5510, w5511, w5512, w5513, w5514, w5515, w5516, w5517, w5518, w5519, w5520, w5521, w5522, w5523, w5524, w5525, w5526, w5527, w5528, w5529, w5530, w5531, w5532, w5533, w5534, w5535, w5536, w5537, w5538, w5539, w5540, w5541, w5542, w5543, w5544, w5545, w5546, w5547, w5548, w5549, w5550, w5551, w5552, w5553, w5554, w5555, w5556, w5557, w5558, w5559, w5560, w5561, w5562, w5563, w5564, w5565, w5566, w5567, w5568, w5569, w5570, w5571, w5572, w5573, w5574, w5575, w5576, w5577, w5578, w5579, w5580, w5581, w5582, w5583, w5584, w5585, w5586, w5587, w5588, w5589, w5590, w5591, w5592, w5593, w5594, w5595, w5596, w5597, w5598, w5599, w5600, w5601, w5602, w5603, w5604, w5605, w5606, w5607, w5608, w5609, w5610, w5611, w5612, w5613, w5614, w5615, w5616, w5617, w5618, w5619, w5620, w5621, w5622, w5623, w5624, w5625, w5626, w5627, w5628, w5629, w5630, w5631, w5632, w5633, w5634, w5635, w5636, w5637, w5638, w5639, w5640, w5641, w5642, w5643, w5644, w5645, w5646, w5647, w5648, w5649, w5650, w5651, w5652, w5653, w5654, w5655, w5656, w5657, w5658, w5659, w5660, w5661, w5662, w5663, w5664, w5665, w5666, w5667, w5668, w5669, w5670, w5671, w5672, w5673, w5674, w5675, w5676, w5677, w5678, w5679, w5680, w5681, w5682, w5683, w5684, w5685, w5686, w5687, w5688, w5689, w5690, w5691, w5692, w5693, w5694, w5695, w5696, w5697, w5698, w5699, w5700, w5701, w5702, w5703, w5704, w5705, w5706, w5707, w5708, w5709, w5710, w5711, w5712, w5713, w5714, w5715, w5716, w5717, w5718, w5719, w5720, w5721, w5722, w5723, w5724, w5725, w5726, w5727, w5728, w5729, w5730, w5731, w5732, w5733, w5734, w5735, w5736, w5737, w5738, w5739, w5740, w5741, w5742, w5743, w5744, w5745, w5746, w5747, w5748, w5749, w5750, w5751, w5752, w5753, w5754, w5755, w5756, w5757, w5758, w5759, w5760, w5761, w5762, w5763, w5764, w5765, w5766, w5767, w5768, w5769, w5770, w5771, w5772, w5773, w5774, w5775, w5776, w5777, w5778, w5779, w5780, w5781, w5782, w5783, w5784, w5785, w5786, w5787, w5788, w5789, w5790, w5791, w5792, w5793, w5794, w5795, w5796, w5797, w5798, w5799, w5800, w5801, w5802, w5803, w5804, w5805, w5806, w5807, w5808, w5809, w5810, w5811, w5812, w5813, w5814, w5815, w5816, w5817, w5818, w5819, w5820, w5821, w5822, w5823, w5824, w5825, w5826, w5827, w5828, w5829, w5830, w5831, w5832, w5833, w5834, w5835, w5836, w5837, w5838, w5839, w5840, w5841, w5842, w5843, w5844, w5845, w5846, w5847, w5848, w5849, w5850, w5851, w5852, w5853, w5854, w5855, w5856, w5857, w5858, w5859, w5860, w5861, w5862, w5863, w5864, w5865, w5866, w5867, w5868, w5869, w5870, w5871, w5872, w5873, w5874, w5875, w5876, w5877, w5878, w5879, w5880, w5881, w5882, w5883, w5884, w5885, w5886, w5887, w5888, w5889, w5890, w5891, w5892, w5893, w5894, w5895, w5896, w5897, w5898, w5899, w5900, w5901, w5902, w5903, w5904, w5905, w5906, w5907, w5908, w5909, w5910, w5911, w5912, w5913, w5914, w5915, w5916, w5917, w5918, w5919, w5920, w5921, w5922, w5923, w5924, w5925, w5926, w5927, w5928, w5929, w5930, w5931, w5932, w5933, w5934, w5935, w5936, w5937, w5938, w5939, w5940, w5941, w5942, w5943, w5944, w5945, w5946, w5947, w5948, w5949, w5950, w5951, w5952, w5953, w5954, w5955, w5956, w5957, w5958, w5959, w5960, w5961, w5962, w5963, w5964, w5965, w5966, w5967, w5968, w5969, w5970, w5971, w5972, w5973, w5974, w5975, w5976, w5977, w5978, w5979, w5980, w5981, w5982, w5983, w5984, w5985, w5986, w5987, w5988, w5989, w5990, w5991, w5992, w5993, w5994, w5995, w5996, w5997, w5998, w5999, w6000, w6001, w6002, w6003, w6004, w6005, w6006, w6007, w6008, w6009, w6010, w6011, w6012, w6013, w6014, w6015, w6016, w6017, w6018, w6019, w6020, w6021, w6022, w6023, w6024, w6025, w6026, w6027, w6028, w6029, w6030, w6031, w6032, w6033, w6034, w6035, w6036, w6037, w6038, w6039, w6040, w6041, w6042, w6043, w6044, w6045, w6046, w6047, w6048, w6049, w6050, w6051, w6052, w6053, w6054, w6055, w6056, w6057, w6058, w6059, w6060, w6061, w6062, w6063, w6064, w6065, w6066, w6067, w6068, w6069, w6070, w6071, w6072, w6073, w6074, w6075, w6076, w6077, w6078, w6079, w6080, w6081, w6082, w6083, w6084, w6085, w6086, w6087, w6088, w6089, w6090, w6091, w6092, w6093, w6094, w6095, w6096, w6097, w6098, w6099, w6100, w6101, w6102, w6103, w6104, w6105, w6106, w6107, w6108, w6109, w6110, w6111, w6112, w6113, w6114, w6115, w6116, w6117, w6118, w6119, w6120, w6121, w6122, w6123, w6124, w6125, w6126, w6127, w6128, w6129, w6130, w6131, w6132, w6133, w6134, w6135, w6136, w6137, w6138, w6139, w6140, w6141, w6142, w6143, w6144, w6145, w6146, w6147, w6148, w6149, w6150, w6151, w6152, w6153, w6154, w6155, w6156, w6157, w6158, w6159, w6160, w6161, w6162, w6163, w6164, w6165, w6166, w6167, w6168, w6169, w6170, w6171, w6172, w6173, w6174, w6175, w6176, w6177, w6178, w6179, w6180, w6181, w6182, w6183, w6184, w6185, w6186, w6187, w6188, w6189, w6190, w6191, w6192, w6193, w6194, w6195, w6196, w6197, w6198, w6199, w6200, w6201, w6202, w6203, w6204, w6205, w6206, w6207, w6208, w6209, w6210, w6211, w6212, w6213, w6214, w6215, w6216, w6217, w6218, w6219, w6220, w6221, w6222, w6223, w6224, w6225, w6226, w6227, w6228, w6229, w6230, w6231, w6232, w6233, w6234, w6235, w6236, w6237, w6238, w6239, w6240, w6241, w6242, w6243, w6244, w6245, w6246, w6247, w6248, w6249, w6250, w6251, w6252, w6253, w6254, w6255, w6256, w6257, w6258, w6259, w6260, w6261, w6262, w6263, w6264, w6265, w6266, w6267, w6268, w6269, w6270, w6271, w6272, w6273, w6274, w6275, w6276, w6277, w6278, w6279, w6280, w6281, w6282, w6283, w6284, w6285, w6286, w6287, w6288, w6289, w6290, w6291, w6292, w6293, w6294, w6295, w6296, w6297, w6298, w6299, w6300, w6301, w6302, w6303, w6304, w6305, w6306, w6307, w6308, w6309, w6310, w6311, w6312, w6313, w6314, w6315, w6316, w6317, w6318, w6319, w6320, w6321, w6322, w6323, w6324, w6325, w6326, w6327, w6328, w6329, w6330, w6331, w6332, w6333, w6334, w6335, w6336, w6337, w6338, w6339, w6340, w6341, w6342, w6343, w6344, w6345, w6346, w6347, w6348, w6349, w6350, w6351, w6352, w6353, w6354, w6355, w6356, w6357, w6358, w6359, w6360, w6361, w6362, w6363, w6364, w6365, w6366, w6367, w6368, w6369, w6370, w6371, w6372, w6373, w6374, w6375, w6376, w6377, w6378, w6379, w6380, w6381, w6382, w6383, w6384, w6385, w6386, w6387, w6388, w6389, w6390, w6391, w6392, w6393, w6394, w6395, w6396, w6397, w6398, w6399, w6400, w6401, w6402, w6403, w6404, w6405, w6406, w6407, w6408, w6409, w6410, w6411, w6412, w6413, w6414, w6415, w6416, w6417, w6418, w6419, w6420, w6421, w6422, w6423, w6424, w6425, w6426, w6427, w6428, w6429, w6430, w6431, w6432, w6433, w6434, w6435, w6436, w6437, w6438, w6439, w6440, w6441, w6442, w6443, w6444, w6445, w6446, w6447, w6448, w6449, w6450, w6451, w6452, w6453, w6454, w6455, w6456, w6457, w6458, w6459, w6460, w6461, w6462, w6463, w6464, w6465, w6466, w6467, w6468, w6469, w6470, w6471, w6472, w6473, w6474, w6475, w6476, w6477, w6478, w6479, w6480, w6481, w6482, w6483, w6484, w6485, w6486, w6487, w6488, w6489, w6490, w6491, w6492, w6493, w6494, w6495, w6496, w6497, w6498, w6499, w6500, w6501, w6502, w6503, w6504, w6505, w6506, w6507, w6508, w6509, w6510, w6511, w6512, w6513, w6514, w6515, w6516, w6517, w6518, w6519, w6520, w6521, w6522, w6523, w6524, w6525, w6526, w6527, w6528, w6529, w6530, w6531, w6532, w6533, w6534, w6535, w6536, w6537, w6538, w6539, w6540, w6541, w6542, w6543, w6544, w6545, w6546, w6547, w6548, w6549, w6550, w6551, w6552, w6553, w6554, w6555, w6556, w6557, w6558, w6559, w6560, w6561, w6562, w6563, w6564, w6565, w6566, w6567, w6568, w6569, w6570, w6571, w6572, w6573, w6574, w6575, w6576, w6577, w6578, w6579, w6580, w6581, w6582, w6583, w6584, w6585, w6586, w6587, w6588, w6589, w6590, w6591, w6592, w6593, w6594, w6595, w6596, w6597, w6598, w6599, w6600, w6601, w6602, w6603, w6604, w6605, w6606, w6607, w6608, w6609, w6610, w6611, w6612, w6613, w6614, w6615, w6616, w6617, w6618, w6619, w6620, w6621, w6622, w6623, w6624, w6625, w6626, w6627, w6628, w6629, w6630, w6631, w6632, w6633, w6634, w6635, w6636, w6637, w6638, w6639, w6640, w6641, w6642, w6643, w6644, w6645, w6646, w6647, w6648, w6649, w6650, w6651, w6652, w6653, w6654, w6655, w6656, w6657, w6658, w6659, w6660, w6661, w6662, w6663, w6664, w6665, w6666, w6667, w6668, w6669, w6670, w6671, w6672, w6673, w6674, w6675, w6676, w6677, w6678, w6679, w6680, w6681, w6682, w6683, w6684, w6685, w6686, w6687, w6688, w6689, w6690, w6691, w6692, w6693, w6694, w6695, w6696, w6697, w6698, w6699, w6700, w6701, w6702, w6703, w6704, w6705, w6706, w6707, w6708, w6709, w6710, w6711, w6712, w6713, w6714, w6715, w6716, w6717, w6718, w6719, w6720, w6721, w6722, w6723, w6724, w6725, w6726, w6727, w6728, w6729, w6730, w6731, w6732, w6733, w6734, w6735, w6736, w6737, w6738, w6739, w6740, w6741, w6742, w6743, w6744, w6745, w6746, w6747, w6748, w6749, w6750, w6751, w6752, w6753, w6754, w6755, w6756, w6757, w6758, w6759, w6760, w6761, w6762, w6763, w6764, w6765, w6766, w6767, w6768, w6769, w6770, w6771, w6772, w6773, w6774, w6775, w6776, w6777, w6778, w6779, w6780, w6781, w6782, w6783, w6784, w6785, w6786, w6787, w6788, w6789, w6790, w6791, w6792, w6793, w6794, w6795, w6796, w6797, w6798, w6799, w6800, w6801, w6802, w6803, w6804, w6805, w6806, w6807, w6808, w6809, w6810, w6811, w6812, w6813, w6814, w6815, w6816, w6817, w6818, w6819, w6820, w6821, w6822, w6823, w6824, w6825, w6826, w6827, w6828, w6829, w6830, w6831, w6832, w6833, w6834, w6835, w6836, w6837, w6838, w6839, w6840, w6841, w6842, w6843, w6844, w6845, w6846, w6847, w6848, w6849, w6850, w6851, w6852, w6853, w6854, w6855, w6856, w6857, w6858, w6859, w6860, w6861, w6862, w6863, w6864, w6865, w6866, w6867, w6868, w6869, w6870, w6871, w6872, w6873, w6874, w6875, w6876, w6877, w6878, w6879, w6880, w6881, w6882, w6883, w6884, w6885, w6886, w6887, w6888, w6889, w6890, w6891, w6892, w6893, w6894, w6895, w6896, w6897, w6898, w6899, w6900, w6901, w6902, w6903, w6904, w6905, w6906, w6907, w6908, w6909, w6910, w6911, w6912, w6913, w6914, w6915, w6916, w6917, w6918, w6919, w6920, w6921, w6922, w6923, w6924, w6925, w6926, w6927, w6928, w6929, w6930, w6931, w6932, w6933, w6934, w6935, w6936, w6937, w6938, w6939, w6940, w6941, w6942, w6943, w6944, w6945, w6946, w6947, w6948, w6949, w6950, w6951, w6952, w6953, w6954, w6955, w6956, w6957, w6958, w6959, w6960, w6961, w6962, w6963, w6964, w6965, w6966, w6967, w6968, w6969, w6970, w6971, w6972, w6973, w6974, w6975, w6976, w6977, w6978, w6979, w6980, w6981, w6982, w6983, w6984, w6985, w6986, w6987, w6988, w6989, w6990, w6991, w6992, w6993, w6994, w6995, w6996, w6997, w6998, w6999, w7000, w7001, w7002, w7003, w7004, w7005, w7006, w7007, w7008, w7009, w7010, w7011, w7012, w7013, w7014, w7015, w7016, w7017, w7018, w7019, w7020, w7021, w7022, w7023, w7024, w7025, w7026, w7027, w7028, w7029, w7030, w7031, w7032, w7033, w7034, w7035, w7036, w7037, w7038, w7039, w7040, w7041, w7042, w7043, w7044, w7045, w7046, w7047, w7048, w7049, w7050, w7051, w7052, w7053, w7054, w7055, w7056, w7057, w7058, w7059, w7060, w7061, w7062, w7063, w7064, w7065, w7066, w7067, w7068, w7069, w7070, w7071, w7072, w7073, w7074, w7075, w7076, w7077, w7078, w7079, w7080, w7081, w7082, w7083, w7084, w7085, w7086, w7087, w7088, w7089, w7090, w7091, w7092, w7093, w7094, w7095, w7096, w7097, w7098, w7099, w7100, w7101, w7102, w7103, w7104, w7105, w7106, w7107, w7108, w7109, w7110, w7111, w7112, w7113, w7114, w7115, w7116, w7117, w7118, w7119, w7120, w7121, w7122, w7123, w7124, w7125, w7126, w7127, w7128, w7129, w7130, w7131, w7132, w7133, w7134, w7135, w7136, w7137, w7138, w7139, w7140, w7141, w7142, w7143, w7144, w7145, w7146, w7147, w7148, w7149, w7150, w7151, w7152, w7153, w7154, w7155, w7156, w7157, w7158, w7159, w7160, w7161, w7162, w7163, w7164, w7165, w7166, w7167, w7168, w7169, w7170, w7171, w7172, w7173, w7174, w7175, w7176, w7177, w7178, w7179, w7180, w7181, w7182, w7183, w7184, w7185, w7186, w7187, w7188, w7189, w7190, w7191, w7192, w7193, w7194, w7195, w7196, w7197, w7198, w7199, w7200, w7201, w7202, w7203, w7204, w7205, w7206, w7207, w7208, w7209, w7210, w7211, w7212, w7213, w7214, w7215, w7216, w7217, w7218, w7219, w7220, w7221, w7222, w7223, w7224, w7225, w7226, w7227, w7228, w7229, w7230, w7231, w7232, w7233, w7234, w7235, w7236, w7237, w7238, w7239, w7240, w7241, w7242, w7243, w7244, w7245, w7246, w7247, w7248, w7249, w7250, w7251, w7252, w7253, w7254, w7255, w7256, w7257, w7258, w7259, w7260, w7261, w7262, w7263, w7264, w7265, w7266, w7267, w7268, w7269, w7270, w7271, w7272, w7273, w7274, w7275, w7276, w7277, w7278, w7279, w7280, w7281, w7282, w7283, w7284, w7285, w7286, w7287, w7288, w7289, w7290, w7291, w7292, w7293, w7294, w7295, w7296, w7297, w7298, w7299, w7300, w7301, w7302, w7303, w7304, w7305, w7306, w7307, w7308, w7309, w7310, w7311, w7312, w7313, w7314, w7315, w7316, w7317, w7318, w7319, w7320, w7321, w7322, w7323, w7324, w7325, w7326, w7327, w7328, w7329, w7330, w7331, w7332, w7333, w7334, w7335, w7336, w7337, w7338, w7339, w7340, w7341, w7342, w7343, w7344, w7345, w7346, w7347, w7348, w7349, w7350, w7351, w7352, w7353, w7354, w7355, w7356, w7357, w7358, w7359, w7360, w7361, w7362, w7363, w7364, w7365, w7366, w7367, w7368, w7369, w7370, w7371, w7372, w7373, w7374, w7375, w7376, w7377, w7378, w7379, w7380, w7381, w7382, w7383, w7384, w7385, w7386, w7387, w7388, w7389, w7390, w7391, w7392, w7393, w7394, w7395, w7396, w7397, w7398, w7399, w7400, w7401, w7402, w7403, w7404, w7405, w7406, w7407, w7408, w7409, w7410, w7411, w7412, w7413, w7414, w7415, w7416, w7417, w7418, w7419, w7420, w7421, w7422, w7423, w7424, w7425, w7426, w7427, w7428, w7429, w7430, w7431, w7432, w7433, w7434, w7435, w7436, w7437, w7438, w7439, w7440, w7441, w7442, w7443, w7444, w7445, w7446, w7447, w7448, w7449, w7450, w7451, w7452, w7453, w7454, w7455, w7456, w7457, w7458, w7459, w7460, w7461, w7462, w7463, w7464, w7465, w7466, w7467, w7468, w7469, w7470, w7471, w7472, w7473, w7474, w7475, w7476, w7477, w7478, w7479, w7480, w7481, w7482, w7483, w7484, w7485, w7486, w7487, w7488, w7489, w7490, w7491, w7492, w7493, w7494, w7495, w7496, w7497, w7498, w7499, w7500, w7501, w7502, w7503, w7504, w7505, w7506, w7507, w7508, w7509, w7510, w7511, w7512, w7513, w7514, w7515, w7516, w7517, w7518, w7519, w7520, w7521, w7522, w7523, w7524, w7525, w7526, w7527, w7528, w7529, w7530, w7531, w7532, w7533, w7534, w7535, w7536, w7537, w7538, w7539, w7540, w7541, w7542, w7543, w7544, w7545, w7546, w7547, w7548, w7549, w7550, w7551, w7552, w7553, w7554, w7555, w7556, w7557, w7558, w7559, w7560, w7561, w7562, w7563, w7564, w7565, w7566, w7567, w7568, w7569, w7570, w7571, w7572, w7573, w7574, w7575, w7576, w7577, w7578, w7579, w7580, w7581, w7582, w7583, w7584, w7585, w7586, w7587, w7588, w7589, w7590, w7591, w7592, w7593, w7594, w7595, w7596, w7597, w7598, w7599, w7600, w7601, w7602, w7603, w7604, w7605, w7606, w7607, w7608, w7609, w7610, w7611, w7612, w7613, w7614, w7615, w7616, w7617, w7618, w7619, w7620, w7621, w7622, w7623, w7624, w7625, w7626, w7627, w7628, w7629, w7630, w7631, w7632, w7633, w7634, w7635, w7636, w7637, w7638, w7639, w7640, w7641, w7642, w7643, w7644, w7645, w7646, w7647, w7648, w7649, w7650, w7651, w7652, w7653, w7654, w7655, w7656, w7657, w7658, w7659, w7660, w7661, w7662, w7663, w7664, w7665, w7666, w7667, w7668, w7669, w7670, w7671, w7672, w7673, w7674, w7675, w7676, w7677, w7678, w7679, w7680, w7681, w7682, w7683, w7684, w7685, w7686, w7687, w7688, w7689, w7690, w7691, w7692, w7693, w7694, w7695, w7696, w7697, w7698, w7699, w7700, w7701, w7702, w7703, w7704, w7705, w7706, w7707, w7708, w7709, w7710, w7711, w7712, w7713, w7714, w7715, w7716, w7717, w7718, w7719, w7720, w7721, w7722, w7723, w7724, w7725, w7726, w7727, w7728, w7729, w7730, w7731, w7732, w7733, w7734, w7735, w7736, w7737, w7738, w7739, w7740, w7741, w7742, w7743, w7744, w7745, w7746, w7747, w7748, w7749, w7750, w7751, w7752, w7753, w7754, w7755, w7756, w7757, w7758, w7759, w7760, w7761, w7762, w7763, w7764, w7765, w7766, w7767, w7768, w7769, w7770, w7771, w7772, w7773, w7774, w7775, w7776, w7777, w7778, w7779, w7780, w7781, w7782, w7783, w7784, w7785, w7786, w7787, w7788, w7789, w7790, w7791, w7792, w7793, w7794, w7795, w7796, w7797, w7798, w7799, w7800, w7801, w7802, w7803, w7804, w7805, w7806, w7807, w7808, w7809, w7810, w7811, w7812, w7813, w7814, w7815, w7816, w7817, w7818, w7819, w7820, w7821, w7822, w7823, w7824, w7825, w7826, w7827, w7828, w7829, w7830, w7831, w7832, w7833, w7834, w7835, w7836, w7837, w7838, w7839, w7840, w7841, w7842, w7843, w7844, w7845, w7846, w7847, w7848, w7849, w7850, w7851, w7852, w7853, w7854, w7855, w7856, w7857, w7858, w7859, w7860, w7861, w7862, w7863, w7864, w7865, w7866, w7867, w7868, w7869, w7870, w7871, w7872, w7873, w7874, w7875, w7876, w7877, w7878, w7879, w7880, w7881, w7882, w7883, w7884, w7885, w7886, w7887, w7888, w7889, w7890, w7891, w7892, w7893, w7894, w7895, w7896, w7897, w7898, w7899, w7900, w7901, w7902, w7903, w7904, w7905, w7906, w7907, w7908, w7909, w7910, w7911, w7912, w7913, w7914, w7915, w7916, w7917, w7918, w7919, w7920, w7921, w7922, w7923, w7924, w7925, w7926, w7927, w7928, w7929, w7930, w7931, w7932, w7933, w7934, w7935, w7936, w7937, w7938, w7939, w7940, w7941, w7942, w7943, w7944, w7945, w7946, w7947, w7948, w7949, w7950, w7951, w7952, w7953, w7954, w7955, w7956, w7957, w7958, w7959, w7960, w7961, w7962, w7963, w7964, w7965, w7966, w7967, w7968, w7969, w7970, w7971, w7972, w7973, w7974, w7975, w7976, w7977, w7978, w7979, w7980, w7981, w7982, w7983, w7984, w7985, w7986, w7987, w7988, w7989, w7990, w7991, w7992, w7993, w7994, w7995, w7996, w7997, w7998, w7999, w8000, w8001, w8002, w8003, w8004, w8005, w8006, w8007, w8008, w8009, w8010, w8011, w8012, w8013, w8014, w8015, w8016, w8017, w8018, w8019, w8020, w8021, w8022, w8023, w8024, w8025, w8026, w8027, w8028, w8029, w8030, w8031, w8032, w8033, w8034, w8035, w8036, w8037, w8038, w8039, w8040, w8041, w8042, w8043, w8044, w8045, w8046, w8047, w8048, w8049, w8050, w8051, w8052, w8053, w8054, w8055, w8056, w8057, w8058, w8059, w8060, w8061, w8062, w8063, w8064, w8065, w8066, w8067, w8068, w8069, w8070, w8071, w8072, w8073, w8074, w8075, w8076, w8077, w8078, w8079, w8080, w8081, w8082, w8083, w8084, w8085, w8086, w8087, w8088, w8089, w8090, w8091, w8092, w8093, w8094, w8095, w8096, w8097, w8098, w8099, w8100, w8101, w8102, w8103, w8104, w8105, w8106, w8107, w8108, w8109, w8110, w8111, w8112, w8113, w8114, w8115, w8116, w8117, w8118, w8119, w8120, w8121, w8122, w8123, w8124, w8125, w8126, w8127, w8128, w8129, w8130, w8131, w8132, w8133, w8134, w8135, w8136, w8137, w8138, w8139, w8140, w8141, w8142, w8143, w8144, w8145, w8146, w8147, w8148, w8149, w8150, w8151, w8152, w8153, w8154, w8155, w8156, w8157, w8158, w8159, w8160, w8161, w8162, w8163, w8164, w8165, w8166, w8167, w8168, w8169, w8170, w8171, w8172, w8173, w8174, w8175, w8176, w8177, w8178, w8179, w8180, w8181, w8182, w8183, w8184, w8185, w8186, w8187, w8188, w8189, w8190, w8191, w8192, w8193, w8194, w8195, w8196, w8197, w8198, w8199, w8200, w8201, w8202, w8203, w8204, w8205, w8206, w8207, w8208, w8209, w8210, w8211, w8212, w8213, w8214, w8215, w8216, w8217, w8218, w8219, w8220, w8221, w8222, w8223, w8224, w8225, w8226, w8227, w8228, w8229, w8230, w8231, w8232, w8233, w8234, w8235, w8236, w8237, w8238, w8239, w8240, w8241, w8242, w8243, w8244, w8245, w8246, w8247, w8248, w8249, w8250, w8251, w8252, w8253, w8254, w8255, w8256, w8257, w8258, w8259, w8260, w8261, w8262, w8263, w8264, w8265, w8266, w8267, w8268, w8269, w8270, w8271, w8272, w8273, w8274, w8275, w8276, w8277, w8278, w8279, w8280, w8281, w8282, w8283, w8284, w8285, w8286, w8287, w8288, w8289, w8290, w8291, w8292, w8293, w8294, w8295, w8296, w8297, w8298, w8299, w8300, w8301, w8302, w8303, w8304, w8305, w8306, w8307, w8308, w8309, w8310, w8311, w8312, w8313, w8314, w8315, w8316, w8317, w8318, w8319, w8320, w8321, w8322, w8323, w8324, w8325, w8326, w8327, w8328, w8329, w8330, w8331, w8332, w8333, w8334, w8335, w8336, w8337, w8338, w8339, w8340, w8341, w8342, w8343, w8344, w8345, w8346, w8347, w8348, w8349, w8350, w8351, w8352, w8353, w8354, w8355, w8356, w8357, w8358, w8359, w8360, w8361, w8362, w8363, w8364, w8365, w8366, w8367, w8368, w8369, w8370, w8371, w8372, w8373, w8374, w8375, w8376, w8377, w8378, w8379, w8380, w8381, w8382, w8383, w8384, w8385, w8386, w8387, w8388, w8389, w8390, w8391, w8392, w8393, w8394, w8395, w8396, w8397, w8398, w8399, w8400, w8401, w8402, w8403, w8404, w8405, w8406, w8407, w8408, w8409, w8410, w8411, w8412, w8413, w8414, w8415, w8416, w8417, w8418, w8419, w8420, w8421, w8422, w8423, w8424, w8425, w8426, w8427, w8428, w8429, w8430, w8431, w8432, w8433, w8434, w8435, w8436, w8437, w8438, w8439, w8440, w8441, w8442, w8443, w8444, w8445, w8446, w8447, w8448, w8449, w8450, w8451, w8452, w8453, w8454, w8455, w8456, w8457, w8458, w8459, w8460, w8461, w8462, w8463, w8464, w8465, w8466, w8467, w8468, w8469, w8470, w8471, w8472, w8473, w8474, w8475, w8476, w8477, w8478, w8479, w8480, w8481, w8482, w8483, w8484, w8485, w8486, w8487, w8488, w8489, w8490, w8491, w8492, w8493, w8494, w8495, w8496, w8497, w8498, w8499, w8500, w8501, w8502, w8503, w8504, w8505, w8506, w8507, w8508, w8509, w8510, w8511, w8512, w8513, w8514, w8515, w8516, w8517, w8518, w8519, w8520, w8521, w8522, w8523, w8524, w8525, w8526, w8527, w8528, w8529, w8530, w8531, w8532, w8533, w8534, w8535, w8536, w8537, w8538, w8539, w8540, w8541, w8542, w8543, w8544, w8545, w8546, w8547, w8548, w8549, w8550, w8551, w8552, w8553, w8554, w8555, w8556, w8557, w8558, w8559, w8560, w8561, w8562, w8563, w8564, w8565, w8566, w8567, w8568, w8569, w8570, w8571, w8572, w8573, w8574, w8575, w8576, w8577, w8578, w8579, w8580, w8581, w8582, w8583, w8584, w8585, w8586, w8587, w8588, w8589, w8590, w8591, w8592, w8593, w8594, w8595, w8596, w8597, w8598, w8599, w8600, w8601, w8602, w8603, w8604, w8605, w8606, w8607, w8608, w8609, w8610, w8611, w8612, w8613, w8614, w8615, w8616, w8617, w8618, w8619, w8620, w8621, w8622, w8623, w8624, w8625, w8626, w8627, w8628, w8629, w8630, w8631, w8632, w8633, w8634, w8635, w8636, w8637, w8638, w8639, w8640, w8641, w8642, w8643, w8644, w8645, w8646, w8647, w8648, w8649, w8650, w8651, w8652, w8653, w8654, w8655, w8656, w8657, w8658, w8659, w8660, w8661, w8662, w8663, w8664, w8665, w8666, w8667, w8668, w8669, w8670, w8671, w8672, w8673, w8674, w8675, w8676, w8677, w8678, w8679, w8680, w8681, w8682, w8683, w8684, w8685, w8686, w8687, w8688, w8689, w8690, w8691, w8692, w8693, w8694, w8695, w8696, w8697, w8698, w8699, w8700, w8701, w8702, w8703, w8704, w8705, w8706, w8707, w8708, w8709, w8710, w8711, w8712, w8713, w8714, w8715, w8716, w8717, w8718, w8719, w8720, w8721, w8722, w8723, w8724, w8725, w8726, w8727, w8728, w8729, w8730, w8731, w8732, w8733, w8734, w8735, w8736, w8737, w8738, w8739, w8740, w8741, w8742, w8743, w8744, w8745, w8746, w8747, w8748, w8749, w8750, w8751, w8752, w8753, w8754, w8755, w8756, w8757, w8758, w8759, w8760, w8761, w8762, w8763, w8764, w8765, w8766, w8767, w8768, w8769, w8770, w8771, w8772, w8773, w8774, w8775, w8776, w8777, w8778, w8779, w8780, w8781, w8782, w8783, w8784, w8785, w8786, w8787, w8788, w8789, w8790, w8791, w8792, w8793, w8794, w8795, w8796, w8797, w8798, w8799, w8800, w8801, w8802, w8803, w8804, w8805, w8806, w8807, w8808, w8809, w8810, w8811, w8812, w8813, w8814, w8815, w8816, w8817, w8818, w8819, w8820, w8821, w8822, w8823, w8824, w8825, w8826, w8827, w8828, w8829, w8830, w8831, w8832, w8833, w8834, w8835, w8836, w8837, w8838, w8839, w8840, w8841, w8842, w8843, w8844, w8845, w8846, w8847, w8848, w8849, w8850, w8851, w8852, w8853, w8854, w8855, w8856, w8857, w8858, w8859, w8860, w8861, w8862, w8863, w8864, w8865, w8866, w8867, w8868, w8869, w8870, w8871, w8872, w8873, w8874, w8875, w8876, w8877, w8878, w8879, w8880, w8881, w8882, w8883, w8884, w8885, w8886, w8887, w8888, w8889, w8890, w8891, w8892, w8893, w8894, w8895, w8896, w8897, w8898, w8899, w8900, w8901, w8902, w8903, w8904, w8905, w8906, w8907, w8908, w8909, w8910, w8911, w8912, w8913, w8914, w8915, w8916, w8917, w8918, w8919, w8920, w8921, w8922, w8923, w8924, w8925, w8926, w8927, w8928, w8929, w8930, w8931, w8932, w8933, w8934, w8935, w8936, w8937, w8938, w8939, w8940, w8941, w8942, w8943, w8944, w8945, w8946, w8947, w8948, w8949, w8950, w8951, w8952, w8953, w8954, w8955, w8956, w8957, w8958, w8959, w8960, w8961, w8962, w8963, w8964, w8965, w8966, w8967, w8968, w8969, w8970, w8971, w8972, w8973, w8974, w8975, w8976, w8977, w8978, w8979, w8980, w8981, w8982, w8983, w8984, w8985, w8986, w8987, w8988, w8989, w8990, w8991, w8992, w8993, w8994, w8995, w8996, w8997, w8998, w8999, w9000, w9001, w9002, w9003, w9004, w9005, w9006, w9007, w9008, w9009, w9010, w9011, w9012, w9013, w9014, w9015, w9016, w9017, w9018, w9019, w9020, w9021, w9022, w9023, w9024, w9025, w9026, w9027, w9028, w9029, w9030, w9031, w9032, w9033, w9034, w9035, w9036, w9037, w9038, w9039, w9040, w9041, w9042, w9043, w9044, w9045, w9046, w9047, w9048, w9049, w9050, w9051, w9052, w9053, w9054, w9055, w9056, w9057, w9058, w9059, w9060, w9061, w9062, w9063, w9064, w9065, w9066, w9067, w9068, w9069, w9070, w9071, w9072, w9073, w9074, w9075, w9076, w9077, w9078, w9079, w9080, w9081, w9082, w9083, w9084, w9085, w9086, w9087, w9088, w9089, w9090, w9091, w9092, w9093, w9094, w9095, w9096, w9097, w9098, w9099, w9100, w9101, w9102, w9103, w9104, w9105, w9106, w9107, w9108, w9109, w9110, w9111, w9112, w9113, w9114, w9115, w9116, w9117, w9118, w9119, w9120, w9121, w9122, w9123, w9124, w9125, w9126, w9127, w9128, w9129, w9130, w9131, w9132, w9133, w9134, w9135, w9136, w9137, w9138, w9139, w9140, w9141, w9142, w9143, w9144, w9145, w9146, w9147, w9148, w9149, w9150, w9151, w9152, w9153, w9154, w9155, w9156, w9157, w9158, w9159, w9160, w9161, w9162, w9163, w9164, w9165, w9166, w9167, w9168, w9169, w9170, w9171, w9172, w9173, w9174, w9175, w9176, w9177, w9178, w9179, w9180, w9181, w9182, w9183, w9184, w9185, w9186, w9187, w9188, w9189, w9190, w9191, w9192, w9193, w9194, w9195, w9196, w9197, w9198, w9199, w9200, w9201, w9202, w9203, w9204, w9205, w9206, w9207, w9208, w9209, w9210, w9211, w9212, w9213, w9214, w9215, w9216, w9217, w9218, w9219, w9220, w9221, w9222, w9223, w9224, w9225, w9226, w9227, w9228, w9229, w9230, w9231, w9232, w9233, w9234, w9235, w9236, w9237, w9238, w9239, w9240, w9241, w9242, w9243, w9244, w9245, w9246, w9247, w9248, w9249, w9250, w9251, w9252, w9253, w9254, w9255, w9256, w9257, w9258, w9259, w9260, w9261, w9262, w9263, w9264, w9265, w9266, w9267, w9268, w9269, w9270, w9271, w9272, w9273, w9274, w9275, w9276, w9277, w9278, w9279, w9280, w9281, w9282, w9283, w9284, w9285, w9286, w9287, w9288, w9289, w9290, w9291, w9292, w9293, w9294, w9295, w9296, w9297, w9298, w9299, w9300, w9301, w9302, w9303, w9304, w9305, w9306, w9307, w9308, w9309, w9310, w9311, w9312, w9313, w9314, w9315, w9316, w9317, w9318, w9319, w9320, w9321, w9322, w9323, w9324, w9325, w9326, w9327, w9328, w9329, w9330, w9331, w9332, w9333, w9334, w9335, w9336, w9337, w9338, w9339, w9340, w9341, w9342, w9343, w9344, w9345, w9346, w9347, w9348, w9349, w9350, w9351, w9352, w9353, w9354, w9355, w9356, w9357, w9358, w9359, w9360, w9361, w9362, w9363, w9364, w9365, w9366, w9367, w9368, w9369, w9370, w9371, w9372, w9373, w9374, w9375, w9376, w9377, w9378, w9379, w9380, w9381, w9382, w9383, w9384, w9385, w9386, w9387, w9388, w9389, w9390, w9391, w9392, w9393, w9394, w9395, w9396, w9397, w9398, w9399, w9400, w9401, w9402, w9403, w9404, w9405, w9406, w9407, w9408, w9409, w9410, w9411, w9412, w9413, w9414, w9415, w9416, w9417, w9418, w9419, w9420, w9421, w9422, w9423, w9424, w9425, w9426, w9427, w9428, w9429, w9430, w9431, w9432, w9433, w9434, w9435, w9436, w9437, w9438, w9439, w9440, w9441, w9442, w9443, w9444, w9445, w9446, w9447, w9448, w9449, w9450, w9451, w9452, w9453, w9454, w9455, w9456, w9457, w9458, w9459, w9460, w9461, w9462, w9463, w9464, w9465, w9466, w9467, w9468, w9469, w9470, w9471, w9472, w9473, w9474, w9475, w9476, w9477, w9478, w9479, w9480, w9481, w9482, w9483, w9484, w9485, w9486, w9487, w9488, w9489, w9490, w9491, w9492, w9493, w9494, w9495, w9496, w9497, w9498, w9499, w9500, w9501, w9502, w9503, w9504, w9505, w9506, w9507, w9508, w9509, w9510, w9511, w9512, w9513, w9514, w9515, w9516, w9517, w9518, w9519, w9520, w9521, w9522, w9523, w9524, w9525, w9526, w9527, w9528, w9529, w9530, w9531, w9532, w9533, w9534, w9535, w9536, w9537, w9538, w9539, w9540, w9541, w9542, w9543, w9544, w9545, w9546, w9547, w9548, w9549, w9550, w9551, w9552, w9553, w9554, w9555, w9556, w9557, w9558, w9559, w9560, w9561, w9562, w9563, w9564, w9565, w9566, w9567, w9568, w9569, w9570, w9571, w9572, w9573, w9574, w9575, w9576, w9577, w9578, w9579, w9580, w9581, w9582, w9583, w9584, w9585, w9586, w9587, w9588, w9589, w9590, w9591, w9592, w9593, w9594, w9595, w9596, w9597, w9598, w9599, w9600, w9601, w9602, w9603, w9604, w9605, w9606, w9607, w9608, w9609, w9610, w9611, w9612, w9613, w9614, w9615, w9616, w9617, w9618, w9619, w9620, w9621, w9622, w9623, w9624, w9625, w9626, w9627, w9628, w9629, w9630, w9631, w9632, w9633, w9634, w9635, w9636, w9637, w9638, w9639, w9640, w9641, w9642, w9643, w9644, w9645, w9646, w9647, w9648, w9649, w9650, w9651, w9652, w9653, w9654, w9655, w9656, w9657, w9658, w9659, w9660, w9661, w9662, w9663, w9664, w9665, w9666, w9667, w9668, w9669, w9670, w9671, w9672, w9673, w9674, w9675, w9676, w9677, w9678, w9679, w9680, w9681, w9682, w9683, w9684, w9685, w9686, w9687, w9688, w9689, w9690, w9691, w9692, w9693, w9694, w9695, w9696, w9697, w9698, w9699, w9700, w9701, w9702, w9703, w9704, w9705, w9706, w9707, w9708, w9709, w9710, w9711, w9712, w9713, w9714, w9715, w9716, w9717, w9718, w9719, w9720, w9721, w9722, w9723, w9724, w9725, w9726, w9727, w9728, w9729, w9730, w9731, w9732, w9733, w9734, w9735, w9736, w9737, w9738, w9739, w9740, w9741, w9742, w9743, w9744, w9745, w9746, w9747, w9748, w9749, w9750, w9751, w9752, w9753, w9754, w9755, w9756, w9757, w9758, w9759, w9760, w9761, w9762, w9763, w9764, w9765, w9766, w9767, w9768, w9769, w9770, w9771, w9772, w9773, w9774, w9775, w9776, w9777, w9778, w9779, w9780, w9781, w9782, w9783, w9784, w9785, w9786, w9787, w9788, w9789, w9790, w9791, w9792, w9793, w9794, w9795, w9796, w9797, w9798, w9799, w9800, w9801, w9802, w9803, w9804, w9805, w9806, w9807, w9808, w9809, w9810, w9811, w9812, w9813, w9814, w9815, w9816, w9817, w9818, w9819, w9820, w9821, w9822, w9823, w9824, w9825, w9826, w9827, w9828, w9829, w9830, w9831, w9832, w9833, w9834, w9835, w9836, w9837, w9838, w9839, w9840, w9841, w9842, w9843, w9844, w9845, w9846, w9847, w9848, w9849, w9850, w9851, w9852, w9853, w9854, w9855, w9856, w9857, w9858, w9859, w9860, w9861, w9862, w9863, w9864, w9865, w9866, w9867, w9868, w9869, w9870, w9871, w9872, w9873, w9874, w9875, w9876, w9877, w9878, w9879, w9880, w9881, w9882, w9883, w9884, w9885, w9886, w9887, w9888, w9889, w9890, w9891, w9892, w9893, w9894, w9895, w9896, w9897, w9898, w9899, w9900, w9901, w9902, w9903, w9904, w9905, w9906, w9907, w9908, w9909, w9910, w9911, w9912, w9913, w9914, w9915, w9916, w9917, w9918, w9919, w9920, w9921, w9922, w9923, w9924, w9925, w9926, w9927, w9928, w9929, w9930, w9931, w9932, w9933, w9934, w9935, w9936, w9937, w9938, w9939, w9940, w9941, w9942, w9943, w9944, w9945, w9946, w9947, w9948, w9949, w9950, w9951, w9952, w9953, w9954, w9955, w9956, w9957, w9958, w9959, w9960, w9961, w9962, w9963, w9964, w9965, w9966, w9967, w9968, w9969, w9970, w9971, w9972, w9973, w9974, w9975, w9976, w9977, w9978, w9979, w9980, w9981, w9982, w9983, w9984, w9985, w9986, w9987, w9988, w9989, w9990, w9991, w9992, w9993, w9994, w9995, w9996, w9997, w9998, w9999, w10000, w10001, w10002, w10003, w10004, w10005, w10006, w10007, w10008, w10009, w10010, w10011, w10012, w10013, w10014, w10015, w10016, w10017, w10018, w10019, w10020, w10021, w10022, w10023, w10024, w10025, w10026, w10027, w10028, w10029, w10030, w10031, w10032, w10033, w10034, w10035, w10036, w10037, w10038, w10039, w10040, w10041, w10042, w10043, w10044, w10045, w10046, w10047, w10048, w10049, w10050, w10051, w10052, w10053, w10054, w10055, w10056, w10057, w10058, w10059, w10060, w10061, w10062, w10063, w10064, w10065, w10066, w10067, w10068, w10069, w10070, w10071, w10072, w10073, w10074, w10075, w10076, w10077, w10078, w10079, w10080, w10081, w10082, w10083, w10084, w10085, w10086, w10087, w10088, w10089, w10090, w10091, w10092, w10093, w10094, w10095, w10096, w10097, w10098, w10099, w10100, w10101, w10102, w10103, w10104, w10105, w10106, w10107, w10108, w10109, w10110, w10111, w10112, w10113, w10114, w10115, w10116, w10117, w10118, w10119, w10120, w10121, w10122, w10123, w10124, w10125, w10126, w10127, w10128, w10129, w10130, w10131, w10132, w10133, w10134, w10135, w10136, w10137, w10138, w10139, w10140, w10141, w10142, w10143, w10144, w10145, w10146, w10147, w10148, w10149, w10150, w10151, w10152, w10153, w10154, w10155, w10156, w10157, w10158, w10159, w10160, w10161, w10162, w10163, w10164, w10165, w10166, w10167, w10168, w10169, w10170, w10171, w10172, w10173, w10174, w10175, w10176, w10177, w10178, w10179, w10180, w10181, w10182, w10183, w10184, w10185, w10186, w10187, w10188, w10189, w10190, w10191, w10192, w10193, w10194, w10195, w10196, w10197, w10198, w10199, w10200, w10201, w10202, w10203, w10204, w10205, w10206, w10207, w10208, w10209, w10210, w10211, w10212, w10213, w10214, w10215, w10216, w10217, w10218, w10219, w10220, w10221, w10222, w10223, w10224, w10225, w10226, w10227, w10228, w10229, w10230, w10231, w10232, w10233, w10234, w10235, w10236, w10237, w10238, w10239, w10240, w10241, w10242, w10243, w10244, w10245, w10246, w10247, w10248, w10249, w10250, w10251, w10252, w10253, w10254, w10255, w10256, w10257, w10258, w10259, w10260, w10261, w10262, w10263, w10264, w10265, w10266, w10267, w10268, w10269, w10270, w10271, w10272, w10273, w10274, w10275, w10276, w10277, w10278, w10279, w10280, w10281, w10282, w10283, w10284, w10285, w10286, w10287, w10288, w10289, w10290, w10291, w10292, w10293, w10294, w10295, w10296, w10297, w10298, w10299, w10300, w10301, w10302, w10303, w10304, w10305, w10306, w10307, w10308, w10309, w10310, w10311, w10312, w10313, w10314, w10315, w10316, w10317, w10318, w10319, w10320, w10321, w10322, w10323, w10324, w10325, w10326, w10327, w10328, w10329, w10330, w10331, w10332, w10333, w10334, w10335, w10336, w10337, w10338, w10339, w10340, w10341, w10342, w10343, w10344, w10345, w10346, w10347, w10348, w10349, w10350, w10351, w10352, w10353, w10354, w10355, w10356, w10357, w10358, w10359, w10360, w10361, w10362, w10363, w10364, w10365, w10366, w10367, w10368, w10369, w10370, w10371, w10372, w10373, w10374, w10375, w10376, w10377, w10378, w10379, w10380, w10381, w10382, w10383, w10384, w10385, w10386, w10387, w10388, w10389, w10390, w10391, w10392, w10393, w10394, w10395, w10396, w10397, w10398, w10399, w10400, w10401, w10402, w10403, w10404, w10405, w10406, w10407, w10408, w10409, w10410, w10411, w10412, w10413, w10414, w10415, w10416, w10417, w10418, w10419, w10420, w10421, w10422, w10423, w10424, w10425, w10426, w10427, w10428, w10429, w10430, w10431, w10432, w10433, w10434, w10435, w10436, w10437, w10438, w10439, w10440, w10441, w10442, w10443, w10444, w10445, w10446, w10447, w10448, w10449, w10450, w10451, w10452, w10453, w10454, w10455, w10456, w10457, w10458, w10459, w10460, w10461, w10462, w10463, w10464, w10465, w10466, w10467, w10468, w10469, w10470, w10471, w10472, w10473, w10474, w10475, w10476, w10477, w10478, w10479, w10480, w10481, w10482, w10483, w10484, w10485, w10486, w10487, w10488, w10489, w10490, w10491, w10492, w10493, w10494, w10495, w10496, w10497, w10498, w10499, w10500, w10501, w10502, w10503, w10504, w10505, w10506, w10507, w10508, w10509, w10510, w10511, w10512, w10513, w10514, w10515, w10516, w10517, w10518, w10519, w10520, w10521, w10522, w10523, w10524, w10525, w10526, w10527, w10528, w10529, w10530, w10531, w10532, w10533, w10534, w10535, w10536, w10537, w10538, w10539, w10540, w10541, w10542, w10543, w10544, w10545, w10546, w10547, w10548, w10549, w10550, w10551, w10552, w10553, w10554, w10555, w10556, w10557, w10558, w10559, w10560, w10561, w10562, w10563, w10564, w10565, w10566, w10567, w10568, w10569, w10570, w10571, w10572, w10573, w10574, w10575, w10576, w10577, w10578, w10579, w10580, w10581, w10582, w10583, w10584, w10585, w10586, w10587, w10588, w10589, w10590, w10591, w10592, w10593, w10594, w10595, w10596, w10597, w10598, w10599, w10600, w10601, w10602, w10603, w10604, w10605, w10606, w10607, w10608, w10609, w10610, w10611, w10612, w10613, w10614, w10615, w10616, w10617, w10618, w10619, w10620, w10621, w10622, w10623, w10624, w10625, w10626, w10627, w10628, w10629, w10630, w10631, w10632, w10633, w10634, w10635, w10636, w10637, w10638, w10639, w10640, w10641, w10642, w10643, w10644, w10645, w10646, w10647, w10648, w10649, w10650, w10651, w10652, w10653, w10654, w10655, w10656, w10657, w10658, w10659, w10660, w10661, w10662, w10663, w10664, w10665, w10666, w10667, w10668, w10669, w10670, w10671, w10672, w10673, w10674, w10675, w10676, w10677, w10678, w10679, w10680, w10681, w10682, w10683, w10684, w10685, w10686, w10687, w10688, w10689, w10690, w10691, w10692, w10693, w10694, w10695, w10696, w10697, w10698, w10699, w10700, w10701, w10702, w10703, w10704, w10705, w10706, w10707, w10708, w10709, w10710, w10711, w10712, w10713, w10714, w10715, w10716, w10717, w10718, w10719, w10720, w10721, w10722, w10723, w10724, w10725, w10726, w10727, w10728, w10729, w10730, w10731, w10732, w10733, w10734, w10735, w10736, w10737, w10738, w10739, w10740, w10741, w10742, w10743, w10744, w10745, w10746, w10747, w10748, w10749, w10750, w10751, w10752, w10753, w10754, w10755, w10756, w10757, w10758, w10759, w10760, w10761, w10762, w10763, w10764, w10765, w10766, w10767, w10768, w10769, w10770, w10771, w10772, w10773, w10774, w10775, w10776, w10777, w10778, w10779, w10780, w10781, w10782, w10783, w10784, w10785, w10786, w10787, w10788, w10789, w10790, w10791, w10792, w10793, w10794, w10795, w10796, w10797, w10798, w10799, w10800, w10801, w10802, w10803, w10804, w10805, w10806, w10807, w10808, w10809, w10810, w10811, w10812, w10813, w10814, w10815, w10816, w10817, w10818, w10819, w10820, w10821, w10822, w10823, w10824, w10825, w10826, w10827, w10828, w10829, w10830, w10831, w10832, w10833, w10834, w10835, w10836, w10837, w10838, w10839, w10840, w10841, w10842, w10843, w10844, w10845, w10846, w10847, w10848, w10849, w10850, w10851, w10852, w10853, w10854, w10855, w10856, w10857, w10858, w10859, w10860, w10861, w10862, w10863, w10864, w10865, w10866, w10867, w10868, w10869, w10870, w10871, w10872, w10873, w10874, w10875, w10876, w10877, w10878, w10879, w10880, w10881, w10882, w10883, w10884, w10885, w10886, w10887, w10888, w10889, w10890, w10891, w10892, w10893, w10894, w10895, w10896, w10897, w10898, w10899, w10900, w10901, w10902, w10903, w10904, w10905, w10906, w10907, w10908, w10909, w10910, w10911, w10912, w10913, w10914, w10915, w10916, w10917, w10918, w10919, w10920, w10921, w10922, w10923, w10924, w10925, w10926, w10927, w10928, w10929, w10930, w10931, w10932, w10933, w10934, w10935, w10936, w10937, w10938, w10939, w10940, w10941, w10942, w10943, w10944, w10945, w10946, w10947, w10948, w10949, w10950, w10951, w10952, w10953, w10954, w10955, w10956, w10957, w10958, w10959, w10960, w10961, w10962, w10963, w10964, w10965, w10966, w10967, w10968, w10969, w10970, w10971, w10972, w10973, w10974, w10975, w10976, w10977, w10978, w10979, w10980, w10981, w10982, w10983, w10984, w10985, w10986, w10987, w10988, w10989, w10990, w10991, w10992, w10993, w10994, w10995, w10996, w10997, w10998, w10999, w11000, w11001, w11002, w11003, w11004, w11005, w11006, w11007, w11008, w11009, w11010, w11011, w11012, w11013, w11014, w11015, w11016, w11017, w11018, w11019, w11020, w11021, w11022, w11023, w11024, w11025, w11026, w11027, w11028, w11029, w11030, w11031, w11032, w11033, w11034, w11035, w11036, w11037, w11038, w11039, w11040, w11041, w11042, w11043, w11044, w11045, w11046, w11047, w11048, w11049, w11050, w11051, w11052, w11053, w11054, w11055, w11056, w11057, w11058, w11059, w11060, w11061, w11062, w11063, w11064, w11065, w11066, w11067, w11068, w11069, w11070, w11071, w11072, w11073, w11074, w11075, w11076, w11077, w11078, w11079, w11080, w11081, w11082, w11083, w11084, w11085, w11086, w11087, w11088, w11089, w11090, w11091, w11092, w11093, w11094, w11095, w11096, w11097, w11098, w11099, w11100, w11101, w11102, w11103, w11104, w11105, w11106, w11107, w11108, w11109, w11110, w11111, w11112, w11113, w11114, w11115, w11116, w11117, w11118, w11119, w11120, w11121, w11122, w11123, w11124, w11125, w11126, w11127, w11128, w11129, w11130, w11131, w11132, w11133, w11134, w11135, w11136, w11137, w11138, w11139, w11140, w11141, w11142, w11143, w11144, w11145, w11146, w11147, w11148, w11149, w11150, w11151, w11152, w11153, w11154, w11155, w11156, w11157, w11158, w11159, w11160, w11161, w11162, w11163, w11164, w11165, w11166, w11167, w11168, w11169, w11170, w11171, w11172, w11173, w11174, w11175, w11176, w11177, w11178, w11179, w11180, w11181, w11182, w11183, w11184, w11185, w11186, w11187, w11188, w11189, w11190, w11191, w11192, w11193, w11194, w11195, w11196, w11197, w11198, w11199, w11200, w11201, w11202, w11203, w11204, w11205, w11206, w11207, w11208, w11209, w11210, w11211, w11212, w11213, w11214, w11215, w11216, w11217, w11218, w11219, w11220, w11221, w11222, w11223, w11224, w11225, w11226, w11227, w11228, w11229, w11230, w11231, w11232, w11233, w11234, w11235, w11236, w11237, w11238, w11239, w11240, w11241, w11242, w11243, w11244, w11245, w11246, w11247, w11248, w11249, w11250, w11251, w11252, w11253, w11254, w11255, w11256, w11257, w11258, w11259, w11260, w11261, w11262, w11263, w11264, w11265, w11266, w11267, w11268, w11269, w11270, w11271, w11272, w11273, w11274, w11275, w11276, w11277, w11278, w11279, w11280, w11281, w11282, w11283, w11284, w11285, w11286, w11287, w11288, w11289, w11290, w11291, w11292, w11293, w11294, w11295, w11296, w11297, w11298, w11299, w11300, w11301, w11302, w11303, w11304, w11305, w11306, w11307, w11308, w11309, w11310, w11311, w11312, w11313, w11314, w11315, w11316, w11317, w11318, w11319, w11320, w11321, w11322, w11323, w11324, w11325, w11326, w11327, w11328, w11329, w11330, w11331, w11332, w11333, w11334, w11335, w11336, w11337, w11338, w11339, w11340, w11341, w11342, w11343, w11344, w11345, w11346, w11347, w11348, w11349, w11350, w11351, w11352, w11353, w11354, w11355, w11356, w11357, w11358, w11359, w11360, w11361, w11362, w11363, w11364, w11365, w11366, w11367, w11368, w11369, w11370, w11371, w11372, w11373, w11374, w11375, w11376, w11377, w11378, w11379, w11380, w11381, w11382, w11383, w11384, w11385, w11386, w11387, w11388, w11389, w11390, w11391, w11392, w11393, w11394, w11395, w11396, w11397, w11398, w11399, w11400, w11401, w11402, w11403, w11404, w11405, w11406, w11407, w11408, w11409, w11410, w11411, w11412, w11413, w11414, w11415, w11416, w11417, w11418, w11419, w11420, w11421, w11422, w11423, w11424, w11425, w11426, w11427, w11428, w11429, w11430, w11431, w11432, w11433, w11434, w11435, w11436, w11437, w11438, w11439, w11440, w11441, w11442, w11443, w11444, w11445, w11446, w11447, w11448, w11449, w11450, w11451, w11452, w11453, w11454, w11455, w11456, w11457, w11458, w11459, w11460, w11461, w11462, w11463, w11464, w11465, w11466, w11467, w11468, w11469, w11470, w11471, w11472, w11473, w11474, w11475, w11476, w11477, w11478, w11479, w11480, w11481, w11482, w11483, w11484, w11485, w11486, w11487, w11488, w11489, w11490, w11491, w11492, w11493, w11494, w11495, w11496, w11497, w11498, w11499, w11500, w11501, w11502, w11503, w11504, w11505, w11506, w11507, w11508, w11509, w11510, w11511, w11512, w11513, w11514, w11515, w11516, w11517, w11518, w11519, w11520, w11521, w11522, w11523, w11524, w11525, w11526, w11527, w11528, w11529, w11530, w11531, w11532, w11533, w11534, w11535, w11536, w11537, w11538, w11539, w11540, w11541, w11542, w11543, w11544, w11545, w11546, w11547, w11548, w11549, w11550, w11551, w11552, w11553, w11554, w11555, w11556, w11557, w11558, w11559, w11560, w11561, w11562, w11563, w11564, w11565, w11566, w11567, w11568, w11569, w11570, w11571, w11572, w11573, w11574, w11575, w11576, w11577, w11578, w11579, w11580, w11581, w11582, w11583, w11584, w11585, w11586, w11587, w11588, w11589, w11590, w11591, w11592, w11593, w11594, w11595, w11596, w11597, w11598, w11599, w11600, w11601, w11602, w11603, w11604, w11605, w11606, w11607, w11608, w11609, w11610, w11611, w11612, w11613, w11614, w11615, w11616, w11617, w11618, w11619, w11620, w11621, w11622, w11623, w11624, w11625, w11626, w11627, w11628, w11629, w11630, w11631, w11632, w11633, w11634, w11635, w11636, w11637, w11638, w11639, w11640, w11641, w11642, w11643, w11644, w11645, w11646, w11647, w11648, w11649, w11650, w11651, w11652, w11653, w11654, w11655, w11656, w11657, w11658, w11659, w11660, w11661, w11662, w11663, w11664, w11665, w11666, w11667, w11668, w11669, w11670, w11671, w11672, w11673, w11674, w11675, w11676, w11677, w11678, w11679, w11680, w11681, w11682, w11683, w11684, w11685, w11686, w11687, w11688, w11689, w11690, w11691, w11692, w11693, w11694, w11695, w11696, w11697, w11698, w11699, w11700, w11701, w11702, w11703, w11704, w11705, w11706, w11707, w11708, w11709, w11710, w11711, w11712, w11713, w11714, w11715, w11716, w11717, w11718, w11719, w11720, w11721, w11722, w11723, w11724, w11725, w11726, w11727, w11728, w11729, w11730, w11731, w11732, w11733, w11734, w11735, w11736, w11737, w11738, w11739, w11740, w11741, w11742, w11743, w11744, w11745, w11746, w11747, w11748, w11749, w11750, w11751, w11752, w11753, w11754, w11755, w11756, w11757, w11758, w11759, w11760, w11761, w11762, w11763, w11764, w11765, w11766, w11767, w11768, w11769, w11770, w11771, w11772, w11773, w11774, w11775, w11776, w11777, w11778, w11779, w11780, w11781, w11782, w11783, w11784, w11785, w11786, w11787, w11788, w11789, w11790, w11791, w11792, w11793, w11794, w11795, w11796, w11797, w11798, w11799, w11800, w11801, w11802, w11803, w11804, w11805, w11806, w11807, w11808, w11809, w11810, w11811, w11812, w11813, w11814, w11815, w11816, w11817, w11818, w11819, w11820, w11821, w11822, w11823, w11824, w11825, w11826, w11827, w11828, w11829, w11830, w11831, w11832, w11833, w11834, w11835, w11836, w11837, w11838, w11839, w11840, w11841, w11842, w11843, w11844, w11845, w11846, w11847, w11848, w11849, w11850, w11851, w11852, w11853, w11854, w11855, w11856, w11857, w11858, w11859, w11860, w11861, w11862, w11863, w11864, w11865, w11866, w11867, w11868, w11869, w11870, w11871, w11872, w11873, w11874, w11875, w11876, w11877, w11878, w11879, w11880, w11881, w11882, w11883, w11884, w11885, w11886, w11887, w11888, w11889, w11890, w11891, w11892, w11893, w11894, w11895, w11896, w11897, w11898, w11899, w11900, w11901, w11902, w11903, w11904, w11905, w11906, w11907, w11908, w11909, w11910, w11911, w11912, w11913, w11914, w11915, w11916, w11917, w11918, w11919, w11920, w11921, w11922, w11923, w11924, w11925, w11926, w11927, w11928, w11929, w11930, w11931, w11932, w11933, w11934, w11935, w11936, w11937, w11938, w11939, w11940, w11941, w11942, w11943, w11944, w11945, w11946, w11947, w11948, w11949, w11950, w11951, w11952, w11953, w11954, w11955, w11956, w11957, w11958, w11959, w11960, w11961, w11962, w11963, w11964, w11965, w11966, w11967, w11968, w11969, w11970, w11971, w11972, w11973, w11974, w11975, w11976, w11977, w11978, w11979, w11980, w11981, w11982, w11983, w11984, w11985, w11986, w11987, w11988, w11989, w11990, w11991, w11992, w11993, w11994, w11995, w11996, w11997, w11998, w11999, w12000, w12001, w12002, w12003, w12004, w12005, w12006, w12007, w12008, w12009, w12010, w12011, w12012, w12013, w12014, w12015, w12016, w12017, w12018, w12019, w12020, w12021, w12022, w12023, w12024, w12025, w12026, w12027, w12028, w12029, w12030, w12031, w12032, w12033, w12034, w12035, w12036, w12037, w12038, w12039, w12040, w12041, w12042, w12043, w12044, w12045, w12046, w12047, w12048, w12049, w12050, w12051, w12052, w12053, w12054, w12055, w12056, w12057, w12058, w12059, w12060, w12061, w12062, w12063, w12064, w12065, w12066, w12067, w12068, w12069, w12070, w12071, w12072, w12073, w12074, w12075, w12076, w12077, w12078, w12079, w12080, w12081, w12082, w12083, w12084, w12085, w12086, w12087, w12088, w12089, w12090, w12091, w12092, w12093, w12094, w12095, w12096, w12097, w12098, w12099, w12100, w12101, w12102, w12103, w12104, w12105, w12106, w12107, w12108, w12109, w12110, w12111, w12112, w12113, w12114, w12115, w12116, w12117, w12118, w12119, w12120, w12121, w12122, w12123, w12124, w12125, w12126, w12127, w12128, w12129, w12130, w12131, w12132, w12133, w12134, w12135, w12136, w12137, w12138, w12139, w12140, w12141, w12142, w12143, w12144, w12145, w12146, w12147, w12148, w12149, w12150, w12151, w12152, w12153, w12154, w12155, w12156, w12157, w12158, w12159, w12160, w12161, w12162, w12163, w12164, w12165, w12166, w12167, w12168, w12169, w12170, w12171, w12172, w12173, w12174, w12175, w12176, w12177, w12178, w12179, w12180, w12181, w12182, w12183, w12184, w12185, w12186, w12187, w12188, w12189, w12190, w12191, w12192, w12193, w12194, w12195, w12196, w12197, w12198, w12199, w12200, w12201, w12202, w12203, w12204, w12205, w12206, w12207, w12208, w12209, w12210, w12211, w12212, w12213, w12214, w12215, w12216, w12217, w12218, w12219, w12220, w12221, w12222, w12223, w12224, w12225, w12226, w12227, w12228, w12229, w12230, w12231, w12232, w12233, w12234, w12235, w12236, w12237, w12238, w12239, w12240, w12241, w12242, w12243, w12244, w12245, w12246, w12247, w12248, w12249, w12250, w12251, w12252, w12253, w12254, w12255, w12256, w12257, w12258, w12259, w12260, w12261, w12262, w12263, w12264, w12265, w12266, w12267, w12268, w12269, w12270, w12271, w12272, w12273, w12274, w12275, w12276, w12277, w12278, w12279, w12280, w12281, w12282, w12283, w12284, w12285, w12286, w12287, w12288, w12289, w12290, w12291, w12292, w12293, w12294, w12295, w12296, w12297, w12298, w12299, w12300, w12301, w12302, w12303, w12304, w12305, w12306, w12307, w12308, w12309, w12310, w12311, w12312, w12313, w12314, w12315, w12316, w12317, w12318, w12319, w12320, w12321, w12322, w12323, w12324, w12325, w12326, w12327, w12328, w12329, w12330, w12331, w12332, w12333, w12334, w12335, w12336, w12337, w12338, w12339, w12340, w12341, w12342, w12343, w12344, w12345, w12346, w12347, w12348, w12349, w12350, w12351, w12352, w12353, w12354, w12355, w12356, w12357, w12358, w12359, w12360, w12361, w12362, w12363, w12364, w12365, w12366, w12367, w12368, w12369, w12370, w12371, w12372, w12373, w12374, w12375, w12376, w12377, w12378, w12379, w12380, w12381, w12382, w12383, w12384, w12385, w12386, w12387, w12388, w12389, w12390, w12391, w12392, w12393, w12394, w12395, w12396, w12397, w12398, w12399, w12400, w12401, w12402, w12403, w12404, w12405, w12406, w12407, w12408, w12409, w12410, w12411, w12412, w12413, w12414, w12415, w12416, w12417, w12418, w12419, w12420, w12421, w12422, w12423, w12424, w12425, w12426, w12427, w12428, w12429, w12430, w12431, w12432, w12433, w12434, w12435, w12436, w12437, w12438, w12439, w12440, w12441, w12442, w12443, w12444, w12445, w12446, w12447, w12448, w12449, w12450, w12451, w12452, w12453, w12454, w12455, w12456, w12457, w12458, w12459, w12460, w12461, w12462, w12463, w12464, w12465, w12466, w12467, w12468, w12469, w12470, w12471, w12472, w12473, w12474, w12475, w12476, w12477, w12478, w12479, w12480, w12481, w12482, w12483, w12484, w12485, w12486, w12487, w12488, w12489, w12490, w12491, w12492, w12493, w12494, w12495, w12496, w12497, w12498, w12499, w12500, w12501, w12502, w12503, w12504, w12505, w12506, w12507, w12508, w12509, w12510, w12511, w12512, w12513, w12514, w12515, w12516, w12517, w12518, w12519, w12520, w12521, w12522, w12523, w12524, w12525, w12526, w12527, w12528, w12529, w12530, w12531, w12532, w12533, w12534, w12535, w12536, w12537, w12538, w12539, w12540, w12541, w12542, w12543, w12544, w12545, w12546, w12547, w12548, w12549, w12550, w12551, w12552, w12553, w12554, w12555, w12556, w12557, w12558, w12559, w12560, w12561, w12562, w12563, w12564, w12565, w12566, w12567, w12568, w12569, w12570, w12571, w12572, w12573, w12574, w12575, w12576, w12577, w12578, w12579, w12580, w12581, w12582, w12583, w12584, w12585, w12586, w12587, w12588, w12589, w12590, w12591, w12592, w12593, w12594, w12595, w12596, w12597, w12598, w12599, w12600, w12601, w12602, w12603, w12604, w12605, w12606, w12607, w12608, w12609, w12610, w12611, w12612, w12613, w12614, w12615, w12616, w12617, w12618, w12619, w12620, w12621, w12622, w12623, w12624, w12625, w12626, w12627, w12628, w12629, w12630, w12631, w12632, w12633, w12634, w12635, w12636, w12637, w12638, w12639, w12640, w12641, w12642, w12643, w12644, w12645, w12646, w12647, w12648, w12649, w12650, w12651, w12652, w12653, w12654, w12655, w12656, w12657, w12658, w12659, w12660, w12661, w12662, w12663, w12664, w12665, w12666, w12667, w12668, w12669, w12670, w12671, w12672, w12673, w12674, w12675, w12676, w12677, w12678, w12679, w12680, w12681, w12682, w12683, w12684, w12685, w12686, w12687, w12688, w12689, w12690, w12691, w12692, w12693, w12694, w12695, w12696, w12697, w12698, w12699, w12700, w12701, w12702, w12703, w12704, w12705, w12706, w12707, w12708, w12709, w12710, w12711, w12712, w12713, w12714, w12715, w12716, w12717, w12718, w12719, w12720, w12721, w12722, w12723, w12724, w12725, w12726, w12727, w12728, w12729, w12730, w12731, w12732, w12733, w12734, w12735, w12736, w12737, w12738, w12739, w12740, w12741, w12742, w12743, w12744, w12745, w12746, w12747, w12748, w12749, w12750, w12751, w12752, w12753, w12754, w12755, w12756, w12757, w12758, w12759, w12760, w12761, w12762, w12763, w12764, w12765, w12766, w12767, w12768, w12769, w12770, w12771, w12772, w12773, w12774, w12775, w12776, w12777, w12778, w12779, w12780, w12781, w12782, w12783, w12784, w12785, w12786, w12787, w12788, w12789, w12790, w12791, w12792, w12793, w12794, w12795, w12796, w12797, w12798, w12799, w12800, w12801, w12802, w12803, w12804, w12805, w12806, w12807, w12808, w12809, w12810, w12811, w12812, w12813, w12814, w12815, w12816, w12817, w12818, w12819, w12820, w12821, w12822, w12823, w12824, w12825, w12826, w12827, w12828, w12829, w12830, w12831, w12832, w12833, w12834, w12835, w12836, w12837, w12838, w12839, w12840, w12841, w12842, w12843, w12844, w12845, w12846, w12847, w12848, w12849, w12850, w12851, w12852, w12853, w12854, w12855, w12856, w12857, w12858, w12859, w12860, w12861, w12862, w12863, w12864, w12865, w12866, w12867, w12868, w12869, w12870, w12871, w12872, w12873, w12874, w12875, w12876, w12877, w12878, w12879, w12880, w12881, w12882, w12883, w12884, w12885, w12886, w12887, w12888, w12889, w12890, w12891, w12892, w12893, w12894, w12895, w12896, w12897, w12898, w12899, w12900, w12901, w12902, w12903, w12904, w12905, w12906, w12907, w12908, w12909, w12910, w12911, w12912, w12913, w12914, w12915, w12916, w12917, w12918, w12919, w12920, w12921, w12922, w12923, w12924, w12925, w12926, w12927, w12928, w12929, w12930, w12931, w12932, w12933, w12934, w12935, w12936, w12937, w12938, w12939, w12940, w12941, w12942, w12943, w12944, w12945, w12946, w12947, w12948, w12949, w12950, w12951, w12952, w12953, w12954, w12955, w12956, w12957, w12958, w12959, w12960, w12961, w12962, w12963, w12964, w12965, w12966, w12967, w12968, w12969, w12970, w12971, w12972, w12973, w12974, w12975, w12976, w12977, w12978, w12979, w12980, w12981, w12982, w12983, w12984, w12985, w12986, w12987, w12988, w12989, w12990, w12991, w12992, w12993, w12994, w12995, w12996, w12997, w12998, w12999, w13000, w13001, w13002, w13003, w13004, w13005, w13006, w13007, w13008, w13009, w13010, w13011, w13012, w13013, w13014, w13015, w13016, w13017, w13018, w13019, w13020, w13021, w13022, w13023, w13024, w13025, w13026, w13027, w13028, w13029, w13030, w13031, w13032, w13033, w13034, w13035, w13036, w13037, w13038, w13039, w13040, w13041, w13042, w13043, w13044, w13045, w13046, w13047, w13048, w13049, w13050, w13051, w13052, w13053, w13054, w13055, w13056, w13057, w13058, w13059, w13060, w13061, w13062, w13063, w13064, w13065, w13066, w13067, w13068, w13069, w13070, w13071, w13072, w13073, w13074, w13075, w13076, w13077, w13078, w13079, w13080, w13081, w13082, w13083, w13084, w13085, w13086, w13087, w13088, w13089, w13090, w13091, w13092, w13093, w13094, w13095, w13096, w13097, w13098, w13099, w13100, w13101, w13102, w13103, w13104, w13105, w13106, w13107, w13108, w13109, w13110, w13111, w13112, w13113, w13114, w13115, w13116, w13117, w13118, w13119, w13120, w13121, w13122, w13123, w13124, w13125, w13126, w13127, w13128, w13129, w13130, w13131, w13132, w13133, w13134, w13135, w13136, w13137, w13138, w13139, w13140, w13141, w13142, w13143, w13144, w13145, w13146, w13147, w13148, w13149, w13150, w13151, w13152, w13153, w13154, w13155, w13156, w13157, w13158, w13159, w13160, w13161, w13162, w13163, w13164, w13165, w13166, w13167, w13168, w13169, w13170, w13171, w13172, w13173, w13174, w13175, w13176, w13177, w13178, w13179, w13180, w13181, w13182, w13183, w13184, w13185, w13186, w13187, w13188, w13189, w13190, w13191, w13192, w13193, w13194, w13195, w13196, w13197, w13198, w13199, w13200, w13201, w13202, w13203, w13204, w13205, w13206, w13207, w13208, w13209, w13210, w13211, w13212, w13213, w13214, w13215, w13216, w13217, w13218, w13219, w13220, w13221, w13222, w13223, w13224, w13225, w13226, w13227, w13228, w13229, w13230, w13231, w13232, w13233, w13234, w13235, w13236, w13237, w13238, w13239, w13240, w13241, w13242, w13243, w13244, w13245, w13246, w13247, w13248, w13249, w13250, w13251, w13252, w13253, w13254, w13255, w13256, w13257, w13258, w13259, w13260, w13261, w13262, w13263, w13264, w13265, w13266, w13267, w13268, w13269, w13270, w13271, w13272, w13273, w13274, w13275, w13276, w13277, w13278, w13279, w13280, w13281, w13282, w13283, w13284, w13285, w13286, w13287, w13288, w13289, w13290, w13291, w13292, w13293, w13294, w13295, w13296, w13297, w13298, w13299, w13300, w13301, w13302, w13303, w13304, w13305, w13306, w13307, w13308, w13309, w13310, w13311, w13312, w13313, w13314, w13315, w13316, w13317, w13318, w13319, w13320, w13321, w13322, w13323, w13324, w13325, w13326, w13327, w13328, w13329, w13330, w13331, w13332, w13333, w13334, w13335, w13336, w13337, w13338, w13339, w13340, w13341, w13342, w13343, w13344, w13345, w13346, w13347, w13348, w13349, w13350, w13351, w13352, w13353, w13354, w13355, w13356, w13357, w13358, w13359, w13360, w13361, w13362, w13363, w13364, w13365, w13366, w13367, w13368, w13369, w13370, w13371, w13372, w13373, w13374, w13375, w13376, w13377, w13378, w13379, w13380, w13381, w13382, w13383, w13384, w13385, w13386, w13387, w13388, w13389, w13390, w13391, w13392, w13393, w13394, w13395, w13396, w13397, w13398, w13399, w13400, w13401, w13402, w13403, w13404, w13405, w13406, w13407, w13408, w13409, w13410, w13411, w13412, w13413, w13414, w13415, w13416, w13417, w13418, w13419, w13420, w13421, w13422, w13423, w13424, w13425, w13426, w13427, w13428, w13429, w13430, w13431, w13432, w13433, w13434, w13435, w13436, w13437, w13438, w13439, w13440, w13441, w13442, w13443, w13444, w13445, w13446, w13447, w13448, w13449, w13450, w13451, w13452, w13453, w13454, w13455, w13456, w13457, w13458, w13459, w13460, w13461, w13462, w13463, w13464, w13465, w13466, w13467, w13468, w13469, w13470, w13471, w13472, w13473, w13474, w13475, w13476, w13477, w13478, w13479, w13480, w13481, w13482, w13483, w13484, w13485, w13486, w13487, w13488, w13489, w13490, w13491, w13492, w13493, w13494, w13495, w13496, w13497, w13498, w13499, w13500, w13501, w13502, w13503, w13504, w13505, w13506, w13507, w13508, w13509, w13510, w13511, w13512, w13513, w13514, w13515, w13516, w13517, w13518, w13519, w13520, w13521, w13522, w13523, w13524, w13525, w13526, w13527, w13528, w13529, w13530, w13531, w13532, w13533, w13534, w13535, w13536, w13537, w13538, w13539, w13540, w13541, w13542, w13543, w13544, w13545, w13546, w13547, w13548, w13549, w13550, w13551, w13552, w13553, w13554, w13555, w13556, w13557, w13558, w13559, w13560, w13561, w13562, w13563, w13564, w13565, w13566, w13567, w13568, w13569, w13570, w13571, w13572, w13573, w13574, w13575, w13576, w13577, w13578, w13579, w13580, w13581, w13582, w13583, w13584, w13585, w13586, w13587, w13588, w13589, w13590, w13591, w13592, w13593, w13594, w13595, w13596, w13597, w13598, w13599, w13600, w13601, w13602, w13603, w13604, w13605, w13606, w13607, w13608, w13609, w13610, w13611, w13612, w13613, w13614, w13615, w13616, w13617, w13618, w13619, w13620, w13621, w13622, w13623, w13624, w13625, w13626, w13627, w13628, w13629, w13630, w13631, w13632, w13633, w13634, w13635, w13636, w13637, w13638, w13639, w13640, w13641, w13642, w13643, w13644, w13645, w13646, w13647, w13648, w13649, w13650, w13651, w13652, w13653, w13654, w13655, w13656, w13657, w13658, w13659, w13660, w13661, w13662, w13663, w13664, w13665, w13666, w13667, w13668, w13669, w13670, w13671, w13672, w13673, w13674, w13675, w13676, w13677, w13678, w13679, w13680, w13681, w13682, w13683, w13684, w13685, w13686, w13687, w13688, w13689, w13690, w13691, w13692, w13693, w13694, w13695, w13696, w13697, w13698, w13699, w13700, w13701, w13702, w13703, w13704, w13705, w13706, w13707, w13708, w13709, w13710, w13711, w13712, w13713, w13714, w13715, w13716, w13717, w13718, w13719, w13720, w13721, w13722, w13723, w13724, w13725, w13726, w13727, w13728, w13729, w13730, w13731, w13732, w13733, w13734, w13735, w13736, w13737, w13738, w13739, w13740, w13741, w13742, w13743, w13744, w13745, w13746, w13747, w13748, w13749, w13750, w13751, w13752, w13753, w13754, w13755, w13756, w13757, w13758, w13759, w13760, w13761, w13762, w13763, w13764, w13765, w13766, w13767, w13768, w13769, w13770, w13771, w13772, w13773, w13774, w13775, w13776, w13777, w13778, w13779, w13780, w13781, w13782, w13783, w13784, w13785, w13786, w13787, w13788, w13789, w13790, w13791, w13792, w13793, w13794, w13795, w13796, w13797, w13798, w13799, w13800, w13801, w13802, w13803, w13804, w13805, w13806, w13807, w13808, w13809, w13810, w13811, w13812, w13813, w13814, w13815, w13816, w13817, w13818, w13819, w13820, w13821, w13822, w13823, w13824, w13825, w13826, w13827, w13828, w13829, w13830, w13831, w13832, w13833, w13834, w13835, w13836, w13837, w13838, w13839, w13840, w13841, w13842, w13843, w13844, w13845, w13846, w13847, w13848, w13849, w13850, w13851, w13852, w13853, w13854, w13855, w13856, w13857, w13858, w13859, w13860, w13861, w13862, w13863, w13864, w13865, w13866, w13867, w13868, w13869, w13870, w13871, w13872, w13873, w13874, w13875, w13876, w13877, w13878, w13879, w13880, w13881, w13882, w13883, w13884, w13885, w13886, w13887, w13888, w13889, w13890, w13891, w13892, w13893, w13894, w13895, w13896, w13897, w13898, w13899, w13900, w13901, w13902, w13903, w13904, w13905, w13906, w13907, w13908, w13909, w13910, w13911, w13912, w13913, w13914, w13915, w13916, w13917, w13918, w13919, w13920, w13921, w13922, w13923, w13924, w13925, w13926, w13927, w13928, w13929, w13930, w13931, w13932, w13933, w13934, w13935, w13936, w13937, w13938, w13939, w13940, w13941, w13942, w13943, w13944, w13945, w13946, w13947, w13948, w13949, w13950, w13951, w13952, w13953, w13954, w13955, w13956, w13957, w13958, w13959, w13960, w13961, w13962, w13963, w13964, w13965, w13966, w13967, w13968, w13969, w13970, w13971, w13972, w13973, w13974, w13975, w13976, w13977, w13978, w13979, w13980, w13981, w13982, w13983, w13984, w13985, w13986, w13987, w13988, w13989, w13990, w13991, w13992, w13993, w13994, w13995, w13996, w13997, w13998, w13999, w14000, w14001, w14002, w14003, w14004, w14005, w14006, w14007, w14008, w14009, w14010, w14011, w14012, w14013, w14014, w14015, w14016, w14017, w14018, w14019, w14020, w14021, w14022, w14023, w14024, w14025, w14026, w14027, w14028, w14029, w14030, w14031, w14032, w14033, w14034, w14035, w14036, w14037, w14038, w14039, w14040, w14041, w14042, w14043, w14044, w14045, w14046, w14047, w14048, w14049, w14050, w14051, w14052, w14053, w14054, w14055, w14056, w14057, w14058, w14059, w14060, w14061, w14062, w14063, w14064, w14065, w14066, w14067, w14068, w14069, w14070, w14071, w14072, w14073, w14074, w14075, w14076, w14077, w14078, w14079, w14080, w14081, w14082, w14083, w14084, w14085, w14086, w14087, w14088, w14089, w14090, w14091, w14092, w14093, w14094, w14095, w14096, w14097, w14098, w14099, w14100, w14101, w14102, w14103, w14104, w14105, w14106, w14107, w14108, w14109, w14110, w14111, w14112, w14113, w14114, w14115, w14116, w14117, w14118, w14119, w14120, w14121, w14122, w14123, w14124, w14125, w14126, w14127, w14128, w14129, w14130, w14131, w14132, w14133, w14134, w14135, w14136, w14137, w14138, w14139, w14140, w14141, w14142, w14143, w14144, w14145, w14146, w14147, w14148, w14149, w14150, w14151, w14152, w14153, w14154, w14155, w14156, w14157, w14158, w14159, w14160, w14161, w14162, w14163, w14164, w14165, w14166, w14167, w14168, w14169, w14170, w14171, w14172, w14173, w14174, w14175, w14176, w14177, w14178, w14179, w14180, w14181, w14182, w14183, w14184, w14185, w14186, w14187, w14188, w14189, w14190, w14191, w14192, w14193, w14194, w14195, w14196, w14197, w14198, w14199, w14200, w14201, w14202, w14203, w14204, w14205, w14206, w14207, w14208, w14209, w14210, w14211, w14212, w14213, w14214, w14215, w14216, w14217, w14218, w14219, w14220, w14221, w14222, w14223, w14224, w14225, w14226, w14227, w14228, w14229, w14230, w14231, w14232, w14233, w14234, w14235, w14236, w14237, w14238, w14239, w14240, w14241, w14242, w14243, w14244, w14245, w14246, w14247, w14248, w14249, w14250, w14251, w14252, w14253, w14254, w14255, w14256, w14257, w14258, w14259, w14260, w14261, w14262, w14263, w14264, w14265, w14266, w14267, w14268, w14269, w14270, w14271, w14272, w14273, w14274, w14275, w14276, w14277, w14278, w14279, w14280, w14281, w14282, w14283, w14284, w14285, w14286, w14287, w14288, w14289, w14290, w14291, w14292, w14293, w14294, w14295, w14296, w14297, w14298, w14299, w14300, w14301, w14302, w14303, w14304, w14305, w14306, w14307, w14308, w14309, w14310, w14311, w14312, w14313, w14314, w14315, w14316, w14317, w14318, w14319, w14320, w14321, w14322, w14323, w14324, w14325, w14326, w14327, w14328, w14329, w14330, w14331, w14332, w14333, w14334, w14335, w14336, w14337, w14338, w14339, w14340, w14341, w14342, w14343, w14344, w14345, w14346, w14347, w14348, w14349, w14350, w14351, w14352, w14353, w14354, w14355, w14356, w14357, w14358, w14359, w14360, w14361, w14362, w14363, w14364, w14365, w14366, w14367, w14368, w14369, w14370, w14371, w14372, w14373, w14374, w14375, w14376, w14377, w14378, w14379, w14380, w14381, w14382, w14383, w14384, w14385, w14386, w14387, w14388, w14389, w14390, w14391, w14392, w14393, w14394, w14395, w14396, w14397, w14398, w14399, w14400, w14401, w14402, w14403, w14404, w14405, w14406, w14407, w14408, w14409, w14410, w14411, w14412, w14413, w14414, w14415, w14416, w14417, w14418, w14419, w14420, w14421, w14422, w14423, w14424, w14425, w14426, w14427, w14428, w14429, w14430, w14431, w14432, w14433, w14434, w14435, w14436, w14437, w14438, w14439, w14440, w14441, w14442, w14443, w14444, w14445, w14446, w14447, w14448, w14449, w14450, w14451, w14452, w14453, w14454, w14455, w14456, w14457, w14458, w14459, w14460, w14461, w14462, w14463, w14464, w14465, w14466, w14467, w14468, w14469, w14470, w14471, w14472, w14473, w14474, w14475, w14476, w14477, w14478, w14479, w14480, w14481, w14482, w14483, w14484, w14485, w14486, w14487, w14488, w14489, w14490, w14491, w14492, w14493, w14494, w14495, w14496, w14497, w14498, w14499, w14500, w14501, w14502, w14503, w14504, w14505, w14506, w14507, w14508, w14509, w14510, w14511, w14512, w14513, w14514, w14515, w14516, w14517, w14518, w14519, w14520, w14521, w14522, w14523, w14524, w14525, w14526, w14527, w14528, w14529, w14530, w14531, w14532, w14533, w14534, w14535, w14536, w14537, w14538, w14539, w14540, w14541, w14542, w14543, w14544, w14545, w14546, w14547, w14548, w14549, w14550, w14551, w14552, w14553, w14554, w14555, w14556, w14557, w14558, w14559, w14560, w14561, w14562, w14563, w14564, w14565, w14566, w14567, w14568, w14569, w14570, w14571, w14572, w14573, w14574, w14575, w14576, w14577, w14578, w14579, w14580, w14581, w14582, w14583, w14584, w14585, w14586, w14587, w14588, w14589, w14590, w14591, w14592, w14593, w14594, w14595, w14596, w14597, w14598, w14599, w14600, w14601, w14602, w14603, w14604, w14605, w14606, w14607, w14608, w14609, w14610, w14611, w14612, w14613, w14614, w14615, w14616, w14617, w14618, w14619, w14620, w14621, w14622, w14623, w14624, w14625, w14626, w14627, w14628, w14629, w14630, w14631, w14632, w14633, w14634, w14635, w14636, w14637, w14638, w14639, w14640, w14641, w14642, w14643, w14644, w14645, w14646, w14647, w14648, w14649, w14650, w14651, w14652, w14653, w14654, w14655, w14656, w14657, w14658, w14659, w14660, w14661, w14662, w14663, w14664, w14665, w14666, w14667, w14668, w14669, w14670, w14671;
assign w0 = ~w12825 & w10256;
assign w1 = w4213 & w12868;
assign w2 = (~w10926 & ~w8659) | (~w10926 & w4511) | (~w8659 & w4511);
assign w3 = w3383 & ~w11516;
assign w4 = w14280 & w2938;
assign w5 = ~w5522 & ~w11934;
assign w6 = ~w5005 & w10483;
assign w7 = (~w6387 & w11354) | (~w6387 & w8029) | (w11354 & w8029);
assign w8 = ~w2387 & ~w9940;
assign w9 = (w10704 & ~w12614) | (w10704 & w4825) | (~w12614 & w4825);
assign w10 = ~w5997 & w3656;
assign w11 = ~w5 & ~w13429;
assign w12 = (~w10075 & w499) | (~w10075 & w13848) | (w499 & w13848);
assign w13 = (~w8396 & w1426) | (~w8396 & w11591) | (w1426 & w11591);
assign w14 = ~w8171 & ~w4269;
assign w15 = ~w11117 & w3017;
assign w16 = w7889 & w3963;
assign w17 = ~w9000 & w5452;
assign w18 = w8186 & w9092;
assign w19 = ~w5422 & w3645;
assign w20 = w12122 & w14327;
assign w21 = ~w14054 & w12107;
assign w22 = (~w14114 & w6712) | (~w14114 & w6884) | (w6712 & w6884);
assign w23 = (~w2599 & ~w8389) | (~w2599 & w2215) | (~w8389 & w2215);
assign w24 = (w7123 & w10061) | (w7123 & ~w2362) | (w10061 & ~w2362);
assign w25 = w8626 & ~w9244;
assign w26 = (w9541 & w2740) | (w9541 & w9778) | (w2740 & w9778);
assign w27 = ~w1542 & ~w12591;
assign w28 = ~w6689 & w3288;
assign w29 = ~w1166 & w199;
assign w30 = w1270 & ~w13807;
assign w31 = ~w7455 & w10075;
assign w32 = (~w9608 & w14112) | (~w9608 & w12507) | (w14112 & w12507);
assign w33 = ~w10602 & ~w8122;
assign w34 = ~w3410 & w12047;
assign w35 = ~w4261 & w13431;
assign w36 = ~w8691 & ~w10408;
assign w37 = ~w1840 & ~w9523;
assign w38 = w8450 & w14181;
assign w39 = w33 & w5975;
assign w40 = w13713 & w3734;
assign w41 = (w5952 & w3093) | (w5952 & w10527) | (w3093 & w10527);
assign w42 = ~w8009 & ~w13981;
assign w43 = (w6708 & w13742) | (w6708 & w2075) | (w13742 & w2075);
assign w44 = w3927 & w4947;
assign w45 = b71 & a71;
assign w46 = (~w4287 & w2971) | (~w4287 & ~w7644) | (w2971 & ~w7644);
assign w47 = (w10637 & w9700) | (w10637 & w307) | (w9700 & w307);
assign w48 = w11628 & w9481;
assign w49 = w4819 & w11071;
assign w50 = ~b12 & ~a12;
assign w51 = ~w7376 & w10075;
assign w52 = ~w7437 & w1692;
assign w53 = (w378 & w14599) | (w378 & w9729) | (w14599 & w9729);
assign w54 = w183 & w14072;
assign w55 = w13360 & ~w1919;
assign w56 = (~w14463 & w11182) | (~w14463 & w13433) | (w11182 & w13433);
assign w57 = w8195 & w11190;
assign w58 = (w1758 & ~w9608) | (w1758 & w5659) | (~w9608 & w5659);
assign w59 = (w5115 & w12810) | (w5115 & w5310) | (w12810 & w5310);
assign w60 = (w6502 & ~w4213) | (w6502 & w6322) | (~w4213 & w6322);
assign w61 = ~w1588 & w9604;
assign w62 = w6101 & w14389;
assign w63 = (w8 & w13819) | (w8 & w14455) | (w13819 & w14455);
assign w64 = ~w13222 & ~w2850;
assign w65 = w9655 & w1387;
assign w66 = w10676 & ~w14070;
assign w67 = w2291 & ~w12893;
assign w68 = w8589 & ~w9411;
assign w69 = ~w829 & w7914;
assign w70 = (w10254 & w2966) | (w10254 & w715) | (w2966 & w715);
assign w71 = (~w1520 & w1490) | (~w1520 & w10971) | (w1490 & w10971);
assign w72 = ~w9083 & ~w12580;
assign w73 = (~w1162 & w12326) | (~w1162 & w12628) | (w12326 & w12628);
assign w74 = w9999 & ~w11629;
assign w75 = (~w1873 & w7630) | (~w1873 & w5307) | (w7630 & w5307);
assign w76 = (w13896 & w6506) | (w13896 & w2022) | (w6506 & w2022);
assign w77 = ~w852 & ~w3025;
assign w78 = (w4359 & w4512) | (w4359 & w113) | (w4512 & w113);
assign w79 = (w6819 & w12596) | (w6819 & ~w11732) | (w12596 & ~w11732);
assign w80 = ~w10435 & w7516;
assign w81 = (w10997 & w13122) | (w10997 & w617) | (w13122 & w617);
assign w82 = ~w9086 & w7796;
assign w83 = ~w11298 & ~w4267;
assign w84 = ~w8220 & w11983;
assign w85 = w3914 & w11902;
assign w86 = ~w14565 & ~w810;
assign w87 = (w13713 & ~w7464) | (w13713 & w4466) | (~w7464 & w4466);
assign w88 = w2387 & w9940;
assign w89 = (~w14395 & w2500) | (~w14395 & w5262) | (w2500 & w5262);
assign w90 = ~w1563 & w4587;
assign w91 = (w2698 & w5875) | (w2698 & w7901) | (w5875 & w7901);
assign w92 = ~w11572 & ~w5677;
assign w93 = (w6970 & w8821) | (w6970 & ~w3798) | (w8821 & ~w3798);
assign w94 = (w6427 & w7741) | (w6427 & w14261) | (w7741 & w14261);
assign w95 = ~w5495 & ~w2782;
assign w96 = w1925 & ~w6755;
assign w97 = w11746 & w9603;
assign w98 = w12271 & w10317;
assign w99 = (~w1694 & w7376) | (~w1694 & w4862) | (w7376 & w4862);
assign w100 = (~w13256 & w4982) | (~w13256 & w12247) | (w4982 & w12247);
assign w101 = ~w7253 & ~w527;
assign w102 = (~w3550 & w7564) | (~w3550 & w7176) | (w7564 & w7176);
assign w103 = (w6885 & w7419) | (w6885 & w12536) | (w7419 & w12536);
assign w104 = w3563 & ~w9121;
assign w105 = w11097 & ~w1821;
assign w106 = ~w8512 & w12533;
assign w107 = ~w2680 & ~w10075;
assign w108 = w499 & ~w6935;
assign w109 = w11049 & ~w3427;
assign w110 = w636 & ~w3963;
assign w111 = ~w2926 & w2986;
assign w112 = ~w13713 & w1114;
assign w113 = w5294 & w4359;
assign w114 = ~w13256 & ~w3587;
assign w115 = ~w12659 & ~w1533;
assign w116 = ~w7452 & w3904;
assign w117 = w7453 & w3904;
assign w118 = ~w5522 & ~w13323;
assign w119 = w11395 & w5397;
assign w120 = (w10123 & w14025) | (w10123 & w14522) | (w14025 & w14522);
assign w121 = w7001 & w7670;
assign w122 = (~w2159 & w2144) | (~w2159 & w3179) | (w2144 & w3179);
assign w123 = ~w3098 & ~w8975;
assign w124 = ~w11261 & w9448;
assign w125 = w9613 & ~w6442;
assign w126 = w9480 & ~w11031;
assign w127 = ~w13451 & w3988;
assign w128 = ~w10257 & w3754;
assign w129 = w3576 & ~w4841;
assign w130 = ~w6427 & w9471;
assign w131 = ~w10244 & ~w2552;
assign w132 = (w13323 & ~w5731) | (w13323 & w13855) | (~w5731 & w13855);
assign w133 = ~w8086 & w3557;
assign w134 = w4359 & ~w5664;
assign w135 = w10676 & w9938;
assign w136 = w5732 & w10855;
assign w137 = ~w3751 & ~w8120;
assign w138 = ~w5089 & ~w6312;
assign w139 = (~w1639 & ~w10923) | (~w1639 & ~w12154) | (~w10923 & ~w12154);
assign w140 = w7712 & w11791;
assign w141 = w6641 & w11099;
assign w142 = b96 & a96;
assign w143 = (~w2663 & w8742) | (~w2663 & w13281) | (w8742 & w13281);
assign w144 = (~w13654 & w8495) | (~w13654 & w8126) | (w8495 & w8126);
assign w145 = ~w922 & w3611;
assign w146 = ~w3151 & w13887;
assign w147 = (~w217 & ~w10482) | (~w217 & w7036) | (~w10482 & w7036);
assign w148 = (w7922 & w14176) | (w7922 & w9575) | (w14176 & w9575);
assign w149 = ~w5619 & w3574;
assign w150 = w607 & ~w646;
assign w151 = w5732 & w11395;
assign w152 = ~w14184 & ~w1101;
assign w153 = w6097 & w11552;
assign w154 = (w7041 & w2854) | (w7041 & w4684) | (w2854 & w4684);
assign w155 = w8396 & ~w7889;
assign w156 = w360 & ~w13820;
assign w157 = ~w2570 & ~w9939;
assign w158 = ~w4756 & w12080;
assign w159 = ~w4575 & ~w5982;
assign w160 = (w13713 & ~w7464) | (w13713 & w14151) | (~w7464 & w14151);
assign w161 = ~w14441 & w7069;
assign w162 = w4484 & ~w6964;
assign w163 = w7365 & w8992;
assign w164 = ~w2680 & w5196;
assign w165 = w9433 & ~w7423;
assign w166 = ~w8019 & ~w5282;
assign w167 = ~w12903 & w13414;
assign w168 = w7670 & w3194;
assign w169 = ~w7782 & w8881;
assign w170 = ~w71 & w11660;
assign w171 = w11355 | ~w9989;
assign w172 = w741 & w12932;
assign w173 = ~w9244 & w6381;
assign w174 = w2881 & ~w12182;
assign w175 = ~a127 & ~b127;
assign w176 = w7177 & ~w12778;
assign w177 = ~w2572 & w10277;
assign w178 = w1876 & w9542;
assign w179 = (~w10850 & ~w8556) | (~w10850 & ~w7690) | (~w8556 & ~w7690);
assign w180 = ~w13324 & w14653;
assign w181 = ~w11905 & w3169;
assign w182 = (w11416 & w1685) | (w11416 & w5802) | (w1685 & w5802);
assign w183 = ~w2839 & ~w5305;
assign w184 = w4367 & ~w10584;
assign w185 = ~w13854 & ~w1809;
assign w186 = w9995 & w12706;
assign w187 = w12038 & w4195;
assign w188 = ~w11811 & ~w2417;
assign w189 = ~w636 & w3963;
assign w190 = ~w5521 & ~w8327;
assign w191 = w11726 & ~w6211;
assign w192 = (~w11838 & w13597) | (~w11838 & w2934) | (w13597 & w2934);
assign w193 = ~w11080 & ~w7146;
assign w194 = ~w14195 & w5127;
assign w195 = ~w13126 & ~w2823;
assign w196 = ~w7662 & w8992;
assign w197 = w5865 & ~w4494;
assign w198 = w12371 & ~w3904;
assign w199 = w3611 & w9265;
assign w200 = ~w7369 & ~w14614;
assign w201 = (~w11483 & w9621) | (~w11483 & w2184) | (w9621 & w2184);
assign w202 = w8426 | w3452;
assign w203 = ~w6436 & ~w2941;
assign w204 = w2737 & w665;
assign w205 = ~w2250 & ~w2828;
assign w206 = ~w1343 & ~w13534;
assign w207 = (~w1260 & ~w9541) | (~w1260 & w14584) | (~w9541 & w14584);
assign w208 = w13426 & w12642;
assign w209 = w13189 & ~w10699;
assign w210 = ~w4050 & w3110;
assign w211 = ~w4032 & w199;
assign w212 = (~w7515 & w10724) | (~w7515 & w24) | (w10724 & w24);
assign w213 = ~w6735 & ~w1990;
assign w214 = w5613 & w11506;
assign w215 = w13282 & w13854;
assign w216 = ~w4665 & ~w5844;
assign w217 = ~w3885 & ~w325;
assign w218 = ~w14072 & ~w3435;
assign w219 = ~w142 & ~w5761;
assign w220 = w11934 & w7889;
assign w221 = ~w12464 & w12893;
assign w222 = (w5927 & w12864) | (w5927 & w9709) | (w12864 & w9709);
assign w223 = (w9264 & w14664) | (w9264 & w8132) | (w14664 & w8132);
assign w224 = ~w922 & w247;
assign w225 = (w13924 & ~w4032) | (w13924 & w709) | (~w4032 & w709);
assign w226 = (~w254 & w5847) | (~w254 & w7055) | (w5847 & w7055);
assign w227 = w1186 & ~w11434;
assign w228 = (w8176 & w13858) | (w8176 & w12297) | (w13858 & w12297);
assign w229 = ~w4810 & ~w406;
assign w230 = ~w10191 & w7882;
assign w231 = ~w5447 & ~w11238;
assign w232 = (~w7684 & w6623) | (~w7684 & w10667) | (w6623 & w10667);
assign w233 = ~w4921 & w3600;
assign w234 = w880 & w6704;
assign w235 = ~b41 & ~a41;
assign w236 = ~w4078 & w14212;
assign w237 = (~w11756 & w14506) | (~w11756 & w12588) | (w14506 & w12588);
assign w238 = (~w7589 & w9213) | (~w7589 & w1233) | (w9213 & w1233);
assign w239 = ~w3963 & ~w2509;
assign w240 = ~w5664 & ~w6141;
assign w241 = w6979 & ~w4290;
assign w242 = (w976 & w8515) | (w976 & ~w8444) | (w8515 & ~w8444);
assign w243 = w8072 & w3373;
assign w244 = ~w13182 & ~w1487;
assign w245 = w347 & ~w1929;
assign w246 = w9534 & w9950;
assign w247 = w10045 & w14048;
assign w248 = ~w5461 & w7432;
assign w249 = w4467 & ~w4170;
assign w250 = (w14346 & w9746) | (w14346 & ~w5007) | (w9746 & ~w5007);
assign w251 = (w5828 & w3485) | (w5828 & w9733) | (w3485 & w9733);
assign w252 = (w6230 & w5543) | (w6230 & w8260) | (w5543 & w8260);
assign w253 = ~w12483 & ~w11959;
assign w254 = w11949 & ~w11373;
assign w255 = (w11993 & w2754) | (w11993 & ~w1430) | (w2754 & ~w1430);
assign w256 = (~w13375 & ~w5498) | (~w13375 & w9403) | (~w5498 & w9403);
assign w257 = (~w5237 & w6633) | (~w5237 & w3397) | (w6633 & w3397);
assign w258 = (w12135 & w7645) | (w12135 & w1092) | (w7645 & w1092);
assign w259 = ~w11817 & w1272;
assign w260 = (~w3075 & w9252) | (~w3075 & w14303) | (w9252 & w14303);
assign w261 = w7244 & w7670;
assign w262 = w13358 & ~w4111;
assign w263 = ~w1873 & w13863;
assign w264 = (w13980 & w7123) | (w13980 & w10061) | (w7123 & w10061);
assign w265 = ~w6975 & ~w13902;
assign w266 = w1692 & ~w2783;
assign w267 = w7596 & w7969;
assign w268 = w647 & ~w3827;
assign w269 = w11732 & w14506;
assign w270 = (w3957 & ~w13282) | (w3957 & w12058) | (~w13282 & w12058);
assign w271 = (~w6462 & w6024) | (~w6462 & w10401) | (w6024 & w10401);
assign w272 = (~w11261 & w1363) | (~w11261 & w10723) | (w1363 & w10723);
assign w273 = ~w2317 & w13138;
assign w274 = ~w9805 & ~w6817;
assign w275 = (w12376 & w3624) | (w12376 & w3837) | (w3624 & w3837);
assign w276 = w4561 & ~w7566;
assign w277 = w3035 & w5784;
assign w278 = ~w14038 & ~w8013;
assign w279 = w11899 & ~w6250;
assign w280 = (w11385 & w5958) | (w11385 & w6909) | (w5958 & w6909);
assign w281 = w2302 & w5616;
assign w282 = (~w11973 & w5653) | (~w11973 & w14014) | (w5653 & w14014);
assign w283 = w6190 & w4111;
assign w284 = ~w10343 & w12460;
assign w285 = ~w7376 & ~w11411;
assign w286 = w5522 & w5761;
assign w287 = ~w5827 & w137;
assign w288 = ~w7267 & ~w993;
assign w289 = (w14463 & w5646) | (w14463 & w823) | (w5646 & w823);
assign w290 = (w9528 & w523) | (w9528 & w11984) | (w523 & w11984);
assign w291 = ~w8694 & w10808;
assign w292 = w8964 & ~w2571;
assign w293 = ~w7867 & ~w10317;
assign w294 = ~w6573 & ~w2064;
assign w295 = ~w2752 & ~w1766;
assign w296 = (w11708 & w2226) | (w11708 & w9785) | (w2226 & w9785);
assign w297 = w11488 & ~w4541;
assign w298 = ~w3611 & ~w9583;
assign w299 = (w1150 & w7150) | (w1150 & w6452) | (w7150 & w6452);
assign w300 = w554 & ~w12731;
assign w301 = w3563 & w9623;
assign w302 = (w217 & ~w6879) | (w217 & w2457) | (~w6879 & w2457);
assign w303 = ~w4921 & w398;
assign w304 = (~w8019 & w6374) | (~w8019 & w6498) | (w6374 & w6498);
assign w305 = ~w12427 & w5819;
assign w306 = w10568 & w5945;
assign w307 = (w14048 & ~w189) | (w14048 & w8075) | (~w189 & w8075);
assign w308 = (~w5622 & ~w4318) | (~w5622 & w13309) | (~w4318 & w13309);
assign w309 = ~b61 & ~a61;
assign w310 = ~w5490 & ~w12807;
assign w311 = ~w13282 & w13946;
assign w312 = (~w6716 & ~w956) | (~w6716 & w6394) | (~w956 & w6394);
assign w313 = ~w10435 & w6252;
assign w314 = (~w6637 & w2958) | (~w6637 & w2793) | (w2958 & w2793);
assign w315 = ~w10390 & w13039;
assign w316 = (w346 & w7318) | (w346 & ~w8282) | (w7318 & ~w8282);
assign w317 = (w6267 & w2953) | (w6267 & w5662) | (w2953 & w5662);
assign w318 = ~w9871 & ~w6986;
assign w319 = (w12406 & w1560) | (w12406 & w13112) | (w1560 & w13112);
assign w320 = ~w6927 & ~w2698;
assign w321 = ~w10041 & ~w7997;
assign w322 = w5741 & w9296;
assign w323 = (~w4989 & ~w12121) | (~w4989 & w3797) | (~w12121 & w3797);
assign w324 = (w1785 & w1932) | (w1785 & w9175) | (w1932 & w9175);
assign w325 = ~w3742 & ~w9788;
assign w326 = ~w13873 & w5664;
assign w327 = (~w1795 & w14664) | (~w1795 & w10798) | (w14664 & w10798);
assign w328 = w14306 & ~w8646;
assign w329 = ~w1563 & w13854;
assign w330 = ~w11302 & w4626;
assign w331 = (~w6426 & w5848) | (~w6426 & w9489) | (w5848 & w9489);
assign w332 = ~w2386 & ~w3927;
assign w333 = (~w13628 & w5867) | (~w13628 & w12796) | (w5867 & w12796);
assign w334 = w1957 & w8729;
assign w335 = (w2287 & w1920) | (w2287 & w14272) | (w1920 & w14272);
assign w336 = ~w12271 & ~w7445;
assign w337 = ~w14491 & w9183;
assign w338 = ~w2029 & w3589;
assign w339 = ~w9717 & w1305;
assign w340 = (w14074 & w14650) | (w14074 & w13311) | (w14650 & w13311);
assign w341 = w9817 & w5593;
assign w342 = ~w3903 & ~w12974;
assign w343 = ~w3751 & ~w9949;
assign w344 = (w14215 & w13596) | (w14215 & w1933) | (w13596 & w1933);
assign w345 = w13600 & ~w13134;
assign w346 = (w2445 & w12769) | (w2445 & w7518) | (w12769 & w7518);
assign w347 = w14486 & w9817;
assign w348 = w3201 & ~w11018;
assign w349 = w761 & ~w10854;
assign w350 = (w4561 & w10633) | (w4561 & w276) | (w10633 & w276);
assign w351 = ~w12798 & w2707;
assign w352 = ~w10618 & w8993;
assign w353 = (~w9798 & ~w2823) | (~w9798 & ~w6994) | (~w2823 & ~w6994);
assign w354 = (~w8282 & w6994) | (~w8282 & w2445) | (w6994 & w2445);
assign w355 = ~w6583 & w7713;
assign w356 = (~w1442 & w11429) | (~w1442 & w9089) | (w11429 & w9089);
assign w357 = (w4245 & w2027) | (w4245 & w13280) | (w2027 & w13280);
assign w358 = w7697 & w3978;
assign w359 = w12087 & w1965;
assign w360 = w2603 & w7317;
assign w361 = (w1507 & w12499) | (w1507 & w3061) | (w12499 & w3061);
assign w362 = (~w2698 & w1570) | (~w2698 & ~w3262) | (w1570 & ~w3262);
assign w363 = (~w1843 & w7689) | (~w1843 & w3811) | (w7689 & w3811);
assign w364 = ~b30 & ~a30;
assign w365 = (w11634 & w5259) | (w11634 & w14568) | (w5259 & w14568);
assign w366 = ~w4780 & w14659;
assign w367 = ~w142 & ~w1062;
assign w368 = (~w3721 & w9862) | (~w3721 & w5996) | (w9862 & w5996);
assign w369 = w3924 | w11732;
assign w370 = (w9510 & w5119) | (w9510 & w8692) | (w5119 & w8692);
assign w371 = (~w3904 & ~w10862) | (~w3904 & ~w14539) | (~w10862 & ~w14539);
assign w372 = w2751 & ~w3803;
assign w373 = (w4679 & w7265) | (w4679 & w12075) | (w7265 & w12075);
assign w374 = ~w7834 & ~w4193;
assign w375 = (~w6929 & w9970) | (~w6929 & w1615) | (w9970 & w1615);
assign w376 = (~w7962 & w2656) | (~w7962 & w9071) | (w2656 & w9071);
assign w377 = ~w183 & w7642;
assign w378 = (~w8130 & w7473) | (~w8130 & w8614) | (w7473 & w8614);
assign w379 = w7168 & ~w14268;
assign w380 = (~w5932 & w14051) | (~w5932 & ~w10117) | (w14051 & ~w10117);
assign w381 = (~w2655 & w10632) | (~w2655 & w10899) | (w10632 & w10899);
assign w382 = ~w4751 & w9938;
assign w383 = w11745 & w4458;
assign w384 = ~w12240 & w7684;
assign w385 = ~w6244 & w6179;
assign w386 = ~w11962 & w5150;
assign w387 = ~w12393 & ~w8033;
assign w388 = w11648 & ~w5340;
assign w389 = (w11925 & w650) | (w11925 & w10565) | (w650 & w10565);
assign w390 = (w6739 & ~w10263) | (w6739 & w14559) | (~w10263 & w14559);
assign w391 = w3039 & ~w12398;
assign w392 = ~w1799 & ~w7670;
assign w393 = ~w3012 & w7914;
assign w394 = ~w7369 & ~w3427;
assign w395 = (w5593 & w13947) | (w5593 & w7895) | (w13947 & w7895);
assign w396 = w7500 & ~w3657;
assign w397 = w3893 & ~w5344;
assign w398 = ~w12271 & w6014;
assign w399 = (~w14396 & w3458) | (~w14396 & w10160) | (w3458 & w10160);
assign w400 = w14594 & w12789;
assign w401 = w7794 & w2334;
assign w402 = (~w7737 & w1556) | (~w7737 & w749) | (w1556 & w749);
assign w403 = ~w13349 & w2687;
assign w404 = w6675 & w11474;
assign w405 = w13154 & w4873;
assign w406 = (~w7521 & w8565) | (~w7521 & w3859) | (w8565 & w3859);
assign w407 = ~w646 & w1799;
assign w408 = ~w11576 & w12357;
assign w409 = (w10317 & w13152) | (w10317 & w4455) | (w13152 & w4455);
assign w410 = ~w607 & ~w2701;
assign w411 = ~w4700 & ~w3427;
assign w412 = (~w4129 & w8226) | (~w4129 & w8222) | (w8226 & w8222);
assign w413 = w9423 & w2798;
assign w414 = (w13987 & w5449) | (w13987 & w14035) | (w5449 & w14035);
assign w415 = (~w5243 & w3146) | (~w5243 & w6935) | (w3146 & w6935);
assign w416 = w12662 & ~w8769;
assign w417 = w10676 & w3611;
assign w418 = w9349 & ~w9298;
assign w419 = ~w11547 & w8973;
assign w420 = (~w12889 & w1954) | (~w12889 & w3810) | (w1954 & w3810);
assign w421 = w11328 & w4361;
assign w422 = w7704 & ~w8512;
assign w423 = w7674 & w2072;
assign w424 = w13905 & ~w8667;
assign w425 = (w11318 & w3438) | (w11318 & w12376) | (w3438 & w12376);
assign w426 = ~w3288 & ~w11117;
assign w427 = ~w3765 & ~w7195;
assign w428 = (w5654 & w314) | (w5654 & ~w12376) | (w314 & ~w12376);
assign w429 = w8964 & w5284;
assign w430 = (w7114 & w13487) | (w7114 & ~w1467) | (w13487 & ~w1467);
assign w431 = ~w5827 & w12482;
assign w432 = w830 & w6166;
assign w433 = w809 & w2937;
assign w434 = (w9015 & w8226) | (w9015 & w12840) | (w8226 & w12840);
assign w435 = w13452 & ~w8629;
assign w436 = ~w8512 & w14528;
assign w437 = w13190 & ~w2748;
assign w438 = w5604 & ~w7768;
assign w439 = (~w8943 & w9872) | (~w8943 & w3300) | (w9872 & w3300);
assign w440 = ~w12271 & w13531;
assign w441 = ~w4512 & w12690;
assign w442 = w13443 & w10412;
assign w443 = ~w14465 & ~w5432;
assign w444 = ~w14558 & ~w14231;
assign w445 = (~w14659 & ~w10778) | (~w14659 & w9088) | (~w10778 & w9088);
assign w446 = ~w10654 & ~w8211;
assign w447 = (~w3602 & w8071) | (~w3602 & w5315) | (w8071 & w5315);
assign w448 = (~w6381 & w8234) | (~w6381 & w8987) | (w8234 & w8987);
assign w449 = w11405 & ~w11343;
assign w450 = (~w803 & w6113) | (~w803 & w13114) | (w6113 & w13114);
assign w451 = ~w12460 & ~w10114;
assign w452 = (w4855 & w14342) | (w4855 & ~w5620) | (w14342 & ~w5620);
assign w453 = ~w1668 & w3200;
assign w454 = (w9329 & ~w2) | (w9329 & ~w11756) | (~w2 & ~w11756);
assign w455 = ~w14227 & ~w3435;
assign w456 = w1607 & ~w13917;
assign w457 = (w1236 & ~w13027) | (w1236 & ~w1362) | (~w13027 & ~w1362);
assign w458 = w3914 & ~w14512;
assign w459 = w5515 & w9524;
assign w460 = w8665 & w12656;
assign w461 = (~w4515 & w2162) | (~w4515 & w8607) | (w2162 & w8607);
assign w462 = ~w5522 & ~w10182;
assign w463 = w608 & w7317;
assign w464 = ~w1257 & ~w11003;
assign w465 = ~w13864 & w11117;
assign w466 = w11835 & ~w2656;
assign w467 = ~w326 & w3487;
assign w468 = ~w10334 & ~w3693;
assign w469 = (w8399 & ~w4545) | (w8399 & ~w996) | (~w4545 & ~w996);
assign w470 = (~w14227 & w13222) | (~w14227 & w5569) | (w13222 & w5569);
assign w471 = w9788 & ~w6500;
assign w472 = (~w14141 & w9863) | (~w14141 & w714) | (w9863 & w714);
assign w473 = ~b82 & ~a82;
assign w474 = (~w1785 & w293) | (~w1785 & w9166) | (w293 & w9166);
assign w475 = b49 & a49;
assign w476 = w4109 & w5976;
assign w477 = (w10551 & w922) | (w10551 & w13831) | (w922 & w13831);
assign w478 = w192 & ~w9093;
assign w479 = w6538 & ~w9400;
assign w480 = ~w9608 & ~w1166;
assign w481 = ~w1805 & ~w1712;
assign w482 = w5177 & w5556;
assign w483 = w9827 & w10116;
assign w484 = ~w8840 & w10839;
assign w485 = ~w7488 & w6690;
assign w486 = w7498 & w12436;
assign w487 = w4213 & w8977;
assign w488 = ~w13321 & w8105;
assign w489 = ~w2941 & ~w690;
assign w490 = (~w10926 & w977) | (~w10926 & w8238) | (w977 & w8238);
assign w491 = ~w8001 & ~w8893;
assign w492 = ~w11547 & w4232;
assign w493 = ~w12121 & ~w13445;
assign w494 = (~w4697 & w4975) | (~w4697 & w3420) | (w4975 & w3420);
assign w495 = (w11978 & w4544) | (w11978 & ~w12937) | (w4544 & ~w12937);
assign w496 = ~w404 & w4994;
assign w497 = (w3400 & w12424) | (w3400 & w13500) | (w12424 & w13500);
assign w498 = ~w12452 & w11181;
assign w499 = ~w8035 & ~w2680;
assign w500 = ~w2675 & ~w475;
assign w501 = ~w11233 & w10372;
assign w502 = w9226 & ~w5664;
assign w503 = ~w14034 & w47;
assign w504 = ~w13324 & w14496;
assign w505 = ~w12481 & w9284;
assign w506 = ~w9296 & ~w10180;
assign w507 = (w7911 & w619) | (w7911 & w13818) | (w619 & w13818);
assign w508 = (~w13008 & w9506) | (~w13008 & w6750) | (w9506 & w6750);
assign w509 = w7400 & ~w7452;
assign w510 = ~w8234 & w608;
assign w511 = (w8030 & w14158) | (w8030 & w11398) | (w14158 & w11398);
assign w512 = (~w13587 & w2641) | (~w13587 & w14666) | (w2641 & w14666);
assign w513 = ~w8440 & w12241;
assign w514 = (~w11385 & w1996) | (~w11385 & w6901) | (w1996 & w6901);
assign w515 = w9518 & w2348;
assign w516 = ~w1563 & w11810;
assign w517 = (w1518 & w7092) | (w1518 & w2413) | (w7092 & w2413);
assign w518 = (~w10613 & w5025) | (~w10613 & w14381) | (w5025 & w14381);
assign w519 = w3914 & ~w5568;
assign w520 = w9518 & ~w2017;
assign w521 = ~w12808 & w1760;
assign w522 = w2320 & w6845;
assign w523 = (w3694 & w1254) | (w3694 & w1888) | (w1254 & w1888);
assign w524 = (~w7914 & ~w183) | (~w7914 & w12098) | (~w183 & w12098);
assign w525 = (~w9305 & w371) | (~w9305 & w9829) | (w371 & w9829);
assign w526 = (~w3325 & w1785) | (~w3325 & w4486) | (w1785 & w4486);
assign w527 = ~w706 & w3963;
assign w528 = (w13331 & w11593) | (w13331 & w2898) | (w11593 & w2898);
assign w529 = w4905 & ~w14317;
assign w530 = w7668 & w9748;
assign w531 = (w8234 & w11187) | (w8234 & w249) | (w11187 & w249);
assign w532 = (w11045 & ~w7137) | (w11045 & w6150) | (~w7137 & w6150);
assign w533 = (~w6583 & w2272) | (~w6583 & w9619) | (w2272 & w9619);
assign w534 = w10290 & ~w5556;
assign w535 = (~w3550 & w7397) | (~w3550 & w9973) | (w7397 & w9973);
assign w536 = (~w10477 & w9694) | (~w10477 & w8274) | (w9694 & w8274);
assign w537 = w10564 & ~w13058;
assign w538 = (w6502 & ~w1563) | (w6502 & w13416) | (~w1563 & w13416);
assign w539 = ~w5811 & w14259;
assign w540 = ~w11817 & ~w7365;
assign w541 = w14545 & w4615;
assign w542 = ~w1840 & w3524;
assign w543 = w14086 & ~w895;
assign w544 = w6436 & w2851;
assign w545 = w5213 & w5482;
assign w546 = ~w11117 & w5126;
assign w547 = w10872 & w10514;
assign w548 = ~w4780 & w5906;
assign w549 = w14302 & w8827;
assign w550 = (w1805 & w4050) | (w1805 & w10492) | (w4050 & w10492);
assign w551 = ~w7212 & w11689;
assign w552 = (~w9541 & w6288) | (~w9541 & w4282) | (w6288 & w4282);
assign w553 = (w12138 & w10384) | (w12138 & ~w8444) | (w10384 & ~w8444);
assign w554 = w7157 & ~w11213;
assign w555 = w497 & w12015;
assign w556 = ~w12475 & w4601;
assign w557 = (~w13654 & w10785) | (~w13654 & w14397) | (w10785 & w14397);
assign w558 = (~w11597 & w6615) | (~w11597 & w5180) | (w6615 & w5180);
assign w559 = w10020 & w12698;
assign w560 = ~w13854 & ~w12170;
assign w561 = w4213 & ~w10423;
assign w562 = w10036 & w9032;
assign w563 = ~w8328 & ~w6763;
assign w564 = (~w8827 & ~w953) | (~w8827 & w7959) | (~w953 & w7959);
assign w565 = ~w6321 & w878;
assign w566 = ~w4241 & w8250;
assign w567 = (w3853 & w14604) | (w3853 & ~w12293) | (w14604 & ~w12293);
assign w568 = w3289 & w14074;
assign w569 = ~w3483 & ~w13095;
assign w570 = (w9881 & w1438) | (w9881 & ~w2670) | (w1438 & ~w2670);
assign w571 = w10082 & w3963;
assign w572 = w5715 & w5900;
assign w573 = ~w2701 & ~w9256;
assign w574 = (w13743 & w4779) | (w13743 & w1480) | (w4779 & w1480);
assign w575 = (~w4479 & w12071) | (~w4479 & w9239) | (w12071 & w9239);
assign w576 = w13924 & ~w11395;
assign w577 = ~w12819 & w6763;
assign w578 = ~w13094 & w7829;
assign w579 = (~w10116 & w10301) | (~w10116 & w12553) | (w10301 & w12553);
assign w580 = ~w13349 & w8596;
assign w581 = w13929 & w3172;
assign w582 = ~w12528 & w2159;
assign w583 = w2701 & ~w2448;
assign w584 = w5103 & ~w447;
assign w585 = w7968 & w6908;
assign w586 = w226 & w9074;
assign w587 = ~w8234 & ~w3526;
assign w588 = w11420 & w5233;
assign w589 = (w6209 & w9262) | (w6209 & w2835) | (w9262 & w2835);
assign w590 = (~w13375 & ~w5498) | (~w13375 & ~w8282) | (~w5498 & ~w8282);
assign w591 = ~w9608 & w11223;
assign w592 = w9243 & ~w2386;
assign w593 = w12713 & ~w10962;
assign w594 = ~w4889 & w4546;
assign w595 = (w6724 & w6181) | (w6724 & w6790) | (w6181 & w6790);
assign w596 = w11068 & ~w14340;
assign w597 = ~w4050 & w812;
assign w598 = ~w5178 & ~w4291;
assign w599 = (w1274 & ~w183) | (w1274 & w10750) | (~w183 & w10750);
assign w600 = (~w3727 & ~w4858) | (~w3727 & w9498) | (~w4858 & w9498);
assign w601 = ~w6006 & w10615;
assign w602 = w2128 & w6522;
assign w603 = ~w11882 & ~w8197;
assign w604 = ~w5300 & w14605;
assign w605 = (w4976 & w12917) | (w4976 & w3999) | (w12917 & w3999);
assign w606 = w11309 & ~w13977;
assign w607 = b94 & a94;
assign w608 = ~w4312 & ~w12112;
assign w609 = ~w1563 & ~w6187;
assign w610 = (w10560 & ~w2555) | (w10560 & w7292) | (~w2555 & w7292);
assign w611 = (~w3550 & w3824) | (~w3550 & w7382) | (w3824 & w7382);
assign w612 = (w6979 & w9136) | (w6979 & w8243) | (w9136 & w8243);
assign w613 = ~w2928 & w10773;
assign w614 = w14062 & ~w13835;
assign w615 = (~w3550 & w11876) | (~w3550 & w1611) | (w11876 & w1611);
assign w616 = ~w9846 & ~w12732;
assign w617 = w2656 & w10997;
assign w618 = w6167 & ~w8287;
assign w619 = w10123 & w10385;
assign w620 = w3958 & ~w3734;
assign w621 = ~w309 & ~w8827;
assign w622 = w12460 & w1821;
assign w623 = ~w12460 & ~w11360;
assign w624 = w8171 & ~w11216;
assign w625 = w3904 & w9499;
assign w626 = w10676 & w2680;
assign w627 = (w3219 & w2317) | (w3219 & w981) | (w2317 & w981);
assign w628 = (~w13178 & w1510) | (~w13178 & w10741) | (w1510 & w10741);
assign w629 = w9252 & w1293;
assign w630 = w12170 & ~w1692;
assign w631 = (w3036 & w13324) | (w3036 & w1410) | (w13324 & w1410);
assign w632 = ~w11008 & ~w13717;
assign w633 = ~w1182 & ~w275;
assign w634 = w9252 & ~w1206;
assign w635 = (w10946 & w1846) | (w10946 & w2088) | (w1846 & w2088);
assign w636 = ~w142 & ~w10334;
assign w637 = w14640 & ~w5761;
assign w638 = ~w5562 & w5288;
assign w639 = (w990 & w9485) | (w990 & w14164) | (w9485 & w14164);
assign w640 = w10941 & w10182;
assign w641 = (~w9227 & w2175) | (~w9227 & w10608) | (w2175 & w10608);
assign w642 = (~w999 & w3953) | (~w999 & w3134) | (w3953 & w3134);
assign w643 = (w2936 & w5060) | (w2936 & ~w3957) | (w5060 & ~w3957);
assign w644 = w3550 & w902;
assign w645 = (~w224 & w2578) | (~w224 & w13453) | (w2578 & w13453);
assign w646 = ~w6538 & ~w10949;
assign w647 = w1821 & ~w12614;
assign w648 = (w14074 & w7522) | (w14074 & w2240) | (w7522 & w2240);
assign w649 = ~w9264 & ~w3546;
assign w650 = ~w10689 & w2381;
assign w651 = (w9305 & w986) | (w9305 & w9739) | (w986 & w9739);
assign w652 = ~w7722 & ~w7962;
assign w653 = ~w11246 & w1059;
assign w654 = ~w218 & w6301;
assign w655 = ~w1986 & ~w14266;
assign w656 = ~w13878 & ~w9642;
assign w657 = w7022 & ~w3427;
assign w658 = w1821 & ~w8992;
assign w659 = w3823 & w10366;
assign w660 = ~w6580 & ~w9846;
assign w661 = ~w5018 & w695;
assign w662 = ~w1782 & w7857;
assign w663 = w10517 & ~w12604;
assign w664 = ~w4311 & ~w802;
assign w665 = (~w2044 & ~w13019) | (~w2044 & w13474) | (~w13019 & w13474);
assign w666 = (~w7754 & w10350) | (~w7754 & w21) | (w10350 & w21);
assign w667 = w7941 & ~w8929;
assign w668 = (~w13344 & w12798) | (~w13344 & w3991) | (w12798 & w3991);
assign w669 = ~w9086 & ~w1305;
assign w670 = w5604 & w8919;
assign w671 = ~w1047 & w1953;
assign w672 = (~w4627 & w7545) | (~w4627 & ~w9872) | (w7545 & ~w9872);
assign w673 = ~w13697 & w6584;
assign w674 = (w2409 & ~w13262) | (w2409 & w9446) | (~w13262 & w9446);
assign w675 = ~w14387 & ~w12052;
assign w676 = ~w13462 & w6158;
assign w677 = (w6486 & w9450) | (w6486 & w10963) | (w9450 & w10963);
assign w678 = (~w4030 & w5758) | (~w4030 & w2418) | (w5758 & w2418);
assign w679 = (w3215 & w14664) | (w3215 & w947) | (w14664 & w947);
assign w680 = w9541 & ~w3056;
assign w681 = w9776 & ~w716;
assign w682 = w14019 & w4049;
assign w683 = (~w9608 & w1331) | (~w9608 & w6133) | (w1331 & w6133);
assign w684 = ~w5852 & w7668;
assign w685 = (w5184 & w10242) | (w5184 & w13910) | (w10242 & w13910);
assign w686 = ~w318 & ~w7212;
assign w687 = (~w13596 & w4099) | (~w13596 & w3084) | (w4099 & w3084);
assign w688 = (w14594 & w3371) | (w14594 & w10154) | (w3371 & w10154);
assign w689 = ~w1139 & w10930;
assign w690 = ~w12148 & ~w8768;
assign w691 = w7001 & w4458;
assign w692 = w5996 | w9862;
assign w693 = ~w5294 & ~w6795;
assign w694 = ~w9298 & w3730;
assign w695 = ~w165 & ~w14471;
assign w696 = (w4354 & w12878) | (w4354 & w14506) | (w12878 & w14506);
assign w697 = (w3039 & ~w7630) | (w3039 & w7324) | (~w7630 & w7324);
assign w698 = (w11708 & w8900) | (w11708 & w2170) | (w8900 & w2170);
assign w699 = (~w4512 & w8965) | (~w4512 & w13415) | (w8965 & w13415);
assign w700 = w2712 & w1892;
assign w701 = w3224 & w10511;
assign w702 = (~w12537 & w1927) | (~w12537 & w12794) | (w1927 & w12794);
assign w703 = w9480 & ~w3904;
assign w704 = (w4771 & w13432) | (w4771 & ~w12376) | (w13432 & ~w12376);
assign w705 = (w5950 & w10791) | (w5950 & w11696) | (w10791 & w11696);
assign w706 = b105 & a105;
assign w707 = (~w1086 & w11548) | (~w1086 & w6200) | (w11548 & w6200);
assign w708 = ~w13423 & ~w9296;
assign w709 = w13924 & ~w5406;
assign w710 = w9268 & ~w1883;
assign w711 = ~w3578 & ~w5444;
assign w712 = (~w9296 & w9146) | (~w9296 & w8617) | (w9146 & w8617);
assign w713 = (w52 & w5947) | (w52 & w1028) | (w5947 & w1028);
assign w714 = (~w10119 & ~w12240) | (~w10119 & w9863) | (~w12240 & w9863);
assign w715 = w3012 & w10254;
assign w716 = ~w11940 & ~w2646;
assign w717 = (w2150 & w13825) | (w2150 & ~w4783) | (w13825 & ~w4783);
assign w718 = ~w3325 & ~w8742;
assign w719 = w5412 & ~w7732;
assign w720 = w11682 & w6896;
assign w721 = ~w3038 & ~w6572;
assign w722 = w3161 & ~w13258;
assign w723 = w11871 & ~w5994;
assign w724 = w8018 & w7317;
assign w725 = (w1190 & w2901) | (w1190 & w3296) | (w2901 & w3296);
assign w726 = (w1634 & w2525) | (w1634 & ~w12376) | (w2525 & ~w12376);
assign w727 = (w2924 & ~w4999) | (w2924 & w8446) | (~w4999 & w8446);
assign w728 = w13620 & ~w10689;
assign w729 = (~w10023 & w3721) | (~w10023 & w11759) | (w3721 & w11759);
assign w730 = w13275 & ~w4198;
assign w731 = (w6879 & w11712) | (w6879 & w6802) | (w11712 & w6802);
assign w732 = (w967 & w300) | (w967 & w3274) | (w300 & w3274);
assign w733 = (~w2655 & w5903) | (~w2655 & w9140) | (w5903 & w9140);
assign w734 = (w7914 & ~w14396) | (w7914 & w6174) | (~w14396 & w6174);
assign w735 = w13704 & w3173;
assign w736 = w2611 & w14113;
assign w737 = w5288 & w8459;
assign w738 = (~w2951 & w6345) | (~w2951 & w5827) | (w6345 & w5827);
assign w739 = ~w11785 & w10246;
assign w740 = (~w556 & w7692) | (~w556 & w11774) | (w7692 & w11774);
assign w741 = w1402 & w12439;
assign w742 = w14395 & w10290;
assign w743 = w10708 & ~w13400;
assign w744 = w7142 & w9104;
assign w745 = w2680 & ~w8769;
assign w746 = (~w7906 & w3767) | (~w7906 & w1951) | (w3767 & w1951);
assign w747 = (w749 & w10767) | (w749 & w11073) | (w10767 & w11073);
assign w748 = w10704 & ~w6845;
assign w749 = w13126 & w10486;
assign w750 = ~w10703 & ~w5217;
assign w751 = ~w3157 & w3904;
assign w752 = w12655 & w1676;
assign w753 = w5794 | w7220;
assign w754 = (~w1789 & w2145) | (~w1789 & w2249) | (w2145 & w2249);
assign w755 = (w7267 & ~w11459) | (w7267 & w13087) | (~w11459 & w13087);
assign w756 = (~w302 & w8678) | (~w302 & w11837) | (w8678 & w11837);
assign w757 = (~w5785 & ~w4336) | (~w5785 & w7405) | (~w4336 & w7405);
assign w758 = w724 & w11613;
assign w759 = w8546 & w8682;
assign w760 = w5132 & ~w4257;
assign w761 = w13452 & ~w8305;
assign w762 = ~w6176 & w9120;
assign w763 = ~w1873 & w12893;
assign w764 = (w2211 & w12969) | (w2211 & w4917) | (w12969 & w4917);
assign w765 = w12577 & ~w13854;
assign w766 = (~w5406 & w8191) | (~w5406 & ~w4334) | (w8191 & ~w4334);
assign w767 = w7652 & ~w3704;
assign w768 = ~w11138 & w13118;
assign w769 = (~w10023 & w5655) | (~w10023 & w6618) | (w5655 & w6618);
assign w770 = w12958 & w8389;
assign w771 = ~w3774 & ~w10042;
assign w772 = ~w13451 & ~w4202;
assign w773 = w9458 & w9341;
assign w774 = w2656 & ~w3823;
assign w775 = ~w6597 & w8606;
assign w776 = (~w1712 & w10304) | (~w1712 & w11864) | (w10304 & w11864);
assign w777 = w2493 & w6384;
assign w778 = w6665 & w217;
assign w779 = (~w4127 & w12003) | (~w4127 & w7996) | (w12003 & w7996);
assign w780 = ~w14043 & ~w3112;
assign w781 = ~w9608 & w11943;
assign w782 = (w8007 & w2124) | (w8007 & w7073) | (w2124 & w7073);
assign w783 = (w9921 & w153) | (w9921 & w12484) | (w153 & w12484);
assign w784 = (~w9151 & w7182) | (~w9151 & w13015) | (w7182 & w13015);
assign w785 = ~w2317 & w2430;
assign w786 = w8553 & w10352;
assign w787 = w3759 & ~w4341;
assign w788 = (~w13685 & w14357) | (~w13685 & w428) | (w14357 & w428);
assign w789 = (w10966 & w3726) | (w10966 & w5642) | (w3726 & w5642);
assign w790 = w10338 & w9711;
assign w791 = w6436 & w1087;
assign w792 = w9518 & ~w11950;
assign w793 = (w2599 & ~w9059) | (w2599 & w10313) | (~w9059 & w10313);
assign w794 = w10013 & ~w706;
assign w795 = ~w1472 & ~w7058;
assign w796 = w1518 & ~w5497;
assign w797 = (~w5823 & ~w8572) | (~w5823 & w1407) | (~w8572 & w1407);
assign w798 = ~w7373 & w12775;
assign w799 = w3124 & ~w3904;
assign w800 = ~w1563 & w563;
assign w801 = w8830 & w227;
assign w802 = (w13531 & w12980) | (w13531 & w12346) | (w12980 & w12346);
assign w803 = b56 & a56;
assign w804 = ~w15 & ~w10959;
assign w805 = ~w1552 & w11721;
assign w806 = ~w13451 & ~w50;
assign w807 = ~w3717 & w10880;
assign w808 = (~w142 & ~w6500) | (~w142 & w6872) | (~w6500 & w6872);
assign w809 = w10290 & w10700;
assign w810 = w5103 & ~w4978;
assign w811 = ~w7764 & w10763;
assign w812 = ~w13222 & w14072;
assign w813 = ~w11216 & ~w2387;
assign w814 = (~w2922 & ~w4103) | (~w2922 & w5429) | (~w4103 & w5429);
assign w815 = w3550 & w5658;
assign w816 = (w3904 & ~w3224) | (w3904 & w13200) | (~w3224 & w13200);
assign w817 = w5265 & ~w10450;
assign w818 = w7296 & w5532;
assign w819 = (w6219 & w4520) | (w6219 & w13772) | (w4520 & w13772);
assign w820 = ~w3590 & ~w13861;
assign w821 = ~w9672 & w8080;
assign w822 = (~w8226 & w12925) | (~w8226 & w13678) | (w12925 & w13678);
assign w823 = (~w6825 & w3480) | (~w6825 & w6264) | (w3480 & w6264);
assign w824 = ~w4700 & w11861;
assign w825 = w14400 & w8687;
assign w826 = w13357 & ~w5630;
assign w827 = ~w6461 & ~w10212;
assign w828 = (w13531 & w5702) | (w13531 & w5980) | (w5702 & w5980);
assign w829 = ~b54 & ~a54;
assign w830 = w2618 & w1780;
assign w831 = w10713 & w9400;
assign w832 = (w12988 & w13700) | (w12988 & w8337) | (w13700 & w8337);
assign w833 = (~w4587 & ~w9748) | (~w4587 & w3474) | (~w9748 & w3474);
assign w834 = (w5756 & w12928) | (w5756 & w9152) | (w12928 & w9152);
assign w835 = w25 & w2491;
assign w836 = ~w7630 & ~w5333;
assign w837 = (w10248 & w2910) | (w10248 & w5146) | (w2910 & w5146);
assign w838 = w4153 & w10597;
assign w839 = ~w5599 & ~w28;
assign w840 = ~w8475 & ~w2433;
assign w841 = w14412 & w7841;
assign w842 = w3137 & ~w13323;
assign w843 = ~w7857 & w4961;
assign w844 = ~w11040 & w1852;
assign w845 = w7213 & ~w4191;
assign w846 = (w2670 & w9730) | (w2670 & w747) | (w9730 & w747);
assign w847 = w3562 & ~w14385;
assign w848 = w1756 & w5348;
assign w849 = (~w695 & ~w8484) | (~w695 & w5622) | (~w8484 & w5622);
assign w850 = (w10367 & w6660) | (w10367 & w6295) | (w6660 & w6295);
assign w851 = ~w982 & w12311;
assign w852 = ~b67 & ~a67;
assign w853 = (w13685 & w8685) | (w13685 & w7972) | (w8685 & w7972);
assign w854 = ~w6336 & w9673;
assign w855 = (w10966 & w11913) | (w10966 & w789) | (w11913 & w789);
assign w856 = (~w10719 & w2673) | (~w10719 & w7158) | (w2673 & w7158);
assign w857 = w11759 & w1317;
assign w858 = ~w13652 & w9242;
assign w859 = ~w11642 & ~w14445;
assign w860 = ~w12225 & w6123;
assign w861 = w1802 & w646;
assign w862 = (~w7429 & w3155) | (~w7429 & w10420) | (w3155 & w10420);
assign w863 = ~w6538 & ~w6580;
assign w864 = (w13288 & w2562) | (w13288 & ~w2670) | (w2562 & ~w2670);
assign w865 = (w5767 & w1986) | (w5767 & w4383) | (w1986 & w4383);
assign w866 = (w6425 & ~w474) | (w6425 & w6036) | (~w474 & w6036);
assign w867 = ~w4431 & ~w4111;
assign w868 = (~w6041 & w4099) | (~w6041 & w1034) | (w4099 & w1034);
assign w869 = (w7240 & w5869) | (w7240 & w5861) | (w5869 & w5861);
assign w870 = ~w5532 & ~w2492;
assign w871 = (w453 & ~w9320) | (w453 & w8349) | (~w9320 & w8349);
assign w872 = ~w71 & w482;
assign w873 = ~w6442 & ~w4483;
assign w874 = ~w13297 & w6689;
assign w875 = (w2181 & w6380) | (w2181 & w2148) | (w6380 & w2148);
assign w876 = ~w12548 & ~w11989;
assign w877 = (w4796 & w11681) | (w4796 & w9926) | (w11681 & w9926);
assign w878 = ~w11447 & ~w9408;
assign w879 = (~w9480 & w6689) | (~w9480 & w8619) | (w6689 & w8619);
assign w880 = (w10045 & ~w9541) | (w10045 & w7946) | (~w9541 & w7946);
assign w881 = (~w2941 & ~w1087) | (~w2941 & w203) | (~w1087 & w203);
assign w882 = w7886 & ~w11666;
assign w883 = (~w7962 & w13122) | (~w7962 & w376) | (w13122 & w376);
assign w884 = ~b80 & ~a80;
assign w885 = ~w7226 & ~w14340;
assign w886 = w7317 & w2171;
assign w887 = (~w11810 & w9608) | (~w11810 & w6012) | (w9608 & w6012);
assign w888 = w10784 & ~w14028;
assign w889 = ~w9890 & w13040;
assign w890 = ~w10408 & w12642;
assign w891 = w13767 & w2084;
assign w892 = ~w11228 & w4129;
assign w893 = w1986 & w13628;
assign w894 = b59 & a59;
assign w895 = w10422 & w2157;
assign w896 = ~b126 & ~a126;
assign w897 = (~w5070 & w2559) | (~w5070 & w10650) | (w2559 & w10650);
assign w898 = w13412 & w6898;
assign w899 = (w2150 & w13825) | (w2150 & ~w9215) | (w13825 & ~w9215);
assign w900 = w8873 & ~w11732;
assign w901 = ~w5830 & ~w3316;
assign w902 = ~w4780 & ~w11068;
assign w903 = w8154 & ~w1298;
assign w904 = (w8769 & w6412) | (w8769 & w10840) | (w6412 & w10840);
assign w905 = w7190 & ~w9087;
assign w906 = (w1457 & w236) | (w1457 & w14074) | (w236 & w14074);
assign w907 = ~w13839 & w6785;
assign w908 = ~w166 & w5005;
assign w909 = (~w4938 & w5086) | (~w4938 & w8541) | (w5086 & w8541);
assign w910 = w7349 & w8537;
assign w911 = w6391 & w3527;
assign w912 = w13344 & ~w8475;
assign w913 = w14417 & ~w309;
assign w914 = w12330 & ~w3122;
assign w915 = w5778 & w1062;
assign w916 = ~w2264 & w6257;
assign w917 = (~w3823 & w4099) | (~w3823 & w774) | (w4099 & w774);
assign w918 = (~w1469 & w13904) | (~w1469 & ~w6563) | (w13904 & ~w6563);
assign w919 = (~w439 & w14435) | (~w439 & w9958) | (w14435 & w9958);
assign w920 = (w4099 & w4581) | (w4099 & w7446) | (w4581 & w7446);
assign w921 = w14396 & w9225;
assign w922 = ~w6601 & ~w9526;
assign w923 = (~w7080 & w2470) | (~w7080 & w5673) | (w2470 & w5673);
assign w924 = w7681 & ~w3963;
assign w925 = ~w4158 & w11884;
assign w926 = w5998 & ~w6170;
assign w927 = (w1704 & w13859) | (w1704 & ~w2595) | (w13859 & ~w2595);
assign w928 = ~w468 & w4337;
assign w929 = (w12656 & w13507) | (w12656 & ~w12553) | (w13507 & ~w12553);
assign w930 = ~w4688 & w14038;
assign w931 = w1813 & w12510;
assign w932 = (w14087 & w8868) | (w14087 & w5417) | (w8868 & w5417);
assign w933 = ~w14253 & w616;
assign w934 = w3516 & w14523;
assign w935 = ~w12003 & w11532;
assign w936 = ~w71 & w6136;
assign w937 = (~w10820 & ~w3316) | (~w10820 & w13108) | (~w3316 & w13108);
assign w938 = w3944 & w13857;
assign w939 = (w5901 & w11852) | (w5901 & w12513) | (w11852 & w12513);
assign w940 = w10523 & w13839;
assign w941 = ~w3098 & ~w3885;
assign w942 = ~w813 & w13013;
assign w943 = ~w2660 & w6040;
assign w944 = (~w2159 & w9608) | (~w2159 & w14669) | (w9608 & w14669);
assign w945 = (~w12480 & ~w6691) | (~w12480 & ~w11165) | (~w6691 & ~w11165);
assign w946 = (w2476 & w3884) | (w2476 & w10428) | (w3884 & w10428);
assign w947 = (w3550 & w6447) | (w3550 & w5886) | (w6447 & w5886);
assign w948 = w4905 & ~w8858;
assign w949 = ~w8423 & ~w9705;
assign w950 = ~w2464 & ~w2941;
assign w951 = ~w7834 & w4253;
assign w952 = (~w11261 & w8999) | (~w11261 & w6590) | (w8999 & w6590);
assign w953 = ~w12371 & ~w3175;
assign w954 = w2656 & w3602;
assign w955 = ~w3506 & ~w3976;
assign w956 = w3175 & ~w13465;
assign w957 = w5272 & w12097;
assign w958 = w13323 & w8253;
assign w959 = w12088 & w2363;
assign w960 = ~w2736 & ~w3045;
assign w961 = w8681 & ~w13085;
assign w962 = (w7082 & w10569) | (w7082 & w13829) | (w10569 & w13829);
assign w963 = w1166 & w8827;
assign w964 = ~w10298 & ~w190;
assign w965 = ~w7418 & w12764;
assign w966 = ~w10468 & ~w972;
assign w967 = w13872 & ~w3320;
assign w968 = w9499 & ~w6297;
assign w969 = ~w2144 & w8734;
assign w970 = ~w5140 & w6888;
assign w971 = (~w2663 & ~w12893) | (~w2663 & w13281) | (~w12893 & w13281);
assign w972 = (w10463 & w9487) | (w10463 & w5617) | (w9487 & w5617);
assign w973 = ~w14224 & ~w6929;
assign w974 = ~w5559 & w8078;
assign w975 = ~w5363 & w10795;
assign w976 = (w6935 & w11191) | (w6935 & w9749) | (w11191 & w9749);
assign w977 = (~w12528 & ~w6699) | (~w12528 & w582) | (~w6699 & w582);
assign w978 = ~w12543 & w10481;
assign w979 = ~w7001 & ~w13323;
assign w980 = w607 & ~w10182;
assign w981 = w1563 & w3219;
assign w982 = (~w1821 & w5395) | (~w1821 & w14006) | (w5395 & w14006);
assign w983 = w840 & w11760;
assign w984 = ~w142 & ~w13839;
assign w985 = ~w9533 & ~w11550;
assign w986 = ~w9708 & w6849;
assign w987 = ~w12543 & w2083;
assign w988 = ~w3379 & ~w5766;
assign w989 = ~w13810 & w12763;
assign w990 = w4855 & ~w14398;
assign w991 = ~w2887 & w7911;
assign w992 = (~w6716 & ~w227) | (~w6716 & w6713) | (~w227 & w6713);
assign w993 = ~w8475 & w11287;
assign w994 = ~w12929 & w3221;
assign w995 = (w4511 & w13397) | (w4511 & w2825) | (w13397 & w2825);
assign w996 = (~w7639 & w5229) | (~w7639 & w1228) | (w5229 & w1228);
assign w997 = (w4354 & w12878) | (w4354 & w12588) | (w12878 & w12588);
assign w998 = (w8584 & w10467) | (w8584 & ~w3226) | (w10467 & ~w3226);
assign w999 = w3215 & w4541;
assign w1000 = w7113 & w3098;
assign w1001 = w7587 & w14026;
assign w1002 = w12483 & ~w5068;
assign w1003 = ~w2218 & w6967;
assign w1004 = w11041 & w10140;
assign w1005 = w2065 & ~w9211;
assign w1006 = w14087 & ~w5328;
assign w1007 = w4287 & w608;
assign w1008 = (w7082 & w14288) | (w7082 & w851) | (w14288 & w851);
assign w1009 = w12112 & w10872;
assign w1010 = w2159 & ~w6889;
assign w1011 = (~w11031 & w9389) | (~w11031 & w5827) | (w9389 & w5827);
assign w1012 = ~w183 & ~w2567;
assign w1013 = (~w9747 & w2617) | (~w9747 & w6619) | (w2617 & w6619);
assign w1014 = (~w4607 & w10776) | (~w4607 & w2447) | (w10776 & w2447);
assign w1015 = ~w7490 & ~w1221;
assign w1016 = ~w12065 & ~w8827;
assign w1017 = ~w5294 & ~w11878;
assign w1018 = (~w8451 & w1191) | (~w8451 & w3579) | (w1191 & w3579);
assign w1019 = w3526 & ~w9805;
assign w1020 = ~w2210 & w6321;
assign w1021 = ~w2500 & ~w7821;
assign w1022 = ~w3170 & ~w7705;
assign w1023 = ~w3823 & ~w7423;
assign w1024 = w14295 & ~w13065;
assign w1025 = (w6802 & w3896) | (w6802 & w702) | (w3896 & w702);
assign w1026 = (~w2655 & w6565) | (~w2655 & w7153) | (w6565 & w7153);
assign w1027 = ~w852 & ~w13733;
assign w1028 = ~w6783 & w9486;
assign w1029 = ~w9283 & w7483;
assign w1030 = ~w5294 & w9713;
assign w1031 = ~w12569 & w6795;
assign w1032 = w1498 & w7526;
assign w1033 = (~w8614 & w6754) | (~w8614 & w7039) | (w6754 & w7039);
assign w1034 = w2656 & ~w6041;
assign w1035 = (~w13685 & w14362) | (~w13685 & w2043) | (w14362 & w2043);
assign w1036 = ~w3036 & ~w12819;
assign w1037 = w8666 & w8860;
assign w1038 = w10431 & w13793;
assign w1039 = ~w13902 & ~w7461;
assign w1040 = ~w9960 & ~w10641;
assign w1041 = w10491 & w2300;
assign w1042 = ~w7668 & w1805;
assign w1043 = (w11708 & w1353) | (w11708 & ~w14375) | (w1353 & ~w14375);
assign w1044 = ~w491 & w14601;
assign w1045 = w3904 & ~w13410;
assign w1046 = (~w463 & ~w11147) | (~w463 & w6956) | (~w11147 & w6956);
assign w1047 = (~w3034 & w4381) | (~w3034 & w2235) | (w4381 & w2235);
assign w1048 = (w894 & w2463) | (w894 & w5375) | (w2463 & w5375);
assign w1049 = ~w9432 & w11668;
assign w1050 = w5481 & w14631;
assign w1051 = ~w3914 & w12620;
assign w1052 = ~w5693 & ~w10145;
assign w1053 = ~w5525 & w2312;
assign w1054 = ~w7085 & w588;
assign w1055 = w14116 & ~w5270;
assign w1056 = ~w4158 & w11203;
assign w1057 = w7857 & w957;
assign w1058 = ~w5005 & ~w13820;
assign w1059 = ~w2353 & ~w5843;
assign w1060 = w5697 & w6310;
assign w1061 = w11661 & w466;
assign w1062 = ~w12604 & ~w9480;
assign w1063 = (~w591 & ~w13219) | (~w591 & w887) | (~w13219 & w887);
assign w1064 = ~w2425 & ~w7085;
assign w1065 = w3963 & w13726;
assign w1066 = w14302 & w11902;
assign w1067 = w5522 & w8396;
assign w1068 = ~w4992 & w11798;
assign w1069 = ~w13256 & w13980;
assign w1070 = ~w13740 & ~w12492;
assign w1071 = w12271 & w12868;
assign w1072 = (w13771 & w7797) | (w13771 & w7849) | (w7797 & w7849);
assign w1073 = (w1267 & w14245) | (w1267 & w12226) | (w14245 & w12226);
assign w1074 = (w2275 & w1135) | (w2275 & w2801) | (w1135 & w2801);
assign w1075 = w505 & w6689;
assign w1076 = ~w3786 & w7213;
assign w1077 = w8464 | w7762;
assign w1078 = ~w10450 & ~w4464;
assign w1079 = ~w4473 & ~w8285;
assign w1080 = w7645 & ~w10682;
assign w1081 = (w3334 & w14355) | (w3334 & w318) | (w14355 & w318);
assign w1082 = w6035 & w3530;
assign w1083 = ~w922 & w569;
assign w1084 = (~w13281 & w763) | (~w13281 & w9261) | (w763 & w9261);
assign w1085 = (w5399 & w3616) | (w5399 & w10979) | (w3616 & w10979);
assign w1086 = ~w6577 & ~w1303;
assign w1087 = (~w12604 & w13730) | (~w12604 & w663) | (w13730 & w663);
assign w1088 = w4525 & ~w8839;
assign w1089 = (~w3550 & w8982) | (~w3550 & w10374) | (w8982 & w10374);
assign w1090 = w7587 & ~w5057;
assign w1091 = w10326 & ~w11168;
assign w1092 = ~w5732 & w12135;
assign w1093 = ~w11745 & ~w2729;
assign w1094 = w21 & w256;
assign w1095 = w8929 & ~w125;
assign w1096 = b87 & a87;
assign w1097 = w6739 & ~w6790;
assign w1098 = ~w1348 & w786;
assign w1099 = (w5742 & w12499) | (w5742 & w3312) | (w12499 & w3312);
assign w1100 = (~w1712 & w3879) | (~w1712 & w4874) | (w3879 & w4874);
assign w1101 = b11 & a11;
assign w1102 = (w3631 & w5477) | (w3631 & w7124) | (w5477 & w7124);
assign w1103 = w8754 & ~w1096;
assign w1104 = ~w12553 & w12662;
assign w1105 = w12088 & ~w6301;
assign w1106 = w13796 & w13634;
assign w1107 = ~a93 & w12460;
assign w1108 = w11364 & ~w6064;
assign w1109 = ~w8234 & w13115;
assign w1110 = w6282 & w12593;
assign w1111 = ~w9801 & w791;
assign w1112 = (w3994 & w9047) | (w3994 & w14644) | (w9047 & w14644);
assign w1113 = (w5316 & w6426) | (w5316 & w9382) | (w6426 & w9382);
assign w1114 = w3734 & w10514;
assign w1115 = ~w12167 & ~w1993;
assign w1116 = ~w1748 & w8469;
assign w1117 = w433 & ~w13815;
assign w1118 = ~w12057 & ~w6081;
assign w1119 = ~w7244 & ~w6689;
assign w1120 = w5103 & ~w6860;
assign w1121 = w7100 & ~w6889;
assign w1122 = w1729 & w2909;
assign w1123 = ~w10343 & w6318;
assign w1124 = w13733 & ~w3717;
assign w1125 = w607 & w10699;
assign w1126 = (w13169 & w13844) | (w13169 & w3215) | (w13844 & w3215);
assign w1127 = w3550 & w6108;
assign w1128 = w14396 & w382;
assign w1129 = w5778 & ~w4178;
assign w1130 = w3007 & ~w9246;
assign w1131 = w13599 & ~w6342;
assign w1132 = ~w6358 & ~w12949;
assign w1133 = w3755 & ~w10305;
assign w1134 = w10225 & w8900;
assign w1135 = (~w6886 & w4512) | (~w6886 & w2917) | (w4512 & w2917);
assign w1136 = ~w14302 & w5732;
assign w1137 = (~w11699 & w12592) | (~w11699 & w5839) | (w12592 & w5839);
assign w1138 = ~w11225 & w13833;
assign w1139 = w13189 & ~w8396;
assign w1140 = w3175 & w7794;
assign w1141 = w7794 & w7218;
assign w1142 = ~w1625 & ~w7783;
assign w1143 = ~w1082 & w14476;
assign w1144 = (~w5993 & w5188) | (~w5993 & w9649) | (w5188 & w9649);
assign w1145 = w7794 & w1695;
assign w1146 = w1570 | ~w2698;
assign w1147 = w10114 & w10122;
assign w1148 = w3288 & ~w10182;
assign w1149 = w9708 & w11128;
assign w1150 = ~w7783 & ~w2538;
assign w1151 = ~w4700 & w13937;
assign w1152 = w7213 & w6505;
assign w1153 = (w9817 & w6986) | (w9817 & w6869) | (w6986 & w6869);
assign w1154 = (w14449 & w7386) | (w14449 & w6205) | (w7386 & w6205);
assign w1155 = (~w1049 & w14053) | (~w1049 & w2863) | (w14053 & w2863);
assign w1156 = (w13771 & w3588) | (w13771 & w5706) | (w3588 & w5706);
assign w1157 = w3508 & ~w2599;
assign w1158 = ~w2144 & w13669;
assign w1159 = (w13792 & w176) | (w13792 & w11645) | (w176 & w11645);
assign w1160 = (~w2939 & w3641) | (~w2939 & w2418) | (w3641 & w2418);
assign w1161 = w9685 & w8462;
assign w1162 = (w254 & w6285) | (w254 & w7916) | (w6285 & w7916);
assign w1163 = w13764 & ~w9638;
assign w1164 = (w8451 & w4871) | (w8451 & w12502) | (w4871 & w12502);
assign w1165 = w5515 & ~w9460;
assign w1166 = ~w1758 & ~w8105;
assign w1167 = w11482 & ~w1561;
assign w1168 = (w8327 & w1349) | (w8327 & w13664) | (w1349 & w13664);
assign w1169 = w5422 & w5785;
assign w1170 = (~w5952 & w6173) | (~w5952 & w10714) | (w6173 & w10714);
assign w1171 = ~w5860 & ~w11488;
assign w1172 = (~w12958 & w14) | (~w12958 & w5386) | (w14 & w5386);
assign w1173 = ~w3448 & w13260;
assign w1174 = ~w10757 & w3963;
assign w1175 = ~w13713 & w11744;
assign w1176 = (~w6301 & w6266) | (~w6301 & w1105) | (w6266 & w1105);
assign w1177 = w11127 & w11922;
assign w1178 = w5115 & ~w532;
assign w1179 = ~w2845 & w4807;
assign w1180 = w14622 & w5687;
assign w1181 = ~w11732 | w10917;
assign w1182 = (w2670 & w8723) | (w2670 & w11143) | (w8723 & w11143);
assign w1183 = w7794 & ~w10017;
assign w1184 = w7512 & w10346;
assign w1185 = w11533 & ~w13820;
assign w1186 = ~w3885 & w7376;
assign w1187 = ~w7782 & w4313;
assign w1188 = (w5794 & w4756) | (w5794 & w7220) | (w4756 & w7220);
assign w1189 = ~w4850 & w7471;
assign w1190 = ~w7690 & w11559;
assign w1191 = (w10625 & w9747) | (w10625 & w5423) | (w9747 & w5423);
assign w1192 = (w5845 & w9756) | (w5845 & w551) | (w9756 & w551);
assign w1193 = ~w7437 & w13953;
assign w1194 = (w8584 & ~w2289) | (w8584 & w10467) | (~w2289 & w10467);
assign w1195 = ~w5742 & ~w3663;
assign w1196 = w3944 & w10393;
assign w1197 = ~w10675 & w9940;
assign w1198 = w9055 & ~w11211;
assign w1199 = w9366 & ~w10145;
assign w1200 = ~w9582 & w4961;
assign w1201 = (~w9305 & w5508) | (~w9305 & w9234) | (w5508 & w9234);
assign w1202 = (~w8295 & ~w1362) | (~w8295 & w9351) | (~w1362 & w9351);
assign w1203 = w3717 & ~w10483;
assign w1204 = (~w3550 & w2322) | (~w3550 & w10940) | (w2322 & w10940);
assign w1205 = ~w2135 & ~w7630;
assign w1206 = ~w2147 & ~w6951;
assign w1207 = (w10477 & w4921) | (w10477 & w3718) | (w4921 & w3718);
assign w1208 = (w12568 & w8747) | (w12568 & w13377) | (w8747 & w13377);
assign w1209 = (w13136 & w4724) | (w13136 & w14611) | (w4724 & w14611);
assign w1210 = ~w7018 & ~w8077;
assign w1211 = ~w1166 & ~w12915;
assign w1212 = (~w4587 & ~w7342) | (~w4587 & w9100) | (~w7342 & w9100);
assign w1213 = ~w1388 & w3531;
assign w1214 = (~w11185 & w6210) | (~w11185 & w4802) | (w6210 & w4802);
assign w1215 = w13103 & w3128;
assign w1216 = w9949 & w11117;
assign w1217 = ~w803 & w12569;
assign w1218 = w7324 & w3039;
assign w1219 = w5526 & w4892;
assign w1220 = ~w13943 & w10057;
assign w1221 = b45 & a45;
assign w1222 = ~w2689 & w1289;
assign w1223 = (w7708 & w12159) | (w7708 & w13091) | (w12159 & w13091);
assign w1224 = ~w11949 & ~w1840;
assign w1225 = ~w1782 & ~w8019;
assign w1226 = w5282 & w968;
assign w1227 = ~w9541 & w11377;
assign w1228 = (~w50 & w9324) | (~w50 & w14226) | (w9324 & w14226);
assign w1229 = ~w884 & ~w4359;
assign w1230 = w9944 & w4419;
assign w1231 = ~w4029 & w14083;
assign w1232 = (w12460 & ~w6506) | (w12460 & w7358) | (~w6506 & w7358);
assign w1233 = (w5110 & w5235) | (w5110 & ~w2582) | (w5235 & ~w2582);
assign w1234 = ~w12505 & w1637;
assign w1235 = ~w13531 & ~w9226;
assign w1236 = (w14512 & w9012) | (w14512 & w4773) | (w9012 & w4773);
assign w1237 = (~w2675 & w9747) | (~w2675 & w2241) | (w9747 & w2241);
assign w1238 = w14417 & w12065;
assign w1239 = w3563 | w217;
assign w1240 = w6219 & ~w4312;
assign w1241 = (~w965 & w3232) | (~w965 & w3617) | (w3232 & w3617);
assign w1242 = (~w7645 & w7688) | (~w7645 & w1468) | (w7688 & w1468);
assign w1243 = (w12142 & w14439) | (w12142 & w8282) | (w14439 & w8282);
assign w1244 = ~w8234 & w1821;
assign w1245 = (w11500 & w7342) | (w11500 & w4394) | (w7342 & w4394);
assign w1246 = w9846 & w7670;
assign w1247 = w6572 & w7423;
assign w1248 = (~w12569 & w7531) | (~w12569 & w4964) | (w7531 & w4964);
assign w1249 = (w4239 & w7440) | (w4239 & w217) | (w7440 & w217);
assign w1250 = ~w6052 & ~w8639;
assign w1251 = w12859 & w4091;
assign w1252 = w2050 & w7350;
assign w1253 = ~w8906 & ~w764;
assign w1254 = ~w9747 & w5412;
assign w1255 = ~w13620 & w1712;
assign w1256 = ~w10441 & ~w9211;
assign w1257 = (w11117 & w10486) | (w11117 & w11464) | (w10486 & w11464);
assign w1258 = w2698 & w1855;
assign w1259 = w9645 & w4765;
assign w1260 = w5767 & w14486;
assign w1261 = w4934 & w13948;
assign w1262 = (~w654 & ~w10712) | (~w654 & w347) | (~w10712 & w347);
assign w1263 = ~w12170 & ~w13531;
assign w1264 = w12170 & w7722;
assign w1265 = ~w1384 & w9316;
assign w1266 = w13839 & w2851;
assign w1267 = (~w7234 & w6555) | (~w7234 & w7810) | (w6555 & w7810);
assign w1268 = (w2598 & ~w5253) | (w2598 & w5951) | (~w5253 & w5951);
assign w1269 = w10037 & ~w11383;
assign w1270 = (~w5490 & w14538) | (~w5490 & w11624) | (w14538 & w11624);
assign w1271 = (~w5753 & w12010) | (~w5753 & w9665) | (w12010 & w9665);
assign w1272 = (w3812 & ~w7365) | (w3812 & w12988) | (~w7365 & w12988);
assign w1273 = (~w12915 & w10462) | (~w12915 & w5589) | (w10462 & w5589);
assign w1274 = w1873 & w9087;
assign w1275 = ~w6663 & w13022;
assign w1276 = ~w10245 & w14525;
assign w1277 = w3540 & ~w11589;
assign w1278 = (w3435 & w183) | (w3435 & w2443) | (w183 & w2443);
assign w1279 = w6918 & ~w8279;
assign w1280 = (w6802 & w2131) | (w6802 & w14117) | (w2131 & w14117);
assign w1281 = (w7243 & w1495) | (w7243 & ~w13309) | (w1495 & ~w13309);
assign w1282 = (w3502 & w2029) | (w3502 & w8995) | (w2029 & w8995);
assign w1283 = (~w11345 & w5224) | (~w11345 & w7980) | (w5224 & w7980);
assign w1284 = w3550 & w564;
assign w1285 = ~w11897 & ~w2295;
assign w1286 = w13993 & w4193;
assign w1287 = w9940 & w8513;
assign w1288 = (~w9305 & w4775) | (~w9305 & w3193) | (w4775 & w3193);
assign w1289 = w9837 & w2897;
assign w1290 = w12464 & w12398;
assign w1291 = w4312 & w4287;
assign w1292 = ~w2463 & w10543;
assign w1293 = w5778 & w719;
assign w1294 = ~w6439 & w8537;
assign w1295 = ~w443 & w1804;
assign w1296 = w12271 & w11902;
assign w1297 = ~w9066 & w4219;
assign w1298 = (w12112 & w3122) | (w12112 & w8626) | (w3122 & w8626);
assign w1299 = w1845 & ~w11117;
assign w1300 = (w3615 & ~w7662) | (w3615 & w12446) | (~w7662 & w12446);
assign w1301 = ~w644 & ~w3479;
assign w1302 = ~w183 & w5906;
assign w1303 = ~w8226 & w12827;
assign w1304 = (~w1642 & w4050) | (~w1642 & w2981) | (w4050 & w2981);
assign w1305 = b7 & a7;
assign w1306 = (~w14395 & ~w8389) | (~w14395 & w5225) | (~w8389 & w5225);
assign w1307 = ~w9805 & ~w6533;
assign w1308 = w8253 & w646;
assign w1309 = w9602 & w2580;
assign w1310 = w3956 & ~w9614;
assign w1311 = w8459 & ~w6234;
assign w1312 = ~w7914 & ~w3885;
assign w1313 = w8900 & ~w11096;
assign w1314 = ~w3139 & w2466;
assign w1315 = ~w7958 & ~w2683;
assign w1316 = (w11201 & w667) | (w11201 & w12436) | (w667 & w12436);
assign w1317 = ~w7905 & w4657;
assign w1318 = (~w6362 & w12478) | (~w6362 & w12006) | (w12478 & w12006);
assign w1319 = (~w8171 & w4182) | (~w8171 & ~w10272) | (w4182 & ~w10272);
assign w1320 = (w8168 & w8522) | (w8168 & w3789) | (w8522 & w3789);
assign w1321 = w7794 & w5325;
assign w1322 = ~w1758 & ~w10334;
assign w1323 = (~w9093 & w12644) | (~w9093 & w478) | (w12644 & w478);
assign w1324 = w9454 & ~w3830;
assign w1325 = w607 & ~w6500;
assign w1326 = w10396 & w8591;
assign w1327 = w4307 & ~w9506;
assign w1328 = (~w4512 & w14219) | (~w4512 & w1736) | (w14219 & w1736);
assign w1329 = ~w12514 & w7721;
assign w1330 = w3449 & w6382;
assign w1331 = w3039 & w1506;
assign w1332 = ~w12481 & w13839;
assign w1333 = w11184 & w5420;
assign w1334 = (w1416 & w6276) | (w1416 & w8228) | (w6276 & w8228);
assign w1335 = ~w10517 & w11899;
assign w1336 = ~w9284 & w2941;
assign w1337 = w7747 & w13575;
assign w1338 = (w3727 & ~w1900) | (w3727 & w4118) | (~w1900 & w4118);
assign w1339 = (w4545 & w4082) | (w4545 & w5011) | (w4082 & w5011);
assign w1340 = ~w3435 & w8886;
assign w1341 = ~w834 & ~w5764;
assign w1342 = (w10115 & w14018) | (w10115 & w8590) | (w14018 & w8590);
assign w1343 = ~w5522 & ~w4458;
assign w1344 = ~w10847 & w12883;
assign w1345 = ~w13222 & w13733;
assign w1346 = (~w1171 & w13122) | (~w1171 & w12887) | (w13122 & w12887);
assign w1347 = w841 & w7841;
assign w1348 = (w5090 & w220) | (w5090 & w8194) | (w220 & w8194);
assign w1349 = ~w5419 & w11454;
assign w1350 = ~w3484 & w9771;
assign w1351 = (~w142 & ~w3550) | (~w142 & w14491) | (~w3550 & w14491);
assign w1352 = ~w11444 & w3142;
assign w1353 = (~w5483 & w296) | (~w5483 & w12402) | (w296 & w12402);
assign w1354 = (~w6825 & w3480) | (~w6825 & w926) | (w3480 & w926);
assign w1355 = w4322 & w5912;
assign w1356 = (w9244 & w12060) | (w9244 & w5439) | (w12060 & w5439);
assign w1357 = ~w8290 & ~w13820;
assign w1358 = ~w7000 & ~w10703;
assign w1359 = (w13287 & w1971) | (w13287 & w11813) | (w1971 & w11813);
assign w1360 = ~w5879 & ~w11476;
assign w1361 = ~w1563 & w3717;
assign w1362 = ~w8791 & ~w4607;
assign w1363 = w6427 & ~w2410;
assign w1364 = w7013 & w11117;
assign w1365 = (~w13462 & w8965) | (~w13462 & w2690) | (w8965 & w2690);
assign w1366 = (w7417 & w10563) | (w7417 & ~w2362) | (w10563 & ~w2362);
assign w1367 = w5489 & w4237;
assign w1368 = ~w9786 & w1070;
assign w1369 = ~w9097 & ~w5113;
assign w1370 = ~w2256 & ~w9464;
assign w1371 = ~w6897 & w2171;
assign w1372 = ~w1812 & w10765;
assign w1373 = (~w8534 & w10732) | (~w8534 & w13316) | (w10732 & w13316);
assign w1374 = ~w4043 & ~w7949;
assign w1375 = w7973 & w1000;
assign w1376 = ~w12163 & ~w612;
assign w1377 = (~w10884 & ~w9249) | (~w10884 & w8447) | (~w9249 & w8447);
assign w1378 = w2451 & w9690;
assign w1379 = (w5020 & w11562) | (w5020 & w12303) | (w11562 & w12303);
assign w1380 = w7267 & w11507;
assign w1381 = w7808 & w5223;
assign w1382 = ~w5522 & ~w7670;
assign w1383 = w9454 & w4375;
assign w1384 = w5772 & ~w13864;
assign w1385 = (~w2998 & w4099) | (~w2998 & w11120) | (w4099 & w11120);
assign w1386 = (~w8540 & w9012) | (~w8540 & w2426) | (w9012 & w2426);
assign w1387 = ~w3025 & ~w3215;
assign w1388 = (~w4796 & w1692) | (~w4796 & w11636) | (w1692 & w11636);
assign w1389 = w9087 & w9938;
assign w1390 = w4191 & w5634;
assign w1391 = w10221 & ~w3904;
assign w1392 = ~w9608 & w11489;
assign w1393 = w11500 & w13008;
assign w1394 = (~w4287 & w2971) | (~w4287 & ~w7999) | (w2971 & ~w7999);
assign w1395 = ~w1821 & ~w13976;
assign w1396 = ~w4958 & ~w12542;
assign w1397 = ~w14141 & w7366;
assign w1398 = ~w4099 & w6348;
assign w1399 = ~w12240 & w6113;
assign w1400 = (w8497 & w1741) | (w8497 & w12376) | (w1741 & w12376);
assign w1401 = w1323 & ~w2743;
assign w1402 = ~w2837 & w13211;
assign w1403 = w5532 & ~w4127;
assign w1404 = ~w7261 & ~w14412;
assign w1405 = (~w6233 & w10652) | (~w6233 & w13273) | (w10652 & w13273);
assign w1406 = ~w9781 & ~w13408;
assign w1407 = ~w10748 & ~w5823;
assign w1408 = ~w2858 & w12311;
assign w1409 = (w2331 & w8087) | (w2331 & w6802) | (w8087 & w6802);
assign w1410 = w3914 & w3036;
assign w1411 = w10725 & w3564;
assign w1412 = w5788 & ~w14584;
assign w1413 = ~w10190 & ~w8703;
assign w1414 = w5015 & ~w8598;
assign w1415 = (~w1199 & w13462) | (~w1199 & w13385) | (w13462 & w13385);
assign w1416 = (~w7538 & ~w7240) | (~w7538 & ~w9096) | (~w7240 & ~w9096);
assign w1417 = ~w1821 & w12460;
assign w1418 = ~w10942 & ~w3049;
assign w1419 = ~w10435 & w13945;
assign w1420 = (w347 & ~w1712) | (w347 & w4047) | (~w1712 & w4047);
assign w1421 = (w9305 & w1316) | (w9305 & w1670) | (w1316 & w1670);
assign w1422 = (~w11488 & w2500) | (~w11488 & w10498) | (w2500 & w10498);
assign w1423 = w3786 & w9296;
assign w1424 = ~w5867 & ~w2850;
assign w1425 = ~w13378 & w13648;
assign w1426 = w8335 & w1225;
assign w1427 = (w3452 & w8426) | (w3452 & ~w12376) | (w8426 & ~w12376);
assign w1428 = (~w9138 & w9747) | (~w9138 & w13171) | (w9747 & w13171);
assign w1429 = w7505 & w13086;
assign w1430 = ~w4084 & w5043;
assign w1431 = ~w1166 & w12868;
assign w1432 = w9817 & ~w10301;
assign w1433 = ~w11375 & w616;
assign w1434 = (~w11313 & ~w7248) | (~w11313 & w10990) | (~w7248 & w10990);
assign w1435 = ~w7954 & ~w6381;
assign w1436 = (~w318 & w2470) | (~w318 & w8814) | (w2470 & w8814);
assign w1437 = w607 & w5282;
assign w1438 = (w4370 & w7201) | (w4370 & w8228) | (w7201 & w8228);
assign w1439 = ~w7001 & ~w3727;
assign w1440 = (~w5528 & w6915) | (~w5528 & w8930) | (w6915 & w8930);
assign w1441 = ~w240 & w2669;
assign w1442 = ~w12170 & w13873;
assign w1443 = w4006 & ~w2221;
assign w1444 = (w8106 & w12235) | (w8106 & w12907) | (w12235 & w12907);
assign w1445 = ~w10042 & ~w3380;
assign w1446 = w3858 & ~w3026;
assign w1447 = w8430 & w14201;
assign w1448 = ~w12591 & w2456;
assign w1449 = w4433 & w8631;
assign w1450 = w12550 & ~w4304;
assign w1451 = w13357 & ~w725;
assign w1452 = (w12210 & ~w12312) | (w12210 & w11782) | (~w12312 & w11782);
assign w1453 = ~w12240 & w3098;
assign w1454 = (w3388 & w14586) | (w3388 & w8282) | (w14586 & w8282);
assign w1455 = ~w10523 & ~w13590;
assign w1456 = w12771 | w1455;
assign w1457 = ~w12546 & w2536;
assign w1458 = (w1274 & ~w12240) | (w1274 & w3750) | (~w12240 & w3750);
assign w1459 = (~w13135 & ~w1868) | (~w13135 & w3225) | (~w1868 & w3225);
assign w1460 = w11755 & w5578;
assign w1461 = (~w7782 & w1371) | (~w7782 & w3749) | (w1371 & w3749);
assign w1462 = ~w1563 & w2425;
assign w1463 = ~w922 & w13328;
assign w1464 = ~w12976 & w10994;
assign w1465 = w14276 & w12642;
assign w1466 = w4359 & ~w9244;
assign w1467 = (w13018 & w7566) | (w13018 & w5413) | (w7566 & w5413);
assign w1468 = w12460 & w8724;
assign w1469 = ~w884 & w3823;
assign w1470 = ~w3716 & w8888;
assign w1471 = (w2403 & w10738) | (w2403 & w3838) | (w10738 & w3838);
assign w1472 = w5842 & w8719;
assign w1473 = ~w8171 & w1156;
assign w1474 = ~b97 & ~a97;
assign w1475 = w1773 & w650;
assign w1476 = w14555 & w9768;
assign w1477 = ~w8226 & w12126;
assign w1478 = w10036 & w2698;
assign w1479 = w9170 & w7936;
assign w1480 = ~w11261 & w10936;
assign w1481 = ~w934 & ~w712;
assign w1482 = w2680 & w8900;
assign w1483 = ~w4315 & ~w13439;
assign w1484 = w8737 | w12332;
assign w1485 = ~w11287 & w14499;
assign w1486 = (~w4512 & w8331) | (~w4512 & w9561) | (w8331 & w9561);
assign w1487 = ~w3243 & ~w13875;
assign w1488 = (~w235 & w1722) | (~w235 & w7312) | (w1722 & w7312);
assign w1489 = ~w12858 & w6008;
assign w1490 = w1140 & w13299;
assign w1491 = ~w2045 & w858;
assign w1492 = ~w2217 & w12038;
assign w1493 = w10757 & ~w988;
assign w1494 = ~w8234 & w3508;
assign w1495 = ~w7217 & w11336;
assign w1496 = (w11753 & w6243) | (w11753 & w9079) | (w6243 & w9079);
assign w1497 = w8931 & w13994;
assign w1498 = w12575 & w14504;
assign w1499 = ~w8226 & w13480;
assign w1500 = ~w9613 & ~w873;
assign w1501 = ~w1503 & w4204;
assign w1502 = (w7082 & w13267) | (w7082 & w13505) | (w13267 & w13505);
assign w1503 = ~w4033 & w7111;
assign w1504 = (~w5094 & ~w10123) | (~w5094 & w10579) | (~w10123 & w10579);
assign w1505 = (~w806 & w10126) | (~w806 & w3145) | (w10126 & w3145);
assign w1506 = w3038 & ~w8827;
assign w1507 = ~w852 & ~w9227;
assign w1508 = ~w5624 & ~w14125;
assign w1509 = w11041 & ~w9961;
assign w1510 = ~w13208 & w12575;
assign w1511 = ~w13277 & ~w11587;
assign w1512 = w14382 & ~w3209;
assign w1513 = ~w6339 & ~w410;
assign w1514 = ~w2463 & w14299;
assign w1515 = w11997 & w1707;
assign w1516 = ~b34 & ~a34;
assign w1517 = w6190 & w5218;
assign w1518 = ~w4610 & ~w13841;
assign w1519 = ~w5702 & w5826;
assign w1520 = ~w5522 & w3427;
assign w1521 = ~w4099 & w7208;
assign w1522 = w11906 & ~w12945;
assign w1523 = ~w12656 & w12936;
assign w1524 = w9748 & ~w8477;
assign w1525 = (w4622 & w7470) | (w4622 & ~w7031) | (w7470 & ~w7031);
assign w1526 = w9123 & ~w5449;
assign w1527 = ~w2742 & ~w13181;
assign w1528 = (~w9012 & w4083) | (~w9012 & w4351) | (w4083 & w4351);
assign w1529 = ~w7376 & ~w3175;
assign w1530 = ~w640 & ~w9952;
assign w1531 = ~w10040 & w3377;
assign w1532 = ~w4117 & ~w9253;
assign w1533 = (w9305 & w5404) | (w9305 & w1339) | (w5404 & w1339);
assign w1534 = ~w12450 & w8369;
assign w1535 = ~w1119 & ~w2014;
assign w1536 = w309 & ~w12065;
assign w1537 = (~w3502 & w1166) | (~w3502 & w8085) | (w1166 & w8085);
assign w1538 = w13229 & w1489;
assign w1539 = w14395 & ~w2118;
assign w1540 = ~w6135 & ~w7889;
assign w1541 = w7486 & ~w5282;
assign w1542 = (~w5635 & ~w5708) | (~w5635 & w1112) | (~w5708 & w1112);
assign w1543 = (~w3893 & w1712) | (~w3893 & w7678) | (w1712 & w7678);
assign w1544 = ~w1797 & ~w14388;
assign w1545 = b53 & ~w13282;
assign w1546 = (w9305 & w8383) | (w9305 & w3571) | (w8383 & w3571);
assign w1547 = w11583 & ~w7062;
assign w1548 = (w4479 & w1856) | (w4479 & w11501) | (w1856 & w11501);
assign w1549 = (w1114 & w9541) | (w1114 & w112) | (w9541 & w112);
assign w1550 = w8346 & w8563;
assign w1551 = (w7457 & w4108) | (w7457 & w12523) | (w4108 & w12523);
assign w1552 = ~w5556 & w6632;
assign w1553 = (w7406 & w13623) | (w7406 & w6966) | (w13623 & w6966);
assign w1554 = (w12170 & w4512) | (w12170 & w9135) | (w4512 & w9135);
assign w1555 = (w6716 & ~w12464) | (w6716 & w11103) | (~w12464 & w11103);
assign w1556 = (w10523 & ~w7737) | (w10523 & ~w11586) | (~w7737 & ~w11586);
assign w1557 = ~w3885 & ~w5778;
assign w1558 = ~w1563 & ~w9004;
assign w1559 = ~w11429 & ~w3209;
assign w1560 = (~w10213 & w9963) | (~w10213 & ~w1928) | (w9963 & ~w1928);
assign w1561 = w5867 & ~w6554;
assign w1562 = ~w10084 & ~w6458;
assign w1563 = ~w3346 & ~w3542;
assign w1564 = ~w829 & w13620;
assign w1565 = w5020 & w3801;
assign w1566 = w13924 & w5914;
assign w1567 = ~w14302 & ~w13481;
assign w1568 = ~w14660 & w10807;
assign w1569 = w10317 & w7376;
assign w1570 = ~w9032 & ~w2698;
assign w1571 = (w8168 & w2003) | (w8168 & w4940) | (w2003 & w4940);
assign w1572 = (~w13587 & w13060) | (~w13587 & w8485) | (w13060 & w8485);
assign w1573 = (w6387 & w9437) | (w6387 & w3731) | (w9437 & w3731);
assign w1574 = w9560 & w4927;
assign w1575 = ~w5867 & ~w1052;
assign w1576 = (w12952 & w9174) | (w12952 & ~w12293) | (w9174 & ~w12293);
assign w1577 = ~w254 & w3013;
assign w1578 = ~w4500 & ~w8099;
assign w1579 = w5805 & ~w10105;
assign w1580 = ~w9087 & w9430;
assign w1581 = w5757 & w6721;
assign w1582 = w6093 & ~w13350;
assign w1583 = (w5952 & w568) | (w5952 & w14289) | (w568 & w14289);
assign w1584 = w6739 & w7690;
assign w1585 = (~w1665 & w6239) | (~w1665 & w2657) | (w6239 & w2657);
assign w1586 = w11023 & ~w3781;
assign w1587 = ~w3502 & ~w8512;
assign w1588 = ~w9150 & w13662;
assign w1589 = ~w9608 & w8342;
assign w1590 = (w11211 & w2147) | (w11211 & w4292) | (w2147 & w4292);
assign w1591 = w187 & w9077;
assign w1592 = (~w4545 & w12501) | (~w4545 & w4675) | (w12501 & w4675);
assign w1593 = (w3556 & w12145) | (w3556 & w9034) | (w12145 & w9034);
assign w1594 = (~w378 & w368) | (~w378 & w10232) | (w368 & w10232);
assign w1595 = (w11327 & w13213) | (w11327 & w2457) | (w13213 & w2457);
assign w1596 = (w9608 & w12236) | (w9608 & w2862) | (w12236 & w2862);
assign w1597 = w11070 & w8872;
assign w1598 = ~w4700 & w13323;
assign w1599 = ~w4401 & ~w3098;
assign w1600 = w1607 & w10532;
assign w1601 = w11560 & ~w3427;
assign w1602 = ~w5867 & w6542;
assign w1603 = (~w326 & w467) | (~w326 & w4346) | (w467 & w4346);
assign w1604 = (~w14463 & w1526) | (~w14463 & w4306) | (w1526 & w4306);
assign w1605 = (~w5532 & w13122) | (~w5532 & w2796) | (w13122 & w2796);
assign w1606 = w6436 & ~w12642;
assign w1607 = w8886 & w7135;
assign w1608 = ~w8742 & ~w9006;
assign w1609 = w1087 & ~w2096;
assign w1610 = w2924 & w13210;
assign w1611 = ~w5035 & ~w13820;
assign w1612 = (~w4612 & ~w9537) | (~w4612 & w12092) | (~w9537 & w12092);
assign w1613 = ~w13526 & ~w2663;
assign w1614 = ~w5852 & ~b93;
assign w1615 = ~w3957 & ~w6929;
assign w1616 = ~w10766 & w12443;
assign w1617 = ~w183 & w9226;
assign w1618 = w967 & ~w11986;
assign w1619 = (~w3025 & w3906) | (~w3025 & w11732) | (w3906 & w11732);
assign w1620 = (~w3098 & ~w1140) | (~w3098 & w13667) | (~w1140 & w13667);
assign w1621 = (~w1498 & w14141) | (~w1498 & w14032) | (w14141 & w14032);
assign w1622 = ~w10483 & ~w2142;
assign w1623 = ~w7455 & ~w911;
assign w1624 = ~w9607 & w4541;
assign w1625 = (~w2081 & w12122) | (~w2081 & w12720) | (w12122 & w12720);
assign w1626 = w3809 & w11708;
assign w1627 = ~w9012 & w3213;
assign w1628 = ~w8977 & ~w1340;
assign w1629 = ~w1503 & w11725;
assign w1630 = ~w7213 & ~w11560;
assign w1631 = w9679 & ~w4447;
assign w1632 = (~w2858 & w4099) | (~w2858 & w10489) | (w4099 & w10489);
assign w1633 = w3943 & ~w6387;
assign w1634 = (w378 & w13539) | (w378 & w8798) | (w13539 & w8798);
assign w1635 = ~w12240 & w7668;
assign w1636 = (~w11629 & ~w11202) | (~w11629 & w74) | (~w11202 & w74);
assign w1637 = (~w7782 & w12058) | (~w7782 & w270) | (w12058 & w270);
assign w1638 = ~w11726 & ~w5738;
assign w1639 = w7400 & ~w7410;
assign w1640 = (w6637 & w2659) | (w6637 & w5019) | (w2659 & w5019);
assign w1641 = (~w12231 & w14369) | (~w12231 & w11110) | (w14369 & w11110);
assign w1642 = ~w4190 & ~w7513;
assign w1643 = (~w142 & ~w2701) | (~w142 & w6872) | (~w2701 & w6872);
assign w1644 = w4221 & w6315;
assign w1645 = w10872 & ~w6281;
assign w1646 = ~w2922 & ~w8047;
assign w1647 = (~w2335 & w5916) | (~w2335 & w6202) | (w5916 & w6202);
assign w1648 = (~w11321 & w2568) | (~w11321 & w2969) | (w2568 & w2969);
assign w1649 = (w3508 & ~w6391) | (w3508 & w5472) | (~w6391 & w5472);
assign w1650 = (~w6162 & w6723) | (~w6162 & w10953) | (w6723 & w10953);
assign w1651 = w279 & w1997;
assign w1652 = ~w2464 & ~w11031;
assign w1653 = w3714 & ~w5664;
assign w1654 = ~w10334 & ~w14285;
assign w1655 = w12088 & w2680;
assign w1656 = w75 & ~w2619;
assign w1657 = ~w11081 & w2847;
assign w1658 = (~w12893 & w298) | (~w12893 & w67) | (w298 & w67);
assign w1659 = w14491 & ~w3963;
assign w1660 = ~w80 & ~w1624;
assign w1661 = (~w8327 & w2054) | (~w8327 & w8251) | (w2054 & w8251);
assign w1662 = (w9227 & w12041) | (w9227 & w12713) | (w12041 & w12713);
assign w1663 = (~w9305 & w9082) | (~w9305 & w12975) | (w9082 & w12975);
assign w1664 = ~w7931 & w10080;
assign w1665 = (w13531 & w11261) | (w13531 & w9483) | (w11261 & w9483);
assign w1666 = ~w2844 & ~w9506;
assign w1667 = ~b1 & ~a1;
assign w1668 = w12481 & w1062;
assign w1669 = ~w2218 & w7777;
assign w1670 = (w8405 & w12916) | (w8405 & w3196) | (w12916 & w3196);
assign w1671 = w10174 & w7709;
assign w1672 = w7681 & w11934;
assign w1673 = w5005 & ~w8262;
assign w1674 = w386 & w8048;
assign w1675 = w211 & w5865;
assign w1676 = ~w916 & ~w1418;
assign w1677 = w7354 & ~w13854;
assign w1678 = ~w14664 & w615;
assign w1679 = ~w12893 & w9286;
assign w1680 = ~w1540 & w5785;
assign w1681 = ~w7447 & ~w5560;
assign w1682 = ~b110 & ~a110;
assign w1683 = (~w9713 & ~w9013) | (~w9713 & w10228) | (~w9013 & w10228);
assign w1684 = ~w14500 & ~w7909;
assign w1685 = ~w6309 & w3752;
assign w1686 = w7612 & ~w2311;
assign w1687 = w1186 & w5884;
assign w1688 = ~w11429 & w9565;
assign w1689 = (~w9928 & w8163) | (~w9928 & w12937) | (w8163 & w12937);
assign w1690 = ~w11004 & w5470;
assign w1691 = ~w118 & ~w5652;
assign w1692 = ~w2094 & ~w1204;
assign w1693 = w12662 & w4334;
assign w1694 = ~w4714 & ~w892;
assign w1695 = ~w1382 & ~w10474;
assign w1696 = ~w4050 & w4382;
assign w1697 = ~w5191 & ~w5633;
assign w1698 = ~w13122 & ~w6242;
assign w1699 = ~w8035 & ~w5693;
assign w1700 = ~w7645 & ~w9107;
assign w1701 = ~w2317 & w516;
assign w1702 = w3502 & ~w852;
assign w1703 = ~w7904 & w5963;
assign w1704 = (~w10923 & w6847) | (~w10923 & w8496) | (w6847 & w8496);
assign w1705 = w10124 & w35;
assign w1706 = ~w10517 & ~w11861;
assign w1707 = (w4855 & ~w2500) | (w4855 & w11365) | (~w2500 & w11365);
assign w1708 = w13628 & w2962;
assign w1709 = ~w13349 & w12707;
assign w1710 = (~w12807 & w10858) | (~w12807 & w310) | (w10858 & w310);
assign w1711 = w14293 & ~w10245;
assign w1712 = ~w2176 & ~w397;
assign w1713 = w3914 & ~w6045;
assign w1714 = w8047 & w1036;
assign w1715 = w14545 & ~w13922;
assign w1716 = w8949 & w6464;
assign w1717 = w7159 & ~w12431;
assign w1718 = ~w3969 & w4960;
assign w1719 = ~w254 & w2597;
assign w1720 = (~w3158 & ~w9748) | (~w3158 & w4932) | (~w9748 & w4932);
assign w1721 = (w3973 & w13067) | (w3973 & ~w9034) | (w13067 & ~w9034);
assign w1722 = (~w235 & w12664) | (~w235 & w13249) | (w12664 & w13249);
assign w1723 = (w2116 & w1652) | (w2116 & w2724) | (w1652 & w2724);
assign w1724 = ~w13668 & w8812;
assign w1725 = w12433 & ~w7005;
assign w1726 = ~w11049 & w5634;
assign w1727 = ~w8171 & ~w10925;
assign w1728 = (w11500 & w5294) | (w11500 & w6831) | (w5294 & w6831);
assign w1729 = w3242 & w8786;
assign w1730 = ~w5091 & ~w13422;
assign w1731 = (w11744 & w10790) | (w11744 & w2767) | (w10790 & w2767);
assign w1732 = (w9952 & w6250) | (w9952 & w6337) | (w6250 & w6337);
assign w1733 = ~w1491 & ~w9224;
assign w1734 = w5282 & w7889;
assign w1735 = w7981 & ~w3289;
assign w1736 = (w12879 & ~w5294) | (w12879 & w14219) | (~w5294 & w14219);
assign w1737 = (w13685 & w8764) | (w13685 & w6998) | (w8764 & w6998);
assign w1738 = w9646 & ~w3427;
assign w1739 = ~w13713 & w9724;
assign w1740 = (~w7082 & w163) | (~w7082 & w3108) | (w163 & w3108);
assign w1741 = (w10115 & w9783) | (w10115 & w11609) | (w9783 & w11609);
assign w1742 = ~w254 & w2661;
assign w1743 = (~w2073 & ~w988) | (~w2073 & w3766) | (~w988 & w3766);
assign w1744 = ~w9682 & ~w1820;
assign w1745 = ~w4033 & ~w2941;
assign w1746 = ~w2463 & w7408;
assign w1747 = w8431 & w8647;
assign w1748 = ~w10334 & ~w7661;
assign w1749 = ~w12951 & w9069;
assign w1750 = w14178 & ~w4987;
assign w1751 = w473 & ~w9541;
assign w1752 = ~w12479 & ~w13547;
assign w1753 = w3944 & ~w4893;
assign w1754 = w12464 & w8827;
assign w1755 = w14444 & w1020;
assign w1756 = ~w6583 & ~w11361;
assign w1757 = (~w5243 & w3146) | (~w5243 & ~w7644) | (w3146 & ~w7644);
assign w1758 = ~w4700 & w12460;
assign w1759 = (w5414 & w7533) | (w5414 & ~w12376) | (w7533 & ~w12376);
assign w1760 = w12943 & w14280;
assign w1761 = w4503 & ~w2493;
assign w1762 = ~w607 & ~w11861;
assign w1763 = ~w331 & ~w6733;
assign w1764 = w7493 & w2393;
assign w1765 = (w11067 & w4489) | (w11067 & ~w11429) | (w4489 & ~w11429);
assign w1766 = (~w8459 & w8294) | (~w8459 & w4192) | (w8294 & w4192);
assign w1767 = w1772 & w1006;
assign w1768 = (w13332 & ~w10239) | (w13332 & w8202) | (~w10239 & w8202);
assign w1769 = ~w6836 & ~w2564;
assign w1770 = w1114 & w11744;
assign w1771 = (w6563 & w12862) | (w6563 & w10240) | (w12862 & w10240);
assign w1772 = (w7966 & ~w1697) | (w7966 & w9270) | (~w1697 & w9270);
assign w1773 = (w9803 & w2741) | (w9803 & w650) | (w2741 & w650);
assign w1774 = (w12856 & w10462) | (w12856 & w12561) | (w10462 & w12561);
assign w1775 = ~w9601 & ~w9198;
assign w1776 = w11275 & w6997;
assign w1777 = (w4073 & w3934) | (w4073 & ~w2868) | (w3934 & ~w2868);
assign w1778 = (w11803 & w3272) | (w11803 & w10780) | (w3272 & w10780);
assign w1779 = w5556 & ~w6542;
assign w1780 = w9679 & ~w2208;
assign w1781 = (w11417 & w13122) | (w11417 & w2265) | (w13122 & w2265);
assign w1782 = w7305 & ~w8396;
assign w1783 = w100 & ~w10399;
assign w1784 = w13452 & ~w2983;
assign w1785 = w1116 & ~w12033;
assign w1786 = ~w1821 & w10551;
assign w1787 = w2938 & w2493;
assign w1788 = ~w2660 & ~w4499;
assign w1789 = (~w5845 & w11240) | (~w5845 & w5857) | (w11240 & w5857);
assign w1790 = ~w4460 & ~w5303;
assign w1791 = w12577 & ~w215;
assign w1792 = w13830 & ~w3842;
assign w1793 = w10951 & ~w14517;
assign w1794 = ~w12065 & ~w621;
assign w1795 = (~w7190 & ~w9672) | (~w7190 & w5307) | (~w9672 & w5307);
assign w1796 = w6113 & ~w5664;
assign w1797 = w6113 & ~w5845;
assign w1798 = (~w2762 & w3982) | (~w2762 & w5538) | (w3982 & w5538);
assign w1799 = (~w6080 & w1335) | (~w6080 & w8529) | (w1335 & w8529);
assign w1800 = ~w9256 & ~w13652;
assign w1801 = (~w1362 & w13278) | (~w1362 & w12750) | (w13278 & w12750);
assign w1802 = b106 & a106;
assign w1803 = ~w4429 & w7142;
assign w1804 = w11364 & ~w3017;
assign w1805 = ~w12662 & ~w11159;
assign w1806 = (w3740 & w7562) | (w3740 & w11180) | (w7562 & w11180);
assign w1807 = ~w1828 & w12382;
assign w1808 = ~w11429 & w8958;
assign w1809 = (~w10704 & w2270) | (~w10704 & w12365) | (w2270 & w12365);
assign w1810 = (w14259 & ~w5189) | (w14259 & w539) | (~w5189 & w539);
assign w1811 = w607 & w1062;
assign w1812 = (~w12416 & w8755) | (~w12416 & w3565) | (w8755 & w3565);
assign w1813 = ~w2848 & w7674;
assign w1814 = ~w5219 & w1486;
assign w1815 = ~w8110 & w4071;
assign w1816 = w10045 & w13341;
assign w1817 = w2135 & w7722;
assign w1818 = ~w11547 & w7155;
assign w1819 = ~w309 & ~w4017;
assign w1820 = ~w2317 & w1361;
assign w1821 = ~b93 & ~a93;
assign w1822 = ~w719 & w13981;
assign w1823 = ~w13152 & w4935;
assign w1824 = w13423 & ~w1540;
assign w1825 = ~w2933 & ~w10514;
assign w1826 = ~w5177 & w2320;
assign w1827 = (w804 & w1969) | (w804 & w7321) | (w1969 & w7321);
assign w1828 = ~w10930 & ~w10195;
assign w1829 = w5867 & w13713;
assign w1830 = (~w7782 & w7539) | (~w7782 & w4880) | (w7539 & w4880);
assign w1831 = w14526 & w7645;
assign w1832 = (~w8937 & w11521) | (~w8937 & w766) | (w11521 & w766);
assign w1833 = ~w10547 & w6376;
assign w1834 = w5397 & w14417;
assign w1835 = (w13755 & w9639) | (w13755 & w4051) | (w9639 & w4051);
assign w1836 = w7668 & ~w5845;
assign w1837 = (w9541 & w4577) | (w9541 & w1412) | (w4577 & w1412);
assign w1838 = ~b109 & ~a109;
assign w1839 = ~w12088 & w11193;
assign w1840 = ~w5271 & ~w2859;
assign w1841 = ~w499 & w8769;
assign w1842 = ~w12958 & ~w2387;
assign w1843 = (~w4739 & w4638) | (~w4739 & w13478) | (w4638 & w13478);
assign w1844 = ~w254 & w11595;
assign w1845 = ~w7369 & ~w8253;
assign w1846 = ~w4881 & ~w6975;
assign w1847 = ~w8388 & ~w6716;
assign w1848 = (w4996 & ~w6755) | (w4996 & w292) | (~w6755 & w292);
assign w1849 = (w6802 & w5727) | (w6802 & w13984) | (w5727 & w13984);
assign w1850 = w2310 | w4432;
assign w1851 = (~w13685 & w3860) | (~w13685 & w7802) | (w3860 & w7802);
assign w1852 = (w5865 & ~w9541) | (w5865 & w5690) | (~w9541 & w5690);
assign w1853 = (~w10722 & w12626) | (~w10722 & w1999) | (w12626 & w1999);
assign w1854 = w5522 & w6689;
assign w1855 = w1498 & w10590;
assign w1856 = w3153 & w14579;
assign w1857 = w4269 & ~w2387;
assign w1858 = ~w8422 & w10281;
assign w1859 = (w11655 & w12347) | (w11655 & ~w9034) | (w12347 & ~w9034);
assign w1860 = w7464 & ~w4287;
assign w1861 = w13190 & ~w5079;
assign w1862 = ~w10075 & ~w7851;
assign w1863 = (w7578 & w8770) | (w7578 & w1689) | (w8770 & w1689);
assign w1864 = ~w12606 & w8356;
assign w1865 = ~w4309 & w11594;
assign w1866 = ~w10853 & w1240;
assign w1867 = (w3682 & w5609) | (w3682 & w1262) | (w5609 & w1262);
assign w1868 = w4399 & w7295;
assign w1869 = ~w5845 & ~w2858;
assign w1870 = ~w11745 & ~w13937;
assign w1871 = ~w10523 & w12545;
assign w1872 = (~w4134 & w2306) | (~w4134 & w12820) | (w2306 & w12820);
assign w1873 = ~w7190 & ~w13565;
assign w1874 = ~w980 & ~w5882;
assign w1875 = (w8106 & w9312) | (w8106 & w8866) | (w9312 & w8866);
assign w1876 = (w2816 & w3709) | (w2816 & w12978) | (w3709 & w12978);
assign w1877 = ~w12757 & w537;
assign w1878 = ~w4213 & ~w13152;
assign w1879 = (w10162 & w10123) | (w10162 & w13000) | (w10123 & w13000);
assign w1880 = ~w11197 & ~w938;
assign w1881 = w9133 & w496;
assign w1882 = ~w3233 & w8334;
assign w1883 = ~w9986 & ~w6530;
assign w1884 = (w9454 & ~w1518) | (w9454 & w12965) | (~w1518 & w12965);
assign w1885 = w12656 & w4787;
assign w1886 = ~w4111 & w12047;
assign w1887 = ~w2358 & ~w356;
assign w1888 = ~w10286 & w3694;
assign w1889 = ~w3682 & ~w11750;
assign w1890 = (w3764 & w5562) | (w3764 & w8365) | (w5562 & w8365);
assign w1891 = (~w217 & ~w4757) | (~w217 & w7036) | (~w4757 & w7036);
assign w1892 = w8057 & w1401;
assign w1893 = (w4363 & w11919) | (w4363 & w904) | (w11919 & w904);
assign w1894 = w2656 & ~w7879;
assign w1895 = (w8459 & w1629) | (w8459 & w6843) | (w1629 & w6843);
assign w1896 = w7888 & w11466;
assign w1897 = (w13013 & ~w1156) | (w13013 & w942) | (~w1156 & w942);
assign w1898 = w8389 & ~w10903;
assign w1899 = (w8205 & w4921) | (w8205 & w2681) | (w4921 & w2681);
assign w1900 = ~w3164 & ~w3949;
assign w1901 = ~w13118 & w2788;
assign w1902 = (~w8938 & ~w10737) | (~w8938 & w13220) | (~w10737 & w13220);
assign w1903 = w9672 & ~w7630;
assign w1904 = w6785 & ~w1601;
assign w1905 = w12459 & ~w616;
assign w1906 = ~b7 & ~a7;
assign w1907 = ~w7376 & ~w4671;
assign w1908 = w6584 & a53;
assign w1909 = ~w974 & ~w6840;
assign w1910 = w227 & w1091;
assign w1911 = (w9608 & w10546) | (w9608 & w10319) | (w10546 & w10319);
assign w1912 = ~w922 & w7772;
assign w1913 = (~w9608 & w3417) | (~w9608 & w2151) | (w3417 & w2151);
assign w1914 = ~w10334 & ~w6620;
assign w1915 = (~w8937 & w3413) | (~w8937 & w11554) | (w3413 & w11554);
assign w1916 = w12531 & w14502;
assign w1917 = (~w11613 & w12985) | (~w11613 & w183) | (w12985 & w183);
assign w1918 = ~w12452 & w8379;
assign w1919 = ~w6542 & w10295;
assign w1920 = w12516 & ~w930;
assign w1921 = (~w13306 & w4952) | (~w13306 & ~w1503) | (w4952 & ~w1503);
assign w1922 = ~w5867 & ~w9156;
assign w1923 = w10223 & ~w11902;
assign w1924 = (~w302 & w2534) | (~w302 & w8500) | (w2534 & w8500);
assign w1925 = ~w2029 & w8823;
assign w1926 = ~w12658 & ~w1016;
assign w1927 = (w14527 & w3421) | (w14527 & w9403) | (w3421 & w9403);
assign w1928 = ~w533 & w4655;
assign w1929 = ~w13336 & ~w10874;
assign w1930 = ~w254 & w6037;
assign w1931 = ~w4158 & w9177;
assign w1932 = w11264 & w2592;
assign w1933 = w8171 & w14215;
assign w1934 = w3950 & w6053;
assign w1935 = w12296 & ~w6247;
assign w1936 = w12359 & w7157;
assign w1937 = ~w4213 & ~w536;
assign w1938 = (w12896 & w12027) | (w12896 & w9034) | (w12027 & w9034);
assign w1939 = ~w7749 & ~w1701;
assign w1940 = w9306 & ~w1149;
assign w1941 = ~w12240 & w6716;
assign w1942 = (w12038 & w5553) | (w12038 & w1492) | (w5553 & w1492);
assign w1943 = w8110 & ~w3904;
assign w1944 = ~w2610 & w9607;
assign w1945 = w2747 & w6471;
assign w1946 = ~w493 & ~w6266;
assign w1947 = ~w13635 & w723;
assign w1948 = (w4987 & w9735) | (w4987 & w55) | (w9735 & w55);
assign w1949 = ~w13854 & ~w10704;
assign w1950 = w13189 & w9638;
assign w1951 = w14227 & ~w7906;
assign w1952 = (w992 & ~w1190) | (w992 & ~w6716) | (~w1190 & ~w6716);
assign w1953 = ~w10235 & w2651;
assign w1954 = w8367 & w4987;
assign w1955 = ~w1068 & ~w2460;
assign w1956 = w8878 & w1115;
assign w1957 = ~w13234 & ~w134;
assign w1958 = ~w922 & w3717;
assign w1959 = (~w9733 & w6994) | (~w9733 & w2445) | (w6994 & w2445);
assign w1960 = ~w7525 & w857;
assign w1961 = w13197 & ~w11031;
assign w1962 = w10224 & ~w9226;
assign w1963 = w3553 & ~w11809;
assign w1964 = ~w4921 & w5933;
assign w1965 = w1283 & ~w11117;
assign w1966 = ~w922 & w6652;
assign w1967 = (~w12170 & ~w10676) | (~w12170 & w13953) | (~w10676 & w13953);
assign w1968 = ~w3508 & w499;
assign w1969 = ~w1802 & w11117;
assign w1970 = w4193 & ~w1335;
assign w1971 = (w503 & w4067) | (w503 & w7326) | (w4067 & w7326);
assign w1972 = ~w8937 & w8218;
assign w1973 = (~w7914 & w11658) | (~w7914 & w1312) | (w11658 & w1312);
assign w1974 = (w2218 & w4745) | (w2218 & w7563) | (w4745 & w7563);
assign w1975 = w12569 & w6784;
assign w1976 = (w5491 & w6848) | (w5491 & w2457) | (w6848 & w2457);
assign w1977 = ~w9015 & ~w8085;
assign w1978 = w1263 & w14395;
assign w1979 = w2096 & w8676;
assign w1980 = ~w6761 & ~w7808;
assign w1981 = (w11416 & w10718) | (w11416 & w11270) | (w10718 & w11270);
assign w1982 = ~w11429 & w6680;
assign w1983 = ~w10772 & w3074;
assign w1984 = w7459 & ~w8347;
assign w1985 = w2526 & ~w11981;
assign w1986 = w9170 & w13988;
assign w1987 = w3098 & w13873;
assign w1988 = (~w13587 & w10929) | (~w13587 & w13052) | (w10929 & w13052);
assign w1989 = ~w7082 & ~w3233;
assign w1990 = ~w607 & w11031;
assign w1991 = ~w142 & ~w11117;
assign w1992 = w10949 & w14253;
assign w1993 = w8280 & ~w12642;
assign w1994 = (~w3615 & w11278) | (~w3615 & w3209) | (w11278 & w3209);
assign w1995 = (~w12506 & ~w6689) | (~w12506 & w6357) | (~w6689 & w6357);
assign w1996 = (~w12209 & w11529) | (~w12209 & w12627) | (w11529 & w12627);
assign w1997 = ~w3431 & ~w12787;
assign w1998 = ~w11057 & ~w10527;
assign w1999 = (~w4159 & w5521) | (~w4159 & w12106) | (w5521 & w12106);
assign w2000 = w1756 & w8459;
assign w2001 = (w11261 & w14562) | (w11261 & w3059) | (w14562 & w3059);
assign w2002 = ~w14141 & w10159;
assign w2003 = ~w6798 & w12324;
assign w2004 = w3751 & ~w11117;
assign w2005 = w4559 & w13005;
assign w2006 = (~w3230 & w13654) | (~w3230 & w512) | (w13654 & w512);
assign w2007 = w2316 & w9009;
assign w2008 = ~w1979 & ~w13751;
assign w2009 = (w9805 & w10462) | (w9805 & w5801) | (w10462 & w5801);
assign w2010 = (w7757 & w10418) | (w7757 & w318) | (w10418 & w318);
assign w2011 = (w11500 & w13008) | (w11500 & w2440) | (w13008 & w2440);
assign w2012 = w2135 & w249;
assign w2013 = ~w11084 & ~w10222;
assign w2014 = w7244 & w6689;
assign w2015 = w2268 & ~w4992;
assign w2016 = w6845 & ~w7288;
assign w2017 = w4558 & w10480;
assign w2018 = ~w5230 & w5514;
assign w2019 = ~w12735 & w3599;
assign w2020 = ~w3175 & ~w8992;
assign w2021 = (w5901 & w14234) | (w5901 & w3080) | (w14234 & w3080);
assign w2022 = ~w10435 & w9469;
assign w2023 = w820 & w6804;
assign w2024 = (~w12955 & ~w13654) | (~w12955 & w13497) | (~w13654 & w13497);
assign w2025 = ~w9837 & w11724;
assign w2026 = ~w1650 & ~w1440;
assign w2027 = w7822 & ~w9378;
assign w2028 = w5102 & w4001;
assign w2029 = (~w12192 & w2144) | (~w12192 & w5336) | (w2144 & w5336);
assign w2030 = w3914 & ~w5673;
assign w2031 = ~w8448 & w4533;
assign w2032 = w11488 & w1712;
assign w2033 = w11031 & w10568;
assign w2034 = w13827 & w2698;
assign w2035 = ~w3942 & w7162;
assign w2036 = b110 & a110;
assign w2037 = w9004 & w12662;
assign w2038 = ~w3717 & ~w10880;
assign w2039 = w13526 & ~w7423;
assign w2040 = (~w5936 & w9564) | (~w5936 & w4444) | (w9564 & w4444);
assign w2041 = ~w8760 & w760;
assign w2042 = ~w2864 & w11606;
assign w2043 = (w12476 & w7581) | (w12476 & ~w12376) | (w7581 & ~w12376);
assign w2044 = ~w11176 & w13492;
assign w2045 = ~w10354 & w4458;
assign w2046 = w12982 & ~w7217;
assign w2047 = ~w8786 & w6201;
assign w2048 = (~w10272 & ~w4656) | (~w10272 & ~w7464) | (~w4656 & ~w7464);
assign w2049 = w9506 | ~w13008;
assign w2050 = w4221 & ~w7431;
assign w2051 = w12688 & ~w14392;
assign w2052 = w12621 & ~w2362;
assign w2053 = (w4723 & w836) | (w4723 & w2560) | (w836 & w2560);
assign w2054 = w5419 & ~w11454;
assign w2055 = w4836 & w2270;
assign w2056 = w1062 & ~w7075;
assign w2057 = w10545 & ~w11723;
assign w2058 = ~w1563 & w3508;
assign w2059 = w7721 & w23;
assign w2060 = ~w13942 & ~w6429;
assign w2061 = (w11661 & ~w1703) | (w11661 & w4737) | (~w1703 & w4737);
assign w2062 = (w4795 & w436) | (w4795 & ~w4799) | (w436 & ~w4799);
assign w2063 = ~w11246 & ~w2353;
assign w2064 = (w3023 & w1433) | (w3023 & w8750) | (w1433 & w8750);
assign w2065 = (w9646 & w845) | (w9646 & w2399) | (w845 & w2399);
assign w2066 = w3288 & ~w13323;
assign w2067 = ~w3444 & ~w8612;
assign w2068 = ~w5936 & w6433;
assign w2069 = w2583 & w5201;
assign w2070 = ~w13839 & ~w6436;
assign w2071 = (w12568 & w7021) | (w12568 & w6029) | (w7021 & w6029);
assign w2072 = ~w2848 & ~w11325;
assign w2073 = ~w7244 & ~w2701;
assign w2074 = ~w13011 & w9285;
assign w2075 = w10181 & w363;
assign w2076 = ~w1890 & ~w3370;
assign w2077 = ~w13249 & w2605;
assign w2078 = (w6310 & w12154) | (w6310 & ~w4754) | (w12154 & ~w4754);
assign w2079 = ~w5522 & w11861;
assign w2080 = (w2175 & w14322) | (w2175 & w9966) | (w14322 & w9966);
assign w2081 = ~b37 & ~a37;
assign w2082 = ~w4312 & ~w6219;
assign w2083 = w2753 & w11531;
assign w2084 = (~w10245 & w5881) | (~w10245 & w961) | (w5881 & w961);
assign w2085 = w167 & w6603;
assign w2086 = ~w11649 & ~w10601;
assign w2087 = ~w8367 & w2119;
assign w2088 = ~w4881 & w8785;
assign w2089 = ~w2486 & w3802;
assign w2090 = (~w5932 & w14051) | (~w5932 & ~w347) | (w14051 & ~w347);
assign w2091 = w13313 & w6757;
assign w2092 = w6291 & w11163;
assign w2093 = w7489 & w6445;
assign w2094 = (w3550 & w6455) | (w3550 & w13820) | (w6455 & w13820);
assign w2095 = w2228 & ~w3727;
assign w2096 = ~w10180 & w14569;
assign w2097 = w10439 & w12989;
assign w2098 = w7045 & w13041;
assign w2099 = w4647 & ~w3746;
assign w2100 = (~w1849 & w12190) | (~w1849 & w7118) | (w12190 & w7118);
assign w2101 = ~w10935 & w13730;
assign w2102 = w10036 & w8018;
assign w2103 = (~w14302 & w3817) | (~w14302 & w11620) | (w3817 & w11620);
assign w2104 = w13209 & w12139;
assign w2105 = (w7235 & w1613) | (w7235 & w12702) | (w1613 & w12702);
assign w2106 = (~w14395 & w13222) | (~w14395 & w5262) | (w13222 & w5262);
assign w2107 = w14087 & w4584;
assign w2108 = ~w10245 & w8917;
assign w2109 = (~w11261 & w1260) | (~w11261 & w6527) | (w1260 & w6527);
assign w2110 = w9004 & w11732;
assign w2111 = (~w2310 & w1084) | (~w2310 & w12971) | (w1084 & w12971);
assign w2112 = w697 & ~w6795;
assign w2113 = (~w13008 & w11261) | (~w13008 & w3940) | (w11261 & w3940);
assign w2114 = ~w8215 & w12043;
assign w2115 = w4100 & ~w959;
assign w2116 = (~w6975 & w8785) | (~w6975 & w10946) | (w8785 & w10946);
assign w2117 = ~w11745 & ~w646;
assign w2118 = w953 & w11538;
assign w2119 = w10605 & ~w3502;
assign w2120 = ~w8455 & w14578;
assign w2121 = ~w2946 & ~w13296;
assign w2122 = (~w5052 & w12951) | (~w5052 & w3862) | (w12951 & w3862);
assign w2123 = ~w450 & ~w5674;
assign w2124 = (~w7754 & w10350) | (~w7754 & w6994) | (w10350 & w6994);
assign w2125 = ~w3786 & w12173;
assign w2126 = ~w1419 & ~w12475;
assign w2127 = w10461 & w2629;
assign w2128 = w12102 & w12073;
assign w2129 = ~w11261 & w3294;
assign w2130 = w4700 & w3904;
assign w2131 = (~w12537 & w6079) | (~w12537 & w316) | (w6079 & w316);
assign w2132 = w9368 | w2849;
assign w2133 = w10676 & w5482;
assign w2134 = (w4127 & ~w12240) | (w4127 & w7877) | (~w12240 & w7877);
assign w2135 = ~w10704 & ~w803;
assign w2136 = ~w3209 & w4855;
assign w2137 = w5767 & w9265;
assign w2138 = (w10689 & w8766) | (w10689 & w7398) | (w8766 & w7398);
assign w2139 = w772 & ~w996;
assign w2140 = ~w1862 & ~w7455;
assign w2141 = (w11385 & w10307) | (w11385 & w11749) | (w10307 & w11749);
assign w2142 = w3435 & w3309;
assign w2143 = w13105 & ~w13585;
assign w2144 = w5468 & ~w5266;
assign w2145 = w11124 & w2492;
assign w2146 = w13172 & w10386;
assign w2147 = ~w235 & w7295;
assign w2148 = (w659 & w3505) | (w659 & w14002) | (w3505 & w14002);
assign w2149 = (~w14054 & w13227) | (~w14054 & w13307) | (w13227 & w13307);
assign w2150 = ~w12856 & w652;
assign w2151 = (w11708 & w3809) | (w11708 & ~w7853) | (w3809 & ~w7853);
assign w2152 = w11971 & ~w14060;
assign w2153 = ~w7415 & w11400;
assign w2154 = ~w11487 & w14070;
assign w2155 = ~w5480 & w3640;
assign w2156 = w3373 & w1243;
assign w2157 = w13830 & ~w9800;
assign w2158 = w7376 & w6542;
assign w2159 = b72 & a72;
assign w2160 = ~w3215 & ~w3717;
assign w2161 = ~w1828 & w10977;
assign w2162 = ~w10545 & ~w4515;
assign w2163 = ~w1142 & w8266;
assign w2164 = w9672 & w7645;
assign w2165 = ~w9545 & ~w5406;
assign w2166 = (~w4373 & w6367) | (~w4373 & w8593) | (w6367 & w8593);
assign w2167 = (w9364 & w6994) | (w9364 & w2445) | (w6994 & w2445);
assign w2168 = w6478 & ~w10380;
assign w2169 = (~w8659 & w8742) | (~w8659 & w4259) | (w8742 & w4259);
assign w2170 = ~w894 & w11708;
assign w2171 = w8584 & ~w2933;
assign w2172 = w8589 & ~w7348;
assign w2173 = ~w9852 & ~w10924;
assign w2174 = w8463 & ~w8651;
assign w2175 = w5675 & ~w13794;
assign w2176 = ~w3582 & ~w11546;
assign w2177 = w1285 & w11727;
assign w2178 = (w6617 & ~w12271) | (w6617 & w4627) | (~w12271 & w4627);
assign w2179 = w716 & ~w1351;
assign w2180 = (~w9688 & ~w14174) | (~w9688 & ~w9062) | (~w14174 & ~w9062);
assign w2181 = w11759 & w2;
assign w2182 = (w3144 & w2978) | (w3144 & ~w2576) | (w2978 & ~w2576);
assign w2183 = (w3776 & w13972) | (w3776 & w7990) | (w13972 & w7990);
assign w2184 = w13325 & w7716;
assign w2185 = w7806 & w910;
assign w2186 = w14178 & w5406;
assign w2187 = ~w11312 & w14336;
assign w2188 = (~w2060 & w1837) | (~w2060 & w26) | (w1837 & w26);
assign w2189 = b10 & a10;
assign w2190 = (w7085 & w2463) | (w7085 & w14608) | (w2463 & w14608);
assign w2191 = (~w5243 & w3146) | (~w5243 & ~w1583) | (w3146 & ~w1583);
assign w2192 = (~w6381 & w11429) | (~w6381 & w10848) | (w11429 & w10848);
assign w2193 = w10876 & ~w12292;
assign w2194 = ~w4764 & w14079;
assign w2195 = ~w8997 & w6127;
assign w2196 = w1798 & w3401;
assign w2197 = w12119 & w11186;
assign w2198 = (~w11487 & w3439) | (~w11487 & ~w9042) | (w3439 & ~w9042);
assign w2199 = ~w13306 & w9623;
assign w2200 = (~w11915 & w2874) | (~w11915 & w10405) | (w2874 & w10405);
assign w2201 = (~w3550 & w11875) | (~w3550 & w1357) | (w11875 & w1357);
assign w2202 = b42 & a42;
assign w2203 = ~w10514 & w4190;
assign w2204 = ~w770 & ~w14011;
assign w2205 = (~w10514 & w8234) | (~w10514 & w1825) | (w8234 & w1825);
assign w2206 = ~w8226 & w12134;
assign w2207 = ~w13583 & w6570;
assign w2208 = ~w10448 & ~w3622;
assign w2209 = w14396 & w3936;
assign w2210 = (~w7082 & w196) | (~w7082 & w6806) | (w196 & w6806);
assign w2211 = (w14194 & w9269) | (w14194 & w8165) | (w9269 & w8165);
assign w2212 = (w8916 & w13520) | (w8916 & w5450) | (w13520 & w5450);
assign w2213 = w6885 & ~w6500;
assign w2214 = w3550 & w8360;
assign w2215 = ~w10075 & ~w2599;
assign w2216 = (~w2317 & w13416) | (~w2317 & w538) | (w13416 & w538);
assign w2217 = (w5767 & ~w4171) | (w5767 & w1260) | (~w4171 & w1260);
assign w2218 = w5740 & ~w7279;
assign w2219 = w7592 | ~w2948;
assign w2220 = ~w4213 & w4359;
assign w2221 = (w8725 & w8548) | (w8725 & w6996) | (w8548 & w6996);
assign w2222 = w2433 & ~w6689;
assign w2223 = w3124 & ~w2701;
assign w2224 = (w12589 & w12897) | (w12589 & ~w6730) | (w12897 & ~w6730);
assign w2225 = (w8613 & w12161) | (w8613 & w2239) | (w12161 & w2239);
assign w2226 = (w11708 & ~w6992) | (w11708 & w8022) | (~w6992 & w8022);
assign w2227 = ~w11757 & ~w2228;
assign w2228 = ~b123 & ~a123;
assign w2229 = w5741 & w11117;
assign w2230 = w10225 & ~w10483;
assign w2231 = w13576 & w11276;
assign w2232 = w3447 & w12988;
assign w2233 = ~w7754 & w5224;
assign w2234 = (w3364 & w5877) | (w3364 & ~w5319) | (w5877 & ~w5319);
assign w2235 = ~w12642 & ~w9894;
assign w2236 = ~w2159 & w5767;
assign w2237 = (~w4420 & ~w1489) | (~w4420 & w9205) | (~w1489 & w9205);
assign w2238 = (w7567 & w12275) | (w7567 & ~w14534) | (w12275 & ~w14534);
assign w2239 = w1810 & w8613;
assign w2240 = (~w9138 & w9747) | (~w9138 & w10974) | (w9747 & w10974);
assign w2241 = w3289 & ~w2675;
assign w2242 = w3550 & w2702;
assign w2243 = ~w14659 & ~w6441;
assign w2244 = (w8389 & w12466) | (w8389 & w1600) | (w12466 & w1600);
assign w2245 = ~w8951 & w9398;
assign w2246 = (w13872 & w10847) | (w13872 & ~w2362) | (w10847 & ~w2362);
assign w2247 = w2698 & w4473;
assign w2248 = w7213 & w6885;
assign w2249 = (w2492 & w11124) | (w2492 & w5073) | (w11124 & w5073);
assign w2250 = ~w2175 & w12397;
assign w2251 = w813 & ~w10675;
assign w2252 = (w14146 & w13317) | (w14146 & w5038) | (w13317 & w5038);
assign w2253 = (~w10123 & w7748) | (~w10123 & w11625) | (w7748 & w11625);
assign w2254 = ~w9673 & w6657;
assign w2255 = (w2354 & w14371) | (w2354 & w6310) | (w14371 & w6310);
assign w2256 = w8574 & ~w4459;
assign w2257 = ~w2029 & w14292;
assign w2258 = ~w254 & w10076;
assign w2259 = ~w14302 & w3215;
assign w2260 = (~w4162 & w1612) | (~w4162 & ~w12376) | (w1612 & ~w12376);
assign w2261 = ~w3759 & ~w12685;
assign w2262 = (w1235 & w2358) | (w1235 & w9155) | (w2358 & w9155);
assign w2263 = (~w302 & w11709) | (~w302 & w12565) | (w11709 & w12565);
assign w2264 = (w9952 & ~w8790) | (w9952 & w5158) | (~w8790 & w5158);
assign w2265 = w2656 & w11417;
assign w2266 = w14033 & ~w3268;
assign w2267 = (~w268 & w11227) | (~w268 & w3648) | (w11227 & w3648);
assign w2268 = ~w11934 & w9716;
assign w2269 = (w8399 & ~w4545) | (w8399 & ~w2287) | (~w4545 & ~w2287);
assign w2270 = ~w3098 & ~w2320;
assign w2271 = ~w265 & w5676;
assign w2272 = ~w4483 & ~w8096;
assign w2273 = ~w4808 & ~w8867;
assign w2274 = ~w9586 & ~w10932;
assign w2275 = ~w5818 & w14308;
assign w2276 = ~w3341 & w5749;
assign w2277 = (~w2317 & w5873) | (~w2317 & w4226) | (w5873 & w4226);
assign w2278 = (w4538 & w12531) | (w4538 & w2587) | (w12531 & w2587);
assign w2279 = ~w12240 & w4299;
assign w2280 = (w12138 & w10384) | (w12138 & ~w10023) | (w10384 & ~w10023);
assign w2281 = w7052 & w8530;
assign w2282 = w4866 & w689;
assign w2283 = (w347 & ~w12295) | (w347 & w12963) | (~w12295 & w12963);
assign w2284 = w12575 & w12135;
assign w2285 = ~w8285 & ~w4028;
assign w2286 = w12485 & ~w2815;
assign w2287 = (~w50 & w9324) | (~w50 & w3145) | (w9324 & w3145);
assign w2288 = ~w12170 & ~w2135;
assign w2289 = ~w10219 & ~w3254;
assign w2290 = ~w10534 & w1633;
assign w2291 = b70 & a70;
assign w2292 = (w11861 & w432) | (w11861 & w7422) | (w432 & w7422);
assign w2293 = (w12460 & w13587) | (w12460 & w14572) | (w13587 & w14572);
assign w2294 = w12334 & ~w11608;
assign w2295 = w4270 & ~w10699;
assign w2296 = w3128 & w6829;
assign w2297 = ~w4756 & ~w3242;
assign w2298 = (w5662 & w13532) | (w5662 & w7002) | (w13532 & w7002);
assign w2299 = (w6586 & ~w11780) | (w6586 & w7098) | (~w11780 & w7098);
assign w2300 = ~w707 & w14537;
assign w2301 = w6746 & ~w5973;
assign w2302 = ~w2889 & w14161;
assign w2303 = (w8937 & w6401) | (w8937 & w2198) | (w6401 & w2198);
assign w2304 = w14306 & w5374;
assign w2305 = (~w4071 & ~w11586) | (~w4071 & w3583) | (~w11586 & w3583);
assign w2306 = ~w7633 & w9623;
assign w2307 = w11441 & ~w4517;
assign w2308 = (w5952 & w8303) | (w5952 & w5474) | (w8303 & w5474);
assign w2309 = ~w2203 & ~w6435;
assign w2310 = (w378 & w3721) | (w378 & w2181) | (w3721 & w2181);
assign w2311 = (~w8992 & w7082) | (~w8992 & w12311) | (w7082 & w12311);
assign w2312 = ~w8683 & w6857;
assign w2313 = (w6113 & w10197) | (w6113 & w12150) | (w10197 & w12150);
assign w2314 = w499 & ~w10075;
assign w2315 = (~w10590 & w7488) | (~w10590 & w12383) | (w7488 & w12383);
assign w2316 = (~w1362 & w3472) | (~w1362 & w4532) | (w3472 & w4532);
assign w2317 = ~w1321 & w14238;
assign w2318 = ~w12856 & ~w1552;
assign w2319 = ~w7132 & w10957;
assign w2320 = b54 & a54;
assign w2321 = w258 & ~w5728;
assign w2322 = (~w3963 & w11940) | (~w3963 & w1659) | (w11940 & w1659);
assign w2323 = ~w803 & w13620;
assign w2324 = w6989 & w13105;
assign w2325 = w2369 & w152;
assign w2326 = (~w14340 & w596) | (~w14340 & ~w6010) | (w596 & ~w6010);
assign w2327 = (~w2655 & w10167) | (~w2655 & w3014) | (w10167 & w3014);
assign w2328 = (~w5161 & w31) | (~w5161 & w2140) | (w31 & w2140);
assign w2329 = (w2655 & w6957) | (w2655 & w12863) | (w6957 & w12863);
assign w2330 = w9503 & w7272;
assign w2331 = w13590 & w3492;
assign w2332 = b73 & a73;
assign w2333 = ~w14504 & w3826;
assign w2334 = ~w4993 & ~w1854;
assign w2335 = ~w12958 & ~w5002;
assign w2336 = w4751 & ~w9219;
assign w2337 = ~w12255 & w12558;
assign w2338 = w183 & w5225;
assign w2339 = ~w2013 & ~w13123;
assign w2340 = w1840 & ~w4303;
assign w2341 = w3334 & w10068;
assign w2342 = w7167 & w2700;
assign w2343 = (w6207 & w5668) | (w6207 & ~w9096) | (w5668 & ~w9096);
assign w2344 = ~w14227 & ~w13694;
assign w2345 = ~w3157 & w6500;
assign w2346 = ~w14094 & w13552;
assign w2347 = w5294 & ~w2422;
assign w2348 = (w9304 & w1256) | (w9304 & w2836) | (w1256 & w2836);
assign w2349 = w9694 & ~w6716;
assign w2350 = (~w2680 & w4032) | (~w2680 & w5243) | (w4032 & w5243);
assign w2351 = cin & w9546;
assign w2352 = ~w10334 & ~w8302;
assign w2353 = ~w8328 & ~w11817;
assign w2354 = w1895 & ~w14324;
assign w2355 = ~w10949 & ~w11871;
assign w2356 = ~w2949 & ~w9580;
assign w2357 = w8253 & w11861;
assign w2358 = (w11429 & w1994) | (w11429 & w7396) | (w1994 & w7396);
assign w2359 = w2873 & ~w1252;
assign w2360 = w8769 & ~w6384;
assign w2361 = ~w5709 & w11453;
assign w2362 = ~w4982 & ~w5014;
assign w2363 = ~w13915 & w5854;
assign w2364 = (w6722 & w11834) | (w6722 & w12551) | (w11834 & w12551);
assign w2365 = (~w13802 & ~w9541) | (~w13802 & w5519) | (~w9541 & w5519);
assign w2366 = ~w14125 & w13684;
assign w2367 = (~w7012 & w13918) | (~w7012 & w2416) | (w13918 & w2416);
assign w2368 = w3963 & ~w11013;
assign w2369 = ~b10 & ~a10;
assign w2370 = w5593 & w13946;
assign w2371 = (~w11294 & ~w14414) | (~w11294 & w13773) | (~w14414 & w13773);
assign w2372 = ~w10761 & ~w10518;
assign w2373 = ~w13713 & w11037;
assign w2374 = ~w852 & w9227;
assign w2375 = w3047 & w8981;
assign w2376 = ~w3790 & ~w10669;
assign w2377 = w13197 & ~w5760;
assign w2378 = (w2717 & w6560) | (w2717 & ~w1563) | (w6560 & ~w1563);
assign w2379 = w10769 & ~w8824;
assign w2380 = ~w5619 & w12578;
assign w2381 = w13620 & ~w3098;
assign w2382 = (~w11936 & w3707) | (~w11936 & w11777) | (w3707 & w11777);
assign w2383 = w11458 & w7343;
assign w2384 = (~w11429 & w11716) | (~w11429 & w4690) | (w11716 & w4690);
assign w2385 = ~w3885 & w13306;
assign w2386 = w2076 & w10885;
assign w2387 = ~b90 & ~a90;
assign w2388 = w8871 & w12642;
assign w2389 = (~w10123 & w44) | (~w10123 & w5614) | (w44 & w5614);
assign w2390 = w13867 & ~w6381;
assign w2391 = w5177 & b93;
assign w2392 = (w6802 & w2404) | (w6802 & w355) | (w2404 & w355);
assign w2393 = w2872 & w3734;
assign w2394 = ~w3067 & ~w13607;
assign w2395 = ~w607 & w9788;
assign w2396 = (w869 & w8714) | (w869 & ~w9034) | (w8714 & ~w9034);
assign w2397 = w2433 & ~w7670;
assign w2398 = ~w4033 & ~w7013;
assign w2399 = w1152 & w9646;
assign w2400 = ~w1840 & ~w3024;
assign w2401 = ~w10941 & w9679;
assign w2402 = (~w7654 & ~w3846) | (~w7654 & ~w5662) | (~w3846 & ~w5662);
assign w2403 = w8905 & w1934;
assign w2404 = (w10808 & w5487) | (w10808 & w10984) | (w5487 & w10984);
assign w2405 = (w13860 & ~w10500) | (w13860 & w14458) | (~w10500 & w14458);
assign w2406 = w852 & ~w77;
assign w2407 = w8183 & w4458;
assign w2408 = ~w10676 & w8827;
assign w2409 = ~w8543 & ~w9661;
assign w2410 = ~b75 & ~a75;
assign w2411 = w13404 | ~w6266;
assign w2412 = (w12091 & w12308) | (w12091 & w12214) | (w12308 & w12214);
assign w2413 = (w2544 & ~w7342) | (w2544 & w7092) | (~w7342 & w7092);
assign w2414 = w7498 & ~w7077;
assign w2415 = ~w13011 & w4338;
assign w2416 = (~w5845 & w1258) | (~w5845 & w7011) | (w1258 & w7011);
assign w2417 = w7193 & w7628;
assign w2418 = ~w13636 & ~w9963;
assign w2419 = (w13924 & w5479) | (w13924 & w7975) | (w5479 & w7975);
assign w2420 = (w4363 & w5048) | (w4363 & w5361) | (w5048 & w5361);
assign w2421 = w12237 & ~w290;
assign w2422 = w5036 & w3958;
assign w2423 = w2656 & w4299;
assign w2424 = w3576 & w5746;
assign w2425 = ~w12958 & ~w813;
assign w2426 = ~w6451 & ~w8540;
assign w2427 = ~w71 & w11627;
assign w2428 = (~w14072 & w11635) | (~w14072 & w8371) | (w11635 & w8371);
assign w2429 = w5177 & w2569;
assign w2430 = ~w1563 & ~w6632;
assign w2431 = ~w4213 & w9871;
assign w2432 = w4286 & w12788;
assign w2433 = b113 & a113;
assign w2434 = w1472 & ~w12744;
assign w2435 = w9032 & ~w12061;
assign w2436 = w6104 & w9054;
assign w2437 = (~w1712 & w10764) | (~w1712 & w11953) | (w10764 & w11953);
assign w2438 = w351 & ~w10835;
assign w2439 = ~w14526 & ~w8171;
assign w2440 = b93 & w11500;
assign w2441 = w14347 | w13834;
assign w2442 = (w9156 & ~w9452) | (w9156 & w4849) | (~w9452 & w4849);
assign w2443 = w2428 & w3435;
assign w2444 = w9946 & ~w12560;
assign w2445 = w21 & ~w5498;
assign w2446 = w9495 & w7455;
assign w2447 = (w3734 & w10265) | (w3734 & ~w8791) | (w10265 & ~w8791);
assign w2448 = ~w7335 & ~w3251;
assign w2449 = (~w142 & ~w8459) | (~w142 & w6872) | (~w8459 & w6872);
assign w2450 = ~w3288 & w3162;
assign w2451 = ~w6696 & w141;
assign w2452 = w6045 & ~w9898;
assign w2453 = (~w5556 & w13222) | (~w5556 & w14395) | (w13222 & w14395);
assign w2454 = w4845 & w11117;
assign w2455 = (~w888 & ~w11481) | (~w888 & w12718) | (~w11481 & w12718);
assign w2456 = ~w1935 & w13655;
assign w2457 = (w217 & ~w11138) | (w217 & w7696) | (~w11138 & w7696);
assign w2458 = ~w1524 & ~w9220;
assign w2459 = ~w5294 & w8390;
assign w2460 = ~w7625 & w4975;
assign w2461 = (w13357 & w2115) | (w13357 & w2908) | (w2115 & w2908);
assign w2462 = ~w12271 & ~w2123;
assign w2463 = w167 & ~w1145;
assign w2464 = w4105 & w1283;
assign w2465 = ~w1712 & w5904;
assign w2466 = ~w11005 & ~w6856;
assign w2467 = ~w5522 & w7794;
assign w2468 = ~w5867 & w12039;
assign w2469 = ~w14629 & ~w12378;
assign w2470 = ~w4299 & ~w10590;
assign w2471 = ~w3914 & w12398;
assign w2472 = ~w1062 & w8713;
assign w2473 = w1790 & ~w6410;
assign w2474 = ~w5219 & w4997;
assign w2475 = (~w14300 & w8433) | (~w14300 & w12977) | (w8433 & w12977);
assign w2476 = ~w533 & ~w8768;
assign w2477 = ~w13733 & ~w3611;
assign w2478 = w6938 & w12114;
assign w2479 = w12709 & ~w1999;
assign w2480 = (~w4184 & w10529) | (~w4184 & w14143) | (w10529 & w14143);
assign w2481 = w8459 & ~w2941;
assign w2482 = ~w14302 & ~w6795;
assign w2483 = ~w6750 & w9672;
assign w2484 = w229 & w1481;
assign w2485 = w5422 & w10618;
assign w2486 = w3767 & w8516;
assign w2487 = (w8964 & w1848) | (w8964 & ~w536) | (w1848 & ~w536);
assign w2488 = (~w11013 & ~w4361) | (~w11013 & w6145) | (~w4361 & w6145);
assign w2489 = ~w4032 & ~w7762;
assign w2490 = ~w6935 & w2314;
assign w2491 = (~w13253 & ~w11439) | (~w13253 & ~w1416) | (~w11439 & ~w1416);
assign w2492 = ~w2121 & ~w7878;
assign w2493 = (~w9244 & w9338) | (~w9244 & w1466) | (w9338 & w1466);
assign w2494 = (~w2065 & w11647) | (~w2065 & w2842) | (w11647 & w2842);
assign w2495 = ~w1107 & ~w1468;
assign w2496 = w14053 & ~w1049;
assign w2497 = ~w6526 & ~w1035;
assign w2498 = ~w4099 & w9017;
assign w2499 = w9428 & w10419;
assign w2500 = ~w1151 & ~w6085;
assign w2501 = ~w10757 & ~w8475;
assign w2502 = (~w9853 & w4924) | (~w9853 & ~w11933) | (w4924 & ~w11933);
assign w2503 = ~w5098 & ~w2291;
assign w2504 = w9940 & w9378;
assign w2505 = (~w13107 & ~w10123) | (~w13107 & w1304) | (~w10123 & w1304);
assign w2506 = w9484 & w2635;
assign w2507 = (~w2655 & w6197) | (~w2655 & w10911) | (w6197 & w10911);
assign w2508 = ~w9871 & ~w6889;
assign w2509 = ~b115 & ~a115;
assign w2510 = (~w14343 & w12984) | (~w14343 & w415) | (w12984 & w415);
assign w2511 = ~w3734 & ~w12776;
assign w2512 = (~w2167 & w1018) | (~w2167 & w10759) | (w1018 & w10759);
assign w2513 = ~w13668 & w9032;
assign w2514 = w3611 & ~w12614;
assign w2515 = w6936 & ~w4931;
assign w2516 = (~w12286 & w381) | (~w12286 & w3455) | (w381 & w3455);
assign w2517 = w12609 & ~w9832;
assign w2518 = (w3435 & w13587) | (w3435 & w1278) | (w13587 & w1278);
assign w2519 = w7621 & w6626;
assign w2520 = (w3626 & w5698) | (w3626 & w1416) | (w5698 & w1416);
assign w2521 = ~w6378 & ~w9660;
assign w2522 = (~w3633 & ~w8181) | (~w3633 & w12389) | (~w8181 & w12389);
assign w2523 = ~w12112 & ~w5845;
assign w2524 = ~w14667 & ~w6460;
assign w2525 = (~w5569 & w13595) | (~w5569 & w9749) | (w13595 & w9749);
assign w2526 = w3065 & w1690;
assign w2527 = ~w10013 & ~w8280;
assign w2528 = (~w11756 & w6754) | (~w11756 & w7039) | (w6754 & w7039);
assign w2529 = w11481 & ~w8364;
assign w2530 = ~w7542 & w7914;
assign w2531 = ~w8955 & ~w5006;
assign w2532 = (w4239 & w7440) | (w4239 & w2457) | (w7440 & w2457);
assign w2533 = w10663 & w11594;
assign w2534 = (w9467 & w3783) | (w9467 & w2670) | (w3783 & w2670);
assign w2535 = (w5070 & w13157) | (w5070 & w12274) | (w13157 & w12274);
assign w2536 = ~w4134 & ~w4078;
assign w2537 = w13073 & w4989;
assign w2538 = ~w14064 & w3199;
assign w2539 = ~w3038 & w7968;
assign w2540 = (w14254 & w4149) | (w14254 & w236) | (w4149 & w236);
assign w2541 = (w14028 & ~w11481) | (w14028 & w2494) | (~w11481 & w2494);
assign w2542 = (w4193 & ~w8790) | (w4193 & w11792) | (~w8790 & w11792);
assign w2543 = w3914 & w218;
assign w2544 = ~w2425 & ~w2710;
assign w2545 = w5294 & ~w3958;
assign w2546 = (w5662 & w6354) | (w5662 & w7102) | (w6354 & w7102);
assign w2547 = w4798 & ~w1445;
assign w2548 = ~w4464 & w1470;
assign w2549 = ~w8213 & ~w4585;
assign w2550 = ~w2500 & w3508;
assign w2551 = w12569 & ~w5571;
assign w2552 = (w13685 & w11230) | (w13685 & w12894) | (w11230 & w12894);
assign w2553 = w3751 & ~w2941;
assign w2554 = w13937 & w3885;
assign w2555 = ~w3209 & w10516;
assign w2556 = ~w71 & w3311;
assign w2557 = ~w5842 & w13982;
assign w2558 = (w10997 & w12499) | (w10997 & w11485) | (w12499 & w11485);
assign w2559 = w2261 & ~w10339;
assign w2560 = ~w7630 & w2569;
assign w2561 = ~w11395 & ~w3502;
assign w2562 = (w2343 & w12610) | (w2343 & w8228) | (w12610 & w8228);
assign w2563 = ~w6750 & w6421;
assign w2564 = w1760 & w10036;
assign w2565 = (w227 & w614) | (w227 & w10821) | (w614 & w10821);
assign w2566 = ~w7001 & ~w6689;
assign w2567 = w10119 & w2858;
assign w2568 = w10368 | ~w14390;
assign w2569 = ~w7365 & ~w3321;
assign w2570 = w607 & ~w13937;
assign w2571 = (w2144 & w12837) | (w2144 & w3881) | (w12837 & w3881);
assign w2572 = ~w5660 & ~w5178;
assign w2573 = ~w4787 & w9541;
assign w2574 = ~w12121 & ~w2850;
assign w2575 = w6041 & w6886;
assign w2576 = (w3017 & w3137) | (w3017 & w14481) | (w3137 & w14481);
assign w2577 = ~w3790 & w10997;
assign w2578 = ~w1972 & ~w2206;
assign w2579 = w3153 & ~w3412;
assign w2580 = w12253 & w7559;
assign w2581 = w4525 & w13283;
assign w2582 = w12632 & ~w8381;
assign w2583 = ~w4508 & w11219;
assign w2584 = ~w12148 & ~w2272;
assign w2585 = w3215 & w6230;
assign w2586 = ~w13737 & w6574;
assign w2587 = w1061 & w4256;
assign w2588 = w3540 & ~w13271;
assign w2589 = ~w2032 & ~w6906;
assign w2590 = ~w7645 & w6206;
assign w2591 = (~w9672 & ~w9898) | (~w9672 & w6889) | (~w9898 & w6889);
assign w2592 = ~w6651 & w3337;
assign w2593 = w5140 | ~w3289;
assign w2594 = w1581 & ~w5907;
assign w2595 = (~w9403 & w8282) | (~w9403 & w12154) | (w8282 & w12154);
assign w2596 = w2749 & w6722;
assign w2597 = ~w1840 & ~w11068;
assign w2598 = (w2289 & ~w4867) | (w2289 & w10871) | (~w4867 & w10871);
assign w2599 = ~w10075 & ~w884;
assign w2600 = w5794 & ~w10213;
assign w2601 = w12918 & w7130;
assign w2602 = w11330 & ~w7557;
assign w2603 = w9465 & w9183;
assign w2604 = w8390 & w4796;
assign w2605 = ~w4881 & ~w2202;
assign w2606 = w10378 & ~w10377;
assign w2607 = w6044 & ~w7815;
assign w2608 = ~w408 & w3168;
assign w2609 = (w11803 & w3998) | (w11803 & w13912) | (w3998 & w13912);
assign w2610 = w11068 & w3767;
assign w2611 = ~w4122 & w8214;
assign w2612 = (~w8130 & w11867) | (~w8130 & w8771) | (w11867 & w8771);
assign w2613 = w3007 & ~w12120;
assign w2614 = w153 & w10217;
assign w2615 = (w6802 & w11156) | (w6802 & w1863) | (w11156 & w1863);
assign w2616 = (w4511 & w1181) | (w4511 & w9600) | (w1181 & w9600);
assign w2617 = ~w4071 & ~w3361;
assign w2618 = w11364 & ~w443;
assign w2619 = ~w5559 & w8757;
assign w2620 = ~w7756 & w8550;
assign w2621 = w12879 & w5360;
assign w2622 = ~w7859 & ~w6744;
assign w2623 = w8626 & ~w884;
assign w2624 = ~w1542 & w4210;
assign w2625 = (w11902 & w13462) | (w11902 & w1066) | (w13462 & w1066);
assign w2626 = ~w6538 & w5156;
assign w2627 = w9482 & w12642;
assign w2628 = (w14121 & w5466) | (w14121 & w3955) | (w5466 & w3955);
assign w2629 = ~w2877 & ~w994;
assign w2630 = ~w917 & ~w11706;
assign w2631 = w10699 & w13837;
assign w2632 = (w11708 & ~w1840) | (w11708 & w8331) | (~w1840 & w8331);
assign w2633 = w6562 & w10353;
assign w2634 = w480 & ~w8065;
assign w2635 = w12934 & w13776;
assign w2636 = (w8584 & w4512) | (w8584 & w5181) | (w4512 & w5181);
assign w2637 = ~w1322 & w4523;
assign w2638 = ~w12879 & w12656;
assign w2639 = w9713 & w8769;
assign w2640 = (w10317 & w2175) | (w10317 & w11653) | (w2175 & w11653);
assign w2641 = ~w12716 & w7662;
assign w2642 = w7794 & w6000;
assign w2643 = (w6542 & w12003) | (w6542 & w6870) | (w12003 & w6870);
assign w2644 = w10853 & ~w3044;
assign w2645 = w552 & w12127;
assign w2646 = (w6952 & w4658) | (w6952 & w5722) | (w4658 & w5722);
assign w2647 = w12615 & ~w14564;
assign w2648 = ~w3761 & w13776;
assign w2649 = (~w10234 & w12555) | (~w10234 & w3618) | (w12555 & w3618);
assign w2650 = (w12482 & w9614) | (w12482 & w431) | (w9614 & w431);
assign w2651 = w12195 & w11883;
assign w2652 = ~w6366 & w2119;
assign w2653 = (~w142 & ~w9296) | (~w142 & w6872) | (~w9296 & w6872);
assign w2654 = w2701 & w8045;
assign w2655 = (~w6426 & w13454) | (~w6426 & w13889) | (w13454 & w13889);
assign w2656 = ~w8662 & ~w11941;
assign w2657 = w2129 & ~w1665;
assign w2658 = w142 & ~w3904;
assign w2659 = (w8623 & w11826) | (w8623 & w6060) | (w11826 & w6060);
assign w2660 = ~w9012 & w2960;
assign w2661 = ~w1840 & w13713;
assign w2662 = w2024 & ~w2006;
assign w2663 = ~w2332 & ~w2508;
assign w2664 = ~w11745 & ~w13323;
assign w2665 = (w3727 & w6324) | (w3727 & w840) | (w6324 & w840);
assign w2666 = w3373 & ~w9403;
assign w2667 = w11779 & ~w4565;
assign w2668 = (~w8436 & w14211) | (~w8436 & w4476) | (w14211 & w4476);
assign w2669 = w334 & w9555;
assign w2670 = (w6802 & w13871) | (w6802 & w4342) | (w13871 & w4342);
assign w2671 = w11236 & w4142;
assign w2672 = (w3039 & ~w985) | (w3039 & w11341) | (~w985 & w11341);
assign w2673 = w10165 & w5319;
assign w2674 = ~w7744 & ~w12296;
assign w2675 = b48 & a48;
assign w2676 = ~w6461 & ~w11484;
assign w2677 = ~w14553 & ~w2822;
assign w2678 = ~w12355 & w6971;
assign w2679 = w3914 & ~w12060;
assign w2680 = b79 & a79;
assign w2681 = w12271 & w8205;
assign w2682 = ~w5778 & w13839;
assign w2683 = (~w3333 & w12855) | (~w3333 & w266) | (w12855 & w266);
assign w2684 = ~w1811 & ~w14155;
assign w2685 = w8988 & w11820;
assign w2686 = ~w5644 & w8028;
assign w2687 = ~w5294 & w7772;
assign w2688 = w10331 & w4666;
assign w2689 = w12458 & ~w8015;
assign w2690 = ~w4989 & w8147;
assign w2691 = (~w2270 & ~w14542) | (~w2270 & ~w4339) | (~w14542 & ~w4339);
assign w2692 = w6929 & ~w5694;
assign w2693 = (w5952 & w13696) | (w5952 & w1576) | (w13696 & w1576);
assign w2694 = (w1705 & w14196) | (w1705 & w2487) | (w14196 & w2487);
assign w2695 = ~w13122 & w5645;
assign w2696 = ~w11492 & ~w3916;
assign w2697 = ~w3962 & w13752;
assign w2698 = w2599 & w9032;
assign w2699 = w6279 & w27;
assign w2700 = (w13924 & ~w8769) | (w13924 & w576) | (~w8769 & w576);
assign w2701 = ~w8782 & ~w896;
assign w2702 = ~w3790 & w7772;
assign w2703 = ~w7312 & w5575;
assign w2704 = (w8513 & w387) | (w8513 & w10537) | (w387 & w10537);
assign w2705 = w6391 & w10728;
assign w2706 = (w2181 & w14284) | (w2181 & w7509) | (w14284 & w7509);
assign w2707 = ~w2036 & ~w14614;
assign w2708 = w3124 & w394;
assign w2709 = (w12138 & w7579) | (w12138 & w3249) | (w7579 & w3249);
assign w2710 = w10675 & w9838;
assign w2711 = ~w4820 & w14459;
assign w2712 = ~w13194 & w5064;
assign w2713 = (~w9614 & w1310) | (~w9614 & w9721) | (w1310 & w9721);
assign w2714 = w11708 & ~w8953;
assign w2715 = w9226 & w9748;
assign w2716 = (w13870 & w9556) | (w13870 & w6263) | (w9556 & w6263);
assign w2717 = w2137 & w14486;
assign w2718 = w6521 & w7751;
assign w2719 = ~w10675 & ~w12589;
assign w2720 = ~w14011 & w7782;
assign w2721 = (w339 & w10521) | (w339 & ~w13409) | (w10521 & ~w13409);
assign w2722 = ~w12460 & w7660;
assign w2723 = ~w7120 & w7728;
assign w2724 = ~w2464 & ~w8809;
assign w2725 = ~w569 & w531;
assign w2726 = w2656 & w2425;
assign w2727 = w10346 & w14652;
assign w2728 = w2913 & w9385;
assign w2729 = ~w12809 & ~w14588;
assign w2730 = ~w13297 & ~w5937;
assign w2731 = ~w12240 & w10075;
assign w2732 = ~w12306 & ~w691;
assign w2733 = (~w5482 & w13749) | (~w5482 & ~w112) | (w13749 & ~w112);
assign w2734 = w7875 & ~w9294;
assign w2735 = ~w12146 & ~w2991;
assign w2736 = ~w2317 & w4640;
assign w2737 = ~w7845 & w12244;
assign w2738 = (~w6802 & w6160) | (~w6802 & w3009) | (w6160 & w3009);
assign w2739 = w646 & w2501;
assign w2740 = w9839 & w1260;
assign w2741 = ~w10689 & ~w3885;
assign w2742 = ~w5559 & w7964;
assign w2743 = (w9093 & w13074) | (w9093 & w2016) | (w13074 & w2016);
assign w2744 = (w7914 & w9012) | (w7914 & w7825) | (w9012 & w7825);
assign w2745 = ~w6620 & ~w9444;
assign w2746 = ~w4312 & w12112;
assign w2747 = (~w11429 & w10745) | (~w11429 & w5445) | (w10745 & w5445);
assign w2748 = w10889 & w6610;
assign w2749 = w13919 & w10888;
assign w2750 = ~w6697 & w3039;
assign w2751 = b30 & a30;
assign w2752 = w9284 & w5912;
assign w2753 = ~w6034 & ~w10870;
assign w2754 = ~w1730 & w11993;
assign w2755 = w9788 & ~w2701;
assign w2756 = (~w3885 & ~w325) | (~w3885 & w3563) | (~w325 & w3563);
assign w2757 = ~w12023 & ~w9194;
assign w2758 = ~w260 & ~w12642;
assign w2759 = ~w13426 & ~w11031;
assign w2760 = ~w11003 & ~w11303;
assign w2761 = w183 & ~w7662;
assign w2762 = b22 & a22;
assign w2763 = w14650 | w13311;
assign w2764 = w3288 & ~w5761;
assign w2765 = (w9032 & w4473) | (w9032 & w6927) | (w4473 & w6927);
assign w2766 = ~w2218 & w384;
assign w2767 = w13013 & ~w11109;
assign w2768 = (w7567 & w12275) | (w7567 & ~w5662) | (w12275 & ~w5662);
assign w2769 = (w7612 & w1771) | (w7612 & w3494) | (w1771 & w3494);
assign w2770 = (w9702 & w6630) | (w9702 & ~w4736) | (w6630 & ~w4736);
assign w2771 = ~w14410 & w5017;
assign w2772 = w9287 & w11427;
assign w2773 = ~w2762 & ~w13872;
assign w2774 = (~w11429 & w8498) | (~w11429 & w13602) | (w8498 & w13602);
assign w2775 = w6128 & ~w7022;
assign w2776 = w7376 & w13565;
assign w2777 = w11583 & ~w9724;
assign w2778 = (~w10435 & w521) | (~w10435 & w8933) | (w521 & w8933);
assign w2779 = ~w10077 & w14649;
assign w2780 = (~w13620 & w12206) | (~w13620 & ~w3564) | (w12206 & ~w3564);
assign w2781 = w6083 & ~w11028;
assign w2782 = ~w71 & w2429;
assign w2783 = ~w463 & ~w13125;
assign w2784 = ~w1609 & w6334;
assign w2785 = w14470 & ~w13902;
assign w2786 = (~w918 & w14424) | (~w918 & w1686) | (w14424 & w1686);
assign w2787 = ~w13349 & w10642;
assign w2788 = ~w217 & w7914;
assign w2789 = (w1264 & w11429) | (w1264 & w10743) | (w11429 & w10743);
assign w2790 = w14592 & ~w13674;
assign w2791 = ~w9861 & w8443;
assign w2792 = w2656 & w10853;
assign w2793 = (w79 & w6789) | (w79 & ~w237) | (w6789 & ~w237);
assign w2794 = (~w12875 & w10829) | (~w12875 & w3762) | (w10829 & w3762);
assign w2795 = ~w9118 & ~w4804;
assign w2796 = w2656 & ~w5532;
assign w2797 = (w11925 & w7565) | (w11925 & w14315) | (w7565 & w14315);
assign w2798 = ~w6237 & ~w12342;
assign w2799 = (w12473 & w4608) | (w12473 & w1230) | (w4608 & w1230);
assign w2800 = (w10551 & w8937) | (w10551 & w477) | (w8937 & w477);
assign w2801 = (~w2575 & w4512) | (~w2575 & w3445) | (w4512 & w3445);
assign w2802 = w13652 & w2701;
assign w2803 = (w12077 & ~w7616) | (w12077 & w8510) | (~w7616 & w8510);
assign w2804 = w3828 & w11411;
assign w2805 = w10136 | ~w4007;
assign w2806 = w5949 & w329;
assign w2807 = (w4103 & w5254) | (w4103 & w8064) | (w5254 & w8064);
assign w2808 = ~w1534 & ~w1022;
assign w2809 = ~w843 & w9782;
assign w2810 = (w14543 & w12345) | (w14543 & w3846) | (w12345 & w3846);
assign w2811 = w3435 & ~w12993;
assign w2812 = (w8437 & w1088) | (w8437 & w2581) | (w1088 & w2581);
assign w2813 = (w5574 & w8199) | (w5574 & w3028) | (w8199 & w3028);
assign w2814 = ~w9927 & w4458;
assign w2815 = w848 & w11821;
assign w2816 = ~w2824 & ~w1753;
assign w2817 = ~w2500 & w545;
assign w2818 = w14518 & ~w2857;
assign w2819 = w10807 & ~w3404;
assign w2820 = w4190 & w8018;
assign w2821 = (~w8018 & w5702) | (~w8018 & w11406) | (w5702 & w11406);
assign w2822 = ~w1308 & w1784;
assign w2823 = ~w6536 & w9139;
assign w2824 = ~w7630 & ~w11218;
assign w2825 = w8873 & ~w9655;
assign w2826 = w4213 & w4587;
assign w2827 = (~w2422 & w13349) | (~w2422 & w2347) | (w13349 & w2347);
assign w2828 = ~w13324 & w4326;
assign w2829 = w14640 & ~w6689;
assign w2830 = ~w4700 & w8396;
assign w2831 = w1646 & ~w12776;
assign w2832 = ~w4920 & ~w7700;
assign w2833 = ~w1524 & ~w5114;
assign w2834 = (w12125 & ~w9298) | (w12125 & ~w9794) | (~w9298 & ~w9794);
assign w2835 = w325 & w2385;
assign w2836 = ~w10441 & w8777;
assign w2837 = w4877 & ~w10762;
assign w2838 = w2237 & w9971;
assign w2839 = ~w142 & ~w6500;
assign w2840 = ~w607 & w12642;
assign w2841 = ~w2509 & w646;
assign w2842 = w14028 & ~w14372;
assign w2843 = w1838 & ~w2036;
assign w2844 = ~w1870 & ~w505;
assign w2845 = w2888 & ~w13359;
assign w2846 = ~w4836 & w8827;
assign w2847 = w3401 & ~w13258;
assign w2848 = (w2982 & w8699) | (w2982 & w252) | (w8699 & w252);
assign w2849 = ~w1380 & ~w9907;
assign w2850 = (~w1821 & w6763) | (~w1821 & w3614) | (w6763 & w3614);
assign w2851 = ~w10221 & ~w6689;
assign w2852 = w11171 & w6774;
assign w2853 = w11578 | w12460;
assign w2854 = (w12 & w7455) | (w12 & w3639) | (w7455 & w3639);
assign w2855 = w3661 & ~w10483;
assign w2856 = w4756 & w2600;
assign w2857 = w6562 & ~w11536;
assign w2858 = (~w6572 & w14417) | (~w6572 & w6359) | (w14417 & w6359);
assign w2859 = ~w142 & ~w2941;
assign w2860 = ~w1113 & ~w11612;
assign w2861 = ~w4479 & w6503;
assign w2862 = (w1166 & w1580) | (w1166 & w12236) | (w1580 & w12236);
assign w2863 = (w5127 & w3465) | (w5127 & w194) | (w3465 & w194);
assign w2864 = ~b43 & ~a43;
assign w2865 = ~w11997 & w6949;
assign w2866 = (w699 & w14596) | (w699 & w9053) | (w14596 & w9053);
assign w2867 = (w6949 & ~w11158) | (w6949 & w11958) | (~w11158 & w11958);
assign w2868 = w11755 & w4943;
assign w2869 = ~w1431 & ~w5105;
assign w2870 = (w14648 & w4101) | (w14648 & w11850) | (w4101 & w11850);
assign w2871 = w11899 & w12460;
assign w2872 = ~w11905 & ~w9465;
assign w2873 = ~w8158 & w11607;
assign w2874 = (w5794 & w4756) | (w5794 & w2600) | (w4756 & w2600);
assign w2875 = ~w3435 & ~w3044;
assign w2876 = w9917 & w11336;
assign w2877 = w6328 & ~w11375;
assign w2878 = (w13899 & w7860) | (w13899 & ~w12376) | (w7860 & ~w12376);
assign w2879 = (w6683 & w2262) | (w6683 & w4096) | (w2262 & w4096);
assign w2880 = (~w6381 & w13282) | (~w6381 & w8987) | (w13282 & w8987);
assign w2881 = w4997 & w14401;
assign w2882 = w10676 & w4627;
assign w2883 = w13451 & w4202;
assign w2884 = w8713 & w9921;
assign w2885 = (w13168 & w1072) | (w13168 & ~w9591) | (w1072 & ~w9591);
assign w2886 = (w12209 & w10294) | (w12209 & w12408) | (w10294 & w12408);
assign w2887 = (w309 & w4050) | (w309 & w13608) | (w4050 & w13608);
assign w2888 = ~w10774 & ~w6377;
assign w2889 = ~w164 & w14406;
assign w2890 = ~w6929 & w1658;
assign w2891 = ~w2159 & ~w45;
assign w2892 = w3734 & w13485;
assign w2893 = ~w13852 & ~w13001;
assign w2894 = (w3550 & w13711) | (w3550 & w13738) | (w13711 & w13738);
assign w2895 = ~w479 & ~w4542;
assign w2896 = w11340 & w10169;
assign w2897 = w11754 & w3314;
assign w2898 = (~w10618 & w11337) | (~w10618 & ~w1928) | (w11337 & ~w1928);
assign w2899 = w8005 & w4740;
assign w2900 = w9612 & ~w6362;
assign w2901 = ~w12028 & w3968;
assign w2902 = (w7644 & w7522) | (w7644 & w2240) | (w7522 & w2240);
assign w2903 = ~w6485 & w13434;
assign w2904 = (~w9541 & w1885) | (~w9541 & w7928) | (w1885 & w7928);
assign w2905 = ~w4473 & ~w10203;
assign w2906 = ~w5935 & ~w2053;
assign w2907 = (~w10435 & w11365) | (~w10435 & w8625) | (w11365 & w8625);
assign w2908 = ~w14217 & w13357;
assign w2909 = w5052 & w5422;
assign w2910 = w12531 & w5163;
assign w2911 = (~w10855 & w13324) | (~w10855 & w11935) | (w13324 & w11935);
assign w2912 = w13542 & ~w4886;
assign w2913 = ~w6072 & ~w3567;
assign w2914 = ~w5317 & ~w8929;
assign w2915 = ~w6032 & ~w4611;
assign w2916 = w10290 & w13629;
assign w2917 = w5294 & ~w6886;
assign w2918 = (~w4287 & w2971) | (~w4287 & ~w14074) | (w2971 & ~w14074);
assign w2919 = ~w4050 & w10623;
assign w2920 = w6224 & w9921;
assign w2921 = (~w11861 & w8511) | (~w11861 & w1384) | (w8511 & w1384);
assign w2922 = b91 & a91;
assign w2923 = ~w9046 & w10426;
assign w2924 = ~w6561 & ~w11452;
assign w2925 = (w853 & w12576) | (w853 & w5380) | (w12576 & w5380);
assign w2926 = (w3067 & w2049) | (w3067 & w10443) | (w2049 & w10443);
assign w2927 = w829 & ~w9748;
assign w2928 = ~w14291 & ~w9613;
assign w2929 = (w1036 & w2175) | (w1036 & w9677) | (w2175 & w9677);
assign w2930 = w9780 & w4855;
assign w2931 = (~w4099 & w3408) | (~w4099 & w8082) | (w3408 & w8082);
assign w2932 = ~w12982 & ~w2039;
assign w2933 = ~b87 & ~a87;
assign w2934 = ~w2808 & ~w11838;
assign w2935 = ~w8900 & ~w9449;
assign w2936 = ~w11909 & ~w1507;
assign w2937 = ~w3619 & ~w5800;
assign w2938 = ~w12943 & ~w1229;
assign w2939 = (~w1928 & w10688) | (~w1928 & w13331) | (w10688 & w13331);
assign w2940 = w2320 & ~w13854;
assign w2941 = ~w1802 & ~w3288;
assign w2942 = ~w1712 & w7009;
assign w2943 = ~w10204 & w8245;
assign w2944 = w5294 & ~w5002;
assign w2945 = ~w13687 & ~w6417;
assign w2946 = ~w3425 & w956;
assign w2947 = ~w7267 & w14031;
assign w2948 = ~w14664 & w2201;
assign w2949 = ~w10410 & w9541;
assign w2950 = w3852 & w6433;
assign w2951 = b33 & a33;
assign w2952 = ~w3906 & ~w13946;
assign w2953 = ~w3587 & ~w11437;
assign w2954 = ~w1465 & ~w6874;
assign w2955 = ~w11745 & ~w11117;
assign w2956 = ~w607 & ~w12460;
assign w2957 = w2656 & w2938;
assign w2958 = (w79 & w6789) | (w79 & ~w5530) | (w6789 & ~w5530);
assign w2959 = w11583 & ~w11037;
assign w2960 = ~w5867 & w12856;
assign w2961 = ~w12543 & w4711;
assign w2962 = ~w2159 & ~w2332;
assign w2963 = (w13379 & w7938) | (w13379 & w13291) | (w7938 & w13291);
assign w2964 = w1498 & ~w852;
assign w2965 = ~w641 & ~w2911;
assign w2966 = ~w468 & w1643;
assign w2967 = (w10664 & ~w4843) | (w10664 & w14655) | (~w4843 & w14655);
assign w2968 = w6421 & w4541;
assign w2969 = (~w14390 & w10368) | (~w14390 & ~w8589) | (w10368 & ~w8589);
assign w2970 = (w14646 & ~w4336) | (w14646 & w14413) | (~w4336 & w14413);
assign w2971 = (~w4287 & w7464) | (~w4287 & w9884) | (w7464 & w9884);
assign w2972 = (w13089 & w8289) | (w13089 & w7805) | (w8289 & w7805);
assign w2973 = ~w2380 & w3287;
assign w2974 = (~w2159 & w8893) | (~w2159 & w7080) | (w8893 & w7080);
assign w2975 = ~w9921 & w12826;
assign w2976 = (w2284 & w13152) | (w2284 & w11388) | (w13152 & w11388);
assign w2977 = (w12330 & w6803) | (w12330 & w6219) | (w6803 & w6219);
assign w2978 = ~w861 & w12141;
assign w2979 = ~w1699 & w7226;
assign w2980 = w7349 & ~w7185;
assign w2981 = ~w4637 & ~w1642;
assign w2982 = (~w10245 & w3069) | (~w10245 & w2435) | (w3069 & w2435);
assign w2983 = w1838 & ~w646;
assign w2984 = ~w11932 & w12573;
assign w2985 = ~w7228 & ~w12849;
assign w2986 = ~w2386 & w11500;
assign w2987 = (w4352 & ~w3264) | (w4352 & w9185) | (~w3264 & w9185);
assign w2988 = ~w3733 & ~w4464;
assign w2989 = w9672 & w14335;
assign w2990 = (w9734 & w8829) | (w9734 & w7514) | (w8829 & w7514);
assign w2991 = (~w9198 & w13363) | (~w9198 & w1775) | (w13363 & w1775);
assign w2992 = w4989 & ~w3785;
assign w2993 = ~w10519 | ~w5282;
assign w2994 = ~w12656 & ~w13114;
assign w2995 = (~w8843 & ~w1794) | (~w8843 & w5228) | (~w1794 & w5228);
assign w2996 = w13344 & ~w3727;
assign w2997 = w6556 & w4408;
assign w2998 = ~w13526 & ~w7080;
assign w2999 = (w14009 & w13493) | (w14009 & w10406) | (w13493 & w10406);
assign w3000 = (~w6266 & w9012) | (~w6266 & w10989) | (w9012 & w10989);
assign w3001 = w13734 & w13873;
assign w3002 = (w637 & ~w349) | (w637 & w3118) | (~w349 & w3118);
assign w3003 = (w534 & w4411) | (w534 & w3564) | (w4411 & w3564);
assign w3004 = (w14074 & w160) | (w14074 & w87) | (w160 & w87);
assign w3005 = ~w11057 & ~w5119;
assign w3006 = (w1359 & w4463) | (w1359 & w3939) | (w4463 & w3939);
assign w3007 = w10689 & w12569;
assign w3008 = ~w12807 & ~w9043;
assign w3009 = (w11472 & w10905) | (w11472 & w12537) | (w10905 & w12537);
assign w3010 = ~w1199 & w9541;
assign w3011 = w10045 & w13551;
assign w3012 = ~w3693 & ~w5782;
assign w3013 = ~w1840 & w12893;
assign w3014 = (w3442 & w897) | (w3442 & ~w996) | (w897 & ~w996);
assign w3015 = ~w4033 & w7132;
assign w3016 = w11680 & ~w833;
assign w3017 = (~w1802 & w10039) | (~w1802 & w7171) | (w10039 & w7171);
assign w3018 = w874 & ~w8603;
assign w3019 = b86 & a86;
assign w3020 = w3550 & ~w4780;
assign w3021 = (w13713 & w14289) | (w13713 & w12831) | (w14289 & w12831);
assign w3022 = ~w14302 & w3098;
assign w3023 = ~w12193 & w14260;
assign w3024 = (~w4359 & w7851) | (~w4359 & w11074) | (w7851 & w11074);
assign w3025 = b67 & a67;
assign w3026 = (w13219 & w10392) | (w13219 & w12035) | (w10392 & w12035);
assign w3027 = w9944 & ~w7590;
assign w3028 = ~w2492 & ~w11958;
assign w3029 = (~w11738 & ~w6432) | (~w11738 & w4673) | (~w6432 & w4673);
assign w3030 = (~w9107 & w10964) | (~w9107 & w1700) | (w10964 & w1700);
assign w3031 = ~w9918 & ~w6954;
assign w3032 = ~w7376 & ~w3508;
assign w3033 = w6287 & w5183;
assign w3034 = ~w14570 & ~w14361;
assign w3035 = ~w6553 & w7349;
assign w3036 = ~b91 & ~a91;
assign w3037 = ~w2454 & ~w12873;
assign w3038 = ~w12398 & ~w5732;
assign w3039 = w14660 & w3158;
assign w3040 = ~w4970 & w4851;
assign w3041 = w8396 & w1367;
assign w3042 = w11236 & w3181;
assign w3043 = w7470 & w4622;
assign w3044 = w3392 & ~w70;
assign w3045 = ~w5702 & w7778;
assign w3046 = ~w7426 & ~w6925;
assign w3047 = w2126 & w4705;
assign w3048 = ~w708 & ~w11042;
assign w3049 = ~w2947 & w10066;
assign w3050 = (w6306 & w7986) | (w6306 & w4025) | (w7986 & w4025);
assign w3051 = ~w12240 & w9433;
assign w3052 = (~w13135 & ~w1868) | (~w13135 & ~w1928) | (~w1868 & ~w1928);
assign w3053 = ~w2463 & w6878;
assign w3054 = w6651 & w13713;
assign w3055 = (w3289 & ~w5783) | (w3289 & w4415) | (~w5783 & w4415);
assign w3056 = ~w13077 & ~w3964;
assign w3057 = ~w10786 & w6428;
assign w3058 = w9389 & ~w11031;
assign w3059 = (~w4233 & w13651) | (~w4233 & w8234) | (w13651 & w8234);
assign w3060 = ~w3914 & w8390;
assign w3061 = w10676 & w1507;
assign w3062 = ~w3894 & ~w11004;
assign w3063 = ~w2100 & ~w5639;
assign w3064 = w5867 & ~w12338;
assign w3065 = w11357 & ~w3894;
assign w3066 = ~w5292 & ~w9697;
assign w3067 = (~w8196 & w4050) | (~w8196 & w12099) | (w4050 & w12099);
assign w3068 = (~w6929 & w8636) | (~w6929 & w1615) | (w8636 & w1615);
assign w3069 = ~w884 & w9032;
assign w3070 = w7412 & w9188;
assign w3071 = (~w5365 & w13501) | (~w5365 & w12940) | (w13501 & w12940);
assign w3072 = ~w3069 & w4026;
assign w3073 = (w13532 & w7002) | (w13532 & w8405) | (w7002 & w8405);
assign w3074 = ~w8244 & ~w9814;
assign w3075 = ~b47 & ~a47;
assign w3076 = (~w7926 & w12123) | (~w7926 & w10053) | (w12123 & w10053);
assign w3077 = ~w142 & ~w12642;
assign w3078 = w2083 & w2757;
assign w3079 = (w4627 & w12980) | (w4627 & w3376) | (w12980 & w3376);
assign w3080 = (w259 & w10896) | (w259 & w8337) | (w10896 & w8337);
assign w3081 = ~w922 & w5178;
assign w3082 = (~w5406 & w8191) | (~w5406 & ~w9004) | (w8191 & ~w9004);
assign w3083 = w11779 & w9707;
assign w3084 = w2656 & ~w13596;
assign w3085 = w13794 & ~w9989;
assign w3086 = (w12460 & w8234) | (w12460 & w1417) | (w8234 & w1417);
assign w3087 = ~w13713 & ~w12330;
assign w3088 = (w3745 & w11982) | (w3745 & w13746) | (w11982 & w13746);
assign w3089 = (~w1986 & w446) | (~w1986 & w6587) | (w446 & w6587);
assign w3090 = w14373 & ~w748;
assign w3091 = w3917 & ~w3500;
assign w3092 = w13799 & w1877;
assign w3093 = (w9510 & w5119) | (w9510 & ~w12293) | (w5119 & ~w12293);
assign w3094 = w6325 & w9288;
assign w3095 = (w8228 & w9034) | (w8228 & w217) | (w9034 & w217);
assign w3096 = w9623 & ~w11031;
assign w3097 = ~w4719 & ~w7698;
assign w3098 = b53 & a53;
assign w3099 = w9284 & w6500;
assign w3100 = w3175 & w2954;
assign w3101 = ~w7488 & w14047;
assign w3102 = w12589 & ~w1114;
assign w3103 = ~w13530 & ~w13491;
assign w3104 = w3338 & w854;
assign w3105 = (~w9608 & w1626) | (~w9608 & w9581) | (w1626 & w9581);
assign w3106 = (w1190 & w5719) | (w1190 & w4519) | (w5719 & w4519);
assign w3107 = w8183 & w2701;
assign w3108 = w7365 & ~w12311;
assign w3109 = w8154 & ~w11951;
assign w3110 = ~w13222 & ~w3699;
assign w3111 = w9949 & w2941;
assign w3112 = ~w858 & ~w3727;
assign w3113 = (w3036 & w12980) | (w3036 & w5832) | (w12980 & w5832);
assign w3114 = w13244 & ~w9860;
assign w3115 = ~w12891 & w13446;
assign w3116 = w13743 & w9110;
assign w3117 = ~w5522 & ~w5282;
assign w3118 = w7267 & w637;
assign w3119 = (~w11973 & w1731) | (~w11973 & w1897) | (w1731 & w1897);
assign w3120 = w13839 & w12545;
assign w3121 = w3734 & w8018;
assign w3122 = w12112 & ~w6219;
assign w3123 = ~w13944 & ~w1318;
assign w3124 = (~w3251 & w8719) | (~w3251 & w8566) | (w8719 & w8566);
assign w3125 = w11500 & w10997;
assign w3126 = w2464 & ~w12642;
assign w3127 = ~w1669 & ~w2002;
assign w3128 = (~w183 & ~w13587) | (~w183 & w6923) | (~w13587 & w6923);
assign w3129 = (~w7042 & w2080) | (~w7042 & w10760) | (w2080 & w10760);
assign w3130 = ~b125 & ~a125;
assign w3131 = ~w254 & w37;
assign w3132 = w1368 & w10261;
assign w3133 = w14648 & ~w1549;
assign w3134 = (w10435 & w12279) | (w10435 & w13484) | (w12279 & w13484);
assign w3135 = ~w6135 & ~w7305;
assign w3136 = w13733 & w3957;
assign w3137 = w4193 & w2101;
assign w3138 = w3577 & w14531;
assign w3139 = w11458 & ~w8781;
assign w3140 = w3385 | ~w1260;
assign w3141 = (w14462 & w12122) | (w14462 & w4057) | (w12122 & w4057);
assign w3142 = ~w4820 & ~w5053;
assign w3143 = (w9021 & ~w13401) | (w9021 & w11339) | (~w13401 & w11339);
assign w3144 = w12141 & w14420;
assign w3145 = w14226 & ~w14643;
assign w3146 = w8035 & ~w5243;
assign w3147 = ~w7541 & ~w2093;
assign w3148 = w4836 & w6113;
assign w3149 = w844 & w4818;
assign w3150 = w4449 & ~w10122;
assign w3151 = (~w6563 & w13803) | (~w6563 & w12307) | (w13803 & w12307);
assign w3152 = (w4855 & w5490) | (w4855 & w14342) | (w5490 & w14342);
assign w3153 = w5004 & w8708;
assign w3154 = w9977 & w11575;
assign w3155 = (w9547 & w1942) | (w9547 & w12000) | (w1942 & w12000);
assign w3156 = (w8900 & w13964) | (w8900 & w7795) | (w13964 & w7795);
assign w3157 = w1935 & ~w5209;
assign w3158 = ~w8512 & ~w6572;
assign w3159 = ~b40 & ~a40;
assign w3160 = (~w5193 & ~w6167) | (~w5193 & w9405) | (~w6167 & w9405);
assign w3161 = w5605 & w2928;
assign w3162 = w9679 & w14183;
assign w3163 = (w5651 & w2716) | (w5651 & w2990) | (w2716 & w2990);
assign w3164 = ~w9498 & ~w13492;
assign w3165 = ~w12317 & w3767;
assign w3166 = w12371 & ~w11861;
assign w3167 = (w1013 & w4285) | (w1013 & ~w7999) | (w4285 & ~w7999);
assign w3168 = ~w14478 & ~w14152;
assign w3169 = (w10172 & w9892) | (w10172 & w8228) | (w9892 & w8228);
assign w3170 = w1087 & w1606;
assign w3171 = ~w12378 & w11288;
assign w3172 = (~w3128 & w2049) | (~w3128 & w508) | (w2049 & w508);
assign w3173 = ~w3815 & ~w13387;
assign w3174 = w11586 & w7474;
assign w3175 = ~w4700 & ~w142;
assign w3176 = ~w7348 & w2632;
assign w3177 = (~w10139 & w345) | (~w10139 & w5486) | (w345 & w5486);
assign w3178 = w3288 & ~w7670;
assign w3179 = (~w2159 & w4032) | (~w2159 & w14486) | (w4032 & w14486);
assign w3180 = (w4361 & w10572) | (w4361 & w14576) | (w10572 & w14576);
assign w3181 = ~w1516 & ~w5224;
assign w3182 = ~w142 & ~w13323;
assign w3183 = (w4787 & ~w3044) | (w4787 & w5873) | (~w3044 & w5873);
assign w3184 = ~w4751 & w4425;
assign w3185 = ~w12121 & w8521;
assign w3186 = ~w3674 | ~w5694;
assign w3187 = w5865 & ~w3502;
assign w3188 = ~w10997 & ~w12911;
assign w3189 = ~w1795 & w13820;
assign w3190 = (w12642 & ~w635) | (w12642 & w7117) | (~w635 & w7117);
assign w3191 = w10629 & w6041;
assign w3192 = w2031 & w4003;
assign w3193 = (w9027 & w7917) | (w9027 & w2402) | (w7917 & w2402);
assign w3194 = w2729 & w13323;
assign w3195 = (~w11634 & w5277) | (~w11634 & w10908) | (w5277 & w10908);
assign w3196 = (w11201 & w667) | (w11201 & ~w7077) | (w667 & ~w7077);
assign w3197 = w3330 & w10903;
assign w3198 = (w1712 & w12265) | (w1712 & w2733) | (w12265 & w2733);
assign w3199 = w4203 & w9237;
assign w3200 = w13730 & w14569;
assign w3201 = w12464 & ~w2067;
assign w3202 = w1710 & w878;
assign w3203 = w12232 & w12812;
assign w3204 = w1452 & ~w1460;
assign w3205 = (w14514 & w6546) | (w14514 & w9295) | (w6546 & w9295);
assign w3206 = (w13168 & w1072) | (w13168 & ~w3095) | (w1072 & ~w3095);
assign w3207 = (w8130 & w10209) | (w8130 & w11970) | (w10209 & w11970);
assign w3208 = ~w1322 & w5621;
assign w3209 = ~w984 & ~w5582;
assign w3210 = w3963 & ~w13370;
assign w3211 = ~w13368 & w1622;
assign w3212 = w12438 & ~w5693;
assign w3213 = ~w5867 & ~w11068;
assign w3214 = ~w11975 & w3465;
assign w3215 = b68 & a68;
assign w3216 = w6836 & w4541;
assign w3217 = (~w10483 & w6805) | (~w10483 & w6702) | (w6805 & w6702);
assign w3218 = ~w905 & ~w7367;
assign w3219 = b93 & a93;
assign w3220 = ~w210 & w4516;
assign w3221 = w3963 & ~w11954;
assign w3222 = ~w12121 & ~w5137;
assign w3223 = w11613 & ~w8374;
assign w3224 = (~w7754 & w11796) | (~w7754 & w7672) | (w11796 & w7672);
assign w3225 = w8740 & w6910;
assign w3226 = (~w1096 & w4032) | (~w1096 & w3359) | (w4032 & w3359);
assign w3227 = w5853 & w10965;
assign w3228 = (~w5918 & w5673) | (~w5918 & w7955) | (w5673 & w7955);
assign w3229 = ~w10078 & ~w9517;
assign w3230 = (~w7662 & w13587) | (~w7662 & w2761) | (w13587 & w2761);
assign w3231 = ~w5218 & w13358;
assign w3232 = w8169 & ~w12764;
assign w3233 = w3201 & ~w13382;
assign w3234 = (~w4632 & w10640) | (~w4632 & w7745) | (w10640 & w7745);
assign w3235 = ~w12997 & w2800;
assign w3236 = w11613 & w5513;
assign w3237 = (w10687 & w2156) | (w10687 & w9928) | (w2156 & w9928);
assign w3238 = w9471 & ~w273;
assign w3239 = ~w11351 & ~w10250;
assign w3240 = ~w9713 & ~w7065;
assign w3241 = (~w1052 & w13324) | (~w1052 & w5205) | (w13324 & w5205);
assign w3242 = ~w235 & ~w4881;
assign w3243 = ~w4213 & ~w12980;
assign w3244 = ~w6453 & w13373;
assign w3245 = ~w13300 & ~w6867;
assign w3246 = (~w756 & w12781) | (~w756 & ~w2263) | (w12781 & ~w2263);
assign w3247 = w6980 & w1968;
assign w3248 = ~w9747 & w9356;
assign w3249 = (w14455 & w8337) | (w14455 & w10384) | (w8337 & w10384);
assign w3250 = ~w13306 & ~w9121;
assign w3251 = b107 & a107;
assign w3252 = w5932 & w1692;
assign w3253 = ~w6795 & w5247;
assign w3254 = ~w14664 & w8944;
assign w3255 = w7001 & w3727;
assign w3256 = ~w13521 & ~w13423;
assign w3257 = (~w9305 & w13458) | (~w9305 & w2517) | (w13458 & w2517);
assign w3258 = (w1842 & w7548) | (w1842 & w1578) | (w7548 & w1578);
assign w3259 = (w5952 & w8271) | (w5952 & w352) | (w8271 & w352);
assign w3260 = w6293 & ~w13980;
assign w3261 = w4835 & ~w13606;
assign w3262 = ~w3209 & w884;
assign w3263 = w12642 & w1115;
assign w3264 = (~w9305 & w2818) | (~w9305 & w3343) | (w2818 & w3343);
assign w3265 = (~w5070 & w11157) | (~w5070 & w14341) | (w11157 & w14341);
assign w3266 = (~w9364 & w9733) | (~w9364 & w2595) | (w9733 & w2595);
assign w3267 = w6279 & w2624;
assign w3268 = w7889 & w10699;
assign w3269 = w5761 & w9792;
assign w3270 = (~w3502 & w9608) | (~w3502 & w1537) | (w9608 & w1537);
assign w3271 = ~w1260 & w5537;
assign w3272 = w1705 & w569;
assign w3273 = ~w5620 & w10997;
assign w3274 = ~w7890 & w967;
assign w3275 = w8920 & ~w857;
assign w3276 = w10315 & w14597;
assign w3277 = w7085 & w4405;
assign w3278 = ~w9609 & w8026;
assign w3279 = (w6572 & w2500) | (w6572 & w13766) | (w2500 & w13766);
assign w3280 = ~w2175 & w3440;
assign w3281 = ~w14622 & ~w13635;
assign w3282 = ~w12762 & w4790;
assign w3283 = w4319 & w5243;
assign w3284 = ~w7607 & ~w14560;
assign w3285 = ~w5156 & ~w7322;
assign w3286 = (~w14048 & ~w4317) | (~w14048 & ~w5435) | (~w4317 & ~w5435);
assign w3287 = w3727 & ~w9480;
assign w3288 = ~b106 & ~a106;
assign w3289 = (~w3786 & w11442) | (~w3786 & w9911) | (w11442 & w9911);
assign w3290 = (w2611 & w7870) | (w2611 & w7353) | (w7870 & w7353);
assign w3291 = (w719 & w634) | (w719 & w7614) | (w634 & w7614);
assign w3292 = (~w11855 & w9608) | (~w11855 & w8471) | (w9608 & w8471);
assign w3293 = (~w12884 & w5671) | (~w12884 & w14472) | (w5671 & w14472);
assign w3294 = ~w8234 & ~w1263;
assign w3295 = w9854 & w9989;
assign w3296 = w3968 & ~w9380;
assign w3297 = w11169 & w6504;
assign w3298 = (w2648 & w3418) | (w2648 & w9484) | (w3418 & w9484);
assign w3299 = w48 & ~w3085;
assign w3300 = (~w2492 & w13958) | (~w2492 & w1432) | (w13958 & w1432);
assign w3301 = w10483 & ~w1172;
assign w3302 = ~w607 & ~w13839;
assign w3303 = ~w13769 & ~w4782;
assign w3304 = (w10079 & w3598) | (w10079 & w12861) | (w3598 & w12861);
assign w3305 = ~w5852 & w13854;
assign w3306 = ~w71 & w2391;
assign w3307 = ~w3934 & w12149;
assign w3308 = w1498 & w7877;
assign w3309 = (w2962 & ~w9159) | (w2962 & w4048) | (~w9159 & w4048);
assign w3310 = w9284 & w1062;
assign w3311 = w5177 & w6421;
assign w3312 = w10676 & w5742;
assign w3313 = ~w14000 & w6476;
assign w3314 = w12415 & ~w4023;
assign w3315 = w8871 & w14501;
assign w3316 = ~w896 & w3727;
assign w3317 = ~w309 & ~w1171;
assign w3318 = w347 & ~w45;
assign w3319 = (w12666 & w2766) | (w12666 & w10620) | (w2766 & w10620);
assign w3320 = w3587 & ~w9412;
assign w3321 = ~w2922 & ~w8328;
assign w3322 = ~w4836 & w884;
assign w3323 = w11586 & ~w10486;
assign w3324 = ~w4780 & ~w11827;
assign w3325 = w14504 & w9265;
assign w3326 = (~w13620 & w12206) | (~w13620 & w3209) | (w12206 & w3209);
assign w3327 = ~w11642 & ~w5594;
assign w3328 = ~w9543 & ~w11985;
assign w3329 = w12709 & ~w12106;
assign w3330 = (w6301 & w13848) | (w6301 & w7485) | (w13848 & w7485);
assign w3331 = w14557 & ~w688;
assign w3332 = w4787 & ~w2320;
assign w3333 = ~w4842 & ~w6379;
assign w3334 = ~w7190 & w12060;
assign w3335 = (~w11385 & w41) | (~w11385 & w7275) | (w41 & w7275);
assign w3336 = w36 & w2773;
assign w3337 = ~w2933 & ~w8171;
assign w3338 = ~w4246 & w10638;
assign w3339 = ~w14640 & ~w7670;
assign w3340 = (w6042 & w14479) | (w6042 & w10438) | (w14479 & w10438);
assign w3341 = ~w5779 & w6051;
assign w3342 = (~w7630 & w1903) | (~w7630 & w11909) | (w1903 & w11909);
assign w3343 = w14518 & ~w10624;
assign w3344 = w552 & w13355;
assign w3345 = ~w9625 & ~w1080;
assign w3346 = ~w4700 & w10182;
assign w3347 = (w6219 & w4520) | (w6219 & w3702) | (w4520 & w3702);
assign w3348 = ~w8567 & ~w7611;
assign w3349 = (w12636 & w227) | (w12636 & w13152) | (w227 & w13152);
assign w3350 = w3137 & w15;
assign w3351 = ~w922 & w10225;
assign w3352 = w7669 & ~w8363;
assign w3353 = w7970 & w10515;
assign w3354 = w2698 & ~w12416;
assign w3355 = (~w13685 & w12198) | (~w13685 & w4916) | (w12198 & w4916);
assign w3356 = w3015 & w139;
assign w3357 = ~w2751 & w12152;
assign w3358 = ~w7376 & w12893;
assign w3359 = w3971 & ~w1096;
assign w3360 = w4598 & w11446;
assign w3361 = ~w8110 & ~w475;
assign w3362 = w11613 & w10042;
assign w3363 = w1332 & w6689;
assign w3364 = w7726 & ~w6542;
assign w3365 = w3885 & w3904;
assign w3366 = ~w7794 & w8528;
assign w3367 = w235 & ~w1540;
assign w3368 = w8733 & w6826;
assign w3369 = ~w11735 & w12589;
assign w3370 = (w4859 & w1609) | (w4859 & w11841) | (w1609 & w11841);
assign w3371 = (~w9762 & w8136) | (~w9762 & w11348) | (w8136 & w11348);
assign w3372 = (w7433 & w8089) | (w7433 & w515) | (w8089 & w515);
assign w3373 = w9211 & w2909;
assign w3374 = w8345 & w5177;
assign w3375 = (w12915 & ~w12278) | (w12915 & w9784) | (~w12278 & w9784);
assign w3376 = w4213 & w4627;
assign w3377 = (w11117 & ~w9163) | (w11117 & w4152) | (~w9163 & w4152);
assign w3378 = (~w3317 & w6491) | (~w3317 & ~w2632) | (w6491 & ~w2632);
assign w3379 = ~w7001 & ~w2701;
assign w3380 = w724 & w8285;
assign w3381 = (w6293 & w7515) | (w6293 & w4413) | (w7515 & w4413);
assign w3382 = (~w5568 & w13324) | (~w5568 & w519) | (w13324 & w519);
assign w3383 = (~w2159 & w6699) | (~w2159 & w12528) | (w6699 & w12528);
assign w3384 = w95 & w11009;
assign w3385 = ~w5767 & ~w1260;
assign w3386 = ~w10523 & ~w475;
assign w3387 = ~w13587 & w4554;
assign w3388 = ~w4741 & w13985;
assign w3389 = (w1859 & w5815) | (w1859 & w2670) | (w5815 & w2670);
assign w3390 = ~w12240 & ~w7097;
assign w3391 = w9055 & w12301;
assign w3392 = ~w3012 & ~w928;
assign w3393 = w11533 & ~w5247;
assign w3394 = (w11902 & w12980) | (w11902 & w10770) | (w12980 & w10770);
assign w3395 = ~w10503 & ~w5227;
assign w3396 = w3146 | ~w5243;
assign w3397 = w11164 & ~w12549;
assign w3398 = w10290 & w1707;
assign w3399 = (~w12239 & w13724) | (~w12239 & w3591) | (w13724 & w3591);
assign w3400 = w3904 & w11861;
assign w3401 = (~w9613 & w5317) | (~w9613 & w12630) | (w5317 & w12630);
assign w3402 = ~w3133 & w736;
assign w3403 = ~w343 & ~w2713;
assign w3404 = (w8106 & w233) | (w8106 & w14384) | (w233 & w14384);
assign w3405 = ~w13321 & w2839;
assign w3406 = w3038 & ~w6572;
assign w3407 = w9480 & ~w7889;
assign w3408 = ~w1919 & ~w10295;
assign w3409 = (w8424 & w1409) | (w8424 & w11881) | (w1409 & w11881);
assign w3410 = (~w6580 & w11871) | (~w6580 & w8304) | (w11871 & w8304);
assign w3411 = (w4362 & ~w9915) | (w4362 & w11322) | (~w9915 & w11322);
assign w3412 = w5515 & w10176;
assign w3413 = w8191 & ~w5406;
assign w3414 = (~w13685 & w11220) | (~w13685 & w726) | (w11220 & w726);
assign w3415 = w12088 & w4658;
assign w3416 = ~w9116 & ~w8775;
assign w3417 = (w11708 & w3809) | (w11708 & w894) | (w3809 & w894);
assign w3418 = (w13776 & w2648) | (w13776 & ~w6920) | (w2648 & ~w6920);
assign w3419 = ~w10997 & w11744;
assign w3420 = w11798 & ~w4697;
assign w3421 = ~w14054 & w7189;
assign w3422 = ~w6696 & ~w7202;
assign w3423 = (w7782 & w5120) | (w7782 & w14232) | (w5120 & w14232);
assign w3424 = ~w6700 & ~w7087;
assign w3425 = w14276 & w10699;
assign w3426 = ~w5867 & ~w13953;
assign w3427 = ~w1838 & ~w8253;
assign w3428 = (~w6802 & w13690) | (~w6802 & w5377) | (w13690 & w5377);
assign w3429 = w9256 & ~w2228;
assign w3430 = w3483 & w9004;
assign w3431 = ~w1474 & w11861;
assign w3432 = ~w11487 & w3526;
assign w3433 = ~w3219 & ~w12958;
assign w3434 = (w13196 & w9815) | (w13196 & w9714) | (w9815 & w9714);
assign w3435 = (~w14227 & w12317) | (~w14227 & w13529) | (w12317 & w13529);
assign w3436 = (~w62 & w9993) | (~w62 & w12692) | (w9993 & w12692);
assign w3437 = ~w183 & w12170;
assign w3438 = (w9873 & w9640) | (w9873 & ~w3885) | (w9640 & ~w3885);
assign w3439 = w7762 & ~w11487;
assign w3440 = ~w3914 & ~w13073;
assign w3441 = ~w10676 & w12170;
assign w3442 = ~w10433 & w2559;
assign w3443 = ~w6377 & w7701;
assign w3444 = ~w11198 & ~w11117;
assign w3445 = w5294 & ~w2575;
assign w3446 = ~w14662 & ~w12378;
assign w3447 = ~w10675 & ~w11216;
assign w3448 = ~w8459 & ~w9348;
assign w3449 = ~w1785 & w6582;
assign w3450 = w9851 & ~w7210;
assign w3451 = ~w5522 & ~w9296;
assign w3452 = (w9749 & w10499) | (w9749 & w2328) | (w10499 & w2328);
assign w3453 = (w2655 & w1505) | (w2655 & w10194) | (w1505 & w10194);
assign w3454 = (~w2850 & w4512) | (~w2850 & w11851) | (w4512 & w11851);
assign w3455 = (~w13980 & w2773) | (~w13980 & w12824) | (w2773 & w12824);
assign w3456 = w9296 & w1062;
assign w3457 = w6358 & w8769;
assign w3458 = w8904 | ~w9454;
assign w3459 = (w852 & w7488) | (w852 & w6609) | (w7488 & w6609);
assign w3460 = (w1849 & w856) | (w1849 & w6768) | (w856 & w6768);
assign w3461 = (~w10450 & w1470) | (~w10450 & w817) | (w1470 & w817);
assign w3462 = (~w10669 & w13152) | (~w10669 & w11839) | (w13152 & w11839);
assign w3463 = ~w2352 & w9358;
assign w3464 = (w378 & w8983) | (w378 & w10310) | (w8983 & w10310);
assign w3465 = (~w91 & w11132) | (~w91 & w3981) | (w11132 & w3981);
assign w3466 = w1563 & w1821;
assign w3467 = ~w13744 & w7634;
assign w3468 = w11273 & w11658;
assign w3469 = (~w706 & w8294) | (~w706 & w794) | (w8294 & w794);
assign w3470 = w922 & w11395;
assign w3471 = w5156 & w14447;
assign w3472 = ~w7141 & w1236;
assign w3473 = (~w10946 & w12710) | (~w10946 & w3800) | (w12710 & w3800);
assign w3474 = (w813 & w1172) | (w813 & w4574) | (w1172 & w4574);
assign w3475 = (w11287 & w4357) | (w11287 & w3926) | (w4357 & w3926);
assign w3476 = w9912 | ~w7637;
assign w3477 = (w14346 & w9746) | (w14346 & ~w3266) | (w9746 & ~w3266);
assign w3478 = (w14664 & w7570) | (w14664 & w2770) | (w7570 & w2770);
assign w3479 = w3550 & w9051;
assign w3480 = w3181 & ~w6825;
assign w3481 = ~w8239 & w10488;
assign w3482 = w11441 & ~w5678;
assign w3483 = w6542 & ~w5860;
assign w3484 = ~w3568 & ~w9412;
assign w3485 = (~w10318 & w3323) | (~w10318 & w11036) | (w3323 & w11036);
assign w3486 = ~w13268 & w11239;
assign w3487 = ~w12613 & w12268;
assign w3488 = ~w8937 & w13289;
assign w3489 = (~w13521 & w12571) | (~w13521 & w749) | (w12571 & w749);
assign w3490 = (~w6802 & w2255) | (~w6802 & w8467) | (w2255 & w8467);
assign w3491 = ~w14629 & ~w3181;
assign w3492 = (~w7737 & ~w11586) | (~w7737 & w14443) | (~w11586 & w14443);
assign w3493 = (w4587 & w13152) | (w4587 & w2826) | (w13152 & w2826);
assign w3494 = ~w5490 & w7612;
assign w3495 = (~w6426 & w9028) | (~w6426 & w2721) | (w9028 & w2721);
assign w3496 = ~w3034 & w4371;
assign w3497 = (w12376 & w186) | (w12376 & w10268) | (w186 & w10268);
assign w3498 = w13591 & w7675;
assign w3499 = w5389 & w7023;
assign w3500 = (w10123 & w9683) | (w10123 & w7339) | (w9683 & w7339);
assign w3501 = ~w6886 & w13381;
assign w3502 = b66 & a66;
assign w3503 = w12732 & ~w8304;
assign w3504 = w2797 & w5776;
assign w3505 = ~w5161 & w3191;
assign w3506 = (~w6816 & w12980) | (~w6816 & w6916) | (w12980 & w6916);
assign w3507 = (~w101 & w14001) | (~w101 & w11889) | (w14001 & w11889);
assign w3508 = ~b79 & ~a79;
assign w3509 = (~w6045 & w2175) | (~w6045 & w1713) | (w2175 & w1713);
assign w3510 = w14309 & ~w13621;
assign w3511 = w12783 & w13463;
assign w3512 = ~w13971 & w10699;
assign w3513 = ~w8171 & w4706;
assign w3514 = (w11610 & w4526) | (w11610 & w9488) | (w4526 & w9488);
assign w3515 = ~w5178 & w8419;
assign w3516 = (~w12464 & ~w7218) | (~w12464 & w5037) | (~w7218 & w5037);
assign w3517 = w5040 & w13037;
assign w3518 = w9147 & ~w7188;
assign w3519 = w11708 & ~w12054;
assign w3520 = (~w7654 & ~w3846) | (~w7654 & ~w14534) | (~w3846 & ~w14534);
assign w3521 = (w2116 & w10588) | (w2116 & w8689) | (w10588 & w8689);
assign w3522 = (~w4291 & w12003) | (~w4291 & w12230) | (w12003 & w12230);
assign w3523 = ~w11905 & w4456;
assign w3524 = ~w11488 & ~w11108;
assign w3525 = (w6423 & w10528) | (w6423 & w1976) | (w10528 & w1976);
assign w3526 = ~w8893 & w13838;
assign w3527 = ~w142 & ~w12943;
assign w3528 = ~w9252 & w1062;
assign w3529 = w10880 & ~w8080;
assign w3530 = ~w16 & ~w9716;
assign w3531 = (w3039 & ~w1692) | (w3039 & w6728) | (~w1692 & w6728);
assign w3532 = ~w142 & ~b78;
assign w3533 = w10241 & w5135;
assign w3534 = ~w770 & w2720;
assign w3535 = w1014 & w4333;
assign w3536 = ~w1452 & ~w11836;
assign w3537 = (w8614 & w4590) | (w8614 & w2) | (w4590 & w2);
assign w3538 = ~w13587 & w1302;
assign w3539 = ~w11462 & w13885;
assign w3540 = w3982 & ~w5014;
assign w3541 = (~w11211 & ~w13885) | (~w11211 & ~w9139) | (~w13885 & ~w9139);
assign w3542 = ~w142 & ~w10182;
assign w3543 = ~w12291 & w2838;
assign w3544 = ~w2223 & ~w14591;
assign w3545 = (~w3550 & w9974) | (~w3550 & w12016) | (w9974 & w12016);
assign w3546 = ~w9012 & w11114;
assign w3547 = ~w12273 & ~w1930;
assign w3548 = ~w1712 & ~w14548;
assign w3549 = w4140 & ~w4155;
assign w3550 = ~w9422 & ~w1029;
assign w3551 = (~w12992 & w1351) | (~w12992 & w5475) | (w1351 & w5475);
assign w3552 = ~w1434 & ~w12288;
assign w3553 = ~w14571 & ~w13943;
assign w3554 = w922 & ~w12988;
assign w3555 = ~w13720 & ~w9230;
assign w3556 = (~w5385 & w7709) | (~w5385 & ~w4709) | (w7709 & ~w4709);
assign w3557 = w12488 & ~w10004;
assign w3558 = w5177 & w3219;
assign w3559 = w11431 & w9286;
assign w3560 = ~w8648 & w11199;
assign w3561 = w1821 & w876;
assign w3562 = w7135 & ~w4340;
assign w3563 = ~w13306 & ~w3885;
assign w3564 = w12464 & ~w3209;
assign w3565 = w11680 & ~w3424;
assign w3566 = w5490 & w11123;
assign w3567 = ~w14569 & ~w9812;
assign w3568 = ~b21 & ~a21;
assign w3569 = w14396 & w14304;
assign w3570 = w10339 & w8013;
assign w3571 = (w4545 & w11229) | (w4545 & w5512) | (w11229 & w5512);
assign w3572 = (w6183 & w495) | (w6183 & w12966) | (w495 & w12966);
assign w3573 = w12567 & w6845;
assign w3574 = w10300 & w13839;
assign w3575 = w10224 & w11655;
assign w3576 = ~w9244 & w1764;
assign w3577 = w7042 & ~w12726;
assign w3578 = (w14390 & w12499) | (w14390 & w14595) | (w12499 & w14595);
assign w3579 = (w10625 & w11149) | (w10625 & ~w2305) | (w11149 & ~w2305);
assign w3580 = ~w4158 & w10705;
assign w3581 = (w13227 & w4741) | (w13227 & w3015) | (w4741 & w3015);
assign w3582 = ~w8254 & w3690;
assign w3583 = ~w12131 & ~w4071;
assign w3584 = (~w12893 & w11635) | (~w12893 & w8974) | (w11635 & w8974);
assign w3585 = ~w9751 & w10902;
assign w3586 = w10431 & ~w11757;
assign w3587 = ~b20 & ~a20;
assign w3588 = w13596 & ~w8419;
assign w3589 = ~w12553 & ~w1608;
assign w3590 = w607 & ~w2941;
assign w3591 = ~w13522 & w10915;
assign w3592 = ~w3675 & ~w6740;
assign w3593 = w9163 & w8618;
assign w3594 = ~w5787 & ~w2558;
assign w3595 = w9073 & w1033;
assign w3596 = w2155 & w12717;
assign w3597 = ~w1738 & ~w13463;
assign w3598 = (w4202 & w2883) | (w4202 & ~w50) | (w2883 & ~w50);
assign w3599 = ~w6876 & ~w11225;
assign w3600 = ~w12271 & w1794;
assign w3601 = (~w2310 & w12474) | (~w2310 & w3143) | (w12474 & w3143);
assign w3602 = ~w3219 & ~w2850;
assign w3603 = ~w13521 & ~w4881;
assign w3604 = ~w9810 & w14519;
assign w3605 = ~w6542 & ~w7962;
assign w3606 = ~w3493 & ~w3771;
assign w3607 = (~w14455 & ~w8337) | (~w14455 & w7644) | (~w8337 & w7644);
assign w3608 = w8769 & w5630;
assign w3609 = ~w13526 & w3823;
assign w3610 = ~w4700 & w11031;
assign w3611 = ~b69 & ~a69;
assign w3612 = (~w7690 & w6947) | (~w7690 & w6531) | (w6947 & w6531);
assign w3613 = ~w1766 & ~w9078;
assign w3614 = w8328 & ~w1821;
assign w3615 = ~w803 & w12656;
assign w3616 = (w3635 & w4149) | (w3635 & w13713) | (w4149 & w13713);
assign w3617 = w8169 & ~w6770;
assign w3618 = ~w10234 & ~w6130;
assign w3619 = ~w3724 & w12171;
assign w3620 = (w653 & w4551) | (w653 & ~w5570) | (w4551 & ~w5570);
assign w3621 = w4809 & w1913;
assign w3622 = ~w10941 & w11861;
assign w3623 = ~w1096 & ~w12958;
assign w3624 = w8232 & ~w8347;
assign w3625 = ~w10978 & ~w12238;
assign w3626 = (w14313 & w3247) | (w14313 & w8605) | (w3247 & w8605);
assign w3627 = w4855 & w13824;
assign w3628 = (w8584 & w12614) | (w8584 & w2171) | (w12614 & w2171);
assign w3629 = (w6502 & ~w9541) | (w6502 & w6322) | (~w9541 & w6322);
assign w3630 = (~w2655 & w438) | (~w2655 & w670) | (w438 & w670);
assign w3631 = (~w9305 & w10238) | (~w9305 & w2078) | (w10238 & w2078);
assign w3632 = (~w852 & w10605) | (~w852 & w1702) | (w10605 & w1702);
assign w3633 = (~w3613 & w12453) | (~w3613 & w12254) | (w12453 & w12254);
assign w3634 = w1332 & w7667;
assign w3635 = (w5952 & w3004) | (w5952 & w3021) | (w3004 & w3021);
assign w3636 = ~w14276 & ~w9283;
assign w3637 = ~w2218 & w8478;
assign w3638 = (w7809 & w5318) | (w7809 & w8614) | (w5318 & w8614);
assign w3639 = ~w4359 & w6061;
assign w3640 = (w11416 & w1600) | (w11416 & w5051) | (w1600 & w5051);
assign w3641 = ~w13636 & w10213;
assign w3642 = ~w3768 & w1234;
assign w3643 = ~w3137 & w14021;
assign w3644 = ~w4158 & w10266;
assign w3645 = w6975 & ~w5785;
assign w3646 = w3682 & w1627;
assign w3647 = ~w4921 & w5469;
assign w3648 = (w10483 & w1057) | (w10483 & w8913) | (w1057 & w8913);
assign w3649 = (w10736 & w10117) | (w10736 & w4781) | (w10117 & w4781);
assign w3650 = ~w13754 & ~w9199;
assign w3651 = w4270 & w6689;
assign w3652 = w4449 & ~w1147;
assign w3653 = (w3292 & ~w13219) | (w3292 & w4035) | (~w13219 & w4035);
assign w3654 = ~w9793 & ~w3725;
assign w3655 = ~w14166 & w13127;
assign w3656 = ~w3101 & ~w8628;
assign w3657 = (w1711 & w12795) | (w1711 & w4179) | (w12795 & w4179);
assign w3658 = w7594 & ~w2379;
assign w3659 = ~w8819 & w3806;
assign w3660 = w13937 & ~w217;
assign w3661 = w3502 & w5865;
assign w3662 = ~w6135 & w8396;
assign w3663 = w7886 & w6251;
assign w3664 = (~w4938 & w13319) | (~w4938 & w14516) | (w13319 & w14516);
assign w3665 = ~w14045 & ~w1553;
assign w3666 = ~w80 & ~w5129;
assign w3667 = w7625 & w11508;
assign w3668 = ~w8182 & w14404;
assign w3669 = (w9442 & w9624) | (w9442 & ~w12036) | (w9624 & ~w12036);
assign w3670 = w8788 & ~w622;
assign w3671 = (~w2500 & w5454) | (~w2500 & w14654) | (w5454 & w14654);
assign w3672 = ~w4119 & ~w4124;
assign w3673 = ~w13282 & w2370;
assign w3674 = ~w14390 & w5694;
assign w3675 = (w9305 & w486) | (w9305 & w5695) | (w486 & w5695);
assign w3676 = ~w4033 & w10923;
assign w3677 = (w1378 & w10877) | (w1378 & ~w81) | (w10877 & ~w81);
assign w3678 = w12437 & w9599;
assign w3679 = w10290 & ~w1261;
assign w3680 = ~w11333 & w7012;
assign w3681 = ~w4447 & w14021;
assign w3682 = (~w9012 & w6010) | (~w9012 & w8653) | (w6010 & w8653);
assign w3683 = (w13924 & ~w8234) | (w13924 & w709) | (~w8234 & w709);
assign w3684 = w4798 & ~w10148;
assign w3685 = (~w563 & w2001) | (~w563 & w13061) | (w2001 & w13061);
assign w3686 = w7697 & w12676;
assign w3687 = ~w4129 & ~w11940;
assign w3688 = w8201 & w6539;
assign w3689 = ~w13587 & w7954;
assign w3690 = w3175 & ~w3166;
assign w3691 = ~w1194 & w1430;
assign w3692 = (~w894 & w5867) | (~w894 & w7962) | (w5867 & w7962);
assign w3693 = ~w4700 & w2701;
assign w3694 = w11041 & w14179;
assign w3695 = (w3655 & w14017) | (w3655 & w9392) | (w14017 & w9392);
assign w3696 = (w10409 & w9748) | (w10409 & w12483) | (w9748 & w12483);
assign w3697 = ~w13122 & w8869;
assign w3698 = w12656 & w2323;
assign w3699 = ~w3906 & ~w11438;
assign w3700 = ~w14574 & ~w7247;
assign w3701 = w2486 & w13137;
assign w3702 = (w5768 & w13772) | (w5768 & w11037) | (w13772 & w11037);
assign w3703 = ~w13222 & w9226;
assign w3704 = (~w1949 & w4512) | (~w1949 & w9186) | (w4512 & w9186);
assign w3705 = ~w13282 & w7668;
assign w3706 = (w7722 & w1817) | (w7722 & w11278) | (w1817 & w11278);
assign w3707 = ~w3289 | ~w12125;
assign w3708 = (w7082 & w11832) | (w7082 & w14467) | (w11832 & w14467);
assign w3709 = (~w5227 & w13503) | (~w5227 & w3395) | (w13503 & w3395);
assign w3710 = (~w3747 & ~w13254) | (~w3747 & w12348) | (~w13254 & w12348);
assign w3711 = ~w2468 & ~w9454;
assign w3712 = (w2648 & w3418) | (w2648 & w405) | (w3418 & w405);
assign w3713 = ~w6239 & w6365;
assign w3714 = ~w5395 & ~w2232;
assign w3715 = ~w9165 & w4724;
assign w3716 = w13438 & w10050;
assign w3717 = b69 & a69;
assign w3718 = w12271 & w10477;
assign w3719 = w12531 & w14050;
assign w3720 = (~w2950 & ~w8356) | (~w2950 & w8740) | (~w8356 & w8740);
assign w3721 = (w11759 & ~w9983) | (w11759 & w5155) | (~w9983 & w5155);
assign w3722 = ~w14570 & w7478;
assign w3723 = w5099 & ~w6236;
assign w3724 = ~w2218 & w5536;
assign w3725 = (~w6802 & w14156) | (~w6802 & w10797) | (w14156 & w10797);
assign w3726 = ~w1048 & w1365;
assign w3727 = ~w10820 & ~w175;
assign w3728 = w772 & ~w2287;
assign w3729 = ~w1062 & ~w3963;
assign w3730 = (~w1221 & w12922) | (~w1221 & w4223) | (w12922 & w4223);
assign w3731 = w12701 & w11076;
assign w3732 = w309 & w4855;
assign w3733 = w11364 & w4039;
assign w3734 = ~w3019 & ~w8754;
assign w3735 = ~w5294 & w3215;
assign w3736 = w2065 & ~w3427;
assign w3737 = w9015 & ~w3025;
assign w3738 = w3128 & w7915;
assign w3739 = (w9663 & w2520) | (w9663 & w7568) | (w2520 & w7568);
assign w3740 = ~w9141 & ~w209;
assign w3741 = ~w7348 & w8331;
assign w3742 = ~b51 & ~a51;
assign w3743 = ~b53 & w13852;
assign w3744 = ~w9552 & w13954;
assign w3745 = (~w4325 & w12456) | (~w4325 & w2182) | (w12456 & w2182);
assign w3746 = ~w10185 & w10230;
assign w3747 = ~w7650 & w12693;
assign w3748 = (w8130 & w6019) | (w8130 & w12096) | (w6019 & w12096);
assign w3749 = ~w6897 & w4728;
assign w3750 = ~w2332 & w1274;
assign w3751 = ~b32 & ~a32;
assign w3752 = w4405 & ~w10916;
assign w3753 = (w11993 & w2754) | (w11993 & ~w3691) | (w2754 & ~w3691);
assign w3754 = w21 & w2147;
assign w3755 = ~w1369 & ~w6844;
assign w3756 = ~w12728 & ~w7424;
assign w3757 = (w9862 & w5996) | (w9862 & ~w11759) | (w5996 & ~w11759);
assign w3758 = (w6276 & w5492) | (w6276 & w10034) | (w5492 & w10034);
assign w3759 = b16 & a16;
assign w3760 = w3015 & ~w6310;
assign w3761 = (w3057 & w6709) | (w3057 & w12375) | (w6709 & w12375);
assign w3762 = w305 & ~w9184;
assign w3763 = w9704 & ~w3602;
assign w3764 = ~w10941 & w10645;
assign w3765 = ~w12252 & w1733;
assign w3766 = w3963 & ~w2073;
assign w3767 = ~w2410 & ~w14072;
assign w3768 = ~w11095 & w4308;
assign w3769 = w10704 & w4541;
assign w3770 = ~w3736 & w1090;
assign w3771 = (~w2544 & w12980) | (~w2544 & w8137) | (w12980 & w8137);
assign w3772 = (~w12537 & w13340) | (~w12537 & w13642) | (w13340 & w13642);
assign w3773 = (~w10331 & w7376) | (~w10331 & w10021) | (w7376 & w10021);
assign w3774 = ~w13222 & w13300;
assign w3775 = ~w922 & ~w4021;
assign w3776 = (w6637 & w5256) | (w6637 & w454) | (w5256 & w454);
assign w3777 = ~w6080 & ~w3727;
assign w3778 = w1574 & w3499;
assign w3779 = (~w10966 & ~w4103) | (~w10966 & w2190) | (~w4103 & w2190);
assign w3780 = w3038 & w8512;
assign w3781 = w7559 & ~w2678;
assign w3782 = w1016 & ~w5732;
assign w3783 = (w13193 & w7598) | (w13193 & ~w8228) | (w7598 & ~w8228);
assign w3784 = w3128 & w2483;
assign w3785 = ~w13073 & w3007;
assign w3786 = b47 & a47;
assign w3787 = (w11385 & w8385) | (w11385 & w12641) | (w8385 & w12641);
assign w3788 = w8459 & w2941;
assign w3789 = (~w888 & w2455) | (~w888 & w13486) | (w2455 & w13486);
assign w3790 = w7376 & w953;
assign w3791 = ~w8937 & w4086;
assign w3792 = ~w8234 & w199;
assign w3793 = (~w7085 & w12121) | (~w7085 & w1064) | (w12121 & w1064);
assign w3794 = ~w8991 & w8276;
assign w3795 = (~w6018 & ~w12153) | (~w6018 & w7999) | (~w12153 & w7999);
assign w3796 = (~w4287 & w2971) | (~w4287 & ~w4007) | (w2971 & ~w4007);
assign w3797 = ~w6542 & ~w4989;
assign w3798 = w3015 & ~w1639;
assign w3799 = (w5687 & ~w2912) | (w5687 & w1180) | (~w2912 & w1180);
assign w3800 = (w2941 & w4902) | (w2941 & ~w8785) | (w4902 & ~w8785);
assign w3801 = w13967 & w1882;
assign w3802 = w12708 & w9886;
assign w3803 = ~b31 & ~a31;
assign w3804 = ~w12988 & ~w2922;
assign w3805 = (~w6889 & w1121) | (~w6889 & ~w4174) | (w1121 & ~w4174);
assign w3806 = ~w12798 & w6280;
assign w3807 = ~w4921 & w5416;
assign w3808 = w1805 & ~w6818;
assign w3809 = w7962 & w11708;
assign w3810 = w8367 & w7482;
assign w3811 = (~w12842 & w7689) | (~w12842 & w4792) | (w7689 & w4792);
assign w3812 = ~w7365 & w2922;
assign w3813 = (~a93 & w4158) | (~a93 & w4000) | (w4158 & w4000);
assign w3814 = (w6886 & w2251) | (w6886 & w4646) | (w2251 & w4646);
assign w3815 = w3671 & w6251;
assign w3816 = w457 & w11530;
assign w3817 = (w2962 & w1708) | (w2962 & ~w14486) | (w1708 & ~w14486);
assign w3818 = (~w5569 & w13595) | (~w5569 & ~w13526) | (w13595 & ~w13526);
assign w3819 = ~w544 & ~w1075;
assign w3820 = (~w9672 & w5867) | (~w9672 & w5123) | (w5867 & w5123);
assign w3821 = (w7376 & w11198) | (w7376 & w11279) | (w11198 & w11279);
assign w3822 = (w6572 & w7488) | (w6572 & w3279) | (w7488 & w3279);
assign w3823 = (~w3508 & w6935) | (~w3508 & w8967) | (w6935 & w8967);
assign w3824 = w2320 & ~w5247;
assign w3825 = w10561 & w2544;
assign w3826 = ~w2514 & ~w1203;
assign w3827 = ~w7050 & ~w13515;
assign w3828 = ~w198 & w12618;
assign w3829 = ~w12483 & ~w10409;
assign w3830 = (~w10853 & w13222) | (~w10853 & w14162) | (w13222 & w14162);
assign w3831 = (~w11185 & w7274) | (~w11185 & w2963) | (w7274 & w2963);
assign w3832 = w13857 & ~w8992;
assign w3833 = w2964 | w1498;
assign w3834 = (~w6825 & w3480) | (~w6825 & w5657) | (w3480 & w5657);
assign w3835 = ~w10252 & w13335;
assign w3836 = ~w4312 & w7317;
assign w3837 = (w514 & w3624) | (w514 & w5359) | (w3624 & w5359);
assign w3838 = w8905 & w12250;
assign w3839 = ~w4966 & w4364;
assign w3840 = ~w7043 & ~w3901;
assign w3841 = (~w1627 & ~w1362) | (~w1627 & w3892) | (~w1362 & w3892);
assign w3842 = (w5070 & w7992) | (w5070 & w3932) | (w7992 & w3932);
assign w3843 = ~w10462 & w5248;
assign w3844 = w11747 & ~w6220;
assign w3845 = ~w7717 & ~w2384;
assign w3846 = w13872 & w2953;
assign w3847 = (w3446 & w3491) | (w3446 & w2469) | (w3491 & w2469);
assign w3848 = b53 & ~w10768;
assign w3849 = w6930 & w9566;
assign w3850 = (w8512 & w14661) | (w8512 & w3209) | (w14661 & w3209);
assign w3851 = ~w14227 & ~w12438;
assign w3852 = ~w5936 & ~w14291;
assign w3853 = (w1455 & w12771) | (w1455 & w10958) | (w12771 & w10958);
assign w3854 = (~w14395 & w12240) | (~w14395 & w5262) | (w12240 & w5262);
assign w3855 = ~w13282 & w2387;
assign w3856 = w13545 & ~w7551;
assign w3857 = ~w3044 & ~w9100;
assign w3858 = w10047 & w8527;
assign w3859 = w6556 & ~w7521;
assign w3860 = w7460 | w9698;
assign w3861 = w8911 & w9436;
assign w3862 = w8778 & ~w5052;
assign w3863 = ~w2070 & ~w10619;
assign w3864 = ~w607 & w6500;
assign w3865 = w4586 & w12614;
assign w3866 = w3135 | ~w7305;
assign w3867 = w14302 & ~w10247;
assign w3868 = ~w14469 & w9454;
assign w3869 = (~w341 & w1929) | (~w341 & w5992) | (w1929 & w5992);
assign w3870 = w9454 & w10853;
assign w3871 = w4787 & w5285;
assign w3872 = ~w13880 & ~w5710;
assign w3873 = w9694 & ~w5744;
assign w3874 = (w7734 & w8614) | (w7734 & w6819) | (w8614 & w6819);
assign w3875 = w13732 & w14021;
assign w3876 = ~w3309 & ~w3044;
assign w3877 = w8094 & w3671;
assign w3878 = (~w6427 & w12416) | (~w6427 & w6541) | (w12416 & w6541);
assign w3879 = w9454 & w5105;
assign w3880 = w11702 & ~w11553;
assign w3881 = (w7762 & w9866) | (w7762 & ~w225) | (w9866 & ~w225);
assign w3882 = ~w3325 & ~w12700;
assign w3883 = ~w9141 & w11904;
assign w3884 = w8909 & ~w5946;
assign w3885 = b52 & a52;
assign w3886 = ~w10334 & ~w3610;
assign w3887 = w9952 & w6064;
assign w3888 = w12271 & w5660;
assign w3889 = (~w8130 & w11514) | (~w8130 & w11237) | (w11514 & w11237);
assign w3890 = ~w1785 & w7352;
assign w3891 = ~w8330 & w3524;
assign w3892 = (~w9672 & w9012) | (~w9672 & w3820) | (w9012 & w3820);
assign w3893 = w7794 & ~w11546;
assign w3894 = ~w2317 & w4439;
assign w3895 = w1152 & w11049;
assign w3896 = (~w9928 & w1927) | (~w9928 & w12794) | (w1927 & w12794);
assign w3897 = ~w10462 & w5546;
assign w3898 = w4186 & w7622;
assign w3899 = (w9831 & ~w630) | (w9831 & w2948) | (~w630 & w2948);
assign w3900 = (w7889 & w8019) | (w7889 & w1734) | (w8019 & w1734);
assign w3901 = ~w8475 & w13323;
assign w3902 = ~w5157 & w3227;
assign w3903 = ~w2218 & w10617;
assign w3904 = ~w14614 & ~w13344;
assign w3905 = ~w11256 & w400;
assign w3906 = ~w3025 & ~w10855;
assign w3907 = (~w10923 & w3760) | (~w10923 & w3798) | (w3760 & w3798);
assign w3908 = ~w4236 & ~w6094;
assign w3909 = (w2116 & w2759) | (w2116 & w7016) | (w2759 & w7016);
assign w3910 = ~w6238 & ~w3495;
assign w3911 = (~w2857 & ~w10624) | (~w2857 & ~w9305) | (~w10624 & ~w9305);
assign w3912 = ~w10855 & w1387;
assign w3913 = w11855 & ~w1620;
assign w3914 = ~w1598 & ~w3182;
assign w3915 = (w1013 & w4285) | (w1013 & ~w14074) | (w4285 & ~w14074);
assign w3916 = ~w14141 & w11903;
assign w3917 = ~w1696 & ~w10927;
assign w3918 = (w694 & w10958) | (w694 & w8692) | (w10958 & w8692);
assign w3919 = (w5675 & w227) | (w5675 & w2175) | (w227 & w2175);
assign w3920 = (w9305 & w13961) | (w9305 & w13822) | (w13961 & w13822);
assign w3921 = ~w142 & w9244;
assign w3922 = ~w7013 & w4033;
assign w3923 = (~w5694 & ~w3674) | (~w5694 & w4796) | (~w3674 & w4796);
assign w3924 = ~w4080 & w1587;
assign w3925 = ~w13721 & w4518;
assign w3926 = (~w9719 & w28) | (~w9719 & w12933) | (w28 & w12933);
assign w3927 = w12460 & w2076;
assign w3928 = ~w1864 & w11055;
assign w3929 = (~w2445 & w1169) | (~w2445 & w11816) | (w1169 & w11816);
assign w3930 = (w4353 & ~w7725) | (w4353 & w8610) | (~w7725 & w8610);
assign w3931 = (~w343 & w9614) | (~w343 & w12046) | (w9614 & w12046);
assign w3932 = (~w4515 & w8693) | (~w4515 & w8607) | (w8693 & w8607);
assign w3933 = (w8 & w13819) | (w8 & w8337) | (w13819 & w8337);
assign w3934 = w11043 & w4073;
assign w3935 = ~w2705 & w11146;
assign w3936 = ~w4751 & w1395;
assign w3937 = w141 & w3422;
assign w3938 = ~w10334 & ~w3346;
assign w3939 = (w3753 & w255) | (w3753 & ~w13524) | (w255 & ~w13524);
assign w3940 = ~w1244 & ~w13008;
assign w3941 = w13189 & ~w5282;
assign w3942 = w10477 & w7423;
assign w3943 = ~w6741 & w1133;
assign w3944 = ~w5559 & ~w12464;
assign w3945 = w4058 & ~w6737;
assign w3946 = w2480 & w12678;
assign w3947 = (~w11934 & w5701) | (~w11934 & w4911) | (w5701 & w4911);
assign w3948 = (w4756 & w14151) | (w4756 & w4466) | (w14151 & w4466);
assign w3949 = ~w4501 & w4962;
assign w3950 = ~w6920 & w2506;
assign w3951 = w5732 & w6230;
assign w3952 = w7896 & w3349;
assign w3953 = (w5694 & ~w2692) | (w5694 & ~w3957) | (~w2692 & ~w3957);
assign w3954 = (~w8294 & w8016) | (~w8294 & w2527) | (w8016 & w2527);
assign w3955 = ~w4914 & w14121;
assign w3956 = ~w6583 & ~w690;
assign w3957 = w14504 & w10880;
assign w3958 = (~w1096 & w13214) | (~w1096 & w1103) | (w13214 & w1103);
assign w3959 = (w10457 & w2152) | (w10457 & w6894) | (w2152 & w6894);
assign w3960 = (w9305 & w10844) | (w9305 & w12494) | (w10844 & w12494);
assign w3961 = ~w4213 & w569;
assign w3962 = w7263 & w8865;
assign w3963 = ~w7001 & ~w7244;
assign w3964 = w9805 & w5788;
assign w3965 = w1867 & w1362;
assign w3966 = ~w12958 & w11500;
assign w3967 = ~w892 & w11034;
assign w3968 = ~w10740 & w2420;
assign w3969 = (~w5841 & w6587) | (~w5841 & w655) | (w6587 & w655);
assign w3970 = ~w4700 & w11117;
assign w3971 = ~w8754 & ~w2933;
assign w3972 = (w13899 & ~w11925) | (w13899 & w5713) | (~w11925 & w5713);
assign w3973 = (w9096 & w6950) | (w9096 & w6284) | (w6950 & w6284);
assign w3974 = (~w318 & w11516) | (~w318 & ~w4709) | (w11516 & ~w4709);
assign w3975 = (w12646 & w7427) | (w12646 & w9117) | (w7427 & w9117);
assign w3976 = (~w7122 & w13152) | (~w7122 & w11235) | (w13152 & w11235);
assign w3977 = ~w7962 & ~w894;
assign w3978 = w14086 & ~w8267;
assign w3979 = (~w5702 & w105) | (~w5702 & w7254) | (w105 & w7254);
assign w3980 = (w6542 & w10462) | (w6542 & w11024) | (w10462 & w11024);
assign w3981 = (~w6700 & w6192) | (~w6700 & ~w6427) | (w6192 & ~w6427);
assign w3982 = ~w13256 & ~w9412;
assign w3983 = (w7376 & w11198) | (w7376 & w14218) | (w11198 & w14218);
assign w3984 = (w3386 & w3730) | (w3386 & w11392) | (w3730 & w11392);
assign w3985 = (~w7962 & w3914) | (~w7962 & w3605) | (w3914 & w3605);
assign w3986 = ~w12664 & w7306;
assign w3987 = w7681 & ~w8253;
assign w3988 = ~w4688 & ~w14639;
assign w3989 = (w11138 & w3660) | (w11138 & w5501) | (w3660 & w5501);
assign w3990 = w6433 & ~w14291;
assign w3991 = ~w13344 & ~w2707;
assign w3992 = (w9871 & w10462) | (w9871 & w12333) | (w10462 & w12333);
assign w3993 = w12460 & ~w11804;
assign w3994 = ~w13183 & ~w20;
assign w3995 = ~w10695 & ~w10142;
assign w3996 = ~w8791 & ~w10712;
assign w3997 = ~w9145 & ~w6406;
assign w3998 = (~w2144 & w11930) | (~w2144 & w998) | (w11930 & w998);
assign w3999 = ~w5490 & w14004;
assign w4000 = ~w4836 & ~a93;
assign w4001 = w9235 & ~w13441;
assign w4002 = w2228 & w3727;
assign w4003 = ~w3770 & w3374;
assign w4004 = w4233 & w9361;
assign w4005 = (w2697 & w685) | (w2697 & w7078) | (w685 & w7078);
assign w4006 = w4589 & w2207;
assign w4007 = (w12125 & ~w9298) | (w12125 & w11936) | (~w9298 & w11936);
assign w4008 = w5140 & ~w5664;
assign w4009 = w12915 & w10423;
assign w4010 = (w9305 & w6643) | (w9305 & w12712) | (w6643 & w12712);
assign w4011 = w7794 & w206;
assign w4012 = ~w9648 & w13765;
assign w4013 = w6750 & w3025;
assign w4014 = ~w607 & ~w5282;
assign w4015 = b53 & ~w7645;
assign w4016 = (w13210 & w1535) | (w13210 & w9347) | (w1535 & w9347);
assign w4017 = ~w309 & ~w11488;
assign w4018 = (w9254 & w10589) | (w9254 & w871) | (w10589 & w871);
assign w4019 = w11948 & w9807;
assign w4020 = ~w2392 & ~w1604;
assign w4021 = (~w8035 & ~w11583) | (~w8035 & w4839) | (~w11583 & w4839);
assign w4022 = w719 & ~w1540;
assign w4023 = w3128 & w4616;
assign w4024 = ~w5852 & w13857;
assign w4025 = w10146 & w11621;
assign w4026 = (~w9244 & ~w14280) | (~w9244 & w4229) | (~w14280 & w4229);
assign w4027 = (w10711 & w4582) | (w10711 & w1959) | (w4582 & w1959);
assign w4028 = (w4473 & w10778) | (w4473 & w13708) | (w10778 & w13708);
assign w4029 = ~w1379 & w1755;
assign w4030 = (~w1928 & w6656) | (~w1928 & w13331) | (w6656 & w13331);
assign w4031 = w5030 & w10721;
assign w4032 = ~w9342 & ~w8302;
assign w4033 = ~b29 & ~a29;
assign w4034 = (~w13521 & w12571) | (~w13521 & w10486) | (w12571 & w10486);
assign w4035 = (w9608 & w9830) | (w9608 & w11778) | (w9830 & w11778);
assign w4036 = w8871 & ~w3251;
assign w4037 = (w11385 & w2886) | (w11385 & w8054) | (w2886 & w8054);
assign w4038 = w11899 & ~w1979;
assign w4039 = ~w12798 & ~w13053;
assign w4040 = (w14048 & w5325) | (w14048 & w5222) | (w5325 & w5222);
assign w4041 = ~w13226 & w9710;
assign w4042 = w499 & w10993;
assign w4043 = ~w2218 & w1453;
assign w4044 = (~w5785 & w9139) | (~w5785 & w6994) | (w9139 & w6994);
assign w4045 = (~w11429 & w2964) | (~w11429 & w10982) | (w2964 & w10982);
assign w4046 = (w5863 & w9965) | (w5863 & w6524) | (w9965 & w6524);
assign w4047 = ~w3025 & w347;
assign w4048 = w11431 & w2962;
assign w4049 = (w11500 & w4512) | (w11500 & w1728) | (w4512 & w1728);
assign w4050 = w4572 & ~w10809;
assign w4051 = ~w8897 & w13755;
assign w4052 = ~w4858 | ~w3727;
assign w4053 = (~w3334 & ~w14355) | (~w3334 & w10033) | (~w14355 & w10033);
assign w4054 = w2432 & w12504;
assign w4055 = ~w9370 & w2367;
assign w4056 = ~w4607 & w3996;
assign w4057 = ~w8785 & w14462;
assign w4058 = w8624 & w7869;
assign w4059 = (w2922 & w13152) | (w2922 & w4201) | (w13152 & w4201);
assign w4060 = ~w614 & w8306;
assign w4061 = (w14215 & w1156) | (w14215 & w1933) | (w1156 & w1933);
assign w4062 = ~w6542 & ~w7722;
assign w4063 = (w6935 & w11191) | (w6935 & w9707) | (w11191 & w9707);
assign w4064 = w13919 & ~w13120;
assign w4065 = ~w4820 & w2879;
assign w4066 = (w10045 & w4387) | (w10045 & w4032) | (w4387 & w4032);
assign w4067 = (w713 & w3899) | (w713 & w6402) | (w3899 & w6402);
assign w4068 = w2872 & ~w9244;
assign w4069 = (~w8085 & w9608) | (~w8085 & w10133) | (w9608 & w10133);
assign w4070 = w10900 & ~w11134;
assign w4071 = ~b48 & ~a48;
assign w4072 = w11456 & ~w8296;
assign w4073 = (~w8183 & ~w12312) | (~w8183 & w10195) | (~w12312 & w10195);
assign w4074 = (w1513 & w2966) | (w1513 & w6096) | (w2966 & w6096);
assign w4075 = w6446 & ~w3904;
assign w4076 = (w6651 & ~w8285) | (w6651 & w9308) | (~w8285 & w9308);
assign w4077 = ~w13349 & w693;
assign w4078 = ~w9623 & ~w5741;
assign w4079 = ~w10590 & ~w5733;
assign w4080 = ~w12398 & ~w5692;
assign w4081 = w8234 & w2410;
assign w4082 = w4453 & w8580;
assign w4083 = ~w1171 & w5357;
assign w4084 = ~w5002 & w1692;
assign w4085 = w1540 & ~w827;
assign w4086 = ~w922 & ~w10178;
assign w4087 = w1572 & ~w9637;
assign w4088 = (w4233 & w12078) | (w4233 & w14484) | (w12078 & w14484);
assign w4089 = ~w703 & w2377;
assign w4090 = ~w8484 & w11582;
assign w4091 = (~w7637 & w9912) | (~w7637 & ~w9592) | (w9912 & ~w9592);
assign w4092 = ~w11215 & ~w1196;
assign w4093 = w9219 & ~w5208;
assign w4094 = w8347 & w13540;
assign w4095 = w2578 & w8817;
assign w4096 = (w6683 & w11429) | (w6683 & w9072) | (w11429 & w9072);
assign w4097 = w6368 & ~w2699;
assign w4098 = ~w13189 & w2732;
assign w4099 = w10326 & ~w13877;
assign w4100 = ~w12380 & w8799;
assign w4101 = ~w8769 & w8171;
assign w4102 = ~w2109 & ~w3573;
assign w4103 = ~w13071 & ~w7626;
assign w4104 = ~w14099 & ~w9310;
assign w4105 = ~w14137 & w13228;
assign w4106 = ~w12240 & w7338;
assign w4107 = w11085 & w9534;
assign w4108 = w1770 & w9724;
assign w4109 = w7968 & ~w676;
assign w4110 = ~w3914 & ~w2175;
assign w4111 = ~w979 & ~w8842;
assign w4112 = (w10685 & w8998) | (w10685 & ~w11185) | (w8998 & ~w11185);
assign w4113 = ~w6559 & w10125;
assign w4114 = ~w7076 & ~w9808;
assign w4115 = w9122 & ~w13293;
assign w4116 = ~w3632 & ~w8992;
assign w4117 = (w1692 & w3433) | (w1692 & w8237) | (w3433 & w8237);
assign w4118 = ~w2996 & w3727;
assign w4119 = w3550 & w7584;
assign w4120 = ~w43 & w1768;
assign w4121 = ~w498 & w9176;
assign w4122 = w2922 & ~w8769;
assign w4123 = (~w5952 & w2297) | (~w5952 & w8261) | (w2297 & w8261);
assign w4124 = w3550 & w7987;
assign w4125 = (~w7534 & w9578) | (~w7534 & w6535) | (w9578 & w6535);
assign w4126 = ~w932 & w10206;
assign w4127 = w3038 & w8085;
assign w4128 = (w11418 & w10344) | (w11418 & w11523) | (w10344 & w11523);
assign w4129 = ~w7365 & ~w1821;
assign w4130 = (w3957 & w5602) | (w3957 & ~w8675) | (w5602 & ~w8675);
assign w4131 = (w7457 & w2373) | (w7457 & w1175) | (w2373 & w1175);
assign w4132 = ~w12856 & w4062;
assign w4133 = ~w11462 & ~w4881;
assign w4134 = ~w8110 & ~w500;
assign w4135 = w3019 & ~w2933;
assign w4136 = (~w9170 & w10094) | (~w9170 & w8791) | (w10094 & w8791);
assign w4137 = ~w9626 & w7328;
assign w4138 = w1274 & w9817;
assign w4139 = ~w5294 & w13733;
assign w4140 = ~w11243 & w9840;
assign w4141 = (w2655 & w14242) | (w2655 & w3304) | (w14242 & w3304);
assign w4142 = ~w12108 & w11561;
assign w4143 = (~w3916 & w2867) | (~w3916 & w2696) | (w2867 & w2696);
assign w4144 = w13650 & ~w14643;
assign w4145 = ~w2872 & w8456;
assign w4146 = w4962 & ~w10013;
assign w4147 = w14015 & w11117;
assign w4148 = (~w13906 & w5968) | (~w13906 & w11825) | (w5968 & w11825);
assign w4149 = (w12406 & w4007) | (w12406 & w7644) | (w4007 & w7644);
assign w4150 = (~w10015 & w4686) | (~w10015 & w7378) | (w4686 & w7378);
assign w4151 = ~w10893 & w5557;
assign w4152 = w12901 & w11117;
assign w4153 = w11070 & ~w8268;
assign w4154 = (w6500 & w12783) | (w6500 & w11767) | (w12783 & w11767);
assign w4155 = ~w8520 & ~w4297;
assign w4156 = ~w8582 & ~w13365;
assign w4157 = ~w7205 & ~w8339;
assign w4158 = w12618 & w11596;
assign w4159 = b3 & a3;
assign w4160 = w1274 & w14486;
assign w4161 = (~w1260 & w12003) | (~w1260 & w10260) | (w12003 & w10260);
assign w4162 = w9537 & w6769;
assign w4163 = w7935 & ~w9336;
assign w4164 = w3751 & w8120;
assign w4165 = ~w11395 & ~w14417;
assign w4166 = w6485 & w6845;
assign w4167 = (~w6113 & w11159) | (~w6113 & w7710) | (w11159 & w7710);
assign w4168 = w9284 & w12642;
assign w4169 = ~w4863 & ~w2682;
assign w4170 = w11488 & ~w8827;
assign w4171 = ~w7537 & ~w3992;
assign w4172 = (~w11579 & w13343) | (~w11579 & w11911) | (w13343 & w11911);
assign w4173 = w4105 & ~w5785;
assign w4174 = w10966 & ~w6448;
assign w4175 = ~w13587 & w11267;
assign w4176 = ~w10860 & w8381;
assign w4177 = w9265 & w9658;
assign w4178 = ~w475 & w8713;
assign w4179 = ~w10245 & w1931;
assign w4180 = w4506 & w13395;
assign w4181 = (w2936 & w5060) | (w2936 & ~w14224) | (w5060 & ~w14224);
assign w4182 = ~w8171 & w10675;
assign w4183 = ~w8356 & ~w2950;
assign w4184 = ~w2125 & ~w42;
assign w4185 = w11500 & ~w10925;
assign w4186 = (~w7143 & ~w1476) | (~w7143 & w1641) | (~w1476 & w1641);
assign w4187 = w6042 & w4933;
assign w4188 = (w7295 & w4399) | (w7295 & w5506) | (w4399 & w5506);
assign w4189 = ~w11183 & ~w7178;
assign w4190 = ~w3019 & ~w10872;
assign w4191 = ~w2864 & w4203;
assign w4192 = w10013 & ~w8459;
assign w4193 = w12479 & ~w9090;
assign w4194 = w13056 & w762;
assign w4195 = w12090 & w2366;
assign w4196 = ~w4921 & w6617;
assign w4197 = ~w1166 & w5759;
assign w4198 = (w9226 & w11429) | (w9226 & w6131) | (w11429 & w6131);
assign w4199 = ~w5743 & ~w3427;
assign w4200 = ~w5845 & w7526;
assign w4201 = w4213 & w2922;
assign w4202 = ~w14038 & ~w4688;
assign w4203 = w3256 & w1015;
assign w4204 = ~w4881 & ~w8786;
assign w4205 = (~w14463 & w10634) | (~w14463 & w13811) | (w10634 & w13811);
assign w4206 = w7080 & ~w7423;
assign w4207 = ~w7572 & ~w3647;
assign w4208 = (w9831 & ~w630) | (w9831 & ~w2219) | (~w630 & ~w2219);
assign w4209 = ~w10997 & ~w10277;
assign w4210 = (~w14150 & w4421) | (~w14150 & w1448) | (w4421 & w1448);
assign w4211 = (~w7325 & w9250) | (~w7325 & w6039) | (w9250 & w6039);
assign w4212 = w13519 & ~w12915;
assign w4213 = ~w14285 & ~w219;
assign w4214 = w9323 & ~w8587;
assign w4215 = w5231 & w13895;
assign w4216 = ~w4268 & ~w557;
assign w4217 = (w13732 & w7867) | (w13732 & w8505) | (w7867 & w8505);
assign w4218 = (~w3611 & ~w14504) | (~w3611 & w7411) | (~w14504 & w7411);
assign w4219 = w3802 & ~w9162;
assign w4220 = ~w7219 & w1545;
assign w4221 = (~w597 & ~w10123) | (~w597 & w14264) | (~w10123 & w14264);
assign w4222 = ~w3730 & ~w7490;
assign w4223 = w13423 & ~w1221;
assign w4224 = (w3550 & w9615) | (w3550 & w1539) | (w9615 & w1539);
assign w4225 = ~w6302 & w11469;
assign w4226 = (w4787 & ~w1563) | (w4787 & w5873) | (~w1563 & w5873);
assign w4227 = (~w7180 & w9945) | (~w7180 & w14359) | (w9945 & w14359);
assign w4228 = ~w5559 & w6809;
assign w4229 = ~w12943 & ~w9244;
assign w4230 = (w6502 & ~w12271) | (w6502 & w13416) | (~w12271 & w13416);
assign w4231 = ~w3803 & ~w8768;
assign w4232 = ~w14412 & ~w4707;
assign w4233 = w1842 & w11500;
assign w4234 = (~w1862 & ~w5161) | (~w1862 & w10075) | (~w5161 & w10075);
assign w4235 = ~w2228 & ~w4458;
assign w4236 = (~w14028 & ~w4018) | (~w14028 & w888) | (~w4018 & w888);
assign w4237 = w1062 & ~w7889;
assign w4238 = (~w5385 & w7709) | (~w5385 & ~w9512) | (w7709 & ~w9512);
assign w4239 = (w6366 & w7585) | (w6366 & w9034) | (w7585 & w9034);
assign w4240 = ~w10256 & ~w1540;
assign w4241 = w3243 & ~w2995;
assign w4242 = (~w9412 & w11437) | (~w9412 & w3320) | (w11437 & w3320);
assign w4243 = w922 & w11159;
assign w4244 = (w968 & w12314) | (w968 & w1226) | (w12314 & w1226);
assign w4245 = ~w5425 & ~w14052;
assign w4246 = (~w3121 & ~w8900) | (~w3121 & w9241) | (~w8900 & w9241);
assign w4247 = (w10950 & w11967) | (w10950 & w13012) | (w11967 & w13012);
assign w4248 = (~w2410 & ~w6845) | (~w2410 & w10901) | (~w6845 & w10901);
assign w4249 = (~w2144 & w9238) | (~w2144 & w4443) | (w9238 & w4443);
assign w4250 = (~w9733 & w9364) | (~w9733 & w9403) | (w9364 & w9403);
assign w4251 = (~w2655 & w2139) | (~w2655 & w3728) | (w2139 & w3728);
assign w4252 = w9170 & w6266;
assign w4253 = w9679 & ~w8985;
assign w4254 = w10291 & ~w11838;
assign w4255 = w7645 & ~w5332;
assign w4256 = (~w11167 & w9563) | (~w11167 & w1698) | (w9563 & w1698);
assign w4257 = w4633 & w5591;
assign w4258 = ~w4836 & w12170;
assign w4259 = (~w12893 & w8742) | (~w12893 & w11759) | (w8742 & w11759);
assign w4260 = (w8127 & w6443) | (w8127 & w11413) | (w6443 & w11413);
assign w4261 = (w5860 & w2029) | (w5860 & w13390) | (w2029 & w13390);
assign w4262 = ~w9259 & w13038;
assign w4263 = ~w10334 & ~w6601;
assign w4264 = ~w13847 & ~w1026;
assign w4265 = w854 & w1718;
assign w4266 = ~w7914 & ~w3098;
assign w4267 = ~w9608 & w1431;
assign w4268 = ~w2296 & w12412;
assign w4269 = b89 & a89;
assign w4270 = ~b99 & ~a99;
assign w4271 = (w11500 & w10483) | (w11500 & w3966) | (w10483 & w3966);
assign w4272 = (w3885 & w11855) | (w3885 & w11853) | (w11855 & w11853);
assign w4273 = (w844 & w12053) | (w844 & w6086) | (w12053 & w6086);
assign w4274 = ~w3845 & w12859;
assign w4275 = (w6888 & ~w7347) | (w6888 & w10348) | (~w7347 & w10348);
assign w4276 = (~w5246 & w13388) | (~w5246 & w3805) | (w13388 & w3805);
assign w4277 = ~w9715 & w3564;
assign w4278 = ~w7760 & w8123;
assign w4279 = ~w5724 & w5236;
assign w4280 = ~w5707 & w890;
assign w4281 = (w13105 & ~w13585) | (w13105 & w2324) | (~w13585 & w2324);
assign w4282 = w10045 & w6861;
assign w4283 = w10378 & ~w2773;
assign w4284 = w3744 & w9212;
assign w4285 = w2617 & ~w1237;
assign w4286 = ~w13691 & w14540;
assign w4287 = ~w13713 & ~w14526;
assign w4288 = ~w9244 & ~w13445;
assign w4289 = (w5156 & w13837) | (w5156 & w2626) | (w13837 & w2626);
assign w4290 = (~w3742 & w5394) | (~w3742 & w11833) | (w5394 & w11833);
assign w4291 = ~w5005 & ~w622;
assign w4292 = w6951 & w11211;
assign w4293 = ~w4355 & w10710;
assign w4294 = ~w8488 & w5195;
assign w4295 = ~w13349 & w8492;
assign w4296 = w7244 & w2729;
assign w4297 = ~w13726 & w1743;
assign w4298 = ~w4780 & ~w5755;
assign w4299 = w9583 & w5593;
assign w4300 = (~w10522 & w11803) | (~w10522 & w9236) | (w11803 & w9236);
assign w4301 = ~w10497 & w6003;
assign w4302 = w13017 & ~w4805;
assign w4303 = ~w7336 & w7646;
assign w4304 = ~w5702 & w9585;
assign w4305 = w1758 & w325;
assign w4306 = w9123 & ~w13572;
assign w4307 = w8047 & ~w1997;
assign w4308 = (~w77 & w7782) | (~w77 & w9968) | (w7782 & w9968);
assign w4309 = w12846 & w7619;
assign w4310 = w6927 & w5490;
assign w4311 = (w12662 & w13152) | (w12662 & w9631) | (w13152 & w9631);
assign w4312 = b84 & a84;
assign w4313 = ~w13282 & ~w3823;
assign w4314 = ~w12572 & ~w9766;
assign w4315 = ~w12506 & ~w2701;
assign w4316 = w7776 & ~w12496;
assign w4317 = w227 & w4040;
assign w4318 = w9447 & ~w14296;
assign w4319 = w5243 & w10668;
assign w4320 = ~w2849 & w13499;
assign w4321 = w12721 & ~w4721;
assign w4322 = b99 & a99;
assign w4323 = ~w10909 & w12679;
assign w4324 = ~w8149 & ~w166;
assign w4325 = ~w407 & ~w4715;
assign w4326 = ~w3914 & w6542;
assign w4327 = (w6861 & ~w5325) | (w6861 & w6393) | (~w5325 & w6393);
assign w4328 = (w1607 & ~w3044) | (w1607 & w6887) | (~w3044 & w6887);
assign w4329 = w14302 & ~w2493;
assign w4330 = w4071 & ~w475;
assign w4331 = (~w11031 & w1609) | (~w11031 & w126) | (w1609 & w126);
assign w4332 = (w12569 & w8803) | (w12569 & ~w7527) | (w8803 & ~w7527);
assign w4333 = w8018 & w13435;
assign w4334 = (w922 & w913) | (w922 & w8709) | (w913 & w8709);
assign w4335 = ~w11150 & ~w8976;
assign w4336 = ~w8778 & ~w6975;
assign w4337 = w1643 & ~w7794;
assign w4338 = (~w9614 & w6345) | (~w9614 & w738) | (w6345 & w738);
assign w4339 = ~w8113 & w3563;
assign w4340 = w6391 & w7924;
assign w4341 = ~w7447 & ~w4515;
assign w4342 = (~w13375 & ~w5498) | (~w13375 & ~w3266) | (~w5498 & ~w3266);
assign w4343 = w10116 & w12543;
assign w4344 = (w12209 & w12293) | (w12209 & w9877) | (w12293 & w9877);
assign w4345 = ~w2410 & ~w9087;
assign w4346 = (w8602 & ~w1543) | (w8602 & w14119) | (~w1543 & w14119);
assign w4347 = (w7062 & ~w10630) | (w7062 & w819) | (~w10630 & w819);
assign w4348 = (~w14629 & ~w3181) | (~w14629 & w11288) | (~w3181 & w11288);
assign w4349 = w8120 & w13011;
assign w4350 = ~w12121 & w12398;
assign w4351 = (~w5867 & w3317) | (~w5867 & w5964) | (w3317 & w5964);
assign w4352 = (~w13183 & w11877) | (~w13183 & w7720) | (w11877 & w7720);
assign w4353 = (~w2372 & w7136) | (~w2372 & w8575) | (w7136 & w8575);
assign w4354 = ~w12575 & w3906;
assign w4355 = (w3121 & w1831) | (w3121 & w10253) | (w1831 & w10253);
assign w4356 = (w13587 & w5225) | (w13587 & w2338) | (w5225 & w2338);
assign w4357 = w11287 & w11977;
assign w4358 = w11041 & ~w322;
assign w4359 = ~b81 & ~a81;
assign w4360 = w5243 & w8977;
assign w4361 = ~w9820 & ~w3339;
assign w4362 = (~w6777 & w9879) | (~w6777 & w10149) | (w9879 & w10149);
assign w4363 = ~w4388 & ~w416;
assign w4364 = w13224 & ~w3399;
assign w4365 = w11280 & ~w2813;
assign w4366 = ~w4607 & w13248;
assign w4367 = ~w2498 & w9425;
assign w4368 = ~w2858 & ~w8992;
assign w4369 = (~w4050 & w5999) | (~w4050 & w6767) | (w5999 & w6767);
assign w4370 = (w1416 & w6088) | (w1416 & w8458) | (w6088 & w8458);
assign w4371 = ~w3722 & ~w10603;
assign w4372 = w7132 & w7951;
assign w4373 = ~w5816 & ~w13082;
assign w4374 = w5969 | ~w2870;
assign w4375 = ~w2680 & ~w1199;
assign w4376 = w5693 & w12614;
assign w4377 = (w11138 & w6209) | (w11138 & w589) | (w6209 & w589);
assign w4378 = w719 & w1062;
assign w4379 = w4855 & w2589;
assign w4380 = ~w7040 & w2283;
assign w4381 = ~w12642 & w4033;
assign w4382 = ~w13222 & w2425;
assign w4383 = w10116 & w5767;
assign w4384 = ~w13714 & w12309;
assign w4385 = ~w14302 & ~w13462;
assign w4386 = w11759 & ~w10926;
assign w4387 = ~w13531 & w10045;
assign w4388 = w13531 & ~w9541;
assign w4389 = (~w9932 & w9608) | (~w9932 & w12093) | (w9608 & w12093);
assign w4390 = ~w13300 & ~w608;
assign w4391 = (w2798 & w413) | (w2798 & ~w9755) | (w413 & ~w9755);
assign w4392 = w14417 & ~w1536;
assign w4393 = (w12460 & w11578) | (w12460 & w8791) | (w11578 & w8791);
assign w4394 = w11959 & w11500;
assign w4395 = w2680 & w6845;
assign w4396 = (~w3963 & w110) | (~w3963 & w11940) | (w110 & w11940);
assign w4397 = w10676 & w2410;
assign w4398 = ~w1709 & ~w12668;
assign w4399 = ~w2605 & w7295;
assign w4400 = ~w1840 & w542;
assign w4401 = ~w9788 & ~w6716;
assign w4402 = (w1949 & w12842) | (w1949 & w7583) | (w12842 & w7583);
assign w4403 = ~w1563 & ~w10702;
assign w4404 = w11161 | w1564;
assign w4405 = w11500 & ~w622;
assign w4406 = w9574 & w7507;
assign w4407 = (~w142 & ~w11031) | (~w142 & w6872) | (~w11031 & w6872);
assign w4408 = w11041 & ~w14616;
assign w4409 = w9345 & w9340;
assign w4410 = (w9541 & w5573) | (w9541 & w6386) | (w5573 & w6386);
assign w4411 = (w10290 & ~w9715) | (w10290 & w534) | (~w9715 & w534);
assign w4412 = (~w4287 & w183) | (~w4287 & w10335) | (w183 & w10335);
assign w4413 = w2362 & w6293;
assign w4414 = ~w13282 & ~w1027;
assign w4415 = w4756 & w3289;
assign w4416 = (w12776 & w13102) | (w12776 & w2141) | (w13102 & w2141);
assign w4417 = ~w2585 & ~w10524;
assign w4418 = ~w14178 & w8367;
assign w4419 = w4283 & w3997;
assign w4420 = ~w7762 & ~w12614;
assign w4421 = ~w12591 & ~w109;
assign w4422 = ~w6232 & ~w2327;
assign w4423 = w3632 & ~w4127;
assign w4424 = ~w10629 & w2493;
assign w4425 = ~w6281 & ~w5036;
assign w4426 = (w2169 & w1613) | (w2169 & w12702) | (w1613 & w12702);
assign w4427 = w3277 & w4405;
assign w4428 = ~w7376 & ~w13531;
assign w4429 = (w829 & w254) | (w829 & w6523) | (w254 & w6523);
assign w4430 = (w1678 & w4965) | (w1678 & ~w10774) | (w4965 & ~w10774);
assign w4431 = (~w6190 & w4848) | (~w6190 & w8060) | (w4848 & w8060);
assign w4432 = w11759 & w3537;
assign w4433 = w7489 & w10686;
assign w4434 = w2954 & w3001;
assign w4435 = w14096 | w717;
assign w4436 = (~w14528 & w12595) | (~w14528 & w7209) | (w12595 & w7209);
assign w4437 = ~w11196 & ~w10289;
assign w4438 = (w6299 & w2102) | (w6299 & w11331) | (w2102 & w11331);
assign w4439 = ~w1563 & ~w11732;
assign w4440 = w7131 & w11393;
assign w4441 = ~w13854 & ~w13620;
assign w4442 = w2723 & ~w13798;
assign w4443 = (~w9921 & ~w4032) | (~w9921 & w9238) | (~w4032 & w9238);
assign w4444 = w8929 & ~w5936;
assign w4445 = w6584 & w7914;
assign w4446 = ~w1609 & w7468;
assign w4447 = w9952 & w2096;
assign w4448 = (~w1260 & w1692) | (~w1260 & w14584) | (w1692 & w14584);
assign w4449 = w12987 & w752;
assign w4450 = w14512 & ~w3019;
assign w4451 = (w514 & w14044) | (w514 & w9521) | (w14044 & w9521);
assign w4452 = w3175 & ~w7196;
assign w4453 = ~w7022 & ~w12315;
assign w4454 = (w11979 & w12289) | (w11979 & w14123) | (w12289 & w14123);
assign w4455 = w4213 & w10317;
assign w4456 = (w10172 & w9892) | (w10172 & w9034) | (w9892 & w9034);
assign w4457 = w7811 & ~w2850;
assign w4458 = ~w13297 & ~w13900;
assign w4459 = w10 & w735;
assign w4460 = w10853 & w8900;
assign w4461 = ~w9134 & w13444;
assign w4462 = ~w5521 & ~w11454;
assign w4463 = w255 | w3753;
assign w4464 = ~w4930 & w11208;
assign w4465 = ~w2115 & w14217;
assign w4466 = (w13713 & ~w10143) | (w13713 & w3289) | (~w10143 & w3289);
assign w4467 = ~w12065 & ~w11395;
assign w4468 = (w5449 & w14422) | (w5449 & w946) | (w14422 & w946);
assign w4469 = w6467 & ~w12905;
assign w4470 = (~w4017 & w13282) | (~w4017 & w1819) | (w13282 & w1819);
assign w4471 = w7621 & w14656;
assign w4472 = w1114 & w1007;
assign w4473 = (~w3508 & ~w6301) | (~w3508 & w11493) | (~w6301 & w11493);
assign w4474 = ~w2844 & w13008;
assign w4475 = (~w4670 & w7907) | (~w4670 & w6715) | (w7907 & w6715);
assign w4476 = (w12409 & w4852) | (w12409 & w10220) | (w4852 & w10220);
assign w4477 = ~w9788 & ~w13839;
assign w4478 = ~w7963 & ~w11955;
assign w4479 = (w13871 & w8185) | (w13871 & w731) | (w8185 & w731);
assign w4480 = ~w3747 & ~w11154;
assign w4481 = (~w10116 & ~w3671) | (~w10116 & w10301) | (~w3671 & w10301);
assign w4482 = (w13508 & w10464) | (w13508 & w3634) | (w10464 & w3634);
assign w4483 = b26 & a26;
assign w4484 = ~w9822 & ~w7873;
assign w4485 = (~w5050 & w5178) | (~w5050 & w8584) | (w5178 & w8584);
assign w4486 = ~w13832 & ~w3325;
assign w4487 = ~w2509 & ~w5644;
assign w4488 = w1802 & ~w8280;
assign w4489 = ~w11429 & w9196;
assign w4490 = (w4018 & w12651) | (w4018 & w1320) | (w12651 & w1320);
assign w4491 = w7469 & ~w14110;
assign w4492 = w12271 & ~w11228;
assign w4493 = (w12868 & w4921) | (w12868 & w1071) | (w4921 & w1071);
assign w4494 = ~w5683 & w6413;
assign w4495 = w13161 & ~w6686;
assign w4496 = w6064 & w4458;
assign w4497 = ~w12459 & ~w12165;
assign w4498 = ~w5288 & w3427;
assign w4499 = ~w9012 & w1602;
assign w4500 = ~w14526 & ~w6952;
assign w4501 = ~w7349 & ~w8819;
assign w4502 = w13929 & ~w7151;
assign w4503 = ~w473 & ~w11905;
assign w4504 = w13126 & w5825;
assign w4505 = ~w3203 & w427;
assign w4506 = w634 & ~w11808;
assign w4507 = ~w9608 & w6055;
assign w4508 = (w5676 & w9552) | (w5676 & w2271) | (w9552 & w2271);
assign w4509 = w706 & w8396;
assign w4510 = (w5186 & w4194) | (w5186 & ~w6507) | (w4194 & ~w6507);
assign w4511 = (~w7296 & w1238) | (~w7296 & w4392) | (w1238 & w4392);
assign w4512 = w5463 & ~w13790;
assign w4513 = w13728 & w1618;
assign w4514 = w922 & ~w10507;
assign w4515 = ~b17 & ~a17;
assign w4516 = (~w3215 & w4050) | (~w3215 & w12792) | (w4050 & w12792);
assign w4517 = ~w11570 & ~w11772;
assign w4518 = (w7787 & w14274) | (w7787 & w6919) | (w14274 & w6919);
assign w4519 = w9989 & w13611;
assign w4520 = ~w8626 & w6219;
assign w4521 = ~w3593 & w12647;
assign w4522 = ~w4688 & ~w7833;
assign w4523 = (~w142 & ~w12460) | (~w142 & w6872) | (~w12460 & w6872);
assign w4524 = (w6714 & w7333) | (w6714 & w12892) | (w7333 & w12892);
assign w4525 = (w12569 & w6230) | (w12569 & w1217) | (w6230 & w1217);
assign w4526 = w4252 & w6266;
assign w4527 = (w8937 & w8709) | (w8937 & w4334) | (w8709 & w4334);
assign w4528 = w6328 & ~w7308;
assign w4529 = (~w6186 & w5204) | (~w6186 & w3029) | (w5204 & w3029);
assign w4530 = ~w7390 & ~w2662;
assign w4531 = (~w5291 & ~w13084) | (~w5291 & w8928) | (~w13084 & w8928);
assign w4532 = ~w7141 & ~w13027;
assign w4533 = w8975 & ~w2791;
assign w4534 = w5490 & ~w686;
assign w4535 = w14302 & ~w3435;
assign w4536 = w14342 & w4855;
assign w4537 = w13953 & ~w9880;
assign w4538 = ~w5373 & w1061;
assign w4539 = ~w10343 & w3819;
assign w4540 = (w6423 & w1249) | (w6423 & w2532) | (w1249 & w2532);
assign w4541 = (~w5852 & w5804) | (~w5852 & w10389) | (w5804 & w10389);
assign w4542 = w10949 & w12165;
assign w4543 = w6953 & w3436;
assign w4544 = w8339 & ~w10573;
assign w4545 = (w5070 & w11723) | (w5070 & w8607) | (w11723 & w8607);
assign w4546 = ~w6026 & w8386;
assign w4547 = ~w11952 & w8177;
assign w4548 = ~w607 & w7670;
assign w4549 = ~w5522 & ~w1540;
assign w4550 = ~w10155 & w13605;
assign w4551 = w2063 & ~w13569;
assign w4552 = ~w6868 & ~w13856;
assign w4553 = w7681 & ~w5282;
assign w4554 = ~w183 & w13713;
assign w4555 = w12385 & ~w4353;
assign w4556 = ~w9805 & ~w13077;
assign w4557 = ~w7982 & ~w7550;
assign w4558 = ~w9569 & ~w9304;
assign w4559 = w2137 & w10087;
assign w4560 = w8183 & w6689;
assign w4561 = w4151 & w3030;
assign w4562 = ~w5105 & w4389;
assign w4563 = ~w3803 & ~w8459;
assign w4564 = ~w2315 & ~w7280;
assign w4565 = (w2493 & ~w3823) | (w2493 & w1787) | (~w3823 & w1787);
assign w4566 = (~w13587 & w2638) | (~w13587 & w12981) | (w2638 & w12981);
assign w4567 = ~w13222 & ~w13873;
assign w4568 = (w3795 & w7945) | (w3795 & w10593) | (w7945 & w10593);
assign w4569 = w14482 & w525;
assign w4570 = (w1503 & w3261) | (w1503 & w7341) | (w3261 & w7341);
assign w4571 = w13733 & ~w1692;
assign w4572 = ~w11342 & w11291;
assign w4573 = ~w9623 & w7633;
assign w4574 = w2387 & w813;
assign w4575 = w3550 & w366;
assign w4576 = (w10915 & w13327) | (w10915 & w2424) | (w13327 & w2424);
assign w4577 = w5788 & w1260;
assign w4578 = (w13595 & w3818) | (w13595 & ~w2663) | (w3818 & ~w2663);
assign w4579 = (w8010 & w8519) | (w8010 & ~w14455) | (w8519 & ~w14455);
assign w4580 = ~w9921 & ~w3098;
assign w4581 = (w1498 & w1855) | (w1498 & w4299) | (w1855 & w4299);
assign w4582 = ~w195 & w11389;
assign w4583 = w11458 & ~w2303;
assign w4584 = (~w14512 & w10483) | (~w14512 & w10363) | (w10483 & w10363);
assign w4585 = w8389 & ~w6045;
assign w4586 = w10477 & w12614;
assign w4587 = ~w2387 & ~w1172;
assign w4588 = w3671 & ~w5255;
assign w4589 = w6697 & w8843;
assign w4590 = (~w10926 & ~w8659) | (~w10926 & w14417) | (~w8659 & w14417);
assign w4591 = w3550 & w8828;
assign w4592 = (~w3460 & w55) | (~w3460 & w9098) | (w55 & w9098);
assign w4593 = (w2485 & w6893) | (w2485 & w5785) | (w6893 & w5785);
assign w4594 = (~w14564 & w6754) | (~w14564 & w7039) | (w6754 & w7039);
assign w4595 = w10916 & ~w8389;
assign w4596 = w10676 & w40;
assign w4597 = (w9200 & w12499) | (w9200 & w10673) | (w12499 & w10673);
assign w4598 = w8000 & w11622;
assign w4599 = w13635 & w11309;
assign w4600 = ~w10334 & ~w13723;
assign w4601 = (~w14395 & w10435) | (~w14395 & w8278) | (w10435 & w8278);
assign w4602 = w8620 & ~w555;
assign w4603 = (~w11973 & w3620) | (~w11973 & w11963) | (w3620 & w11963);
assign w4604 = w9623 & ~w11117;
assign w4605 = ~w4948 & ~w13778;
assign w4606 = w6716 & w2144;
assign w4607 = (~w12338 & w9012) | (~w12338 & w3064) | (w9012 & w3064);
assign w4608 = (w9305 & w317) | (w9305 & w9771) | (w317 & w9771);
assign w4609 = w1274 & ~w10301;
assign w4610 = w4667 & ~w3044;
assign w4611 = ~w759 & ~w11260;
assign w4612 = ~w9262 & ~w3821;
assign w4613 = w3336 | w1344;
assign w4614 = (~w9364 & w5169) | (~w9364 & w9441) | (w5169 & w9441);
assign w4615 = ~w4154 & w1122;
assign w4616 = ~w6750 & w8512;
assign w4617 = w12216 & ~w12642;
assign w4618 = ~w14614 & w5590;
assign w4619 = ~w12240 & w884;
assign w4620 = (w12893 & w2962) | (w12893 & w5424) | (w2962 & w5424);
assign w4621 = ~w14664 & w1089;
assign w4622 = w10483 & ~w11299;
assign w4623 = w3550 & w2376;
assign w4624 = (w1949 & w7988) | (w1949 & w11162) | (w7988 & w11162);
assign w4625 = ~w2915 & w14210;
assign w4626 = w7392 & w39;
assign w4627 = ~w8035 & ~w6935;
assign w4628 = ~w11980 & ~w7297;
assign w4629 = w10906 & ~w7335;
assign w4630 = ~w3409 & ~w850;
assign w4631 = ~w607 & ~w2729;
assign w4632 = (~w12464 & ~w213) | (~w12464 & w5037) | (~w213 & w5037);
assign w4633 = ~w12926 & w11927;
assign w4634 = ~w5604 & w7768;
assign w4635 = ~w7782 & w8838;
assign w4636 = w791 & w5983;
assign w4637 = ~w13222 & w40;
assign w4638 = w13206 & w9921;
assign w4639 = ~w13421 & ~w1502;
assign w4640 = ~w1563 & w10225;
assign w4641 = w5522 & w646;
assign w4642 = w3550 & w13913;
assign w4643 = w1498 & w4127;
assign w4644 = ~w4158 & w5986;
assign w4645 = w2433 & ~w2701;
assign w4646 = w813 & w4706;
assign w4647 = w9970 & w11632;
assign w4648 = ~w71 & w12906;
assign w4649 = ~w3885 & w13839;
assign w4650 = w9321 & ~w12960;
assign w4651 = ~w12464 & w9608;
assign w4652 = w4189 & ~w2421;
assign w4653 = w5127 & ~w11975;
assign w4654 = (~w8483 & w11262) | (~w8483 & w837) | (w11262 & w837);
assign w4655 = w7111 & w5870;
assign w4656 = ~w5482 & ~w6171;
assign w4657 = ~w4620 & w2610;
assign w4658 = w6219 & w4503;
assign w4659 = w8790 & w10944;
assign w4660 = ~w13587 & w1012;
assign w4661 = w10676 & w3906;
assign w4662 = (w10625 & w11149) | (w10625 & ~w5895) | (w11149 & ~w5895);
assign w4663 = (~w3717 & w1387) | (~w3717 & w1124) | (w1387 & w1124);
assign w4664 = (~w2270 & ~w14542) | (~w2270 & w3885) | (~w14542 & w3885);
assign w4665 = (w3714 & w4921) | (w3714 & w8547) | (w4921 & w8547);
assign w4666 = w12294 & w13978;
assign w4667 = w12483 & w9932;
assign w4668 = ~w3958 & w2171;
assign w4669 = w9788 & w11861;
assign w4670 = ~w13843 & w2195;
assign w4671 = ~w5556 & ~w894;
assign w4672 = ~w4050 & w1345;
assign w4673 = (~w11738 & ~w6229) | (~w11738 & w11623) | (~w6229 & w11623);
assign w4674 = w7267 & w2829;
assign w4675 = (w14472 & w5671) | (w14472 & ~w14534) | (w5671 & ~w14534);
assign w4676 = ~w3938 & w10074;
assign w4677 = (~w8100 & w7799) | (~w8100 & ~w4218) | (w7799 & ~w4218);
assign w4678 = ~w14275 & ~w5794;
assign w4679 = (~w10433 & w9106) | (~w10433 & w7250) | (w9106 & w7250);
assign w4680 = ~w4700 & w7670;
assign w4681 = (w6267 & w2953) | (w6267 & w8580) | (w2953 & w8580);
assign w4682 = (w12589 & w9081) | (w12589 & ~w112) | (w9081 & ~w112);
assign w4683 = (w5532 & w818) | (w5532 & ~w14271) | (w818 & ~w14271);
assign w4684 = ~w4359 & w13772;
assign w4685 = (w5732 & w12499) | (w5732 & w7658) | (w12499 & w7658);
assign w4686 = w1570 & ~w2698;
assign w4687 = ~w14302 & w6716;
assign w4688 = b13 & a13;
assign w4689 = w14278 & ~w10432;
assign w4690 = (w4127 & ~w3209) | (w4127 & w11716) | (~w3209 & w11716);
assign w4691 = ~w8108 & ~w3018;
assign w4692 = (w12344 & w5161) | (w12344 & w14551) | (w5161 & w14551);
assign w4693 = ~w4700 & w10699;
assign w4694 = (w1849 & w4112) | (w1849 & w9662) | (w4112 & w9662);
assign w4695 = w805 & w10210;
assign w4696 = (w6410 & w1313) | (w6410 & w8407) | (w1313 & w8407);
assign w4697 = w7154 & w1062;
assign w4698 = w10136 | ~w7999;
assign w4699 = ~w10930 & ~w2984;
assign w4700 = ~b96 & ~a96;
assign w4701 = w10847 & w13872;
assign w4702 = ~w3914 & w473;
assign w4703 = (w3364 & w5877) | (w3364 & ~w9709) | (w5877 & ~w9709);
assign w4704 = w9172 & w8353;
assign w4705 = ~w6511 & ~w11888;
assign w4706 = w1096 & ~w10675;
assign w4707 = b6 & a6;
assign w4708 = (w1498 & w2964) | (w1498 & ~w8992) | (w2964 & ~w8992);
assign w4709 = (w9512 & ~w7482) | (w9512 & w9668) | (~w7482 & w9668);
assign w4710 = w13222 & ~w7437;
assign w4711 = ~w14294 & ~w9216;
assign w4712 = w5522 & ~w3904;
assign w4713 = (w10872 & w3122) | (w10872 & w12518) | (w3122 & w12518);
assign w4714 = ~w6605 & w10009;
assign w4715 = w646 & w13508;
assign w4716 = w7794 & w213;
assign w4717 = w1150 & w629;
assign w4718 = ~w6190 & w5282;
assign w4719 = w3550 & w9189;
assign w4720 = (~w10590 & w2470) | (~w10590 & w3209) | (w2470 & w3209);
assign w4721 = (w7428 & ~w9475) | (w7428 & w7364) | (~w9475 & w7364);
assign w4722 = w4339 & ~w3885;
assign w4723 = ~w11703 & w10058;
assign w4724 = ~w14620 & ~w9964;
assign w4725 = (~w11052 & ~w6138) | (~w11052 & w1747) | (~w6138 & w1747);
assign w4726 = (~w9012 & w6156) | (~w9012 & w2892) | (w6156 & w2892);
assign w4727 = ~w12121 & ~w3526;
assign w4728 = (w8584 & ~w13282) | (w8584 & w2171) | (~w13282 & w2171);
assign w4729 = (~w6301 & w2175) | (~w6301 & w6613) | (w2175 & w6613);
assign w4730 = w4587 & w11500;
assign w4731 = ~w1390 & ~w5244;
assign w4732 = ~w3219 & w12460;
assign w4733 = ~w4744 & ~w4255;
assign w4734 = w7070 & w12425;
assign w4735 = (~w6716 & ~w9715) | (~w6716 & w7914) | (~w9715 & w7914);
assign w4736 = (~w3550 & w13745) | (~w3550 & w14016) | (w13745 & w14016);
assign w4737 = w1521 & w11661;
assign w4738 = w6716 & w9921;
assign w4739 = ~b53 & ~w12204;
assign w4740 = (~w13469 & w6688) | (~w13469 & w10934) | (w6688 & w10934);
assign w4741 = ~w8120 & w13227;
assign w4742 = w5865 & w4491;
assign w4743 = ~w7483 & ~w12377;
assign w4744 = ~w254 & w6764;
assign w4745 = (~w13526 & w2998) | (~w13526 & ~w3750) | (w2998 & ~w3750);
assign w4746 = w8737 & w490;
assign w4747 = (~w11915 & w9773) | (~w11915 & w2600) | (w9773 & w2600);
assign w4748 = (w12224 & w14282) | (w12224 & w9029) | (w14282 & w9029);
assign w4749 = ~w5231 & w8120;
assign w4750 = (~w3734 & w922) | (~w3734 & w620) | (w922 & w620);
assign w4751 = w3550 & w5531;
assign w4752 = w7719 & w10692;
assign w4753 = ~w1129 & w9417;
assign w4754 = ~w2362 & ~w7515;
assign w4755 = w5135 & w8870;
assign w4756 = w5575 & ~w12825;
assign w4757 = w11041 & w13566;
assign w4758 = ~w6764 & ~w724;
assign w4759 = (~w3537 & w263) | (~w3537 & w10387) | (w263 & w10387);
assign w4760 = ~w2097 & w6403;
assign w4761 = ~w5741 & ~w1540;
assign w4762 = w13459 & w14519;
assign w4763 = w5936 & w2928;
assign w4764 = ~w10334 & ~w9823;
assign w4765 = (~w13587 & w12098) | (~w13587 & w524) | (w12098 & w524);
assign w4766 = ~w13282 & ~w6981;
assign w4767 = (~w3549 & w9887) | (~w3549 & w11100) | (w9887 & w11100);
assign w4768 = (w8778 & w12597) | (w8778 & w4188) | (w12597 & w4188);
assign w4769 = w5060 | w2936;
assign w4770 = ~w4783 | ~w9215;
assign w4771 = (w6873 & w9217) | (w6873 & w8614) | (w9217 & w8614);
assign w4772 = (w13576 & w9745) | (w13576 & w13024) | (w9745 & w13024);
assign w4773 = ~w6151 & w14512;
assign w4774 = (~w6700 & w6192) | (~w6700 & ~w7526) | (w6192 & ~w7526);
assign w4775 = (w9027 & w7917) | (w9027 & w11413) | (w7917 & w11413);
assign w4776 = (w2485 & w6893) | (w2485 & ~w9139) | (w6893 & ~w9139);
assign w4777 = ~w2159 & w14504;
assign w4778 = (w167 & w227) | (w167 & w2463) | (w227 & w2463);
assign w4779 = (w852 & w6845) | (w852 & w8957) | (w6845 & w8957);
assign w4780 = w7376 & w1140;
assign w4781 = ~w8111 & w10736;
assign w4782 = ~w14187 & w11719;
assign w4783 = (w5744 & w13172) | (w5744 & ~w3885) | (w13172 & ~w3885);
assign w4784 = (~w10923 & w8150) | (~w10923 & w5868) | (w8150 & w5868);
assign w4785 = (w7273 & w6416) | (w7273 & w246) | (w6416 & w246);
assign w4786 = ~w10669 & ~w7630;
assign w4787 = w14395 & w7962;
assign w4788 = ~w12519 & w2649;
assign w4789 = ~w1563 & w4288;
assign w4790 = w4405 & ~w14124;
assign w4791 = w12464 & ~w11117;
assign w4792 = (~w7782 & w5226) | (~w7782 & w12187) | (w5226 & w12187);
assign w4793 = w9912 & ~w2789;
assign w4794 = (~w5002 & w4512) | (~w5002 & w2944) | (w4512 & w2944);
assign w4795 = ~w7482 & w5793;
assign w4796 = w3038 & w12135;
assign w4797 = w3121 & w4216;
assign w4798 = ~w1563 & ~w2317;
assign w4799 = w9034 | w8228;
assign w4800 = w9679 & w10182;
assign w4801 = (w5860 & w13152) | (w5860 & w8310) | (w13152 & w8310);
assign w4802 = (w6107 & w1473) | (w6107 & ~w13292) | (w1473 & ~w13292);
assign w4803 = ~w14007 & w5735;
assign w4804 = ~w2357 & w10306;
assign w4805 = w2463 & w6958;
assign w4806 = w7317 & w8285;
assign w4807 = (w3531 & w223) | (w3531 & w1213) | (w223 & w1213);
assign w4808 = ~w12662 & w7926;
assign w4809 = (~w9608 & w11349) | (~w9608 & w2613) | (w11349 & w2613);
assign w4810 = ~w5001 & ~w7521;
assign w4811 = ~w9719 & w8335;
assign w4812 = ~w8694 & w12407;
assign w4813 = w14585 & w6671;
assign w4814 = (w894 & w12499) | (w894 & w8557) | (w12499 & w8557);
assign w4815 = ~w3450 & w3688;
assign w4816 = (w13987 & w13572) | (w13987 & w14035) | (w13572 & w14035);
assign w4817 = ~w8225 & ~w9032;
assign w4818 = (w2165 & w2342) | (w2165 & w10810) | (w2342 & w10810);
assign w4819 = (w4318 & w849) | (w4318 & w14171) | (w849 & w14171);
assign w4820 = ~w7580 & w4793;
assign w4821 = (w4607 & w5806) | (w4607 & w4136) | (w5806 & w4136);
assign w4822 = w10592 & ~w2284;
assign w4823 = w10704 & w10708;
assign w4824 = w13526 & ~w5845;
assign w4825 = w10689 & w10704;
assign w4826 = ~w12121 & w2425;
assign w4827 = (w9766 & w4438) | (w9766 & w7029) | (w4438 & w7029);
assign w4828 = (w4855 & w14342) | (w4855 & ~w6750) | (w14342 & ~w6750);
assign w4829 = ~w6033 & ~w10118;
assign w4830 = (w13580 & w9991) | (w13580 & w7601) | (w9991 & w7601);
assign w4831 = ~w3885 & w12460;
assign w4832 = w7620 & w11549;
assign w4833 = ~w5058 & w1720;
assign w4834 = w13328 & ~w2492;
assign w4835 = ~w6442 & w690;
assign w4836 = ~w2658 & ~w2130;
assign w4837 = ~w183 & w1821;
assign w4838 = w5535 & ~w12882;
assign w4839 = w3851 & ~w8035;
assign w4840 = ~w7259 & ~w10187;
assign w4841 = w4032 & w473;
assign w4842 = ~w14664 & w4736;
assign w4843 = (~w12574 & w1356) | (~w12574 & w5849) | (w1356 & w5849);
assign w4844 = (w3550 & w6914) | (w3550 & w11125) | (w6914 & w11125);
assign w4845 = (~w4033 & w690) | (~w4033 & w11000) | (w690 & w11000);
assign w4846 = (~w10590 & ~w9748) | (~w10590 & w2470) | (~w9748 & w2470);
assign w4847 = w1274 & w10116;
assign w4848 = ~w10757 & ~w10949;
assign w4849 = w13445 & w9156;
assign w4850 = (w3289 & ~w5238) | (w3289 & w12396) | (~w5238 & w12396);
assign w4851 = w4563 & ~w10781;
assign w4852 = (~w10884 & w1377) | (~w10884 & w11724) | (w1377 & w11724);
assign w4853 = (w12776 & w13482) | (w12776 & w9736) | (w13482 & w9736);
assign w4854 = w13411 & ~w385;
assign w4855 = w4467 & w14417;
assign w4856 = ~w9482 & ~w11764;
assign w4857 = ~w533 & ~w6500;
assign w4858 = w14614 & w3727;
assign w4859 = ~w7889 & ~w9211;
assign w4860 = w8663 & ~w6152;
assign w4861 = ~w3883 & w4279;
assign w4862 = (w7376 & w1569) | (w7376 & w892) | (w1569 & w892);
assign w4863 = ~w13839 & ~w9861;
assign w4864 = (~w6795 & w12499) | (~w6795 & w5838) | (w12499 & w5838);
assign w4865 = w5948 & ~w5761;
assign w4866 = ~w8934 & w9503;
assign w4867 = (~w3478 & w12957) | (~w3478 & w8209) | (w12957 & w8209);
assign w4868 = w8239 & w10141;
assign w4869 = (~w1362 & w6419) | (~w1362 & w5152) | (w6419 & w5152);
assign w4870 = w10398 & w3606;
assign w4871 = ~w9747 & w9138;
assign w4872 = ~w11038 & w5390;
assign w4873 = w12833 & w6351;
assign w4874 = w9454 & w112;
assign w4875 = ~w9608 & w8316;
assign w4876 = (w758 & w1245) | (w758 & w13107) | (w1245 & w13107);
assign w4877 = (~w6230 & w7688) | (~w6230 & w1468) | (w7688 & w1468);
assign w4878 = (w1658 & ~w6929) | (w1658 & w7610) | (~w6929 & w7610);
assign w4879 = ~w11500 & w10;
assign w4880 = ~w11025 & ~w9005;
assign w4881 = b41 & a41;
assign w4882 = ~w581 & w2668;
assign w4883 = w14640 & ~w13323;
assign w4884 = w5761 & w4458;
assign w4885 = ~w5412 & ~w4134;
assign w4886 = (w4041 & w6635) | (w4041 & w11090) | (w6635 & w11090);
assign w4887 = ~w4810 & ~w7371;
assign w4888 = w13594 & ~w7640;
assign w4889 = (w7812 & ~w4569) | (w7812 & w7934) | (~w4569 & w7934);
assign w4890 = w880 & w7856;
assign w4891 = ~w12065 & w683;
assign w4892 = ~w11200 & ~w81;
assign w4893 = ~w40 & ~w1007;
assign w4894 = w11264 & w9001;
assign w4895 = ~w10590 & ~w2423;
assign w4896 = w9715 & w3025;
assign w4897 = (w11606 & w2605) | (w11606 & ~w8133) | (w2605 & ~w8133);
assign w4898 = ~w4570 & w14612;
assign w4899 = (w13685 & w12423) | (w13685 & w8514) | (w12423 & w8514);
assign w4900 = ~w1111 & w2521;
assign w4901 = ~w4992 & w9716;
assign w4902 = w4881 & w2941;
assign w4903 = (w12642 & w5562) | (w12642 & w7558) | (w5562 & w7558);
assign w4904 = ~w4110 & ~w8891;
assign w4905 = w6125 & w10804;
assign w4906 = w13892 & w730;
assign w4907 = ~w6749 & w6854;
assign w4908 = ~w6281 & w7317;
assign w4909 = w2608 & w9420;
assign w4910 = ~w3914 & w803;
assign w4911 = w1828 & ~w11934;
assign w4912 = w7385 & w5350;
assign w4913 = ~w13769 & ~w5134;
assign w4914 = ~w3756 & w780;
assign w4915 = ~w142 & ~w2729;
assign w4916 = (w2071 & w12197) | (w2071 & ~w12376) | (w12197 & ~w12376);
assign w4917 = w12385 & ~w5210;
assign w4918 = (~w4099 & w6469) | (~w4099 & w11695) | (w6469 & w11695);
assign w4919 = (~w4453 & w14421) | (~w4453 & w12203) | (w14421 & w12203);
assign w4920 = w1087 & w12648;
assign w4921 = w1116 & ~w13557;
assign w4922 = ~w1840 & ~w7100;
assign w4923 = w3904 & ~w1756;
assign w4924 = ~w14567 & ~w9853;
assign w4925 = (w8551 & ~w2167) | (w8551 & ~w9403) | (~w2167 & ~w9403);
assign w4926 = w3944 & ~w6260;
assign w4927 = ~w12094 & ~w744;
assign w4928 = (~w218 & w10540) | (~w218 & w9426) | (w10540 & w9426);
assign w4929 = (~w1955 & w8608) | (~w1955 & ~w682) | (w8608 & ~w682);
assign w4930 = ~w12167 & w1299;
assign w4931 = ~w9494 & w3627;
assign w4932 = w8512 & ~w3158;
assign w4933 = ~w13903 & ~w11584;
assign w4934 = (~w10189 & ~w10123) | (~w10189 & w8945) | (~w10123 & w8945);
assign w4935 = ~w4213 & w10621;
assign w4936 = (w12499 & w12645) | (w12499 & w1975) | (w12645 & w1975);
assign w4937 = ~w3100 & ~w8234;
assign w4938 = (w2029 & w6611) | (w2029 & w9113) | (w6611 & w9113);
assign w4939 = w10773 & w7719;
assign w4940 = ~w6798 & w12089;
assign w4941 = (~w8645 & w2871) | (~w8645 & w4038) | (w2871 & w4038);
assign w4942 = (w8389 & w1393) | (w8389 & w2011) | (w1393 & w2011);
assign w4943 = (w13492 & w4052) | (w13492 & w600) | (w4052 & w600);
assign w4944 = w12135 & w2798;
assign w4945 = w4310 & w14061;
assign w4946 = w12414 & w2876;
assign w4947 = (w9273 & w4050) | (w9273 & w6089) | (w4050 & w6089);
assign w4948 = w616 & ~w2732;
assign w4949 = w14590 & w12522;
assign w4950 = ~w12939 & ~w13709;
assign w4951 = ~w3435 & ~w2492;
assign w4952 = (~w13306 & w12922) | (~w13306 & w10375) | (w12922 & w10375);
assign w4953 = ~w2643 & w698;
assign w4954 = w6299 & w11613;
assign w4955 = ~w12271 & ~w14430;
assign w4956 = (w13064 & w8299) | (w13064 & w1503) | (w8299 & w1503);
assign w4957 = w10666 & ~w2844;
assign w4958 = ~w9788 & ~w9211;
assign w4959 = w7216 & ~w12927;
assign w4960 = ~w5509 & w3338;
assign w4961 = ~w7335 & ~w10906;
assign w4962 = ~w7681 & ~w7305;
assign w4963 = w3128 & w14250;
assign w4964 = w2656 & w10295;
assign w4965 = ~w14664 & w102;
assign w4966 = w7837 & w7027;
assign w4967 = w8707 & ~w4212;
assign w4968 = w12868 & ~w8992;
assign w4969 = (~w1260 & w4921) | (~w1260 & w6645) | (w4921 & w6645);
assign w4970 = w10781 & ~w12267;
assign w4971 = ~w5522 & ~w5761;
assign w4972 = (w13893 & ~w5783) | (w13893 & w2308) | (~w5783 & w2308);
assign w4973 = w2173 & ~w14504;
assign w4974 = ~w5807 & ~w1163;
assign w4975 = ~w10986 & w3662;
assign w4976 = (~w3700 & w593) | (~w3700 & w14466) | (w593 & w14466);
assign w4977 = (~w7022 & w6128) | (~w7022 & ~w12463) | (w6128 & ~w12463);
assign w4978 = ~w1007 & ~w12779;
assign w4979 = w14246 & w11086;
assign w4980 = w7641 & ~w623;
assign w4981 = w8286 & w3127;
assign w4982 = ~w3587 & w7157;
assign w4983 = (w1663 & w2512) | (w1663 & w4662) | (w2512 & w4662);
assign w4984 = (w9541 & w4363) | (w9541 & w2573) | (w4363 & w2573);
assign w4985 = ~w183 & w8972;
assign w4986 = ~w1261 & w11306;
assign w4987 = ~w5406 & w4467;
assign w4988 = ~w922 & w5482;
assign w4989 = (~w894 & w7722) | (~w894 & w9880) | (w7722 & w9880);
assign w4990 = (~w1842 & w13282) | (~w1842 & w11890) | (w13282 & w11890);
assign w4991 = ~w11284 & ~w12109;
assign w4992 = ~w9925 & ~w10180;
assign w4993 = ~w5522 & ~w6689;
assign w4994 = (~w13587 & w2964) | (~w13587 & w13718) | (w2964 & w13718);
assign w4995 = (~w7439 & w2496) | (~w7439 & w1155) | (w2496 & w1155);
assign w4996 = ~w2144 & w2489;
assign w4997 = (~w13349 & w1217) | (~w13349 & w5383) | (w1217 & w5383);
assign w4998 = w3154 & w11662;
assign w4999 = ~w9595 & w7044;
assign w5000 = (w1489 & ~w11715) | (w1489 & w1538) | (~w11715 & w1538);
assign w5001 = ~w217 & w9296;
assign w5002 = (~w2387 & w3447) | (~w2387 & w1857) | (w3447 & w1857);
assign w5003 = w10676 & w3508;
assign w5004 = ~w2099 & w14265;
assign w5005 = (~w3219 & w3321) | (~w3219 & w9291) | (w3321 & w9291);
assign w5006 = ~w14577 & ~w1127;
assign w5007 = (~w9364 & w5476) | (~w9364 & w9733) | (w5476 & w9733);
assign w5008 = (~w326 & w467) | (~w326 & w11153) | (w467 & w11153);
assign w5009 = ~w2751 & w7951;
assign w5010 = ~w2762 & ~w9324;
assign w5011 = ~w14421 & w6254;
assign w5012 = ~w254 & w2400;
assign w5013 = w13930 & ~w10010;
assign w5014 = w12315 & ~w3587;
assign w5015 = (w10689 & w10245) | (w10689 & w11710) | (w10245 & w11710);
assign w5016 = w12121 & w473;
assign w5017 = (w1699 & w12614) | (w1699 & w5087) | (w12614 & w5087);
assign w5018 = ~w14178 & ~w7423;
assign w5019 = (w11418 & w13205) | (w11418 & w8585) | (w13205 & w8585);
assign w5020 = (w13268 & w4404) | (w13268 & w14188) | (w4404 & w14188);
assign w5021 = ~w9788 & w2701;
assign w5022 = ~w11256 & ~w10416;
assign w5023 = ~w5599 & ~w12933;
assign w5024 = (~w9614 & w3058) | (~w9614 & w1011) | (w3058 & w1011);
assign w5025 = (~w5657 & w11288) | (~w5657 & w4348) | (w11288 & w4348);
assign w5026 = (w1607 & w8389) | (w1607 & w6887) | (w8389 & w6887);
assign w5027 = (w14453 & w4234) | (w14453 & ~w7549) | (w4234 & ~w7549);
assign w5028 = w12868 & w12311;
assign w5029 = ~w9732 & w7068;
assign w5030 = ~w1808 & ~w8845;
assign w5031 = w533 & ~w5449;
assign w5032 = w13935 & ~w14511;
assign w5033 = ~w142 & w5522;
assign w5034 = (~w4050 & w9791) | (~w4050 & w13849) | (w9791 & w13849);
assign w5035 = ~w894 & ~w12065;
assign w5036 = (~w4312 & w6219) | (~w4312 & w7665) | (w6219 & w7665);
assign w5037 = ~w7794 & ~w12464;
assign w5038 = (w952 & w13743) | (w952 & w6948) | (w13743 & w6948);
assign w5039 = (w10708 & ~w1544) | (w10708 & w7994) | (~w1544 & w7994);
assign w5040 = w11459 & ~w392;
assign w5041 = ~w4213 & w3098;
assign w5042 = (w6103 & w13449) | (w6103 & w12116) | (w13449 & w12116);
assign w5043 = w9373 & ~w4621;
assign w5044 = w13579 & w681;
assign w5045 = w10993 & w6932;
assign w5046 = ~w703 & w3200;
assign w5047 = w14030 & ~w3234;
assign w5048 = (w10553 & w4410) | (w10553 & ~w2365) | (w4410 & ~w2365);
assign w5049 = ~w922 & ~w3958;
assign w5050 = ~w1291 & ~w5178;
assign w5051 = ~w13917 & w12466;
assign w5052 = ~w5785 & ~w6975;
assign w5053 = w1559 & ~w2262;
assign w5054 = (w5952 & w1188) | (w5952 & w2200) | (w1188 & w2200);
assign w5055 = w7109 & w7739;
assign w5056 = ~w9608 & w4197;
assign w5057 = (w13463 & w634) | (w13463 & w3511) | (w634 & w3511);
assign w5058 = ~w71 & w13048;
assign w5059 = w11638 & w14340;
assign w5060 = (~w11909 & ~w6929) | (~w11909 & w2936) | (~w6929 & w2936);
assign w5061 = (~w13092 & w8348) | (~w13092 & w4495) | (w8348 & w4495);
assign w5062 = w10211 & ~w1801;
assign w5063 = ~w2701 & ~w2527;
assign w5064 = ~w11929 & ~w13510;
assign w5065 = ~w1201 & ~w1421;
assign w5066 = w13854 & ~w10704;
assign w5067 = ~w8100 & ~w10590;
assign w5068 = ~w10514 & a87;
assign w5069 = ~w14133 & ~w5577;
assign w5070 = ~w127 & ~w8899;
assign w5071 = w9268 & w5669;
assign w5072 = w12371 & ~w13839;
assign w5073 = (w8512 & w2492) | (w8512 & w12637) | (w2492 & w12637);
assign w5074 = (w4607 & w2853) | (w4607 & w4393) | (w2853 & w4393);
assign w5075 = (~w11385 & w10340) | (~w11385 & w2540) | (w10340 & w2540);
assign w5076 = (~w11091 & w11896) | (~w11091 & w12784) | (w11896 & w12784);
assign w5077 = w14451 & w3856;
assign w5078 = ~w7962 & w8427;
assign w5079 = ~w1148 & w10889;
assign w5080 = w14015 & ~w9480;
assign w5081 = w13159 & w13673;
assign w5082 = (w11590 & w3342) | (w11590 & w9947) | (w3342 & w9947);
assign w5083 = (w11429 & w3326) | (w11429 & w2780) | (w3326 & w2780);
assign w5084 = (w10923 & w5009) | (w10923 & w5954) | (w5009 & w5954);
assign w5085 = ~w5628 & w1271;
assign w5086 = (~w4032 & w11914) | (~w4032 & w11487) | (w11914 & w11487);
assign w5087 = ~w7226 & w1699;
assign w5088 = ~w6912 & w7183;
assign w5089 = ~w5664 & w11083;
assign w5090 = ~w6135 & ~w10986;
assign w5091 = ~w2850 & w1692;
assign w5092 = (w6390 & ~w6579) | (w6390 & ~w11005) | (~w6579 & ~w11005);
assign w5093 = w5845 & ~w6292;
assign w5094 = ~w4050 & w9535;
assign w5095 = w13665 & w12614;
assign w5096 = w5015 & w10282;
assign w5097 = w7808 & w7814;
assign w5098 = w3717 & ~w9583;
assign w5099 = ~w8429 & w11029;
assign w5100 = ~w9373 & w10496;
assign w5101 = w7769 & w1636;
assign w5102 = w4031 & ~w7320;
assign w5103 = ~w12240 & ~w14141;
assign w5104 = w9544 & w10365;
assign w5105 = w1114 & w4287;
assign w5106 = ~w566 & ~w8483;
assign w5107 = w7001 & ~w5761;
assign w5108 = ~b33 & ~a33;
assign w5109 = (~w142 & ~w4458) | (~w142 & w6872) | (~w4458 & w6872);
assign w5110 = (w1378 & w10877) | (w1378 & w1219) | (w10877 & w1219);
assign w5111 = (w5662 & w5965) | (w5662 & w1024) | (w5965 & w1024);
assign w5112 = (w13685 & w3504) | (w13685 & w10598) | (w3504 & w10598);
assign w5113 = ~w7244 & ~w5761;
assign w5114 = w10664 & w9748;
assign w5115 = ~w8055 & w10049;
assign w5116 = ~w7897 & w10345;
assign w5117 = (~w996 & w6185) | (~w996 & w11019) | (w6185 & w11019);
assign w5118 = ~w1522 & w10469;
assign w5119 = ~w9298 & w14136;
assign w5120 = (~w7338 & w7169) | (~w7338 & w6572) | (w7169 & w6572);
assign w5121 = ~w11210 & ~w7761;
assign w5122 = (w5756 & w7413) | (w5756 & w4785) | (w7413 & w4785);
assign w5123 = w11068 & ~w9672;
assign w5124 = (w11456 & w13424) | (w11456 & ~w13355) | (w13424 & ~w13355);
assign w5125 = (w3602 & w10462) | (w3602 & w11740) | (w10462 & w11740);
assign w5126 = ~w13423 & ~w235;
assign w5127 = ~w91 & w8456;
assign w5128 = ~w3869 & ~w375;
assign w5129 = (~w10435 & w6010) | (~w10435 & w11672) | (w6010 & w11672);
assign w5130 = (~w10075 & w4360) | (~w10075 & w13559) | (w4360 & w13559);
assign w5131 = ~w9066 & w5290;
assign w5132 = w10765 & w8735;
assign w5133 = w14364 & w12660;
assign w5134 = w8512 & ~w3044;
assign w5135 = ~w3048 & w13967;
assign w5136 = w13743 & w10008;
assign w5137 = ~w4627 & ~w9805;
assign w5138 = (~w13292 & w2885) | (~w13292 & w7730) | (w2885 & w7730);
assign w5139 = w10880 & ~w3611;
assign w5140 = w13713 & w1114;
assign w5141 = ~w10361 & ~w6198;
assign w5142 = (w9644 & w11601) | (w9644 & w4756) | (w11601 & w4756);
assign w5143 = w12544 & w13059;
assign w5144 = (~w1227 & w4984) | (~w1227 & w12843) | (w4984 & w12843);
assign w5145 = ~w409 & ~w3394;
assign w5146 = w8534 & w1443;
assign w5147 = w1208 | w5159;
assign w5148 = ~w14287 & w9456;
assign w5149 = w4323 & ~w12727;
assign w5150 = w7223 & ~w8688;
assign w5151 = (w9716 & ~w11508) | (w9716 & w4901) | (~w11508 & w4901);
assign w5152 = (~w12575 & w9012) | (~w12575 & w13660) | (w9012 & w13660);
assign w5153 = ~w14395 & w4671;
assign w5154 = (w2979 & w6780) | (w2979 & w7549) | (w6780 & w7549);
assign w5155 = ~w11732 & w11759;
assign w5156 = w8396 & w5282;
assign w5157 = ~w11987 & ~w13116;
assign w5158 = w8748 & w9952;
assign w5159 = w10184 & ~w10540;
assign w5160 = (~w9989 & w11673) | (~w9989 & w9431) | (w11673 & w9431);
assign w5161 = (w499 & w14343) | (w499 & w108) | (w14343 & w108);
assign w5162 = ~w5093 & ~w9228;
assign w5163 = w7794 & ~w7881;
assign w5164 = w2578 & w14583;
assign w5165 = w12760 & w9757;
assign w5166 = (w8584 & w6521) | (w8584 & w13236) | (w6521 & w13236);
assign w5167 = (~w14454 & w1362) | (~w14454 & w11277) | (w1362 & w11277);
assign w5168 = w9428 & w10128;
assign w5169 = (w11870 & w11206) | (w11870 & w6310) | (w11206 & w6310);
assign w5170 = (~w10711 & ~w4582) | (~w10711 & ~w13984) | (~w4582 & ~w13984);
assign w5171 = (w10551 & w5294) | (w10551 & w13831) | (w5294 & w13831);
assign w5172 = (~w6802 & w13770) | (~w6802 & w10577) | (w13770 & w10577);
assign w5173 = ~w14015 & w11899;
assign w5174 = ~w12252 & ~w1491;
assign w5175 = ~w11075 & w3275;
assign w5176 = w6176 & ~w14054;
assign w5177 = ~w12785 & ~w13927;
assign w5178 = ~w11216 & ~w14;
assign w5179 = w334 & w484;
assign w5180 = w13732 & ~w11597;
assign w5181 = (w8584 & w5294) | (w8584 & w2171) | (w5294 & w2171);
assign w5182 = (~w14486 & w4032) | (~w14486 & w5656) | (w4032 & w5656);
assign w5183 = ~w11701 & ~w12137;
assign w5184 = w5550 & ~w9232;
assign w5185 = ~w5560 & ~w9263;
assign w5186 = (w762 & w13056) | (w762 & ~w3181) | (w13056 & ~w3181);
assign w5187 = w12464 & w829;
assign w5188 = w12295 & w5664;
assign w5189 = w11364 & w61;
assign w5190 = (~w142 & ~w1062) | (~w142 & w6872) | (~w1062 & w6872);
assign w5191 = ~w6041 & w12614;
assign w5192 = (~w2218 & w3750) | (~w2218 & w1458) | (w3750 & w1458);
assign w5193 = (w7906 & w5559) | (w7906 & w8671) | (w5559 & w8671);
assign w5194 = (w1190 & w13031) | (w1190 & w3299) | (w13031 & w3299);
assign w5195 = ~w2036 & ~w2701;
assign w5196 = (w6301 & ~w1340) | (w6301 & w11788) | (~w1340 & w11788);
assign w5197 = w12604 & w11031;
assign w5198 = w569 & w2035;
assign w5199 = ~w8791 & w2719;
assign w5200 = ~w13189 & ~w8727;
assign w5201 = ~w9711 & ~w5707;
assign w5202 = w4219 & w5131;
assign w5203 = ~w5522 & ~w10699;
assign w5204 = w11900 & w12639;
assign w5205 = w3914 & ~w1052;
assign w5206 = ~w5194 & w1053;
assign w5207 = w13596 & w2592;
assign w5208 = w9921 & w6575;
assign w5209 = w8694 & w8297;
assign w5210 = (~w2299 & w3930) | (~w2299 & w13933) | (w3930 & w13933);
assign w5211 = ~w2035 & w6473;
assign w5212 = ~w6352 & ~w8093;
assign w5213 = ~w8171 & ~w10675;
assign w5214 = ~w5522 & ~w8396;
assign w5215 = ~w14072 & w2811;
assign w5216 = w1507 & ~w7630;
assign w5217 = ~w9480 & w6689;
assign w5218 = ~w2566 & ~w7370;
assign w5219 = (w894 & w13349) | (w894 & w7081) | (w13349 & w7081);
assign w5220 = ~w14647 & w7017;
assign w5221 = w2387 & ~w2922;
assign w5222 = ~w7794 & w14048;
assign w5223 = w11287 & w13323;
assign w5224 = ~w2951 & ~w10309;
assign w5225 = ~w5556 & ~w14395;
assign w5226 = w10708 & ~w7561;
assign w5227 = ~w9244 & ~w8626;
assign w5228 = (~w1794 & w12175) | (~w1794 & ~w6697) | (w12175 & ~w6697);
assign w5229 = w9324 & ~w50;
assign w5230 = ~w11500 & w11420;
assign w5231 = (~w3751 & w7111) | (~w3751 & w8272) | (w7111 & w8272);
assign w5232 = (~w445 & ~w2243) | (~w445 & ~w7047) | (~w2243 & ~w7047);
assign w5233 = ~w10186 & ~w8090;
assign w5234 = w7401 & ~w12543;
assign w5235 = (w8501 & w8932) | (w8501 & w3677) | (w8932 & w3677);
assign w5236 = w3586 & w6965;
assign w5237 = ~w1740 & w13710;
assign w5238 = w13967 & ~w12487;
assign w5239 = (w4405 & w3277) | (w4405 & ~w1386) | (w3277 & ~w1386);
assign w5240 = w607 & ~w1540;
assign w5241 = (~w2463 & w7574) | (~w2463 & w2621) | (w7574 & w2621);
assign w5242 = w7662 & ~w8499;
assign w5243 = ~w3508 & ~w2680;
assign w5244 = w9212 & w3427;
assign w5245 = w7669 & w14514;
assign w5246 = w8978 & ~w7693;
assign w5247 = w3963 & ~w14491;
assign w5248 = ~w10676 & w3441;
assign w5249 = (w1033 & w9073) | (w1033 & w12376) | (w9073 & w12376);
assign w5250 = ~w5829 & ~w12183;
assign w5251 = w13459 & ~w13630;
assign w5252 = w9453 & ~w6889;
assign w5253 = ~w11302 & w7392;
assign w5254 = ~w13462 & w7145;
assign w5255 = (w2142 & w2315) | (w2142 & w9865) | (w2315 & w9865);
assign w5256 = (w9329 & ~w2) | (w9329 & ~w14564) | (~w2 & ~w14564);
assign w5257 = ~w10403 & w12469;
assign w5258 = ~w7792 & ~w9459;
assign w5259 = (w12761 & w6221) | (w12761 & w8228) | (w6221 & w8228);
assign w5260 = (w12774 & ~w6787) | (w12774 & ~w11986) | (~w6787 & ~w11986);
assign w5261 = ~w7488 & w1021;
assign w5262 = ~w9226 & ~w14395;
assign w5263 = ~w7317 & w7165;
assign w5264 = ~w3427 & ~w9498;
assign w5265 = (w15 & w14046) | (w15 & w3350) | (w14046 & w3350);
assign w5266 = w7794 & ~w14563;
assign w5267 = ~w569 & ~w10621;
assign w5268 = (w11902 & w13324) | (w11902 & w85) | (w13324 & w85);
assign w5269 = (~w9305 & w4260) | (~w9305 & w14165) | (w4260 & w14165);
assign w5270 = ~w7191 & w634;
assign w5271 = ~w4700 & w2941;
assign w5272 = w3456 & ~w6684;
assign w5273 = (~w8374 & ~w4092) | (~w8374 & w3223) | (~w4092 & w3223);
assign w5274 = ~w8248 & ~w13640;
assign w5275 = w3957 & w7357;
assign w5276 = ~w6027 & ~w4641;
assign w5277 = (w835 & w10734) | (w835 & ~w8228) | (w10734 & ~w8228);
assign w5278 = (w11594 & ~w5351) | (w11594 & w7937) | (~w5351 & w7937);
assign w5279 = ~w3851 & w11583;
assign w5280 = w2387 & ~w12614;
assign w5281 = ~w4714 & w10782;
assign w5282 = ~w9846 & ~w10082;
assign w5283 = w12429 & ~w13423;
assign w5284 = (~w2029 & w4457) | (~w2029 & w13698) | (w4457 & w13698);
assign w5285 = w12656 & ~w2320;
assign w5286 = ~w14227 & ~w2680;
assign w5287 = (~w934 & w10468) | (~w934 & w10838) | (w10468 & w10838);
assign w5288 = ~w12604 & ~w7335;
assign w5289 = w12135 & w3406;
assign w5290 = w8562 & w955;
assign w5291 = ~w13095 & ~w7423;
assign w5292 = w13598 & w11381;
assign w5293 = (w4784 & w11133) | (w4784 & ~w8282) | (w11133 & ~w8282);
assign w5294 = ~w6069 & ~w2830;
assign w5295 = w3682 & ~w3892;
assign w5296 = ~w4921 & w440;
assign w5297 = w7743 & ~w11942;
assign w5298 = w5890 & w9770;
assign w5299 = (w11159 & w8937) | (w11159 & w4243) | (w8937 & w4243);
assign w5300 = w509 & w10918;
assign w5301 = (~w4312 & ~w9183) | (~w4312 & w10945) | (~w9183 & w10945);
assign w5302 = ~w3498 & ~w11408;
assign w5303 = ~w12003 & w493;
assign w5304 = ~w12199 & ~w7091;
assign w5305 = ~w4700 & w6500;
assign w5306 = ~w9432 & w12624;
assign w5307 = ~w7190 & ~w1873;
assign w5308 = (w4021 & ~w1986) | (w4021 & w11096) | (~w1986 & w11096);
assign w5309 = w3914 & ~w14425;
assign w5310 = ~w11045 & w5115;
assign w5311 = ~w13222 & ~w9036;
assign w5312 = ~w260 & ~w2941;
assign w5313 = ~w7794 & w11855;
assign w5314 = ~w13730 & ~w4458;
assign w5315 = ~w7886 & ~w12992;
assign w5316 = ~w14412 & ~w7841;
assign w5317 = ~w10408 & ~w6433;
assign w5318 = (w4511 & w721) | (w4511 & w9799) | (w721 & w9799);
assign w5319 = (~w2381 & ~w8499) | (~w2381 & ~w217) | (~w8499 & ~w217);
assign w5320 = w14072 & ~w12438;
assign w5321 = w318 & w12543;
assign w5322 = ~a53 & ~w7606;
assign w5323 = (w4127 & w11716) | (w4127 & ~w8992) | (w11716 & ~w8992);
assign w5324 = (w5070 & w9519) | (w5070 & w9962) | (w9519 & w9962);
assign w5325 = ~w462 & ~w9031;
assign w5326 = ~w3209 & w5906;
assign w5327 = ~w3926 & w8558;
assign w5328 = w4312 & ~w10483;
assign w5329 = (w9932 & w13152) | (w9932 & w12835) | (w13152 & w12835);
assign w5330 = ~w254 & w5478;
assign w5331 = (w2374 & w6366) | (w2374 & w12595) | (w6366 & w12595);
assign w5332 = ~w5178 & ~w5513;
assign w5333 = (~w1096 & w3321) | (~w1096 & w6112) | (w3321 & w6112);
assign w5334 = w2060 & ~w2639;
assign w5335 = ~w1023 & ~w12802;
assign w5336 = w4032 & ~w12192;
assign w5337 = (w10551 & w1692) | (w10551 & w1786) | (w1692 & w1786);
assign w5338 = ~w12481 & ~w4458;
assign w5339 = ~w12158 & ~w150;
assign w5340 = (~w8440 & w7094) | (~w8440 & w3880) | (w7094 & w3880);
assign w5341 = ~w7819 & ~w11887;
assign w5342 = ~w5742 & ~w12866;
assign w5343 = ~w10077 & w6985;
assign w5344 = ~w6193 & ~w2079;
assign w5345 = w12714 & w10081;
assign w5346 = ~w12609 & ~w4515;
assign w5347 = ~w5522 & ~w13937;
assign w5348 = w12267 & w14389;
assign w5349 = w14504 & w9013;
assign w5350 = (w10123 & w5720) | (w10123 & w4876) | (w5720 & w4876);
assign w5351 = ~w2359 & w4309;
assign w5352 = w7673 & ~w12420;
assign w5353 = w2509 & w1743;
assign w5354 = ~w2463 & w3022;
assign w5355 = (~w9226 & ~w1885) | (~w9226 & w9976) | (~w1885 & w9976);
assign w5356 = w12528 & ~w10033;
assign w5357 = w621 & ~w309;
assign w5358 = (w12589 & w6384) | (w12589 & w3102) | (w6384 & w3102);
assign w5359 = (~w8347 & w8232) | (~w8347 & ~w9262) | (w8232 & ~w9262);
assign w5360 = (w12569 & ~w14302) | (w12569 & w1217) | (~w14302 & w1217);
assign w5361 = (w10553 & w4410) | (w10553 & ~w2904) | (w4410 & ~w2904);
assign w5362 = w13924 & ~w5860;
assign w5363 = ~w7444 & w8438;
assign w5364 = ~w1727 & ~w12746;
assign w5365 = (w8019 & w7967) | (w8019 & w9275) | (w7967 & w9275);
assign w5366 = ~w327 & w14645;
assign w5367 = w13008 & w876;
assign w5368 = (~w4679 & w14461) | (~w4679 & w1783) | (w14461 & w1783);
assign w5369 = w3550 & w12725;
assign w5370 = ~w3629 & w9849;
assign w5371 = w5626 & ~w2370;
assign w5372 = w2114 & w6311;
assign w5373 = (~w3007 & w11167) | (~w3007 & w6242) | (w11167 & w6242);
assign w5374 = ~w3920 & w3368;
assign w5375 = w14302 & w894;
assign w5376 = ~w4050 & w5311;
assign w5377 = (w3521 & w13098) | (w3521 & ~w3356) | (w13098 & ~w3356);
assign w5378 = ~w4751 & ~w6795;
assign w5379 = ~w10824 & ~w7261;
assign w5380 = (~w2168 & w13184) | (~w2168 & w1548) | (w13184 & w1548);
assign w5381 = (w11983 & w2515) | (w11983 & w84) | (w2515 & w84);
assign w5382 = w4299 & w12311;
assign w5383 = (w12569 & ~w5294) | (w12569 & w1217) | (~w5294 & w1217);
assign w5384 = ~w14486 & ~w2159;
assign w5385 = w12575 & w1507;
assign w5386 = w11216 & ~w12958;
assign w5387 = (~w10676 & w3441) | (~w10676 & ~w10987) | (w3441 & ~w10987);
assign w5388 = w4171 & w1508;
assign w5389 = ~w14607 & w8887;
assign w5390 = w114 & w3484;
assign w5391 = (w659 & w3505) | (w659 & ~w7549) | (w3505 & ~w7549);
assign w5392 = (w11261 & w369) | (w11261 & w7119) | (w369 & w7119);
assign w5393 = ~w6823 & ~w8038;
assign w5394 = w7981 & ~w3835;
assign w5395 = ~w3036 & ~w10247;
assign w5396 = ~w14215 & w9478;
assign w5397 = ~w6572 & ~w12398;
assign w5398 = w12943 & ~w3508;
assign w5399 = (~w5783 & w4466) | (~w5783 & w3948) | (w4466 & w3948);
assign w5400 = (w9921 & ~w11084) | (w9921 & w2920) | (~w11084 & w2920);
assign w5401 = (w12285 & w6517) | (w12285 & w9984) | (w6517 & w9984);
assign w5402 = (~w142 & ~w10182) | (~w142 & w6872) | (~w10182 & w6872);
assign w5403 = (~w13772 & w12995) | (~w13772 & w8600) | (w12995 & w8600);
assign w5404 = w4453 & w5662;
assign w5405 = w8513 & ~w2372;
assign w5406 = ~b63 & ~a63;
assign w5407 = (w807 & w10926) | (w807 & w14128) | (w10926 & w14128);
assign w5408 = (w13136 & w4724) | (w13136 & w2861) | (w4724 & w2861);
assign w5409 = w7942 & w11947;
assign w5410 = (w4050 & w8805) | (w4050 & w5572) | (w8805 & w5572);
assign w5411 = w10198 & ~w6381;
assign w5412 = ~w4071 & ~w8110;
assign w5413 = ~w4561 & w13018;
assign w5414 = (w9749 & w2667) | (w9749 & w8979) | (w2667 & w8979);
assign w5415 = ~w922 & w2159;
assign w5416 = ~w12271 & w5406;
assign w5417 = w12614 & ~w9326;
assign w5418 = w9990 & w4041;
assign w5419 = ~w4159 & ~w13610;
assign w5420 = ~w11155 & ~w13490;
assign w5421 = ~w6583 & ~w9949;
assign w5422 = ~w14470 & ~w13902;
assign w5423 = w500 & w1815;
assign w5424 = w6889 & w12893;
assign w5425 = w10317 & w2492;
assign w5426 = (~w3550 & w3393) | (~w3550 & w1185) | (w3393 & w1185);
assign w5427 = ~w5172 & ~w289;
assign w5428 = ~w11701 & w526;
assign w5429 = w7085 & w6858;
assign w5430 = ~w3960 & ~w10168;
assign w5431 = ~w7919 & ~w8696;
assign w5432 = ~w1802 & w11861;
assign w5433 = (w1849 & w14615) | (w1849 & w1214) | (w14615 & w1214);
assign w5434 = w10290 & ~w5262;
assign w5435 = ~w12452 & w2069;
assign w5436 = (~w8973 & w6720) | (~w8973 & ~w11448) | (w6720 & ~w11448);
assign w5437 = w14396 & w3184;
assign w5438 = (w12332 & w11923) | (w12332 & ~w10023) | (w11923 & ~w10023);
assign w5439 = w7190 & w9244;
assign w5440 = ~w1333 & w6738;
assign w5441 = ~w8226 & w14394;
assign w5442 = ~w13587 & w1617;
assign w5443 = (w6266 & w4252) | (w6266 & w3963) | (w4252 & w3963);
assign w5444 = ~w10231 & w12261;
assign w5445 = (w7811 & w6240) | (w7811 & w3564) | (w6240 & w3564);
assign w5446 = ~w3885 & w3427;
assign w5447 = w616 & ~w12165;
assign w5448 = ~w2218 & w10316;
assign w5449 = ~w6656 & w7271;
assign w5450 = w11750 & ~w10279;
assign w5451 = ~w14072 & ~w7906;
assign w5452 = (~w10123 & w3220) | (~w10123 & w11797) | (w3220 & w11797);
assign w5453 = ~w12980 & w7264;
assign w5454 = ~w7606 & ~w5347;
assign w5455 = w1096 & ~w2933;
assign w5456 = w14215 & ~w12589;
assign w5457 = ~w4627 & w923;
assign w5458 = (~w14128 & w13255) | (~w14128 & w5929) | (w13255 & w5929);
assign w5459 = ~w7449 & ~w5433;
assign w5460 = ~w5867 & ~w8707;
assign w5461 = w3944 & ~w13265;
assign w5462 = w848 & ~w1864;
assign w5463 = ~w7542 & w4452;
assign w5464 = ~w7190 & ~w2410;
assign w5465 = (w3039 & ~w5867) | (w3039 & w6728) | (~w5867 & w6728);
assign w5466 = w14447 & ~w7687;
assign w5467 = ~w5294 & ~w9784;
assign w5468 = ~w2352 & w2449;
assign w5469 = ~w12271 & w2410;
assign w5470 = ~w2138 & ~w785;
assign w5471 = ~w7855 & w11263;
assign w5472 = w142 & w3508;
assign w5473 = ~w10023 & w4305;
assign w5474 = (~w11915 & w2856) | (~w11915 & w13784) | (w2856 & w13784);
assign w5475 = ~w882 & ~w12992;
assign w5476 = (~w9403 & w8282) | (~w9403 & w6310) | (w8282 & w6310);
assign w5477 = w4173 & w6308;
assign w5478 = ~w1840 & w9301;
assign w5479 = (~w8937 & w1566) | (~w8937 & w8393) | (w1566 & w8393);
assign w5480 = ~w12816 & w13204;
assign w5481 = w2035 & w14550;
assign w5482 = ~w1096 & ~w3971;
assign w5483 = (w14463 & w10613) | (w14463 & w12638) | (w10613 & w12638);
assign w5484 = (w9007 & w3391) | (w9007 & w5007) | (w3391 & w5007);
assign w5485 = w10975 & w1144;
assign w5486 = (~w10139 & ~w7399) | (~w10139 & w10147) | (~w7399 & w10147);
assign w5487 = ~w6583 & w7410;
assign w5488 = (w1640 & w7129) | (w1640 & w12376) | (w7129 & w12376);
assign w5489 = ~w4322 & w9296;
assign w5490 = (~w8992 & w3700) | (~w8992 & w2020) | (w3700 & w2020);
assign w5491 = (w5331 & w4436) | (w5331 & w9034) | (w4436 & w9034);
assign w5492 = (w1770 & w8235) | (w1770 & w7062) | (w8235 & w7062);
assign w5493 = (~w7782 & w886) | (~w7782 & w7174) | (w886 & w7174);
assign w5494 = w11275 & w11367;
assign w5495 = w563 & w9748;
assign w5496 = ~w607 & ~w10699;
assign w5497 = ~w10856 & ~w2104;
assign w5498 = w11475 & ~w4741;
assign w5499 = (w2975 & w3207) | (w2975 & w12376) | (w3207 & w12376);
assign w5500 = w1342 & w6195;
assign w5501 = (~w10023 & w2554) | (~w10023 & w3660) | (w2554 & w3660);
assign w5502 = (~w4856 & w12515) | (~w4856 & w3190) | (w12515 & w3190);
assign w5503 = w12315 & w3904;
assign w5504 = ~w4900 & w4942;
assign w5505 = ~w4080 & ~w8085;
assign w5506 = ~w3986 & ~w235;
assign w5507 = (~w10434 & ~w6701) | (~w10434 & w12570) | (~w6701 & w12570);
assign w5508 = (w10832 & w8627) | (w10832 & ~w13980) | (w8627 & ~w13980);
assign w5509 = ~w12322 & w4161;
assign w5510 = w12240 & w6572;
assign w5511 = w13175 & ~w7256;
assign w5512 = (~w14421 & w2775) | (~w14421 & w4977) | (w2775 & w4977);
assign w5513 = w5213 & w5660;
assign w5514 = w14091 & w8023;
assign w5515 = ~w11152 & w8357;
assign w5516 = ~w4158 & w14008;
assign w5517 = w13800 & ~w1905;
assign w5518 = (~w12915 & w13519) | (~w12915 & ~w5867) | (w13519 & ~w5867);
assign w5519 = w4787 & ~w12170;
assign w5520 = ~w4032 & w3508;
assign w5521 = ~w5851 & ~w11454;
assign w5522 = ~b94 & ~a94;
assign w5523 = (w14463 & w11347) | (w14463 & w6862) | (w11347 & w6862);
assign w5524 = (w13685 & w4406) | (w13685 & w14106) | (w4406 & w14106);
assign w5525 = (w11617 & w4689) | (w11617 & w14057) | (w4689 & w14057);
assign w5526 = ~w12682 & w7885;
assign w5527 = (~w14600 & w9470) | (~w14600 & w222) | (w9470 & w222);
assign w5528 = (~w4097 & w6481) | (~w4097 & w13274) | (w6481 & w13274);
assign w5529 = (~w10541 & w7194) | (~w10541 & w13577) | (w7194 & w13577);
assign w5530 = (~w14564 & w14506) | (~w14564 & w12588) | (w14506 & w12588);
assign w5531 = ~w4700 & w488;
assign w5532 = (~w3025 & w7704) | (~w3025 & w3737) | (w7704 & w3737);
assign w5533 = w4787 & ~w4363;
assign w5534 = w4503 & ~w4565;
assign w5535 = ~w3434 & ~w13959;
assign w5536 = ~w12240 & w5556;
assign w5537 = ~w8907 & ~w6792;
assign w5538 = w3568 & ~w2762;
assign w5539 = w9989 & w14167;
assign w5540 = ~w1616 & ~w11518;
assign w5541 = (~w10520 & w7971) | (~w10520 & w8397) | (w7971 & w8397);
assign w5542 = (~w14486 & w2144) | (~w14486 & w5182) | (w2144 & w5182);
assign w5543 = w1760 & w6230;
assign w5544 = (w9757 & ~w13320) | (w9757 & w5165) | (~w13320 & w5165);
assign w5545 = w14614 & ~w11013;
assign w5546 = (~w12499 & w6600) | (~w12499 & w5387) | (w6600 & w5387);
assign w5547 = ~w4080 & ~w119;
assign w5548 = w13452 & ~w11654;
assign w5549 = ~w2698 & w3154;
assign w5550 = ~w11588 & w7061;
assign w5551 = ~w7940 & w573;
assign w5552 = w6630 & w9702;
assign w5553 = (~w628 & w8144) | (~w628 & w1793) | (w8144 & w1793);
assign w5554 = ~w3885 & w2701;
assign w5555 = ~w6275 & w2655;
assign w5556 = b58 & a58;
assign w5557 = w12681 & w11061;
assign w5558 = ~w13462 & w5649;
assign w5559 = ~w2467 & ~w6298;
assign w5560 = b18 & a18;
assign w5561 = w8412 & w3564;
assign w5562 = ~w2101 & w5912;
assign w5563 = (~w4512 & w893) | (~w4512 & w9178) | (w893 & w9178);
assign w5564 = ~w12867 & ~w7037;
assign w5565 = w9623 & ~w12642;
assign w5566 = w11510 & ~w5454;
assign w5567 = (w12605 & w14154) | (w12605 & ~w14182) | (w14154 & ~w14182);
assign w5568 = (~w473 & w3024) | (~w473 & w13759) | (w3024 & w13759);
assign w5569 = ~w14072 & ~w14227;
assign w5570 = (w10277 & ~w11744) | (w10277 & w177) | (~w11744 & w177);
assign w5571 = w10823 & ~w5167;
assign w5572 = (w2858 & w2567) | (w2858 & w13608) | (w2567 & w13608);
assign w5573 = ~w569 & w249;
assign w5574 = ~w12081 & w9377;
assign w5575 = ~w11462 & ~w12664;
assign w5576 = ~w8098 & ~w3302;
assign w5577 = ~w10221 & w2701;
assign w5578 = ~w8476 & ~w6118;
assign w5579 = w3098 & w9715;
assign w5580 = ~w11997 & ~w10290;
assign w5581 = ~w14141 & w8470;
assign w5582 = ~w4700 & w13839;
assign w5583 = w11821 & w5462;
assign w5584 = ~w14153 & w444;
assign w5585 = w10961 & ~w3209;
assign w5586 = ~w3751 & w11031;
assign w5587 = (w4679 & w1277) | (w4679 & w2588) | (w1277 & w2588);
assign w5588 = (w10123 & w11311) | (w10123 & w9413) | (w11311 & w9413);
assign w5589 = w10676 & ~w12915;
assign w5590 = ~w1682 & ~w13344;
assign w5591 = ~w11412 & w8702;
assign w5592 = w8328 & w11817;
assign w5593 = w13838 & w2891;
assign w5594 = (w11803 & w6543) | (w11803 & w13326) | (w6543 & w13326);
assign w5595 = (w6719 & ~w3708) | (w6719 & w9094) | (~w3708 & w9094);
assign w5596 = ~w1065 & w9699;
assign w5597 = w8572 & w10421;
assign w5598 = w8819 & ~w10699;
assign w5599 = w12479 & w3017;
assign w5600 = (w12398 & w10462) | (w12398 & w9943) | (w10462 & w9943);
assign w5601 = ~w2223 & ~w10802;
assign w5602 = w3038 & w3957;
assign w5603 = (w9831 & ~w630) | (w9831 & ~w10214) | (~w630 & ~w10214);
assign w5604 = ~w2369 & ~w2189;
assign w5605 = ~w6433 & ~w5936;
assign w5606 = (~w14600 & w11592) | (~w14600 & w5208) | (w11592 & w5208);
assign w5607 = ~w7546 & ~w3863;
assign w5608 = ~w4963 & w13514;
assign w5609 = ~w10712 & ~w654;
assign w5610 = w5643 & w2704;
assign w5611 = (w857 & w1960) | (w857 & w13860) | (w1960 & w13860);
assign w5612 = ~w7438 & ~w6049;
assign w5613 = w5412 & w260;
assign w5614 = w3927 & ~w12703;
assign w5615 = w4417 & w10665;
assign w5616 = w8931 & w1301;
assign w5617 = ~w5343 & w10463;
assign w5618 = (w13873 & ~w4803) | (w13873 & w4434) | (~w4803 & w4434);
assign w5619 = ~w7000 & ~w9122;
assign w5620 = w3550 & w11353;
assign w5621 = w4523 & w7376;
assign w5622 = w852 & ~w7423;
assign w5623 = w2671 & w926;
assign w5624 = (~w14070 & w10462) | (~w14070 & w66) | (w10462 & w66);
assign w5625 = (w6397 & w13329) | (w6397 & w8892) | (w13329 & w8892);
assign w5626 = (~w6889 & w13838) | (~w6889 & w1010) | (w13838 & w1010);
assign w5627 = ~w10278 & w1267;
assign w5628 = w3104 & ~w14071;
assign w5629 = w7486 & w12705;
assign w5630 = ~w8153 & w5144;
assign w5631 = w13219 & ~w11692;
assign w5632 = ~w9914 & w13217;
assign w5633 = ~w5036 & w10483;
assign w5634 = ~w3159 & w1729;
assign w5635 = ~w109 & ~w12407;
assign w5636 = ~w7315 & w11450;
assign w5637 = (w13595 & w3818) | (w13595 & w971) | (w3818 & w971);
assign w5638 = w9623 & ~w9296;
assign w5639 = (~w13685 & w4435) | (~w13685 & w9033) | (w4435 & w9033);
assign w5640 = (~w445 & ~w2243) | (~w445 & w6753) | (~w2243 & w6753);
assign w5641 = ~w9012 & w6451;
assign w5642 = ~w2463 & w2482;
assign w5643 = ~w12070 & w501;
assign w5644 = ~w5200 & ~w7776;
assign w5645 = ~w2656 & w803;
assign w5646 = (w10613 & w1354) | (w10613 & w3834) | (w1354 & w3834);
assign w5647 = ~w4834 & ~w2523;
assign w5648 = ~w2230 & ~w12680;
assign w5649 = ~w14302 & w12398;
assign w5650 = (~w9305 & w2402) | (~w9305 & w11413) | (w2402 & w11413);
assign w5651 = (w10574 & w13951) | (w10574 & w13731) | (w13951 & w13731);
assign w5652 = w5522 & w13323;
assign w5653 = (w11768 & w8536) | (w11768 & ~w5570) | (w8536 & ~w5570);
assign w5654 = (w2616 & w3874) | (w2616 & w11010) | (w3874 & w11010);
assign w5655 = w7794 & w8615;
assign w5656 = ~w9871 & ~w14486;
assign w5657 = (w5998 & w9614) | (w5998 & w11545) | (w9614 & w11545);
assign w5658 = ~w4780 & w10409;
assign w5659 = w12464 & w1758;
assign w5660 = ~w2933 & ~w6651;
assign w5661 = w8234 & w9871;
assign w5662 = (~w8399 & w8336) | (~w8399 & w8323) | (w8336 & w8323);
assign w5663 = (~w10514 & w11261) | (~w10514 & w2205) | (w11261 & w2205);
assign w5664 = ~w2176 & ~w7714;
assign w5665 = w8796 & ~w2870;
assign w5666 = ~w11429 & w3262;
assign w5667 = (~w5189 & w11287) | (~w5189 & w3475) | (w11287 & w3475);
assign w5668 = (w7709 & w6470) | (w7709 & w8219) | (w6470 & w8219);
assign w5669 = w7034 & ~w4102;
assign w5670 = w6084 & ~w10317;
assign w5671 = ~w114 & w7022;
assign w5672 = ~w4312 & w7727;
assign w5673 = ~w7080 & ~w9433;
assign w5674 = w4738 & w10045;
assign w5675 = ~w10454 & w13167;
assign w5676 = w11211 & ~w235;
assign w5677 = ~w1474 & w10699;
assign w5678 = ~w13563 & ~w4631;
assign w5679 = w11041 & ~w2229;
assign w5680 = (~w3608 & w826) | (~w3608 & w1451) | (w826 & w1451);
assign w5681 = ~w11560 & w719;
assign w5682 = w3075 & ~w9296;
assign w5683 = (w8085 & w7873) | (w8085 & w13238) | (w7873 & w13238);
assign w5684 = w4299 & ~w8992;
assign w5685 = ~w12980 & w1937;
assign w5686 = ~w2941 & ~w5879;
assign w5687 = ~w12800 & ~w8654;
assign w5688 = ~w2144 & w7238;
assign w5689 = (w12330 & ~w3122) | (w12330 & w6803) | (~w3122 & w6803);
assign w5690 = ~w9015 & w5865;
assign w5691 = ~w10523 & ~w11560;
assign w5692 = ~w8512 & ~w5732;
assign w5693 = ~b78 & ~a78;
assign w5694 = ~w1507 & ~w136;
assign w5695 = (w8405 & w6392) | (w8405 & w2414) | (w6392 & w2414);
assign w5696 = w4270 & ~w5282;
assign w5697 = ~w7410 & w8247;
assign w5698 = (w1968 & w6980) | (w1968 & w7062) | (w6980 & w7062);
assign w5699 = (w5977 & w2916) | (w5977 & w5008) | (w2916 & w5008);
assign w5700 = ~w13349 & w3735;
assign w5701 = w840 & ~w668;
assign w5702 = ~w5949 & w14238;
assign w5703 = ~w922 & w3508;
assign w5704 = ~w1992 & ~w11569;
assign w5705 = w7084 & w12140;
assign w5706 = w13596 & ~w10031;
assign w5707 = (~w8691 & w13872) | (~w8691 & w12177) | (w13872 & w12177);
assign w5708 = w2909 & ~w5814;
assign w5709 = ~w1629 & ~w6727;
assign w5710 = ~w3469 & w12370;
assign w5711 = w791 & w1766;
assign w5712 = w9226 & ~w5845;
assign w5713 = w5817 | w13899;
assign w5714 = ~w9253 & w3186;
assign w5715 = (w5788 & ~w2060) | (w5788 & w9839) | (~w2060 & w9839);
assign w5716 = ~w9454 & ~w10778;
assign w5717 = ~w5732 & w8085;
assign w5718 = (w6739 & w1960) | (w6739 & w390) | (w1960 & w390);
assign w5719 = w7914 & w10465;
assign w5720 = (w758 & w1245) | (w758 & ~w1304) | (w1245 & ~w1304);
assign w5721 = ~w6500 & w5915;
assign w5722 = w4312 & w6952;
assign w5723 = (~w341 & w254) | (~w341 & w12066) | (w254 & w12066);
assign w5724 = (~w7244 & ~w863) | (~w7244 & w7736) | (~w863 & w7736);
assign w5725 = ~w7030 & ~w3898;
assign w5726 = (w12799 & w6863) | (w12799 & w9473) | (w6863 & w9473);
assign w5727 = (~w12537 & w1094) | (~w12537 & w354) | (w1094 & w354);
assign w5728 = (~w1844 & w14269) | (~w1844 & w13614) | (w14269 & w13614);
assign w5729 = ~w183 & w4299;
assign w5730 = w7111 & w11410;
assign w5731 = w11364 & ~w13866;
assign w5732 = b65 & a65;
assign w5733 = w3914 & w4299;
assign w5734 = ~w12167 & w12869;
assign w5735 = (~w8234 & ~w11261) | (~w8234 & w9671) | (~w11261 & w9671);
assign w5736 = w9672 & w8389;
assign w5737 = w1507 & w6929;
assign w5738 = w11202 & ~w9999;
assign w5739 = w10045 & w11592;
assign w5740 = ~w7303 & w7007;
assign w5741 = b50 & a50;
assign w5742 = (~w1821 & w577) | (~w1821 & w10317) | (w577 & w10317);
assign w5743 = w533 & w10781;
assign w5744 = w2270 & w2135;
assign w5745 = (w7455 & w5294) | (w7455 & w10892) | (w5294 & w10892);
assign w5746 = (~w14425 & w2175) | (~w14425 & w5309) | (w2175 & w5309);
assign w5747 = (w13733 & w10462) | (w13733 & w13777) | (w10462 & w13777);
assign w5748 = w6478 & w178;
assign w5749 = ~w7845 & w602;
assign w5750 = ~w2539 & w4944;
assign w5751 = (~w8793 & w5490) | (~w8793 & w8474) | (w5490 & w8474);
assign w5752 = ~w12619 & w9095;
assign w5753 = (w13405 & w5143) | (w13405 & w10583) | (w5143 & w10583);
assign w5754 = ~b36 & ~a36;
assign w5755 = ~w8827 & w10423;
assign w5756 = (w6802 & w927) | (w6802 & w10878) | (w927 & w10878);
assign w5757 = (~w8761 & ~w12666) | (~w8761 & w14521) | (~w12666 & w14521);
assign w5758 = ~w13636 & w5891;
assign w5759 = ~w5732 & ~w10423;
assign w5760 = w12604 & w3904;
assign w5761 = ~w10354 & ~w2228;
assign w5762 = ~w9940 & w10398;
assign w5763 = ~w13222 & w7668;
assign w5764 = (w4149 & w13301) | (w4149 & w4568) | (w13301 & w4568);
assign w5765 = ~w11462 & w3224;
assign w5766 = w7001 & w2701;
assign w5767 = w9817 & w1873;
assign w5768 = (~w12943 & w12) | (~w12943 & w6061) | (w12 & w6061);
assign w5769 = (w6886 & w5213) | (w6886 & w3513) | (w5213 & w3513);
assign w5770 = (~w10719 & w6594) | (~w10719 & w13999) | (w6594 & w13999);
assign w5771 = ~w9539 & w990;
assign w5772 = ~w5741 & ~w13306;
assign w5773 = (w5952 & w753) | (w5952 & w8686) | (w753 & w8686);
assign w5774 = w1842 & ~w12958;
assign w5775 = (~w10245 & w5824) | (~w10245 & w3701) | (w5824 & w3701);
assign w5776 = (w14360 & w9311) | (w14360 & w4783) | (w9311 & w4783);
assign w5777 = ~w12249 & w891;
assign w5778 = (~w9788 & w8113) | (~w9788 & w6474) | (w8113 & w6474);
assign w5779 = ~w7742 & w13203;
assign w5780 = ~w13839 & w11442;
assign w5781 = ~w13282 & ~w7782;
assign w5782 = ~w142 & ~w2701;
assign w5783 = (~w4336 & w13364) | (~w4336 & w1488) | (w13364 & w1488);
assign w5784 = ~w13188 & ~w8019;
assign w5785 = ~b38 & ~a38;
assign w5786 = (w5483 & w13455) | (w5483 & w2970) | (w13455 & w2970);
assign w5787 = (~w2544 & w10462) | (~w2544 & w11130) | (w10462 & w11130);
assign w5788 = w13694 & w5569;
assign w5789 = ~w12483 & w4870;
assign w5790 = w3963 & ~w10182;
assign w5791 = ~w10182 & ~w11745;
assign w5792 = w9015 & ~w852;
assign w5793 = w14178 & ~w8512;
assign w5794 = w12922 & ~w9296;
assign w5795 = ~w9012 & w1424;
assign w5796 = (w7062 & w2854) | (w7062 & w4684) | (w2854 & w4684);
assign w5797 = ~w9741 & w453;
assign w5798 = w9268 & w13142;
assign w5799 = ~w3036 & w8513;
assign w5800 = ~w12879 & w342;
assign w5801 = w10676 & w9805;
assign w5802 = ~w6309 & w4790;
assign w5803 = w4658 & w12899;
assign w5804 = ~w4632 & ~w10017;
assign w5805 = w11047 & w6960;
assign w5806 = w10094 | ~w9170;
assign w5807 = ~w10757 & w646;
assign w5808 = (w829 & w5559) | (w829 & w5187) | (w5559 & w5187);
assign w5809 = (~w11067 & w9656) | (~w11067 & w8815) | (w9656 & w8815);
assign w5810 = w12809 & w6689;
assign w5811 = (w9719 & w839) | (w9719 & w5023) | (w839 & w5023);
assign w5812 = ~w6116 & ~w13218;
assign w5813 = w7794 & ~w5276;
assign w5814 = ~w2361 & w13072;
assign w5815 = (w11655 & w12347) | (w11655 & ~w8228) | (w12347 & ~w8228);
assign w5816 = (w13395 & ~w9878) | (w13395 & w4180) | (~w9878 & w4180);
assign w5817 = ~w3175 & w8728;
assign w5818 = ~w4512 & w7088;
assign w5819 = w12691 & w7349;
assign w5820 = (w1164 & w4107) | (w1164 & w2167) | (w4107 & w2167);
assign w5821 = ~w11261 & w13809;
assign w5822 = w5257 & ~w3849;
assign w5823 = w10773 & w6438;
assign w5824 = w2486 & w9350;
assign w5825 = w6459 & w7295;
assign w5826 = ~w1563 & w40;
assign w5827 = ~w690 & w5421;
assign w5828 = (w353 & w3323) | (w353 & w11036) | (w3323 & w11036);
assign w5829 = (~w9305 & w13347) | (~w9305 & w10816) | (w13347 & w10816);
assign w5830 = ~w8782 & ~w3727;
assign w5831 = ~w5989 & ~w4915;
assign w5832 = w4213 & w3036;
assign w5833 = ~w7863 & ~w10193;
assign w5834 = ~w7040 & ~w4813;
assign w5835 = ~w11395 & ~w3158;
assign w5836 = ~w12129 & ~w2745;
assign w5837 = w8391 & w13124;
assign w5838 = w10676 & ~w6795;
assign w5839 = w13535 & w10557;
assign w5840 = ~w8006 & ~w7523;
assign w5841 = w11810 & w8900;
assign w5842 = ~w7305 & ~w3288;
assign w5843 = ~w3036 & w8047;
assign w5844 = (~w11228 & w1785) | (~w11228 & w4492) | (w1785 & w4492);
assign w5845 = ~w2121 & ~w1717;
assign w5846 = w7163 & ~w6062;
assign w5847 = ~b93 & a93;
assign w5848 = w798 & ~w4232;
assign w5849 = ~w9805 & ~w4288;
assign w5850 = w8742 & w5247;
assign w5851 = b2 & a2;
assign w5852 = ~w3610 & ~w13921;
assign w5853 = w9163 & ~w12343;
assign w5854 = w10822 & w9452;
assign w5855 = w12107 & w3427;
assign w5856 = (~w993 & w1295) | (~w993 & w288) | (w1295 & w288);
assign w5857 = ~w10855 & ~w5845;
assign w5858 = (w2670 & w13965) | (w2670 & w14477) | (w13965 & w14477);
assign w5859 = (w254 & w4769) | (w254 & w4181) | (w4769 & w4181);
assign w5860 = b60 & a60;
assign w5861 = (w5385 & w5139) | (w5385 & w6644) | (w5139 & w6644);
assign w5862 = w3885 & ~w11861;
assign w5863 = w13939 & w10156;
assign w5864 = w6425 & w12654;
assign w5865 = w1387 & w1027;
assign w5866 = ~w14302 & ~w7236;
assign w5867 = ~w367 & ~w13723;
assign w5868 = w13227 & w12673;
assign w5869 = w10880 & w4709;
assign w5870 = ~w4033 & ~w8768;
assign w5871 = w12724 & w14302;
assign w5872 = w6588 & ~b53;
assign w5873 = ~w12662 & w4787;
assign w5874 = ~w13677 & w3615;
assign w5875 = ~w1785 & w12339;
assign w5876 = ~w12635 & ~w8854;
assign w5877 = ~w10165 & w3364;
assign w5878 = ~w1540 & ~w757;
assign w5879 = (~w12464 & ~w820) | (~w12464 & w5037) | (~w820 & w5037);
assign w5880 = w12124 & ~w11126;
assign w5881 = w7135 & w13694;
assign w5882 = ~w607 & w10182;
assign w5883 = ~w11013 & ~w10182;
assign w5884 = ~w5214 & ~w1067;
assign w5885 = ~w8234 & w2933;
assign w5886 = w3963 & w6670;
assign w5887 = ~w4721 & ~w10308;
assign w5888 = w5207 | w5769;
assign w5889 = ~w183 & ~w2428;
assign w5890 = (~w8646 & w5374) | (~w8646 & w2987) | (w5374 & w2987);
assign w5891 = ~w2605 & ~w11606;
assign w5892 = w6087 & w661;
assign w5893 = w1909 & w14100;
assign w5894 = (w1274 & ~w12457) | (w1274 & w7552) | (~w12457 & w7552);
assign w5895 = (w9950 & w9534) | (w9950 & w1959) | (w9534 & w1959);
assign w5896 = ~w10939 & ~w14132;
assign w5897 = w7533 | w5414;
assign w5898 = ~w3633 & ~w13475;
assign w5899 = ~w5644 & w2841;
assign w5900 = ~w207 & ~w2356;
assign w5901 = w10384 | w12138;
assign w5902 = ~w3044 & ~w1212;
assign w5903 = w10072 & ~w3145;
assign w5904 = w4823 & w10290;
assign w5905 = (~w10719 & w11592) | (~w10719 & w5208) | (w11592 & w5208);
assign w5906 = w4359 & w14280;
assign w5907 = ~w14141 & w4106;
assign w5908 = (w3538 & w11579) | (w3538 & w3128) | (w11579 & w3128);
assign w5909 = ~w12980 & w2220;
assign w5910 = ~w2144 & w6928;
assign w5911 = w10036 & w7636;
assign w5912 = (~w9480 & w14569) | (~w9480 & w5080) | (w14569 & w5080);
assign w5913 = ~w12583 & w1476;
assign w5914 = (w6502 & w13416) | (w6502 & ~w922) | (w13416 & ~w922);
assign w5915 = (~w7058 & ~w11272) | (~w7058 & w795) | (~w11272 & w795);
assign w5916 = (~w40 & ~w14659) | (~w40 & w10868) | (~w14659 & w10868);
assign w5917 = (w7722 & w1817) | (w7722 & ~w3615) | (w1817 & ~w3615);
assign w5918 = (w7082 & w5684) | (w7082 & w5382) | (w5684 & w5382);
assign w5919 = ~w10997 & ~w6251;
assign w5920 = ~w2677 & w4316;
assign w5921 = ~w13222 & w1821;
assign w5922 = ~w13733 & w3025;
assign w5923 = ~w5974 & w2244;
assign w5924 = ~w12464 & w12856;
assign w5925 = (w12460 & ~w3671) | (w12460 & w4732) | (~w3671 & w4732);
assign w5926 = (~w10272 & ~w4656) | (~w10272 & w3289) | (~w4656 & w3289);
assign w5927 = ~w7726 & w1919;
assign w5928 = ~w3710 & ~w9129;
assign w5929 = ~w491 & ~w11002;
assign w5930 = w6972 & ~w5810;
assign w5931 = (w1939 & w14084) | (w1939 & w9303) | (w14084 & w9303);
assign w5932 = ~w14227 & ~w3767;
assign w5933 = (w6617 & ~w12271) | (w6617 & w12616) | (~w12271 & w12616);
assign w5934 = ~w607 & ~w3727;
assign w5935 = w3944 & ~w7686;
assign w5936 = ~b24 & ~a24;
assign w5937 = ~w10354 & ~w13900;
assign w5938 = w2101 & ~w10182;
assign w5939 = (w10045 & ~w12614) | (w10045 & w7946) | (~w12614 & w7946);
assign w5940 = (~w5952 & ~w568) | (~w5952 & w6146) | (~w568 & w6146);
assign w5941 = w11925 & w7260;
assign w5942 = ~w7782 & w4414;
assign w5943 = w4965 & w1678;
assign w5944 = ~w10674 & w12582;
assign w5945 = ~w5785 & ~w235;
assign w5946 = ~w7013 & ~w2751;
assign w5947 = ~w6783 & w1692;
assign w5948 = b120 & a120;
assign w5949 = w7794 & w1874;
assign w5950 = ~w4504 & w7577;
assign w5951 = ~w11566 & w2598;
assign w5952 = ~w8778 & ~w12951;
assign w5953 = w1871 & w10486;
assign w5954 = ~w3015 & w5009;
assign w5955 = w12716 & w1217;
assign w5956 = ~w1900 & w11495;
assign w5957 = (w11613 & w6299) | (w11613 & w8018) | (w6299 & w8018);
assign w5958 = (~w5952 & w7876) | (~w5952 & w4698) | (w7876 & w4698);
assign w5959 = (w8827 & w13462) | (w8827 & w549) | (w13462 & w549);
assign w5960 = (w3963 & ~w5489) | (w3963 & w12534) | (~w5489 & w12534);
assign w5961 = (~w3537 & w692) | (~w3537 & w3757) | (w692 & w3757);
assign w5962 = ~w5453 & w2976;
assign w5963 = (~w4918 & w11167) | (~w4918 & w10891) | (w11167 & w10891);
assign w5964 = ~w1171 & w621;
assign w5965 = w14295 & ~w8649;
assign w5966 = (w12656 & w8665) | (w12656 & ~w6750) | (w8665 & ~w6750);
assign w5967 = ~w7880 & w14305;
assign w5968 = w9776 & ~w1623;
assign w5969 = w8802 & w5665;
assign w5970 = (w2701 & w3586) | (w2701 & w2802) | (w3586 & w2802);
assign w5971 = ~w9012 & w3426;
assign w5972 = (~w6218 & ~w5490) | (~w6218 & w13110) | (~w5490 & w13110);
assign w5973 = w5306 & w7454;
assign w5974 = ~w5736 & ~w9889;
assign w5975 = ~w4571 & ~w679;
assign w5976 = ~w12749 & ~w4385;
assign w5977 = (~w10299 & w9352) | (~w10299 & w2465) | (w9352 & w2465);
assign w5978 = w4193 & w3017;
assign w5979 = ~w383 & ~w9479;
assign w5980 = w1563 & w13531;
assign w5981 = w12483 & ~w10800;
assign w5982 = w3550 & w8175;
assign w5983 = ~w11031 & ~w11693;
assign w5984 = ~w3632 & ~w5664;
assign w5985 = w4573 & ~w10379;
assign w5986 = w4836 & w5227;
assign w5987 = w11031 & w9482;
assign w5988 = w9424 & w12176;
assign w5989 = ~w4700 & w2729;
assign w5990 = (w694 & w10958) | (w694 & w9721) | (w10958 & w9721);
assign w5991 = (w9512 & w9668) | (w9512 & ~w4987) | (w9668 & ~w4987);
assign w5992 = ~w347 & ~w341;
assign w5993 = w4379 & w7277;
assign w5994 = w13189 & ~w10757;
assign w5995 = w1535 & w1246;
assign w5996 = (~w14486 & w6699) | (~w14486 & w9862) | (w6699 & w9862);
assign w5997 = (~w2844 & ~w5925) | (~w2844 & w8658) | (~w5925 & w8658);
assign w5998 = ~w3751 & w13227;
assign w5999 = ~w185 & w7437;
assign w6000 = ~w4548 & ~w10869;
assign w6001 = w5505 & w12588;
assign w6002 = (w6637 & w2647) | (w6637 & w10337) | (w2647 & w10337);
assign w6003 = ~w10130 & ~w3460;
assign w6004 = w3914 & w10997;
assign w6005 = ~w668 & w11463;
assign w6006 = (w3671 & w12319) | (w3671 & w6142) | (w12319 & w6142);
assign w6007 = (w12170 & w4158) | (w12170 & w4258) | (w4158 & w4258);
assign w6008 = (w13924 & ~w12614) | (w13924 & w709) | (~w12614 & w709);
assign w6009 = (~w12406 & w1757) | (~w12406 & w9691) | (w1757 & w9691);
assign w6010 = w2486 & w1873;
assign w6011 = (~w14455 & ~w8337) | (~w14455 & w1583) | (~w8337 & w1583);
assign w6012 = (~w11810 & w1166) | (~w11810 & w9430) | (w1166 & w9430);
assign w6013 = (w8135 & w14416) | (w8135 & ~w5595) | (w14416 & ~w5595);
assign w6014 = w9015 & w5865;
assign w6015 = w2470 | ~w10590;
assign w6016 = (~w3759 & w7362) | (~w3759 & w9106) | (w7362 & w9106);
assign w6017 = w419 & ~w6265;
assign w6018 = ~w9747 & w7981;
assign w6019 = w2975 & w11970;
assign w6020 = w3738 & w7458;
assign w6021 = ~w6230 & ~w14642;
assign w6022 = ~w1785 & w8643;
assign w6023 = (w2979 & w6780) | (w2979 & ~w9749) | (w6780 & ~w9749);
assign w6024 = ~w3067 & w13162;
assign w6025 = (w878 & ~w6321) | (w878 & w10288) | (~w6321 & w10288);
assign w6026 = (w10795 & w10550) | (w10795 & w975) | (w10550 & w975);
assign w6027 = ~w5522 & ~w646;
assign w6028 = (~w2670 & w7677) | (~w2670 & w13362) | (w7677 & w13362);
assign w6029 = ~w491 & ~w7695;
assign w6030 = (w6195 & w1342) | (w6195 & w12376) | (w1342 & w12376);
assign w6031 = (w5601 & w14328) | (w5601 & w3954) | (w14328 & w3954);
assign w6032 = (w6427 & w10570) | (w6427 & w94) | (w10570 & w94);
assign w6033 = (~w3631 & w7147) | (~w3631 & w5293) | (w7147 & w5293);
assign w6034 = w13526 & w9748;
assign w6035 = w7857 & ~w6164;
assign w6036 = ~w9653 & w6425;
assign w6037 = ~w1840 & ~w560;
assign w6038 = ~w12609 & w9263;
assign w6039 = w10526 & ~w7325;
assign w6040 = (~w894 & w9012) | (~w894 & w3692) | (w9012 & w3692);
assign w6041 = (~w6281 & w4503) | (~w6281 & w11535) | (w4503 & w11535);
assign w6042 = ~w1415 & ~w6468;
assign w6043 = (w13685 & w5500) | (w13685 & w6030) | (w5500 & w6030);
assign w6044 = (~w254 & w8331) | (~w254 & w2632) | (w8331 & w2632);
assign w6045 = ~w8100 & ~w9672;
assign w6046 = ~w13063 & w8109;
assign w6047 = ~w3694 & ~w1540;
assign w6048 = w8512 & ~w12398;
assign w6049 = ~w4512 & w10024;
assign w6050 = w11779 & ~w4424;
assign w6051 = ~w13528 & w13019;
assign w6052 = w13854 & ~w9748;
assign w6053 = w2283 & w5834;
assign w6054 = (w8713 & w9809) | (w8713 & w2472) | (w9809 & w2472);
assign w6055 = ~w1166 & w9015;
assign w6056 = (~w11091 & w7028) | (~w11091 & w10413) | (w7028 & w10413);
assign w6057 = (~w10722 & w12626) | (~w10722 & w12106) | (w12626 & w12106);
assign w6058 = (~w2386 & w9243) | (~w2386 & w332) | (w9243 & w332);
assign w6059 = (~w10514 & w922) | (~w10514 & w12248) | (w922 & w12248);
assign w6060 = (w1619 & w14613) | (w1619 & w4354) | (w14613 & w4354);
assign w6061 = w884 & ~w12943;
assign w6062 = ~w6113 & w1263;
assign w6063 = (~w6929 & w254) | (~w6929 & w973) | (w254 & w973);
assign w6064 = w5842 & ~w794;
assign w6065 = ~w5702 & w800;
assign w6066 = w6080 & ~w7335;
assign w6067 = ~w7670 & ~w13862;
assign w6068 = ~w4270 & w506;
assign w6069 = ~w142 & ~w8396;
assign w6070 = (~w14463 & w4510) | (~w14463 & w7891) | (w4510 & w7891);
assign w6071 = w4573 & ~w10286;
assign w6072 = ~w13730 & ~w13963;
assign w6073 = ~w12569 & w10295;
assign w6074 = (w1362 & w5295) | (w1362 & w3646) | (w5295 & w3646);
assign w6075 = ~w2252 & w13785;
assign w6076 = w1828 & w14532;
assign w6077 = ~w8367 & w10605;
assign w6078 = (w2608 & w3043) | (w2608 & w1525) | (w3043 & w1525);
assign w6079 = (w346 & w7318) | (w346 & w9403) | (w7318 & w9403);
assign w6080 = ~b103 & ~a103;
assign w6081 = ~w11665 & w2434;
assign w6082 = w4254 & ~w13221;
assign w6083 = w5192 & ~w12110;
assign w6084 = w6391 & w6703;
assign w6085 = ~w142 & ~w13937;
assign w6086 = ~w9541 & ~w3439;
assign w6087 = ~w4782 & w4913;
assign w6088 = (w2620 & w5215) | (w2620 & ~w318) | (w5215 & ~w318);
assign w6089 = ~w64 & w9273;
assign w6090 = ~w11204 & ~w12002;
assign w6091 = (w3853 & w14604) | (w3853 & ~w11915) | (w14604 & ~w11915);
assign w6092 = w5944 & w12467;
assign w6093 = w9092 & w13444;
assign w6094 = w4433 & w11637;
assign w6095 = w14554 & w6427;
assign w6096 = w3012 & w1513;
assign w6097 = ~w5072 & ~w4743;
assign w6098 = (~w13462 & w8331) | (~w13462 & w8147) | (w8331 & w8147);
assign w6099 = ~w5747 & ~w13681;
assign w6100 = w9622 & ~w3687;
assign w6101 = w7019 & w2163;
assign w6102 = ~w3355 & ~w12521;
assign w6103 = ~w3218 & ~w14355;
assign w6104 = ~w13312 & w12392;
assign w6105 = w13606 & ~w3990;
assign w6106 = ~w8586 & ~w6669;
assign w6107 = (w7727 & w5888) | (w7727 & w8406) | (w5888 & w8406);
assign w6108 = ~w4780 & ~w10423;
assign w6109 = (~w14600 & w7225) | (~w14600 & w2062) | (w7225 & w2062);
assign w6110 = w7914 & w10414;
assign w6111 = ~w8200 & w5930;
assign w6112 = w7365 & ~w1096;
assign w6113 = ~w10704 & ~w13873;
assign w6114 = w10241 & ~w12480;
assign w6115 = ~w8791 & w7772;
assign w6116 = (w11634 & w5726) | (w11634 & w5042) | (w5726 & w5042);
assign w6117 = (~w2493 & ~w4424) | (~w2493 & ~w5161) | (~w4424 & ~w5161);
assign w6118 = ~w11934 & ~w10324;
assign w6119 = ~w6750 & ~w14088;
assign w6120 = ~w4504 & w4617;
assign w6121 = (~w2317 & w576) | (~w2317 & w8074) | (w576 & w8074);
assign w6122 = w607 & w9211;
assign w6123 = (w171 & w9819) | (w171 & w1896) | (w9819 & w1896);
assign w6124 = w7864 & ~w5862;
assign w6125 = (w719 & w4506) | (w719 & w9843) | (w4506 & w9843);
assign w6126 = ~w3963 & w3503;
assign w6127 = ~w8332 & ~w1074;
assign w6128 = w12315 & ~w7022;
assign w6129 = (w12776 & w939) | (w12776 & w6314) | (w939 & w6314);
assign w6130 = (w9753 & w6046) | (w9753 & w8577) | (w6046 & w8577);
assign w6131 = w3209 & w9226;
assign w6132 = (w6267 & w2953) | (w6267 & w14534) | (w2953 & w14534);
assign w6133 = w7529 & ~w963;
assign w6134 = ~w5522 & ~w12642;
assign w6135 = ~b102 & ~a102;
assign w6136 = w5177 & w2680;
assign w6137 = w3828 & ~w285;
assign w6138 = (~w8431 & w2698) | (~w8431 & w7526) | (w2698 & w7526);
assign w6139 = w8836 & ~b53;
assign w6140 = ~w13908 & w6900;
assign w6141 = (w5664 & w2326) | (w5664 & w13016) | (w2326 & w13016);
assign w6142 = ~w6949 & w3671;
assign w6143 = w9923 & ~w5058;
assign w6144 = w4033 & ~w11117;
assign w6145 = ~w11013 & ~w1838;
assign w6146 = ~w3289 | ~w7999;
assign w6147 = w3502 & w8900;
assign w6148 = w10301 | ~w10116;
assign w6149 = (w9510 & w5119) | (w9510 & w9721) | (w5119 & w9721);
assign w6150 = ~w12810 & w11045;
assign w6151 = ~w5867 & ~w5568;
assign w6152 = (~w5212 & w562) | (~w5212 & w1478) | (w562 & w1478);
assign w6153 = w8073 & w1220;
assign w6154 = ~w3195 & ~w3497;
assign w6155 = (w803 & ~w6113) | (w803 & w6921) | (~w6113 & w6921);
assign w6156 = w8018 & w12525;
assign w6157 = w5294 & ~w5005;
assign w6158 = ~w14302 & w8390;
assign w6159 = ~w11559 & ~w498;
assign w6160 = (w11472 & w10905) | (w11472 & w9928) | (w10905 & w9928);
assign w6161 = ~w309 & ~w7296;
assign w6162 = ~w8449 & w10083;
assign w6163 = w607 & w12460;
assign w6164 = w6135 & ~w3963;
assign w6165 = w13374 & ~w11179;
assign w6166 = ~w4447 & ~w1732;
assign w6167 = ~w6638 & ~w9191;
assign w6168 = (~w13349 & w7324) | (~w13349 & w12350) | (w7324 & w12350);
assign w6169 = ~w6800 & w7886;
assign w6170 = (~w9949 & w10781) | (~w9949 & w7947) | (w10781 & w7947);
assign w6171 = w6651 & ~w10143;
assign w6172 = w558 & w11250;
assign w6173 = ~w1015 & ~w14074;
assign w6174 = w3208 & w8008;
assign w6175 = ~w2332 & w12060;
assign w6176 = ~w12908 & ~w5754;
assign w6177 = ~w1949 & ~w2270;
assign w6178 = (~w7488 & w11365) | (~w7488 & w1707) | (w11365 & w1707);
assign w6179 = (~w4017 & w7782) | (~w4017 & w4470) | (w7782 & w4470);
assign w6180 = (w11753 & w6243) | (w11753 & w217) | (w6243 & w217);
assign w6181 = (w10500 & w3070) | (w10500 & w7629) | (w3070 & w7629);
assign w6182 = w9055 & ~w13885;
assign w6183 = (~w6802 & w12537) | (~w6802 & w9928) | (w12537 & w9928);
assign w6184 = ~w7782 & w11112;
assign w6185 = ~w12516 & w930;
assign w6186 = w8832 & ~w1231;
assign w6187 = (w9181 & ~w1874) | (w9181 & w6564) | (~w1874 & w6564);
assign w6188 = w1597 & ~w822;
assign w6189 = ~w14337 & w10048;
assign w6190 = b117 & a117;
assign w6191 = ~w1474 & w2729;
assign w6192 = ~w6700 & w4021;
assign w6193 = w5522 & ~w11861;
assign w6194 = ~w5223 & ~w4883;
assign w6195 = (w13334 & w6457) | (w13334 & ~w9749) | (w6457 & ~w9749);
assign w6196 = w3435 & ~w5321;
assign w6197 = ~w10509 & ~w12740;
assign w6198 = ~w475 & w13839;
assign w6199 = ~w11775 & ~w412;
assign w6200 = (w12062 & w3488) | (w12062 & w7200) | (w3488 & w7200);
assign w6201 = ~w4881 & w235;
assign w6202 = ~w11959 & ~w2335;
assign w6203 = w153 & ~w4169;
assign w6204 = w3401 & ~w3904;
assign w6205 = ~w7488 & w6139;
assign w6206 = (b53 & w1840) | (b53 & w3098) | (w1840 & w3098);
assign w6207 = (~w5385 & w3559) | (~w5385 & w13489) | (w3559 & w13489);
assign w6208 = ~w11583 & w499;
assign w6209 = ~w3885 & w325;
assign w6210 = (w6107 & w1473) | (w6107 & ~w9591) | (w1473 & ~w9591);
assign w6211 = ~w11793 & w14118;
assign w6212 = b53 & w8836;
assign w6213 = ~w10205 & ~w12991;
assign w6214 = w2332 & ~w13565;
assign w6215 = (w8018 & w1519) | (w8018 & w11937) | (w1519 & w11937);
assign w6216 = ~w5867 & w13733;
assign w6217 = ~w6972 & ~w8603;
assign w6218 = ~w8171 & w11264;
assign w6219 = ~w9244 & ~w9465;
assign w6220 = w3587 & ~w11117;
assign w6221 = (w12786 & w11966) | (w12786 & w4131) | (w11966 & w4131);
assign w6222 = (w13548 & w2612) | (w13548 & ~w12376) | (w2612 & ~w12376);
assign w6223 = (~w2386 & w592) | (~w2386 & ~w10656) | (w592 & ~w10656);
assign w6224 = ~w3886 & w6607;
assign w6225 = (~w7490 & w9298) | (~w7490 & w4222) | (w9298 & w4222);
assign w6226 = (w1114 & w13462) | (w1114 & w6730) | (w13462 & w6730);
assign w6227 = w12569 & ~w12170;
assign w6228 = ~w10225 & w422;
assign w6229 = (~w6567 & w6013) | (~w6567 & w10233) | (w6013 & w10233);
assign w6230 = w14293 & ~w2804;
assign w6231 = ~w1712 & ~w12331;
assign w6232 = (w2655 & w10097) | (w2655 & w7989) | (w10097 & w7989);
assign w6233 = w1096 & ~w8389;
assign w6234 = (~w3885 & w4178) | (~w3885 & w1557) | (w4178 & w1557);
assign w6235 = ~w7244 & ~w2729;
assign w6236 = (~w5845 & w14485) | (~w5845 & w8578) | (w14485 & w8578);
assign w6237 = (~w13445 & w13462) | (~w13445 & w10236) | (w13462 & w10236);
assign w6238 = (w6426 & w14095) | (w6426 & w1818) | (w14095 & w1818);
assign w6239 = ~w7256 & w6845;
assign w6240 = (~w2850 & ~w9715) | (~w2850 & w7811) | (~w9715 & w7811);
assign w6241 = w638 & w8878;
assign w6242 = ~w12569 & ~w3007;
assign w6243 = (~w10016 & ~w5242) | (~w10016 & w6155) | (~w5242 & w6155);
assign w6244 = w11488 & w8389;
assign w6245 = (~w14664 & w718) | (~w14664 & w3882) | (w718 & w3882);
assign w6246 = (w11734 & w5438) | (w11734 & w11857) | (w5438 & w11857);
assign w6247 = w3751 & ~w2951;
assign w6248 = (~w8104 & w14320) | (~w8104 & w12399) | (w14320 & w12399);
assign w6249 = w9016 & w13672;
assign w6250 = ~w1706 & ~w10846;
assign w6251 = w7085 & w10042;
assign w6252 = ~w5852 & ~w11068;
assign w6253 = ~w7808 & w10182;
assign w6254 = ~w12463 & w4453;
assign w6255 = (w11817 & w2317) | (w11817 & w11344) | (w2317 & w11344);
assign w6256 = ~w2144 & w5520;
assign w6257 = w2729 & ~w4447;
assign w6258 = w3175 & w3098;
assign w6259 = ~w7132 & w11251;
assign w6260 = (w10423 & ~w697) | (w10423 & w4009) | (~w697 & w4009);
assign w6261 = (~w7488 & w10969) | (~w7488 & w1515) | (w10969 & w1515);
assign w6262 = (w12088 & w1482) | (w12088 & w12699) | (w1482 & w12699);
assign w6263 = w12654 & w6636;
assign w6264 = (~w2939 & w9571) | (~w2939 & w14438) | (w9571 & w14438);
assign w6265 = w7373 & w7796;
assign w6266 = w7455 & w13544;
assign w6267 = (~w3587 & w6128) | (~w3587 & w7597) | (w6128 & w7597);
assign w6268 = (w9316 & w14460) | (w9316 & w8864) | (w14460 & w8864);
assign w6269 = (w7455 & w4512) | (w7455 & w5745) | (w4512 & w5745);
assign w6270 = (w6939 & w6319) | (w6939 & w12742) | (w6319 & w12742);
assign w6271 = ~w7782 & w311;
assign w6272 = ~w9643 & w12369;
assign w6273 = ~w7276 & ~w3427;
assign w6274 = w11492 & ~w1195;
assign w6275 = w1906 & ~w9902;
assign w6276 = (~w4709 & ~w7538) | (~w4709 & ~w7240) | (~w7538 & ~w7240);
assign w6277 = ~w13526 & w5626;
assign w6278 = w6697 & ~w12914;
assign w6279 = ~w11815 & w1001;
assign w6280 = w2707 & ~w7369;
assign w6281 = ~b84 & ~a84;
assign w6282 = w8721 & w11676;
assign w6283 = ~w12271 & w9805;
assign w6284 = (w7240 & w9018) | (w7240 & w3) | (w9018 & w3);
assign w6285 = w5768 & w13570;
assign w6286 = w607 & ~w9296;
assign w6287 = w4207 & w6213;
assign w6288 = w10045 & ~w2270;
assign w6289 = (~w14040 & ~w5946) | (~w14040 & ~w8768) | (~w5946 & ~w8768);
assign w6290 = (w5626 & w12420) | (w5626 & w14432) | (w12420 & w14432);
assign w6291 = w2377 & w5046;
assign w6292 = ~w2335 & ~w9833;
assign w6293 = w3982 & ~w3568;
assign w6294 = w1015 & ~w13521;
assign w6295 = (w5952 & w567) | (w5952 & w6091) | (w567 & w6091);
assign w6296 = ~w4266 & w11592;
assign w6297 = w7369 & w5282;
assign w6298 = ~w607 & ~w7794;
assign w6299 = w3121 & w11613;
assign w6300 = ~w4158 & w12379;
assign w6301 = (~w8035 & ~w1699) | (~w8035 & w14505) | (~w1699 & w14505);
assign w6302 = w3957 & ~w8636;
assign w6303 = (w3638 & w11046) | (w3638 & ~w12376) | (w11046 & ~w12376);
assign w6304 = ~w4836 & w6542;
assign w6305 = w4142 & w3042;
assign w6306 = (w606 & w5967) | (w606 & w10476) | (w5967 & w10476);
assign w6307 = ~w12128 | w8326;
assign w6308 = (w8551 & ~w2167) | (w8551 & w8282) | (~w2167 & w8282);
assign w6309 = w2544 & ~w7331;
assign w6310 = w2773 & w6883;
assign w6311 = (w4442 & ~w14042) | (w4442 & w9293) | (~w14042 & w9293);
assign w6312 = ~w1712 & w3529;
assign w6313 = (~w2870 & w5969) | (~w2870 & ~w13973) | (w5969 & ~w13973);
assign w6314 = (w2309 & w14442) | (w2309 & w280) | (w14442 & w280);
assign w6315 = ~w7431 & ~w5094;
assign w6316 = ~w1563 & w6014;
assign w6317 = ~w7722 & w9694;
assign w6318 = w11500 & w7715;
assign w6319 = ~w11064 & ~w10365;
assign w6320 = (w5342 & w8604) | (w5342 & w6756) | (w8604 & w6756);
assign w6321 = ~w11021 & w3152;
assign w6322 = w6502 & ~w10477;
assign w6323 = w3730 & w2077;
assign w6324 = w8183 & w3727;
assign w6325 = w12460 & w2522;
assign w6326 = ~w13540 & w7914;
assign w6327 = w12041 & w9227;
assign w6328 = ~w6235 & ~w4296;
assign w6329 = (w11908 & w6762) | (w11908 & w12495) | (w6762 & w12495);
assign w6330 = w12482 & w9949;
assign w6331 = (w14593 & w9271) | (w14593 & w4250) | (w9271 & w4250);
assign w6332 = (w12799 & w9112) | (w12799 & w1551) | (w9112 & w1551);
assign w6333 = ~w5052 & ~w7066;
assign w6334 = w7276 & ~w8459;
assign w6335 = w14325 & w3594;
assign w6336 = ~w6262 & w13826;
assign w6337 = ~w11899 & w9952;
assign w6338 = ~w7898 & ~w13901;
assign w6339 = w607 & w2701;
assign w6340 = w6932 & w499;
assign w6341 = (~w8973 & w6720) | (~w8973 & w7155) | (w6720 & w7155);
assign w6342 = (~w12642 & w8715) | (~w12642 & w2758) | (w8715 & w2758);
assign w6343 = w9813 & w12461;
assign w6344 = w1116 & ~w5813;
assign w6345 = ~w12482 & ~w2951;
assign w6346 = ~w12972 & w14206;
assign w6347 = (w1208 & w53) | (w1208 & ~w8444) | (w53 & ~w8444);
assign w6348 = ~w2656 & w12170;
assign w6349 = w5213 & w2933;
assign w6350 = (w8977 & w13152) | (w8977 & w487) | (w13152 & w487);
assign w6351 = (~w5664 & ~w3198) | (~w5664 & w4008) | (~w3198 & w4008);
assign w6352 = ~w14141 & w4619;
assign w6353 = ~w10549 & ~w2896;
assign w6354 = ~w3484 & w6267;
assign w6355 = w1535 & ~w14173;
assign w6356 = (w2040 & w14221) | (w2040 & ~w4754) | (w14221 & ~w4754);
assign w6357 = w13297 & ~w12506;
assign w6358 = ~w7906 & ~w3851;
assign w6359 = w11395 & ~w6572;
assign w6360 = (~w14512 & w2175) | (~w14512 & w458) | (w2175 & w458);
assign w6361 = ~w6436 & ~w14133;
assign w6362 = (~w13324 & w2470) | (~w13324 & w4079) | (w2470 & w4079);
assign w6363 = ~w3699 & ~w1692;
assign w6364 = ~w894 & ~w10295;
assign w6365 = ~w2129 & w11470;
assign w6366 = (w8367 & w7482) | (w8367 & w4418) | (w7482 & w4418);
assign w6367 = (w3128 & w13683) | (w3128 & ~w10994) | (w13683 & ~w10994);
assign w6368 = (w3192 & w14306) | (w3192 & w9770) | (w14306 & w9770);
assign w6369 = (~w12776 & w13447) | (~w12776 & w6937) | (w13447 & w6937);
assign w6370 = w7844 & w281;
assign w6371 = (w6572 & w7782) | (w6572 & w10667) | (w7782 & w10667);
assign w6372 = (~w5537 & w7375) | (~w5537 & w9763) | (w7375 & w9763);
assign w6373 = ~w10483 & ~w11732;
assign w6374 = w3135 & ~w7305;
assign w6375 = ~w10517 & w2101;
assign w6376 = (~w12055 & w8108) | (~w12055 & w13006) | (w8108 & w13006);
assign w6377 = ~w12915 & ~w1692;
assign w6378 = w5912 & w13638;
assign w6379 = w473 & w1692;
assign w6380 = (w659 & w3505) | (w659 & w9707) | (w3505 & w9707);
assign w6381 = w2872 & w9183;
assign w6382 = (~w227 & ~w9989) | (~w227 & ~w14514) | (~w9989 & ~w14514);
assign w6383 = w7051 & w7337;
assign w6384 = w12330 & ~w2603;
assign w6385 = ~cin & ~w9546;
assign w6386 = ~w569 & w11187;
assign w6387 = ~w3002 & ~w3269;
assign w6388 = (~w6802 & w8020) | (~w6802 & w11214) | (w8020 & w11214);
assign w6389 = w8299 & w13064;
assign w6390 = (w11395 & w8937) | (w11395 & w3470) | (w8937 & w3470);
assign w6391 = ~w607 & ~w14276;
assign w6392 = w7498 & ~w10052;
assign w6393 = ~w7794 & w6861;
assign w6394 = ~w14249 & ~w6716;
assign w6395 = (w5002 & ~w7811) | (w5002 & w14487) | (~w7811 & w14487);
assign w6396 = ~w3252 & ~w13155;
assign w6397 = (w2038 & ~w8655) | (w2038 & w13044) | (~w8655 & w13044);
assign w6398 = w12814 & w859;
assign w6399 = w4605 & ~w9493;
assign w6400 = (w11712 & w7842) | (w11712 & w9826) | (w7842 & w9826);
assign w6401 = (~w11487 & w3439) | (~w11487 & ~w3187) | (w3439 & ~w3187);
assign w6402 = (w9831 & ~w630) | (w9831 & ~w7592) | (~w630 & ~w7592);
assign w6403 = w10054 & ~w214;
assign w6404 = ~w8059 & ~w5529;
assign w6405 = (w5406 & w7423) | (w5406 & w2186) | (w7423 & w2186);
assign w6406 = ~w9412 & ~w2762;
assign w6407 = ~w2381 & w1919;
assign w6408 = ~w10435 & w4024;
assign w6409 = ~w12048 & w3544;
assign w6410 = (w10116 & w5841) | (w10116 & w14266) | (w5841 & w14266);
assign w6411 = (~w9012 & w4427) | (~w9012 & w8453) | (w4427 & w8453);
assign w6412 = ~w8380 & ~w9226;
assign w6413 = ~w6147 & w779;
assign w6414 = (~w11608 & ~w5771) | (~w11608 & w2294) | (~w5771 & w2294);
assign w6415 = ~w5702 & w4789;
assign w6416 = (~w9747 & w11917) | (~w9747 & w7273) | (w11917 & w7273);
assign w6417 = ~w8937 & w14230;
assign w6418 = w7794 & w5564;
assign w6419 = (w9012 & w12823) | (w9012 & w10332) | (w12823 & w10332);
assign w6420 = ~w10486 & w3730;
assign w6421 = ~w5406 & ~w4467;
assign w6422 = w4032 & w829;
assign w6423 = (~w5727 & w5170) | (~w5727 & w12999) | (w5170 & w12999);
assign w6424 = ~w12050 & ~w7627;
assign w6425 = w2978 & w4217;
assign w6426 = (w8327 & w6057) | (w8327 & w1853) | (w6057 & w1853);
assign w6427 = w9032 & w13544;
assign w6428 = (w12460 & w1712) | (w12460 & w4732) | (w1712 & w4732);
assign w6429 = w11810 & w8769;
assign w6430 = (w4364 & ~w9119) | (w4364 & w3839) | (~w9119 & w3839);
assign w6431 = ~w11031 & ~w4632;
assign w6432 = ~w6676 & w1184;
assign w6433 = b24 & a24;
assign w6434 = w4349 & ~w8809;
assign w6435 = w10514 & ~w4190;
assign w6436 = ~w11745 & ~w12481;
assign w6437 = (~w14048 & ~w4317) | (~w14048 & ~w11559) | (~w4317 & ~w11559);
assign w6438 = w7719 & ~w3427;
assign w6439 = (~w7369 & w6668) | (~w7369 & w7643) | (w6668 & w7643);
assign w6440 = ~w5959 & w12017;
assign w6441 = (w4375 & w10778) | (w4375 & w1383) | (w10778 & w1383);
assign w6442 = ~b26 & ~a26;
assign w6443 = w1500 & w3720;
assign w6444 = ~w1785 & w8701;
assign w6445 = w10686 & ~w12634;
assign w6446 = ~w751 & ~w14065;
assign w6447 = w3215 & w5247;
assign w6448 = (w13462 & w12724) | (w13462 & w5871) | (w12724 & w5871);
assign w6449 = ~w11475 & w6176;
assign w6450 = ~w13587 & w4837;
assign w6451 = ~w5867 & w2335;
assign w6452 = (w6885 & ~w8097) | (w6885 & w2248) | (~w8097 & w2248);
assign w6453 = (~w8253 & ~w3427) | (~w8253 & w3987) | (~w3427 & w3987);
assign w6454 = w7794 & w7881;
assign w6455 = ~w11940 & w5247;
assign w6456 = w14302 & ~w8573;
assign w6457 = (~w2599 & w5161) | (~w2599 & w1157) | (w5161 & w1157);
assign w6458 = (w1849 & w9681) | (w1849 & w5138) | (w9681 & w5138);
assign w6459 = ~w2202 & ~w12429;
assign w6460 = (w1849 & w13787) | (w1849 & w3831) | (w13787 & w3831);
assign w6461 = ~w10252 & ~w9287;
assign w6462 = (w7047 & ~w6753) | (w7047 & ~w10123) | (~w6753 & ~w10123);
assign w6463 = ~w1080 & w7480;
assign w6464 = ~w4729 & ~w3241;
assign w6465 = ~w1166 & ~w14070;
assign w6466 = ~w9480 & ~w7000;
assign w6467 = ~w13688 & w9059;
assign w6468 = (~w8573 & w2463) | (~w8573 & w6456) | (w2463 & w6456);
assign w6469 = ~w14633 & ~w10295;
assign w6470 = w11431 & w1679;
assign w6471 = ~w11429 & w9953;
assign w6472 = ~w5294 & ~w13940;
assign w6473 = (~w852 & w621) | (~w852 & w8635) | (w621 & w8635);
assign w6474 = w13306 & ~w9788;
assign w6475 = (~w8052 & w7781) | (~w8052 & w10063) | (w7781 & w10063);
assign w6476 = (~w10435 & w14358) | (~w10435 & w10208) | (w14358 & w10208);
assign w6477 = ~w11956 & w9551;
assign w6478 = w11346 & w2906;
assign w6479 = ~w12759 & w3126;
assign w6480 = (w5697 & w3676) | (w5697 & w12154) | (w3676 & w12154);
assign w6481 = w1550 & w3267;
assign w6482 = (~w7912 & w5956) | (~w7912 & w14063) | (w5956 & w14063);
assign w6483 = ~w71 & w6661;
assign w6484 = (w9021 & w4565) | (w9021 & w11339) | (w4565 & w11339);
assign w6485 = w3717 & w9265;
assign w6486 = w10993 & ~w499;
assign w6487 = ~w13282 & w9040;
assign w6488 = w9145 & ~w3427;
assign w6489 = ~w6398 & w7624;
assign w6490 = w9509 & ~w4868;
assign w6491 = w4989 & ~w3317;
assign w6492 = ~w8013 & ~w8370;
assign w6493 = w956 & w14249;
assign w6494 = (w9981 & w13076) | (w9981 & w4321) | (w13076 & w4321);
assign w6495 = w309 & ~w1016;
assign w6496 = (~w10272 & w14289) | (~w10272 & w2048) | (w14289 & w2048);
assign w6497 = ~w2569 & w11817;
assign w6498 = (~w7305 & w3135) | (~w7305 & ~w5282) | (w3135 & ~w5282);
assign w6499 = w12240 & w6889;
assign w6500 = ~w3251 & ~w8280;
assign w6501 = w1565 & w2735;
assign w6502 = w4017 & w1016;
assign w6503 = w10014 & w825;
assign w6504 = ~w2634 & ~w5631;
assign w6505 = (~w12429 & w2605) | (~w12429 & w6775) | (w2605 & w6775);
assign w6506 = ~w5852 & ~w10435;
assign w6507 = (~w4030 & w9571) | (~w4030 & w14438) | (w9571 & w14438);
assign w6508 = (~w6755 & w11803) | (~w6755 & w1925) | (w11803 & w1925);
assign w6509 = ~w14437 & ~w4774;
assign w6510 = w10271 & ~w1970;
assign w6511 = ~w1805 & w4541;
assign w6512 = (w13834 & w14347) | (w13834 & w8923) | (w14347 & w8923);
assign w6513 = ~w9912 & w5083;
assign w6514 = ~w4050 & w5921;
assign w6515 = ~w3878 & ~w12986;
assign w6516 = (w5406 & w5702) | (w5406 & w12686) | (w5702 & w12686);
assign w6517 = w2941 & w11764;
assign w6518 = (~w5406 & w12614) | (~w5406 & w8442) | (w12614 & w8442);
assign w6519 = (~w4127 & w13587) | (~w4127 & w8968) | (w13587 & w8968);
assign w6520 = w11117 & w9015;
assign w6521 = ~w10980 & ~w11166;
assign w6522 = ~w449 & ~w2044;
assign w6523 = w1840 & w829;
assign w6524 = (w12817 & w7268) | (w12817 & w1725) | (w7268 & w1725);
assign w6525 = (~w5428 & ~w7282) | (~w5428 & w14111) | (~w7282 & w14111);
assign w6526 = (~w3460 & w1948) | (~w3460 & w9272) | (w1948 & w9272);
assign w6527 = w2236 & ~w5661;
assign w6528 = ~w3017 & ~w5761;
assign w6529 = ~w5884 & ~w12531;
assign w6530 = ~w6986 & w6845;
assign w6531 = w10968 & ~w7899;
assign w6532 = (~w6750 & w11638) | (~w6750 & w7442) | (w11638 & w7442);
assign w6533 = ~w3526 & w1260;
assign w6534 = w4832 & ~w9030;
assign w6535 = (w3459 & ~w13594) | (w3459 & w3822) | (~w13594 & w3822);
assign w6536 = ~w5676 & w7655;
assign w6537 = w8389 & ~w9050;
assign w6538 = ~b116 & ~a116;
assign w6539 = w9063 & w11801;
assign w6540 = (w11730 & w13263) | (w11730 & w14180) | (w13263 & w14180);
assign w6541 = ~w2698 & ~w6427;
assign w6542 = ~b59 & ~a59;
assign w6543 = (~w2144 & w1655) | (~w2144 & w10502) | (w1655 & w10502);
assign w6544 = ~w12121 & w13300;
assign w6545 = w4349 & ~w11031;
assign w6546 = w9997 & w227;
assign w6547 = w1541 & ~w7623;
assign w6548 = (~w7630 & w4786) | (~w7630 & ~w6596) | (w4786 & ~w6596);
assign w6549 = (w890 & w4280) | (w890 & w2362) | (w4280 & w2362);
assign w6550 = ~w10395 & ~w546;
assign w6551 = ~w8254 & w7914;
assign w6552 = ~w12836 & ~w5112;
assign w6553 = w706 & w11934;
assign w6554 = w11855 & w560;
assign w6555 = w12717 & ~w12262;
assign w6556 = ~w7981 & ~w13864;
assign w6557 = (w11400 & ~w5040) | (w11400 & w2153) | (~w5040 & w2153);
assign w6558 = w7794 & ~w2745;
assign w6559 = w11880 & ~w9002;
assign w6560 = w2137 & ~w2159;
assign w6561 = w12809 & w13323;
assign w6562 = ~w12685 & w554;
assign w6563 = ~w2698 & ~w11830;
assign w6564 = ~w7794 & w9181;
assign w6565 = (w152 & w2325) | (w152 & w14643) | (w2325 & w14643);
assign w6566 = w1949 & ~w5808;
assign w6567 = (w878 & w565) | (w878 & w13504) | (w565 & w13504);
assign w6568 = (w10115 & w5154) | (w10115 & w2979) | (w5154 & w2979);
assign w6569 = ~w9788 & ~w12460;
assign w6570 = ~w3462 & ~w9045;
assign w6571 = (~w9591 & ~w13292) | (~w9591 & ~w11185) | (~w13292 & ~w11185);
assign w6572 = ~b64 & ~a64;
assign w6573 = (w3023 & w8402) | (w3023 & w4528) | (w8402 & w4528);
assign w6574 = (~w254 & w8231) | (~w254 & w2098) | (w8231 & w2098);
assign w6575 = (w3098 & ~w4266) | (w3098 & ~w217) | (~w4266 & ~w217);
assign w6576 = ~w4287 & ~w14526;
assign w6577 = ~w8937 & w9466;
assign w6578 = ~w11547 & w7796;
assign w6579 = ~w922 & ~w8937;
assign w6580 = ~b117 & ~a117;
assign w6581 = w1766 & ~w13197;
assign w6582 = w247 & ~w12271;
assign w6583 = b28 & a28;
assign w6584 = (~w142 & ~w1540) | (~w142 & w6872) | (~w1540 & w6872);
assign w6585 = ~w13459 & w8135;
assign w6586 = (~w7012 & w2698) | (~w7012 & w7526) | (w2698 & w7526);
assign w6587 = ~w10116 & ~w1986;
assign w6588 = ~w3886 & w10424;
assign w6589 = (w217 & ~w9262) | (w217 & w1239) | (~w9262 & w1239);
assign w6590 = (~w536 & ~w8234) | (~w536 & w8999) | (~w8234 & w8999);
assign w6591 = ~w13810 & w6178;
assign w6592 = w4572 & w13093;
assign w6593 = w13344 & ~w5282;
assign w6594 = (w1919 & w5927) | (w1919 & ~w10341) | (w5927 & ~w10341);
assign w6595 = ~w4603 & ~w12845;
assign w6596 = (w8827 & w5559) | (w8827 & w1754) | (w5559 & w1754);
assign w6597 = ~w8785 & w4142;
assign w6598 = (~w10272 & w10196) | (~w10272 & w10596) | (w10196 & w10596);
assign w6599 = w5257 & ~w6188;
assign w6600 = (~w10676 & w3441) | (~w10676 & w2135) | (w3441 & w2135);
assign w6601 = ~w4700 & w11934;
assign w6602 = (w13168 & w1072) | (w13168 & ~w13292) | (w1072 & ~w13292);
assign w6603 = ~w13279 & ~w5354;
assign w6604 = ~w1166 & w9805;
assign w6605 = ~w1642 & w9468;
assign w6606 = w10459 & w10631;
assign w6607 = w4407 & ~a53;
assign w6608 = w5794 | w9773;
assign w6609 = w2500 & w852;
assign w6610 = ~w11001 & ~w1148;
assign w6611 = w10928 | ~w3325;
assign w6612 = w3128 & w6119;
assign w6613 = w3914 & ~w6301;
assign w6614 = w3289 & w10286;
assign w6615 = ~w8882 & ~w5938;
assign w6616 = ~w9841 & ~w12822;
assign w6617 = ~w12271 & w4288;
assign w6618 = w2467 & ~w217;
assign w6619 = ~w3361 & w11194;
assign w6620 = ~w4700 & w5282;
assign w6621 = ~w12271 & ~w14103;
assign w6622 = ~w11298 & w4389;
assign w6623 = w6949 & ~w7684;
assign w6624 = (~w464 & ~w1940) | (~w464 & w7345) | (~w1940 & w7345);
assign w6625 = ~w238 & w9182;
assign w6626 = (w4787 & w6845) | (w4787 & w5873) | (w6845 & w5873);
assign w6627 = ~w14494 & ~w2814;
assign w6628 = w8871 & w3904;
assign w6629 = ~w12271 & w9713;
assign w6630 = ~w3019 & ~w13132;
assign w6631 = (~w9733 & w9364) | (~w9733 & ~w8282) | (w9364 & ~w8282);
assign w6632 = ~w803 & ~w12662;
assign w6633 = w11164 & ~w1008;
assign w6634 = w12344 & ~w8031;
assign w6635 = w9796 & w10713;
assign w6636 = (~w12944 & w14436) | (~w12944 & w7003) | (w14436 & w7003);
assign w6637 = (w8130 & w4783) | (w8130 & w9215) | (w4783 & w9215);
assign w6638 = ~w5559 & w9935;
assign w6639 = ~w1206 & w13885;
assign w6640 = ~w6165 & ~w4636;
assign w6641 = w4605 & ~w9309;
assign w6642 = (w12553 & w14487) | (w12553 & w9576) | (w14487 & w9576);
assign w6643 = (w13980 & w10715) | (w13980 & w13261) | (w10715 & w13261);
assign w6644 = w10880 & w4218;
assign w6645 = ~w8021 & ~w1260;
assign w6646 = ~w13300 & ~w563;
assign w6647 = w7794 & ~w1695;
assign w6648 = w12983 & w8443;
assign w6649 = w4213 & w218;
assign w6650 = (~w7085 & w12003) | (~w7085 & w3793) | (w12003 & w3793);
assign w6651 = ~w3019 & ~w1096;
assign w6652 = w5482 & w8584;
assign w6653 = w14619 & w9067;
assign w6654 = w7794 & w5884;
assign w6655 = (w1785 & w3087) | (w1785 & w12964) | (w3087 & w12964);
assign w6656 = ~w3846 & w3225;
assign w6657 = w10742 & ~w9816;
assign w6658 = ~w13940 & w5045;
assign w6659 = w4870 & w14367;
assign w6660 = (~w5783 & w1456) | (~w5783 & w12719) | (w1456 & w12719);
assign w6661 = w5177 & ~w5532;
assign w6662 = (~w7719 & w651) | (~w7719 & w11787) | (w651 & w11787);
assign w6663 = ~w2144 & w13950;
assign w6664 = ~w5786 & ~w2738;
assign w6665 = w7483 & w8975;
assign w6666 = ~w4921 & w8041;
assign w6667 = (w7636 & w5911) | (w7636 & w2824) | (w5911 & w2824);
assign w6668 = ~w1802 & ~w3251;
assign w6669 = w4288 & ~w5845;
assign w6670 = w142 & w3215;
assign w6671 = ~w12290 & ~w481;
assign w6672 = w9202 & ~w3904;
assign w6673 = (w7567 & w12275) | (w7567 & ~w8580) | (w12275 & ~w8580);
assign w6674 = (~w5282 & ~w10519) | (~w5282 & ~w3900) | (~w10519 & ~w3900);
assign w6675 = (~w9396 & ~w13654) | (~w9396 & w2518) | (~w13654 & w2518);
assign w6676 = w13239 & ~w11308;
assign w6677 = (~w1957 & w776) | (~w1957 & w1100) | (w776 & w1100);
assign w6678 = (w12589 & w9081) | (w12589 & ~w5105) | (w9081 & ~w5105);
assign w6679 = w646 & w8396;
assign w6680 = (w11675 & ~w3209) | (w11675 & w12398) | (~w3209 & w12398);
assign w6681 = ~w13587 & w11748;
assign w6682 = w6845 & ~w8319;
assign w6683 = ~w7301 & w13842;
assign w6684 = w4322 & w5282;
assign w6685 = w6301 & ~w10853;
assign w6686 = (w894 & ~w3550) | (w894 & w2118) | (~w3550 & w2118);
assign w6687 = (w12706 & w9995) | (w12706 & ~w9262) | (w9995 & ~w9262);
assign w6688 = w8352 | w11708;
assign w6689 = ~w12506 & ~w3130;
assign w6690 = ~w2500 & w4;
assign w6691 = ~w4678 & ~w7205;
assign w6692 = ~w2222 & ~w4560;
assign w6693 = ~w2719 & ~w12136;
assign w6694 = ~w2144 & w1675;
assign w6695 = ~w8229 & ~w73;
assign w6696 = ~w4098 & ~w14399;
assign w6697 = ~w4801 & w6821;
assign w6698 = w11357 & w8741;
assign w6699 = w11431 & ~w5098;
assign w6700 = w14280 & w10853;
assign w6701 = w8201 & w9063;
assign w6702 = ~w2270 & ~w10483;
assign w6703 = ~w142 & ~w2922;
assign w6704 = w7914 & w10183;
assign w6705 = ~w14088 & ~w12144;
assign w6706 = ~w6758 & w12689;
assign w6707 = ~w13387 & ~w11959;
assign w6708 = w7823 & w1040;
assign w6709 = w13732 & w9218;
assign w6710 = w2680 & w1229;
assign w6711 = ~b53 & w4303;
assign w6712 = (w5795 & w1362) | (w5795 & w9515) | (w1362 & w9515);
assign w6713 = (~w6716 & w1914) | (~w6716 & w1847) | (w1914 & w1847);
assign w6714 = (~w11031 & w6170) | (~w11031 & w9389) | (w6170 & w9389);
assign w6715 = (w2636 & w10064) | (w2636 & w8554) | (w10064 & w8554);
assign w6716 = ~b53 & ~a53;
assign w6717 = w10290 & ~w3619;
assign w6718 = ~w191 & w14233;
assign w6719 = ~w10828 & ~w10948;
assign w6720 = w11547 & ~w8973;
assign w6721 = ~w9502 & ~w3319;
assign w6722 = ~w4588 & w9144;
assign w6723 = (w876 & ~w9443) | (w876 & w10113) | (~w9443 & w10113);
assign w6724 = w499 & w10263;
assign w6725 = ~w14533 & w5892;
assign w6726 = ~w12586 & ~w12174;
assign w6727 = w12267 & w1756;
assign w6728 = ~w8827 & w3039;
assign w6729 = (~w7879 & w4099) | (~w7879 & w1894) | (w4099 & w1894);
assign w6730 = (w1114 & w14302) | (w1114 & w112) | (w14302 & w112);
assign w6731 = ~w8298 & ~w3257;
assign w6732 = (w7645 & w10320) | (w7645 & w2495) | (w10320 & w2495);
assign w6733 = (w6426 & w6808) | (w6426 & w7600) | (w6808 & w7600);
assign w6734 = (w1573 & w5418) | (w1573 & w13066) | (w5418 & w13066);
assign w6735 = w607 & ~w11031;
assign w6736 = (w9938 & w12499) | (w9938 & w135) | (w12499 & w135);
assign w6737 = ~w5082 & w248;
assign w6738 = ~w8061 & w11831;
assign w6739 = (w1199 & w2623) | (w1199 & w11105) | (w2623 & w11105);
assign w6740 = (~w9305 & w7340) | (~w9305 & w6944) | (w7340 & w6944);
assign w6741 = (w951 & w11687) | (w951 & w10163) | (w11687 & w10163);
assign w6742 = (~w9805 & ~w9013) | (~w9805 & w1019) | (~w9013 & w1019);
assign w6743 = ~w13993 & w13732;
assign w6744 = w9284 & w3904;
assign w6745 = ~w2500 & w9226;
assign w6746 = w7282 & w7071;
assign w6747 = (w4692 & w6634) | (w4692 & ~w14564) | (w6634 & ~w14564);
assign w6748 = w10422 & ~w12765;
assign w6749 = w5556 & w8389;
assign w6750 = w3550 & w9439;
assign w6751 = w12059 & w11066;
assign w6752 = (w2161 & w11247) | (w2161 & w14331) | (w11247 & w14331);
assign w6753 = ~w4050 & w13496;
assign w6754 = w5835 & ~w14417;
assign w6755 = (w11395 & w2029) | (w11395 & w13144) | (w2029 & w13144);
assign w6756 = w12460 & w9330;
assign w6757 = (w1274 & w4585) | (w1274 & w4635) | (w4585 & w4635);
assign w6758 = ~w7435 & w306;
assign w6759 = ~w4099 & w9933;
assign w6760 = w14178 & ~w7482;
assign w6761 = w1838 & ~w6689;
assign w6762 = w1190 & w1910;
assign w6763 = ~w3036 & ~w7365;
assign w6764 = ~w1840 & ~w8258;
assign w6765 = w11456 & ~w3011;
assign w6766 = ~w935 & w7497;
assign w6767 = ~w185 & ~w4710;
assign w6768 = (~w14600 & w2673) | (~w14600 & w7158) | (w2673 & w7158);
assign w6769 = ~b53 & ~w7854;
assign w6770 = (w4541 & ~w642) | (w4541 & w9137) | (~w642 & w9137);
assign w6771 = (~w7630 & w6298) | (~w7630 & w3366) | (w6298 & w3366);
assign w6772 = ~w8491 & ~w11515;
assign w6773 = w4213 & w3611;
assign w6774 = ~w11581 & w989;
assign w6775 = w11606 & ~w12429;
assign w6776 = ~w2144 & w211;
assign w6777 = w7576 & ~w12384;
assign w6778 = (w4268 & w3993) | (w4268 & w2293) | (w3993 & w2293);
assign w6779 = ~w5852 & w5227;
assign w6780 = (~w1699 & w14343) | (~w1699 & w2979) | (w14343 & w2979);
assign w6781 = (~w2698 & ~w4541) | (~w2698 & w320) | (~w4541 & w320);
assign w6782 = w2337 & ~w2143;
assign w6783 = (w803 & w14664) | (w803 & w4844) | (w14664 & w4844);
assign w6784 = (~w803 & w11482) | (~w803 & w10676) | (w11482 & w10676);
assign w6785 = w13590 & w9138;
assign w6786 = ~w13080 & ~w8947;
assign w6787 = ~w10339 & ~w6492;
assign w6788 = ~w3914 & w14390;
assign w6789 = w12596 | w6819;
assign w6790 = ~w857 & w6724;
assign w6791 = w3128 & w2563;
assign w6792 = ~w13349 & w1030;
assign w6793 = ~w12493 & w7121;
assign w6794 = w6558 & w11461;
assign w6795 = (~w12065 & w1171) | (~w12065 & w1536) | (w1171 & w1536);
assign w6796 = w6405 & ~w5622;
assign w6797 = (~w8659 & w977) | (~w8659 & w8238) | (w977 & w8238);
assign w6798 = (~w5483 & w11384) | (~w5483 & w5878) | (w11384 & w5878);
assign w6799 = (w302 & w10458) | (w302 & w7262) | (w10458 & w7262);
assign w6800 = ~w1062 & ~w10864;
assign w6801 = ~w8052 & ~w3105;
assign w6802 = (w9305 & w4754) | (w9305 & w13980) | (w4754 & w13980);
assign w6803 = w12330 & ~w12112;
assign w6804 = w7794 & ~w11476;
assign w6805 = (~w10044 & w8595) | (~w10044 & w1952) | (w8595 & w1952);
assign w6806 = ~w7662 & ~w12311;
assign w6807 = w10676 & w7772;
assign w6808 = (~w12775 & w10188) | (~w12775 & w4232) | (w10188 & w4232);
assign w6809 = ~w12464 & w13733;
assign w6810 = ~w11745 & ~w7670;
assign w6811 = ~w12606 & w4812;
assign w6812 = ~w3555 & ~w12147;
assign w6813 = ~w11810 & ~w9938;
assign w6814 = (w13462 & w8143) | (w13462 & w10258) | (w8143 & w10258);
assign w6815 = w13099 & w12425;
assign w6816 = ~w11487 & ~w12471;
assign w6817 = ~w3526 & w2236;
assign w6818 = w1263 & w4441;
assign w6819 = ~w14504 & w5922;
assign w6820 = ~w2036 & ~w3904;
assign w6821 = (~w12980 & w6322) | (~w12980 & w60) | (w6322 & w60);
assign w6822 = (~w3611 & w4218) | (~w3611 & ~w3556) | (w4218 & ~w3556);
assign w6823 = w1087 & ~w3904;
assign w6824 = ~w2433 & ~w5761;
assign w6825 = ~w14054 & ~w11345;
assign w6826 = (w3401 & ~w8572) | (w3401 & w2196) | (~w8572 & w2196);
assign w6827 = (w4204 & w1501) | (w4204 & ~w1928) | (w1501 & ~w1928);
assign w6828 = (w6500 & w5562) | (w6500 & w8003) | (w5562 & w8003);
assign w6829 = ~w6750 & w3125;
assign w6830 = (w12305 & w5088) | (w12305 & w13165) | (w5088 & w13165);
assign w6831 = ~w2387 & w11500;
assign w6832 = (w9912 & w1982) | (w9912 & w1688) | (w1982 & w1688);
assign w6833 = ~w4158 & w8042;
assign w6834 = w12091 & w6409;
assign w6835 = ~w5240 & ~w14589;
assign w6836 = (~w5036 & w10143) | (~w5036 & w8806) | (w10143 & w8806);
assign w6837 = (~w10182 & w12167) | (~w10182 & w7694) | (w12167 & w7694);
assign w6838 = ~w8937 & w1912;
assign w6839 = w2656 & w852;
assign w6840 = w894 & ~w7630;
assign w6841 = (~w77 & w2406) | (~w77 & ~w2656) | (w2406 & ~w2656);
assign w6842 = ~w12609 & w2162;
assign w6843 = w12267 & w2000;
assign w6844 = ~w6824 & w3210;
assign w6845 = (~w8234 & w12652) | (~w8234 & w4937) | (w12652 & w4937);
assign w6846 = ~w1563 & ~w4676;
assign w6847 = ~w5498 & ~w13375;
assign w6848 = (w5331 & w4436) | (w5331 & w8228) | (w4436 & w8228);
assign w6849 = (~w10688 & ~w6656) | (~w10688 & w5662) | (~w6656 & w5662);
assign w6850 = ~w1523 & w9130;
assign w6851 = (w12569 & w8803) | (w12569 & ~w13621) | (w8803 & ~w13621);
assign w6852 = ~w6663 & ~w969;
assign w6853 = w1764 & w14016;
assign w6854 = w12918 & w2985;
assign w6855 = w11680 & ~w13998;
assign w6856 = ~w8937 & w10735;
assign w6857 = w10328 & w2672;
assign w6858 = ~w8171 & ~w2922;
assign w6859 = (w10997 & w2175) | (w10997 & w6004) | (w2175 & w6004);
assign w6860 = (~w3602 & w8071) | (~w3602 & ~w12992) | (w8071 & ~w12992);
assign w6861 = ~w829 & ~w2270;
assign w6862 = (~w4030 & w6389) | (~w4030 & w4956) | (w6389 & w4956);
assign w6863 = (w6103 & w13449) | (w6103 & w9034) | (w13449 & w9034);
assign w6864 = (w7343 & w7635) | (w7343 & w3791) | (w7635 & w3791);
assign w6865 = (w8637 & w2415) | (w8637 & ~w12638) | (w2415 & ~w12638);
assign w6866 = (~w3317 & w6491) | (~w3317 & ~w8331) | (w6491 & ~w8331);
assign w6867 = w724 & w608;
assign w6868 = ~b53 & ~w6588;
assign w6869 = w9871 & w9817;
assign w6870 = w12121 & w6542;
assign w6871 = ~w5263 & w11047;
assign w6872 = ~w14276 & ~w142;
assign w6873 = (w8873 & ~w14506) | (w8873 & w900) | (~w14506 & w900);
assign w6874 = w12371 & ~w12642;
assign w6875 = ~w1152 & ~w3904;
assign w6876 = w6820 & ~w8488;
assign w6877 = ~w3734 & w6886;
assign w6878 = ~w14302 & w2680;
assign w6879 = (w10711 & w4582) | (w10711 & w21) | (w4582 & w21);
assign w6880 = ~w12003 & w3222;
assign w6881 = w14403 & ~w1983;
assign w6882 = (~w12642 & ~w8740) | (~w12642 & w8925) | (~w8740 & w8925);
assign w6883 = w5317 & w2928;
assign w6884 = ~w5074 & ~w14114;
assign w6885 = w9861 & w9646;
assign w6886 = (~w2933 & w10872) | (~w2933 & w4135) | (w10872 & w4135);
assign w6887 = w1607 & ~w14227;
assign w6888 = (~w10675 & w3971) | (~w10675 & w4706) | (w3971 & w4706);
assign w6889 = ~b73 & ~a73;
assign w6890 = (~w5702 & w7603) | (~w5702 & w2378) | (w7603 & w2378);
assign w6891 = ~w5294 & ~w2135;
assign w6892 = (w7556 & w7465) | (w7556 & w3514) | (w7465 & w3514);
assign w6893 = ~w1540 & w2485;
assign w6894 = w11971 & ~w14483;
assign w6895 = w10568 & ~w11764;
assign w6896 = w265 & w2605;
assign w6897 = ~w5482 & ~w40;
assign w6898 = w13197 & w2481;
assign w6899 = w7875 & ~w11940;
assign w6900 = w2316 & ~w6074;
assign w6901 = (~w14463 & w9404) | (~w14463 & w8789) | (w9404 & w8789);
assign w6902 = (w1746 & w11268) | (w1746 & w4174) | (w11268 & w4174);
assign w6903 = ~w12723 & ~w13345;
assign w6904 = ~w2463 & w1136;
assign w6905 = ~w12003 & w8053;
assign w6906 = w309 & w5664;
assign w6907 = w8131 & w9041;
assign w6908 = ~w676 & ~w12749;
assign w6909 = (~w12406 & w8329) | (~w12406 & w2805) | (w8329 & w2805);
assign w6910 = ~w6433 & ~w125;
assign w6911 = w5505 & w14506;
assign w6912 = w9119 & ~w7101;
assign w6913 = ~w1474 & w11117;
assign w6914 = w803 & w5247;
assign w6915 = w2602 & ~w2041;
assign w6916 = w4213 & ~w6816;
assign w6917 = ~w13768 & ~w11539;
assign w6918 = (~w3550 & w13166) | (~w3550 & w156) | (w13166 & w156);
assign w6919 = (w1190 & w7015) | (w1190 & w9989) | (w7015 & w9989);
assign w6920 = w7395 & ~w8178;
assign w6921 = w10689 & w803;
assign w6922 = ~w10675 & w10122;
assign w6923 = w12464 & ~w183;
assign w6924 = (w9378 & ~w2372) | (w9378 & w2504) | (~w2372 & w2504);
assign w6925 = (~w12776 & w8673) | (~w12776 & w10701) | (w8673 & w10701);
assign w6926 = ~w12506 & ~w8782;
assign w6927 = w10075 & w9032;
assign w6928 = w211 & w11487;
assign w6929 = w12575 & w3957;
assign w6930 = w11371 & w2173;
assign w6931 = w12385 & ~w8610;
assign w6932 = w499 & ~w5693;
assign w6933 = w2332 & ~w2492;
assign w6934 = w8791 & w10916;
assign w6935 = (~w5693 & w5451) | (~w5693 & w3212) | (w5451 & w3212);
assign w6936 = w10371 & w5431;
assign w6937 = (w5952 & w340) | (w5952 & w6496) | (w340 & w6496);
assign w6938 = ~w9280 & ~w13649;
assign w6939 = ~w5268 & ~w2640;
assign w6940 = w14408 & w3787;
assign w6941 = w2941 & w4845;
assign w6942 = w7794 & w9957;
assign w6943 = w5911 | w7636;
assign w6944 = (w7515 & w6991) | (w7515 & w6549) | (w6991 & w6549);
assign w6945 = (w8513 & w11360) | (w8513 & w10537) | (w11360 & w10537);
assign w6946 = w2320 & w7630;
assign w6947 = (w10968 & w6181) | (w10968 & w5175) | (w6181 & w5175);
assign w6948 = ~w11261 & w13115;
assign w6949 = (~w8512 & w4467) | (~w8512 & w8017) | (w4467 & w8017);
assign w6950 = w3383 & ~w10033;
assign w6951 = w2202 & ~w2864;
assign w6952 = ~w6281 & ~w13713;
assign w6953 = w4300 & w7615;
assign w6954 = (~w9305 & w3260) | (~w9305 & w3381) | (w3260 & w3381);
assign w6955 = (w5961 & w1594) | (w5961 & w12376) | (w1594 & w12376);
assign w6956 = ~w13665 & ~w463;
assign w6957 = w10509 & w7115;
assign w6958 = w10704 & ~w12170;
assign w6959 = w12483 & w5105;
assign w6960 = ~w5263 & ~w7149;
assign w6961 = ~w5294 & ~w1442;
assign w6962 = (~w8513 & ~w12271) | (~w8513 & w10626) | (~w12271 & w10626);
assign w6963 = w10880 & w9159;
assign w6964 = w14390 & w8900;
assign w6965 = w5282 & ~w2228;
assign w6966 = ~w1530 & w7406;
assign w6967 = ~w12240 & ~w3435;
assign w6968 = ~w3006 & ~w12511;
assign w6969 = w3914 & ~w10813;
assign w6970 = ~w3751 & w12087;
assign w6971 = (w11934 & ~w10562) | (w11934 & w12540) | (~w10562 & w12540);
assign w6972 = w13323 & w5761;
assign w6973 = (w10470 & ~w12755) | (w10470 & w9354) | (~w12755 & w9354);
assign w6974 = (~w5243 & w3146) | (~w5243 & ~w12125) | (w3146 & ~w12125);
assign w6975 = b38 & a38;
assign w6976 = (~w11211 & ~w13885) | (~w11211 & w5785) | (~w13885 & w5785);
assign w6977 = w183 & w6716;
assign w6978 = w2982 & w12025;
assign w6979 = ~w928 & w393;
assign w6980 = ~w11583 & w1968;
assign w6981 = w7169 | ~w7338;
assign w6982 = (w13020 & w8762) | (w13020 & w12376) | (w8762 & w12376);
assign w6983 = ~w12589 & w8769;
assign w6984 = (w8288 & w8670) | (w8288 & w832) | (w8670 & w832);
assign w6985 = w2653 & a53;
assign w6986 = (~w2159 & w11431) | (~w2159 & w12528) | (w11431 & w12528);
assign w6987 = (~w1260 & w3385) | (~w1260 & w14669) | (w3385 & w14669);
assign w6988 = ~w13627 & ~w8597;
assign w6989 = ~w7242 & w1985;
assign w6990 = (~w756 & w12781) | (~w756 & ~w4694) | (w12781 & ~w4694);
assign w6991 = w4280 | w890;
assign w6992 = ~w845 & w10073;
assign w6993 = w8613 & ~w7346;
assign w6994 = w21 & ~w13375;
assign w6995 = ~w7348 & w11604;
assign w6996 = (w1190 & w3952) | (w1190 & w9989) | (w3952 & w9989);
assign w6997 = (w18 & w9092) | (w18 & ~w13920) | (w9092 & ~w13920);
assign w6998 = (w11273 & w13372) | (w11273 & w12376) | (w13372 & w12376);
assign w6999 = (~w13222 & w742) | (~w13222 & w5434) | (w742 & w5434);
assign w7000 = ~w14015 & ~w12604;
assign w7001 = ~b119 & ~a119;
assign w7002 = w5707 & ~w9996;
assign w7003 = w6425 & w324;
assign w7004 = w6176 & ~w12839;
assign w7005 = ~w705 & ~w7333;
assign w7006 = (~w9608 & w5045) | (~w9608 & w8581) | (w5045 & w8581);
assign w7007 = (~w142 & w3727) | (~w142 & w6872) | (w3727 & w6872);
assign w7008 = (w3538 & w11579) | (w3538 & w1724) | (w11579 & w1724);
assign w7009 = ~w107 & ~w884;
assign w7010 = w6935 & ~w1862;
assign w7011 = ~w2470 & w11286;
assign w7012 = ~w7420 & ~w8170;
assign w7013 = b29 & a29;
assign w7014 = ~w142 & w12065;
assign w7015 = w6603 & w4778;
assign w7016 = ~w13426 & ~w8809;
assign w7017 = w2850 & ~w10393;
assign w7018 = (w1663 & w9617) | (w1663 & w251) | (w9617 & w251);
assign w7019 = w2909 & ~w1150;
assign w7020 = (~w473 & ~w5016) | (~w473 & ~w12003) | (~w5016 & ~w12003);
assign w7021 = ~w491 & ~w5407;
assign w7022 = ~b19 & ~a19;
assign w7023 = ~w5401 & ~w8640;
assign w7024 = (~w14395 & w7488) | (~w14395 & w89) | (w7488 & w89);
assign w7025 = w10037 & ~w13748;
assign w7026 = ~w5448 & ~w5581;
assign w7027 = w13396 & ~w12625;
assign w7028 = (~w6276 & w8300) | (~w6276 & w9416) | (w8300 & w9416);
assign w7029 = (w12801 & w11331) | (w12801 & w8948) | (w11331 & w8948);
assign w7030 = ~w192 & ~w12644;
assign w7031 = (~w10483 & w9) | (~w10483 & w13716) | (w9 & w13716);
assign w7032 = w5669 & w8961;
assign w7033 = w6346 & w1414;
assign w7034 = (w10116 & w6845) | (w10116 & w14655) | (w6845 & w14655);
assign w7035 = w808 & ~w471;
assign w7036 = ~w6556 & ~w217;
assign w7037 = w607 & ~w6689;
assign w7038 = ~w7670 & ~w6627;
assign w7039 = w5835 & ~w4511;
assign w7040 = ~w13628 & w10274;
assign w7041 = w9607 & w14313;
assign w7042 = ~w9906 & ~w9659;
assign w7043 = ~w11013 & ~w13323;
assign w7044 = ~w14535 & ~w12105;
assign w7045 = w10993 & w13026;
assign w7046 = w8584 & ~w10006;
assign w7047 = (~w10853 & w4050) | (~w10853 & w3830) | (w4050 & w3830);
assign w7048 = ~w11924 & ~w9396;
assign w7049 = w8572 & w10748;
assign w7050 = ~w3667 & w13883;
assign w7051 = ~w8960 & ~w7232;
assign w7052 = ~w6712 & w5074;
assign w7053 = ~w3348 & w13143;
assign w7054 = ~w4416 & ~w365;
assign w7055 = (~b93 & ~w1840) | (~b93 & w5847) | (~w1840 & w5847);
assign w7056 = w2800 & ~w6199;
assign w7057 = ~w1789 & w8680;
assign w7058 = ~w3288 & ~w8719;
assign w7059 = ~w12271 & w10621;
assign w7060 = ~w3914 & w11835;
assign w7061 = (~w14216 & w12277) | (~w14216 & w4742) | (w12277 & w4742);
assign w7062 = (w11516 & w11037) | (w11516 & w9724) | (w11037 & w9724);
assign w7063 = w10277 & ~w3515;
assign w7064 = (~w4464 & w7179) | (~w4464 & w2988) | (w7179 & w2988);
assign w7065 = w7772 & w1260;
assign w7066 = ~w8778 & ~w7312;
assign w7067 = ~w3759 & w4341;
assign w7068 = (~w894 & w9608) | (~w894 & w7853) | (w9608 & w7853);
assign w7069 = w11880 & w4088;
assign w7070 = (~w6215 & w8490) | (~w6215 & w13235) | (w8490 & w13235);
assign w7071 = w12936 & w6917;
assign w7072 = ~w7908 & w8161;
assign w7073 = (~w9733 & w9364) | (~w9733 & ~w2595) | (w9364 & ~w2595);
assign w7074 = ~w11500 & w5005;
assign w7075 = ~w14015 & ~w14569;
assign w7076 = (~w8080 & w13122) | (~w8080 & w9299) | (w13122 & w9299);
assign w7077 = w8740 & ~w3846;
assign w7078 = (w13752 & w13910) | (w13752 & w13035) | (w13910 & w13035);
assign w7079 = ~w1437 & ~w4014;
assign w7080 = ~w2159 & ~w13838;
assign w7081 = w5294 & w894;
assign w7082 = (~w4780 & w3700) | (~w4780 & w10962) | (w3700 & w10962);
assign w7083 = ~w14276 & ~w3098;
assign w7084 = w8663 & w7575;
assign w7085 = w14215 & w1842;
assign w7086 = (~w14504 & w12003) | (~w14504 & w12598) | (w12003 & w12598);
assign w7087 = ~w6301 & w6427;
assign w7088 = ~w5294 & w6281;
assign w7089 = (w347 & w13928) | (w347 & w5330) | (w13928 & w5330);
assign w7090 = ~w10309 & w4741;
assign w7091 = w894 & ~w6230;
assign w7092 = w2544 & ~w14659;
assign w7093 = (w11500 & w1692) | (w11500 & w6831) | (w1692 & w6831);
assign w7094 = w11702 & ~w1540;
assign w7095 = ~w1102 & ~w12946;
assign w7096 = ~w13954 & w3427;
assign w7097 = w1805 & ~w7684;
assign w7098 = ~w9720 & w10135;
assign w7099 = (w13192 & ~w13320) | (w13192 & w8155) | (~w13320 & w8155);
assign w7100 = (~w13946 & ~w6929) | (~w13946 & w2952) | (~w6929 & w2952);
assign w7101 = w3138 & w3123;
assign w7102 = ~w3484 & w2953;
assign w7103 = (~w13219 & w1911) | (~w13219 & w4069) | (w1911 & w4069);
assign w7104 = ~w6538 & ~w4848;
assign w7105 = ~w3659 & ~w2161;
assign w7106 = ~w5604 & ~w8919;
assign w7107 = (~w6637 & w13266) | (~w6637 & w13536) | (w13266 & w13536);
assign w7108 = w10653 & ~w11795;
assign w7109 = (~w13219 & w6622) | (~w13219 & w83) | (w6622 & w83);
assign w7110 = w330 & w4838;
assign w7111 = ~w364 & ~w3803;
assign w7112 = w14344 & w13355;
assign w7113 = ~w13321 & w9342;
assign w7114 = (~w8851 & ~w161) | (~w8851 & w13795) | (~w161 & w13795);
assign w7115 = (~w8899 & w5070) | (~w8899 & w2287) | (w5070 & w2287);
assign w7116 = ~w3015 & w7951;
assign w7117 = ~w10568 & w12642;
assign w7118 = (w10719 & w11688) | (w10719 & w10635) | (w11688 & w10635);
assign w7119 = (w11732 & w3924) | (w11732 & w8234) | (w3924 & w8234);
assign w7120 = ~w9482 & w2941;
assign w7121 = w14417 & w12662;
assign w7122 = ~w10225 & ~w3661;
assign w7123 = ~w2762 & w13872;
assign w7124 = w4173 & w4925;
assign w7125 = ~w7244 & ~w3727;
assign w7126 = w14498 & w7267;
assign w7127 = (w6802 & w2502) | (w6802 & w11015) | (w2502 & w11015);
assign w7128 = ~w10309 & w13227;
assign w7129 = (~w8614 & w696) | (~w8614 & w997) | (w696 & w997);
assign w7130 = (~w10290 & ~w8389) | (~w10290 & w5580) | (~w8389 & w5580);
assign w7131 = w6093 & w8926;
assign w7132 = ~w364 & ~w2751;
assign w7133 = w13564 & ~w12181;
assign w7134 = ~w9004 & ~w3044;
assign w7135 = w499 & w9366;
assign w7136 = w9378 & w8513;
assign w7137 = w14019 & ~w8410;
assign w7138 = ~w4553 & w9207;
assign w7139 = w3568 & ~w11747;
assign w7140 = (w659 & w3505) | (w659 & w4426) | (w3505 & w4426);
assign w7141 = ~w9012 & w1575;
assign w7142 = (w1949 & w7645) | (w1949 & w12854) | (w7645 & w12854);
assign w7143 = ~w14369 & w5663;
assign w7144 = ~w6855 & w2458;
assign w7145 = ~w14302 & w3036;
assign w7146 = (w14463 & w4816) | (w14463 & w414) | (w4816 & w414);
assign w7147 = (w4784 & w11133) | (w4784 & w9403) | (w11133 & w9403);
assign w7148 = w5030 & w4150;
assign w7149 = w7165 & w2390;
assign w7150 = ~w8097 & w6885;
assign w7151 = w3128 & w7192;
assign w7152 = w9554 & w257;
assign w7153 = (w152 & w2325) | (w152 & w7639) | (w2325 & w7639);
assign w7154 = ~w14015 & w14569;
assign w7155 = (w7796 & w82) | (w7796 & w13409) | (w82 & w13409);
assign w7156 = (w3973 & w13067) | (w3973 & ~w8228) | (w13067 & ~w8228);
assign w7157 = ~w12463 & ~w7022;
assign w7158 = w10165 & w9709;
assign w7159 = w7794 & ~w13296;
assign w7160 = (~w13628 & w5294) | (~w13628 & w12796) | (w5294 & w12796);
assign w7161 = ~w5203 & ~w9706;
assign w7162 = (w6502 & ~w3044) | (w6502 & w13416) | (~w3044 & w13416);
assign w7163 = ~w2500 & w1805;
assign w7164 = w1802 & w7670;
assign w7165 = w7255 & w12462;
assign w7166 = (w13502 & w9598) | (w13502 & w11141) | (w9598 & w11141);
assign w7167 = w11232 & w2700;
assign w7168 = ~w4623 & ~w13147;
assign w7169 = w2858 & ~w7338;
assign w7170 = ~w4846 & ~w12168;
assign w7171 = w7305 & ~w1802;
assign w7172 = w13452 & ~w10956;
assign w7173 = ~w9480 & w2701;
assign w7174 = w7317 & w4728;
assign w7175 = (~w14526 & w183) | (~w14526 & w4287) | (w183 & w4287);
assign w7176 = (w12065 & ~w3963) | (w12065 & w7014) | (~w3963 & w7014);
assign w7177 = ~w8780 & w172;
assign w7178 = w5556 & w3671;
assign w7179 = ~w1827 & ~w13187;
assign w7180 = (w13406 & w14621) | (w13406 & w11490) | (w14621 & w11490);
assign w7181 = w7013 & w12642;
assign w7182 = (w13047 & w6092) | (w13047 & w7983) | (w6092 & w7983);
assign w7183 = w3552 & w4364;
assign w7184 = ~w7782 & w11026;
assign w7185 = w706 & w10699;
assign w7186 = (w3039 & w8900) | (w3039 & w7324) | (w8900 & w7324);
assign w7187 = (~w7806 & w3348) | (~w7806 & w10175) | (w3348 & w10175);
assign w7188 = ~w2701 & ~w901;
assign w7189 = (w6176 & w4741) | (w6176 & w6449) | (w4741 & w6449);
assign w7190 = b74 & a74;
assign w7191 = ~w12664 & ~w12825;
assign w7192 = ~w6750 & ~w13853;
assign w7193 = ~w10992 & ~w6385;
assign w7194 = ~w4939 & w9075;
assign w7195 = ~w5097 & ~w10478;
assign w7196 = w12371 & ~w8396;
assign w7197 = ~w13153 & ~w9675;
assign w7198 = (~w68 & w1648) | (~w68 & w12044) | (w1648 & w12044);
assign w7199 = ~w7001 & ~w7670;
assign w7200 = w10116 & w9938;
assign w7201 = (w6276 & w6088) | (w6276 & w8458) | (w6088 & w8458);
assign w7202 = ~w14005 & w7286;
assign w7203 = (w11327 & w13213) | (w11327 & w217) | (w13213 & w217);
assign w7204 = w12603 & ~w4756;
assign w7205 = ~w2864 & ~w9296;
assign w7206 = ~w6588 & w9712;
assign w7207 = ~w13324 & w2471;
assign w7208 = ~w2656 & w1130;
assign w7209 = w2374 & ~w6077;
assign w7210 = ~w10099 & w6725;
assign w7211 = ~w9043 & w10858;
assign w7212 = w10590 & ~w8080;
assign w7213 = w11442 & ~w8034;
assign w7214 = ~w607 & ~w9211;
assign w7215 = (w6117 & w9279) | (w6117 & w5534) | (w9279 & w5534);
assign w7216 = w12457 & w57;
assign w7217 = (~w10590 & w7423) | (~w10590 & w2470) | (w7423 & w2470);
assign w7218 = ~w6286 & ~w7788;
assign w7219 = ~w13697 & w1908;
assign w7220 = (w4756 & w11205) | (w4756 & w2600) | (w11205 & w2600);
assign w7221 = ~w1062 & w10441;
assign w7222 = ~w5702 & w2058;
assign w7223 = w5731 & ~w2066;
assign w7224 = w3325 & w6228;
assign w7225 = (w4795 & w436) | (w4795 & ~w3095) | (w436 & ~w3095);
assign w7226 = ~w12438 & ~w5451;
assign w7227 = (~w2933 & w1642) | (~w2933 & w5455) | (w1642 & w5455);
assign w7228 = w11997 & w8389;
assign w7229 = ~w11117 & ~w6614;
assign w7230 = w10290 & ~w5225;
assign w7231 = ~w6442 & w1756;
assign w7232 = ~w13324 & w14480;
assign w7233 = ~w4477 & ~w4649;
assign w7234 = w610 & w5102;
assign w7235 = (~w10926 & w8742) | (~w10926 & w4259) | (w8742 & w4259);
assign w7236 = ~w14072 & ~w3508;
assign w7237 = w7493 & w4068;
assign w7238 = ~w4032 & w9871;
assign w7239 = (w4627 & w91) | (w4627 & w12616) | (w91 & w12616);
assign w7240 = (~w3611 & ~w7709) | (~w3611 & w4218) | (~w7709 & w4218);
assign w7241 = w128 & w10338;
assign w7242 = (w14185 & w2972) | (w14185 & w4748) | (w2972 & w4748);
assign w7243 = ~w8484 & w2046;
assign w7244 = b119 & a119;
assign w7245 = w1491 & ~w3194;
assign w7246 = ~w12653 & ~w11504;
assign w7247 = ~w3636 & ~w11117;
assign w7248 = ~w14186 & w2478;
assign w7249 = w4312 & ~w13713;
assign w7250 = ~w3759 & ~w11723;
assign w7251 = w8737 & ~w3383;
assign w7252 = w10409 & w8115;
assign w7253 = ~w7305 & ~w3963;
assign w7254 = w11097 & ~w3466;
assign w7255 = ~w12870 & ~w11526;
assign w7256 = (~w12662 & w2135) | (~w12662 & w12191) | (w2135 & w12191);
assign w7257 = ~w12003 & w7679;
assign w7258 = ~w14141 & w10018;
assign w7259 = (~w3704 & w4295) | (~w3704 & w767) | (w4295 & w767);
assign w7260 = w8105 & w2722;
assign w7261 = ~b5 & ~a5;
assign w7262 = (w4454 & w14587) | (w4454 & w14182) | (w14587 & w14182);
assign w7263 = ~w12001 & w10321;
assign w7264 = ~w4213 & w12398;
assign w7265 = ~w4453 & ~w12884;
assign w7266 = (~w1955 & w8608) | (~w1955 & ~w9248) | (w8608 & ~w9248);
assign w7267 = ~w12167 & w1845;
assign w7268 = w12433 & ~w13786;
assign w7269 = ~w2317 & w4403;
assign w7270 = ~w4376 & ~w9085;
assign w7271 = ~w9708 & ~w12148;
assign w7272 = ~w1517 & w4016;
assign w7273 = w4078 & w4134;
assign w7274 = (~w6276 & w1547) | (~w6276 & w11314) | (w1547 & w11314);
assign w7275 = (w12406 & w6149) | (w12406 & w370) | (w6149 & w370);
assign w7276 = ~w9480 & ~w10013;
assign w7277 = w14271 & ~w10119;
assign w7278 = w9809 & w9211;
assign w7279 = w9388 & ~w8776;
assign w7280 = w3025 & ~w3671;
assign w7281 = (w2548 & w817) | (w2548 & w1078) | (w817 & w1078);
assign w7282 = ~w11449 & w2819;
assign w7283 = ~w1557 & ~w0;
assign w7284 = ~w10245 & w4644;
assign w7285 = w1041 & w9490;
assign w7286 = w4599 & w10342;
assign w7287 = ~w5620 & w11810;
assign w7288 = ~w6700 & ~w8421;
assign w7289 = ~w12148 & w11933;
assign w7290 = (w5863 & w9965) | (w5863 & w10806) | (w9965 & w10806);
assign w7291 = (w1479 & w11638) | (w1479 & w812) | (w11638 & w812);
assign w7292 = w11429 & w10560;
assign w7293 = (w3039 & w6230) | (w3039 & w7324) | (w6230 & w7324);
assign w7294 = w4598 & ~w6698;
assign w7295 = ~w11606 & ~w2864;
assign w7296 = (~w11488 & w11604) | (~w11488 & w8852) | (w11604 & w8852);
assign w7297 = ~w3885 & w1062;
assign w7298 = w10091 & ~w1159;
assign w7299 = (w1559 & w13303) | (w1559 & w6705) | (w13303 & w6705);
assign w7300 = w13935 & w14077;
assign w7301 = ~w12545 & w10388;
assign w7302 = (w3388 & w14586) | (w3388 & ~w9403) | (w14586 & ~w9403);
assign w7303 = ~w10334 & ~w8338;
assign w7304 = (~w4783 & ~w8130) | (~w4783 & w4770) | (~w8130 & w4770);
assign w7305 = ~b105 & ~a105;
assign w7306 = ~w11462 & ~w6975;
assign w7307 = ~w6776 & ~w338;
assign w7308 = w723 & ~w10713;
assign w7309 = ~w13963 & ~w9812;
assign w7310 = w8819 & ~w8396;
assign w7311 = w10824 & ~w1404;
assign w7312 = ~w2674 & w2650;
assign w7313 = ~w1166 & w14659;
assign w7314 = ~w770 & w10400;
assign w7315 = ~w8440 & w13230;
assign w7316 = (w8085 & w3914) | (w8085 & w5717) | (w3914 & w5717);
assign w7317 = w4287 & w3734;
assign w7318 = (w4044 & w10988) | (w4044 & w3539) | (w10988 & w3539);
assign w7319 = w8768 & w10781;
assign w7320 = w9912 & ~w10894;
assign w7321 = ~w1802 & w14356;
assign w7322 = w5282 & w7001;
assign w7323 = (~w4545 & w6673) | (~w4545 & w2238) | (w6673 & w2238);
assign w7324 = ~w12065 & w3039;
assign w7325 = (w9927 & ~w1800) | (w9927 & w14524) | (~w1800 & w14524);
assign w7326 = (~w9223 & w5603) | (~w9223 & w4208) | (w5603 & w4208);
assign w7327 = (w8584 & w10467) | (w8584 & w8734) | (w10467 & w8734);
assign w7328 = w1387 & w7704;
assign w7329 = w5490 & ~w3369;
assign w7330 = (w1315 & ~w5253) | (w1315 & w10558) | (~w5253 & w10558);
assign w7331 = w12868 & w12483;
assign w7332 = ~w2267 & w4324;
assign w7333 = ~w11663 & w5987;
assign w7334 = w2578 & w8937;
assign w7335 = b104 & a104;
assign w7336 = ~w10334 & ~w5271;
assign w7337 = ~w180 & ~w3280;
assign w7338 = ~w3502 & ~w10605;
assign w7339 = ~w4050 & w9998;
assign w7340 = (w890 & w4280) | (w890 & ~w13980) | (w4280 & ~w13980);
assign w7341 = ~w509 & w1503;
assign w7342 = w7085 & w724;
assign w7343 = w12257 & ~w434;
assign w7344 = w6603 & ~w8313;
assign w7345 = ~w4752 & ~w464;
assign w7346 = ~w9954 & w14241;
assign w7347 = w6226 & ~w1514;
assign w7348 = (~w6542 & w1235) | (~w6542 & w1779) | (w1235 & w1779);
assign w7349 = w2941 & w6500;
assign w7350 = w1504 & ~w8704;
assign w7351 = ~w1423 & ~w3289;
assign w7352 = ~w12271 & w12662;
assign w7353 = w8769 & ~w10173;
assign w7354 = (~w9219 & ~w14396) | (~w9219 & w2336) | (~w14396 & w2336);
assign w7355 = w9854 & w227;
assign w7356 = ~w2676 & w4085;
assign w7357 = w12575 & ~w852;
assign w7358 = w5220 & w12460;
assign w7359 = (~w11385 & w13460) | (~w11385 & w13023) | (w13460 & w13023);
assign w7360 = (w9503 & ~w6938) | (w9503 & w13043) | (~w6938 & w13043);
assign w7361 = ~w781 & w4651;
assign w7362 = w8370 & ~w10339;
assign w7363 = (w13937 & w3989) | (w13937 & w11712) | (w3989 & w11712);
assign w7364 = w11843 & w7428;
assign w7365 = ~b92 & ~a92;
assign w7366 = ~w12240 & w9226;
assign w7367 = ~w7190 & w9087;
assign w7368 = (w10317 & w2463) | (w10317 & w9282) | (w2463 & w9282);
assign w7369 = b108 & a108;
assign w7370 = w7001 & w6689;
assign w7371 = ~w5638 & w4358;
assign w7372 = ~w1177 & w7512;
assign w7373 = ~b6 & ~a6;
assign w7374 = ~w10699 & w7486;
assign w7375 = w5563 | w1986;
assign w7376 = ~w607 & ~w5522;
assign w7377 = w1173 & ~w10525;
assign w7378 = (w11429 & w1146) | (w11429 & w362) | (w1146 & w362);
assign w7379 = w8390 & w4127;
assign w7380 = w536 & w13531;
assign w7381 = ~w10309 & ~w13227;
assign w7382 = (w2320 & ~w3963) | (w2320 & w10103) | (~w3963 & w10103);
assign w7383 = ~w10245 & w12767;
assign w7384 = ~w3159 & ~w9211;
assign w7385 = ~w2386 & ~w2926;
assign w7386 = ~b53 & w1816;
assign w7387 = ~w8226 & w4988;
assign w7388 = w13095 & w12914;
assign w7389 = (w1935 & w5270) | (w1935 & w11823) | (w5270 & w11823);
assign w7390 = (~w13654 & w4356) | (~w13654 & w13179) | (w4356 & w13179);
assign w7391 = w607 & w8459;
assign w7392 = ~w12212 & w6892;
assign w7393 = w3017 & ~w4458;
assign w7394 = w9176 & w6159;
assign w7395 = w14492 & w10842;
assign w7396 = (~w3615 & w11278) | (~w3615 & ~w3564) | (w11278 & ~w3564);
assign w7397 = ~w9454 & ~w9052;
assign w7398 = w2806 & w10689;
assign w7399 = ~w7913 & ~w6482;
assign w7400 = ~w6583 & ~w7013;
assign w7401 = w3435 & ~w1389;
assign w7402 = (w3025 & ~w3128) | (w3025 & w4013) | (~w3128 & w4013);
assign w7403 = w9949 & w12642;
assign w7404 = w5166 & ~w11039;
assign w7405 = w7312 & ~w5785;
assign w7406 = w6064 & w10182;
assign w7407 = (w922 & w1962) | (w922 & w11822) | (w1962 & w11822);
assign w7408 = ~w14302 & w2332;
assign w7409 = ~w3914 & w3317;
assign w7410 = w690 & ~w2272;
assign w7411 = w3215 & ~w3611;
assign w7412 = w11497 & w8160;
assign w7413 = (w7273 & w6416) | (w7273 & w7664) | (w6416 & w7664);
assign w7414 = ~w5852 & w3136;
assign w7415 = (w13508 & w1631) | (w13508 & w3681) | (w1631 & w3681);
assign w7416 = ~w9762 & w10590;
assign w7417 = ~w5936 & w13960;
assign w7418 = ~w8425 & w603;
assign w7419 = w1150 & w2248;
assign w7420 = w3508 & ~w5845;
assign w7421 = ~w6993 & w7740;
assign w7422 = (w11861 & w13413) | (w11861 & w11565) | (w13413 & w11565);
assign w7423 = ~w4074 & w3392;
assign w7424 = w3316 & ~w1995;
assign w7425 = ~w3723 & w5162;
assign w7426 = (w1849 & w5076) | (w1849 & w8684) | (w5076 & w8684);
assign w7427 = ~w12148 & w2272;
assign w7428 = (~w12400 & w4691) | (~w12400 & w11271) | (w4691 & w11271);
assign w7429 = (w1223 & w13974) | (w1223 & w2899) | (w13974 & w2899);
assign w7430 = w2858 & ~w9040;
assign w7431 = ~w3067 & w7287;
assign w7432 = w618 & ~w245;
assign w7433 = (w9304 & w14138) | (w9304 & w3678) | (w14138 & w3678);
assign w7434 = (w2410 & w11261) | (w2410 & w4081) | (w11261 & w4081);
assign w7435 = ~w21 & w4105;
assign w7436 = ~w522 & w5618;
assign w7437 = (~w13854 & w11855) | (~w13854 & w2940) | (w11855 & w2940);
assign w7438 = ~w13349 & w7865;
assign w7439 = (~w10709 & w14023) | (~w10709 & w4196) | (w14023 & w4196);
assign w7440 = (w6366 & w7585) | (w6366 & w8228) | (w7585 & w8228);
assign w7441 = w2320 & w560;
assign w7442 = w9170 & w4319;
assign w7443 = w2656 & ~w11108;
assign w7444 = (~w12122 & w6672) | (~w12122 & w8382) | (w6672 & w8382);
assign w7445 = ~w8362 & ~w5739;
assign w7446 = (w1498 & w1855) | (w1498 & w2423) | (w1855 & w2423);
assign w7447 = b17 & a17;
assign w7448 = (w6117 & w3083) | (w6117 & w2667) | (w3083 & w2667);
assign w7449 = ~w5213 & w12804;
assign w7450 = w2288 & w8900;
assign w7451 = ~w12481 & w3727;
assign w7452 = w8096 & ~w8768;
assign w7453 = w8713 & w6785;
assign w7454 = ~w12844 & ~w3033;
assign w7455 = ~w4359 & ~w12943;
assign w7456 = (w154 & w5796) | (w154 & w8461) | (w5796 & w8461);
assign w7457 = (w13772 & w11160) | (w13772 & w5689) | (w11160 & w5689);
assign w7458 = w8450 & w11065;
assign w7459 = ~w13306 & ~w8113;
assign w7460 = (w7774 & w13549) | (w7774 & ~w6637) | (w13549 & ~w6637);
assign w7461 = (w9896 & ~w4336) | (w9896 & w13242) | (~w4336 & w13242);
assign w7462 = ~w13908 & w11537;
assign w7463 = ~w5789 & w11517;
assign w7464 = ~w14659 & ~w1866;
assign w7465 = w4252 | w6266;
assign w7466 = (w9015 & w2144) | (w9015 & w12328) | (w2144 & w12328);
assign w7467 = w230 & w9989;
assign w7468 = ~w9480 & ~w1540;
assign w7469 = (~w11261 & w709) | (~w11261 & w3683) | (w709 & w3683);
assign w7470 = w10483 & w5860;
assign w7471 = ~w1540 & ~w12216;
assign w7472 = w4452 & w2530;
assign w7473 = (w14564 & w11756) | (w14564 & ~w9215) | (w11756 & ~w9215);
assign w7474 = w12131 & ~w10486;
assign w7475 = w3215 & w7645;
assign w7476 = (w5865 & ~w4032) | (w5865 & w5690) | (~w4032 & w5690);
assign w7477 = ~w6268 & ~w11512;
assign w7478 = ~w125 & ~w9046;
assign w7479 = ~w673 & ~w13282;
assign w7480 = (~w1016 & w254) | (~w1016 & w1926) | (w254 & w1926);
assign w7481 = w14147 & w11467;
assign w7482 = w4987 & ~w11655;
assign w7483 = ~w14276 & w3175;
assign w7484 = ~w13900 & ~w6689;
assign w7485 = ~w10075 & ~w11493;
assign w7486 = (~w10032 & w840) | (~w10032 & w8040) | (w840 & w8040);
assign w7487 = ~w14227 & w14072;
assign w7488 = w11510 & ~w14243;
assign w7489 = w9320 & w13578;
assign w7490 = ~b45 & ~a45;
assign w7491 = ~w7207 & w9920;
assign w7492 = w11968 & ~w11773;
assign w7493 = w12330 & w6952;
assign w7494 = w8390 & ~w11636;
assign w7495 = w3922 | ~w7013;
assign w7496 = ~w607 & w11934;
assign w7497 = ~w4887 & w2779;
assign w7498 = w6882 & w7957;
assign w7499 = w790 & w13860;
assign w7500 = w5615 & w8675;
assign w7501 = w7244 & w13323;
assign w7502 = w7662 & w10430;
assign w7503 = w8878 & ~w6828;
assign w7504 = (~w358 & ~w14321) | (~w358 & ~w9305) | (~w14321 & ~w9305);
assign w7505 = (w12533 & w10123) | (w12533 & w106) | (w10123 & w106);
assign w7506 = w11783 & w9703;
assign w7507 = (~w8614 & w6911) | (~w8614 & w6001) | (w6911 & w6001);
assign w7508 = w11906 & w6153;
assign w7509 = (w14453 & w4234) | (w14453 & w14002) | (w4234 & w14002);
assign w7510 = (~w6929 & w10435) | (~w6929 & w12299) | (w10435 & w12299);
assign w7511 = (w2396 & w9131) | (w2396 & w2670) | (w9131 & w2670);
assign w7512 = w10531 & ~w14519;
assign w7513 = ~w4312 & w13214;
assign w7514 = w5864 & w11460;
assign w7515 = (w4679 & w13813) | (w4679 & w10399) | (w13813 & w10399);
assign w7516 = ~w5852 & ~w8898;
assign w7517 = ~w10729 & ~w9038;
assign w7518 = (w9139 & w10988) | (w9139 & w3539) | (w10988 & w3539);
assign w7519 = w5108 & ~w2951;
assign w7520 = (w3039 & w7324) | (w3039 & ~w8791) | (w7324 & ~w8791);
assign w7521 = ~w11198 & ~w9296;
assign w7522 = w9747 & ~w9138;
assign w7523 = (~w8327 & w3329) | (~w8327 & w2479) | (w3329 & w2479);
assign w7524 = w8026 & w10713;
assign w7525 = ~w12228 & w7412;
assign w7526 = w9032 & w10313;
assign w7527 = w13658 & w6028;
assign w7528 = ~w10755 & ~w7741;
assign w7529 = w3038 & w3039;
assign w7530 = w3508 & w9748;
assign w7531 = w14633 & ~w12569;
assign w7532 = ~w7376 & ~w9694;
assign w7533 = (w2310 & w7448) | (w2310 & w9365) | (w7448 & w9365);
assign w7534 = w3671 & ~w5532;
assign w7535 = w11287 & w646;
assign w7536 = (w10210 & w805) | (w10210 & w894) | (w805 & w894);
assign w7537 = (w2159 & w12499) | (w2159 & w13476) | (w12499 & w13476);
assign w7538 = (~w3611 & w5385) | (~w3611 & w4218) | (w5385 & w4218);
assign w7539 = ~w11025 & ~w829;
assign w7540 = (w6310 & w5697) | (w6310 & ~w4033) | (w5697 & ~w4033);
assign w7541 = w7489 & ~w13383;
assign w7542 = w14276 & w8396;
assign w7543 = w2933 & ~w8171;
assign w7544 = (w13924 & w5479) | (w13924 & ~w4527) | (w5479 & ~w4527);
assign w7545 = (w5845 & w5457) | (w5845 & w3115) | (w5457 & w3115);
assign w7546 = ~w1332 & ~w13753;
assign w7547 = ~w2033 & w6714;
assign w7548 = w922 & w1842;
assign w7549 = (~w9707 & ~w14002) | (~w9707 & ~w3721) | (~w14002 & ~w3721);
assign w7550 = ~w5559 & w10436;
assign w7551 = ~w3217 & w13509;
assign w7552 = (w4478 & w6814) | (w4478 & w14618) | (w6814 & w14618);
assign w7553 = ~w13938 & ~w8992;
assign w7554 = (~w6101 & w8079) | (~w6101 & w10369) | (w8079 & w10369);
assign w7555 = (~w13222 & w3750) | (~w13222 & w4138) | (w3750 & w4138);
assign w7556 = ~w1052 & w1692;
assign w7557 = w1372 & ~w10505;
assign w7558 = ~w5288 & w12642;
assign w7559 = w12860 & w6772;
assign w7560 = (w4204 & w1501) | (w4204 & w13331) | (w1501 & w13331);
assign w7561 = w1949 & w829;
assign w7562 = w10699 & ~w8831;
assign w7563 = (~w13526 & w2998) | (~w13526 & ~w1458) | (w2998 & ~w1458);
assign w7564 = w12065 & ~w5247;
assign w7565 = (w14360 & w9311) | (w14360 & w5744) | (w9311 & w5744);
assign w7566 = w11743 & w11694;
assign w7567 = (~w11747 & w4242) | (~w11747 & w7139) | (w4242 & w7139);
assign w7568 = (w8228 & w9034) | (w8228 & w2457) | (w9034 & w2457);
assign w7569 = ~w341 & w1301;
assign w7570 = w6630 | w9702;
assign w7571 = (~w11744 & w344) | (~w11744 & w8241) | (w344 & w8241);
assign w7572 = ~w1785 & w14670;
assign w7573 = w6502 & w5000;
assign w7574 = w12879 & w1217;
assign w7575 = w5212 & w14228;
assign w7576 = ~w7524 & ~w933;
assign w7577 = w12216 & ~w11031;
assign w7578 = (w1871 & ~w11586) | (w1871 & w5953) | (~w11586 & w5953);
assign w7579 = w8337 | w14455;
assign w7580 = (~w11416 & w5917) | (~w11416 & w3706) | (w5917 & w3706);
assign w7581 = (w9095 & w5752) | (w9095 & w378) | (w5752 & w378);
assign w7582 = (~w7423 & w11577) | (~w7423 & w8739) | (w11577 & w8739);
assign w7583 = (w7782 & w7561) | (w7782 & w10347) | (w7561 & w10347);
assign w7584 = (w13733 & ~w1140) | (w13733 & w11659) | (~w1140 & w11659);
assign w7585 = w8367 & ~w14528;
assign w7586 = ~w7630 & w12620;
assign w7587 = ~w10218 & ~w9676;
assign w7588 = w8085 & w12398;
assign w7589 = w12632 & ~w4176;
assign w7590 = w533 & w3401;
assign w7591 = ~w9368 & ~w5920;
assign w7592 = (w10704 & w14664) | (w10704 & w14475) | (w14664 & w14475);
assign w7593 = w12642 & w4483;
assign w7594 = w10491 & ~w14190;
assign w7595 = (~w4341 & ~w8399) | (~w4341 & w787) | (~w8399 & w787);
assign w7596 = (~w4363 & w10356) | (~w4363 & w7112) | (w10356 & w7112);
assign w7597 = w13256 & ~w3587;
assign w7598 = (~w6276 & w2010) | (~w6276 & w11534) | (w2010 & w11534);
assign w7599 = ~w11571 & w9704;
assign w7600 = (~w12775 & w10188) | (~w12775 & w13409) | (w10188 & w13409);
assign w7601 = (w3758 & w6332) | (w3758 & w9034) | (w6332 & w9034);
assign w7602 = w1441 & w12909;
assign w7603 = w6560 & w2717;
assign w7604 = ~w3426 & ~w8362;
assign w7605 = ~w2175 & w1051;
assign w7606 = (~w12464 & ~w157) | (~w12464 & w5037) | (~w157 & w5037);
assign w7607 = w3094 & w6718;
assign w7608 = (w13654 & w1988) | (w13654 & w4566) | (w1988 & w4566);
assign w7609 = (w10477 & w5702) | (w10477 & w7817) | (w5702 & w7817);
assign w7610 = ~w3906 & w1658;
assign w7611 = ~w13850 & w239;
assign w7612 = ~w7329 & ~w13295;
assign w7613 = ~w2762 & w5317;
assign w7614 = w12783 & w719;
assign w7615 = ~w4606 & w11188;
assign w7616 = ~w4959 & w6249;
assign w7617 = (w14340 & w12980) | (w14340 & w13361) | (w12980 & w13361);
assign w7618 = w1062 & ~w1590;
assign w7619 = ~w14199 & ~w271;
assign w7620 = (~w7784 & w2419) | (~w7784 & w7544) | (w2419 & w7544);
assign w7621 = ~w8923 & w14146;
assign w7622 = w13949 & w11720;
assign w7623 = w10930 & ~w6593;
assign w7624 = w2609 & w11718;
assign w7625 = ~w10935 & ~w9333;
assign w7626 = (~w10223 & w13462) | (~w10223 & w9579) | (w13462 & w9579);
assign w7627 = (~w11511 & w6490) | (~w11511 & w9633) | (w6490 & w9633);
assign w7628 = ~w1667 & ~w13240;
assign w7629 = w7525 & ~w12736;
assign w7630 = ~w2467 & ~w13386;
assign w7631 = (w2680 & w12499) | (w2680 & w626) | (w12499 & w626);
assign w7632 = ~w1949 & ~w14542;
assign w7633 = ~w3742 & ~w13306;
assign w7634 = (~w1086 & w4343) | (~w1086 & w865) | (w4343 & w865);
assign w7635 = ~w8937 & w3351;
assign w7636 = ~w8754 & w8018;
assign w7637 = (w11429 & w11558) | (w11429 & w13616) | (w11558 & w13616);
assign w7638 = w2912 & w3281;
assign w7639 = w6275 & w14643;
assign w7640 = (w6277 & w2315) | (w6277 & w8095) | (w2315 & w8095);
assign w7641 = (w13508 & w11175) | (w13508 & w3875) | (w11175 & w3875);
assign w7642 = w12464 & w8972;
assign w7643 = w8280 & ~w7369;
assign w7644 = (w13331 & w2834) | (w13331 & w9331) | (w2834 & w9331);
assign w7645 = (~w1840 & w1360) | (~w1840 & w1224) | (w1360 & w1224);
assign w7646 = w14075 & a53;
assign w7647 = (~w14560 & w9530) | (~w14560 & w3284) | (w9530 & w3284);
assign w7648 = w10545 & ~w8607;
assign w7649 = ~w10116 & ~w4648;
assign w7650 = w3550 & w14536;
assign w7651 = w11451 & ~w1471;
assign w7652 = ~w4512 & w6961;
assign w7653 = (~w10484 & ~w4114) | (~w10484 & w920) | (~w4114 & w920);
assign w7654 = w13872 & w6267;
assign w7655 = ~w13249 & ~w4881;
assign w7656 = (w8827 & w12003) | (w8827 & w12539) | (w12003 & w12539);
assign w7657 = w654 & ~w11089;
assign w7658 = w10676 & w5732;
assign w7659 = ~w11505 & ~w4718;
assign w7660 = ~w142 & ~w3885;
assign w7661 = ~w4700 & w646;
assign w7662 = (~w12170 & w13873) | (~w12170 & w6958) | (w13873 & w6958);
assign w7663 = ~w13473 & w11656;
assign w7664 = (w9950 & w9534) | (w9950 & w21) | (w9534 & w21);
assign w7665 = w11905 & ~w4312;
assign w7666 = w8355 & w13461;
assign w7667 = ~w4458 & w9679;
assign w7668 = ~w12662 & ~w1263;
assign w7669 = w1544 & ~w9687;
assign w7670 = ~w5948 & ~w9927;
assign w7671 = ~w6572 & ~w3158;
assign w7672 = ~w12107 & ~w7754;
assign w7673 = ~w8460 & w13675;
assign w7674 = w6343 & w10198;
assign w7675 = ~w1134 & ~w7257;
assign w7676 = ~w3734 & ~w12138;
assign w7677 = w4755 | w9680;
assign w7678 = (~w2320 & w11546) | (~w2320 & w13029) | (w11546 & w13029);
assign w7679 = ~w12121 & w11487;
assign w7680 = w7528 & ~w4888;
assign w7681 = ~b108 & ~a108;
assign w7682 = w2135 & w11187;
assign w7683 = ~w6147 & w8816;
assign w7684 = ~w9015 & ~w7704;
assign w7685 = w4425 & w5105;
assign w7686 = ~w563 & ~w7252;
assign w7687 = ~w831 & w231;
assign w7688 = w12460 & ~w7746;
assign w7689 = w10708 & ~w1949;
assign w7690 = (w9305 & w2298) | (w9305 & w3073) | (w2298 & w3073);
assign w7691 = (~w2794 & w3239) | (~w2794 & w13851) | (w3239 & w13851);
assign w7692 = w10708 & ~w7839;
assign w7693 = (~w2508 & w13462) | (~w2508 & w13477) | (w13462 & w13477);
assign w7694 = ~w1845 & ~w10182;
assign w7695 = (w807 & w8659) | (w807 & w14128) | (w8659 & w14128);
assign w7696 = w13118 | w217;
assign w7697 = ~w8956 & w11619;
assign w7698 = w3550 & w548;
assign w7699 = (w7757 & w10418) | (w7757 & ~w10033) | (w10418 & ~w10033);
assign w7700 = w5912 & w3099;
assign w7701 = (~w14664 & w1031) | (~w14664 & w3545) | (w1031 & w3545);
assign w7702 = w7771 & w14446;
assign w7703 = w10831 & w216;
assign w7704 = ~w5732 & ~w3502;
assign w7705 = w5912 & w4168;
assign w7706 = w6190 & ~w9846;
assign w7707 = (w3914 & w9289) | (w3914 & w9857) | (w9289 & w9857);
assign w7708 = ~w11762 & w13956;
assign w7709 = w5759 & ~w5385;
assign w7710 = ~w13531 & ~w13114;
assign w7711 = ~w1805 & w8389;
assign w7712 = ~w13349 & w6891;
assign w7713 = (w7410 & w10808) | (w7410 & ~w12154) | (w10808 & ~w12154);
assign w7714 = w3893 & ~w13550;
assign w7715 = w11817 & w12460;
assign w7716 = w10012 & ~w5705;
assign w7717 = (~w11429 & w5585) | (~w11429 & w11265) | (w5585 & w11265);
assign w7718 = ~w13521 & w11117;
assign w7719 = ~w12148 & ~w8096;
assign w7720 = ~w5823 & ~w4199;
assign w7721 = ~w1898 & w632;
assign w7722 = ~w12662 & ~w5556;
assign w7723 = (w11997 & w9748) | (w11997 & w8146) | (w9748 & w8146);
assign w7724 = ~w10221 & ~w3727;
assign w7725 = ~w13130 & w7425;
assign w7726 = (w4671 & w1805) | (w4671 & w5153) | (w1805 & w5153);
assign w7727 = (~w5768 & w3122) | (~w5768 & w13247) | (w3122 & w13247);
assign w7728 = ~w14102 & ~w11115;
assign w7729 = (w11925 & w9229) | (w11925 & w1475) | (w9229 & w1475);
assign w7730 = (~w10719 & w3206) | (~w10719 & w13888) | (w3206 & w13888);
assign w7731 = (w12337 & w9039) | (w12337 & w5952) | (w9039 & w5952);
assign w7732 = w3075 & ~w2675;
assign w7733 = (~w10462 & w13953) | (~w10462 & w1967) | (w13953 & w1967);
assign w7734 = (w6819 & w12596) | (w6819 & ~w269) | (w12596 & ~w269);
assign w7735 = ~w6889 & w14423;
assign w7736 = w7001 & ~w7244;
assign w7737 = ~w10523 & ~w12545;
assign w7738 = ~w11991 & w9742;
assign w7739 = ~w5437 & ~w13689;
assign w7740 = w7428 & w8914;
assign w7741 = w8977 & w3671;
assign w7742 = w5044 & ~w10302;
assign w7743 = ~w7450 & ~w935;
assign w7744 = w12107 & ~w11796;
assign w7745 = w10054 & w6431;
assign w7746 = b93 & ~a93;
assign w7747 = ~w14489 & ~w8990;
assign w7748 = (w4050 & w5225) | (w4050 & w10825) | (w5225 & w10825);
assign w7749 = ~w5702 & w8142;
assign w7750 = w10241 & ~w6691;
assign w7751 = ~w8937 & w9897;
assign w7752 = ~w9769 & w5643;
assign w7753 = w10676 & w12620;
assign w7754 = b37 & a37;
assign w7755 = ~w11079 & w348;
assign w7756 = w3334 & w11297;
assign w7757 = (w8886 & w7756) | (w8886 & w1340) | (w7756 & w1340);
assign w7758 = b93 & w4541;
assign w7759 = ~w7542 & w12417;
assign w7760 = w4114 & w13436;
assign w7761 = (w2938 & w4099) | (w2938 & w2957) | (w4099 & w2957);
assign w7762 = (~w9015 & w5397) | (~w9015 & w7874) | (w5397 & w7874);
assign w7763 = w13845 & w11170;
assign w7764 = ~w5997 & ~w13586;
assign w7765 = (w11934 & w10397) | (w11934 & w8256) | (w10397 & w8256);
assign w7766 = ~w7882 & w7914;
assign w7767 = ~w3276 & w7970;
assign w7768 = b9 & a9;
assign w7769 = w12814 & w3327;
assign w7770 = w9788 & w3366;
assign w7771 = w14235 & w10900;
assign w7772 = ~w12893 & ~w11431;
assign w7773 = (~w12543 & w12614) | (~w12543 & w14208) | (w12614 & w14208);
assign w7774 = (w14573 & w4132) | (w14573 & w10280) | (w4132 & w10280);
assign w7775 = (~w177 & w4209) | (~w177 & w3419) | (w4209 & w3419);
assign w7776 = w10182 & w11934;
assign w7777 = ~w12240 & w3025;
assign w7778 = ~w1563 & w11487;
assign w7779 = ~w9224 & ~w9557;
assign w7780 = (w4692 & w6634) | (w4692 & w7549) | (w6634 & w7549);
assign w7781 = (~w13219 & w5029) | (~w13219 & w14345) | (w5029 & w14345);
assign w7782 = w673 & ~w8046;
assign w7783 = w13914 & w8459;
assign w7784 = ~w11458 & ~w7975;
assign w7785 = ~w3017 & ~w2729;
assign w7786 = ~w6305 & w775;
assign w7787 = w6603 & w2463;
assign w7788 = ~w607 & w9296;
assign w7789 = ~w14407 & ~w8036;
assign w7790 = w6270 & w8672;
assign w7791 = (~w7546 & w11957) | (~w7546 & ~w3564) | (w11957 & ~w3564);
assign w7792 = (w1849 & w10495) | (w1849 & w6109) | (w10495 & w6109);
assign w7793 = w1838 & ~w2729;
assign w7794 = ~w14276 & ~w12371;
assign w7795 = ~w6795 & w8900;
assign w7796 = ~w1305 & ~w9902;
assign w7797 = ~w3019 & w4713;
assign w7798 = w2275 & w4658;
assign w7799 = ~w6963 & ~w8100;
assign w7800 = ~w607 & w4458;
assign w7801 = w7295 & ~w2077;
assign w7802 = (w9698 & w7460) | (w9698 & ~w12376) | (w7460 & ~w12376);
assign w7803 = (w13357 & ~w14012) | (w13357 & w2461) | (~w14012 & w2461);
assign w7804 = ~w13346 & w12755;
assign w7805 = w4798 & ~w13622;
assign w7806 = ~w6126 & w5596;
assign w7807 = w4213 & w3717;
assign w7808 = (~w1838 & w9421) | (~w1838 & w8418) | (w9421 & w8418);
assign w7809 = ~w13558 & w721;
assign w7810 = ~w12262 & w3596;
assign w7811 = ~w2850 & ~w10916;
assign w7812 = w6446 & w10907;
assign w7813 = (w12483 & w5746) | (w12483 & w10915) | (w5746 & w10915);
assign w7814 = w11287 & w4458;
assign w7815 = w894 & ~w7645;
assign w7816 = ~w7276 & ~w12642;
assign w7817 = w1563 & w10477;
assign w7818 = ~w4998 & w11121;
assign w7819 = ~w9925 & w9204;
assign w7820 = w9296 & w8621;
assign w7821 = ~w13526 & ~w11350;
assign w7822 = ~w2984 & ~w14049;
assign w7823 = ~w12842 & w12404;
assign w7824 = (~w7765 & ~w1098) | (~w7765 & w10920) | (~w1098 & w10920);
assign w7825 = (w7914 & w5867) | (w7914 & w10622) | (w5867 & w10622);
assign w7826 = ~w13636 & ~w235;
assign w7827 = (~w12776 & w13447) | (~w12776 & w4149) | (w13447 & w4149);
assign w7828 = ~w5676 & w11477;
assign w7829 = ~w13177 & ~w13442;
assign w7830 = (w2144 & w2411) | (w2144 & w11828) | (w2411 & w11828);
assign w7831 = (w14087 & w3301) | (w14087 & w13207) | (w3301 & w13207);
assign w7832 = w2475 & w10275;
assign w7833 = w13451 & ~w14038;
assign w7834 = w6080 & ~w5761;
assign w7835 = (w4432 & w2310) | (w4432 & ~w8444) | (w2310 & ~w8444);
assign w7836 = ~w2628 & w7072;
assign w7837 = (~w6362 & ~w10328) | (~w6362 & w2900) | (~w10328 & w2900);
assign w7838 = (w7114 & w13487) | (w7114 & ~w12104) | (w13487 & ~w12104);
assign w7839 = w8705 & ~w3313;
assign w7840 = ~w2866 & w5632;
assign w7841 = ~w4707 & ~w7373;
assign w7842 = (w1859 & w5815) | (w1859 & ~w217) | (w5815 & ~w217);
assign w7843 = (w14028 & w2541) | (w14028 & w3669) | (w2541 & w3669);
assign w7844 = ~w10919 & ~w2242;
assign w7845 = w4384 & w3551;
assign w7846 = (w10117 & w4056) | (w10117 & w10680) | (w4056 & w10680);
assign w7847 = (w5062 & w2551) | (w5062 & w12881) | (w2551 & w12881);
assign w7848 = (w13349 & w13149) | (w13349 & w8387) | (w13149 & w8387);
assign w7849 = ~w6803 & w13461;
assign w7850 = ~w12656 & w803;
assign w7851 = ~w3508 & ~w884;
assign w7852 = (~w142 & ~w5761) | (~w142 & w6872) | (~w5761 & w6872);
assign w7853 = (~w894 & w1166) | (~w894 & w7962) | (w1166 & w7962);
assign w7854 = (w1858 & w523) | (w1858 & w11573) | (w523 & w11573);
assign w7855 = (w6572 & w14141) | (w6572 & w5510) | (w14141 & w5510);
assign w7856 = (w7914 & ~w227) | (w7914 & w12302) | (~w227 & w12302);
assign w7857 = w9211 & w11031;
assign w7858 = ~w12271 & w13328;
assign w7859 = w6436 & ~w3904;
assign w7860 = w5817 & ~w11925;
assign w7861 = w6683 & ~w9870;
assign w7862 = w6161 & ~w7296;
assign w7863 = (w1849 & w5905) | (w1849 & w5606) | (w5905 & w5606);
assign w7864 = w7376 & ~w4669;
assign w7865 = ~w5294 & w5732;
assign w7866 = (~w2320 & ~w4032) | (~w2320 & w9921) | (~w4032 & w9921);
assign w7867 = ~w2117 & ~w12390;
assign w7868 = ~w7144 & w3696;
assign w7869 = w3160 & ~w12677;
assign w7870 = w8769 & w10317;
assign w7871 = ~w12394 & w12742;
assign w7872 = (~w14523 & w12003) | (~w14523 & w10199) | (w12003 & w10199);
assign w7873 = w5732 & w8900;
assign w7874 = w5732 & ~w9015;
assign w7875 = ~w636 & ~w3727;
assign w7876 = w10136 | ~w14074;
assign w7877 = ~w8512 & w4127;
assign w7878 = w7159 & w7161;
assign w7879 = (~w13526 & ~w12543) | (~w13526 & w2998) | (~w12543 & w2998);
assign w7880 = ~w7099 & ~w5544;
assign w7881 = ~w4971 & ~w286;
assign w7882 = (~w142 & ~w2729) | (~w142 & w6872) | (~w2729 & w6872);
assign w7883 = w3914 & w7080;
assign w7884 = (~w12042 & ~w13219) | (~w12042 & w8070) | (~w13219 & w8070);
assign w7885 = (~w4099 & w8579) | (~w4099 & w8902) | (w8579 & w8902);
assign w7886 = w11817 & w11500;
assign w7887 = w5867 & w13565;
assign w7888 = w609 & w14603;
assign w7889 = b102 & a102;
assign w7890 = ~w12315 & w3982;
assign w7891 = (w5186 & w4194) | (w5186 & ~w6264) | (w4194 & ~w6264);
assign w7892 = (w14514 & w12118) | (w14514 & w5539) | (w12118 & w5539);
assign w7893 = w8315 & ~w3560;
assign w7894 = w8389 & w4473;
assign w7895 = ~w7782 & w3673;
assign w7896 = ~w8124 & ~w9787;
assign w7897 = (w10916 & w4607) | (w10916 & w6934) | (w4607 & w6934);
assign w7898 = ~w1294 & w6005;
assign w7899 = (~w10500 & w5611) | (~w10500 & w12694) | (w5611 & w12694);
assign w7900 = (w9608 & w9003) | (w9608 & w6987) | (w9003 & w6987);
assign w7901 = ~w4921 & w2034;
assign w7902 = (~w11519 & w12524) | (~w11519 & w1043) | (w12524 & w1043);
assign w7903 = ~w2803 & w3411;
assign w7904 = (~w11167 & w8940) | (~w11167 & w9844) | (w8940 & w9844);
assign w7905 = w4137 & ~w10661;
assign w7906 = ~b77 & ~a77;
assign w7907 = (w2636 & w8997) | (w2636 & w8398) | (w8997 & w8398);
assign w7908 = ~w723 & w9400;
assign w7909 = (w9305 & w1069) | (w9305 & w5368) | (w1069 & w5368);
assign w7910 = ~w9715 & ~w13389;
assign w7911 = (~w3067 & w4536) | (~w3067 & w452) | (w4536 & w452);
assign w7912 = (w8326 & ~w12128) | (w8326 & ~w2868) | (~w12128 & ~w2868);
assign w7913 = (~w1777 & w1338) | (~w1777 & w3307) | (w1338 & w3307);
assign w7914 = ~w3098 & ~w6716;
assign w7915 = ~w6750 & w12662;
assign w7916 = w5768 & w8377;
assign w7917 = (w13331 & w1459) | (w13331 & w3052) | (w1459 & w3052);
assign w7918 = (~w6266 & w13404) | (~w6266 & w2350) | (w13404 & w2350);
assign w7919 = (w9536 & w12086) | (w9536 & w10731) | (w12086 & w10731);
assign w7920 = ~w13222 & ~w5371;
assign w7921 = ~w1241 & w4868;
assign w7922 = w9861 & ~w12983;
assign w7923 = ~w2922 & w8047;
assign w7924 = ~w142 & w7906;
assign w7925 = ~w12856 & ~w7962;
assign w7926 = w3550 & w3324;
assign w7927 = w724 & w6381;
assign w7928 = w4787 & w8454;
assign w7929 = (w122 & ~w5688) | (w122 & ~w11803) | (~w5688 & ~w11803);
assign w7930 = ~w3816 & w10442;
assign w7931 = w4425 & w8389;
assign w7932 = (w10290 & ~w13222) | (w10290 & w7230) | (~w13222 & w7230);
assign w7933 = w14626 & w2473;
assign w7934 = ~w1546 & w10571;
assign w7935 = (~w11488 & w7488) | (~w11488 & w1422) | (w7488 & w1422);
assign w7936 = w5243 & w5569;
assign w7937 = w2873 & w2533;
assign w7938 = (w2777 & w2959) | (w2777 & w9096) | (w2959 & w9096);
assign w7939 = ~w7794 & w2395;
assign w7940 = ~w14588 & ~w13793;
assign w7941 = ~w5936 & ~w2928;
assign w7942 = (~w7103 & ~w3858) | (~w7103 & w13403) | (~w3858 & w13403);
assign w7943 = w3904 & w7376;
assign w7944 = w7808 & w11287;
assign w7945 = w11422 & w5952;
assign w7946 = ~w829 & w10045;
assign w7947 = w3803 & ~w9949;
assign w7948 = w1741 & w8497;
assign w7949 = ~w14141 & w1941;
assign w7950 = w14271 & ~w8996;
assign w7951 = ~w3803 & ~w11361;
assign w7952 = (~w3508 & ~w953) | (~w3508 & w3032) | (~w953 & w3032);
assign w7953 = w3550 & w12797;
assign w7954 = ~w183 & w14659;
assign w7955 = ~w7080 & ~w12891;
assign w7956 = (w12135 & ~w13398) | (w12135 & w4796) | (~w13398 & w4796);
assign w7957 = w3161 & ~w8691;
assign w7958 = (w1764 & w6379) | (w1764 & w9527) | (w6379 & w9527);
assign w7959 = ~w7376 & ~w8827;
assign w7960 = ~w5177 & ~w8085;
assign w7961 = ~w12003 & w11289;
assign w7962 = ~w6542 & ~w894;
assign w7963 = ~w13462 & w10445;
assign w7964 = ~w12464 & w1821;
assign w7965 = ~w7089 & w13725;
assign w7966 = (w7317 & w12614) | (w7317 & w4908) | (w12614 & w4908);
assign w7967 = ~w5562 & w10691;
assign w7968 = ~w5558 & ~w6904;
assign w7969 = w2307 & w9989;
assign w7970 = ~w14376 & w9049;
assign w7971 = w13612 & w14256;
assign w7972 = (w12172 & w9463) | (w12172 & w12376) | (w9463 & w12376);
assign w7973 = ~w4700 & w3550;
assign w7974 = ~w11415 & ~w11603;
assign w7975 = ~w8937 & w9632;
assign w7976 = ~w12753 & ~w56;
assign w7977 = ~w1166 & ~w11457;
assign w7978 = w6135 & ~w11934;
assign w7979 = ~w13349 & w14220;
assign w7980 = w1516 & ~w11345;
assign w7981 = ~w9623 & w5412;
assign w7982 = w6566 & w8549;
assign w7983 = (w13047 & ~w10845) | (w13047 & w12967) | (~w10845 & w12967);
assign w7984 = w8920 & ~w2179;
assign w7985 = (w3017 & w13623) | (w3017 & w5978) | (w13623 & w5978);
assign w7986 = w7670 & w14097;
assign w7987 = (w3215 & ~w953) | (w3215 & w10417) | (~w953 & w10417);
assign w7988 = ~w607 & ~w3904;
assign w7989 = (w10449 & w5324) | (w10449 & w2287) | (w5324 & w2287);
assign w7990 = w8762 & w13329;
assign w7991 = w2225 & w13049;
assign w7992 = (~w4515 & w8693) | (~w4515 & w11723) | (w8693 & w11723);
assign w7993 = ~w13222 & ~w4050;
assign w7994 = w12879 & w10708;
assign w7995 = (w3192 & w14456) | (w3192 & w5298) | (w14456 & w5298);
assign w7996 = (~w4127 & w12121) | (~w4127 & w11224) | (w12121 & w11224);
assign w7997 = ~w9296 & w9925;
assign w7998 = (w9989 & w4095) | (w9989 & w7334) | (w4095 & w7334);
assign w7999 = (~w11915 & w12125) | (~w11915 & w10779) | (w12125 & w10779);
assign w8000 = (~w1939 & w10116) | (~w1939 & w1986) | (w10116 & w1986);
assign w8001 = ~w9583 & ~w13628;
assign w8002 = (w5243 & w7936) | (w5243 & ~w5569) | (w7936 & ~w5569);
assign w8003 = ~w5288 & w6500;
assign w8004 = w13222 & w6572;
assign w8005 = (~w5078 & w7708) | (~w5078 & w8359) | (w7708 & w8359);
assign w8006 = (w8327 & w12166) | (w8327 & w9930) | (w12166 & w9930);
assign w8007 = (~w5498 & w10350) | (~w5498 & w666) | (w10350 & w666);
assign w8008 = ~w11893 & w7914;
assign w8009 = (w1540 & w7981) | (w1540 & w9522) | (w7981 & w9522);
assign w8010 = w1646 & ~w12988;
assign w8011 = (~w13008 & w9506) | (~w13008 & w12553) | (w9506 & w12553);
assign w8012 = w11779 & ~w2493;
assign w8013 = ~b14 & ~a14;
assign w8014 = ~w1025 & ~w6070;
assign w8015 = w10967 & w4335;
assign w8016 = w2701 & ~w8294;
assign w8017 = w5406 & ~w8512;
assign w8018 = w10514 & w5213;
assign w8019 = ~w10906 & w10039;
assign w8020 = (w5084 & w3357) | (w5084 & w6310) | (w3357 & w6310);
assign w8021 = ~w12271 & w13761;
assign w8022 = w1062 & w11708;
assign w8023 = (w8890 & w11845) | (w8890 & w12358) | (w11845 & w12358);
assign w8024 = ~w8760 & w5132;
assign w8025 = w5884 & w9989;
assign w8026 = ~w10490 & ~w261;
assign w8027 = w4380 & w3950;
assign w8028 = ~w2509 & ~w7486;
assign w8029 = w5761 & ~w10851;
assign w8030 = (w3586 & ~w9197) | (w3586 & w12032) | (~w9197 & w12032);
assign w8031 = ~w2938 & w3823;
assign w8032 = (w13434 & ~w13219) | (w13434 & w2903) | (~w13219 & w2903);
assign w8033 = w2096 & w8863;
assign w8034 = w13521 & ~w7490;
assign w8035 = b78 & a78;
assign w8036 = w10042 & w8900;
assign w8037 = ~w881 & ~w11564;
assign w8038 = w5912 & w3904;
assign w8039 = ~w8049 & ~w12535;
assign w8040 = w8183 & ~w10032;
assign w8041 = ~w12271 & ~w7762;
assign w8042 = w4836 & ~w12915;
assign w8043 = (~w3158 & w183) | (~w3158 & w4932) | (w183 & w4932);
assign w8044 = w1098 & w3235;
assign w8045 = ~w8475 & ~w5545;
assign w8046 = w7794 & w6835;
assign w8047 = ~w8328 & ~w7365;
assign w8048 = w9679 & w8813;
assign w8049 = ~w607 & w5761;
assign w8050 = w5781 & ~w3423;
assign w8051 = ~w297 & w2907;
assign w8052 = ~w9608 & w1211;
assign w8053 = ~w12121 & w8390;
assign w8054 = (w14463 & w1160) | (w14463 & w678) | (w1160 & w678);
assign w8055 = w8831 & w8396;
assign w8056 = w12922 & ~w6951;
assign w8057 = w5913 & ~w5798;
assign w8058 = w5556 & ~w1712;
assign w8059 = (w9075 & w4923) | (w9075 & w1045) | (w4923 & w1045);
assign w8060 = w6538 & ~w6190;
assign w8061 = ~w6832 & w3845;
assign w8062 = (~w10435 & w9516) | (~w10435 & w14192) | (w9516 & w14192);
assign w8063 = ~w6436 & ~w3427;
assign w8064 = ~w13462 & w1567;
assign w8065 = (~w1862 & ~w7006) | (~w1862 & w7010) | (~w7006 & w7010);
assign w8066 = w11482 & w6554;
assign w8067 = ~w1139 & w4866;
assign w8068 = ~w7013 & w2941;
assign w8069 = w2711 & ~w3335;
assign w8070 = w1608 & ~w12042;
assign w8071 = ~w1727 & ~w3602;
assign w8072 = ~w14137 & ~w21;
assign w8073 = (~w10525 & ~w6953) | (~w10525 & w7377) | (~w6953 & w7377);
assign w8074 = (w13924 & ~w1563) | (w13924 & w576) | (~w1563 & w576);
assign w8075 = w14048 & w11940;
assign w8076 = ~w7464 & ~w5140;
assign w8077 = (~w4149 & w1170) | (~w4149 & w12245) | (w1170 & w12245);
assign w8078 = ~w12464 & w6542;
assign w8079 = (w1293 & w4717) | (w1293 & ~w1055) | (w4717 & ~w1055);
assign w8080 = (~w3717 & ~w14504) | (~w3717 & w2160) | (~w14504 & w2160);
assign w8081 = (~w254 & w13078) | (~w254 & w11685) | (w13078 & w11685);
assign w8082 = (~w1919 & ~w2656) | (~w1919 & w3408) | (~w2656 & w3408);
assign w8083 = w11118 & ~w8103;
assign w8084 = ~w3180 & ~w10104;
assign w8085 = ~w3502 & ~w9015;
assign w8086 = (~w6781 & w14549) | (~w6781 & w11319) | (w14549 & w11319);
assign w8087 = w13590 & w402;
assign w8088 = ~w4050 & w4567;
assign w8089 = w8246 & w11295;
assign w8090 = ~w5702 & w1462;
assign w8091 = (w5282 & w968) | (w5282 & w10716) | (w968 & w10716);
assign w8092 = ~w3038 & w5612;
assign w8093 = ~w2218 & w2731;
assign w8094 = ~w473 & ~w2493;
assign w8095 = ~w9433 & w6277;
assign w8096 = b27 & a27;
assign w8097 = w14116 & ~w3895;
assign w8098 = w607 & w13839;
assign w8099 = ~w4269 & ~w3447;
assign w8100 = ~w11431 & w9159;
assign w8101 = ~w2371 & ~w11032;
assign w8102 = ~w4835 & w116;
assign w8103 = (w13565 & ~w3550) | (w13565 & w8994) | (~w3550 & w8994);
assign w8104 = (~w12464 & ~w13805) | (~w12464 & w9951) | (~w13805 & w9951);
assign w8105 = ~w142 & ~w12460;
assign w8106 = ~w1207 & w13986;
assign w8107 = ~w12240 & w3019;
assign w8108 = w7484 & ~w6217;
assign w8109 = w10315 & w13886;
assign w8110 = ~b49 & ~a49;
assign w8111 = (~w13628 & w9012) | (~w13628 & w333) | (w9012 & w333);
assign w8112 = w7847 & ~w14145;
assign w8113 = ~w9623 & ~w3742;
assign w8114 = (~w5243 & w3146) | (~w5243 & w9298) | (w3146 & w9298);
assign w8115 = w11500 & ~w6888;
assign w8116 = w8475 & w6689;
assign w8117 = (w3721 & w8129) | (w3721 & w7251) | (w8129 & w7251);
assign w8118 = w3550 & w13573;
assign w8119 = w260 & ~w11031;
assign w8120 = ~w5108 & ~w2951;
assign w8121 = w13084 & ~w7217;
assign w8122 = ~w1692 & ~w10410;
assign w8123 = w7653 & ~w2961;
assign w8124 = ~w12980 & w12242;
assign w8125 = (~w3727 & w1900) | (~w3727 & w2996) | (w1900 & w2996);
assign w8126 = ~w4175 & ~w5442;
assign w8127 = w1500 & w4183;
assign w8128 = w7447 & w11117;
assign w8129 = w8737 & ~w12528;
assign w8130 = w13140 & ~w1254;
assign w8131 = ~w8959 & ~w4493;
assign w8132 = (w3550 & w11323) | (w3550 & w13314) | (w11323 & w13314);
assign w8133 = ~w235 & ~w11606;
assign w8134 = ~w6388 & ~w10788;
assign w8135 = ~w9435 & w12832;
assign w8136 = ~w12614 & w13526;
assign w8137 = w4213 & ~w2544;
assign w8138 = w13604 & w520;
assign w8139 = w8827 & ~w11395;
assign w8140 = (~w1404 & w6426) | (~w1404 & w7311) | (w6426 & w7311);
assign w8141 = ~w4023 & w8936;
assign w8142 = ~w1563 & w2410;
assign w8143 = w1274 & w14307;
assign w8144 = w10951 & ~w3325;
assign w8145 = ~w12121 & w9015;
assign w8146 = ~w11604 & w11108;
assign w8147 = (w11708 & ~w14302) | (w11708 & w8331) | (~w14302 & w8331);
assign w8148 = (~w2039 & w7735) | (~w2039 & w2932) | (w7735 & w2932);
assign w8149 = (w5282 & w843) | (w5282 & w10827) | (w843 & w10827);
assign w8150 = ~w10309 & w3581;
assign w8151 = (w7317 & w5294) | (w7317 & w3836) | (w5294 & w3836);
assign w8152 = ~w3738 & ~w7608;
assign w8153 = (w1190 & w12007) | (w1190 & w267) | (w12007 & w267);
assign w8154 = w12330 & w1114;
assign w8155 = w2401 & w13192;
assign w8156 = ~w4592 & ~w1851;
assign w8157 = ~w7100 & w3020;
assign w8158 = w1644 & ~w10027;
assign w8159 = ~w1434 & ~w14036;
assign w8160 = w4137 & w14430;
assign w8161 = ~w4497 & w3963;
assign w8162 = ~w9875 & ~w2529;
assign w8163 = (~w353 & w10318) | (~w353 & w9403) | (w10318 & w9403);
assign w8164 = w5231 & w13426;
assign w8165 = ~w11428 & w14194;
assign w8166 = w12135 & ~w2685;
assign w8167 = w13432 | w4771;
assign w8168 = (~w6802 & w3266) | (~w6802 & w5007) | (w3266 & w5007);
assign w8169 = w1660 & w10323;
assign w8170 = w2680 & ~w2492;
assign w8171 = b88 & a88;
assign w8172 = w11108 & w8737;
assign w8173 = w5532 & w6572;
assign w8174 = ~w9871 & w12528;
assign w8175 = ~w3790 & ~w5301;
assign w8176 = ~w11429 & w9584;
assign w8177 = w10285 & w3498;
assign w8178 = (w11264 & ~w1712) | (w11264 & w6218) | (~w1712 & w6218);
assign w8179 = (~w10116 & w2492) | (~w10116 & w10301) | (w2492 & w10301);
assign w8180 = w10265 & w13485;
assign w8181 = w11500 & ~w13643;
assign w8182 = w3671 & ~w7401;
assign w8183 = ~b113 & ~a113;
assign w8184 = (w9023 & w1376) | (w9023 & w49) | (w1376 & w49);
assign w8185 = (w6879 & w11712) | (w6879 & w4342) | (w11712 & w4342);
assign w8186 = (~w4099 & w8716) | (~w4099 & w10215) | (w8716 & w10215);
assign w8187 = w505 & w3727;
assign w8188 = w7109 & w399;
assign w8189 = (~w2467 & ~w10436) | (~w2467 & w13879) | (~w10436 & w13879);
assign w8190 = (w9007 & w3391) | (w9007 & w3266) | (w3391 & w3266);
assign w8191 = ~w10477 & ~w5406;
assign w8192 = (~w10123 & w10873) | (~w10123 & w10110) | (w10873 & w10110);
assign w8193 = w4153 & w1314;
assign w8194 = w11934 & ~w1367;
assign w8195 = ~w12040 & ~w9811;
assign w8196 = w12464 & ~w13222;
assign w8197 = w6506 & ~w14566;
assign w8198 = w12528 & ~w11516;
assign w8199 = ~w2492 & ~w6949;
assign w8200 = w14588 & ~w6689;
assign w8201 = w13201 & ~w11858;
assign w8202 = ~w674 & w13332;
assign w8203 = (w2035 & ~w4531) | (w2035 & w5198) | (~w4531 & w5198);
assign w8204 = (w6935 & w11191) | (w6935 & w14002) | (w11191 & w14002);
assign w8205 = w6281 & w4287;
assign w8206 = w10676 & w8390;
assign w8207 = ~w8874 & w282;
assign w8208 = ~w14302 & w3508;
assign w8209 = (w1692 & w1279) | (w1692 & w9203) | (w1279 & w9203);
assign w8210 = ~w10153 & ~w12923;
assign w8211 = (w2410 & w10462) | (w2410 & w4397) | (w10462 & w4397);
assign w8212 = w5412 & ~w3289;
assign w8213 = ~w7782 & w13055;
assign w8214 = (w8513 & w9541) | (w8513 & w5799) | (w9541 & w5799);
assign w8215 = ~w14607 & ~w7738;
assign w8216 = ~w3088 & ~w3163;
assign w8217 = w8737 & w6797;
assign w8218 = ~w922 & w3098;
assign w8219 = (w10174 & w13975) | (w10174 & w3559) | (w13975 & w3559);
assign w8220 = (w8859 & w5923) | (w8859 & w2091) | (w5923 & w2091);
assign w8221 = ~w5620 & w9672;
assign w8222 = w922 & ~w4129;
assign w8223 = w7369 & w3963;
assign w8224 = (~w11108 & w4099) | (~w11108 & w7443) | (w4099 & w7443);
assign w8225 = ~w13282 & ~w13938;
assign w8226 = w8817 & ~w6942;
assign w8227 = w13650 & ~w7639;
assign w8228 = (w1171 & ~w11699) | (w1171 & w10557) | (~w11699 & w10557);
assign w8229 = (w13263 & w8340) | (w13263 & w5012) | (w8340 & w5012);
assign w8230 = w9219 & ~w6296;
assign w8231 = w7045 & w6340;
assign w8232 = (~w1254 & w1984) | (~w1254 & w9727) | (w1984 & w9727);
assign w8233 = w10898 & w7789;
assign w8234 = ~w12671 & ~w3077;
assign w8235 = (w13772 & w903) | (w13772 & w3109) | (w903 & w3109);
assign w8236 = ~w13991 & w6168;
assign w8237 = (~w3219 & ~w2850) | (~w3219 & w3433) | (~w2850 & w3433);
assign w8238 = (~w12528 & ~w3383) | (~w12528 & w11759) | (~w3383 & w11759);
assign w8239 = (w11329 & ~w12488) | (w11329 & w4827) | (~w12488 & w4827);
assign w8240 = (~w4287 & w1860) | (~w4287 & w10384) | (w1860 & w10384);
assign w8241 = (w13596 & w1933) | (w13596 & w5456) | (w1933 & w5456);
assign w8242 = ~w5177 & w11488;
assign w8243 = w4290 & w6979;
assign w8244 = (~w4458 & ~w4193) | (~w4458 & w5314) | (~w4193 & w5314);
assign w8245 = (w12569 & ~w7630) | (w12569 & w1217) | (~w7630 & w1217);
assign w8246 = (w3067 & w8954) | (w3067 & w13021) | (w8954 & w13021);
assign w8247 = w7400 & ~w4033;
assign w8248 = ~w5823 & ~w1106;
assign w8249 = ~w11189 & w14089;
assign w8250 = ~w8889 & w11062;
assign w8251 = w5419 & w4462;
assign w8252 = (~w6266 & w12003) | (~w6266 & w1946) | (w12003 & w1946);
assign w8253 = b109 & a109;
assign w8254 = w14276 & w11861;
assign w8255 = (~w3139 & w12687) | (~w3139 & w5092) | (w12687 & w5092);
assign w8256 = (w11934 & w4501) | (w11934 & w1672) | (w4501 & w1672);
assign w8257 = w14263 & ~w9815;
assign w8258 = (~w11216 & w6888) | (~w11216 & w624) | (w6888 & w624);
assign w8259 = w8576 & ~w2089;
assign w8260 = (~w13645 & w6230) | (~w13645 & w5130) | (w6230 & w5130);
assign w8261 = ~w4756 & w12874;
assign w8262 = w12958 & w11500;
assign w8263 = w3786 & w11117;
assign w8264 = ~w5620 & ~w5694;
assign w8265 = ~w12315 & ~w300;
assign w8266 = w14116 & ~w11092;
assign w8267 = w10422 & w1792;
assign w8268 = ~w5299 & w1477;
assign w8269 = w2656 & w10409;
assign w8270 = w13576 & w8535;
assign w8271 = ~w10618 & w12428;
assign w8272 = w11361 & ~w3751;
assign w8273 = ~w6993 & w12008;
assign w8274 = w894 & ~w10477;
assign w8275 = ~w11222 & w13647;
assign w8276 = ~w2807 & w3517;
assign w8277 = ~w10824 & ~w10722;
assign w8278 = (~w14395 & w5852) | (~w14395 & w5262) | (w5852 & w5262);
assign w8279 = (w3550 & w13820) | (w3550 & w5247) | (w13820 & w5247);
assign w8280 = ~b107 & ~a107;
assign w8281 = ~w9708 & ~w6656;
assign w8282 = ~w5231 & ~w9403;
assign w8283 = ~w4050 & w3774;
assign w8284 = (w2535 & w7595) | (w2535 & w996) | (w7595 & w996);
assign w8285 = w9183 & w13328;
assign w8286 = ~w9628 & ~w11938;
assign w8287 = w7190 & ~w7630;
assign w8288 = (w11385 & w5940) | (w11385 & w13898) | (w5940 & w13898);
assign w8289 = ~w2317 & w1558;
assign w8290 = (~w803 & w1809) | (~w803 & w10754) | (w1809 & w10754);
assign w8291 = ~w4215 & ~w359;
assign w8292 = w10001 & w601;
assign w8293 = (~w7782 & w4668) | (~w7782 & w11301) | (w4668 & w11301);
assign w8294 = (~w7335 & w12479) | (~w7335 & w6066) | (w12479 & w6066);
assign w8295 = ~w9012 & w1922;
assign w8296 = ~w11855 & w10045;
assign w8297 = w12714 & ~w2951;
assign w8298 = (w9305 & w10314) | (w9305 & w10747) | (w10314 & w10747);
assign w8299 = (w137 & w9614) | (w137 & w287) | (w9614 & w287);
assign w8300 = (w6486 & w9450) | (w6486 & ~w7062) | (w9450 & ~w7062);
assign w8301 = ~w142 & ~w7670;
assign w8302 = ~w4700 & w8459;
assign w8303 = w4756 & w7220;
assign w8304 = w10949 & ~w6580;
assign w8305 = w8253 & w5761;
assign w8306 = ~w6420 & w2772;
assign w8307 = ~w1624 & w3666;
assign w8308 = w13654 & ~w4172;
assign w8309 = w5867 & w3977;
assign w8310 = w4213 & w5860;
assign w8311 = (w12406 & w6827) | (w12406 & w7560) | (w6827 & w7560);
assign w8312 = w5490 & ~w8814;
assign w8313 = w7914 & ~w14302;
assign w8314 = w8584 & w7317;
assign w8315 = w6475 & w1446;
assign w8316 = ~w1166 & w4359;
assign w8317 = ~w1280 & ~w8493;
assign w8318 = w9809 & w12340;
assign w8319 = (~w13743 & w10151) | (~w13743 & w11865) | (w10151 & w11865);
assign w8320 = w13439 & ~w13146;
assign w8321 = (w12088 & ~w6042) | (w12088 & w12074) | (~w6042 & w12074);
assign w8322 = (~w4709 & w6207) | (~w4709 & w3559) | (w6207 & w3559);
assign w8323 = (w12884 & w8580) | (w12884 & w3759) | (w8580 & w3759);
assign w8324 = ~w10781 & w13495;
assign w8325 = ~w13188 & w3035;
assign w8326 = (w14532 & w5701) | (w14532 & w6076) | (w5701 & w6076);
assign w8327 = (~w13240 & ~w7193) | (~w13240 & w9440) | (~w7193 & w9440);
assign w8328 = b92 & a92;
assign w8329 = w10136 | ~w7644;
assign w8330 = ~w10600 & ~w12208;
assign w8331 = w11708 & ~w6542;
assign w8332 = (w2275 & w8630) | (w2275 & w2827) | (w8630 & w2827);
assign w8333 = ~w2507 & ~w2329;
assign w8334 = ~w7082 & w3585;
assign w8335 = w7349 & ~w4509;
assign w8336 = w8580 | w12884;
assign w8337 = (w7464 & w14455) | (w7464 & w8479) | (w14455 & w8479);
assign w8338 = ~w4700 & ~w3727;
assign w8339 = ~w2864 & w6459;
assign w8340 = (w13263 & w12220) | (w13263 & w6658) | (w12220 & w6658);
assign w8341 = ~w9004 & w225;
assign w8342 = ~w1166 & w9871;
assign w8343 = (w683 & w13219) | (w683 & w4891) | (w13219 & w4891);
assign w8344 = ~w12394 & w6319;
assign w8345 = ~w2927 & ~w11285;
assign w8346 = ~w2715 & ~w872;
assign w8347 = ~w3885 & ~w9788;
assign w8348 = w13161 & w4224;
assign w8349 = (w453 & w9012) | (w453 & w5797) | (w9012 & w5797);
assign w8350 = ~w2081 & ~w13564;
assign w8351 = ~w2427 & ~w8656;
assign w8352 = (w11708 & w10676) | (w11708 & w9376) | (w10676 & w9376);
assign w8353 = w13694 & w11940;
assign w8354 = (~w14395 & w183) | (~w14395 & w5262) | (w183 & w5262);
assign w8355 = ~w12330 & w13461;
assign w8356 = ~w8929 & w3852;
assign w8357 = w4647 & ~w4926;
assign w8358 = ~w8638 & ~w5524;
assign w8359 = ~w13469 & ~w5078;
assign w8360 = w1949 & w10708;
assign w8361 = ~w14389 & w8459;
assign w8362 = ~w2323 & w13953;
assign w8363 = w11673 & ~w11242;
assign w8364 = ~w7221 & w8792;
assign w8365 = ~w10691 & w3764;
assign w8366 = w11441 & w4517;
assign w8367 = ~w8512 & w3038;
assign w8368 = ~w12601 & w9627;
assign w8369 = (w1115 & ~w12649) | (w1115 & w3263) | (~w12649 & w3263);
assign w8370 = ~b15 & ~a15;
assign w8371 = w9453 & ~w14072;
assign w8372 = (w3090 & w9743) | (w3090 & w11599) | (w9743 & w11599);
assign w8373 = ~w10824 & w1404;
assign w8374 = w3019 & w7630;
assign w8375 = ~w9657 & w2999;
assign w8376 = ~w9253 & w223;
assign w8377 = ~w5045 | ~w4042;
assign w8378 = ~w2968 & ~w12758;
assign w8379 = w2583 & ~w10793;
assign w8380 = w4787 & ~w13953;
assign w8381 = w13223 & w4440;
assign w8382 = (~w3904 & w9202) | (~w3904 & w8785) | (w9202 & w8785);
assign w8383 = (~w7022 & w6128) | (~w7022 & w5662) | (w6128 & w5662);
assign w8384 = ~w13152 & w3961;
assign w8385 = (~w5952 & w1998) | (~w5952 & w14434) | (w1998 & w14434);
assign w8386 = w6346 & w5096;
assign w8387 = (~w6716 & w7472) | (~w6716 & w5294) | (w7472 & w5294);
assign w8388 = (~w142 & ~w5282) | (~w142 & w6872) | (~w5282 & w6872);
assign w8389 = (~w13282 & w11848) | (~w13282 & w7479) | (w11848 & w7479);
assign w8390 = ~w8512 & ~w14178;
assign w8391 = ~w1048 & w11746;
assign w8392 = ~w13636 & ~w11606;
assign w8393 = w6502 & w5362;
assign w8394 = ~w10645 & ~w3777;
assign w8395 = ~w9845 & ~w12121;
assign w8396 = ~w6190 & ~w6580;
assign w8397 = w13612 & w12745;
assign w8398 = ~w6127 & w2636;
assign w8399 = (w12685 & ~w11723) | (w12685 & ~w10433) | (~w11723 & ~w10433);
assign w8400 = w7645 & ~w13352;
assign w8401 = ~w6500 & ~w9315;
assign w8402 = w6328 & w10713;
assign w8403 = ~w4190 & w11959;
assign w8404 = ~w13423 & ~w11117;
assign w8405 = (w4545 & w8580) | (w4545 & w14534) | (w8580 & w14534);
assign w8406 = (w5769 & w5207) | (w5769 & ~w12330) | (w5207 & ~w12330);
assign w8407 = w8900 & ~w5308;
assign w8408 = ~w3665 & ~w13407;
assign w8409 = ~w12738 & ~w12223;
assign w8410 = ~w10696 & ~w3454;
assign w8411 = w12460 & ~w9660;
assign w8412 = ~w9715 & w9672;
assign w8413 = w675 & w10095;
assign w8414 = w6189 & ~w14225;
assign w8415 = w12636 & w7896;
assign w8416 = w1764 & w13665;
assign w8417 = ~w12509 & w8878;
assign w8418 = w7369 & ~w1838;
assign w8419 = ~w5660 & w6803;
assign w8420 = ~w217 & w1540;
assign w8421 = w6427 & ~w4021;
assign w8422 = ~w10334 & ~w1151;
assign w8423 = (w6802 & w782) | (w6802 & w3772) | (w782 & w3772);
assign w8424 = (w10318 & ~w353) | (w10318 & ~w5007) | (~w353 & ~w5007);
assign w8425 = (w3957 & w999) | (w3957 & w13437) | (w999 & w13437);
assign w8426 = ~w7455 & w14270;
assign w8427 = ~w4814 & ~w3980;
assign w8428 = (w2040 & w14221) | (w2040 & ~w13980) | (w14221 & ~w13980);
assign w8429 = w1642 & ~w2492;
assign w8430 = w14129 & ~w828;
assign w8431 = ~w7631 & ~w12227;
assign w8432 = (w302 & w570) | (w302 & w8526) | (w570 & w8526);
assign w8433 = ~w6083 & ~w1003;
assign w8434 = ~w5297 & w10787;
assign w8435 = ~w13587 & w13014;
assign w8436 = ~w1835 & w1222;
assign w8437 = ~w8839 & ~w8720;
assign w8438 = w1122 & ~w816;
assign w8439 = w1373 & w13923;
assign w8440 = ~w4115 & ~w2973;
assign w8441 = (w11594 & w2359) | (w11594 & w1865) | (w2359 & w1865);
assign w8442 = (~w5406 & w621) | (~w5406 & w10538) | (w621 & w10538);
assign w8443 = ~w9788 & ~w3427;
assign w8444 = ~w9262 & w4952;
assign w8445 = ~w6135 & w5282;
assign w8446 = w262 & w2924;
assign w8447 = ~w6778 & ~w10884;
assign w8448 = ~w5778 & w5446;
assign w8449 = ~w13880 & w3315;
assign w8450 = (w3128 & w4536) | (w3128 & w4828) | (w4536 & w4828);
assign w8451 = (w10486 & w9798) | (w10486 & w749) | (w9798 & w749);
assign w8452 = ~w922 & w1821;
assign w8453 = (w4405 & w3277) | (w4405 & w6451) | (w3277 & w6451);
assign w8454 = w12656 & ~w12170;
assign w8455 = (w2317 & w8709) | (w2317 & w12704) | (w8709 & w12704);
assign w8456 = ~w12876 & w10591;
assign w8457 = (w7267 & ~w7223) | (w7267 & w7126) | (~w7223 & w7126);
assign w8458 = (w2620 & w5215) | (w2620 & w11516) | (w5215 & w11516);
assign w8459 = ~w706 & ~w7305;
assign w8460 = w12415 & w8141;
assign w8461 = (w1416 & w6276) | (w1416 & w9034) | (w6276 & w9034);
assign w8462 = w7813 & ~w13378;
assign w8463 = w4458 & w6689;
assign w8464 = ~w8512 & w7762;
assign w8465 = w12135 & w2531;
assign w8466 = w991 & ~w2253;
assign w8467 = (w2354 & w14371) | (w2354 & w12154) | (w14371 & w12154);
assign w8468 = w8465 & w9505;
assign w8469 = (~w142 & ~w646) | (~w142 & w6872) | (~w646 & w6872);
assign w8470 = ~w12240 & w2425;
assign w8471 = w1166 & ~w11855;
assign w8472 = ~w11959 & ~w4587;
assign w8473 = (~w724 & w254) | (~w724 & w4758) | (w254 & w4758);
assign w8474 = w7365 & ~w8793;
assign w8475 = b112 & a112;
assign w8476 = w11934 & ~w200;
assign w8477 = ~w4472 & w970;
assign w8478 = ~w12240 & w4473;
assign w8479 = w3447 & w4656;
assign w8480 = ~w12003 & w10043;
assign w8481 = ~w12429 & w4203;
assign w8482 = ~w7437 & ~w12170;
assign w8483 = w13923 & ~w2290;
assign w8484 = ~w1498 & w695;
assign w8485 = (w9032 & w3069) | (w9032 & ~w183) | (w3069 & ~w183);
assign w8486 = ~w5898 & w7647;
assign w8487 = ~w2252 & w14216;
assign w8488 = ~w1838 & ~w1845;
assign w8489 = w4105 & w10256;
assign w8490 = (~w6215 & w4390) | (~w6215 & w3245) | (w4390 & w3245);
assign w8491 = w10032 & ~w988;
assign w8492 = ~w5294 & w2320;
assign w8493 = (w1039 & w3259) | (w1039 & w11258) | (w3259 & w11258);
assign w8494 = ~w5701 & w1807;
assign w8495 = ~w4175 & w13246;
assign w8496 = (~w13375 & ~w5498) | (~w13375 & w3015) | (~w5498 & w3015);
assign w8497 = (w11106 & w14229) | (w11106 & ~w9749) | (w14229 & ~w9749);
assign w8498 = w9060 & ~w3209;
assign w8499 = w13620 & w4266;
assign w8500 = (w9467 & w3783) | (w9467 & ~w14182) | (w3783 & ~w14182);
assign w8501 = (w12768 & w5494) | (w12768 & w1776) | (w5494 & w1776);
assign w8502 = ~w6889 & ~w10861;
assign w8503 = ~w1358 & w879;
assign w8504 = ~w6946 & ~w14556;
assign w8505 = w12460 & w13732;
assign w8506 = (w976 & w8515) | (w976 & ~w10023) | (w8515 & ~w10023);
assign w8507 = (w8389 & w13979) | (w8389 & w8759) | (w13979 & w8759);
assign w8508 = w12943 & ~w7645;
assign w8509 = w3963 & w5545;
assign w8510 = w12077 & w13030;
assign w8511 = w7459 & ~w11861;
assign w8512 = b64 & a64;
assign w8513 = w8047 & w11817;
assign w8514 = (w4759 & w2111) | (w4759 & w12376) | (w2111 & w12376);
assign w8515 = (w378 & w11178) | (w378 & w11305) | (w11178 & w11305);
assign w8516 = ~w9453 & ~w14227;
assign w8517 = w12662 & w9921;
assign w8518 = ~w235 & w8786;
assign w8519 = w1646 & ~w13700;
assign w8520 = ~w3503 & ~w988;
assign w8521 = w3508 & w12088;
assign w8522 = (~w888 & w2455) | (~w888 & w3669) | (w2455 & w3669);
assign w8523 = (w7914 & w13479) | (w7914 & w11705) | (w13479 & w11705);
assign w8524 = (w7757 & w10418) | (w7757 & w9096) | (w10418 & w9096);
assign w8525 = w11722 & ~w11098;
assign w8526 = (w9881 & w1438) | (w9881 & w14182) | (w1438 & w14182);
assign w8527 = ~w921 & ~w5056;
assign w8528 = ~w607 & ~w3098;
assign w8529 = ~w4193 & ~w6080;
assign w8530 = (~w5641 & ~w1362) | (~w5641 & w1386) | (~w1362 & w1386);
assign w8531 = w7270 & ~w2771;
assign w8532 = w1486 & ~w1554;
assign w8533 = w2406 & ~w77;
assign w8534 = w9323 & w5202;
assign w8535 = (w3727 & w10648) | (w3727 & w9294) | (w10648 & w9294);
assign w8536 = ~w1714 & ~w13569;
assign w8537 = w625 & w13003;
assign w8538 = ~w3914 & w8827;
assign w8539 = ~w7149 & w8883;
assign w8540 = ~w2387 & ~w9838;
assign w8541 = (~w4032 & w11914) | (~w4032 & w5910) | (w11914 & w5910);
assign w8542 = ~w1497 & w4480;
assign w8543 = (w13854 & w7782) | (w13854 & w215) | (w7782 & w215);
assign w8544 = w5301 & ~w13333;
assign w8545 = ~w12018 & w7733;
assign w8546 = ~w3877 & ~w485;
assign w8547 = w12271 & w3714;
assign w8548 = (w1190 & w3952) | (w1190 & w8415) | (w3952 & w8415);
assign w8549 = (~w9921 & ~w7630) | (~w9921 & w13957) | (~w7630 & w13957);
assign w8550 = w3435 & ~w14072;
assign w8551 = (~w6994 & ~w2445) | (~w6994 & w9733) | (~w2445 & w9733);
assign w8552 = w3671 & ~w3808;
assign w8553 = ~w11800 & w8325;
assign w8554 = ~w11783 & w2636;
assign w8555 = ~w10917 & w1387;
assign w8556 = w10653 & w790;
assign w8557 = w10676 & w894;
assign w8558 = (w1540 & w8503) | (w1540 & w10093) | (w8503 & w10093);
assign w8559 = ~w9810 & ~w13630;
assign w8560 = w6889 & w7423;
assign w8561 = w8253 & w2729;
assign w8562 = ~w11641 & ~w13782;
assign w8563 = ~w530 & ~w11421;
assign w8564 = w13594 & ~w1647;
assign w8565 = w6461 & w2125;
assign w8566 = w3288 & ~w3251;
assign w8567 = ~w2686 & w1174;
assign w8568 = (~w1190 & w12260) | (~w1190 & w12364) | (w12260 & w12364);
assign w8569 = ~w9226 & w10290;
assign w8570 = ~w10245 & w3580;
assign w8571 = (~w12569 & w14633) | (~w12569 & w6073) | (w14633 & w6073);
assign w8572 = w13399 & ~w6488;
assign w8573 = ~w2680 & w6301;
assign w8574 = ~w7764 & ~w4879;
assign w8575 = w9378 & w1287;
assign w8576 = w13774 & ~w10264;
assign w8577 = ~w7767 & w9753;
assign w8578 = w7513 & w1645;
assign w8579 = (w12460 & w2850) | (w12460 & w10916) | (w2850 & w10916);
assign w8580 = ~w12463 & ~w11213;
assign w8581 = w4042 & ~w12557;
assign w8582 = (~w3631 & w11790) | (~w3631 & w6331) | (w11790 & w6331);
assign w8583 = (w11097 & w12766) | (w11097 & w13190) | (w12766 & w13190);
assign w8584 = w5213 & w14215;
assign w8585 = (w4354 & w12878) | (w4354 & w9655) | (w12878 & w9655);
assign w8586 = w6700 & ~w2492;
assign w8587 = ~w12282 & w10170;
assign w8588 = w12609 & ~w14634;
assign w8589 = ~w10644 & w7293;
assign w8590 = (w13334 & w6457) | (w13334 & w7549) | (w6457 & w7549);
assign w8591 = (w9804 & ~w2709) | (w9804 & ~w12776) | (~w2709 & ~w12776);
assign w8592 = ~w142 & ~w1540;
assign w8593 = (w3128 & w13683) | (w3128 & ~w8861) | (w13683 & ~w8861);
assign w8594 = ~w607 & ~w8459;
assign w8595 = ~w1190 & w992;
assign w8596 = ~w5294 & w2680;
assign w8597 = (~w8067 & w8753) | (~w8067 & w8810) | (w8753 & w8810);
assign w8598 = ~w4753 & w148;
assign w8599 = (w9541 & w7224) | (w9541 & w5988) | (w7224 & w5988);
assign w8600 = w12112 & w2082;
assign w8601 = w4178 & w5446;
assign w8602 = w2320 & ~w1712;
assign w8603 = ~w10354 & ~w2227;
assign w8604 = w12460 & ~w7546;
assign w8605 = (w1968 & w6980) | (w1968 & w9607) | (w6980 & w9607);
assign w8606 = ~w243 & ~w11249;
assign w8607 = ~w12685 & ~w7362;
assign w8608 = ~w11338 & w12022;
assign w8609 = (~w14325 & w284) | (~w14325 & w1123) | (w284 & w1123);
assign w8610 = w6924 & w5405;
assign w8611 = w3215 & w14504;
assign w8612 = ~w217 & w11117;
assign w8613 = w14172 & w12587;
assign w8614 = (w14564 & w11756) | (w14564 & ~w4783) | (w11756 & ~w4783);
assign w8615 = ~w5522 & w3885;
assign w8616 = (~w3242 & w14159) | (~w3242 & w7312) | (w14159 & w7312);
assign w8617 = (~w9296 & w4134) | (~w9296 & w9618) | (w4134 & w9618);
assign w8618 = ~w12343 & ~w4105;
assign w8619 = ~w10517 & ~w9480;
assign w8620 = w10794 & ~w14127;
assign w8621 = ~w750 & w11352;
assign w8622 = w3963 & ~w7125;
assign w8623 = (~w14417 & ~w4511) | (~w14417 & ~w14564) | (~w4511 & ~w14564);
assign w8624 = ~w13503 & w8681;
assign w8625 = (w4855 & ~w5852) | (w4855 & w11365) | (~w5852 & w11365);
assign w8626 = ~w4359 & ~w473;
assign w8627 = (w2928 & w9564) | (w2928 & w9764) | (w9564 & w9764);
assign w8628 = w2569 & w3671;
assign w8629 = w1838 & ~w4458;
assign w8630 = (~w3958 & w13349) | (~w3958 & w2545) | (w13349 & w2545);
assign w8631 = w7902 & w8112;
assign w8632 = ~w5620 & ~w6949;
assign w8633 = (~w9012 & w11341) | (~w9012 & w13747) | (w11341 & w13747);
assign w8634 = w3373 & w12142;
assign w8635 = w12065 & ~w852;
assign w8636 = ~w5700 & ~w14580;
assign w8637 = (w6170 & w10129) | (w6170 & w2074) | (w10129 & w2074);
assign w8638 = (~w302 & w14330) | (~w302 & w5567) | (w14330 & w5567);
assign w8639 = (w10704 & w71) | (w10704 & w9492) | (w71 & w9492);
assign w8640 = (~w2941 & w6706) | (~w2941 & w5312) | (w6706 & w5312);
assign w8641 = (w12910 & w11912) | (w12910 & w10678) | (w11912 & w10678);
assign w8642 = w14629 & ~w9302;
assign w8643 = ~w12271 & w3661;
assign w8644 = ~w13462 & w10327;
assign w8645 = w13751 & ~w12460;
assign w8646 = w3911 & w9474;
assign w8647 = ~w14610 & ~w11052;
assign w8648 = (~w13854 & w3653) | (~w13854 & w1677) | (w3653 & w1677);
assign w8649 = ~w3997 & ~w2953;
assign w8650 = (~w595 & w1584) | (~w595 & w14329) | (w1584 & w14329);
assign w8651 = w10354 & w3727;
assign w8652 = (w12896 & w12027) | (w12896 & w8228) | (w12027 & w8228);
assign w8653 = w14335 & ~w7887;
assign w8654 = (~w3194 & w9250) | (~w3194 & w10453) | (w9250 & w10453);
assign w8655 = w2477 & ~w3912;
assign w8656 = w9748 & ~w3913;
assign w8657 = w3963 & w13635;
assign w8658 = ~w7488 & w4957;
assign w8659 = w11732 & w65;
assign w8660 = ~w563 & w12460;
assign w8661 = w4349 & ~w2004;
assign w8662 = ~w4700 & w4458;
assign w8663 = w4437 & w86;
assign w8664 = ~w4019 & w208;
assign w8665 = ~w3098 & w12656;
assign w8666 = (w10290 & ~w10659) | (w10290 & w742) | (~w10659 & w742);
assign w8667 = (w5574 & w1869) | (w5574 & w10991) | (w1869 & w10991);
assign w8668 = w10370 & w4328;
assign w8669 = w3649 & ~w4869;
assign w8670 = (w12988 & w13700) | (w12988 & w14455) | (w13700 & w14455);
assign w8671 = w12464 & w7906;
assign w8672 = w13290 & ~w9940;
assign w8673 = (w6598 & w5396) | (w6598 & w12376) | (w5396 & w12376);
assign w8674 = w12852 & w9332;
assign w8675 = ~w3951 & ~w8570;
assign w8676 = w10182 & ~w1474;
assign w8677 = (w12170 & w13462) | (w12170 & w13823) | (w13462 & w13823);
assign w8678 = (w13391 & w9103) | (w13391 & w2670) | (w9103 & w2670);
assign w8679 = w2752 & w3764;
assign w8680 = (~w4127 & w2492) | (~w4127 & w1403) | (w2492 & w1403);
assign w8681 = ~w12438 & w7135;
assign w8682 = ~w10610 & ~w9179;
assign w8683 = w11628 & w11248;
assign w8684 = (~w11185 & w11896) | (~w11185 & w12784) | (w11896 & w12784);
assign w8685 = w9463 & w12172;
assign w8686 = (~w11915 & w8846) | (~w11915 & w6608) | (w8846 & w6608);
assign w8687 = (~w11138 & w778) | (~w11138 & w9334) | (w778 & w9334);
assign w8688 = ~w13508 & w13323;
assign w8689 = ~w10358 & w6545;
assign w8690 = w7794 & w8039;
assign w8691 = ~b23 & ~a23;
assign w8692 = ~w1503 | w13331;
assign w8693 = w3759 & ~w4515;
assign w8694 = ~w1503 & ~w372;
assign w8695 = (w14528 & w2119) | (w14528 & w2087) | (w2119 & w2087);
assign w8696 = (w9536 & w11252) | (w9536 & w8050) | (w11252 & w8050);
assign w8697 = (w7784 & w12076) | (w7784 & w11842) | (w12076 & w11842);
assign w8698 = ~w8773 & w12084;
assign w8699 = w5543 & w6230;
assign w8700 = (w2166 & w1259) | (w2166 & w11683) | (w1259 & w11683);
assign w8701 = ~w12271 & ~w11732;
assign w8702 = w13692 & ~w8969;
assign w8703 = (w6657 & w12004) | (w6657 & w2254) | (w12004 & w2254);
assign w8704 = ~w4050 & w7920;
assign w8705 = ~w13541 & ~w3769;
assign w8706 = ~w11261 & w10312;
assign w8707 = w10423 & ~w3906;
assign w8708 = ~w1165 & ~w459;
assign w8709 = w14417 & ~w12493;
assign w8710 = (~w7026 & w1120) | (~w7026 & w584) | (w1120 & w584);
assign w8711 = ~w3611 & ~w14504;
assign w8712 = w8894 & w3564;
assign w8713 = w4078 & w7633;
assign w8714 = (w9096 & w5861) | (w9096 & w10887) | (w5861 & w10887);
assign w8715 = (~w6758 & w2627) | (~w6758 & w9267) | (w2627 & w9267);
assign w8716 = (w6281 & ~w7085) | (w6281 & w10284) | (~w7085 & w10284);
assign w8717 = ~w9494 & ~w4907;
assign w8718 = (w5243 & w7936) | (w5243 & w14227) | (w7936 & w14227);
assign w8719 = ~w706 & ~w1802;
assign w8720 = ~w12972 & w5015;
assign w8721 = (w6832 & w3476) | (w6832 & w4091) | (w3476 & w4091);
assign w8722 = ~w5177 & w3025;
assign w8723 = (~w3885 & w4377) | (~w3885 & w6879) | (w4377 & w6879);
assign w8724 = ~w7746 & ~b93;
assign w8725 = w7896 & w13152;
assign w8726 = w9461 & w1209;
assign w8727 = ~w2433 & ~w10032;
assign w8728 = ~w12371 & ~w9788;
assign w8729 = ~w2942 & ~w11101;
assign w8730 = (w4692 & w6634) | (w4692 & ~w11756) | (w6634 & ~w11756);
assign w8731 = (w2272 & w12646) | (w2272 & w6310) | (w12646 & w6310);
assign w8732 = ~w142 & ~w9211;
assign w8733 = ~w13183 & w5743;
assign w8734 = ~w4032 & w5482;
assign w8735 = ~w1812 & w3078;
assign w8736 = ~w14437 & ~w13618;
assign w8737 = ~w9871 & ~w9817;
assign w8738 = (~w4363 & w13355) | (~w4363 & w12127) | (w13355 & w12127);
assign w8739 = w10045 & w10357;
assign w8740 = (~w10408 & w6406) | (~w10408 & w14636) | (w6406 & w14636);
assign w8741 = ~w2284 & w6090;
assign w8742 = ~w6699 & ~w12893;
assign w8743 = w8589 & w11321;
assign w8744 = w4322 & ~w6689;
assign w8745 = w3852 & w4835;
assign w8746 = ~w1742 & ~w2258;
assign w8747 = (w4386 & w14059) | (w4386 & w5159) | (w14059 & w5159);
assign w8748 = w10517 & ~w2729;
assign w8749 = ~w5562 & w737;
assign w8750 = ~w11375 & ~w1905;
assign w8751 = w13854 & ~w9486;
assign w8752 = w10014 & w2273;
assign w8753 = ~w8396 & ~w7104;
assign w8754 = ~b86 & ~a86;
assign w8755 = w11680 & ~w12045;
assign w8756 = (w1849 & w6056) | (w1849 & w677) | (w6056 & w677);
assign w8757 = ~w12464 & ~w7190;
assign w8758 = ~w10517 & ~w13730;
assign w8759 = w5178 & w8389;
assign w8760 = w10107 & ~w12276;
assign w8761 = w10700 & w472;
assign w8762 = (~w8614 & w5625) | (~w8614 & w10921) | (w5625 & w10921);
assign w8763 = w2583 & ~w9711;
assign w8764 = (w11925 & w1973) | (w11925 & w3468) | (w1973 & w3468);
assign w8765 = ~w14028 & ~w1829;
assign w8766 = ~w2317 & w6846;
assign w8767 = w3721 & ~w10023;
assign w8768 = ~b28 & ~a28;
assign w8769 = ~w12497 & ~w8366;
assign w8770 = (w1871 & w13310) | (w1871 & w749) | (w13310 & w749);
assign w8771 = w14624 & w4664;
assign w8772 = (w6464 & ~w3129) | (w6464 & w1716) | (~w3129 & w1716);
assign w8773 = w6391 & w3532;
assign w8774 = ~w142 & ~w10699;
assign w8775 = (~w3612 & w204) | (~w3612 & w2276) | (w204 & w2276);
assign w8776 = w5522 & ~w3727;
assign w8777 = w9212 & w11976;
assign w8778 = ~w9374 & w8350;
assign w8779 = w5178 & w4233;
assign w8780 = w423 & ~w5777;
assign w8781 = (w8937 & w11822) | (w8937 & w7407) | (w11822 & w7407);
assign w8782 = b126 & a126;
assign w8783 = ~w8937 & w10753;
assign w8784 = w11137 & w793;
assign w8785 = (~w7754 & w12095) | (~w7754 & w9357) | (w12095 & w9357);
assign w8786 = ~w2202 & ~w11606;
assign w8787 = ~w9550 & w10818;
assign w8788 = (~w8328 & ~w12460) | (~w8328 & w10507) | (~w12460 & w10507);
assign w8789 = (w4030 & w10726) | (w4030 & w1921) | (w10726 & w1921);
assign w8790 = w11899 & ~w12388;
assign w8791 = w3550 & w10895;
assign w8792 = w14246 & w6054;
assign w8793 = (w8047 & w10247) | (w8047 & w12211) | (w10247 & w12211);
assign w8794 = (~w4545 & w12075) | (~w4545 & w4919) | (w12075 & w4919);
assign w8795 = ~w14510 & ~w11920;
assign w8796 = (~w844 & w10109) | (~w844 & w11144) | (w10109 & w11144);
assign w8797 = w3627 & w8717;
assign w8798 = (w3721 & w14665) | (w3721 & w5637) | (w14665 & w5637);
assign w8799 = (w14648 & w2442) | (w14648 & w9856) | (w2442 & w9856);
assign w8800 = ~w922 & w3036;
assign w8801 = w5294 & w12943;
assign w8802 = w2188 & ~w4273;
assign w8803 = w12569 & ~w9921;
assign w8804 = (w12332 & w3464) | (w12332 & w1484) | (w3464 & w1484);
assign w8805 = (w2858 & w2567) | (w2858 & w309) | (w2567 & w309);
assign w8806 = ~w13713 & ~w11372;
assign w8807 = (~w1362 & w10226) | (~w1362 & w3000) | (w10226 & w3000);
assign w8808 = ~w5737 & w10132;
assign w8809 = w4881 & w11031;
assign w8810 = ~w8396 & w10137;
assign w8811 = ~w12216 & ~w2941;
assign w8812 = w9032 & w11910;
assign w8813 = ~w9190 & w2193;
assign w8814 = w8080 & ~w318;
assign w8815 = ~w7717 & ~w8176;
assign w8816 = ~w12663 & ~w6905;
assign w8817 = ~w4263 & w11445;
assign w8818 = ~w8140 & ~w8885;
assign w8819 = ~w8280 & ~w6668;
assign w8820 = (w6572 & w2492) | (w6572 & w8173) | (w2492 & w8173);
assign w8821 = ~w5231 & w6970;
assign w8822 = (~w10023 & w4432) | (~w10023 & w2181) | (w4432 & w2181);
assign w8823 = ~w12553 & ~w11732;
assign w8824 = w8044 & w889;
assign w8825 = (~w3387 & ~w13654) | (~w3387 & w13758) | (~w13654 & w13758);
assign w8826 = w10290 & w11365;
assign w8827 = ~b62 & ~a62;
assign w8828 = (~w9694 & ~w1140) | (~w9694 & w7532) | (~w1140 & w7532);
assign w8829 = w5864 & ~w6907;
assign w8830 = w7159 & ~w7161;
assign w8831 = ~w14202 & ~w3806;
assign w8832 = ~w6676 & w2727;
assign w8833 = ~w4830 & ~w6129;
assign w8834 = w3823 & ~w5059;
assign w8835 = ~w2431 & w2236;
assign w8836 = ~w2500 & w1816;
assign w8837 = ~w254 & w4400;
assign w8838 = ~w13282 & w14380;
assign w8839 = (w12170 & w10245) | (w12170 & w6007) | (w10245 & w6007);
assign w8840 = w4627 & ~w5664;
assign w8841 = w1096 & ~w10483;
assign w8842 = w7001 & w13323;
assign w8843 = w4787 & w664;
assign w8844 = ~w1839 & w1884;
assign w8845 = ~w11429 & w5326;
assign w8846 = w5794 | w2600;
assign w8847 = w11683 & ~w10192;
assign w8848 = (w1938 & w8652) | (w1938 & ~w2670) | (w8652 & ~w2670);
assign w8849 = (w5105 & w815) | (w5105 & w6959) | (w815 & w6959);
assign w8850 = ~w9608 & w6465;
assign w8851 = ~w6241 & w13173;
assign w8852 = w10477 & ~w11488;
assign w8853 = ~w5852 & ~w10119;
assign w8854 = ~w1579 & w862;
assign w8855 = w5348 & w4231;
assign w8856 = w1821 & w12311;
assign w8857 = w7886 & ~w7026;
assign w8858 = w10910 & ~w4513;
assign w8859 = (w5593 & w3642) | (w5593 & w395) | (w3642 & w395);
assign w8860 = w5574 & ~w1805;
assign w8861 = w541 & w1464;
assign w8862 = w4655 & w14389;
assign w8863 = w5761 & ~w1474;
assign w8864 = (w9316 & w11737) | (w9316 & w1265) | (w11737 & w1265);
assign w8865 = (~w6342 & w7436) | (~w6342 & w1131) | (w7436 & w1131);
assign w8866 = ~w1785 & w11257;
assign w8867 = w14207 & w2214;
assign w8868 = w12614 & ~w5002;
assign w8869 = ~w2656 & w11488;
assign w8870 = (~w8896 & w6114) | (~w8896 & w7750) | (w6114 & w7750);
assign w8871 = (~w8280 & w5842) | (~w8280 & w4488) | (w5842 & w4488);
assign w8872 = ~w11005 & ~w3139;
assign w8873 = ~w9015 & ~w77;
assign w8874 = (~w6984 & w2831) | (~w6984 & w13601) | (w2831 & w13601);
assign w8875 = ~w13302 & w8396;
assign w8876 = (~w922 & w3775) | (~w922 & w9938) | (w3775 & w9938);
assign w8877 = ~w9805 & w2486;
assign w8878 = w13197 & w3788;
assign w8879 = w12958 & ~w3036;
assign w8880 = w9349 & ~w10486;
assign w8881 = ~w13282 & w309;
assign w8882 = w2096 & w10182;
assign w8883 = ~w3089 & w6138;
assign w8884 = (~w846 & w6940) | (~w846 & w14374) | (w6940 & w14374);
assign w8885 = ~w6426 & w8373;
assign w8886 = ~w14072 & w13694;
assign w8887 = w13566 & w14497;
assign w8888 = w10959 & w9952;
assign w8889 = (w1878 & w11994) | (w1878 & w1823) | (w11994 & w1823);
assign w8890 = w13190 & w1553;
assign w8891 = w4076 & w14193;
assign w8892 = (~w4511 & w8555) | (~w4511 & w65) | (w8555 & w65);
assign w8893 = w9583 & w13628;
assign w8894 = ~w9715 & w10075;
assign w8895 = w8253 & w4458;
assign w8896 = (~w11606 & w9798) | (~w11606 & w10573) | (w9798 & w10573);
assign w8897 = ~w8700 & w10914;
assign w8898 = ~w14340 & ~w13077;
assign w8899 = ~w14639 & ~w278;
assign w8900 = (~w12121 & w9487) | (~w12121 & w8395) | (w9487 & w8395);
assign w8901 = ~w7344 & w97;
assign w8902 = w12460 & ~w954;
assign w8903 = (w14543 & w12345) | (w14543 & w7654) | (w12345 & w7654);
assign w8904 = ~w4425 & ~w9454;
assign w8905 = w13533 & w11574;
assign w8906 = (~w2984 & ~w1806) | (~w2984 & w4699) | (~w1806 & w4699);
assign w8907 = ~w4512 & w1017;
assign w8908 = w7069 & ~w4293;
assign w8909 = ~w364 & ~w7951;
assign w8910 = (w8512 & w14661) | (w8512 & ~w3564) | (w14661 & ~w3564);
assign w8911 = ~w13947 & ~w6271;
assign w8912 = w4253 & w374;
assign w8913 = w11508 & w14671;
assign w8914 = ~w8941 & w2330;
assign w8915 = w10467 & w8584;
assign w8916 = (~w4607 & w1218) | (~w4607 & w7520) | (w1218 & w7520);
assign w8917 = ~w4158 & w13002;
assign w8918 = w852 & w5845;
assign w8919 = w6275 & ~w7768;
assign w8920 = w4704 & w4928;
assign w8921 = ~w12575 & w9655;
assign w8922 = (~w9688 & ~w14174) | (~w9688 & w6256) | (~w14174 & w6256);
assign w8923 = (w10477 & w11261) | (w10477 & w9143) | (w11261 & w9143);
assign w8924 = ~w9259 & ~w11960;
assign w8925 = w6406 & ~w12642;
assign w8926 = w9472 & w11968;
assign w8927 = (w13331 & w11337) | (w13331 & w2898) | (w11337 & w2898);
assign w8928 = (w12914 & w7423) | (w12914 & w7388) | (w7423 & w7388);
assign w8929 = w8691 & ~w6433;
assign w8930 = w2602 & ~w8024;
assign w8931 = w159 & w3097;
assign w8932 = w10877 & w1378;
assign w8933 = (w1760 & ~w12808) | (w1760 & w4024) | (~w12808 & w4024);
assign w8934 = w10032 & w8396;
assign w8935 = (w7272 & w5995) | (w7272 & w6355) | (w5995 & w6355);
assign w8936 = (~w3158 & w13587) | (~w3158 & w8043) | (w13587 & w8043);
assign w8937 = w8817 & ~w14068;
assign w8938 = ~w4607 & w5199;
assign w8939 = (w12614 & w4586) | (w12614 & w12233) | (w4586 & w12233);
assign w8940 = w13148 & ~w9266;
assign w8941 = ~w11934 & w14172;
assign w8942 = ~w6135 & ~w8396;
assign w8943 = ~w4824 & ~w4951;
assign w8944 = ~w8279 & ~w14425;
assign w8945 = (~w5556 & w4050) | (~w5556 & w2453) | (w4050 & w2453);
assign w8946 = w4515 & ~w11117;
assign w8947 = w11757 & ~w2701;
assign w8948 = w10036 & w6299;
assign w8949 = ~w14335 & w7042;
assign w8950 = ~w13874 & w8411;
assign w8951 = w474 & w9653;
assign w8952 = ~w569 & w2012;
assign w8953 = w1140 & w2158;
assign w8954 = w13199 | w7914;
assign w8955 = (~w6929 & w3672) | (~w6929 & w1615) | (w3672 & w1615);
assign w8956 = ~w4521 & ~w1531;
assign w8957 = w12575 & w852;
assign w8958 = ~w3209 & w14659;
assign w8959 = (w5660 & w1785) | (w5660 & w3888) | (w1785 & w3888);
assign w8960 = ~w2175 & w4910;
assign w8961 = w9268 & ~w9543;
assign w8962 = w6889 & w9748;
assign w8963 = ~w11069 & w978;
assign w8964 = ~w4032 & ~w2144;
assign w8965 = ~w4989 & w8331;
assign w8966 = ~w5282 & w4431;
assign w8967 = ~w3508 & ~w499;
assign w8968 = (~w4127 & w183) | (~w4127 & w4423) | (w183 & w4423);
assign w8969 = ~w14395 & w8346;
assign w8970 = (~w10483 & w4324) | (~w10483 & w9931) | (w4324 & w9931);
assign w8971 = ~w1474 & w13323;
assign w8972 = w3885 & w6500;
assign w8973 = ~w7768 & ~w14130;
assign w8974 = w9453 & ~w12893;
assign w8975 = w7914 & w7376;
assign w8976 = w11579 & ~w6290;
assign w8977 = w12438 & w1699;
assign w8978 = (~w13462 & w3817) | (~w13462 & w2103) | (w3817 & w2103);
assign w8979 = (~w5161 & w8012) | (~w5161 & w6050) | (w8012 & w6050);
assign w8980 = w5867 & w8827;
assign w8981 = w8705 & w5400;
assign w8982 = ~w1172 & ~w5247;
assign w8983 = (w2 & w977) | (w2 & w8238) | (w977 & w8238);
assign w8984 = (w13562 & w2368) | (w13562 & w8509) | (w2368 & w8509);
assign w8985 = w10941 & w5761;
assign w8986 = (w9300 & ~w4557) | (w9300 & w13727) | (~w4557 & w13727);
assign w8987 = ~w608 & ~w6381;
assign w8988 = w5612 & ~w1709;
assign w8989 = (~w3325 & w11261) | (~w3325 & w13176) | (w11261 & w13176);
assign w8990 = w2320 & ~w6845;
assign w8991 = ~w3779 & ~w814;
assign w8992 = ~w1991 & ~w3970;
assign w8993 = ~w13902 & ~w9896;
assign w8994 = w1140 & w2776;
assign w8995 = w12553 & w3502;
assign w8996 = ~w13907 & ~w13555;
assign w8997 = w10566 & ~w8784;
assign w8998 = (w6822 & w11873) | (w6822 & w8198) | (w11873 & w8198);
assign w8999 = ~w536 & ~w10477;
assign w9000 = ~w3067 & w8264;
assign w9001 = ~w8171 & w8513;
assign w9002 = ~w6732 & w10883;
assign w9003 = (~w1260 & w3385) | (~w1260 & ~w2159) | (w3385 & ~w2159);
assign w9004 = (~w11395 & w14430) | (~w11395 & w8139) | (w14430 & w8139);
assign w9005 = w13282 & w829;
assign w9006 = w3325 & w10225;
assign w9007 = (~w4044 & w1198) | (~w4044 & w6182) | (w1198 & w6182);
assign w9008 = (w3615 & w8499) | (w3615 & w11615) | (w8499 & w11615);
assign w9009 = (~w11750 & w3841) | (~w11750 & w1889) | (w3841 & w1889);
assign w9010 = ~w13010 & w11732;
assign w9011 = w13780 & ~a53;
assign w9012 = w12472 & ~w9593;
assign w9013 = (w2236 & w12980) | (w2236 & w8835) | (w12980 & w8835);
assign w9014 = ~w2701 & w8280;
assign w9015 = ~b66 & ~a66;
assign w9016 = ~w2807 & ~w8991;
assign w9017 = ~w2656 & w6572;
assign w9018 = w3383 & w318;
assign w9019 = ~w12271 & w11395;
assign w9020 = ~w575 & ~w10007;
assign w9021 = ~w9465 & ~w9183;
assign w9022 = ~w13321 & w367;
assign w9023 = (~w308 & w4946) | (~w308 & w9824) | (w4946 & w9824);
assign w9024 = w13839 & ~w5338;
assign w9025 = ~w5021 & ~w2755;
assign w9026 = w9846 & ~w3963;
assign w9027 = (w13331 & w9520) | (w13331 & w3052) | (w9520 & w3052);
assign w9028 = (w339 & w10521) | (w339 & ~w4232) | (w10521 & ~w4232);
assign w9029 = w14185 & w2120;
assign w9030 = (w8697 & w12687) | (w8697 & w8255) | (w12687 & w8255);
assign w9031 = w5522 & w10182;
assign w9032 = w7455 & w14280;
assign w9033 = (w717 & w14096) | (w717 & ~w12376) | (w14096 & ~w12376);
assign w9034 = w1171 & ~w14140;
assign w9035 = ~w2799 & ~w12169;
assign w9036 = w2567 | w2858;
assign w9037 = w6343 & w5411;
assign w9038 = (~w4099 & w3829) | (~w4099 & w10362) | (w3829 & w10362);
assign w9039 = w4204 & ~w11915;
assign w9040 = ~w5860 & ~w10224;
assign w9041 = ~w1899 & ~w6655;
assign w9042 = (w5865 & ~w922) | (w5865 & w3187) | (~w922 & w3187);
assign w9043 = (w7082 & w5323) | (w7082 & w13962) | (w5323 & w13962);
assign w9044 = ~w3914 & w12065;
assign w9045 = (~w10423 & w12980) | (~w10423 & w561) | (w12980 & w561);
assign w9046 = ~w6442 & w3852;
assign w9047 = ~w5635 & ~w3427;
assign w9048 = (w8827 & w4158) | (w8827 & w2846) | (w4158 & w2846);
assign w9049 = w7006 & w5788;
assign w9050 = w3435 & ~w4473;
assign w9051 = ~w3790 & w9672;
assign w9052 = w9183 & w142;
assign w9053 = (~w5219 & w12124) | (~w5219 & w4077) | (w12124 & w4077);
assign w9054 = ~w13198 & w8641;
assign w9055 = ~w11462 & w3242;
assign w9056 = (w4127 & w2656) | (w4127 & w7877) | (w2656 & w7877);
assign w9057 = ~w10182 & w6145;
assign w9058 = w13156 & w6525;
assign w9059 = ~w580 & ~w13788;
assign w9060 = ~w9715 & ~w5301;
assign w9061 = (~w5783 & w5773) | (~w5783 & w5054) | (w5773 & w5054);
assign w9062 = (~w2680 & w2144) | (~w2680 & w2350) | (w2144 & w2350);
assign w9063 = w796 & w10259;
assign w9064 = w9183 & ~w4359;
assign w9065 = ~w7031 & ~w5939;
assign w9066 = ~w1878 & ~w1683;
assign w9067 = (w4894 & ~w5055) | (w4894 & w32) | (~w5055 & w32);
assign w9068 = ~w10594 & ~w12830;
assign w9069 = ~w8778 & w3986;
assign w9070 = w9672 & w4541;
assign w9071 = w6542 & ~w7962;
assign w9072 = w3209 & w6683;
assign w9073 = (w6637 & w2528) | (w6637 & w4594) | (w2528 & w4594);
assign w9074 = w3872 & w8037;
assign w9075 = ~w12556 & ~w8102;
assign w9076 = (~w1362 & w6110) | (~w1362 & w2744) | (w6110 & w2744);
assign w9077 = w9455 & w11758;
assign w9078 = w8459 & ~w1200;
assign w9079 = (w217 & ~w11138) | (w217 & w6589) | (~w11138 & w6589);
assign w9080 = (~w1712 & w9868) | (~w1712 & w1327) | (w9868 & w1327);
assign w9081 = w9776 & w12589;
assign w9082 = (w2595 & w5476) | (w2595 & ~w13980) | (w5476 & ~w13980);
assign w9083 = (w11634 & w7456) | (w11634 & w14080) | (w7456 & w14080);
assign w9084 = (w12915 & w9784) | (w12915 & ~w2170) | (w9784 & ~w2170);
assign w9085 = w8035 & w10483;
assign w9086 = ~w7373 & ~w1906;
assign w9087 = ~w2410 & ~w9453;
assign w9088 = ~w4375 & ~w14659;
assign w9089 = w3209 & ~w1442;
assign w9090 = w12604 & ~w6135;
assign w9091 = (w5845 & w8918) | (w5845 & w8820) | (w8918 & w8820);
assign w9092 = ~w687 & ~w12034;
assign w9093 = (w2698 & w4395) | (w2698 & w8706) | (w4395 & w8706);
assign w9094 = w9842 & w6719;
assign w9095 = ~w8827 & ~w14660;
assign w9096 = (w12889 & w5991) | (w12889 & w4709) | (w5991 & w4709);
assign w9097 = ~w7001 & w5761;
assign w9098 = (w13360 & w7726) | (w13360 & w55) | (w7726 & w55);
assign w9099 = w7198 & w396;
assign w9100 = ~w4587 & ~w4425;
assign w9101 = ~w11218 & w8900;
assign w9102 = w7740 & w8273;
assign w9103 = (~w13633 & w11426) | (~w13633 & ~w8228) | (w11426 & ~w8228);
assign w9104 = (~w254 & w9238) | (~w254 & w10088) | (w9238 & w10088);
assign w9105 = w9904 & w10708;
assign w9106 = ~w3759 & w12685;
assign w9107 = ~w254 & w4922;
assign w9108 = ~w494 & w8942;
assign w9109 = w813 & w10925;
assign w9110 = (w6845 & w2967) | (w6845 & w13322) | (w2967 & w13322);
assign w9111 = ~w12121 & w7588;
assign w9112 = (w1770 & w8235) | (w1770 & w11037) | (w8235 & w11037);
assign w9113 = (~w3325 & w10928) | (~w3325 & w12553) | (w10928 & w12553);
assign w9114 = (~w1260 & w3385) | (~w1260 & ~w8342) | (w3385 & ~w8342);
assign w9115 = ~w142 & ~w11861;
assign w9116 = (~w14513 & ~w8368) | (~w14513 & w511) | (~w8368 & w511);
assign w9117 = ~w12148 & w6310;
assign w9118 = ~w993 & ~w11829;
assign w9119 = (~w8772 & w1425) | (~w8772 & w1161) | (w1425 & w1161);
assign w9120 = ~w11345 & w14054;
assign w9121 = w5741 & ~w9623;
assign w9122 = ~w12604 & ~w3727;
assign w9123 = ~w10692 & ~w2584;
assign w9124 = (~w1037 & w12953) | (~w1037 & w4365) | (w12953 & w4365);
assign w9125 = ~w9912 & ~w12816;
assign w9126 = (w1768 & w1571) | (w1768 & w4120) | (w1571 & w4120);
assign w9127 = (w10855 & w11433) | (w10855 & w12913) | (w11433 & w12913);
assign w9128 = ~w6752 & ~w3941;
assign w9129 = (~w11173 & w10662) | (~w11173 & w12733) | (w10662 & w12733);
assign w9130 = w8106 & w4787;
assign w9131 = (w869 & w8714) | (w869 & ~w8228) | (w8714 & ~w8228);
assign w9132 = (w6423 & w10329) | (w6423 & w3739) | (w10329 & w3739);
assign w9133 = ~w14552 & w14258;
assign w9134 = (w4658 & ~w5121) | (w4658 & w3415) | (~w5121 & w3415);
assign w9135 = w5294 & w12170;
assign w9136 = (w7690 & w4121) | (w7690 & w7394) | (w4121 & w7394);
assign w9137 = w11909 & w4541;
assign w9138 = ~w2675 & ~w4071;
assign w9139 = ~w4105 & ~w5785;
assign w9140 = w10072 & ~w10079;
assign w9141 = w10032 & w10699;
assign w9142 = w12065 & w3039;
assign w9143 = w8234 & w10477;
assign w9144 = w759 & w7680;
assign w9145 = ~b22 & ~a22;
assign w9146 = w13376 & w7351;
assign w9147 = ~w2095 & w2174;
assign w9148 = w7347 & w3517;
assign w9149 = w2762 & w3427;
assign w9150 = ~w1802 & w8019;
assign w9151 = (w9126 & w5381) | (w9126 & w12657) | (w5381 & w12657);
assign w9152 = (w7664 & w6071) | (w7664 & w11939) | (w6071 & w11939);
assign w9153 = ~w7804 & w4602;
assign w9154 = (w11734 & w10069) | (w11734 & w6347) | (w10069 & w6347);
assign w9155 = w560 & w1235;
assign w9156 = (~w13713 & w12112) | (~w13713 & w7249) | (w12112 & w7249);
assign w9157 = w7794 & w9410;
assign w9158 = ~w3216 & ~w14168;
assign w9159 = ~w2159 & w13838;
assign w9160 = ~w12749 & ~w6440;
assign w9161 = ~w11333 & w2492;
assign w9162 = ~w3243 & ~w6742;
assign w9163 = w2485 & ~w13342;
assign w9164 = w4836 & w3501;
assign w9165 = ~w8752 & w5061;
assign w9166 = ~w7867 & ~w98;
assign w9167 = ~w9608 & w6604;
assign w9168 = (~w1586 & w9887) | (~w1586 & w4767) | (w9887 & w4767);
assign w9169 = w7709 | ~w5385;
assign w9170 = w13694 & w1699;
assign w9171 = (w13654 & w38) | (w13654 & w6791) | (w38 & w6791);
assign w9172 = ~w8698 & w10090;
assign w9173 = ~w5294 & w3508;
assign w9174 = ~w5691 & ~w6225;
assign w9175 = w6218 & w3888;
assign w9176 = ~w1918 & w4060;
assign w9177 = w4836 & w8390;
assign w9178 = w1986 & ~w7160;
assign w9179 = ~w7488 & w2550;
assign w9180 = ~w4865 & ~w7670;
assign w9181 = ~w2320 & ~w11855;
assign w9182 = (~w3937 & w3765) | (~w3937 & w7779) | (w3765 & w7779);
assign w9183 = ~w4312 & ~w6281;
assign w9184 = (w13552 & w11369) | (w13552 & w9274) | (w11369 & w9274);
assign w9185 = w13356 & w797;
assign w9186 = (~w1949 & w5294) | (~w1949 & w13075) | (w5294 & w13075);
assign w9187 = ~w1048 & w13243;
assign w9188 = ~w12228 & ~w13860;
assign w9189 = ~w3790 & ~w4026;
assign w9190 = ~w7172 & ~w6194;
assign w9191 = ~w7630 & w11533;
assign w9192 = ~w10075 & ~w11551;
assign w9193 = w1208 | w14059;
assign w9194 = (w9748 & w10364) | (w9748 & w9629) | (w10364 & w9629);
assign w9195 = w2954 & w6258;
assign w9196 = (~w10200 & w2136) | (~w10200 & w13858) | (w2136 & w13858);
assign w9197 = (~w5948 & ~w3285) | (~w5948 & w11432) | (~w3285 & w11432);
assign w9198 = ~w1257 & w2760;
assign w9199 = (~w12992 & w7026) | (~w12992 & w5315) | (w7026 & w5315);
assign w9200 = ~w8754 & ~w13214;
assign w9201 = ~w12924 & ~w6640;
assign w9202 = ~w9855 & ~w3904;
assign w9203 = (~w8279 & w6918) | (~w8279 & w473) | (w6918 & w473);
assign w9204 = ~w10180 & ~w3963;
assign w9205 = w6518 & ~w4420;
assign w9206 = (~w12807 & w11078) | (~w12807 & w10552) | (w11078 & w10552);
assign w9207 = (w8149 & w2993) | (w8149 & w6674) | (w2993 & w6674);
assign w9208 = ~w2787 & w6269;
assign w9209 = (w2144 & w11131) | (w2144 & w7918) | (w11131 & w7918);
assign w9210 = ~w2705 & w14651;
assign w9211 = ~w10941 & ~w6080;
assign w9212 = w4203 & w1729;
assign w9213 = (w5110 & w5235) | (w5110 & w9797) | (w5235 & w9797);
assign w9214 = w10437 & w1936;
assign w9215 = (w5744 & w13172) | (w5744 & w4339) | (w13172 & w4339);
assign w9216 = (w11350 & w4099) | (w11350 & w12584) | (w4099 & w12584);
assign w9217 = (w8873 & ~w11732) | (w8873 & w995) | (~w11732 & w995);
assign w9218 = w830 & w1651;
assign w9219 = ~w13854 & w1809;
assign w9220 = w1114 & w10036;
assign w9221 = w5422 & ~w4044;
assign w9222 = ~w12553 & ~w598;
assign w9223 = (~w52 & w14657) | (~w52 & w8751) | (w14657 & w8751);
assign w9224 = ~w2045 & ~w4235;
assign w9225 = ~w4751 & ~w5547;
assign w9226 = ~b58 & ~a58;
assign w9227 = ~w3502 & ~w3025;
assign w9228 = w2492 & ~w5919;
assign w9229 = w1773 & w10565;
assign w9230 = w8294 & w799;
assign w9231 = (w3671 & w4643) | (w3671 & w3308) | (w4643 & w3308);
assign w9232 = (w13613 & w6075) | (w13613 & w8487) | (w6075 & w8487);
assign w9233 = w9211 & w3291;
assign w9234 = (w10832 & w8627) | (w10832 & ~w4754) | (w8627 & ~w4754);
assign w9235 = (~w12816 & ~w7299) | (~w12816 & w9125) | (~w7299 & w9125);
assign w9236 = (~w2144 & w9921) | (~w2144 & w7866) | (w9921 & w7866);
assign w9237 = ~w2864 & ~w8459;
assign w9238 = ~w9921 & ~w829;
assign w9239 = (w8230 & w4093) | (w8230 & w768) | (w4093 & w768);
assign w9240 = ~w12121 & w7811;
assign w9241 = ~w7636 & ~w3121;
assign w9242 = ~w9256 & ~w10354;
assign w9243 = ~w3067 & w12526;
assign w9244 = b82 & a82;
assign w9245 = (w13452 & w983) | (w13452 & w12455) | (w983 & w12455);
assign w9246 = ~w6113 & ~w9290;
assign w9247 = (~w1518 & w3857) | (~w1518 & w5902) | (w3857 & w5902);
assign w9248 = ~w14024 & w682;
assign w9249 = w11733 & w4502;
assign w9250 = w5761 & ~w12421;
assign w9251 = w9461 & w5408;
assign w9252 = w12545 & ~w4223;
assign w9253 = ~w14664 & ~w8279;
assign w9254 = w2281 & w1902;
assign w9255 = w1842 & w3447;
assign w9256 = b122 & a122;
assign w9257 = w2656 & ~w6949;
assign w9258 = w7084 & w11918;
assign w9259 = ~w2627 & ~w6120;
assign w9260 = ~w11700 & ~w11245;
assign w9261 = ~w1873 & w2663;
assign w9262 = (~w9623 & w4134) | (~w9623 & w9121) | (w4134 & w9121);
assign w9263 = w7447 & ~w4515;
assign w9264 = w5732 & w12135;
assign w9265 = w10880 & w13628;
assign w9266 = (w4989 & w6242) | (w4989 & w2537) | (w6242 & w2537);
assign w9267 = w6120 & ~w6758;
assign w9268 = (w4395 & w13617) | (w4395 & w12600) | (w13617 & w12600);
assign w9269 = (w12101 & ~w12156) | (w12101 & w14039) | (~w12156 & w14039);
assign w9270 = (w12614 & w9737) | (w12614 & w10976) | (w9737 & w10976);
assign w9271 = (w8786 & w11650) | (w8786 & w10318) | (w11650 & w10318);
assign w9272 = (w4987 & w9735) | (w4987 & w9098) | (w9735 & w9098);
assign w9273 = ~w8328 & ~w577;
assign w9274 = ~w3331 & w13552;
assign w9275 = ~w14033 & w8019;
assign w9276 = w11759 & ~w8659;
assign w9277 = ~w4780 & w3602;
assign w9278 = w4114 & ~w12374;
assign w9279 = w4503 & w9707;
assign w9280 = w10032 & ~w4111;
assign w9281 = (~w7623 & w2161) | (~w7623 & w6547) | (w2161 & w6547);
assign w9282 = w14302 & w10317;
assign w9283 = ~w5522 & ~w12371;
assign w9284 = ~w1474 & ~w10221;
assign w9285 = w7519 | ~w2951;
assign w9286 = ~w12893 & w3611;
assign w9287 = w12545 & ~w3075;
assign w9288 = ~w13659 & ~w10606;
assign w9289 = w9170 & w12060;
assign w9290 = w6716 & w13620;
assign w9291 = w7365 & ~w3219;
assign w9292 = ~w7508 & w5118;
assign w9293 = w7127 & w4442;
assign w9294 = w6391 & w5033;
assign w9295 = w9997 & w9989;
assign w9296 = ~w10517 & ~w14015;
assign w9297 = w2701 & w3251;
assign w9298 = ~w13423 & w4399;
assign w9299 = w2656 & ~w8080;
assign w9300 = w6566 & w8504;
assign w9301 = w12893 & w347;
assign w9302 = w14054 & ~w11117;
assign w9303 = ~w14578 & w1939;
assign w9304 = ~w9233 & ~w1005;
assign w9305 = (w2655 & w2287) | (w2655 & w996) | (w2287 & w996);
assign w9306 = ~w6144 & w14663;
assign w9307 = w142 & w803;
assign w9308 = ~w7317 & w6651;
assign w9309 = w8657 & ~w13876;
assign w9310 = ~cin & w10992;
assign w9311 = (w6364 & w2313) | (w6364 & w9790) | (w2313 & w9790);
assign w9312 = ~w1785 & w7059;
assign w9313 = ~w8226 & w14352;
assign w9314 = ~w13946 & w11068;
assign w9315 = w7133 & ~w12629;
assign w9316 = ~w7459 & w11861;
assign w9317 = w1697 & ~w5095;
assign w9318 = ~w8644 & ~w1292;
assign w9319 = w11670 & ~w5768;
assign w9320 = (~w14114 & w5116) | (~w14114 & w22) | (w5116 & w22);
assign w9321 = ~w6 & w11751;
assign w9322 = w8465 & w3891;
assign w9323 = w6659 & w244;
assign w9324 = w1101 & ~w50;
assign w9325 = w9817 & w11516;
assign w9326 = w6886 & w5002;
assign w9327 = ~w4921 & w2178;
assign w9328 = ~w9168 & ~w14638;
assign w9329 = w14506 & w11002;
assign w9330 = (w11429 & w10947) | (w11429 & w7791) | (w10947 & w7791);
assign w9331 = (w12125 & ~w9298) | (w12125 & w13269) | (~w9298 & w13269);
assign w9332 = ~w3689 & ~w8308;
assign w9333 = w9284 & ~w4270;
assign w9334 = w6665 & w10054;
assign w9335 = w3734 & ~w14491;
assign w9336 = ~w7488 & w13828;
assign w9337 = ~w10483 & ~w2110;
assign w9338 = ~w10075 & ~w12943;
assign w9339 = w1250 & w7689;
assign w9340 = w8740 & ~w11117;
assign w9341 = w8335 & w662;
assign w9342 = ~w142 & ~w8459;
assign w9343 = w4503 & ~w4424;
assign w9344 = w2332 & ~w9817;
assign w9345 = (~w13256 & w12359) | (~w13256 & w11437) | (w12359 & w11437);
assign w9346 = ~w4464 & ~w11212;
assign w9347 = ~w6580 & w13210;
assign w9348 = (~w9788 & w12983) | (~w9788 & w13034) | (w12983 & w13034);
assign w9349 = ~w9794 & w3289;
assign w9350 = w1873 & ~w7190;
assign w9351 = (w9776 & w9012) | (w9776 & w13467) | (w9012 & w13467);
assign w9352 = w10290 & w10708;
assign w9353 = w6135 & ~w10699;
assign w9354 = w13346 & w10470;
assign w9355 = ~w14486 & ~w4259;
assign w9356 = w5412 & w5778;
assign w9357 = w5754 & ~w7754;
assign w9358 = w2449 & w8975;
assign w9359 = w3717 & w8900;
assign w9360 = (~w7455 & w1166) | (~w7455 & w12979) | (w1166 & w12979);
assign w9361 = (~w4269 & ~w1840) | (~w4269 & w14215) | (~w1840 & w14215);
assign w9362 = ~w4595 & w6184;
assign w9363 = (w13685 & w12947) | (w13685 & w6955) | (w12947 & w6955);
assign w9364 = w3015 & ~w10923;
assign w9365 = w11779 & w13401;
assign w9366 = ~w5693 & ~w3508;
assign w9367 = ~w10339 & w14038;
assign w9368 = ~w4974 & ~w5899;
assign w9369 = ~w3734 & w14151;
assign w9370 = (~w1789 & w10886) | (~w1789 & w9091) | (w10886 & w9091);
assign w9371 = ~w7814 & ~w9901;
assign w9372 = (~w5601 & w9297) | (~w5601 & w583) | (w9297 & w583);
assign w9373 = (w5341 & w12451) | (w5341 & w9606) | (w12451 & w9606);
assign w9374 = w8785 & ~w12122;
assign w9375 = ~w13282 & w8099;
assign w9376 = ~w14048 & w11708;
assign w9377 = (w4855 & ~w2492) | (w4855 & w14342) | (~w2492 & w14342);
assign w9378 = w10830 & w11324;
assign w9379 = w5852 & w13565;
assign w9380 = w7596 & ~w7467;
assign w9381 = w6436 & w7724;
assign w9382 = ~w5379 & w5316;
assign w9383 = w6230 & ~w2591;
assign w9384 = w2656 & w5742;
assign w9385 = ~w10841 & ~w6361;
assign w9386 = (~w3885 & w4339) | (~w3885 & w13140) | (w4339 & w13140);
assign w9387 = ~w283 & w1610;
assign w9388 = w7794 & ~w10643;
assign w9389 = w3751 & ~w11031;
assign w9390 = w705 & w5024;
assign w9391 = (w5977 & w2916) | (w5977 & w1603) | (w2916 & w1603);
assign w9392 = ~w10349 & w4543;
assign w9393 = ~w6820 & ~w4618;
assign w9394 = w2544 & ~w12483;
assign w9395 = w10032 & ~w5218;
assign w9396 = ~w13587 & w5889;
assign w9397 = ~w11924 & w2518;
assign w9398 = (w6218 & ~w12944) | (w6218 & w324) | (~w12944 & w324);
assign w9399 = ~w4700 & w9211;
assign w9400 = (~w7125 & ~w12165) | (~w7125 & w8622) | (~w12165 & w8622);
assign w9401 = w509 & w5345;
assign w9402 = ~w6856 & w838;
assign w9403 = ~w3751 & ~w12087;
assign w9404 = (w2939 & w10726) | (w2939 & w1921) | (w10726 & w1921);
assign w9405 = w2486 & ~w5193;
assign w9406 = w2656 & w7227;
assign w9407 = (w14038 & ~w7833) | (w14038 & ~w9324) | (~w7833 & ~w9324);
assign w9408 = (w7082 & w4368) | (w7082 & w1408) | (w4368 & w1408);
assign w9409 = ~w5522 & w3904;
assign w9410 = ~w12300 & ~w14081;
assign w9411 = ~w11799 & ~w12403;
assign w9412 = b21 & a21;
assign w9413 = (~w4050 & w14244) | (~w4050 & w7291) | (w14244 & w7291);
assign w9414 = w8412 & ~w3209;
assign w9415 = ~w13511 & w12754;
assign w9416 = (w6486 & w9450) | (w6486 & w14353) | (w9450 & w14353);
assign w9417 = ~w1293 & w3904;
assign w9418 = ~w7484 & ~w874;
assign w9419 = w8931 & w2302;
assign w9420 = ~w7031 & ~w12362;
assign w9421 = ~w8280 & ~w7681;
assign w9422 = ~w6391 & w953;
assign w9423 = (w6042 & w3053) | (w6042 & w11316) | (w3053 & w11316);
assign w9424 = ~w10225 & w3325;
assign w9425 = (w4127 & w13122) | (w4127 & w9056) | (w13122 & w9056);
assign w9426 = ~w2610 & ~w218;
assign w9427 = ~w2625 & ~w7368;
assign w9428 = (~w9714 & w12772) | (~w9714 & w8257) | (w12772 & w8257);
assign w9429 = w13276 & w6106;
assign w9430 = w12317 & ~w2410;
assign w9431 = ~w2492 & w312;
assign w9432 = w6287 & w4969;
assign w9433 = ~w5098 & ~w12895;
assign w9434 = w607 & ~w12642;
assign w9435 = ~w10590 & ~w5918;
assign w9436 = ~w11095 & ~w5942;
assign w9437 = ~w10251 & w11309;
assign w9438 = (~w8179 & ~w8943) | (~w8179 & w10536) | (~w8943 & w10536);
assign w9439 = ~w4700 & w3405;
assign w9440 = ~w7628 & ~w13240;
assign w9441 = (w11870 & w11206) | (w11870 & ~w3798) | (w11206 & ~w3798);
assign w9442 = w13914 & w7618;
assign w9443 = w12460 & ~w14297;
assign w9444 = ~w142 & ~w5282;
assign w9445 = (w13635 & ~w12165) | (w13635 & w8657) | (~w12165 & w8657);
assign w9446 = ~w3946 & w2409;
assign w9447 = (~w852 & ~w3044) | (~w852 & w77) | (~w3044 & w77);
assign w9448 = ~w8234 & w4190;
assign w9449 = ~w12003 & w9240;
assign w9450 = w10993 & ~w6208;
assign w9451 = (~w2951 & w7519) | (~w2951 & w3751) | (w7519 & w3751);
assign w9452 = ~w1751 & w14160;
assign w9453 = b75 & a75;
assign w9454 = w9183 & w4658;
assign w9455 = w11602 & w13208;
assign w9456 = (~w254 & w6227) | (~w254 & w11281) | (w6227 & w11281);
assign w9457 = (w1842 & w922) | (w1842 & w10070) | (w922 & w10070);
assign w9458 = (~w5090 & w155) | (~w5090 & w3041) | (w155 & w3041);
assign w9459 = (w13685 & w3595) | (w13685 & w5249) | (w3595 & w5249);
assign w9460 = w13821 & w13741;
assign w9461 = ~w10756 & w13581;
assign w9462 = (w9921 & w2614) | (w9921 & ~w11416) | (w2614 & ~w11416);
assign w9463 = (w10707 & w6771) | (w10707 & w11925) | (w6771 & w11925);
assign w9464 = (w4625 & ~w2364) | (w4625 & w11290) | (~w2364 & w11290);
assign w9465 = b83 & a83;
assign w9466 = ~w922 & w11810;
assign w9467 = (w13193 & w7598) | (w13193 & ~w9034) | (w7598 & ~w9034);
assign w9468 = ~w1096 & ~w1009;
assign w9469 = w4024 & ~w13668;
assign w9470 = (w5927 & w12864) | (w5927 & w5319) | (w12864 & w5319);
assign w9471 = ~w6415 & ~w9905;
assign w9472 = w4711 & ~w12554;
assign w9473 = (w6103 & w13449) | (w6103 & w12786) | (w13449 & w12786);
assign w9474 = w14518 & w7049;
assign w9475 = ~w8935 & w1833;
assign w9476 = w2728 & w13197;
assign w9477 = ~w12271 & ~w10471;
assign w9478 = (~w7464 & w1319) | (~w7464 & w12222) | (w1319 & w12222);
assign w9479 = ~w9284 & ~w14058;
assign w9480 = ~b101 & ~a101;
assign w9481 = w14278 & w5675;
assign w9482 = w827 & ~w14267;
assign w9483 = w8234 & w13531;
assign w9484 = (~w14492 & w2437) | (~w14492 & w9080) | (w2437 & w9080);
assign w9485 = ~w71 & w12931;
assign w9486 = ~w14664 & w611;
assign w9487 = ~w3516 & ~w3451;
assign w9488 = (~w1351 & w7465) | (~w1351 & w5443) | (w7465 & w5443);
assign w9489 = w798 & ~w13409;
assign w9490 = (w12532 & w9402) | (w12532 & w8193) | (w9402 & w8193);
assign w9491 = w3024 & ~w14659;
assign w9492 = ~w5177 & w10704;
assign w9493 = ~w13762 & w4289;
assign w9494 = w6854 & w1306;
assign w9495 = (~w14385 & ~w9172) | (~w14385 & w847) | (~w9172 & w847);
assign w9496 = ~w14509 & w1904;
assign w9497 = ~w12762 & w3752;
assign w9498 = ~w7369 & ~w9421;
assign w9499 = w3427 & w11117;
assign w9500 = (~w6500 & w7922) | (~w6500 & w2213) | (w7922 & w2213);
assign w9501 = w5294 & w8827;
assign w9502 = (w5471 & ~w4143) | (w5471 & w14126) | (~w4143 & w14126);
assign w9503 = w4848 & w11871;
assign w9504 = w13531 & w7423;
assign w9505 = ~w8330 & ~w379;
assign w9506 = ~b93 & ~w13008;
assign w9507 = ~w9012 & w6216;
assign w9508 = ~w12266 & w5962;
assign w9509 = (w10488 & w133) | (w10488 & w3481) | (w133 & w3481);
assign w9510 = w12125 & w5780;
assign w9511 = ~w1118 & w13045;
assign w9512 = w12575 & w10855;
assign w9513 = (~w9817 & w3209) | (~w9817 & w9344) | (w3209 & w9344);
assign w9514 = (w11037 & w9724) | (w11037 & ~w9096) | (w9724 & ~w9096);
assign w9515 = ~w9012 & w13926;
assign w9516 = w347 & w13628;
assign w9517 = w10523 & w8459;
assign w9518 = ~w8088 & w8246;
assign w9519 = w10339 & ~w2261;
assign w9520 = ~w1868 & ~w13135;
assign w9521 = (w6023 & w14602) | (w6023 & ~w9262) | (w14602 & ~w9262);
assign w9522 = w13864 & w1540;
assign w9523 = w2850 & ~w9570;
assign w9524 = w5893 & ~w2943;
assign w9525 = ~w6203 & w10690;
assign w9526 = ~w142 & ~w11934;
assign w9527 = ~w14664 & w12316;
assign w9528 = ~w8422 & w9011;
assign w9529 = (w1013 & w4285) | (w1013 & ~w4007) | (w4285 & ~w4007);
assign w9530 = (w5118 & w3695) | (w5118 & w9292) | (w3695 & w9292);
assign w9531 = ~w10935 & w3963;
assign w9532 = (w11895 & ~w5174) | (w11895 & ~w6627) | (~w5174 & ~w6627);
assign w9533 = ~w2175 & w9044;
assign w9534 = (~w195 & w11657) | (~w195 & w2305) | (w11657 & w2305);
assign w9535 = ~w13222 & w13526;
assign w9536 = (w4127 & w8389) | (w4127 & w7877) | (w8389 & w7877);
assign w9537 = (w1816 & w14449) | (w1816 & w13703) | (w14449 & w13703);
assign w9538 = (w10115 & w5154) | (w10115 & w6780) | (w5154 & w6780);
assign w9539 = w309 & ~w9748;
assign w9540 = w9788 & ~w3904;
assign w9541 = ~w12497 & ~w3482;
assign w9542 = w1880 & ~w12529;
assign w9543 = ~w4166 & w8989;
assign w9544 = ~w2664 & ~w8971;
assign w9545 = (w8769 & ~w3629) | (w8769 & w11585) | (~w3629 & w11585);
assign w9546 = a0 & b0;
assign w9547 = w2225 & w6494;
assign w9548 = ~w9265 & w11371;
assign w9549 = ~w1114 & ~w1071;
assign w9550 = (~w11803 & w9209) | (~w11803 & w7830) | (w9209 & w7830);
assign w9551 = ~w3457 & w13657;
assign w9552 = (w7754 & w12825) | (w7754 & w12318) | (w12825 & w12318);
assign w9553 = (~w6542 & w12620) | (~w6542 & w12547) | (w12620 & w12547);
assign w9554 = (~w7064 & ~w5237) | (~w7064 & w9577) | (~w5237 & w9577);
assign w9555 = ~w8840 & ~w6231;
assign w9556 = w12654 & w866;
assign w9557 = (w6399 & w9532) | (w6399 & w14191) | (w9532 & w14191);
assign w9558 = ~w1276 & ~w9383;
assign w9559 = w8294 & w9716;
assign w9560 = w3345 & ~w8400;
assign w9561 = (w11708 & ~w5294) | (w11708 & w8331) | (~w5294 & w8331);
assign w9562 = (w13288 & w2562) | (w13288 & w14182) | (w2562 & w14182);
assign w9563 = ~w13122 & w3007;
assign w9564 = ~w10847 & w7613;
assign w9565 = (w11675 & ~w3209) | (w11675 & w10607) | (~w3209 & w10607);
assign w9566 = ~w6864 & ~w4583;
assign w9567 = w10974 & ~w9298;
assign w9568 = ~w1802 & ~w5842;
assign w9569 = ~w12825 & w12622;
assign w9570 = w2387 & w11500;
assign w9571 = w5657 & w926;
assign w9572 = ~w922 & ~w5050;
assign w9573 = (~w7784 & w1915) | (~w7784 & w1832) | (w1915 & w1832);
assign w9574 = (w6637 & w11425) | (w6637 & w4128) | (w11425 & w4128);
assign w9575 = (w7376 & w7943) | (w7376 & w6885) | (w7943 & w6885);
assign w9576 = w5002 & ~w7811;
assign w9577 = ~w5751 & ~w7064;
assign w9578 = ~w13594 & w3459;
assign w9579 = w14302 & ~w10223;
assign w9580 = w8742 & w8769;
assign w9581 = (w11708 & w3809) | (w11708 & w11489) | (w3809 & w11489);
assign w9582 = w10645 & ~w10013;
assign w9583 = ~b70 & ~a70;
assign w9584 = ~w3209 & w3732;
assign w9585 = ~w1563 & w4627;
assign w9586 = w10116 & ~w1086;
assign w9587 = ~w11243 & w10336;
assign w9588 = (~w12958 & w1842) | (~w12958 & ~w4032) | (w1842 & ~w4032);
assign w9589 = w7526 & w1855;
assign w9590 = ~w12321 & ~w3038;
assign w9591 = (w6276 & w7041) | (w6276 & w7062) | (w7041 & w7062);
assign w9592 = (w11429 & w3850) | (w11429 & w8910) | (w3850 & w8910);
assign w9593 = w7794 & ~w2684;
assign w9594 = ~w387 & w5145;
assign w9595 = w1246 & w12047;
assign w9596 = ~w3790 & ~w6795;
assign w9597 = (~w1362 & w943) | (~w1362 & w1788) | (w943 & w1788);
assign w9598 = (w8515 & w3396) | (w8515 & w11664) | (w3396 & w11664);
assign w9599 = w4284 & w7278;
assign w9600 = ~w11732 | ~w9655;
assign w9601 = w5825 & ~w6550;
assign w9602 = w9153 & ~w6834;
assign w9603 = ~w1048 & w5241;
assign w9604 = ~w6761 & w5548;
assign w9605 = w9265 & ~w10485;
assign w9606 = w1143 & w5341;
assign w9607 = (~w12438 & w3435) | (~w12438 & w5320) | (w3435 & w5320);
assign w9608 = w2637 & ~w13004;
assign w9609 = (w723 & w14253) | (w723 & w1947) | (w14253 & w1947);
assign w9610 = ~w13938 & w12311;
assign w9611 = w5322 & w6212;
assign w9612 = w7491 & w7197;
assign w9613 = b25 & a25;
assign w9614 = ~w3803 & ~w10781;
assign w9615 = w14395 & ~w894;
assign w9616 = w3550 & w9277;
assign w9617 = (~w12056 & w3323) | (~w12056 & w11036) | (w3323 & w11036);
assign w9618 = w5741 & ~w9296;
assign w9619 = w12148 & ~w6583;
assign w9620 = w7772 & w6230;
assign w9621 = w4949 & ~w11145;
assign w9622 = (~w10317 & ~w14515) | (~w10317 & w5670) | (~w14515 & w5670);
assign w9623 = ~b50 & ~a50;
assign w9624 = w10849 & ~w6639;
assign w9625 = ~w254 & w12658;
assign w9626 = ~w12321 & w5397;
assign w9627 = w5937 & w937;
assign w9628 = ~w2218 & w11728;
assign w9629 = w7080 & w9748;
assign w9630 = (w10210 & w805) | (w10210 & w11489) | (w805 & w11489);
assign w9631 = w4213 & w12662;
assign w9632 = ~w922 & ~w9004;
assign w9633 = w9509 & ~w7921;
assign w9634 = ~w2397 & ~w13992;
assign w9635 = ~w7681 & w13562;
assign w9636 = w2606 & w12566;
assign w9637 = (w14072 & w13587) | (w14072 & w54) | (w13587 & w54);
assign w9638 = (~w10757 & w8727) | (~w10757 & w5994) | (w8727 & w5994);
assign w9639 = (w12441 & w9035) | (w12441 & w9847) | (w9035 & w9847);
assign w9640 = (w10386 & ~w4167) | (w10386 & w2146) | (~w4167 & w2146);
assign w9641 = ~w6250 & w11646;
assign w9642 = (w8650 & w13736) | (w8650 & w99) | (w13736 & w99);
assign w9643 = ~w8507 & w10845;
assign w9644 = w1872 & ~w12153;
assign w9645 = (w3128 & w460) | (w3128 & w5966) | (w460 & w5966);
assign w9646 = (~w475 & w13335) | (~w475 & w4330) | (w13335 & w4330);
assign w9647 = (w1842 & w8226) | (w1842 & w13483) | (w8226 & w13483);
assign w9648 = (w13685 & w7729) | (w13685 & w10803) | (w7729 & w10803);
assign w9649 = w12295 & ~w5984;
assign w9650 = ~w5522 & w2701;
assign w9651 = w9328 & w8184;
assign w9652 = (w11791 & ~w4840) | (w11791 & w140) | (~w4840 & w140);
assign w9653 = (~w4921 & w10626) | (~w4921 & w6962) | (w10626 & w6962);
assign w9654 = w1389 & ~w10483;
assign w9655 = ~w5732 & ~w5397;
assign w9656 = ~w7717 & ~w4855;
assign w9657 = (~w1460 & w3947) | (~w1460 & w3204) | (w3947 & w3204);
assign w9658 = (w9013 & ~w8562) | (w9013 & w5349) | (~w8562 & w5349);
assign w9659 = (w5932 & w13324) | (w5932 & w10582) | (w13324 & w10582);
assign w9660 = ~w9801 & ~w4446;
assign w9661 = w10704 & ~w8389;
assign w9662 = (w10685 & w8998) | (w10685 & ~w11091) | (w8998 & ~w11091);
assign w9663 = (w3626 & w5698) | (w3626 & w6276) | (w5698 & w6276);
assign w9664 = ~w7981 & w465;
assign w9665 = (~w1413 & w11496) | (~w1413 & w8210) | (w11496 & w8210);
assign w9666 = ~w2762 & w50;
assign w9667 = ~w2656 & w14227;
assign w9668 = ~w8367 & w9512;
assign w9669 = ~w7244 & ~w13323;
assign w9670 = ~w5412 & ~w475;
assign w9671 = ~w6716 & ~w8234;
assign w9672 = ~w6889 & ~w2962;
assign w9673 = ~w10071 & w14301;
assign w9674 = ~w325 & ~w3885;
assign w9675 = ~w2175 & w6788;
assign w9676 = ~w3597 & ~w9496;
assign w9677 = w3914 & w1036;
assign w9678 = (~w11973 & w7775) | (~w11973 & w3188) | (w7775 & w3188);
assign w9679 = w11031 & w8459;
assign w9680 = w945 & w3533;
assign w9681 = (~w11091 & w2885) | (~w11091 & w6602) | (w2885 & w6602);
assign w9682 = ~w5702 & w10998;
assign w9683 = w7085 & ~w11241;
assign w9684 = (w3040 & w9982) | (w3040 & ~w5031) | (w9982 & ~w5031);
assign w9685 = w3576 & ~w10775;
assign w9686 = ~w8100 & w12420;
assign w9687 = w6716 & ~w5845;
assign w9688 = (~w10853 & ~w6266) | (~w10853 & w6685) | (~w6266 & w6685);
assign w9689 = ~w1563 & w6700;
assign w9690 = w4505 & ~w12508;
assign w9691 = (~w11936 & w6974) | (~w11936 & w8114) | (w6974 & w8114);
assign w9692 = w12088 & ~w5243;
assign w9693 = w9861 & ~w9211;
assign w9694 = ~w9226 & ~w6542;
assign w9695 = w12079 & ~w11147;
assign w9696 = ~w13587 & w12014;
assign w9697 = (~w4479 & w9942) | (~w4479 & w14255) | (w9942 & w14255);
assign w9698 = (w7774 & w13549) | (w7774 & ~w4783) | (w13549 & ~w4783);
assign w9699 = ~w571 & ~w9026;
assign w9700 = (w14048 & ~w189) | (w14048 & w9731) | (~w189 & w9731);
assign w9701 = (w11604 & w2313) | (w11604 & w6995) | (w2313 & w6995);
assign w9702 = (~w3019 & ~w11147) | (~w3019 & w4450) | (~w11147 & w4450);
assign w9703 = ~w3068 & ~w8092;
assign w9704 = ~w10864 & ~w7309;
assign w9705 = (~w14463 & w12930) | (~w14463 & w11509) | (w12930 & w11509);
assign w9706 = w5522 & w10699;
assign w9707 = (w13281 & w3584) | (w13281 & w1613) | (w3584 & w1613);
assign w9708 = (~w125 & ~w9046) | (~w125 & w1095) | (~w9046 & w1095);
assign w9709 = ~w8499 & ~w2381;
assign w9710 = (w5156 & w9796) | (w5156 & w2626) | (w9796 & w2626);
assign w9711 = ~w8929 & ~w7613;
assign w9712 = b53 & ~w5852;
assign w9713 = w1873 & w9672;
assign w9714 = (~w1692 & w6363) | (~w1692 & w223) | (w6363 & w223);
assign w9715 = w12377 & ~w3636;
assign w9716 = (~w7889 & w7000) | (~w7889 & w3407) | (w7000 & w3407);
assign w9717 = ~w11547 & ~w9902;
assign w9718 = (w12915 & w9784) | (w12915 & ~w11708) | (w9784 & ~w11708);
assign w9719 = ~w7305 & ~w843;
assign w9720 = (w8943 & w10581) | (w8943 & w672) | (w10581 & w672);
assign w9721 = ~w1503 | ~w1928;
assign w9722 = w4425 & w6230;
assign w9723 = ~w11012 & w2781;
assign w9724 = w9607 & ~w13518;
assign w9725 = (~w5607 & ~w6320) | (~w5607 & w14349) | (~w6320 & w14349);
assign w9726 = (w5768 & w13772) | (w5768 & w9724) | (w13772 & w9724);
assign w9727 = (~w8347 & w1984) | (~w8347 & w13140) | (w1984 & w13140);
assign w9728 = w6436 & ~w1062;
assign w9729 = (w14059 & w5159) | (w14059 & w2181) | (w5159 & w2181);
assign w9730 = (w749 & w10767) | (w749 & w9139) | (w10767 & w9139);
assign w9731 = w14048 & w9294;
assign w9732 = ~w9608 & w7977;
assign w9733 = (~w9403 & w8282) | (~w9403 & ~w3798) | (w8282 & ~w3798);
assign w9734 = w11460 & ~w14433;
assign w9735 = ~w621 & w4987;
assign w9736 = (w8288 & w63) | (w8288 & w3933) | (w63 & w3933);
assign w9737 = w4658 & w7317;
assign w9738 = (w4187 & ~w14279) | (w4187 & w12585) | (~w14279 & w12585);
assign w9739 = (w8405 & w12184) | (w8405 & w8281) | (w12184 & w8281);
assign w9740 = w6558 & ~w7079;
assign w9741 = ~w5867 & w545;
assign w9742 = (~w5879 & w1891) | (~w5879 & w5686) | (w1891 & w5686);
assign w9743 = ~w13599 & ~w7436;
assign w9744 = ~w5948 & ~w2729;
assign w9745 = (~w10637 & w2734) | (~w10637 & w6899) | (w2734 & w6899);
assign w9746 = (w10318 & w4034) | (w10318 & w3489) | (w4034 & w3489);
assign w9747 = ~w9287 & w13394;
assign w9748 = ~w1490 & w5177;
assign w9749 = (w12568 & w2105) | (w12568 & w4426) | (w2105 & w4426);
assign w9750 = ~w11796 & w5855;
assign w9751 = w3075 & ~w11117;
assign w9752 = ~w14302 & w14390;
assign w9753 = w11846 & w3297;
assign w9754 = w533 & ~w13572;
assign w9755 = ~w3340 & w8321;
assign w9756 = w6301 & w1436;
assign w9757 = ~w3288 & ~w2729;
assign w9758 = (w3611 & w10462) | (w3611 & w417) | (w10462 & w417);
assign w9759 = (w11855 & ~w5325) | (w11855 & w5313) | (~w5325 & w5313);
assign w9760 = ~w1821 & w6845;
assign w9761 = w5522 & w5282;
assign w9762 = ~w9654 & w7773;
assign w9763 = (w1986 & w5563) | (w1986 & w403) | (w5563 & w403);
assign w9764 = ~w12821 & w2928;
assign w9765 = ~w1712 & w4823;
assign w9766 = w3019 & w4541;
assign w9767 = ~w4512 & w6472;
assign w9768 = ~w11868 & ~w13402;
assign w9769 = ~w12460 & ~w387;
assign w9770 = (w11815 & w14306) | (w11815 & w9339) | (w14306 & w9339);
assign w9771 = (w4545 & w4681) | (w4545 & w6132) | (w4681 & w6132);
assign w9772 = ~w13158 & w7569;
assign w9773 = w5794 & w11606;
assign w9774 = w7025 & w11053;
assign w9775 = ~w4607 & w12284;
assign w9776 = (~w14526 & w5036) | (~w14526 & w11372) | (w5036 & w11372);
assign w9777 = (w10123 & w5232) | (w10123 & w5640) | (w5232 & w5640);
assign w9778 = w9839 & ~w14584;
assign w9779 = w14278 & w3919;
assign w9780 = w4367 & w10555;
assign w9781 = w2433 & ~w13323;
assign w9782 = ~w7305 & w3963;
assign w9783 = (w11106 & w14229) | (w11106 & ~w378) | (w14229 & ~w378);
assign w9784 = w7348 & w12915;
assign w9785 = w4336 & w2703;
assign w9786 = ~w12135 & w5615;
assign w9787 = ~w13152 & w5041;
assign w9788 = ~b52 & ~a52;
assign w9789 = (w6215 & w7269) | (w6215 & w2547) | (w7269 & w2547);
assign w9790 = ~w7348 & w6364;
assign w9791 = w13844 & w13169;
assign w9792 = (w11287 & ~w761) | (w11287 & w7944) | (~w761 & w7944);
assign w9793 = (~w12406 & w3403) | (~w12406 & w12263) | (w3403 & w12263);
assign w9794 = ~w13423 & ~w12922;
assign w9795 = ~w11926 & w7503;
assign w9796 = ~w5113 & ~w13546;
assign w9797 = w2278 & ~w6329;
assign w9798 = ~w6536 & ~w5785;
assign w9799 = ~w6572 & w9590;
assign w9800 = (w10433 & w13715) | (w10433 & w7992) | (w13715 & w7992);
assign w9801 = ~w5562 & w13513;
assign w9802 = ~w1247 & ~w12919;
assign w9803 = w13620 & w1599;
assign w9804 = (w3055 & w6011) | (w3055 & w10000) | (w6011 & w10000);
assign w9805 = ~w7190 & ~w12060;
assign w9806 = (~w2218 & w14342) | (~w2218 & w10479) | (w14342 & w10479);
assign w9807 = ~w13233 & ~w5231;
assign w9808 = (w9433 & w4099) | (w9433 & w14452) | (w4099 & w14452);
assign w9809 = (~w475 & w3835) | (~w475 & w9670) | (w3835 & w9670);
assign w9810 = ~w12351 & w3686;
assign w9811 = w4109 & w9160;
assign w9812 = ~w10517 & w2701;
assign w9813 = ~w12811 & ~w14507;
assign w9814 = (w4458 & ~w9952) | (w4458 & w13641) | (~w9952 & w13641);
assign w9815 = (~w1692 & w6363) | (~w1692 & w8390) | (w6363 & w8390);
assign w9816 = ~w6375 & ~w6068;
assign w9817 = ~w6889 & ~w2332;
assign w9818 = ~w13668 & w11910;
assign w9819 = (w13180 & ~w14514) | (w13180 & w7888) | (~w14514 & w7888);
assign w9820 = ~w11287 & w7670;
assign w9821 = w8409 & ~w3209;
assign w9822 = ~w12003 & w4350;
assign w9823 = ~w4700 & w6689;
assign w9824 = w12414 & w4090;
assign w9825 = w3438 & w11318;
assign w9826 = (w1859 & w5815) | (w1859 & ~w2457) | (w5815 & ~w2457);
assign w9827 = ~w12121 & w2410;
assign w9828 = ~w4836 & w7906;
assign w9829 = (~w3904 & ~w10862) | (~w3904 & ~w2633) | (~w10862 & ~w2633);
assign w9830 = w13620 & ~w11855;
assign w9831 = w1692 & w12170;
assign w9832 = (w5070 & w14003) | (w5070 & w461) | (w14003 & w461);
assign w9833 = w7085 & w6349;
assign w9834 = w8847 & w12485;
assign w9835 = w12664 & w3427;
assign w9836 = ~w5353 & w12082;
assign w9837 = ~w13163 & w8674;
assign w9838 = ~w4269 & ~w12958;
assign w9839 = w9087 & w5788;
assign w9840 = (~w988 & w1038) | (~w988 & w559) | (w1038 & w559);
assign w9841 = (w13580 & w3523) | (w13580 & w181) | (w3523 & w181);
assign w9842 = w5556 & ~w5490;
assign w9843 = (w719 & w12783) | (w719 & w13626) | (w12783 & w13626);
assign w9844 = w13148 & ~w2992;
assign w9845 = ~w10077 & w2653;
assign w9846 = ~b118 & ~a118;
assign w9847 = ~w2799 & w9834;
assign w9848 = ~w1614 & ~w13008;
assign w9849 = (w9541 & w11187) | (w9541 & w249) | (w11187 & w249);
assign w9850 = ~w12459 & ~w14253;
assign w9851 = (w4318 & w13051) | (w4318 & w1281) | (w13051 & w1281);
assign w9852 = ~w8226 & w145;
assign w9853 = ~w11891 & ~w6941;
assign w9854 = w7794 & ~w11;
assign w9855 = ~w2081 & ~w3159;
assign w9856 = ~w9541 & w14648;
assign w9857 = w9170 & w6175;
assign w9858 = w10391 & w7056;
assign w9859 = ~w9004 & w709;
assign w9860 = (~w8431 & w8736) | (~w8431 & w6509) | (w8736 & w6509);
assign w9861 = (~w3885 & w5772) | (~w3885 & w10046) | (w5772 & w10046);
assign w9862 = ~w14486 & w12893;
assign w9863 = ~w10119 & w309;
assign w9864 = (~w2228 & w13652) | (~w2228 & w3429) | (w13652 & w3429);
assign w9865 = w3309 & w10733;
assign w9866 = w8442 & w7762;
assign w9867 = w5560 & ~w12463;
assign w9868 = w4307 & w13008;
assign w9869 = (~w7962 & w13324) | (~w7962 & w3985) | (w13324 & w3985);
assign w9870 = ~w907 & w12599;
assign w9871 = ~b72 & ~a72;
assign w9872 = (~w2492 & w11974) | (~w2492 & w14575) | (w11974 & w14575);
assign w9873 = (w10386 & ~w4167) | (w10386 & w10559) | (~w4167 & w10559);
assign w9874 = ~w1559 & w7861;
assign w9875 = ~w9012 & w14149;
assign w9876 = (w13896 & w6506) | (w13896 & ~w13668) | (w6506 & ~w13668);
assign w9877 = ~w2674 & w7204;
assign w9878 = w14545 & ~w4154;
assign w9879 = w10512 & w8084;
assign w9880 = ~w894 & w9226;
assign w9881 = (w4370 & w7201) | (w4370 & w9034) | (w7201 & w9034);
assign w9882 = w1257 & w4483;
assign w9883 = w13973 & w3149;
assign w9884 = ~w4287 & ~w3289;
assign w9885 = w10032 & w5282;
assign w9886 = ~w11172 & ~w7617;
assign w9887 = (w6973 & ~w7804) | (w6973 & ~w11186) | (~w7804 & ~w11186);
assign w9888 = w6572 & ~w5732;
assign w9889 = (~w7782 & w9817) | (~w7782 & w10026) | (w9817 & w10026);
assign w9890 = ~w8226 & w8800;
assign w9891 = (w1593 & w11060) | (w1593 & w2457) | (w11060 & w2457);
assign w9892 = (w1416 & w14415) | (w1416 & w4347) | (w14415 & w4347);
assign w9893 = w13189 & w1535;
assign w9894 = ~w6442 & ~w4033;
assign w9895 = ~w14395 & w14585;
assign w9896 = ~w14470 & ~w5785;
assign w9897 = ~w922 & w4485;
assign w9898 = w5593 & w11909;
assign w9899 = (~w9087 & w1166) | (~w9087 & w4345) | (w1166 & w4345);
assign w9900 = w1274 & w10647;
assign w9901 = w14640 & ~w4458;
assign w9902 = b8 & a8;
assign w9903 = (~w6949 & w13122) | (~w6949 & w9257) | (w13122 & w9257);
assign w9904 = (~w7782 & w765) | (~w7782 & w1791) | (w765 & w1791);
assign w9905 = ~w2317 & w9689;
assign w9906 = (w218 & w2175) | (w218 & w2543) | (w2175 & w2543);
assign w9907 = w7808 & w7535;
assign w9908 = ~w2228 & w4458;
assign w9909 = ~w8900 & ~w2323;
assign w9910 = w3963 & ~w6692;
assign w9911 = w11560 & ~w3786;
assign w9912 = (~w11429 & w10660) | (~w11429 & w4277) | (w10660 & w4277);
assign w9913 = ~w8561 & w11364;
assign w9914 = (w1814 & w13936) | (w1814 & w13471) | (w13936 & w13471);
assign w9915 = w12077 & w10706;
assign w9916 = ~w870 & w2492;
assign w9917 = w11722 & ~w9937;
assign w9918 = (w9305 & w1350) | (w9305 & w2546) | (w1350 & w2546);
assign w9919 = w5569 & w9817;
assign w9920 = (w8085 & w2175) | (w8085 & w7316) | (w2175 & w7316);
assign w9921 = ~w829 & ~w2320;
assign w9922 = (w10210 & w805) | (w10210 & ~w7853) | (w805 & ~w7853);
assign w9923 = (~w6483 & w9127) | (~w6483 & w13419) | (w9127 & w13419);
assign w9924 = w3153 & w9300;
assign w9925 = ~w4322 & w6436;
assign w9926 = (~w10435 & w12449) | (~w10435 & w10817) | (w12449 & w10817);
assign w9927 = ~b120 & ~a120;
assign w9928 = (~w3798 & w12154) | (~w3798 & ~w9364) | (w12154 & ~w9364);
assign w9929 = ~w3815 & w6707;
assign w9930 = (~w8277 & w11209) | (~w8277 & w1999) | (w11209 & w1999);
assign w9931 = ~w8149 & w908;
assign w9932 = ~w2933 & ~w3958;
assign w9933 = ~w2656 & w309;
assign w9934 = (w1300 & w9008) | (w1300 & w6589) | (w9008 & w6589);
assign w9935 = ~w12464 & ~w746;
assign w9936 = ~w14098 & ~w6933;
assign w9937 = ~w14105 & ~w9025;
assign w9938 = w2332 & w1873;
assign w9939 = ~w607 & w13937;
assign w9940 = ~w3036 & ~w2922;
assign w9941 = (w8288 & w14234) | (w8288 & w3080) | (w14234 & w3080);
assign w9942 = (w1300 & w9008) | (w1300 & w217) | (w9008 & w217);
assign w9943 = w10676 & w12398;
assign w9944 = w8855 & w12695;
assign w9945 = (w7907 & w12287) | (w7907 & w12640) | (w12287 & w12640);
assign w9946 = ~w867 & ~w34;
assign w9947 = (~w7630 & w1903) | (~w7630 & w341) | (w1903 & w341);
assign w9948 = (w5626 & w2470) | (w5626 & w14432) | (w2470 & w14432);
assign w9949 = b32 & a32;
assign w9950 = (~w4071 & w8451) | (~w4071 & w2305) | (w8451 & w2305);
assign w9951 = w9434 & ~w12464;
assign w9952 = w10645 & ~w3407;
assign w9953 = ~w3209 & ~w5607;
assign w9954 = w11013 & ~w6689;
assign w9955 = w9678 & ~w1326;
assign w9956 = (~w9454 & w9012) | (~w9454 & w3711) | (w9012 & w3711);
assign w9957 = ~w7496 & ~w12756;
assign w9958 = w7012 & w1192;
assign w9959 = ~w14078 & w8067;
assign w9960 = w11863 & ~w13113;
assign w9961 = w5741 & w11031;
assign w9962 = ~w2261 & ~w7362;
assign w9963 = (~w10213 & w11606) | (~w10213 & ~w1503) | (w11606 & ~w1503);
assign w9964 = (~w3672 & w14541) | (~w3672 & w10120) | (w14541 & w10120);
assign w9965 = ~w5133 & w5863;
assign w9966 = w9170 | w7707;
assign w9967 = (w2396 & w9131) | (w2396 & ~w14182) | (w9131 & ~w14182);
assign w9968 = (~w77 & w13282) | (~w77 & w13911) | (w13282 & w13911);
assign w9969 = ~w13282 & w884;
assign w9970 = ~w4228 & ~w14010;
assign w9971 = w3826 & w5648;
assign w9972 = ~w13733 & ~w14504;
assign w9973 = ~w9454 & ~w10201;
assign w9974 = ~w12569 & ~w11494;
assign w9975 = ~w12773 & w2925;
assign w9976 = ~w10754 & w13881;
assign w9977 = ~w11691 & ~w5441;
assign w9978 = w1772 & w2107;
assign w9979 = (~w12011 & w815) | (~w12011 & w11022) | (w815 & w11022);
assign w9980 = ~w11356 & w1498;
assign w9981 = ~w4721 & ~w8609;
assign w9982 = w14314 & ~w7319;
assign w9983 = w1387 & w14506;
assign w9984 = (w2941 & ~w6895) | (w2941 & w3473) | (~w6895 & w3473);
assign w9985 = (~w10462 & w1193) | (~w10462 & w14418) | (w1193 & w14418);
assign w9986 = ~w11261 & w587;
assign w9987 = (w7914 & w6124) | (w7914 & w6326) | (w6124 & w6326);
assign w9988 = ~w13544 & w334;
assign w9989 = (w227 & w1918) | (w227 & w2565) | (w1918 & w2565);
assign w9990 = ~w3755 & w4041;
assign w9991 = (w3758 & w6332) | (w3758 & w8228) | (w6332 & w8228);
assign w9992 = w11116 & w8018;
assign w9993 = (~w6101 & w299) | (~w6101 & w103) | (w299 & w103);
assign w9994 = (w11456 & w13424) | (w11456 & ~w12127) | (w13424 & ~w12127);
assign w9995 = (w10115 & w7780) | (w10115 & w14429) | (w7780 & w14429);
assign w9996 = ~w9412 & ~w6267;
assign w9997 = ~w6344 & w6582;
assign w9998 = w3774 & w7085;
assign w9999 = (~w1158 & ~w11803) | (~w1158 & w10330) | (~w11803 & w10330);
assign w10000 = (w12406 & w3607) | (w12406 & w11374) | (w3607 & w11374);
assign w10001 = ~w7534 & ~w12422;
assign w10002 = (~w10435 & w4954) | (~w10435 & w11765) | (w4954 & w11765);
assign w10003 = (w10687 & w2156) | (w10687 & w12537) | (w2156 & w12537);
assign w10004 = (~w6781 & w9876) | (~w6781 & w76) | (w9876 & w76);
assign w10005 = (~w5070 & w2057) | (~w5070 & w7648) | (w2057 & w7648);
assign w10006 = ~w9200 & ~w7317;
assign w10007 = (~w13685 & w3889) | (~w13685 & w6222) | (w3889 & w6222);
assign w10008 = ~w4843 & w10664;
assign w10009 = ~w3602 & w9109;
assign w10010 = w146 & w12361;
assign w10011 = w9925 & w7085;
assign w10012 = ~w4860 & w14056;
assign w10013 = ~b104 & ~a104;
assign w10014 = w13092 & ~w13670;
assign w10015 = (~w11429 & w13232) | (~w11429 & w8712) | (w13232 & w8712);
assign w10016 = ~w10689 & w6113;
assign w10017 = ~w5522 & ~w11031;
assign w10018 = ~w12240 & ~w3823;
assign w10019 = w9503 & ~w9281;
assign w10020 = ~w12809 & w10431;
assign w10021 = (w7376 & w1569) | (w7376 & ~w12294) | (w1569 & ~w12294);
assign w10022 = w7348 & w11108;
assign w10023 = (~w4134 & w2199) | (~w4134 & w3250) | (w2199 & w3250);
assign w10024 = ~w5294 & w12398;
assign w10025 = ~w201 & ~w3177;
assign w10026 = (~w2332 & ~w13282) | (~w2332 & w9817) | (~w13282 & w9817);
assign w10027 = (w1274 & w11894) | (w1274 & w11671) | (w11894 & w11671);
assign w10028 = w4809 & w3105;
assign w10029 = ~w5294 & w693;
assign w10030 = w13533 & w8027;
assign w10031 = ~w5660 & w914;
assign w10032 = b114 & a114;
assign w10033 = (~w318 & w11516) | (~w318 & ~w7538) | (w11516 & ~w7538);
assign w10034 = (w1770 & w8235) | (w1770 & w7041) | (w8235 & w7041);
assign w10035 = w6558 & ~w11461;
assign w10036 = w2872 & w7493;
assign w10037 = ~w12121 & ~w12003;
assign w10038 = (~w13953 & w2144) | (~w13953 & w14022) | (w2144 & w14022);
assign w10039 = ~w7335 & ~w706;
assign w10040 = ~w13249 & ~w5676;
assign w10041 = w9284 & w7154;
assign w10042 = w1096 & w5213;
assign w10043 = ~w12121 & ~w4893;
assign w10044 = w12129 & w9989;
assign w10045 = w1949 & w10689;
assign w10046 = w3742 & ~w3885;
assign w10047 = (~w4507 & ~w13219) | (~w4507 & w3270) | (~w13219 & w3270);
assign w10048 = ~w843 & w10960;
assign w10049 = ~w1138 & w2282;
assign w10050 = ~w13993 & ~w2096;
assign w10051 = ~w5013 & w4529;
assign w10052 = w8740 & ~w7654;
assign w10053 = w8975 & w8517;
assign w10054 = (~w9262 & w9674) | (~w9262 & w2756) | (w9674 & w2756);
assign w10055 = (w6542 & w4158) | (w6542 & w6304) | (w4158 & w6304);
assign w10056 = w11137 & ~w9208;
assign w10057 = (w2144 & w13582) | (w2144 & w4066) | (w13582 & w4066);
assign w10058 = w10409 & w11500;
assign w10059 = w13805 & ~w9434;
assign w10060 = ~w8159 & ~w6830;
assign w10061 = ~w2762 & w10847;
assign w10062 = ~w7982 & w8189;
assign w10063 = (~w13219 & w6801) | (~w13219 & w11736) | (w6801 & w11736);
assign w10064 = w4225 & w12352;
assign w10065 = w5825 & w14262;
assign w10066 = w14640 & ~w2729;
assign w10067 = (w12021 & ~w1878) | (w12021 & ~w5909) | (~w1878 & ~w5909);
assign w10068 = ~w9817 & w3767;
assign w10069 = (w1208 & w53) | (w1208 & ~w10023) | (w53 & ~w10023);
assign w10070 = w1842 & ~w8099;
assign w10071 = ~w12962 & w6650;
assign w10072 = ~w1101 & w806;
assign w10073 = ~w4756 & w1729;
assign w10074 = w5402 & ~w10704;
assign w10075 = b80 & a80;
assign w10076 = ~w1840 & w14659;
assign w10077 = ~w10334 & ~w13722;
assign w10078 = w11560 & ~w8459;
assign w10079 = w14226 & ~w7639;
assign w10080 = (~w6381 & w7782) | (~w6381 & w2880) | (w7782 & w2880);
assign w10081 = ~w2951 & ~w2751;
assign w10082 = b118 & a118;
assign w10083 = ~w12509 & ~w13428;
assign w10084 = (w1085 & w2511) | (w1085 & w12430) | (w2511 & w12430);
assign w10085 = w1881 & w5352;
assign w10086 = (w3334 & w14355) | (w3334 & ~w11516) | (w14355 & ~w11516);
assign w10087 = w14504 & w14486;
assign w10088 = (~w9921 & ~w1840) | (~w9921 & w9238) | (~w1840 & w9238);
assign w10089 = ~w10658 & w11812;
assign w10090 = ~w1649 & w13894;
assign w10091 = (~w12727 & ~w1402) | (~w12727 & w5149) | (~w1402 & w5149);
assign w10092 = ~w7450 & w6766;
assign w10093 = w750 & w1540;
assign w10094 = w6301 & ~w9170;
assign w10095 = w3427 & w12642;
assign w10096 = (w7782 & w12117) | (w7782 & w232) | (w12117 & w232);
assign w10097 = (w10449 & w5324) | (w10449 & w996) | (w5324 & w996);
assign w10098 = (~w6889 & w11635) | (~w6889 & w5252) | (w11635 & w5252);
assign w10099 = (~w3044 & w8203) | (~w3044 & w7134) | (w8203 & w7134);
assign w10100 = w4372 & ~w11292;
assign w10101 = w4262 & ~w3675;
assign w10102 = ~w1166 & ~w2154;
assign w10103 = ~w142 & w2320;
assign w10104 = ~w13452 & w4361;
assign w10105 = w4725 & w3114;
assign w10106 = ~w7782 & w6487;
assign w10107 = ~w11412 & w4633;
assign w10108 = w14276 & w3904;
assign w10109 = (w3325 & w8769) | (w3325 & w9424) | (w8769 & w9424);
assign w10110 = (~w10778 & w5716) | (~w10778 & ~w6753) | (w5716 & ~w6753);
assign w10111 = ~w2500 & ~w3632;
assign w10112 = w6230 & w5364;
assign w10113 = w9748 & w3561;
assign w10114 = ~w1093 & ~w6191;
assign w10115 = (~w9707 & ~w14002) | (~w9707 & ~w2181) | (~w14002 & ~w2181);
assign w10116 = w5569 & w9170;
assign w10117 = ~w4607 & w6115;
assign w10118 = (~w14463 & w6865) | (~w14463 & w12281) | (w6865 & w12281);
assign w10119 = (~w309 & w10224) | (~w309 & w13470) | (w10224 & w13470);
assign w10120 = w12920 & ~w11126;
assign w10121 = ~w11544 & w6519;
assign w10122 = ~w451 & w4659;
assign w10123 = ~w5620 & ~w3067;
assign w10124 = ~w6755 & w12968;
assign w10125 = (w350 & w7838) | (w350 & w430) | (w7838 & w430);
assign w10126 = w1101 & ~w806;
assign w10127 = ~w855 & w585;
assign w10128 = ~w13959 & w2888;
assign w10129 = ~w13011 & w9451;
assign w10130 = w14395 & ~w1805;
assign w10131 = ~w9772 & w8083;
assign w10132 = w14286 & ~w2332;
assign w10133 = (~w8085 & w1166) | (~w8085 & w1977) | (w1166 & w1977);
assign w10134 = w8769 & ~w777;
assign w10135 = (~w7012 & w4200) | (~w7012 & w12083) | (w4200 & w12083);
assign w10136 = w7464 | w2593;
assign w10137 = w7486 & ~w7104;
assign w10138 = ~w6988 & ~w4227;
assign w10139 = ~w2628 & ~w7481;
assign w10140 = w7376 & ~w5741;
assign w10141 = w10089 & ~w8307;
assign w10142 = ~w13122 & w10972;
assign w10143 = ~w13713 & w14526;
assign w10144 = w1507 & w6230;
assign w10145 = w7906 & ~w8035;
assign w10146 = w13635 & w3023;
assign w10147 = ~w7836 & ~w10139;
assign w10148 = (~w14578 & w10595) | (~w14578 & w3240) | (w10595 & w3240);
assign w10149 = ~w11874 & ~w6777;
assign w10150 = w5040 & w4980;
assign w10151 = w1673 & ~w8779;
assign w10152 = ~w10339 & w3988;
assign w10153 = ~w12003 & w4727;
assign w10154 = w3211 & w14594;
assign w10155 = (w10123 & w10171) | (w10123 & w2919) | (w10171 & w2919);
assign w10156 = (w12764 & ~w14364) | (w12764 & w10983) | (~w14364 & w10983);
assign w10157 = ~w4158 & w11254;
assign w10158 = w3154 & w2945;
assign w10159 = ~w12240 & w852;
assign w10160 = (~w9454 & w8904) | (~w9454 & w4751) | (w8904 & w4751);
assign w10161 = w10669 & ~w3039;
assign w10162 = (~w4050 & w743) | (~w4050 & w10333) | (w743 & w10333);
assign w10163 = w5761 & ~w3887;
assign w10164 = (~w5556 & w183) | (~w5556 & w14395) | (w183 & w14395);
assign w10165 = ~w6113 & w1978;
assign w10166 = ~w1774 & ~w13033;
assign w10167 = (w3442 & w897) | (w3442 & ~w2287) | (w897 & ~w2287);
assign w10168 = (~w9305 & w8428) | (~w9305 & w6356) | (w8428 & w6356);
assign w10169 = (w1288 & ~w11385) | (w1288 & ~w13561) | (~w11385 & ~w13561);
assign w10170 = w8259 & w13544;
assign w10171 = (~w4050 & w3870) | (~w4050 & w1324) | (w3870 & w1324);
assign w10172 = (w12786 & w3347) | (w12786 & w13068) | (w3347 & w13068);
assign w10173 = w10247 & ~w10317;
assign w10174 = ~w3215 & w14504;
assign w10175 = ~w13143 & ~w7806;
assign w10176 = w5893 & w11129;
assign w10177 = ~w2553 & w11640;
assign w10178 = w11732 & ~w10225;
assign w10179 = w3958 & w1172;
assign w10180 = w10221 & ~w4322;
assign w10181 = ~w9661 & w9904;
assign w10182 = ~w8183 & ~w2433;
assign w10183 = w2307 & w227;
assign w10184 = ~w9087 & w11068;
assign w10185 = (w12398 & w5559) | (w12398 & w1290) | (w5559 & w1290);
assign w10186 = ~w2317 & w90;
assign w10187 = w1328 & ~w7848;
assign w10188 = w7373 & ~w12775;
assign w10189 = ~w4050 & w3703;
assign w10190 = ~w9816 & w321;
assign w10191 = ~w10334 & ~w5989;
assign w10192 = (w6500 & w5583) | (w6500 & w2345) | (w5583 & w2345);
assign w10193 = (w13685 & w3748) | (w13685 & w5499) | (w3748 & w5499);
assign w10194 = (~w806 & w10126) | (~w806 & w10079) | (w10126 & w10079);
assign w10195 = ~w8183 & ~w840;
assign w10196 = ~w14215 & ~w8171;
assign w10197 = w7722 & ~w803;
assign w10198 = ~w9722 & ~w10796;
assign w10199 = w12121 & ~w14523;
assign w10200 = (w2858 & ~w13892) | (w2858 & w7430) | (~w13892 & w7430);
assign w10201 = ~w11940 & w337;
assign w10202 = (w7578 & w8770) | (w7578 & w10318) | (w8770 & w10318);
assign w10203 = w1607 & w455;
assign w10204 = (w12170 & w5559) | (w12170 & w14635) | (w5559 & w14635);
assign w10205 = ~w4921 & w6283;
assign w10206 = w11751 & w8970;
assign w10207 = w5522 & ~w2701;
assign w10208 = (w1949 & ~w5852) | (w1949 & w14358) | (~w5852 & w14358);
assign w10209 = (w4580 & w14108) | (w4580 & ~w3885) | (w14108 & ~w3885);
assign w10210 = w3809 & w2318;
assign w10211 = (w1362 & w12729) | (w1362 & w8633) | (w12729 & w8633);
assign w10212 = ~w10486 & ~w5283;
assign w10213 = ~w11606 & ~w2605;
assign w10214 = (~w2948 & w7592) | (~w2948 & w6783) | (w7592 & w6783);
assign w10215 = w6281 & ~w8269;
assign w10216 = ~w9200 & ~w10866;
assign w10217 = ~w5141 & w2884;
assign w10218 = ~w6648 & ~w8601;
assign w10219 = w12868 & w1692;
assign w10220 = (~w10884 & w1377) | (~w10884 & w10085) | (w1377 & w10085);
assign w10221 = ~b98 & ~a98;
assign w10222 = (~b53 & w6506) | (~b53 & w5872) | (w6506 & w5872);
assign w10223 = (~w3036 & w813) | (~w3036 & w8879) | (w813 & w8879);
assign w10224 = ~w6542 & ~w10477;
assign w10225 = ~w13733 & ~w1387;
assign w10226 = ~w6266 & w1236;
assign w10227 = ~w6301 & ~w13820;
assign w10228 = ~w7772 & ~w9713;
assign w10229 = ~w11577 & ~w14312;
assign w10230 = (w12135 & ~w7630) | (w12135 & w1092) | (~w7630 & w1092);
assign w10231 = ~w10462 & w2408;
assign w10232 = (~w2 & w5996) | (~w2 & w9355) | (w5996 & w9355);
assign w10233 = (w8135 & w14416) | (w8135 & ~w6025) | (w14416 & ~w6025);
assign w10234 = w11169 & ~w6653;
assign w10235 = ~w3034 & ~w4752;
assign w10236 = w14302 & ~w13445;
assign w10237 = ~w11652 & ~w11739;
assign w10238 = (w6310 & w12154) | (w6310 & ~w13980) | (w12154 & ~w13980);
assign w10239 = (w10708 & w6708) | (w10708 & w363) | (w6708 & w363);
assign w10240 = (w10903 & w3197) | (w10903 & ~w4310) | (w3197 & ~w4310);
assign w10241 = ~w1423 & w13376;
assign w10242 = w7032 & w10472;
assign w10243 = ~w12341 & w1540;
assign w10244 = (~w302 & w3389) | (~w302 & w6400) | (w3389 & w6400);
assign w10245 = ~w7988 & w6137;
assign w10246 = w8849 & w8542;
assign w10247 = (~w2922 & w9838) | (~w2922 & w5221) | (w9838 & w5221);
assign w10248 = w8534 & w4006;
assign w10249 = (~w11385 & w2693) | (~w11385 & w4205) | (w2693 & w4205);
assign w10250 = w10019 & w9128;
assign w10251 = w11013 & ~w5761;
assign w10252 = w10523 & ~w3075;
assign w10253 = ~w254 & w13294;
assign w10254 = ~w10207 & ~w9650;
assign w10255 = ~w5607 & w7342;
assign w10256 = ~w12664 & w4133;
assign w10257 = ~w5998 & w1283;
assign w10258 = w1274 & w13516;
assign w10259 = ~w9247 & w12477;
assign w10260 = ~w14281 & ~w1260;
assign w10261 = (~w5615 & w10513) | (~w5615 & w4130) | (w10513 & w4130);
assign w10262 = ~w3119 & ~w4853;
assign w10263 = (w9607 & w10540) | (w9607 & w1944) | (w10540 & w1944);
assign w10264 = ~w9170 & w12708;
assign w10265 = ~w14526 & w3734;
assign w10266 = w4836 & ~w2850;
assign w10267 = w419 & ~w7796;
assign w10268 = (w514 & w186) | (w514 & w6687) | (w186 & w6687);
assign w10269 = ~w7782 & w3705;
assign w10270 = w10676 & w1096;
assign w10271 = ~w3137 & ~w11861;
assign w10272 = ~w5482 & ~w3054;
assign w10273 = w9170 & w3283;
assign w10274 = ~w13170 & ~w11605;
assign w10275 = w4981 & ~w77;
assign w10276 = (w7082 & w7553) | (w7082 & w9610) | (w7553 & w9610);
assign w10277 = ~w12868 & w9255;
assign w10278 = w610 & w2028;
assign w10279 = (w9012 & w12435) | (w9012 & w4967) | (w12435 & w4967);
assign w10280 = ~w11604 & w14573;
assign w10281 = w13780 & a53;
assign w10282 = ~w13588 & w11945;
assign w10283 = (w11902 & w4921) | (w11902 & w1296) | (w4921 & w1296);
assign w10284 = w8171 & w6281;
assign w10285 = w7683 & w162;
assign w10286 = (~w5741 & w500) | (~w5741 & w10379) | (w500 & w10379);
assign w10287 = w7993 & ~w5410;
assign w10288 = w878 & w6719;
assign w10289 = ~w14141 & w12243;
assign w10290 = w7962 & w10295;
assign w10291 = (w12460 & w11261) | (w12460 & w3086) | (w11261 & w3086);
assign w10292 = ~w12460 & ~w92;
assign w10293 = ~w14239 & ~w3630;
assign w10294 = (w10758 & w7826) | (w10758 & w3641) | (w7826 & w3641);
assign w10295 = ~w5860 & ~w10477;
assign w10296 = (w2535 & w7595) | (w2535 & w2287) | (w7595 & w2287);
assign w10297 = w6391 & ~w13620;
assign w10298 = w5521 & w8327;
assign w10299 = w1255 & ~w1796;
assign w10300 = (~w9480 & w3727) | (~w9480 & w8619) | (w3727 & w8619);
assign w10301 = ~w13682 & ~w10116;
assign w10302 = ~w535 & w2446;
assign w10303 = (w10711 & w4582) | (w10711 & w2167) | (w4582 & w2167);
assign w10304 = w5803 & w5105;
assign w10305 = (~w5761 & w8912) | (~w5761 & w6528) | (w8912 & w6528);
assign w10306 = ~w12217 & w13452;
assign w10307 = (~w5952 & w2918) | (~w5952 & w1394) | (w2918 & w1394);
assign w10308 = w6871 & w8539;
assign w10309 = b34 & a34;
assign w10310 = (~w12528 & ~w3383) | (~w12528 & w3721) | (~w3383 & w3721);
assign w10311 = ~w12094 & w9560;
assign w10312 = w1494 & w2698;
assign w10313 = w5243 & w2599;
assign w10314 = (~w4679 & w5346) | (~w4679 & w6038) | (w5346 & w6038);
assign w10315 = w1063 & w13304;
assign w10316 = ~w12240 & w10997;
assign w10317 = ~w1821 & ~w10507;
assign w10318 = (w2445 & w9798) | (w2445 & w2823) | (w9798 & w2823);
assign w10319 = w1166 & w10546;
assign w10320 = ~w1107 & ~w7688;
assign w10321 = ~w5502 & w3713;
assign w10322 = ~w11401 & w10806;
assign w10323 = ~w9070 & ~w313;
assign w10324 = ~w7681 & ~w13344;
assign w10325 = (~w13462 & w5358) | (~w13462 & w2224) | (w5358 & w2224);
assign w10326 = ~w13251 & w5109;
assign w10327 = ~w14302 & w473;
assign w10328 = ~w13756 & w2965;
assign w10329 = (w9663 & w2520) | (w9663 & w3095) | (w2520 & w3095);
assign w10330 = w7401 & ~w1158;
assign w10331 = ~w1096 & ~w1642;
assign w10332 = w5867 & w12823;
assign w10333 = w10708 & ~w14464;
assign w10334 = ~w12371 & ~w4700;
assign w10335 = ~w13713 & ~w4287;
assign w10336 = w9840 & w6679;
assign w10337 = w12615 & ~w11756;
assign w10338 = w1503 & w8745;
assign w10339 = b15 & a15;
assign w10340 = (w14254 & w4149) | (w14254 & w1457) | (w4149 & w1457);
assign w10341 = ~w11699 | ~w11399;
assign w10342 = ~w12948 & ~w11366;
assign w10343 = ~w1266 & ~w3363;
assign w10344 = w5505 & ~w10917;
assign w10345 = (w1362 & w5239) | (w1362 & w6411) | (w5239 & w6411);
assign w10346 = ~w1177 & ~w12196;
assign w10347 = w13282 & w7561;
assign w10348 = w9156 & w6888;
assign w10349 = w8459 & ~w7554;
assign w10350 = w14137 & ~w7754;
assign w10351 = w13282 & ~w13206;
assign w10352 = w7857 & ~w7978;
assign w10353 = (w12774 & ~w6787) | (w12774 & ~w13270) | (~w6787 & ~w13270);
assign w10354 = b123 & a123;
assign w10355 = (~w8636 & w7979) | (~w8636 & w5880) | (w7979 & w5880);
assign w10356 = w14344 & w12127;
assign w10357 = w9921 & ~w6716;
assign w10358 = ~w12087 & w5586;
assign w10359 = ~w254 & w14224;
assign w10360 = ~w6888 & w9541;
assign w10361 = ~w8110 & ~w13839;
assign w10362 = ~w12483 & ~w8269;
assign w10363 = ~w4312 & ~w14512;
assign w10364 = (w9748 & w12891) | (w9748 & w11468) | (w12891 & w11468);
assign w10365 = (w13732 & w9544) | (w13732 & w8505) | (w9544 & w8505);
assign w10366 = ~w2938 & w6041;
assign w10367 = (w12406 & w5990) | (w12406 & w3918) | (w5990 & w3918);
assign w10368 = w4989 & ~w14390;
assign w10369 = (w1293 & w4717) | (w1293 & w7389) | (w4717 & w7389);
assign w10370 = (w5497 & w14402) | (w5497 & w4054) | (w14402 & w4054);
assign w10371 = w2549 & w3861;
assign w10372 = w4253 & w13527;
assign w10373 = w1942 & w9547;
assign w10374 = ~w1172 & ~w13820;
assign w10375 = w13423 & ~w13306;
assign w10376 = ~w217 & ~w2941;
assign w10377 = w2762 & w3904;
assign w10378 = w36 & w5605;
assign w10379 = ~w5741 & w8110;
assign w10380 = w5273 & w11770;
assign w10381 = ~w9362 & w8950;
assign w10382 = w5950 & w6714;
assign w10383 = w9429 & w4353;
assign w10384 = (w2105 & w7140) | (w2105 & w11819) | (w7140 & w11819);
assign w10385 = ~w3067 & w8632;
assign w10386 = ~w12662 & ~w14395;
assign w10387 = ~w1873 & w13969;
assign w10388 = ~w10523 & ~w13839;
assign w10389 = ~w13916 & ~w5852;
assign w10390 = ~w11500 & w95;
assign w10391 = w1098 & ~w12997;
assign w10392 = (w13219 & w13380) | (w13219 & w13440) | (w13380 & w13440);
assign w10393 = w11500 & w2425;
assign w10394 = ~w6258 & ~w8992;
assign w10395 = w11117 & w3603;
assign w10396 = ~w5178 & ~w1842;
assign w10397 = w8325 & ~w9719;
assign w10398 = ~w3113 & ~w4059;
assign w10399 = ~w12621 & ~w9263;
assign w10400 = (~w1842 & w7782) | (~w1842 & w4990) | (w7782 & w4990);
assign w10401 = w10123 & ~w2285;
assign w10402 = (w8408 & w8583) | (w8408 & w13931) | (w8583 & w13931);
assign w10403 = w11371 & w4973;
assign w10404 = ~w7488 & w5846;
assign w10405 = (w5794 & w4756) | (w5794 & w9773) | (w4756 & w9773);
assign w10406 = (~w2379 & ~w13457) | (~w2379 & w3658) | (~w13457 & w3658);
assign w10407 = (w9328 & ~w4815) | (w9328 & w9651) | (~w4815 & w9651);
assign w10408 = b23 & a23;
assign w10409 = ~w8171 & w7085;
assign w10410 = ~w199 & w3526;
assign w10411 = (w3906 & w10462) | (w3906 & w4661) | (w10462 & w4661);
assign w10412 = ~w12489 & ~w5960;
assign w10413 = (w6486 & w9450) | (w6486 & ~w13292) | (w9450 & ~w13292);
assign w10414 = (~w8362 & w9012) | (~w8362 & w7604) | (w9012 & w7604);
assign w10415 = ~w4032 & w13531;
assign w10416 = (~w408 & w3865) | (~w408 & w8939) | (w3865 & w8939);
assign w10417 = ~w7376 & w3215;
assign w10418 = w8886 & ~w2811;
assign w10419 = ~w13959 & w3443;
assign w10420 = (w9547 & ~w11996) | (w9547 & w10373) | (~w11996 & w10373);
assign w10421 = w10748 & w12315;
assign w10422 = w12269 & w9214;
assign w10423 = (~w12398 & w14178) | (~w12398 & w6048) | (w14178 & w6048);
assign w10424 = w4407 & a53;
assign w10425 = (w11031 & w9403) | (w11031 & w10999) | (w9403 & w10999);
assign w10426 = ~w125 & ~w4483;
assign w10427 = ~w13321 & w8732;
assign w10428 = w8909 & ~w14040;
assign w10429 = ~w2470 & w1032;
assign w10430 = (~w803 & ~w13620) | (~w803 & w11618) | (~w13620 & w11618);
assign w10431 = ~w9927 & ~w14588;
assign w10432 = (w12569 & ~w7051) | (w12569 & w3007) | (~w7051 & w3007);
assign w10433 = (~w8370 & w278) | (~w8370 & w14122) | (w278 & w14122);
assign w10434 = w13201 & ~w10370;
assign w10435 = w13916 & ~w4716;
assign w10436 = (~w8975 & ~w7630) | (~w8975 & w123) | (~w7630 & w123);
assign w10437 = ~w8128 & ~w8946;
assign w10438 = ~w13462 & w5866;
assign w10439 = w5613 & w7283;
assign w10440 = ~w142 & ~w9296;
assign w10441 = w9809 & ~w5681;
assign w10442 = ~w8807 & ~w9956;
assign w10443 = (~w13008 & w9506) | (~w13008 & w5620) | (w9506 & w5620);
assign w10444 = (w12893 & ~w1140) | (w12893 & w3358) | (~w1140 & w3358);
assign w10445 = ~w14302 & w13733;
assign w10446 = w2337 & w860;
assign w10447 = ~w10435 & w8853;
assign w10448 = ~w6080 & ~w11861;
assign w10449 = (~w2261 & w10433) | (~w2261 & w9519) | (w10433 & w9519);
assign w10450 = w11212 & w11035;
assign w10451 = ~w7790 & w1674;
assign w10452 = (~w9087 & w9608) | (~w9087 & w9899) | (w9608 & w9899);
assign w10453 = w10526 & ~w3194;
assign w10454 = ~w10334 & ~w1598;
assign w10455 = ~w10757 & ~w10699;
assign w10456 = (w14028 & w2541) | (w14028 & w13486) | (w2541 & w13486);
assign w10457 = (w3372 & w11370) | (w3372 & w13195) | (w11370 & w13195);
assign w10458 = (w4454 & w14587) | (w4454 & ~w2670) | (w14587 & ~w2670);
assign w10459 = w9525 & w10744;
assign w10460 = ~w11479 & w13624;
assign w10461 = w11013 & ~w2729;
assign w10462 = w2194 & ~w6418;
assign w10463 = b53 & ~w12121;
assign w10464 = w1332 & w9679;
assign w10465 = w10035 & w227;
assign w10466 = (w13461 & w8355) | (w13461 & w12112) | (w8355 & w12112);
assign w10467 = w10514 & w8584;
assign w10468 = ~b53 & ~w7872;
assign w10469 = ~w1638 & w11087;
assign w10470 = ~w6689 & ~w1483;
assign w10471 = w13095 & w14430;
assign w10472 = (w3592 & w12590) | (w3592 & w10101) | (w12590 & w10101);
assign w10473 = (~w3550 & w12847) | (~w3550 & w1058) | (w12847 & w1058);
assign w10474 = w5522 & w7670;
assign w10475 = w4487 & w8984;
assign w10476 = w1418 & w606;
assign w10477 = ~b60 & ~a60;
assign w10478 = w7267 & w9901;
assign w10479 = (w4855 & ~w12240) | (w4855 & w14342) | (~w12240 & w14342);
assign w10480 = w7786 & ~w5623;
assign w10481 = ~w11847 & ~w11626;
assign w10482 = ~w3096 & w1509;
assign w10483 = ~w5836 & ~w6794;
assign w10484 = (~w4099 & w2470) | (~w4099 & w4895) | (w2470 & w4895);
assign w10485 = ~w14163 & ~w9758;
assign w10486 = ~w13423 & w7295;
assign w10487 = w1555 & ~w10962;
assign w10488 = w8101 & w1232;
assign w10489 = w2656 & ~w2858;
assign w10490 = ~w7244 & ~w7670;
assign w10491 = w9647 & w10612;
assign w10492 = (w1805 & w13222) | (w1805 & w1042) | (w13222 & w1042);
assign w10493 = w1607 & ~w12564;
assign w10494 = ~a117 & ~w7244;
assign w10495 = (~w10719 & w7225) | (~w10719 & w2062) | (w7225 & w2062);
assign w10496 = w3507 & w11093;
assign w10497 = (w13685 & w9825) | (w13685 & w425) | (w9825 & w425);
assign w10498 = w10119 & ~w11488;
assign w10499 = ~w2490 & w2140;
assign w10500 = ~w7108 & w4760;
assign w10501 = w8964 & ~w11520;
assign w10502 = (~w4032 & w1655) | (~w4032 & w9692) | (w1655 & w9692);
assign w10503 = ~w2680 & ~w9366;
assign w10504 = ~w2509 & ~w11013;
assign w10505 = ~w987 & w13775;
assign w10506 = (w10290 & w9748) | (w10290 & w11686) | (w9748 & w11686);
assign w10507 = ~w8328 & ~w3219;
assign w10508 = w10676 & w3215;
assign w10509 = ~w8370 & ~w10339;
assign w10510 = (w2116 & w6545) | (w2116 & w6434) | (w6545 & w6434);
assign w10511 = ~w11462 & w6500;
assign w10512 = (w4599 & w2488) | (w4599 & w11283) | (w2488 & w11283);
assign w10513 = w5602 | w3957;
assign w10514 = ~w1096 & ~w2933;
assign w10515 = ~w8032 & w5865;
assign w10516 = (w11416 & w14508) | (w11416 & w11503) | (w14508 & w11503);
assign w10517 = ~b100 & ~a100;
assign w10518 = w1036 & w2492;
assign w10519 = w706 & w5282;
assign w10520 = (~w1663 & w4027) | (~w1663 & w10303) | (w4027 & w10303);
assign w10521 = ~w9717 & ~w669;
assign w10522 = (w829 & w2144) | (w829 & w6422) | (w2144 & w6422);
assign w10523 = b46 & a46;
assign w10524 = ~w10245 & w10157;
assign w10525 = (w11803 & w13712) | (w11803 & w4249) | (w13712 & w4249);
assign w10526 = ~w5761 & w1800;
assign w10527 = (w9510 & w5119) | (w9510 & ~w11915) | (w5119 & ~w11915);
assign w10528 = (w5491 & w6848) | (w5491 & w217) | (w6848 & w217);
assign w10529 = (~w1540 & ~w13981) | (~w1540 & w4022) | (~w13981 & w4022);
assign w10530 = ~w3536 & w7824;
assign w10531 = w5237 & ~w5972;
assign w10532 = ~w14227 & w1274;
assign w10533 = w92 & w9378;
assign w10534 = w7752 & ~w9594;
assign w10535 = (w13685 & w2183) | (w13685 & w6982) | (w2183 & w6982);
assign w10536 = (~w2492 & w4847) | (~w2492 & w4609) | (w4847 & w4609);
assign w10537 = w12460 & w8513;
assign w10538 = w12065 & ~w5406;
assign w10539 = w7365 & ~w5664;
assign w10540 = ~w8742 & ~w9672;
assign w10541 = w5348 & w3904;
assign w10542 = (w10551 & w13349) | (w10551 & w5171) | (w13349 & w5171);
assign w10543 = ~w14302 & w9244;
assign w10544 = ~w7605 & ~w504;
assign w10545 = ~w3759 & ~w7447;
assign w10546 = ~w8085 & ~w3502;
assign w10547 = ~w10431 & w6689;
assign w10548 = ~w2974 & w10098;
assign w10549 = (w6802 & w250) | (w6802 & w3477) | (w250 & w3477);
assign w10550 = w6446 & ~w6404;
assign w10551 = w9284 & w6436;
assign w10552 = ~w5490 & ~w14055;
assign w10553 = (w9541 & w12851) | (w9541 & w8952) | (w12851 & w8952);
assign w10554 = w9306 & w3037;
assign w10555 = ~w6759 & ~w3697;
assign w10556 = ~w5761 & ~w11745;
assign w10557 = ~w1919 & w1171;
assign w10558 = w5081 & w1315;
assign w10559 = w5744 & w10386;
assign w10560 = ~w10015 & ~w5666;
assign w10561 = (w6886 & ~w1007) | (w6886 & w6877) | (~w1007 & w6877);
assign w10562 = ~w4645 & ~w3107;
assign w10563 = ~w9564 & w12821;
assign w10564 = ~w7765 & ~w13997;
assign w10565 = w1599 & w728;
assign w10566 = ~w10056 & w7798;
assign w10567 = w4564 & ~w4125;
assign w10568 = w2485 & w5825;
assign w10569 = w4472 & ~w8992;
assign w10570 = ~w4481 & ~w3668;
assign w10571 = w10907 & w4075;
assign w10572 = w7670 & w8475;
assign w10573 = ~w10256 & w8133;
assign w10574 = w11761 & w2301;
assign w10575 = ~w4512 & w12612;
assign w10576 = (~w6377 & w5943) | (~w6377 & w4430) | (w5943 & w4430);
assign w10577 = (w7302 & w1454) | (w7302 & w12537) | (w1454 & w12537);
assign w10578 = (w6276 & w1153) | (w6276 & w9325) | (w1153 & w9325);
assign w10579 = w2452 & ~w5094;
assign w10580 = (w1457 & w236) | (w1457 & w7999) | (w236 & w7999);
assign w10581 = (~w4627 & w7545) | (~w4627 & ~w3300) | (w7545 & ~w3300);
assign w10582 = w3914 & w5932;
assign w10583 = (w13059 & w12544) | (w13059 & w8434) | (w12544 & w8434);
assign w10584 = ~w9903 & ~w1632;
assign w10585 = w7022 & w4515;
assign w10586 = w7786 & ~w10973;
assign w10587 = (w6502 & ~w4032) | (w6502 & w6322) | (~w4032 & w6322);
assign w10588 = ~w10358 & w6434;
assign w10589 = ~w9320 & w453;
assign w10590 = w10880 & w5593;
assign w10591 = (w7493 & w4921) | (w7493 & w14142) | (w4921 & w14142);
assign w10592 = ~w2855 & ~w14393;
assign w10593 = (w5952 & w11422) | (w5952 & w1872) | (w11422 & w1872);
assign w10594 = (w2655 & w8284) | (w2655 & w10296) | (w8284 & w10296);
assign w10595 = ~w9713 & ~w10812;
assign w10596 = ~w14215 & w4182;
assign w10597 = w8872 & w645;
assign w10598 = (w5776 & w2797) | (w5776 & w12376) | (w2797 & w12376);
assign w10599 = (w9340 & ~w12269) | (w9340 & w4409) | (~w12269 & w4409);
assign w10600 = (~w5732 & ~w7168) | (~w5732 & w3782) | (~w7168 & w3782);
assign w10601 = w3288 & ~w4458;
assign w10602 = (w8742 & w14664) | (w8742 & w12700) | (w14664 & w12700);
assign w10603 = ~w12642 & ~w6105;
assign w10604 = ~w1346 & ~w8224;
assign w10605 = ~w12398 & ~w9015;
assign w10606 = (w11718 & w2257) | (w11718 & w10952) | (w2257 & w10952);
assign w10607 = ~w3502 & w12398;
assign w10608 = w3914 & ~w9227;
assign w10609 = (~w3019 & w11443) | (~w3019 & ~w14526) | (w11443 & ~w14526);
assign w10610 = w8967 & w3671;
assign w10611 = w6301 & ~w6700;
assign w10612 = ~w12413 & ~w7404;
assign w10613 = w1503 & ~w4030;
assign w10614 = (w11429 & w6015) | (w11429 & w4720) | (w6015 & w4720);
assign w10615 = (~w9336 & ~w6591) | (~w9336 & w4163) | (~w6591 & w4163);
assign w10616 = ~w9725 & ~w1073;
assign w10617 = ~w12240 & w4441;
assign w10618 = ~w11462 & ~w3159;
assign w10619 = ~w9284 & w13839;
assign w10620 = ~w2218 & w3390;
assign w10621 = ~w8827 & ~w14430;
assign w10622 = w13953 & w7914;
assign w10623 = w13496 & w9454;
assign w10624 = w6562 & ~w12650;
assign w10625 = ~w8110 & w500;
assign w10626 = ~w8513 & ~w11902;
assign w10627 = ~w1785 & w9019;
assign w10628 = (w2194 & w12531) | (w2194 & w12499) | (w12531 & w12499);
assign w10629 = (~w3508 & w1229) | (~w3508 & w5398) | (w1229 & w5398);
assign w10630 = (~w6219 & ~w4520) | (~w6219 & ~w5768) | (~w4520 & ~w5768);
assign w10631 = ~w6513 & w1887;
assign w10632 = ~w2762 & ~w996;
assign w10633 = (w3778 & w11731) | (w3778 & w11844) | (w11731 & w11844);
assign w10634 = (w12952 & w9174) | (w12952 & ~w12638) | (w9174 & ~w12638);
assign w10635 = w3364 & ~w2673;
assign w10636 = w3601 & w13932;
assign w10637 = w10500 & w179;
assign w10638 = w7020 & w11044;
assign w10639 = (w1362 & w14427) | (w1362 & w9775) | (w14427 & w9775);
assign w10640 = w11031 & w147;
assign w10641 = ~w4739 & ~w10649;
assign w10642 = ~w5294 & w10075;
assign w10643 = ~w5522 & w3727;
assign w10644 = (w8827 & w10245) | (w8827 & w9048) | (w10245 & w9048);
assign w10645 = ~w6135 & ~w6080;
assign w10646 = ~w2317 & w11315;
assign w10647 = ~w12893 & w14486;
assign w10648 = w636 & w3727;
assign w10649 = (w1545 & w11848) | (w1545 & w4220) | (w11848 & w4220);
assign w10650 = w2261 & w7362;
assign w10651 = (w4855 & w11067) | (w4855 & w8176) | (w11067 & w8176);
assign w10652 = w9375 & ~w13282;
assign w10653 = w10439 & w128;
assign w10654 = (w11810 & w12499) | (w11810 & w12503) | (w12499 & w12503);
assign w10655 = w4786 & ~w7630;
assign w10656 = w2926 & ~w6514;
assign w10657 = ~w1474 & w7670;
assign w10658 = ~w6408 & w6781;
assign w10659 = ~w5712 & ~w13676;
assign w10660 = ~w9715 & ~w3209;
assign w10661 = ~w11148 & w1834;
assign w10662 = w739 & ~w9251;
assign w10663 = (w13086 & ~w17) | (w13086 & w1429) | (~w17 & w1429);
assign w10664 = (~w9244 & w12574) | (~w9244 & w4288) | (w12574 & w4288);
assign w10665 = ~w2108 & ~w10144;
assign w10666 = ~w2500 & w1821;
assign w10667 = w13282 & w6572;
assign w10668 = ~w14227 & ~w10075;
assign w10669 = (~w5732 & w12321) | (~w5732 & w9888) | (w12321 & w9888);
assign w10670 = w1710 & w565;
assign w10671 = ~w2279 & ~w10590;
assign w10672 = w10045 & w7914;
assign w10673 = w10676 & w9200;
assign w10674 = ~w1898 & w12696;
assign w10675 = ~b88 & ~a88;
assign w10676 = ~w9823 & ~w14135;
assign w10677 = (~w7057 & w11333) | (~w7057 & w12020) | (w11333 & w12020);
assign w10678 = ~w10150 & w12910;
assign w10679 = ~w10245 & w3644;
assign w10680 = ~w4607 & w11107;
assign w10681 = ~w5852 & w2820;
assign w10682 = ~w12065 & w10669;
assign w10683 = w13857 & w12311;
assign w10684 = (w13572 & w14422) | (w13572 & w946) | (w14422 & w946);
assign w10685 = (w9096 & w5356) | (w9096 & w14029) | (w5356 & w14029);
assign w10686 = w3957 & w10943;
assign w10687 = (w14439 & w2666) | (w14439 & w8634) | (w2666 & w8634);
assign w10688 = ~w7654 & w3225;
assign w10689 = ~w803 & ~w12170;
assign w10690 = (~w5579 & ~w11429) | (~w5579 & w4735) | (~w11429 & w4735);
assign w10691 = ~w12604 & ~w7889;
assign w10692 = ~w6583 & ~w8768;
assign w10693 = (~w7296 & ~w183) | (~w7296 & w6161) | (~w183 & w6161);
assign w10694 = w1712 & ~w7950;
assign w10695 = ~w2656 & ~w4099;
assign w10696 = (~w5005 & w13349) | (~w5005 & w6157) | (w13349 & w6157);
assign w10697 = ~w3799 & w12411;
assign w10698 = (w608 & w10462) | (w608 & w13032) | (w10462 & w13032);
assign w10699 = ~w10757 & ~w2509;
assign w10700 = w5471 & w11158;
assign w10701 = (w6598 & w5396) | (w6598 & ~w5901) | (w5396 & ~w5901);
assign w10702 = ~w10042 & ~w8285;
assign w10703 = ~w12604 & ~w6689;
assign w10704 = b55 & a55;
assign w10705 = w4836 & w12398;
assign w10706 = w57 & w13131;
assign w10707 = (~w7630 & w7770) | (~w7630 & w7939) | (w7770 & w7939);
assign w10708 = w10689 & w12656;
assign w10709 = w12538 & ~w7239;
assign w10710 = ~w4255 & w8473;
assign w10711 = w3248 & w8451;
assign w10712 = w14286 & w654;
assign w10713 = ~w10082 & ~w660;
assign w10714 = ~w1015 & ~w7999;
assign w10715 = (w10773 & w613) | (w10773 & w7417) | (w613 & w7417);
assign w10716 = ~w13562 & w5282;
assign w10717 = (w3039 & w10676) | (w3039 & w7324) | (w10676 & w7324);
assign w10718 = w10255 & w3752;
assign w10719 = w768 & ~w10711;
assign w10720 = w11177 & w2881;
assign w10721 = ~w2774 & ~w14632;
assign w10722 = b4 & a4;
assign w10723 = w6427 & ~w4081;
assign w10724 = w10061 & w7123;
assign w10725 = ~w9715 & w11488;
assign w10726 = w4952 | ~w13306;
assign w10727 = (~w9525 & w783) | (~w9525 & w9462) | (w783 & w9462);
assign w10728 = ~w142 & w13713;
assign w10729 = w8926 & w1582;
assign w10730 = ~w7681 & ~w4501;
assign w10731 = w8389 & ~w10096;
assign w10732 = w7463 & ~w12266;
assign w10733 = w3435 & w8080;
assign w10734 = w25 & ~w12661;
assign w10735 = ~w922 & ~w12669;
assign w10736 = w347 & w3682;
assign w10737 = (w1362 & w4726) | (w1362 & w11094) | (w4726 & w11094);
assign w10738 = (~w7477 & w5699) | (~w7477 & w9391) | (w5699 & w9391);
assign w10739 = (w7911 & w5376) | (w7911 & w10287) | (w5376 & w10287);
assign w10740 = (~w4363 & w2645) | (~w4363 & w3344) | (w2645 & w3344);
assign w10741 = (w12575 & w1510) | (w12575 & w7956) | (w1510 & w7956);
assign w10742 = (w12460 & w2935) | (w12460 & w11771) | (w2935 & w11771);
assign w10743 = w3209 & w1264;
assign w10744 = (~w11429 & w9821) | (~w11429 & w11082) | (w9821 & w11082);
assign w10745 = (w7811 & w6240) | (w7811 & ~w3209) | (w6240 & ~w3209);
assign w10746 = (~w8667 & ~w11916) | (~w8667 & w424) | (~w11916 & w424);
assign w10747 = (w4545 & w5346) | (w4545 & w6842) | (w5346 & w6842);
assign w10748 = ~w657 & w5390;
assign w10749 = ~w13189 & w10699;
assign w10750 = w1274 & ~w6889;
assign w10751 = ~w8857 & w11901;
assign w10752 = ~w8937 & w5049;
assign w10753 = ~w922 & w6700;
assign w10754 = w13854 & ~w803;
assign w10755 = ~w7488 & w14554;
assign w10756 = (w3020 & w9322) | (w3020 & w8157) | (w9322 & w8157);
assign w10757 = b115 & a115;
assign w10758 = (~w11606 & w10213) | (~w11606 & ~w4756) | (w10213 & ~w4756);
assign w10759 = (w10625 & w11149) | (w10625 & ~w9534) | (w11149 & ~w9534);
assign w10760 = (w9170 & w13284) | (w9170 & w12726) | (w13284 & w12726);
assign w10761 = w3036 & w5845;
assign w10762 = (~w10245 & w5847) | (~w10245 & w11678) | (w5847 & w11678);
assign w10763 = w1764 & ~w9929;
assign w10764 = ~w1997 & w13008;
assign w10765 = w3384 & w12454;
assign w10766 = w2606 & w11677;
assign w10767 = (w10486 & w749) | (w10486 & ~w6536) | (w749 & ~w6536);
assign w10768 = w3690 & w6551;
assign w10769 = ~w9858 & w10530;
assign w10770 = w4213 & w11902;
assign w10771 = w1840 & w4359;
assign w10772 = ~w14058 & w9024;
assign w10773 = ~w14291 & w873;
assign w10774 = (~w6795 & w14664) | (~w6795 & w11435) | (w14664 & w11435);
assign w10775 = ~w6360 & ~w3382;
assign w10776 = w10265 & w3734;
assign w10777 = w6623 | ~w7684;
assign w10778 = w2698 & w6381;
assign w10779 = ~w9794 & ~w9298;
assign w10780 = (~w9010 & w96) | (~w9010 & w6508) | (w96 & w6508);
assign w10781 = (~w11361 & w5946) | (~w11361 & w12791) | (w5946 & w12791);
assign w10782 = w13978 & ~w892;
assign w10783 = (~w13219 & w4562) | (~w13219 & w12815) | (w4562 & w12815);
assign w10784 = w10221 & ~w1062;
assign w10785 = (w13587 & w6576) | (w13587 & w12838) | (w6576 & w12838);
assign w10786 = w1821 & ~w5664;
assign w10787 = w4953 & w11053;
assign w10788 = (w14463 & w4468) | (w14463 & w10684) | (w4468 & w10684);
assign w10789 = w2519 & w1585;
assign w10790 = w13013 & ~w3814;
assign w10791 = ~w6758 & ~w2033;
assign w10792 = ~w11440 & w7035;
assign w10793 = w8745 & w5730;
assign w10794 = w3963 & w10562;
assign w10795 = ~w14248 & ~w13680;
assign w10796 = ~w10245 & w925;
assign w10797 = (w93 & w12527) | (w93 & w12154) | (w12527 & w12154);
assign w10798 = (w3550 & w11824) | (w3550 & w3189) | (w11824 & w3189);
assign w10799 = (w4325 & w10937) | (w4325 & w4320) | (w10937 & w4320);
assign w10800 = (~w10514 & ~w3914) | (~w10514 & w5068) | (~w3914 & w5068);
assign w10801 = (w11870 & w11206) | (w11870 & w12154) | (w11206 & w12154);
assign w10802 = w8871 & w2701;
assign w10803 = (w1773 & w389) | (w1773 & w12376) | (w389 & w12376);
assign w10804 = w3157 & ~w3928;
assign w10805 = w3081 & w9572;
assign w10806 = w10290 & w740;
assign w10807 = w13191 & w11380;
assign w10808 = (w690 & ~w9708) | (w690 & w7410) | (~w9708 & w7410);
assign w10809 = w7794 & ~w13448;
assign w10810 = (w2700 & w7167) | (w2700 & ~w5370) | (w7167 & ~w5370);
assign w10811 = ~w6163 & ~w2956;
assign w10812 = w7772 & w2236;
assign w10813 = ~w8100 & w821;
assign w10814 = (~w4756 & w1868) | (~w4756 & w12597) | (w1868 & w12597);
assign w10815 = (w5026 & w7894) | (w5026 & w6537) | (w7894 & w6537);
assign w10816 = (w7515 & w4613) | (w7515 & w12336) | (w4613 & w12336);
assign w10817 = w4796 & ~w12970;
assign w10818 = w12543 & ~w12828;
assign w10819 = ~w8561 & ~w7808;
assign w10820 = a127 & b127;
assign w10821 = ~w12559 & w227;
assign w10822 = ~w14283 & ~w745;
assign w10823 = (~w5971 & ~w1362) | (~w5971 & w10414) | (~w1362 & w10414);
assign w10824 = ~b4 & ~a4;
assign w10825 = w13222 & w5225;
assign w10826 = w9511 & ~w6812;
assign w10827 = w7305 & w5282;
assign w10828 = ~w7296 & w5490;
assign w10829 = w305 & ~w2346;
assign w10830 = w13501 & ~w10292;
assign w10831 = ~w10283 & w474;
assign w10832 = (w2928 & ~w13960) | (w2928 & w4763) | (~w13960 & w4763);
assign w10833 = ~w2500 & w4299;
assign w10834 = ~w10119 & ~w8992;
assign w10835 = w968 & ~w4553;
assign w10836 = ~w6799 & ~w788;
assign w10837 = ~w13924 & w13191;
assign w10838 = w972 & ~w934;
assign w10839 = (~w9170 & w1712) | (~w9170 & w10094) | (w1712 & w10094);
assign w10840 = ~w8380 & ~w9880;
assign w10841 = ~w9284 & ~w5577;
assign w10842 = ~w1653 & ~w12335;
assign w10843 = (w13932 & w3601) | (w13932 & w12376) | (w3601 & w12376);
assign w10844 = (w5662 & w2810) | (w5662 & w8903) | (w2810 & w8903);
assign w10845 = (w2204 & ~w1405) | (w2204 & w3534) | (~w1405 & w3534);
assign w10846 = ~w14015 & w11861;
assign w10847 = ~w3982 & w13872;
assign w10848 = ~w8958 & ~w6381;
assign w10849 = w1062 & w13914;
assign w10850 = w10439 & w7241;
assign w10851 = ~w1802 & ~w8475;
assign w10852 = w12609 & ~w13763;
assign w10853 = ~w4359 & ~w9338;
assign w10854 = w1838 & ~w5761;
assign w10855 = ~w9015 & ~w852;
assign w10856 = w13209 & w11300;
assign w10857 = w8110 & ~w6500;
assign w10858 = (~w7082 & w6327) | (~w7082 & w1662) | (w6327 & w1662);
assign w10859 = w2656 & w4473;
assign w10860 = ~w2061 & w2930;
assign w10861 = ~w2218 & w12304;
assign w10862 = (w3904 & w300) | (w3904 & w5503) | (w300 & w5503);
assign w10863 = w2608 & w9065;
assign w10864 = ~w13101 & ~w7173;
assign w10865 = ~w6043 & ~w8756;
assign w10866 = w10872 & ~w5301;
assign w10867 = w13604 & w792;
assign w10868 = ~w10265 & ~w40;
assign w10869 = w607 & ~w7670;
assign w10870 = ~w71 & w10879;
assign w10871 = w14664 & w2289;
assign w10872 = ~w13713 & ~w8754;
assign w10873 = (~w10778 & w5716) | (~w10778 & w7047) | (w5716 & w7047);
assign w10874 = w7772 & ~w7630;
assign w10875 = ~w1642 & ~w4806;
assign w10876 = w11309 & ~w3840;
assign w10877 = ~w7663 & w1378;
assign w10878 = (w1704 & w13859) | (w1704 & ~w5476) | (w13859 & ~w5476);
assign w10879 = w5177 & ~w3435;
assign w10880 = ~w2291 & ~w9583;
assign w10881 = (w10923 & w1060) | (w10923 & w7540) | (w1060 & w7540);
assign w10882 = w1283 & w12087;
assign w10883 = ~w3131 & ~w11269;
assign w10884 = ~w11362 & ~w14273;
assign w10885 = ~w8679 & ~w14120;
assign w10886 = w8918 & w5845;
assign w10887 = (~w7709 & w5139) | (~w7709 & w6644) | (w5139 & w6644);
assign w10888 = ~w12237 & ~w1154;
assign w10889 = w11364 & ~w11376;
assign w10890 = (w7762 & w8464) | (w7762 & w1563) | (w8464 & w1563);
assign w10891 = (w4099 & w8571) | (w4099 & w1248) | (w8571 & w1248);
assign w10892 = ~w884 & w7455;
assign w10893 = (w3957 & w7475) | (w3957 & w10359) | (w7475 & w10359);
assign w10894 = (~w11416 & w2905) | (~w11416 & w12853) | (w2905 & w12853);
assign w10895 = ~w4700 & w9022;
assign w10896 = (w13700 & w540) | (w13700 & w13392) | (w540 & w13392);
assign w10897 = w12330 & ~w8626;
assign w10898 = ~w12872 & ~w12962;
assign w10899 = (~w3145 & w9666) | (~w3145 & w5010) | (w9666 & w5010);
assign w10900 = ~w1831 & w8746;
assign w10901 = w6813 & ~w2410;
assign w10902 = w12173 & ~w8263;
assign w10903 = ~w1760 & ~w4425;
assign w10904 = ~w6135 & w11934;
assign w10905 = (w3929 & w9221) | (w3929 & ~w9403) | (w9221 & ~w9403);
assign w10906 = w10941 & ~w10013;
assign w10907 = w10795 & w11231;
assign w10908 = (w835 & w10734) | (w835 & ~w9034) | (w10734 & ~w9034);
assign w10909 = (w6230 & w2495) | (w6230 & w10320) | (w2495 & w10320);
assign w10910 = w11055 & w13264;
assign w10911 = ~w10509 & ~w7115;
assign w10912 = (~w13685 & w8167) | (~w13685 & w704) | (w8167 & w704);
assign w10913 = ~w4780 & w2425;
assign w10914 = w144 & w8152;
assign w10915 = (w13324 & w1002) | (w13324 & w5981) | (w1002 & w5981);
assign w10916 = w3219 & w12460;
assign w10917 = (w11395 & w5397) | (w11395 & w151) | (w5397 & w151);
assign w10918 = ~w2941 & ~w4483;
assign w10919 = w3550 & w10444;
assign w10920 = ~w12623 & ~w7765;
assign w10921 = (w6397 & w13329) | (w6397 & w9983) | (w13329 & w9983);
assign w10922 = (w996 & w1920) | (w996 & w14272) | (w1920 & w14272);
assign w10923 = (w9708 & w14623) | (w9708 & w1639) | (w14623 & w1639);
assign w10924 = ~w8937 & w1958;
assign w10925 = ~w2933 & ~w10675;
assign w10926 = w11732 & w8555;
assign w10927 = ~w3067 & w3273;
assign w10928 = ~w6485 & ~w3325;
assign w10929 = (w12656 & ~w12879) | (w12656 & w11123) | (~w12879 & w11123);
assign w10930 = w11861 & w10182;
assign w10931 = ~w11505 & w3410;
assign w10932 = w11458 & ~w11383;
assign w10933 = ~w5122 & ~w5075;
assign w10934 = (w11708 & w8352) | (w11708 & ~w8545) | (w8352 & ~w8545);
assign w10935 = w12481 & ~w4270;
assign w10936 = ~w8234 & ~w2477;
assign w10937 = ~w2849 & w11140;
assign w10938 = w6927 & ~w1469;
assign w10939 = ~w607 & w8396;
assign w10940 = ~w3963 & ~w142;
assign w10941 = b103 & a103;
assign w10942 = ~w13989 & w13145;
assign w10943 = ~w12938 & w8669;
assign w10944 = ~w8748 & w13732;
assign w10945 = ~w9465 & ~w4312;
assign w10946 = ~w12901 & ~w6975;
assign w10947 = (~w7546 & w11957) | (~w7546 & w3209) | (w11957 & w3209);
assign w10948 = (w7082 & w10834) | (w7082 & w12030) | (w10834 & w12030);
assign w10949 = b116 & a116;
assign w10950 = w1509 & w11473;
assign w10951 = w5388 & ~w9605;
assign w10952 = ~w2029 & w9222;
assign w10953 = ~w13952 & ~w6162;
assign w10954 = (w12330 & w6803) | (w12330 & w4520) | (w6803 & w4520);
assign w10955 = w7886 & w2335;
assign w10956 = w1838 & ~w13323;
assign w10957 = (w533 & w7495) | (w533 & w11251) | (w7495 & w11251);
assign w10958 = ~w1221 & w12125;
assign w10959 = w11117 & w6064;
assign w10960 = ~w7305 & w10699;
assign w10961 = ~w9715 & ~w5532;
assign w10962 = (~w3175 & ~w1140) | (~w3175 & w1529) | (~w1140 & w1529);
assign w10963 = (w13983 & ~w13292) | (w13983 & ~w11185) | (~w13292 & ~w11185);
assign w10964 = (~w7475 & w643) | (~w7475 & w5859) | (w643 & w5859);
assign w10965 = w7004 & w8642;
assign w10966 = ~w14302 & ~w2463;
assign w10967 = w6675 & ~w3784;
assign w10968 = (w4148 & w12961) | (w4148 & w7984) | (w12961 & w7984);
assign w10969 = w11997 & w11365;
assign w10970 = w8246 & w12069;
assign w10971 = w4780 & ~w1520;
assign w10972 = ~w2656 & w3502;
assign w10973 = w2671 & w5657;
assign w10974 = w3289 & ~w9138;
assign w10975 = (~w7950 & w12201) | (~w7950 & w10694) | (w12201 & w10694);
assign w10976 = w4658 & w4908;
assign w10977 = ~w13189 & w5282;
assign w10978 = (~w3427 & w1609) | (~w3427 & w6273) | (w1609 & w6273);
assign w10979 = (w3635 & w4149) | (w3635 & ~w7464) | (w4149 & ~w7464);
assign w10980 = (~w3734 & w8937) | (~w3734 & w4750) | (w8937 & w4750);
assign w10981 = w7001 & w2729;
assign w10982 = (w1498 & ~w3209) | (w1498 & w2964) | (~w3209 & w2964);
assign w10983 = w8051 & w12764;
assign w10984 = ~w6583 & ~w6310;
assign w10985 = (~w999 & w1615) | (~w999 & w7510) | (w1615 & w7510);
assign w10986 = ~w6466 & ~w3456;
assign w10987 = w10676 & ~w2135;
assign w10988 = ~w11462 & w11211;
assign w10989 = ~w6151 & ~w6266;
assign w10990 = w1886 & ~w11313;
assign w10991 = ~w5845 & ~w2567;
assign w10992 = ~a0 & ~b0;
assign w10993 = ~w10075 & w7851;
assign w10994 = w7376 & w10792;
assign w10995 = w7754 & ~w5785;
assign w10996 = w13728 & w12793;
assign w10997 = w5178 & w1842;
assign w10998 = ~w1563 & w3611;
assign w10999 = w5231 & w11031;
assign w11000 = w6583 & ~w4033;
assign w11001 = ~w10182 & w10517;
assign w11002 = w1387 & w11732;
assign w11003 = w8056 & ~w11117;
assign w11004 = w14578 & ~w13353;
assign w11005 = ~w8937 & w1083;
assign w11006 = w13398 & ~w14311;
assign w11007 = w7376 & ~w4628;
assign w11008 = ~w7782 & w8225;
assign w11009 = ~w3016 & ~w12229;
assign w11010 = (w7734 & w8614) | (w7734 & w12596) | (w8614 & w12596);
assign w11011 = w5569 & ~w9453;
assign w11012 = ~w9628 & w1621;
assign w11013 = ~b112 & ~a112;
assign w11014 = ~w7953 & ~w8118;
assign w11015 = (~w9853 & w4924) | (~w9853 & ~w8731) | (w4924 & ~w8731);
assign w11016 = w1772 & w13305;
assign w11017 = w7401 & w14208;
assign w11018 = (w11117 & w8565) | (w11117 & w9664) | (w8565 & w9664);
assign w11019 = w12059 & ~w7833;
assign w11020 = ~w6758 & w7547;
assign w11021 = (~w7082 & w14450) | (~w7082 & w12935) | (w14450 & w12935);
assign w11022 = w12483 & ~w12011;
assign w11023 = ~w9836 & w9587;
assign w11024 = w10676 & w6542;
assign w11025 = (~w12464 & ~w6835) | (~w12464 & w5037) | (~w6835 & w5037);
assign w11026 = ~w13282 & ~w3609;
assign w11027 = (~w2060 & w12865) | (~w2060 & w680) | (w12865 & w680);
assign w11028 = (~w10590 & w14141) | (~w10590 & w10671) | (w14141 & w10671);
assign w11029 = (w11959 & w5845) | (w11959 & w8403) | (w5845 & w8403);
assign w11030 = w13805 & ~w6134;
assign w11031 = ~w7335 & ~w10013;
assign w11032 = w4541 & ~w13151;
assign w11033 = ~w6459 & w14275;
assign w11034 = (~w4714 & w13978) | (~w4714 & w2688) | (w13978 & w2688);
assign w11035 = ~w6913 & ~w2955;
assign w11036 = w11586 & ~w749;
assign w11037 = w9607 & ~w2341;
assign w11038 = w9145 & ~w3904;
assign w11039 = ~w7387 & ~w10752;
assign w11040 = w3502 & w8769;
assign w11041 = w325 & w3563;
assign w11042 = ~w13521 & w9296;
assign w11043 = ~w4501 & w4146;
assign w11044 = w7237 & ~w10190;
assign w11045 = ~w13070 & ~w13;
assign w11046 = (w7809 & w5318) | (w7809 & w378) | (w5318 & w378);
assign w11047 = w8609 & ~w12741;
assign w11048 = ~w169 & ~w10106;
assign w11049 = (~w11462 & w265) | (~w11462 & w12829) | (w265 & w12829);
assign w11050 = w9318 & w6381;
assign w11051 = (~w10813 & w2175) | (~w10813 & w6969) | (w2175 & w6969);
assign w11052 = (w4288 & w10462) | (w4288 & w12904) | (w10462 & w12904);
assign w11053 = ~w7656 & w7186;
assign w11054 = (~w11030 & ~w6248) | (~w11030 & w12366) | (~w6248 & w12366);
assign w11055 = ~w3261 & w9401;
assign w11056 = w8657 & ~w9634;
assign w11057 = (w12545 & ~w6785) | (w12545 & w3120) | (~w6785 & w3120);
assign w11058 = (~w7464 & w13695) | (~w7464 & w9369) | (w13695 & w9369);
assign w11059 = ~w5837 & w3375;
assign w11060 = (w3556 & w12145) | (w3556 & w8228) | (w12145 & w8228);
assign w11061 = ~w13928 & ~w1577;
assign w11062 = (w3039 & w11862) | (w3039 & w2750) | (w11862 & w2750);
assign w11063 = ~w2931 & w883;
assign w11064 = ~w842 & ~w13100;
assign w11065 = (~w13587 & w11686) | (~w13587 & w13046) | (w11686 & w13046);
assign w11066 = (~w3145 & w11119) | (~w3145 & w9407) | (w11119 & w9407);
assign w11067 = (~w11429 & w11679) | (~w11429 & w1411) | (w11679 & w1411);
assign w11068 = (~w13565 & w2508) | (~w13565 & w6214) | (w2508 & w6214);
assign w11069 = w1274 & ~w4639;
assign w11070 = (~w7975 & w4527) | (~w7975 & w7784) | (w4527 & w7784);
assign w11071 = w1050 & ~w12163;
assign w11072 = ~w4899 & w13150;
assign w11073 = (~w5785 & w9139) | (~w5785 & w21) | (w9139 & w21);
assign w11074 = w10075 & ~w4359;
assign w11075 = (~w1351 & ~w4148) | (~w1351 & w2179) | (~w4148 & w2179);
assign w11076 = w11088 & ~w10251;
assign w11077 = ~w2590 & ~w3743;
assign w11078 = ~w5490 & w3025;
assign w11079 = (w3585 & w11763) | (w3585 & w7229) | (w11763 & w7229);
assign w11080 = (~w6802 & w10881) | (~w6802 & w6480) | (w10881 & w6480);
assign w11081 = ~w2362 & w5707;
assign w11082 = w8409 & w3564;
assign w11083 = ~w12895 & w2503;
assign w11084 = (w9712 & w5804) | (w9712 & w7206) | (w5804 & w7206);
assign w11085 = ~w9747 & ~w2675;
assign w11086 = ~w13215 & ~w915;
assign w11087 = ~w1282 & w3664;
assign w11088 = ~w2764 & w11309;
assign w11089 = w9672 & w6010;
assign w11090 = w9796 & ~w7308;
assign w11091 = (w14600 & w4799) | (w14600 & w3095) | (w4799 & w3095);
assign w11092 = w8459 & ~w3224;
assign w11093 = (w910 & w7053) | (w910 & w2185) | (w7053 & w2185);
assign w11094 = (~w9012 & w12990) | (~w9012 & w8180) | (w12990 & w8180);
assign w11095 = ~w1387 & w8389;
assign w11096 = w4021 & ~w9938;
assign w11097 = ~w1485 & ~w14157;
assign w11098 = ~w14105 & ~w5554;
assign w11099 = ~w11525 & ~w6627;
assign w11100 = (w6973 & ~w7804) | (w6973 & ~w2197) | (~w7804 & ~w2197);
assign w11101 = w1862 & ~w5664;
assign w11102 = ~w966 & w2484;
assign w11103 = w11117 & w6716;
assign w11104 = (w12943 & w13349) | (w12943 & w8801) | (w13349 & w8801);
assign w11105 = w8626 & w11921;
assign w11106 = ~w13694 & w7487;
assign w11107 = ~w8791 & ~w654;
assign w11108 = ~w10477 & ~w309;
assign w11109 = w13596 & w11557;
assign w11110 = ~w5663 & ~w12231;
assign w11111 = (~w11147 & w12079) | (~w11147 & ~w4842) | (w12079 & ~w4842);
assign w11112 = ~w13282 & ~w2850;
assign w11113 = (w8405 & w5965) | (w8405 & w1024) | (w5965 & w1024);
assign w11114 = ~w5867 & ~w3699;
assign w11115 = (~w2941 & w12759) | (~w2941 & w950) | (w12759 & w950);
assign w11116 = ~w1563 & w1642;
assign w11117 = ~w2036 & ~w1682;
assign w11118 = w11638 & w14335;
assign w11119 = (w14038 & ~w7833) | (w14038 & w50) | (~w7833 & w50);
assign w11120 = w2656 & ~w2998;
assign w11121 = (w7493 & ~w9977) | (w7493 & w10036) | (~w9977 & w10036);
assign w11122 = ~w607 & ~w3427;
assign w11123 = w12656 & w803;
assign w11124 = w3025 & w2492;
assign w11125 = w3963 & w9307;
assign w11126 = (~w11909 & w1615) | (~w11909 & w2936) | (w1615 & w2936);
assign w11127 = w7612 & ~w14247;
assign w11128 = ~w4483 & ~w11117;
assign w11129 = ~w11616 & ~w1205;
assign w11130 = w10676 & ~w2544;
assign w11131 = (~w6266 & w13404) | (~w6266 & ~w2680) | (w13404 & ~w2680);
assign w11132 = w6192 & ~w6700;
assign w11133 = (~w9733 & w7128) | (~w9733 & w7090) | (w7128 & w7090);
assign w11134 = ~w8508 & w8081;
assign w11135 = (w536 & ~w13084) | (w536 & w13250) | (~w13084 & w13250);
assign w11136 = (~w8100 & w7799) | (~w8100 & w3611) | (w7799 & w3611);
assign w11137 = ~w11104 & ~w78;
assign w11138 = ~w11244 & w6018;
assign w11139 = w11272 & w1472;
assign w11140 = w6064 & w646;
assign w11141 = (~w3055 & w2191) | (~w3055 & w6009) | (w2191 & w6009);
assign w11142 = w3288 & ~w646;
assign w11143 = (~w3885 & w4377) | (~w3885 & w11712) | (w4377 & w11712);
assign w11144 = (w3325 & w8769) | (w3325 & w8599) | (w8769 & w8599);
assign w11145 = w7084 & w7832;
assign w11146 = w8018 & w9335;
assign w11147 = w14280 & w1764;
assign w11148 = ~w11108 & w14430;
assign w11149 = w9747 & w10625;
assign w11150 = ~w9686 & w6612;
assign w11151 = ~w5691 & ~w12157;
assign w11152 = (w2112 & w10655) | (w2112 & w6548) | (w10655 & w6548);
assign w11153 = (w8602 & ~w1543) | (w8602 & w9987) | (~w1543 & w9987);
assign w11154 = w159 & ~w6381;
assign w11155 = w11416 & w7910;
assign w11156 = (~w5007 & w10202) | (~w5007 & w11928) | (w10202 & w11928);
assign w11157 = (w11213 & w14421) | (w11213 & ~w11723) | (w14421 & ~w11723);
assign w11158 = ~w13639 & w9806;
assign w11159 = w803 & ~w13531;
assign w11160 = (~w3122 & w10897) | (~w3122 & w6803) | (w10897 & w6803);
assign w11161 = w7914 & w1564;
assign w11162 = w11855 & w1949;
assign w11163 = ~w14351 & ~w1391;
assign w11164 = (w12460 & ~w5490) | (w12460 & w4732) | (~w5490 & w4732);
assign w11165 = (~w11606 & w2823) | (~w11606 & w10573) | (w2823 & w10573);
assign w11166 = (~w10514 & w8937) | (~w10514 & w6059) | (w8937 & w6059);
assign w11167 = ~w2695 & ~w1398;
assign w11168 = w7794 & ~w206;
assign w11169 = ~w14316 & ~w2209;
assign w11170 = ~w3178 & ~w6064;
assign w11171 = w13430 & w10567;
assign w11172 = (w218 & w13152) | (w218 & w6649) | (w13152 & w6649);
assign w11173 = (~w13685 & w3972) | (~w13685 & w2878) | (w3972 & w2878);
assign w11174 = (~w8226 & w10805) | (~w8226 & w11786) | (w10805 & w11786);
assign w11175 = w13732 & w9679;
assign w11176 = ~w1200 & w5842;
assign w11177 = ~w5219 & w8532;
assign w11178 = (w2181 & w4063) | (w2181 & w8204) | (w4063 & w8204);
assign w11179 = ~w2752 & ~w5983;
assign w11180 = w12155 & w3740;
assign w11181 = w2583 & w8929;
assign w11182 = (~w13572 & w6259) | (~w13572 & w2319) | (w6259 & w2319);
assign w11183 = ~w7488 & w6745;
assign w11184 = ~w6832 & w5809;
assign w11185 = (w10719 & w4799) | (w10719 & w3095) | (w4799 & w3095);
assign w11186 = w4884 & w6786;
assign w11187 = w4467 & ~w11488;
assign w11188 = ~w2029 & ~w1375;
assign w11189 = w5040 & w14189;
assign w11190 = w4187 & w5750;
assign w11191 = ~w14343 & w6935;
assign w11192 = w9623 & ~w2941;
assign w11193 = ~w14366 & ~w2644;
assign w11194 = ~w4071 & w2675;
assign w11195 = ~w1384 & w325;
assign w11196 = ~w2218 & w8107;
assign w11197 = ~w7630 & w6927;
assign w11198 = ~w9788 & ~w3563;
assign w11199 = (w13219 & w10028) | (w13219 & w3621) | (w10028 & w3621);
assign w11200 = (w2425 & w4099) | (w2425 & w2726) | (w4099 & w2726);
assign w11201 = ~w2928 & w2068;
assign w11202 = ~w9550 & ~w12828;
assign w11203 = w4836 & ~w885;
assign w11204 = ~w5702 & w6316;
assign w11205 = w5794 & w4897;
assign w11206 = ~w9403 & w4749;
assign w11207 = w3461 & w9346;
assign w11208 = w4039 & ~w14495;
assign w11209 = w13610 & ~w8277;
assign w11210 = (w10853 & w13122) | (w10853 & w2792) | (w13122 & w2792);
assign w11211 = ~w14470 & ~w3159;
assign w11212 = w13438 & w6743;
assign w11213 = w4515 & ~w5560;
assign w11214 = (w5084 & w3357) | (w5084 & w12154) | (w3357 & w12154);
assign w11215 = ~w7630 & w4730;
assign w11216 = ~b89 & ~a89;
assign w11217 = w14051 | ~w5932;
assign w11218 = (w5036 & w10609) | (w5036 & w12581) | (w10609 & w12581);
assign w11219 = w6323 & w11796;
assign w11220 = w2525 | w1634;
assign w11221 = (~w12003 & w9553) | (~w12003 & w323) | (w9553 & w323);
assign w11222 = w830 & w6510;
assign w11223 = ~w1166 & w2410;
assign w11224 = ~w9015 & ~w4127;
assign w11225 = w4618 & ~w6453;
assign w11226 = w1607 & ~w3435;
assign w11227 = w7857 & w3827;
assign w11228 = (~w2922 & w1172) | (~w2922 & w3804) | (w1172 & w3804);
assign w11229 = (~w7022 & w6128) | (~w7022 & w8580) | (w6128 & w8580);
assign w11230 = w6002 & w12185;
assign w11231 = ~w5540 & w9075;
assign w11232 = ~w8442 & ~w9541;
assign w11233 = ~w13257 & ~w13632;
assign w11234 = w3991 & ~w10699;
assign w11235 = w4213 & ~w7122;
assign w11236 = w6825 & w6176;
assign w11237 = w13548 | w11867;
assign w11238 = ~w11992 & ~w12432;
assign w11239 = (~w8992 & w3700) | (~w8992 & w10394) | (w3700 & w10394);
assign w11240 = (w12398 & ~w2492) | (w12398 & w7588) | (~w2492 & w7588);
assign w11241 = (~w10042 & w4050) | (~w10042 & w771) | (w4050 & w771);
assign w11242 = w6493 & w227;
assign w11243 = w9846 & ~w1743;
assign w11244 = w11586 & w12131;
assign w11245 = (w13685 & w10636) | (w13685 & w10843) | (w10636 & w10843);
assign w11246 = (w11817 & w577) | (w11817 & w5592) | (w577 & w5592);
assign w11247 = (w5282 & w9885) | (w5282 & w14614) | (w9885 & w14614);
assign w11248 = w14278 & ~w7060;
assign w11249 = ~w11049 & w7384;
assign w11250 = ~w13623 & ~w640;
assign w11251 = (~w7013 & w3922) | (~w7013 & w8768) | (w3922 & w8768);
assign w11252 = ~w7782 & w4766;
assign w11253 = w1563 & w3430;
assign w11254 = w4836 & w13733;
assign w11255 = ~w11261 & w5885;
assign w11256 = w9971 & w4822;
assign w11257 = ~w12271 & ~w5267;
assign w11258 = (w5650 & w528) | (w5650 & w8927) | (w528 & w8927);
assign w11259 = w8825 & w5608;
assign w11260 = ~w3877 & w12405;
assign w11261 = w3100 & ~w10059;
assign w11262 = w13351 & w5106;
assign w11263 = (~w2218 & w7877) | (~w2218 & w2134) | (w7877 & w2134);
assign w11264 = w7085 & w1197;
assign w11265 = w10961 & w3564;
assign w11266 = (~w4587 & w10216) | (~w4587 & w8472) | (w10216 & w8472);
assign w11267 = ~w183 & w13531;
assign w11268 = w10966 & ~w8808;
assign w11269 = ~w9273 & w7645;
assign w11270 = w10255 & w4790;
assign w11271 = w6111 & ~w12400;
assign w11272 = ~w10013 & ~w8294;
assign w11273 = (~w7914 & w11658) | (~w7914 & ~w3885) | (w11658 & ~w3885);
assign w11274 = (~w6640 & w7758) | (~w6640 & w9201) | (w7758 & w9201);
assign w11275 = w5526 & ~w11200;
assign w11276 = (w3727 & w10648) | (w3727 & w11940) | (w10648 & w11940);
assign w11277 = (~w9012 & w8066) | (~w9012 & w1167) | (w8066 & w1167);
assign w11278 = (~w3615 & w9715) | (~w3615 & w12998) | (w9715 & w12998);
assign w11279 = w13937 & w7376;
assign w11280 = ~w1789 & ~w870;
assign w11281 = (w12569 & ~w1840) | (w12569 & w6227) | (~w1840 & w6227);
assign w11282 = ~w9952 & ~w10941;
assign w11283 = w7670 & w4599;
assign w11284 = ~w2029 & w14440;
assign w11285 = (w2320 & w71) | (w2320 & w1826) | (w71 & w1826);
assign w11286 = w1498 & w2698;
assign w11287 = (~w11013 & w5590) | (~w11013 & w5545) | (w5590 & w5545);
assign w11288 = ~w14629 & ~w14662;
assign w11289 = ~w12121 & w3508;
assign w11290 = w13653 & w4625;
assign w11291 = (~w142 & ~w9211) | (~w142 & w6872) | (~w9211 & w6872);
assign w11292 = ~w8068 & ~w1745;
assign w11293 = ~w8475 & ~w3963;
assign w11294 = ~w13374 & ~w5983;
assign w11295 = ~w8088 & w12437;
assign w11296 = w14137 & w13227;
assign w11297 = ~w9817 & ~w2410;
assign w11298 = ~w9608 & w7313;
assign w11299 = ~w2320 & ~w5860;
assign w11300 = w7599 & w7423;
assign w11301 = ~w3958 & w4728;
assign w11302 = w13159 & ~w5366;
assign w11303 = ~w7718 & ~w8404;
assign w11304 = (~w1692 & w3923) | (~w1692 & w13615) | (w3923 & w13615);
assign w11305 = (w6935 & w11191) | (w6935 & ~w7549) | (w11191 & ~w7549);
assign w11306 = w991 & w120;
assign w11307 = w5178 & ~w13651;
assign w11308 = ~w8963 & w12132;
assign w11309 = w10182 & w3963;
assign w11310 = ~w277 & w6439;
assign w11311 = (~w4050 & w11742) | (~w4050 & w11567) | (w11742 & w11567);
assign w11312 = w1730 & ~w7093;
assign w11313 = (~w727 & w11326) | (~w727 & w11872) | (w11326 & w11872);
assign w11314 = (w11583 & ~w14313) | (w11583 & w12391) | (~w14313 & w12391);
assign w11315 = ~w1563 & w8967;
assign w11316 = ~w2463 & w14200;
assign w11317 = w9558 & ~w11325;
assign w11318 = (w9873 & w9640) | (w9873 & w11925) | (w9640 & w11925);
assign w11319 = w4541 & w2778;
assign w11320 = ~w6339 & ~w10207;
assign w11321 = w11708 & w5304;
assign w11322 = w3925 & w4362;
assign w11323 = w9264 & w5247;
assign w11324 = w2266 & w2177;
assign w11325 = (w1711 & w6978) | (w1711 & w7284) | (w6978 & w7284);
assign w11326 = w9946 & ~w7360;
assign w11327 = (w10578 & w12973) | (w10578 & w9034) | (w12973 & w9034);
assign w11328 = ~w11056 & ~w9850;
assign w11329 = (w9766 & w5957) | (w9766 & w10002) | (w5957 & w10002);
assign w11330 = ~w11528 & w315;
assign w11331 = w10036 & w11613;
assign w11332 = (~w11408 & w197) | (~w11408 & w5302) | (w197 & w5302);
assign w11333 = w9438 & ~w14354;
assign w11334 = (w10318 & ~w353) | (w10318 & w7073) | (~w353 & w7073);
assign w11335 = w6105 & ~w464;
assign w11336 = w12982 & ~w695;
assign w11337 = ~w1503 & ~w10618;
assign w11338 = (~w12958 & ~w14024) | (~w12958 & w3623) | (~w14024 & w3623);
assign w11339 = ~w4503 & w9021;
assign w11340 = ~w3256 & ~w12429;
assign w11341 = w1016 & w3039;
assign w11342 = ~w10334 & ~w9399;
assign w11343 = (w5912 & ~w7625) | (w5912 & w1355) | (~w7625 & w1355);
assign w11344 = (w11817 & w1563) | (w11817 & w6497) | (w1563 & w6497);
assign w11345 = b35 & a35;
assign w11346 = w1527 & w4092;
assign w11347 = (~w2939 & w6389) | (~w2939 & w4956) | (w6389 & w4956);
assign w11348 = ~w12614 & ~w10548;
assign w11349 = w12569 & w13677;
assign w11350 = w6889 & w1274;
assign w11351 = ~w8966 & ~w10931;
assign w11352 = ~w8744 & ~w3651;
assign w11353 = ~w4700 & w10427;
assign w11354 = w5761 & w8475;
assign w11355 = w7794 & ~w5325;
assign w11356 = (w3025 & w71) | (w3025 & w8722) | (w71 & w8722);
assign w11357 = w1744 & w960;
assign w11358 = w3917 & w2505;
assign w11359 = (w9608 & w3140) | (w9608 & w9114) | (w3140 & w9114);
assign w11360 = ~w6810 & ~w10657;
assign w11361 = b31 & a31;
assign w11362 = ~w14222 & ~w9795;
assign w11363 = w12121 & ~w1442;
assign w11364 = w6500 & w12642;
assign w11365 = w4855 & ~w309;
assign w11366 = w8475 & w4458;
assign w11367 = w9092 | w18;
assign w11368 = ~w1540 & ~w3645;
assign w11369 = w3905 & ~w3543;
assign w11370 = (~w6802 & w3237) | (~w6802 & w10003) | (w3237 & w10003);
assign w11371 = w8795 & w12256;
assign w11372 = w6281 & ~w14526;
assign w11373 = w7794 & w820;
assign w11374 = (~w14455 & ~w8337) | (~w14455 & w4007) | (~w8337 & w4007);
assign w11375 = ~w14378 & ~w10981;
assign w11376 = w1802 & w10182;
assign w11377 = (~w4363 & ~w9994) | (~w4363 & ~w5124) | (~w9994 & ~w5124);
assign w11378 = ~w5852 & w1007;
assign w11379 = (w8450 & w6681) | (w8450 & w4660) | (w6681 & w4660);
assign w11380 = ~w3807 & ~w10627;
assign w11381 = (~w13685 & w7304) | (~w13685 & w11854) | (w7304 & w11854);
assign w11382 = ~w9284 & w3427;
assign w11383 = (~w4627 & ~w1986) | (~w4627 & w5137) | (~w1986 & w5137);
assign w11384 = (w5952 & w1680) | (w5952 & w11368) | (w1680 & w11368);
assign w11385 = ~w4756 & w5783;
assign w11386 = ~w2355 & w8396;
assign w11387 = ~w14028 & ~w13713;
assign w11388 = ~w13609 & w2284;
assign w11389 = w10486 & w3248;
assign w11390 = w2629 & w13320;
assign w11391 = w5548 & w1980;
assign w11392 = ~w12545 & w3386;
assign w11393 = ~w13350 & w9278;
assign w11394 = ~w12606 & ~w12617;
assign w11395 = b63 & a63;
assign w11396 = ~w5090 & w13443;
assign w11397 = ~w9620 & ~w12734;
assign w11398 = ~w14513 & w9864;
assign w11399 = w10165 & ~w2381;
assign w11400 = ~w7763 & w12594;
assign w11401 = ~w14204 & w2375;
assign w11402 = ~w4700 & w1540;
assign w11403 = w654 & ~w2989;
assign w11404 = w12464 & ~w5934;
assign w11405 = w13492 & w9559;
assign w11406 = w1563 & ~w8018;
assign w11407 = ~w5584 & w10250;
assign w11408 = ~w9359 & w7086;
assign w11409 = ~w1062 & ~w8758;
assign w11410 = ~w4033 & ~w3751;
assign w11411 = ~w4712 & ~w9409;
assign w11412 = w9923 & w4833;
assign w11413 = (~w4545 & w13543) | (~w4545 & w3520) | (w13543 & w3520);
assign w11414 = ~w6855 & w2833;
assign w11415 = (~w2655 & w6751) | (~w2655 & w5117) | (w6751 & w5117);
assign w11416 = (~w3209 & ~w11429) | (~w3209 & w3564) | (~w11429 & w3564);
assign w11417 = (~w6219 & w2603) | (~w6219 & w11741) | (w2603 & w11741);
assign w11418 = (~w14417 & ~w4511) | (~w14417 & ~w11756) | (~w4511 & ~w11756);
assign w11419 = w9454 & w1623;
assign w11420 = ~w6065 & w6255;
assign w11421 = ~w71 & w13128;
assign w11422 = (w14074 & w11601) | (w14074 & w9644) | (w11601 & w9644);
assign w11423 = w6861 & w3790;
assign w11424 = w4431 & ~w13358;
assign w11425 = (w8623 & w10344) | (w8623 & w11523) | (w10344 & w11523);
assign w11426 = (~w6276 & w1081) | (~w6276 & w10086) | (w1081 & w10086);
assign w11427 = w5412 & w8113;
assign w11428 = w10746 & w9124;
assign w11429 = w6097 & ~w13367;
assign w11430 = ~w14578 & ~w11937;
assign w11431 = ~w2291 & ~w45;
assign w11432 = w13160 & ~w5948;
assign w11433 = (~w8085 & w71) | (~w8085 & w7960) | (w71 & w7960);
assign w11434 = (w325 & w5394) | (w325 & w11195) | (w5394 & w11195);
assign w11435 = (w3550 & w3253) | (w3550 & w11494) | (w3253 & w11494);
assign w11436 = ~w9608 & w10102;
assign w11437 = ~w13256 & w7022;
assign w11438 = w12398 & w12135;
assign w11439 = (w5768 & w13772) | (w5768 & w7041) | (w13772 & w7041);
assign w11440 = ~w10334 & ~w5305;
assign w11441 = w7794 & ~w5831;
assign w11442 = ~w1221 & ~w10523;
assign w11443 = w13713 & ~w3019;
assign w11444 = w10631 & ~w10727;
assign w11445 = (~w142 & ~w11934) | (~w142 & w6872) | (~w11934 & w6872);
assign w11446 = w1447 & ~w6698;
assign w11447 = ~w6949 & w5490;
assign w11448 = (~w7796 & ~w82) | (~w7796 & ~w4232) | (~w82 & ~w4232);
assign w11449 = (w14195 & w1444) | (w14195 & w1875) | (w1444 & w1875);
assign w11450 = w11031 & ~w12356;
assign w11451 = ~w14383 & w11478;
assign w11452 = w14588 & ~w13323;
assign w11453 = w13686 & w14389;
assign w11454 = ~b2 & ~a2;
assign w11455 = ~w10941 & w11117;
assign w11456 = w10224 & w8442;
assign w11457 = ~w12856 & ~w1264;
assign w11458 = ~w922 & ~w8226;
assign w11459 = ~w3178 & w13845;
assign w11460 = (~w8951 & ~w7703) | (~w8951 & w2245) | (~w7703 & w2245);
assign w11461 = ~w3117 & ~w9761;
assign w11462 = b40 & a40;
assign w11463 = w9638 & w11293;
assign w11464 = w5283 & w11117;
assign w11465 = w3671 & ~w11266;
assign w11466 = (~w12886 & w3286) | (~w12886 & w6437) | (w3286 & w6437);
assign w11467 = w14121 & ~w12019;
assign w11468 = w9433 & ~w2470;
assign w11469 = w5537 & ~w403;
assign w11470 = w12173 & w14627;
assign w11471 = w1268 & w7330;
assign w11472 = (w3929 & w9221) | (w3929 & w8282) | (w9221 & w8282);
assign w11473 = ~w3096 & w12173;
assign w11474 = ~w3784 & w2332;
assign w11475 = ~w10309 & ~w11345;
assign w11476 = ~w5522 & ~w2941;
assign w11477 = ~w13249 & w1540;
assign w11478 = (~w2795 & ~w10030) | (~w2795 & w13121) | (~w10030 & w13121);
assign w11479 = ~w12563 & w130;
assign w11480 = w6266 & ~w8531;
assign w11481 = ~w4607 & ~w4979;
assign w11482 = w1809 & ~w803;
assign w11483 = ~w12751 & w2594;
assign w11484 = ~w1824 & w5238;
assign w11485 = w10676 & w10997;
assign w11486 = w8234 & w9015;
assign w11487 = ~w3215 & ~w1027;
assign w11488 = b61 & a61;
assign w11489 = ~w1166 & w6542;
assign w11490 = ~w12448 & w13406;
assign w11491 = ~w8552 & ~w10404;
assign w11492 = ~w12240 & ~w2218;
assign w11493 = w2680 & ~w3508;
assign w11494 = ~w6795 & w13820;
assign w11495 = ~w2996 & ~w3727;
assign w11496 = ~w4265 & ~w1413;
assign w11497 = w11604 & ~w6317;
assign w11498 = w1705 & ~w1963;
assign w11499 = w10075 & ~w6230;
assign w11500 = w9940 & w8047;
assign w11501 = w3153 & w8986;
assign w11502 = ~w14141 & w1635;
assign w11503 = (~w3823 & ~w3609) | (~w3823 & w456) | (~w3609 & w456);
assign w11504 = (~w6802 & w5484) | (~w6802 & w8190) | (w5484 & w8190);
assign w11505 = ~w6580 & ~w5282;
assign w11506 = w5778 & ~w12216;
assign w11507 = w14640 & ~w646;
assign w11508 = ~w5696 & w5272;
assign w11509 = (w3847 & w3171) | (w3847 & ~w6264) | (w3171 & ~w6264);
assign w11510 = ~w8422 & w13780;
assign w11511 = (w10322 & w4046) | (w10322 & w7290) | (w4046 & w7290);
assign w11512 = (~w14460 & w8511) | (~w14460 & w11674) | (w8511 & w11674);
assign w11513 = (w1164 & w4107) | (w1164 & w1959) | (w4107 & w1959);
assign w11514 = w13548 | w8771;
assign w11515 = w13189 & w1743;
assign w11516 = ~w6963 & ~w318;
assign w11517 = ~w5762 & w5610;
assign w11518 = ~w9636 & w6204;
assign w11519 = w8162 & w9076;
assign w11520 = (w2029 & w6395) | (w2029 & w6642) | (w6395 & w6642);
assign w11521 = (w12493 & w13348) | (w12493 & w11639) | (w13348 & w11639);
assign w11522 = (~w10688 & ~w6656) | (~w10688 & w8405) | (~w6656 & w8405);
assign w11523 = w5505 & w9655;
assign w11524 = (w13595 & w3818) | (w13595 & w13281) | (w3818 & w13281);
assign w11525 = ~w11871 & w13837;
assign w11526 = (w5482 & w10462) | (w5482 & w2133) | (w10462 & w2133);
assign w11527 = ~w11197 & ~w2698;
assign w11528 = w3384 & ~w7868;
assign w11529 = (w4756 & w10726) | (w4756 & w11644) | (w10726 & w11644);
assign w11530 = ~w7141 & w4821;
assign w11531 = ~w170 & ~w8962;
assign w11532 = ~w12121 & ~w13953;
assign w11533 = ~w14072 & ~w8516;
assign w11534 = (w7757 & w10418) | (w7757 & ~w11516) | (w10418 & ~w11516);
assign w11535 = w9465 & ~w6281;
assign w11536 = ~w10339 & ~w10433;
assign w11537 = (~w4781 & w11898) | (~w4781 & w380) | (w11898 & w380);
assign w11538 = w7376 & w894;
assign w11539 = ~w1785 & w336;
assign w11540 = ~w4032 & w13957;
assign w11541 = w11046 | w3638;
assign w11542 = (w3025 & ~w14055) | (w3025 & w9227) | (~w14055 & w9227);
assign w11543 = (~w6802 & w12770) | (~w6802 & w4614) | (w12770 & w4614);
assign w11544 = w3128 & w14488;
assign w11545 = ~w5827 & w5998;
assign w11546 = ~w9115 & ~w824;
assign w11547 = ~b8 & ~a8;
assign w11548 = w3488 & w12062;
assign w11549 = (w7343 & w9573) | (w7343 & w2383) | (w9573 & w2383);
assign w11550 = ~w13324 & w8538;
assign w11551 = (~w884 & w9366) | (~w884 & w11921) | (w9366 & w11921);
assign w11552 = w8975 & ~w7233;
assign w11553 = w149 & w10243;
assign w11554 = (~w922 & w3413) | (~w922 & w3082) | (w3413 & w3082);
assign w11555 = w10676 & w3717;
assign w11556 = ~w3092 & ~w2379;
assign w11557 = w5660 & w813;
assign w11558 = (w3025 & w4896) | (w3025 & w3209) | (w4896 & w3209);
assign w11559 = ~w12452 & w8763;
assign w11560 = ~b46 & ~a46;
assign w11561 = w7384 & w2909;
assign w11562 = w1989 & ~w7755;
assign w11563 = ~w5523 & ~w11543;
assign w11564 = (w2941 & ~w5912) | (w2941 & w1336) | (~w5912 & w1336);
assign w11565 = ~w7808 & w11861;
assign w11566 = w39 & ~w12575;
assign w11567 = w9170 & w12325;
assign w11568 = (w11261 & w14326) | (w11261 & w12607) | (w14326 & w12607);
assign w11569 = w6538 & ~w8026;
assign w11570 = ~w5522 & ~w2729;
assign w11571 = w2913 & ~w12426;
assign w11572 = ~w11745 & ~w10699;
assign w11573 = w3821 & w1858;
assign w11574 = w14027 & ~w9895;
assign w11575 = ~w1499 & ~w8783;
assign w11576 = w3483 & w12614;
assign w11577 = w9921 & w10045;
assign w11578 = (w12460 & w5005) | (w12460 & w622) | (w5005 & w622);
assign w11579 = ~w183 & ~w13587;
assign w11580 = (w4987 & w7482) | (w4987 & ~w12889) | (w7482 & ~w12889);
assign w11581 = ~w7178 & w7024;
assign w11582 = w12982 & w9917;
assign w11583 = ~w7906 & w1699;
assign w11584 = (~w3435 & w2463) | (~w3435 & w4535) | (w2463 & w4535);
assign w11585 = w5860 & w8769;
assign w11586 = ~w11033 & w6294;
assign w11587 = (~w12376 & w8804) | (~w12376 & w6246) | (w8804 & w6246);
assign w11588 = (w14216 & w13869) | (w14216 & w13779) | (w13869 & w13779);
assign w11589 = w4982 & ~w5185;
assign w11590 = w11643 & ~w1929;
assign w11591 = (~w8396 & ~w3806) | (~w8396 & w7310) | (~w3806 & w7310);
assign w11592 = w9921 & w3098;
assign w11593 = (~w10618 & w11337) | (~w10618 & w3225) | (w11337 & w3225);
assign w11594 = (~w3091 & w111) | (~w3091 & w4912) | (w111 & w4912);
assign w11595 = ~w1840 & ~w10423;
assign w11596 = ~w198 & ~w7794;
assign w11597 = w14015 & w10182;
assign w11598 = ~w13733 & ~w12575;
assign w11599 = w1337 & w3090;
assign w11600 = (w6473 & w11135) | (w6473 & w5211) | (w11135 & w5211);
assign w11601 = w1872 & ~w6018;
assign w11602 = w10485 & w6099;
assign w11603 = (w2655 & w335) | (w2655 & w10922) | (w335 & w10922);
assign w11604 = ~w894 & ~w5860;
assign w11605 = w12893 & ~w5664;
assign w11606 = ~b42 & ~a42;
assign w11607 = ~w8192 & w5588;
assign w11608 = ~w2858 & w9748;
assign w11609 = (w11106 & w14229) | (w11106 & w7549) | (w14229 & w7549);
assign w11610 = (~w3550 & w12748) | (~w3550 & w10227) | (w12748 & w10227);
assign w11611 = ~w4983 & ~w12850;
assign w11612 = (~w6426 & w1347) | (~w6426 & w14448) | (w1347 & w14448);
assign w11613 = w11500 & w7085;
assign w11614 = w217 & w12642;
assign w11615 = ~w7662 & w3615;
assign w11616 = ~w5559 & w13702;
assign w11617 = w985 & w3103;
assign w11618 = w3098 & ~w803;
assign w11619 = ~w10554 & ~w8291;
assign w11620 = (w2962 & w1708) | (w2962 & ~w10647) | (w1708 & ~w10647);
assign w11621 = ~w2629 & w7670;
assign w11622 = (w6890 & ~w1744) | (w6890 & w13090) | (~w1744 & w13090);
assign w11623 = (w7152 & w4762) | (w7152 & w5251) | (w4762 & w5251);
assign w11624 = (w1235 & w12998) | (w1235 & w14350) | (w12998 & w14350);
assign w11625 = (~w14395 & w4050) | (~w14395 & w2106) | (w4050 & w2106);
assign w11626 = (w7082 & w13996) | (w7082 & w13025) | (w13996 & w13025);
assign w11627 = w5177 & ~w2270;
assign w11628 = w11617 & w6383;
assign w11629 = w8964 & ~w14426;
assign w11630 = w13111 & w3650;
assign w11631 = ~w5218 & w1535;
assign w11632 = ~w14020 & ~w5216;
assign w11633 = ~w13531 & w536;
assign w11634 = (~w2670 & w14182) | (~w2670 & w302) | (w14182 & w302);
assign w11635 = ~w13565 & ~w2410;
assign w11636 = ~w11438 & ~w4796;
assign w11637 = w7847 & w7902;
assign w11638 = w5243 & w9170;
assign w11639 = (~w5406 & w8191) | (~w5406 & ~w14417) | (w8191 & ~w14417);
assign w11640 = w4349 & ~w3111;
assign w11641 = (w3611 & w12980) | (w3611 & w6773) | (w12980 & w6773);
assign w11642 = ~w2029 & w12490;
assign w11643 = w347 & w11909;
assign w11644 = (~w13306 & w4952) | (~w13306 & w235) | (w4952 & w235);
assign w11645 = w7177 & ~w12902;
assign w11646 = w11899 & w13732;
assign w11647 = w14028 & w12959;
assign w11648 = ~w8125 & w2868;
assign w11649 = w1802 & w4458;
assign w11650 = ~w10256 & w8518;
assign w11651 = w3550 & w2577;
assign w11652 = w12987 & ~w3050;
assign w11653 = w3914 & w10317;
assign w11654 = w8253 & w6689;
assign w11655 = ~w309 & w1016;
assign w11656 = w14203 & w12813;
assign w11657 = ~w4071 & ~w3174;
assign w11658 = w9788 & ~w7914;
assign w11659 = ~w7376 & w13733;
assign w11660 = w5177 & w2332;
assign w11661 = ~w11063 & w10604;
assign w11662 = w2945 & ~w5243;
assign w11663 = ~w10791 & w3909;
assign w11664 = (w9749 & w415) | (w9749 & w2510) | (w415 & w2510);
assign w11665 = w10013 & ~w3904;
assign w11666 = ~w8540 & w11940;
assign w11667 = (w13311 & w14650) | (w13311 & w4756) | (w14650 & w4756);
assign w11668 = w12624 & ~w12844;
assign w11669 = ~w1609 & w14139;
assign w11670 = (w9454 & w13152) | (w9454 & w3868) | (w13152 & w3868);
assign w11671 = (~w4050 & w4138) | (~w4050 & w7555) | (w4138 & w7555);
assign w11672 = w14335 & ~w9379;
assign w11673 = ~w6716 & ~w2492;
assign w11674 = (~w11737 & w8511) | (~w11737 & w2921) | (w8511 & w2921);
assign w11675 = ~w3209 & ~w10855;
assign w11676 = (w12859 & w6832) | (w12859 & w4274) | (w6832 & w4274);
assign w11677 = ~w11038 & ~w967;
assign w11678 = ~b93 & ~w3813;
assign w11679 = w10725 & ~w3209;
assign w11680 = w5177 & ~w71;
assign w11681 = w8512 & w4541;
assign w11682 = w5765 & w14419;
assign w11683 = ~w14240 & w9645;
assign w11684 = ~w8253 & ~w8475;
assign w11685 = w9454 & ~w10771;
assign w11686 = w10290 & ~w309;
assign w11687 = w5761 & ~w6064;
assign w11688 = w3364 & w10341;
assign w11689 = ~w318 & w6301;
assign w11690 = w6324 & w3727;
assign w11691 = ~w8937 & w1463;
assign w11692 = (~w12949 & ~w7006) | (~w12949 & w1132) | (~w7006 & w1132);
assign w11693 = ~w6080 & ~w12479;
assign w11694 = (~w13674 & ~w10311) | (~w13674 & w2790) | (~w10311 & w2790);
assign w11695 = ~w14633 & ~w4964;
assign w11696 = ~w1723 & w5950;
assign w11697 = ~w7423 & w7379;
assign w11698 = ~w12677 & w5128;
assign w11699 = w10165 & ~w8499;
assign w11700 = (w11973 & w5672) | (w11973 & w5403) | (w5672 & w5403);
assign w11701 = ~w4921 & w13671;
assign w11702 = ~w8394 & ~w1752;
assign w11703 = (w10675 & w5559) | (w10675 & w12711) | (w5559 & w12711);
assign w11704 = w5741 & w2941;
assign w11705 = ~w7376 & w7914;
assign w11706 = (w4473 & w13122) | (w4473 & w10859) | (w13122 & w10859);
assign w11707 = w967 & w8356;
assign w11708 = w1171 & w11108;
assign w11709 = (w1721 & w7156) | (w1721 & w2670) | (w7156 & w2670);
assign w11710 = ~w13237 & w10689;
assign w11711 = ~w4751 & w12943;
assign w11712 = w4582 & w10711;
assign w11713 = (w13426 & ~w10177) | (w13426 & w8164) | (~w10177 & w8164);
assign w11714 = (~w803 & w183) | (~w803 & w10689) | (w183 & w10689);
assign w11715 = ~w14478 & ~w408;
assign w11716 = w4127 & ~w6572;
assign w11717 = w14251 & w3147;
assign w11718 = w8181 & ~w4991;
assign w11719 = ~w10605 & ~w7423;
assign w11720 = ~w192 & ~w2001;
assign w11721 = ~w12856 & w11708;
assign w11722 = w2966 & w11320;
assign w11723 = w10339 & ~w12685;
assign w11724 = ~w11259 & w4797;
assign w11725 = ~w372 & ~w11361;
assign w11726 = ~w14474 & w8787;
assign w11727 = w13937 & w3456;
assign w11728 = ~w12240 & ~w8080;
assign w11729 = (~w7515 & w12834) | (~w7515 & w1366) | (w12834 & w1366);
assign w11730 = (~w254 & w3741) | (~w254 & w3176) | (w3741 & w3176);
assign w11731 = w3547 & ~w2114;
assign w11732 = (~w3502 & w5692) | (~w3502 & w10607) | (w5692 & w10607);
assign w11733 = ~w9696 & ~w2296;
assign w11734 = (w5483 & w4344) | (w5483 & w11385) | (w4344 & w11385);
assign w11735 = w14526 & w1114;
assign w11736 = ~w8052 & ~w1913;
assign w11737 = w6125 & ~w720;
assign w11738 = (~w14519 & ~w7152) | (~w14519 & w13630) | (~w7152 & w13630);
assign w11739 = (~w11818 & w7803) | (~w11818 & w5680) | (w7803 & w5680);
assign w11740 = w10676 & w3602;
assign w11741 = w2872 & ~w6219;
assign w11742 = w9170 & w8718;
assign w11743 = ~w6463 & w2321;
assign w11744 = (w5768 & w2977) | (w5768 & w10954) | (w2977 & w10954);
assign w11745 = b97 & a97;
assign w11746 = w6098 & ~w8677;
assign w11747 = ~w2762 & ~w9145;
assign w11748 = ~w183 & ~w2858;
assign w11749 = (~w12406 & w46) | (~w12406 & w3796) | (w46 & w3796);
assign w11750 = ~w5867 & ~w9012;
assign w11751 = ~w3827 & ~w13592;
assign w11752 = ~w2284 & w14334;
assign w11753 = ~w10016 & ~w7502;
assign w11754 = ~w9171 & ~w11379;
assign w11755 = w10930 & w9499;
assign w11756 = ~w2313 & w10022;
assign w11757 = ~b122 & ~a122;
assign w11758 = w13398 & w12643;
assign w11759 = ~w3912 & w12895;
assign w11760 = ~w8183 & ~w8253;
assign w11761 = ~w1330 & ~w3205;
assign w11762 = (w9985 & w3843) | (w9985 & w3897) | (w3843 & w3897);
assign w11763 = ~w11117 & ~w10286;
assign w11764 = ~w9747 & ~w1076;
assign w11765 = (w11613 & w6299) | (w11613 & w10681) | (w6299 & w10681);
assign w11766 = ~w9988 & ~w5179;
assign w11767 = ~w3386 & w6500;
assign w11768 = ~w1714 & ~w5843;
assign w11769 = w6580 & ~w12047;
assign w11770 = (w1753 & w6943) | (w1753 & w6667) | (w6943 & w6667);
assign w11771 = w3522 & w12460;
assign w11772 = w5522 & w2729;
assign w11773 = (w1607 & w13122) | (w1607 & w14668) | (w13122 & w14668);
assign w11774 = ~w3047 & ~w556;
assign w11775 = (~w10507 & w8937) | (~w10507 & w4514) | (w8937 & w4514);
assign w11776 = w2433 & ~w4458;
assign w11777 = ~w3289 | w9298;
assign w11778 = w1166 & w9830;
assign w11779 = ~w473 & ~w2872;
assign w11780 = (w919 & w9161) | (w919 & w3680) | (w9161 & w3680);
assign w11781 = ~w1015 & ~w4756;
assign w11782 = ~w840 & w12210;
assign w11783 = ~w3271 & w6372;
assign w11784 = ~w3914 & w3025;
assign w11785 = w9419 & ~w10131;
assign w11786 = (w9572 & w3081) | (w9572 & w1966) | (w3081 & w1966);
assign w11787 = w4483 & ~w7719;
assign w11788 = w5693 & w6301;
assign w11789 = w13506 & ~w4796;
assign w11790 = (w14593 & w9271) | (w14593 & w6631) | (w9271 & w6631);
assign w11791 = w8532 & w2474;
assign w11792 = w8748 & w4193;
assign w11793 = ~w2144 & w909;
assign w11794 = ~w5724 & w7808;
assign w11795 = ~w4570 & w10882;
assign w11796 = (~w12908 & w11475) | (~w12908 & w12419) | (w11475 & w12419);
assign w11797 = ~w210 & ~w4672;
assign w11798 = w9716 & ~w8396;
assign w11799 = ~w10245 & w6833;
assign w11800 = w2268 & ~w4697;
assign w11801 = w8148 & ~w2875;
assign w11802 = (~w4050 & w1126) | (~w4050 & w13631) | (w1126 & w13631);
assign w11803 = ~w12553 & ~w2029;
assign w11804 = ~w13587 & w13069;
assign w11805 = ~w10826 & ~w2019;
assign w11806 = (~w4780 & w10913) | (~w4780 & w12782) | (w10913 & w12782);
assign w11807 = ~w9247 & w796;
assign w11808 = ~w2202 & w0;
assign w11809 = ~w10038 & w13890;
assign w11810 = ~w2410 & ~w12317;
assign w11811 = ~w7193 & ~w7628;
assign w11812 = (w13970 & w4541) | (w13970 & w5881) | (w4541 & w5881);
assign w11813 = w330 & w2499;
assign w11814 = (w11803 & w2180) | (w11803 & w8922) | (w2180 & w8922);
assign w11815 = w8345 & ~w8351;
assign w11816 = (w5422 & w4105) | (w5422 & w1169) | (w4105 & w1169);
assign w11817 = ~w1821 & ~w3219;
assign w11818 = ~w13693 & w14205;
assign w11819 = (w659 & w3505) | (w659 & w12568) | (w3505 & w12568);
assign w11820 = ~w12668 & ~w8236;
assign w11821 = w6500 & ~w11394;
assign w11822 = w10224 & ~w13117;
assign w11823 = ~w14116 & w1935;
assign w11824 = ~w1795 & w5247;
assign w11825 = w9776 & ~w11419;
assign w11826 = (w1619 & w8921) | (w1619 & w4354) | (w8921 & w4354);
assign w11827 = w1263 & ~w10754;
assign w11828 = (~w6266 & w13404) | (~w6266 & ~w5520) | (w13404 & ~w5520);
assign w11829 = ~w11861 & ~w3991;
assign w11830 = (w7082 & w3832) | (w7082 & w10683) | (w3832 & w10683);
assign w11831 = (w6832 & w1251) | (w6832 & w13523) | (w1251 & w13523);
assign w11832 = (w10290 & w8569) | (w10290 & ~w8992) | (w8569 & ~w8992);
assign w11833 = ~w1384 & ~w3742;
assign w11834 = w2260 & w4064;
assign w11835 = w7914 & w12879;
assign w11836 = w3947 & w11310;
assign w11837 = (w13391 & w9103) | (w13391 & ~w14182) | (w9103 & ~w14182);
assign w11838 = ~w1534 & ~w9415;
assign w11839 = w4213 & ~w10669;
assign w11840 = (w3537 & w8767) | (w3537 & w729) | (w8767 & w729);
assign w11841 = ~w14139 & w4859;
assign w11842 = (w8937 & w6793) | (w8937 & w1693) | (w6793 & w1693);
assign w11843 = (w7272 & w3231) | (w7272 & w13202) | (w3231 & w13202);
assign w11844 = w3547 & w1574;
assign w11845 = ~w2008 & w13190;
assign w11846 = ~w4875 & w5055;
assign w11847 = ~w3435 & w5490;
assign w11848 = ~w11025 & ~w4549;
assign w11849 = (w14463 & w12562) | (w14463 & w9684) | (w12562 & w9684);
assign w11850 = ~w8769 & ~w2439;
assign w11851 = w5294 & ~w2850;
assign w11852 = w14442 | w2309;
assign w11853 = w2320 & w3885;
assign w11854 = (~w4783 & ~w6637) | (~w4783 & ~w12376) | (~w6637 & ~w12376);
assign w11855 = ~w6716 & ~w829;
assign w11856 = (w6719 & w13504) | (w6719 & w5595) | (w13504 & w5595);
assign w11857 = (w12332 & w11923) | (w12332 & ~w8444) | (w11923 & ~w8444);
assign w11858 = ~w10856 & ~w517;
assign w11859 = ~w5691 & w7490;
assign w11860 = ~w11057 & ~w9510;
assign w11861 = ~w8475 & ~w11013;
assign w11862 = ~w8384 & ~w5685;
assign w11863 = ~w6047 & w2480;
assign w11864 = w5803 & w112;
assign w11865 = w1673 & ~w11307;
assign w11866 = w8018 & ~w13713;
assign w11867 = w14624 & w2691;
assign w11868 = w9200 & w6845;
assign w11869 = w10300 & ~w5489;
assign w11870 = (w8120 & w12087) | (w8120 & w4164) | (w12087 & w4164);
assign w11871 = ~w2509 & ~w6538;
assign w11872 = ~w13789 & ~w727;
assign w11873 = ~w6986 & w8174;
assign w11874 = w11328 & w13009;
assign w11875 = ~w8290 & ~w5247;
assign w11876 = ~w5035 & ~w5247;
assign w11877 = ~w5823 & w3427;
assign w11878 = ~w9805 & ~w13761;
assign w11879 = ~w1661 & ~w1168;
assign w11880 = (w9074 & ~w1242) | (w9074 & w586) | (~w1242 & w586);
assign w11881 = (w2331 & w8087) | (w2331 & w11334) | (w8087 & w11334);
assign w11882 = w7772 & w4541;
assign w11883 = ~w12373 & w4372;
assign w11884 = w4836 & w608;
assign w11885 = (w6939 & w7871) | (w6939 & w8344) | (w7871 & w8344);
assign w11886 = ~w11462 & ~w5785;
assign w11887 = ~w9333 & w9531;
assign w11888 = ~w10435 & w684;
assign w11889 = w442 & ~w101;
assign w11890 = ~w2387 & ~w1842;
assign w11891 = w509 & w489;
assign w11892 = (w14302 & w4160) | (w14302 & w9900) | (w4160 & w9900);
assign w11893 = ~w6569 & ~w4831;
assign w11894 = ~w3067 & w8221;
assign w11895 = (~w3194 & w12252) | (~w3194 & w7245) | (w12252 & w7245);
assign w11896 = (w7571 & w4061) | (w7571 & ~w9591) | (w4061 & ~w9591);
assign w11897 = w4322 & w10699;
assign w11898 = (~w3682 & w11217) | (~w3682 & w2090) | (w11217 & w2090);
assign w11899 = w1062 & w1540;
assign w11900 = w6501 & w7504;
assign w11901 = ~w6274 & w513;
assign w11902 = ~w3219 & ~w4129;
assign w11903 = ~w12240 & w4165;
assign w11904 = w4848 & ~w7244;
assign w11905 = ~b83 & ~a83;
assign w11906 = ~w1778 & ~w2694;
assign w11907 = ~w3957 & w10647;
assign w11908 = w10326 & w9989;
assign w11909 = w3717 & w10880;
assign w11910 = w9032 & ~w10075;
assign w11911 = w4026 & ~w2765;
assign w11912 = ~w11360 & w9427;
assign w11913 = w11746 & w9187;
assign w11914 = ~w4032 & ~w14070;
assign w11915 = ~w4756 & w5506;
assign w11916 = w5574 & w8666;
assign w11917 = w4078 & ~w8110;
assign w11918 = w2475 & ~w9723;
assign w11919 = (w8769 & w5355) | (w8769 & w12631) | (w5355 & w12631);
assign w11920 = ~w8226 & w13308;
assign w11921 = w2680 & ~w884;
assign w11922 = ~w9220 & ~w962;
assign w11923 = (w8983 & w8117) | (w8983 & w7107) | (w8117 & w7107);
assign w11924 = (~w13587 & w10750) | (~w13587 & w599) | (w10750 & w599);
assign w11925 = (~w1254 & w4722) | (~w1254 & w9386) | (w4722 & w9386);
assign w11926 = (~w6500 & w1609) | (~w6500 & w13701) | (w1609 & w13701);
assign w11927 = w7170 & w9980;
assign w11928 = (w7578 & w8770) | (w7578 & ~w353) | (w8770 & ~w353);
assign w11929 = w5669 & w710;
assign w11930 = (w8584 & w10467) | (w8584 & w1096) | (w10467 & w1096);
assign w11931 = ~w10906 & ~w9582;
assign w11932 = ~w1828 & w10749;
assign w11933 = (w2272 & w12646) | (w2272 & w12154) | (w12646 & w12154);
assign w11934 = ~w10032 & ~w13189;
assign w11935 = w3914 & ~w10855;
assign w11936 = (~w9794 & w13269) | (~w9794 & ~w1928) | (w13269 & ~w1928);
assign w11937 = ~w2317 & w9992;
assign w11938 = ~w14141 & w3051;
assign w11939 = (~w9747 & w5985) | (~w9747 & w6071) | (w5985 & w6071);
assign w11940 = w6391 & ~w142;
assign w11941 = ~w142 & ~w4458;
assign w11942 = ~w9909 & ~w12806;
assign w11943 = ~w1166 & ~w13873;
assign w11944 = ~w2009 & ~w6736;
assign w11945 = (w12941 & w117) | (w12941 & w13806) | (w117 & w13806);
assign w11946 = ~w7806 & ~w6338;
assign w11947 = ~w3276 & w3353;
assign w11948 = w4349 & ~w7403;
assign w11949 = ~w7336 & w14075;
assign w11950 = w4558 & w10586;
assign w11951 = w3122 & w12112;
assign w11952 = (w11053 & w3156) | (w11053 & w9774) | (w3156 & w9774);
assign w11953 = ~w1997 & ~w9506;
assign w11954 = ~w2433 & ~w2729;
assign w11955 = ~w2463 & w2259;
assign w11956 = w5715 & ~w5334;
assign w11957 = w9715 & ~w7546;
assign w11958 = w7296 & w6949;
assign w11959 = w7085 & w8018;
assign w11960 = ~w6479 & ~w8664;
assign w11961 = w473 & ~w9465;
assign w11962 = ~w1799 & ~w13323;
assign w11963 = (w653 & w4551) | (w653 & ~w12911) | (w4551 & ~w12911);
assign w11964 = (~w6750 & w2513) | (~w6750 & w9818) | (w2513 & w9818);
assign w11965 = ~w142 & w3727;
assign w11966 = (w7457 & w1739) | (w7457 & w1175) | (w1739 & w1175);
assign w11967 = w11031 & ~w11764;
assign w11968 = w5121 & w2630;
assign w11969 = (~w5783 & w2763) | (~w5783 & w11667) | (w2763 & w11667);
assign w11970 = (w4580 & w14108) | (w4580 & w4339) | (w14108 & w4339);
assign w11971 = w17 & w13955;
assign w11972 = (w7751 & w6521) | (w7751 & ~w8937) | (w6521 & ~w8937);
assign w11973 = (w1849 & w6571) | (w1849 & w12395) | (w6571 & w12395);
assign w11974 = w4138 & w10116;
assign w11975 = (w91 & w9327) | (w91 & w1964) | (w9327 & w1964);
assign w11976 = ~w2864 & ~w9211;
assign w11977 = w10645 & w6064;
assign w11978 = w6459 & w2042;
assign w11979 = (w11580 & w4238) | (w11580 & w14069) | (w4238 & w14069);
assign w11980 = ~w9788 & ~w1062;
assign w11981 = ~w5702 & w12608;
assign w11982 = (w9368 & w5920) | (w9368 & w2132) | (w5920 & w2132);
assign w11983 = w9643 & w13707;
assign w11984 = w3821 & w9528;
assign w11985 = ~w574 & ~w13584;
assign w11986 = w3988 & w9367;
assign w11987 = ~w13895 & ~w1965;
assign w11988 = (w40 & w10462) | (w40 & w4596) | (w10462 & w4596);
assign w11989 = (~w3427 & ~w1087) | (~w3427 & w8063) | (~w1087 & w8063);
assign w11990 = w10545 & w12685;
assign w11991 = ~w13118 & w10376;
assign w11992 = ~w5948 & ~w3727;
assign w11993 = (w10496 & w2187) | (w10496 & w5100) | (w2187 & w5100);
assign w11994 = w8843 & w6278;
assign w11995 = ~w7659 & ~w7691;
assign w11996 = w10308 & ~w1591;
assign w11997 = ~w10477 & ~w11604;
assign w11998 = w13256 & w11117;
assign w11999 = (w378 & w11840) | (w378 & w8822) | (w11840 & w8822);
assign w12000 = w7991 & w5887;
assign w12001 = w8924 & ~w671;
assign w12002 = ~w2317 & w12188;
assign w12003 = w9845 & ~w1141;
assign w12004 = ~w12444 & w8233;
assign w12005 = w4385 & w4187;
assign w12006 = (~w5673 & w13324) | (~w5673 & w2030) | (w13324 & w2030);
assign w12007 = w8738 & w234;
assign w12008 = w5189 & w5327;
assign w12009 = ~w4721 & ~w9102;
assign w12010 = w11496 & ~w1413;
assign w12011 = ~w5660 & ~w11735;
assign w12012 = ~w142 & ~w646;
assign w12013 = w5166 & ~w5549;
assign w12014 = ~w183 & w10393;
assign w12015 = ~w3244 & ~w4294;
assign w12016 = ~w12569 & ~w3253;
assign w12017 = (~w2463 & w7324) | (~w2463 & w14658) | (w7324 & w14658);
assign w12018 = (~w2135 & w12499) | (~w2135 & w10987) | (w12499 & w10987);
assign w12019 = ~w7908 & w12633;
assign w12020 = w439 & ~w7057;
assign w12021 = (w4425 & w13152) | (w4425 & w14339) | (w13152 & w14339);
assign w12022 = w12124 & ~w1955;
assign w12023 = w11680 & ~w12381;
assign w12024 = ~w10402 & ~w12031;
assign w12025 = (~w11551 & w6230) | (~w11551 & w9192) | (w6230 & w9192);
assign w12026 = ~w5555 & ~w14209;
assign w12027 = (~w8100 & w7799) | (~w8100 & w1416) | (w7799 & w1416);
assign w12028 = w8738 & w4890;
assign w12029 = w818 | w5532;
assign w12030 = ~w10119 & w12311;
assign w12031 = (~w4281 & w10446) | (~w4281 & w6782) | (w10446 & w6782);
assign w12032 = w571 & w3586;
assign w12033 = w7794 & w5276;
assign w12034 = (w7227 & w13122) | (w7227 & w9406) | (w13122 & w9406);
assign w12035 = w14396 & w5378;
assign w12036 = (~w5785 & w9139) | (~w5785 & w2445) | (w9139 & w2445);
assign w12037 = (w1949 & ~w6137) | (w1949 & w4624) | (~w6137 & w4624);
assign w12038 = w446 & w11944;
assign w12039 = w473 & w6381;
assign w12040 = (~w6929 & w4478) | (~w6929 & w1615) | (w4478 & w1615);
assign w12041 = ~w5732 & w9227;
assign w12042 = ~w9608 & w29;
assign w12043 = w1803 & w11077;
assign w12044 = ~w6230 & ~w68;
assign w12045 = (~w6700 & w6541) | (~w6700 & w10611) | (w6541 & w10611);
assign w12046 = ~w3956 & ~w343;
assign w12047 = ~w9669 & ~w7501;
assign w12048 = (~w5601 & w9014) | (~w5601 & w5063) | (w9014 & w5063);
assign w12049 = w14382 & w3564;
assign w12050 = ~w2371 & ~w11274;
assign w12051 = ~w1878 & w12021;
assign w12052 = w3251 & w3904;
assign w12053 = ~w9541 & w11487;
assign w12054 = ~w2250 & w9869;
assign w12055 = ~w13793 & ~w6689;
assign w12056 = (w10318 & ~w353) | (w10318 & w9364) | (~w353 & w9364);
assign w12057 = ~w6628 & ~w799;
assign w12058 = w3957 & ~w13733;
assign w12059 = ~w4688 & ~w12516;
assign w12060 = ~w6889 & ~w13565;
assign w12061 = (w884 & w4158) | (w884 & w3322) | (w4158 & w3322);
assign w12062 = ~w8937 & w8876;
assign w12063 = (~w3698 & ~w5490) | (~w3698 & ~w12656) | (~w5490 & ~w12656);
assign w12064 = ~w5294 & ~w5196;
assign w12065 = b62 & a62;
assign w12066 = ~w2597 & ~w341;
assign w12067 = ~w855 & w476;
assign w12068 = w3734 & w142;
assign w12069 = ~w8088 & ~w2394;
assign w12070 = ~w13732 & ~w6903;
assign w12071 = w4093 & w8230;
assign w12072 = ~w5294 & ~w12915;
assign w12073 = ~w14513 & w1807;
assign w12074 = w9170 & w12088;
assign w12075 = ~w4453 & ~w8580;
assign w12076 = (w12662 & w8937) | (w12662 & w13781) | (w8937 & w13781);
assign w12077 = (w9054 & ~w3794) | (w9054 & w2436) | (~w3794 & w2436);
assign w12078 = w5178 & w7645;
assign w12079 = ~w1764 & ~w11147;
assign w12080 = (~w4336 & ~w3242) | (~w4336 & w8616) | (~w3242 & w8616);
assign w12081 = w309 & w5845;
assign w12082 = (~w10699 & w988) | (~w10699 & w10455) | (w988 & w10455);
assign w12083 = ~w5845 & w2698;
assign w12084 = ~w1699 & w5243;
assign w12085 = ~w11313 & ~w11885;
assign w12086 = w8389 & ~w10777;
assign w12087 = ~w372 & w12714;
assign w12088 = w2599 & w7455;
assign w12089 = (~w2445 & w4593) | (~w2445 & w4776) | (w4593 & w4776);
assign w12090 = w4171 & ~w5624;
assign w12091 = ~w9372 & w4286;
assign w12092 = (~w4612 & w7854) | (~w4612 & w13637) | (w7854 & w13637);
assign w12093 = ~w1431 & ~w9932;
assign w12094 = (~w7815 & w8837) | (~w7815 & w6540) | (w8837 & w6540);
assign w12095 = ~w11345 & ~w12908;
assign w12096 = w2975 & w10209;
assign w12097 = ~w5696 & w10551;
assign w12098 = ~w7914 & ~w6716;
assign w12099 = w13222 & ~w8196;
assign w12100 = (~w7296 & w6161) | (~w7296 & ~w13222) | (w6161 & ~w13222);
assign w12101 = w11916 & w5039;
assign w12102 = w5590 & w13619;
assign w12103 = ~w7296 & w4541;
assign w12104 = w13018 & w5372;
assign w12105 = ~w13323 & ~w13793;
assign w12106 = ~w4159 & w11454;
assign w12107 = ~w5754 & ~w2081;
assign w12108 = w2081 & w11049;
assign w12109 = (~w2144 & w5774) | (~w2144 & w9588) | (w5774 & w9588);
assign w12110 = (w6889 & w14141) | (w6889 & w6499) | (w14141 & w6499);
assign w12111 = ~w3453 & ~w733;
assign w12112 = ~w11905 & ~w6281;
assign w12113 = ~w4900 & ~w10381;
assign w12114 = ~w727 & w2444;
assign w12115 = (w6845 & w8314) | (w6845 & w7046) | (w8314 & w7046);
assign w12116 = (w12786 & w12799) | (w12786 & w8228) | (w12799 & w8228);
assign w12117 = (~w7684 & w6623) | (~w7684 & w6572) | (w6623 & w6572);
assign w12118 = w7914 & w801;
assign w12119 = ~w5970 & ~w5551;
assign w12120 = w1166 & w13854;
assign w12121 = ~w13722 & ~w10440;
assign w12122 = ~w1516 & w11236;
assign w12123 = w8975 & w9921;
assign w12124 = ~w5294 & ~w13349;
assign w12125 = ~w9794 & ~w10486;
assign w12126 = ~w922 & ~w6062;
assign w12127 = (~w13802 & ~w8769) | (~w13802 & w3332) | (~w8769 & w3332);
assign w12128 = ~w1828 & ~w5701;
assign w12129 = ~w1914 & w8388;
assign w12130 = ~w7800 & ~w12283;
assign w12131 = ~w10523 & ~w3786;
assign w12132 = (w14061 & ~w6563) | (w14061 & w4945) | (~w6563 & w4945);
assign w12133 = w12353 & w6169;
assign w12134 = ~w922 & w6716;
assign w12135 = w8085 & w77;
assign w12136 = ~w6888 & ~w11940;
assign w12137 = ~w1608 & w14195;
assign w12138 = (w378 & w875) | (w378 & w5391) | (w875 & w5391);
assign w12139 = ~w11571 & w3763;
assign w12140 = w2475 & w4981;
assign w12141 = w11364 & ~w11142;
assign w12142 = w11236 & w7381;
assign w12143 = w10423 & w12398;
assign w12144 = ~w8100 & w2470;
assign w12145 = (w420 & w9169) | (w420 & w4238) | (w9169 & w4238);
assign w12146 = w7697 & w6624;
assign w12147 = w4089 & w5393;
assign w12148 = ~b27 & ~a27;
assign w12149 = (w12312 & w11690) | (w12312 & w2665) | (w11690 & w2665);
assign w12150 = w7722 & w13114;
assign w12151 = w7645 & ~w8544;
assign w12152 = (w7951 & w1639) | (w7951 & w7116) | (w1639 & w7116);
assign w12153 = ~w9747 & w1735;
assign w12154 = w2928 & w9564;
assign w12155 = (~w10699 & w11225) | (~w10699 & w11234) | (w11225 & w11234);
assign w12156 = (~w5160 & w3352) | (~w5160 & w5245) | (w3352 & w5245);
assign w12157 = w1221 & ~w7490;
assign w12158 = ~w607 & w646;
assign w12159 = (w11708 & ~w8427) | (w11708 & w3809) | (~w8427 & w3809);
assign w12160 = w2410 & w5788;
assign w12161 = w5667 & w12213;
assign w12162 = ~w572 & w6477;
assign w12163 = ~w9136 & w12683;
assign w12164 = w7794 & w14493;
assign w12165 = ~w1439 & ~w3255;
assign w12166 = (~w8277 & w11209) | (~w8277 & w12106) | (w11209 & w12106);
assign w12167 = w3251 & w12642;
assign w12168 = w852 & ~w9748;
assign w12169 = w10378 & w2516;
assign w12170 = ~b56 & ~a56;
assign w12171 = (~w14395 & w14141) | (~w14395 & w3854) | (w14141 & w3854);
assign w12172 = (w10707 & w6771) | (w10707 & ~w3885) | (w6771 & ~w3885);
assign w12173 = w9138 & w3361;
assign w12174 = ~w4883 & ~w1381;
assign w12175 = w4167 & ~w1794;
assign w12176 = w7704 & ~w3780;
assign w12177 = w2762 & ~w8691;
assign w12178 = w6143 & w6414;
assign w12179 = (~w9305 & w2768) | (~w9305 & w7323) | (w2768 & w7323);
assign w12180 = (w9457 & w3258) | (w9457 & ~w8584) | (w3258 & ~w8584);
assign w12181 = w9949 & ~w5108;
assign w12182 = ~w11434 & w1687;
assign w12183 = (w9305 & w5111) | (w9305 & w11113) | (w5111 & w11113);
assign w12184 = ~w9708 & ~w10688;
assign w12185 = w12615 & ~w8614;
assign w12186 = w10277 & ~w12942;
assign w12187 = (w10708 & ~w13282) | (w10708 & w5226) | (~w13282 & w5226);
assign w12188 = ~w1563 & w3661;
assign w12189 = ~w4214 & w8439;
assign w12190 = (w14600 & w2234) | (w14600 & w4703) | (w2234 & w4703);
assign w12191 = w12170 & ~w12662;
assign w12192 = w12464 & ~w4032;
assign w12193 = w10949 & w11375;
assign w12194 = w5778 & w9211;
assign w12195 = w11948 & w12442;
assign w12196 = (w605 & w310) | (w605 & w9206) | (w310 & w9206);
assign w12197 = (~w12215 & w5458) | (~w12215 & w1044) | (w5458 & w1044);
assign w12198 = w12197 | w2071;
assign w12199 = (w6542 & w10245) | (w6542 & w10055) | (w10245 & w10055);
assign w12200 = (~w1589 & ~w13219) | (~w1589 & w944) | (~w13219 & w944);
assign w12201 = (~w4379 & w12029) | (~w4379 & w4683) | (w12029 & w4683);
assign w12202 = (~w4989 & w14664) | (~w4989 & w2894) | (w14664 & w2894);
assign w12203 = w12463 & ~w4453;
assign w12204 = (~w13206 & w7782) | (~w13206 & w10351) | (w7782 & w10351);
assign w12205 = (w12868 & w12980) | (w12868 & w1) | (w12980 & w1);
assign w12206 = (~w13620 & ~w953) | (~w13620 & w10297) | (~w953 & w10297);
assign w12207 = ~w6912 & w3552;
assign w12208 = (~w7168 & w12920) | (~w7168 & w1284) | (w12920 & w1284);
assign w12209 = (~w235 & w5506) | (~w235 & w8778) | (w5506 & w8778);
assign w12210 = ~w8183 & w11934;
assign w12211 = w3036 & w8047;
assign w12212 = (~w6379 & w9695) | (~w6379 & w11111) | (w9695 & w11111);
assign w12213 = ~w11391 & w6689;
assign w12214 = (~w2701 & w12308) | (~w2701 & w6031) | (w12308 & w6031);
assign w12215 = (w6637 & w237) | (w6637 & w5530) | (w237 & w5530);
assign w12216 = w3289 & w8056;
assign w12217 = w1838 & ~w11861;
assign w12218 = (~w6802 & w7289) | (~w6802 & w3975) | (w7289 & w3975);
assign w12219 = ~w8330 & w8465;
assign w12220 = ~w13940 & w4042;
assign w12221 = w10045 & w69;
assign w12222 = (~w8171 & w4182) | (~w8171 & ~w4656) | (w4182 & ~w4656);
assign w12223 = ~w13839 & ~w9646;
assign w12224 = ~w536 & w14129;
assign w12225 = w9759 & w6382;
assign w12226 = (w1267 & w5440) | (w1267 & w5627) | (w5440 & w5627);
assign w12227 = (w3508 & w10462) | (w3508 & w5003) | (w10462 & w5003);
assign w12228 = w4167 & w3873;
assign w12229 = w2425 & w9748;
assign w12230 = ~w2574 & ~w4291;
assign w12231 = (~w6381 & w11261) | (~w6381 & w448) | (w11261 & w448);
assign w12232 = w11364 & w2086;
assign w12233 = (w13531 & w12614) | (w13531 & w7380) | (w12614 & w7380);
assign w12234 = (w7999 & w7522) | (w7999 & w2240) | (w7522 & w2240);
assign w12235 = ~w4921 & w4955;
assign w12236 = ~w9087 & ~w11810;
assign w12237 = (w6212 & ~w5566) | (w6212 & w9611) | (~w5566 & w9611);
assign w12238 = (w3427 & w5562) | (w3427 & w4498) | (w5562 & w4498);
assign w12239 = (w2544 & w3825) | (w2544 & ~w5746) | (w3825 & ~w5746);
assign w12240 = ~w8338 & ~w11965;
assign w12241 = w11702 & ~w12841;
assign w12242 = ~w4213 & w6716;
assign w12243 = ~w12240 & w4190;
assign w12244 = ~w449 & w2128;
assign w12245 = w5783 & w11781;
assign w12246 = ~w724 & w6343;
assign w12247 = w5014 & ~w13256;
assign w12248 = w2933 & ~w10514;
assign w12249 = w7829 & ~w5775;
assign w12250 = w8027 & w10290;
assign w12251 = w9541 & w11902;
assign w12252 = ~w12421 & w9908;
assign w12253 = ~w3549 & ~w12119;
assign w12254 = (~w13197 & w9078) | (~w13197 & w6581) | (w9078 & w6581);
assign w12255 = ~w10460 & w4734;
assign w12256 = ~w6838 & ~w9313;
assign w12257 = (~w8937 & w3187) | (~w8937 & w9042) | (w3187 & w9042);
assign w12258 = w12716 & w5360;
assign w12259 = w3098 & w3044;
assign w12260 = w11177 & w174;
assign w12261 = (w3039 & w12499) | (w3039 & w10717) | (w12499 & w10717);
assign w12262 = w10721 & w7148;
assign w12263 = (~w8692 & w8324) | (~w8692 & w3931) | (w8324 & w3931);
assign w12264 = ~w13880 & w4036;
assign w12265 = (~w5482 & w13749) | (~w5482 & ~w5105) | (w13749 & ~w5105);
assign w12266 = w4870 & w13757;
assign w12267 = w7132 & w2398;
assign w12268 = (~w10768 & ~w5664) | (~w10768 & w3848) | (~w5664 & w3848);
assign w12269 = w13560 & w3844;
assign w12270 = ~w10837 & ~w11752;
assign w12271 = ~w12012 & ~w7661;
assign w12272 = (w2788 & w11138) | (w2788 & w1901) | (w11138 & w1901);
assign w12273 = ~w2135 & w7645;
assign w12274 = ~w4341 & ~w7250;
assign w12275 = (~w6267 & w7139) | (~w6267 & w14104) | (w7139 & w14104);
assign w12276 = ~w639 & w12178;
assign w12277 = (~w11261 & w5690) | (~w11261 & w13884) | (w5690 & w13884);
assign w12278 = ~w1048 & w6098;
assign w12279 = ~w2692 | w5694;
assign w12280 = ~w10182 & w5978;
assign w12281 = (w8637 & w2415) | (w8637 & ~w10613) | (w2415 & ~w10613);
assign w12282 = w1297 & ~w4177;
assign w12283 = w607 & ~w4458;
assign w12284 = ~w8791 & ~w10669;
assign w12285 = ~w7120 & ~w14102;
assign w12286 = (~w7515 & w4701) | (~w7515 & w2246) | (w4701 & w2246);
assign w12287 = (w59 & w1178) | (w59 & ~w4929) | (w1178 & ~w4929);
assign w12288 = (w7813 & w6859) | (w7813 & w4904) | (w6859 & w4904);
assign w12289 = ~w14140 & w12592;
assign w12290 = w7668 & ~w5664;
assign w12291 = (w1489 & w6373) | (w1489 & w9337) | (w6373 & w9337);
assign w12292 = w11287 & w958;
assign w12293 = ~w4756 & ~w235;
assign w12294 = (~w9465 & w2493) | (~w9465 & w11961) | (w2493 & w11961);
assign w12295 = w10274 & w138;
assign w12296 = (w13227 & w21) | (w13227 & w11296) | (w21 & w11296);
assign w12297 = ~w3209 & ~w10200;
assign w12298 = w5626 & ~w12891;
assign w12299 = ~w7414 & ~w6929;
assign w12300 = ~w607 & w13323;
assign w12301 = (~w2445 & w6976) | (~w2445 & w3541) | (w6976 & w3541);
assign w12302 = (w7914 & w10191) | (w7914 & w7766) | (w10191 & w7766);
assign w12303 = ~w3486 & w5020;
assign w12304 = ~w12240 & ~w2142;
assign w12305 = (w1053 & w1916) | (w1053 & w5206) | (w1916 & w5206);
assign w12306 = ~w7001 & ~w4458;
assign w12307 = (w10276 & w2311) | (w10276 & w13904) | (w2311 & w13904);
assign w12308 = ~w8045 & ~w2701;
assign w12309 = w9925 & w11405;
assign w12310 = ~w7390 & w7458;
assign w12311 = w4791 & ~w8992;
assign w12312 = (w11013 & ~w5545) | (w11013 & ~w13562) | (~w5545 & ~w13562);
assign w12313 = w14302 & ~w2428;
assign w12314 = (w8149 & w3866) | (w8149 & w304) | (w3866 & w304);
assign w12315 = b19 & a19;
assign w12316 = (~w3550 & w6853) | (~w3550 & w14013) | (w6853 & w14013);
assign w12317 = ~w7190 & ~w9453;
assign w12318 = w12664 & w7754;
assign w12319 = ~w13810 & w6261;
assign w12320 = w1257 & ~w2923;
assign w12321 = ~w11395 & ~w8512;
assign w12322 = w8900 & w12567;
assign w12323 = ~w1924 & ~w14609;
assign w12324 = (w2485 & w6893) | (w2485 & ~w4044) | (w6893 & ~w4044);
assign w12325 = (~w13222 & w8718) | (~w13222 & w8002) | (w8718 & w8002);
assign w12326 = w7645 & ~w5768;
assign w12327 = w2817 & w7085;
assign w12328 = w4032 & w9015;
assign w12329 = ~w12468 & ~w11681;
assign w12330 = ~w4312 & ~w14526;
assign w12331 = (w5664 & w11403) | (w5664 & w7657) | (w11403 & w7657);
assign w12332 = (w12568 & w4746) | (w12568 & w8217) | (w4746 & w8217);
assign w12333 = w10676 & w9871;
assign w12334 = (~w11488 & ~w9748) | (~w11488 & w10498) | (~w9748 & w10498);
assign w12335 = w5395 & ~w1712;
assign w12336 = (w1344 & w3336) | (w1344 & w2362) | (w3336 & w2362);
assign w12337 = (w4204 & w4756) | (w4204 & w2047) | (w4756 & w2047);
assign w12338 = w12464 & ~w5867;
assign w12339 = ~w12271 & w2680;
assign w12340 = w9211 & w8713;
assign w12341 = ~w7724 & ~w7451;
assign w12342 = (~w2493 & w2463) | (~w2493 & w4329) | (w2463 & w4329);
assign w12343 = w5785 & ~w11117;
assign w12344 = ~w14280 & ~w10853;
assign w12345 = ~w8740 & w14543;
assign w12346 = w4213 & w13531;
assign w12347 = ~w7726 & w3575;
assign w12348 = ~w13141 & ~w3747;
assign w12349 = (~w4050 & w7862) | (~w4050 & w12100) | (w7862 & w12100);
assign w12350 = (w3039 & ~w5294) | (w3039 & w7324) | (~w5294 & w7324);
assign w12351 = (w9305 & w6748) | (w9305 & w12780) | (w6748 & w12780);
assign w12352 = ~w441 & ~w10355;
assign w12353 = (w13197 & ~w7599) | (w13197 & w9476) | (~w7599 & w9476);
assign w12354 = (~w318 & w8814) | (~w318 & ~w10590) | (w8814 & ~w10590);
assign w12355 = ~w3963 & w988;
assign w12356 = ~w3777 & ~w13547;
assign w12357 = ~w13095 & ~w10483;
assign w12358 = ~w2008 & w14045;
assign w12359 = ~w5560 & ~w12315;
assign w12360 = ~w12512 & ~w7556;
assign w12361 = w14107 & w2769;
assign w12362 = ~w11855 & ~w12614;
assign w12363 = w9412 & ~w3568;
assign w12364 = w10720 & ~w8025;
assign w12365 = w829 & ~w10704;
assign w12366 = w14582 & ~w11030;
assign w12367 = ~w2019 & ~w2622;
assign w12368 = (~w5664 & w6929) | (~w5664 & w5275) | (w6929 & w5275);
assign w12369 = w14257 & w13047;
assign w12370 = ~w7305 & ~w2941;
assign w12371 = ~b95 & ~a95;
assign w12372 = ~w1397 & ~w11502;
assign w12373 = w4845 & w7593;
assign w12374 = (w852 & w4099) | (w852 & w6839) | (w4099 & w6839);
assign w12375 = w830 & w9641;
assign w12376 = (w4149 & w3055) | (w4149 & w1583) | (w3055 & w1583);
assign w12377 = ~w13839 & w3175;
assign w12378 = ~w5754 & ~w12095;
assign w12379 = w4836 & w2335;
assign w12380 = (w9452 & w2360) | (w9452 & w10134) | (w2360 & w10134);
assign w12381 = (~w9748 & w12354) | (~w9748 & w1436) | (w12354 & w1436);
assign w12382 = ~w13189 & ~w2509;
assign w12383 = ~w10833 & ~w10590;
assign w12384 = w5156 & w5704;
assign w12385 = w357 & w13941;
assign w12386 = w3020 & ~w8834;
assign w12387 = ~w1568 & w12270;
assign w12388 = w14015 & w2729;
assign w12389 = ~w11284 & ~w3633;
assign w12390 = ~w1474 & w646;
assign w12391 = ~w9607 & w11583;
assign w12392 = (w4103 & w4275) | (w4103 & w12848) | (w4275 & w12848);
assign w12393 = w2101 & w10556;
assign w12394 = w8513 & w10365;
assign w12395 = (~w9591 & ~w13292) | (~w9591 & ~w11091) | (~w13292 & ~w11091);
assign w12396 = w1824 & w3289;
assign w12397 = ~w3914 & w894;
assign w12398 = ~b65 & ~a65;
assign w12399 = w12642 & ~w8104;
assign w12400 = ~w4458 & ~w9418;
assign w12401 = (~w10483 & w8886) | (~w10483 & w5788) | (w8886 & w5788);
assign w12402 = (w11708 & w2226) | (w11708 & w1749) | (w2226 & w1749);
assign w12403 = ~w6795 & w6230;
assign w12404 = w1830 & ~w13057;
assign w12405 = (~w2698 & w7488) | (~w2698 & w13042) | (w7488 & w13042);
assign w12406 = (~w9305 & ~w6849) | (~w9305 & ~w11522) | (~w6849 & ~w11522);
assign w12407 = (w3427 & w12825) | (w3427 & w9835) | (w12825 & w9835);
assign w12408 = (w12951 & w3641) | (w12951 & w14237) | (w3641 & w14237);
assign w12409 = (w11724 & w2689) | (w11724 & w2025) | (w2689 & w2025);
assign w12410 = (~w5952 & w3915) | (~w5952 & w3167) | (w3915 & w3167);
assign w12411 = (~w8483 & ~w12189) | (~w8483 & w4654) | (~w12189 & w4654);
assign w12412 = (w13587 & w13868) | (w13587 & w1917) | (w13868 & w1917);
assign w12413 = (w11174 & w2718) | (w11174 & w11972) | (w2718 & w11972);
assign w12414 = w5481 & w8121;
assign w12415 = ~w8435 & ~w11544;
assign w12416 = ~w936 & ~w7530;
assign w12417 = ~w3098 & w7794;
assign w12418 = (~w3963 & w110) | (~w3963 & w9294) | (w110 & w9294);
assign w12419 = w14054 & ~w12908;
assign w12420 = (~w10590 & w13587) | (~w10590 & w13679) | (w13587 & w13679);
assign w12421 = w1800 & ~w3194;
assign w12422 = ~w7488 & w10111;
assign w12423 = w2111 & w4759;
assign w12424 = ~w5195 & ~w13373;
assign w12425 = ~w9789 & w588;
assign w12426 = w13839 & ~w5069;
assign w12427 = (w4324 & w4650) | (w4324 & w7332) | (w4650 & w7332);
assign w12428 = (~w13902 & ~w3645) | (~w13902 & w2785) | (~w3645 & w2785);
assign w12429 = b43 & a43;
assign w12430 = (w12857 & w11058) | (w12857 & w7676) | (w11058 & w7676);
assign w12431 = ~w1125 & ~w5496;
assign w12432 = ~w9927 & w3727;
assign w12433 = ~w2013 & ~w5047;
assign w12434 = w6599 & w6534;
assign w12435 = w8707 & ~w5518;
assign w12436 = (~w10052 & ~w7077) | (~w10052 & w5662) | (~w7077 & w5662);
assign w12437 = w8713 & w6592;
assign w12438 = b77 & a77;
assign w12439 = (w11500 & ~w9813) | (w11500 & w11613) | (~w9813 & w11613);
assign w12440 = ~w9583 & ~w12893;
assign w12441 = w8847 & w2286;
assign w12442 = ~w13233 & ~w7181;
assign w12443 = w8356 & w3904;
assign w12444 = ~w4246 & ~w13185;
assign w12445 = (w4425 & w12499) | (w4425 & w13512) | (w12499 & w13512);
assign w12446 = w2381 & w3615;
assign w12447 = (w12398 & w1840) | (w12398 & w12143) | (w1840 & w12143);
assign w12448 = ~w9652 & w7840;
assign w12449 = w12135 & w13924;
assign w12450 = ~w13880 & w2388;
assign w12451 = ~w11396 & w2809;
assign w12452 = ~w6247 & ~w4898;
assign w12453 = ~w2784 & ~w8749;
assign w12454 = ~w3354 & w11414;
assign w12455 = w9057 & w13452;
assign w12456 = (w3144 & w2978) | (w3144 & ~w3017) | (w2978 & ~w3017);
assign w12457 = (~w7693 & w4174) | (~w7693 & w5246) | (w4174 & w5246);
assign w12458 = ~w404 & w9133;
assign w12459 = ~w9141 & w4848;
assign w12460 = ~w11745 & ~w1474;
assign w12461 = ~w7383 & ~w10112;
assign w12462 = ~w11988 & ~w4597;
assign w12463 = ~b18 & ~a18;
assign w12464 = w7376 & w7794;
assign w12465 = ~w7359 & ~w13417;
assign w12466 = w1607 & w1274;
assign w12467 = ~w2059 & ~w1664;
assign w12468 = ~w10435 & w13537;
assign w12469 = ~w9548 & w3467;
assign w12470 = (w4127 & ~w1712) | (w4127 & w7877) | (~w1712 & w7877);
assign w12471 = w1387 & w5792;
assign w12472 = ~w4600 & w5190;
assign w12473 = w9944 & w4283;
assign w12474 = w9021 & ~w7215;
assign w12475 = w5556 & w4541;
assign w12476 = (w9095 & w5752) | (w9095 & w8614) | (w5752 & w8614);
assign w12477 = w11193 & w5335;
assign w12478 = (w7080 & w13324) | (w7080 & w7883) | (w13324 & w7883);
assign w12479 = ~w7889 & ~w10941;
assign w12480 = ~w4678 & w4157;
assign w12481 = b98 & a98;
assign w12482 = ~w3751 & ~w5108;
assign w12483 = w7085 & w5213;
assign w12484 = w10217 | w9921;
assign w12485 = ~w4373 & w1215;
assign w12486 = w2569 & w6230;
assign w12487 = w13521 & w1540;
assign w12488 = w4314 & w9158;
assign w12489 = (~w3963 & ~w7154) | (~w3963 & w3729) | (~w7154 & w3729);
assign w12490 = ~w12553 & ~w10875;
assign w12491 = (w876 & w3306) | (w876 & w5367) | (w3306 & w5367);
assign w12492 = ~w12575 & w4417;
assign w12493 = w309 & w1016;
assign w12494 = (w8405 & w2810) | (w8405 & w8903) | (w2810 & w8903);
assign w12495 = (w1910 & w1190) | (w1910 & ~w11168) | (w1190 & ~w11168);
assign w12496 = ~w2739 & ~w13083;
assign w12497 = ~w230 & ~w5831;
assign w12498 = (w1746 & w11268) | (w1746 & ~w7693) | (w11268 & ~w7693);
assign w12499 = w2194 & ~w401;
assign w12500 = w10407 & w5507;
assign w12501 = (~w8580 & w5671) | (~w8580 & w14472) | (w5671 & w14472);
assign w12502 = w11085 & w2305;
assign w12503 = w10676 & w11810;
assign w12504 = ~w6800 & w12353;
assign w12505 = w3215 & ~w8389;
assign w12506 = b125 & a125;
assign w12507 = w4894 & ~w9360;
assign w12508 = w14203 & w6881;
assign w12509 = ~w5734 & ~w5264;
assign w12510 = w11317 & w578;
assign w12511 = ~w7187 & ~w11946;
assign w12512 = ~w14664 & w11610;
assign w12513 = (w2309 & w14442) | (w2309 & ~w8076) | (w14442 & ~w8076);
assign w12514 = w10075 & w8389;
assign w12515 = w12642 & w11764;
assign w12516 = ~w14639 & ~w8013;
assign w12517 = (~w302 & w7511) | (~w302 & w9967) | (w7511 & w9967);
assign w12518 = ~w12330 & w10872;
assign w12519 = w6130 & ~w5409;
assign w12520 = ~w7437 & ~w10704;
assign w12521 = (w302 & w864) | (w302 & w9562) | (w864 & w9562);
assign w12522 = ~w9258 & w10012;
assign w12523 = (w9724 & w1770) | (w9724 & w1114) | (w1770 & w1114);
assign w12524 = w1353 | w11708;
assign w12525 = ~w13713 & w3734;
assign w12526 = ~w5620 & w3219;
assign w12527 = (w6970 & w8821) | (w6970 & ~w9364) | (w8821 & ~w9364);
assign w12528 = ~w2159 & w12893;
assign w12529 = (~w7630 & w2247) | (~w7630 & w14093) | (w2247 & w14093);
assign w12530 = w7070 & w6815;
assign w12531 = (w227 & w1190) | (w227 & w9989) | (w1190 & w9989);
assign w12532 = ~w13450 & w12739;
assign w12533 = (~w4050 & w5289) | (~w4050 & w12912) | (w5289 & w12912);
assign w12534 = ~w1062 & w3963;
assign w12535 = w607 & ~w5761;
assign w12536 = w7133 & ~w8097;
assign w12537 = (~w3798 & w6310) | (~w3798 & ~w9364) | (w6310 & ~w9364);
assign w12538 = (w3526 & w5428) | (w3526 & w3432) | (w5428 & w3432);
assign w12539 = w12121 & w8827;
assign w12540 = ~w5790 & w11934;
assign w12541 = w11601 | w9644;
assign w12542 = ~w3885 & w9211;
assign w12543 = w9087 & w5767;
assign w12544 = ~w4547 & w13059;
assign w12545 = ~w7490 & ~w11560;
assign w12546 = ~w9747 & w8212;
assign w12547 = w894 & ~w6542;
assign w12548 = (w3427 & ~w5912) | (w3427 & w11382) | (~w5912 & w11382);
assign w12549 = (w7082 & w658) | (w7082 & w8856) | (w658 & w8856);
assign w12550 = ~w7222 & ~w10646;
assign w12551 = (w6722 & ~w2852) | (w6722 & w2596) | (~w2852 & w2596);
assign w12552 = ~w7376 & w884;
assign w12553 = w3550 & w14625;
assign w12554 = ~w13148 & ~w6196;
assign w12555 = (~w8315 & ~w7893) | (~w8315 & ~w12888) | (~w7893 & ~w12888);
assign w12556 = ~w533 & ~w3904;
assign w12557 = w1166 & w5693;
assign w12558 = ~w1054 & w2018;
assign w12559 = w8306 & ~w9788;
assign w12560 = w3963 & ~w1406;
assign w12561 = w10676 & w12856;
assign w12562 = (w3040 & w9982) | (w3040 & ~w9754) | (w9982 & ~w9754);
assign w12563 = w2698 & ~w12550;
assign w12564 = w12240 & w14227;
assign w12565 = (w1721 & w7156) | (w1721 & ~w14182) | (w7156 & ~w14182);
assign w12566 = ~w11038 & ~w1798;
assign w12567 = w2159 & w5767;
assign w12568 = (w14417 & w4511) | (w14417 & w8614) | (w4511 & w8614);
assign w12569 = w12656 & w14395;
assign w12570 = (w4328 & ~w13201) | (w4328 & w8668) | (~w13201 & w8668);
assign w12571 = w11033 & ~w13521;
assign w12572 = ~w10435 & w13286;
assign w12573 = w3740 & ~w7374;
assign w12574 = w4627 & w6266;
assign w12575 = ~w3215 & ~w13733;
assign w12576 = (~w2168 & w13184) | (~w2168 & w9924) | (w13184 & w9924);
assign w12577 = ~w4240 & ~w7828;
assign w12578 = w10300 & ~w7154;
assign w12579 = ~w8432 & ~w3414;
assign w12580 = (~w13685 & w202) | (~w13685 & w1427) | (w202 & w1427);
assign w12581 = (~w3019 & w11443) | (~w3019 & w11372) | (w11443 & w11372);
assign w12582 = ~w6233 & w5493;
assign w12583 = ~w11261 & w510;
assign w12584 = w2656 & w11350;
assign w12585 = ~w4276 & w12005;
assign w12586 = ~w132 & ~w8457;
assign w12587 = ~w9910 & ~w11631;
assign w12588 = (~w10917 & w9655) | (~w10917 & ~w4511) | (w9655 & ~w4511);
assign w12589 = (~w8171 & w6651) | (~w8171 & w7543) | (w6651 & w7543);
assign w12590 = w4262 & ~w722;
assign w12591 = (w3427 & w9552) | (w3427 & w7096) | (w9552 & w7096);
assign w12592 = w1171 & w13535;
assign w12593 = (w13603 & ~w1352) | (w13603 & w13466) | (~w1352 & w13466);
assign w12594 = w7808 & w7670;
assign w12595 = ~w10605 & w2374;
assign w12596 = w9972 & ~w3906;
assign w12597 = (w7295 & w4399) | (w7295 & ~w235) | (w4399 & ~w235);
assign w12598 = (~w14504 & w12121) | (~w14504 & w8711) | (w12121 & w8711);
assign w12599 = ~w11586 & w12545;
assign w12600 = (w272 & ~w7434) | (w272 & w8706) | (~w7434 & w8706);
assign w12601 = (w4279 & w8494) | (w4279 & w4861) | (w8494 & w4861);
assign w12602 = (~w2168 & ~w5748) | (~w2168 & w13783) | (~w5748 & w13783);
assign w12603 = (~w10781 & w6330) | (~w10781 & w14377) | (w6330 & w14377);
assign w12604 = b101 & a101;
assign w12605 = (w2652 & w8695) | (w2652 & ~w9034) | (w8695 & ~w9034);
assign w12606 = ~w7452 & ~w4835;
assign w12607 = w8234 & w14326;
assign w12608 = ~w1563 & ~w1263;
assign w12609 = ~w12463 & ~w5560;
assign w12610 = (w1671 & w12674) | (w1671 & w8322) | (w12674 & w8322);
assign w12611 = w8328 & ~w1712;
assign w12612 = ~w5294 & w1821;
assign w12613 = b53 & w1712;
assign w12614 = ~w5836 & ~w9740;
assign w12615 = (~w1016 & w7296) | (~w1016 & w6495) | (w7296 & w6495);
assign w12616 = w6427 & w4627;
assign w12617 = ~w6442 & w13796;
assign w12618 = w3175 & ~w10108;
assign w12619 = (~w12065 & w7296) | (~w12065 & w1536) | (w7296 & w1536);
assign w12620 = ~w9226 & ~w7722;
assign w12621 = ~w7022 & ~w12359;
assign w12622 = ~w12664 & w9211;
assign w12623 = ~w13882 & ~w2015;
assign w12624 = (~w4207 & w10116) | (~w4207 & w1986) | (w10116 & w1986);
assign w12625 = ~w2175 & w11784;
assign w12626 = w13610 & ~w10722;
assign w12627 = (~w13306 & w4952) | (~w13306 & ~w9877) | (w4952 & ~w9877);
assign w12628 = w7645 & ~w1628;
assign w12629 = w9614 & w14389;
assign w12630 = w5936 & ~w9613;
assign w12631 = (~w9880 & ~w1885) | (~w9880 & w4537) | (~w1885 & w4537);
assign w12632 = (~w9038 & w4278) | (~w9038 & w7517) | (w4278 & w7517);
assign w12633 = ~w4497 & ~w9445;
assign w12634 = ~w2212 & w12684;
assign w12635 = (w2225 & w12009) | (w2225 & w12921) | (w12009 & w12921);
assign w12636 = ~w1654 & w7852;
assign w12637 = w5532 & w8512;
assign w12638 = w1503 & ~w2939;
assign w12639 = (w7152 & w3604) | (w7152 & w8559) | (w3604 & w8559);
assign w12640 = (w59 & w1178) | (w59 & ~w7266) | (w1178 & ~w7266);
assign w12641 = (~w12406 & w13212) | (~w12406 & w14606) | (w13212 & w14606);
assign w12642 = ~w7369 & ~w7681;
assign w12643 = ~w14311 & ~w3578;
assign w12644 = ~w6682 & w6082;
assign w12645 = (w12569 & w11482) | (w12569 & w1217) | (w11482 & w1217);
assign w12646 = w9708 & w2272;
assign w12647 = w10256 & ~w11117;
assign w12648 = w6436 & ~w6500;
assign w12649 = (w3124 & ~w11272) | (w3124 & w13840) | (~w11272 & w13840);
assign w12650 = (~w10339 & ~w5070) | (~w10339 & w7362) | (~w5070 & w7362);
assign w12651 = (w8168 & w7843) | (w8168 & w10456) | (w7843 & w10456);
assign w12652 = ~w8104 & ~w6134;
assign w12653 = (w5483 & w4123) | (w5483 & w158) | (w4123 & w158);
assign w12654 = ~w7591 & w12715;
assign w12655 = ~w13804 & w11390;
assign w12656 = ~w13531 & ~w12662;
assign w12657 = (w11983 & w14363) | (w11983 & w84) | (w14363 & w84);
assign w12658 = ~w1840 & ~w5755;
assign w12659 = (~w9305 & w373) | (~w9305 & w8794) | (w373 & w8794);
assign w12660 = ~w12103 & ~w10447;
assign w12661 = (w6276 & w11439) | (w6276 & w13253) | (w11439 & w13253);
assign w12662 = b57 & a57;
assign w12663 = ~w12003 & w8145;
assign w12664 = w13902 & ~w3159;
assign w12665 = ~w1799 & ~w4458;
assign w12666 = w10700 & w6717;
assign w12667 = w11357 & w3062;
assign w12668 = ~w4512 & w2459;
assign w12669 = ~w12662 & ~w8362;
assign w12670 = (~w3334 & ~w14355) | (~w3334 & ~w9096) | (~w14355 & ~w9096);
assign w12671 = ~w4700 & w12642;
assign w12672 = w4452 & w7759;
assign w12673 = ~w10309 & ~w8120;
assign w12674 = (~w4709 & w6207) | (~w4709 & w13975) | (w6207 & w13975);
assign w12675 = ~w1737 & ~w5858;
assign w12676 = w10599 & w11335;
assign w12677 = w6167 & w1656;
assign w12678 = w13393 & w10065;
assign w12679 = ~w12486 & ~w10679;
assign w12680 = w11487 & ~w12614;
assign w12681 = ~w2164 & ~w1719;
assign w12682 = (w5742 & w13122) | (w5742 & w9384) | (w13122 & w9384);
assign w12683 = ~w8525 & w241;
assign w12684 = ~w10639 & w7300;
assign w12685 = ~b16 & ~a16;
assign w12686 = w1563 & w5406;
assign w12687 = ~w6579 & w6390;
assign w12688 = (w6423 & w13315) | (w6423 & w9891) | (w13315 & w9891);
assign w12689 = w12216 & ~w4504;
assign w12690 = ~w5294 & ~w4878;
assign w12691 = w7138 & w4244;
assign w12692 = (w8459 & ~w6101) | (w8459 & w8361) | (~w6101 & w8361);
assign w12693 = ~w9616 & ~w7886;
assign w12694 = (w857 & w1960) | (w857 & w14458) | (w1960 & w14458);
assign w12695 = (~w6500 & w4939) | (~w6500 & w4857) | (w4939 & w4857);
assign w12696 = (~w9032 & w7782) | (~w9032 & w4817) | (w7782 & w4817);
assign w12697 = w607 & w3427;
assign w12698 = ~w10082 & ~w5948;
assign w12699 = ~w12003 & w3185;
assign w12700 = (w3550 & w5850) | (w3550 & w13891) | (w5850 & w13891);
assign w12701 = w761 & w13468;
assign w12702 = ~w13526 & w13281;
assign w12703 = ~w4050 & w64;
assign w12704 = (w1563 & w913) | (w1563 & w8709) | (w913 & w8709);
assign w12705 = ~w5282 & w14614;
assign w12706 = (w4692 & w6634) | (w4692 & ~w9749) | (w6634 & ~w9749);
assign w12707 = ~w5294 & w14390;
assign w12708 = ~w3079 & ~w6350;
assign w12709 = ~w13610 & w8277;
assign w12710 = (w2941 & w4902) | (w2941 & w6975) | (w4902 & w6975);
assign w12711 = w12464 & w10675;
assign w12712 = (w10773 & w613) | (w10773 & w11729) | (w613 & w11729);
assign w12713 = (w9015 & ~w12464) | (w9015 & w6520) | (~w12464 & w6520);
assign w12714 = ~w11361 & ~w9949;
assign w12715 = w9679 & ~w4325;
assign w12716 = ~w10754 & ~w2323;
assign w12717 = ~w13995 & w1981;
assign w12718 = w14547 & ~w888;
assign w12719 = (w1455 & w12771) | (w1455 & w4756) | (w12771 & w4756);
assign w12720 = ~w8785 & ~w2081;
assign w12721 = ~w4539 & w7820;
assign w12722 = w9021 & ~w13007;
assign w12723 = w2101 & ~w5761;
assign w12724 = w12893 & w14486;
assign w12725 = (w815 & w14290) | (w815 & w11806) | (w14290 & w11806);
assign w12726 = (~w12060 & w13324) | (~w12060 & w2679) | (w13324 & w2679);
assign w12727 = w11805 & ~w12790;
assign w12728 = w5830 & ~w13925;
assign w12729 = (~w9012 & w6728) | (~w9012 & w5465) | (w6728 & w5465);
assign w12730 = w7376 & w2701;
assign w12731 = ~w3759 & w1681;
assign w12732 = ~w6190 & ~w10082;
assign w12733 = w739 & ~w8726;
assign w12734 = ~w10245 & w5516;
assign w12735 = ~w11117 & ~w9393;
assign w12736 = w10653 & w13554;
assign w12737 = w11405 & w10011;
assign w12738 = w13839 & ~w719;
assign w12739 = (w14514 & w5164) | (w14514 & w7998) | (w5164 & w7998);
assign w12740 = (~w8899 & w5070) | (~w8899 & w996) | (w5070 & w996);
assign w12741 = (~w11959 & w7255) | (~w11959 & w253) | (w7255 & w253);
assign w12742 = ~w11064 & ~w5104;
assign w12743 = (w11037 & w9724) | (w11037 & w10033) | (w9724 & w10033);
assign w12744 = w7335 & w3904;
assign w12745 = ~w781 & ~w13088;
assign w12746 = ~w8171 & w3958;
assign w12747 = w433 & w10708;
assign w12748 = ~w6301 & ~w5247;
assign w12749 = ~w2463 & w9752;
assign w12750 = (~w7962 & w9012) | (~w7962 & w14333) | (w9012 & w14333);
assign w12751 = (w4772 & w12747) | (w4772 & w1117) | (w12747 & w1117);
assign w12752 = ~w4010 & ~w5269;
assign w12753 = (w6802 & w3907) | (w6802 & w3356) | (w3907 & w3356);
assign w12754 = w1956 & ~w4903;
assign w12755 = ~w10470 & ~w8320;
assign w12756 = w607 & ~w11934;
assign w12757 = w1098 & w12623;
assign w12758 = ~w10435 & w14457;
assign w12759 = w9403 & w4349;
assign w12760 = ~w6080 & w9679;
assign w12761 = (w12799 & w4131) | (w12799 & w11966) | (w4131 & w11966);
assign w12762 = ~w10997 & ~w4667;
assign w12763 = (~w7488 & w8826) | (~w7488 & w3398) | (w8826 & w3398);
assign w12764 = (w347 & w11882) | (w347 & w8062) | (w11882 & w8062);
assign w12765 = (~w10433 & w11990) | (~w10433 & w2057) | (w11990 & w2057);
assign w12766 = ~w9245 & w11097;
assign w12767 = ~w4158 & w9164;
assign w12768 = (w13444 & w7492) | (w13444 & w4461) | (w7492 & w4461);
assign w12769 = (w13885 & w11886) | (w13885 & w10988) | (w11886 & w10988);
assign w12770 = (~w9364 & w9441) | (~w9364 & w10801) | (w9441 & w10801);
assign w12771 = ~w12545 & w1455;
assign w12772 = w14263 & ~w13196;
assign w12773 = ~w11817 & w1527;
assign w12774 = (w8013 & w6492) | (w8013 & w3570) | (w6492 & w3570);
assign w12775 = ~w1906 & ~w1305;
assign w12776 = (w11734 & w2280) | (w11734 & w553) | (w2280 & w553);
assign w12777 = (w2144 & w5384) | (w2144 & w13846) | (w5384 & w13846);
assign w12778 = w931 & ~w3132;
assign w12779 = w5227 & w10036;
assign w12780 = w10422 & ~w10005;
assign w12781 = ~w3334 & ~w9817;
assign w12782 = w12483 & ~w13596;
assign w12783 = w12545 & ~w3730;
assign w12784 = (w7571 & w4061) | (w7571 & ~w13292) | (w4061 & ~w13292);
assign w12785 = ~w7483 & w411;
assign w12786 = (~w7240 & w3974) | (~w7240 & w10033) | (w3974 & w10033);
assign w12787 = ~w11745 & ~w11861;
assign w12788 = ~w9372 & ~w12048;
assign w12789 = ~w2333 & w7416;
assign w12790 = w9511 & w2092;
assign w12791 = w364 & ~w11361;
assign w12792 = (~w3215 & w13222) | (~w3215 & w12575) | (w13222 & w12575);
assign w12793 = w967 & ~w13270;
assign w12794 = (w14527 & w3421) | (w14527 & ~w8282) | (w3421 & ~w8282);
assign w12795 = w11321 & w2172;
assign w12796 = w45 & ~w13628;
assign w12797 = (w884 & ~w1140) | (w884 & w12552) | (~w1140 & w12552);
assign w12798 = w8253 & w11117;
assign w12799 = (~w9096 & w10033) | (~w9096 & ~w13379) | (w10033 & ~w13379);
assign w12800 = w4211 & w9180;
assign w12801 = w10681 & ~w10435;
assign w12802 = w4473 & ~w3044;
assign w12803 = w10286 & ~w11198;
assign w12804 = (w11969 & w7827) | (w11969 & w6369) | (w7827 & w6369);
assign w12805 = (~w1559 & w12298) | (~w1559 & w9948) | (w12298 & w9948);
assign w12806 = (~w1442 & w12003) | (~w1442 & w11363) | (w12003 & w11363);
assign w12807 = (w7082 & w4116) | (w7082 & w13719) | (w4116 & w13719);
assign w12808 = w12 & ~w1760;
assign w12809 = b121 & a121;
assign w12810 = (w9341 & w9108) | (w9341 & w773) | (w9108 & w773);
assign w12811 = w8540 & w6230;
assign w12812 = ~w7393 & ~w4496;
assign w12813 = w4482 & w5979;
assign w12814 = (~w11803 & w1275) | (~w11803 & w6852) | (w1275 & w6852);
assign w12815 = (~w5105 & w9608) | (~w5105 & w2869) | (w9608 & w2869);
assign w12816 = (~w11429 & w9414) | (~w11429 & w5561) | (w9414 & w5561);
assign w12817 = (w4524 & w14409) | (w4524 & ~w5483) | (w14409 & ~w5483);
assign w12818 = w1840 & w13565;
assign w12819 = ~w12958 & ~w2922;
assign w12820 = ~w7633 & ~w9121;
assign w12821 = ~w8929 & ~w5936;
assign w12822 = (~w13685 & w5897) | (~w13685 & w1759) | (w5897 & w1759);
assign w12823 = ~w12575 & ~w3215;
assign w12824 = ~w2762 & ~w10847;
assign w12825 = ~w5785 & w11211;
assign w12826 = (~w3098 & ~w4401) | (~w3098 & w941) | (~w4401 & w941);
assign w12827 = ~w922 & w2410;
assign w12828 = (w2029 & w6148) | (w2029 & w579) | (w6148 & w579);
assign w12829 = w14470 & ~w11462;
assign w12830 = w7067 & w13272;
assign w12831 = (w13713 & ~w10143) | (w13713 & ~w7464) | (~w10143 & ~w7464);
assign w12832 = (w7082 & w4708) | (w7082 & w13494) | (w4708 & w13494);
assign w12833 = (w13008 & ~w9506) | (w13008 & ~w1712) | (~w9506 & ~w1712);
assign w12834 = w10563 & w7417;
assign w12835 = w4213 & w9932;
assign w12836 = (w1849 & w5527) | (w1849 & w5770) | (w5527 & w5770);
assign w12837 = (w7762 & w9866) | (w7762 & ~w709) | (w9866 & ~w709);
assign w12838 = w183 & w6576;
assign w12839 = w11345 & w11117;
assign w12840 = w922 & w9015;
assign w12841 = ~w9381 & ~w8187;
assign w12842 = w2320 & ~w8389;
assign w12843 = ~w5533 & w1893;
assign w12844 = ~w6427 & ~w91;
assign w12845 = (w12776 & w2021) | (w12776 & w9941) | (w2021 & w9941);
assign w12846 = w11358 & w4550;
assign w12847 = ~w5005 & ~w5247;
assign w12848 = w4385 & w4103;
assign w12849 = ~w7782 & w14037;
assign w12850 = (w11385 & w12410) | (w11385 & w14365) | (w12410 & w14365);
assign w12851 = ~w569 & w7682;
assign w12852 = w8825 & ~w4963;
assign w12853 = ~w4473 & ~w12890;
assign w12854 = ~w2320 & w1949;
assign w12855 = w1692 & ~w1046;
assign w12856 = ~w5556 & ~w1235;
assign w12857 = (w13713 & w12831) | (w13713 & ~w10384) | (w12831 & ~w10384);
assign w12858 = w11395 & w10483;
assign w12859 = ~w10614 & w4045;
assign w12860 = ~w1493 & ~w5353;
assign w12861 = (w4202 & w2883) | (w4202 & w9324) | (w2883 & w9324);
assign w12862 = w3197 & w10903;
assign w12863 = w10509 & w12740;
assign w12864 = (w1919 & w5927) | (w1919 & w10165) | (w5927 & w10165);
assign w12865 = w9541 & ~w13054;
assign w12866 = (w11416 & w9497) | (w11416 & w3282) | (w9497 & w3282);
assign w12867 = ~w607 & w6689;
assign w12868 = ~w1096 & ~w6886;
assign w12869 = w1845 & ~w1838;
assign w12870 = (w1096 & w12499) | (w1096 & w10270) | (w12499 & w10270);
assign w12871 = ~w8791 & w12620;
assign w12872 = ~w12003 & w4826;
assign w12873 = w509 & ~w11117;
assign w12874 = ~w3986 & ~w3242;
assign w12875 = ~w14094 & w5077;
assign w12876 = ~w1785 & w7858;
assign w12877 = w2372 & w7725;
assign w12878 = ~w12575 & w1619;
assign w12879 = w9921 & w1949;
assign w12880 = (w1938 & w8652) | (w1938 & w14182) | (w8652 & w14182);
assign w12881 = ~w14375 & w5062;
assign w12882 = ~w10576 & w1179;
assign w12883 = ~w2762 & w36;
assign w12884 = (~w12463 & w9263) | (~w12463 & w9867) | (w9263 & w9867);
assign w12885 = (w11138 & w4305) | (w11138 & w5473) | (w4305 & w5473);
assign w12886 = (~w9305 & w5587) | (~w9305 & w13812) | (w5587 & w13812);
assign w12887 = w2656 & ~w1171;
assign w12888 = (~w14131 & w13174) | (~w14131 & w5541) | (w13174 & w5541);
assign w12889 = ~w7726 & w10224;
assign w12890 = ~w13917 & w11226;
assign w12891 = w9433 & w10590;
assign w12892 = (w11020 & w10382) | (w11020 & w11696) | (w10382 & w11696);
assign w12893 = ~b71 & ~a71;
assign w12894 = (w12185 & w6002) | (w12185 & w12376) | (w6002 & w12376);
assign w12895 = ~w9583 & w2477;
assign w12896 = (w3556 & w11136) | (w3556 & w4677) | (w11136 & w4677);
assign w12897 = w6384 & w12589;
assign w12898 = w1555 & w4780;
assign w12899 = w9183 & w7455;
assign w12900 = ~w10182 & w3017;
assign w12901 = (~w5785 & w12107) | (~w5785 & w10995) | (w12107 & w10995);
assign w12902 = (w931 & w9099) | (w931 & w12778) | (w9099 & w12778);
assign w12903 = ~w10334 & ~w4680;
assign w12904 = w10676 & w4288;
assign w12905 = ~w8035 & w9767;
assign w12906 = w5177 & w13682;
assign w12907 = ~w4921 & w9477;
assign w12908 = b36 & a36;
assign w12909 = w7395 & ~w3548;
assign w12910 = w13009 & w421;
assign w12911 = (w13771 & w12186) | (w13771 & w7063) | (w12186 & w7063);
assign w12912 = w4796 & ~w8004;
assign w12913 = ~w12398 & w10855;
assign w12914 = w7256 & ~w7441;
assign w12915 = (~w8827 & w11108) | (~w8827 & w4170) | (w11108 & w4170);
assign w12916 = (w11201 & w667) | (w11201 & ~w10052) | (w667 & ~w10052);
assign w12917 = ~w5490 & w11542;
assign w12918 = ~w6244 & w11048;
assign w12919 = ~w12321 & w3044;
assign w12920 = w3550 & ~w3790;
assign w12921 = ~w4721 & ~w7421;
assign w12922 = ~w12429 & ~w13521;
assign w12923 = ~w6986 & w8900;
assign w12924 = (~w13008 & w10435) | (~w13008 & w9848) | (w10435 & w9848);
assign w12925 = w4787 & ~w13531;
assign w12926 = ~w4127 & w9923;
assign w12927 = (w11059 & w10127) | (w11059 & w12067) | (w10127 & w12067);
assign w12928 = (w246 & w6071) | (w246 & w11939) | (w6071 & w11939);
assign w12929 = ~w8183 & w2729;
assign w12930 = ~w12378 & w518;
assign w12931 = w5177 & w3311;
assign w12932 = ~w9037 & ~w12246;
assign w12933 = (~w6689 & w3017) | (~w6689 & w28) | (w3017 & w28);
assign w12934 = (~w5664 & w14335) | (~w5664 & w6010) | (w14335 & w6010);
assign w12935 = w309 & ~w12311;
assign w12936 = ~w3890 & ~w5296;
assign w12937 = (~w353 & w10318) | (~w353 & ~w8282) | (w10318 & ~w8282);
assign w12938 = w5032 & w11789;
assign w12939 = (~w2389 & w6058) | (~w2389 & w6223) | (w6058 & w6223);
assign w12940 = w2980 & w3512;
assign w12941 = (~w11560 & w4191) | (~w11560 & w1630) | (w4191 & w1630);
assign w12942 = w914 & w2572;
assign w12943 = b81 & a81;
assign w12944 = (~w4921 & w13663) | (~w4921 & w9549) | (w13663 & w9549);
assign w12945 = w4787 & w11498;
assign w12946 = (w5483 & w2122) | (w5483 & w6333) | (w2122 & w6333);
assign w12947 = w1594 & w5961;
assign w12948 = w11013 & ~w4458;
assign w12949 = ~w884 & ~w12;
assign w12950 = w12672 & w1736;
assign w12951 = ~w2674 & w12603;
assign w12952 = (w12125 & w11859) | (w12125 & w11151) | (w11859 & w11151);
assign w12953 = ~w1789 & w9916;
assign w12954 = (w3650 & ~w7084) | (w3650 & w11630) | (~w7084 & w11630);
assign w12955 = ~w13587 & w3437;
assign w12956 = (w13005 & w4559) | (w13005 & ~w1563) | (w4559 & ~w1563);
assign w12957 = (~w8279 & w6918) | (~w8279 & ~w5552) | (w6918 & ~w5552);
assign w12958 = b90 & a90;
assign w12959 = (w1062 & ~w4378) | (w1062 & w3528) | (~w4378 & w3528);
assign w12960 = ~w5280 & w4271;
assign w12961 = w8920 & w1351;
assign w12962 = w4587 & w8900;
assign w12963 = w12368 & w1420;
assign w12964 = w12271 & w3087;
assign w12965 = w7342 & w9454;
assign w12966 = (w11978 & w4544) | (w11978 & ~w8163) | (w4544 & ~w8163);
assign w12967 = w8507 & w13047;
assign w12968 = (~w2144 & w709) | (~w2144 & w225) | (w709 & w225);
assign w12969 = (w7725 & w4555) | (w7725 & w6931) | (w4555 & w6931);
assign w12970 = (~w3158 & w5852) | (~w3158 & w7671) | (w5852 & w7671);
assign w12971 = ~w1873 & ~w143;
assign w12972 = w4441 & w6230;
assign w12973 = (w1416 & w1153) | (w1416 & w9325) | (w1153 & w9325);
assign w12974 = ~w14141 & w1399;
assign w12975 = (w2595 & w5476) | (w2595 & ~w4754) | (w5476 & ~w4754);
assign w12976 = ~w3141 & ~w701;
assign w12977 = w8502 & ~w14300;
assign w12978 = ~w1753 & w14073;
assign w12979 = ~w4359 & ~w7455;
assign w12980 = w12636 & ~w8690;
assign w12981 = (w12656 & w2638) | (w12656 & w3437) | (w2638 & w3437);
assign w12982 = ~w8560 & w13568;
assign w12983 = ~w8110 & w8713;
assign w12984 = w3146 & ~w5243;
assign w12985 = ~w10393 & ~w11613;
assign w12986 = ~w1274 & w2753;
assign w12987 = (~w13862 & w294) | (~w13862 & w6067) | (w294 & w6067);
assign w12988 = ~w2387 & ~w3036;
assign w12989 = w2147 & ~w8489;
assign w12990 = w10265 & w11866;
assign w12991 = ~w1785 & w6629;
assign w12992 = w11817 & w11613;
assign w12993 = w12060 & w5464;
assign w12994 = ~w12194 & ~w9693;
assign w12995 = (w3122 & w13553) | (w3122 & w2746) | (w13553 & w2746);
assign w12996 = ~w8791 & w1507;
assign w12997 = ~w8226 & w8452;
assign w12998 = ~w12656 & ~w3615;
assign w12999 = (~w10711 & ~w4582) | (~w10711 & ~w6802) | (~w4582 & ~w6802);
assign w13000 = w4369 & w10162;
assign w13001 = ~w2023 & w6711;
assign w13002 = w4836 & w3906;
assign w13003 = ~w8223 & ~w924;
assign w13004 = w7794 & ~w10811;
assign w13005 = w2137 & w4777;
assign w13006 = w3018 & ~w12055;
assign w13007 = (~w5161 & w1761) | (~w5161 & w9343) | (w1761 & w9343);
assign w13008 = ~w622 & ~w10916;
assign w13009 = ~w3278 & w7576;
assign w13010 = (~w2144 & w9859) | (~w2144 & w8341) | (w9859 & w8341);
assign w13011 = ~w10309 & ~w1516;
assign w13012 = w8119 & w10950;
assign w13013 = (w9940 & w1172) | (w9940 & w88) | (w1172 & w88);
assign w13014 = ~w183 & ~w3632;
assign w13015 = (w12369 & w6092) | (w12369 & w6272) | (w6092 & w6272);
assign w13016 = (~w14340 & w596) | (~w14340 & ~w14335) | (w596 & ~w14335);
assign w13017 = (~w2463 & w1217) | (~w2463 & w5360) | (w1217 & w5360);
assign w13018 = ~w7965 & w2586;
assign w13019 = ~w13714 & w12737;
assign w13020 = (w2038 & w13329) | (w2038 & w3776) | (w13329 & w3776);
assign w13021 = (w7914 & w13199) | (w7914 & w5620) | (w13199 & w5620);
assign w13022 = (~w1096 & w2144) | (~w1096 & w3226) | (w2144 & w3226);
assign w13023 = (w12406 & w2902) | (w12406 & w1428) | (w2902 & w1428);
assign w13024 = (w10637 & w2231) | (w10637 & w8270) | (w2231 & w8270);
assign w13025 = w13526 & w12311;
assign w13026 = w7367 & w5788;
assign w13027 = ~w9012 & w6151;
assign w13028 = w8743 & ~w7033;
assign w13029 = ~w7794 & ~w2320;
assign w13030 = (w9738 & w2798) | (w9738 & w4391) | (w2798 & w4391);
assign w13031 = w11628 & w9779;
assign w13032 = w10676 & w608;
assign w13033 = (w12620 & w12499) | (w12620 & w7753) | (w12499 & w7753);
assign w13034 = ~w9861 & ~w9788;
assign w13035 = w7032 & w5184;
assign w13036 = ~w12113 & ~w784;
assign w13037 = w7641 & w6945;
assign w13038 = ~w11960 & w3496;
assign w13039 = w12491 & ~w6162;
assign w13040 = (w8047 & w8937) | (w8047 & w14082) | (w8937 & w14082);
assign w13041 = (w499 & w6932) | (w499 & ~w1840) | (w6932 & ~w1840);
assign w13042 = ~w6690 & ~w2698;
assign w13043 = w11934 & w9503;
assign w13044 = w2038 & w11732;
assign w13045 = ~w12735 & w8413;
assign w13046 = (w10290 & ~w183) | (w10290 & w11686) | (~w183 & w11686);
assign w13047 = ~w7314 & w5504;
assign w13048 = w5177 & w8512;
assign w13049 = (w12721 & ~w8609) | (w12721 & w13076) | (~w8609 & w13076);
assign w13050 = w11807 & ~w8844;
assign w13051 = (w7243 & w1495) | (w7243 & w5622) | (w1495 & w5622);
assign w13052 = (w12656 & w2638) | (w12656 & ~w11714) | (w2638 & ~w11714);
assign w13053 = w1838 & ~w11117;
assign w13054 = (~w13077 & ~w9839) | (~w13077 & w4556) | (~w9839 & w4556);
assign w13055 = ~w13282 & ~w5626;
assign w13056 = ~w6176 & ~w11345;
assign w13057 = ~w8420 & w3983;
assign w13058 = (~w12819 & w8937) | (~w12819 & w13646) | (w8937 & w13646);
assign w13059 = w11332 & w9265;
assign w13060 = w3069 & w9032;
assign w13061 = w5002 & ~w563;
assign w13062 = w12672 & w14219;
assign w13063 = (~w8032 & w11436) | (~w8032 & w8850) | (w11436 & w8850);
assign w13064 = ~w6170 & w137;
assign w13065 = ~w3997 & ~w6267;
assign w13066 = (w4041 & w9990) | (w4041 & ~w7) | (w9990 & ~w7);
assign w13067 = (w6822 & w9018) | (w6822 & w3) | (w9018 & w3);
assign w13068 = (w6219 & w4520) | (w6219 & w9726) | (w4520 & w9726);
assign w13069 = ~w183 & ~w6646;
assign w13070 = (w8396 & w4811) | (w8396 & w8875) | (w4811 & w8875);
assign w13071 = (~w10247 & w2463) | (~w10247 & w3867) | (w2463 & w3867);
assign w13072 = (w3427 & w1935) | (w3427 & w9750) | (w1935 & w9750);
assign w13073 = ~w4441 & ~w1987;
assign w13074 = w6845 & ~w6192;
assign w13075 = w560 & ~w1949;
assign w13076 = w6335 & w12721;
assign w13077 = w14072 & w13694;
assign w13078 = w4658 & w9064;
assign w13079 = ~w2311 & ~w3566;
assign w13080 = w9256 & w2701;
assign w13081 = w142 & ~w12371;
assign w13082 = ~w1715 & w9500;
assign w13083 = ~w646 & w10504;
assign w13084 = ~w9504 & w3183;
assign w13085 = (w7906 & w4158) | (w7906 & w9828) | (w4158 & w9828);
assign w13086 = (w10123 & w11802) | (w10123 & w5034) | (w11802 & w5034);
assign w13087 = w3017 & w7267;
assign w13088 = ~w4651 & w12885;
assign w13089 = ~w13095 & w14129;
assign w13090 = (~w5702 & w2005) | (~w5702 & w12956) | (w2005 & w12956);
assign w13091 = w11708 & w8359;
assign w13092 = ~w4591 & ~w4642;
assign w13093 = w7376 & ~w1396;
assign w13094 = w347 & ~w11397;
assign w13095 = ~w5556 & w11604;
assign w13096 = ~w6064 & w2729;
assign w13097 = (~w9141 & w2732) | (~w9141 & w12459) | (w2732 & w12459);
assign w13098 = w10510 & ~w10425;
assign w13099 = w1450 & w3238;
assign w13100 = w4447 & w13323;
assign w13101 = ~w12604 & ~w2701;
assign w13102 = (w12138 & ~w4287) | (w12138 & w8240) | (~w4287 & w8240);
assign w13103 = ~w3027 & ~w8401;
assign w13104 = ~w12380 & ~w11027;
assign w13105 = ~w14530 & w12530;
assign w13106 = ~w10249 & ~w2615;
assign w13107 = ~w4050 & w4637;
assign w13108 = w6926 & ~w10820;
assign w13109 = ~w3289 | ~w7644;
assign w13110 = ~w11264 & ~w6218;
assign w13111 = (~w2218 & w6887) | (~w2218 & w10493) | (w6887 & w10493);
assign w13112 = (~w10213 & w9963) | (~w10213 & w13331) | (w9963 & w13331);
assign w13113 = ~w7356 & w13245;
assign w13114 = w12170 & ~w803;
assign w13115 = ~w8234 & ~w8442;
assign w13116 = ~w1216 & w8661;
assign w13117 = w9226 & w7962;
assign w13118 = (~w4134 & w301) | (~w4134 & w104) | (w301 & w104);
assign w13119 = w8122 & ~w4448;
assign w13120 = (w2670 & w14503) | (w2670 & w7363) | (w14503 & w7363);
assign w13121 = w5485 & ~w2795;
assign w13122 = w10326 & ~w4011;
assign w13123 = w14030 & w4247;
assign w13124 = w4302 & ~w1442;
assign w13125 = (w13665 & w11147) | (w13665 & w8416) | (w11147 & w8416);
assign w13126 = ~w235 & ~w10256;
assign w13127 = (w6953 & w7554) | (w6953 & w14148) | (w7554 & w14148);
assign w13128 = w5177 & ~w1805;
assign w13129 = ~w142 & w884;
assign w13130 = ~w2872 & w13276;
assign w13131 = w12457 & w8901;
assign w13132 = w1764 & ~w14512;
assign w13133 = ~w4607 & w12871;
assign w13134 = ~w8710 & w10751;
assign w13135 = (w7295 & w4399) | (w7295 & w1503) | (w4399 & w1503);
assign w13136 = (w4724 & ~w12219) | (w4724 & w3715) | (~w12219 & w3715);
assign w13137 = (~w4158 & w9350) | (~w4158 & w14090) | (w9350 & w14090);
assign w13138 = ~w1563 & w5279;
assign w13139 = (w9457 & w3258) | (w9457 & ~w13236) | (w3258 & ~w13236);
assign w13140 = w10286 & ~w13306;
assign w13141 = ~w9616 & ~w7650;
assign w13142 = w7034 & ~w4248;
assign w13143 = w6679 & w9699;
assign w13144 = w12553 & w11395;
assign w13145 = w11287 & w2729;
assign w13146 = ~w2730 & ~w4884;
assign w13147 = w3550 & w4298;
assign w13148 = ~w13122 & ~w2656;
assign w13149 = w7472 | ~w6716;
assign w13150 = (w14617 & w6990) | (w14617 & w3246) | (w6990 & w3246);
assign w13151 = w13976 & ~w3362;
assign w13152 = w12636 & ~w6454;
assign w13153 = ~w13324 & w3060;
assign w13154 = (~w1997 & w4307) | (~w1997 & ~w14492) | (w4307 & ~w14492);
assign w13155 = ~w14664 & w5426;
assign w13156 = w1049 & w12387;
assign w13157 = ~w4341 & ~w6016;
assign w13158 = w347 & ~w7844;
assign w13159 = w12360 & w6396;
assign w13160 = (~w7244 & ~w5282) | (~w7244 & w10494) | (~w5282 & w10494);
assign w13161 = (w3550 & w8331) | (w3550 & w2714) | (w8331 & w2714);
assign w13162 = ~w5620 & ~w13760;
assign w13163 = (w11964 & w7008) | (w11964 & w5908) | (w7008 & w5908);
assign w13164 = ~w9132 & ~w7166;
assign w13165 = w12207 & w6430;
assign w13166 = w360 & ~w5247;
assign w13167 = (~w142 & ~w13323) | (~w142 & w6872) | (~w13323 & w6872);
assign w13168 = (w10630 & w7666) | (w10630 & w10466) | (w7666 & w10466);
assign w13169 = w9265 & w10087;
assign w13170 = w7772 & ~w1712;
assign w13171 = (w11936 & w13706) | (w11936 & w9567) | (w13706 & w9567);
assign w13172 = ~w4401 & w5744;
assign w13173 = w3872 & ~w898;
assign w13174 = w13612 & w7361;
assign w13175 = (~w13531 & ~w953) | (~w13531 & w4428) | (~w953 & w4428);
assign w13176 = ~w3792 & ~w3325;
assign w13177 = ~w10245 & w1056;
assign w13178 = w11006 & w711;
assign w13179 = (~w14395 & w13587) | (~w14395 & w8354) | (w13587 & w8354);
assign w13180 = w7888 & ~w4317;
assign w13181 = w3219 & ~w7630;
assign w13182 = (w9319 & w12051) | (w9319 & w10067) | (w12051 & w10067);
assign w13183 = ~w9374 & ~w7133;
assign w13184 = (~w2168 & w2579) | (~w2168 & w12602) | (w2579 & w12602);
assign w13185 = ~w8480 & ~w9101;
assign w13186 = w6572 & w5664;
assign w13187 = (w804 & w426) | (w804 & w2450) | (w426 & w2450);
assign w13188 = w7305 & ~w11934;
assign w13189 = ~b114 & ~a114;
assign w13190 = ~w6253 & ~w6837;
assign w13191 = ~w6444 & ~w6666;
assign w13192 = ~w1802 & w2729;
assign w13193 = (w13379 & w8524) | (w13379 & w7699) | (w8524 & w7699);
assign w13194 = w5071 & w3328;
assign w13195 = (w5483 & w10867) | (w5483 & w8138) | (w10867 & w8138);
assign w13196 = (~w1692 & w2604) | (~w1692 & w7494) | (w2604 & w7494);
assign w13197 = w10645 & w12479;
assign w13198 = ~w6557 & ~w8249;
assign w13199 = w13620 & w7914;
assign w13200 = w11462 & w3904;
assign w13201 = ~w2412 & w1309;
assign w13202 = ~w5218 & ~w11424;
assign w13203 = (w3550 & w3935) | (w3550 & w9210) | (w3935 & w9210);
assign w13204 = (~w9817 & w11429) | (~w9817 & w9513) | (w11429 & w9513);
assign w13205 = (w4354 & w12878) | (w4354 & ~w10917) | (w12878 & ~w10917);
assign w13206 = ~w13697 & w4445;
assign w13207 = w10483 & ~w10179;
assign w13208 = ~w361 & ~w10411;
assign w13209 = (w12460 & w3044) | (w12460 & w11578) | (w3044 & w11578);
assign w13210 = w5282 & w7670;
assign w13211 = ~w10826 & w12367;
assign w13212 = ~w11057 & ~w6149;
assign w13213 = (w10578 & w12973) | (w10578 & w8228) | (w12973 & w8228);
assign w13214 = ~w14526 & ~w3019;
assign w13215 = w9861 & ~w1062;
assign w13216 = (w12920 & w9979) | (w12920 & w11651) | (w9979 & w11651);
assign w13217 = w5612 & w4398;
assign w13218 = (~w12376 & w13808) | (~w12376 & w9154) | (w13808 & w9154);
assign w13219 = w14396 & ~w4751;
assign w13220 = w1202 & ~w8938;
assign w13221 = w13743 & ~w3685;
assign w13222 = ~w8732 & ~w9399;
assign w13223 = ~w1605 & w14391;
assign w13224 = w6270 & w13290;
assign w13225 = ~w3151 & w3494;
assign w13226 = w10949 & ~w13800;
assign w13227 = ~w5108 & ~w1516;
assign w13228 = ~w7754 & ~w6975;
assign w13229 = (w4787 & ~w10483) | (w4787 & w5873) | (~w10483 & w5873);
assign w13230 = w12241 & ~w12460;
assign w13231 = w5294 & ~w1172;
assign w13232 = w8894 & ~w3209;
assign w13233 = w3751 & ~w12642;
assign w13234 = w12943 & ~w1712;
assign w13235 = (~w1519 & w2821) | (~w1519 & w11430) | (w2821 & w11430);
assign w13236 = ~w8226 & w1966;
assign w13237 = ~w4158 & w3148;
assign w13238 = ~w12003 & w9111;
assign w13239 = (w1771 & w2786) | (w1771 & w13225) | (w2786 & w13225);
assign w13240 = b1 & a1;
assign w13241 = w4408 & ~w5565;
assign w13242 = w7312 & w9896;
assign w13243 = (~w2463 & w5955) | (~w2463 & w12258) | (w5955 & w12258);
assign w13244 = w7165 & w13867;
assign w13245 = ~w42 & ~w1189;
assign w13246 = (~w5556 & w13587) | (~w5556 & w10164) | (w13587 & w10164);
assign w13247 = w12112 & ~w4520;
assign w13248 = ~w8791 & w9142;
assign w13249 = w11462 & ~w235;
assign w13250 = ~w450 & w11633;
assign w13251 = ~w10334 & ~w8662;
assign w13252 = ~w12517 & ~w10535;
assign w13253 = (w5768 & w13772) | (w5768 & w7062) | (w13772 & w7062);
assign w13254 = ~w5369 & ~w13216;
assign w13255 = ~w491 & ~w807;
assign w13256 = b20 & a20;
assign w13257 = ~w10517 & ~w5761;
assign w13258 = w5707 & ~w1798;
assign w13259 = (w5918 & w8312) | (w5918 & w4534) | (w8312 & w4534);
assign w13260 = w3463 & ~w1311;
assign w13261 = (w10773 & w613) | (w10773 & w10563) | (w613 & w10563);
assign w13262 = (w1949 & w1843) | (w1949 & w4402) | (w1843 & w4402);
assign w13263 = ~w1840 & ~w254;
assign w13264 = ~w732 & w7613;
assign w13265 = (w11068 & ~w341) | (w11068 & w9314) | (~w341 & w9314);
assign w13266 = w4132 & w8172;
assign w13267 = w6889 & ~w8992;
assign w13268 = (~w3700 & w10487) | (~w3700 & w12898) | (w10487 & w12898);
assign w13269 = ~w9794 & ~w1503;
assign w13270 = w10152 & ~w7833;
assign w13271 = w4982 & ~w11213;
assign w13272 = (~w2655 & w2269) | (~w2655 & w469) | (w2269 & w469);
assign w13273 = (~w13282 & w9375) | (~w13282 & w1461) | (w9375 & w1461);
assign w13274 = w1550 & ~w7995;
assign w13275 = (~w11429 & w14198) | (~w11429 & w3003) | (w14198 & w3003);
assign w13276 = w5099 & w5647;
assign w13277 = (w6423 & w7203) | (w6423 & w1595) | (w7203 & w1595);
assign w13278 = (w9012 & w3977) | (w9012 & w8309) | (w3977 & w8309);
assign w13279 = ~w13462 & w4687;
assign w13280 = w7822 & ~w10533;
assign w13281 = w9672 & ~w2663;
assign w13282 = ~w11402 & ~w8592;
assign w13283 = ~w6021 & w12037;
assign w13284 = (w2175 & w9289) | (w2175 & w7707) | (w9289 & w7707);
assign w13285 = ~w12808 | w1760;
assign w13286 = ~w5852 & w4190;
assign w13287 = w330 & w5168;
assign w13288 = (w2343 & w12610) | (w2343 & w9034) | (w12610 & w9034);
assign w13289 = (~w922 & w3775) | (~w922 & w1986) | (w3775 & w1986);
assign w13290 = ~w631 & ~w2929;
assign w13291 = (w2777 & w2959) | (w2777 & ~w10033) | (w2959 & ~w10033);
assign w13292 = (~w13379 & w9514) | (~w13379 & w12743) | (w9514 & w12743);
assign w13293 = ~w5619 & w11869;
assign w13294 = w2661 & w3121;
assign w13295 = (w7082 & w4968) | (w7082 & w5028) | (w4968 & w5028);
assign w13296 = ~w8774 & ~w4693;
assign w13297 = ~b124 & ~a124;
assign w13298 = ~w6662 & ~w12218;
assign w13299 = ~w12697 & ~w11122;
assign w13300 = ~w8171 & ~w6888;
assign w13301 = (~w5783 & w12541) | (~w5783 & w5142) | (w12541 & w5142);
assign w13302 = ~w4501 & w9635;
assign w13303 = ~w14088 & ~w5067;
assign w13304 = ~w1128 & ~w9167;
assign w13305 = w1006 & ~w9317;
assign w13306 = b51 & a51;
assign w13307 = w10309 & ~w14054;
assign w13308 = ~w922 & w9871;
assign w13309 = w6087 & w6796;
assign w13310 = ~w11586 & w1871;
assign w13311 = (~w10272 & ~w7464) | (~w10272 & w14197) | (~w7464 & w14197);
assign w13312 = ~w10966 & ~w10325;
assign w13313 = w5026 & ~w5974;
assign w13314 = w9264 & w13820;
assign w13315 = (w1593 & w11060) | (w1593 & w217) | (w11060 & w217);
assign w13316 = w7463 & w9508;
assign w13317 = ~w11261 & w1109;
assign w13318 = w13197 & ~w5197;
assign w13319 = (~w2144 & w5690) | (~w2144 & w7476) | (w5690 & w7476);
assign w13320 = ~w13096 & ~w7785;
assign w13321 = w7376 & w13081;
assign w13322 = (w10664 & ~w4843) | (w10664 & w10116) | (~w4843 & w10116);
assign w13323 = ~w11757 & ~w9256;
assign w13324 = w5675 & ~w9157;
assign w13325 = ~w9258 & w14590;
assign w13326 = ~w2144 & w13801;
assign w13327 = w3576 & w12483;
assign w13328 = ~w11905 & ~w6219;
assign w13329 = ~w8655 & w2038;
assign w13330 = ~w10970 & w1879;
assign w13331 = w9708 & ~w1928;
assign w13332 = ~w7711 & ~w10269;
assign w13333 = w9244 & w6381;
assign w13334 = ~w2599 & ~w3823;
assign w13335 = ~w3786 & ~w2675;
assign w13336 = ~w5559 & w221;
assign w13337 = (w12909 & ~w13533) | (w12909 & w7602) | (~w13533 & w7602);
assign w13338 = w12667 & ~w7242;
assign w13339 = w8519 & w8010;
assign w13340 = (w8007 & w2124) | (w8007 & w9403) | (w2124 & w9403);
assign w13341 = w9921 & w12656;
assign w13342 = w6975 & w11117;
assign w13343 = (w4026 & w3330) | (w4026 & w3072) | (w3330 & w3072);
assign w13344 = ~b111 & ~a111;
assign w13345 = w2096 & w5761;
assign w13346 = w4315 & ~w2730;
assign w13347 = (w1344 & w3336) | (w1344 & ~w13980) | (w3336 & ~w13980);
assign w13348 = w8191 | ~w5406;
assign w13349 = w5463 & ~w6654;
assign w13350 = (~w4711 & w1385) | (~w4711 & w6729) | (w1385 & w6729);
assign w13351 = w8534 & w6570;
assign w13352 = (w254 & w6866) | (w254 & w3378) | (w6866 & w3378);
assign w13353 = (w2317 & w1077) | (w2317 & w10890) | (w1077 & w10890);
assign w13354 = ~w7348 & ~w1692;
assign w13355 = (~w8769 & w1885) | (~w8769 & w3871) | (w1885 & w3871);
assign w13356 = (w3427 & ~w4199) | (w3427 & ~w13183) | (~w4199 & ~w13183);
assign w13357 = (w13865 & w3150) | (w13865 & w3652) | (w3150 & w3652);
assign w13358 = w10082 & w7670;
assign w13359 = (w11708 & ~w1692) | (w11708 & w8331) | (~w1692 & w8331);
assign w13360 = ~w5860 & w4017;
assign w13361 = w4213 & w14340;
assign w13362 = (w9680 & w4755) | (w9680 & ~w21) | (w4755 & ~w21);
assign w13363 = ~w8956 & ~w3902;
assign w13364 = w1722 | ~w235;
assign w13365 = (~w11385 & w7731) | (~w11385 & w8311) | (w7731 & w8311);
assign w13366 = w7129 & w1640;
assign w13367 = w7794 & ~w5576;
assign w13368 = (w12614 & w5234) | (w12614 & w11017) | (w5234 & w11017);
assign w13369 = (w7458 & ~w144) | (w7458 & w6020) | (~w144 & w6020);
assign w13370 = ~w8183 & w5761;
assign w13371 = ~w2311 & ~w13259;
assign w13372 = (~w7914 & w11658) | (~w7914 & w11925) | (w11658 & w11925);
assign w13373 = ~w1682 & w2701;
assign w13374 = (~w7335 & w9582) | (~w7335 & w4629) | (w9582 & w4629);
assign w13375 = w11475 & ~w13227;
assign w13376 = w12173 & ~w5682;
assign w13377 = (w9276 & w14059) | (w9276 & w5159) | (w14059 & w5159);
assign w13378 = ~w13324 & w4702;
assign w13379 = (w318 & ~w11516) | (w318 & w7240) | (~w11516 & w7240);
assign w13380 = (~w9608 & w7536) | (~w9608 & w9922) | (w7536 & w9922);
assign w13381 = ~w1096 & w5213;
assign w13382 = ~w4604 & w5679;
assign w13383 = (w2007 & w7462) | (w2007 & w6140) | (w7462 & w6140);
assign w13384 = ~w10986 & w10904;
assign w13385 = w14302 & ~w1199;
assign w13386 = w5522 & ~w7794;
assign w13387 = ~w7488 & w12327;
assign w13388 = (~w6889 & w1121) | (~w6889 & w7693) | (w1121 & w7693);
assign w13389 = (w6949 & ~w13892) | (w6949 & w2865) | (~w13892 & w2865);
assign w13390 = w12553 & w5860;
assign w13391 = (~w13633 & w11426) | (~w13633 & ~w9034) | (w11426 & ~w9034);
assign w13392 = ~w11817 & w3812;
assign w13393 = ~w6047 & w11484;
assign w13394 = ~w10252 & ~w3786;
assign w13395 = (w6500 & w1129) | (w6500 & w13574) | (w1129 & w13574);
assign w13396 = (w13324 & w3833) | (w13324 & w13661) | (w3833 & w13661);
assign w13397 = w8873 & w10917;
assign w13398 = ~w4685 & ~w5600;
assign w13399 = w10378 & ~w9149;
assign w13400 = (~w10704 & w9181) | (~w10704 & w5066) | (w9181 & w5066);
assign w13401 = (~w4565 & w6117) | (~w4565 & w14002) | (w6117 & w14002);
assign w13402 = w4425 & w6845;
assign w13403 = w8343 & ~w7103;
assign w13404 = ~w12088 & ~w6266;
assign w13405 = (w3510 & w4332) | (w3510 & w6851) | (w4332 & w6851);
assign w13406 = w8166 & w7506;
assign w13407 = w4941 & w6172;
assign w13408 = w8183 & w13323;
assign w13409 = ~w5379 & w4232;
assign w13410 = w13796 & w7231;
assign w13411 = ~w6371 & w9536;
assign w13412 = ~w1609 & w7276;
assign w13413 = ~w443 & w1108;
assign w13414 = (~w142 & ~w7670) | (~w142 & w6872) | (~w7670 & w6872);
assign w13415 = ~w4989 & w9561;
assign w13416 = ~w5860 & w6502;
assign w13417 = (~w1663 & w11513) | (~w1663 & w5820) | (w11513 & w5820);
assign w13418 = w7453 & ~w10857;
assign w13419 = ~w9748 & ~w6483;
assign w13420 = w12240 & w309;
assign w13421 = w2332 & w5490;
assign w13422 = ~w14664 & w10473;
assign w13423 = ~b44 & ~a44;
assign w13424 = (w9541 & w4072) | (w9541 & w6765) | (w4072 & w6765);
assign w13425 = ~w5559 & w5924;
assign w13426 = w12901 & w2149;
assign w13427 = ~w10863 & w7573;
assign w13428 = ~w11139 & w2708;
assign w13429 = w5522 & w11934;
assign w13430 = (w1498 & ~w10001) | (w1498 & w9231) | (~w10001 & w9231);
assign w13431 = (~w2144 & w6322) | (~w2144 & w10587) | (w6322 & w10587);
assign w13432 = (w6873 & w9217) | (w6873 & w378) | (w9217 & w378);
assign w13433 = (~w5449 & w6259) | (~w5449 & w2319) | (w6259 & w2319);
assign w13434 = (~w3325 & w9608) | (~w3325 & w14332) | (w9608 & w14332);
assign w13435 = (~w9012 & w11387) | (~w9012 & w8765) | (w11387 & w8765);
assign w13436 = ~w12374 & w14177;
assign w13437 = ~w10435 & w7414;
assign w13438 = w11899 & ~w4147;
assign w13439 = ~w3130 & w2701;
assign w13440 = (~w9608 & w4695) | (~w9608 & w9630) | (w4695 & w9630);
assign w13441 = w1559 & ~w12805;
assign w13442 = w218 & w6230;
assign w13443 = ~w16 & w6035;
assign w13444 = ~w868 & ~w1781;
assign w13445 = (~w473 & w1229) | (~w473 & w13759) | (w1229 & w13759);
assign w13446 = ~w7080 & ~w4627;
assign w13447 = (~w10272 & w2048) | (~w10272 & ~w5901) | (w2048 & ~w5901);
assign w13448 = ~w6122 & ~w7214;
assign w13449 = ~w3218 & ~w3334;
assign w13450 = (w14514 & w7355) | (w14514 & w3295) | (w7355 & w3295);
assign w13451 = b12 & a12;
assign w13452 = w5590 & w2707;
assign w13453 = ~w11577 & ~w224;
assign w13454 = (w6017 & w10267) | (w6017 & ~w4232) | (w10267 & ~w4232);
assign w13455 = (~w5952 & w14646) | (~w5952 & w19) | (w14646 & w19);
assign w13456 = w2812 & w13028;
assign w13457 = w3092 & w5822;
assign w13458 = (w8399 & w10852) | (w8399 & w8588) | (w10852 & w8588);
assign w13459 = (w7211 & w310) | (w7211 & w3008) | (w310 & w3008);
assign w13460 = (w5952 & w648) | (w5952 & w12234) | (w648 & w12234);
assign w13461 = w10872 & ~w3019;
assign w13462 = w167 & ~w2642;
assign w13463 = w719 & w3427;
assign w13464 = (~w5934 & w9388) | (~w5934 & w11404) | (w9388 & w11404);
assign w13465 = w12371 & ~w10699;
assign w13466 = w6606 & w13603;
assign w13467 = ~w1922 & w9776;
assign w13468 = ~w10854 & w11364;
assign w13469 = w8427 & w10166;
assign w13470 = w5860 & ~w309;
assign w13471 = ~w4512 & w5467;
assign w13472 = ~w6266 & w10775;
assign w13473 = ~w7886 & w5526;
assign w13474 = w13528 & ~w2044;
assign w13475 = ~w295 & ~w14213;
assign w13476 = w10676 & w2159;
assign w13477 = w14302 & ~w2508;
assign w13478 = (w9921 & w4638) | (w9921 & ~w10649) | (w4638 & ~w10649);
assign w13479 = ~w9540 & ~w3365;
assign w13480 = ~w922 & w4288;
assign w13481 = ~w10675 & ~w3036;
assign w13482 = (w5901 & w63) | (w5901 & w3933) | (w63 & w3933);
assign w13483 = (~w6521 & w12180) | (~w6521 & w13139) | (w12180 & w13139);
assign w13484 = (w5694 & ~w2692) | (w5694 & ~w7414) | (~w2692 & ~w7414);
assign w13485 = (w8018 & ~w5867) | (w8018 & w11866) | (~w5867 & w11866);
assign w13486 = (w9442 & w9624) | (w9442 & ~w4044) | (w9624 & ~w4044);
assign w13487 = (~w8851 & ~w13644) | (~w8851 & w7702) | (~w13644 & w7702);
assign w13488 = ~w11905 & w7493;
assign w13489 = w13975 & ~w4218;
assign w13490 = (w228 & w13836) | (w228 & w1765) | (w13836 & w1765);
assign w13491 = ~w2175 & w7409;
assign w13492 = ~w7369 & w3124;
assign w13493 = (~w2379 & w7594) | (~w2379 & w11556) | (w7594 & w11556);
assign w13494 = (w1498 & w2964) | (w1498 & w12311) | (w2964 & w12311);
assign w13495 = ~w3803 & ~w343;
assign w13496 = ~w13222 & w2938;
assign w13497 = (~w803 & w13587) | (~w803 & w11714) | (w13587 & w11714);
assign w13498 = ~w8895 & w435;
assign w13499 = ~w1631 & w11140;
assign w13500 = w11117 & w3400;
assign w13501 = ~w13971 & w2980;
assign w13502 = (w11734 & w8506) | (w11734 & w242) | (w8506 & w242);
assign w13503 = ~w938 & w11527;
assign w13504 = (~w13807 & w13079) | (~w13807 & w30) | (w13079 & w30);
assign w13505 = w6889 & w12311;
assign w13506 = (~w3546 & ~w1362) | (~w3546 & w649) | (~w1362 & w649);
assign w13507 = ~w2288 & w12656;
assign w13508 = (~w10941 & w5173) | (~w10941 & w11282) | (w5173 & w11282);
assign w13509 = w4909 & ~w3106;
assign w13510 = (w9268 & w5136) | (w9268 & w3116) | (w5136 & w3116);
assign w13511 = (~w12642 & w1609) | (~w12642 & w7816) | (w1609 & w7816);
assign w13512 = w10676 & w4425;
assign w13513 = ~w12604 & w1540;
assign w13514 = (~w6381 & w13587) | (~w6381 & w1435) | (w13587 & w1435);
assign w13515 = ~w5282 & w5151;
assign w13516 = (w14302 & w14307) | (w14302 & w11907) | (w14307 & w11907);
assign w13517 = (w4679 & w3293) | (w4679 & w12501) | (w3293 & w12501);
assign w13518 = w3767 & w3334;
assign w13519 = ~w8827 & ~w12915;
assign w13520 = ~w9012 & w5460;
assign w13521 = b44 & a44;
assign w13522 = ~w3914 & ~w13324;
assign w13523 = w12859 & w3476;
assign w13524 = ~w7110 & w11471;
assign w13525 = w10265 & ~w9156;
assign w13526 = ~w9453 & ~w11635;
assign w13527 = ~w7834 & w11899;
assign w13528 = ~w1351 & ~w6693;
assign w13529 = w2410 & ~w14227;
assign w13530 = ~w13324 & w14598;
assign w13531 = ~b57 & ~a57;
assign w13532 = w5707 & ~w4242;
assign w13533 = w6677 & w11766;
assign w13534 = w5522 & w4458;
assign w13535 = ~w8611 & ~w14348;
assign w13536 = w8737 & w11756;
assign w13537 = ~w5852 & w6572;
assign w13538 = (w2544 & w10561) | (w2544 & w9394) | (w10561 & w9394);
assign w13539 = (w13797 & w4578) | (w13797 & w11524) | (w4578 & w11524);
assign w13540 = ~w6193 & ~w14252;
assign w13541 = ~w10435 & w3305;
assign w13542 = ~w4865 & w4211;
assign w13543 = (~w7654 & ~w3846) | (~w7654 & ~w8580) | (~w3846 & ~w8580);
assign w13544 = w7851 & w107;
assign w13545 = w400 & w5022;
assign w13546 = w7244 & w5761;
assign w13547 = ~w10941 & w3727;
assign w13548 = (w7632 & w4272) | (w7632 & w14319) | (w4272 & w14319);
assign w13549 = w14573 & ~w9701;
assign w13550 = w13540 & ~w1762;
assign w13551 = ~w829 & ~w11855;
assign w13552 = ~w11016 & w4126;
assign w13553 = ~w4312 & w8626;
assign w13554 = w10338 & w13860;
assign w13555 = ~w6949 & ~w1712;
assign w13556 = w3160 & w8624;
assign w13557 = w7794 & w5339;
assign w13558 = w12321 & ~w14417;
assign w13559 = ~w12 & ~w10075;
assign w13560 = w3484 & ~w11998;
assign w13561 = (w9877 & w10814) | (w9877 & w4768) | (w10814 & w4768);
assign w13562 = w5590 & ~w2843;
assign w13563 = w607 & w2729;
assign w13564 = ~w12378 & w2233;
assign w13565 = ~b74 & ~a74;
assign w13566 = ~w11192 & ~w11704;
assign w13567 = ~w10523 & w13335;
assign w13568 = (w1274 & ~w3044) | (w1274 & w3750) | (~w3044 & w3750);
assign w13569 = w10997 & w5843;
assign w13570 = (~w4042 & ~w5045) | (~w4042 & w1840) | (~w5045 & w1840);
assign w13571 = ~w9363 & w14041;
assign w13572 = ~w10688 & w7271;
assign w13573 = (w10075 & ~w953) | (w10075 & w51) | (~w953 & w51);
assign w13574 = w1293 & w6500;
assign w13575 = w4803 & ~w11054;
assign w13576 = w7914 & w10708;
assign w13577 = ~w8855 & ~w10541;
assign w13578 = w3535 & w7930;
assign w13579 = (~w1623 & ~w11419) | (~w1623 & ~w13906) | (~w11419 & ~w13906);
assign w13580 = (w217 & w6423) | (w217 & w2457) | (w6423 & w2457);
assign w13581 = ~w8468 & w6370;
assign w13582 = w4387 | w10045;
assign w13583 = (~w14312 & w7896) | (~w14312 & w10229) | (w7896 & w10229);
assign w13584 = w6845 & ~w4663;
assign w13585 = (~w13338 & w7294) | (~w13338 & w3360) | (w7294 & w3360);
assign w13586 = (w3671 & w4474) | (w3671 & w1666) | (w4474 & w1666);
assign w13587 = w13750 & ~w12164;
assign w13588 = ~w3984 & w3904;
assign w13589 = w13800 & w616;
assign w13590 = ~w3075 & ~w3786;
assign w13591 = ~w13735 & ~w9359;
assign w13592 = ~w2850 & w12614;
assign w13593 = w3684 & w8000;
assign w13594 = ~w2500 & ~w7488;
assign w13595 = w11810 & ~w5569;
assign w13596 = (~w10675 & w6886) | (~w10675 & w4706) | (w6886 & w4706);
assign w13597 = ~w9760 & w2113;
assign w13598 = (~w6113 & w7850) | (~w6113 & w2994) | (w7850 & w2994);
assign w13599 = (~w13854 & w8990) | (~w13854 & w11568) | (w8990 & w11568);
assign w13600 = w5636 & w388;
assign w13601 = (~w3249 & w14473) | (~w3249 & w13966) | (w14473 & w13966);
assign w13602 = w9060 & w3564;
assign w13603 = (w730 & w10651) | (w730 & w4906) | (w10651 & w4906);
assign w13604 = (w12437 & w2348) | (w12437 & w7433) | (w2348 & w7433);
assign w13605 = (~w8283 & ~w10123) | (~w8283 & w11241) | (~w10123 & w11241);
assign w13606 = ~w9613 & ~w4483;
assign w13607 = w6592 & w12994;
assign w13608 = w13222 & w309;
assign w13609 = ~w4213 & w5732;
assign w13610 = ~b3 & ~a3;
assign w13611 = w6558 & w14468;
assign w13612 = ~w3569 & w734;
assign w13613 = (~w14146 & w2441) | (~w14146 & w6512) | (w2441 & w6512);
assign w13614 = (w12398 & w254) | (w12398 & w12447) | (w254 & w12447);
assign w13615 = (~w5694 & ~w3674) | (~w5694 & ~w11636) | (~w3674 & ~w11636);
assign w13616 = (w3025 & w4896) | (w3025 & ~w3564) | (w4896 & ~w3564);
assign w13617 = (w272 & ~w7434) | (w272 & w2698) | (~w7434 & w2698);
assign w13618 = (~w6700 & w6192) | (~w6700 & ~w2698) | (w6192 & ~w2698);
assign w13619 = w5236 & w11794;
assign w13620 = ~w2320 & ~w10704;
assign w13621 = w13658 & ~w11102;
assign w13622 = (w3430 & w5702) | (w3430 & w11253) | (w5702 & w11253);
assign w13623 = ~w12760 & ~w4800;
assign w13624 = (w6381 & w6215) | (w6381 & w7927) | (w6215 & w7927);
assign w13625 = ~w4982 & w3540;
assign w13626 = ~w13567 & w719;
assign w13627 = ~w9959 & w11386;
assign w13628 = ~w12893 & ~w45;
assign w13629 = (w10708 & w9765) | (w10708 & w1796) | (w9765 & w1796);
assign w13630 = (~w11212 & w7064) | (~w11212 & w11207) | (w7064 & w11207);
assign w13631 = (w13169 & w13844) | (w13169 & ~w12792) | (w13844 & ~w12792);
assign w13632 = ~w14015 & w5761;
assign w13633 = (~w13379 & w12670) | (~w13379 & w4053) | (w12670 & w4053);
assign w13634 = ~w6442 & w3427;
assign w13635 = w11934 & w10699;
assign w13636 = ~w2864 & ~w12429;
assign w13637 = b53 & ~w4612;
assign w13638 = w9284 & w1540;
assign w13639 = (w309 & w14141) | (w309 & w13420) | (w14141 & w13420);
assign w13640 = (w8356 & ~w13399) | (w8356 & w11707) | (~w13399 & w11707);
assign w13641 = ~w14569 & w4458;
assign w13642 = (w8007 & w2124) | (w8007 & ~w8282) | (w2124 & ~w8282);
assign w13643 = (w2029 & w2049) | (w2029 & w8011) | (w2049 & w8011);
assign w13644 = ~w14441 & w8908;
assign w13645 = w12 & ~w4360;
assign w13646 = w922 & ~w12819;
assign w13647 = ~w9118 & ~w5856;
assign w13648 = w4576 & ~w13472;
assign w13649 = w13189 & w12047;
assign w13650 = ~w2369 & ~w152;
assign w13651 = ~w9570 & ~w4233;
assign w13652 = w12809 & ~w11757;
assign w13653 = w11171 & ~w8292;
assign w13654 = ~w6750 & w3128;
assign w13655 = ~w7744 & ~w109;
assign w13656 = (w4127 & w9802) | (w4127 & w11697) | (w9802 & w11697);
assign w13657 = ~w3010 & ~w1841;
assign w13658 = (~w5287 & w7743) | (~w5287 & w10092) | (w7743 & w10092);
assign w13659 = (w11718 & w429) | (w11718 & w10501) | (w429 & w10501);
assign w13660 = (~w12575 & w5867) | (~w12575 & w11598) | (w5867 & w11598);
assign w13661 = (w1498 & w2964) | (w1498 & w3914) | (w2964 & w3914);
assign w13662 = ~w9568 & w6689;
assign w13663 = ~w1114 & ~w12868;
assign w13664 = ~w5419 & ~w4462;
assign w13665 = ~w12943 & ~w3024;
assign w13666 = ~w11255 & ~w124;
assign w13667 = ~w7376 & ~w3098;
assign w13668 = (~w884 & w1199) | (~w884 & w11921) | (w1199 & w11921);
assign w13669 = ~w4032 & ~w7821;
assign w13670 = w3550 & w5511;
assign w13671 = ~w12271 & w199;
assign w13672 = w9148 & w11050;
assign w13673 = (~w4448 & ~w6245) | (~w4448 & w13119) | (~w6245 & w13119);
assign w13674 = (~w7475 & w1615) | (~w7475 & w6063) | (w1615 & w6063);
assign w13675 = ~w10121 & ~w7402;
assign w13676 = w5556 & ~w2492;
assign w13677 = ~w13854 & w10689;
assign w13678 = (w4787 & ~w922) | (w4787 & w12925) | (~w922 & w12925);
assign w13679 = ~w5729 & ~w10590;
assign w13680 = ~w4506 & w3904;
assign w13681 = (w3215 & w12499) | (w3215 & w10508) | (w12499 & w10508);
assign w13682 = w14227 & w9170;
assign w13683 = (~w13587 & w4985) | (~w13587 & w377) | (w4985 & w377);
assign w13684 = ~w1273 & ~w4864;
assign w13685 = ~w9262 & w514;
assign w13686 = ~w10309 & w11236;
assign w13687 = ~w8226 & w5703;
assign w13688 = ~w13349 & w12064;
assign w13689 = w14396 & w11711;
assign w13690 = (w3521 & w13098) | (w3521 & ~w3907) | (w13098 & ~w3907);
assign w13691 = ~w1472 & ~w5601;
assign w13692 = w990 & w10506;
assign w13693 = w12162 & w9883;
assign w13694 = ~w12438 & ~w7906;
assign w13695 = ~w3734 & w13713;
assign w13696 = (w12952 & w9174) | (w12952 & ~w11915) | (w9174 & ~w11915);
assign w13697 = ~w10334 & ~w11402;
assign w13698 = (~w2850 & w7811) | (~w2850 & ~w12553) | (w7811 & ~w12553);
assign w13699 = ~w3137 & ~w2729;
assign w13700 = ~w1172 & w12988;
assign w13701 = ~w7276 & ~w6500;
assign w13702 = ~w12464 & ~w560;
assign w13703 = ~w7488 & w8836;
assign w13704 = ~w11465 & ~w8564;
assign w13705 = ~w3572 & ~w4037;
assign w13706 = w10974 & w12125;
assign w13707 = w1329 & ~w10815;
assign w13708 = w9454 & w4473;
assign w13709 = (~w3959 & w8441) | (~w3959 & w5278) | (w8441 & w5278);
assign w13710 = (~w622 & w5490) | (~w622 & w3670) | (w5490 & w3670);
assign w13711 = ~w4989 & w5247;
assign w13712 = ~w2144 & w11540;
assign w13713 = ~b85 & ~a85;
assign w13714 = ~w1351 & ~w6100;
assign w13715 = (~w4515 & w8693) | (~w4515 & ~w12685) | (w8693 & ~w12685);
assign w13716 = ~w6632 & ~w10483;
assign w13717 = ~w7782 & w9969;
assign w13718 = (w1498 & ~w183) | (w1498 & w2964) | (~w183 & w2964);
assign w13719 = ~w3632 & w12311;
assign w13720 = ~w11931 & w6628;
assign w13721 = w12531 & w6647;
assign w13722 = ~w4700 & w9296;
assign w13723 = ~w4700 & w1062;
assign w13724 = ~w13522 & ~w13538;
assign w13725 = ~w2164 & w5723;
assign w13726 = (~w9846 & w863) | (~w9846 & w7706) | (w863 & w7706);
assign w13727 = w14379 & w9300;
assign w13728 = w6562 & ~w6787;
assign w13729 = w9541 & ~w1923;
assign w13730 = ~w4322 & ~w14015;
assign w13731 = w4995 & ~w9058;
assign w13732 = w13839 & w13937;
assign w13733 = ~b68 & ~a68;
assign w13734 = w3175 & w7914;
assign w13735 = ~w12003 & w14076;
assign w13736 = (~w1694 & w4862) | (~w1694 & w3773) | (w4862 & w3773);
assign w13737 = (w13565 & w254) | (w13565 & w12818) | (w254 & w12818);
assign w13738 = ~w4989 & w13820;
assign w13739 = (~w13685 & w11541) | (~w13685 & w6303) | (w11541 & w6303);
assign w13740 = (~w341 & w11397) | (~w341 & w5992) | (w11397 & w5992);
assign w13741 = (w11708 & ~w1909) | (w11708 & w3809) | (~w1909 & w3809);
assign w13742 = ~w9661 & w9105;
assign w13743 = ~w8234 & ~w11261;
assign w13744 = ~w14486 & w8795;
assign w13745 = w9244 & ~w5247;
assign w13746 = (w9368 & ~w7591) | (w9368 & ~w10799) | (~w7591 & ~w10799);
assign w13747 = w7324 & ~w8980;
assign w13748 = (~w8900 & w9718) | (~w8900 & w9084) | (w9718 & w9084);
assign w13749 = ~w14659 & ~w5482;
assign w13750 = ~w11440 & w808;
assign w13751 = w2101 & w5791;
assign w13752 = (w8372 & w4471) | (w8372 & w10789) | (w4471 & w10789);
assign w13753 = ~w10221 & ~w13839;
assign w13754 = ~w3734 & w4437;
assign w13755 = (w13369 & w12310) | (w13369 & w4530) | (w12310 & w4530);
assign w13756 = ~w3038 & w7491;
assign w13757 = w14367 & ~w5105;
assign w13758 = (~w14526 & w13587) | (~w14526 & w7175) | (w13587 & w7175);
assign w13759 = w12943 & ~w473;
assign w13760 = (~w8285 & ~w10778) | (~w8285 & w1079) | (~w10778 & w1079);
assign w13761 = w9871 & w5767;
assign w13762 = w10949 & w2732;
assign w13763 = w9263 | ~w4515;
assign w13764 = ~w2509 & ~w646;
assign w13765 = (~w4479 & w6180) | (~w4479 & w1496) | (w6180 & w1496);
assign w13766 = w3632 & w6572;
assign w13767 = ~w11499 & w2982;
assign w13768 = ~w4921 & w2462;
assign w13769 = ~w5532 & ~w3044;
assign w13770 = (w7302 & w1454) | (w7302 & w9928) | (w1454 & w9928);
assign w13771 = w8626 & ~w13772;
assign w13772 = ~w14092 & w5768;
assign w13773 = w4331 & ~w11294;
assign w13774 = w11670 & ~w5909;
assign w13775 = ~w7649 & w6515;
assign w13776 = ~w2292 & w8275;
assign w13777 = w10676 & w13733;
assign w13778 = w10713 & w13837;
assign w13779 = ~w6845 & ~w2561;
assign w13780 = (~w142 & ~w13937) | (~w142 & w6872) | (~w13937 & w6872);
assign w13781 = (w12662 & w922) | (w12662 & w2037) | (w922 & w2037);
assign w13782 = (w3717 & w13152) | (w3717 & w7807) | (w13152 & w7807);
assign w13783 = w3945 & ~w2168;
assign w13784 = w4756 & w9773;
assign w13785 = ~w6845 & ~w5821;
assign w13786 = ~w10791 & w3428;
assign w13787 = (~w11091 & w7274) | (~w11091 & w2963) | (w7274 & w2963);
assign w13788 = ~w4512 & w9173;
assign w13789 = w9387 & ~w11769;
assign w13790 = w7794 & w5896;
assign w13791 = ~w12464 & w3906;
assign w13792 = ~w594 & w13456;
assign w13793 = ~w5948 & ~w12809;
assign w13794 = w7794 & w1691;
assign w13795 = w10710 & w14109;
assign w13796 = w7719 & w13606;
assign w13797 = (w2 & w8742) | (w2 & w4259) | (w8742 & w4259);
assign w13798 = w2941 & ~w11713;
assign w13799 = ~w9858 & ~w3536;
assign w13800 = ~w9097 & ~w5107;
assign w13801 = ~w4032 & w8521;
assign w13802 = ~w4787 & ~w1885;
assign w13803 = (w10276 & w2311) | (w10276 & ~w1469) | (w2311 & ~w1469);
assign w13804 = ~w2542 & w13699;
assign w13805 = w7794 & ~w2840;
assign w13806 = w7453 & ~w1943;
assign w13807 = ~w7722 & w5490;
assign w13808 = (w2310 & w9193) | (w2310 & w5147) | (w9193 & w5147);
assign w13809 = ~w8234 & ~w7762;
assign w13810 = w11488 & ~w3671;
assign w13811 = (w12952 & w9174) | (w12952 & ~w10613) | (w9174 & ~w10613);
assign w13812 = (w3540 & w3265) | (w3540 & w13625) | (w3265 & w13625);
assign w13813 = (w4515 & w12359) | (w4515 & w10585) | (w12359 & w10585);
assign w13814 = ~w9842 & ~w12063;
assign w13815 = w342 & w1374;
assign w13816 = w9181 & w4780;
assign w13817 = (w6410 & w6880) | (w6410 & w1269) | (w6880 & w1269);
assign w13818 = (w10385 & w10123) | (w10385 & w12349) | (w10123 & w12349);
assign w13819 = ~w1172 & w8;
assign w13820 = w3963 & w142;
assign w13821 = w697 & ~w6596;
assign w13822 = (w8405 & w7049) | (w8405 & w5597) | (w7049 & w5597);
assign w13823 = w14302 & w12170;
assign w13824 = ~w2601 & w4854;
assign w13825 = ~w2313 & w7925;
assign w13826 = ~w4460 & w8252;
assign w13827 = ~w12271 & w3508;
assign w13828 = ~w2500 & ~w2858;
assign w13829 = w4472 & w12311;
assign w13830 = ~w4483 & w3401;
assign w13831 = ~w3219 & w10551;
assign w13832 = ~w12271 & w6485;
assign w13833 = ~w3991 & ~w8396;
assign w13834 = (w11261 & w5573) | (w11261 & w2725) | (w5573 & w2725);
assign w13835 = ~w2674 & w14214;
assign w13836 = w4489 & w11067;
assign w13837 = ~w14310 & ~w14628;
assign w13838 = ~w12893 & ~w9871;
assign w13839 = ~w4322 & ~w4270;
assign w13840 = ~w1472 & w3124;
assign w13841 = w7331 & ~w7423;
assign w13842 = w6785 & ~w940;
assign w13843 = w10566 & w4469;
assign w13844 = w12575 & w13169;
assign w13845 = w11364 & ~w7164;
assign w13846 = w4032 & w5384;
assign w13847 = (w2655 & w4144) | (w2655 & w8227) | (w4144 & w8227);
assign w13848 = w3508 & ~w10075;
assign w13849 = (w13169 & w13844) | (w13169 & w1345) | (w13844 & w1345);
assign w13850 = (w9638 & w1828) | (w9638 & w1950) | (w1828 & w1950);
assign w13851 = ~w11351 & ~w11407;
assign w13852 = (~w4303 & w254) | (~w4303 & w2340) | (w254 & w2340);
assign w13853 = w1673 & ~w3236;
assign w13854 = ~b55 & ~a55;
assign w13855 = w6064 & w13323;
assign w13856 = w213 & w1183;
assign w13857 = w884 & w9032;
assign w13858 = ~w3209 & ~w7430;
assign w13859 = (~w13375 & ~w5498) | (~w13375 & ~w9733) | (~w5498 & ~w9733);
assign w13860 = w4167 & w2349;
assign w13861 = ~w607 & w2941;
assign w13862 = ~w9744 & ~w10020;
assign w13863 = (~w971 & ~w143) | (~w971 & ~w11759) | (~w143 & ~w11759);
assign w13864 = w475 & ~w9623;
assign w13865 = ~w14544 & ~w3290;
assign w13866 = w1802 & w13323;
assign w13867 = ~w10698 & ~w12445;
assign w13868 = w12985 | ~w11613;
assign w13869 = ~w6845 & w3502;
assign w13870 = ~w7703 & ~w8951;
assign w13871 = (~w12537 & w256) | (~w12537 & w590) | (w256 & w590);
assign w13872 = ~w3568 & ~w9145;
assign w13873 = ~w829 & ~w13854;
assign w13874 = w4291 & w8389;
assign w13875 = (~w14659 & ~w11670) | (~w14659 & w9491) | (~w11670 & w9491);
assign w13876 = ~w11776 & ~w2407;
assign w13877 = w7794 & w12130;
assign w13878 = (~w8650 & w3967) | (~w8650 & w5281) | (w3967 & w5281);
assign w13879 = w5559 & ~w2467;
assign w13880 = (w13982 & w1200) | (w13982 & w2557) | (w1200 & w2557);
assign w13881 = ~w12170 & ~w9226;
assign w13882 = ~w7625 & w13384;
assign w13883 = ~w10986 & w8445;
assign w13884 = (w5865 & ~w8234) | (w5865 & w5690) | (~w8234 & w5690);
assign w13885 = ~w5422 & w11211;
assign w13886 = w12200 & w7884;
assign w13887 = w4639 & w10481;
assign w13888 = (w13168 & w1072) | (w13168 & ~w4799) | (w1072 & ~w4799);
assign w13889 = (w6017 & w10267) | (w6017 & ~w13409) | (w10267 & ~w13409);
assign w13890 = (~w2029 & w13507) | (~w2029 & w929) | (w13507 & w929);
assign w13891 = w8742 & w13820;
assign w13892 = w14660 & w6502;
assign w13893 = (w5952 & w4747) | (w5952 & w7220) | (w4747 & w7220);
assign w13894 = ~w2680 & w2599;
assign w13895 = w2149 & w11117;
assign w13896 = ~w10435 & w6779;
assign w13897 = ~w3602 & ~w10955;
assign w13898 = (~w12406 & w13109) | (~w12406 & w2382) | (w13109 & w2382);
assign w13899 = w5817 & w3885;
assign w13900 = b124 & a124;
assign w13901 = ~w14277 & w10475;
assign w13902 = b39 & a39;
assign w13903 = (~w2428 & w13462) | (~w2428 & w12313) | (w13462 & w12313);
assign w13904 = w5490 & w10938;
assign w13905 = w10659 & ~w1836;
assign w13906 = (w3550 & w10201) | (w3550 & w9052) | (w10201 & w9052);
assign w13907 = ~w2858 & ~w5664;
assign w13908 = (w4781 & w3965) | (w4781 & w7846) | (w3965 & w7846);
assign w13909 = w1114 & w3087;
assign w13910 = w7032 & w5550;
assign w13911 = w1027 & ~w77;
assign w13912 = (~w2144 & w8915) | (~w2144 & w7327) | (w8915 & w7327);
assign w13913 = (~w4671 & ~w953) | (~w4671 & w1907) | (~w953 & w1907);
assign w13914 = ~w7801 & w8481;
assign w13915 = ~w1699 & w13657;
assign w13916 = ~w3886 & w4407;
assign w13917 = w9715 & w14227;
assign w13918 = (~w5845 & w9589) | (~w5845 & w10429) | (w9589 & w10429);
assign w13919 = w11491 & w4652;
assign w13920 = w7513 & w547;
assign w13921 = ~w142 & ~w11031;
assign w13922 = w1152 & ~w1726;
assign w13923 = w14318 & w6734;
assign w13924 = w3158 & w3038;
assign w13925 = ~w1995 & ~w8463;
assign w13926 = ~w5867 & w7811;
assign w13927 = w3427 & w636;
assign w13928 = w7772 & w7645;
assign w13929 = ~w11362 & ~w6450;
assign w13930 = ~w6676 & w7372;
assign w13931 = (w11097 & w12766) | (w11097 & w14085) | (w12766 & w14085);
assign w13932 = (~w9749 & w6484) | (~w9749 & w12722) | (w6484 & w12722);
assign w13933 = (w4353 & ~w12877) | (w4353 & w10383) | (~w12877 & w10383);
assign w13934 = w11814 & w11803;
assign w13935 = (~w9507 & ~w1362) | (~w9507 & w14581) | (~w1362 & w14581);
assign w13936 = ~w4512 & w12072;
assign w13937 = ~w12481 & ~w10221;
assign w13938 = ~w5227 & ~w608;
assign w13939 = ~w10985 & w877;
assign w13940 = w6935 & ~w12160;
assign w13941 = (~w14225 & ~w3071) | (~w14225 & w8414) | (~w3071 & w8414);
assign w13942 = w2410 & w9541;
assign w13943 = ~w2029 & w1104;
assign w13944 = (~w6362 & w11051) | (~w6362 & w3509) | (w11051 & w3509);
assign w13945 = ~w5852 & w9226;
assign w13946 = ~w2291 & ~w298;
assign w13947 = w11909 & w8389;
assign w13948 = (~w14428 & ~w10123) | (~w14428 & w550) | (~w10123 & w550);
assign w13949 = (w8584 & ~w14555) | (w8584 & w12115) | (~w14555 & w12115);
assign w13950 = ~w4032 & w13525;
assign w13951 = w4995 & ~w5973;
assign w13952 = w8417 & w3625;
assign w13953 = ~w12170 & ~w10754;
assign w13954 = ~w11462 & ~w12429;
assign w13955 = ~w507 & ~w10739;
assign w13956 = (w12569 & ~w8545) | (w12569 & w4936) | (~w8545 & w4936);
assign w13957 = ~w2320 & ~w9921;
assign w13958 = w9170 & w9919;
assign w13959 = (w11304 & w5714) | (w11304 & w8376) | (w5714 & w8376);
assign w13960 = (~w8929 & ~w2773) | (~w8929 & w2914) | (~w2773 & w2914);
assign w13961 = (w5662 & w7049) | (w5662 & w5597) | (w7049 & w5597);
assign w13962 = (w4127 & w11716) | (w4127 & w12311) | (w11716 & w12311);
assign w13963 = ~w14015 & ~w2701;
assign w13964 = w698 & w11221;
assign w13965 = (w2788 & w11712) | (w2788 & w12272) | (w11712 & w12272);
assign w13966 = (w8010 & w8519) | (w8010 & ~w12138) | (w8519 & ~w12138);
assign w13967 = w1015 & w5691;
assign w13968 = w2653 & w7914;
assign w13969 = ~w143 | ~w971;
assign w13970 = ~w7906 & w7135;
assign w13971 = w7305 & ~w10699;
assign w13972 = w8762 & w2038;
assign w13973 = w8799 & w13104;
assign w13974 = ~w3719 & w10628;
assign w13975 = w11431 & ~w12893;
assign w13976 = (w5005 & ~w4587) | (w5005 & w7074) | (~w4587 & w7074);
assign w13977 = w8475 & w2729;
assign w13978 = ~w10317 & ~w7376;
assign w13979 = ~w6233 & w8293;
assign w13980 = (~w2362 & w9832) | (~w2362 & w2052) | (w9832 & w2052);
assign w13981 = ~w4134 & w4761;
assign w13982 = ~w3288 & w8719;
assign w13983 = (~w6276 & w14353) | (~w6276 & ~w7062) | (w14353 & ~w7062);
assign w13984 = (~w3266 & w6994) | (~w3266 & w2445) | (w6994 & w2445);
assign w13985 = w11475 & ~w14054;
assign w13986 = (~w1785 & w13416) | (~w1785 & w4230) | (w13416 & w4230);
assign w13987 = ~w8768 & ~w2398;
assign w13988 = w5569 & w9087;
assign w13989 = w14031 & w10819;
assign w13990 = ~w10605 & w3995;
assign w13991 = (w8827 & w4512) | (w8827 & w9501) | (w4512 & w9501);
assign w13992 = w8183 & w7670;
assign w13993 = w10517 & ~w11117;
assign w13994 = (~w2698 & w11014) | (~w2698 & w1570) | (w11014 & w1570);
assign w13995 = ~w2774 & w2192;
assign w13996 = w13526 & ~w8992;
assign w13997 = (~w12988 & w8226) | (~w12988 & w3554) | (w8226 & w3554);
assign w13998 = w12011 & ~w7685;
assign w13999 = (w1919 & w5927) | (w1919 & w2673) | (w5927 & w2673);
assign w14000 = w2320 & ~w4541;
assign w14001 = ~w12451 & ~w1143;
assign w14002 = ~w13526 & w143;
assign w14003 = (~w4515 & w2162) | (~w4515 & w11723) | (w2162 & w11723);
assign w14004 = (w3025 & ~w14055) | (w3025 & w12041) | (~w14055 & w12041);
assign w14005 = ~w9371 & ~w13498;
assign w14006 = w2232 & ~w1821;
assign w14007 = ~w12652 & w9195;
assign w14008 = w4836 & w12893;
assign w14009 = (w1041 & ~w12434) | (w1041 & w7285) | (~w12434 & w7285);
assign w14010 = w3215 & ~w7630;
assign w14011 = ~w7782 & w3855;
assign w14012 = (~w12162 & w4374) | (~w12162 & w6313) | (w4374 & w6313);
assign w14013 = w1764 & w13745;
assign w14014 = (w11768 & w8536) | (w11768 & ~w12911) | (w8536 & ~w12911);
assign w14015 = b100 & a100;
assign w14016 = (w9244 & ~w3963) | (w9244 & w3921) | (~w3963 & w3921);
assign w14017 = ~w11849 & ~w3490;
assign w14018 = (w13334 & w6457) | (w13334 & ~w378) | (w6457 & ~w378);
assign w14019 = ~w10575 & w10542;
assign w14020 = ~w5559 & w13791;
assign w14021 = ~w7670 & w9679;
assign w14022 = w4032 & ~w13953;
assign w14023 = ~w4921 & ~w12271;
assign w14024 = ~w14338 & ~w4794;
assign w14025 = (~w4050 & w742) | (~w4050 & w6999) | (w742 & w6999);
assign w14026 = ~w4731 & w1949;
assign w14027 = w14271 & w4379;
assign w14028 = ~w2056 & ~w11409;
assign w14029 = (w7240 & w11873) | (w7240 & w8198) | (w11873 & w8198);
assign w14030 = (~w13856 & ~w6506) | (~w13856 & w4552) | (~w6506 & w4552);
assign w14031 = w13452 & ~w7793;
assign w14032 = ~w3051 & ~w1498;
assign w14033 = w7857 & ~w9353;
assign w14034 = (w10637 & w12418) | (w10637 & w4396) | (w12418 & w4396);
assign w14035 = ~w533 & w13987;
assign w14036 = w12085 & w10451;
assign w14037 = ~w13282 & w9226;
assign w14038 = ~b13 & ~a13;
assign w14039 = w7892 & w12101;
assign w14040 = w4033 & w5946;
assign w14041 = (w302 & w8848) | (w302 & w12880) | (w8848 & w12880);
assign w14042 = (w14605 & w651) | (w14605 & w604) | (w651 & w604);
assign w14043 = (w3727 & w12421) | (w3727 & w4002) | (w12421 & w4002);
assign w14044 = w14602 & w6023;
assign w14045 = (w13623 & w12900) | (w13623 & w12280) | (w12900 & w12280);
assign w14046 = (w4193 & ~w13438) | (w4193 & w1286) | (~w13438 & w1286);
assign w14047 = ~w2500 & w563;
assign w14048 = w7914 & w9921;
assign w14049 = (~w10699 & ~w3806) | (~w10699 & w5598) | (~w3806 & w5598);
assign w14050 = w7794 & ~w2334;
assign w14051 = w1658 & ~w5932;
assign w14052 = w5845 & w11902;
assign w14053 = (w3214 & w194) | (w3214 & w4653) | (w194 & w4653);
assign w14054 = ~b35 & ~a35;
assign w14055 = ~w8512 & ~w3025;
assign w14056 = ~w10139 & w13600;
assign w14057 = ~w3519 & w11617;
assign w14058 = ~w10221 & w4458;
assign w14059 = w10184 & ~w4620;
assign w14060 = w8466 & w3679;
assign w14061 = (w1607 & w5490) | (w1607 & w6887) | (w5490 & w6887);
assign w14062 = ~w4508 & w6323;
assign w14063 = ~w3727 & ~w6307;
assign w14064 = w6505 & ~w5634;
assign w14065 = ~w9315 & ~w3904;
assign w14066 = w4055 & ~w754;
assign w14067 = ~w4005 & w700;
assign w14068 = w7794 & w11;
assign w14069 = (~w5385 & w7709) | (~w5385 & ~w9668) | (w7709 & ~w9668);
assign w14070 = (~w12893 & ~w13628) | (~w12893 & w12440) | (~w13628 & w12440);
assign w14071 = w7933 & w14561;
assign w14072 = ~b76 & ~a76;
assign w14073 = ~w2824 & ~w3944;
assign w14074 = (~w12293 & w12125) | (~w12293 & w10779) | (w12125 & w10779);
assign w14075 = (~w142 & ~w2941) | (~w142 & w6872) | (~w2941 & w6872);
assign w14076 = ~w12121 & w3611;
assign w14077 = ~w14511 & ~w4366;
assign w14078 = ~w13189 & ~w1828;
assign w14079 = (~w142 & ~w6689) | (~w142 & w6872) | (~w6689 & w6872);
assign w14080 = (w154 & w5796) | (w154 & w1334) | (w5796 & w1334);
assign w14081 = w607 & ~w13323;
assign w14082 = (w8047 & w922) | (w8047 & w7923) | (w922 & w7923);
assign w14083 = (w11856 & w3202) | (w11856 & w10670) | (w3202 & w10670);
assign w14084 = (~w14578 & w274) | (~w14578 & w1307) | (w274 & w1307);
assign w14085 = (w7985 & w437) | (w7985 & w1861) | (w437 & w1861);
assign w14086 = (~w1657 & w9882) | (~w1657 & w12320) | (w9882 & w12320);
assign w14087 = ~w8841 & w3628;
assign w14088 = ~w8100 & w8080;
assign w14089 = w755 & ~w7670;
assign w14090 = (~w7190 & w1873) | (~w7190 & w4836) | (w1873 & w4836);
assign w14091 = ~w627 & w3979;
assign w14092 = w11583 & w7851;
assign w14093 = w1760 & ~w7630;
assign w14094 = (w10483 & w9978) | (w10483 & w7831) | (w9978 & w7831);
assign w14095 = (w82 & w492) | (w82 & w6578) | (w492 & w6578);
assign w14096 = (~w8130 & w899) | (~w8130 & w717) | (w899 & w717);
assign w14097 = w10146 & ~w2127;
assign w14098 = w6889 & ~w5845;
assign w14099 = w7193 & ~w2351;
assign w14100 = ~w7586 & ~w13425;
assign w14101 = (w5246 & w12498) | (w5246 & w6902) | (w12498 & w6902);
assign w14102 = (~w2941 & w4504) | (~w2941 & w8811) | (w4504 & w8811);
assign w14103 = w536 & ~w1794;
assign w14104 = ~w11747 & ~w12363;
assign w14105 = ~w1186 & ~w12730;
assign w14106 = (w7507 & w9574) | (w7507 & w12376) | (w9574 & w12376);
assign w14107 = (~w13259 & w3228) | (~w13259 & w13371) | (w3228 & w13371);
assign w14108 = ~w9921 & w1599;
assign w14109 = ~w4355 & ~w8851;
assign w14110 = (w9015 & w11261) | (w9015 & w11486) | (w11261 & w11486);
assign w14111 = w6850 & ~w5428;
assign w14112 = w4894 & w7455;
assign w14113 = (w10122 & w9541) | (w10122 & w6922) | (w9541 & w6922);
assign w14114 = ~w9728 & ~w3310;
assign w14115 = ~w3724 & w12372;
assign w14116 = w6785 & w3229;
assign w14117 = (w346 & w7318) | (w346 & ~w3266) | (w7318 & ~w3266);
assign w14118 = w7929 & w7307;
assign w14119 = ~w4094 & w9987;
assign w14120 = w791 & w4859;
assign w14121 = (~w7188 & w3756) | (~w7188 & w3518) | (w3756 & w3518);
assign w14122 = w14639 & ~w8370;
assign w14123 = w13535 & w3556;
assign w14124 = w9715 & w10916;
assign w14125 = (w7772 & w12499) | (w7772 & w6807) | (w12499 & w6807);
assign w14126 = w6572 & w5471;
assign w14127 = ~w3400 & w2654;
assign w14128 = ~w8655 & w807;
assign w14129 = ~w7609 & w2216;
assign w14130 = ~b9 & ~a9;
assign w14131 = (w13685 & w5941) | (w13685 & w14236) | (w5941 & w14236);
assign w14132 = w607 & ~w8396;
assign w14133 = ~w12481 & ~w2701;
assign w14134 = ~w12179 & ~w14641;
assign w14135 = ~w142 & ~w6689;
assign w14136 = w3730 & w10388;
assign w14137 = w12908 & ~w2081;
assign w14138 = w6592 & w8318;
assign w14139 = ~w9480 & ~w6135;
assign w14140 = w10165 & w6407;
assign w14141 = w5740 & ~w13464;
assign w14142 = (w7493 & w12271) | (w7493 & w13488) | (w12271 & w13488);
assign w14143 = ~w1822 & ~w14323;
assign w14144 = w2081 & ~w3427;
assign w14145 = w14375 & w11519;
assign w14146 = (w6502 & w6845) | (w6502 & w13416) | (w6845 & w13416);
assign w14147 = w3471 & w2895;
assign w14148 = ~w8459 & w6953;
assign w14149 = ~w5867 & w829;
assign w14150 = ~w5274 & w6811;
assign w14151 = ~w10143 & w13713;
assign w14152 = ~w11827 & ~w12614;
assign w14153 = ~w2438 & w7105;
assign w14154 = (w2652 & w8695) | (w2652 & ~w8228) | (w8695 & ~w8228);
assign w14155 = ~w607 & ~w1062;
assign w14156 = (w93 & w12527) | (w93 & w6310) | (w12527 & w6310);
assign w14157 = w5883 & ~w14640;
assign w14158 = ~w14513 & ~w2228;
assign w14159 = ~w5575 & ~w3242;
assign w14160 = (w6381 & w8769) | (w6381 & w173) | (w8769 & w173);
assign w14161 = ~w12386 & w11014;
assign w14162 = ~w2938 & ~w10853;
assign w14163 = (w3717 & w12499) | (w3717 & w11555) | (w12499 & w11555);
assign w14164 = (w7723 & w11680) | (w7723 & w2556) | (w11680 & w2556);
assign w14165 = (w8127 & w6443) | (w8127 & w2402) | (w6443 & w2402);
assign w14166 = ~w8459 & ~w9993;
assign w14167 = w7159 & w14529;
assign w14168 = ~w10435 & w11378;
assign w14169 = ~w5725 & ~w14067;
assign w14170 = w2656 & w1389;
assign w14171 = (~w695 & ~w8484) | (~w695 & ~w13309) | (~w8484 & ~w13309);
assign w14172 = ~w9893 & ~w9395;
assign w14173 = w3410 & ~w1246;
assign w14174 = ~w10853 & ~w1176;
assign w14175 = w7453 & w6500;
assign w14176 = w7943 | w7376;
assign w14177 = (~w13122 & w8533) | (~w13122 & w6841) | (w8533 & w6841);
assign w14178 = ~w5406 & ~w6572;
assign w14179 = w7376 & ~w9623;
assign w14180 = ~w254 & w542;
assign w14181 = (~w13587 & w6161) | (~w13587 & w10693) | (w6161 & w10693);
assign w14182 = (w217 & ~w11712) | (w217 & w2457) | (~w11712 & w2457);
assign w14183 = ~w6080 & ~w11117;
assign w14184 = ~b11 & ~a11;
assign w14185 = ~w6516 & w6121;
assign w14186 = w8813 & ~w6726;
assign w14187 = w3502 & w3044;
assign w14188 = (w1564 & w11161) | (w1564 & ~w11239) | (w11161 & ~w11239);
assign w14189 = (w13508 & w14411) | (w13508 & w3643) | (w14411 & w3643);
assign w14190 = w12013 & w7818;
assign w14191 = (w11895 & ~w5174) | (w11895 & w7038) | (~w5174 & w7038);
assign w14192 = (~w5852 & w3318) | (~w5852 & w9516) | (w3318 & w9516);
assign w14193 = ~w13909 & ~w10997;
assign w14194 = w10677 & w14066;
assign w14195 = ~w12271 & ~w1785;
assign w14196 = w1848 & w8964;
assign w14197 = ~w4656 & ~w10272;
assign w14198 = (w534 & w4411) | (w534 & ~w3209) | (w4411 & ~w3209);
assign w14199 = w7993 & w9777;
assign w14200 = ~w14302 & ~w5286;
assign w14201 = w2277 & w14185;
assign w14202 = ~w14614 & ~w13562;
assign w14203 = w12232 & ~w12665;
assign w14204 = ~w5047 & w2339;
assign w14205 = w4465 & w14012;
assign w14206 = w6137 & w8523;
assign w14207 = ~w11423 & ~w13816;
assign w14208 = ~w11350 & ~w12543;
assign w14209 = (w6426 & w5436) | (w6426 & w6341) | (w5436 & w6341);
assign w14210 = ~w4879 & w811;
assign w14211 = w1377 & ~w10884;
assign w14212 = (~w4134 & w9747) | (~w4134 & w4885) | (w9747 & w4885);
assign w14213 = ~w9078 & ~w5711;
assign w14214 = w11211 & w5945;
assign w14215 = ~w11216 & ~w4269;
assign w14216 = (~w5821 & w5392) | (~w5821 & w13785) | (w5392 & w13785);
assign w14217 = w7085 & w3402;
assign w14218 = w1540 & w7376;
assign w14219 = w12879 & ~w6716;
assign w14220 = ~w5294 & ~w5060;
assign w14221 = ~w5936 & ~w13960;
assign w14222 = ~w12264 & ~w5721;
assign w14223 = w8105 & w11925;
assign w14224 = ~w1840 & w3136;
assign w14225 = w10699 & ~w13302;
assign w14226 = ~w2369 & ~w14184;
assign w14227 = b76 & a76;
assign w14228 = ~w3637 & ~w7258;
assign w14229 = w2344 & ~w3165;
assign w14230 = ~w922 & w2680;
assign w14231 = ~w13302 & w8091;
assign w14232 = (~w7338 & w7169) | (~w7338 & w10667) | (w7169 & w10667);
assign w14233 = ~w13934 & w5101;
assign w14234 = (w259 & w10896) | (w259 & w14455) | (w10896 & w14455);
assign w14235 = w4733 & ~w12151;
assign w14236 = (w2722 & w14223) | (w2722 & w12376) | (w14223 & w12376);
assign w14237 = (~w4756 & w8392) | (~w4756 & w3641) | (w8392 & w3641);
assign w14238 = ~w3938 & w5402;
assign w14239 = (w2655 & w4634) | (w2655 & w7106) | (w4634 & w7106);
assign w14240 = (w6716 & w13587) | (w6716 & w6977) | (w13587 & w6977);
assign w14241 = w11309 & ~w8116;
assign w14242 = (w4202 & w2883) | (w4202 & w2287) | (w2883 & w2287);
assign w14243 = w7794 & w157;
assign w14244 = w11638 & w1479;
assign w14245 = ~w8884 & w1110;
assign w14246 = w12472 & w11007;
assign w14247 = w7685 & w5490;
assign w14248 = (~w3904 & w1726) | (~w3904 & w6875) | (w1726 & w6875);
assign w14249 = (~w3098 & ~w10699) | (~w3098 & w7083) | (~w10699 & w7083);
assign w14250 = ~w6750 & ~w5301;
assign w14251 = (~w1449 & w4490) | (~w1449 & w3908) | (w4490 & w3908);
assign w14252 = w607 & w11861;
assign w14253 = ~w7199 & ~w121;
assign w14254 = (w5952 & w906) | (w5952 & w10580) | (w906 & w10580);
assign w14255 = (~w11138 & w9942) | (~w11138 & w9934) | (w9942 & w9934);
assign w14256 = ~w781 & ~w58;
assign w14257 = (w5026 & w1187) | (w5026 & w7184) | (w1187 & w7184);
assign w14258 = w14630 & w4087;
assign w14259 = (w2829 & ~w9604) | (w2829 & w4674) | (~w9604 & w4674);
assign w14260 = (w5156 & w6328) | (w5156 & w2626) | (w6328 & w2626);
assign w14261 = ~w7488 & w6095;
assign w14262 = ~w14490 & ~w3367;
assign w14263 = ~w12202 & ~w13354;
assign w14264 = (~w14227 & w4050) | (~w14227 & w470) | (w4050 & w470);
assign w14265 = w13556 & w11698;
assign w14266 = ~w12003 & w483;
assign w14267 = w10040 & w6505;
assign w14268 = w3550 & w9596;
assign w14269 = (~w3039 & ~w7645) | (~w3039 & w10161) | (~w7645 & w10161);
assign w14270 = (w378 & w2706) | (w378 & w5027) | (w2706 & w5027);
assign w14271 = ~w13186 & w12470;
assign w14272 = w12516 & ~w4522;
assign w14273 = ~w14222 & ~w2832;
assign w14274 = (w1190 & w7015) | (w1190 & w2085) | (w7015 & w2085);
assign w14275 = ~w2864 & ~w13423;
assign w14276 = b95 & a95;
assign w14277 = ~w10730 & w8537;
assign w14278 = w205 & w10544;
assign w14279 = w5894 & ~w14101;
assign w14280 = ~w9244 & ~w473;
assign w14281 = ~w12121 & w13761;
assign w14282 = w14185 & w14578;
assign w14283 = w3508 & ~w9541;
assign w14284 = (w14453 & w4234) | (w14453 & w9707) | (w4234 & w9707);
assign w14285 = ~w4700 & w5761;
assign w14286 = ~w7772 & ~w11909;
assign w14287 = w803 & ~w7645;
assign w14288 = ~w982 & ~w8992;
assign w14289 = (~w11915 & w8880) | (~w11915 & w418) | (w8880 & w418);
assign w14290 = (~w4780 & w10913) | (~w4780 & ~w13596) | (w10913 & ~w13596);
assign w14291 = ~b25 & ~a25;
assign w14292 = ~w12553 & w4291;
assign w14293 = ~w4158 & w4836;
assign w14294 = (w1389 & w13122) | (w1389 & w14170) | (w13122 & w14170);
assign w14295 = ~w36 & ~w2773;
assign w14296 = w3303 & ~w13656;
assign w14297 = ~w71 & w3558;
assign w14298 = ~w3525 & ~w10912;
assign w14299 = ~w14302 & w14526;
assign w14300 = w5103 & ~w1974;
assign w14301 = (w8900 & w1393) | (w8900 & w2011) | (w1393 & w2011);
assign w14302 = ~w4680 & ~w8301;
assign w14303 = ~w12131 & ~w3075;
assign w14304 = ~w4751 & ~w13620;
assign w14305 = w14031 & w9913;
assign w14306 = w1250 & w10708;
assign w14307 = ~w3957 & w14486;
assign w14308 = (w7317 & w13349) | (w7317 & w8151) | (w13349 & w8151);
assign w14309 = (w319 & w4972) | (w319 & w9061) | (w4972 & w9061);
assign w14310 = ~w7244 & ~w4458;
assign w14311 = (w8390 & w10462) | (w8390 & w8206) | (w10462 & w8206);
assign w14312 = w247 & ~w4213;
assign w14313 = (~w2341 & ~w13518) | (~w2341 & ~w318) | (~w13518 & ~w318);
assign w14314 = ~w4970 & w4563;
assign w14315 = (w14360 & w9311) | (w14360 & w13172) | (w9311 & w13172);
assign w14316 = w480 & ~w13897;
assign w14317 = w10910 & ~w10996;
assign w14318 = w5687 & ~w7638;
assign w14319 = ~w9181 & w6177;
assign w14320 = (~w11198 & ~w13241) | (~w11198 & w12803) | (~w13241 & w12803);
assign w14321 = w7697 & w543;
assign w14322 = w9170 | w9289;
assign w14323 = ~w1004 & w1540;
assign w14324 = ~w8694 & w7410;
assign w14325 = ~w1099 & ~w5125;
assign w14326 = ~w13854 & w829;
assign w14327 = (w14389 & w9614) | (w14389 & w8862) | (w9614 & w8862);
assign w14328 = (~w8294 & w8016) | (~w8294 & ~w8280) | (w8016 & ~w8280);
assign w14329 = (w2405 & w1097) | (w2405 & w5718) | (w1097 & w5718);
assign w14330 = (w12605 & w14154) | (w12605 & w2670) | (w14154 & w2670);
assign w14331 = (w5282 & w9885) | (w5282 & w5629) | (w9885 & w5629);
assign w14332 = ~w29 & ~w3325;
assign w14333 = (~w7962 & w5867) | (~w7962 & w3605) | (w5867 & w3605);
assign w14334 = ~w6022 & ~w303;
assign w14335 = ~w7190 & w2486;
assign w14336 = w5337 & ~w1532;
assign w14337 = ~w11669 & w2266;
assign w14338 = (~w1172 & w13349) | (~w1172 & w13231) | (w13349 & w13231);
assign w14339 = w4213 & w4425;
assign w14340 = w2410 & w5569;
assign w14341 = (w11213 & w14421) | (w11213 & ~w8607) | (w14421 & ~w8607);
assign w14342 = ~w11488 & w4855;
assign w14343 = ~w11810 & w3851;
assign w14344 = (~w9541 & w10672) | (~w9541 & w12221) | (w10672 & w12221);
assign w14345 = ~w9732 & ~w1392;
assign w14346 = (~w353 & w4034) | (~w353 & w3489) | (w4034 & w3489);
assign w14347 = (w11261 & w249) | (w11261 & w531) | (w249 & w531);
assign w14348 = ~w3215 & ~w14504;
assign w14349 = (w6471 & w182) | (w6471 & w1945) | (w182 & w1945);
assign w14350 = w13677 & w1235;
assign w14351 = w12481 & w3904;
assign w14352 = ~w922 & ~w14070;
assign w14353 = (~w11037 & ~w9724) | (~w11037 & w318) | (~w9724 & w318);
assign w14354 = w8943 & w9936;
assign w14355 = ~w9817 & w3334;
assign w14356 = w9679 & w11455;
assign w14357 = w314 | w5654;
assign w14358 = w1949 & ~w829;
assign w14359 = (w4475 & w12287) | (w4475 & w12640) | (w12287 & w12640);
assign w14360 = w6364 & ~w4132;
assign w14361 = w4845 & w12642;
assign w14362 = w7581 | w12476;
assign w14363 = w6936 & ~w8797;
assign w14364 = w12329 & w8378;
assign w14365 = (~w12406 & w14368) | (~w12406 & w9529) | (w14368 & w9529);
assign w14366 = w2938 & ~w7423;
assign w14367 = ~w5329 & ~w12205;
assign w14368 = (w1013 & w4285) | (w1013 & ~w7644) | (w4285 & ~w7644);
assign w14369 = w1096 & w6845;
assign w14370 = ~w4540 & ~w13739;
assign w14371 = w1895 & ~w291;
assign w14372 = w9252 & w4378;
assign w14373 = (~w11261 & w13677) | (~w11261 & w14405) | (w13677 & w14405);
assign w14374 = ~w11444 & w8069;
assign w14375 = ~w13133 & w9597;
assign w14376 = (~w13219 & w1596) | (~w13219 & w10452) | (w1596 & w10452);
assign w14377 = w12482 & ~w7947;
assign w14378 = ~w7001 & ~w2729;
assign w14379 = (w11138 & w6618) | (w11138 & w769) | (w6618 & w769);
assign w14380 = ~w5626 & w1274;
assign w14381 = (~w926 & w11288) | (~w926 & w4348) | (w11288 & w4348);
assign w14382 = ~w9715 & ~w4026;
assign w14383 = (~w13337 & w3298) | (~w13337 & w3712) | (w3298 & w3712);
assign w14384 = ~w4921 & w6621;
assign w14385 = w6391 & w13129;
assign w14386 = w12464 & ~w1166;
assign w14387 = w8280 & ~w3904;
assign w14388 = w4441 & ~w2492;
assign w14389 = w343 & w8120;
assign w14390 = ~w6572 & ~w12321;
assign w14391 = ~w184 & ~w13990;
assign w14392 = (w13685 & w13366) | (w13685 & w5488) | (w13366 & w5488);
assign w14393 = w6014 & ~w12614;
assign w14394 = ~w922 & w11905;
assign w14395 = ~w5556 & ~w9226;
assign w14396 = (~w1166 & ~w9608) | (~w1166 & w14386) | (~w9608 & w14386);
assign w14397 = (~w4287 & w13587) | (~w4287 & w4412) | (w13587 & w4412);
assign w14398 = (w11488 & w71) | (w11488 & w8242) | (w71 & w8242);
assign w14399 = ~w2631 & w13097;
assign w14400 = (w9921 & ~w7926) | (w9921 & w8517) | (~w7926 & w8517);
assign w14401 = (~w4512 & w13062) | (~w4512 & w12950) | (w13062 & w12950);
assign w14402 = w2432 & w12133;
assign w14403 = (w9679 & w13508) | (w9679 & w7667) | (w13508 & w7667);
assign w14404 = ~w12543 & ~w5261;
assign w14405 = (w10689 & ~w8234) | (w10689 & w13677) | (~w8234 & w13677);
assign w14406 = w3550 & w7952;
assign w14407 = ~w12003 & w6544;
assign w14408 = ~w11444 & w4065;
assign w14409 = (w5024 & w7333) | (w5024 & w9390) | (w7333 & w9390);
assign w14410 = w12438 & ~w10483;
assign w14411 = ~w3137 & w9679;
assign w14412 = b5 & a5;
assign w14413 = w7312 & w14646;
assign w14414 = (~w5562 & w1961) | (~w5562 & w13318) | (w1961 & w13318);
assign w14415 = (w7041 & ~w10630) | (w7041 & w819) | (~w10630 & w819);
assign w14416 = w8135 & ~w1710;
assign w14417 = ~w8827 & ~w5406;
assign w14418 = (~w10676 & w8482) | (~w10676 & w1193) | (w8482 & w1193);
assign w14419 = ~w12783 & w13567;
assign w14420 = ~w861 & w646;
assign w14421 = (~w5560 & w10545) | (~w5560 & w11213) | (w10545 & w11213);
assign w14422 = w8909 & w6289;
assign w14423 = ~w4206 & ~w3876;
assign w14424 = w7612 & ~w10276;
assign w14425 = ~w1096 & ~w13909;
assign w14426 = w13445 & ~w12574;
assign w14427 = w8916 & w1528;
assign w14428 = ~w4050 & w5763;
assign w14429 = (w6637 & w6747) | (w6637 & w8730) | (w6747 & w8730);
assign w14430 = ~w11488 & ~w12065;
assign w14431 = ~w4251 & ~w4141;
assign w14432 = ~w9433 & w5626;
assign w14433 = w7703 & ~w4145;
assign w14434 = ~w11057 & ~w3093;
assign w14435 = w7012 & w6301;
assign w14436 = w6425 & w6218;
assign w14437 = ~w10676 & ~w12499;
assign w14438 = (w926 & w5657) | (w926 & w1503) | (w5657 & w1503);
assign w14439 = w13686 & ~w4741;
assign w14440 = ~w12553 & w12958;
assign w14441 = w14235 & w4070;
assign w14442 = ~w10265 & w2309;
assign w14443 = (w10523 & ~w7737) | (w10523 & w10486) | (~w7737 & w10486);
assign w14444 = w3708 & w13814;
assign w14445 = (~w2144 & w11147) | (~w2144 & w129) | (w11147 & w129);
assign w14446 = w6695 & ~w8851;
assign w14447 = (w3194 & w11238) | (w3194 & w168) | (w11238 & w168);
assign w14448 = (w7841 & w841) | (w7841 & w5379) | (w841 & w5379);
assign w14449 = w3671 & ~w9528;
assign w14450 = w309 & w8992;
assign w14451 = ~w6078 & w13427;
assign w14452 = w2656 & w9433;
assign w14453 = ~w1862 & ~w2490;
assign w14454 = (~w6554 & w9012) | (~w6554 & w1561) | (w9012 & w1561);
assign w14455 = w3447 & w10272;
assign w14456 = (w2987 & w328) | (w2987 & w2304) | (w328 & w2304);
assign w14457 = ~w5852 & w4165;
assign w14458 = w10653 & w7499;
assign w14459 = (w7861 & w2262) | (w7861 & w9874) | (w2262 & w9874);
assign w14460 = (w9305 & w529) | (w9305 & w948) | (w529 & w948);
assign w14461 = w100 & ~w13813;
assign w14462 = w9855 & ~w6500;
assign w14463 = (w9305 & w5662) | (w9305 & w8405) | (w5662 & w8405);
assign w14464 = w13222 & w12520;
assign w14465 = ~w3288 & ~w11861;
assign w14466 = w12713 & w4780;
assign w14467 = (w10290 & w8569) | (w10290 & w12311) | (w8569 & w12311);
assign w14468 = ~w11461 & w7914;
assign w14469 = ~w4213 & w12943;
assign w14470 = ~b39 & ~a39;
assign w14471 = ~w8080 & ~w3044;
assign w14472 = ~w114 & ~w6128;
assign w14473 = (~w8337 & w13339) | (~w8337 & w4579) | (w13339 & w4579);
assign w14474 = (~w11803 & w12777) | (~w11803 & w5542) | (w12777 & w5542);
assign w14475 = ~w2201 & w10704;
assign w14476 = w8019 & ~w3963;
assign w14477 = (w2788 & w6879) | (w2788 & w12272) | (w6879 & w12272);
assign w14478 = ~w536 & ~w12614;
assign w14479 = ~w13462 & w8208;
assign w14480 = ~w3914 & w12170;
assign w14481 = ~w9679 & w3017;
assign w14482 = w2606 & w4872;
assign w14483 = (w11306 & w13330) | (w11306 & w4986) | (w13330 & w4986);
assign w14484 = (~w254 & w11613) | (~w254 & w4004) | (w11613 & w4004);
assign w14485 = w7513 & w10872;
assign w14486 = ~w2159 & ~w9871;
assign w14487 = w5002 & w2850;
assign w14488 = ~w6750 & ~w5532;
assign w14489 = (w829 & w11261) | (w829 & w14637) | (w11261 & w14637);
assign w14490 = w4881 & w1540;
assign w14491 = w4700 & ~w142;
assign w14492 = ~w12611 & ~w10539;
assign w14493 = ~w3864 & ~w1325;
assign w14494 = ~w5948 & ~w4458;
assign w14495 = w11117 & w7808;
assign w14496 = ~w3914 & w12856;
assign w14497 = w11041 & w12173;
assign w14498 = w3017 & ~w13323;
assign w14499 = ~w8183 & w840;
assign w14500 = (~w9305 & w13517) | (~w9305 & w1592) | (w13517 & w1592);
assign w14501 = ~w7681 & w3427;
assign w14502 = w7794 & ~w1691;
assign w14503 = (w13937 & w3989) | (w13937 & w6879) | (w3989 & w6879);
assign w14504 = ~w3611 & ~w3717;
assign w14505 = ~w12438 & ~w8035;
assign w14506 = (~w10917 & w9655) | (~w10917 & ~w14417) | (w9655 & ~w14417);
assign w14507 = ~w10245 & w6300;
assign w14508 = (~w3823 & ~w3609) | (~w3823 & w6887) | (~w3609 & w6887);
assign w14509 = w10523 & w3427;
assign w14510 = ~w8937 & w5415;
assign w14511 = ~w4607 & w12996;
assign w14512 = ~w10853 & ~w6710;
assign w14513 = ~w7424 & w937;
assign w14514 = (w11559 & w12886) | (w11559 & w5435) | (w12886 & w5435);
assign w14515 = ~w9940 & w8513;
assign w14516 = ~w7466 & w6694;
assign w14517 = ~w11602 & w3325;
assign w14518 = w1106 & w8265;
assign w14519 = ~w7064 & ~w7281;
assign w14520 = (w11734 & w11999) | (w11734 & w7835) | (w11999 & w7835);
assign w14521 = w14115 & ~w8761;
assign w14522 = (~w4050 & w7230) | (~w4050 & w7932) | (w7230 & w7932);
assign w14523 = ~w10077 & w13968;
assign w14524 = w5761 & w9927;
assign w14525 = w14293 & ~w13265;
assign w14526 = b85 & a85;
assign w14527 = ~w13375 & w5176;
assign w14528 = (w12889 & w1750) | (w12889 & w6760) | (w1750 & w6760);
assign w14529 = ~w7161 & w7914;
assign w14530 = (w8000 & ~w5931) | (w8000 & w13593) | (~w5931 & w13593);
assign w14531 = w6464 & w10775;
assign w14532 = w10039 & w6439;
assign w14533 = ~w7423 & ~w11600;
assign w14534 = ~w12463 & ~w14421;
assign w14535 = ~w10431 & w13323;
assign w14536 = ~w3790 & w5742;
assign w14537 = w10158 & w2274;
assign w14538 = w1235 & ~w5874;
assign w14539 = w6562 & w5260;
assign w14540 = w10095 & w497;
assign w14541 = w12920 & ~w5060;
assign w14542 = w9788 & w2270;
assign w14543 = ~w8691 & ~w5605;
assign w14544 = (w2611 & w12251) | (w2611 & w13729) | (w12251 & w13729);
assign w14545 = (w12941 & w14175) | (w12941 & w13418) | (w14175 & w13418);
assign w14546 = (~w3215 & w5867) | (~w3215 & w12575) | (w5867 & w12575);
assign w14547 = (~w14372 & ~w2065) | (~w14372 & w12959) | (~w2065 & w12959);
assign w14548 = (w1712 & w6678) | (w1712 & w4682) | (w6678 & w4682);
assign w14549 = w4541 & w13285;
assign w14550 = w7582 & ~w12259;
assign w14551 = ~w10629 & w12344;
assign w14552 = (~w13654 & w9397) | (~w13654 & w7048) | (w9397 & w7048);
assign w14553 = ~w11507 & ~w7535;
assign w14554 = ~w2500 & w4627;
assign w14555 = ~w14369 & w13666;
assign w14556 = w12464 & w4738;
assign w14557 = w1767 & w11480;
assign w14558 = ~w2161 & ~w1541;
assign w14559 = ~w499 & w6739;
assign w14560 = w3094 & ~w6489;
assign w14561 = ~w13817 & ~w4696;
assign w14562 = w13651 | ~w4233;
assign w14563 = ~w7391 & ~w8594;
assign w14564 = w11108 & w4132;
assign w14565 = w11492 & ~w1769;
assign w14566 = (w1658 & w3699) | (w1658 & w2890) | (w3699 & w2890);
assign w14567 = ~w12148 & w10692;
assign w14568 = (w12761 & w6221) | (w12761 & w9034) | (w6221 & w9034);
assign w14569 = ~w4270 & ~w10517;
assign w14570 = w509 & ~w12642;
assign w14571 = ~w2144 & w10415;
assign w14572 = (w12460 & w183) | (w12460 & w8660) | (w183 & w8660);
assign w14573 = ~w10477 & ~w4017;
assign w14574 = w3636 & w11117;
assign w14575 = w4138 & ~w10301;
assign w14576 = w7670 & ~w11684;
assign w14577 = (~w12398 & w4623) | (~w12398 & w391) | (w4623 & w391);
assign w14578 = ~w1563 & ~w5702;
assign w14579 = w9300 & ~w10062;
assign w14580 = ~w4512 & w4139;
assign w14581 = (~w3215 & w9012) | (~w3215 & w14546) | (w9012 & w14546);
assign w14582 = (w12642 & w2997) | (w12642 & w11614) | (w2997 & w11614);
assign w14583 = (w8937 & w8817) | (w8937 & w227) | (w8817 & w227);
assign w14584 = ~w13761 & ~w1260;
assign w14585 = ~w8058 & ~w502;
assign w14586 = ~w14054 & w13375;
assign w14587 = (w11979 & w1137) | (w11979 & w14123) | (w1137 & w14123);
assign w14588 = ~b121 & ~a121;
assign w14589 = ~w607 & w1540;
assign w14590 = w8018 & w12954;
assign w14591 = ~w11931 & w10802;
assign w14592 = w2607 & w5148;
assign w14593 = (w8786 & w11650) | (w8786 & ~w353) | (w11650 & ~w353);
assign w14594 = w7270 & w12401;
assign w14595 = w10676 & w14390;
assign w14596 = ~w13349 & w10029;
assign w14597 = (~w13219 & w7900) | (~w13219 & w11359) | (w7900 & w11359);
assign w14598 = ~w3914 & w3524;
assign w14599 = (w14059 & w5159) | (w14059 & w3721) | (w5159 & w3721);
assign w14600 = w768 & ~w4582;
assign w14601 = w8655 | ~w807;
assign w14602 = (~w378 & w6568) | (~w378 & w9538) | (w6568 & w9538);
assign w14603 = w10045 & ~w4327;
assign w14604 = (w1455 & w12771) | (w1455 & w694) | (w12771 & w694);
assign w14605 = w10177 & w10100;
assign w14606 = (~w8692 & w11860) | (~w8692 & w3005) | (w11860 & w3005);
assign w14607 = ~w4015 & w2893;
assign w14608 = w14302 & w7085;
assign w14609 = (w13685 & w7948) | (w13685 & w1400) | (w7948 & w1400);
assign w14610 = (w4627 & w10462) | (w4627 & w2882) | (w10462 & w2882);
assign w14611 = w10014 & w3076;
assign w14612 = w8297 & ~w9614;
assign w14613 = ~w12575 & ~w10917;
assign w14614 = b111 & a111;
assign w14615 = (~w11091 & w6210) | (~w11091 & w4802) | (w6210 & w4802);
assign w14616 = w5741 & w12642;
assign w14617 = (~w12376 & w1850) | (~w12376 & w14520) | (w1850 & w14520);
assign w14618 = (w13462 & w4160) | (w13462 & w11892) | (w4160 & w11892);
assign w14619 = ~w10783 & ~w8188;
assign w14620 = w3957 & ~w3672;
assign w14621 = ~w6529 & w8568;
assign w14622 = (w4041 & w13589) | (w4041 & w5517) | (w13589 & w5517);
assign w14623 = w7400 & ~w690;
assign w14624 = ~w1949 & ~w9181;
assign w14625 = ~w4700 & w7113;
assign w14626 = ~w7961 & ~w1482;
assign w14627 = ~w11030 & w13241;
assign w14628 = w7244 & w4458;
assign w14629 = ~w7754 & ~w2081;
assign w14630 = (w3128 & w10273) | (w3128 & w6532) | (w10273 & w6532);
assign w14631 = w8121 & w12982;
assign w14632 = (~w11429 & w1512) | (~w11429 & w12049) | (w1512 & w12049);
assign w14633 = ~w12856 & w1919;
assign w14634 = (~w4515 & w9263) | (~w4515 & w3759) | (w9263 & w3759);
assign w14635 = w12464 & w12170;
assign w14636 = w9145 & ~w10408;
assign w14637 = w8234 & w829;
assign w14638 = w8201 & w13050;
assign w14639 = b14 & a14;
assign w14640 = (~w8475 & w2707) | (~w8475 & w912) | (w2707 & w912);
assign w14641 = (w9305 & w264) | (w9305 & w212) | (w264 & w212);
assign w14642 = ~w4158 & w2055;
assign w14643 = ~w2189 & ~w7768;
assign w14644 = ~w5635 & w14144;
assign w14645 = (w2486 & w1692) | (w2486 & w8877) | (w1692 & w8877);
assign w14646 = ~w5422 & ~w5785;
assign w14647 = w10409 & w4185;
assign w14648 = ~w10360 & ~w6983;
assign w14649 = w2653 & w8975;
assign w14650 = (~w10272 & ~w7464) | (~w10272 & w5926) | (~w7464 & w5926);
assign w14651 = w8018 & w12068;
assign w14652 = w7512 & w6585;
assign w14653 = ~w3914 & ~w9246;
assign w14654 = ~w11510 & ~w2500;
assign w14655 = w9170 & w11011;
assign w14656 = w6626 & ~w1665;
assign w14657 = w13854 & ~w1692;
assign w14658 = (w3039 & ~w14302) | (w3039 & w7324) | (~w14302 & w7324);
assign w14659 = ~w4312 & ~w6041;
assign w14660 = ~w5406 & ~w11395;
assign w14661 = (w8512 & w12637) | (w8512 & w9715) | (w12637 & w9715);
assign w14662 = ~w14054 & ~w5754;
assign w14663 = w4372 & ~w1364;
assign w14664 = (~w3550 & w10940) | (~w3550 & w1659) | (w10940 & w1659);
assign w14665 = (w13595 & w3818) | (w13595 & w143) | (w3818 & w143);
assign w14666 = ~w12716 & ~w2761;
assign w14667 = (w12376 & w14044) | (w12376 & w4451) | (w14044 & w4451);
assign w14668 = ~w9667 & w1607;
assign w14669 = (~w2159 & w1166) | (~w2159 & w14486) | (w1166 & w14486);
assign w14670 = ~w12271 & w11810;
assign w14671 = w13831 & w7857;
assign one = 1;
assign s0 = w4104;// level 5
assign s1 = w188;// level 5
assign s2 = ~w964;// level 6
assign s3 = w11879;// level 6
assign s4 = w5840;// level 6
assign s5 = w8818;// level 7
assign s6 = w2860;// level 7
assign s7 = w1763;// level 7
assign s8 = ~w3910;// level 7
assign s9 = w12026;// level 8
assign s10 = ~w10293;// level 8
assign s11 = ~w4264;// level 8
assign s12 = ~w12111;// level 8
assign s13 = w14431;// level 8
assign s14 = w7974;// level 8
assign s15 = w8333;// level 8
assign s16 = ~w4422;// level 8
assign s17 = ~w9068;// level 9
assign s18 = ~w6731;// level 9
assign s19 = w115;// level 9
assign s20 = w1684;// level 9
assign s21 = ~w3031;// level 9
assign s22 = w14134;// level 9
assign s23 = ~w5250;// level 9
assign s24 = ~w5430;// level 9
assign s25 = ~w5065;// level 9
assign s26 = w12752;// level 10
assign s27 = ~w13298;// level 10
assign s28 = w4020;// level 10
assign s29 = ~w193;// level 10
assign s30 = w7976;// level 10
assign s31 = ~w8134;// level 10
assign s32 = ~w3654;// level 10
assign s33 = ~w11563;// level 10
assign s34 = w4829;// level 10
assign s35 = ~w5427;// level 10
assign s36 = w8014;// level 10
assign s37 = w949;// level 11
assign s38 = ~w7095;// level 11
assign s39 = ~w6664;// level 11
assign s40 = w8317;// level 11
assign s41 = ~w7246;// level 11
assign s42 = w4156;// level 11
assign s43 = ~w13705;// level 11
assign s44 = w6353;// level 12
assign s45 = ~w1210;// level 11
assign s46 = w13106;// level 11
assign s47 = w4630;// level 11
assign s48 = w12465;// level 11
assign s49 = ~w11611;// level 11
assign s50 = w10933;// level 12
assign s51 = w1341;// level 11
assign s52 = w633;// level 13
assign s53 = w12675;// level 13
assign s54 = w5833;// level 13
assign s55 = ~w9020;// level 13
assign s56 = w4012;// level 13
assign s57 = ~w3066;// level 14
assign s58 = w4301;// level 13
assign s59 = ~w3063;// level 13
assign s60 = w6552;// level 13
assign s61 = ~w8156;// level 13
assign s62 = w131;// level 13
assign s63 = ~w2497;// level 13
assign s64 = w5258;// level 13
assign s65 = ~w14370;// level 13
assign s66 = w8358;// level 13
assign s67 = ~w14298;// level 13
assign s68 = w2051;// level 13
assign s69 = ~w10836;// level 13
assign s70 = w13252;// level 13
assign s71 = ~w6102;// level 13
assign s72 = w13571;// level 13
assign s73 = ~w1511;// level 13
assign s74 = w11072;// level 14
assign s75 = ~w5812;// level 13
assign s76 = ~w12579;// level 13
assign s77 = w12323;// level 13
assign s78 = w2524;// level 14
assign s79 = ~w13164;// level 13
assign s80 = w10865;// level 13
assign s81 = ~w72;// level 13
assign s82 = w6154;// level 13
assign s83 = ~w6616;// level 13
assign s84 = w9260;// level 13
assign s85 = ~w7054;// level 13
assign s86 = w1562;// level 14
assign s87 = ~w8833;// level 13
assign s88 = w5459;// level 15
assign s89 = w3046;// level 13
assign s90 = w9955;// level 14
assign s91 = ~w10262;// level 13
assign s92 = w8207;// level 14
assign s93 = ~w6595;// level 13
assign s94 = w656;// level 14
assign s95 = ~w9975;// level 17
assign s96 = w5928;// level 17
assign s97 = ~w4788;// level 17
assign s98 = w1370;// level 17
assign s99 = w10616;// level 16
assign s100 = w5085;// level 18
assign s101 = w11717;// level 18
assign s102 = w13036;// level 18
assign s103 = w4950;// level 17
assign s104 = ~w6424;// level 17
assign s105 = ~w8486;// level 19
assign s106 = w4113;// level 17
assign s107 = ~w4882;// level 17
assign s108 = ~w14169;// level 17
assign s109 = w2026;// level 17
assign s110 = w10051;// level 16
assign s111 = w7298;// level 18
assign s112 = w7651;// level 17
assign s113 = w12024;// level 17
assign s114 = w8375;// level 17
assign s115 = w1253;// level 18
assign s116 = ~w8216;// level 17
assign s117 = ~w10138;// level 17
assign s118 = w11995;// level 19
assign s119 = ~w6968;// level 18
assign s120 = w7903;// level 17
assign s121 = w10237;// level 18
assign s122 = w10060;// level 17
assign s123 = ~w10697;// level 18
assign s124 = w6625;// level 17
assign s125 = w5876;// level 18
assign s126 = w12500;// level 18
assign s127 = ~w10025;// level 17
assign s128 = ~w3416;// level 14
endmodule
