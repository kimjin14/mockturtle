module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 ;
  wire n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 ;
  assign n61 = x20 | x21 ;
  assign n62 = x22 | n61 ;
  assign n63 = x23 & n62 ;
  assign n64 = x24 & n63 ;
  assign n65 = x25 | x26 ;
  assign n66 = x27 & x28 ;
  assign n67 = n65 & n66 ;
  assign n68 = x29 & n67 ;
  assign n69 = x26 & x27 ;
  assign n70 = x28 & x29 ;
  assign n71 = n69 & n70 ;
  assign n72 = ( n64 & n68 ) | ( n64 & n71 ) | ( n68 & n71 ) ;
  assign n73 = x21 | x22 ;
  assign n74 = x23 & x24 ;
  assign n75 = n73 & n74 ;
  assign n76 = ( n68 & n71 ) | ( n68 & n75 ) | ( n71 & n75 ) ;
  assign n77 = x17 | x18 ;
  assign n78 = x9 | x10 ;
  assign n79 = x11 & n78 ;
  assign n80 = x12 | n79 ;
  assign n81 = x13 | n80 ;
  assign n82 = x14 | n81 ;
  assign n83 = ~x14 & n82 ;
  assign n84 = ( ~n81 & n82 ) | ( ~n81 & n83 ) | ( n82 & n83 ) ;
  assign n85 = ( x14 & n80 ) | ( x14 & ~n84 ) | ( n80 & ~n84 ) ;
  assign n86 = x15 & n85 ;
  assign n87 = x16 & x17 ;
  assign n88 = x18 | n87 ;
  assign n89 = ( n77 & n86 ) | ( n77 & n88 ) | ( n86 & n88 ) ;
  assign n90 = x19 & n89 ;
  assign n91 = ( n72 & n76 ) | ( n72 & n90 ) | ( n76 & n90 ) ;
  assign n92 = x27 & n65 ;
  assign n93 = ( n64 & n69 ) | ( n64 & n92 ) | ( n69 & n92 ) ;
  assign n94 = ( n69 & n75 ) | ( n69 & n92 ) | ( n75 & n92 ) ;
  assign n95 = ( n90 & n93 ) | ( n90 & n94 ) | ( n93 & n94 ) ;
  assign n96 = x27 | n65 ;
  assign n97 = x26 | x27 ;
  assign n98 = ( n64 & n96 ) | ( n64 & n97 ) | ( n96 & n97 ) ;
  assign n99 = ( n75 & n96 ) | ( n75 & n97 ) | ( n96 & n97 ) ;
  assign n100 = ( n90 & n98 ) | ( n90 & n99 ) | ( n98 & n99 ) ;
  assign n101 = ~n95 & n100 ;
  assign n102 = x28 & ~n69 ;
  assign n103 = x28 & ~n92 ;
  assign n104 = ( ~n64 & n102 ) | ( ~n64 & n103 ) | ( n102 & n103 ) ;
  assign n105 = ( ~n75 & n102 ) | ( ~n75 & n103 ) | ( n102 & n103 ) ;
  assign n106 = ( ~n90 & n104 ) | ( ~n90 & n105 ) | ( n104 & n105 ) ;
  assign n107 = ~x28 & n69 ;
  assign n108 = ( ~x28 & n92 ) | ( ~x28 & n103 ) | ( n92 & n103 ) ;
  assign n109 = ( n64 & n107 ) | ( n64 & n108 ) | ( n107 & n108 ) ;
  assign n110 = ( n75 & n107 ) | ( n75 & n108 ) | ( n107 & n108 ) ;
  assign n111 = ( n90 & n109 ) | ( n90 & n110 ) | ( n109 & n110 ) ;
  assign n112 = n106 | n111 ;
  assign n113 = n101 | n112 ;
  assign n114 = ~x9 & n91 ;
  assign n115 = ( n91 & n113 ) | ( n91 & n114 ) | ( n113 & n114 ) ;
  assign n116 = x1 | x2 ;
  assign n117 = x3 | x4 ;
  assign n118 = n116 | n117 ;
  assign n119 = x5 | x6 ;
  assign n120 = x7 | n119 ;
  assign n121 = n118 | n120 ;
  assign n122 = x9 & x10 ;
  assign n123 = n78 & ~n122 ;
  assign n124 = ~x8 & n123 ;
  assign n125 = ~n121 & n124 ;
  assign n126 = x11 | n78 ;
  assign n127 = ~n79 & n126 ;
  assign n128 = x11 & x12 ;
  assign n129 = n78 & n128 ;
  assign n130 = n80 & ~n129 ;
  assign n131 = ~n127 & n130 ;
  assign n132 = n125 & n131 ;
  assign n133 = x13 & n80 ;
  assign n134 = n81 & ~n133 ;
  assign n135 = ~n84 & n134 ;
  assign n136 = n132 & n135 ;
  assign n137 = x16 | n86 ;
  assign n138 = x16 & n86 ;
  assign n139 = n137 & ~n138 ;
  assign n140 = x15 & ~n86 ;
  assign n141 = ( n85 & ~n86 ) | ( n85 & n140 ) | ( ~n86 & n140 ) ;
  assign n142 = n139 & ~n141 ;
  assign n143 = n136 & n142 ;
  assign n144 = x19 | n77 ;
  assign n145 = ( x19 & n88 ) | ( x19 & n144 ) | ( n88 & n144 ) ;
  assign n146 = ( n86 & n144 ) | ( n86 & n145 ) | ( n144 & n145 ) ;
  assign n147 = ~n90 & n146 ;
  assign n148 = ( x17 & n86 ) | ( x17 & n87 ) | ( n86 & n87 ) ;
  assign n149 = x18 & n148 ;
  assign n150 = n89 & ~n149 ;
  assign n151 = x17 | n137 ;
  assign n152 = ~x17 & n151 ;
  assign n153 = ( ~n137 & n151 ) | ( ~n137 & n152 ) | ( n151 & n152 ) ;
  assign n154 = n150 & ~n153 ;
  assign n155 = ~n147 & n154 ;
  assign n156 = n143 & n155 ;
  assign n157 = ( n62 & n73 ) | ( n62 & n90 ) | ( n73 & n90 ) ;
  assign n158 = x20 & n90 ;
  assign n159 = x21 & n158 ;
  assign n160 = x21 & ~n159 ;
  assign n161 = ( x22 & n158 ) | ( x22 & n160 ) | ( n158 & n160 ) ;
  assign n162 = n157 & ~n161 ;
  assign n163 = x20 & ~n158 ;
  assign n164 = ( n90 & ~n158 ) | ( n90 & n163 ) | ( ~n158 & n163 ) ;
  assign n165 = ( n158 & ~n159 ) | ( n158 & n160 ) | ( ~n159 & n160 ) ;
  assign n166 = ~n164 & n165 ;
  assign n167 = n162 & n166 ;
  assign n168 = n156 & n167 ;
  assign n169 = x23 & n73 ;
  assign n170 = ( n63 & n90 ) | ( n63 & n169 ) | ( n90 & n169 ) ;
  assign n171 = x23 | n73 ;
  assign n172 = n61 | n171 ;
  assign n173 = ( n90 & n171 ) | ( n90 & n172 ) | ( n171 & n172 ) ;
  assign n174 = ~n170 & n173 ;
  assign n175 = x24 & n170 ;
  assign n176 = x24 & ~n175 ;
  assign n177 = ( n170 & ~n175 ) | ( n170 & n176 ) | ( ~n175 & n176 ) ;
  assign n178 = n174 | n177 ;
  assign n179 = ( x26 & n64 ) | ( x26 & n65 ) | ( n64 & n65 ) ;
  assign n180 = ( x26 & n65 ) | ( x26 & n75 ) | ( n65 & n75 ) ;
  assign n181 = ( n90 & n179 ) | ( n90 & n180 ) | ( n179 & n180 ) ;
  assign n182 = x25 & x26 ;
  assign n183 = ( n64 & n75 ) | ( n64 & n90 ) | ( n75 & n90 ) ;
  assign n184 = n182 & n183 ;
  assign n185 = n181 & ~n184 ;
  assign n186 = x25 & n183 ;
  assign n187 = x25 & ~n186 ;
  assign n188 = ( n183 & ~n186 ) | ( n183 & n187 ) | ( ~n186 & n187 ) ;
  assign n189 = n185 & ~n188 ;
  assign n190 = ~n178 & n189 ;
  assign n191 = ( n115 & n168 ) | ( n115 & n190 ) | ( n168 & n190 ) ;
  assign n192 = ( n91 & n115 ) | ( n91 & ~n191 ) | ( n115 & ~n191 ) ;
  assign n193 = ~x29 & n67 ;
  assign n194 = x28 & ~x29 ;
  assign n195 = n69 & n194 ;
  assign n196 = ( n64 & n193 ) | ( n64 & n195 ) | ( n193 & n195 ) ;
  assign n197 = ( n75 & n193 ) | ( n75 & n195 ) | ( n193 & n195 ) ;
  assign n198 = ( n90 & n196 ) | ( n90 & n197 ) | ( n196 & n197 ) ;
  assign n199 = x29 & ~n67 ;
  assign n200 = ( x29 & ~n69 ) | ( x29 & n107 ) | ( ~n69 & n107 ) ;
  assign n201 = ( ~n64 & n199 ) | ( ~n64 & n200 ) | ( n199 & n200 ) ;
  assign n202 = ( ~n75 & n199 ) | ( ~n75 & n200 ) | ( n199 & n200 ) ;
  assign n203 = ( ~n90 & n201 ) | ( ~n90 & n202 ) | ( n201 & n202 ) ;
  assign n204 = n198 | n203 ;
  assign n205 = ~x9 & n204 ;
  assign n206 = n101 & n112 ;
  assign n207 = n205 & n206 ;
  assign n208 = ~n185 & n188 ;
  assign n209 = n177 & n208 ;
  assign n210 = n207 & n209 ;
  assign n211 = ~n162 & n174 ;
  assign n212 = n164 & ~n165 ;
  assign n213 = n211 & n212 ;
  assign n214 = n147 & n213 ;
  assign n215 = ~n150 & n153 ;
  assign n216 = ~n139 & n141 ;
  assign n217 = n215 & n216 ;
  assign n218 = n84 & ~n134 ;
  assign n219 = ~n130 & n218 ;
  assign n220 = n217 & n219 ;
  assign n221 = n214 & n220 ;
  assign n222 = n210 & n221 ;
  assign n223 = x0 | n91 ;
  assign n224 = x8 & ~n123 ;
  assign n225 = n127 & n224 ;
  assign n226 = x6 & x7 ;
  assign n227 = x5 & n226 ;
  assign n228 = x4 & n227 ;
  assign n229 = x3 & n228 ;
  assign n230 = n225 & n229 ;
  assign n231 = x1 & x2 ;
  assign n232 = n230 & n231 ;
  assign n233 = ( n91 & n223 ) | ( n91 & n232 ) | ( n223 & n232 ) ;
  assign n234 = ( n91 & n222 ) | ( n91 & n233 ) | ( n222 & n233 ) ;
  assign n235 = ~n192 & n234 ;
  assign n236 = x50 | x51 ;
  assign n237 = x52 | n236 ;
  assign n238 = x53 & n237 ;
  assign n239 = x54 & n238 ;
  assign n240 = x56 & x57 ;
  assign n241 = x58 & x59 ;
  assign n242 = n240 & n241 ;
  assign n243 = x55 | x56 ;
  assign n244 = x57 & n243 ;
  assign n245 = ( n241 & n242 ) | ( n241 & n244 ) | ( n242 & n244 ) ;
  assign n246 = ( n239 & n242 ) | ( n239 & n245 ) | ( n242 & n245 ) ;
  assign n247 = x51 | x52 ;
  assign n248 = x53 & x54 ;
  assign n249 = n247 & n248 ;
  assign n250 = ( n242 & n245 ) | ( n242 & n249 ) | ( n245 & n249 ) ;
  assign n251 = x47 | x48 ;
  assign n252 = x39 | x40 ;
  assign n253 = x41 & n252 ;
  assign n254 = x42 | n253 ;
  assign n255 = x43 | n254 ;
  assign n256 = x44 | n255 ;
  assign n257 = ~x44 & n256 ;
  assign n258 = ( ~n255 & n256 ) | ( ~n255 & n257 ) | ( n256 & n257 ) ;
  assign n259 = ( x44 & n254 ) | ( x44 & ~n258 ) | ( n254 & ~n258 ) ;
  assign n260 = x45 & n259 ;
  assign n261 = x46 & x47 ;
  assign n262 = x48 | n261 ;
  assign n263 = ( n251 & n260 ) | ( n251 & n262 ) | ( n260 & n262 ) ;
  assign n264 = x49 & n263 ;
  assign n265 = ( n246 & n250 ) | ( n246 & n264 ) | ( n250 & n264 ) ;
  assign n266 = x0 & ~n265 ;
  assign n267 = ~n192 & n266 ;
  assign n268 = x58 & ~n240 ;
  assign n269 = x58 & ~n244 ;
  assign n270 = ( ~n239 & n268 ) | ( ~n239 & n269 ) | ( n268 & n269 ) ;
  assign n271 = ( ~n249 & n268 ) | ( ~n249 & n269 ) | ( n268 & n269 ) ;
  assign n272 = ( ~n264 & n270 ) | ( ~n264 & n271 ) | ( n270 & n271 ) ;
  assign n273 = ~x58 & n240 ;
  assign n274 = ( ~x58 & n244 ) | ( ~x58 & n269 ) | ( n244 & n269 ) ;
  assign n275 = ( n239 & n273 ) | ( n239 & n274 ) | ( n273 & n274 ) ;
  assign n276 = ( n249 & n273 ) | ( n249 & n274 ) | ( n273 & n274 ) ;
  assign n277 = ( n264 & n275 ) | ( n264 & n276 ) | ( n275 & n276 ) ;
  assign n278 = n272 | n277 ;
  assign n279 = x30 & ~x39 ;
  assign n280 = x59 & n279 ;
  assign n281 = n278 & n280 ;
  assign n282 = ( x56 & n239 ) | ( x56 & n243 ) | ( n239 & n243 ) ;
  assign n283 = ( x56 & n243 ) | ( x56 & n249 ) | ( n243 & n249 ) ;
  assign n284 = ( n264 & n282 ) | ( n264 & n283 ) | ( n282 & n283 ) ;
  assign n285 = ( n239 & n249 ) | ( n239 & n264 ) | ( n249 & n264 ) ;
  assign n286 = x55 & x56 ;
  assign n287 = n285 & n286 ;
  assign n288 = n284 & ~n287 ;
  assign n289 = ( n239 & n240 ) | ( n239 & n244 ) | ( n240 & n244 ) ;
  assign n290 = ( n240 & n244 ) | ( n240 & n249 ) | ( n244 & n249 ) ;
  assign n291 = ( n264 & n289 ) | ( n264 & n290 ) | ( n289 & n290 ) ;
  assign n292 = x57 | n243 ;
  assign n293 = x56 | x57 ;
  assign n294 = ( n239 & n292 ) | ( n239 & n293 ) | ( n292 & n293 ) ;
  assign n295 = ( n249 & n292 ) | ( n249 & n293 ) | ( n292 & n293 ) ;
  assign n296 = ( n264 & n294 ) | ( n264 & n295 ) | ( n294 & n295 ) ;
  assign n297 = ~n291 & n296 ;
  assign n298 = ~n288 & n297 ;
  assign n299 = n281 & n298 ;
  assign n300 = x53 & n247 ;
  assign n301 = ( n238 & n264 ) | ( n238 & n300 ) | ( n264 & n300 ) ;
  assign n302 = x53 | n247 ;
  assign n303 = n236 | n302 ;
  assign n304 = ( n264 & n302 ) | ( n264 & n303 ) | ( n302 & n303 ) ;
  assign n305 = ~n301 & n304 ;
  assign n306 = x55 & n285 ;
  assign n307 = x55 & ~n306 ;
  assign n308 = ( n285 & ~n306 ) | ( n285 & n307 ) | ( ~n306 & n307 ) ;
  assign n309 = x54 & n301 ;
  assign n310 = x54 & ~n309 ;
  assign n311 = ( n301 & ~n309 ) | ( n301 & n310 ) | ( ~n309 & n310 ) ;
  assign n312 = n308 & n311 ;
  assign n313 = n305 & n312 ;
  assign n314 = n299 & n313 ;
  assign n315 = ( x47 & n260 ) | ( x47 & n261 ) | ( n260 & n261 ) ;
  assign n316 = x48 & n315 ;
  assign n317 = n263 & ~n316 ;
  assign n318 = x49 | n251 ;
  assign n319 = ( x49 & n262 ) | ( x49 & n318 ) | ( n262 & n318 ) ;
  assign n320 = ( n260 & n318 ) | ( n260 & n319 ) | ( n318 & n319 ) ;
  assign n321 = ~n264 & n320 ;
  assign n322 = x50 & n264 ;
  assign n323 = x50 & ~n322 ;
  assign n324 = ( n264 & ~n322 ) | ( n264 & n323 ) | ( ~n322 & n323 ) ;
  assign n325 = ~n247 & n324 ;
  assign n326 = n321 & n325 ;
  assign n327 = ~n317 & n326 ;
  assign n328 = n314 & n327 ;
  assign n329 = x41 | n252 ;
  assign n330 = ~n253 & n329 ;
  assign n331 = x41 & x42 ;
  assign n332 = n252 & n331 ;
  assign n333 = n254 & ~n332 ;
  assign n334 = x43 & n254 ;
  assign n335 = n255 & ~n334 ;
  assign n336 = x46 | n260 ;
  assign n337 = x46 & n260 ;
  assign n338 = n336 & ~n337 ;
  assign n339 = x47 | n336 ;
  assign n340 = ~x47 & n339 ;
  assign n341 = ( ~n336 & n339 ) | ( ~n336 & n340 ) | ( n339 & n340 ) ;
  assign n342 = ~n338 & n341 ;
  assign n343 = x45 & ~n260 ;
  assign n344 = ( n259 & ~n260 ) | ( n259 & n343 ) | ( ~n260 & n343 ) ;
  assign n345 = n342 & n344 ;
  assign n346 = n258 & n345 ;
  assign n347 = ~n335 & n346 ;
  assign n348 = ~n333 & n347 ;
  assign n349 = n330 & n348 ;
  assign n350 = n328 & n349 ;
  assign n351 = n278 | n297 ;
  assign n352 = ~x39 & n265 ;
  assign n353 = ( n265 & n351 ) | ( n265 & n352 ) | ( n351 & n352 ) ;
  assign n354 = x31 | x32 ;
  assign n355 = x33 | x34 ;
  assign n356 = n354 | n355 ;
  assign n357 = x35 | x36 ;
  assign n358 = x37 | n357 ;
  assign n359 = n356 | n358 ;
  assign n360 = x39 & x40 ;
  assign n361 = n252 & ~n360 ;
  assign n362 = ~x38 & n361 ;
  assign n363 = ~n359 & n362 ;
  assign n364 = ~n330 & n333 ;
  assign n365 = n363 & n364 ;
  assign n366 = ~n258 & n335 ;
  assign n367 = n365 & n366 ;
  assign n368 = n338 & ~n344 ;
  assign n369 = n367 & n368 ;
  assign n370 = n317 & ~n341 ;
  assign n371 = ~n321 & n370 ;
  assign n372 = n369 & n371 ;
  assign n373 = x51 & n322 ;
  assign n374 = x51 & ~n373 ;
  assign n375 = ( n322 & ~n373 ) | ( n322 & n374 ) | ( ~n373 & n374 ) ;
  assign n376 = ~n324 & n375 ;
  assign n377 = ~x52 & n376 ;
  assign n378 = n372 & n377 ;
  assign n379 = n305 | n311 ;
  assign n380 = n288 & ~n308 ;
  assign n381 = ~n379 & n380 ;
  assign n382 = ( n353 & n378 ) | ( n353 & n381 ) | ( n378 & n381 ) ;
  assign n383 = ( n265 & n353 ) | ( n265 & ~n382 ) | ( n353 & ~n382 ) ;
  assign n384 = x38 & ~n361 ;
  assign n385 = x37 & n384 ;
  assign n386 = x36 & n385 ;
  assign n387 = x35 & n386 ;
  assign n388 = x34 & n387 ;
  assign n389 = x33 & n388 ;
  assign n390 = x32 & n389 ;
  assign n391 = x31 & n390 ;
  assign n392 = n383 | n391 ;
  assign n393 = ( n350 & n383 ) | ( n350 & n392 ) | ( n383 & n392 ) ;
  assign n394 = x0 | x30 ;
  assign n395 = n265 & n394 ;
  assign n396 = n393 | n395 ;
  assign n397 = n234 & n396 ;
  assign n398 = ( n192 & ~n267 ) | ( n192 & n397 ) | ( ~n267 & n397 ) ;
  assign n399 = x0 & x30 ;
  assign n400 = ( n265 & n383 ) | ( n265 & n399 ) | ( n383 & n399 ) ;
  assign n401 = n235 & n400 ;
  assign y0 = ~n235 ;
  assign y1 = ~n398 ;
  assign y2 = n401 ;
  assign y3 = 1'b0 ;
  assign y4 = 1'b0 ;
  assign y5 = 1'b0 ;
  assign y6 = 1'b0 ;
  assign y7 = 1'b0 ;
  assign y8 = 1'b0 ;
  assign y9 = 1'b0 ;
  assign y10 = 1'b0 ;
  assign y11 = 1'b0 ;
  assign y12 = 1'b0 ;
  assign y13 = 1'b0 ;
  assign y14 = 1'b0 ;
  assign y15 = 1'b0 ;
  assign y16 = 1'b0 ;
  assign y17 = 1'b0 ;
  assign y18 = 1'b0 ;
  assign y19 = 1'b0 ;
  assign y20 = 1'b0 ;
  assign y21 = 1'b0 ;
  assign y22 = 1'b0 ;
  assign y23 = 1'b0 ;
  assign y24 = 1'b0 ;
  assign y25 = 1'b0 ;
  assign y26 = 1'b0 ;
  assign y27 = 1'b0 ;
  assign y28 = 1'b0 ;
  assign y29 = 1'b0 ;
endmodule
