//Written by the Majority Logic Package Fri Nov 14 22:11:54 2014
module top (
            pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09, pi10, pi11, pi12, pi13, pi14, pi15, pi16, pi17, pi18, pi19, pi20, pi21, pi22, pi23, pi24, pi25, pi26, pi27, pi28, pi29, pi30, pi31, pi32, pi33, pi34, pi35, pi36, pi37, pi38, pi39, pi40, pi41, pi42, pi43, pi44, pi45, pi46, pi47, pi48, pi49, pi50, pi51, pi52, pi53, pi54, pi55, pi56, pi57, pi58, pi59, pi60, pi61, pi62, pi63, pi64, pi65, pi66, pi67, pi68, pi69, pi70, pi71, pi72, pi73, pi74, pi75, pi76, pi77, pi78, pi79, pi80, pi81, pi82, pi83, pi84, pi85, pi86, pi87, pi88, pi89, pi90, pi91, pi92, pi93, pi94, pi95, 
            po00, po01, po02, po03, po04, po05, po06, po07, po08, po09, po10, po11, po12, po13, po14, po15, po16, po17, po18, po19, po20, po21, po22, po23, po24, po25, po26, po27, po28, po29, po30, po31);
input pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09, pi10, pi11, pi12, pi13, pi14, pi15, pi16, pi17, pi18, pi19, pi20, pi21, pi22, pi23, pi24, pi25, pi26, pi27, pi28, pi29, pi30, pi31, pi32, pi33, pi34, pi35, pi36, pi37, pi38, pi39, pi40, pi41, pi42, pi43, pi44, pi45, pi46, pi47, pi48, pi49, pi50, pi51, pi52, pi53, pi54, pi55, pi56, pi57, pi58, pi59, pi60, pi61, pi62, pi63, pi64, pi65, pi66, pi67, pi68, pi69, pi70, pi71, pi72, pi73, pi74, pi75, pi76, pi77, pi78, pi79, pi80, pi81, pi82, pi83, pi84, pi85, pi86, pi87, pi88, pi89, pi90, pi91, pi92, pi93, pi94, pi95;
output po00, po01, po02, po03, po04, po05, po06, po07, po08, po09, po10, po11, po12, po13, po14, po15, po16, po17, po18, po19, po20, po21, po22, po23, po24, po25, po26, po27, po28, po29, po30, po31;
wire one, w0, w1, w2, w3, w4, w5, w6, w7, w8, w9, w10, w11, w12, w13, w14, w15, w16, w17, w18, w19, w20, w21, w22, w23, w24, w25, w26, w27, w28, w29, w30, w31, w32, w33, w34, w35, w36, w37, w38, w39, w40, w41, w42, w43, w44, w45, w46, w47, w48, w49, w50, w51, w52, w53, w54, w55, w56, w57, w58, w59, w60, w61, w62, w63, w64, w65, w66, w67, w68, w69, w70, w71, w72, w73, w74, w75, w76, w77, w78, w79, w80, w81, w82, w83, w84, w85, w86, w87, w88, w89, w90, w91, w92, w93, w94, w95, w96, w97, w98, w99, w100, w101, w102, w103, w104, w105, w106, w107, w108, w109, w110, w111, w112, w113, w114, w115, w116, w117, w118, w119, w120, w121, w122, w123, w124, w125, w126, w127, w128, w129, w130, w131, w132, w133, w134, w135, w136, w137, w138, w139, w140, w141, w142, w143, w144, w145, w146, w147, w148, w149, w150, w151, w152, w153, w154, w155, w156, w157, w158, w159, w160, w161, w162, w163, w164, w165, w166, w167, w168, w169, w170, w171, w172, w173, w174, w175, w176, w177, w178, w179, w180, w181, w182, w183, w184, w185, w186, w187, w188, w189, w190, w191, w192, w193, w194, w195, w196, w197, w198, w199, w200, w201, w202, w203, w204, w205, w206, w207, w208, w209, w210, w211, w212, w213, w214, w215, w216, w217, w218, w219, w220, w221, w222, w223, w224, w225, w226, w227, w228, w229, w230, w231, w232, w233, w234, w235, w236, w237, w238, w239, w240, w241, w242, w243, w244, w245, w246, w247, w248, w249, w250, w251, w252, w253, w254, w255, w256, w257, w258, w259, w260, w261, w262, w263, w264, w265, w266, w267, w268, w269, w270, w271, w272, w273, w274, w275, w276, w277, w278, w279, w280, w281, w282, w283, w284, w285, w286, w287, w288, w289, w290, w291, w292, w293, w294, w295, w296, w297, w298, w299, w300, w301, w302, w303, w304, w305, w306, w307, w308, w309, w310, w311, w312, w313, w314, w315, w316, w317, w318, w319, w320, w321, w322, w323, w324, w325, w326, w327, w328, w329, w330, w331, w332, w333, w334, w335, w336, w337, w338, w339, w340, w341, w342, w343, w344, w345, w346, w347, w348, w349, w350, w351, w352, w353, w354, w355, w356, w357, w358, w359, w360, w361, w362, w363, w364, w365, w366, w367, w368, w369, w370, w371, w372, w373, w374, w375, w376, w377, w378, w379, w380, w381, w382, w383, w384, w385, w386, w387, w388, w389, w390, w391, w392, w393, w394, w395, w396, w397, w398, w399, w400, w401, w402, w403, w404, w405, w406, w407, w408, w409, w410, w411, w412, w413, w414, w415, w416, w417, w418, w419, w420, w421, w422, w423, w424, w425, w426, w427, w428, w429, w430, w431, w432, w433, w434, w435, w436, w437, w438, w439, w440, w441, w442, w443, w444, w445, w446, w447, w448, w449, w450, w451, w452, w453, w454, w455, w456, w457, w458, w459, w460, w461, w462, w463, w464, w465, w466, w467, w468, w469, w470, w471, w472, w473, w474, w475, w476, w477, w478, w479, w480, w481, w482, w483, w484, w485, w486, w487, w488, w489, w490, w491, w492, w493, w494, w495, w496, w497, w498, w499, w500, w501, w502, w503, w504, w505, w506, w507, w508, w509, w510, w511, w512, w513, w514, w515, w516, w517, w518, w519, w520, w521, w522, w523, w524, w525, w526, w527, w528, w529, w530, w531, w532, w533, w534, w535, w536, w537, w538, w539, w540, w541, w542, w543, w544, w545, w546, w547, w548, w549, w550, w551, w552, w553, w554, w555, w556, w557, w558, w559, w560, w561, w562, w563, w564, w565, w566, w567, w568, w569, w570, w571, w572, w573, w574, w575, w576, w577, w578, w579, w580, w581, w582, w583, w584, w585, w586, w587, w588, w589, w590, w591, w592, w593, w594, w595, w596, w597, w598, w599, w600, w601, w602, w603, w604, w605, w606, w607, w608, w609, w610, w611, w612, w613, w614, w615, w616, w617, w618, w619, w620, w621, w622, w623, w624, w625, w626, w627, w628, w629, w630, w631, w632, w633, w634, w635, w636, w637, w638, w639, w640, w641, w642, w643, w644, w645, w646, w647, w648, w649, w650, w651, w652, w653, w654, w655, w656, w657, w658, w659, w660, w661, w662, w663, w664, w665, w666, w667, w668, w669, w670, w671, w672, w673, w674, w675, w676, w677, w678, w679, w680, w681, w682, w683, w684, w685, w686, w687, w688, w689, w690, w691, w692, w693, w694, w695, w696, w697, w698, w699, w700, w701, w702, w703, w704, w705, w706, w707, w708, w709, w710, w711, w712, w713, w714, w715, w716, w717, w718, w719, w720, w721, w722, w723, w724, w725, w726, w727, w728, w729, w730, w731, w732, w733, w734, w735, w736, w737, w738, w739, w740, w741, w742, w743, w744, w745, w746, w747, w748, w749, w750, w751, w752, w753, w754, w755, w756, w757, w758, w759, w760, w761, w762, w763, w764, w765, w766, w767, w768, w769, w770, w771, w772, w773, w774, w775, w776, w777, w778, w779, w780, w781, w782, w783, w784, w785, w786, w787, w788, w789, w790, w791, w792, w793, w794, w795, w796, w797, w798, w799, w800, w801, w802, w803, w804, w805, w806, w807, w808, w809, w810, w811, w812, w813, w814, w815, w816, w817, w818, w819, w820, w821, w822, w823, w824, w825, w826, w827, w828, w829, w830, w831, w832, w833, w834, w835, w836, w837, w838, w839, w840, w841, w842, w843, w844, w845, w846, w847, w848, w849, w850, w851, w852, w853, w854, w855, w856, w857, w858, w859, w860, w861, w862, w863, w864, w865, w866, w867, w868, w869, w870, w871, w872, w873, w874, w875, w876, w877, w878, w879, w880, w881, w882, w883, w884, w885, w886, w887, w888, w889, w890, w891, w892, w893, w894, w895, w896, w897, w898, w899, w900, w901, w902, w903, w904, w905, w906, w907, w908, w909, w910, w911, w912, w913, w914, w915, w916, w917, w918, w919, w920, w921, w922, w923, w924, w925, w926, w927, w928, w929, w930, w931, w932, w933, w934, w935, w936, w937, w938, w939, w940, w941, w942, w943, w944, w945, w946, w947, w948, w949, w950, w951, w952, w953, w954, w955, w956, w957, w958, w959, w960, w961, w962, w963, w964, w965, w966, w967, w968, w969, w970, w971, w972, w973, w974, w975, w976, w977, w978, w979, w980, w981, w982, w983, w984, w985, w986, w987, w988, w989, w990, w991, w992, w993, w994, w995, w996, w997, w998, w999, w1000, w1001, w1002, w1003, w1004, w1005, w1006, w1007, w1008, w1009, w1010, w1011, w1012, w1013, w1014, w1015, w1016, w1017, w1018, w1019, w1020, w1021, w1022, w1023, w1024, w1025, w1026, w1027, w1028, w1029, w1030, w1031, w1032, w1033, w1034, w1035, w1036, w1037, w1038, w1039, w1040, w1041, w1042, w1043, w1044, w1045, w1046, w1047, w1048, w1049, w1050, w1051, w1052, w1053, w1054, w1055, w1056, w1057, w1058, w1059, w1060, w1061, w1062, w1063, w1064, w1065, w1066, w1067, w1068, w1069, w1070, w1071, w1072, w1073, w1074, w1075, w1076, w1077, w1078, w1079, w1080, w1081, w1082, w1083, w1084, w1085, w1086, w1087, w1088, w1089, w1090, w1091, w1092, w1093, w1094, w1095, w1096, w1097, w1098, w1099, w1100, w1101, w1102, w1103, w1104, w1105, w1106, w1107, w1108, w1109, w1110, w1111, w1112, w1113, w1114, w1115, w1116, w1117, w1118, w1119, w1120, w1121, w1122, w1123, w1124, w1125, w1126, w1127, w1128, w1129, w1130, w1131, w1132, w1133, w1134, w1135, w1136, w1137, w1138, w1139, w1140, w1141, w1142, w1143, w1144, w1145, w1146, w1147, w1148, w1149, w1150, w1151, w1152, w1153, w1154, w1155, w1156, w1157, w1158, w1159, w1160, w1161, w1162, w1163, w1164, w1165, w1166, w1167, w1168, w1169, w1170, w1171, w1172, w1173, w1174, w1175, w1176, w1177, w1178, w1179, w1180, w1181, w1182, w1183, w1184, w1185, w1186, w1187, w1188, w1189, w1190, w1191, w1192, w1193, w1194, w1195, w1196, w1197, w1198, w1199, w1200, w1201, w1202, w1203, w1204, w1205, w1206, w1207, w1208, w1209, w1210, w1211, w1212, w1213, w1214, w1215, w1216, w1217, w1218, w1219, w1220, w1221, w1222, w1223, w1224, w1225, w1226, w1227, w1228, w1229, w1230, w1231, w1232, w1233, w1234, w1235, w1236, w1237, w1238, w1239, w1240, w1241, w1242, w1243, w1244, w1245, w1246, w1247, w1248, w1249, w1250, w1251, w1252, w1253, w1254, w1255, w1256, w1257, w1258, w1259, w1260, w1261, w1262, w1263, w1264, w1265, w1266, w1267, w1268, w1269, w1270, w1271, w1272, w1273, w1274, w1275, w1276, w1277, w1278, w1279, w1280, w1281, w1282, w1283, w1284, w1285, w1286, w1287, w1288, w1289, w1290, w1291, w1292, w1293, w1294, w1295, w1296, w1297, w1298, w1299, w1300, w1301, w1302, w1303, w1304, w1305, w1306, w1307, w1308, w1309, w1310, w1311, w1312, w1313, w1314, w1315, w1316, w1317, w1318, w1319, w1320, w1321, w1322, w1323, w1324, w1325, w1326, w1327, w1328, w1329, w1330, w1331, w1332, w1333, w1334, w1335, w1336, w1337, w1338, w1339, w1340, w1341, w1342, w1343, w1344, w1345, w1346, w1347, w1348, w1349, w1350, w1351, w1352, w1353, w1354, w1355, w1356, w1357, w1358, w1359, w1360, w1361, w1362, w1363, w1364, w1365, w1366, w1367, w1368, w1369, w1370, w1371, w1372, w1373, w1374, w1375, w1376, w1377, w1378, w1379, w1380, w1381, w1382, w1383, w1384, w1385, w1386, w1387, w1388, w1389, w1390, w1391, w1392, w1393, w1394, w1395, w1396, w1397, w1398, w1399, w1400, w1401, w1402, w1403, w1404, w1405, w1406, w1407, w1408, w1409, w1410, w1411, w1412, w1413, w1414, w1415, w1416, w1417, w1418, w1419, w1420, w1421, w1422, w1423, w1424, w1425, w1426, w1427, w1428, w1429, w1430, w1431, w1432, w1433, w1434, w1435, w1436, w1437, w1438, w1439, w1440, w1441, w1442, w1443, w1444, w1445, w1446, w1447, w1448, w1449, w1450, w1451, w1452, w1453, w1454, w1455, w1456, w1457, w1458, w1459, w1460, w1461, w1462, w1463, w1464, w1465, w1466, w1467, w1468, w1469, w1470, w1471, w1472, w1473, w1474, w1475, w1476, w1477, w1478, w1479, w1480, w1481, w1482, w1483, w1484, w1485, w1486, w1487, w1488, w1489, w1490, w1491, w1492, w1493, w1494, w1495, w1496, w1497, w1498, w1499, w1500, w1501, w1502, w1503, w1504, w1505, w1506, w1507, w1508, w1509, w1510, w1511, w1512, w1513, w1514, w1515, w1516, w1517, w1518, w1519, w1520, w1521, w1522, w1523, w1524, w1525, w1526, w1527, w1528, w1529, w1530, w1531, w1532, w1533, w1534, w1535, w1536, w1537, w1538, w1539, w1540, w1541, w1542, w1543, w1544, w1545, w1546, w1547, w1548, w1549, w1550, w1551, w1552, w1553, w1554, w1555, w1556, w1557, w1558, w1559, w1560, w1561, w1562, w1563, w1564, w1565, w1566, w1567, w1568, w1569, w1570, w1571, w1572, w1573, w1574, w1575, w1576, w1577, w1578, w1579, w1580, w1581, w1582, w1583, w1584, w1585, w1586, w1587, w1588, w1589, w1590, w1591, w1592, w1593, w1594, w1595, w1596, w1597, w1598, w1599, w1600, w1601, w1602, w1603, w1604, w1605, w1606, w1607, w1608, w1609, w1610, w1611, w1612, w1613, w1614, w1615, w1616, w1617, w1618, w1619, w1620, w1621, w1622, w1623, w1624, w1625, w1626, w1627, w1628, w1629, w1630, w1631, w1632, w1633, w1634, w1635, w1636, w1637, w1638, w1639, w1640, w1641, w1642, w1643, w1644, w1645, w1646, w1647, w1648, w1649, w1650, w1651, w1652, w1653, w1654, w1655, w1656, w1657, w1658, w1659, w1660, w1661, w1662, w1663, w1664, w1665, w1666, w1667, w1668, w1669, w1670, w1671, w1672, w1673, w1674, w1675, w1676, w1677, w1678, w1679, w1680, w1681, w1682, w1683, w1684, w1685, w1686, w1687, w1688, w1689, w1690, w1691, w1692, w1693, w1694, w1695, w1696, w1697, w1698, w1699, w1700, w1701, w1702, w1703, w1704, w1705, w1706, w1707, w1708, w1709, w1710, w1711, w1712, w1713, w1714, w1715, w1716, w1717, w1718, w1719, w1720, w1721, w1722, w1723, w1724, w1725, w1726, w1727, w1728, w1729, w1730, w1731, w1732, w1733, w1734, w1735, w1736, w1737, w1738, w1739, w1740, w1741, w1742, w1743, w1744, w1745, w1746, w1747, w1748, w1749, w1750, w1751, w1752, w1753, w1754, w1755, w1756, w1757, w1758, w1759, w1760, w1761, w1762, w1763, w1764, w1765, w1766, w1767, w1768, w1769, w1770, w1771, w1772, w1773, w1774, w1775, w1776, w1777, w1778, w1779, w1780, w1781, w1782, w1783, w1784, w1785, w1786, w1787, w1788, w1789, w1790, w1791, w1792, w1793, w1794, w1795, w1796, w1797, w1798, w1799, w1800, w1801, w1802, w1803, w1804, w1805, w1806, w1807, w1808, w1809, w1810, w1811, w1812, w1813, w1814, w1815, w1816, w1817, w1818, w1819, w1820, w1821, w1822, w1823, w1824, w1825, w1826, w1827, w1828, w1829, w1830, w1831, w1832, w1833, w1834, w1835, w1836, w1837, w1838, w1839, w1840, w1841, w1842, w1843, w1844, w1845, w1846, w1847, w1848, w1849, w1850, w1851, w1852, w1853, w1854, w1855, w1856, w1857, w1858, w1859, w1860, w1861, w1862, w1863, w1864, w1865, w1866, w1867, w1868, w1869, w1870, w1871, w1872, w1873, w1874, w1875, w1876, w1877, w1878, w1879, w1880, w1881, w1882, w1883, w1884, w1885, w1886, w1887, w1888, w1889, w1890, w1891, w1892, w1893, w1894, w1895, w1896, w1897, w1898, w1899, w1900, w1901, w1902, w1903, w1904, w1905, w1906, w1907, w1908, w1909, w1910, w1911, w1912, w1913, w1914, w1915, w1916, w1917, w1918, w1919, w1920, w1921, w1922, w1923, w1924, w1925, w1926, w1927, w1928, w1929, w1930, w1931, w1932, w1933, w1934, w1935, w1936, w1937;
assign w0 = ~w1337 & ~w1536;
assign w1 = ~w820 & ~w1771;
assign w2 = (w1751 & w1200) | (w1751 & w904) | (w1200 & w904);
assign w3 = (w1358 & w270) | (w1358 & w194) | (w270 & w194);
assign w4 = (pi77 & w399) | (pi77 & w836) | (w399 & w836);
assign w5 = (w1358 & w239) | (w1358 & w917) | (w239 & w917);
assign w6 = w1199 & ~w1326;
assign w7 = (w987 & w1492) | (w987 & w462) | (w1492 & w462);
assign w8 = (w1209 & w382) | (w1209 & ~w1600) | (w382 & ~w1600);
assign w9 = (~w1021 & w973) | (~w1021 & w1145) | (w973 & w1145);
assign w10 = ~w1886 & ~w455;
assign w11 = ~pi92 & ~w722;
assign w12 = ~w121 & ~w628;
assign w13 = w1207 & w1701;
assign w14 = pi56 & w1262;
assign w15 = ~w925 & w1881;
assign w16 = ~w501 & ~w202;
assign w17 = (w1304 & w1392) | (w1304 & ~w1021) | (w1392 & ~w1021);
assign w18 = (w1737 & w204) | (w1737 & w1358) | (w204 & w1358);
assign w19 = (w1633 & w1420) | (w1633 & ~w247) | (w1420 & ~w247);
assign w20 = w290 & ~w610;
assign w21 = pi78 & ~pi79;
assign w22 = w1760 & ~w1500;
assign w23 = w854 & w869;
assign w24 = (w937 & w1441) | (w937 & ~w1351) | (w1441 & ~w1351);
assign w25 = ~pi32 & ~w1231;
assign w26 = w1337 & ~w1248;
assign w27 = ~w1594 & ~w1573;
assign w28 = w1737 & w1176;
assign w29 = (w59 & w1905) | (w59 & w1520) | (w1905 & w1520);
assign w30 = (~w105 & w548) | (~w105 & ~w1500) | (w548 & ~w1500);
assign w31 = w1309 & ~w1816;
assign w32 = ~w334 & ~w1434;
assign w33 = (w48 & w1555) | (w48 & w268) | (w1555 & w268);
assign w34 = w1841 & ~w434;
assign w35 = w1510 & ~w1902;
assign w36 = (w1803 & w257) | (w1803 & w864) | (w257 & w864);
assign w37 = w366 & ~w507;
assign w38 = (~w576 & w886) | (~w576 & w446) | (w886 & w446);
assign w39 = (w1272 & w1531) | (w1272 & w647) | (w1531 & w647);
assign w40 = pi53 & ~w941;
assign w41 = ~w883 & ~w970;
assign w42 = pi00 & ~w959;
assign w43 = ~pi81 & ~pi82;
assign w44 = (w1491 & w3) | (w1491 & w78) | (w3 & w78);
assign w45 = ~w51 & w1113;
assign w46 = ~w487 & w1205;
assign w47 = (w1491 & w1025) | (w1491 & w1897) | (w1025 & w1897);
assign w48 = (w247 & w429) | (w247 & w738) | (w429 & w738);
assign w49 = ~w1764 & ~w1111;
assign w50 = (w1856 & w1447) | (w1856 & w350) | (w1447 & w350);
assign w51 = (w1540 & w1866) | (w1540 & w1256) | (w1866 & w1256);
assign w52 = (w1817 & w1518) | (w1817 & w667) | (w1518 & w667);
assign w53 = (w1805 & w375) | (w1805 & ~w694) | (w375 & ~w694);
assign w54 = (w525 & w442) | (w525 & w865) | (w442 & w865);
assign w55 = w173 & ~pi47;
assign w56 = ~w1771 & w820;
assign w57 = (~w247 & w368) | (~w247 & w1088) | (w368 & w1088);
assign w58 = ~w1649 & ~w1017;
assign w59 = (w1142 & w615) | (w1142 & w1313) | (w615 & w1313);
assign w60 = pi30 & pi31;
assign w61 = (w424 & w1327) | (w424 & w48) | (w1327 & w48);
assign w62 = (w694 & w151) | (w694 & w559) | (w151 & w559);
assign w63 = w69 & w1307;
assign w64 = (~w723 & w780) | (~w723 & w1891) | (w780 & w1891);
assign w65 = (w1540 & w1124) | (w1540 & w1705) | (w1124 & w1705);
assign w66 = (w997 & w469) | (w997 & w62) | (w469 & w62);
assign w67 = ~w924 & ~w980;
assign w68 = (w1193 & w1045) | (w1193 & ~w865) | (w1045 & ~w865);
assign w69 = ~w1261 & w72;
assign w70 = (~pi92 & w1335) | (~pi92 & w923) | (w1335 & w923);
assign w71 = ~w1510 & ~pi77;
assign w72 = ~w1622 & ~pi17;
assign w73 = (w1437 & w386) | (w1437 & w16) | (w386 & w16);
assign w74 = w1575 & pi47;
assign w75 = (~w1491 & w17) | (~w1491 & w409) | (w17 & w409);
assign w76 = (w1669 & w614) | (w1669 & ~w48) | (w614 & ~w48);
assign w77 = (w576 & w1683) | (w576 & w283) | (w1683 & w283);
assign w78 = (w48 & w270) | (w48 & w194) | (w270 & w194);
assign w79 = (~w1575 & w1889) | (~w1575 & w316) | (w1889 & w316);
assign w80 = ~w1593 & ~w729;
assign w81 = (pi26 & w1496) | (pi26 & w724) | (w1496 & w724);
assign w82 = w390 & ~w1930;
assign w83 = (~w1147 & w839) | (~w1147 & w1475) | (w839 & w1475);
assign w84 = w877 & ~pi03;
assign w85 = w1886 & ~pi74;
assign w86 = ~w399 & ~w812;
assign w87 = (w1443 & ~w758) | (w1443 & ~w1549) | (~w758 & ~w1549);
assign w88 = (w568 & w1120) | (w568 & w1013) | (w1120 & w1013);
assign w89 = pi42 & pi43;
assign w90 = pi36 & pi37;
assign w91 = w1446 & w1247;
assign w92 = (~w1915 & w475) | (~w1915 & w815) | (w475 & w815);
assign w93 = ~pi36 & pi37;
assign w94 = w992 & pi11;
assign w95 = (~w304 & w370) | (~w304 & w1387) | (w370 & w1387);
assign w96 = (w1715 & w771) | (w1715 & w1003) | (w771 & w1003);
assign w97 = (~w105 & w548) | (~w105 & w1708) | (w548 & w1708);
assign w98 = (w869 & ~w419) | (w869 & w181) | (~w419 & w181);
assign w99 = (w1156 & w1610) | (w1156 & ~w1358) | (w1610 & ~w1358);
assign w100 = ~w1838 & ~w526;
assign w101 = ~w60 & ~w1915;
assign w102 = ~w1766 & ~w1810;
assign w103 = ~w66 & ~w1107;
assign w104 = ~w1310 & ~w1011;
assign w105 = ~w398 & ~w43;
assign w106 = ~w1804 & w799;
assign w107 = (w1888 & w25) | (w1888 & ~w1480) | (w25 & ~w1480);
assign w108 = (~w1 & w1251) | (~w1 & w1065) | (w1251 & w1065);
assign w109 = (~w1499 & w1850) | (~w1499 & w969) | (w1850 & w969);
assign w110 = (w415 & w309) | (w415 & ~w1773) | (w309 & ~w1773);
assign w111 = ~w1246 & w387;
assign w112 = pi12 & ~pi13;
assign w113 = (w578 & w750) | (w578 & ~w1358) | (w750 & ~w1358);
assign w114 = (~w1207 & w1788) | (~w1207 & ~w1915) | (w1788 & ~w1915);
assign w115 = (w997 & w1026) | (w997 & w1373) | (w1026 & w1373);
assign w116 = (w1491 & w1079) | (w1491 & w1191) | (w1079 & w1191);
assign w117 = (w636 & w406) | (w636 & ~w1849) | (w406 & ~w1849);
assign w118 = (~pi47 & w286) | (~pi47 & w1395) | (w286 & w1395);
assign w119 = ~w992 & ~w1499;
assign w120 = (~w958 & w777) | (~w958 & w1185) | (w777 & w1185);
assign w121 = pi14 & w580;
assign w122 = w1326 & w664;
assign w123 = ~w1178 & ~w132;
assign w124 = (~w1856 & w1818) | (~w1856 & ~w1858) | (w1818 & ~w1858);
assign w125 = (w1138 & w74) | (w1138 & w1440) | (w74 & w1440);
assign w126 = (~w1491 & w1075) | (~w1491 & w1405) | (w1075 & w1405);
assign w127 = (~w925 & w1288) | (~w925 & w15) | (w1288 & w15);
assign w128 = (w1650 & w662) | (w1650 & w1027) | (w662 & w1027);
assign w129 = (w350 & w661) | (w350 & w769) | (w661 & w769);
assign w130 = (~w854 & w419) | (~w854 & w1672) | (w419 & w1672);
assign w131 = (~w858 & w430) | (~w858 & w602) | (w430 & w602);
assign w132 = ~pi93 & ~pi94;
assign w133 = (w1491 & w1444) | (w1491 & w562) | (w1444 & w562);
assign w134 = ~w778 & ~pi68;
assign w135 = ~pi90 & ~pi91;
assign w136 = w157 & ~pi80;
assign w137 = (~pi83 & w105) | (~pi83 & w1890) | (w105 & w1890);
assign w138 = ~w1858 & ~w453;
assign w139 = ~w812 & pi77;
assign w140 = (~w1491 & w1233) | (~w1491 & w57) | (w1233 & w57);
assign w141 = w1858 & ~w814;
assign w142 = (~w1817 & w1384) | (~w1817 & w1112) | (w1384 & w1112);
assign w143 = w896 & w756;
assign w144 = w1147 & pi59;
assign w145 = ~w160 & ~w46;
assign w146 = (~w924 & w991) | (~w924 & w1000) | (w991 & w1000);
assign w147 = (w27 & w1883) | (w27 & w422) | (w1883 & w422);
assign w148 = ~w128 & ~w735;
assign w149 = (~w805 & w1854) | (~w805 & w452) | (w1854 & w452);
assign w150 = pi65 & w1557;
assign w151 = (~w665 & w794) | (~w665 & w1351) | (w794 & w1351);
assign w152 = (w1031 & w155) | (w1031 & w433) | (w155 & w433);
assign w153 = (w1773 & w1142) | (w1773 & w48) | (w1142 & w48);
assign w154 = ~w855 & w123;
assign w155 = ~pi62 & w796;
assign w156 = (pi77 & w399) | (pi77 & w1411) | (w399 & w1411);
assign w157 = ~w963 & ~w21;
assign w158 = ~w43 & w398;
assign w159 = (w1491 & w637) | (w1491 & w1604) | (w637 & w1604);
assign w160 = (pi29 & w487) | (pi29 & w2) | (w487 & w2);
assign w161 = (~w104 & w1378) | (~w104 & w1130) | (w1378 & w1130);
assign w162 = (w291 & w1159) | (w291 & w720) | (w1159 & w720);
assign w163 = pi90 & ~pi91;
assign w164 = w1931 & pi38;
assign w165 = (~w694 & w1631) | (~w694 & w1917) | (w1631 & w1917);
assign w166 = (~w325 & ~w915) | (~w325 & w504) | (~w915 & w504);
assign w167 = (w1351 & w454) | (w1351 & w233) | (w454 & w233);
assign w168 = ~w526 & ~w688;
assign w169 = w812 & w696;
assign w170 = w1259 & ~w89;
assign w171 = ~w334 & w1011;
assign w172 = (~w48 & w572) | (~w48 & w1609) | (w572 & w1609);
assign w173 = ~pi42 & ~pi43;
assign w174 = (~w1773 & w97) | (~w1773 & w1370) | (w97 & w1370);
assign w175 = (~w1773 & w745) | (~w1773 & w1887) | (w745 & w1887);
assign w176 = (pi62 & w931) | (pi62 & w1484) | (w931 & w1484);
assign w177 = w1066 & pi65;
assign w178 = (w549 & w774) | (w549 & ~w751) | (w774 & ~w751);
assign w179 = (w1715 & w362) | (w1715 & w1743) | (w362 & w1743);
assign w180 = (~w220 & w383) | (~w220 & w1090) | (w383 & w1090);
assign w181 = (pi59 & w648) | (pi59 & w674) | (w648 & w674);
assign w182 = w967 & ~w1347;
assign w183 = w1340 & ~pi03;
assign w184 = ~w1829 & w994;
assign w185 = ~w181 & ~w1548;
assign w186 = ~w761 & ~w390;
assign w187 = ~w292 & ~w1102;
assign w188 = w1640 & ~w658;
assign w189 = ~pi95 & w801;
assign w190 = ~w554 & w238;
assign w191 = (~w1310 & w1713) | (~w1310 & w870) | (w1713 & w870);
assign w192 = (w1584 & w1227) | (w1584 & w671) | (w1227 & w671);
assign w193 = ~w1011 & ~w547;
assign w194 = (w1142 & w1398) | (w1142 & w73) | (w1398 & w73);
assign w195 = ~w999 & ~w1158;
assign w196 = (w59 & w609) | (w59 & w189) | (w609 & w189);
assign w197 = w929 & w160;
assign w198 = (~w504 & w957) | (~w504 & w775) | (w957 & w775);
assign w199 = (~w743 & w517) | (~w743 & w1242) | (w517 & w1242);
assign w200 = ~w1160 & pi92;
assign w201 = pi65 & w1737;
assign w202 = ~w1589 & w1902;
assign w203 = (w1491 & w1739) | (w1491 & w1679) | (w1739 & w1679);
assign w204 = w1066 & w1737;
assign w205 = (~w958 & w777) | (~w958 & ~w1247) | (w777 & ~w1247);
assign w206 = ~w1074 & ~w1644;
assign w207 = ~w526 & ~w1755;
assign w208 = (w1138 & w1329) | (w1138 & w918) | (w1329 & w918);
assign w209 = (~w1715 & w1204) | (~w1715 & w198) | (w1204 & w198);
assign w210 = ~w1781 & ~w1217;
assign w211 = ~w1678 & ~pi41;
assign w212 = (w485 & w1607) | (w485 & w721) | (w1607 & w721);
assign w213 = (~w1533 & ~w658) | (~w1533 & ~w504) | (~w658 & ~w504);
assign w214 = ~pi84 & pi85;
assign w215 = ~w1881 & ~w1288;
assign w216 = ~w1616 & w1536;
assign w217 = (~w1491 & w236) | (~w1491 & w587) | (w236 & w587);
assign w218 = w1353 & w692;
assign w219 = w1318 & ~w1431;
assign w220 = (~w389 & w946) | (~w389 & w1274) | (w946 & w1274);
assign w221 = (w597 & w523) | (w597 & ~w1358) | (w523 & ~w1358);
assign w222 = ~w931 & w1349;
assign w223 = ~w1826 & w351;
assign w224 = (pi86 & w344) | (pi86 & w1896) | (w344 & w1896);
assign w225 = (w504 & w1821) | (w504 & w1910) | (w1821 & w1910);
assign w226 = ~w1480 & w731;
assign w227 = ~w365 & ~w354;
assign w228 = pi03 & pi04;
assign w229 = (w731 & w1624) | (w731 & w1480) | (w1624 & w1480);
assign w230 = (~pi41 & ~w896) | (~pi41 & w211) | (~w896 & w211);
assign w231 = pi42 & ~pi43;
assign w232 = (~w1199 & ~w739) | (~w1199 & w1900) | (~w739 & w1900);
assign w233 = ~w277 & ~w1077;
assign w234 = (w405 & w1434) | (w405 & w784) | (w1434 & w784);
assign w235 = ~w223 & ~w1356;
assign w236 = (w1515 & w598) | (w1515 & ~w1138) | (w598 & ~w1138);
assign w237 = ~w395 & ~w1493;
assign w238 = ~pi21 & ~pi22;
assign w239 = (w1773 & w726) | (w1773 & w473) | (w726 & w473);
assign w240 = (w1021 & w380) | (w1021 & w340) | (w380 & w340);
assign w241 = (w1491 & w1588) | (w1491 & w1267) | (w1588 & w1267);
assign w242 = ~w402 & w1390;
assign w243 = (w137 & w386) | (w137 & ~w1708) | (w386 & ~w1708);
assign w244 = ~w89 & ~w173;
assign w245 = (~w1817 & w1723) | (~w1817 & w1139) | (w1723 & w1139);
assign w246 = (~w389 & w466) | (~w389 & w1035) | (w466 & w1035);
assign w247 = (w146 & w67) | (w146 & w1527) | (w67 & w1527);
assign w248 = pi59 & ~w621;
assign w249 = ~w215 & ~w546;
assign w250 = (~pi29 & w1266) | (~pi29 & ~w1326) | (w1266 & ~w1326);
assign w251 = ~w109 & w318;
assign w252 = (~w694 & w1501) | (~w694 & w1180) | (w1501 & w1180);
assign w253 = ~w972 & w1466;
assign w254 = pi09 & pi10;
assign w255 = (~w1028 & w301) | (~w1028 & w1254) | (w301 & w1254);
assign w256 = (~w90 & w1098) | (~w90 & w423) | (w1098 & w423);
assign w257 = ~w733 & ~w498;
assign w258 = (w1540 & w107) | (w1540 & w1655) | (w107 & w1655);
assign w259 = (pi47 & ~w1575) | (pi47 & w125) | (~w1575 & w125);
assign w260 = ~pi50 & ~w982;
assign w261 = ~w319 & ~w297;
assign w262 = ~w1326 & ~w361;
assign w263 = (w128 & w1105) | (w128 & w1223) | (w1105 & w1223);
assign w264 = w1725 & ~w59;
assign w265 = (~w247 & w973) | (~w247 & w1145) | (w973 & w1145);
assign w266 = pi29 & ~w1332;
assign w267 = ~w1919 & ~w1106;
assign w268 = (w1201 & w1647) | (w1201 & w27) | (w1647 & w27);
assign w269 = w1693 & w1049;
assign w270 = (w1773 & w1398) | (w1773 & w73) | (w1398 & w73);
assign w271 = ~w1657 & w1733;
assign w272 = (~pi53 & ~w1) | (~pi53 & w1404) | (~w1 & w1404);
assign w273 = ~w1100 & ~w1553;
assign w274 = pi74 & w10;
assign w275 = ~w181 & w1792;
assign w276 = w838 & w943;
assign w277 = ~w1424 & ~w1018;
assign w278 = (~w1007 & ~w1387) | (~w1007 & ~w521) | (~w1387 & ~w521);
assign w279 = pi72 & ~pi73;
assign w280 = (w1501 & w1180) | (w1501 & ~w1849) | (w1180 & ~w1849);
assign w281 = ~w746 & w1851;
assign w282 = (~w1491 & w961) | (~w1491 & w964) | (w961 & w964);
assign w283 = pi95 & w801;
assign w284 = (w1412 & w109) | (w1412 & w717) | (w109 & w717);
assign w285 = (w27 & w661) | (w27 & w769) | (w661 & w769);
assign w286 = (~w1491 & w616) | (~w1491 & w79) | (w616 & w79);
assign w287 = pi71 & w1414;
assign w288 = ~pi86 & w1513;
assign w289 = (pi89 & ~w273) | (pi89 & w1348) | (~w273 & w1348);
assign w290 = pi57 & pi58;
assign w291 = (w389 & w1561) | (w389 & w998) | (w1561 & w998);
assign w292 = ~w1188 & ~w1481;
assign w293 = w840 & ~w1858;
assign w294 = ~w1768 & ~w305;
assign w295 = ~w1838 & ~w1757;
assign w296 = ~w1278 & ~w400;
assign w297 = (~pi41 & w508) | (~pi41 & w47) | (w508 & w47);
assign w298 = (w1575 & w693) | (w1575 & w1138) | (w693 & w1138);
assign w299 = (~pi71 & ~w1856) | (~pi71 & w1675) | (~w1856 & w1675);
assign w300 = (~w1708 & w386) | (~w1708 & w137) | (w386 & w137);
assign w301 = (~w1307 & w534) | (~w1307 & w852) | (w534 & w852);
assign w302 = (w1523 & w1126) | (w1523 & ~w498) | (w1126 & ~w498);
assign w303 = ~pi42 & pi43;
assign w304 = ~w1361 & ~w393;
assign w305 = (~w1665 & w1809) | (~w1665 & w1598) | (w1809 & w1598);
assign w306 = pi74 & ~w10;
assign w307 = (w1142 & w4) | (w1142 & w156) | (w4 & w156);
assign w308 = w1587 & ~w751;
assign w309 = ~pi80 & ~w413;
assign w310 = (~pi80 & w985) | (~pi80 & w654) | (w985 & w654);
assign w311 = (w1491 & w18) | (w1491 & w1597) | (w18 & w1597);
assign w312 = pi68 & w806;
assign w313 = ~w639 & w245;
assign w314 = (~pi92 & w1335) | (~pi92 & w1522) | (w1335 & w1522);
assign w315 = (w324 & w781) | (w324 & w803) | (w781 & w803);
assign w316 = (~w173 & w875) | (~w173 & w1704) | (w875 & w1704);
assign w317 = ~w594 & ~w508;
assign w318 = ~w992 & ~w1412;
assign w319 = pi41 & w317;
assign w320 = (~w220 & ~w1190) | (~w220 & ~w879) | (~w1190 & ~w879);
assign w321 = (w105 & w1465) | (w105 & w1128) | (w1465 & w1128);
assign w322 = (~w1817 & w1692) | (~w1817 & w1793) | (w1692 & w1793);
assign w323 = ~w1657 & w1359;
assign w324 = (~w1751 & w1355) | (~w1751 & w1243) | (w1355 & w1243);
assign w325 = (w591 & w522) | (w591 & w98) | (w522 & w98);
assign w326 = (w48 & w239) | (w48 & w917) | (w239 & w917);
assign w327 = (~w1033 & w1103) | (~w1033 & w510) | (w1103 & w510);
assign w328 = ~pi44 & w1916;
assign w329 = (w1682 & w30) | (w1682 & w378) | (w30 & w378);
assign w330 = ~w273 & pi89;
assign w331 = (w1751 & w1932) | (w1751 & w623) | (w1932 & w623);
assign w332 = w1694 & ~w444;
assign w333 = (w1142 & w300) | (w1142 & w950) | (w300 & w950);
assign w334 = (w388 & w1722) | (w388 & w1786) | (w1722 & w1786);
assign w335 = ~w403 & w451;
assign w336 = (w220 & w831) | (w220 & w617) | (w831 & w617);
assign w337 = w36 & pi20;
assign w338 = w1886 & pi74;
assign w339 = w1207 & pi35;
assign w340 = w1 & w668;
assign w341 = (w845 & w1063) | (w845 & w1773) | (w1063 & w1773);
assign w342 = (w887 & w825) | (w887 & w1600) | (w825 & w1600);
assign w343 = (pi71 & w916) | (pi71 & ~w1856) | (w916 & ~w1856);
assign w344 = ~w43 & ~w517;
assign w345 = ~w1354 & w1867;
assign w346 = w778 & ~pi68;
assign w347 = (~w1668 & w486) | (~w1668 & w694) | (w486 & w694);
assign w348 = (w414 & w1547) | (w414 & ~w694) | (w1547 & ~w694);
assign w349 = (w974 & w560) | (w974 & w1032) | (w560 & w1032);
assign w350 = (~w1594 & w1894) | (~w1594 & w371) | (w1894 & w371);
assign w351 = (w1540 & w535) | (w1540 & w884) | (w535 & w884);
assign w352 = ~w951 & w953;
assign w353 = w1106 & ~w1345;
assign w354 = (~w1885 & w1753) | (~w1885 & w24) | (w1753 & w24);
assign w355 = (~w1491 & w1116) | (~w1491 & w1084) | (w1116 & w1084);
assign w356 = (w997 & w1681) | (w997 & w1505) | (w1681 & w1505);
assign w357 = ~w1469 & ~w1286;
assign w358 = (w1817 & w813) | (w1817 & w1346) | (w813 & w1346);
assign w359 = (~w576 & w989) | (~w576 & w1873) | (w989 & w1873);
assign w360 = w135 & ~w805;
assign w361 = ~pi27 & ~pi28;
assign w362 = (w1653 & w1245) | (w1653 & w1935) | (w1245 & w1935);
assign w363 = (~w1596 & w263) | (~w1596 & w1761) | (w263 & w1761);
assign w364 = ~w1750 & ~pi89;
assign w365 = ~w111 & ~w1583;
assign w366 = ~pi18 & ~pi19;
assign w367 = (~w896 & w1436) | (~w896 & w1937) | (w1436 & w1937);
assign w368 = (~w971 & w673) | (~w971 & w584) | (w673 & w584);
assign w369 = (w1386 & w260) | (w1386 & ~w1138) | (w260 & ~w1138);
assign w370 = w1450 & ~w304;
assign w371 = w910 & ~w1594;
assign w372 = (w1078 & w560) | (w1078 & w1032) | (w560 & w1032);
assign w373 = (w52 & w1664) | (w52 & w322) | (w1664 & w322);
assign w374 = w687 & ~w1254;
assign w375 = (~w439 & w182) | (~w439 & w1807) | (w182 & w1807);
assign w376 = ~w1199 & ~w983;
assign w377 = ~w808 & ~w1605;
assign w378 = (~w105 & w548) | (~w105 & w1760) | (w548 & w1760);
assign w379 = ~w376 & w663;
assign w380 = w1 & pi53;
assign w381 = ~w251 & ~w284;
assign w382 = ~pi38 & ~w644;
assign w383 = (w1744 & w823) | (w1744 & ~w521) | (w823 & ~w521);
assign w384 = ~w1275 & ~w1121;
assign w385 = (pi44 & w1050) | (pi44 & w1311) | (w1050 & w1311);
assign w386 = w105 & ~pi83;
assign w387 = (w1462 & w330) | (w1462 & w1208) | (w330 & w1208);
assign w388 = (w1878 & w1442) | (w1878 & w1740) | (w1442 & w1740);
assign w389 = (~w255 & w618) | (~w255 & w1875) | (w618 & w1875);
assign w390 = (w1179 & w689) | (w1179 & w927) | (w689 & w927);
assign w391 = ~w731 & pi29;
assign w392 = ~w896 & ~pi41;
assign w393 = (~pi50 & w403) | (~pi50 & w1022) | (w403 & w1022);
assign w394 = w1552 & ~pi50;
assign w395 = (w997 & w1503) | (w997 & w1658) | (w1503 & w1658);
assign w396 = (w1142 & w321) | (w1142 & w776) | (w321 & w776);
assign w397 = w1221 & ~w16;
assign w398 = pi81 & pi82;
assign w399 = w1236 & ~w812;
assign w400 = (~w997 & w793) | (~w997 & w161) | (w793 & w161);
assign w401 = w1305 & ~w737;
assign w402 = (~w1363 & w1828) | (~w1363 & w126) | (w1828 & w126);
assign w403 = (~w1491 & w1580) | (~w1491 & w695) | (w1580 & w695);
assign w404 = ~w787 & w287;
assign w405 = (pi74 & w402) | (pi74 & w1153) | (w402 & w1153);
assign w406 = w532 & ~w1584;
assign w407 = (w232 & w376) | (w232 & ~w1167) | (w376 & ~w1167);
assign w408 = ~w1510 & ~w1589;
assign w409 = (w1304 & w1392) | (w1304 & ~w247) | (w1392 & ~w247);
assign w410 = pi39 & pi40;
assign w411 = ~w42 & ~w1634;
assign w412 = pi41 & w896;
assign w413 = ~w157 & ~w202;
assign w414 = (~w1584 & w873) | (~w1584 & w912) | (w873 & w912);
assign w415 = (~pi80 & w1296) | (~pi80 & w136) | (w1296 & w136);
assign w416 = (~w145 & w1825) | (~w145 & w281) | (w1825 & w281);
assign w417 = ~w377 & ~w1167;
assign w418 = ~w336 & ~w1291;
assign w419 = w1548 & ~w869;
assign w420 = (w960 & w833) | (w960 & ~w521) | (w833 & ~w521);
assign w421 = (~w1470 & w1528) | (~w1470 & w640) | (w1528 & w640);
assign w422 = w1856 & w1646;
assign w423 = w857 & ~w90;
assign w424 = ~w443 & w134;
assign w425 = (w1684 & w897) | (w1684 & w971) | (w897 & w971);
assign w426 = (~w1491 & w1477) | (~w1491 & w1252) | (w1477 & w1252);
assign w427 = (~w247 & w851) | (~w247 & w272) | (w851 & w272);
assign w428 = w1656 & pi56;
assign w429 = (w1002 & w1173) | (w1002 & w971) | (w1173 & w971);
assign w430 = ~w534 & w900;
assign w431 = ~w1576 & w75;
assign w432 = w1093 & w746;
assign w433 = (w971 & w1380) | (w971 & w247) | (w1380 & w247);
assign w434 = ~w1928 & ~w1450;
assign w435 = ~w173 & ~pi47;
assign w436 = (w576 & w1905) | (w576 & w1520) | (w1905 & w1520);
assign w437 = w1737 & w177;
assign w438 = (w909 & w14) | (w909 & w1021) | (w14 & w1021);
assign w439 = (w842 & w1885) | (w842 & w751) | (w1885 & w751);
assign w440 = ~w985 & w1040;
assign w441 = (~w576 & w1770) | (~w576 & w1717) | (w1770 & w1717);
assign w442 = ~pi32 & w1231;
assign w443 = ~w910 & ~w1894;
assign w444 = ~w90 & ~w1678;
assign w445 = pi38 & ~w644;
assign w446 = (~pi89 & ~w273) | (~pi89 & w364) | (~w273 & w364);
assign w447 = (~w1021 & w851) | (~w1021 & w272) | (w851 & w272);
assign w448 = ~w334 & w547;
assign w449 = (~w1682 & w1776) | (~w1682 & w1194) | (w1776 & w1194);
assign w450 = ~w854 & ~w1919;
assign w451 = (~w1491 & w369) | (~w1491 & w1903) | (w369 & w1903);
assign w452 = w1553 & ~w805;
assign w453 = ~pi69 & ~pi70;
assign w454 = ~w277 & ~w1799;
assign w455 = ~w453 & w814;
assign w456 = (w1142 & w1260) | (w1142 & w1601) | (w1260 & w1601);
assign w457 = (w1122 & w1562) | (w1122 & w576) | (w1562 & w576);
assign w458 = (w175 & w542) | (w175 & ~w48) | (w542 & ~w48);
assign w459 = (~w1591 & w373) | (~w1591 & w1226) | (w373 & w1226);
assign w460 = (w1514 & w1797) | (w1514 & w1720) | (w1797 & w1720);
assign w461 = w262 & ~w865;
assign w462 = (w1529 & w979) | (w1529 & w1560) | (w979 & w1560);
assign w463 = (w48 & w1089) | (w48 & w456) | (w1089 & w456);
assign w464 = (w576 & w59) | (w576 & w48) | (w59 & w48);
assign w465 = ~w1162 & w827;
assign w466 = (~w1923 & ~w1229) | (~w1923 & w1274) | (~w1229 & w1274);
assign w467 = (~w325 & ~w915) | (~w325 & w1618) | (~w915 & w1618);
assign w468 = w1339 & ~w1358;
assign w469 = (w151 & w559) | (w151 & w1849) | (w559 & w1849);
assign w470 = w36 & ~pi20;
assign w471 = (w504 & w1067) | (w504 & w613) | (w1067 & w613);
assign w472 = (w530 & w1525) | (w530 & w102) | (w1525 & w102);
assign w473 = (w1214 & w1842) | (w1214 & w16) | (w1842 & w16);
assign w474 = pi45 & pi46;
assign w475 = w1585 & ~w1915;
assign w476 = (w1443 & ~w758) | (w1443 & ~w1431) | (~w758 & ~w1431);
assign w477 = ~w914 & ~w692;
assign w478 = ~w90 & ~w1674;
assign w479 = (pi89 & w1909) | (pi89 & w1879) | (w1909 & w1879);
assign w480 = (~pi56 & w1576) | (~pi56 & w760) | (w1576 & w760);
assign w481 = (w549 & w774) | (w549 & ~w1351) | (w774 & ~w1351);
assign w482 = w157 & pi80;
assign w483 = w992 & ~pi11;
assign w484 = (w1438 & w725) | (w1438 & w86) | (w725 & w86);
assign w485 = ~w1836 & w763;
assign w486 = w1011 & ~w1668;
assign w487 = (~w1540 & w229) | (~w1540 & w1332) | (w229 & w1332);
assign w488 = (~w1358 & w1312) | (~w1358 & w585) | (w1312 & w585);
assign w489 = (w1740 & w898) | (w1740 & w1680) | (w898 & w1680);
assign w490 = (~w52 & w358) | (~w52 & w988) | (w358 & w988);
assign w491 = (~w450 & w1319) | (~w450 & w1640) | (w1319 & w1640);
assign w492 = (w1209 & w382) | (w1209 & ~w1410) | (w382 & ~w1410);
assign w493 = (~w1618 & w1819) | (~w1618 & w188) | (w1819 & w188);
assign w494 = w934 & w1163;
assign w495 = (w574 & w895) | (w574 & w1400) | (w895 & w1400);
assign w496 = ~w173 & ~w1132;
assign w497 = w814 & ~w1510;
assign w498 = (~w1616 & ~w1103) | (~w1616 & w862) | (~w1103 & w862);
assign w499 = (~w1138 & w1046) | (~w1138 & w699) | (w1046 & w699);
assign w500 = (w1163 & w150) | (w1163 & w494) | (w150 & w494);
assign w501 = pi78 & pi79;
assign w502 = (~w1491 & w889) | (~w1491 & w1483) | (w889 & w1483);
assign w503 = ~w1746 & ~w524;
assign w504 = (w1053 & w1653) | (w1053 & w1387) | (w1653 & w1387);
assign w505 = ~w805 & ~w135;
assign w506 = (~w59 & w989) | (~w59 & w1873) | (w989 & w1873);
assign w507 = pi18 & pi19;
assign w508 = (w682 & w570) | (w682 & w367) | (w570 & w367);
assign w509 = ~w855 & w1210;
assign w510 = w1616 & ~w1033;
assign w511 = w1500 & pi83;
assign w512 = (w123 & w855) | (w123 & w716) | (w855 & w716);
assign w513 = (w389 & w1904) | (w389 & w1137) | (w1904 & w1137);
assign w514 = ~w1656 & ~pi56;
assign w515 = pi83 & ~w396;
assign w516 = (pi74 & w1273) | (pi74 & w338) | (w1273 & w338);
assign w517 = w1500 & ~w398;
assign w518 = (w597 & w523) | (w597 & ~w48) | (w523 & ~w48);
assign w519 = ~w534 & ~w680;
assign w520 = (w1036 & w274) | (w1036 & w350) | (w274 & w350);
assign w521 = (w295 & w1175) | (w295 & w1431) | (w1175 & w1431);
assign w522 = ~w419 | w869;
assign w523 = pi68 & ~w806;
assign w524 = (~w997 & w348) | (~w997 & w1425) | (w348 & w1425);
assign w525 = ~w1820 & w1154;
assign w526 = ~w508 & w1545;
assign w527 = (w576 & w1490) | (w576 & w479) | (w1490 & w479);
assign w528 = ~pi24 & pi25;
assign w529 = ~w41 & pi32;
assign w530 = (w295 & w1175) | (w295 & w1549) | (w1175 & w1549);
assign w531 = w1749 & ~w1533;
assign w532 = ~w390 & ~w148;
assign w533 = ~w685 & ~w600;
assign w534 = (~w1393 & w1869) | (~w1393 & w1422) | (w1869 & w1422);
assign w535 = (w1712 & w445) | (w1712 & ~w1410) | (w445 & ~w1410);
assign w536 = (w1715 & w710) | (w1715 & w187) | (w710 & w187);
assign w537 = ~w1851 | w1083;
assign w538 = (w1007 & w1387) | (w1007 & w530) | (w1387 & w530);
assign w539 = (~w1354 & w913) | (~w1354 & w1519) | (w913 & w1519);
assign w540 = (w1125 & w1016) | (w1125 & ~w683) | (w1016 & ~w683);
assign w541 = ~w1236 & pi77;
assign w542 = (~w1142 & w745) | (~w1142 & w1887) | (w745 & w1887);
assign w543 = ~w882 & ~w792;
assign w544 = pi92 & ~w722;
assign w545 = (~w1726 & w1324) | (~w1726 & w1550) | (w1324 & w1550);
assign w546 = (~w547 & ~w1011) | (~w547 & w925) | (~w1011 & w925);
assign w547 = ~w402 & w1730;
assign w548 = w501 & ~w105;
assign w549 = (~w186 & w1847) | (~w186 & w1429) | (w1847 & w1429);
assign w550 = ~pi04 & pi05;
assign w551 = w69 & ~w1198;
assign w552 = ~pi54 & pi55;
assign w553 = w1319 & ~w450;
assign w554 = ~w528 & ~w1846;
assign w555 = (w424 & w1327) | (w424 & w1358) | (w1327 & w1358);
assign w556 = ~w303 & ~w231;
assign w557 = w398 & ~w1750;
assign w558 = w1657 & w1396;
assign w559 = (~w665 & w794) | (~w665 & w751) | (w794 & w751);
assign w560 = (pi86 & ~w1726) | (pi86 & w1637) | (~w1726 & w1637);
assign w561 = (~w244 & w1129) | (~w244 & w1704) | (w1129 & w1704);
assign w562 = (pi47 & w1889) | (pi47 & w1300) | (w1889 & w1300);
assign w563 = ~w1096 & ~w162;
assign w564 = (w1491 & w328) | (w1491 & w1224) | (w328 & w1224);
assign w565 = (~w273 & w1909) | (~w273 & w1081) | (w1909 & w1081);
assign w566 = (~pi68 & w981) | (~pi68 & w1471) | (w981 & w1471);
assign w567 = w486 & ~w1668;
assign w568 = ~w1005 & w1023;
assign w569 = ~w1354 & w1412;
assign w570 = (~w896 & w1436) | (~w896 & ~w1678) | (w1436 & ~w1678);
assign w571 = (~w1668 & w486) | (~w1668 & ~w1310) | (w486 & ~w1310);
assign w572 = (~w27 & w940) | (~w27 & w299) | (w940 & w299);
assign w573 = (w352 & w1918) | (w352 & w1527) | (w1918 & w1527);
assign w574 = (w48 & w1620) | (w48 & w1295) | (w1620 & w1295);
assign w575 = w635 & ~pi08;
assign w576 = (w1773 & w615) | (w1773 & w1313) | (w615 & w1313);
assign w577 = (~w1491 & w1152) | (~w1491 & w966) | (w1152 & w966);
assign w578 = (w1700 & w1279) | (w1700 & ~w1142) | (w1279 & ~w1142);
assign w579 = (pi92 & w1298) | (pi92 & w1004) | (w1298 & w1004);
assign w580 = ~w1754 & ~w822;
assign w581 = (w1358 & w1089) | (w1358 & w456) | (w1089 & w456);
assign w582 = (w137 & w386) | (w137 & ~w22) | (w386 & ~w22);
assign w583 = (~pi26 & w986) | (~pi26 & w1435) | (w986 & w1435);
assign w584 = (~pi59 & ~w1684) | (~pi59 & w859) | (~w1684 & w859);
assign w585 = (~pi65 & ~w1737) | (~pi65 & w868) | (~w1737 & w868);
assign w586 = (w1287 & w232) | (w1287 & w955) | (w232 & w955);
assign w587 = (w1515 & w598) | (w1515 & ~w1527) | (w598 & ~w1527);
assign w588 = (w1064 & w1388) | (w1064 & w1413) | (w1388 & w1413);
assign w589 = ~w1033 & ~w1536;
assign w590 = (w481 & w178) | (w481 & ~w694) | (w178 & ~w694);
assign w591 = (~w431 & ~w1792) | (~w431 & w646) | (~w1792 & w646);
assign w592 = (w1491 & w1759) | (w1491 & w678) | (w1759 & w678);
assign w593 = w1552 & pi50;
assign w594 = (w896 & w1491) | (w896 & w1812) | (w1491 & w1812);
assign w595 = (~w1286 & w109) | (~w1286 & w1203) | (w109 & w1203);
assign w596 = (w1927 & w990) | (w1927 & w48) | (w990 & w48);
assign w597 = (pi68 & w443) | (pi68 & w906) | (w443 & w906);
assign w598 = pi50 & ~w982;
assign w599 = (w1633 & w1420) | (w1633 & ~w1021) | (w1420 & ~w1021);
assign w600 = (~w608 & w704) | (~w608 & w1472) | (w704 & w1472);
assign w601 = (~w1412 & w655) | (~w1412 & w558) | (w655 & w558);
assign w602 = (w1307 & w1028) | (w1307 & w63) | (w1028 & w63);
assign w603 = (w754 & w1381) | (w754 & ~w1078) | (w1381 & ~w1078);
assign w604 = (w59 & w314) | (w59 & w70) | (w314 & w70);
assign w605 = (w576 & w289) | (w576 & w1366) | (w289 & w1366);
assign w606 = (~pi95 & w1140) | (~pi95 & w149) | (w1140 & w149);
assign w607 = w207 & ~w530;
assign w608 = ~w1592 & ~w1732;
assign w609 = ~pi95 & w512;
assign w610 = ~w737 & ~w1066;
assign w611 = (~w888 & ~w50) | (~w888 & ~w48) | (~w50 & ~w48);
assign w612 = (pi95 & w1467) | (pi95 & w716) | (w1467 & w716);
assign w613 = (~w1794 & w1117) | (~w1794 & w658) | (w1117 & w658);
assign w614 = (w788 & w1785) | (w788 & ~w350) | (w1785 & ~w350);
assign w615 = (w199 & w773) | (w199 & w1128) | (w773 & w1128);
assign w616 = (~w1575 & w1889) | (~w1575 & w1385) | (w1889 & w1385);
assign w617 = (~w1006 & w1806) | (~w1006 & w530) | (w1806 & w530);
assign w618 = ~w1377 & w1198;
assign w619 = w1771 & ~w1360;
assign w620 = (w1817 & w77) | (w1817 & w826) | (w77 & w826);
assign w621 = (w1021 & w425) | (w1021 & w1913) | (w425 & w1913);
assign w622 = (w1276 & w110) | (w1276 & ~w1358) | (w110 & ~w1358);
assign w623 = ~w376 & w1334;
assign w624 = ~w405 & ~w547;
assign w625 = ~w1552 & ~pi50;
assign w626 = ~w1382 & w1083;
assign w627 = ~w1622 & pi17;
assign w628 = ~pi14 & ~w580;
assign w629 = ~w556 & pi44;
assign w630 = ~w501 & ~w1500;
assign w631 = (~w59 & w886) | (~w59 & w446) | (w886 & w446);
assign w632 = ~w893 & ~w1382;
assign w633 = ~w1621 & ~w1685;
assign w634 = ~w867 & w697;
assign w635 = pi00 & pi01;
assign w636 = (~w1885 & w902) | (~w1885 & w1787) | (w902 & w1787);
assign w637 = (w1021 & w1051) | (w1021 & w1403) | (w1051 & w1403);
assign w638 = ~w1345 & ~w540;
assign w639 = (~w1817 & w976) | (~w1817 & w1745) | (w976 & w1745);
assign w640 = w812 & w139;
assign w641 = w847 & ~w692;
assign w642 = (w1731 & w1628) | (w1731 & w1462) | (w1628 & w1462);
assign w643 = pi04 & ~pi05;
assign w644 = ~w1931 & ~w1674;
assign w645 = (w1817 & w1871) | (w1817 & w1511) | (w1871 & w1511);
assign w646 = ~w431 & w1320;
assign w647 = (w1817 & w604) | (w1817 & w1202) | (w604 & w1202);
assign w648 = (~w1491 & w1426) | (~w1491 & w1859) | (w1426 & w1859);
assign w649 = (w220 & w1265) | (w220 & w1565) | (w1265 & w1565);
assign w650 = ~w1539 & pi86;
assign w651 = (w48 & w1563) | (w48 & w307) | (w1563 & w307);
assign w652 = ~w1160 & ~pi92;
assign w653 = ~w1535 & ~w1936;
assign w654 = (w1491 & w1615) | (w1491 & w1627) | (w1615 & w1627);
assign w655 = ~w1781 & ~w1649;
assign w656 = w1858 & pi71;
assign w657 = (pi68 & w867) | (pi68 & w116) | (w867 & w116);
assign w658 = ~w181 & ~w646;
assign w659 = (~w1540 & w1758) | (~w1540 & w1486) | (w1758 & w1486);
assign w660 = (~w232 & w1266) | (~w232 & w250) | (w1266 & w250);
assign w661 = w1856 & pi71;
assign w662 = (w1817 & w372) | (w1817 & w349) | (w372 & w349);
assign w663 = ~w894 & ~pi26;
assign w664 = ~w1135 & pi29;
assign w665 = ~w1629 & ~w310;
assign w666 = (w222 & w1735) | (w222 & w1651) | (w1735 & w1651);
assign w667 = (w59 & w1780) | (w59 & w1691) | (w1780 & w1691);
assign w668 = w809 & pi53;
assign w669 = (~w505 & w1335) | (~w505 & w1725) | (w1335 & w1725);
assign w670 = (~w1817 & w1149) | (~w1817 & w1625) | (w1149 & w1625);
assign w671 = (~w1542 & w762) | (~w1542 & w1237) | (w762 & w1237);
assign w672 = w138 & ~w27;
assign w673 = ~w1684 & ~pi59;
assign w674 = (w1491 & w1763) | (w1491 & w1857) | (w1763 & w1857);
assign w675 = (w192 & w1827) | (w192 & w694) | (w1827 & w694);
assign w676 = pi44 & w1916;
assign w677 = (~pi08 & ~w1686) | (~pi08 & w795) | (~w1686 & w795);
assign w678 = (w974 & w1078) | (w974 & w48) | (w1078 & w48);
assign w679 = (~w52 & w1086) | (~w52 & w620) | (w1086 & w620);
assign w680 = ~pi11 & ~w381;
assign w681 = (pi11 & w109) | (pi11 & w94) | (w109 & w94);
assign w682 = (w1540 & w748) | (w1540 & w1863) | (w748 & w1863);
assign w683 = (w1185 & w130) | (w1185 & w658) | (w130 & w658);
assign w684 = (w1773 & w321) | (w1773 & w776) | (w321 & w776);
assign w685 = ~w968 & ~w1239;
assign w686 = (w714 & w333) | (w714 & w1358) | (w333 & w1358);
assign w687 = ~w69 & ~w1377;
assign w688 = ~w764 & w426;
assign w689 = (w1491 & w686) | (w1491 & w947) | (w686 & w947);
assign w690 = w1476 & ~w694;
assign w691 = (w1751 & w1235) | (w1751 & w767) | (w1235 & w767);
assign w692 = (pi35 & w928) | (pi35 & w659) | (w928 & w659);
assign w693 = w173 & w1575;
assign w694 = (w1636 & w191) | (w1636 & w1666) | (w191 & w1666);
assign w695 = (~w1464 & w977) | (~w1464 & w1069) | (w977 & w1069);
assign w696 = w1510 & ~pi77;
assign w697 = (~w1491 & w221) | (~w1491 & w518) | (w221 & w518);
assign w698 = (~w1491 & w1488) | (~w1491 & w1161) | (w1488 & w1161);
assign w699 = (~pi47 & ~w1575) | (~pi47 & w435) | (~w1575 & w435);
assign w700 = (w960 & w833) | (w960 & ~w530) | (w833 & ~w530);
assign w701 = (w576 & w1502) | (w576 & w612) | (w1502 & w612);
assign w702 = w1639 & ~pi23;
assign w703 = w373 & w1718;
assign w704 = (pi03 & w1238) | (pi03 & w1521) | (w1238 & w1521);
assign w705 = (~w1540 & w1507) | (~w1540 & w711) | (w1507 & w711);
assign w706 = (w1021 & w1258) | (w1021 & w1784) | (w1258 & w1784);
assign w707 = (w59 & w289) | (w59 & w1366) | (w289 & w1366);
assign w708 = ~w1594 & ~w1858;
assign w709 = w1199 & ~w238;
assign w710 = (w1007 & w1368) | (w1007 & w785) | (w1368 & w785);
assign w711 = (w1277 & w1494) | (w1277 & w865) | (w1494 & w865);
assign w712 = (~w1540 & w1282) | (~w1540 & w1677) | (w1282 & w1677);
assign w713 = (~w911 & w1338) | (~w911 & w1387) | (w1338 & w1387);
assign w714 = (w1773 & w243) | (w1773 & w582) | (w243 & w582);
assign w715 = (w1036 & w274) | (w1036 & w27) | (w274 & w27);
assign w716 = ~w805 & ~w1322;
assign w717 = w992 & w1412;
assign w718 = w632 & ~w618;
assign w719 = w839 & ~w1147;
assign w720 = (~w100 & w1506) | (~w100 & w849) | (w1506 & w849);
assign w721 = (w1347 & w1237) | (w1347 & w1584) | (w1237 & w1584);
assign w722 = ~w1160 & ~w1322;
assign w723 = (~w1326 & w983) | (~w1326 & w6) | (w983 & w6);
assign w724 = (~w1803 & w1670) | (~w1803 & w407) | (w1670 & w407);
assign w725 = (pi77 & w812) | (pi77 & w541) | (w812 & w541);
assign w726 = (w1214 & w1842) | (w1214 & w1128) | (w1842 & w1128);
assign w727 = ~w869 & ~w1163;
assign w728 = (w461 & w114) | (w461 & w1172) | (w114 & w1172);
assign w729 = ~w228 & ~w635;
assign w730 = ~w1195 & ~w1875;
assign w731 = ~w1585 & ~w361;
assign w732 = w1684 & w1369;
assign w733 = ~w507 & ~w366;
assign w734 = (~w304 & w370) | (~w304 & w1007) | (w370 & w1007);
assign w735 = ~w639 & w1271;
assign w736 = w1656 & ~pi56;
assign w737 = pi60 & pi61;
assign w738 = (w1002 & w1173) | (w1002 & w1380) | (w1173 & w1380);
assign w739 = w507 & ~w366;
assign w740 = (~w220 & w1076) | (~w220 & w219) | (w1076 & w219);
assign w741 = ~w1792 & ~w431;
assign w742 = ~w465 & ~w1800;
assign w743 = pi84 & pi85;
assign w744 = ~w782 & w335;
assign w745 = w1550 & ~w1128;
assign w746 = ~w986 & w1371;
assign w747 = (~pi74 & w402) | (~pi74 & w1893) | (w402 & w1893);
assign w748 = w1752 & ~w1410;
assign w749 = (w222 & w1735) | (w222 & w433) | (w1735 & w433);
assign w750 = (w1700 & w1279) | (w1700 & ~w1773) | (w1279 & ~w1773);
assign w751 = ~w334 & ~w925;
assign w752 = w254 & ~w1536;
assign w753 = (w175 & w542) | (w175 & ~w1358) | (w542 & ~w1358);
assign w754 = (~pi86 & w344) | (~pi86 & w1024) | (w344 & w1024);
assign w755 = w384 & ~pi62;
assign w756 = w1678 & pi41;
assign w757 = ~w712 & w1430;
assign w758 = w914 & ~w1443;
assign w759 = (~w261 & w1146) | (~w261 & ~w476) | (w1146 & ~w476);
assign w760 = (w1491 & w828) | (w1491 & w834) | (w828 & w834);
assign w761 = (pi83 & w1775) | (pi83 & w861) | (w1775 & w861);
assign w762 = w1105 & ~w1542;
assign w763 = w1718 | ~w1591;
assign w764 = (~w1491 & w1676) | (~w1491 & w561) | (w1676 & w561);
assign w765 = (w974 & w1813) | (w974 & w1574) | (w1813 & w1574);
assign w766 = ~w649 & ~w740;
assign w767 = ~w731 & w660;
assign w768 = (w1479 & w872) | (w1479 & w9) | (w872 & w9);
assign w769 = w1856 & w656;
assign w770 = pi95 & ~w512;
assign w771 = (~w1263 & w500) | (~w1263 & w467) | (w500 & w467);
assign w772 = ~w764 & w1898;
assign w773 = ~w743 & ~w158;
assign w774 = w1847 & ~w186;
assign w775 = (~w185 & w1719) | (~w185 & w741) | (w1719 & w741);
assign w776 = (w105 & w1465) | (w105 & w16) | (w1465 & w16);
assign w777 = w1919 & ~w958;
assign w778 = ~w1924 & ~w1357;
assign w779 = ~w1061 & ~w891;
assign w780 = w731 & ~pi29;
assign w781 = (w1540 & w266) | (w1540 & w933) | (w266 & w933);
assign w782 = (pi53 & w1814) | (pi53 & w1577) | (w1814 & w1577);
assign w783 = w1906 & ~w1142;
assign w784 = w334 & w405;
assign w785 = ~w292 & ~w1177;
assign w786 = ~w1826 & w1497;
assign w787 = (w1643 & w124) | (w1643 & w1663) | (w124 & w1663);
assign w788 = (~pi74 & w1273) | (~pi74 & w85) | (w1273 & w85);
assign w789 = (~pi86 & w639) | (~pi86 & w1914) | (w639 & w1914);
assign w790 = (w59 & w1490) | (w59 & w479) | (w1490 & w479);
assign w791 = w1860 & ~w1471;
assign w792 = ~pi03 & pi04;
assign w793 = (~w104 & w1378) | (~w104 & w1774) | (w1378 & w1774);
assign w794 = (w1434 & w1629) | (w1434 & w892) | (w1629 & w892);
assign w795 = ~w543 & w575;
assign w796 = ~w384 & ~w1645;
assign w797 = (w1715 & w1512) | (w1715 & w471) | (w1512 & w471);
assign w798 = ~w96 & ~w890;
assign w799 = (~w1851 & w1083) | (~w1851 & ~w618) | (w1083 & ~w618);
assign w800 = (~w1817 & w1234) | (~w1817 & w515) | (w1234 & w515);
assign w801 = (w123 & w855) | (w123 & w149) | (w855 & w149);
assign w802 = (~pi03 & w1611) | (~pi03 & w84) | (w1611 & w84);
assign w803 = (w1540 & w1449) | (w1540 & w901) | (w1449 & w901);
assign w804 = (~pi77 & ~w812) | (~pi77 & w71) | (~w812 & w71);
assign w805 = pi90 & pi91;
assign w806 = ~w778 & ~w1573;
assign w807 = (~w366 & w739) | (~w366 & w1167) | (w739 & w1167);
assign w808 = ~pi18 & pi19;
assign w809 = ~pi48 & ~pi49;
assign w810 = (w1491 & w1308) | (w1491 & w596) | (w1308 & w596);
assign w811 = (w1476 & w540) | (w1476 & w1094) | (w540 & w1094);
assign w812 = ~w1902 & ~w1589;
assign w813 = (w576 & w606) | (w576 & w1659) | (w606 & w1659);
assign w814 = pi69 & pi70;
assign w815 = w262 & ~w1480;
assign w816 = w877 & pi03;
assign w817 = ~w286 & w698;
assign w818 = pi48 & ~pi49;
assign w819 = (~w1 & w1251) | (~w1 & ~w809) | (w1251 & ~w809);
assign w820 = pi51 & pi52;
assign w821 = (w1845 & w269) | (w1845 & ~w1606) | (w269 & ~w1606);
assign w822 = (~w0 & w595) | (~w0 & w1041) | (w595 & w1041);
assign w823 = w34 & ~w434;
assign w824 = ~pi77 & w812;
assign w825 = w1207 & ~pi35;
assign w826 = (w59 & w1683) | (w59 & w283) | (w1683 & w283);
assign w827 = ~w36 & pi20;
assign w828 = (w866 & w1832) | (w866 & w1021) | (w1832 & w1021);
assign w829 = ~w1408 & ~w131;
assign w830 = w786 & ~w1838;
assign w831 = (~w1006 & w1806) | (~w1006 & w521) | (w1806 & w521);
assign w832 = ~w1309 & ~w335;
assign w833 = w1143 & ~w1007;
assign w834 = (w866 & w1832) | (w866 & w247) | (w1832 & w247);
assign w835 = w820 & ~w1926;
assign w836 = w812 & w1654;
assign w837 = w786 & ~w914;
assign w838 = ~w228 & ~w1593;
assign w839 = w820 & ~w1147;
assign w840 = w1901 & ~w1858;
assign w841 = pi86 & ~w1726;
assign w842 = ~w761 & ~w1799;
assign w843 = w496 & ~w1138;
assign w844 = (w504 & w1666) | (w504 & w683) | (w1666 & w683);
assign w845 = ~w1296 & w1516;
assign w846 = w1686 & w1619;
assign w847 = ~w51 & w258;
assign w848 = (w247 & w1258) | (w247 & w1784) | (w1258 & w1784);
assign w849 = ~w914 & ~w786;
assign w850 = (w1491 & w412) | (w1491 & w143) | (w412 & w143);
assign w851 = ~w1 & ~pi53;
assign w852 = w680 & ~w1307;
assign w853 = ~w757 & ~w1211;
assign w854 = (pi65 & w1474) | (pi65 & w203) | (w1474 & w203);
assign w855 = w135 & w123;
assign w856 = ~w949 & ~w1389;
assign w857 = ~pi33 & ~pi34;
assign w858 = ~w1028 & ~w69;
assign w859 = ~w1147 & ~pi59;
assign w860 = w453 & ~w1236;
assign w861 = (w1491 & w5) | (w1491 & w326) | (w5 & w326);
assign w862 = w1033 & ~w1616;
assign w863 = ~pi05 & ~w276;
assign w864 = ~w733 & ~w1925;
assign w865 = ~w1135 & ~w709;
assign w866 = ~w1092 & w514;
assign w867 = (~w708 & w1471) | (~w708 & w1643) | (w1471 & w1643);
assign w868 = ~w1066 & ~pi65;
assign w869 = (pi62 & w948) | (pi62 & w1728) | (w948 & w1728);
assign w870 = w1106 & ~w1310;
assign w871 = ~w232 & w663;
assign w872 = (~w1737 & w1508) | (~w1737 & ~w1066) | (w1508 & ~w1066);
assign w873 = w263 & ~w1596;
assign w874 = (~w1540 & w956) | (~w1540 & w54) | (w956 & w54);
assign w875 = w410 & ~w173;
assign w876 = pi86 & w1513;
assign w877 = pi01 & pi02;
assign w878 = ~pi00 & ~pi01;
assign w879 = (w1618 & w504) | (w1618 & w530) | (w504 & w530);
assign w880 = ~pi90 & pi91;
assign w881 = w1678 & ~w410;
assign w882 = pi03 & ~pi04;
assign w883 = ~pi30 & pi31;
assign w884 = (w1712 & w445) | (w1712 & ~w1600) | (w445 & ~w1600);
assign w885 = ~w1656 & pi56;
assign w886 = ~w273 & ~pi89;
assign w887 = w1207 & w1880;
assign w888 = (w1856 & w1447) | (w1856 & w27) | (w1447 & w27);
assign w889 = (w1546 & w1769) | (w1546 & ~w433) | (w1769 & ~w433);
assign w890 = (~w1715 & w1419) | (~w1715 & w1253) | (w1419 & w1253);
assign w891 = (~w936 & w821) | (~w936 & w1556) | (w821 & w1556);
assign w892 = w310 & w1434;
assign w893 = (pi23 & w1748) | (pi23 & w1581) | (w1748 & w1581);
assign w894 = ~w1135 & ~w1326;
assign w895 = w975 & w1491;
assign w896 = ~w410 & ~w1259;
assign w897 = w1147 & w1684;
assign w898 = (~w812 & w399) | (~w812 & w1878) | (w399 & w1878);
assign w899 = (~w220 & w420) | (~w220 & w700) | (w420 & w700);
assign w900 = ~w680 & ~w944;
assign w901 = ~w1624 & w226;
assign w902 = w532 & ~w751;
assign w903 = ~w1540 & w702;
assign w904 = (w1218 & w391) | (w1218 & w1168) | (w391 & w1168);
assign w905 = (w578 & w750) | (w578 & ~w48) | (w750 & ~w48);
assign w906 = w778 & pi68;
assign w907 = ~w1353 & ~w847;
assign w908 = (~w1058 & w197) | (~w1058 & w1316) | (w197 & w1316);
assign w909 = ~w1092 & w885;
assign w910 = ~pi63 & ~pi64;
assign w911 = ~w1578 & ~w480;
assign w912 = (~w1596 & w263) | (~w1596 & w1587) | (w263 & w1587);
assign w913 = (~w1412 & w1232) | (~w1412 & w271) | (w1232 & w271);
assign w914 = ~w928 & w65;
assign w915 = (w869 & ~w419) | (w869 & ~w658) | (~w419 & ~w658);
assign w916 = (w1491 & w1796) | (w1491 & w1080) | (w1796 & w1080);
assign w917 = (w1142 & w726) | (w1142 & w473) | (w726 & w473);
assign w918 = w1575 & w55;
assign w919 = ~w361 & w1585;
assign w920 = ~w195 & ~w80;
assign w921 = pi54 & ~pi55;
assign w922 = (~w1930 & w82) | (~w1930 & w751) | (w82 & w751);
assign w923 = ~pi92 & w722;
assign w924 = pi48 & pi49;
assign w925 = ~w547 & w405;
assign w926 = ~pi92 & ~w505;
assign w927 = (w1817 & w449) | (w1817 & w253) | (w449 & w253);
assign w928 = (w1540 & w728) | (w1540 & w1765) | (w728 & w1765);
assign w929 = ~w46 & ~w847;
assign w930 = (w1618 & w1821) | (w1618 & w1910) | (w1821 & w1910);
assign w931 = ~w1305 & ~w1791;
assign w932 = (~w366 & w739) | (~w366 & w327) | (w739 & w327);
assign w933 = (~w1624 & w1087) | (~w1624 & w391) | (w1087 & w391);
assign w934 = (~pi65 & w1474) | (~pi65 & w241) | (w1474 & w241);
assign w935 = ~w109 & w1187;
assign w936 = (w997 & w694) | (w997 & w1849) | (w694 & w1849);
assign w937 = ~w735 & w128;
assign w938 = ~w679 & ~w1269;
assign w939 = ~w179 & ~w1839;
assign w940 = ~w1856 & ~pi71;
assign w941 = (w1069 & w819) | (w1069 & w108) | (w819 & w108);
assign w942 = (~w1930 & w82) | (~w1930 & w1584) | (w82 & w1584);
assign w943 = pi02 & ~w878;
assign w944 = ~pi14 & w580;
assign w945 = ~w365 & ~w1001;
assign w946 = (~w160 & w1811) | (~w160 & w626) | (w1811 & w626);
assign w947 = (w714 & w333) | (w714 & w48) | (w333 & w48);
assign w948 = (~w1491 & w1899) | (~w1491 & w1166) | (w1899 & w1166);
assign w949 = (w1715 & w205) | (w1715 & w1148) | (w205 & w1148);
assign w950 = (~w22 & w386) | (~w22 & w137) | (w386 & w137);
assign w951 = ~w1132 & ~w991;
assign w952 = (~w1596 & w263) | (~w1596 & ~w1885) | (w263 & ~w1885);
assign w953 = ~w1552 & pi50;
assign w954 = (~w48 & w1312) | (~w48 & w585) | (w1312 & w585);
assign w955 = w1326 & w1287;
assign w956 = (w525 & w442) | (w525 & w1480) | (w442 & w1480);
assign w957 = w1719 & ~w185;
assign w958 = ~w634 & ~w1336;
assign w959 = ~w877 & ~w1340;
assign w960 = w1143 & ~w1387;
assign w961 = (w176 & w1342) | (w176 & ~w433) | (w1342 & ~w433);
assign w962 = w1221 & ~w1128;
assign w963 = ~pi78 & pi79;
assign w964 = (w176 & w1342) | (w176 & ~w1651) | (w1342 & ~w1651);
assign w965 = ~w157 & pi80;
assign w966 = (~w48 & w293) | (~w48 & w1724) | (w293 & w1724);
assign w967 = ~w1105 & ~w1150;
assign w968 = ~w550 & ~w643;
assign w969 = w228 & ~w1499;
assign w970 = pi30 & ~pi31;
assign w971 = (~w1360 & w1852) | (~w1360 & w619) | (w1852 & w619);
assign w972 = (w1708 & w22) | (w1708 & ~w1773) | (w22 & ~w1773);
assign w973 = w1241 & ~w971;
assign w974 = (w1128 & w16) | (w1128 & w1142) | (w16 & w1142);
assign w975 = (w1358 & w147) | (w1358 & w1054) | (w147 & w1054);
assign w976 = (~w1726 & w1324) | (~w1726 & w175) | (w1324 & w175);
assign w977 = w474 & ~w1464;
assign w978 = (~w1491 & w248) | (~w1491 & w1445) | (w248 & w1445);
assign w979 = ~pi38 & w644;
assign w980 = ~w1132 & w474;
assign w981 = (w1491 & w555) | (w1491 & w61) | (w555 & w61);
assign w982 = ~w1552 & ~w980;
assign w983 = ~w238 & ~w366;
assign w984 = (~pi44 & w764) | (~pi44 & w564) | (w764 & w564);
assign w985 = (~w1491 & w113) | (~w1491 & w905) | (w113 & w905);
assign w986 = (~w1540 & w190) | (~w1540 & w1330) | (w190 & w1330);
assign w987 = (w1480 & w865) | (w1480 & ~w1540) | (w865 & ~w1540);
assign w988 = (w1817 & w1057) | (w1817 & w196) | (w1057 & w196);
assign w989 = w509 & ~w149;
assign w990 = (w1321 & w1802) | (w1321 & w1773) | (w1802 & w1773);
assign w991 = w173 & ~w474;
assign w992 = pi06 & pi07;
assign w993 = (w1805 & w375) | (w1805 & ~w1849) | (w375 & ~w1849);
assign w994 = (~w799 & w1907) | (~w799 & ~w255) | (w1907 & ~w255);
assign w995 = ~w1635 & ~w539;
assign w996 = pi80 & ~w413;
assign w997 = (w220 & w1190) | (w220 & w879) | (w1190 & w879);
assign w998 = (~w1549 & ~w1431) | (~w1549 & ~w946) | (~w1431 & ~w946);
assign w999 = ~pi06 & pi07;
assign w1000 = w1132 & ~w924;
assign w1001 = (~w1885 & w1661) | (~w1885 & w1753) | (w1661 & w1753);
assign w1002 = (~w737 & w1791) | (~w737 & w401) | (w1791 & w401);
assign w1003 = (~w1263 & w500) | (~w1263 & w166) | (w500 & w166);
assign w1004 = (w1817 & w457) | (w1817 & w1517) | (w457 & w1517);
assign w1005 = ~w857 & ~w1098;
assign w1006 = ~w772 & ~w984;
assign w1007 = (~w1928 & w1613) | (~w1928 & w1015) | (w1613 & w1015);
assign w1008 = ~w46 & ~w907;
assign w1009 = w1360 & ~w1684;
assign w1010 = ~pi08 & w1412;
assign w1011 = ~w787 & w1421;
assign w1012 = ~w1725 & ~w1100;
assign w1013 = (~w60 & w1473) | (~w60 & w1402) | (w1473 & w1402);
assign w1014 = pi36 & ~pi37;
assign w1015 = w688 & ~w1928;
assign w1016 = ~w1106 & ~w1713;
assign w1017 = ~pi08 & w1657;
assign w1018 = (~pi83 & w1775) | (~pi83 & w44) | (w1775 & w44);
assign w1019 = (w1491 & w676) | (w1491 & w1864) | (w676 & w1864);
assign w1020 = ~w315 & ~w1093;
assign w1021 = (w146 & w67) | (w146 & w1138) | (w67 & w1138);
assign w1022 = (w1491 & w1830) | (w1491 & w1244) | (w1830 & w1244);
assign w1023 = ~w1931 & pi38;
assign w1024 = w1539 & ~pi86;
assign w1025 = ~pi41 & w896;
assign w1026 = (w167 & w1823) | (w167 & w1849) | (w1823 & w1849);
assign w1027 = (w1817 & w1707) | (w1817 & w765) | (w1707 & w765);
assign w1028 = pi17 & ~w1579;
assign w1029 = (~pi32 & w51) | (~pi32 & w874) | (w51 & w874);
assign w1030 = ~w1614 & ~w1131;
assign w1031 = ~w931 & w1855;
assign w1032 = (pi86 & w1513) | (pi86 & w841) | (w1513 & w841);
assign w1033 = ~pi15 & ~pi16;
assign w1034 = (w1491 & w573) | (w1491 & w1662) | (w573 & w1662);
assign w1035 = (~w1923 & ~w1229) | (~w1923 & w946) | (~w1229 & w946);
assign w1036 = ~w1273 & w1714;
assign w1037 = ~w36 & ~pi20;
assign w1038 = (~w1491 & w427) | (~w1491 & w447) | (w427 & w447);
assign w1039 = (w1358 & w1563) | (w1358 & w307) | (w1563 & w307);
assign w1040 = (~w1491 & w622) | (~w1491 & w1182) | (w622 & w1182);
assign w1041 = w254 & ~w0;
assign w1042 = w273 & ~pi89;
assign w1043 = (w1495 & w544) | (w1495 & ~w1289) | (w544 & ~w1289);
assign w1044 = w1750 & pi89;
assign w1045 = pi32 & ~w1231;
assign w1046 = ~w1575 & ~pi47;
assign w1047 = w1684 & pi59;
assign w1048 = ~w1478 & ~w209;
assign w1049 = ~w938 & ~w1568;
assign w1050 = ~w1259 & ~w881;
assign w1051 = w1 & ~pi53;
assign w1052 = w1446 & ~w844;
assign w1053 = ~w782 & ~w1566;
assign w1054 = (w350 & w1883) | (w350 & w422) | (w1883 & w422);
assign w1055 = ~w210 & ~w1228;
assign w1056 = (~w1423 & w1196) | (~w1423 & w946) | (w1196 & w946);
assign w1057 = (w576 & w609) | (w576 & w189) | (w609 & w189);
assign w1058 = ~w1382 & ~w1851;
assign w1059 = w138 & ~w350;
assign w1060 = (w1917 & w1631) | (w1917 & ~w1849) | (w1631 & ~w1849);
assign w1061 = (w936 & w1225) | (w936 & w212) | (w1225 & w212);
assign w1062 = w1639 & pi23;
assign w1063 = ~pi80 & w413;
assign w1064 = (w255 & w718) | (w255 & w1219) | (w718 & w1219);
assign w1065 = w474 & ~w809;
assign w1066 = ~pi60 & ~pi61;
assign w1067 = (~w1794 & w1117) | (~w1794 & w1533) | (w1117 & w1533);
assign w1068 = (w987 & w88) | (w987 & w1220) | (w88 & w1220);
assign w1069 = w496 & ~w1527;
assign w1070 = (w657 & ~w1713) | (w657 & ~w1666) | (~w1713 & ~w1666);
assign w1071 = (w971 & w1047) | (w971 & w1638) | (w1047 & w1638);
assign w1072 = ~pi01 & pi02;
assign w1073 = (w247 & w380) | (w247 & w340) | (w380 & w340);
assign w1074 = ~w853 & w246;
assign w1075 = (w672 & w1059) | (w672 & ~w1358) | (w1059 & ~w1358);
assign w1076 = w1318 & ~w1549;
assign w1077 = (~w440 & ~w1434) | (~w440 & w1799) | (~w1434 & w1799);
assign w1078 = (w1128 & w16) | (w1128 & w1773) | (w16 & w1773);
assign w1079 = (w1882 & w312) | (w1882 & w1358) | (w312 & w1358);
assign w1080 = (w285 & w129) | (w285 & w48) | (w129 & w48);
assign w1081 = w557 & ~w1750;
assign w1082 = (w1626 & w531) | (w1626 & w320) | (w531 & w320);
assign w1083 = ~w1748 & w1551;
assign w1084 = w1815 & ~w247;
assign w1085 = (~w1926 & w835) | (~w1926 & w1475) | (w835 & w1475);
assign w1086 = (w1817 & w701) | (w1817 & w1641) | (w701 & w1641);
assign w1087 = pi29 & ~w1480;
assign w1088 = (~w1380 & w673) | (~w1380 & w584) | (w673 & w584);
assign w1089 = (w1773 & w1260) | (w1773 & w1601) | (w1260 & w1601);
assign w1090 = (w1744 & w823) | (w1744 & ~w530) | (w823 & ~w530);
assign w1091 = (~w1236 & w141) | (~w1236 & w860) | (w141 & w860);
assign w1092 = ~w1771 & ~w1852;
assign w1093 = (~pi29 & w487) | (~pi29 & w691) | (w487 & w691);
assign w1094 = ~w624 & w1908;
assign w1095 = pi08 & w1657;
assign w1096 = (w220 & w1706) | (w220 & w759) | (w1706 & w759);
assign w1097 = ~w1184 & ~w1364;
assign w1098 = w1915 & ~w1694;
assign w1099 = (w1479 & w872) | (w1479 & w265) | (w872 & w265);
assign w1100 = pi87 & pi88;
assign w1101 = w1160 & ~pi92;
assign w1102 = (w1566 & w1177) | (w1566 & ~w1387) | (w1177 & ~w1387);
assign w1103 = w1337 & ~w1536;
assign w1104 = ~w115 & ~w1433;
assign w1105 = ~w1246 & w1407;
assign w1106 = (~w1643 & w1608) | (~w1643 & w791) | (w1608 & w791);
assign w1107 = (~w997 & w252) | (~w997 & w280) | (w252 & w280);
assign w1108 = ~w1703 & ~w1383;
assign w1109 = (w1718 & w490) | (w1718 & w703) | (w490 & w703);
assign w1110 = (w247 & w425) | (w247 & w1913) | (w425 & w1913);
assign w1111 = (~w997 & w811) | (~w997 & w690) | (w811 & w690);
assign w1112 = ~pi95 & w1783;
assign w1113 = (w1540 & w1299) | (w1540 & w68) | (w1299 & w68);
assign w1114 = (w256 & w478) | (w256 & w1600) | (w478 & w1600);
assign w1115 = (~w742 & w255) | (~w742 & w1206) | (w255 & w1206);
assign w1116 = w1815 & ~w1021;
assign w1117 = w1548 & ~w1794;
assign w1118 = (w1885 & w922) | (w1885 & w1876) | (w922 & w1876);
assign w1119 = (w1523 & w1126) | (w1523 & ~w1925) | (w1126 & ~w1925);
assign w1120 = pi38 & w644;
assign w1121 = pi60 & ~pi61;
assign w1122 = ~w1415 & w200;
assign w1123 = (~pi03 & w1238) | (~pi03 & w183) | (w1238 & w183);
assign w1124 = (~w1410 & w1427) | (~w1410 & w1151) | (w1427 & w1151);
assign w1125 = ~w1106 & w657;
assign w1126 = ~w1639 & w507;
assign w1127 = pi01 & ~pi02;
assign w1128 = (~w501 & w35) | (~w501 & w1570) | (w35 & w1570);
assign w1129 = w410 & ~w244;
assign w1130 = w267 & ~w1666;
assign w1131 = w1572 & w1325;
assign w1132 = ~pi45 & ~pi46;
assign w1133 = ~pi72 & pi73;
assign w1134 = (~w888 & ~w50) | (~w888 & ~w1358) | (~w50 & ~w1358);
assign w1135 = pi24 & pi25;
assign w1136 = pi53 & ~w1283;
assign w1137 = w1008 & ~w1274;
assign w1138 = ~w89 & ~w1240;
assign w1139 = (w224 & w1834) | (w224 & ~w1078) | (w1834 & ~w1078);
assign w1140 = (~pi95 & w855) | (~pi95 & w1344) | (w855 & w1344);
assign w1141 = w687 & w1028;
assign w1142 = (w1091 & w1333) | (w1091 & w350) | (w1333 & w350);
assign w1143 = ~w1450 & ~w335;
assign w1144 = ~w105 & ~w1760;
assign w1145 = w1241 & ~w1380;
assign w1146 = (w786 & w319) | (w786 & w1833) | (w319 & w1833);
assign w1147 = ~pi54 & ~pi55;
assign w1148 = (~w213 & w120) | (~w213 & w1306) | (w120 & w1306);
assign w1149 = (w1181 & w11) | (w1181 & ~w576) | (w11 & ~w576);
assign w1150 = ~w579 & ~w1718;
assign w1151 = (~pi35 & ~w1207) | (~pi35 & w1174) | (~w1207 & w1174);
assign w1152 = (~w1358 & w293) | (~w1358 & w1724) | (w293 & w1724);
assign w1153 = (w1491 & w1538) | (w1491 & w1157) | (w1538 & w1157);
assign w1154 = ~w41 & ~pi32;
assign w1155 = (~w576 & w1468) | (~w576 & w669) | (w1468 & w669);
assign w1156 = (~pi68 & w443) | (~pi68 & w346) | (w443 & w346);
assign w1157 = (w48 & w520) | (w48 & w715) | (w520 & w715);
assign w1158 = pi06 & ~pi07;
assign w1159 = w1506 & ~w100;
assign w1160 = ~w880 & ~w163;
assign w1161 = pi47 & ~w1554;
assign w1162 = (~w1803 & w1922) | (~w1803 & w417) | (w1922 & w417);
assign w1163 = ~w948 & w502;
assign w1164 = w290 & ~w1066;
assign w1165 = (pi80 & w985) | (pi80 & w810) | (w985 & w810);
assign w1166 = (~w610 & w20) | (~w610 & w265) | (w20 & w265);
assign w1167 = ~w1033 & ~w216;
assign w1168 = ~w731 & w1270;
assign w1169 = (w1491 & w152) | (w1491 & w1230) | (w152 & w1230);
assign w1170 = (~w59 & w1468) | (~w59 & w669) | (w1468 & w669);
assign w1171 = (w1491 & w40) | (w1491 & w1136) | (w40 & w1136);
assign w1172 = (~w1207 & w1788) | (~w1207 & w475) | (w1788 & w475);
assign w1173 = ~w737 & ~w1645;
assign w1174 = ~w1915 & ~pi35;
assign w1175 = (~w1838 & w758) | (~w1838 & w830) | (w758 & w830);
assign w1176 = w1066 & ~pi65;
assign w1177 = (~w335 & ~w1450) | (~w335 & w1566) | (~w1450 & w1566);
assign w1178 = pi93 & pi94;
assign w1179 = (~w1470 & w962) | (~w1470 & w397) | (w962 & w397);
assign w1180 = w1343 & ~w751;
assign w1181 = (~pi92 & w1415) | (~pi92 & w1101) | (w1415 & w1101);
assign w1182 = (w1276 & w110) | (w1276 & ~w48) | (w110 & ~w48);
assign w1183 = (pi47 & ~w1575) | (pi47 & w1300) | (~w1575 & w1300);
assign w1184 = ~w1261 & w627;
assign w1185 = ~w854 & ~w1458;
assign w1186 = (~w1491 & w499) | (~w1491 & w1795) | (w499 & w1795);
assign w1187 = ~w992 & ~pi11;
assign w1188 = (w355 & w1171) | (w355 & w1428) | (w1171 & w1428);
assign w1189 = (~pi68 & w981) | (~pi68 & ~w708) | (w981 & ~w708);
assign w1190 = (w1618 & w504) | (w1618 & w521) | (w504 & w521);
assign w1191 = (w1882 & w312) | (w1882 & w48) | (w312 & w48);
assign w1192 = ~w1748 & w1590;
assign w1193 = (pi32 & w1820) | (pi32 & w1365) | (w1820 & w1365);
assign w1194 = ~w548 & w1144;
assign w1195 = ~w1192 & ~w1782;
assign w1196 = w46 & ~w1423;
assign w1197 = (w1892 & w288) | (w1892 & w1078) | (w288 & w1078);
assign w1198 = (pi20 & w1162) | (pi20 & w337) | (w1162 & w337);
assign w1199 = pi21 & pi22;
assign w1200 = (w723 & w391) | (w723 & w1168) | (w391 & w1168);
assign w1201 = ~w1273 & w1920;
assign w1202 = (w576 & w314) | (w576 & w70) | (w314 & w70);
assign w1203 = w992 & ~w1286;
assign w1204 = (~w1618 & w957) | (~w1618 & w775) | (w957 & w775);
assign w1205 = (~w1751 & w64) | (~w1751 & w1417) | (w64 & w1417);
assign w1206 = (w69 & w1800) | (w69 & w1687) | (w1800 & w1687);
assign w1207 = ~w1694 & ~w857;
assign w1208 = (pi89 & ~w273) | (pi89 & w1406) | (~w273 & w1406);
assign w1209 = (~pi38 & w1005) | (~pi38 & w1317) | (w1005 & w1317);
assign w1210 = w123 & pi95;
assign w1211 = (~pi35 & w928) | (~pi35 & w1612) | (w928 & w1612);
assign w1212 = ~w731 & w1266;
assign w1213 = (w783 & w1280) | (w783 & ~w1358) | (w1280 & ~w1358);
assign w1214 = w105 & pi83;
assign w1215 = ~w1165 & ~w440;
assign w1216 = w835 & ~w1926;
assign w1217 = ~w1095 & ~w1843;
assign w1218 = ~w1326 & ~w232;
assign w1219 = w632 & ~w1875;
assign w1220 = (w568 & w1120) | (w568 & w1560) | (w1120 & w1560);
assign w1221 = ~w1500 & ~pi83;
assign w1222 = (~w1423 & w1196) | (~w1423 & w1274) | (w1196 & w1274);
assign w1223 = w460 & w128;
assign w1224 = ~w1050 & w1695;
assign w1225 = (w485 & w1607) | (w485 & w1606) | (w1607 & w1606);
assign w1226 = w490 & ~w1591;
assign w1227 = (~w1542 & w762) | (~w1542 & w1347) | (w762 & w1347);
assign w1228 = w1781 & ~w58;
assign w1229 = (~w847 & ~w46) | (~w847 & w1923) | (~w46 & w1923);
assign w1230 = (w1031 & w155) | (w1031 & w1651) | (w155 & w1651);
assign w1231 = ~w41 & ~w919;
assign w1232 = w1781 & ~w1017;
assign w1233 = (~w1021 & w368) | (~w1021 & w1088) | (w368 & w1088);
assign w1234 = pi83 & ~w684;
assign w1235 = (w723 & w1716) | (w723 & w1212) | (w1716 & w1212);
assign w1236 = pi72 & pi73;
assign w1237 = (~w937 & w1250) | (~w937 & w1257) | (w1250 & w1257);
assign w1238 = ~pi00 & ~w877;
assign w1239 = ~w1870 & ~w1123;
assign w1240 = ~w1259 & w410;
assign w1241 = ~w1147 & ~w1305;
assign w1242 = w43 & ~w743;
assign w1243 = (w664 & w232) | (w664 & w122) | (w232 & w122);
assign w1244 = (w1652 & w1498) | (w1652 & w1138) | (w1498 & w1138);
assign w1245 = (~w911 & w1338) | (~w911 & w1007) | (w1338 & w1007);
assign w1246 = (~w592 & w1848) | (~w592 & w565) | (w1848 & w565);
assign w1247 = (~w1666 & ~w683) | (~w1666 & ~w1618) | (~w683 & ~w1618);
assign w1248 = ~w1616 & ~w1033;
assign w1249 = (~w1684 & w1009) | (~w1684 & w719) | (w1009 & w719);
assign w1250 = ~w460 & w735;
assign w1251 = w924 & ~w1;
assign w1252 = (~pi44 & w1050) | (~pi44 & w1487) | (w1050 & w1487);
assign w1253 = (w213 & w553) | (w213 & w491) | (w553 & w491);
assign w1254 = w944 & ~w1028;
assign w1255 = (w783 & w1280) | (w783 & ~w48) | (w1280 & ~w48);
assign w1256 = (~w101 & w1801) | (~w101 & w461) | (w1801 & w461);
assign w1257 = ~w460 & w390;
assign w1258 = (w971 & w1459) | (w971 & w732) | (w1459 & w732);
assign w1259 = ~pi39 & ~pi40;
assign w1260 = (pi77 & ~w812) | (pi77 & w836) | (~w812 & w836);
assign w1261 = (~w1803 & w1290) | (~w1803 & w1457) | (w1290 & w1457);
assign w1262 = ~w1656 & ~w56;
assign w1263 = ~w150 & ~w934;
assign w1264 = (w551 & w537) | (w551 & w1331) | (w537 & w1331);
assign w1265 = (~w235 & w1558) | (~w235 & w1549) | (w1558 & w1549);
assign w1266 = w1135 & ~pi29;
assign w1267 = (w48 & w1281) | (w48 & w28) | (w1281 & w28);
assign w1268 = (~w997 & w1460) | (~w997 & w117) | (w1460 & w117);
assign w1269 = (w52 & w142) | (w52 & w642) | (w142 & w642);
assign w1270 = w1135 & pi29;
assign w1271 = (~w1817 & w1453) | (~w1817 & w603) | (w1453 & w603);
assign w1272 = (~w1817 & w1454) | (~w1817 & w264) | (w1454 & w264);
assign w1273 = ~w453 & ~w141;
assign w1274 = (~w160 & w1811) | (~w160 & w1058) | (w1811 & w1058);
assign w1275 = ~pi60 & pi61;
assign w1276 = (w415 & w309) | (w415 & ~w1142) | (w309 & ~w1142);
assign w1277 = ~w1820 & w529;
assign w1278 = (w997 & w638) | (w997 & w1824) | (w638 & w1824);
assign w1279 = (~w630 & w1711) | (~w630 & w408) | (w1711 & w408);
assign w1280 = w1906 & ~w1773;
assign w1281 = w1737 & ~pi65;
assign w1282 = (w1207 & w1541) | (w1207 & w1600) | (w1541 & w1600);
assign w1283 = (w843 & w819) | (w843 & w108) | (w819 & w108);
assign w1284 = (~pi62 & w948) | (~pi62 & w1169) | (w948 & w1169);
assign w1285 = w809 & ~pi53;
assign w1286 = ~pi09 & ~pi10;
assign w1287 = ~w1135 & ~pi29;
assign w1288 = (~w388 & w421) | (~w388 & w484) | (w421 & w484);
assign w1289 = (w1491 & w1673) | (w1491 & w464) | (w1673 & w464);
assign w1290 = w1248 & w1536;
assign w1291 = (~w220 & w1544) | (~w220 & w607) | (w1544 & w607);
assign w1292 = pi84 & ~pi85;
assign w1293 = w1838 & w1443;
assign w1294 = (pi77 & ~w812) | (pi77 & w1906) | (~w812 & w1906);
assign w1295 = (~pi71 & w1646) | (~pi71 & w27) | (w1646 & w27);
assign w1296 = ~w1589 & ~w35;
assign w1297 = w929 & ~w946;
assign w1298 = (~w1817 & w1170) | (~w1817 & w1155) | (w1170 & w1155);
assign w1299 = (w1193 & w1045) | (w1193 & ~w1480) | (w1045 & ~w1480);
assign w1300 = (w1527 & w74) | (w1527 & w1440) | (w74 & w1440);
assign w1301 = (w746 & w315) | (w746 & w432) | (w315 & w432);
assign w1302 = ~w356 & ~w1268;
assign w1303 = ~w1451 & ~w184;
assign w1304 = (~pi56 & w1092) | (~pi56 & w736) | (w1092 & w736);
assign w1305 = ~pi57 & ~pi58;
assign w1306 = (~w958 & w777) | (~w958 & w130) | (w777 & w130);
assign w1307 = pi14 & ~w580;
assign w1308 = (w1927 & w990) | (w1927 & w1358) | (w990 & w1358);
assign w1309 = (pi50 & w403) | (pi50 & w1034) | (w403 & w1034);
assign w1310 = (w577 & w343) | (w577 & w1314) | (w343 & w1314);
assign w1311 = w556 & pi44;
assign w1312 = ~w1737 & ~pi65;
assign w1313 = (w199 & w773) | (w199 & w16) | (w773 & w16);
assign w1314 = (pi71 & w916) | (pi71 & w1818) | (w916 & w1818);
assign w1315 = ~pi02 & ~w635;
assign w1316 = w929 & ~w1811;
assign w1317 = w1931 & ~pi38;
assign w1318 = (~w914 & w1443) | (~w914 & w837) | (w1443 & w837);
assign w1319 = (w869 & w1919) | (w869 & w23) | (w1919 & w23);
assign w1320 = (pi56 & w1576) | (pi56 & w1397) | (w1576 & w1397);
assign w1321 = ~w1296 & w965;
assign w1322 = ~w1553 & w1100;
assign w1323 = ~w746 & ~w1083;
assign w1324 = w398 & ~w1726;
assign w1325 = (w278 & ~w538) | (w278 & ~w220) | (~w538 & ~w220);
assign w1326 = ~pi24 & ~pi25;
assign w1327 = ~pi68 & w806;
assign w1328 = ~w536 & ~w1489;
assign w1329 = w1575 & ~pi47;
assign w1330 = ~w554 & ~w709;
assign w1331 = (w1083 & ~w1851) | (w1083 & w1377) | (~w1851 & w1377);
assign w1332 = (w731 & w1624) | (w731 & w865) | (w1624 & w865);
assign w1333 = ~w1236 & ~w455;
assign w1334 = ~w894 & pi26;
assign w1335 = w1100 & ~w505;
assign w1336 = (w1643 & w1189) | (w1643 & w566) | (w1189 & w566);
assign w1337 = pi12 & pi13;
assign w1338 = (w1792 & w1578) | (w1792 & w1362) | (w1578 & w1362);
assign w1339 = ~w1066 & ~w910;
assign w1340 = ~pi01 & ~pi02;
assign w1341 = w173 & pi47;
assign w1342 = pi62 & ~w796;
assign w1343 = ~w1434 & ~w1215;
assign w1344 = ~w123 & ~pi95;
assign w1345 = ~w404 & ~w1738;
assign w1346 = (w59 & w606) | (w59 & w1659) | (w606 & w1659);
assign w1347 = ~w460 & ~w937;
assign w1348 = w273 & w1044;
assign w1349 = ~w384 & pi62;
assign w1350 = (~w1470 & w1530) | (~w1470 & w804) | (w1530 & w804);
assign w1351 = (~w925 & w448) | (~w925 & w171) | (w448 & w171);
assign w1352 = w1324 & ~w1726;
assign w1353 = (pi32 & w51) | (pi32 & w705) | (w51 & w705);
assign w1354 = ~w681 & ~w935;
assign w1355 = w664 & ~w723;
assign w1356 = (~pi38 & w1826) | (~pi38 & w7) | (w1826 & w7);
assign w1357 = pi66 & ~pi67;
assign w1358 = (w1021 & w429) | (w1021 & w738) | (w429 & w738);
assign w1359 = pi08 & w1412;
assign w1360 = pi54 & pi55;
assign w1361 = ~w403 & w217;
assign w1362 = w480 & w1792;
assign w1363 = ~w1236 & ~w1510;
assign w1364 = ~pi17 & ~w1579;
assign w1365 = w41 & pi32;
assign w1366 = (pi89 & ~w273) | (pi89 & w1879) | (~w273 & w1879);
assign w1367 = ~w1931 & ~pi38;
assign w1368 = ~w292 & ~w1566;
assign w1369 = w1147 & ~pi59;
assign w1370 = (~w105 & w548) | (~w105 & w22) | (w548 & w22);
assign w1371 = (~pi26 & w1372) | (~pi26 & w724) | (w1372 & w724);
assign w1372 = w894 & ~pi26;
assign w1373 = (w167 & w1823) | (w167 & w694) | (w1823 & w694);
assign w1374 = w1377 & ~w69;
assign w1375 = w679 & w579;
assign w1376 = ~w1115 & ~w1543;
assign w1377 = ~w1162 & w1037;
assign w1378 = w657 & ~w104;
assign w1379 = ~w1298 & w1043;
assign w1380 = ~w1360 & ~w56;
assign w1381 = ~pi86 & ~w1513;
assign w1382 = (pi26 & w986) | (pi26 & w331) | (w986 & w331);
assign w1383 = (~pi59 & w648) | (~pi59 & w1595) | (w648 & w1595);
assign w1384 = ~pi95 & w441;
assign w1385 = w875 & ~w173;
assign w1386 = (~pi50 & w951) | (~pi50 & w394) | (w951 & w394);
assign w1387 = ~w1928 & ~w1853;
assign w1388 = (~w1020 & w1301) | (~w1020 & ~w1382) | (w1301 & ~w1382);
assign w1389 = (~w1715 & w91) | (~w1715 & w1052) | (w91 & w1052);
assign w1390 = (w516 & w306) | (w516 & w1740) | (w306 & w1740);
assign w1391 = w46 & ~w1353;
assign w1392 = ~pi56 & ~w1262;
assign w1393 = pi11 & w381;
assign w1394 = (w220 & w1632) | (w220 & w472) | (w1632 & w472);
assign w1395 = (w1491 & w1933) | (w1491 & w208) | (w1933 & w208);
assign w1396 = ~pi08 & ~w1412;
assign w1397 = (w1491 & w438) | (w1491 & w1452) | (w438 & w1452);
assign w1398 = (w1437 & w386) | (w1437 & w1128) | (w386 & w1128);
assign w1399 = (w530 & w734) | (w530 & w95) | (w734 & w95);
assign w1400 = (w1491 & w975) | (w1491 & w1856) | (w975 & w1856);
assign w1401 = (~w1248 & w26) | (~w1248 & ~w1536) | (w26 & ~w1536);
assign w1402 = w361 & ~w60;
assign w1403 = w1 & w1285;
assign w1404 = ~w809 & ~pi53;
assign w1405 = (w672 & w1059) | (w672 & ~w48) | (w1059 & ~w48);
assign w1406 = ~w1750 & pi89;
assign w1407 = (~w1817 & w38) | (~w1817 & w631) | (w38 & w631);
assign w1408 = (~w1097 & w301) | (~w1097 & w1564) | (w301 & w1564);
assign w1409 = w160 & w1382;
assign w1410 = (w1013 & w1560) | (w1013 & w865) | (w1560 & w865);
assign w1411 = w812 & pi77;
assign w1412 = ~w254 & ~w1286;
assign w1413 = (~w1020 & w1301) | (~w1020 & w1083) | (w1301 & w1083);
assign w1414 = (~w1491 & w1134) | (~w1491 & w611) | (w1134 & w611);
assign w1415 = ~w1553 & ~w1854;
assign w1416 = ~w119 & ~w1689;
assign w1417 = (~pi29 & w731) | (~pi29 & w586) | (w731 & w586);
assign w1418 = ~w1320 & ~w431;
assign w1419 = (~w450 & w1319) | (~w450 & w493) | (w1319 & w493);
assign w1420 = pi56 & ~w1262;
assign w1421 = (~w1491 & w1911) | (~w1491 & w172) | (w1911 & w172);
assign w1422 = w677 & ~w1393;
assign w1423 = ~w45 & ~w1029;
assign w1424 = ~w1775 & w800;
assign w1425 = (w414 & w1547) | (w414 & ~w1849) | (w1547 & ~w1849);
assign w1426 = (~w1021 & w1671) | (~w1021 & w1249) | (w1671 & w1249);
assign w1427 = ~w1207 & ~pi35;
assign w1428 = (w1491 & w1463) | (w1491 & w1526) | (w1463 & w1526);
assign w1429 = ~w1434 & ~w440;
assign w1430 = pi35 & ~w928;
assign w1431 = (~w692 & w1391) | (~w692 & w641) | (w1391 & w641);
assign w1432 = (~w389 & w1222) | (~w389 & w1056) | (w1222 & w1056);
assign w1433 = (~w997 & w1571) | (~w997 & w590) | (w1571 & w590);
assign w1434 = ~w489 & w1350;
assign w1435 = (w1751 & w871) | (w1751 & w379) | (w871 & w379);
assign w1436 = w90 & ~w896;
assign w1437 = w105 & w1884;
assign w1438 = (~w1491 & w1213) | (~w1491 & w1255) | (w1213 & w1255);
assign w1439 = ~w1639 & ~pi23;
assign w1440 = w1575 & w1341;
assign w1441 = (~w735 & ~w390) | (~w735 & w937) | (~w390 & w937);
assign w1442 = (~w1510 & w497) | (~w1510 & w138) | (w497 & w138);
assign w1443 = (pi38 & w1826) | (pi38 & w1068) | (w1826 & w1068);
assign w1444 = (pi47 & w1889) | (pi47 & w125) | (w1889 & w125);
assign w1445 = pi59 & ~w1110;
assign w1446 = (~w1919 & w657) | (~w1919 & w1729) | (w657 & w1729);
assign w1447 = w1858 & w1856;
assign w1448 = (~w1491 & w1385) | (~w1491 & w316) | (w1385 & w316);
assign w1449 = w731 & ~w1332;
assign w1450 = ~w286 & w1186;
assign w1451 = (w255 & w106) | (w255 & w1734) | (w106 & w1734);
assign w1452 = (w909 & w14) | (w909 & w247) | (w14 & w247);
assign w1453 = (w754 & w1381) | (w754 & ~w974) | (w1381 & ~w974);
assign w1454 = w1725 & ~w576;
assign w1455 = w1339 & ~w48;
assign w1456 = ~w588 & ~w1798;
assign w1457 = w1248 & ~w1103;
assign w1458 = ~w1163 & w869;
assign w1459 = w1684 & ~pi59;
assign w1460 = (w636 & w406) | (w636 & ~w694) | (w406 & ~w694);
assign w1461 = (~w69 & w1198) | (~w69 & w1374) | (w1198 & w1374);
assign w1462 = (~w1491 & ~w1673) | (~w1491 & ~w464) | (~w1673 & ~w464);
assign w1463 = ~w1 & ~w941;
assign w1464 = ~w924 & ~w809;
assign w1465 = w1500 & w105;
assign w1466 = ~w548 & ~w105;
assign w1467 = (pi95 & w855) | (pi95 & w1865) | (w855 & w1865);
assign w1468 = w1335 & ~w505;
assign w1469 = ~w992 & ~w254;
assign w1470 = (w1491 & w1822) | (w1491 & w153) | (w1822 & w153);
assign w1471 = w1901 & ~w708;
assign w1472 = w802 & ~w608;
assign w1473 = w1326 & ~w1585;
assign w1474 = (~w1491 & w768) | (~w1491 & w1099) | (w768 & w1099);
assign w1475 = ~w809 & ~w1771;
assign w1476 = ~w1011 & ~w624;
assign w1477 = ~pi44 & ~w1916;
assign w1478 = (w1715 & w930) | (w1715 & w225) | (w930 & w225);
assign w1479 = (~w1737 & w1508) | (~w1737 & w1164) | (w1508 & w1164);
assign w1480 = ~w1135 & w238;
assign w1481 = (~pi53 & w1814) | (~pi53 & w159) | (w1814 & w159);
assign w1482 = ~w1539 & ~pi86;
assign w1483 = (w1546 & w1769) | (w1546 & ~w1651) | (w1769 & ~w1651);
assign w1484 = w384 & pi62;
assign w1485 = (~w1491 & w488) | (~w1491 & w954) | (w488 & w954);
assign w1486 = (w339 & w13) | (w339 & w1410) | (w13 & w1410);
assign w1487 = w556 & ~pi44;
assign w1488 = pi47 & ~w298;
assign w1489 = (~w1816 & w31) | (~w1816 & w899) | (w31 & w899);
assign w1490 = (pi89 & w1909) | (pi89 & w1348) | (w1909 & w1348);
assign w1491 = (~w1540 & w1537) | (~w1540 & w1114) | (w1537 & w1114);
assign w1492 = (w1529 & w979) | (w1529 & w1013) | (w979 & w1013);
assign w1493 = (~w997 & w165) | (~w997 & w1060) | (w165 & w1060);
assign w1494 = pi32 & w1231;
assign w1495 = (pi92 & w1415) | (pi92 & w1835) | (w1415 & w1835);
assign w1496 = w894 & pi26;
assign w1497 = (w1540 & w492) | (w1540 & w8) | (w492 & w8);
assign w1498 = ~pi50 & w982;
assign w1499 = ~pi06 & ~pi07;
assign w1500 = ~pi78 & ~pi79;
assign w1501 = w1343 & ~w1351;
assign w1502 = (pi95 & w1467) | (pi95 & w149) | (w1467 & w149);
assign w1503 = (w249 & w127) | (w249 & w1849) | (w127 & w1849);
assign w1504 = (w845 & w1063) | (w845 & w1142) | (w1063 & w1142);
assign w1505 = (w1118 & w942) | (w1118 & w1849) | (w942 & w1849);
assign w1506 = (w1443 & w526) | (w1443 & w1293) | (w526 & w1293);
assign w1507 = (w1277 & w1494) | (w1277 & w1480) | (w1494 & w1480);
assign w1508 = w737 & ~w1737;
assign w1509 = (~w477 & w1779) | (~w477 & w1297) | (w1779 & w1297);
assign w1510 = ~pi72 & ~pi73;
assign w1511 = (w59 & w1042) | (w59 & w1872) | (w1042 & w1872);
assign w1512 = (w1618 & w613) | (w1618 & w1067) | (w613 & w1067);
assign w1513 = ~w1539 & ~w158;
assign w1514 = (~w592 & w1081) | (~w592 & w1741) | (w1081 & w1741);
assign w1515 = (pi50 & w951) | (pi50 & w593) | (w951 & w593);
assign w1516 = ~w157 & ~pi80;
assign w1517 = (w1122 & w1562) | (w1122 & w59) | (w1562 & w59);
assign w1518 = (w576 & w1780) | (w576 & w1691) | (w1780 & w1691);
assign w1519 = (w655 & w569) | (w655 & w345) | (w569 & w345);
assign w1520 = (~pi92 & w722) | (~pi92 & w926) | (w722 & w926);
assign w1521 = w1340 & pi03;
assign w1522 = ~w1415 & w652;
assign w1523 = ~w1639 & ~w37;
assign w1524 = (w1491 & w259) | (w1491 & w1183) | (w259 & w1183);
assign w1525 = ~w1766 & ~w1853;
assign w1526 = ~w1 & ~w1283;
assign w1527 = (~w89 & w881) | (~w89 & w170) | (w881 & w170);
assign w1528 = w812 & w1294;
assign w1529 = ~w1005 & w1367;
assign w1530 = ~w812 & ~pi77;
assign w1531 = (w1817 & w29) | (w1817 & w436) | (w29 & w436);
assign w1532 = (~w145 & w1825) | (~w145 & w1323) | (w1825 & w1323);
assign w1533 = (~w646 & w1778) | (~w646 & w275) | (w1778 & w275);
assign w1534 = (w192 & w1827) | (w192 & w1849) | (w1827 & w1849);
assign w1535 = ~w109 & w1709;
assign w1536 = ~pi12 & ~pi13;
assign w1537 = (w256 & w478) | (w256 & w1410) | (w478 & w1410);
assign w1538 = (w1358 & w520) | (w1358 & w715) | (w520 & w715);
assign w1539 = ~w214 & ~w1292;
assign w1540 = (w1803 & w932) | (w1803 & w807) | (w932 & w807);
assign w1541 = w1915 & w1207;
assign w1542 = ~w1379 & ~w39;
assign w1543 = ~w255 & w1461;
assign w1544 = w207 & ~w521;
assign w1545 = (~w1491 & w392) | (~w1491 & w230) | (w392 & w230);
assign w1546 = (~pi62 & w931) | (~pi62 & w755) | (w931 & w755);
assign w1547 = (w308 & w363) | (w308 & w952) | (w363 & w952);
assign w1548 = ~w648 & w140;
assign w1549 = ~w692 & ~w1923;
assign w1550 = ~w1500 & ~w43;
assign w1551 = (~pi23 & w1540) | (~pi23 & w1439) | (w1540 & w1439);
assign w1552 = ~w1702 & ~w818;
assign w1553 = ~pi87 & ~pi88;
assign w1554 = (w1575 & w693) | (w1575 & w1527) | (w693 & w1527);
assign w1555 = (w1201 & w1647) | (w1201 & w350) | (w1647 & w350);
assign w1556 = (w1845 & w269) | (w1845 & ~w721) | (w269 & ~w721);
assign w1557 = ~w311 & ~w1474;
assign w1558 = (w914 & w1356) | (w914 & w1667) | (w1356 & w1667);
assign w1559 = (~w1021 & w1216) | (~w1021 & w1085) | (w1216 & w1085);
assign w1560 = ~w60 & ~w919;
assign w1561 = (~w1549 & ~w1431) | (~w1549 & ~w1274) | (~w1431 & ~w1274);
assign w1562 = pi92 & w722;
assign w1563 = (w1773 & w4) | (w1773 & w156) | (w4 & w156);
assign w1564 = w944 & ~w1097;
assign w1565 = (~w235 & w1558) | (~w235 & w1431) | (w1558 & w1431);
assign w1566 = ~w335 & w1309;
assign w1567 = ~w782 & w1450;
assign w1568 = w1718 & ~w579;
assign w1569 = (w1470 & w824) | (w1470 & w169) | (w824 & w169);
assign w1570 = w1589 & ~w501;
assign w1571 = (w481 & w178) | (w481 & ~w1849) | (w178 & ~w1849);
assign w1572 = ~w1450 & ~w832;
assign w1573 = ~w910 & w1901;
assign w1574 = (pi86 & w1324) | (pi86 & w876) | (w1324 & w876);
assign w1575 = ~w474 & ~w1132;
assign w1576 = (~w1491 & w1582) | (~w1491 & w1559) | (w1582 & w1559);
assign w1577 = (w1491 & w240) | (w1491 & w1073) | (w240 & w1073);
assign w1578 = ~w1576 & w1710;
assign w1579 = ~w1261 & ~w1622;
assign w1580 = (~w1464 & w977) | (~w1464 & w843) | (w977 & w843);
assign w1581 = ~w1540 & w1062;
assign w1582 = (~w247 & w1216) | (~w247 & w1085) | (w1216 & w1085);
assign w1583 = (~pi89 & w1246) | (~pi89 & w645) | (w1246 & w645);
assign w1584 = (w842 & w1885) | (w842 & w1351) | (w1885 & w1351);
assign w1585 = pi27 & pi28;
assign w1586 = ~w1394 & ~w180;
assign w1587 = ~w390 & ~w735;
assign w1588 = (w1358 & w1281) | (w1358 & w28) | (w1281 & w28);
assign w1589 = ~pi75 & ~pi76;
assign w1590 = (pi23 & w1540) | (pi23 & w1623) | (w1540 & w1623);
assign w1591 = w579 & ~w1718;
assign w1592 = pi04 & pi05;
assign w1593 = ~pi03 & ~pi04;
assign w1594 = pi66 & pi67;
assign w1595 = (w1491 & w848) | (w1491 & w706) | (w848 & w706);
assign w1596 = ~w460 & ~w1105;
assign w1597 = (w1737 & w204) | (w1737 & w48) | (w204 & w48);
assign w1598 = (~w301 & w1141) | (~w301 & w374) | (w1141 & w374);
assign w1599 = ~w1307 & ~w944;
assign w1600 = (w1013 & w1560) | (w1013 & w1480) | (w1560 & w1480);
assign w1601 = (pi77 & ~w812) | (pi77 & w1411) | (~w812 & w1411);
assign w1602 = (~w350 & ~w27) | (~w350 & ~w1358) | (~w27 & ~w1358);
assign w1603 = pi95 & ~w801;
assign w1604 = (w247 & w1051) | (w247 & w1403) | (w1051 & w1403);
assign w1605 = pi18 & ~pi19;
assign w1606 = (w1347 & w1237) | (w1347 & w439) | (w1237 & w439);
assign w1607 = (w459 & w1109) | (w459 & w1105) | (w1109 & w1105);
assign w1608 = w1860 & w708;
assign w1609 = (~w350 & w940) | (~w350 & w299) | (w940 & w299);
assign w1610 = ~pi68 & ~w806;
assign w1611 = pi00 & ~w1340;
assign w1612 = (~w1540 & w342) | (~w1540 & w1837) | (w342 & w1837);
assign w1613 = w526 & ~w1841;
assign w1614 = (w220 & w1727) | (w220 & w1399) | (w1727 & w1399);
assign w1615 = (w1358 & w341) | (w1358 & w1504) | (w341 & w1504);
assign w1616 = pi15 & pi16;
assign w1617 = (w1929 & w996) | (w1929 & ~w1470) | (w996 & ~w1470);
assign w1618 = (w1053 & w1653) | (w1053 & w1007) | (w1653 & w1007);
assign w1619 = (pi08 & w543) | (pi08 & w1877) | (w543 & w1877);
assign w1620 = (~pi71 & w1646) | (~pi71 & w350) | (w1646 & w350);
assign w1621 = (w997 & w675) | (w997 & w1534) | (w675 & w1534);
assign w1622 = (w595 & w1401) | (w595 & w1790) | (w1401 & w1790);
assign w1623 = ~w1639 & pi23;
assign w1624 = w1326 & w731;
assign w1625 = (w1181 & w11) | (w1181 & ~w59) | (w11 & ~w59);
assign w1626 = w1749 & ~w658;
assign w1627 = (w48 & w341) | (w48 & w1504) | (w341 & w1504);
assign w1628 = ~pi95 & ~w801;
assign w1629 = ~w985 & w1617;
assign w1630 = ~pi12 & pi13;
assign w1631 = w234 & ~w32;
assign w1632 = (w521 & w1525) | (w521 & w102) | (w1525 & w102);
assign w1633 = (pi56 & w1092) | (pi56 & w428) | (w1092 & w428);
assign w1634 = ~pi00 & ~w1874;
assign w1635 = ~w653 & ~w1698;
assign w1636 = ~w1310 & ~w1125;
assign w1637 = ~w344 & w650;
assign w1638 = w1684 & w144;
assign w1639 = ~w1199 & ~w238;
assign w1640 = ~w1548 & ~w1163;
assign w1641 = (w59 & w1502) | (w59 & w612) | (w1502 & w612);
assign w1642 = ~w543 & w635;
assign w1643 = (~w1491 & w468) | (~w1491 & w1455) | (w468 & w1455);
assign w1644 = (w389 & w1509) | (w389 & w1861) | (w1509 & w1861);
assign w1645 = ~w1305 & w290;
assign w1646 = w1858 & ~pi71;
assign w1647 = ~pi74 & w10;
assign w1648 = ~w105 & w1500;
assign w1649 = pi08 & ~w1657;
assign w1650 = (~w1491 & w753) | (~w1491 & w458) | (w753 & w458);
assign w1651 = (w971 & w1380) | (w971 & w1021) | (w1380 & w1021);
assign w1652 = ~w951 & w625;
assign w1653 = (~w1566 & w744) | (~w1566 & w1567) | (w744 & w1567);
assign w1654 = w1510 & pi77;
assign w1655 = (w1888 & w25) | (w1888 & ~w865) | (w25 & ~w865);
assign w1656 = ~w552 & ~w921;
assign w1657 = ~w1416 & ~w920;
assign w1658 = (w249 & w127) | (w249 & w694) | (w127 & w694);
assign w1659 = (~pi95 & w1140) | (~pi95 & w716) | (w1140 & w716);
assign w1660 = ~w1432 & ~w513;
assign w1661 = (w937 & w1441) | (w937 & ~w751) | (w1441 & ~w751);
assign w1662 = (w352 & w1918) | (w352 & w1138) | (w1918 & w1138);
assign w1663 = (~w1856 & w1818) | (~w1856 & w840) | (w1818 & w840);
assign w1664 = (~w1817 & w359) | (~w1817 & w506) | (w359 & w506);
assign w1665 = ~w893 & ~w1083;
assign w1666 = (w1185 & w130) | (w1185 & w1533) | (w130 & w1533);
assign w1667 = w223 & w914;
assign w1668 = ~w242 & ~w747;
assign w1669 = (w788 & w1785) | (w788 & ~w27) | (w1785 & ~w27);
assign w1670 = (w232 & w376) | (w232 & ~w327) | (w376 & ~w327);
assign w1671 = (~w1684 & w1009) | (~w1684 & w83) | (w1009 & w83);
assign w1672 = w1163 & ~w854;
assign w1673 = (w576 & w59) | (w576 & w1358) | (w59 & w1358);
assign w1674 = ~w857 & w1694;
assign w1675 = ~w1858 & ~pi71;
assign w1676 = w1129 & ~w244;
assign w1677 = (w1207 & w1541) | (w1207 & w1410) | (w1541 & w1410);
assign w1678 = ~pi36 & ~pi37;
assign w1679 = (w437 & w201) | (w437 & w48) | (w201 & w48);
assign w1680 = (~w812 & w399) | (~w812 & w1442) | (w399 & w1442);
assign w1681 = (w1118 & w942) | (w1118 & w694) | (w942 & w694);
assign w1682 = w408 & ~w1142;
assign w1683 = pi95 & w512;
assign w1684 = ~w290 & ~w1305;
assign w1685 = (~w997 & w53) | (~w997 & w993) | (w53 & w993);
assign w1686 = ~w863 & ~w1697;
assign w1687 = w465 & w69;
assign w1688 = ~w778 & pi68;
assign w1689 = ~w228 & ~w1850;
assign w1690 = (w1358 & w1555) | (w1358 & w268) | (w1555 & w268);
assign w1691 = (~w805 & w360) | (~w805 & w1012) | (w360 & w1012);
assign w1692 = (w770 & w1603) | (w770 & ~w576) | (w1603 & ~w576);
assign w1693 = (w579 & w1269) | (w579 & w1375) | (w1269 & w1375);
assign w1694 = pi33 & pi34;
assign w1695 = ~w556 & ~pi44;
assign w1696 = ~w1630 & ~w112;
assign w1697 = ~w838 & ~w1934;
assign w1698 = ~w601 & ~w1747;
assign w1699 = w41 & ~pi32;
assign w1700 = w1711 & ~w630;
assign w1701 = w1915 & pi35;
assign w1702 = ~pi48 & pi49;
assign w1703 = ~w648 & w978;
assign w1704 = ~w1678 & ~w1259;
assign w1705 = (~w1600 & w1427) | (~w1600 & w1151) | (w1427 & w1151);
assign w1706 = (~w261 & w1146) | (~w261 & ~w87) | (w1146 & ~w87);
assign w1707 = (w1078 & w1813) | (w1078 & w1574) | (w1813 & w1574);
assign w1708 = (~w1500 & w1760) | (~w1500 & w408) | (w1760 & w408);
assign w1709 = ~w992 & pi11;
assign w1710 = (~w1491 & w599) | (~w1491 & w19) | (w599 & w19);
assign w1711 = w1902 & ~w630;
assign w1712 = (pi38 & w1005) | (pi38 & w164) | (w1005 & w164);
assign w1713 = w1919 & ~w657;
assign w1714 = ~w1886 & pi74;
assign w1715 = (w220 & w530) | (w220 & w521) | (w530 & w521);
assign w1716 = ~w731 & ~pi29;
assign w1717 = w154 & ~w716;
assign w1718 = ~w1298 & w670;
assign w1719 = w1320 & ~w185;
assign w1720 = (w1817 & w790) | (w1817 & w527) | (w790 & w527);
assign w1721 = (~w540 & w567) | (~w540 & w571) | (w567 & w571);
assign w1722 = (w1491 & w581) | (w1491 & w463) | (w581 & w463);
assign w1723 = (w224 & w1834) | (w224 & ~w974) | (w1834 & ~w974);
assign w1724 = (~w1858 & w840) | (~w1858 & w1339) | (w840 & w1339);
assign w1725 = ~w1750 & ~w1553;
assign w1726 = ~w743 & ~w1750;
assign w1727 = (w521 & w734) | (w521 & w95) | (w734 & w95);
assign w1728 = (w1491 & w749) | (w1491 & w666) | (w749 & w666);
assign w1729 = w1106 & ~w1919;
assign w1730 = (~w1491 & w1736) | (~w1491 & w76) | (w1736 & w76);
assign w1731 = ~pi95 & ~w512;
assign w1732 = ~pi04 & ~pi05;
assign w1733 = pi08 & ~w1412;
assign w1734 = ~w1804 & w1264;
assign w1735 = pi62 & w796;
assign w1736 = (w1669 & w614) | (w1669 & ~w1358) | (w614 & ~w1358);
assign w1737 = ~w1901 & ~w910;
assign w1738 = (~pi71 & w787) | (~pi71 & w495) | (w787 & w495);
assign w1739 = (w437 & w201) | (w437 & w1358) | (w201 & w1358);
assign w1740 = (~w1491 & w1602) | (~w1491 & w1912) | (w1602 & w1912);
assign w1741 = (~w1750 & w557) | (~w1750 & w1550) | (w557 & w1550);
assign w1742 = pi44 & ~w1916;
assign w1743 = (w1653 & w713) | (w1653 & w1935) | (w713 & w1935);
assign w1744 = (~w434 & w34) | (~w434 & w168) | (w34 & w168);
assign w1745 = (~w974 & w1352) | (~w974 & w545) | (w1352 & w545);
assign w1746 = (w936 & w945) | (w936 & w227) | (w945 & w227);
assign w1747 = (w1412 & w1232) | (w1412 & w323) | (w1232 & w323);
assign w1748 = (w1803 & w302) | (w1803 & w1119) | (w302 & w1119);
assign w1749 = ~w1548 & ~w727;
assign w1750 = ~pi84 & ~pi85;
assign w1751 = (w1803 & w1167) | (w1803 & w327) | (w1167 & w327);
assign w1752 = ~w1915 & ~w857;
assign w1753 = (w937 & w1441) | (w937 & ~w842) | (w1441 & ~w842);
assign w1754 = ~w1803 & ~w1696;
assign w1755 = ~w1841 & ~w688;
assign w1756 = w761 & w1165;
assign w1757 = ~w786 & w1443;
assign w1758 = (w339 & w13) | (w339 & w1600) | (w13 & w1600);
assign w1759 = (w974 & w1078) | (w974 & w1358) | (w1078 & w1358);
assign w1760 = w1902 & ~w1500;
assign w1761 = w1587 & ~w842;
assign w1762 = (w1380 & w1047) | (w1380 & w1638) | (w1047 & w1638);
assign w1763 = (w247 & w1071) | (w247 & w1762) | (w1071 & w1762);
assign w1764 = (w997 & w1721) | (w997 & w347) | (w1721 & w347);
assign w1765 = (~w1207 & w1788) | (~w1207 & w92) | (w1788 & w92);
assign w1766 = ~w817 & ~w118;
assign w1767 = ~w948 & w282;
assign w1768 = (w255 & w1840) | (w255 & w730) | (w1840 & w730);
assign w1769 = ~pi62 & ~w796;
assign w1770 = w154 & ~w149;
assign w1771 = ~pi51 & ~pi52;
assign w1772 = ~w1792 & ~w1418;
assign w1773 = (w1091 & w1333) | (w1091 & w27) | (w1333 & w27);
assign w1774 = w267 & ~w683;
assign w1775 = (w329 & w174) | (w329 & ~w1817) | (w174 & ~w1817);
assign w1776 = ~w548 & w1648;
assign w1777 = (w1892 & w288) | (w1892 & w974) | (w288 & w974);
assign w1778 = ~w181 & w431;
assign w1779 = (w1353 & w914) | (w1353 & w218) | (w914 & w218);
assign w1780 = (~w805 & w360) | (~w805 & ~w1100) | (w360 & ~w1100);
assign w1781 = ~w1642 & w1686;
assign w1782 = (~pi23 & w1748) | (~pi23 & w903) | (w1748 & w903);
assign w1783 = (~w59 & w1770) | (~w59 & w1717) | (w1770 & w1717);
assign w1784 = (w1380 & w1459) | (w1380 & w732) | (w1459 & w732);
assign w1785 = ~pi74 & ~w10;
assign w1786 = (w1491 & w1039) | (w1491 & w651) | (w1039 & w651);
assign w1787 = w532 & ~w842;
assign w1788 = w60 & ~w1207;
assign w1789 = ~w1844 & ~w1921;
assign w1790 = (~w1248 & w26) | (~w1248 & w752) | (w26 & w752);
assign w1791 = w1147 & ~w290;
assign w1792 = ~w1814 & w1038;
assign w1793 = (w770 & w1603) | (w770 & ~w59) | (w1603 & ~w59);
assign w1794 = ~w1767 & ~w1284;
assign w1795 = (~w1527 & w1046) | (~w1527 & w699) | (w1046 & w699);
assign w1796 = (w285 & w129) | (w285 & w1358) | (w129 & w1358);
assign w1797 = (w1817 & w707) | (w1817 & w605) | (w707 & w605);
assign w1798 = (w389 & w1532) | (w389 & w416) | (w1532 & w416);
assign w1799 = ~w440 & w1165;
assign w1800 = (~pi20 & w1162) | (~pi20 & w470) | (w1162 & w470);
assign w1801 = w1585 & ~w101;
assign w1802 = pi80 & w413;
assign w1803 = (~w1286 & w109) | (~w1286 & w357) | (w109 & w357);
assign w1804 = ~w1868 & ~w583;
assign w1805 = (~w1584 & w182) | (~w1584 & w1807) | (w182 & w1807);
assign w1806 = w526 & ~w1006;
assign w1807 = w967 & ~w1237;
assign w1808 = w1678 & ~pi41;
assign w1809 = w1198 & ~w1665;
assign w1810 = ~w688 & ~w1613;
assign w1811 = w746 & ~w160;
assign w1812 = w1678 & w896;
assign w1813 = (pi86 & w1324) | (pi86 & w1637) | (w1324 & w1637);
assign w1814 = (~w1491 & w1283) | (~w1491 & w941) | (w1283 & w941);
assign w1815 = ~w809 & pi53;
assign w1816 = ~w782 & ~w1792;
assign w1817 = (w1491 & w48) | (w1491 & w1358) | (w48 & w1358);
assign w1818 = w1594 & ~w1856;
assign w1819 = w1640 & ~w1533;
assign w1820 = ~w361 & ~w1473;
assign w1821 = ~w1108 & ~w646;
assign w1822 = (w1773 & w1142) | (w1773 & w1358) | (w1142 & w1358);
assign w1823 = (w751 & w454) | (w751 & w233) | (w454 & w233);
assign w1824 = (~w1345 & ~w1070) | (~w1345 & w353) | (~w1070 & w353);
assign w1825 = (w1382 & w46) | (w1382 & w1409) | (w46 & w1409);
assign w1826 = (~w444 & w682) | (~w444 & w332) | (w682 & w332);
assign w1827 = (w439 & w1227) | (w439 & w671) | (w1227 & w671);
assign w1828 = w814 & ~w1363;
assign w1829 = ~w1382 & ~w746;
assign w1830 = (w1652 & w1498) | (w1652 & w1527) | (w1498 & w1527);
assign w1831 = ~w797 & ~w1082;
assign w1832 = ~pi56 & w1262;
assign w1833 = w297 & w786;
assign w1834 = pi86 & ~w1513;
assign w1835 = w1160 & pi92;
assign w1836 = ~w373 & ~w490;
assign w1837 = (w887 & w825) | (w887 & w1410) | (w825 & w1410);
assign w1838 = (pi41 & w508) | (pi41 & w850) | (w508 & w850);
assign w1839 = w1772 & w320;
assign w1840 = ~w1195 & ~w618;
assign w1841 = (pi44 & w764) | (pi44 & w1019) | (w764 & w1019);
assign w1842 = w105 & w511;
assign w1843 = ~pi08 & ~w1657;
assign w1844 = ~w519 & ~w12;
assign w1845 = (w1049 & w1693) | (w1049 & ~w1105) | (w1693 & ~w1105);
assign w1846 = pi24 & ~pi25;
assign w1847 = (w1165 & w390) | (w1165 & w1756) | (w390 & w1756);
assign w1848 = (~w273 & w1909) | (~w273 & w1741) | (w1909 & w1741);
assign w1849 = ~w1310 & ~w540;
assign w1850 = ~w1593 & w635;
assign w1851 = w893 & ~w1083;
assign w1852 = w809 & ~w820;
assign w1853 = ~w688 & w1841;
assign w1854 = w1750 & ~w1100;
assign w1855 = ~w384 & ~pi62;
assign w1856 = ~w814 & ~w453;
assign w1857 = (w1021 & w1071) | (w1021 & w1762) | (w1071 & w1762);
assign w1858 = ~pi66 & ~pi67;
assign w1859 = (~w247 & w1671) | (~w247 & w1249) | (w1671 & w1249);
assign w1860 = (~w1491 & w99) | (~w1491 & w1895) | (w99 & w1895);
assign w1861 = (~w477 & w1779) | (~w477 & w908) | (w1779 & w908);
assign w1862 = w1750 & ~pi89;
assign w1863 = w1752 & ~w1600;
assign w1864 = ~w1050 & w629;
assign w1865 = ~w123 & pi95;
assign w1866 = (~w101 & w1801) | (~w101 & w815) | (w1801 & w815);
assign w1867 = w1657 & w1010;
assign w1868 = ~w986 & w81;
assign w1869 = w1657 & ~w846;
assign w1870 = (pi03 & w1611) | (pi03 & w816) | (w1611 & w816);
assign w1871 = (w576 & w1042) | (w576 & w1872) | (w1042 & w1872);
assign w1872 = w273 & w1862;
assign w1873 = w509 & ~w716;
assign w1874 = ~w1072 & ~w1127;
assign w1875 = (~w1377 & w1198) | (~w1377 & w687) | (w1198 & w687);
assign w1876 = (~w1930 & w82) | (~w1930 & w842) | (w82 & w842);
assign w1877 = ~w635 & pi08;
assign w1878 = w497 & ~w1510;
assign w1879 = w273 & pi89;
assign w1880 = w1915 & ~pi35;
assign w1881 = (~pi77 & w489) | (~pi77 & w1569) | (w489 & w1569);
assign w1882 = ~w443 & w1688;
assign w1883 = w1856 & ~pi71;
assign w1884 = w1500 & ~pi83;
assign w1885 = ~w761 & ~w1077;
assign w1886 = ~w1133 & ~w279;
assign w1887 = w1550 & ~w16;
assign w1888 = (~pi32 & w1820) | (~pi32 & w1699) | (w1820 & w1699);
assign w1889 = w89 & ~w1575;
assign w1890 = ~w501 & ~pi83;
assign w1891 = (~pi29 & w731) | (~pi29 & w1287) | (w731 & w1287);
assign w1892 = ~w344 & w1482;
assign w1893 = (w1491 & w1690) | (w1491 & w33) | (w1690 & w33);
assign w1894 = w1066 & ~w1901;
assign w1895 = (w1156 & w1610) | (w1156 & ~w48) | (w1610 & ~w48);
assign w1896 = w1539 & pi86;
assign w1897 = w896 & w1808;
assign w1898 = (~w1491 & w1742) | (~w1491 & w385) | (w1742 & w385);
assign w1899 = (~w610 & w20) | (~w610 & w9) | (w20 & w9);
assign w1900 = w238 & ~w1199;
assign w1901 = pi63 & pi64;
assign w1902 = pi75 & pi76;
assign w1903 = (w1386 & w260) | (w1386 & ~w1527) | (w260 & ~w1527);
assign w1904 = w1008 & ~w946;
assign w1905 = (~pi92 & ~w505) | (~pi92 & w1522) | (~w505 & w1522);
assign w1906 = ~w1510 & pi77;
assign w1907 = (w1851 & ~w1083) | (w1851 & w1875) | (~w1083 & w1875);
assign w1908 = ~w1011 & w1310;
assign w1909 = w743 & ~w273;
assign w1910 = ~w1108 & ~w591;
assign w1911 = (~w1358 & w572) | (~w1358 & w1609) | (w572 & w1609);
assign w1912 = (~w350 & ~w27) | (~w350 & ~w48) | (~w27 & ~w48);
assign w1913 = (w1684 & w897) | (w1684 & w1380) | (w897 & w1380);
assign w1914 = (w1817 & w1777) | (w1817 & w1197) | (w1777 & w1197);
assign w1915 = ~pi30 & ~pi31;
assign w1916 = ~w556 & ~w1240;
assign w1917 = (~w32 & w234) | (~w32 & w193) | (w234 & w193);
assign w1918 = pi50 & w982;
assign w1919 = ~w1474 & w1485;
assign w1920 = ~w1886 & ~pi74;
assign w1921 = w519 & ~w1599;
assign w1922 = ~w377 & ~w327;
assign w1923 = ~w847 & w1353;
assign w1924 = ~pi66 & pi67;
assign w1925 = ~w1616 & ~w589;
assign w1926 = ~w1360 & ~w1147;
assign w1927 = (w1321 & w1802) | (w1321 & w1142) | (w1802 & w1142);
assign w1928 = (w1448 & w1524) | (w1448 & w133) | (w1524 & w133);
assign w1929 = (pi80 & w1296) | (pi80 & w482) | (w1296 & w482);
assign w1930 = ~w313 & ~w789;
assign w1931 = ~w93 & ~w1014;
assign w1932 = ~w232 & w1334;
assign w1933 = (w1527 & w1329) | (w1527 & w918) | (w1329 & w918);
assign w1934 = ~w878 & ~w1315;
assign w1935 = (~w911 & w1338) | (~w911 & w1053) | (w1338 & w1053);
assign w1936 = (~pi11 & w109) | (~pi11 & w483) | (w109 & w483);
assign w1937 = w1694 & ~w1678;
assign one = 1;
assign po00 = ~w411;// level 4
assign po01 = ~w533;// level 6
assign po02 = ~w1055;// level 9
assign po03 = ~w995;// level 11
assign po04 = ~w1789;// level 11
assign po05 = ~w829;// level 11
assign po06 = ~w1376;// level 12
assign po07 = ~w294;// level 12
assign po08 = ~w1303;// level 13
assign po09 = ~w1456;// level 13
assign po10 = ~w1660;// level 13
assign po11 = ~w206;// level 14
assign po12 = ~w766;// level 14
assign po13 = ~w563;// level 14
assign po14 = ~w418;// level 14
assign po15 = ~w1586;// level 14
assign po16 = ~w1030;// level 15
assign po17 = ~w1328;// level 15
assign po18 = ~w939;// level 15
assign po19 = ~w1048;// level 15
assign po20 = ~w1831;// level 15
assign po21 = ~w798;// level 15
assign po22 = ~w856;// level 15
assign po23 = ~w296;// level 15
assign po24 = ~w49;// level 15
assign po25 = ~w237;// level 16
assign po26 = ~w103;// level 16
assign po27 = ~w1104;// level 16
assign po28 = ~w1302;// level 16
assign po29 = ~w503;// level 16
assign po30 = ~w633;// level 16
assign po31 = ~w779;// level 16
endmodule
