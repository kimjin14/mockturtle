module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 , x147 , x148 , x149 , x150 , x151 , x152 , x153 , x154 , x155 , x156 , x157 , x158 , x159 , x160 , x161 , x162 , x163 , x164 , x165 , x166 , x167 , x168 , x169 , x170 , x171 , x172 , x173 , x174 , x175 , x176 , x177 , x178 , x179 , x180 , x181 , x182 , x183 , x184 , x185 , x186 , x187 , x188 , x189 , x190 , x191 , x192 , x193 , x194 , x195 , x196 , x197 , x198 , x199 , x200 , x201 , x202 , x203 , x204 , x205 , x206 , x207 , x208 , x209 , x210 , x211 , x212 , x213 , x214 , x215 , x216 , x217 , x218 , x219 , x220 , x221 , x222 , x223 , x224 , x225 , x226 , x227 , x228 , x229 , x230 , x231 , x232 , x233 , x234 , x235 , x236 , x237 , x238 , x239 , x240 , x241 , x242 , x243 , x244 , x245 , x246 , x247 , x248 , x249 , x250 , x251 , x252 , x253 , x254 , x255 , x256 , x257 , x258 , x259 , x260 , x261 , x262 , x263 , x264 , x265 , x266 , x267 , x268 , x269 , x270 , x271 , x272 , x273 , x274 , x275 , x276 , x277 , x278 , x279 , x280 , x281 , x282 , x283 , x284 , x285 , x286 , x287 , x288 , x289 , x290 , x291 , x292 , x293 , x294 , x295 , x296 , x297 , x298 , x299 , x300 , x301 , x302 , x303 , x304 , x305 , x306 , x307 , x308 , x309 , x310 , x311 , x312 , x313 , x314 , x315 , x316 , x317 , x318 , x319 , x320 , x321 , x322 , x323 , x324 , x325 , x326 , x327 , x328 , x329 , x330 , x331 , x332 , x333 , x334 , x335 , x336 , x337 , x338 , x339 , x340 , x341 , x342 , x343 , x344 , x345 , x346 , x347 , x348 , x349 , x350 , x351 , x352 , x353 , x354 , x355 , x356 , x357 , x358 , x359 , x360 , x361 , x362 , x363 , x364 , x365 , x366 , x367 , x368 , x369 , x370 , x371 , x372 , x373 , x374 , x375 , x376 , x377 , x378 , x379 , x380 , x381 , x382 , x383 , x384 , x385 , x386 , x387 , x388 , x389 , x390 , x391 , x392 , x393 , x394 , x395 , x396 , x397 , x398 , x399 , x400 , x401 , x402 , x403 , x404 , x405 , x406 , x407 , x408 , x409 , x410 , x411 , x412 , x413 , x414 , x415 , x416 , x417 , x418 , x419 , x420 , x421 , x422 , x423 , x424 , x425 , x426 , x427 , x428 , x429 , x430 , x431 , x432 , x433 , x434 , x435 , x436 , x437 , x438 , x439 , x440 , x441 , x442 , x443 , x444 , x445 , x446 , x447 , x448 , x449 , x450 , x451 , x452 , x453 , x454 , x455 , x456 , x457 , x458 , x459 , x460 , x461 , x462 , x463 , x464 , x465 , x466 , x467 , x468 , x469 , x470 , x471 , x472 , x473 , x474 , x475 , x476 , x477 , x478 , x479 , x480 , x481 , x482 , x483 , x484 , x485 , x486 , x487 , x488 , x489 , x490 , x491 , x492 , x493 , x494 , x495 , x496 , x497 , x498 , x499 , x500 , x501 , x502 , x503 , x504 , x505 , x506 , x507 , x508 , x509 , x510 , x511 , x512 , x513 , x514 , x515 , x516 , x517 , x518 , x519 , x520 , x521 , x522 , x523 , x524 , x525 , x526 , x527 , x528 , x529 , x530 , x531 , x532 , x533 , x534 , x535 , x536 , x537 , x538 , x539 , x540 , x541 , x542 , x543 , x544 , x545 , x546 , x547 , x548 , x549 , x550 , x551 , x552 , x553 , x554 , x555 , x556 , x557 , x558 , x559 , x560 , x561 , x562 , x563 , x564 , x565 , x566 , x567 , x568 , x569 , x570 , x571 , x572 , x573 , x574 , x575 , x576 , x577 , x578 , x579 , x580 , x581 , x582 , x583 , x584 , x585 , x586 , x587 , x588 , x589 , x590 , x591 , x592 , x593 , x594 , x595 , x596 , x597 , x598 , x599 , x600 , x601 , x602 , x603 , x604 , x605 , x606 , x607 , x608 , x609 , x610 , x611 , x612 , x613 , x614 , x615 , x616 , x617 , x618 , x619 , x620 , x621 , x622 , x623 , x624 , x625 , x626 , x627 , x628 , x629 , x630 , x631 , x632 , x633 , x634 , x635 , x636 , x637 , x638 , x639 , x640 , x641 , x642 , x643 , x644 , x645 , x646 , x647 , x648 , x649 , x650 , x651 , x652 , x653 , x654 , x655 , x656 , x657 , x658 , x659 , x660 , x661 , x662 , x663 , x664 , x665 , x666 , x667 , x668 , x669 , x670 , x671 , x672 , x673 , x674 , x675 , x676 , x677 , x678 , x679 , x680 , x681 , x682 , x683 , x684 , x685 , x686 , x687 , x688 , x689 , x690 , x691 , x692 , x693 , x694 , x695 , x696 , x697 , x698 , x699 , x700 , x701 , x702 , x703 , x704 , x705 , x706 , x707 , x708 , x709 , x710 , x711 , x712 , x713 , x714 , x715 , x716 , x717 , x718 , x719 , x720 , x721 , x722 , x723 , x724 , x725 , x726 , x727 , x728 , x729 , x730 , x731 , x732 , x733 , x734 , x735 , x736 , x737 , x738 , x739 , x740 , x741 , x742 , x743 , x744 , x745 , x746 , x747 , x748 , x749 , x750 , x751 , x752 , x753 , x754 , x755 , x756 , x757 , x758 , x759 , x760 , x761 , x762 , x763 , x764 , x765 , x766 , x767 , x768 , x769 , x770 , x771 , x772 , x773 , x774 , x775 , x776 , x777 , x778 , x779 , x780 , x781 , x782 , x783 , x784 , x785 , x786 , x787 , x788 , x789 , x790 , x791 , x792 , x793 , x794 , x795 , x796 , x797 , x798 , x799 , x800 , x801 , x802 , x803 , x804 , x805 , x806 , x807 , x808 , x809 , x810 , x811 , x812 , x813 , x814 , x815 , x816 , x817 , x818 , x819 , x820 , x821 , x822 , x823 , x824 , x825 , x826 , x827 , x828 , x829 , x830 , x831 , x832 , x833 , x834 , x835 , x836 , x837 , x838 , x839 , x840 , x841 , x842 , x843 , x844 , x845 , x846 , x847 , x848 , x849 , x850 , x851 , x852 , x853 , x854 , x855 , x856 , x857 , x858 , x859 , x860 , x861 , x862 , x863 , x864 , x865 , x866 , x867 , x868 , x869 , x870 , x871 , x872 , x873 , x874 , x875 , x876 , x877 , x878 , x879 , x880 , x881 , x882 , x883 , x884 , x885 , x886 , x887 , x888 , x889 , x890 , x891 , x892 , x893 , x894 , x895 , x896 , x897 , x898 , x899 , x900 , x901 , x902 , x903 , x904 , x905 , x906 , x907 , x908 , x909 , x910 , x911 , x912 , x913 , x914 , x915 , x916 , x917 , x918 , x919 , x920 , x921 , x922 , x923 , x924 , x925 , x926 , x927 , x928 , x929 , x930 , x931 , x932 , x933 , x934 , x935 , x936 , x937 , x938 , x939 , x940 , x941 , x942 , x943 , x944 , x945 , x946 , x947 , x948 , x949 , x950 , x951 , x952 , x953 , x954 , x955 , x956 , x957 , x958 , x959 , x960 , x961 , x962 , x963 , x964 , x965 , x966 , x967 , x968 , x969 , x970 , x971 , x972 , x973 , x974 , x975 , x976 , x977 , x978 , x979 , x980 , x981 , x982 , x983 , x984 , x985 , x986 , x987 , x988 , x989 , x990 , x991 , x992 , x993 , x994 , x995 , x996 , x997 , x998 , x999 , x1000 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 , x147 , x148 , x149 , x150 , x151 , x152 , x153 , x154 , x155 , x156 , x157 , x158 , x159 , x160 , x161 , x162 , x163 , x164 , x165 , x166 , x167 , x168 , x169 , x170 , x171 , x172 , x173 , x174 , x175 , x176 , x177 , x178 , x179 , x180 , x181 , x182 , x183 , x184 , x185 , x186 , x187 , x188 , x189 , x190 , x191 , x192 , x193 , x194 , x195 , x196 , x197 , x198 , x199 , x200 , x201 , x202 , x203 , x204 , x205 , x206 , x207 , x208 , x209 , x210 , x211 , x212 , x213 , x214 , x215 , x216 , x217 , x218 , x219 , x220 , x221 , x222 , x223 , x224 , x225 , x226 , x227 , x228 , x229 , x230 , x231 , x232 , x233 , x234 , x235 , x236 , x237 , x238 , x239 , x240 , x241 , x242 , x243 , x244 , x245 , x246 , x247 , x248 , x249 , x250 , x251 , x252 , x253 , x254 , x255 , x256 , x257 , x258 , x259 , x260 , x261 , x262 , x263 , x264 , x265 , x266 , x267 , x268 , x269 , x270 , x271 , x272 , x273 , x274 , x275 , x276 , x277 , x278 , x279 , x280 , x281 , x282 , x283 , x284 , x285 , x286 , x287 , x288 , x289 , x290 , x291 , x292 , x293 , x294 , x295 , x296 , x297 , x298 , x299 , x300 , x301 , x302 , x303 , x304 , x305 , x306 , x307 , x308 , x309 , x310 , x311 , x312 , x313 , x314 , x315 , x316 , x317 , x318 , x319 , x320 , x321 , x322 , x323 , x324 , x325 , x326 , x327 , x328 , x329 , x330 , x331 , x332 , x333 , x334 , x335 , x336 , x337 , x338 , x339 , x340 , x341 , x342 , x343 , x344 , x345 , x346 , x347 , x348 , x349 , x350 , x351 , x352 , x353 , x354 , x355 , x356 , x357 , x358 , x359 , x360 , x361 , x362 , x363 , x364 , x365 , x366 , x367 , x368 , x369 , x370 , x371 , x372 , x373 , x374 , x375 , x376 , x377 , x378 , x379 , x380 , x381 , x382 , x383 , x384 , x385 , x386 , x387 , x388 , x389 , x390 , x391 , x392 , x393 , x394 , x395 , x396 , x397 , x398 , x399 , x400 , x401 , x402 , x403 , x404 , x405 , x406 , x407 , x408 , x409 , x410 , x411 , x412 , x413 , x414 , x415 , x416 , x417 , x418 , x419 , x420 , x421 , x422 , x423 , x424 , x425 , x426 , x427 , x428 , x429 , x430 , x431 , x432 , x433 , x434 , x435 , x436 , x437 , x438 , x439 , x440 , x441 , x442 , x443 , x444 , x445 , x446 , x447 , x448 , x449 , x450 , x451 , x452 , x453 , x454 , x455 , x456 , x457 , x458 , x459 , x460 , x461 , x462 , x463 , x464 , x465 , x466 , x467 , x468 , x469 , x470 , x471 , x472 , x473 , x474 , x475 , x476 , x477 , x478 , x479 , x480 , x481 , x482 , x483 , x484 , x485 , x486 , x487 , x488 , x489 , x490 , x491 , x492 , x493 , x494 , x495 , x496 , x497 , x498 , x499 , x500 , x501 , x502 , x503 , x504 , x505 , x506 , x507 , x508 , x509 , x510 , x511 , x512 , x513 , x514 , x515 , x516 , x517 , x518 , x519 , x520 , x521 , x522 , x523 , x524 , x525 , x526 , x527 , x528 , x529 , x530 , x531 , x532 , x533 , x534 , x535 , x536 , x537 , x538 , x539 , x540 , x541 , x542 , x543 , x544 , x545 , x546 , x547 , x548 , x549 , x550 , x551 , x552 , x553 , x554 , x555 , x556 , x557 , x558 , x559 , x560 , x561 , x562 , x563 , x564 , x565 , x566 , x567 , x568 , x569 , x570 , x571 , x572 , x573 , x574 , x575 , x576 , x577 , x578 , x579 , x580 , x581 , x582 , x583 , x584 , x585 , x586 , x587 , x588 , x589 , x590 , x591 , x592 , x593 , x594 , x595 , x596 , x597 , x598 , x599 , x600 , x601 , x602 , x603 , x604 , x605 , x606 , x607 , x608 , x609 , x610 , x611 , x612 , x613 , x614 , x615 , x616 , x617 , x618 , x619 , x620 , x621 , x622 , x623 , x624 , x625 , x626 , x627 , x628 , x629 , x630 , x631 , x632 , x633 , x634 , x635 , x636 , x637 , x638 , x639 , x640 , x641 , x642 , x643 , x644 , x645 , x646 , x647 , x648 , x649 , x650 , x651 , x652 , x653 , x654 , x655 , x656 , x657 , x658 , x659 , x660 , x661 , x662 , x663 , x664 , x665 , x666 , x667 , x668 , x669 , x670 , x671 , x672 , x673 , x674 , x675 , x676 , x677 , x678 , x679 , x680 , x681 , x682 , x683 , x684 , x685 , x686 , x687 , x688 , x689 , x690 , x691 , x692 , x693 , x694 , x695 , x696 , x697 , x698 , x699 , x700 , x701 , x702 , x703 , x704 , x705 , x706 , x707 , x708 , x709 , x710 , x711 , x712 , x713 , x714 , x715 , x716 , x717 , x718 , x719 , x720 , x721 , x722 , x723 , x724 , x725 , x726 , x727 , x728 , x729 , x730 , x731 , x732 , x733 , x734 , x735 , x736 , x737 , x738 , x739 , x740 , x741 , x742 , x743 , x744 , x745 , x746 , x747 , x748 , x749 , x750 , x751 , x752 , x753 , x754 , x755 , x756 , x757 , x758 , x759 , x760 , x761 , x762 , x763 , x764 , x765 , x766 , x767 , x768 , x769 , x770 , x771 , x772 , x773 , x774 , x775 , x776 , x777 , x778 , x779 , x780 , x781 , x782 , x783 , x784 , x785 , x786 , x787 , x788 , x789 , x790 , x791 , x792 , x793 , x794 , x795 , x796 , x797 , x798 , x799 , x800 , x801 , x802 , x803 , x804 , x805 , x806 , x807 , x808 , x809 , x810 , x811 , x812 , x813 , x814 , x815 , x816 , x817 , x818 , x819 , x820 , x821 , x822 , x823 , x824 , x825 , x826 , x827 , x828 , x829 , x830 , x831 , x832 , x833 , x834 , x835 , x836 , x837 , x838 , x839 , x840 , x841 , x842 , x843 , x844 , x845 , x846 , x847 , x848 , x849 , x850 , x851 , x852 , x853 , x854 , x855 , x856 , x857 , x858 , x859 , x860 , x861 , x862 , x863 , x864 , x865 , x866 , x867 , x868 , x869 , x870 , x871 , x872 , x873 , x874 , x875 , x876 , x877 , x878 , x879 , x880 , x881 , x882 , x883 , x884 , x885 , x886 , x887 , x888 , x889 , x890 , x891 , x892 , x893 , x894 , x895 , x896 , x897 , x898 , x899 , x900 , x901 , x902 , x903 , x904 , x905 , x906 , x907 , x908 , x909 , x910 , x911 , x912 , x913 , x914 , x915 , x916 , x917 , x918 , x919 , x920 , x921 , x922 , x923 , x924 , x925 , x926 , x927 , x928 , x929 , x930 , x931 , x932 , x933 , x934 , x935 , x936 , x937 , x938 , x939 , x940 , x941 , x942 , x943 , x944 , x945 , x946 , x947 , x948 , x949 , x950 , x951 , x952 , x953 , x954 , x955 , x956 , x957 , x958 , x959 , x960 , x961 , x962 , x963 , x964 , x965 , x966 , x967 , x968 , x969 , x970 , x971 , x972 , x973 , x974 , x975 , x976 , x977 , x978 , x979 , x980 , x981 , x982 , x983 , x984 , x985 , x986 , x987 , x988 , x989 , x990 , x991 , x992 , x993 , x994 , x995 , x996 , x997 , x998 , x999 , x1000 ;
  output y0 ;
  wire n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , n3931 , n3932 , n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , n3940 , n3941 , n3942 , n3943 , n3944 , n3945 , n3946 , n3947 , n3948 , n3949 , n3950 , n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , n3970 , n3971 , n3972 , n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , n3980 , n3981 , n3982 , n3983 , n3984 , n3985 , n3986 , n3987 , n3988 , n3989 , n3990 , n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , n4000 , n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , n4009 , n4010 , n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , n4019 , n4020 , n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , n4029 , n4030 , n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , n4039 , n4040 , n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4049 , n4050 , n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , n4059 , n4060 , n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , n4070 , n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , n4079 , n4080 , n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , n4089 , n4090 , n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , n4097 , n4098 , n4099 , n4100 , n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , n4109 , n4110 , n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , n4119 , n4120 , n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , n4129 , n4130 , n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , n4139 , n4140 , n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , n4150 , n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , n4159 , n4160 , n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , n4169 , n4170 , n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , n4179 , n4180 , n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , n4189 , n4190 , n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , n4197 , n4198 , n4199 , n4200 , n4201 , n4202 , n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , n4209 , n4210 , n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , n4217 , n4218 , n4219 , n4220 , n4221 , n4222 , n4223 , n4224 , n4225 , n4226 , n4227 , n4228 , n4229 , n4230 , n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , n4237 , n4238 , n4239 , n4240 , n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , n4247 , n4248 , n4249 , n4250 , n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , n4259 , n4260 , n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , n4269 , n4270 , n4271 , n4272 , n4273 , n4274 , n4275 , n4276 , n4277 , n4278 , n4279 , n4280 , n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , n4289 , n4290 , n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , n4299 , n4300 , n4301 , n4302 , n4303 , n4304 , n4305 , n4306 , n4307 , n4308 , n4309 , n4310 , n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , n4319 , n4320 , n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , n4329 , n4330 , n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , n4340 , n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , n4349 , n4350 , n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , n4360 , n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , n4370 , n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , n4380 , n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , n4390 , n4391 , n4392 , n4393 , n4394 , n4395 , n4396 , n4397 , n4398 , n4399 , n4400 , n4401 , n4402 , n4403 , n4404 , n4405 , n4406 , n4407 , n4408 , n4409 , n4410 , n4411 , n4412 , n4413 , n4414 , n4415 , n4416 , n4417 , n4418 , n4419 , n4420 , n4421 , n4422 , n4423 , n4424 , n4425 , n4426 , n4427 , n4428 , n4429 , n4430 , n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , n4437 , n4438 , n4439 , n4440 , n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , n4449 , n4450 , n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , n4459 , n4460 , n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , n4469 , n4470 , n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , n4479 , n4480 , n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , n4487 , n4488 , n4489 , n4490 , n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , n4497 , n4498 , n4499 , n4500 , n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , n4509 , n4510 , n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , n4519 , n4520 , n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , n4529 , n4530 , n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , n4537 , n4538 , n4539 , n4540 , n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , n4547 , n4548 , n4549 , n4550 , n4551 , n4552 , n4553 , n4554 , n4555 , n4556 , n4557 , n4558 , n4559 , n4560 , n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , n4567 , n4568 , n4569 , n4570 , n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , n4579 , n4580 , n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , n4589 , n4590 , n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , n4597 , n4598 , n4599 , n4600 , n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , n4607 , n4608 , n4609 , n4610 , n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , n4617 , n4618 , n4619 , n4620 , n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , n4627 , n4628 , n4629 , n4630 , n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , n4637 , n4638 , n4639 , n4640 , n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , n4647 , n4648 , n4649 , n4650 , n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , n4657 , n4658 , n4659 , n4660 , n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , n4669 , n4670 , n4671 , n4672 , n4673 , n4674 , n4675 , n4676 , n4677 , n4678 , n4679 , n4680 , n4681 , n4682 , n4683 , n4684 , n4685 , n4686 , n4687 , n4688 , n4689 , n4690 , n4691 , n4692 , n4693 , n4694 , n4695 , n4696 , n4697 , n4698 , n4699 , n4700 , n4701 , n4702 , n4703 , n4704 , n4705 , n4706 , n4707 , n4708 , n4709 , n4710 , n4711 , n4712 , n4713 , n4714 , n4715 , n4716 , n4717 , n4718 , n4719 , n4720 , n4721 , n4722 , n4723 , n4724 , n4725 , n4726 , n4727 , n4728 , n4729 , n4730 , n4731 , n4732 , n4733 , n4734 , n4735 , n4736 , n4737 , n4738 , n4739 , n4740 , n4741 , n4742 , n4743 , n4744 , n4745 , n4746 , n4747 , n4748 , n4749 , n4750 , n4751 , n4752 , n4753 , n4754 , n4755 , n4756 , n4757 , n4758 , n4759 , n4760 , n4761 , n4762 , n4763 , n4764 , n4765 , n4766 , n4767 , n4768 , n4769 , n4770 , n4771 , n4772 , n4773 , n4774 , n4775 , n4776 , n4777 , n4778 , n4779 , n4780 , n4781 , n4782 , n4783 , n4784 , n4785 , n4786 , n4787 , n4788 , n4789 , n4790 , n4791 , n4792 , n4793 , n4794 , n4795 , n4796 , n4797 , n4798 , n4799 , n4800 , n4801 , n4802 , n4803 , n4804 , n4805 , n4806 , n4807 , n4808 , n4809 , n4810 , n4811 , n4812 , n4813 , n4814 , n4815 , n4816 , n4817 , n4818 , n4819 , n4820 , n4821 , n4822 , n4823 , n4824 , n4825 , n4826 , n4827 , n4828 , n4829 , n4830 , n4831 , n4832 , n4833 , n4834 , n4835 , n4836 , n4837 , n4838 , n4839 , n4840 , n4841 , n4842 , n4843 , n4844 , n4845 , n4846 , n4847 , n4848 , n4849 , n4850 , n4851 , n4852 , n4853 , n4854 , n4855 , n4856 , n4857 , n4858 , n4859 , n4860 , n4861 , n4862 , n4863 , n4864 , n4865 , n4866 , n4867 , n4868 , n4869 , n4870 , n4871 , n4872 , n4873 , n4874 , n4875 , n4876 , n4877 , n4878 , n4879 , n4880 , n4881 , n4882 , n4883 , n4884 , n4885 , n4886 , n4887 , n4888 , n4889 , n4890 , n4891 , n4892 , n4893 , n4894 , n4895 , n4896 , n4897 , n4898 , n4899 , n4900 , n4901 , n4902 , n4903 , n4904 , n4905 , n4906 , n4907 , n4908 , n4909 , n4910 , n4911 , n4912 , n4913 , n4914 , n4915 , n4916 , n4917 , n4918 , n4919 , n4920 , n4921 , n4922 , n4923 , n4924 , n4925 , n4926 , n4927 , n4928 , n4929 , n4930 , n4931 , n4932 , n4933 , n4934 , n4935 , n4936 , n4937 , n4938 , n4939 , n4940 , n4941 , n4942 , n4943 , n4944 , n4945 , n4946 , n4947 , n4948 , n4949 , n4950 , n4951 , n4952 , n4953 , n4954 , n4955 , n4956 , n4957 , n4958 , n4959 , n4960 , n4961 , n4962 , n4963 , n4964 , n4965 , n4966 , n4967 , n4968 , n4969 , n4970 , n4971 , n4972 , n4973 , n4974 , n4975 , n4976 , n4977 , n4978 , n4979 , n4980 , n4981 , n4982 , n4983 , n4984 , n4985 , n4986 , n4987 , n4988 , n4989 , n4990 , n4991 , n4992 , n4993 , n4994 , n4995 , n4996 , n4997 , n4998 , n4999 , n5000 , n5001 , n5002 , n5003 , n5004 , n5005 , n5006 , n5007 , n5008 , n5009 , n5010 , n5011 , n5012 , n5013 , n5014 , n5015 , n5016 , n5017 , n5018 , n5019 , n5020 , n5021 , n5022 , n5023 , n5024 , n5025 , n5026 , n5027 , n5028 , n5029 , n5030 , n5031 , n5032 , n5033 , n5034 , n5035 , n5036 , n5037 , n5038 , n5039 , n5040 , n5041 , n5042 , n5043 , n5044 , n5045 , n5046 , n5047 , n5048 , n5049 , n5050 , n5051 , n5052 , n5053 , n5054 , n5055 , n5056 , n5057 , n5058 , n5059 , n5060 , n5061 , n5062 , n5063 , n5064 , n5065 , n5066 , n5067 , n5068 , n5069 , n5070 , n5071 , n5072 , n5073 , n5074 , n5075 , n5076 , n5077 , n5078 , n5079 , n5080 , n5081 , n5082 , n5083 , n5084 , n5085 , n5086 , n5087 , n5088 , n5089 , n5090 , n5091 , n5092 , n5093 , n5094 , n5095 , n5096 , n5097 , n5098 , n5099 , n5100 , n5101 , n5102 , n5103 , n5104 , n5105 , n5106 , n5107 , n5108 , n5109 , n5110 , n5111 , n5112 , n5113 , n5114 , n5115 , n5116 , n5117 , n5118 , n5119 , n5120 , n5121 , n5122 , n5123 , n5124 , n5125 , n5126 , n5127 , n5128 , n5129 , n5130 , n5131 , n5132 , n5133 , n5134 , n5135 , n5136 , n5137 , n5138 , n5139 , n5140 , n5141 , n5142 , n5143 , n5144 , n5145 , n5146 , n5147 , n5148 , n5149 , n5150 , n5151 , n5152 , n5153 , n5154 , n5155 , n5156 , n5157 , n5158 , n5159 , n5160 , n5161 , n5162 , n5163 , n5164 , n5165 , n5166 , n5167 , n5168 , n5169 , n5170 , n5171 , n5172 , n5173 , n5174 , n5175 , n5176 , n5177 , n5178 , n5179 , n5180 , n5181 , n5182 , n5183 , n5184 , n5185 , n5186 , n5187 , n5188 , n5189 , n5190 , n5191 , n5192 , n5193 , n5194 , n5195 , n5196 , n5197 , n5198 , n5199 , n5200 , n5201 , n5202 , n5203 , n5204 , n5205 , n5206 , n5207 , n5208 , n5209 , n5210 , n5211 , n5212 , n5213 , n5214 , n5215 , n5216 , n5217 , n5218 , n5219 , n5220 , n5221 , n5222 , n5223 , n5224 , n5225 , n5226 , n5227 , n5228 , n5229 , n5230 , n5231 , n5232 , n5233 , n5234 , n5235 , n5236 , n5237 , n5238 , n5239 , n5240 , n5241 , n5242 , n5243 , n5244 , n5245 , n5246 , n5247 , n5248 , n5249 , n5250 , n5251 , n5252 , n5253 , n5254 , n5255 , n5256 , n5257 , n5258 , n5259 , n5260 , n5261 , n5262 , n5263 , n5264 , n5265 , n5266 , n5267 , n5268 , n5269 , n5270 , n5271 , n5272 , n5273 , n5274 , n5275 , n5276 , n5277 , n5278 , n5279 , n5280 , n5281 , n5282 , n5283 , n5284 , n5285 , n5286 , n5287 , n5288 , n5289 , n5290 , n5291 , n5292 , n5293 , n5294 , n5295 , n5296 , n5297 , n5298 , n5299 , n5300 , n5301 , n5302 , n5303 , n5304 , n5305 , n5306 , n5307 , n5308 , n5309 , n5310 , n5311 , n5312 , n5313 , n5314 , n5315 , n5316 , n5317 , n5318 , n5319 , n5320 , n5321 , n5322 , n5323 , n5324 , n5325 , n5326 , n5327 , n5328 , n5329 , n5330 , n5331 , n5332 , n5333 , n5334 , n5335 , n5336 , n5337 , n5338 , n5339 , n5340 , n5341 , n5342 , n5343 , n5344 , n5345 , n5346 , n5347 , n5348 , n5349 , n5350 , n5351 , n5352 , n5353 , n5354 , n5355 , n5356 , n5357 , n5358 , n5359 , n5360 , n5361 , n5362 , n5363 , n5364 , n5365 , n5366 , n5367 , n5368 , n5369 , n5370 , n5371 , n5372 , n5373 , n5374 , n5375 , n5376 , n5377 , n5378 , n5379 , n5380 , n5381 , n5382 , n5383 , n5384 , n5385 , n5386 , n5387 , n5388 , n5389 , n5390 , n5391 , n5392 , n5393 , n5394 , n5395 , n5396 , n5397 , n5398 , n5399 , n5400 , n5401 , n5402 , n5403 , n5404 , n5405 , n5406 , n5407 , n5408 , n5409 , n5410 , n5411 , n5412 , n5413 , n5414 , n5415 , n5416 , n5417 , n5418 , n5419 , n5420 , n5421 , n5422 , n5423 , n5424 , n5425 , n5426 , n5427 , n5428 , n5429 , n5430 , n5431 , n5432 , n5433 , n5434 , n5435 , n5436 , n5437 , n5438 , n5439 , n5440 , n5441 , n5442 , n5443 , n5444 , n5445 , n5446 , n5447 , n5448 , n5449 , n5450 , n5451 , n5452 , n5453 , n5454 , n5455 , n5456 , n5457 , n5458 , n5459 , n5460 , n5461 , n5462 , n5463 , n5464 , n5465 , n5466 , n5467 , n5468 , n5469 , n5470 , n5471 , n5472 , n5473 , n5474 , n5475 , n5476 , n5477 , n5478 , n5479 , n5480 , n5481 , n5482 , n5483 , n5484 , n5485 , n5486 , n5487 , n5488 , n5489 , n5490 , n5491 , n5492 , n5493 , n5494 , n5495 , n5496 , n5497 , n5498 , n5499 , n5500 , n5501 , n5502 , n5503 , n5504 , n5505 , n5506 , n5507 , n5508 , n5509 , n5510 , n5511 , n5512 , n5513 , n5514 , n5515 , n5516 , n5517 , n5518 , n5519 , n5520 , n5521 , n5522 , n5523 , n5524 , n5525 , n5526 , n5527 , n5528 , n5529 , n5530 , n5531 , n5532 , n5533 , n5534 , n5535 , n5536 , n5537 , n5538 , n5539 , n5540 , n5541 , n5542 , n5543 , n5544 , n5545 , n5546 , n5547 , n5548 , n5549 , n5550 , n5551 , n5552 , n5553 , n5554 , n5555 , n5556 , n5557 , n5558 , n5559 , n5560 , n5561 , n5562 , n5563 , n5564 , n5565 , n5566 , n5567 , n5568 , n5569 , n5570 , n5571 , n5572 , n5573 , n5574 , n5575 , n5576 , n5577 , n5578 , n5579 , n5580 , n5581 , n5582 , n5583 , n5584 , n5585 , n5586 , n5587 , n5588 , n5589 , n5590 , n5591 , n5592 , n5593 , n5594 , n5595 , n5596 , n5597 , n5598 , n5599 , n5600 , n5601 , n5602 , n5603 , n5604 , n5605 , n5606 , n5607 , n5608 , n5609 , n5610 , n5611 , n5612 , n5613 , n5614 , n5615 , n5616 , n5617 , n5618 , n5619 , n5620 , n5621 , n5622 , n5623 , n5624 , n5625 , n5626 , n5627 , n5628 , n5629 , n5630 , n5631 , n5632 , n5633 , n5634 , n5635 , n5636 , n5637 , n5638 , n5639 , n5640 , n5641 , n5642 , n5643 , n5644 , n5645 , n5646 , n5647 , n5648 , n5649 , n5650 , n5651 , n5652 , n5653 , n5654 , n5655 , n5656 , n5657 , n5658 , n5659 , n5660 , n5661 , n5662 , n5663 , n5664 , n5665 , n5666 , n5667 , n5668 , n5669 , n5670 , n5671 , n5672 , n5673 , n5674 , n5675 , n5676 , n5677 , n5678 , n5679 , n5680 , n5681 , n5682 , n5683 , n5684 , n5685 , n5686 , n5687 , n5688 , n5689 , n5690 , n5691 , n5692 , n5693 , n5694 , n5695 , n5696 , n5697 , n5698 , n5699 , n5700 , n5701 , n5702 , n5703 , n5704 , n5705 , n5706 , n5707 , n5708 , n5709 , n5710 , n5711 , n5712 , n5713 , n5714 , n5715 , n5716 , n5717 , n5718 , n5719 , n5720 , n5721 , n5722 , n5723 , n5724 , n5725 , n5726 , n5727 , n5728 , n5729 , n5730 , n5731 , n5732 , n5733 , n5734 , n5735 , n5736 , n5737 , n5738 , n5739 , n5740 , n5741 , n5742 , n5743 , n5744 , n5745 , n5746 , n5747 , n5748 , n5749 , n5750 , n5751 , n5752 , n5753 , n5754 , n5755 , n5756 , n5757 , n5758 , n5759 , n5760 , n5761 , n5762 , n5763 , n5764 , n5765 , n5766 , n5767 , n5768 , n5769 , n5770 , n5771 , n5772 , n5773 , n5774 , n5775 , n5776 , n5777 , n5778 , n5779 , n5780 , n5781 , n5782 , n5783 , n5784 , n5785 , n5786 , n5787 , n5788 , n5789 , n5790 , n5791 , n5792 , n5793 , n5794 , n5795 , n5796 , n5797 , n5798 , n5799 , n5800 , n5801 , n5802 , n5803 , n5804 , n5805 , n5806 , n5807 , n5808 , n5809 , n5810 , n5811 , n5812 , n5813 , n5814 , n5815 , n5816 , n5817 , n5818 , n5819 , n5820 , n5821 , n5822 , n5823 , n5824 , n5825 , n5826 , n5827 , n5828 , n5829 , n5830 , n5831 , n5832 , n5833 , n5834 , n5835 , n5836 , n5837 , n5838 , n5839 , n5840 , n5841 , n5842 , n5843 , n5844 , n5845 , n5846 , n5847 , n5848 , n5849 , n5850 , n5851 , n5852 , n5853 , n5854 , n5855 , n5856 , n5857 , n5858 , n5859 , n5860 , n5861 , n5862 , n5863 , n5864 , n5865 , n5866 , n5867 , n5868 , n5869 , n5870 , n5871 , n5872 , n5873 , n5874 , n5875 , n5876 , n5877 , n5878 , n5879 , n5880 , n5881 , n5882 , n5883 , n5884 , n5885 , n5886 , n5887 , n5888 , n5889 , n5890 , n5891 , n5892 , n5893 , n5894 , n5895 , n5896 , n5897 , n5898 , n5899 , n5900 , n5901 , n5902 , n5903 , n5904 , n5905 , n5906 , n5907 , n5908 , n5909 , n5910 , n5911 , n5912 , n5913 , n5914 , n5915 , n5916 , n5917 , n5918 , n5919 , n5920 , n5921 , n5922 , n5923 , n5924 , n5925 , n5926 , n5927 , n5928 , n5929 , n5930 , n5931 , n5932 , n5933 , n5934 , n5935 , n5936 , n5937 , n5938 , n5939 , n5940 , n5941 , n5942 , n5943 , n5944 , n5945 , n5946 , n5947 , n5948 , n5949 , n5950 , n5951 , n5952 , n5953 , n5954 , n5955 , n5956 , n5957 , n5958 , n5959 , n5960 , n5961 , n5962 , n5963 , n5964 , n5965 , n5966 , n5967 , n5968 , n5969 , n5970 , n5971 , n5972 , n5973 , n5974 , n5975 , n5976 , n5977 , n5978 , n5979 , n5980 , n5981 , n5982 , n5983 , n5984 , n5985 , n5986 , n5987 , n5988 , n5989 , n5990 , n5991 , n5992 , n5993 , n5994 , n5995 , n5996 , n5997 , n5998 , n5999 , n6000 , n6001 , n6002 , n6003 , n6004 , n6005 , n6006 , n6007 , n6008 , n6009 , n6010 , n6011 , n6012 , n6013 , n6014 , n6015 , n6016 , n6017 , n6018 , n6019 , n6020 , n6021 , n6022 , n6023 , n6024 , n6025 , n6026 , n6027 , n6028 , n6029 , n6030 , n6031 , n6032 , n6033 , n6034 , n6035 , n6036 , n6037 , n6038 , n6039 , n6040 , n6041 , n6042 , n6043 , n6044 , n6045 , n6046 , n6047 , n6048 , n6049 , n6050 , n6051 , n6052 , n6053 , n6054 , n6055 , n6056 , n6057 , n6058 , n6059 , n6060 , n6061 , n6062 , n6063 , n6064 , n6065 , n6066 , n6067 , n6068 , n6069 , n6070 , n6071 , n6072 , n6073 , n6074 , n6075 , n6076 , n6077 , n6078 , n6079 , n6080 , n6081 , n6082 , n6083 , n6084 , n6085 , n6086 , n6087 , n6088 , n6089 , n6090 , n6091 , n6092 , n6093 , n6094 , n6095 , n6096 , n6097 , n6098 , n6099 , n6100 , n6101 , n6102 , n6103 , n6104 , n6105 , n6106 , n6107 , n6108 , n6109 , n6110 , n6111 , n6112 , n6113 , n6114 , n6115 , n6116 , n6117 , n6118 , n6119 , n6120 , n6121 , n6122 , n6123 , n6124 , n6125 , n6126 , n6127 , n6128 , n6129 , n6130 , n6131 , n6132 , n6133 , n6134 , n6135 , n6136 , n6137 , n6138 , n6139 , n6140 , n6141 , n6142 , n6143 , n6144 , n6145 , n6146 , n6147 , n6148 , n6149 , n6150 , n6151 , n6152 , n6153 , n6154 , n6155 , n6156 , n6157 , n6158 , n6159 , n6160 , n6161 , n6162 , n6163 , n6164 , n6165 , n6166 , n6167 , n6168 , n6169 , n6170 , n6171 , n6172 , n6173 , n6174 , n6175 , n6176 , n6177 , n6178 , n6179 , n6180 , n6181 , n6182 , n6183 , n6184 , n6185 , n6186 , n6187 , n6188 , n6189 , n6190 , n6191 , n6192 , n6193 , n6194 , n6195 , n6196 , n6197 , n6198 , n6199 , n6200 , n6201 , n6202 , n6203 , n6204 , n6205 , n6206 , n6207 , n6208 , n6209 , n6210 , n6211 , n6212 , n6213 , n6214 , n6215 , n6216 , n6217 , n6218 , n6219 , n6220 , n6221 , n6222 , n6223 , n6224 , n6225 , n6226 , n6227 , n6228 , n6229 , n6230 , n6231 , n6232 , n6233 , n6234 , n6235 , n6236 , n6237 , n6238 , n6239 , n6240 , n6241 , n6242 , n6243 , n6244 , n6245 , n6246 , n6247 , n6248 , n6249 , n6250 , n6251 , n6252 , n6253 , n6254 , n6255 , n6256 , n6257 , n6258 , n6259 , n6260 , n6261 , n6262 , n6263 , n6264 , n6265 , n6266 , n6267 , n6268 , n6269 , n6270 , n6271 , n6272 , n6273 , n6274 , n6275 , n6276 , n6277 , n6278 , n6279 , n6280 , n6281 , n6282 , n6283 , n6284 , n6285 , n6286 , n6287 , n6288 , n6289 , n6290 , n6291 , n6292 , n6293 , n6294 , n6295 , n6296 , n6297 , n6298 , n6299 , n6300 , n6301 , n6302 , n6303 , n6304 , n6305 , n6306 , n6307 , n6308 , n6309 , n6310 , n6311 , n6312 , n6313 , n6314 , n6315 , n6316 , n6317 , n6318 , n6319 , n6320 , n6321 , n6322 , n6323 , n6324 , n6325 , n6326 , n6327 , n6328 , n6329 , n6330 , n6331 , n6332 , n6333 , n6334 , n6335 , n6336 , n6337 , n6338 , n6339 , n6340 , n6341 , n6342 , n6343 , n6344 , n6345 , n6346 , n6347 , n6348 , n6349 , n6350 , n6351 , n6352 , n6353 , n6354 , n6355 , n6356 , n6357 , n6358 , n6359 , n6360 , n6361 , n6362 , n6363 , n6364 , n6365 , n6366 , n6367 , n6368 , n6369 , n6370 , n6371 , n6372 , n6373 , n6374 , n6375 , n6376 , n6377 , n6378 , n6379 , n6380 , n6381 , n6382 , n6383 , n6384 , n6385 , n6386 , n6387 , n6388 , n6389 , n6390 , n6391 , n6392 , n6393 , n6394 , n6395 , n6396 , n6397 , n6398 , n6399 , n6400 , n6401 , n6402 , n6403 , n6404 , n6405 , n6406 , n6407 , n6408 , n6409 , n6410 , n6411 , n6412 , n6413 , n6414 , n6415 , n6416 , n6417 , n6418 , n6419 , n6420 , n6421 , n6422 , n6423 , n6424 , n6425 , n6426 , n6427 , n6428 , n6429 , n6430 , n6431 , n6432 , n6433 , n6434 , n6435 , n6436 , n6437 , n6438 , n6439 , n6440 , n6441 , n6442 , n6443 , n6444 , n6445 , n6446 , n6447 , n6448 , n6449 , n6450 , n6451 , n6452 , n6453 , n6454 , n6455 , n6456 , n6457 , n6458 , n6459 , n6460 , n6461 , n6462 , n6463 , n6464 , n6465 , n6466 , n6467 , n6468 , n6469 , n6470 , n6471 , n6472 , n6473 , n6474 , n6475 , n6476 , n6477 , n6478 , n6479 , n6480 , n6481 , n6482 , n6483 , n6484 , n6485 , n6486 , n6487 , n6488 , n6489 , n6490 , n6491 , n6492 , n6493 , n6494 , n6495 , n6496 , n6497 , n6498 , n6499 , n6500 , n6501 , n6502 , n6503 , n6504 , n6505 , n6506 , n6507 , n6508 , n6509 , n6510 , n6511 , n6512 , n6513 , n6514 , n6515 , n6516 , n6517 , n6518 , n6519 , n6520 , n6521 , n6522 , n6523 , n6524 , n6525 , n6526 , n6527 , n6528 , n6529 , n6530 , n6531 , n6532 , n6533 , n6534 , n6535 , n6536 , n6537 , n6538 , n6539 , n6540 , n6541 , n6542 , n6543 , n6544 , n6545 , n6546 , n6547 , n6548 , n6549 , n6550 , n6551 , n6552 , n6553 , n6554 , n6555 , n6556 , n6557 , n6558 , n6559 , n6560 , n6561 , n6562 , n6563 , n6564 , n6565 , n6566 , n6567 , n6568 , n6569 , n6570 , n6571 , n6572 , n6573 , n6574 , n6575 , n6576 , n6577 , n6578 , n6579 , n6580 , n6581 , n6582 , n6583 , n6584 , n6585 , n6586 , n6587 , n6588 , n6589 , n6590 , n6591 , n6592 , n6593 , n6594 , n6595 , n6596 , n6597 , n6598 , n6599 , n6600 , n6601 , n6602 , n6603 , n6604 , n6605 , n6606 , n6607 , n6608 , n6609 , n6610 , n6611 , n6612 , n6613 , n6614 , n6615 , n6616 , n6617 , n6618 , n6619 , n6620 , n6621 , n6622 , n6623 , n6624 , n6625 , n6626 , n6627 , n6628 , n6629 , n6630 , n6631 , n6632 , n6633 , n6634 , n6635 , n6636 , n6637 , n6638 , n6639 , n6640 , n6641 , n6642 , n6643 , n6644 , n6645 , n6646 , n6647 , n6648 , n6649 , n6650 , n6651 , n6652 , n6653 , n6654 , n6655 , n6656 , n6657 , n6658 , n6659 , n6660 , n6661 , n6662 , n6663 , n6664 , n6665 , n6666 , n6667 , n6668 , n6669 , n6670 , n6671 , n6672 , n6673 , n6674 , n6675 , n6676 , n6677 , n6678 , n6679 , n6680 , n6681 , n6682 , n6683 , n6684 , n6685 , n6686 , n6687 , n6688 , n6689 , n6690 , n6691 , n6692 , n6693 , n6694 , n6695 , n6696 , n6697 , n6698 , n6699 , n6700 , n6701 , n6702 , n6703 , n6704 , n6705 , n6706 , n6707 , n6708 , n6709 , n6710 , n6711 , n6712 , n6713 , n6714 , n6715 , n6716 , n6717 , n6718 , n6719 , n6720 , n6721 , n6722 , n6723 , n6724 , n6725 , n6726 , n6727 , n6728 , n6729 , n6730 , n6731 , n6732 , n6733 , n6734 , n6735 , n6736 , n6737 , n6738 , n6739 , n6740 , n6741 , n6742 , n6743 , n6744 , n6745 , n6746 , n6747 , n6748 , n6749 , n6750 , n6751 , n6752 , n6753 , n6754 , n6755 , n6756 , n6757 , n6758 , n6759 , n6760 , n6761 , n6762 , n6763 , n6764 , n6765 , n6766 , n6767 , n6768 , n6769 , n6770 , n6771 , n6772 , n6773 , n6774 , n6775 , n6776 , n6777 , n6778 , n6779 , n6780 , n6781 , n6782 , n6783 , n6784 , n6785 , n6786 , n6787 , n6788 , n6789 , n6790 , n6791 , n6792 , n6793 , n6794 , n6795 , n6796 , n6797 , n6798 , n6799 , n6800 , n6801 , n6802 , n6803 , n6804 , n6805 , n6806 , n6807 , n6808 , n6809 , n6810 , n6811 , n6812 , n6813 , n6814 , n6815 , n6816 , n6817 , n6818 , n6819 , n6820 , n6821 , n6822 , n6823 , n6824 , n6825 , n6826 , n6827 , n6828 , n6829 , n6830 , n6831 , n6832 , n6833 , n6834 , n6835 , n6836 , n6837 , n6838 , n6839 , n6840 , n6841 , n6842 , n6843 , n6844 , n6845 , n6846 , n6847 , n6848 , n6849 , n6850 , n6851 , n6852 , n6853 , n6854 , n6855 , n6856 , n6857 , n6858 , n6859 , n6860 , n6861 , n6862 , n6863 , n6864 , n6865 , n6866 , n6867 , n6868 , n6869 , n6870 , n6871 , n6872 , n6873 , n6874 , n6875 , n6876 , n6877 , n6878 , n6879 , n6880 , n6881 , n6882 , n6883 , n6884 , n6885 , n6886 , n6887 , n6888 , n6889 , n6890 , n6891 , n6892 , n6893 , n6894 , n6895 , n6896 , n6897 , n6898 , n6899 , n6900 , n6901 , n6902 , n6903 , n6904 , n6905 , n6906 , n6907 , n6908 , n6909 , n6910 , n6911 , n6912 , n6913 , n6914 , n6915 , n6916 , n6917 , n6918 , n6919 , n6920 , n6921 , n6922 , n6923 , n6924 , n6925 , n6926 , n6927 , n6928 , n6929 , n6930 , n6931 , n6932 , n6933 , n6934 , n6935 , n6936 , n6937 , n6938 , n6939 , n6940 , n6941 , n6942 , n6943 , n6944 , n6945 , n6946 , n6947 , n6948 , n6949 , n6950 , n6951 , n6952 , n6953 , n6954 , n6955 , n6956 , n6957 , n6958 , n6959 , n6960 , n6961 , n6962 , n6963 , n6964 , n6965 , n6966 , n6967 , n6968 , n6969 , n6970 , n6971 , n6972 , n6973 , n6974 , n6975 , n6976 , n6977 , n6978 , n6979 , n6980 , n6981 , n6982 , n6983 , n6984 , n6985 , n6986 , n6987 , n6988 , n6989 , n6990 , n6991 , n6992 , n6993 , n6994 , n6995 , n6996 , n6997 , n6998 , n6999 , n7000 , n7001 , n7002 , n7003 , n7004 , n7005 , n7006 , n7007 , n7008 , n7009 , n7010 , n7011 , n7012 , n7013 , n7014 , n7015 , n7016 , n7017 , n7018 , n7019 , n7020 , n7021 , n7022 , n7023 , n7024 , n7025 , n7026 , n7027 , n7028 , n7029 , n7030 , n7031 , n7032 , n7033 , n7034 , n7035 , n7036 , n7037 , n7038 , n7039 , n7040 , n7041 , n7042 , n7043 , n7044 , n7045 , n7046 , n7047 , n7048 , n7049 , n7050 , n7051 , n7052 , n7053 , n7054 , n7055 , n7056 , n7057 , n7058 , n7059 , n7060 , n7061 , n7062 , n7063 , n7064 , n7065 , n7066 , n7067 , n7068 , n7069 , n7070 , n7071 , n7072 , n7073 , n7074 , n7075 , n7076 , n7077 , n7078 , n7079 , n7080 , n7081 , n7082 , n7083 , n7084 , n7085 , n7086 , n7087 , n7088 , n7089 , n7090 , n7091 , n7092 , n7093 , n7094 , n7095 , n7096 , n7097 , n7098 , n7099 , n7100 , n7101 , n7102 , n7103 , n7104 , n7105 , n7106 , n7107 , n7108 , n7109 , n7110 , n7111 , n7112 , n7113 , n7114 , n7115 , n7116 , n7117 , n7118 , n7119 , n7120 , n7121 , n7122 , n7123 , n7124 , n7125 , n7126 , n7127 , n7128 , n7129 , n7130 , n7131 , n7132 , n7133 , n7134 , n7135 , n7136 , n7137 , n7138 , n7139 , n7140 , n7141 , n7142 , n7143 , n7144 , n7145 , n7146 , n7147 , n7148 , n7149 , n7150 , n7151 , n7152 , n7153 , n7154 , n7155 , n7156 , n7157 , n7158 , n7159 , n7160 , n7161 , n7162 , n7163 , n7164 , n7165 , n7166 , n7167 , n7168 , n7169 , n7170 , n7171 , n7172 , n7173 , n7174 , n7175 , n7176 , n7177 , n7178 , n7179 , n7180 , n7181 , n7182 , n7183 , n7184 , n7185 , n7186 , n7187 , n7188 , n7189 , n7190 , n7191 , n7192 , n7193 , n7194 , n7195 , n7196 , n7197 , n7198 , n7199 , n7200 , n7201 , n7202 , n7203 , n7204 , n7205 , n7206 , n7207 , n7208 , n7209 , n7210 , n7211 , n7212 , n7213 , n7214 , n7215 , n7216 , n7217 , n7218 , n7219 , n7220 , n7221 , n7222 , n7223 , n7224 , n7225 , n7226 , n7227 , n7228 , n7229 , n7230 , n7231 , n7232 , n7233 , n7234 , n7235 , n7236 , n7237 , n7238 , n7239 , n7240 , n7241 , n7242 , n7243 , n7244 , n7245 , n7246 , n7247 , n7248 , n7249 , n7250 , n7251 , n7252 , n7253 , n7254 , n7255 , n7256 , n7257 , n7258 , n7259 , n7260 , n7261 , n7262 , n7263 , n7264 , n7265 , n7266 , n7267 , n7268 , n7269 , n7270 , n7271 , n7272 , n7273 , n7274 , n7275 , n7276 , n7277 , n7278 , n7279 , n7280 , n7281 , n7282 , n7283 , n7284 , n7285 , n7286 , n7287 , n7288 , n7289 , n7290 , n7291 , n7292 , n7293 , n7294 , n7295 , n7296 , n7297 , n7298 , n7299 , n7300 , n7301 , n7302 , n7303 , n7304 , n7305 , n7306 , n7307 , n7308 , n7309 , n7310 , n7311 , n7312 , n7313 , n7314 , n7315 , n7316 , n7317 , n7318 , n7319 , n7320 , n7321 , n7322 , n7323 , n7324 , n7325 , n7326 , n7327 , n7328 , n7329 , n7330 , n7331 , n7332 , n7333 , n7334 , n7335 , n7336 , n7337 , n7338 , n7339 , n7340 , n7341 , n7342 , n7343 , n7344 , n7345 , n7346 , n7347 , n7348 , n7349 , n7350 , n7351 , n7352 , n7353 , n7354 , n7355 , n7356 , n7357 , n7358 , n7359 , n7360 , n7361 , n7362 , n7363 , n7364 , n7365 , n7366 , n7367 , n7368 , n7369 , n7370 , n7371 , n7372 , n7373 , n7374 , n7375 , n7376 , n7377 , n7378 , n7379 , n7380 , n7381 , n7382 , n7383 , n7384 , n7385 , n7386 , n7387 , n7388 , n7389 , n7390 , n7391 , n7392 , n7393 , n7394 , n7395 , n7396 , n7397 , n7398 , n7399 , n7400 , n7401 , n7402 , n7403 , n7404 , n7405 , n7406 , n7407 , n7408 , n7409 , n7410 , n7411 , n7412 , n7413 , n7414 , n7415 , n7416 , n7417 , n7418 , n7419 , n7420 , n7421 , n7422 , n7423 , n7424 , n7425 , n7426 , n7427 , n7428 , n7429 , n7430 , n7431 , n7432 , n7433 , n7434 , n7435 , n7436 , n7437 , n7438 , n7439 , n7440 , n7441 , n7442 , n7443 , n7444 , n7445 , n7446 , n7447 , n7448 , n7449 , n7450 , n7451 , n7452 , n7453 , n7454 , n7455 , n7456 , n7457 , n7458 , n7459 , n7460 , n7461 , n7462 , n7463 , n7464 , n7465 , n7466 , n7467 , n7468 , n7469 , n7470 , n7471 , n7472 , n7473 , n7474 , n7475 , n7476 , n7477 , n7478 , n7479 , n7480 , n7481 , n7482 , n7483 , n7484 , n7485 , n7486 , n7487 , n7488 , n7489 , n7490 , n7491 , n7492 , n7493 , n7494 , n7495 , n7496 , n7497 , n7498 , n7499 , n7500 , n7501 , n7502 , n7503 , n7504 , n7505 , n7506 , n7507 , n7508 , n7509 , n7510 , n7511 , n7512 , n7513 , n7514 , n7515 , n7516 , n7517 , n7518 , n7519 , n7520 , n7521 , n7522 , n7523 , n7524 , n7525 , n7526 , n7527 , n7528 , n7529 , n7530 , n7531 , n7532 , n7533 , n7534 , n7535 , n7536 , n7537 , n7538 , n7539 , n7540 , n7541 , n7542 , n7543 , n7544 , n7545 , n7546 , n7547 , n7548 , n7549 , n7550 , n7551 , n7552 , n7553 , n7554 , n7555 , n7556 , n7557 , n7558 , n7559 , n7560 , n7561 , n7562 , n7563 , n7564 , n7565 , n7566 , n7567 , n7568 , n7569 , n7570 , n7571 , n7572 , n7573 , n7574 , n7575 , n7576 , n7577 , n7578 , n7579 , n7580 , n7581 , n7582 , n7583 , n7584 , n7585 , n7586 , n7587 , n7588 , n7589 , n7590 , n7591 , n7592 , n7593 , n7594 , n7595 , n7596 , n7597 , n7598 , n7599 , n7600 , n7601 , n7602 , n7603 , n7604 , n7605 , n7606 , n7607 , n7608 , n7609 , n7610 , n7611 , n7612 , n7613 , n7614 , n7615 , n7616 , n7617 , n7618 , n7619 , n7620 , n7621 , n7622 , n7623 , n7624 , n7625 , n7626 , n7627 , n7628 , n7629 , n7630 , n7631 , n7632 , n7633 , n7634 , n7635 , n7636 , n7637 , n7638 , n7639 , n7640 , n7641 , n7642 , n7643 , n7644 , n7645 , n7646 , n7647 , n7648 , n7649 , n7650 , n7651 , n7652 , n7653 , n7654 , n7655 , n7656 , n7657 , n7658 , n7659 , n7660 , n7661 , n7662 , n7663 , n7664 , n7665 , n7666 , n7667 ;
  assign n1002 = ( x286 & x287 ) | ( x286 & x288 ) | ( x287 & x288 ) ;
  assign n1003 = ( x283 & x284 ) | ( x283 & x285 ) | ( x284 & x285 ) ;
  assign n1004 = ( x283 & ~x284 ) | ( x283 & x285 ) | ( ~x284 & x285 ) ;
  assign n1005 = ( ~x283 & x284 ) | ( ~x283 & n1004 ) | ( x284 & n1004 ) ;
  assign n1006 = ( ~x285 & n1004 ) | ( ~x285 & n1005 ) | ( n1004 & n1005 ) ;
  assign n1007 = ( x286 & ~x287 ) | ( x286 & x288 ) | ( ~x287 & x288 ) ;
  assign n1008 = ( ~x286 & x287 ) | ( ~x286 & n1007 ) | ( x287 & n1007 ) ;
  assign n1009 = ( ~x288 & n1007 ) | ( ~x288 & n1008 ) | ( n1007 & n1008 ) ;
  assign n1010 = n1006 & n1009 ;
  assign n1011 = ( n1002 & n1003 ) | ( n1002 & n1010 ) | ( n1003 & n1010 ) ;
  assign n1012 = ( x292 & x293 ) | ( x292 & x294 ) | ( x293 & x294 ) ;
  assign n1013 = ( x289 & x290 ) | ( x289 & x291 ) | ( x290 & x291 ) ;
  assign n1014 = ( x289 & ~x290 ) | ( x289 & x291 ) | ( ~x290 & x291 ) ;
  assign n1015 = ( ~x289 & x290 ) | ( ~x289 & n1014 ) | ( x290 & n1014 ) ;
  assign n1016 = ( ~x291 & n1014 ) | ( ~x291 & n1015 ) | ( n1014 & n1015 ) ;
  assign n1017 = ( x292 & ~x293 ) | ( x292 & x294 ) | ( ~x293 & x294 ) ;
  assign n1018 = ( ~x292 & x293 ) | ( ~x292 & n1017 ) | ( x293 & n1017 ) ;
  assign n1019 = ( ~x294 & n1017 ) | ( ~x294 & n1018 ) | ( n1017 & n1018 ) ;
  assign n1020 = n1016 & n1019 ;
  assign n1021 = ( n1012 & n1013 ) | ( n1012 & n1020 ) | ( n1013 & n1020 ) ;
  assign n1022 = ( n1003 & n1010 ) | ( n1003 & ~n1011 ) | ( n1010 & ~n1011 ) ;
  assign n1023 = ( n1002 & ~n1011 ) | ( n1002 & n1022 ) | ( ~n1011 & n1022 ) ;
  assign n1024 = ( n1013 & n1020 ) | ( n1013 & ~n1021 ) | ( n1020 & ~n1021 ) ;
  assign n1025 = ( n1012 & ~n1021 ) | ( n1012 & n1024 ) | ( ~n1021 & n1024 ) ;
  assign n1026 = n1011 & n1023 ;
  assign n1027 = n1006 & ~n1009 ;
  assign n1028 = ~n1006 & n1009 ;
  assign n1029 = n1027 | n1028 ;
  assign n1030 = n1016 & ~n1019 ;
  assign n1031 = ~n1016 & n1019 ;
  assign n1032 = n1030 | n1031 ;
  assign n1033 = n1029 & n1032 ;
  assign n1034 = ~n1026 & n1033 ;
  assign n1035 = ( n1023 & n1025 ) | ( n1023 & n1034 ) | ( n1025 & n1034 ) ;
  assign n1036 = ( n1011 & n1021 ) | ( n1011 & n1035 ) | ( n1021 & n1035 ) ;
  assign n1037 = ( x280 & x281 ) | ( x280 & x282 ) | ( x281 & x282 ) ;
  assign n1038 = ( x277 & x278 ) | ( x277 & x279 ) | ( x278 & x279 ) ;
  assign n1039 = ( x277 & ~x278 ) | ( x277 & x279 ) | ( ~x278 & x279 ) ;
  assign n1040 = ( ~x277 & x278 ) | ( ~x277 & n1039 ) | ( x278 & n1039 ) ;
  assign n1041 = ( ~x279 & n1039 ) | ( ~x279 & n1040 ) | ( n1039 & n1040 ) ;
  assign n1042 = ( x280 & ~x281 ) | ( x280 & x282 ) | ( ~x281 & x282 ) ;
  assign n1043 = ( ~x280 & x281 ) | ( ~x280 & n1042 ) | ( x281 & n1042 ) ;
  assign n1044 = ( ~x282 & n1042 ) | ( ~x282 & n1043 ) | ( n1042 & n1043 ) ;
  assign n1045 = n1041 & n1044 ;
  assign n1046 = ( n1037 & n1038 ) | ( n1037 & n1045 ) | ( n1038 & n1045 ) ;
  assign n1047 = ( x274 & x275 ) | ( x274 & x276 ) | ( x275 & x276 ) ;
  assign n1048 = ( x271 & x272 ) | ( x271 & x273 ) | ( x272 & x273 ) ;
  assign n1049 = ( x271 & ~x272 ) | ( x271 & x273 ) | ( ~x272 & x273 ) ;
  assign n1050 = ( ~x271 & x272 ) | ( ~x271 & n1049 ) | ( x272 & n1049 ) ;
  assign n1051 = ( ~x273 & n1049 ) | ( ~x273 & n1050 ) | ( n1049 & n1050 ) ;
  assign n1052 = ( x274 & ~x275 ) | ( x274 & x276 ) | ( ~x275 & x276 ) ;
  assign n1053 = ( ~x274 & x275 ) | ( ~x274 & n1052 ) | ( x275 & n1052 ) ;
  assign n1054 = ( ~x276 & n1052 ) | ( ~x276 & n1053 ) | ( n1052 & n1053 ) ;
  assign n1055 = n1051 & n1054 ;
  assign n1056 = ( n1047 & n1048 ) | ( n1047 & n1055 ) | ( n1048 & n1055 ) ;
  assign n1057 = ( n1048 & n1055 ) | ( n1048 & ~n1056 ) | ( n1055 & ~n1056 ) ;
  assign n1058 = ( n1047 & ~n1056 ) | ( n1047 & n1057 ) | ( ~n1056 & n1057 ) ;
  assign n1059 = n1056 & n1058 ;
  assign n1060 = ( n1038 & n1045 ) | ( n1038 & ~n1046 ) | ( n1045 & ~n1046 ) ;
  assign n1061 = ( n1037 & ~n1046 ) | ( n1037 & n1060 ) | ( ~n1046 & n1060 ) ;
  assign n1062 = n1046 & n1061 ;
  assign n1063 = n1041 & ~n1044 ;
  assign n1064 = ~n1041 & n1044 ;
  assign n1065 = n1063 | n1064 ;
  assign n1066 = n1051 & ~n1054 ;
  assign n1067 = ~n1051 & n1054 ;
  assign n1068 = n1066 | n1067 ;
  assign n1069 = n1065 & n1068 ;
  assign n1070 = ~n1062 & n1069 ;
  assign n1071 = n1061 & n1070 ;
  assign n1072 = ~n1059 & n1071 ;
  assign n1073 = ~n1059 & n1070 ;
  assign n1074 = ~n1061 & n1073 ;
  assign n1075 = ( n1058 & n1061 ) | ( n1058 & n1074 ) | ( n1061 & n1074 ) ;
  assign n1076 = n1072 | n1075 ;
  assign n1077 = ( n1046 & n1056 ) | ( n1046 & n1076 ) | ( n1056 & n1076 ) ;
  assign n1078 = n1036 & n1077 ;
  assign n1079 = n1077 & ~n1078 ;
  assign n1080 = ( n1036 & ~n1078 ) | ( n1036 & n1079 ) | ( ~n1078 & n1079 ) ;
  assign n1081 = n1078 | n1080 ;
  assign n1082 = ( n1058 & n1061 ) | ( n1058 & ~n1073 ) | ( n1061 & ~n1073 ) ;
  assign n1083 = n1058 & ~n1072 ;
  assign n1084 = ( n1061 & ~n1082 ) | ( n1061 & n1083 ) | ( ~n1082 & n1083 ) ;
  assign n1085 = ( n1074 & n1082 ) | ( n1074 & ~n1084 ) | ( n1082 & ~n1084 ) ;
  assign n1086 = n1029 & ~n1032 ;
  assign n1087 = ~n1029 & n1032 ;
  assign n1088 = n1086 | n1087 ;
  assign n1089 = ~n1065 & n1068 ;
  assign n1090 = n1065 & ~n1068 ;
  assign n1091 = n1089 | n1090 ;
  assign n1092 = n1088 & n1091 ;
  assign n1093 = n1025 & n1033 ;
  assign n1094 = n1025 | n1034 ;
  assign n1095 = ( n1023 & n1093 ) | ( n1023 & ~n1094 ) | ( n1093 & ~n1094 ) ;
  assign n1096 = ~n1035 & n1094 ;
  assign n1097 = n1095 | n1096 ;
  assign n1098 = n1092 | n1097 ;
  assign n1099 = n1085 & n1098 ;
  assign n1100 = ( n1092 & n1095 ) | ( n1092 & n1096 ) | ( n1095 & n1096 ) ;
  assign n1101 = n1099 | n1100 ;
  assign n1102 = n1046 & ~n1056 ;
  assign n1103 = ~n1046 & n1056 ;
  assign n1104 = n1102 | n1103 ;
  assign n1105 = n1072 | n1104 ;
  assign n1106 = n1075 | n1105 ;
  assign n1107 = n1076 & n1104 ;
  assign n1108 = n1106 & ~n1107 ;
  assign n1109 = ~n1011 & n1021 ;
  assign n1110 = n1011 & ~n1021 ;
  assign n1111 = n1109 | n1110 ;
  assign n1112 = n1035 & n1111 ;
  assign n1113 = n1035 | n1111 ;
  assign n1114 = ~n1112 & n1113 ;
  assign n1115 = ( n1101 & n1108 ) | ( n1101 & n1114 ) | ( n1108 & n1114 ) ;
  assign n1116 = ( n1078 & n1081 ) | ( n1078 & n1115 ) | ( n1081 & n1115 ) ;
  assign n1117 = ( x310 & x311 ) | ( x310 & x312 ) | ( x311 & x312 ) ;
  assign n1118 = ( x307 & x308 ) | ( x307 & x309 ) | ( x308 & x309 ) ;
  assign n1119 = ( x307 & ~x308 ) | ( x307 & x309 ) | ( ~x308 & x309 ) ;
  assign n1120 = ( ~x307 & x308 ) | ( ~x307 & n1119 ) | ( x308 & n1119 ) ;
  assign n1121 = ( ~x309 & n1119 ) | ( ~x309 & n1120 ) | ( n1119 & n1120 ) ;
  assign n1122 = ( x310 & ~x311 ) | ( x310 & x312 ) | ( ~x311 & x312 ) ;
  assign n1123 = ( ~x310 & x311 ) | ( ~x310 & n1122 ) | ( x311 & n1122 ) ;
  assign n1124 = ( ~x312 & n1122 ) | ( ~x312 & n1123 ) | ( n1122 & n1123 ) ;
  assign n1125 = n1121 & n1124 ;
  assign n1126 = ( n1117 & n1118 ) | ( n1117 & n1125 ) | ( n1118 & n1125 ) ;
  assign n1127 = ( x316 & x317 ) | ( x316 & x318 ) | ( x317 & x318 ) ;
  assign n1128 = ( x313 & x314 ) | ( x313 & x315 ) | ( x314 & x315 ) ;
  assign n1129 = ( x313 & ~x314 ) | ( x313 & x315 ) | ( ~x314 & x315 ) ;
  assign n1130 = ( ~x313 & x314 ) | ( ~x313 & n1129 ) | ( x314 & n1129 ) ;
  assign n1131 = ( ~x315 & n1129 ) | ( ~x315 & n1130 ) | ( n1129 & n1130 ) ;
  assign n1132 = ( x316 & ~x317 ) | ( x316 & x318 ) | ( ~x317 & x318 ) ;
  assign n1133 = ( ~x316 & x317 ) | ( ~x316 & n1132 ) | ( x317 & n1132 ) ;
  assign n1134 = ( ~x318 & n1132 ) | ( ~x318 & n1133 ) | ( n1132 & n1133 ) ;
  assign n1135 = n1131 & n1134 ;
  assign n1136 = ( n1127 & n1128 ) | ( n1127 & n1135 ) | ( n1128 & n1135 ) ;
  assign n1137 = ( n1118 & n1125 ) | ( n1118 & ~n1126 ) | ( n1125 & ~n1126 ) ;
  assign n1138 = ( n1117 & ~n1126 ) | ( n1117 & n1137 ) | ( ~n1126 & n1137 ) ;
  assign n1139 = ( n1128 & n1135 ) | ( n1128 & ~n1136 ) | ( n1135 & ~n1136 ) ;
  assign n1140 = ( n1127 & ~n1136 ) | ( n1127 & n1139 ) | ( ~n1136 & n1139 ) ;
  assign n1141 = n1126 & n1138 ;
  assign n1142 = n1121 & ~n1124 ;
  assign n1143 = ~n1121 & n1124 ;
  assign n1144 = n1142 | n1143 ;
  assign n1145 = n1131 & ~n1134 ;
  assign n1146 = ~n1131 & n1134 ;
  assign n1147 = n1145 | n1146 ;
  assign n1148 = n1144 & n1147 ;
  assign n1149 = ~n1141 & n1148 ;
  assign n1150 = ( n1138 & n1140 ) | ( n1138 & n1149 ) | ( n1140 & n1149 ) ;
  assign n1151 = ( n1126 & n1136 ) | ( n1126 & n1150 ) | ( n1136 & n1150 ) ;
  assign n1152 = ( x298 & x299 ) | ( x298 & x300 ) | ( x299 & x300 ) ;
  assign n1153 = ( x295 & x296 ) | ( x295 & x297 ) | ( x296 & x297 ) ;
  assign n1154 = ( x295 & ~x296 ) | ( x295 & x297 ) | ( ~x296 & x297 ) ;
  assign n1155 = ( ~x295 & x296 ) | ( ~x295 & n1154 ) | ( x296 & n1154 ) ;
  assign n1156 = ( ~x297 & n1154 ) | ( ~x297 & n1155 ) | ( n1154 & n1155 ) ;
  assign n1157 = ( x298 & ~x299 ) | ( x298 & x300 ) | ( ~x299 & x300 ) ;
  assign n1158 = ( ~x298 & x299 ) | ( ~x298 & n1157 ) | ( x299 & n1157 ) ;
  assign n1159 = ( ~x300 & n1157 ) | ( ~x300 & n1158 ) | ( n1157 & n1158 ) ;
  assign n1160 = n1156 & n1159 ;
  assign n1161 = ( n1152 & n1153 ) | ( n1152 & n1160 ) | ( n1153 & n1160 ) ;
  assign n1162 = ( x304 & x305 ) | ( x304 & x306 ) | ( x305 & x306 ) ;
  assign n1163 = ( x301 & x302 ) | ( x301 & x303 ) | ( x302 & x303 ) ;
  assign n1164 = ( x301 & ~x302 ) | ( x301 & x303 ) | ( ~x302 & x303 ) ;
  assign n1165 = ( ~x301 & x302 ) | ( ~x301 & n1164 ) | ( x302 & n1164 ) ;
  assign n1166 = ( ~x303 & n1164 ) | ( ~x303 & n1165 ) | ( n1164 & n1165 ) ;
  assign n1167 = ( x304 & ~x305 ) | ( x304 & x306 ) | ( ~x305 & x306 ) ;
  assign n1168 = ( ~x304 & x305 ) | ( ~x304 & n1167 ) | ( x305 & n1167 ) ;
  assign n1169 = ( ~x306 & n1167 ) | ( ~x306 & n1168 ) | ( n1167 & n1168 ) ;
  assign n1170 = n1166 & n1169 ;
  assign n1171 = ( n1162 & n1163 ) | ( n1162 & n1170 ) | ( n1163 & n1170 ) ;
  assign n1172 = ( n1153 & n1160 ) | ( n1153 & ~n1161 ) | ( n1160 & ~n1161 ) ;
  assign n1173 = ( n1152 & ~n1161 ) | ( n1152 & n1172 ) | ( ~n1161 & n1172 ) ;
  assign n1174 = ( n1163 & n1170 ) | ( n1163 & ~n1171 ) | ( n1170 & ~n1171 ) ;
  assign n1175 = ( n1162 & ~n1171 ) | ( n1162 & n1174 ) | ( ~n1171 & n1174 ) ;
  assign n1176 = n1161 & n1173 ;
  assign n1177 = n1171 & n1175 ;
  assign n1178 = n1156 & ~n1159 ;
  assign n1179 = ~n1156 & n1159 ;
  assign n1180 = n1178 | n1179 ;
  assign n1181 = n1166 & ~n1169 ;
  assign n1182 = ~n1166 & n1169 ;
  assign n1183 = n1181 | n1182 ;
  assign n1184 = n1180 & n1183 ;
  assign n1185 = ~n1177 & n1184 ;
  assign n1186 = ~n1176 & n1185 ;
  assign n1187 = ~n1175 & n1186 ;
  assign n1188 = ( n1173 & n1175 ) | ( n1173 & n1187 ) | ( n1175 & n1187 ) ;
  assign n1189 = n1175 & n1185 ;
  assign n1190 = ~n1176 & n1189 ;
  assign n1191 = n1188 | n1190 ;
  assign n1192 = ( n1161 & n1171 ) | ( n1161 & n1191 ) | ( n1171 & n1191 ) ;
  assign n1193 = ~n1161 & n1171 ;
  assign n1194 = n1161 & ~n1171 ;
  assign n1195 = n1193 | n1194 ;
  assign n1196 = n1190 | n1195 ;
  assign n1197 = n1188 | n1196 ;
  assign n1198 = n1191 & n1195 ;
  assign n1199 = n1197 & ~n1198 ;
  assign n1200 = ~n1126 & n1136 ;
  assign n1201 = n1126 & ~n1136 ;
  assign n1202 = n1200 | n1201 ;
  assign n1203 = n1150 & n1202 ;
  assign n1204 = n1150 | n1202 ;
  assign n1205 = ~n1203 & n1204 ;
  assign n1206 = n1199 | n1205 ;
  assign n1207 = ( n1173 & n1175 ) | ( n1173 & ~n1186 ) | ( n1175 & ~n1186 ) ;
  assign n1208 = n1173 & ~n1190 ;
  assign n1209 = ( n1175 & ~n1207 ) | ( n1175 & n1208 ) | ( ~n1207 & n1208 ) ;
  assign n1210 = ( n1187 & n1207 ) | ( n1187 & ~n1209 ) | ( n1207 & ~n1209 ) ;
  assign n1211 = n1144 & ~n1147 ;
  assign n1212 = ~n1144 & n1147 ;
  assign n1213 = n1211 | n1212 ;
  assign n1214 = n1180 & ~n1183 ;
  assign n1215 = ~n1180 & n1183 ;
  assign n1216 = n1214 | n1215 ;
  assign n1217 = n1213 & n1216 ;
  assign n1218 = n1140 | n1149 ;
  assign n1219 = ~n1150 & n1218 ;
  assign n1220 = n1140 & n1148 ;
  assign n1221 = ( n1138 & ~n1218 ) | ( n1138 & n1220 ) | ( ~n1218 & n1220 ) ;
  assign n1222 = n1219 | n1221 ;
  assign n1223 = n1217 | n1222 ;
  assign n1224 = ( n1217 & n1219 ) | ( n1217 & n1221 ) | ( n1219 & n1221 ) ;
  assign n1225 = ( n1210 & n1223 ) | ( n1210 & n1224 ) | ( n1223 & n1224 ) ;
  assign n1226 = n1206 & n1225 ;
  assign n1227 = n1199 & n1205 ;
  assign n1228 = n1226 | n1227 ;
  assign n1229 = ( n1151 & n1192 ) | ( n1151 & n1228 ) | ( n1192 & n1228 ) ;
  assign n1230 = n1116 & n1229 ;
  assign n1231 = ~n1151 & n1192 ;
  assign n1232 = n1151 & ~n1192 ;
  assign n1233 = n1231 | n1232 ;
  assign n1234 = n1227 | n1233 ;
  assign n1235 = n1226 | n1234 ;
  assign n1236 = n1228 & n1233 ;
  assign n1237 = n1235 & ~n1236 ;
  assign n1238 = n1080 | n1115 ;
  assign n1239 = ~n1080 & n1238 ;
  assign n1240 = ( ~n1115 & n1238 ) | ( ~n1115 & n1239 ) | ( n1238 & n1239 ) ;
  assign n1241 = n1237 | n1240 ;
  assign n1242 = ( n1101 & ~n1108 ) | ( n1101 & n1114 ) | ( ~n1108 & n1114 ) ;
  assign n1243 = ( ~n1101 & n1108 ) | ( ~n1101 & n1242 ) | ( n1108 & n1242 ) ;
  assign n1244 = ( ~n1114 & n1242 ) | ( ~n1114 & n1243 ) | ( n1242 & n1243 ) ;
  assign n1245 = ( ~n1199 & n1205 ) | ( ~n1199 & n1225 ) | ( n1205 & n1225 ) ;
  assign n1246 = ( n1199 & ~n1225 ) | ( n1199 & n1245 ) | ( ~n1225 & n1245 ) ;
  assign n1247 = ( ~n1205 & n1245 ) | ( ~n1205 & n1246 ) | ( n1245 & n1246 ) ;
  assign n1248 = n1213 & ~n1216 ;
  assign n1249 = ~n1213 & n1216 ;
  assign n1250 = n1248 | n1249 ;
  assign n1251 = n1088 & ~n1091 ;
  assign n1252 = ~n1088 & n1091 ;
  assign n1253 = n1251 | n1252 ;
  assign n1254 = n1250 & n1253 ;
  assign n1255 = ~n1217 & n1223 ;
  assign n1256 = ( ~n1222 & n1223 ) | ( ~n1222 & n1255 ) | ( n1223 & n1255 ) ;
  assign n1257 = n1210 & ~n1256 ;
  assign n1258 = ~n1210 & n1256 ;
  assign n1259 = n1257 | n1258 ;
  assign n1260 = ( n1085 & n1092 ) | ( n1085 & ~n1097 ) | ( n1092 & ~n1097 ) ;
  assign n1261 = ( ~n1085 & n1097 ) | ( ~n1085 & n1260 ) | ( n1097 & n1260 ) ;
  assign n1262 = ( ~n1092 & n1260 ) | ( ~n1092 & n1261 ) | ( n1260 & n1261 ) ;
  assign n1263 = ( n1254 & n1259 ) | ( n1254 & n1262 ) | ( n1259 & n1262 ) ;
  assign n1264 = ( n1244 & n1247 ) | ( n1244 & n1263 ) | ( n1247 & n1263 ) ;
  assign n1265 = n1241 & n1264 ;
  assign n1266 = n1237 & n1240 ;
  assign n1267 = n1265 | n1266 ;
  assign n1268 = n1229 & ~n1230 ;
  assign n1269 = ( n1116 & ~n1230 ) | ( n1116 & n1268 ) | ( ~n1230 & n1268 ) ;
  assign n1270 = ( n1081 & n1229 ) | ( n1081 & n1269 ) | ( n1229 & n1269 ) ;
  assign n1271 = ( n1230 & n1267 ) | ( n1230 & n1270 ) | ( n1267 & n1270 ) ;
  assign n1272 = ( x340 & x341 ) | ( x340 & x342 ) | ( x341 & x342 ) ;
  assign n1273 = ( x337 & x338 ) | ( x337 & x339 ) | ( x338 & x339 ) ;
  assign n1274 = ( x337 & ~x338 ) | ( x337 & x339 ) | ( ~x338 & x339 ) ;
  assign n1275 = ( ~x337 & x338 ) | ( ~x337 & n1274 ) | ( x338 & n1274 ) ;
  assign n1276 = ( ~x339 & n1274 ) | ( ~x339 & n1275 ) | ( n1274 & n1275 ) ;
  assign n1277 = ( x340 & ~x341 ) | ( x340 & x342 ) | ( ~x341 & x342 ) ;
  assign n1278 = ( ~x340 & x341 ) | ( ~x340 & n1277 ) | ( x341 & n1277 ) ;
  assign n1279 = ( ~x342 & n1277 ) | ( ~x342 & n1278 ) | ( n1277 & n1278 ) ;
  assign n1280 = n1276 & n1279 ;
  assign n1281 = ( n1272 & n1273 ) | ( n1272 & n1280 ) | ( n1273 & n1280 ) ;
  assign n1282 = ( x331 & ~x332 ) | ( x331 & x333 ) | ( ~x332 & x333 ) ;
  assign n1283 = ( ~x331 & x332 ) | ( ~x331 & n1282 ) | ( x332 & n1282 ) ;
  assign n1284 = ( ~x333 & n1282 ) | ( ~x333 & n1283 ) | ( n1282 & n1283 ) ;
  assign n1285 = ( x334 & ~x335 ) | ( x334 & x336 ) | ( ~x335 & x336 ) ;
  assign n1286 = ( ~x334 & x335 ) | ( ~x334 & n1285 ) | ( x335 & n1285 ) ;
  assign n1287 = ( ~x336 & n1285 ) | ( ~x336 & n1286 ) | ( n1285 & n1286 ) ;
  assign n1288 = n1284 & n1287 ;
  assign n1289 = ( x334 & x335 ) | ( x334 & x336 ) | ( x335 & x336 ) ;
  assign n1290 = ( x331 & x332 ) | ( x331 & x333 ) | ( x332 & x333 ) ;
  assign n1291 = ( n1288 & n1289 ) | ( n1288 & n1290 ) | ( n1289 & n1290 ) ;
  assign n1292 = ( n1273 & n1280 ) | ( n1273 & ~n1281 ) | ( n1280 & ~n1281 ) ;
  assign n1293 = ( n1272 & ~n1281 ) | ( n1272 & n1292 ) | ( ~n1281 & n1292 ) ;
  assign n1294 = ( n1288 & n1290 ) | ( n1288 & ~n1291 ) | ( n1290 & ~n1291 ) ;
  assign n1295 = ( n1289 & ~n1291 ) | ( n1289 & n1294 ) | ( ~n1291 & n1294 ) ;
  assign n1296 = n1291 & n1295 ;
  assign n1297 = n1276 & ~n1279 ;
  assign n1298 = ~n1276 & n1279 ;
  assign n1299 = n1297 | n1298 ;
  assign n1300 = n1284 & ~n1287 ;
  assign n1301 = ~n1284 & n1287 ;
  assign n1302 = n1300 | n1301 ;
  assign n1303 = n1299 & n1302 ;
  assign n1304 = ~n1296 & n1303 ;
  assign n1305 = ( n1293 & n1295 ) | ( n1293 & n1304 ) | ( n1295 & n1304 ) ;
  assign n1306 = ( n1281 & n1291 ) | ( n1281 & n1305 ) | ( n1291 & n1305 ) ;
  assign n1307 = ( x328 & x329 ) | ( x328 & x330 ) | ( x329 & x330 ) ;
  assign n1308 = ( x325 & x326 ) | ( x325 & x327 ) | ( x326 & x327 ) ;
  assign n1309 = ( x325 & ~x326 ) | ( x325 & x327 ) | ( ~x326 & x327 ) ;
  assign n1310 = ( ~x325 & x326 ) | ( ~x325 & n1309 ) | ( x326 & n1309 ) ;
  assign n1311 = ( ~x327 & n1309 ) | ( ~x327 & n1310 ) | ( n1309 & n1310 ) ;
  assign n1312 = ( x328 & ~x329 ) | ( x328 & x330 ) | ( ~x329 & x330 ) ;
  assign n1313 = ( ~x328 & x329 ) | ( ~x328 & n1312 ) | ( x329 & n1312 ) ;
  assign n1314 = ( ~x330 & n1312 ) | ( ~x330 & n1313 ) | ( n1312 & n1313 ) ;
  assign n1315 = n1311 & n1314 ;
  assign n1316 = ( n1307 & n1308 ) | ( n1307 & n1315 ) | ( n1308 & n1315 ) ;
  assign n1317 = ( x322 & x323 ) | ( x322 & x324 ) | ( x323 & x324 ) ;
  assign n1318 = ( x319 & x320 ) | ( x319 & x321 ) | ( x320 & x321 ) ;
  assign n1319 = ( x319 & ~x320 ) | ( x319 & x321 ) | ( ~x320 & x321 ) ;
  assign n1320 = ( ~x319 & x320 ) | ( ~x319 & n1319 ) | ( x320 & n1319 ) ;
  assign n1321 = ( ~x321 & n1319 ) | ( ~x321 & n1320 ) | ( n1319 & n1320 ) ;
  assign n1322 = ( x322 & ~x323 ) | ( x322 & x324 ) | ( ~x323 & x324 ) ;
  assign n1323 = ( ~x322 & x323 ) | ( ~x322 & n1322 ) | ( x323 & n1322 ) ;
  assign n1324 = ( ~x324 & n1322 ) | ( ~x324 & n1323 ) | ( n1322 & n1323 ) ;
  assign n1325 = n1321 & n1324 ;
  assign n1326 = ( n1317 & n1318 ) | ( n1317 & n1325 ) | ( n1318 & n1325 ) ;
  assign n1327 = ( n1318 & n1325 ) | ( n1318 & ~n1326 ) | ( n1325 & ~n1326 ) ;
  assign n1328 = ( n1317 & ~n1326 ) | ( n1317 & n1327 ) | ( ~n1326 & n1327 ) ;
  assign n1329 = n1326 & n1328 ;
  assign n1330 = ( n1308 & n1315 ) | ( n1308 & ~n1316 ) | ( n1315 & ~n1316 ) ;
  assign n1331 = ( n1307 & ~n1316 ) | ( n1307 & n1330 ) | ( ~n1316 & n1330 ) ;
  assign n1332 = n1316 & n1331 ;
  assign n1333 = n1311 & ~n1314 ;
  assign n1334 = ~n1311 & n1314 ;
  assign n1335 = n1333 | n1334 ;
  assign n1336 = n1321 & ~n1324 ;
  assign n1337 = ~n1321 & n1324 ;
  assign n1338 = n1336 | n1337 ;
  assign n1339 = n1335 & n1338 ;
  assign n1340 = ~n1332 & n1339 ;
  assign n1341 = n1331 & n1340 ;
  assign n1342 = ~n1329 & n1341 ;
  assign n1343 = ~n1329 & n1340 ;
  assign n1344 = ~n1331 & n1343 ;
  assign n1345 = ( n1328 & n1331 ) | ( n1328 & n1344 ) | ( n1331 & n1344 ) ;
  assign n1346 = n1342 | n1345 ;
  assign n1347 = ( n1316 & n1326 ) | ( n1316 & n1346 ) | ( n1326 & n1346 ) ;
  assign n1348 = ( n1328 & n1331 ) | ( n1328 & ~n1343 ) | ( n1331 & ~n1343 ) ;
  assign n1349 = n1328 & ~n1342 ;
  assign n1350 = ( n1331 & ~n1348 ) | ( n1331 & n1349 ) | ( ~n1348 & n1349 ) ;
  assign n1351 = ( n1344 & n1348 ) | ( n1344 & ~n1350 ) | ( n1348 & ~n1350 ) ;
  assign n1352 = ~n1299 & n1302 ;
  assign n1353 = n1299 & ~n1302 ;
  assign n1354 = n1352 | n1353 ;
  assign n1355 = ~n1335 & n1338 ;
  assign n1356 = n1335 & ~n1338 ;
  assign n1357 = n1355 | n1356 ;
  assign n1358 = n1354 & n1357 ;
  assign n1359 = n1293 & n1303 ;
  assign n1360 = n1293 | n1304 ;
  assign n1361 = ( n1295 & n1359 ) | ( n1295 & ~n1360 ) | ( n1359 & ~n1360 ) ;
  assign n1362 = ~n1305 & n1360 ;
  assign n1363 = n1361 | n1362 ;
  assign n1364 = n1358 | n1363 ;
  assign n1365 = n1351 & n1364 ;
  assign n1366 = ( n1358 & n1361 ) | ( n1358 & n1362 ) | ( n1361 & n1362 ) ;
  assign n1367 = n1365 | n1366 ;
  assign n1368 = n1316 & ~n1326 ;
  assign n1369 = ~n1316 & n1326 ;
  assign n1370 = n1368 | n1369 ;
  assign n1371 = n1342 | n1370 ;
  assign n1372 = n1345 | n1371 ;
  assign n1373 = n1346 & n1370 ;
  assign n1374 = n1372 & ~n1373 ;
  assign n1375 = ( n1281 & n1291 ) | ( n1281 & ~n1305 ) | ( n1291 & ~n1305 ) ;
  assign n1376 = ( n1281 & ~n1291 ) | ( n1281 & n1305 ) | ( ~n1291 & n1305 ) ;
  assign n1377 = ( ~n1281 & n1375 ) | ( ~n1281 & n1376 ) | ( n1375 & n1376 ) ;
  assign n1378 = ( n1367 & n1374 ) | ( n1367 & n1377 ) | ( n1374 & n1377 ) ;
  assign n1379 = ( n1306 & n1347 ) | ( n1306 & n1378 ) | ( n1347 & n1378 ) ;
  assign n1380 = ( x364 & x365 ) | ( x364 & x366 ) | ( x365 & x366 ) ;
  assign n1381 = ( x361 & x362 ) | ( x361 & x363 ) | ( x362 & x363 ) ;
  assign n1382 = ( x361 & ~x362 ) | ( x361 & x363 ) | ( ~x362 & x363 ) ;
  assign n1383 = ( ~x361 & x362 ) | ( ~x361 & n1382 ) | ( x362 & n1382 ) ;
  assign n1384 = ( ~x363 & n1382 ) | ( ~x363 & n1383 ) | ( n1382 & n1383 ) ;
  assign n1385 = ( x364 & ~x365 ) | ( x364 & x366 ) | ( ~x365 & x366 ) ;
  assign n1386 = ( ~x364 & x365 ) | ( ~x364 & n1385 ) | ( x365 & n1385 ) ;
  assign n1387 = ( ~x366 & n1385 ) | ( ~x366 & n1386 ) | ( n1385 & n1386 ) ;
  assign n1388 = n1384 & n1387 ;
  assign n1389 = ( n1380 & n1381 ) | ( n1380 & n1388 ) | ( n1381 & n1388 ) ;
  assign n1390 = ( x355 & ~x356 ) | ( x355 & x357 ) | ( ~x356 & x357 ) ;
  assign n1391 = ( ~x355 & x356 ) | ( ~x355 & n1390 ) | ( x356 & n1390 ) ;
  assign n1392 = ( ~x357 & n1390 ) | ( ~x357 & n1391 ) | ( n1390 & n1391 ) ;
  assign n1393 = ( x358 & ~x359 ) | ( x358 & x360 ) | ( ~x359 & x360 ) ;
  assign n1394 = ( ~x358 & x359 ) | ( ~x358 & n1393 ) | ( x359 & n1393 ) ;
  assign n1395 = ( ~x360 & n1393 ) | ( ~x360 & n1394 ) | ( n1393 & n1394 ) ;
  assign n1396 = n1392 & n1395 ;
  assign n1397 = ( x358 & x359 ) | ( x358 & x360 ) | ( x359 & x360 ) ;
  assign n1398 = ( x355 & x356 ) | ( x355 & x357 ) | ( x356 & x357 ) ;
  assign n1399 = ( n1396 & n1397 ) | ( n1396 & n1398 ) | ( n1397 & n1398 ) ;
  assign n1400 = ( n1381 & n1388 ) | ( n1381 & ~n1389 ) | ( n1388 & ~n1389 ) ;
  assign n1401 = ( n1380 & ~n1389 ) | ( n1380 & n1400 ) | ( ~n1389 & n1400 ) ;
  assign n1402 = ( n1396 & n1398 ) | ( n1396 & ~n1399 ) | ( n1398 & ~n1399 ) ;
  assign n1403 = ( n1397 & ~n1399 ) | ( n1397 & n1402 ) | ( ~n1399 & n1402 ) ;
  assign n1404 = n1399 & n1403 ;
  assign n1405 = n1392 & ~n1395 ;
  assign n1406 = ~n1392 & n1395 ;
  assign n1407 = n1405 | n1406 ;
  assign n1408 = n1384 & ~n1387 ;
  assign n1409 = ~n1384 & n1387 ;
  assign n1410 = n1408 | n1409 ;
  assign n1411 = ~n1388 & n1410 ;
  assign n1412 = n1407 & n1411 ;
  assign n1413 = ~n1404 & n1412 ;
  assign n1414 = ( n1401 & n1403 ) | ( n1401 & n1413 ) | ( n1403 & n1413 ) ;
  assign n1415 = ( n1389 & n1399 ) | ( n1389 & n1414 ) | ( n1399 & n1414 ) ;
  assign n1416 = ( x343 & ~x344 ) | ( x343 & x345 ) | ( ~x344 & x345 ) ;
  assign n1417 = ( ~x343 & x344 ) | ( ~x343 & n1416 ) | ( x344 & n1416 ) ;
  assign n1418 = ( ~x345 & n1416 ) | ( ~x345 & n1417 ) | ( n1416 & n1417 ) ;
  assign n1419 = ( x346 & ~x347 ) | ( x346 & x348 ) | ( ~x347 & x348 ) ;
  assign n1420 = ( ~x346 & x347 ) | ( ~x346 & n1419 ) | ( x347 & n1419 ) ;
  assign n1421 = ( ~x348 & n1419 ) | ( ~x348 & n1420 ) | ( n1419 & n1420 ) ;
  assign n1422 = n1418 & n1421 ;
  assign n1423 = ( x346 & x347 ) | ( x346 & x348 ) | ( x347 & x348 ) ;
  assign n1424 = ( x343 & x344 ) | ( x343 & x345 ) | ( x344 & x345 ) ;
  assign n1425 = ( n1422 & n1423 ) | ( n1422 & n1424 ) | ( n1423 & n1424 ) ;
  assign n1426 = ( x352 & x353 ) | ( x352 & x354 ) | ( x353 & x354 ) ;
  assign n1427 = ( x349 & x350 ) | ( x349 & x351 ) | ( x350 & x351 ) ;
  assign n1428 = ( x349 & ~x350 ) | ( x349 & x351 ) | ( ~x350 & x351 ) ;
  assign n1429 = ( ~x349 & x350 ) | ( ~x349 & n1428 ) | ( x350 & n1428 ) ;
  assign n1430 = ( ~x351 & n1428 ) | ( ~x351 & n1429 ) | ( n1428 & n1429 ) ;
  assign n1431 = ( x352 & ~x353 ) | ( x352 & x354 ) | ( ~x353 & x354 ) ;
  assign n1432 = ( ~x352 & x353 ) | ( ~x352 & n1431 ) | ( x353 & n1431 ) ;
  assign n1433 = ( ~x354 & n1431 ) | ( ~x354 & n1432 ) | ( n1431 & n1432 ) ;
  assign n1434 = n1430 & n1433 ;
  assign n1435 = ( n1426 & n1427 ) | ( n1426 & n1434 ) | ( n1427 & n1434 ) ;
  assign n1436 = ( n1422 & n1424 ) | ( n1422 & ~n1425 ) | ( n1424 & ~n1425 ) ;
  assign n1437 = ( n1423 & ~n1425 ) | ( n1423 & n1436 ) | ( ~n1425 & n1436 ) ;
  assign n1438 = ( n1427 & n1434 ) | ( n1427 & ~n1435 ) | ( n1434 & ~n1435 ) ;
  assign n1439 = ( n1426 & ~n1435 ) | ( n1426 & n1438 ) | ( ~n1435 & n1438 ) ;
  assign n1440 = n1425 & n1437 ;
  assign n1441 = n1435 & n1439 ;
  assign n1442 = n1418 & ~n1421 ;
  assign n1443 = ~n1418 & n1421 ;
  assign n1444 = n1442 | n1443 ;
  assign n1445 = n1430 & ~n1433 ;
  assign n1446 = ~n1430 & n1433 ;
  assign n1447 = n1445 | n1446 ;
  assign n1448 = n1444 & n1447 ;
  assign n1449 = ~n1441 & n1448 ;
  assign n1450 = ~n1440 & n1449 ;
  assign n1451 = ~n1439 & n1450 ;
  assign n1452 = ( n1437 & n1439 ) | ( n1437 & n1451 ) | ( n1439 & n1451 ) ;
  assign n1453 = n1439 & n1449 ;
  assign n1454 = ~n1440 & n1453 ;
  assign n1455 = n1452 | n1454 ;
  assign n1456 = ( n1425 & n1435 ) | ( n1425 & n1455 ) | ( n1435 & n1455 ) ;
  assign n1457 = ~n1425 & n1435 ;
  assign n1458 = n1425 & ~n1435 ;
  assign n1459 = n1457 | n1458 ;
  assign n1460 = n1454 | n1459 ;
  assign n1461 = n1452 | n1460 ;
  assign n1462 = n1455 & n1459 ;
  assign n1463 = n1461 & ~n1462 ;
  assign n1464 = ( n1389 & n1399 ) | ( n1389 & ~n1414 ) | ( n1399 & ~n1414 ) ;
  assign n1465 = ( n1389 & ~n1399 ) | ( n1389 & n1414 ) | ( ~n1399 & n1414 ) ;
  assign n1466 = ( ~n1389 & n1464 ) | ( ~n1389 & n1465 ) | ( n1464 & n1465 ) ;
  assign n1467 = n1463 | n1466 ;
  assign n1468 = ( n1437 & n1439 ) | ( n1437 & ~n1450 ) | ( n1439 & ~n1450 ) ;
  assign n1469 = n1437 & ~n1454 ;
  assign n1470 = ( n1439 & ~n1468 ) | ( n1439 & n1469 ) | ( ~n1468 & n1469 ) ;
  assign n1471 = ( n1451 & n1468 ) | ( n1451 & ~n1470 ) | ( n1468 & ~n1470 ) ;
  assign n1472 = n1407 & ~n1411 ;
  assign n1473 = ~n1407 & n1411 ;
  assign n1474 = n1472 | n1473 ;
  assign n1475 = n1444 & ~n1447 ;
  assign n1476 = ~n1444 & n1447 ;
  assign n1477 = n1475 | n1476 ;
  assign n1478 = n1474 & n1477 ;
  assign n1479 = n1401 | n1413 ;
  assign n1480 = ~n1414 & n1479 ;
  assign n1481 = n1401 & n1412 ;
  assign n1482 = ( n1403 & ~n1479 ) | ( n1403 & n1481 ) | ( ~n1479 & n1481 ) ;
  assign n1483 = n1480 | n1482 ;
  assign n1484 = n1478 | n1483 ;
  assign n1485 = ( n1478 & n1480 ) | ( n1478 & n1482 ) | ( n1480 & n1482 ) ;
  assign n1486 = ( n1471 & n1484 ) | ( n1471 & n1485 ) | ( n1484 & n1485 ) ;
  assign n1487 = n1467 & n1486 ;
  assign n1488 = n1463 & n1466 ;
  assign n1489 = n1487 | n1488 ;
  assign n1490 = ( n1415 & n1456 ) | ( n1415 & n1489 ) | ( n1456 & n1489 ) ;
  assign n1491 = n1379 & n1490 ;
  assign n1492 = ~n1415 & n1456 ;
  assign n1493 = n1415 & ~n1456 ;
  assign n1494 = n1492 | n1493 ;
  assign n1495 = n1488 | n1494 ;
  assign n1496 = n1487 | n1495 ;
  assign n1497 = n1489 & n1494 ;
  assign n1498 = n1496 & ~n1497 ;
  assign n1499 = ~n1306 & n1347 ;
  assign n1500 = n1306 & ~n1347 ;
  assign n1501 = n1499 | n1500 ;
  assign n1502 = n1378 | n1501 ;
  assign n1503 = ~n1501 & n1502 ;
  assign n1504 = ( ~n1378 & n1502 ) | ( ~n1378 & n1503 ) | ( n1502 & n1503 ) ;
  assign n1505 = n1498 | n1504 ;
  assign n1506 = ( n1367 & ~n1374 ) | ( n1367 & n1377 ) | ( ~n1374 & n1377 ) ;
  assign n1507 = ( ~n1367 & n1374 ) | ( ~n1367 & n1506 ) | ( n1374 & n1506 ) ;
  assign n1508 = ( ~n1377 & n1506 ) | ( ~n1377 & n1507 ) | ( n1506 & n1507 ) ;
  assign n1509 = ( ~n1463 & n1466 ) | ( ~n1463 & n1486 ) | ( n1466 & n1486 ) ;
  assign n1510 = ( n1463 & ~n1486 ) | ( n1463 & n1509 ) | ( ~n1486 & n1509 ) ;
  assign n1511 = ( ~n1466 & n1509 ) | ( ~n1466 & n1510 ) | ( n1509 & n1510 ) ;
  assign n1512 = n1474 & ~n1477 ;
  assign n1513 = ~n1474 & n1477 ;
  assign n1514 = n1512 | n1513 ;
  assign n1515 = n1354 & ~n1357 ;
  assign n1516 = ~n1354 & n1357 ;
  assign n1517 = n1515 | n1516 ;
  assign n1518 = n1514 & n1517 ;
  assign n1519 = ~n1478 & n1484 ;
  assign n1520 = ( ~n1483 & n1484 ) | ( ~n1483 & n1519 ) | ( n1484 & n1519 ) ;
  assign n1521 = n1471 & ~n1520 ;
  assign n1522 = ~n1471 & n1520 ;
  assign n1523 = n1521 | n1522 ;
  assign n1524 = ( n1351 & n1358 ) | ( n1351 & ~n1363 ) | ( n1358 & ~n1363 ) ;
  assign n1525 = ( ~n1351 & n1363 ) | ( ~n1351 & n1524 ) | ( n1363 & n1524 ) ;
  assign n1526 = ( ~n1358 & n1524 ) | ( ~n1358 & n1525 ) | ( n1524 & n1525 ) ;
  assign n1527 = ( n1518 & n1523 ) | ( n1518 & n1526 ) | ( n1523 & n1526 ) ;
  assign n1528 = ( n1508 & n1511 ) | ( n1508 & n1527 ) | ( n1511 & n1527 ) ;
  assign n1529 = n1505 & n1528 ;
  assign n1530 = n1498 & n1504 ;
  assign n1531 = n1529 | n1530 ;
  assign n1532 = n1490 & ~n1491 ;
  assign n1533 = ( n1379 & ~n1491 ) | ( n1379 & n1532 ) | ( ~n1491 & n1532 ) ;
  assign n1534 = n1531 & n1533 ;
  assign n1535 = ( n1490 & n1531 ) | ( n1490 & n1534 ) | ( n1531 & n1534 ) ;
  assign n1536 = n1491 | n1535 ;
  assign n1537 = n1530 | n1533 ;
  assign n1538 = n1529 | n1537 ;
  assign n1539 = ~n1534 & n1538 ;
  assign n1540 = n1266 | n1269 ;
  assign n1541 = n1265 | n1540 ;
  assign n1542 = n1267 & n1269 ;
  assign n1543 = n1541 & ~n1542 ;
  assign n1544 = ( ~n1244 & n1247 ) | ( ~n1244 & n1263 ) | ( n1247 & n1263 ) ;
  assign n1545 = ( n1244 & ~n1263 ) | ( n1244 & n1544 ) | ( ~n1263 & n1544 ) ;
  assign n1546 = ( ~n1247 & n1544 ) | ( ~n1247 & n1545 ) | ( n1544 & n1545 ) ;
  assign n1547 = ( ~n1508 & n1511 ) | ( ~n1508 & n1527 ) | ( n1511 & n1527 ) ;
  assign n1548 = ( n1508 & ~n1527 ) | ( n1508 & n1547 ) | ( ~n1527 & n1547 ) ;
  assign n1549 = ( ~n1511 & n1547 ) | ( ~n1511 & n1548 ) | ( n1547 & n1548 ) ;
  assign n1550 = n1514 & ~n1517 ;
  assign n1551 = ~n1514 & n1517 ;
  assign n1552 = n1550 | n1551 ;
  assign n1553 = n1250 & ~n1253 ;
  assign n1554 = ~n1250 & n1253 ;
  assign n1555 = n1553 | n1554 ;
  assign n1556 = n1552 & n1555 ;
  assign n1557 = ( n1518 & ~n1523 ) | ( n1518 & n1526 ) | ( ~n1523 & n1526 ) ;
  assign n1558 = ( ~n1518 & n1523 ) | ( ~n1518 & n1557 ) | ( n1523 & n1557 ) ;
  assign n1559 = ( ~n1526 & n1557 ) | ( ~n1526 & n1558 ) | ( n1557 & n1558 ) ;
  assign n1560 = ( n1254 & ~n1259 ) | ( n1254 & n1262 ) | ( ~n1259 & n1262 ) ;
  assign n1561 = ( ~n1254 & n1259 ) | ( ~n1254 & n1560 ) | ( n1259 & n1560 ) ;
  assign n1562 = ( ~n1262 & n1560 ) | ( ~n1262 & n1561 ) | ( n1560 & n1561 ) ;
  assign n1563 = ( n1556 & n1559 ) | ( n1556 & n1562 ) | ( n1559 & n1562 ) ;
  assign n1564 = ( n1546 & n1549 ) | ( n1546 & n1563 ) | ( n1549 & n1563 ) ;
  assign n1565 = ( ~n1498 & n1504 ) | ( ~n1498 & n1528 ) | ( n1504 & n1528 ) ;
  assign n1566 = ( n1498 & ~n1528 ) | ( n1498 & n1565 ) | ( ~n1528 & n1565 ) ;
  assign n1567 = ( ~n1504 & n1565 ) | ( ~n1504 & n1566 ) | ( n1565 & n1566 ) ;
  assign n1568 = ( ~n1237 & n1240 ) | ( ~n1237 & n1264 ) | ( n1240 & n1264 ) ;
  assign n1569 = ( n1237 & ~n1264 ) | ( n1237 & n1568 ) | ( ~n1264 & n1568 ) ;
  assign n1570 = ( ~n1240 & n1568 ) | ( ~n1240 & n1569 ) | ( n1568 & n1569 ) ;
  assign n1571 = ( n1564 & n1567 ) | ( n1564 & n1570 ) | ( n1567 & n1570 ) ;
  assign n1572 = ( n1539 & n1543 ) | ( n1539 & n1571 ) | ( n1543 & n1571 ) ;
  assign n1573 = ( n1271 & n1536 ) | ( n1271 & ~n1572 ) | ( n1536 & ~n1572 ) ;
  assign n1574 = ( ~n1536 & n1572 ) | ( ~n1536 & n1573 ) | ( n1572 & n1573 ) ;
  assign n1575 = ( ~n1271 & n1573 ) | ( ~n1271 & n1574 ) | ( n1573 & n1574 ) ;
  assign n1576 = ( x382 & x383 ) | ( x382 & x384 ) | ( x383 & x384 ) ;
  assign n1577 = ( x379 & x380 ) | ( x379 & x381 ) | ( x380 & x381 ) ;
  assign n1578 = ( x379 & ~x380 ) | ( x379 & x381 ) | ( ~x380 & x381 ) ;
  assign n1579 = ( ~x379 & x380 ) | ( ~x379 & n1578 ) | ( x380 & n1578 ) ;
  assign n1580 = ( ~x381 & n1578 ) | ( ~x381 & n1579 ) | ( n1578 & n1579 ) ;
  assign n1581 = ( x382 & ~x383 ) | ( x382 & x384 ) | ( ~x383 & x384 ) ;
  assign n1582 = ( ~x382 & x383 ) | ( ~x382 & n1581 ) | ( x383 & n1581 ) ;
  assign n1583 = ( ~x384 & n1581 ) | ( ~x384 & n1582 ) | ( n1581 & n1582 ) ;
  assign n1584 = n1580 & n1583 ;
  assign n1585 = ( n1576 & n1577 ) | ( n1576 & n1584 ) | ( n1577 & n1584 ) ;
  assign n1586 = ( x388 & x389 ) | ( x388 & x390 ) | ( x389 & x390 ) ;
  assign n1587 = ( x385 & x386 ) | ( x385 & x387 ) | ( x386 & x387 ) ;
  assign n1588 = ( x385 & ~x386 ) | ( x385 & x387 ) | ( ~x386 & x387 ) ;
  assign n1589 = ( ~x385 & x386 ) | ( ~x385 & n1588 ) | ( x386 & n1588 ) ;
  assign n1590 = ( ~x387 & n1588 ) | ( ~x387 & n1589 ) | ( n1588 & n1589 ) ;
  assign n1591 = ( x388 & ~x389 ) | ( x388 & x390 ) | ( ~x389 & x390 ) ;
  assign n1592 = ( ~x388 & x389 ) | ( ~x388 & n1591 ) | ( x389 & n1591 ) ;
  assign n1593 = ( ~x390 & n1591 ) | ( ~x390 & n1592 ) | ( n1591 & n1592 ) ;
  assign n1594 = n1590 & n1593 ;
  assign n1595 = ( n1586 & n1587 ) | ( n1586 & n1594 ) | ( n1587 & n1594 ) ;
  assign n1596 = ( n1577 & n1584 ) | ( n1577 & ~n1585 ) | ( n1584 & ~n1585 ) ;
  assign n1597 = ( n1576 & ~n1585 ) | ( n1576 & n1596 ) | ( ~n1585 & n1596 ) ;
  assign n1598 = ( n1587 & n1594 ) | ( n1587 & ~n1595 ) | ( n1594 & ~n1595 ) ;
  assign n1599 = ( n1586 & ~n1595 ) | ( n1586 & n1598 ) | ( ~n1595 & n1598 ) ;
  assign n1600 = n1585 & n1597 ;
  assign n1601 = n1580 & ~n1583 ;
  assign n1602 = ~n1580 & n1583 ;
  assign n1603 = n1601 | n1602 ;
  assign n1604 = n1590 & ~n1593 ;
  assign n1605 = ~n1590 & n1593 ;
  assign n1606 = n1604 | n1605 ;
  assign n1607 = n1603 & n1606 ;
  assign n1608 = ~n1600 & n1607 ;
  assign n1609 = ( n1597 & n1599 ) | ( n1597 & n1608 ) | ( n1599 & n1608 ) ;
  assign n1610 = ( n1585 & n1595 ) | ( n1585 & n1609 ) | ( n1595 & n1609 ) ;
  assign n1611 = ( x370 & x371 ) | ( x370 & x372 ) | ( x371 & x372 ) ;
  assign n1612 = ( x367 & x368 ) | ( x367 & x369 ) | ( x368 & x369 ) ;
  assign n1613 = ( x367 & ~x368 ) | ( x367 & x369 ) | ( ~x368 & x369 ) ;
  assign n1614 = ( ~x367 & x368 ) | ( ~x367 & n1613 ) | ( x368 & n1613 ) ;
  assign n1615 = ( ~x369 & n1613 ) | ( ~x369 & n1614 ) | ( n1613 & n1614 ) ;
  assign n1616 = ( x370 & ~x371 ) | ( x370 & x372 ) | ( ~x371 & x372 ) ;
  assign n1617 = ( ~x370 & x371 ) | ( ~x370 & n1616 ) | ( x371 & n1616 ) ;
  assign n1618 = ( ~x372 & n1616 ) | ( ~x372 & n1617 ) | ( n1616 & n1617 ) ;
  assign n1619 = n1615 & n1618 ;
  assign n1620 = ( n1611 & n1612 ) | ( n1611 & n1619 ) | ( n1612 & n1619 ) ;
  assign n1621 = ( x376 & x377 ) | ( x376 & x378 ) | ( x377 & x378 ) ;
  assign n1622 = ( x373 & x374 ) | ( x373 & x375 ) | ( x374 & x375 ) ;
  assign n1623 = ( x373 & ~x374 ) | ( x373 & x375 ) | ( ~x374 & x375 ) ;
  assign n1624 = ( ~x373 & x374 ) | ( ~x373 & n1623 ) | ( x374 & n1623 ) ;
  assign n1625 = ( ~x375 & n1623 ) | ( ~x375 & n1624 ) | ( n1623 & n1624 ) ;
  assign n1626 = ( x376 & ~x377 ) | ( x376 & x378 ) | ( ~x377 & x378 ) ;
  assign n1627 = ( ~x376 & x377 ) | ( ~x376 & n1626 ) | ( x377 & n1626 ) ;
  assign n1628 = ( ~x378 & n1626 ) | ( ~x378 & n1627 ) | ( n1626 & n1627 ) ;
  assign n1629 = n1625 & n1628 ;
  assign n1630 = ( n1621 & n1622 ) | ( n1621 & n1629 ) | ( n1622 & n1629 ) ;
  assign n1631 = ( n1612 & n1619 ) | ( n1612 & ~n1620 ) | ( n1619 & ~n1620 ) ;
  assign n1632 = ( n1611 & ~n1620 ) | ( n1611 & n1631 ) | ( ~n1620 & n1631 ) ;
  assign n1633 = n1620 & n1632 ;
  assign n1634 = ( n1622 & n1629 ) | ( n1622 & ~n1630 ) | ( n1629 & ~n1630 ) ;
  assign n1635 = ( n1621 & ~n1630 ) | ( n1621 & n1634 ) | ( ~n1630 & n1634 ) ;
  assign n1636 = n1630 & n1635 ;
  assign n1637 = n1615 & ~n1618 ;
  assign n1638 = ~n1615 & n1618 ;
  assign n1639 = n1637 | n1638 ;
  assign n1640 = n1625 & ~n1628 ;
  assign n1641 = ~n1625 & n1628 ;
  assign n1642 = n1640 | n1641 ;
  assign n1643 = n1639 & n1642 ;
  assign n1644 = ~n1636 & n1643 ;
  assign n1645 = n1635 & n1644 ;
  assign n1646 = ~n1633 & n1645 ;
  assign n1647 = ~n1633 & n1644 ;
  assign n1648 = ~n1635 & n1647 ;
  assign n1649 = ( n1632 & n1635 ) | ( n1632 & n1648 ) | ( n1635 & n1648 ) ;
  assign n1650 = n1646 | n1649 ;
  assign n1651 = ( n1620 & n1630 ) | ( n1620 & n1650 ) | ( n1630 & n1650 ) ;
  assign n1652 = n1610 & n1651 ;
  assign n1653 = n1651 & ~n1652 ;
  assign n1654 = ( n1610 & ~n1652 ) | ( n1610 & n1653 ) | ( ~n1652 & n1653 ) ;
  assign n1655 = n1652 | n1654 ;
  assign n1656 = ( n1632 & n1635 ) | ( n1632 & ~n1647 ) | ( n1635 & ~n1647 ) ;
  assign n1657 = n1632 & ~n1646 ;
  assign n1658 = ( n1635 & ~n1656 ) | ( n1635 & n1657 ) | ( ~n1656 & n1657 ) ;
  assign n1659 = ( n1648 & n1656 ) | ( n1648 & ~n1658 ) | ( n1656 & ~n1658 ) ;
  assign n1660 = n1603 & ~n1606 ;
  assign n1661 = ~n1603 & n1606 ;
  assign n1662 = n1660 | n1661 ;
  assign n1663 = n1639 & ~n1642 ;
  assign n1664 = ~n1639 & n1642 ;
  assign n1665 = n1663 | n1664 ;
  assign n1666 = n1662 & n1665 ;
  assign n1667 = n1599 & n1607 ;
  assign n1668 = n1599 | n1608 ;
  assign n1669 = ( n1597 & n1667 ) | ( n1597 & ~n1668 ) | ( n1667 & ~n1668 ) ;
  assign n1670 = ~n1609 & n1668 ;
  assign n1671 = n1669 | n1670 ;
  assign n1672 = n1666 | n1671 ;
  assign n1673 = n1659 & n1672 ;
  assign n1674 = ( n1666 & n1669 ) | ( n1666 & n1670 ) | ( n1669 & n1670 ) ;
  assign n1675 = n1673 | n1674 ;
  assign n1676 = ~n1620 & n1630 ;
  assign n1677 = n1620 & ~n1630 ;
  assign n1678 = n1676 | n1677 ;
  assign n1679 = n1646 | n1678 ;
  assign n1680 = n1649 | n1679 ;
  assign n1681 = n1650 & n1678 ;
  assign n1682 = n1680 & ~n1681 ;
  assign n1683 = ~n1585 & n1595 ;
  assign n1684 = n1585 & ~n1595 ;
  assign n1685 = n1683 | n1684 ;
  assign n1686 = n1609 & n1685 ;
  assign n1687 = n1609 | n1685 ;
  assign n1688 = ~n1686 & n1687 ;
  assign n1689 = ( n1675 & n1682 ) | ( n1675 & n1688 ) | ( n1682 & n1688 ) ;
  assign n1690 = ( n1652 & n1655 ) | ( n1652 & n1689 ) | ( n1655 & n1689 ) ;
  assign n1691 = ( x403 & ~x404 ) | ( x403 & x405 ) | ( ~x404 & x405 ) ;
  assign n1692 = ( ~x403 & x404 ) | ( ~x403 & n1691 ) | ( x404 & n1691 ) ;
  assign n1693 = ( ~x405 & n1691 ) | ( ~x405 & n1692 ) | ( n1691 & n1692 ) ;
  assign n1694 = ( x406 & ~x407 ) | ( x406 & x408 ) | ( ~x407 & x408 ) ;
  assign n1695 = ( ~x406 & x407 ) | ( ~x406 & n1694 ) | ( x407 & n1694 ) ;
  assign n1696 = ( ~x408 & n1694 ) | ( ~x408 & n1695 ) | ( n1694 & n1695 ) ;
  assign n1697 = n1693 & n1696 ;
  assign n1698 = ( x406 & x407 ) | ( x406 & x408 ) | ( x407 & x408 ) ;
  assign n1699 = ( x403 & x404 ) | ( x403 & x405 ) | ( x404 & x405 ) ;
  assign n1700 = ( n1697 & n1698 ) | ( n1697 & n1699 ) | ( n1698 & n1699 ) ;
  assign n1701 = ( x412 & x413 ) | ( x412 & x414 ) | ( x413 & x414 ) ;
  assign n1702 = ( x409 & x410 ) | ( x409 & x411 ) | ( x410 & x411 ) ;
  assign n1703 = ( x409 & ~x410 ) | ( x409 & x411 ) | ( ~x410 & x411 ) ;
  assign n1704 = ( ~x409 & x410 ) | ( ~x409 & n1703 ) | ( x410 & n1703 ) ;
  assign n1705 = ( ~x411 & n1703 ) | ( ~x411 & n1704 ) | ( n1703 & n1704 ) ;
  assign n1706 = ( x412 & ~x413 ) | ( x412 & x414 ) | ( ~x413 & x414 ) ;
  assign n1707 = ( ~x412 & x413 ) | ( ~x412 & n1706 ) | ( x413 & n1706 ) ;
  assign n1708 = ( ~x414 & n1706 ) | ( ~x414 & n1707 ) | ( n1706 & n1707 ) ;
  assign n1709 = n1705 & n1708 ;
  assign n1710 = ( n1701 & n1702 ) | ( n1701 & n1709 ) | ( n1702 & n1709 ) ;
  assign n1711 = ( n1697 & n1699 ) | ( n1697 & ~n1700 ) | ( n1699 & ~n1700 ) ;
  assign n1712 = ( n1698 & ~n1700 ) | ( n1698 & n1711 ) | ( ~n1700 & n1711 ) ;
  assign n1713 = ( n1702 & n1709 ) | ( n1702 & ~n1710 ) | ( n1709 & ~n1710 ) ;
  assign n1714 = ( n1701 & ~n1710 ) | ( n1701 & n1713 ) | ( ~n1710 & n1713 ) ;
  assign n1715 = n1700 & n1712 ;
  assign n1716 = n1693 & ~n1696 ;
  assign n1717 = ~n1693 & n1696 ;
  assign n1718 = n1716 | n1717 ;
  assign n1719 = n1705 & ~n1708 ;
  assign n1720 = ~n1705 & n1708 ;
  assign n1721 = n1719 | n1720 ;
  assign n1722 = n1718 & n1721 ;
  assign n1723 = ~n1715 & n1722 ;
  assign n1724 = ( n1712 & n1714 ) | ( n1712 & n1723 ) | ( n1714 & n1723 ) ;
  assign n1725 = ( n1700 & n1710 ) | ( n1700 & n1724 ) | ( n1710 & n1724 ) ;
  assign n1726 = ( x391 & ~x392 ) | ( x391 & x393 ) | ( ~x392 & x393 ) ;
  assign n1727 = ( ~x391 & x392 ) | ( ~x391 & n1726 ) | ( x392 & n1726 ) ;
  assign n1728 = ( ~x393 & n1726 ) | ( ~x393 & n1727 ) | ( n1726 & n1727 ) ;
  assign n1729 = ( x394 & ~x395 ) | ( x394 & x396 ) | ( ~x395 & x396 ) ;
  assign n1730 = ( ~x394 & x395 ) | ( ~x394 & n1729 ) | ( x395 & n1729 ) ;
  assign n1731 = ( ~x396 & n1729 ) | ( ~x396 & n1730 ) | ( n1729 & n1730 ) ;
  assign n1732 = n1728 & n1731 ;
  assign n1733 = ( x394 & x395 ) | ( x394 & x396 ) | ( x395 & x396 ) ;
  assign n1734 = ( x391 & x392 ) | ( x391 & x393 ) | ( x392 & x393 ) ;
  assign n1735 = ( n1732 & n1733 ) | ( n1732 & n1734 ) | ( n1733 & n1734 ) ;
  assign n1736 = ( x400 & x401 ) | ( x400 & x402 ) | ( x401 & x402 ) ;
  assign n1737 = ( x397 & x398 ) | ( x397 & x399 ) | ( x398 & x399 ) ;
  assign n1738 = ( x397 & ~x398 ) | ( x397 & x399 ) | ( ~x398 & x399 ) ;
  assign n1739 = ( ~x397 & x398 ) | ( ~x397 & n1738 ) | ( x398 & n1738 ) ;
  assign n1740 = ( ~x399 & n1738 ) | ( ~x399 & n1739 ) | ( n1738 & n1739 ) ;
  assign n1741 = ( x400 & ~x401 ) | ( x400 & x402 ) | ( ~x401 & x402 ) ;
  assign n1742 = ( ~x400 & x401 ) | ( ~x400 & n1741 ) | ( x401 & n1741 ) ;
  assign n1743 = ( ~x402 & n1741 ) | ( ~x402 & n1742 ) | ( n1741 & n1742 ) ;
  assign n1744 = n1740 & n1743 ;
  assign n1745 = ( n1736 & n1737 ) | ( n1736 & n1744 ) | ( n1737 & n1744 ) ;
  assign n1746 = ( n1732 & n1734 ) | ( n1732 & ~n1735 ) | ( n1734 & ~n1735 ) ;
  assign n1747 = ( n1733 & ~n1735 ) | ( n1733 & n1746 ) | ( ~n1735 & n1746 ) ;
  assign n1748 = n1735 & n1747 ;
  assign n1749 = ( n1737 & n1744 ) | ( n1737 & ~n1745 ) | ( n1744 & ~n1745 ) ;
  assign n1750 = ( n1736 & ~n1745 ) | ( n1736 & n1749 ) | ( ~n1745 & n1749 ) ;
  assign n1751 = n1745 & n1750 ;
  assign n1752 = n1728 & ~n1731 ;
  assign n1753 = ~n1728 & n1731 ;
  assign n1754 = n1752 | n1753 ;
  assign n1755 = n1740 & ~n1743 ;
  assign n1756 = ~n1740 & n1743 ;
  assign n1757 = n1755 | n1756 ;
  assign n1758 = n1754 & n1757 ;
  assign n1759 = ~n1751 & n1758 ;
  assign n1760 = n1750 & n1759 ;
  assign n1761 = ~n1748 & n1760 ;
  assign n1762 = ~n1748 & n1759 ;
  assign n1763 = ~n1750 & n1762 ;
  assign n1764 = ( n1747 & n1750 ) | ( n1747 & n1763 ) | ( n1750 & n1763 ) ;
  assign n1765 = n1761 | n1764 ;
  assign n1766 = ( n1735 & n1745 ) | ( n1735 & n1765 ) | ( n1745 & n1765 ) ;
  assign n1767 = ~n1735 & n1745 ;
  assign n1768 = n1735 & ~n1745 ;
  assign n1769 = n1767 | n1768 ;
  assign n1770 = n1761 | n1769 ;
  assign n1771 = n1764 | n1770 ;
  assign n1772 = n1765 & n1769 ;
  assign n1773 = n1771 & ~n1772 ;
  assign n1774 = ( n1700 & n1710 ) | ( n1700 & ~n1724 ) | ( n1710 & ~n1724 ) ;
  assign n1775 = ( ~n1700 & n1710 ) | ( ~n1700 & n1724 ) | ( n1710 & n1724 ) ;
  assign n1776 = ( ~n1710 & n1774 ) | ( ~n1710 & n1775 ) | ( n1774 & n1775 ) ;
  assign n1777 = n1773 | n1776 ;
  assign n1778 = ( n1747 & n1750 ) | ( n1747 & ~n1762 ) | ( n1750 & ~n1762 ) ;
  assign n1779 = n1747 & ~n1761 ;
  assign n1780 = ( n1750 & ~n1778 ) | ( n1750 & n1779 ) | ( ~n1778 & n1779 ) ;
  assign n1781 = ( n1763 & n1778 ) | ( n1763 & ~n1780 ) | ( n1778 & ~n1780 ) ;
  assign n1782 = n1718 & ~n1721 ;
  assign n1783 = ~n1718 & n1721 ;
  assign n1784 = n1782 | n1783 ;
  assign n1785 = n1754 & ~n1757 ;
  assign n1786 = ~n1754 & n1757 ;
  assign n1787 = n1785 | n1786 ;
  assign n1788 = n1784 & n1787 ;
  assign n1789 = n1714 | n1723 ;
  assign n1790 = ~n1724 & n1789 ;
  assign n1791 = n1714 & n1722 ;
  assign n1792 = ( n1712 & ~n1789 ) | ( n1712 & n1791 ) | ( ~n1789 & n1791 ) ;
  assign n1793 = n1790 | n1792 ;
  assign n1794 = n1788 | n1793 ;
  assign n1795 = ( n1788 & n1790 ) | ( n1788 & n1792 ) | ( n1790 & n1792 ) ;
  assign n1796 = ( n1781 & n1794 ) | ( n1781 & n1795 ) | ( n1794 & n1795 ) ;
  assign n1797 = n1777 & n1796 ;
  assign n1798 = n1773 & n1776 ;
  assign n1799 = n1797 | n1798 ;
  assign n1800 = ( n1725 & n1766 ) | ( n1725 & n1799 ) | ( n1766 & n1799 ) ;
  assign n1801 = n1690 & n1800 ;
  assign n1802 = n1800 & ~n1801 ;
  assign n1803 = ( n1690 & ~n1801 ) | ( n1690 & n1802 ) | ( ~n1801 & n1802 ) ;
  assign n1804 = ~n1725 & n1766 ;
  assign n1805 = n1725 & ~n1766 ;
  assign n1806 = n1804 | n1805 ;
  assign n1807 = n1798 | n1806 ;
  assign n1808 = n1797 | n1807 ;
  assign n1809 = n1799 & n1806 ;
  assign n1810 = n1808 & ~n1809 ;
  assign n1811 = n1654 | n1689 ;
  assign n1812 = ~n1654 & n1811 ;
  assign n1813 = ( ~n1689 & n1811 ) | ( ~n1689 & n1812 ) | ( n1811 & n1812 ) ;
  assign n1814 = ( n1675 & ~n1682 ) | ( n1675 & n1688 ) | ( ~n1682 & n1688 ) ;
  assign n1815 = ( ~n1675 & n1682 ) | ( ~n1675 & n1814 ) | ( n1682 & n1814 ) ;
  assign n1816 = ( ~n1688 & n1814 ) | ( ~n1688 & n1815 ) | ( n1814 & n1815 ) ;
  assign n1817 = ( ~n1773 & n1776 ) | ( ~n1773 & n1796 ) | ( n1776 & n1796 ) ;
  assign n1818 = ( n1773 & ~n1796 ) | ( n1773 & n1817 ) | ( ~n1796 & n1817 ) ;
  assign n1819 = ( ~n1776 & n1817 ) | ( ~n1776 & n1818 ) | ( n1817 & n1818 ) ;
  assign n1820 = n1784 & ~n1787 ;
  assign n1821 = ~n1784 & n1787 ;
  assign n1822 = n1820 | n1821 ;
  assign n1823 = n1662 & ~n1665 ;
  assign n1824 = ~n1662 & n1665 ;
  assign n1825 = n1823 | n1824 ;
  assign n1826 = n1822 & n1825 ;
  assign n1827 = ~n1788 & n1794 ;
  assign n1828 = ( ~n1793 & n1794 ) | ( ~n1793 & n1827 ) | ( n1794 & n1827 ) ;
  assign n1829 = n1781 & ~n1828 ;
  assign n1830 = ~n1781 & n1828 ;
  assign n1831 = n1829 | n1830 ;
  assign n1832 = ( n1659 & n1666 ) | ( n1659 & ~n1671 ) | ( n1666 & ~n1671 ) ;
  assign n1833 = ( ~n1659 & n1671 ) | ( ~n1659 & n1832 ) | ( n1671 & n1832 ) ;
  assign n1834 = ( ~n1666 & n1832 ) | ( ~n1666 & n1833 ) | ( n1832 & n1833 ) ;
  assign n1835 = ( n1826 & n1831 ) | ( n1826 & n1834 ) | ( n1831 & n1834 ) ;
  assign n1836 = ( n1816 & n1819 ) | ( n1816 & n1835 ) | ( n1819 & n1835 ) ;
  assign n1837 = ( n1810 & n1813 ) | ( n1810 & n1836 ) | ( n1813 & n1836 ) ;
  assign n1838 = n1803 & n1837 ;
  assign n1839 = n1803 | n1837 ;
  assign n1840 = ~n1838 & n1839 ;
  assign n1841 = ( x442 & x443 ) | ( x442 & x444 ) | ( x443 & x444 ) ;
  assign n1842 = ( x439 & ~x440 ) | ( x439 & x441 ) | ( ~x440 & x441 ) ;
  assign n1843 = ( ~x439 & x440 ) | ( ~x439 & n1842 ) | ( x440 & n1842 ) ;
  assign n1844 = ( ~x441 & n1842 ) | ( ~x441 & n1843 ) | ( n1842 & n1843 ) ;
  assign n1845 = ( x442 & ~x443 ) | ( x442 & x444 ) | ( ~x443 & x444 ) ;
  assign n1846 = ( ~x442 & x443 ) | ( ~x442 & n1845 ) | ( x443 & n1845 ) ;
  assign n1847 = ( ~x444 & n1845 ) | ( ~x444 & n1846 ) | ( n1845 & n1846 ) ;
  assign n1848 = n1844 & n1847 ;
  assign n1849 = ( x439 & x440 ) | ( x439 & x441 ) | ( x440 & x441 ) ;
  assign n1850 = ( n1841 & n1848 ) | ( n1841 & n1849 ) | ( n1848 & n1849 ) ;
  assign n1851 = ( n1848 & n1849 ) | ( n1848 & ~n1850 ) | ( n1849 & ~n1850 ) ;
  assign n1852 = ( n1841 & ~n1850 ) | ( n1841 & n1851 ) | ( ~n1850 & n1851 ) ;
  assign n1853 = ( x448 & x449 ) | ( x448 & x450 ) | ( x449 & x450 ) ;
  assign n1854 = ( x445 & x446 ) | ( x445 & x447 ) | ( x446 & x447 ) ;
  assign n1855 = ( x445 & ~x446 ) | ( x445 & x447 ) | ( ~x446 & x447 ) ;
  assign n1856 = ( ~x445 & x446 ) | ( ~x445 & n1855 ) | ( x446 & n1855 ) ;
  assign n1857 = ( ~x447 & n1855 ) | ( ~x447 & n1856 ) | ( n1855 & n1856 ) ;
  assign n1858 = ( x448 & ~x449 ) | ( x448 & x450 ) | ( ~x449 & x450 ) ;
  assign n1859 = ( ~x448 & x449 ) | ( ~x448 & n1858 ) | ( x449 & n1858 ) ;
  assign n1860 = ( ~x450 & n1858 ) | ( ~x450 & n1859 ) | ( n1858 & n1859 ) ;
  assign n1861 = n1857 & n1860 ;
  assign n1862 = ( n1853 & n1854 ) | ( n1853 & n1861 ) | ( n1854 & n1861 ) ;
  assign n1863 = ( n1854 & n1861 ) | ( n1854 & ~n1862 ) | ( n1861 & ~n1862 ) ;
  assign n1864 = ( n1853 & ~n1862 ) | ( n1853 & n1863 ) | ( ~n1862 & n1863 ) ;
  assign n1865 = n1850 & n1852 ;
  assign n1866 = n1862 & n1864 ;
  assign n1867 = n1844 & ~n1847 ;
  assign n1868 = ~n1844 & n1847 ;
  assign n1869 = n1867 | n1868 ;
  assign n1870 = n1857 & ~n1860 ;
  assign n1871 = ~n1857 & n1860 ;
  assign n1872 = n1870 | n1871 ;
  assign n1873 = n1869 & n1872 ;
  assign n1874 = ~n1866 & n1873 ;
  assign n1875 = ~n1865 & n1874 ;
  assign n1876 = ~n1864 & n1875 ;
  assign n1877 = ( n1852 & n1864 ) | ( n1852 & n1876 ) | ( n1864 & n1876 ) ;
  assign n1878 = n1864 & n1874 ;
  assign n1879 = ~n1865 & n1878 ;
  assign n1880 = ~n1850 & n1862 ;
  assign n1881 = n1850 & ~n1862 ;
  assign n1882 = n1880 | n1881 ;
  assign n1883 = n1879 | n1882 ;
  assign n1884 = n1877 | n1883 ;
  assign n1885 = n1877 | n1879 ;
  assign n1886 = n1882 & n1885 ;
  assign n1887 = n1884 & ~n1886 ;
  assign n1888 = ( x460 & x461 ) | ( x460 & x462 ) | ( x461 & x462 ) ;
  assign n1889 = ( x457 & x458 ) | ( x457 & x459 ) | ( x458 & x459 ) ;
  assign n1890 = ( x457 & ~x458 ) | ( x457 & x459 ) | ( ~x458 & x459 ) ;
  assign n1891 = ( ~x457 & x458 ) | ( ~x457 & n1890 ) | ( x458 & n1890 ) ;
  assign n1892 = ( ~x459 & n1890 ) | ( ~x459 & n1891 ) | ( n1890 & n1891 ) ;
  assign n1893 = ( x460 & ~x461 ) | ( x460 & x462 ) | ( ~x461 & x462 ) ;
  assign n1894 = ( ~x460 & x461 ) | ( ~x460 & n1893 ) | ( x461 & n1893 ) ;
  assign n1895 = ( ~x462 & n1893 ) | ( ~x462 & n1894 ) | ( n1893 & n1894 ) ;
  assign n1896 = n1892 & n1895 ;
  assign n1897 = ( n1888 & n1889 ) | ( n1888 & n1896 ) | ( n1889 & n1896 ) ;
  assign n1898 = ( x451 & ~x452 ) | ( x451 & x453 ) | ( ~x452 & x453 ) ;
  assign n1899 = ( ~x451 & x452 ) | ( ~x451 & n1898 ) | ( x452 & n1898 ) ;
  assign n1900 = ( ~x453 & n1898 ) | ( ~x453 & n1899 ) | ( n1898 & n1899 ) ;
  assign n1901 = ( x454 & ~x455 ) | ( x454 & x456 ) | ( ~x455 & x456 ) ;
  assign n1902 = ( ~x454 & x455 ) | ( ~x454 & n1901 ) | ( x455 & n1901 ) ;
  assign n1903 = ( ~x456 & n1901 ) | ( ~x456 & n1902 ) | ( n1901 & n1902 ) ;
  assign n1904 = n1900 & n1903 ;
  assign n1905 = ( x454 & x455 ) | ( x454 & x456 ) | ( x455 & x456 ) ;
  assign n1906 = ( x451 & x452 ) | ( x451 & x453 ) | ( x452 & x453 ) ;
  assign n1907 = ( n1904 & n1905 ) | ( n1904 & n1906 ) | ( n1905 & n1906 ) ;
  assign n1908 = ( n1889 & n1896 ) | ( n1889 & ~n1897 ) | ( n1896 & ~n1897 ) ;
  assign n1909 = ( n1888 & ~n1897 ) | ( n1888 & n1908 ) | ( ~n1897 & n1908 ) ;
  assign n1910 = ( n1904 & n1906 ) | ( n1904 & ~n1907 ) | ( n1906 & ~n1907 ) ;
  assign n1911 = ( n1905 & ~n1907 ) | ( n1905 & n1910 ) | ( ~n1907 & n1910 ) ;
  assign n1912 = n1907 & n1911 ;
  assign n1913 = n1900 & ~n1903 ;
  assign n1914 = ~n1900 & n1903 ;
  assign n1915 = n1913 | n1914 ;
  assign n1916 = n1892 & ~n1895 ;
  assign n1917 = ~n1892 & n1895 ;
  assign n1918 = n1916 | n1917 ;
  assign n1919 = ~n1896 & n1918 ;
  assign n1920 = n1915 & n1919 ;
  assign n1921 = ~n1912 & n1920 ;
  assign n1922 = ( n1909 & n1911 ) | ( n1909 & n1921 ) | ( n1911 & n1921 ) ;
  assign n1923 = ( n1897 & n1907 ) | ( n1897 & ~n1922 ) | ( n1907 & ~n1922 ) ;
  assign n1924 = ( n1897 & ~n1907 ) | ( n1897 & n1922 ) | ( ~n1907 & n1922 ) ;
  assign n1925 = ( ~n1897 & n1923 ) | ( ~n1897 & n1924 ) | ( n1923 & n1924 ) ;
  assign n1926 = n1887 | n1925 ;
  assign n1927 = ( n1852 & n1864 ) | ( n1852 & ~n1875 ) | ( n1864 & ~n1875 ) ;
  assign n1928 = n1852 & ~n1879 ;
  assign n1929 = ( n1864 & ~n1927 ) | ( n1864 & n1928 ) | ( ~n1927 & n1928 ) ;
  assign n1930 = ( n1876 & n1927 ) | ( n1876 & ~n1929 ) | ( n1927 & ~n1929 ) ;
  assign n1931 = n1915 & ~n1919 ;
  assign n1932 = ~n1915 & n1919 ;
  assign n1933 = n1931 | n1932 ;
  assign n1934 = n1869 & ~n1872 ;
  assign n1935 = ~n1869 & n1872 ;
  assign n1936 = n1934 | n1935 ;
  assign n1937 = n1933 & n1936 ;
  assign n1938 = n1909 | n1921 ;
  assign n1939 = ~n1922 & n1938 ;
  assign n1940 = n1909 & n1920 ;
  assign n1941 = ( n1911 & ~n1938 ) | ( n1911 & n1940 ) | ( ~n1938 & n1940 ) ;
  assign n1942 = n1939 | n1941 ;
  assign n1943 = n1937 | n1942 ;
  assign n1944 = ( n1937 & n1939 ) | ( n1937 & n1941 ) | ( n1939 & n1941 ) ;
  assign n1945 = ( n1930 & n1943 ) | ( n1930 & n1944 ) | ( n1943 & n1944 ) ;
  assign n1946 = n1926 & n1945 ;
  assign n1947 = n1887 & n1925 ;
  assign n1948 = n1946 | n1947 ;
  assign n1949 = ( n1897 & n1907 ) | ( n1897 & n1922 ) | ( n1907 & n1922 ) ;
  assign n1950 = ( n1850 & n1862 ) | ( n1850 & n1885 ) | ( n1862 & n1885 ) ;
  assign n1951 = n1949 & n1950 ;
  assign n1952 = n1950 & ~n1951 ;
  assign n1953 = ( n1949 & ~n1951 ) | ( n1949 & n1952 ) | ( ~n1951 & n1952 ) ;
  assign n1954 = n1948 & n1953 ;
  assign n1955 = n1947 | n1953 ;
  assign n1956 = n1946 | n1955 ;
  assign n1957 = ~n1954 & n1956 ;
  assign n2005 = ( x424 & x425 ) | ( x424 & x426 ) | ( x425 & x426 ) ;
  assign n2006 = ( x421 & x422 ) | ( x421 & x423 ) | ( x422 & x423 ) ;
  assign n2007 = ( x421 & ~x422 ) | ( x421 & x423 ) | ( ~x422 & x423 ) ;
  assign n2008 = ( ~x421 & x422 ) | ( ~x421 & n2007 ) | ( x422 & n2007 ) ;
  assign n2009 = ( ~x423 & n2007 ) | ( ~x423 & n2008 ) | ( n2007 & n2008 ) ;
  assign n2010 = ( x424 & ~x425 ) | ( x424 & x426 ) | ( ~x425 & x426 ) ;
  assign n2011 = ( ~x424 & x425 ) | ( ~x424 & n2010 ) | ( x425 & n2010 ) ;
  assign n2012 = ( ~x426 & n2010 ) | ( ~x426 & n2011 ) | ( n2010 & n2011 ) ;
  assign n2013 = n2009 & n2012 ;
  assign n2014 = ( n2005 & n2006 ) | ( n2005 & n2013 ) | ( n2006 & n2013 ) ;
  assign n2015 = ( n2006 & n2013 ) | ( n2006 & ~n2014 ) | ( n2013 & ~n2014 ) ;
  assign n2016 = ( n2005 & ~n2014 ) | ( n2005 & n2015 ) | ( ~n2014 & n2015 ) ;
  assign n1995 = ( x418 & x419 ) | ( x418 & x420 ) | ( x419 & x420 ) ;
  assign n1996 = ( x415 & x416 ) | ( x415 & x417 ) | ( x416 & x417 ) ;
  assign n1997 = ( x415 & ~x416 ) | ( x415 & x417 ) | ( ~x416 & x417 ) ;
  assign n1998 = ( ~x415 & x416 ) | ( ~x415 & n1997 ) | ( x416 & n1997 ) ;
  assign n1999 = ( ~x417 & n1997 ) | ( ~x417 & n1998 ) | ( n1997 & n1998 ) ;
  assign n2000 = ( x418 & ~x419 ) | ( x418 & x420 ) | ( ~x419 & x420 ) ;
  assign n2001 = ( ~x418 & x419 ) | ( ~x418 & n2000 ) | ( x419 & n2000 ) ;
  assign n2002 = ( ~x420 & n2000 ) | ( ~x420 & n2001 ) | ( n2000 & n2001 ) ;
  assign n2003 = n1999 & n2002 ;
  assign n2004 = ( n1995 & n1996 ) | ( n1995 & n2003 ) | ( n1996 & n2003 ) ;
  assign n2017 = ( n1996 & n2003 ) | ( n1996 & ~n2004 ) | ( n2003 & ~n2004 ) ;
  assign n2018 = ( n1995 & ~n2004 ) | ( n1995 & n2017 ) | ( ~n2004 & n2017 ) ;
  assign n2019 = n2004 & n2018 ;
  assign n2020 = n2014 & n2016 ;
  assign n2021 = n2009 & ~n2012 ;
  assign n2022 = ~n2009 & n2012 ;
  assign n2023 = n2021 | n2022 ;
  assign n2024 = n1999 & ~n2002 ;
  assign n2025 = ~n1999 & n2002 ;
  assign n2026 = n2024 | n2025 ;
  assign n2027 = n2023 & n2026 ;
  assign n2028 = ~n2020 & n2027 ;
  assign n2029 = ~n2019 & n2028 ;
  assign n2031 = ~n2016 & n2029 ;
  assign n2038 = ( n2016 & n2018 ) | ( n2016 & ~n2029 ) | ( n2018 & ~n2029 ) ;
  assign n2030 = n2016 & n2029 ;
  assign n2039 = n2018 & ~n2030 ;
  assign n2040 = ( n2016 & ~n2038 ) | ( n2016 & n2039 ) | ( ~n2038 & n2039 ) ;
  assign n2041 = ( n2031 & n2038 ) | ( n2031 & ~n2040 ) | ( n2038 & ~n2040 ) ;
  assign n1960 = ( x433 & ~x434 ) | ( x433 & x435 ) | ( ~x434 & x435 ) ;
  assign n1961 = ( ~x433 & x434 ) | ( ~x433 & n1960 ) | ( x434 & n1960 ) ;
  assign n1962 = ( ~x435 & n1960 ) | ( ~x435 & n1961 ) | ( n1960 & n1961 ) ;
  assign n1963 = ( x436 & ~x437 ) | ( x436 & x438 ) | ( ~x437 & x438 ) ;
  assign n1964 = ( ~x436 & x437 ) | ( ~x436 & n1963 ) | ( x437 & n1963 ) ;
  assign n1965 = ( ~x438 & n1963 ) | ( ~x438 & n1964 ) | ( n1963 & n1964 ) ;
  assign n1984 = n1962 & ~n1965 ;
  assign n1985 = ~n1962 & n1965 ;
  assign n1986 = n1984 | n1985 ;
  assign n1968 = ( x427 & ~x428 ) | ( x427 & x429 ) | ( ~x428 & x429 ) ;
  assign n1969 = ( ~x427 & x428 ) | ( ~x427 & n1968 ) | ( x428 & n1968 ) ;
  assign n1970 = ( ~x429 & n1968 ) | ( ~x429 & n1969 ) | ( n1968 & n1969 ) ;
  assign n1971 = ( x430 & ~x431 ) | ( x430 & x432 ) | ( ~x431 & x432 ) ;
  assign n1972 = ( ~x430 & x431 ) | ( ~x430 & n1971 ) | ( x431 & n1971 ) ;
  assign n1973 = ( ~x432 & n1971 ) | ( ~x432 & n1972 ) | ( n1971 & n1972 ) ;
  assign n1987 = n1970 & ~n1973 ;
  assign n1988 = ~n1970 & n1973 ;
  assign n1989 = n1987 | n1988 ;
  assign n2042 = ~n1986 & n1989 ;
  assign n2043 = n1986 & ~n1989 ;
  assign n2044 = n2042 | n2043 ;
  assign n2045 = ~n2023 & n2026 ;
  assign n2046 = n2023 & ~n2026 ;
  assign n2047 = n2045 | n2046 ;
  assign n2048 = n2044 & n2047 ;
  assign n1975 = ( x430 & x431 ) | ( x430 & x432 ) | ( x431 & x432 ) ;
  assign n1974 = n1970 & n1973 ;
  assign n1976 = ( x427 & x428 ) | ( x427 & x429 ) | ( x428 & x429 ) ;
  assign n1977 = ( n1974 & n1975 ) | ( n1974 & n1976 ) | ( n1975 & n1976 ) ;
  assign n1980 = ( n1974 & n1976 ) | ( n1974 & ~n1977 ) | ( n1976 & ~n1977 ) ;
  assign n1981 = ( n1975 & ~n1977 ) | ( n1975 & n1980 ) | ( ~n1977 & n1980 ) ;
  assign n1958 = ( x436 & x437 ) | ( x436 & x438 ) | ( x437 & x438 ) ;
  assign n1959 = ( x433 & x434 ) | ( x433 & x435 ) | ( x434 & x435 ) ;
  assign n1966 = n1962 & n1965 ;
  assign n1967 = ( n1958 & n1959 ) | ( n1958 & n1966 ) | ( n1959 & n1966 ) ;
  assign n1978 = ( n1959 & n1966 ) | ( n1959 & ~n1967 ) | ( n1966 & ~n1967 ) ;
  assign n1979 = ( n1958 & ~n1967 ) | ( n1958 & n1978 ) | ( ~n1967 & n1978 ) ;
  assign n1983 = n1967 & n1979 ;
  assign n1990 = n1986 & n1989 ;
  assign n1991 = ~n1983 & n1990 ;
  assign n2049 = n1979 & n1991 ;
  assign n1982 = n1977 & n1981 ;
  assign n1992 = ~n1982 & n1991 ;
  assign n2050 = n1979 | n1992 ;
  assign n2051 = ( n1981 & n2049 ) | ( n1981 & ~n2050 ) | ( n2049 & ~n2050 ) ;
  assign n1993 = ( n1979 & n1981 ) | ( n1979 & n1992 ) | ( n1981 & n1992 ) ;
  assign n2052 = ~n1993 & n2050 ;
  assign n2053 = n2051 | n2052 ;
  assign n2054 = n2048 | n2053 ;
  assign n2055 = n2041 & n2054 ;
  assign n2056 = ( n2048 & n2051 ) | ( n2048 & n2052 ) | ( n2051 & n2052 ) ;
  assign n2057 = n2055 | n2056 ;
  assign n2032 = ( n2016 & n2018 ) | ( n2016 & n2031 ) | ( n2018 & n2031 ) ;
  assign n2058 = ~n2004 & n2014 ;
  assign n2059 = n2004 & ~n2014 ;
  assign n2060 = n2058 | n2059 ;
  assign n2061 = n2030 | n2060 ;
  assign n2062 = n2032 | n2061 ;
  assign n2033 = n2030 | n2032 ;
  assign n2063 = n2033 & n2060 ;
  assign n2064 = n2062 & ~n2063 ;
  assign n2065 = ( n1967 & n1977 ) | ( n1967 & ~n1993 ) | ( n1977 & ~n1993 ) ;
  assign n2066 = ( n1967 & ~n1977 ) | ( n1967 & n1993 ) | ( ~n1977 & n1993 ) ;
  assign n2067 = ( ~n1967 & n2065 ) | ( ~n1967 & n2066 ) | ( n2065 & n2066 ) ;
  assign n2068 = ( n2057 & n2064 ) | ( n2057 & n2067 ) | ( n2064 & n2067 ) ;
  assign n1994 = ( n1967 & n1977 ) | ( n1967 & n1993 ) | ( n1977 & n1993 ) ;
  assign n2034 = ( n2004 & n2014 ) | ( n2004 & n2033 ) | ( n2014 & n2033 ) ;
  assign n2035 = n1994 & n2034 ;
  assign n2036 = n1994 | n2034 ;
  assign n2037 = ~n2035 & n2036 ;
  assign n2069 = n2037 | n2068 ;
  assign n2070 = ~n2037 & n2069 ;
  assign n2071 = ( ~n2068 & n2069 ) | ( ~n2068 & n2070 ) | ( n2069 & n2070 ) ;
  assign n2072 = n1957 | n2071 ;
  assign n2073 = ( n2057 & ~n2064 ) | ( n2057 & n2067 ) | ( ~n2064 & n2067 ) ;
  assign n2074 = ( ~n2057 & n2064 ) | ( ~n2057 & n2073 ) | ( n2064 & n2073 ) ;
  assign n2075 = ( ~n2067 & n2073 ) | ( ~n2067 & n2074 ) | ( n2073 & n2074 ) ;
  assign n2076 = ( ~n1887 & n1925 ) | ( ~n1887 & n1945 ) | ( n1925 & n1945 ) ;
  assign n2077 = ( n1887 & ~n1945 ) | ( n1887 & n2076 ) | ( ~n1945 & n2076 ) ;
  assign n2078 = ( ~n1925 & n2076 ) | ( ~n1925 & n2077 ) | ( n2076 & n2077 ) ;
  assign n2079 = n1933 & ~n1936 ;
  assign n2080 = ~n1933 & n1936 ;
  assign n2081 = n2079 | n2080 ;
  assign n2082 = n2044 & ~n2047 ;
  assign n2083 = ~n2044 & n2047 ;
  assign n2084 = n2082 | n2083 ;
  assign n2085 = n2081 & n2084 ;
  assign n2086 = ~n1937 & n1943 ;
  assign n2087 = ( ~n1942 & n1943 ) | ( ~n1942 & n2086 ) | ( n1943 & n2086 ) ;
  assign n2088 = n1930 & ~n2087 ;
  assign n2089 = ~n1930 & n2087 ;
  assign n2090 = n2088 | n2089 ;
  assign n2091 = ( n2041 & n2048 ) | ( n2041 & ~n2053 ) | ( n2048 & ~n2053 ) ;
  assign n2092 = ( ~n2041 & n2053 ) | ( ~n2041 & n2091 ) | ( n2053 & n2091 ) ;
  assign n2093 = ( ~n2048 & n2091 ) | ( ~n2048 & n2092 ) | ( n2091 & n2092 ) ;
  assign n2094 = ( n2085 & n2090 ) | ( n2085 & n2093 ) | ( n2090 & n2093 ) ;
  assign n2095 = ( n2075 & n2078 ) | ( n2075 & n2094 ) | ( n2078 & n2094 ) ;
  assign n2096 = n2072 & n2095 ;
  assign n2097 = n1957 & n2071 ;
  assign n2098 = n2096 | n2097 ;
  assign n2099 = ( n2035 & n2036 ) | ( n2035 & n2068 ) | ( n2036 & n2068 ) ;
  assign n2100 = n1951 | n1954 ;
  assign n2101 = n2099 & n2100 ;
  assign n2102 = n2100 & ~n2101 ;
  assign n2103 = ( n2099 & ~n2101 ) | ( n2099 & n2102 ) | ( ~n2101 & n2102 ) ;
  assign n2104 = n2098 & n2103 ;
  assign n2105 = n2097 | n2103 ;
  assign n2106 = n2096 | n2105 ;
  assign n2107 = ~n2104 & n2106 ;
  assign n2108 = n1840 | n2107 ;
  assign n2109 = ( ~n1816 & n1819 ) | ( ~n1816 & n1835 ) | ( n1819 & n1835 ) ;
  assign n2110 = ( n1816 & ~n1835 ) | ( n1816 & n2109 ) | ( ~n1835 & n2109 ) ;
  assign n2111 = ( ~n1819 & n2109 ) | ( ~n1819 & n2110 ) | ( n2109 & n2110 ) ;
  assign n2112 = ( ~n2075 & n2078 ) | ( ~n2075 & n2094 ) | ( n2078 & n2094 ) ;
  assign n2113 = ( n2075 & ~n2094 ) | ( n2075 & n2112 ) | ( ~n2094 & n2112 ) ;
  assign n2114 = ( ~n2078 & n2112 ) | ( ~n2078 & n2113 ) | ( n2112 & n2113 ) ;
  assign n2115 = n2081 & ~n2084 ;
  assign n2116 = ~n2081 & n2084 ;
  assign n2117 = n2115 | n2116 ;
  assign n2118 = n1822 & ~n1825 ;
  assign n2119 = ~n1822 & n1825 ;
  assign n2120 = n2118 | n2119 ;
  assign n2121 = n2117 & n2120 ;
  assign n2122 = ( n2085 & ~n2090 ) | ( n2085 & n2093 ) | ( ~n2090 & n2093 ) ;
  assign n2123 = ( ~n2085 & n2090 ) | ( ~n2085 & n2122 ) | ( n2090 & n2122 ) ;
  assign n2124 = ( ~n2093 & n2122 ) | ( ~n2093 & n2123 ) | ( n2122 & n2123 ) ;
  assign n2125 = ( n1826 & ~n1831 ) | ( n1826 & n1834 ) | ( ~n1831 & n1834 ) ;
  assign n2126 = ( ~n1826 & n1831 ) | ( ~n1826 & n2125 ) | ( n1831 & n2125 ) ;
  assign n2127 = ( ~n1834 & n2125 ) | ( ~n1834 & n2126 ) | ( n2125 & n2126 ) ;
  assign n2128 = ( n2121 & n2124 ) | ( n2121 & n2127 ) | ( n2124 & n2127 ) ;
  assign n2129 = ( n2111 & n2114 ) | ( n2111 & n2128 ) | ( n2114 & n2128 ) ;
  assign n2130 = ( ~n1957 & n2071 ) | ( ~n1957 & n2095 ) | ( n2071 & n2095 ) ;
  assign n2131 = ( n1957 & ~n2095 ) | ( n1957 & n2130 ) | ( ~n2095 & n2130 ) ;
  assign n2132 = ( ~n2071 & n2130 ) | ( ~n2071 & n2131 ) | ( n2130 & n2131 ) ;
  assign n2133 = ( ~n1810 & n1813 ) | ( ~n1810 & n1836 ) | ( n1813 & n1836 ) ;
  assign n2134 = ( n1810 & ~n1836 ) | ( n1810 & n2133 ) | ( ~n1836 & n2133 ) ;
  assign n2135 = ( ~n1813 & n2133 ) | ( ~n1813 & n2134 ) | ( n2133 & n2134 ) ;
  assign n2136 = ( n2129 & n2132 ) | ( n2129 & n2135 ) | ( n2132 & n2135 ) ;
  assign n2137 = n2108 & n2136 ;
  assign n2138 = n1840 & n2107 ;
  assign n2139 = ( n1655 & n1800 ) | ( n1655 & n1803 ) | ( n1800 & n1803 ) ;
  assign n2140 = ( n1801 & n1837 ) | ( n1801 & n2139 ) | ( n1837 & n2139 ) ;
  assign n2141 = ( n2098 & n2100 ) | ( n2098 & n2104 ) | ( n2100 & n2104 ) ;
  assign n2142 = n2101 | n2141 ;
  assign n2143 = n2140 & n2142 ;
  assign n2144 = n2142 & ~n2143 ;
  assign n2145 = ( n2140 & ~n2143 ) | ( n2140 & n2144 ) | ( ~n2143 & n2144 ) ;
  assign n2146 = n2138 | n2145 ;
  assign n2147 = n2137 | n2146 ;
  assign n2148 = n2137 | n2138 ;
  assign n2149 = n2145 & n2148 ;
  assign n2150 = n2147 & ~n2149 ;
  assign n2151 = ( n1539 & ~n1543 ) | ( n1539 & n1571 ) | ( ~n1543 & n1571 ) ;
  assign n2152 = ( n1543 & ~n1571 ) | ( n1543 & n2151 ) | ( ~n1571 & n2151 ) ;
  assign n2153 = ( ~n1539 & n2151 ) | ( ~n1539 & n2152 ) | ( n2151 & n2152 ) ;
  assign n2154 = ( ~n1840 & n2107 ) | ( ~n1840 & n2136 ) | ( n2107 & n2136 ) ;
  assign n2155 = ( n1840 & ~n2136 ) | ( n1840 & n2154 ) | ( ~n2136 & n2154 ) ;
  assign n2156 = ( ~n2107 & n2154 ) | ( ~n2107 & n2155 ) | ( n2154 & n2155 ) ;
  assign n2157 = ( ~n1546 & n1549 ) | ( ~n1546 & n1563 ) | ( n1549 & n1563 ) ;
  assign n2158 = ( n1546 & ~n1563 ) | ( n1546 & n2157 ) | ( ~n1563 & n2157 ) ;
  assign n2159 = ( ~n1549 & n2157 ) | ( ~n1549 & n2158 ) | ( n2157 & n2158 ) ;
  assign n2160 = ( ~n2111 & n2114 ) | ( ~n2111 & n2128 ) | ( n2114 & n2128 ) ;
  assign n2161 = ( n2111 & ~n2128 ) | ( n2111 & n2160 ) | ( ~n2128 & n2160 ) ;
  assign n2162 = ( ~n2114 & n2160 ) | ( ~n2114 & n2161 ) | ( n2160 & n2161 ) ;
  assign n2163 = n2117 & ~n2120 ;
  assign n2164 = ~n2117 & n2120 ;
  assign n2165 = n2163 | n2164 ;
  assign n2166 = n1552 & ~n1555 ;
  assign n2167 = ~n1552 & n1555 ;
  assign n2168 = n2166 | n2167 ;
  assign n2169 = n2165 & n2168 ;
  assign n2170 = ~n2121 & n2124 ;
  assign n2171 = n2121 & ~n2124 ;
  assign n2172 = n2170 | n2171 ;
  assign n2173 = n2127 & ~n2172 ;
  assign n2174 = ~n2127 & n2172 ;
  assign n2175 = n2173 | n2174 ;
  assign n2176 = ( n1556 & n1562 ) | ( n1556 & ~n1563 ) | ( n1562 & ~n1563 ) ;
  assign n2177 = ( n1559 & ~n1563 ) | ( n1559 & n2176 ) | ( ~n1563 & n2176 ) ;
  assign n2178 = ( n2169 & n2175 ) | ( n2169 & n2177 ) | ( n2175 & n2177 ) ;
  assign n2179 = ( n2159 & n2162 ) | ( n2159 & n2178 ) | ( n2162 & n2178 ) ;
  assign n2180 = ( n2129 & ~n2132 ) | ( n2129 & n2135 ) | ( ~n2132 & n2135 ) ;
  assign n2181 = ( ~n2129 & n2132 ) | ( ~n2129 & n2180 ) | ( n2132 & n2180 ) ;
  assign n2182 = ( ~n2135 & n2180 ) | ( ~n2135 & n2181 ) | ( n2180 & n2181 ) ;
  assign n2183 = ( n1564 & ~n1567 ) | ( n1564 & n1570 ) | ( ~n1567 & n1570 ) ;
  assign n2184 = ( ~n1564 & n1567 ) | ( ~n1564 & n2183 ) | ( n1567 & n2183 ) ;
  assign n2185 = ( ~n1570 & n2183 ) | ( ~n1570 & n2184 ) | ( n2183 & n2184 ) ;
  assign n2186 = ( n2179 & n2182 ) | ( n2179 & n2185 ) | ( n2182 & n2185 ) ;
  assign n2187 = ( n2153 & n2156 ) | ( n2153 & n2186 ) | ( n2156 & n2186 ) ;
  assign n2188 = ( n1575 & ~n2150 ) | ( n1575 & n2187 ) | ( ~n2150 & n2187 ) ;
  assign n2189 = ( n2150 & ~n2187 ) | ( n2150 & n2188 ) | ( ~n2187 & n2188 ) ;
  assign n2190 = ( ~n1575 & n2188 ) | ( ~n1575 & n2189 ) | ( n2188 & n2189 ) ;
  assign n2191 = ( x106 & x107 ) | ( x106 & x108 ) | ( x107 & x108 ) ;
  assign n2192 = ( x103 & x104 ) | ( x103 & x105 ) | ( x104 & x105 ) ;
  assign n2193 = ( x103 & ~x104 ) | ( x103 & x105 ) | ( ~x104 & x105 ) ;
  assign n2194 = ( ~x103 & x104 ) | ( ~x103 & n2193 ) | ( x104 & n2193 ) ;
  assign n2195 = ( ~x105 & n2193 ) | ( ~x105 & n2194 ) | ( n2193 & n2194 ) ;
  assign n2196 = ( x106 & ~x107 ) | ( x106 & x108 ) | ( ~x107 & x108 ) ;
  assign n2197 = ( ~x106 & x107 ) | ( ~x106 & n2196 ) | ( x107 & n2196 ) ;
  assign n2198 = ( ~x108 & n2196 ) | ( ~x108 & n2197 ) | ( n2196 & n2197 ) ;
  assign n2199 = n2195 & n2198 ;
  assign n2200 = ( n2191 & n2192 ) | ( n2191 & n2199 ) | ( n2192 & n2199 ) ;
  assign n2201 = ( n2192 & n2199 ) | ( n2192 & ~n2200 ) | ( n2199 & ~n2200 ) ;
  assign n2202 = ( n2191 & ~n2200 ) | ( n2191 & n2201 ) | ( ~n2200 & n2201 ) ;
  assign n2203 = ( x112 & x113 ) | ( x112 & x114 ) | ( x113 & x114 ) ;
  assign n2204 = ( x109 & x110 ) | ( x109 & x111 ) | ( x110 & x111 ) ;
  assign n2205 = ( x109 & ~x110 ) | ( x109 & x111 ) | ( ~x110 & x111 ) ;
  assign n2206 = ( ~x109 & x110 ) | ( ~x109 & n2205 ) | ( x110 & n2205 ) ;
  assign n2207 = ( ~x111 & n2205 ) | ( ~x111 & n2206 ) | ( n2205 & n2206 ) ;
  assign n2208 = ( x112 & ~x113 ) | ( x112 & x114 ) | ( ~x113 & x114 ) ;
  assign n2209 = ( ~x112 & x113 ) | ( ~x112 & n2208 ) | ( x113 & n2208 ) ;
  assign n2210 = ( ~x114 & n2208 ) | ( ~x114 & n2209 ) | ( n2208 & n2209 ) ;
  assign n2211 = n2207 & n2210 ;
  assign n2212 = ( n2203 & n2204 ) | ( n2203 & n2211 ) | ( n2204 & n2211 ) ;
  assign n2213 = ( n2204 & n2211 ) | ( n2204 & ~n2212 ) | ( n2211 & ~n2212 ) ;
  assign n2214 = ( n2203 & ~n2212 ) | ( n2203 & n2213 ) | ( ~n2212 & n2213 ) ;
  assign n2215 = n2200 & n2202 ;
  assign n2216 = n2212 & n2214 ;
  assign n2217 = n2195 & ~n2198 ;
  assign n2218 = ~n2195 & n2198 ;
  assign n2219 = n2217 | n2218 ;
  assign n2220 = n2207 & ~n2210 ;
  assign n2221 = ~n2207 & n2210 ;
  assign n2222 = n2220 | n2221 ;
  assign n2223 = n2219 & n2222 ;
  assign n2224 = ~n2216 & n2223 ;
  assign n2225 = ~n2215 & n2224 ;
  assign n2226 = ~n2214 & n2225 ;
  assign n2227 = ( n2202 & n2214 ) | ( n2202 & n2226 ) | ( n2214 & n2226 ) ;
  assign n2228 = n2214 & n2224 ;
  assign n2229 = ~n2215 & n2228 ;
  assign n2230 = ~n2200 & n2212 ;
  assign n2231 = n2200 & ~n2212 ;
  assign n2232 = n2230 | n2231 ;
  assign n2233 = n2229 | n2232 ;
  assign n2234 = n2227 | n2233 ;
  assign n2235 = n2227 | n2229 ;
  assign n2236 = n2232 & n2235 ;
  assign n2237 = n2234 & ~n2236 ;
  assign n2238 = ( x118 & x119 ) | ( x118 & x120 ) | ( x119 & x120 ) ;
  assign n2239 = ( x115 & x116 ) | ( x115 & x117 ) | ( x116 & x117 ) ;
  assign n2240 = ( x115 & ~x116 ) | ( x115 & x117 ) | ( ~x116 & x117 ) ;
  assign n2241 = ( ~x115 & x116 ) | ( ~x115 & n2240 ) | ( x116 & n2240 ) ;
  assign n2242 = ( ~x117 & n2240 ) | ( ~x117 & n2241 ) | ( n2240 & n2241 ) ;
  assign n2243 = ( x118 & ~x119 ) | ( x118 & x120 ) | ( ~x119 & x120 ) ;
  assign n2244 = ( ~x118 & x119 ) | ( ~x118 & n2243 ) | ( x119 & n2243 ) ;
  assign n2245 = ( ~x120 & n2243 ) | ( ~x120 & n2244 ) | ( n2243 & n2244 ) ;
  assign n2246 = n2242 & n2245 ;
  assign n2247 = ( n2238 & n2239 ) | ( n2238 & n2246 ) | ( n2239 & n2246 ) ;
  assign n2248 = ( n2239 & n2246 ) | ( n2239 & ~n2247 ) | ( n2246 & ~n2247 ) ;
  assign n2249 = ( n2238 & ~n2247 ) | ( n2238 & n2248 ) | ( ~n2247 & n2248 ) ;
  assign n2250 = ( x124 & x125 ) | ( x124 & x126 ) | ( x125 & x126 ) ;
  assign n2251 = ( x121 & x122 ) | ( x121 & x123 ) | ( x122 & x123 ) ;
  assign n2252 = ( x121 & ~x122 ) | ( x121 & x123 ) | ( ~x122 & x123 ) ;
  assign n2253 = ( ~x121 & x122 ) | ( ~x121 & n2252 ) | ( x122 & n2252 ) ;
  assign n2254 = ( ~x123 & n2252 ) | ( ~x123 & n2253 ) | ( n2252 & n2253 ) ;
  assign n2255 = ( x124 & ~x125 ) | ( x124 & x126 ) | ( ~x125 & x126 ) ;
  assign n2256 = ( ~x124 & x125 ) | ( ~x124 & n2255 ) | ( x125 & n2255 ) ;
  assign n2257 = ( ~x126 & n2255 ) | ( ~x126 & n2256 ) | ( n2255 & n2256 ) ;
  assign n2258 = n2254 & n2257 ;
  assign n2259 = ( n2250 & n2251 ) | ( n2250 & n2258 ) | ( n2251 & n2258 ) ;
  assign n2260 = ( n2251 & n2258 ) | ( n2251 & ~n2259 ) | ( n2258 & ~n2259 ) ;
  assign n2261 = ( n2250 & ~n2259 ) | ( n2250 & n2260 ) | ( ~n2259 & n2260 ) ;
  assign n2262 = n2247 & n2249 ;
  assign n2263 = n2242 & ~n2245 ;
  assign n2264 = ~n2242 & n2245 ;
  assign n2265 = n2263 | n2264 ;
  assign n2266 = n2254 & ~n2257 ;
  assign n2267 = ~n2254 & n2257 ;
  assign n2268 = n2266 | n2267 ;
  assign n2269 = n2265 & n2268 ;
  assign n2270 = ~n2262 & n2269 ;
  assign n2271 = ( n2249 & n2261 ) | ( n2249 & n2270 ) | ( n2261 & n2270 ) ;
  assign n2272 = ~n2247 & n2259 ;
  assign n2273 = n2247 & ~n2259 ;
  assign n2274 = n2272 | n2273 ;
  assign n2275 = n2271 & n2274 ;
  assign n2276 = n2271 | n2274 ;
  assign n2277 = ~n2275 & n2276 ;
  assign n2278 = n2237 | n2277 ;
  assign n2279 = ( n2202 & n2214 ) | ( n2202 & ~n2225 ) | ( n2214 & ~n2225 ) ;
  assign n2280 = n2202 & ~n2229 ;
  assign n2281 = ( n2214 & ~n2279 ) | ( n2214 & n2280 ) | ( ~n2279 & n2280 ) ;
  assign n2282 = ( n2226 & n2279 ) | ( n2226 & ~n2281 ) | ( n2279 & ~n2281 ) ;
  assign n2283 = n2265 & ~n2268 ;
  assign n2284 = ~n2265 & n2268 ;
  assign n2285 = n2283 | n2284 ;
  assign n2286 = n2219 & ~n2222 ;
  assign n2287 = ~n2219 & n2222 ;
  assign n2288 = n2286 | n2287 ;
  assign n2289 = n2285 & n2288 ;
  assign n2290 = n2261 | n2270 ;
  assign n2291 = ~n2271 & n2290 ;
  assign n2292 = n2261 & n2269 ;
  assign n2293 = ( n2249 & ~n2290 ) | ( n2249 & n2292 ) | ( ~n2290 & n2292 ) ;
  assign n2294 = n2291 | n2293 ;
  assign n2295 = n2289 | n2294 ;
  assign n2296 = ( n2289 & n2291 ) | ( n2289 & n2293 ) | ( n2291 & n2293 ) ;
  assign n2297 = ( n2282 & n2295 ) | ( n2282 & n2296 ) | ( n2295 & n2296 ) ;
  assign n2298 = n2278 & n2297 ;
  assign n2299 = n2237 & n2277 ;
  assign n2300 = ( n2247 & n2259 ) | ( n2247 & n2271 ) | ( n2259 & n2271 ) ;
  assign n2301 = ( n2200 & n2212 ) | ( n2200 & n2235 ) | ( n2212 & n2235 ) ;
  assign n2302 = ~n2300 & n2301 ;
  assign n2303 = n2300 & ~n2301 ;
  assign n2304 = n2302 | n2303 ;
  assign n2305 = n2299 | n2304 ;
  assign n2306 = n2298 | n2305 ;
  assign n2307 = n2298 | n2299 ;
  assign n2308 = n2304 & n2307 ;
  assign n2309 = n2306 & ~n2308 ;
  assign n2345 = ( x88 & x89 ) | ( x88 & x90 ) | ( x89 & x90 ) ;
  assign n2346 = ( x85 & x86 ) | ( x85 & x87 ) | ( x86 & x87 ) ;
  assign n2347 = ( x85 & ~x86 ) | ( x85 & x87 ) | ( ~x86 & x87 ) ;
  assign n2348 = ( ~x85 & x86 ) | ( ~x85 & n2347 ) | ( x86 & n2347 ) ;
  assign n2349 = ( ~x87 & n2347 ) | ( ~x87 & n2348 ) | ( n2347 & n2348 ) ;
  assign n2350 = ( x88 & ~x89 ) | ( x88 & x90 ) | ( ~x89 & x90 ) ;
  assign n2351 = ( ~x88 & x89 ) | ( ~x88 & n2350 ) | ( x89 & n2350 ) ;
  assign n2352 = ( ~x90 & n2350 ) | ( ~x90 & n2351 ) | ( n2350 & n2351 ) ;
  assign n2353 = n2349 & n2352 ;
  assign n2354 = ( n2345 & n2346 ) | ( n2345 & n2353 ) | ( n2346 & n2353 ) ;
  assign n2368 = ( n2346 & n2353 ) | ( n2346 & ~n2354 ) | ( n2353 & ~n2354 ) ;
  assign n2369 = ( n2345 & ~n2354 ) | ( n2345 & n2368 ) | ( ~n2354 & n2368 ) ;
  assign n2355 = ( x82 & x83 ) | ( x82 & x84 ) | ( x83 & x84 ) ;
  assign n2356 = ( x79 & x80 ) | ( x79 & x81 ) | ( x80 & x81 ) ;
  assign n2357 = ( x79 & ~x80 ) | ( x79 & x81 ) | ( ~x80 & x81 ) ;
  assign n2358 = ( ~x79 & x80 ) | ( ~x79 & n2357 ) | ( x80 & n2357 ) ;
  assign n2359 = ( ~x81 & n2357 ) | ( ~x81 & n2358 ) | ( n2357 & n2358 ) ;
  assign n2360 = ( x82 & ~x83 ) | ( x82 & x84 ) | ( ~x83 & x84 ) ;
  assign n2361 = ( ~x82 & x83 ) | ( ~x82 & n2360 ) | ( x83 & n2360 ) ;
  assign n2362 = ( ~x84 & n2360 ) | ( ~x84 & n2361 ) | ( n2360 & n2361 ) ;
  assign n2363 = n2359 & n2362 ;
  assign n2364 = ( n2355 & n2356 ) | ( n2355 & n2363 ) | ( n2356 & n2363 ) ;
  assign n2365 = ( n2356 & n2363 ) | ( n2356 & ~n2364 ) | ( n2363 & ~n2364 ) ;
  assign n2366 = ( n2355 & ~n2364 ) | ( n2355 & n2365 ) | ( ~n2364 & n2365 ) ;
  assign n2367 = n2364 & n2366 ;
  assign n2370 = n2354 & n2369 ;
  assign n2371 = n2349 & ~n2352 ;
  assign n2372 = ~n2349 & n2352 ;
  assign n2373 = n2371 | n2372 ;
  assign n2374 = n2359 & ~n2362 ;
  assign n2375 = ~n2359 & n2362 ;
  assign n2376 = n2374 | n2375 ;
  assign n2377 = n2373 & n2376 ;
  assign n2378 = ~n2370 & n2377 ;
  assign n2381 = ~n2367 & n2378 ;
  assign n2382 = ~n2369 & n2381 ;
  assign n2389 = ( n2366 & n2369 ) | ( n2366 & ~n2381 ) | ( n2369 & ~n2381 ) ;
  assign n2379 = n2369 & n2378 ;
  assign n2380 = ~n2367 & n2379 ;
  assign n2390 = n2366 & ~n2380 ;
  assign n2391 = ( n2369 & ~n2389 ) | ( n2369 & n2390 ) | ( ~n2389 & n2390 ) ;
  assign n2392 = ( n2382 & n2389 ) | ( n2382 & ~n2391 ) | ( n2389 & ~n2391 ) ;
  assign n2312 = ( x91 & ~x92 ) | ( x91 & x93 ) | ( ~x92 & x93 ) ;
  assign n2313 = ( ~x91 & x92 ) | ( ~x91 & n2312 ) | ( x92 & n2312 ) ;
  assign n2314 = ( ~x93 & n2312 ) | ( ~x93 & n2313 ) | ( n2312 & n2313 ) ;
  assign n2315 = ( x94 & ~x95 ) | ( x94 & x96 ) | ( ~x95 & x96 ) ;
  assign n2316 = ( ~x94 & x95 ) | ( ~x94 & n2315 ) | ( x95 & n2315 ) ;
  assign n2317 = ( ~x96 & n2315 ) | ( ~x96 & n2316 ) | ( n2315 & n2316 ) ;
  assign n2335 = n2314 & ~n2317 ;
  assign n2336 = ~n2314 & n2317 ;
  assign n2337 = n2335 | n2336 ;
  assign n2322 = ( x97 & ~x98 ) | ( x97 & x99 ) | ( ~x98 & x99 ) ;
  assign n2323 = ( ~x97 & x98 ) | ( ~x97 & n2322 ) | ( x98 & n2322 ) ;
  assign n2324 = ( ~x99 & n2322 ) | ( ~x99 & n2323 ) | ( n2322 & n2323 ) ;
  assign n2325 = ( x100 & ~x101 ) | ( x100 & x102 ) | ( ~x101 & x102 ) ;
  assign n2326 = ( ~x100 & x101 ) | ( ~x100 & n2325 ) | ( x101 & n2325 ) ;
  assign n2327 = ( ~x102 & n2325 ) | ( ~x102 & n2326 ) | ( n2325 & n2326 ) ;
  assign n2338 = n2324 & ~n2327 ;
  assign n2339 = ~n2324 & n2327 ;
  assign n2340 = n2338 | n2339 ;
  assign n2393 = n2337 & ~n2340 ;
  assign n2394 = ~n2337 & n2340 ;
  assign n2395 = n2393 | n2394 ;
  assign n2396 = ~n2373 & n2376 ;
  assign n2397 = n2373 & ~n2376 ;
  assign n2398 = n2396 | n2397 ;
  assign n2399 = n2395 & n2398 ;
  assign n2310 = ( x94 & x95 ) | ( x94 & x96 ) | ( x95 & x96 ) ;
  assign n2311 = ( x91 & x92 ) | ( x91 & x93 ) | ( x92 & x93 ) ;
  assign n2318 = n2314 & n2317 ;
  assign n2319 = ( n2310 & n2311 ) | ( n2310 & n2318 ) | ( n2311 & n2318 ) ;
  assign n2330 = ( n2311 & n2318 ) | ( n2311 & ~n2319 ) | ( n2318 & ~n2319 ) ;
  assign n2331 = ( n2310 & ~n2319 ) | ( n2310 & n2330 ) | ( ~n2319 & n2330 ) ;
  assign n2320 = ( x100 & x101 ) | ( x100 & x102 ) | ( x101 & x102 ) ;
  assign n2321 = ( x97 & x98 ) | ( x97 & x99 ) | ( x98 & x99 ) ;
  assign n2328 = n2324 & n2327 ;
  assign n2329 = ( n2320 & n2321 ) | ( n2320 & n2328 ) | ( n2321 & n2328 ) ;
  assign n2332 = ( n2321 & n2328 ) | ( n2321 & ~n2329 ) | ( n2328 & ~n2329 ) ;
  assign n2333 = ( n2320 & ~n2329 ) | ( n2320 & n2332 ) | ( ~n2329 & n2332 ) ;
  assign n2341 = n2337 & n2340 ;
  assign n2400 = n2333 & n2341 ;
  assign n2334 = n2319 & n2331 ;
  assign n2342 = ~n2334 & n2341 ;
  assign n2401 = n2333 | n2342 ;
  assign n2402 = ( n2331 & n2400 ) | ( n2331 & ~n2401 ) | ( n2400 & ~n2401 ) ;
  assign n2343 = ( n2331 & n2333 ) | ( n2331 & n2342 ) | ( n2333 & n2342 ) ;
  assign n2403 = ~n2343 & n2401 ;
  assign n2404 = n2402 | n2403 ;
  assign n2405 = n2399 | n2404 ;
  assign n2406 = n2392 & n2405 ;
  assign n2407 = ( n2399 & n2402 ) | ( n2399 & n2403 ) | ( n2402 & n2403 ) ;
  assign n2408 = n2406 | n2407 ;
  assign n2383 = ( n2366 & n2369 ) | ( n2366 & n2382 ) | ( n2369 & n2382 ) ;
  assign n2409 = n2354 & ~n2364 ;
  assign n2410 = ~n2354 & n2364 ;
  assign n2411 = n2409 | n2410 ;
  assign n2412 = n2380 | n2411 ;
  assign n2413 = n2383 | n2412 ;
  assign n2384 = n2380 | n2383 ;
  assign n2414 = n2384 & n2411 ;
  assign n2415 = n2413 & ~n2414 ;
  assign n2416 = ~n2319 & n2329 ;
  assign n2417 = n2319 & ~n2329 ;
  assign n2418 = n2416 | n2417 ;
  assign n2419 = n2343 & n2418 ;
  assign n2420 = n2343 | n2418 ;
  assign n2421 = ~n2419 & n2420 ;
  assign n2422 = ( n2408 & n2415 ) | ( n2408 & n2421 ) | ( n2415 & n2421 ) ;
  assign n2344 = ( n2319 & n2329 ) | ( n2319 & n2343 ) | ( n2329 & n2343 ) ;
  assign n2385 = ( n2354 & n2364 ) | ( n2354 & n2384 ) | ( n2364 & n2384 ) ;
  assign n2386 = n2344 & n2385 ;
  assign n2387 = n2385 & ~n2386 ;
  assign n2388 = ( n2344 & ~n2386 ) | ( n2344 & n2387 ) | ( ~n2386 & n2387 ) ;
  assign n2423 = n2388 | n2422 ;
  assign n2424 = ~n2388 & n2423 ;
  assign n2425 = ( ~n2422 & n2423 ) | ( ~n2422 & n2424 ) | ( n2423 & n2424 ) ;
  assign n2426 = n2309 | n2425 ;
  assign n2427 = ( n2408 & ~n2415 ) | ( n2408 & n2421 ) | ( ~n2415 & n2421 ) ;
  assign n2428 = ( ~n2408 & n2415 ) | ( ~n2408 & n2427 ) | ( n2415 & n2427 ) ;
  assign n2429 = ( ~n2421 & n2427 ) | ( ~n2421 & n2428 ) | ( n2427 & n2428 ) ;
  assign n2430 = ( ~n2237 & n2277 ) | ( ~n2237 & n2297 ) | ( n2277 & n2297 ) ;
  assign n2431 = ( n2237 & ~n2297 ) | ( n2237 & n2430 ) | ( ~n2297 & n2430 ) ;
  assign n2432 = ( ~n2277 & n2430 ) | ( ~n2277 & n2431 ) | ( n2430 & n2431 ) ;
  assign n2433 = n2285 & ~n2288 ;
  assign n2434 = ~n2285 & n2288 ;
  assign n2435 = n2433 | n2434 ;
  assign n2436 = n2395 & ~n2398 ;
  assign n2437 = ~n2395 & n2398 ;
  assign n2438 = n2436 | n2437 ;
  assign n2439 = n2435 & n2438 ;
  assign n2440 = ~n2289 & n2295 ;
  assign n2441 = ( ~n2294 & n2295 ) | ( ~n2294 & n2440 ) | ( n2295 & n2440 ) ;
  assign n2442 = n2282 & ~n2441 ;
  assign n2443 = ~n2282 & n2441 ;
  assign n2444 = n2442 | n2443 ;
  assign n2445 = ( n2392 & n2399 ) | ( n2392 & ~n2404 ) | ( n2399 & ~n2404 ) ;
  assign n2446 = ( ~n2392 & n2404 ) | ( ~n2392 & n2445 ) | ( n2404 & n2445 ) ;
  assign n2447 = ( ~n2399 & n2445 ) | ( ~n2399 & n2446 ) | ( n2445 & n2446 ) ;
  assign n2448 = ( n2439 & n2444 ) | ( n2439 & n2447 ) | ( n2444 & n2447 ) ;
  assign n2449 = ( n2429 & n2432 ) | ( n2429 & n2448 ) | ( n2432 & n2448 ) ;
  assign n2450 = n2426 & n2449 ;
  assign n2451 = n2309 & n2425 ;
  assign n2452 = n2450 | n2451 ;
  assign n2453 = n2386 | n2388 ;
  assign n2454 = ( n2386 & n2422 ) | ( n2386 & n2453 ) | ( n2422 & n2453 ) ;
  assign n2455 = ( n2300 & n2301 ) | ( n2300 & n2307 ) | ( n2301 & n2307 ) ;
  assign n2456 = n2454 & n2455 ;
  assign n2457 = n2455 & ~n2456 ;
  assign n2458 = ( n2454 & ~n2456 ) | ( n2454 & n2457 ) | ( ~n2456 & n2457 ) ;
  assign n2459 = ( n2453 & n2455 ) | ( n2453 & n2458 ) | ( n2455 & n2458 ) ;
  assign n2460 = ( n2452 & n2456 ) | ( n2452 & n2459 ) | ( n2456 & n2459 ) ;
  assign n2461 = ( x142 & x143 ) | ( x142 & x144 ) | ( x143 & x144 ) ;
  assign n2462 = ( x139 & x140 ) | ( x139 & x141 ) | ( x140 & x141 ) ;
  assign n2463 = ( x139 & ~x140 ) | ( x139 & x141 ) | ( ~x140 & x141 ) ;
  assign n2464 = ( ~x139 & x140 ) | ( ~x139 & n2463 ) | ( x140 & n2463 ) ;
  assign n2465 = ( ~x141 & n2463 ) | ( ~x141 & n2464 ) | ( n2463 & n2464 ) ;
  assign n2466 = ( x142 & ~x143 ) | ( x142 & x144 ) | ( ~x143 & x144 ) ;
  assign n2467 = ( ~x142 & x143 ) | ( ~x142 & n2466 ) | ( x143 & n2466 ) ;
  assign n2468 = ( ~x144 & n2466 ) | ( ~x144 & n2467 ) | ( n2466 & n2467 ) ;
  assign n2469 = n2465 & n2468 ;
  assign n2470 = ( n2461 & n2462 ) | ( n2461 & n2469 ) | ( n2462 & n2469 ) ;
  assign n2471 = ( x148 & x149 ) | ( x148 & x150 ) | ( x149 & x150 ) ;
  assign n2472 = ( x145 & x146 ) | ( x145 & x147 ) | ( x146 & x147 ) ;
  assign n2473 = ( x145 & ~x146 ) | ( x145 & x147 ) | ( ~x146 & x147 ) ;
  assign n2474 = ( ~x145 & x146 ) | ( ~x145 & n2473 ) | ( x146 & n2473 ) ;
  assign n2475 = ( ~x147 & n2473 ) | ( ~x147 & n2474 ) | ( n2473 & n2474 ) ;
  assign n2476 = ( x148 & ~x149 ) | ( x148 & x150 ) | ( ~x149 & x150 ) ;
  assign n2477 = ( ~x148 & x149 ) | ( ~x148 & n2476 ) | ( x149 & n2476 ) ;
  assign n2478 = ( ~x150 & n2476 ) | ( ~x150 & n2477 ) | ( n2476 & n2477 ) ;
  assign n2479 = n2475 & n2478 ;
  assign n2480 = ( n2471 & n2472 ) | ( n2471 & n2479 ) | ( n2472 & n2479 ) ;
  assign n2481 = ( n2462 & n2469 ) | ( n2462 & ~n2470 ) | ( n2469 & ~n2470 ) ;
  assign n2482 = ( n2461 & ~n2470 ) | ( n2461 & n2481 ) | ( ~n2470 & n2481 ) ;
  assign n2483 = ( n2472 & n2479 ) | ( n2472 & ~n2480 ) | ( n2479 & ~n2480 ) ;
  assign n2484 = ( n2471 & ~n2480 ) | ( n2471 & n2483 ) | ( ~n2480 & n2483 ) ;
  assign n2485 = n2470 & n2482 ;
  assign n2486 = n2465 & ~n2468 ;
  assign n2487 = ~n2465 & n2468 ;
  assign n2488 = n2486 | n2487 ;
  assign n2489 = n2475 & ~n2478 ;
  assign n2490 = ~n2475 & n2478 ;
  assign n2491 = n2489 | n2490 ;
  assign n2492 = n2488 & n2491 ;
  assign n2493 = ~n2485 & n2492 ;
  assign n2494 = ( n2482 & n2484 ) | ( n2482 & n2493 ) | ( n2484 & n2493 ) ;
  assign n2495 = ( n2470 & n2480 ) | ( n2470 & n2494 ) | ( n2480 & n2494 ) ;
  assign n2496 = ( x136 & x137 ) | ( x136 & x138 ) | ( x137 & x138 ) ;
  assign n2497 = ( x133 & x134 ) | ( x133 & x135 ) | ( x134 & x135 ) ;
  assign n2498 = ( x133 & ~x134 ) | ( x133 & x135 ) | ( ~x134 & x135 ) ;
  assign n2499 = ( ~x133 & x134 ) | ( ~x133 & n2498 ) | ( x134 & n2498 ) ;
  assign n2500 = ( ~x135 & n2498 ) | ( ~x135 & n2499 ) | ( n2498 & n2499 ) ;
  assign n2501 = ( x136 & ~x137 ) | ( x136 & x138 ) | ( ~x137 & x138 ) ;
  assign n2502 = ( ~x136 & x137 ) | ( ~x136 & n2501 ) | ( x137 & n2501 ) ;
  assign n2503 = ( ~x138 & n2501 ) | ( ~x138 & n2502 ) | ( n2501 & n2502 ) ;
  assign n2504 = n2500 & n2503 ;
  assign n2505 = ( n2496 & n2497 ) | ( n2496 & n2504 ) | ( n2497 & n2504 ) ;
  assign n2506 = ( x130 & x131 ) | ( x130 & x132 ) | ( x131 & x132 ) ;
  assign n2507 = ( x127 & x128 ) | ( x127 & x129 ) | ( x128 & x129 ) ;
  assign n2508 = ( x127 & ~x128 ) | ( x127 & x129 ) | ( ~x128 & x129 ) ;
  assign n2509 = ( ~x127 & x128 ) | ( ~x127 & n2508 ) | ( x128 & n2508 ) ;
  assign n2510 = ( ~x129 & n2508 ) | ( ~x129 & n2509 ) | ( n2508 & n2509 ) ;
  assign n2511 = ( x130 & ~x131 ) | ( x130 & x132 ) | ( ~x131 & x132 ) ;
  assign n2512 = ( ~x130 & x131 ) | ( ~x130 & n2511 ) | ( x131 & n2511 ) ;
  assign n2513 = ( ~x132 & n2511 ) | ( ~x132 & n2512 ) | ( n2511 & n2512 ) ;
  assign n2514 = n2510 & n2513 ;
  assign n2515 = ( n2506 & n2507 ) | ( n2506 & n2514 ) | ( n2507 & n2514 ) ;
  assign n2516 = ( n2507 & n2514 ) | ( n2507 & ~n2515 ) | ( n2514 & ~n2515 ) ;
  assign n2517 = ( n2506 & ~n2515 ) | ( n2506 & n2516 ) | ( ~n2515 & n2516 ) ;
  assign n2518 = n2515 & n2517 ;
  assign n2519 = ( n2497 & n2504 ) | ( n2497 & ~n2505 ) | ( n2504 & ~n2505 ) ;
  assign n2520 = ( n2496 & ~n2505 ) | ( n2496 & n2519 ) | ( ~n2505 & n2519 ) ;
  assign n2521 = n2505 & n2520 ;
  assign n2522 = n2500 & ~n2503 ;
  assign n2523 = ~n2500 & n2503 ;
  assign n2524 = n2522 | n2523 ;
  assign n2525 = n2510 & ~n2513 ;
  assign n2526 = ~n2510 & n2513 ;
  assign n2527 = n2525 | n2526 ;
  assign n2528 = n2524 & n2527 ;
  assign n2529 = ~n2521 & n2528 ;
  assign n2530 = n2520 & n2529 ;
  assign n2531 = ~n2518 & n2530 ;
  assign n2532 = ~n2518 & n2529 ;
  assign n2533 = ~n2520 & n2532 ;
  assign n2534 = ( n2517 & n2520 ) | ( n2517 & n2533 ) | ( n2520 & n2533 ) ;
  assign n2535 = n2531 | n2534 ;
  assign n2536 = ( n2505 & n2515 ) | ( n2505 & n2535 ) | ( n2515 & n2535 ) ;
  assign n2537 = ( n2517 & n2520 ) | ( n2517 & ~n2532 ) | ( n2520 & ~n2532 ) ;
  assign n2538 = n2517 & ~n2531 ;
  assign n2539 = ( n2520 & ~n2537 ) | ( n2520 & n2538 ) | ( ~n2537 & n2538 ) ;
  assign n2540 = ( n2533 & n2537 ) | ( n2533 & ~n2539 ) | ( n2537 & ~n2539 ) ;
  assign n2541 = n2488 & ~n2491 ;
  assign n2542 = ~n2488 & n2491 ;
  assign n2543 = n2541 | n2542 ;
  assign n2544 = ~n2524 & n2527 ;
  assign n2545 = n2524 & ~n2527 ;
  assign n2546 = n2544 | n2545 ;
  assign n2547 = n2543 & n2546 ;
  assign n2548 = n2484 & n2492 ;
  assign n2549 = n2484 | n2493 ;
  assign n2550 = ( n2482 & n2548 ) | ( n2482 & ~n2549 ) | ( n2548 & ~n2549 ) ;
  assign n2551 = ~n2494 & n2549 ;
  assign n2552 = n2550 | n2551 ;
  assign n2553 = n2547 | n2552 ;
  assign n2554 = n2540 & n2553 ;
  assign n2555 = ( n2547 & n2550 ) | ( n2547 & n2551 ) | ( n2550 & n2551 ) ;
  assign n2556 = n2554 | n2555 ;
  assign n2557 = n2505 & ~n2515 ;
  assign n2558 = ~n2505 & n2515 ;
  assign n2559 = n2557 | n2558 ;
  assign n2560 = n2531 | n2559 ;
  assign n2561 = n2534 | n2560 ;
  assign n2562 = n2535 & n2559 ;
  assign n2563 = n2561 & ~n2562 ;
  assign n2564 = ~n2470 & n2480 ;
  assign n2565 = n2470 & ~n2480 ;
  assign n2566 = n2564 | n2565 ;
  assign n2567 = n2494 & n2566 ;
  assign n2568 = n2494 | n2566 ;
  assign n2569 = ~n2567 & n2568 ;
  assign n2570 = ( n2556 & n2563 ) | ( n2556 & n2569 ) | ( n2563 & n2569 ) ;
  assign n2571 = ( n2495 & n2536 ) | ( n2495 & n2570 ) | ( n2536 & n2570 ) ;
  assign n2572 = ( x166 & x167 ) | ( x166 & x168 ) | ( x167 & x168 ) ;
  assign n2573 = ( x163 & x164 ) | ( x163 & x165 ) | ( x164 & x165 ) ;
  assign n2574 = ( x163 & ~x164 ) | ( x163 & x165 ) | ( ~x164 & x165 ) ;
  assign n2575 = ( ~x163 & x164 ) | ( ~x163 & n2574 ) | ( x164 & n2574 ) ;
  assign n2576 = ( ~x165 & n2574 ) | ( ~x165 & n2575 ) | ( n2574 & n2575 ) ;
  assign n2577 = ( x166 & ~x167 ) | ( x166 & x168 ) | ( ~x167 & x168 ) ;
  assign n2578 = ( ~x166 & x167 ) | ( ~x166 & n2577 ) | ( x167 & n2577 ) ;
  assign n2579 = ( ~x168 & n2577 ) | ( ~x168 & n2578 ) | ( n2577 & n2578 ) ;
  assign n2580 = n2576 & n2579 ;
  assign n2581 = ( n2572 & n2573 ) | ( n2572 & n2580 ) | ( n2573 & n2580 ) ;
  assign n2582 = ( x172 & x173 ) | ( x172 & x174 ) | ( x173 & x174 ) ;
  assign n2583 = ( x169 & x170 ) | ( x169 & x171 ) | ( x170 & x171 ) ;
  assign n2584 = ( x169 & ~x170 ) | ( x169 & x171 ) | ( ~x170 & x171 ) ;
  assign n2585 = ( ~x169 & x170 ) | ( ~x169 & n2584 ) | ( x170 & n2584 ) ;
  assign n2586 = ( ~x171 & n2584 ) | ( ~x171 & n2585 ) | ( n2584 & n2585 ) ;
  assign n2587 = ( x172 & ~x173 ) | ( x172 & x174 ) | ( ~x173 & x174 ) ;
  assign n2588 = ( ~x172 & x173 ) | ( ~x172 & n2587 ) | ( x173 & n2587 ) ;
  assign n2589 = ( ~x174 & n2587 ) | ( ~x174 & n2588 ) | ( n2587 & n2588 ) ;
  assign n2590 = n2586 & n2589 ;
  assign n2591 = ( n2582 & n2583 ) | ( n2582 & n2590 ) | ( n2583 & n2590 ) ;
  assign n2592 = ( n2573 & n2580 ) | ( n2573 & ~n2581 ) | ( n2580 & ~n2581 ) ;
  assign n2593 = ( n2572 & ~n2581 ) | ( n2572 & n2592 ) | ( ~n2581 & n2592 ) ;
  assign n2594 = ( n2583 & n2590 ) | ( n2583 & ~n2591 ) | ( n2590 & ~n2591 ) ;
  assign n2595 = ( n2582 & ~n2591 ) | ( n2582 & n2594 ) | ( ~n2591 & n2594 ) ;
  assign n2596 = n2581 & n2593 ;
  assign n2597 = n2576 & ~n2579 ;
  assign n2598 = ~n2576 & n2579 ;
  assign n2599 = n2597 | n2598 ;
  assign n2600 = n2586 & ~n2589 ;
  assign n2601 = ~n2586 & n2589 ;
  assign n2602 = n2600 | n2601 ;
  assign n2603 = n2599 & n2602 ;
  assign n2604 = ~n2596 & n2603 ;
  assign n2605 = ( n2593 & n2595 ) | ( n2593 & n2604 ) | ( n2595 & n2604 ) ;
  assign n2606 = ( n2581 & n2591 ) | ( n2581 & n2605 ) | ( n2591 & n2605 ) ;
  assign n2607 = ( x154 & x155 ) | ( x154 & x156 ) | ( x155 & x156 ) ;
  assign n2608 = ( x151 & x152 ) | ( x151 & x153 ) | ( x152 & x153 ) ;
  assign n2609 = ( x151 & ~x152 ) | ( x151 & x153 ) | ( ~x152 & x153 ) ;
  assign n2610 = ( ~x151 & x152 ) | ( ~x151 & n2609 ) | ( x152 & n2609 ) ;
  assign n2611 = ( ~x153 & n2609 ) | ( ~x153 & n2610 ) | ( n2609 & n2610 ) ;
  assign n2612 = ( x154 & ~x155 ) | ( x154 & x156 ) | ( ~x155 & x156 ) ;
  assign n2613 = ( ~x154 & x155 ) | ( ~x154 & n2612 ) | ( x155 & n2612 ) ;
  assign n2614 = ( ~x156 & n2612 ) | ( ~x156 & n2613 ) | ( n2612 & n2613 ) ;
  assign n2615 = n2611 & n2614 ;
  assign n2616 = ( n2607 & n2608 ) | ( n2607 & n2615 ) | ( n2608 & n2615 ) ;
  assign n2617 = ( x160 & x161 ) | ( x160 & x162 ) | ( x161 & x162 ) ;
  assign n2618 = ( x157 & x158 ) | ( x157 & x159 ) | ( x158 & x159 ) ;
  assign n2619 = ( x157 & ~x158 ) | ( x157 & x159 ) | ( ~x158 & x159 ) ;
  assign n2620 = ( ~x157 & x158 ) | ( ~x157 & n2619 ) | ( x158 & n2619 ) ;
  assign n2621 = ( ~x159 & n2619 ) | ( ~x159 & n2620 ) | ( n2619 & n2620 ) ;
  assign n2622 = ( x160 & ~x161 ) | ( x160 & x162 ) | ( ~x161 & x162 ) ;
  assign n2623 = ( ~x160 & x161 ) | ( ~x160 & n2622 ) | ( x161 & n2622 ) ;
  assign n2624 = ( ~x162 & n2622 ) | ( ~x162 & n2623 ) | ( n2622 & n2623 ) ;
  assign n2625 = n2621 & n2624 ;
  assign n2626 = ( n2617 & n2618 ) | ( n2617 & n2625 ) | ( n2618 & n2625 ) ;
  assign n2627 = ( n2608 & n2615 ) | ( n2608 & ~n2616 ) | ( n2615 & ~n2616 ) ;
  assign n2628 = ( n2607 & ~n2616 ) | ( n2607 & n2627 ) | ( ~n2616 & n2627 ) ;
  assign n2629 = ( n2618 & n2625 ) | ( n2618 & ~n2626 ) | ( n2625 & ~n2626 ) ;
  assign n2630 = ( n2617 & ~n2626 ) | ( n2617 & n2629 ) | ( ~n2626 & n2629 ) ;
  assign n2631 = n2616 & n2628 ;
  assign n2632 = n2626 & n2630 ;
  assign n2633 = n2611 & ~n2614 ;
  assign n2634 = ~n2611 & n2614 ;
  assign n2635 = n2633 | n2634 ;
  assign n2636 = n2621 & ~n2624 ;
  assign n2637 = ~n2621 & n2624 ;
  assign n2638 = n2636 | n2637 ;
  assign n2639 = n2635 & n2638 ;
  assign n2640 = ~n2632 & n2639 ;
  assign n2641 = ~n2631 & n2640 ;
  assign n2642 = ~n2630 & n2641 ;
  assign n2643 = ( n2628 & n2630 ) | ( n2628 & n2642 ) | ( n2630 & n2642 ) ;
  assign n2644 = n2630 & n2640 ;
  assign n2645 = ~n2631 & n2644 ;
  assign n2646 = n2643 | n2645 ;
  assign n2647 = ( n2616 & n2626 ) | ( n2616 & n2646 ) | ( n2626 & n2646 ) ;
  assign n2648 = ~n2616 & n2626 ;
  assign n2649 = n2616 & ~n2626 ;
  assign n2650 = n2648 | n2649 ;
  assign n2651 = n2645 | n2650 ;
  assign n2652 = n2643 | n2651 ;
  assign n2653 = n2646 & n2650 ;
  assign n2654 = n2652 & ~n2653 ;
  assign n2655 = ~n2581 & n2591 ;
  assign n2656 = n2581 & ~n2591 ;
  assign n2657 = n2655 | n2656 ;
  assign n2658 = n2605 & n2657 ;
  assign n2659 = n2605 | n2657 ;
  assign n2660 = ~n2658 & n2659 ;
  assign n2661 = n2654 | n2660 ;
  assign n2662 = ( n2628 & n2630 ) | ( n2628 & ~n2641 ) | ( n2630 & ~n2641 ) ;
  assign n2663 = n2628 & ~n2645 ;
  assign n2664 = ( n2630 & ~n2662 ) | ( n2630 & n2663 ) | ( ~n2662 & n2663 ) ;
  assign n2665 = ( n2642 & n2662 ) | ( n2642 & ~n2664 ) | ( n2662 & ~n2664 ) ;
  assign n2666 = n2599 & ~n2602 ;
  assign n2667 = ~n2599 & n2602 ;
  assign n2668 = n2666 | n2667 ;
  assign n2669 = n2635 & ~n2638 ;
  assign n2670 = ~n2635 & n2638 ;
  assign n2671 = n2669 | n2670 ;
  assign n2672 = n2668 & n2671 ;
  assign n2673 = n2595 | n2604 ;
  assign n2674 = ~n2605 & n2673 ;
  assign n2675 = n2595 & n2603 ;
  assign n2676 = ( n2593 & ~n2673 ) | ( n2593 & n2675 ) | ( ~n2673 & n2675 ) ;
  assign n2677 = n2674 | n2676 ;
  assign n2678 = n2672 | n2677 ;
  assign n2679 = ( n2672 & n2674 ) | ( n2672 & n2676 ) | ( n2674 & n2676 ) ;
  assign n2680 = ( n2665 & n2678 ) | ( n2665 & n2679 ) | ( n2678 & n2679 ) ;
  assign n2681 = n2661 & n2680 ;
  assign n2682 = n2654 & n2660 ;
  assign n2683 = n2681 | n2682 ;
  assign n2684 = ( n2606 & n2647 ) | ( n2606 & n2683 ) | ( n2647 & n2683 ) ;
  assign n2685 = n2571 & n2684 ;
  assign n2686 = ~n2606 & n2647 ;
  assign n2687 = n2606 & ~n2647 ;
  assign n2688 = n2686 | n2687 ;
  assign n2689 = n2682 | n2688 ;
  assign n2690 = n2681 | n2689 ;
  assign n2691 = n2683 & n2688 ;
  assign n2692 = n2690 & ~n2691 ;
  assign n2693 = ~n2495 & n2536 ;
  assign n2694 = n2495 & ~n2536 ;
  assign n2695 = n2693 | n2694 ;
  assign n2696 = n2570 | n2695 ;
  assign n2697 = ~n2695 & n2696 ;
  assign n2698 = ( ~n2570 & n2696 ) | ( ~n2570 & n2697 ) | ( n2696 & n2697 ) ;
  assign n2699 = n2692 | n2698 ;
  assign n2700 = ( n2556 & ~n2563 ) | ( n2556 & n2569 ) | ( ~n2563 & n2569 ) ;
  assign n2701 = ( ~n2556 & n2563 ) | ( ~n2556 & n2700 ) | ( n2563 & n2700 ) ;
  assign n2702 = ( ~n2569 & n2700 ) | ( ~n2569 & n2701 ) | ( n2700 & n2701 ) ;
  assign n2703 = ( ~n2654 & n2660 ) | ( ~n2654 & n2680 ) | ( n2660 & n2680 ) ;
  assign n2704 = ( n2654 & ~n2680 ) | ( n2654 & n2703 ) | ( ~n2680 & n2703 ) ;
  assign n2705 = ( ~n2660 & n2703 ) | ( ~n2660 & n2704 ) | ( n2703 & n2704 ) ;
  assign n2706 = n2668 & ~n2671 ;
  assign n2707 = ~n2668 & n2671 ;
  assign n2708 = n2706 | n2707 ;
  assign n2709 = n2543 & ~n2546 ;
  assign n2710 = ~n2543 & n2546 ;
  assign n2711 = n2709 | n2710 ;
  assign n2712 = n2708 & n2711 ;
  assign n2713 = ~n2672 & n2678 ;
  assign n2714 = ( ~n2677 & n2678 ) | ( ~n2677 & n2713 ) | ( n2678 & n2713 ) ;
  assign n2715 = n2665 & ~n2714 ;
  assign n2716 = ~n2665 & n2714 ;
  assign n2717 = n2715 | n2716 ;
  assign n2718 = ( n2540 & n2547 ) | ( n2540 & ~n2552 ) | ( n2547 & ~n2552 ) ;
  assign n2719 = ( ~n2540 & n2552 ) | ( ~n2540 & n2718 ) | ( n2552 & n2718 ) ;
  assign n2720 = ( ~n2547 & n2718 ) | ( ~n2547 & n2719 ) | ( n2718 & n2719 ) ;
  assign n2721 = ( n2712 & n2717 ) | ( n2712 & n2720 ) | ( n2717 & n2720 ) ;
  assign n2722 = ( n2702 & n2705 ) | ( n2702 & n2721 ) | ( n2705 & n2721 ) ;
  assign n2723 = n2699 & n2722 ;
  assign n2724 = n2692 & n2698 ;
  assign n2725 = n2723 | n2724 ;
  assign n2726 = n2684 & ~n2685 ;
  assign n2727 = ( n2571 & ~n2685 ) | ( n2571 & n2726 ) | ( ~n2685 & n2726 ) ;
  assign n2728 = n2725 & n2727 ;
  assign n2729 = ( n2684 & n2725 ) | ( n2684 & n2728 ) | ( n2725 & n2728 ) ;
  assign n2730 = n2685 | n2729 ;
  assign n2731 = n2451 | n2458 ;
  assign n2732 = n2450 | n2731 ;
  assign n2733 = n2452 & n2458 ;
  assign n2734 = n2732 & ~n2733 ;
  assign n2735 = n2724 | n2727 ;
  assign n2736 = n2723 | n2735 ;
  assign n2737 = ~n2728 & n2736 ;
  assign n2738 = ( ~n2429 & n2432 ) | ( ~n2429 & n2448 ) | ( n2432 & n2448 ) ;
  assign n2739 = ( n2429 & ~n2448 ) | ( n2429 & n2738 ) | ( ~n2448 & n2738 ) ;
  assign n2740 = ( ~n2432 & n2738 ) | ( ~n2432 & n2739 ) | ( n2738 & n2739 ) ;
  assign n2741 = ( ~n2702 & n2705 ) | ( ~n2702 & n2721 ) | ( n2705 & n2721 ) ;
  assign n2742 = ( n2702 & ~n2721 ) | ( n2702 & n2741 ) | ( ~n2721 & n2741 ) ;
  assign n2743 = ( ~n2705 & n2741 ) | ( ~n2705 & n2742 ) | ( n2741 & n2742 ) ;
  assign n2744 = n2708 & ~n2711 ;
  assign n2745 = ~n2708 & n2711 ;
  assign n2746 = n2744 | n2745 ;
  assign n2747 = n2435 & ~n2438 ;
  assign n2748 = ~n2435 & n2438 ;
  assign n2749 = n2747 | n2748 ;
  assign n2750 = n2746 & n2749 ;
  assign n2751 = ( n2712 & ~n2717 ) | ( n2712 & n2720 ) | ( ~n2717 & n2720 ) ;
  assign n2752 = ( ~n2712 & n2717 ) | ( ~n2712 & n2751 ) | ( n2717 & n2751 ) ;
  assign n2753 = ( ~n2720 & n2751 ) | ( ~n2720 & n2752 ) | ( n2751 & n2752 ) ;
  assign n2754 = ( n2439 & ~n2444 ) | ( n2439 & n2447 ) | ( ~n2444 & n2447 ) ;
  assign n2755 = ( ~n2439 & n2444 ) | ( ~n2439 & n2754 ) | ( n2444 & n2754 ) ;
  assign n2756 = ( ~n2447 & n2754 ) | ( ~n2447 & n2755 ) | ( n2754 & n2755 ) ;
  assign n2757 = ( n2750 & n2753 ) | ( n2750 & n2756 ) | ( n2753 & n2756 ) ;
  assign n2758 = ( n2740 & n2743 ) | ( n2740 & n2757 ) | ( n2743 & n2757 ) ;
  assign n2759 = ( ~n2692 & n2698 ) | ( ~n2692 & n2722 ) | ( n2698 & n2722 ) ;
  assign n2760 = ( n2692 & ~n2722 ) | ( n2692 & n2759 ) | ( ~n2722 & n2759 ) ;
  assign n2761 = ( ~n2698 & n2759 ) | ( ~n2698 & n2760 ) | ( n2759 & n2760 ) ;
  assign n2762 = ( ~n2309 & n2425 ) | ( ~n2309 & n2449 ) | ( n2425 & n2449 ) ;
  assign n2763 = ( n2309 & ~n2449 ) | ( n2309 & n2762 ) | ( ~n2449 & n2762 ) ;
  assign n2764 = ( ~n2425 & n2762 ) | ( ~n2425 & n2763 ) | ( n2762 & n2763 ) ;
  assign n2765 = ( n2758 & n2761 ) | ( n2758 & n2764 ) | ( n2761 & n2764 ) ;
  assign n2766 = ( n2734 & n2737 ) | ( n2734 & n2765 ) | ( n2737 & n2765 ) ;
  assign n2767 = ( n2460 & n2730 ) | ( n2460 & ~n2766 ) | ( n2730 & ~n2766 ) ;
  assign n2768 = ( ~n2730 & n2766 ) | ( ~n2730 & n2767 ) | ( n2766 & n2767 ) ;
  assign n2769 = ( ~n2460 & n2767 ) | ( ~n2460 & n2768 ) | ( n2767 & n2768 ) ;
  assign n2770 = ( x202 & x203 ) | ( x202 & x204 ) | ( x203 & x204 ) ;
  assign n2771 = ( x199 & ~x200 ) | ( x199 & x201 ) | ( ~x200 & x201 ) ;
  assign n2772 = ( ~x199 & x200 ) | ( ~x199 & n2771 ) | ( x200 & n2771 ) ;
  assign n2773 = ( ~x201 & n2771 ) | ( ~x201 & n2772 ) | ( n2771 & n2772 ) ;
  assign n2774 = ( x202 & ~x203 ) | ( x202 & x204 ) | ( ~x203 & x204 ) ;
  assign n2775 = ( ~x202 & x203 ) | ( ~x202 & n2774 ) | ( x203 & n2774 ) ;
  assign n2776 = ( ~x204 & n2774 ) | ( ~x204 & n2775 ) | ( n2774 & n2775 ) ;
  assign n2777 = n2773 & n2776 ;
  assign n2778 = ( x199 & x200 ) | ( x199 & x201 ) | ( x200 & x201 ) ;
  assign n2779 = ( n2770 & n2777 ) | ( n2770 & n2778 ) | ( n2777 & n2778 ) ;
  assign n2780 = ( n2777 & n2778 ) | ( n2777 & ~n2779 ) | ( n2778 & ~n2779 ) ;
  assign n2781 = ( n2770 & ~n2779 ) | ( n2770 & n2780 ) | ( ~n2779 & n2780 ) ;
  assign n2782 = ( x208 & x209 ) | ( x208 & x210 ) | ( x209 & x210 ) ;
  assign n2783 = ( x205 & x206 ) | ( x205 & x207 ) | ( x206 & x207 ) ;
  assign n2784 = ( x205 & ~x206 ) | ( x205 & x207 ) | ( ~x206 & x207 ) ;
  assign n2785 = ( ~x205 & x206 ) | ( ~x205 & n2784 ) | ( x206 & n2784 ) ;
  assign n2786 = ( ~x207 & n2784 ) | ( ~x207 & n2785 ) | ( n2784 & n2785 ) ;
  assign n2787 = ( x208 & ~x209 ) | ( x208 & x210 ) | ( ~x209 & x210 ) ;
  assign n2788 = ( ~x208 & x209 ) | ( ~x208 & n2787 ) | ( x209 & n2787 ) ;
  assign n2789 = ( ~x210 & n2787 ) | ( ~x210 & n2788 ) | ( n2787 & n2788 ) ;
  assign n2790 = n2786 & n2789 ;
  assign n2791 = ( n2782 & n2783 ) | ( n2782 & n2790 ) | ( n2783 & n2790 ) ;
  assign n2792 = ( n2783 & n2790 ) | ( n2783 & ~n2791 ) | ( n2790 & ~n2791 ) ;
  assign n2793 = ( n2782 & ~n2791 ) | ( n2782 & n2792 ) | ( ~n2791 & n2792 ) ;
  assign n2794 = n2779 & n2781 ;
  assign n2795 = n2791 & n2793 ;
  assign n2796 = n2773 & ~n2776 ;
  assign n2797 = ~n2773 & n2776 ;
  assign n2798 = n2796 | n2797 ;
  assign n2799 = n2786 & ~n2789 ;
  assign n2800 = ~n2786 & n2789 ;
  assign n2801 = n2799 | n2800 ;
  assign n2802 = n2798 & n2801 ;
  assign n2803 = ~n2795 & n2802 ;
  assign n2804 = ~n2794 & n2803 ;
  assign n2805 = ~n2793 & n2804 ;
  assign n2806 = ( n2781 & n2793 ) | ( n2781 & n2805 ) | ( n2793 & n2805 ) ;
  assign n2807 = n2793 & n2803 ;
  assign n2808 = ~n2794 & n2807 ;
  assign n2809 = ~n2779 & n2791 ;
  assign n2810 = n2779 & ~n2791 ;
  assign n2811 = n2809 | n2810 ;
  assign n2812 = n2808 | n2811 ;
  assign n2813 = n2806 | n2812 ;
  assign n2814 = n2806 | n2808 ;
  assign n2815 = n2811 & n2814 ;
  assign n2816 = n2813 & ~n2815 ;
  assign n2817 = ( x220 & x221 ) | ( x220 & x222 ) | ( x221 & x222 ) ;
  assign n2818 = ( x217 & x218 ) | ( x217 & x219 ) | ( x218 & x219 ) ;
  assign n2819 = ( x217 & ~x218 ) | ( x217 & x219 ) | ( ~x218 & x219 ) ;
  assign n2820 = ( ~x217 & x218 ) | ( ~x217 & n2819 ) | ( x218 & n2819 ) ;
  assign n2821 = ( ~x219 & n2819 ) | ( ~x219 & n2820 ) | ( n2819 & n2820 ) ;
  assign n2822 = ( x220 & ~x221 ) | ( x220 & x222 ) | ( ~x221 & x222 ) ;
  assign n2823 = ( ~x220 & x221 ) | ( ~x220 & n2822 ) | ( x221 & n2822 ) ;
  assign n2824 = ( ~x222 & n2822 ) | ( ~x222 & n2823 ) | ( n2822 & n2823 ) ;
  assign n2825 = n2821 & n2824 ;
  assign n2826 = ( n2817 & n2818 ) | ( n2817 & n2825 ) | ( n2818 & n2825 ) ;
  assign n2827 = ( x211 & ~x212 ) | ( x211 & x213 ) | ( ~x212 & x213 ) ;
  assign n2828 = ( ~x211 & x212 ) | ( ~x211 & n2827 ) | ( x212 & n2827 ) ;
  assign n2829 = ( ~x213 & n2827 ) | ( ~x213 & n2828 ) | ( n2827 & n2828 ) ;
  assign n2830 = ( x214 & ~x215 ) | ( x214 & x216 ) | ( ~x215 & x216 ) ;
  assign n2831 = ( ~x214 & x215 ) | ( ~x214 & n2830 ) | ( x215 & n2830 ) ;
  assign n2832 = ( ~x216 & n2830 ) | ( ~x216 & n2831 ) | ( n2830 & n2831 ) ;
  assign n2833 = n2829 & n2832 ;
  assign n2834 = ( x214 & x215 ) | ( x214 & x216 ) | ( x215 & x216 ) ;
  assign n2835 = ( x211 & x212 ) | ( x211 & x213 ) | ( x212 & x213 ) ;
  assign n2836 = ( n2833 & n2834 ) | ( n2833 & n2835 ) | ( n2834 & n2835 ) ;
  assign n2837 = ( n2818 & n2825 ) | ( n2818 & ~n2826 ) | ( n2825 & ~n2826 ) ;
  assign n2838 = ( n2817 & ~n2826 ) | ( n2817 & n2837 ) | ( ~n2826 & n2837 ) ;
  assign n2839 = ( n2833 & n2835 ) | ( n2833 & ~n2836 ) | ( n2835 & ~n2836 ) ;
  assign n2840 = ( n2834 & ~n2836 ) | ( n2834 & n2839 ) | ( ~n2836 & n2839 ) ;
  assign n2841 = n2836 & n2840 ;
  assign n2842 = n2829 & ~n2832 ;
  assign n2843 = ~n2829 & n2832 ;
  assign n2844 = n2842 | n2843 ;
  assign n2845 = n2821 & ~n2824 ;
  assign n2846 = ~n2821 & n2824 ;
  assign n2847 = n2845 | n2846 ;
  assign n2848 = ~n2825 & n2847 ;
  assign n2849 = n2844 & n2848 ;
  assign n2850 = ~n2841 & n2849 ;
  assign n2851 = ( n2838 & n2840 ) | ( n2838 & n2850 ) | ( n2840 & n2850 ) ;
  assign n2852 = ( n2826 & n2836 ) | ( n2826 & ~n2851 ) | ( n2836 & ~n2851 ) ;
  assign n2853 = ( n2826 & ~n2836 ) | ( n2826 & n2851 ) | ( ~n2836 & n2851 ) ;
  assign n2854 = ( ~n2826 & n2852 ) | ( ~n2826 & n2853 ) | ( n2852 & n2853 ) ;
  assign n2855 = n2816 | n2854 ;
  assign n2856 = ( n2781 & n2793 ) | ( n2781 & ~n2804 ) | ( n2793 & ~n2804 ) ;
  assign n2857 = n2781 & ~n2808 ;
  assign n2858 = ( n2793 & ~n2856 ) | ( n2793 & n2857 ) | ( ~n2856 & n2857 ) ;
  assign n2859 = ( n2805 & n2856 ) | ( n2805 & ~n2858 ) | ( n2856 & ~n2858 ) ;
  assign n2860 = n2844 & ~n2848 ;
  assign n2861 = ~n2844 & n2848 ;
  assign n2862 = n2860 | n2861 ;
  assign n2863 = n2798 & ~n2801 ;
  assign n2864 = ~n2798 & n2801 ;
  assign n2865 = n2863 | n2864 ;
  assign n2866 = n2862 & n2865 ;
  assign n2867 = n2838 | n2850 ;
  assign n2868 = ~n2851 & n2867 ;
  assign n2869 = n2838 & n2849 ;
  assign n2870 = ( n2840 & ~n2867 ) | ( n2840 & n2869 ) | ( ~n2867 & n2869 ) ;
  assign n2871 = n2868 | n2870 ;
  assign n2872 = n2866 | n2871 ;
  assign n2873 = ( n2866 & n2868 ) | ( n2866 & n2870 ) | ( n2868 & n2870 ) ;
  assign n2874 = ( n2859 & n2872 ) | ( n2859 & n2873 ) | ( n2872 & n2873 ) ;
  assign n2875 = n2855 & n2874 ;
  assign n2876 = n2816 & n2854 ;
  assign n2877 = ( n2826 & n2836 ) | ( n2826 & n2851 ) | ( n2836 & n2851 ) ;
  assign n2878 = ( n2779 & n2791 ) | ( n2779 & n2814 ) | ( n2791 & n2814 ) ;
  assign n2879 = ~n2877 & n2878 ;
  assign n2880 = n2877 & ~n2878 ;
  assign n2881 = n2879 | n2880 ;
  assign n2882 = n2876 | n2881 ;
  assign n2883 = n2875 | n2882 ;
  assign n2884 = n2875 | n2876 ;
  assign n2885 = n2881 & n2884 ;
  assign n2886 = n2883 & ~n2885 ;
  assign n2922 = ( x184 & x185 ) | ( x184 & x186 ) | ( x185 & x186 ) ;
  assign n2923 = ( x181 & x182 ) | ( x181 & x183 ) | ( x182 & x183 ) ;
  assign n2924 = ( x181 & ~x182 ) | ( x181 & x183 ) | ( ~x182 & x183 ) ;
  assign n2925 = ( ~x181 & x182 ) | ( ~x181 & n2924 ) | ( x182 & n2924 ) ;
  assign n2926 = ( ~x183 & n2924 ) | ( ~x183 & n2925 ) | ( n2924 & n2925 ) ;
  assign n2927 = ( x184 & ~x185 ) | ( x184 & x186 ) | ( ~x185 & x186 ) ;
  assign n2928 = ( ~x184 & x185 ) | ( ~x184 & n2927 ) | ( x185 & n2927 ) ;
  assign n2929 = ( ~x186 & n2927 ) | ( ~x186 & n2928 ) | ( n2927 & n2928 ) ;
  assign n2930 = n2926 & n2929 ;
  assign n2931 = ( n2922 & n2923 ) | ( n2922 & n2930 ) | ( n2923 & n2930 ) ;
  assign n2945 = ( n2923 & n2930 ) | ( n2923 & ~n2931 ) | ( n2930 & ~n2931 ) ;
  assign n2946 = ( n2922 & ~n2931 ) | ( n2922 & n2945 ) | ( ~n2931 & n2945 ) ;
  assign n2932 = ( x178 & x179 ) | ( x178 & x180 ) | ( x179 & x180 ) ;
  assign n2933 = ( x175 & x176 ) | ( x175 & x177 ) | ( x176 & x177 ) ;
  assign n2934 = ( x175 & ~x176 ) | ( x175 & x177 ) | ( ~x176 & x177 ) ;
  assign n2935 = ( ~x175 & x176 ) | ( ~x175 & n2934 ) | ( x176 & n2934 ) ;
  assign n2936 = ( ~x177 & n2934 ) | ( ~x177 & n2935 ) | ( n2934 & n2935 ) ;
  assign n2937 = ( x178 & ~x179 ) | ( x178 & x180 ) | ( ~x179 & x180 ) ;
  assign n2938 = ( ~x178 & x179 ) | ( ~x178 & n2937 ) | ( x179 & n2937 ) ;
  assign n2939 = ( ~x180 & n2937 ) | ( ~x180 & n2938 ) | ( n2937 & n2938 ) ;
  assign n2940 = n2936 & n2939 ;
  assign n2941 = ( n2932 & n2933 ) | ( n2932 & n2940 ) | ( n2933 & n2940 ) ;
  assign n2942 = ( n2933 & n2940 ) | ( n2933 & ~n2941 ) | ( n2940 & ~n2941 ) ;
  assign n2943 = ( n2932 & ~n2941 ) | ( n2932 & n2942 ) | ( ~n2941 & n2942 ) ;
  assign n2944 = n2941 & n2943 ;
  assign n2947 = n2931 & n2946 ;
  assign n2948 = n2926 & ~n2929 ;
  assign n2949 = ~n2926 & n2929 ;
  assign n2950 = n2948 | n2949 ;
  assign n2951 = n2936 & ~n2939 ;
  assign n2952 = ~n2936 & n2939 ;
  assign n2953 = n2951 | n2952 ;
  assign n2954 = n2950 & n2953 ;
  assign n2955 = ~n2947 & n2954 ;
  assign n2958 = ~n2944 & n2955 ;
  assign n2959 = ~n2946 & n2958 ;
  assign n2966 = ( n2943 & n2946 ) | ( n2943 & ~n2958 ) | ( n2946 & ~n2958 ) ;
  assign n2956 = n2946 & n2955 ;
  assign n2957 = ~n2944 & n2956 ;
  assign n2967 = n2943 & ~n2957 ;
  assign n2968 = ( n2946 & ~n2966 ) | ( n2946 & n2967 ) | ( ~n2966 & n2967 ) ;
  assign n2969 = ( n2959 & n2966 ) | ( n2959 & ~n2968 ) | ( n2966 & ~n2968 ) ;
  assign n2889 = ( x187 & ~x188 ) | ( x187 & x189 ) | ( ~x188 & x189 ) ;
  assign n2890 = ( ~x187 & x188 ) | ( ~x187 & n2889 ) | ( x188 & n2889 ) ;
  assign n2891 = ( ~x189 & n2889 ) | ( ~x189 & n2890 ) | ( n2889 & n2890 ) ;
  assign n2892 = ( x190 & ~x191 ) | ( x190 & x192 ) | ( ~x191 & x192 ) ;
  assign n2893 = ( ~x190 & x191 ) | ( ~x190 & n2892 ) | ( x191 & n2892 ) ;
  assign n2894 = ( ~x192 & n2892 ) | ( ~x192 & n2893 ) | ( n2892 & n2893 ) ;
  assign n2912 = n2891 & ~n2894 ;
  assign n2913 = ~n2891 & n2894 ;
  assign n2914 = n2912 | n2913 ;
  assign n2899 = ( x193 & ~x194 ) | ( x193 & x195 ) | ( ~x194 & x195 ) ;
  assign n2900 = ( ~x193 & x194 ) | ( ~x193 & n2899 ) | ( x194 & n2899 ) ;
  assign n2901 = ( ~x195 & n2899 ) | ( ~x195 & n2900 ) | ( n2899 & n2900 ) ;
  assign n2902 = ( x196 & ~x197 ) | ( x196 & x198 ) | ( ~x197 & x198 ) ;
  assign n2903 = ( ~x196 & x197 ) | ( ~x196 & n2902 ) | ( x197 & n2902 ) ;
  assign n2904 = ( ~x198 & n2902 ) | ( ~x198 & n2903 ) | ( n2902 & n2903 ) ;
  assign n2915 = n2901 & ~n2904 ;
  assign n2916 = ~n2901 & n2904 ;
  assign n2917 = n2915 | n2916 ;
  assign n2970 = n2914 & ~n2917 ;
  assign n2971 = ~n2914 & n2917 ;
  assign n2972 = n2970 | n2971 ;
  assign n2973 = ~n2950 & n2953 ;
  assign n2974 = n2950 & ~n2953 ;
  assign n2975 = n2973 | n2974 ;
  assign n2976 = n2972 & n2975 ;
  assign n2887 = ( x190 & x191 ) | ( x190 & x192 ) | ( x191 & x192 ) ;
  assign n2888 = ( x187 & x188 ) | ( x187 & x189 ) | ( x188 & x189 ) ;
  assign n2895 = n2891 & n2894 ;
  assign n2896 = ( n2887 & n2888 ) | ( n2887 & n2895 ) | ( n2888 & n2895 ) ;
  assign n2907 = ( n2888 & n2895 ) | ( n2888 & ~n2896 ) | ( n2895 & ~n2896 ) ;
  assign n2908 = ( n2887 & ~n2896 ) | ( n2887 & n2907 ) | ( ~n2896 & n2907 ) ;
  assign n2897 = ( x196 & x197 ) | ( x196 & x198 ) | ( x197 & x198 ) ;
  assign n2898 = ( x193 & x194 ) | ( x193 & x195 ) | ( x194 & x195 ) ;
  assign n2905 = n2901 & n2904 ;
  assign n2906 = ( n2897 & n2898 ) | ( n2897 & n2905 ) | ( n2898 & n2905 ) ;
  assign n2909 = ( n2898 & n2905 ) | ( n2898 & ~n2906 ) | ( n2905 & ~n2906 ) ;
  assign n2910 = ( n2897 & ~n2906 ) | ( n2897 & n2909 ) | ( ~n2906 & n2909 ) ;
  assign n2918 = n2914 & n2917 ;
  assign n2977 = n2910 & n2918 ;
  assign n2911 = n2896 & n2908 ;
  assign n2919 = ~n2911 & n2918 ;
  assign n2978 = n2910 | n2919 ;
  assign n2979 = ( n2908 & n2977 ) | ( n2908 & ~n2978 ) | ( n2977 & ~n2978 ) ;
  assign n2920 = ( n2908 & n2910 ) | ( n2908 & n2919 ) | ( n2910 & n2919 ) ;
  assign n2980 = ~n2920 & n2978 ;
  assign n2981 = n2979 | n2980 ;
  assign n2982 = n2976 | n2981 ;
  assign n2983 = n2969 & n2982 ;
  assign n2984 = ( n2976 & n2979 ) | ( n2976 & n2980 ) | ( n2979 & n2980 ) ;
  assign n2985 = n2983 | n2984 ;
  assign n2960 = ( n2943 & n2946 ) | ( n2943 & n2959 ) | ( n2946 & n2959 ) ;
  assign n2986 = n2931 & ~n2941 ;
  assign n2987 = ~n2931 & n2941 ;
  assign n2988 = n2986 | n2987 ;
  assign n2989 = n2957 | n2988 ;
  assign n2990 = n2960 | n2989 ;
  assign n2961 = n2957 | n2960 ;
  assign n2991 = n2961 & n2988 ;
  assign n2992 = n2990 & ~n2991 ;
  assign n2993 = ~n2896 & n2906 ;
  assign n2994 = n2896 & ~n2906 ;
  assign n2995 = n2993 | n2994 ;
  assign n2996 = n2920 & n2995 ;
  assign n2997 = n2920 | n2995 ;
  assign n2998 = ~n2996 & n2997 ;
  assign n2999 = ( n2985 & n2992 ) | ( n2985 & n2998 ) | ( n2992 & n2998 ) ;
  assign n2921 = ( n2896 & n2906 ) | ( n2896 & n2920 ) | ( n2906 & n2920 ) ;
  assign n2962 = ( n2931 & n2941 ) | ( n2931 & n2961 ) | ( n2941 & n2961 ) ;
  assign n2963 = n2921 & n2962 ;
  assign n2964 = n2962 & ~n2963 ;
  assign n2965 = ( n2921 & ~n2963 ) | ( n2921 & n2964 ) | ( ~n2963 & n2964 ) ;
  assign n3000 = n2965 | n2999 ;
  assign n3001 = ~n2965 & n3000 ;
  assign n3002 = ( ~n2999 & n3000 ) | ( ~n2999 & n3001 ) | ( n3000 & n3001 ) ;
  assign n3003 = n2886 | n3002 ;
  assign n3004 = ( n2985 & ~n2992 ) | ( n2985 & n2998 ) | ( ~n2992 & n2998 ) ;
  assign n3005 = ( ~n2985 & n2992 ) | ( ~n2985 & n3004 ) | ( n2992 & n3004 ) ;
  assign n3006 = ( ~n2998 & n3004 ) | ( ~n2998 & n3005 ) | ( n3004 & n3005 ) ;
  assign n3007 = ( ~n2816 & n2854 ) | ( ~n2816 & n2874 ) | ( n2854 & n2874 ) ;
  assign n3008 = ( n2816 & ~n2874 ) | ( n2816 & n3007 ) | ( ~n2874 & n3007 ) ;
  assign n3009 = ( ~n2854 & n3007 ) | ( ~n2854 & n3008 ) | ( n3007 & n3008 ) ;
  assign n3010 = n2862 & ~n2865 ;
  assign n3011 = ~n2862 & n2865 ;
  assign n3012 = n3010 | n3011 ;
  assign n3013 = n2972 & ~n2975 ;
  assign n3014 = ~n2972 & n2975 ;
  assign n3015 = n3013 | n3014 ;
  assign n3016 = n3012 & n3015 ;
  assign n3017 = ~n2866 & n2872 ;
  assign n3018 = ( ~n2871 & n2872 ) | ( ~n2871 & n3017 ) | ( n2872 & n3017 ) ;
  assign n3019 = n2859 & ~n3018 ;
  assign n3020 = ~n2859 & n3018 ;
  assign n3021 = n3019 | n3020 ;
  assign n3022 = ( n2969 & n2976 ) | ( n2969 & ~n2981 ) | ( n2976 & ~n2981 ) ;
  assign n3023 = ( ~n2969 & n2981 ) | ( ~n2969 & n3022 ) | ( n2981 & n3022 ) ;
  assign n3024 = ( ~n2976 & n3022 ) | ( ~n2976 & n3023 ) | ( n3022 & n3023 ) ;
  assign n3025 = ( n3016 & n3021 ) | ( n3016 & n3024 ) | ( n3021 & n3024 ) ;
  assign n3026 = ( n3006 & n3009 ) | ( n3006 & n3025 ) | ( n3009 & n3025 ) ;
  assign n3027 = n3003 & n3026 ;
  assign n3028 = n2886 & n3002 ;
  assign n3029 = n2963 | n2965 ;
  assign n3030 = ( n2963 & n2999 ) | ( n2963 & n3029 ) | ( n2999 & n3029 ) ;
  assign n3031 = ( n2877 & n2878 ) | ( n2877 & n2884 ) | ( n2878 & n2884 ) ;
  assign n3032 = n3030 & n3031 ;
  assign n3033 = n3031 & ~n3032 ;
  assign n3034 = ( n3030 & ~n3032 ) | ( n3030 & n3033 ) | ( ~n3032 & n3033 ) ;
  assign n3035 = n3028 | n3034 ;
  assign n3036 = n3027 | n3035 ;
  assign n3037 = n3027 | n3028 ;
  assign n3038 = n3034 & n3037 ;
  assign n3039 = n3036 & ~n3038 ;
  assign n3040 = ( x250 & x251 ) | ( x250 & x252 ) | ( x251 & x252 ) ;
  assign n3041 = ( x247 & ~x248 ) | ( x247 & x249 ) | ( ~x248 & x249 ) ;
  assign n3042 = ( ~x247 & x248 ) | ( ~x247 & n3041 ) | ( x248 & n3041 ) ;
  assign n3043 = ( ~x249 & n3041 ) | ( ~x249 & n3042 ) | ( n3041 & n3042 ) ;
  assign n3044 = ( x250 & ~x251 ) | ( x250 & x252 ) | ( ~x251 & x252 ) ;
  assign n3045 = ( ~x250 & x251 ) | ( ~x250 & n3044 ) | ( x251 & n3044 ) ;
  assign n3046 = ( ~x252 & n3044 ) | ( ~x252 & n3045 ) | ( n3044 & n3045 ) ;
  assign n3047 = n3043 & n3046 ;
  assign n3048 = ( x247 & x248 ) | ( x247 & x249 ) | ( x248 & x249 ) ;
  assign n3049 = ( n3040 & n3047 ) | ( n3040 & n3048 ) | ( n3047 & n3048 ) ;
  assign n3050 = ( n3047 & n3048 ) | ( n3047 & ~n3049 ) | ( n3048 & ~n3049 ) ;
  assign n3051 = ( n3040 & ~n3049 ) | ( n3040 & n3050 ) | ( ~n3049 & n3050 ) ;
  assign n3052 = ( x256 & x257 ) | ( x256 & x258 ) | ( x257 & x258 ) ;
  assign n3053 = ( x253 & x254 ) | ( x253 & x255 ) | ( x254 & x255 ) ;
  assign n3054 = ( x253 & ~x254 ) | ( x253 & x255 ) | ( ~x254 & x255 ) ;
  assign n3055 = ( ~x253 & x254 ) | ( ~x253 & n3054 ) | ( x254 & n3054 ) ;
  assign n3056 = ( ~x255 & n3054 ) | ( ~x255 & n3055 ) | ( n3054 & n3055 ) ;
  assign n3057 = ( x256 & ~x257 ) | ( x256 & x258 ) | ( ~x257 & x258 ) ;
  assign n3058 = ( ~x256 & x257 ) | ( ~x256 & n3057 ) | ( x257 & n3057 ) ;
  assign n3059 = ( ~x258 & n3057 ) | ( ~x258 & n3058 ) | ( n3057 & n3058 ) ;
  assign n3060 = n3056 & n3059 ;
  assign n3061 = ( n3052 & n3053 ) | ( n3052 & n3060 ) | ( n3053 & n3060 ) ;
  assign n3062 = ( n3053 & n3060 ) | ( n3053 & ~n3061 ) | ( n3060 & ~n3061 ) ;
  assign n3063 = ( n3052 & ~n3061 ) | ( n3052 & n3062 ) | ( ~n3061 & n3062 ) ;
  assign n3064 = n3049 & n3051 ;
  assign n3065 = n3061 & n3063 ;
  assign n3066 = n3043 & ~n3046 ;
  assign n3067 = ~n3043 & n3046 ;
  assign n3068 = n3066 | n3067 ;
  assign n3069 = n3056 & ~n3059 ;
  assign n3070 = ~n3056 & n3059 ;
  assign n3071 = n3069 | n3070 ;
  assign n3072 = n3068 & n3071 ;
  assign n3073 = ~n3065 & n3072 ;
  assign n3074 = ~n3064 & n3073 ;
  assign n3075 = ~n3063 & n3074 ;
  assign n3076 = ( n3051 & n3063 ) | ( n3051 & n3075 ) | ( n3063 & n3075 ) ;
  assign n3077 = n3063 & n3073 ;
  assign n3078 = ~n3064 & n3077 ;
  assign n3079 = ~n3049 & n3061 ;
  assign n3080 = n3049 & ~n3061 ;
  assign n3081 = n3079 | n3080 ;
  assign n3082 = n3078 | n3081 ;
  assign n3083 = n3076 | n3082 ;
  assign n3084 = n3076 | n3078 ;
  assign n3085 = n3081 & n3084 ;
  assign n3086 = n3083 & ~n3085 ;
  assign n3087 = ( x268 & x269 ) | ( x268 & x270 ) | ( x269 & x270 ) ;
  assign n3088 = ( x265 & x266 ) | ( x265 & x267 ) | ( x266 & x267 ) ;
  assign n3089 = ( x265 & ~x266 ) | ( x265 & x267 ) | ( ~x266 & x267 ) ;
  assign n3090 = ( ~x265 & x266 ) | ( ~x265 & n3089 ) | ( x266 & n3089 ) ;
  assign n3091 = ( ~x267 & n3089 ) | ( ~x267 & n3090 ) | ( n3089 & n3090 ) ;
  assign n3092 = ( x268 & ~x269 ) | ( x268 & x270 ) | ( ~x269 & x270 ) ;
  assign n3093 = ( ~x268 & x269 ) | ( ~x268 & n3092 ) | ( x269 & n3092 ) ;
  assign n3094 = ( ~x270 & n3092 ) | ( ~x270 & n3093 ) | ( n3092 & n3093 ) ;
  assign n3095 = n3091 & n3094 ;
  assign n3096 = ( n3087 & n3088 ) | ( n3087 & n3095 ) | ( n3088 & n3095 ) ;
  assign n3097 = ( x259 & ~x260 ) | ( x259 & x261 ) | ( ~x260 & x261 ) ;
  assign n3098 = ( ~x259 & x260 ) | ( ~x259 & n3097 ) | ( x260 & n3097 ) ;
  assign n3099 = ( ~x261 & n3097 ) | ( ~x261 & n3098 ) | ( n3097 & n3098 ) ;
  assign n3100 = ( x262 & ~x263 ) | ( x262 & x264 ) | ( ~x263 & x264 ) ;
  assign n3101 = ( ~x262 & x263 ) | ( ~x262 & n3100 ) | ( x263 & n3100 ) ;
  assign n3102 = ( ~x264 & n3100 ) | ( ~x264 & n3101 ) | ( n3100 & n3101 ) ;
  assign n3103 = n3099 & n3102 ;
  assign n3104 = ( x262 & x263 ) | ( x262 & x264 ) | ( x263 & x264 ) ;
  assign n3105 = ( x259 & x260 ) | ( x259 & x261 ) | ( x260 & x261 ) ;
  assign n3106 = ( n3103 & n3104 ) | ( n3103 & n3105 ) | ( n3104 & n3105 ) ;
  assign n3107 = ( n3088 & n3095 ) | ( n3088 & ~n3096 ) | ( n3095 & ~n3096 ) ;
  assign n3108 = ( n3087 & ~n3096 ) | ( n3087 & n3107 ) | ( ~n3096 & n3107 ) ;
  assign n3109 = ( n3103 & n3105 ) | ( n3103 & ~n3106 ) | ( n3105 & ~n3106 ) ;
  assign n3110 = ( n3104 & ~n3106 ) | ( n3104 & n3109 ) | ( ~n3106 & n3109 ) ;
  assign n3111 = n3106 & n3110 ;
  assign n3112 = n3099 & ~n3102 ;
  assign n3113 = ~n3099 & n3102 ;
  assign n3114 = n3112 | n3113 ;
  assign n3115 = n3091 & ~n3094 ;
  assign n3116 = ~n3091 & n3094 ;
  assign n3117 = n3115 | n3116 ;
  assign n3118 = ~n3095 & n3117 ;
  assign n3119 = n3114 & n3118 ;
  assign n3120 = ~n3111 & n3119 ;
  assign n3121 = ( n3108 & n3110 ) | ( n3108 & n3120 ) | ( n3110 & n3120 ) ;
  assign n3122 = ( n3096 & n3106 ) | ( n3096 & ~n3121 ) | ( n3106 & ~n3121 ) ;
  assign n3123 = ( n3096 & ~n3106 ) | ( n3096 & n3121 ) | ( ~n3106 & n3121 ) ;
  assign n3124 = ( ~n3096 & n3122 ) | ( ~n3096 & n3123 ) | ( n3122 & n3123 ) ;
  assign n3125 = n3086 | n3124 ;
  assign n3126 = ( n3051 & n3063 ) | ( n3051 & ~n3074 ) | ( n3063 & ~n3074 ) ;
  assign n3127 = n3051 & ~n3078 ;
  assign n3128 = ( n3063 & ~n3126 ) | ( n3063 & n3127 ) | ( ~n3126 & n3127 ) ;
  assign n3129 = ( n3075 & n3126 ) | ( n3075 & ~n3128 ) | ( n3126 & ~n3128 ) ;
  assign n3130 = n3114 & ~n3118 ;
  assign n3131 = ~n3114 & n3118 ;
  assign n3132 = n3130 | n3131 ;
  assign n3133 = n3068 & ~n3071 ;
  assign n3134 = ~n3068 & n3071 ;
  assign n3135 = n3133 | n3134 ;
  assign n3136 = n3132 & n3135 ;
  assign n3137 = n3108 | n3120 ;
  assign n3138 = ~n3121 & n3137 ;
  assign n3139 = n3108 & n3119 ;
  assign n3140 = ( n3110 & ~n3137 ) | ( n3110 & n3139 ) | ( ~n3137 & n3139 ) ;
  assign n3141 = n3138 | n3140 ;
  assign n3142 = n3136 | n3141 ;
  assign n3143 = ( n3136 & n3138 ) | ( n3136 & n3140 ) | ( n3138 & n3140 ) ;
  assign n3144 = ( n3129 & n3142 ) | ( n3129 & n3143 ) | ( n3142 & n3143 ) ;
  assign n3145 = n3125 & n3144 ;
  assign n3146 = n3086 & n3124 ;
  assign n3147 = ( n3096 & n3106 ) | ( n3096 & n3121 ) | ( n3106 & n3121 ) ;
  assign n3148 = ( n3049 & n3061 ) | ( n3049 & n3084 ) | ( n3061 & n3084 ) ;
  assign n3149 = ~n3147 & n3148 ;
  assign n3150 = n3147 & ~n3148 ;
  assign n3151 = n3149 | n3150 ;
  assign n3152 = n3146 | n3151 ;
  assign n3153 = n3145 | n3152 ;
  assign n3154 = n3145 | n3146 ;
  assign n3155 = n3151 & n3154 ;
  assign n3156 = n3153 & ~n3155 ;
  assign n3192 = ( x232 & x233 ) | ( x232 & x234 ) | ( x233 & x234 ) ;
  assign n3193 = ( x229 & x230 ) | ( x229 & x231 ) | ( x230 & x231 ) ;
  assign n3194 = ( x229 & ~x230 ) | ( x229 & x231 ) | ( ~x230 & x231 ) ;
  assign n3195 = ( ~x229 & x230 ) | ( ~x229 & n3194 ) | ( x230 & n3194 ) ;
  assign n3196 = ( ~x231 & n3194 ) | ( ~x231 & n3195 ) | ( n3194 & n3195 ) ;
  assign n3197 = ( x232 & ~x233 ) | ( x232 & x234 ) | ( ~x233 & x234 ) ;
  assign n3198 = ( ~x232 & x233 ) | ( ~x232 & n3197 ) | ( x233 & n3197 ) ;
  assign n3199 = ( ~x234 & n3197 ) | ( ~x234 & n3198 ) | ( n3197 & n3198 ) ;
  assign n3200 = n3196 & n3199 ;
  assign n3201 = ( n3192 & n3193 ) | ( n3192 & n3200 ) | ( n3193 & n3200 ) ;
  assign n3215 = ( n3193 & n3200 ) | ( n3193 & ~n3201 ) | ( n3200 & ~n3201 ) ;
  assign n3216 = ( n3192 & ~n3201 ) | ( n3192 & n3215 ) | ( ~n3201 & n3215 ) ;
  assign n3202 = ( x226 & x227 ) | ( x226 & x228 ) | ( x227 & x228 ) ;
  assign n3203 = ( x223 & x224 ) | ( x223 & x225 ) | ( x224 & x225 ) ;
  assign n3204 = ( x223 & ~x224 ) | ( x223 & x225 ) | ( ~x224 & x225 ) ;
  assign n3205 = ( ~x223 & x224 ) | ( ~x223 & n3204 ) | ( x224 & n3204 ) ;
  assign n3206 = ( ~x225 & n3204 ) | ( ~x225 & n3205 ) | ( n3204 & n3205 ) ;
  assign n3207 = ( x226 & ~x227 ) | ( x226 & x228 ) | ( ~x227 & x228 ) ;
  assign n3208 = ( ~x226 & x227 ) | ( ~x226 & n3207 ) | ( x227 & n3207 ) ;
  assign n3209 = ( ~x228 & n3207 ) | ( ~x228 & n3208 ) | ( n3207 & n3208 ) ;
  assign n3210 = n3206 & n3209 ;
  assign n3211 = ( n3202 & n3203 ) | ( n3202 & n3210 ) | ( n3203 & n3210 ) ;
  assign n3212 = ( n3203 & n3210 ) | ( n3203 & ~n3211 ) | ( n3210 & ~n3211 ) ;
  assign n3213 = ( n3202 & ~n3211 ) | ( n3202 & n3212 ) | ( ~n3211 & n3212 ) ;
  assign n3214 = n3211 & n3213 ;
  assign n3217 = n3201 & n3216 ;
  assign n3218 = n3196 & ~n3199 ;
  assign n3219 = ~n3196 & n3199 ;
  assign n3220 = n3218 | n3219 ;
  assign n3221 = n3206 & ~n3209 ;
  assign n3222 = ~n3206 & n3209 ;
  assign n3223 = n3221 | n3222 ;
  assign n3224 = n3220 & n3223 ;
  assign n3225 = ~n3217 & n3224 ;
  assign n3228 = ~n3214 & n3225 ;
  assign n3229 = ~n3216 & n3228 ;
  assign n3236 = ( n3213 & n3216 ) | ( n3213 & ~n3228 ) | ( n3216 & ~n3228 ) ;
  assign n3226 = n3216 & n3225 ;
  assign n3227 = ~n3214 & n3226 ;
  assign n3237 = n3213 & ~n3227 ;
  assign n3238 = ( n3216 & ~n3236 ) | ( n3216 & n3237 ) | ( ~n3236 & n3237 ) ;
  assign n3239 = ( n3229 & n3236 ) | ( n3229 & ~n3238 ) | ( n3236 & ~n3238 ) ;
  assign n3159 = ( x241 & ~x242 ) | ( x241 & x243 ) | ( ~x242 & x243 ) ;
  assign n3160 = ( ~x241 & x242 ) | ( ~x241 & n3159 ) | ( x242 & n3159 ) ;
  assign n3161 = ( ~x243 & n3159 ) | ( ~x243 & n3160 ) | ( n3159 & n3160 ) ;
  assign n3162 = ( x244 & ~x245 ) | ( x244 & x246 ) | ( ~x245 & x246 ) ;
  assign n3163 = ( ~x244 & x245 ) | ( ~x244 & n3162 ) | ( x245 & n3162 ) ;
  assign n3164 = ( ~x246 & n3162 ) | ( ~x246 & n3163 ) | ( n3162 & n3163 ) ;
  assign n3182 = n3161 & ~n3164 ;
  assign n3183 = ~n3161 & n3164 ;
  assign n3184 = n3182 | n3183 ;
  assign n3167 = ( x235 & ~x236 ) | ( x235 & x237 ) | ( ~x236 & x237 ) ;
  assign n3168 = ( ~x235 & x236 ) | ( ~x235 & n3167 ) | ( x236 & n3167 ) ;
  assign n3169 = ( ~x237 & n3167 ) | ( ~x237 & n3168 ) | ( n3167 & n3168 ) ;
  assign n3170 = ( x238 & ~x239 ) | ( x238 & x240 ) | ( ~x239 & x240 ) ;
  assign n3171 = ( ~x238 & x239 ) | ( ~x238 & n3170 ) | ( x239 & n3170 ) ;
  assign n3172 = ( ~x240 & n3170 ) | ( ~x240 & n3171 ) | ( n3170 & n3171 ) ;
  assign n3185 = n3169 & ~n3172 ;
  assign n3186 = ~n3169 & n3172 ;
  assign n3187 = n3185 | n3186 ;
  assign n3240 = ~n3184 & n3187 ;
  assign n3241 = n3184 & ~n3187 ;
  assign n3242 = n3240 | n3241 ;
  assign n3243 = ~n3220 & n3223 ;
  assign n3244 = n3220 & ~n3223 ;
  assign n3245 = n3243 | n3244 ;
  assign n3246 = n3242 & n3245 ;
  assign n3174 = ( x238 & x239 ) | ( x238 & x240 ) | ( x239 & x240 ) ;
  assign n3173 = n3169 & n3172 ;
  assign n3175 = ( x235 & x236 ) | ( x235 & x237 ) | ( x236 & x237 ) ;
  assign n3176 = ( n3173 & n3174 ) | ( n3173 & n3175 ) | ( n3174 & n3175 ) ;
  assign n3179 = ( n3173 & n3175 ) | ( n3173 & ~n3176 ) | ( n3175 & ~n3176 ) ;
  assign n3180 = ( n3174 & ~n3176 ) | ( n3174 & n3179 ) | ( ~n3176 & n3179 ) ;
  assign n3157 = ( x244 & x245 ) | ( x244 & x246 ) | ( x245 & x246 ) ;
  assign n3158 = ( x241 & x242 ) | ( x241 & x243 ) | ( x242 & x243 ) ;
  assign n3165 = n3161 & n3164 ;
  assign n3166 = ( n3157 & n3158 ) | ( n3157 & n3165 ) | ( n3158 & n3165 ) ;
  assign n3177 = ( n3158 & n3165 ) | ( n3158 & ~n3166 ) | ( n3165 & ~n3166 ) ;
  assign n3178 = ( n3157 & ~n3166 ) | ( n3157 & n3177 ) | ( ~n3166 & n3177 ) ;
  assign n3188 = n3184 & n3187 ;
  assign n3247 = n3178 & n3188 ;
  assign n3181 = n3176 & n3180 ;
  assign n3189 = ~n3181 & n3188 ;
  assign n3248 = n3178 | n3189 ;
  assign n3249 = ( n3180 & n3247 ) | ( n3180 & ~n3248 ) | ( n3247 & ~n3248 ) ;
  assign n3190 = ( n3178 & n3180 ) | ( n3178 & n3189 ) | ( n3180 & n3189 ) ;
  assign n3250 = ~n3190 & n3248 ;
  assign n3251 = n3249 | n3250 ;
  assign n3252 = n3246 | n3251 ;
  assign n3253 = n3239 & n3252 ;
  assign n3254 = ( n3246 & n3249 ) | ( n3246 & n3250 ) | ( n3249 & n3250 ) ;
  assign n3255 = n3253 | n3254 ;
  assign n3230 = ( n3213 & n3216 ) | ( n3213 & n3229 ) | ( n3216 & n3229 ) ;
  assign n3256 = n3201 & ~n3211 ;
  assign n3257 = ~n3201 & n3211 ;
  assign n3258 = n3256 | n3257 ;
  assign n3259 = n3227 | n3258 ;
  assign n3260 = n3230 | n3259 ;
  assign n3231 = n3227 | n3230 ;
  assign n3261 = n3231 & n3258 ;
  assign n3262 = n3260 & ~n3261 ;
  assign n3263 = ( n3166 & n3176 ) | ( n3166 & ~n3190 ) | ( n3176 & ~n3190 ) ;
  assign n3264 = ( n3166 & ~n3176 ) | ( n3166 & n3190 ) | ( ~n3176 & n3190 ) ;
  assign n3265 = ( ~n3166 & n3263 ) | ( ~n3166 & n3264 ) | ( n3263 & n3264 ) ;
  assign n3266 = ( n3255 & n3262 ) | ( n3255 & n3265 ) | ( n3262 & n3265 ) ;
  assign n3191 = ( n3166 & n3176 ) | ( n3166 & n3190 ) | ( n3176 & n3190 ) ;
  assign n3232 = ( n3201 & n3211 ) | ( n3201 & n3231 ) | ( n3211 & n3231 ) ;
  assign n3233 = ~n3191 & n3232 ;
  assign n3234 = n3191 & ~n3232 ;
  assign n3235 = n3233 | n3234 ;
  assign n3267 = n3235 | n3266 ;
  assign n3268 = ~n3235 & n3267 ;
  assign n3269 = ( ~n3266 & n3267 ) | ( ~n3266 & n3268 ) | ( n3267 & n3268 ) ;
  assign n3270 = n3156 | n3269 ;
  assign n3271 = ( n3255 & ~n3262 ) | ( n3255 & n3265 ) | ( ~n3262 & n3265 ) ;
  assign n3272 = ( ~n3255 & n3262 ) | ( ~n3255 & n3271 ) | ( n3262 & n3271 ) ;
  assign n3273 = ( ~n3265 & n3271 ) | ( ~n3265 & n3272 ) | ( n3271 & n3272 ) ;
  assign n3274 = ( ~n3086 & n3124 ) | ( ~n3086 & n3144 ) | ( n3124 & n3144 ) ;
  assign n3275 = ( n3086 & ~n3144 ) | ( n3086 & n3274 ) | ( ~n3144 & n3274 ) ;
  assign n3276 = ( ~n3124 & n3274 ) | ( ~n3124 & n3275 ) | ( n3274 & n3275 ) ;
  assign n3277 = n3132 & ~n3135 ;
  assign n3278 = ~n3132 & n3135 ;
  assign n3279 = n3277 | n3278 ;
  assign n3280 = n3242 & ~n3245 ;
  assign n3281 = ~n3242 & n3245 ;
  assign n3282 = n3280 | n3281 ;
  assign n3283 = n3279 & n3282 ;
  assign n3284 = ~n3136 & n3142 ;
  assign n3285 = ( ~n3141 & n3142 ) | ( ~n3141 & n3284 ) | ( n3142 & n3284 ) ;
  assign n3286 = n3129 & ~n3285 ;
  assign n3287 = ~n3129 & n3285 ;
  assign n3288 = n3286 | n3287 ;
  assign n3289 = ( n3239 & n3246 ) | ( n3239 & ~n3251 ) | ( n3246 & ~n3251 ) ;
  assign n3290 = ( ~n3239 & n3251 ) | ( ~n3239 & n3289 ) | ( n3251 & n3289 ) ;
  assign n3291 = ( ~n3246 & n3289 ) | ( ~n3246 & n3290 ) | ( n3289 & n3290 ) ;
  assign n3292 = ( n3283 & n3288 ) | ( n3283 & n3291 ) | ( n3288 & n3291 ) ;
  assign n3293 = ( n3273 & n3276 ) | ( n3273 & n3292 ) | ( n3276 & n3292 ) ;
  assign n3294 = n3270 & n3293 ;
  assign n3295 = n3156 & n3269 ;
  assign n3296 = n3294 | n3295 ;
  assign n3297 = ( n3191 & n3232 ) | ( n3191 & n3266 ) | ( n3232 & n3266 ) ;
  assign n3298 = ( n3147 & n3148 ) | ( n3147 & n3154 ) | ( n3148 & n3154 ) ;
  assign n3299 = n3297 & n3298 ;
  assign n3300 = n3298 & ~n3299 ;
  assign n3301 = ( n3297 & ~n3299 ) | ( n3297 & n3300 ) | ( ~n3299 & n3300 ) ;
  assign n3302 = n3296 & n3301 ;
  assign n3303 = n3295 | n3301 ;
  assign n3304 = n3294 | n3303 ;
  assign n3305 = ~n3302 & n3304 ;
  assign n3306 = n3039 | n3305 ;
  assign n3307 = ( ~n3006 & n3009 ) | ( ~n3006 & n3025 ) | ( n3009 & n3025 ) ;
  assign n3308 = ( n3006 & ~n3025 ) | ( n3006 & n3307 ) | ( ~n3025 & n3307 ) ;
  assign n3309 = ( ~n3009 & n3307 ) | ( ~n3009 & n3308 ) | ( n3307 & n3308 ) ;
  assign n3310 = ( ~n3273 & n3276 ) | ( ~n3273 & n3292 ) | ( n3276 & n3292 ) ;
  assign n3311 = ( n3273 & ~n3292 ) | ( n3273 & n3310 ) | ( ~n3292 & n3310 ) ;
  assign n3312 = ( ~n3276 & n3310 ) | ( ~n3276 & n3311 ) | ( n3310 & n3311 ) ;
  assign n3313 = n3279 & ~n3282 ;
  assign n3314 = ~n3279 & n3282 ;
  assign n3315 = n3313 | n3314 ;
  assign n3316 = n3012 & ~n3015 ;
  assign n3317 = ~n3012 & n3015 ;
  assign n3318 = n3316 | n3317 ;
  assign n3319 = n3315 & n3318 ;
  assign n3320 = ( n3283 & ~n3288 ) | ( n3283 & n3291 ) | ( ~n3288 & n3291 ) ;
  assign n3321 = ( ~n3283 & n3288 ) | ( ~n3283 & n3320 ) | ( n3288 & n3320 ) ;
  assign n3322 = ( ~n3291 & n3320 ) | ( ~n3291 & n3321 ) | ( n3320 & n3321 ) ;
  assign n3323 = ( n3016 & ~n3021 ) | ( n3016 & n3024 ) | ( ~n3021 & n3024 ) ;
  assign n3324 = ( ~n3016 & n3021 ) | ( ~n3016 & n3323 ) | ( n3021 & n3323 ) ;
  assign n3325 = ( ~n3024 & n3323 ) | ( ~n3024 & n3324 ) | ( n3323 & n3324 ) ;
  assign n3326 = ( n3319 & n3322 ) | ( n3319 & n3325 ) | ( n3322 & n3325 ) ;
  assign n3327 = ( n3309 & n3312 ) | ( n3309 & n3326 ) | ( n3312 & n3326 ) ;
  assign n3328 = ( ~n3156 & n3269 ) | ( ~n3156 & n3293 ) | ( n3269 & n3293 ) ;
  assign n3329 = ( n3156 & ~n3293 ) | ( n3156 & n3328 ) | ( ~n3293 & n3328 ) ;
  assign n3330 = ( ~n3269 & n3328 ) | ( ~n3269 & n3329 ) | ( n3328 & n3329 ) ;
  assign n3331 = ( ~n2886 & n3002 ) | ( ~n2886 & n3026 ) | ( n3002 & n3026 ) ;
  assign n3332 = ( n2886 & ~n3026 ) | ( n2886 & n3331 ) | ( ~n3026 & n3331 ) ;
  assign n3333 = ( ~n3002 & n3331 ) | ( ~n3002 & n3332 ) | ( n3331 & n3332 ) ;
  assign n3334 = ( n3327 & n3330 ) | ( n3327 & n3333 ) | ( n3330 & n3333 ) ;
  assign n3335 = n3306 & n3334 ;
  assign n3336 = n3039 & n3305 ;
  assign n3337 = ( n3029 & n3031 ) | ( n3029 & n3034 ) | ( n3031 & n3034 ) ;
  assign n3338 = ( n3032 & n3037 ) | ( n3032 & n3337 ) | ( n3037 & n3337 ) ;
  assign n3339 = ( n3296 & n3298 ) | ( n3296 & n3302 ) | ( n3298 & n3302 ) ;
  assign n3340 = n3299 | n3339 ;
  assign n3341 = n3338 & n3340 ;
  assign n3342 = n3340 & ~n3341 ;
  assign n3343 = ( n3338 & ~n3341 ) | ( n3338 & n3342 ) | ( ~n3341 & n3342 ) ;
  assign n3344 = n3336 | n3343 ;
  assign n3345 = n3335 | n3344 ;
  assign n3346 = n3335 | n3336 ;
  assign n3347 = n3343 & n3346 ;
  assign n3348 = n3345 & ~n3347 ;
  assign n3349 = ( ~n2734 & n2737 ) | ( ~n2734 & n2765 ) | ( n2737 & n2765 ) ;
  assign n3350 = ( n2734 & ~n2765 ) | ( n2734 & n3349 ) | ( ~n2765 & n3349 ) ;
  assign n3351 = ( ~n2737 & n3349 ) | ( ~n2737 & n3350 ) | ( n3349 & n3350 ) ;
  assign n3352 = ( ~n3039 & n3305 ) | ( ~n3039 & n3334 ) | ( n3305 & n3334 ) ;
  assign n3353 = ( n3039 & ~n3334 ) | ( n3039 & n3352 ) | ( ~n3334 & n3352 ) ;
  assign n3354 = ( ~n3305 & n3352 ) | ( ~n3305 & n3353 ) | ( n3352 & n3353 ) ;
  assign n3355 = ( ~n2740 & n2743 ) | ( ~n2740 & n2757 ) | ( n2743 & n2757 ) ;
  assign n3356 = ( n2740 & ~n2757 ) | ( n2740 & n3355 ) | ( ~n2757 & n3355 ) ;
  assign n3357 = ( ~n2743 & n3355 ) | ( ~n2743 & n3356 ) | ( n3355 & n3356 ) ;
  assign n3358 = ( ~n3309 & n3312 ) | ( ~n3309 & n3326 ) | ( n3312 & n3326 ) ;
  assign n3359 = ( n3309 & ~n3326 ) | ( n3309 & n3358 ) | ( ~n3326 & n3358 ) ;
  assign n3360 = ( ~n3312 & n3358 ) | ( ~n3312 & n3359 ) | ( n3358 & n3359 ) ;
  assign n3361 = n3315 & ~n3318 ;
  assign n3362 = ~n3315 & n3318 ;
  assign n3363 = n3361 | n3362 ;
  assign n3364 = n2746 & ~n2749 ;
  assign n3365 = ~n2746 & n2749 ;
  assign n3366 = n3364 | n3365 ;
  assign n3367 = n3363 & n3366 ;
  assign n3368 = ~n3319 & n3322 ;
  assign n3369 = n3319 & ~n3322 ;
  assign n3370 = n3368 | n3369 ;
  assign n3371 = n3325 & ~n3370 ;
  assign n3372 = ~n3325 & n3370 ;
  assign n3373 = n3371 | n3372 ;
  assign n3374 = ( n2750 & n2756 ) | ( n2750 & ~n2757 ) | ( n2756 & ~n2757 ) ;
  assign n3375 = ( n2753 & ~n2757 ) | ( n2753 & n3374 ) | ( ~n2757 & n3374 ) ;
  assign n3376 = ( n3367 & n3373 ) | ( n3367 & n3375 ) | ( n3373 & n3375 ) ;
  assign n3377 = ( n3357 & n3360 ) | ( n3357 & n3376 ) | ( n3360 & n3376 ) ;
  assign n3378 = ( n3327 & ~n3330 ) | ( n3327 & n3333 ) | ( ~n3330 & n3333 ) ;
  assign n3379 = ( ~n3327 & n3330 ) | ( ~n3327 & n3378 ) | ( n3330 & n3378 ) ;
  assign n3380 = ( ~n3333 & n3378 ) | ( ~n3333 & n3379 ) | ( n3378 & n3379 ) ;
  assign n3381 = ( n2758 & ~n2761 ) | ( n2758 & n2764 ) | ( ~n2761 & n2764 ) ;
  assign n3382 = ( ~n2758 & n2761 ) | ( ~n2758 & n3381 ) | ( n2761 & n3381 ) ;
  assign n3383 = ( ~n2764 & n3381 ) | ( ~n2764 & n3382 ) | ( n3381 & n3382 ) ;
  assign n3384 = ( n3377 & n3380 ) | ( n3377 & n3383 ) | ( n3380 & n3383 ) ;
  assign n3385 = ( n3351 & n3354 ) | ( n3351 & n3384 ) | ( n3354 & n3384 ) ;
  assign n3386 = ( n2769 & ~n3348 ) | ( n2769 & n3385 ) | ( ~n3348 & n3385 ) ;
  assign n3387 = ( n3348 & ~n3385 ) | ( n3348 & n3386 ) | ( ~n3385 & n3386 ) ;
  assign n3388 = ( ~n2769 & n3386 ) | ( ~n2769 & n3387 ) | ( n3386 & n3387 ) ;
  assign n3389 = ( n3351 & ~n3354 ) | ( n3351 & n3384 ) | ( ~n3354 & n3384 ) ;
  assign n3390 = ( ~n3351 & n3354 ) | ( ~n3351 & n3389 ) | ( n3354 & n3389 ) ;
  assign n3391 = ( ~n3384 & n3389 ) | ( ~n3384 & n3390 ) | ( n3389 & n3390 ) ;
  assign n3392 = ( n2153 & ~n2156 ) | ( n2153 & n2186 ) | ( ~n2156 & n2186 ) ;
  assign n3393 = ( ~n2153 & n2156 ) | ( ~n2153 & n3392 ) | ( n2156 & n3392 ) ;
  assign n3394 = ( ~n2186 & n3392 ) | ( ~n2186 & n3393 ) | ( n3392 & n3393 ) ;
  assign n3395 = ( ~n3357 & n3360 ) | ( ~n3357 & n3376 ) | ( n3360 & n3376 ) ;
  assign n3396 = ( n3357 & ~n3376 ) | ( n3357 & n3395 ) | ( ~n3376 & n3395 ) ;
  assign n3397 = ( ~n3360 & n3395 ) | ( ~n3360 & n3396 ) | ( n3395 & n3396 ) ;
  assign n3398 = ( ~n2159 & n2162 ) | ( ~n2159 & n2178 ) | ( n2162 & n2178 ) ;
  assign n3399 = ( n2159 & ~n2178 ) | ( n2159 & n3398 ) | ( ~n2178 & n3398 ) ;
  assign n3400 = ( ~n2162 & n3398 ) | ( ~n2162 & n3399 ) | ( n3398 & n3399 ) ;
  assign n3401 = n2165 & ~n2168 ;
  assign n3402 = ~n2165 & n2168 ;
  assign n3403 = n3401 | n3402 ;
  assign n3404 = n3363 & ~n3366 ;
  assign n3405 = ~n3363 & n3366 ;
  assign n3406 = n3404 | n3405 ;
  assign n3407 = n3403 & n3406 ;
  assign n3408 = ( n2169 & ~n2175 ) | ( n2169 & n2177 ) | ( ~n2175 & n2177 ) ;
  assign n3409 = ( ~n2169 & n2175 ) | ( ~n2169 & n3408 ) | ( n2175 & n3408 ) ;
  assign n3410 = ( ~n2177 & n3408 ) | ( ~n2177 & n3409 ) | ( n3408 & n3409 ) ;
  assign n3411 = ( n3367 & ~n3373 ) | ( n3367 & n3375 ) | ( ~n3373 & n3375 ) ;
  assign n3412 = ( ~n3367 & n3373 ) | ( ~n3367 & n3411 ) | ( n3373 & n3411 ) ;
  assign n3413 = ( ~n3375 & n3411 ) | ( ~n3375 & n3412 ) | ( n3411 & n3412 ) ;
  assign n3414 = ( n3407 & n3410 ) | ( n3407 & n3413 ) | ( n3410 & n3413 ) ;
  assign n3415 = ( n3397 & n3400 ) | ( n3397 & n3414 ) | ( n3400 & n3414 ) ;
  assign n3416 = ( n2179 & ~n2182 ) | ( n2179 & n2185 ) | ( ~n2182 & n2185 ) ;
  assign n3417 = ( ~n2179 & n2182 ) | ( ~n2179 & n3416 ) | ( n2182 & n3416 ) ;
  assign n3418 = ( ~n2185 & n3416 ) | ( ~n2185 & n3417 ) | ( n3416 & n3417 ) ;
  assign n3419 = ( n3377 & ~n3380 ) | ( n3377 & n3383 ) | ( ~n3380 & n3383 ) ;
  assign n3420 = ( ~n3377 & n3380 ) | ( ~n3377 & n3419 ) | ( n3380 & n3419 ) ;
  assign n3421 = ( ~n3383 & n3419 ) | ( ~n3383 & n3420 ) | ( n3419 & n3420 ) ;
  assign n3422 = ( n3415 & n3418 ) | ( n3415 & n3421 ) | ( n3418 & n3421 ) ;
  assign n3423 = ( n3391 & n3394 ) | ( n3391 & n3422 ) | ( n3394 & n3422 ) ;
  assign n3424 = ( n2190 & n3388 ) | ( n2190 & n3423 ) | ( n3388 & n3423 ) ;
  assign n3425 = n2769 | n3348 ;
  assign n3426 = n3385 & n3425 ;
  assign n3427 = n2769 & n3348 ;
  assign n3428 = n2460 & n2730 ;
  assign n3429 = n2456 | n2685 ;
  assign n3430 = n2459 | n3429 ;
  assign n3431 = ( n2452 & n3429 ) | ( n2452 & n3430 ) | ( n3429 & n3430 ) ;
  assign n3432 = n2729 | n3431 ;
  assign n3433 = ( n2766 & n3428 ) | ( n2766 & n3432 ) | ( n3428 & n3432 ) ;
  assign n3434 = n3032 | n3299 ;
  assign n3435 = n3337 | n3434 ;
  assign n3436 = ( n3037 & n3434 ) | ( n3037 & n3435 ) | ( n3434 & n3435 ) ;
  assign n3437 = n3339 | n3436 ;
  assign n3438 = n3346 & n3437 ;
  assign n3439 = n3341 | n3438 ;
  assign n3440 = n3433 & n3439 ;
  assign n3441 = n3439 & ~n3440 ;
  assign n3442 = ( n3433 & ~n3440 ) | ( n3433 & n3441 ) | ( ~n3440 & n3441 ) ;
  assign n3443 = n3427 | n3442 ;
  assign n3444 = n3426 | n3443 ;
  assign n3445 = n3426 | n3427 ;
  assign n3446 = n3442 & n3445 ;
  assign n3447 = n3444 & ~n3446 ;
  assign n3448 = n1271 & n1536 ;
  assign n3449 = n1230 | n1491 ;
  assign n3450 = n1270 | n3449 ;
  assign n3451 = ( n1267 & n3449 ) | ( n1267 & n3450 ) | ( n3449 & n3450 ) ;
  assign n3452 = n1535 | n3451 ;
  assign n3453 = ( n1572 & n3448 ) | ( n1572 & n3452 ) | ( n3448 & n3452 ) ;
  assign n3454 = n1801 | n2101 ;
  assign n3455 = n2139 | n3454 ;
  assign n3456 = ( n1837 & n3454 ) | ( n1837 & n3455 ) | ( n3454 & n3455 ) ;
  assign n3457 = n2141 | n3456 ;
  assign n3458 = n2148 & n3457 ;
  assign n3459 = n2143 | n3458 ;
  assign n3460 = ( n1575 & n2150 ) | ( n1575 & n2187 ) | ( n2150 & n2187 ) ;
  assign n3461 = ( n3453 & n3459 ) | ( n3453 & ~n3460 ) | ( n3459 & ~n3460 ) ;
  assign n3462 = ( ~n3459 & n3460 ) | ( ~n3459 & n3461 ) | ( n3460 & n3461 ) ;
  assign n3463 = ( ~n3453 & n3461 ) | ( ~n3453 & n3462 ) | ( n3461 & n3462 ) ;
  assign n3464 = n3447 | n3463 ;
  assign n3465 = n3424 & n3464 ;
  assign n3466 = n3447 & n3463 ;
  assign n3467 = n3465 | n3466 ;
  assign n3468 = n2143 | n3448 ;
  assign n3469 = n3452 | n3468 ;
  assign n3470 = ( n1572 & n3468 ) | ( n1572 & n3469 ) | ( n3468 & n3469 ) ;
  assign n3471 = n3458 | n3470 ;
  assign n3472 = n3460 & n3471 ;
  assign n3473 = n3453 & n3459 ;
  assign n3474 = n3440 | n3473 ;
  assign n3475 = n3341 | n3428 ;
  assign n3476 = n3432 | n3475 ;
  assign n3477 = ( n2766 & n3475 ) | ( n2766 & n3476 ) | ( n3475 & n3476 ) ;
  assign n3478 = n3438 | n3477 ;
  assign n3479 = n3474 | n3478 ;
  assign n3480 = ( n3445 & n3474 ) | ( n3445 & n3479 ) | ( n3474 & n3479 ) ;
  assign n3481 = n3472 | n3480 ;
  assign n3482 = n3467 & n3481 ;
  assign n3483 = ( n3440 & n3445 ) | ( n3440 & n3478 ) | ( n3445 & n3478 ) ;
  assign n3484 = n3472 | n3473 ;
  assign n3485 = n3483 & n3484 ;
  assign n3486 = ( x19 & ~x20 ) | ( x19 & x21 ) | ( ~x20 & x21 ) ;
  assign n3487 = ( ~x19 & x20 ) | ( ~x19 & n3486 ) | ( x20 & n3486 ) ;
  assign n3488 = ( ~x21 & n3486 ) | ( ~x21 & n3487 ) | ( n3486 & n3487 ) ;
  assign n3489 = ( x22 & ~x23 ) | ( x22 & x24 ) | ( ~x23 & x24 ) ;
  assign n3490 = ( ~x22 & x23 ) | ( ~x22 & n3489 ) | ( x23 & n3489 ) ;
  assign n3491 = ( ~x24 & n3489 ) | ( ~x24 & n3490 ) | ( n3489 & n3490 ) ;
  assign n3492 = n3488 & n3491 ;
  assign n3493 = ( x22 & x23 ) | ( x22 & x24 ) | ( x23 & x24 ) ;
  assign n3494 = ( x19 & x20 ) | ( x19 & x21 ) | ( x20 & x21 ) ;
  assign n3495 = ( n3492 & n3493 ) | ( n3492 & n3494 ) | ( n3493 & n3494 ) ;
  assign n3496 = ( x28 & x29 ) | ( x28 & x30 ) | ( x29 & x30 ) ;
  assign n3497 = ( x25 & x26 ) | ( x25 & x27 ) | ( x26 & x27 ) ;
  assign n3498 = ( x25 & ~x26 ) | ( x25 & x27 ) | ( ~x26 & x27 ) ;
  assign n3499 = ( ~x25 & x26 ) | ( ~x25 & n3498 ) | ( x26 & n3498 ) ;
  assign n3500 = ( ~x27 & n3498 ) | ( ~x27 & n3499 ) | ( n3498 & n3499 ) ;
  assign n3501 = ( x28 & ~x29 ) | ( x28 & x30 ) | ( ~x29 & x30 ) ;
  assign n3502 = ( ~x28 & x29 ) | ( ~x28 & n3501 ) | ( x29 & n3501 ) ;
  assign n3503 = ( ~x30 & n3501 ) | ( ~x30 & n3502 ) | ( n3501 & n3502 ) ;
  assign n3504 = n3500 & n3503 ;
  assign n3505 = ( n3496 & n3497 ) | ( n3496 & n3504 ) | ( n3497 & n3504 ) ;
  assign n3506 = ( n3492 & n3494 ) | ( n3492 & ~n3495 ) | ( n3494 & ~n3495 ) ;
  assign n3507 = ( n3493 & ~n3495 ) | ( n3493 & n3506 ) | ( ~n3495 & n3506 ) ;
  assign n3508 = ( n3497 & n3504 ) | ( n3497 & ~n3505 ) | ( n3504 & ~n3505 ) ;
  assign n3509 = ( n3496 & ~n3505 ) | ( n3496 & n3508 ) | ( ~n3505 & n3508 ) ;
  assign n3510 = n3495 & n3507 ;
  assign n3511 = n3488 & ~n3491 ;
  assign n3512 = ~n3488 & n3491 ;
  assign n3513 = n3511 | n3512 ;
  assign n3514 = n3500 & ~n3503 ;
  assign n3515 = ~n3500 & n3503 ;
  assign n3516 = n3514 | n3515 ;
  assign n3517 = n3513 & n3516 ;
  assign n3518 = ~n3510 & n3517 ;
  assign n3519 = ( n3507 & n3509 ) | ( n3507 & n3518 ) | ( n3509 & n3518 ) ;
  assign n3520 = ( n3495 & n3505 ) | ( n3495 & n3519 ) | ( n3505 & n3519 ) ;
  assign n3521 = ( x7 & ~x8 ) | ( x7 & x9 ) | ( ~x8 & x9 ) ;
  assign n3522 = ( ~x7 & x8 ) | ( ~x7 & n3521 ) | ( x8 & n3521 ) ;
  assign n3523 = ( ~x9 & n3521 ) | ( ~x9 & n3522 ) | ( n3521 & n3522 ) ;
  assign n3524 = ( x10 & ~x11 ) | ( x10 & x12 ) | ( ~x11 & x12 ) ;
  assign n3525 = ( ~x10 & x11 ) | ( ~x10 & n3524 ) | ( x11 & n3524 ) ;
  assign n3526 = ( ~x12 & n3524 ) | ( ~x12 & n3525 ) | ( n3524 & n3525 ) ;
  assign n3527 = n3523 & n3526 ;
  assign n3528 = ( x10 & x11 ) | ( x10 & x12 ) | ( x11 & x12 ) ;
  assign n3529 = ( x7 & x8 ) | ( x7 & x9 ) | ( x8 & x9 ) ;
  assign n3530 = ( n3527 & n3528 ) | ( n3527 & n3529 ) | ( n3528 & n3529 ) ;
  assign n3531 = ( x16 & x17 ) | ( x16 & x18 ) | ( x17 & x18 ) ;
  assign n3532 = ( x13 & x14 ) | ( x13 & x15 ) | ( x14 & x15 ) ;
  assign n3533 = ( x13 & ~x14 ) | ( x13 & x15 ) | ( ~x14 & x15 ) ;
  assign n3534 = ( ~x13 & x14 ) | ( ~x13 & n3533 ) | ( x14 & n3533 ) ;
  assign n3535 = ( ~x15 & n3533 ) | ( ~x15 & n3534 ) | ( n3533 & n3534 ) ;
  assign n3536 = ( x16 & ~x17 ) | ( x16 & x18 ) | ( ~x17 & x18 ) ;
  assign n3537 = ( ~x16 & x17 ) | ( ~x16 & n3536 ) | ( x17 & n3536 ) ;
  assign n3538 = ( ~x18 & n3536 ) | ( ~x18 & n3537 ) | ( n3536 & n3537 ) ;
  assign n3539 = n3535 & n3538 ;
  assign n3540 = ( n3531 & n3532 ) | ( n3531 & n3539 ) | ( n3532 & n3539 ) ;
  assign n3541 = ( n3527 & n3529 ) | ( n3527 & ~n3530 ) | ( n3529 & ~n3530 ) ;
  assign n3542 = ( n3528 & ~n3530 ) | ( n3528 & n3541 ) | ( ~n3530 & n3541 ) ;
  assign n3543 = n3530 & n3542 ;
  assign n3544 = ( n3532 & n3539 ) | ( n3532 & ~n3540 ) | ( n3539 & ~n3540 ) ;
  assign n3545 = ( n3531 & ~n3540 ) | ( n3531 & n3544 ) | ( ~n3540 & n3544 ) ;
  assign n3546 = n3540 & n3545 ;
  assign n3547 = n3523 & ~n3526 ;
  assign n3548 = ~n3523 & n3526 ;
  assign n3549 = n3547 | n3548 ;
  assign n3550 = n3535 & ~n3538 ;
  assign n3551 = ~n3535 & n3538 ;
  assign n3552 = n3550 | n3551 ;
  assign n3553 = n3549 & n3552 ;
  assign n3554 = ~n3546 & n3553 ;
  assign n3555 = n3545 & n3554 ;
  assign n3556 = ~n3543 & n3555 ;
  assign n3557 = ~n3543 & n3554 ;
  assign n3558 = ~n3545 & n3557 ;
  assign n3559 = ( n3542 & n3545 ) | ( n3542 & n3558 ) | ( n3545 & n3558 ) ;
  assign n3560 = n3556 | n3559 ;
  assign n3561 = ( n3530 & n3540 ) | ( n3530 & n3560 ) | ( n3540 & n3560 ) ;
  assign n3562 = ~n3530 & n3540 ;
  assign n3563 = n3530 & ~n3540 ;
  assign n3564 = n3562 | n3563 ;
  assign n3565 = n3556 | n3564 ;
  assign n3566 = n3559 | n3565 ;
  assign n3567 = n3560 & n3564 ;
  assign n3568 = n3566 & ~n3567 ;
  assign n3569 = ( n3495 & n3505 ) | ( n3495 & ~n3519 ) | ( n3505 & ~n3519 ) ;
  assign n3570 = ( ~n3495 & n3505 ) | ( ~n3495 & n3519 ) | ( n3505 & n3519 ) ;
  assign n3571 = ( ~n3505 & n3569 ) | ( ~n3505 & n3570 ) | ( n3569 & n3570 ) ;
  assign n3572 = ( n3542 & n3545 ) | ( n3542 & ~n3557 ) | ( n3545 & ~n3557 ) ;
  assign n3573 = n3542 & ~n3556 ;
  assign n3574 = ( n3545 & ~n3572 ) | ( n3545 & n3573 ) | ( ~n3572 & n3573 ) ;
  assign n3575 = ( n3558 & n3572 ) | ( n3558 & ~n3574 ) | ( n3572 & ~n3574 ) ;
  assign n3576 = n3513 & ~n3516 ;
  assign n3577 = ~n3513 & n3516 ;
  assign n3578 = n3576 | n3577 ;
  assign n3579 = n3549 & ~n3552 ;
  assign n3580 = ~n3549 & n3552 ;
  assign n3581 = n3579 | n3580 ;
  assign n3582 = n3578 & n3581 ;
  assign n3583 = n3509 | n3518 ;
  assign n3584 = ~n3519 & n3583 ;
  assign n3585 = n3509 & n3517 ;
  assign n3586 = ( n3507 & ~n3583 ) | ( n3507 & n3585 ) | ( ~n3583 & n3585 ) ;
  assign n3587 = n3584 | n3586 ;
  assign n3588 = n3582 | n3587 ;
  assign n3589 = ( n3582 & n3584 ) | ( n3582 & n3586 ) | ( n3584 & n3586 ) ;
  assign n3590 = ( n3575 & n3588 ) | ( n3575 & n3589 ) | ( n3588 & n3589 ) ;
  assign n3591 = ( n3568 & n3571 ) | ( n3568 & n3590 ) | ( n3571 & n3590 ) ;
  assign n3592 = ( n3520 & n3561 ) | ( n3520 & n3591 ) | ( n3561 & n3591 ) ;
  assign n3593 = ( x994 & x995 ) | ( x994 & x996 ) | ( x995 & x996 ) ;
  assign n3594 = ( x991 & x992 ) | ( x991 & x993 ) | ( x992 & x993 ) ;
  assign n3595 = ( x991 & ~x992 ) | ( x991 & x993 ) | ( ~x992 & x993 ) ;
  assign n3596 = ( ~x991 & x992 ) | ( ~x991 & n3595 ) | ( x992 & n3595 ) ;
  assign n3597 = ( ~x993 & n3595 ) | ( ~x993 & n3596 ) | ( n3595 & n3596 ) ;
  assign n3598 = ( x994 & ~x995 ) | ( x994 & x996 ) | ( ~x995 & x996 ) ;
  assign n3599 = ( ~x994 & x995 ) | ( ~x994 & n3598 ) | ( x995 & n3598 ) ;
  assign n3600 = ( ~x996 & n3598 ) | ( ~x996 & n3599 ) | ( n3598 & n3599 ) ;
  assign n3601 = n3597 & n3600 ;
  assign n3602 = ( n3593 & n3594 ) | ( n3593 & n3601 ) | ( n3594 & n3601 ) ;
  assign n3603 = x0 & ~x1 ;
  assign n3604 = ~x0 & x1 ;
  assign n3605 = x2 & ~n3604 ;
  assign n3606 = ~n3603 & n3605 ;
  assign n3607 = ( ~x2 & n3603 ) | ( ~x2 & n3604 ) | ( n3603 & n3604 ) ;
  assign n3608 = n3606 | n3607 ;
  assign n3609 = x6 & n3608 ;
  assign n3610 = ( x0 & x1 ) | ( x0 & x2 ) | ( x1 & x2 ) ;
  assign n3611 = ( x3 & x4 ) | ( x3 & x5 ) | ( x4 & x5 ) ;
  assign n3612 = n3610 & n3611 ;
  assign n3613 = n3611 & ~n3612 ;
  assign n3614 = ( n3610 & ~n3612 ) | ( n3610 & n3613 ) | ( ~n3612 & n3613 ) ;
  assign n3615 = n3609 | n3614 ;
  assign n3616 = ~x6 & n3608 ;
  assign n3617 = ( x3 & ~x4 ) | ( x3 & x5 ) | ( ~x4 & x5 ) ;
  assign n3618 = ( ~x3 & x4 ) | ( ~x3 & n3617 ) | ( x4 & n3617 ) ;
  assign n3619 = ( ~x5 & n3617 ) | ( ~x5 & n3618 ) | ( n3617 & n3618 ) ;
  assign n3620 = x6 & ~n3608 ;
  assign n3621 = ( n3616 & n3619 ) | ( n3616 & n3620 ) | ( n3619 & n3620 ) ;
  assign n3622 = n3615 | n3621 ;
  assign n3623 = ( n3609 & n3614 ) | ( n3609 & n3621 ) | ( n3614 & n3621 ) ;
  assign n3624 = n3622 & ~n3623 ;
  assign n3625 = ( n3616 & n3619 ) | ( n3616 & ~n3620 ) | ( n3619 & ~n3620 ) ;
  assign n3626 = ( n3620 & ~n3621 ) | ( n3620 & n3625 ) | ( ~n3621 & n3625 ) ;
  assign n3627 = ( x997 & ~x998 ) | ( x997 & x999 ) | ( ~x998 & x999 ) ;
  assign n3628 = ( ~x997 & x998 ) | ( ~x997 & n3627 ) | ( x998 & n3627 ) ;
  assign n3629 = ( ~x999 & n3627 ) | ( ~x999 & n3628 ) | ( n3627 & n3628 ) ;
  assign n3630 = n3626 & n3629 ;
  assign n3631 = n3624 | n3630 ;
  assign n3632 = ( x997 & x998 ) | ( x997 & x999 ) | ( x998 & x999 ) ;
  assign n3633 = n3631 & n3632 ;
  assign n3634 = n3612 | n3623 ;
  assign n3635 = n3624 & n3630 ;
  assign n3636 = ~n3634 & n3635 ;
  assign n3637 = ( n3633 & ~n3634 ) | ( n3633 & n3636 ) | ( ~n3634 & n3636 ) ;
  assign n3638 = n3631 & ~n3635 ;
  assign n3639 = n3632 & ~n3638 ;
  assign n3640 = ( ~n3632 & n3638 ) | ( ~n3632 & n3639 ) | ( n3638 & n3639 ) ;
  assign n3641 = ( ~n3631 & n3634 ) | ( ~n3631 & n3640 ) | ( n3634 & n3640 ) ;
  assign n3642 = n3637 | n3641 ;
  assign n3643 = n3602 & n3642 ;
  assign n3644 = ( n3594 & n3601 ) | ( n3594 & ~n3602 ) | ( n3601 & ~n3602 ) ;
  assign n3645 = ( n3593 & ~n3602 ) | ( n3593 & n3644 ) | ( ~n3602 & n3644 ) ;
  assign n3646 = n3597 & ~n3600 ;
  assign n3647 = ~n3597 & n3600 ;
  assign n3648 = n3646 | n3647 ;
  assign n3649 = n3626 | n3629 ;
  assign n3650 = ~n3629 & n3649 ;
  assign n3651 = ( ~n3626 & n3649 ) | ( ~n3626 & n3650 ) | ( n3649 & n3650 ) ;
  assign n3652 = n3648 & n3651 ;
  assign n3653 = n3639 | n3640 ;
  assign n3654 = ( n3645 & n3652 ) | ( n3645 & n3653 ) | ( n3652 & n3653 ) ;
  assign n3655 = ( n3602 & n3643 ) | ( n3602 & n3654 ) | ( n3643 & n3654 ) ;
  assign n3656 = ( n3633 & n3634 ) | ( n3633 & ~n3642 ) | ( n3634 & ~n3642 ) ;
  assign n3657 = n3655 & n3656 ;
  assign n3658 = n3592 & n3657 ;
  assign n3659 = n3655 | n3656 ;
  assign n3660 = ~n3602 & n3642 ;
  assign n3661 = ( n3642 & n3654 ) | ( n3642 & n3660 ) | ( n3654 & n3660 ) ;
  assign n3662 = n3659 | n3661 ;
  assign n3663 = ~n3657 & n3662 ;
  assign n3664 = ( ~n3642 & n3654 ) | ( ~n3642 & n3660 ) | ( n3654 & n3660 ) ;
  assign n3665 = ( n3642 & ~n3661 ) | ( n3642 & n3664 ) | ( ~n3661 & n3664 ) ;
  assign n3666 = ( n3568 & ~n3571 ) | ( n3568 & n3590 ) | ( ~n3571 & n3590 ) ;
  assign n3667 = ( ~n3568 & n3571 ) | ( ~n3568 & n3666 ) | ( n3571 & n3666 ) ;
  assign n3668 = ( ~n3590 & n3666 ) | ( ~n3590 & n3667 ) | ( n3666 & n3667 ) ;
  assign n3669 = n3578 & ~n3581 ;
  assign n3670 = ~n3578 & n3581 ;
  assign n3671 = n3669 | n3670 ;
  assign n3672 = n3648 & ~n3652 ;
  assign n3673 = ( n3651 & ~n3652 ) | ( n3651 & n3672 ) | ( ~n3652 & n3672 ) ;
  assign n3674 = n3671 & n3673 ;
  assign n3675 = ~n3582 & n3588 ;
  assign n3676 = ( ~n3587 & n3588 ) | ( ~n3587 & n3675 ) | ( n3588 & n3675 ) ;
  assign n3677 = n3575 & ~n3676 ;
  assign n3678 = ~n3575 & n3676 ;
  assign n3679 = n3677 | n3678 ;
  assign n3680 = ( n3645 & n3652 ) | ( n3645 & ~n3654 ) | ( n3652 & ~n3654 ) ;
  assign n3681 = ( n3653 & ~n3654 ) | ( n3653 & n3680 ) | ( ~n3654 & n3680 ) ;
  assign n3682 = ( n3674 & n3679 ) | ( n3674 & n3681 ) | ( n3679 & n3681 ) ;
  assign n3683 = ( n3665 & n3668 ) | ( n3665 & n3682 ) | ( n3668 & n3682 ) ;
  assign n3684 = ( n3520 & n3561 ) | ( n3520 & ~n3591 ) | ( n3561 & ~n3591 ) ;
  assign n3685 = ( ~n3561 & n3591 ) | ( ~n3561 & n3684 ) | ( n3591 & n3684 ) ;
  assign n3686 = ( ~n3520 & n3684 ) | ( ~n3520 & n3685 ) | ( n3684 & n3685 ) ;
  assign n3687 = ( n3663 & n3683 ) | ( n3663 & n3686 ) | ( n3683 & n3686 ) ;
  assign n3688 = n3592 | n3657 ;
  assign n3689 = ( n3658 & n3687 ) | ( n3658 & n3688 ) | ( n3687 & n3688 ) ;
  assign n3690 = ( x52 & x53 ) | ( x52 & x54 ) | ( x53 & x54 ) ;
  assign n3691 = ( x49 & x50 ) | ( x49 & x51 ) | ( x50 & x51 ) ;
  assign n3692 = ( x49 & ~x50 ) | ( x49 & x51 ) | ( ~x50 & x51 ) ;
  assign n3693 = ( ~x49 & x50 ) | ( ~x49 & n3692 ) | ( x50 & n3692 ) ;
  assign n3694 = ( ~x51 & n3692 ) | ( ~x51 & n3693 ) | ( n3692 & n3693 ) ;
  assign n3695 = ( x52 & ~x53 ) | ( x52 & x54 ) | ( ~x53 & x54 ) ;
  assign n3696 = ( ~x52 & x53 ) | ( ~x52 & n3695 ) | ( x53 & n3695 ) ;
  assign n3697 = ( ~x54 & n3695 ) | ( ~x54 & n3696 ) | ( n3695 & n3696 ) ;
  assign n3698 = n3694 & n3697 ;
  assign n3699 = ( n3690 & n3691 ) | ( n3690 & n3698 ) | ( n3691 & n3698 ) ;
  assign n3700 = ( x43 & ~x44 ) | ( x43 & x45 ) | ( ~x44 & x45 ) ;
  assign n3701 = ( ~x43 & x44 ) | ( ~x43 & n3700 ) | ( x44 & n3700 ) ;
  assign n3702 = ( ~x45 & n3700 ) | ( ~x45 & n3701 ) | ( n3700 & n3701 ) ;
  assign n3703 = ( x46 & ~x47 ) | ( x46 & x48 ) | ( ~x47 & x48 ) ;
  assign n3704 = ( ~x46 & x47 ) | ( ~x46 & n3703 ) | ( x47 & n3703 ) ;
  assign n3705 = ( ~x48 & n3703 ) | ( ~x48 & n3704 ) | ( n3703 & n3704 ) ;
  assign n3706 = n3702 & n3705 ;
  assign n3707 = ( x46 & x47 ) | ( x46 & x48 ) | ( x47 & x48 ) ;
  assign n3708 = ( x43 & x44 ) | ( x43 & x45 ) | ( x44 & x45 ) ;
  assign n3709 = ( n3706 & n3707 ) | ( n3706 & n3708 ) | ( n3707 & n3708 ) ;
  assign n3710 = ( n3691 & n3698 ) | ( n3691 & ~n3699 ) | ( n3698 & ~n3699 ) ;
  assign n3711 = ( n3690 & ~n3699 ) | ( n3690 & n3710 ) | ( ~n3699 & n3710 ) ;
  assign n3712 = ( n3706 & n3708 ) | ( n3706 & ~n3709 ) | ( n3708 & ~n3709 ) ;
  assign n3713 = ( n3707 & ~n3709 ) | ( n3707 & n3712 ) | ( ~n3709 & n3712 ) ;
  assign n3714 = n3709 & n3713 ;
  assign n3715 = n3694 & ~n3697 ;
  assign n3716 = ~n3694 & n3697 ;
  assign n3717 = n3715 | n3716 ;
  assign n3718 = n3702 & ~n3705 ;
  assign n3719 = ~n3702 & n3705 ;
  assign n3720 = n3718 | n3719 ;
  assign n3721 = n3717 & n3720 ;
  assign n3722 = ~n3714 & n3721 ;
  assign n3723 = ( n3711 & n3713 ) | ( n3711 & n3722 ) | ( n3713 & n3722 ) ;
  assign n3724 = ( n3699 & n3709 ) | ( n3699 & n3723 ) | ( n3709 & n3723 ) ;
  assign n3725 = ( x40 & x41 ) | ( x40 & x42 ) | ( x41 & x42 ) ;
  assign n3726 = ( x37 & x38 ) | ( x37 & x39 ) | ( x38 & x39 ) ;
  assign n3727 = ( x37 & ~x38 ) | ( x37 & x39 ) | ( ~x38 & x39 ) ;
  assign n3728 = ( ~x37 & x38 ) | ( ~x37 & n3727 ) | ( x38 & n3727 ) ;
  assign n3729 = ( ~x39 & n3727 ) | ( ~x39 & n3728 ) | ( n3727 & n3728 ) ;
  assign n3730 = ( x40 & ~x41 ) | ( x40 & x42 ) | ( ~x41 & x42 ) ;
  assign n3731 = ( ~x40 & x41 ) | ( ~x40 & n3730 ) | ( x41 & n3730 ) ;
  assign n3732 = ( ~x42 & n3730 ) | ( ~x42 & n3731 ) | ( n3730 & n3731 ) ;
  assign n3733 = n3729 & n3732 ;
  assign n3734 = ( n3725 & n3726 ) | ( n3725 & n3733 ) | ( n3726 & n3733 ) ;
  assign n3735 = ( x34 & x35 ) | ( x34 & x36 ) | ( x35 & x36 ) ;
  assign n3736 = ( x31 & x32 ) | ( x31 & x33 ) | ( x32 & x33 ) ;
  assign n3737 = ( x31 & ~x32 ) | ( x31 & x33 ) | ( ~x32 & x33 ) ;
  assign n3738 = ( ~x31 & x32 ) | ( ~x31 & n3737 ) | ( x32 & n3737 ) ;
  assign n3739 = ( ~x33 & n3737 ) | ( ~x33 & n3738 ) | ( n3737 & n3738 ) ;
  assign n3740 = ( x34 & ~x35 ) | ( x34 & x36 ) | ( ~x35 & x36 ) ;
  assign n3741 = ( ~x34 & x35 ) | ( ~x34 & n3740 ) | ( x35 & n3740 ) ;
  assign n3742 = ( ~x36 & n3740 ) | ( ~x36 & n3741 ) | ( n3740 & n3741 ) ;
  assign n3743 = n3739 & n3742 ;
  assign n3744 = ( n3735 & n3736 ) | ( n3735 & n3743 ) | ( n3736 & n3743 ) ;
  assign n3745 = ( n3736 & n3743 ) | ( n3736 & ~n3744 ) | ( n3743 & ~n3744 ) ;
  assign n3746 = ( n3735 & ~n3744 ) | ( n3735 & n3745 ) | ( ~n3744 & n3745 ) ;
  assign n3747 = n3744 & n3746 ;
  assign n3748 = ( n3726 & n3733 ) | ( n3726 & ~n3734 ) | ( n3733 & ~n3734 ) ;
  assign n3749 = ( n3725 & ~n3734 ) | ( n3725 & n3748 ) | ( ~n3734 & n3748 ) ;
  assign n3750 = n3734 & n3749 ;
  assign n3751 = n3729 & ~n3732 ;
  assign n3752 = ~n3729 & n3732 ;
  assign n3753 = n3751 | n3752 ;
  assign n3754 = n3739 & ~n3742 ;
  assign n3755 = ~n3739 & n3742 ;
  assign n3756 = n3754 | n3755 ;
  assign n3757 = n3753 & n3756 ;
  assign n3758 = ~n3750 & n3757 ;
  assign n3759 = n3749 & n3758 ;
  assign n3760 = ~n3747 & n3759 ;
  assign n3761 = ~n3747 & n3758 ;
  assign n3762 = ~n3749 & n3761 ;
  assign n3763 = ( n3746 & n3749 ) | ( n3746 & n3762 ) | ( n3749 & n3762 ) ;
  assign n3764 = n3760 | n3763 ;
  assign n3765 = ( n3734 & n3744 ) | ( n3734 & n3764 ) | ( n3744 & n3764 ) ;
  assign n3766 = ( n3746 & n3749 ) | ( n3746 & ~n3761 ) | ( n3749 & ~n3761 ) ;
  assign n3767 = n3746 & ~n3760 ;
  assign n3768 = ( n3749 & ~n3766 ) | ( n3749 & n3767 ) | ( ~n3766 & n3767 ) ;
  assign n3769 = ( n3762 & n3766 ) | ( n3762 & ~n3768 ) | ( n3766 & ~n3768 ) ;
  assign n3770 = ~n3717 & n3720 ;
  assign n3771 = n3717 & ~n3720 ;
  assign n3772 = n3770 | n3771 ;
  assign n3773 = ~n3753 & n3756 ;
  assign n3774 = n3753 & ~n3756 ;
  assign n3775 = n3773 | n3774 ;
  assign n3776 = n3772 & n3775 ;
  assign n3777 = n3711 & n3721 ;
  assign n3778 = n3711 | n3722 ;
  assign n3779 = ( n3713 & n3777 ) | ( n3713 & ~n3778 ) | ( n3777 & ~n3778 ) ;
  assign n3780 = ~n3723 & n3778 ;
  assign n3781 = n3779 | n3780 ;
  assign n3782 = n3776 | n3781 ;
  assign n3783 = n3769 & n3782 ;
  assign n3784 = ( n3776 & n3779 ) | ( n3776 & n3780 ) | ( n3779 & n3780 ) ;
  assign n3785 = n3783 | n3784 ;
  assign n3786 = n3734 & ~n3744 ;
  assign n3787 = ~n3734 & n3744 ;
  assign n3788 = n3786 | n3787 ;
  assign n3789 = n3760 | n3788 ;
  assign n3790 = n3763 | n3789 ;
  assign n3791 = n3764 & n3788 ;
  assign n3792 = n3790 & ~n3791 ;
  assign n3793 = ( n3699 & n3709 ) | ( n3699 & ~n3723 ) | ( n3709 & ~n3723 ) ;
  assign n3794 = ( n3699 & ~n3709 ) | ( n3699 & n3723 ) | ( ~n3709 & n3723 ) ;
  assign n3795 = ( ~n3699 & n3793 ) | ( ~n3699 & n3794 ) | ( n3793 & n3794 ) ;
  assign n3796 = ( n3785 & n3792 ) | ( n3785 & n3795 ) | ( n3792 & n3795 ) ;
  assign n3797 = ( n3724 & n3765 ) | ( n3724 & n3796 ) | ( n3765 & n3796 ) ;
  assign n3798 = ( x76 & x77 ) | ( x76 & x78 ) | ( x77 & x78 ) ;
  assign n3799 = ( x73 & x74 ) | ( x73 & x75 ) | ( x74 & x75 ) ;
  assign n3800 = ( x73 & ~x74 ) | ( x73 & x75 ) | ( ~x74 & x75 ) ;
  assign n3801 = ( ~x73 & x74 ) | ( ~x73 & n3800 ) | ( x74 & n3800 ) ;
  assign n3802 = ( ~x75 & n3800 ) | ( ~x75 & n3801 ) | ( n3800 & n3801 ) ;
  assign n3803 = ( x76 & ~x77 ) | ( x76 & x78 ) | ( ~x77 & x78 ) ;
  assign n3804 = ( ~x76 & x77 ) | ( ~x76 & n3803 ) | ( x77 & n3803 ) ;
  assign n3805 = ( ~x78 & n3803 ) | ( ~x78 & n3804 ) | ( n3803 & n3804 ) ;
  assign n3806 = n3802 & n3805 ;
  assign n3807 = ( n3798 & n3799 ) | ( n3798 & n3806 ) | ( n3799 & n3806 ) ;
  assign n3808 = ( x67 & ~x68 ) | ( x67 & x69 ) | ( ~x68 & x69 ) ;
  assign n3809 = ( ~x67 & x68 ) | ( ~x67 & n3808 ) | ( x68 & n3808 ) ;
  assign n3810 = ( ~x69 & n3808 ) | ( ~x69 & n3809 ) | ( n3808 & n3809 ) ;
  assign n3811 = ( x70 & ~x71 ) | ( x70 & x72 ) | ( ~x71 & x72 ) ;
  assign n3812 = ( ~x70 & x71 ) | ( ~x70 & n3811 ) | ( x71 & n3811 ) ;
  assign n3813 = ( ~x72 & n3811 ) | ( ~x72 & n3812 ) | ( n3811 & n3812 ) ;
  assign n3814 = n3810 & n3813 ;
  assign n3815 = ( x70 & x71 ) | ( x70 & x72 ) | ( x71 & x72 ) ;
  assign n3816 = ( x67 & x68 ) | ( x67 & x69 ) | ( x68 & x69 ) ;
  assign n3817 = ( n3814 & n3815 ) | ( n3814 & n3816 ) | ( n3815 & n3816 ) ;
  assign n3818 = ( n3799 & n3806 ) | ( n3799 & ~n3807 ) | ( n3806 & ~n3807 ) ;
  assign n3819 = ( n3798 & ~n3807 ) | ( n3798 & n3818 ) | ( ~n3807 & n3818 ) ;
  assign n3820 = ( n3814 & n3816 ) | ( n3814 & ~n3817 ) | ( n3816 & ~n3817 ) ;
  assign n3821 = ( n3815 & ~n3817 ) | ( n3815 & n3820 ) | ( ~n3817 & n3820 ) ;
  assign n3822 = n3817 & n3821 ;
  assign n3823 = n3810 & ~n3813 ;
  assign n3824 = ~n3810 & n3813 ;
  assign n3825 = n3823 | n3824 ;
  assign n3826 = n3802 & ~n3805 ;
  assign n3827 = ~n3802 & n3805 ;
  assign n3828 = n3826 | n3827 ;
  assign n3829 = ~n3806 & n3828 ;
  assign n3830 = n3825 & n3829 ;
  assign n3831 = ~n3822 & n3830 ;
  assign n3832 = ( n3819 & n3821 ) | ( n3819 & n3831 ) | ( n3821 & n3831 ) ;
  assign n3833 = ( n3807 & n3817 ) | ( n3807 & n3832 ) | ( n3817 & n3832 ) ;
  assign n3834 = ( x55 & ~x56 ) | ( x55 & x57 ) | ( ~x56 & x57 ) ;
  assign n3835 = ( ~x55 & x56 ) | ( ~x55 & n3834 ) | ( x56 & n3834 ) ;
  assign n3836 = ( ~x57 & n3834 ) | ( ~x57 & n3835 ) | ( n3834 & n3835 ) ;
  assign n3837 = ( x58 & ~x59 ) | ( x58 & x60 ) | ( ~x59 & x60 ) ;
  assign n3838 = ( ~x58 & x59 ) | ( ~x58 & n3837 ) | ( x59 & n3837 ) ;
  assign n3839 = ( ~x60 & n3837 ) | ( ~x60 & n3838 ) | ( n3837 & n3838 ) ;
  assign n3840 = n3836 & n3839 ;
  assign n3841 = ( x58 & x59 ) | ( x58 & x60 ) | ( x59 & x60 ) ;
  assign n3842 = ( x55 & x56 ) | ( x55 & x57 ) | ( x56 & x57 ) ;
  assign n3843 = ( n3840 & n3841 ) | ( n3840 & n3842 ) | ( n3841 & n3842 ) ;
  assign n3844 = ( x64 & x65 ) | ( x64 & x66 ) | ( x65 & x66 ) ;
  assign n3845 = ( x61 & x62 ) | ( x61 & x63 ) | ( x62 & x63 ) ;
  assign n3846 = ( x61 & ~x62 ) | ( x61 & x63 ) | ( ~x62 & x63 ) ;
  assign n3847 = ( ~x61 & x62 ) | ( ~x61 & n3846 ) | ( x62 & n3846 ) ;
  assign n3848 = ( ~x63 & n3846 ) | ( ~x63 & n3847 ) | ( n3846 & n3847 ) ;
  assign n3849 = ( x64 & ~x65 ) | ( x64 & x66 ) | ( ~x65 & x66 ) ;
  assign n3850 = ( ~x64 & x65 ) | ( ~x64 & n3849 ) | ( x65 & n3849 ) ;
  assign n3851 = ( ~x66 & n3849 ) | ( ~x66 & n3850 ) | ( n3849 & n3850 ) ;
  assign n3852 = n3848 & n3851 ;
  assign n3853 = ( n3844 & n3845 ) | ( n3844 & n3852 ) | ( n3845 & n3852 ) ;
  assign n3854 = ( n3840 & n3842 ) | ( n3840 & ~n3843 ) | ( n3842 & ~n3843 ) ;
  assign n3855 = ( n3841 & ~n3843 ) | ( n3841 & n3854 ) | ( ~n3843 & n3854 ) ;
  assign n3856 = ( n3845 & n3852 ) | ( n3845 & ~n3853 ) | ( n3852 & ~n3853 ) ;
  assign n3857 = ( n3844 & ~n3853 ) | ( n3844 & n3856 ) | ( ~n3853 & n3856 ) ;
  assign n3858 = n3843 & n3855 ;
  assign n3859 = n3853 & n3857 ;
  assign n3860 = n3836 & ~n3839 ;
  assign n3861 = ~n3836 & n3839 ;
  assign n3862 = n3860 | n3861 ;
  assign n3863 = n3848 & ~n3851 ;
  assign n3864 = ~n3848 & n3851 ;
  assign n3865 = n3863 | n3864 ;
  assign n3866 = n3862 & n3865 ;
  assign n3867 = ~n3859 & n3866 ;
  assign n3868 = ~n3858 & n3867 ;
  assign n3869 = ~n3857 & n3868 ;
  assign n3870 = ( n3855 & n3857 ) | ( n3855 & n3869 ) | ( n3857 & n3869 ) ;
  assign n3871 = n3857 & n3867 ;
  assign n3872 = ~n3858 & n3871 ;
  assign n3873 = n3870 | n3872 ;
  assign n3874 = ( n3843 & n3853 ) | ( n3843 & n3873 ) | ( n3853 & n3873 ) ;
  assign n3875 = ~n3843 & n3853 ;
  assign n3876 = n3843 & ~n3853 ;
  assign n3877 = n3875 | n3876 ;
  assign n3878 = n3872 | n3877 ;
  assign n3879 = n3870 | n3878 ;
  assign n3880 = n3873 & n3877 ;
  assign n3881 = n3879 & ~n3880 ;
  assign n3882 = ( n3807 & n3817 ) | ( n3807 & ~n3832 ) | ( n3817 & ~n3832 ) ;
  assign n3883 = ( n3807 & ~n3817 ) | ( n3807 & n3832 ) | ( ~n3817 & n3832 ) ;
  assign n3884 = ( ~n3807 & n3882 ) | ( ~n3807 & n3883 ) | ( n3882 & n3883 ) ;
  assign n3885 = n3881 | n3884 ;
  assign n3886 = ( n3855 & n3857 ) | ( n3855 & ~n3868 ) | ( n3857 & ~n3868 ) ;
  assign n3887 = n3855 & ~n3872 ;
  assign n3888 = ( n3857 & ~n3886 ) | ( n3857 & n3887 ) | ( ~n3886 & n3887 ) ;
  assign n3889 = ( n3869 & n3886 ) | ( n3869 & ~n3888 ) | ( n3886 & ~n3888 ) ;
  assign n3890 = n3825 & ~n3829 ;
  assign n3891 = ~n3825 & n3829 ;
  assign n3892 = n3890 | n3891 ;
  assign n3893 = n3862 & ~n3865 ;
  assign n3894 = ~n3862 & n3865 ;
  assign n3895 = n3893 | n3894 ;
  assign n3896 = n3892 & n3895 ;
  assign n3897 = n3819 | n3831 ;
  assign n3898 = ~n3832 & n3897 ;
  assign n3899 = n3819 & n3830 ;
  assign n3900 = ( n3821 & ~n3897 ) | ( n3821 & n3899 ) | ( ~n3897 & n3899 ) ;
  assign n3901 = n3898 | n3900 ;
  assign n3902 = n3896 | n3901 ;
  assign n3903 = ( n3896 & n3898 ) | ( n3896 & n3900 ) | ( n3898 & n3900 ) ;
  assign n3904 = ( n3889 & n3902 ) | ( n3889 & n3903 ) | ( n3902 & n3903 ) ;
  assign n3905 = n3885 & n3904 ;
  assign n3906 = n3881 & n3884 ;
  assign n3907 = n3905 | n3906 ;
  assign n3908 = ( n3833 & n3874 ) | ( n3833 & n3907 ) | ( n3874 & n3907 ) ;
  assign n3909 = n3797 & n3908 ;
  assign n3910 = ~n3833 & n3874 ;
  assign n3911 = n3833 & ~n3874 ;
  assign n3912 = n3910 | n3911 ;
  assign n3913 = n3906 | n3912 ;
  assign n3914 = n3905 | n3913 ;
  assign n3915 = n3907 & n3912 ;
  assign n3916 = n3914 & ~n3915 ;
  assign n3917 = ~n3724 & n3765 ;
  assign n3918 = n3724 & ~n3765 ;
  assign n3919 = n3917 | n3918 ;
  assign n3920 = n3796 | n3919 ;
  assign n3921 = ~n3919 & n3920 ;
  assign n3922 = ( ~n3796 & n3920 ) | ( ~n3796 & n3921 ) | ( n3920 & n3921 ) ;
  assign n3923 = n3916 | n3922 ;
  assign n3924 = ( n3785 & ~n3792 ) | ( n3785 & n3795 ) | ( ~n3792 & n3795 ) ;
  assign n3925 = ( ~n3785 & n3792 ) | ( ~n3785 & n3924 ) | ( n3792 & n3924 ) ;
  assign n3926 = ( ~n3795 & n3924 ) | ( ~n3795 & n3925 ) | ( n3924 & n3925 ) ;
  assign n3927 = ( ~n3881 & n3884 ) | ( ~n3881 & n3904 ) | ( n3884 & n3904 ) ;
  assign n3928 = ( n3881 & ~n3904 ) | ( n3881 & n3927 ) | ( ~n3904 & n3927 ) ;
  assign n3929 = ( ~n3884 & n3927 ) | ( ~n3884 & n3928 ) | ( n3927 & n3928 ) ;
  assign n3930 = n3892 & ~n3895 ;
  assign n3931 = ~n3892 & n3895 ;
  assign n3932 = n3930 | n3931 ;
  assign n3933 = n3772 & ~n3775 ;
  assign n3934 = ~n3772 & n3775 ;
  assign n3935 = n3933 | n3934 ;
  assign n3936 = n3932 & n3935 ;
  assign n3937 = ~n3896 & n3902 ;
  assign n3938 = ( ~n3901 & n3902 ) | ( ~n3901 & n3937 ) | ( n3902 & n3937 ) ;
  assign n3939 = n3889 & ~n3938 ;
  assign n3940 = ~n3889 & n3938 ;
  assign n3941 = n3939 | n3940 ;
  assign n3942 = ( n3769 & n3776 ) | ( n3769 & ~n3781 ) | ( n3776 & ~n3781 ) ;
  assign n3943 = ( ~n3769 & n3781 ) | ( ~n3769 & n3942 ) | ( n3781 & n3942 ) ;
  assign n3944 = ( ~n3776 & n3942 ) | ( ~n3776 & n3943 ) | ( n3942 & n3943 ) ;
  assign n3945 = ( n3936 & n3941 ) | ( n3936 & n3944 ) | ( n3941 & n3944 ) ;
  assign n3946 = ( n3926 & n3929 ) | ( n3926 & n3945 ) | ( n3929 & n3945 ) ;
  assign n3947 = n3923 & n3946 ;
  assign n3948 = n3916 & n3922 ;
  assign n3949 = n3947 | n3948 ;
  assign n3950 = n3908 & ~n3909 ;
  assign n3951 = ( n3797 & ~n3909 ) | ( n3797 & n3950 ) | ( ~n3909 & n3950 ) ;
  assign n3952 = n3949 & n3951 ;
  assign n3953 = ( n3908 & n3949 ) | ( n3908 & n3952 ) | ( n3949 & n3952 ) ;
  assign n3954 = n3909 | n3953 ;
  assign n3955 = n3689 & n3954 ;
  assign n3956 = n3954 & ~n3955 ;
  assign n3957 = ( n3689 & ~n3955 ) | ( n3689 & n3956 ) | ( ~n3955 & n3956 ) ;
  assign n3958 = n3948 | n3951 ;
  assign n3959 = n3947 | n3958 ;
  assign n3960 = ~n3952 & n3959 ;
  assign n3961 = ( ~n3658 & n3687 ) | ( ~n3658 & n3688 ) | ( n3687 & n3688 ) ;
  assign n3962 = ( n3658 & ~n3687 ) | ( n3658 & n3961 ) | ( ~n3687 & n3961 ) ;
  assign n3963 = ( ~n3688 & n3961 ) | ( ~n3688 & n3962 ) | ( n3961 & n3962 ) ;
  assign n3964 = ( ~n3665 & n3668 ) | ( ~n3665 & n3682 ) | ( n3668 & n3682 ) ;
  assign n3965 = ( n3665 & ~n3682 ) | ( n3665 & n3964 ) | ( ~n3682 & n3964 ) ;
  assign n3966 = ( ~n3668 & n3964 ) | ( ~n3668 & n3965 ) | ( n3964 & n3965 ) ;
  assign n3967 = ( ~n3926 & n3929 ) | ( ~n3926 & n3945 ) | ( n3929 & n3945 ) ;
  assign n3968 = ( n3926 & ~n3945 ) | ( n3926 & n3967 ) | ( ~n3945 & n3967 ) ;
  assign n3969 = ( ~n3929 & n3967 ) | ( ~n3929 & n3968 ) | ( n3967 & n3968 ) ;
  assign n3970 = n3932 & ~n3935 ;
  assign n3971 = ~n3932 & n3935 ;
  assign n3972 = n3970 | n3971 ;
  assign n3973 = n3671 | n3673 ;
  assign n3974 = ~n3673 & n3973 ;
  assign n3975 = ( ~n3671 & n3973 ) | ( ~n3671 & n3974 ) | ( n3973 & n3974 ) ;
  assign n3976 = n3972 & n3975 ;
  assign n3977 = ( n3936 & ~n3941 ) | ( n3936 & n3944 ) | ( ~n3941 & n3944 ) ;
  assign n3978 = ( ~n3936 & n3941 ) | ( ~n3936 & n3977 ) | ( n3941 & n3977 ) ;
  assign n3979 = ( ~n3944 & n3977 ) | ( ~n3944 & n3978 ) | ( n3977 & n3978 ) ;
  assign n3980 = ( n3674 & ~n3679 ) | ( n3674 & n3681 ) | ( ~n3679 & n3681 ) ;
  assign n3981 = ( ~n3674 & n3679 ) | ( ~n3674 & n3980 ) | ( n3679 & n3980 ) ;
  assign n3982 = ( ~n3681 & n3980 ) | ( ~n3681 & n3981 ) | ( n3980 & n3981 ) ;
  assign n3983 = ( n3976 & n3979 ) | ( n3976 & n3982 ) | ( n3979 & n3982 ) ;
  assign n3984 = ( n3966 & n3969 ) | ( n3966 & n3983 ) | ( n3969 & n3983 ) ;
  assign n3985 = ( ~n3916 & n3922 ) | ( ~n3916 & n3946 ) | ( n3922 & n3946 ) ;
  assign n3986 = ( n3916 & ~n3946 ) | ( n3916 & n3985 ) | ( ~n3946 & n3985 ) ;
  assign n3987 = ( ~n3922 & n3985 ) | ( ~n3922 & n3986 ) | ( n3985 & n3986 ) ;
  assign n3988 = ( n3663 & n3683 ) | ( n3663 & ~n3687 ) | ( n3683 & ~n3687 ) ;
  assign n3989 = ( n3686 & ~n3687 ) | ( n3686 & n3988 ) | ( ~n3687 & n3988 ) ;
  assign n3990 = ( n3984 & n3987 ) | ( n3984 & n3989 ) | ( n3987 & n3989 ) ;
  assign n3991 = ( n3960 & n3963 ) | ( n3960 & n3990 ) | ( n3963 & n3990 ) ;
  assign n3992 = n3957 & n3991 ;
  assign n3993 = n3957 | n3991 ;
  assign n3994 = ~n3992 & n3993 ;
  assign n3995 = ( x988 & x989 ) | ( x988 & x990 ) | ( x989 & x990 ) ;
  assign n3996 = ( x985 & x986 ) | ( x985 & x987 ) | ( x986 & x987 ) ;
  assign n3997 = ( x985 & ~x986 ) | ( x985 & x987 ) | ( ~x986 & x987 ) ;
  assign n3998 = ( ~x985 & x986 ) | ( ~x985 & n3997 ) | ( x986 & n3997 ) ;
  assign n3999 = ( ~x987 & n3997 ) | ( ~x987 & n3998 ) | ( n3997 & n3998 ) ;
  assign n4000 = ( x988 & ~x989 ) | ( x988 & x990 ) | ( ~x989 & x990 ) ;
  assign n4001 = ( ~x988 & x989 ) | ( ~x988 & n4000 ) | ( x989 & n4000 ) ;
  assign n4002 = ( ~x990 & n4000 ) | ( ~x990 & n4001 ) | ( n4000 & n4001 ) ;
  assign n4003 = n3999 & n4002 ;
  assign n4004 = ( n3995 & n3996 ) | ( n3995 & n4003 ) | ( n3996 & n4003 ) ;
  assign n4005 = ( x979 & ~x980 ) | ( x979 & x981 ) | ( ~x980 & x981 ) ;
  assign n4006 = ( ~x979 & x980 ) | ( ~x979 & n4005 ) | ( x980 & n4005 ) ;
  assign n4007 = ( ~x981 & n4005 ) | ( ~x981 & n4006 ) | ( n4005 & n4006 ) ;
  assign n4008 = ( x982 & ~x983 ) | ( x982 & x984 ) | ( ~x983 & x984 ) ;
  assign n4009 = ( ~x982 & x983 ) | ( ~x982 & n4008 ) | ( x983 & n4008 ) ;
  assign n4010 = ( ~x984 & n4008 ) | ( ~x984 & n4009 ) | ( n4008 & n4009 ) ;
  assign n4011 = n4007 & n4010 ;
  assign n4012 = ( x982 & x983 ) | ( x982 & x984 ) | ( x983 & x984 ) ;
  assign n4013 = ( x979 & x980 ) | ( x979 & x981 ) | ( x980 & x981 ) ;
  assign n4014 = ( n4011 & n4012 ) | ( n4011 & n4013 ) | ( n4012 & n4013 ) ;
  assign n4015 = ( n3996 & n4003 ) | ( n3996 & ~n4004 ) | ( n4003 & ~n4004 ) ;
  assign n4016 = ( n3995 & ~n4004 ) | ( n3995 & n4015 ) | ( ~n4004 & n4015 ) ;
  assign n4017 = ( n4011 & n4013 ) | ( n4011 & ~n4014 ) | ( n4013 & ~n4014 ) ;
  assign n4018 = ( n4012 & ~n4014 ) | ( n4012 & n4017 ) | ( ~n4014 & n4017 ) ;
  assign n4019 = n4014 & n4018 ;
  assign n4020 = n4007 & ~n4010 ;
  assign n4021 = ~n4007 & n4010 ;
  assign n4022 = n4020 | n4021 ;
  assign n4023 = n3999 & ~n4002 ;
  assign n4024 = ~n3999 & n4002 ;
  assign n4025 = n4023 | n4024 ;
  assign n4026 = ~n4003 & n4025 ;
  assign n4027 = n4022 & n4026 ;
  assign n4028 = ~n4019 & n4027 ;
  assign n4029 = ( n4016 & n4018 ) | ( n4016 & n4028 ) | ( n4018 & n4028 ) ;
  assign n4030 = ( n4004 & n4014 ) | ( n4004 & n4029 ) | ( n4014 & n4029 ) ;
  assign n4031 = ( x967 & ~x968 ) | ( x967 & x969 ) | ( ~x968 & x969 ) ;
  assign n4032 = ( ~x967 & x968 ) | ( ~x967 & n4031 ) | ( x968 & n4031 ) ;
  assign n4033 = ( ~x969 & n4031 ) | ( ~x969 & n4032 ) | ( n4031 & n4032 ) ;
  assign n4034 = ( x970 & ~x971 ) | ( x970 & x972 ) | ( ~x971 & x972 ) ;
  assign n4035 = ( ~x970 & x971 ) | ( ~x970 & n4034 ) | ( x971 & n4034 ) ;
  assign n4036 = ( ~x972 & n4034 ) | ( ~x972 & n4035 ) | ( n4034 & n4035 ) ;
  assign n4037 = n4033 & n4036 ;
  assign n4038 = ( x970 & x971 ) | ( x970 & x972 ) | ( x971 & x972 ) ;
  assign n4039 = ( x967 & x968 ) | ( x967 & x969 ) | ( x968 & x969 ) ;
  assign n4040 = ( n4037 & n4038 ) | ( n4037 & n4039 ) | ( n4038 & n4039 ) ;
  assign n4041 = ( x976 & x977 ) | ( x976 & x978 ) | ( x977 & x978 ) ;
  assign n4042 = ( x973 & x974 ) | ( x973 & x975 ) | ( x974 & x975 ) ;
  assign n4043 = ( x973 & ~x974 ) | ( x973 & x975 ) | ( ~x974 & x975 ) ;
  assign n4044 = ( ~x973 & x974 ) | ( ~x973 & n4043 ) | ( x974 & n4043 ) ;
  assign n4045 = ( ~x975 & n4043 ) | ( ~x975 & n4044 ) | ( n4043 & n4044 ) ;
  assign n4046 = ( x976 & ~x977 ) | ( x976 & x978 ) | ( ~x977 & x978 ) ;
  assign n4047 = ( ~x976 & x977 ) | ( ~x976 & n4046 ) | ( x977 & n4046 ) ;
  assign n4048 = ( ~x978 & n4046 ) | ( ~x978 & n4047 ) | ( n4046 & n4047 ) ;
  assign n4049 = n4045 & n4048 ;
  assign n4050 = ( n4041 & n4042 ) | ( n4041 & n4049 ) | ( n4042 & n4049 ) ;
  assign n4051 = ( n4037 & n4039 ) | ( n4037 & ~n4040 ) | ( n4039 & ~n4040 ) ;
  assign n4052 = ( n4038 & ~n4040 ) | ( n4038 & n4051 ) | ( ~n4040 & n4051 ) ;
  assign n4053 = ( n4042 & n4049 ) | ( n4042 & ~n4050 ) | ( n4049 & ~n4050 ) ;
  assign n4054 = ( n4041 & ~n4050 ) | ( n4041 & n4053 ) | ( ~n4050 & n4053 ) ;
  assign n4055 = n4040 & n4052 ;
  assign n4056 = n4050 & n4054 ;
  assign n4057 = n4033 & ~n4036 ;
  assign n4058 = ~n4033 & n4036 ;
  assign n4059 = n4057 | n4058 ;
  assign n4060 = n4045 & ~n4048 ;
  assign n4061 = ~n4045 & n4048 ;
  assign n4062 = n4060 | n4061 ;
  assign n4063 = n4059 & n4062 ;
  assign n4064 = ~n4056 & n4063 ;
  assign n4065 = ~n4055 & n4064 ;
  assign n4066 = ~n4054 & n4065 ;
  assign n4067 = ( n4052 & n4054 ) | ( n4052 & n4066 ) | ( n4054 & n4066 ) ;
  assign n4068 = n4054 & n4064 ;
  assign n4069 = ~n4055 & n4068 ;
  assign n4070 = n4067 | n4069 ;
  assign n4071 = ( n4040 & n4050 ) | ( n4040 & n4070 ) | ( n4050 & n4070 ) ;
  assign n4072 = ~n4040 & n4050 ;
  assign n4073 = n4040 & ~n4050 ;
  assign n4074 = n4072 | n4073 ;
  assign n4075 = n4069 | n4074 ;
  assign n4076 = n4067 | n4075 ;
  assign n4077 = n4070 & n4074 ;
  assign n4078 = n4076 & ~n4077 ;
  assign n4079 = ( n4004 & n4014 ) | ( n4004 & ~n4029 ) | ( n4014 & ~n4029 ) ;
  assign n4080 = ( n4004 & ~n4014 ) | ( n4004 & n4029 ) | ( ~n4014 & n4029 ) ;
  assign n4081 = ( ~n4004 & n4079 ) | ( ~n4004 & n4080 ) | ( n4079 & n4080 ) ;
  assign n4082 = n4078 | n4081 ;
  assign n4083 = ( n4052 & n4054 ) | ( n4052 & ~n4065 ) | ( n4054 & ~n4065 ) ;
  assign n4084 = n4052 & ~n4069 ;
  assign n4085 = ( n4054 & ~n4083 ) | ( n4054 & n4084 ) | ( ~n4083 & n4084 ) ;
  assign n4086 = ( n4066 & n4083 ) | ( n4066 & ~n4085 ) | ( n4083 & ~n4085 ) ;
  assign n4087 = n4022 & ~n4026 ;
  assign n4088 = ~n4022 & n4026 ;
  assign n4089 = n4087 | n4088 ;
  assign n4090 = n4059 & ~n4062 ;
  assign n4091 = ~n4059 & n4062 ;
  assign n4092 = n4090 | n4091 ;
  assign n4093 = n4089 & n4092 ;
  assign n4094 = n4016 | n4028 ;
  assign n4095 = ~n4029 & n4094 ;
  assign n4096 = n4016 & n4027 ;
  assign n4097 = ( n4018 & ~n4094 ) | ( n4018 & n4096 ) | ( ~n4094 & n4096 ) ;
  assign n4098 = n4095 | n4097 ;
  assign n4099 = n4093 | n4098 ;
  assign n4100 = ( n4093 & n4095 ) | ( n4093 & n4097 ) | ( n4095 & n4097 ) ;
  assign n4101 = ( n4086 & n4099 ) | ( n4086 & n4100 ) | ( n4099 & n4100 ) ;
  assign n4102 = n4082 & n4101 ;
  assign n4103 = n4078 & n4081 ;
  assign n4104 = n4102 | n4103 ;
  assign n4105 = ( n4030 & n4071 ) | ( n4030 & n4104 ) | ( n4071 & n4104 ) ;
  assign n4217 = ~n4030 & n4071 ;
  assign n4218 = n4030 & ~n4071 ;
  assign n4219 = n4217 | n4218 ;
  assign n4220 = n4103 | n4219 ;
  assign n4221 = n4102 | n4220 ;
  assign n4222 = n4104 & n4219 ;
  assign n4223 = n4221 & ~n4222 ;
  assign n4141 = ( x952 & x953 ) | ( x952 & x954 ) | ( x953 & x954 ) ;
  assign n4142 = ( x949 & x950 ) | ( x949 & x951 ) | ( x950 & x951 ) ;
  assign n4143 = ( x949 & ~x950 ) | ( x949 & x951 ) | ( ~x950 & x951 ) ;
  assign n4144 = ( ~x949 & x950 ) | ( ~x949 & n4143 ) | ( x950 & n4143 ) ;
  assign n4145 = ( ~x951 & n4143 ) | ( ~x951 & n4144 ) | ( n4143 & n4144 ) ;
  assign n4146 = ( x952 & ~x953 ) | ( x952 & x954 ) | ( ~x953 & x954 ) ;
  assign n4147 = ( ~x952 & x953 ) | ( ~x952 & n4146 ) | ( x953 & n4146 ) ;
  assign n4148 = ( ~x954 & n4146 ) | ( ~x954 & n4147 ) | ( n4146 & n4147 ) ;
  assign n4149 = n4145 & n4148 ;
  assign n4150 = ( n4141 & n4142 ) | ( n4141 & n4149 ) | ( n4142 & n4149 ) ;
  assign n4164 = ( n4142 & n4149 ) | ( n4142 & ~n4150 ) | ( n4149 & ~n4150 ) ;
  assign n4165 = ( n4141 & ~n4150 ) | ( n4141 & n4164 ) | ( ~n4150 & n4164 ) ;
  assign n4151 = ( x946 & x947 ) | ( x946 & x948 ) | ( x947 & x948 ) ;
  assign n4152 = ( x943 & x944 ) | ( x943 & x945 ) | ( x944 & x945 ) ;
  assign n4153 = ( x943 & ~x944 ) | ( x943 & x945 ) | ( ~x944 & x945 ) ;
  assign n4154 = ( ~x943 & x944 ) | ( ~x943 & n4153 ) | ( x944 & n4153 ) ;
  assign n4155 = ( ~x945 & n4153 ) | ( ~x945 & n4154 ) | ( n4153 & n4154 ) ;
  assign n4156 = ( x946 & ~x947 ) | ( x946 & x948 ) | ( ~x947 & x948 ) ;
  assign n4157 = ( ~x946 & x947 ) | ( ~x946 & n4156 ) | ( x947 & n4156 ) ;
  assign n4158 = ( ~x948 & n4156 ) | ( ~x948 & n4157 ) | ( n4156 & n4157 ) ;
  assign n4159 = n4155 & n4158 ;
  assign n4160 = ( n4151 & n4152 ) | ( n4151 & n4159 ) | ( n4152 & n4159 ) ;
  assign n4161 = ( n4152 & n4159 ) | ( n4152 & ~n4160 ) | ( n4159 & ~n4160 ) ;
  assign n4162 = ( n4151 & ~n4160 ) | ( n4151 & n4161 ) | ( ~n4160 & n4161 ) ;
  assign n4163 = n4160 & n4162 ;
  assign n4166 = n4150 & n4165 ;
  assign n4167 = n4145 & ~n4148 ;
  assign n4168 = ~n4145 & n4148 ;
  assign n4169 = n4167 | n4168 ;
  assign n4170 = n4155 & ~n4158 ;
  assign n4171 = ~n4155 & n4158 ;
  assign n4172 = n4170 | n4171 ;
  assign n4173 = n4169 & n4172 ;
  assign n4174 = ~n4166 & n4173 ;
  assign n4177 = ~n4163 & n4174 ;
  assign n4178 = ~n4165 & n4177 ;
  assign n4182 = ( n4162 & n4165 ) | ( n4162 & ~n4177 ) | ( n4165 & ~n4177 ) ;
  assign n4175 = n4165 & n4174 ;
  assign n4176 = ~n4163 & n4175 ;
  assign n4183 = n4162 & ~n4176 ;
  assign n4184 = ( n4165 & ~n4182 ) | ( n4165 & n4183 ) | ( ~n4182 & n4183 ) ;
  assign n4185 = ( n4178 & n4182 ) | ( n4178 & ~n4184 ) | ( n4182 & ~n4184 ) ;
  assign n4108 = ( x955 & ~x956 ) | ( x955 & x957 ) | ( ~x956 & x957 ) ;
  assign n4109 = ( ~x955 & x956 ) | ( ~x955 & n4108 ) | ( x956 & n4108 ) ;
  assign n4110 = ( ~x957 & n4108 ) | ( ~x957 & n4109 ) | ( n4108 & n4109 ) ;
  assign n4111 = ( x958 & ~x959 ) | ( x958 & x960 ) | ( ~x959 & x960 ) ;
  assign n4112 = ( ~x958 & x959 ) | ( ~x958 & n4111 ) | ( x959 & n4111 ) ;
  assign n4113 = ( ~x960 & n4111 ) | ( ~x960 & n4112 ) | ( n4111 & n4112 ) ;
  assign n4131 = n4110 & ~n4113 ;
  assign n4132 = ~n4110 & n4113 ;
  assign n4133 = n4131 | n4132 ;
  assign n4118 = ( x961 & ~x962 ) | ( x961 & x963 ) | ( ~x962 & x963 ) ;
  assign n4119 = ( ~x961 & x962 ) | ( ~x961 & n4118 ) | ( x962 & n4118 ) ;
  assign n4120 = ( ~x963 & n4118 ) | ( ~x963 & n4119 ) | ( n4118 & n4119 ) ;
  assign n4121 = ( x964 & ~x965 ) | ( x964 & x966 ) | ( ~x965 & x966 ) ;
  assign n4122 = ( ~x964 & x965 ) | ( ~x964 & n4121 ) | ( x965 & n4121 ) ;
  assign n4123 = ( ~x966 & n4121 ) | ( ~x966 & n4122 ) | ( n4121 & n4122 ) ;
  assign n4134 = n4120 & ~n4123 ;
  assign n4135 = ~n4120 & n4123 ;
  assign n4136 = n4134 | n4135 ;
  assign n4186 = n4133 & ~n4136 ;
  assign n4187 = ~n4133 & n4136 ;
  assign n4188 = n4186 | n4187 ;
  assign n4189 = ~n4169 & n4172 ;
  assign n4190 = n4169 & ~n4172 ;
  assign n4191 = n4189 | n4190 ;
  assign n4192 = n4188 & n4191 ;
  assign n4106 = ( x958 & x959 ) | ( x958 & x960 ) | ( x959 & x960 ) ;
  assign n4107 = ( x955 & x956 ) | ( x955 & x957 ) | ( x956 & x957 ) ;
  assign n4114 = n4110 & n4113 ;
  assign n4115 = ( n4106 & n4107 ) | ( n4106 & n4114 ) | ( n4107 & n4114 ) ;
  assign n4126 = ( n4107 & n4114 ) | ( n4107 & ~n4115 ) | ( n4114 & ~n4115 ) ;
  assign n4127 = ( n4106 & ~n4115 ) | ( n4106 & n4126 ) | ( ~n4115 & n4126 ) ;
  assign n4116 = ( x964 & x965 ) | ( x964 & x966 ) | ( x965 & x966 ) ;
  assign n4117 = ( x961 & x962 ) | ( x961 & x963 ) | ( x962 & x963 ) ;
  assign n4124 = n4120 & n4123 ;
  assign n4125 = ( n4116 & n4117 ) | ( n4116 & n4124 ) | ( n4117 & n4124 ) ;
  assign n4128 = ( n4117 & n4124 ) | ( n4117 & ~n4125 ) | ( n4124 & ~n4125 ) ;
  assign n4129 = ( n4116 & ~n4125 ) | ( n4116 & n4128 ) | ( ~n4125 & n4128 ) ;
  assign n4137 = n4133 & n4136 ;
  assign n4193 = n4129 & n4137 ;
  assign n4130 = n4115 & n4127 ;
  assign n4138 = ~n4130 & n4137 ;
  assign n4194 = n4129 | n4138 ;
  assign n4195 = ( n4127 & n4193 ) | ( n4127 & ~n4194 ) | ( n4193 & ~n4194 ) ;
  assign n4139 = ( n4127 & n4129 ) | ( n4127 & n4138 ) | ( n4129 & n4138 ) ;
  assign n4196 = ~n4139 & n4194 ;
  assign n4197 = n4195 | n4196 ;
  assign n4198 = n4192 | n4197 ;
  assign n4199 = n4185 & n4198 ;
  assign n4200 = ( n4192 & n4195 ) | ( n4192 & n4196 ) | ( n4195 & n4196 ) ;
  assign n4201 = n4199 | n4200 ;
  assign n4179 = ( n4162 & n4165 ) | ( n4162 & n4178 ) | ( n4165 & n4178 ) ;
  assign n4202 = n4150 & ~n4160 ;
  assign n4203 = ~n4150 & n4160 ;
  assign n4204 = n4202 | n4203 ;
  assign n4205 = n4176 | n4204 ;
  assign n4206 = n4179 | n4205 ;
  assign n4180 = n4176 | n4179 ;
  assign n4207 = n4180 & n4204 ;
  assign n4208 = n4206 & ~n4207 ;
  assign n4209 = ~n4115 & n4125 ;
  assign n4210 = n4115 & ~n4125 ;
  assign n4211 = n4209 | n4210 ;
  assign n4212 = n4139 & n4211 ;
  assign n4213 = n4139 | n4211 ;
  assign n4214 = ~n4212 & n4213 ;
  assign n4215 = ( n4201 & n4208 ) | ( n4201 & n4214 ) | ( n4208 & n4214 ) ;
  assign n4140 = ( n4115 & n4125 ) | ( n4115 & n4139 ) | ( n4125 & n4139 ) ;
  assign n4181 = ( n4150 & n4160 ) | ( n4150 & n4180 ) | ( n4160 & n4180 ) ;
  assign n4224 = ~n4140 & n4181 ;
  assign n4225 = n4140 & ~n4181 ;
  assign n4226 = n4224 | n4225 ;
  assign n4227 = n4215 | n4226 ;
  assign n4228 = ~n4226 & n4227 ;
  assign n4229 = ( ~n4215 & n4227 ) | ( ~n4215 & n4228 ) | ( n4227 & n4228 ) ;
  assign n4230 = ( n4201 & ~n4208 ) | ( n4201 & n4214 ) | ( ~n4208 & n4214 ) ;
  assign n4231 = ( ~n4201 & n4208 ) | ( ~n4201 & n4230 ) | ( n4208 & n4230 ) ;
  assign n4232 = ( ~n4214 & n4230 ) | ( ~n4214 & n4231 ) | ( n4230 & n4231 ) ;
  assign n4233 = ( ~n4078 & n4081 ) | ( ~n4078 & n4101 ) | ( n4081 & n4101 ) ;
  assign n4234 = ( n4078 & ~n4101 ) | ( n4078 & n4233 ) | ( ~n4101 & n4233 ) ;
  assign n4235 = ( ~n4081 & n4233 ) | ( ~n4081 & n4234 ) | ( n4233 & n4234 ) ;
  assign n4236 = n4089 & ~n4092 ;
  assign n4237 = ~n4089 & n4092 ;
  assign n4238 = n4236 | n4237 ;
  assign n4239 = n4188 & ~n4191 ;
  assign n4240 = ~n4188 & n4191 ;
  assign n4241 = n4239 | n4240 ;
  assign n4242 = n4238 & n4241 ;
  assign n4243 = ~n4093 & n4099 ;
  assign n4244 = ( ~n4098 & n4099 ) | ( ~n4098 & n4243 ) | ( n4099 & n4243 ) ;
  assign n4245 = n4086 & ~n4244 ;
  assign n4246 = ~n4086 & n4244 ;
  assign n4247 = n4245 | n4246 ;
  assign n4248 = ( n4185 & n4192 ) | ( n4185 & ~n4197 ) | ( n4192 & ~n4197 ) ;
  assign n4249 = ( ~n4185 & n4197 ) | ( ~n4185 & n4248 ) | ( n4197 & n4248 ) ;
  assign n4250 = ( ~n4192 & n4248 ) | ( ~n4192 & n4249 ) | ( n4248 & n4249 ) ;
  assign n4251 = ( n4242 & n4247 ) | ( n4242 & n4250 ) | ( n4247 & n4250 ) ;
  assign n4252 = ( n4232 & n4235 ) | ( n4232 & n4251 ) | ( n4235 & n4251 ) ;
  assign n4253 = ( n4223 & n4229 ) | ( n4223 & n4252 ) | ( n4229 & n4252 ) ;
  assign n4216 = ( n4140 & n4181 ) | ( n4140 & n4215 ) | ( n4181 & n4215 ) ;
  assign n4254 = ( n4105 & n4216 ) | ( n4105 & ~n4253 ) | ( n4216 & ~n4253 ) ;
  assign n4255 = ( ~n4105 & n4253 ) | ( ~n4105 & n4254 ) | ( n4253 & n4254 ) ;
  assign n4256 = ( ~n4216 & n4254 ) | ( ~n4216 & n4255 ) | ( n4254 & n4255 ) ;
  assign n4257 = ( n4105 & n4253 ) | ( n4105 & ~n4256 ) | ( n4253 & ~n4256 ) ;
  assign n4258 = n3994 | n4257 ;
  assign n4259 = n3993 & n4257 ;
  assign n4260 = ~n3992 & n4259 ;
  assign n4261 = n3960 & ~n3963 ;
  assign n4262 = ~n3960 & n3963 ;
  assign n4263 = n4261 | n4262 ;
  assign n4264 = n3990 | n4263 ;
  assign n4265 = ( ~n4223 & n4229 ) | ( ~n4223 & n4252 ) | ( n4229 & n4252 ) ;
  assign n4266 = ( n4223 & ~n4252 ) | ( n4223 & n4265 ) | ( ~n4252 & n4265 ) ;
  assign n4267 = ( ~n4229 & n4265 ) | ( ~n4229 & n4266 ) | ( n4265 & n4266 ) ;
  assign n4268 = ( ~n4232 & n4235 ) | ( ~n4232 & n4251 ) | ( n4235 & n4251 ) ;
  assign n4269 = ( n4232 & ~n4251 ) | ( n4232 & n4268 ) | ( ~n4251 & n4268 ) ;
  assign n4270 = ( ~n4235 & n4268 ) | ( ~n4235 & n4269 ) | ( n4268 & n4269 ) ;
  assign n4271 = n3972 & ~n3975 ;
  assign n4272 = ~n3972 & n3975 ;
  assign n4273 = n4271 | n4272 ;
  assign n4274 = n4238 & ~n4241 ;
  assign n4275 = ~n4238 & n4241 ;
  assign n4276 = n4274 | n4275 ;
  assign n4277 = n4273 & n4276 ;
  assign n4278 = ~n3976 & n3979 ;
  assign n4279 = n3976 & ~n3979 ;
  assign n4280 = n4278 | n4279 ;
  assign n4281 = n3982 & ~n4280 ;
  assign n4282 = ~n3982 & n4280 ;
  assign n4283 = n4281 | n4282 ;
  assign n4284 = ( n4242 & ~n4247 ) | ( n4242 & n4250 ) | ( ~n4247 & n4250 ) ;
  assign n4285 = ( ~n4242 & n4247 ) | ( ~n4242 & n4284 ) | ( n4247 & n4284 ) ;
  assign n4286 = ( ~n4250 & n4284 ) | ( ~n4250 & n4285 ) | ( n4284 & n4285 ) ;
  assign n4287 = ( n4277 & n4283 ) | ( n4277 & n4286 ) | ( n4283 & n4286 ) ;
  assign n4288 = ( n3966 & ~n3969 ) | ( n3966 & n3983 ) | ( ~n3969 & n3983 ) ;
  assign n4289 = ( ~n3966 & n3969 ) | ( ~n3966 & n4288 ) | ( n3969 & n4288 ) ;
  assign n4290 = ( ~n3983 & n4288 ) | ( ~n3983 & n4289 ) | ( n4288 & n4289 ) ;
  assign n4291 = ( n4270 & n4287 ) | ( n4270 & n4290 ) | ( n4287 & n4290 ) ;
  assign n4292 = ( ~n3984 & n3987 ) | ( ~n3984 & n3989 ) | ( n3987 & n3989 ) ;
  assign n4293 = ( n3984 & ~n3989 ) | ( n3984 & n4292 ) | ( ~n3989 & n4292 ) ;
  assign n4294 = ( ~n3987 & n4292 ) | ( ~n3987 & n4293 ) | ( n4292 & n4293 ) ;
  assign n4295 = ( n4267 & n4291 ) | ( n4267 & n4294 ) | ( n4291 & n4294 ) ;
  assign n4296 = ( n3990 & n4256 ) | ( n3990 & ~n4263 ) | ( n4256 & ~n4263 ) ;
  assign n4297 = ( ~n3990 & n4263 ) | ( ~n3990 & n4296 ) | ( n4263 & n4296 ) ;
  assign n4298 = ( ~n4256 & n4296 ) | ( ~n4256 & n4297 ) | ( n4296 & n4297 ) ;
  assign n4299 = n4295 & n4298 ;
  assign n4300 = ( n3990 & ~n4256 ) | ( n3990 & n4263 ) | ( ~n4256 & n4263 ) ;
  assign n4301 = ( n4264 & n4299 ) | ( n4264 & ~n4300 ) | ( n4299 & ~n4300 ) ;
  assign n4302 = ( n4258 & n4260 ) | ( n4258 & n4301 ) | ( n4260 & n4301 ) ;
  assign n4303 = n3658 | n3909 ;
  assign n4304 = n3688 | n4303 ;
  assign n4305 = ( n3687 & n4303 ) | ( n3687 & n4304 ) | ( n4303 & n4304 ) ;
  assign n4306 = n3953 | n4305 ;
  assign n4307 = n3955 | n4306 ;
  assign n4308 = ( n3955 & n3991 ) | ( n3955 & n4307 ) | ( n3991 & n4307 ) ;
  assign n4309 = n4302 & ~n4308 ;
  assign n4310 = ( x874 & x875 ) | ( x874 & x876 ) | ( x875 & x876 ) ;
  assign n4311 = ( x871 & x872 ) | ( x871 & x873 ) | ( x872 & x873 ) ;
  assign n4312 = ( x871 & ~x872 ) | ( x871 & x873 ) | ( ~x872 & x873 ) ;
  assign n4313 = ( ~x871 & x872 ) | ( ~x871 & n4312 ) | ( x872 & n4312 ) ;
  assign n4314 = ( ~x873 & n4312 ) | ( ~x873 & n4313 ) | ( n4312 & n4313 ) ;
  assign n4315 = ( x874 & ~x875 ) | ( x874 & x876 ) | ( ~x875 & x876 ) ;
  assign n4316 = ( ~x874 & x875 ) | ( ~x874 & n4315 ) | ( x875 & n4315 ) ;
  assign n4317 = ( ~x876 & n4315 ) | ( ~x876 & n4316 ) | ( n4315 & n4316 ) ;
  assign n4318 = n4314 & n4317 ;
  assign n4319 = ( n4310 & n4311 ) | ( n4310 & n4318 ) | ( n4311 & n4318 ) ;
  assign n4320 = ( n4311 & n4318 ) | ( n4311 & ~n4319 ) | ( n4318 & ~n4319 ) ;
  assign n4321 = ( n4310 & ~n4319 ) | ( n4310 & n4320 ) | ( ~n4319 & n4320 ) ;
  assign n4322 = ( x880 & x881 ) | ( x880 & x882 ) | ( x881 & x882 ) ;
  assign n4323 = ( x877 & x878 ) | ( x877 & x879 ) | ( x878 & x879 ) ;
  assign n4324 = ( x877 & ~x878 ) | ( x877 & x879 ) | ( ~x878 & x879 ) ;
  assign n4325 = ( ~x877 & x878 ) | ( ~x877 & n4324 ) | ( x878 & n4324 ) ;
  assign n4326 = ( ~x879 & n4324 ) | ( ~x879 & n4325 ) | ( n4324 & n4325 ) ;
  assign n4327 = ( x880 & ~x881 ) | ( x880 & x882 ) | ( ~x881 & x882 ) ;
  assign n4328 = ( ~x880 & x881 ) | ( ~x880 & n4327 ) | ( x881 & n4327 ) ;
  assign n4329 = ( ~x882 & n4327 ) | ( ~x882 & n4328 ) | ( n4327 & n4328 ) ;
  assign n4330 = n4326 & n4329 ;
  assign n4331 = ( n4322 & n4323 ) | ( n4322 & n4330 ) | ( n4323 & n4330 ) ;
  assign n4332 = ( n4323 & n4330 ) | ( n4323 & ~n4331 ) | ( n4330 & ~n4331 ) ;
  assign n4333 = ( n4322 & ~n4331 ) | ( n4322 & n4332 ) | ( ~n4331 & n4332 ) ;
  assign n4334 = n4319 & n4321 ;
  assign n4335 = n4331 & n4333 ;
  assign n4336 = n4314 & ~n4317 ;
  assign n4337 = ~n4314 & n4317 ;
  assign n4338 = n4336 | n4337 ;
  assign n4339 = n4326 & ~n4329 ;
  assign n4340 = ~n4326 & n4329 ;
  assign n4341 = n4339 | n4340 ;
  assign n4342 = n4338 & n4341 ;
  assign n4343 = ~n4335 & n4342 ;
  assign n4344 = ~n4334 & n4343 ;
  assign n4345 = ~n4333 & n4344 ;
  assign n4346 = ( n4321 & n4333 ) | ( n4321 & n4345 ) | ( n4333 & n4345 ) ;
  assign n4347 = n4333 & n4343 ;
  assign n4348 = ~n4334 & n4347 ;
  assign n4349 = ~n4319 & n4331 ;
  assign n4350 = n4319 & ~n4331 ;
  assign n4351 = n4349 | n4350 ;
  assign n4352 = n4348 | n4351 ;
  assign n4353 = n4346 | n4352 ;
  assign n4354 = n4346 | n4348 ;
  assign n4355 = n4351 & n4354 ;
  assign n4356 = n4353 & ~n4355 ;
  assign n4357 = ( x886 & x887 ) | ( x886 & x888 ) | ( x887 & x888 ) ;
  assign n4358 = ( x883 & x884 ) | ( x883 & x885 ) | ( x884 & x885 ) ;
  assign n4359 = ( x883 & ~x884 ) | ( x883 & x885 ) | ( ~x884 & x885 ) ;
  assign n4360 = ( ~x883 & x884 ) | ( ~x883 & n4359 ) | ( x884 & n4359 ) ;
  assign n4361 = ( ~x885 & n4359 ) | ( ~x885 & n4360 ) | ( n4359 & n4360 ) ;
  assign n4362 = ( x886 & ~x887 ) | ( x886 & x888 ) | ( ~x887 & x888 ) ;
  assign n4363 = ( ~x886 & x887 ) | ( ~x886 & n4362 ) | ( x887 & n4362 ) ;
  assign n4364 = ( ~x888 & n4362 ) | ( ~x888 & n4363 ) | ( n4362 & n4363 ) ;
  assign n4365 = n4361 & n4364 ;
  assign n4366 = ( n4357 & n4358 ) | ( n4357 & n4365 ) | ( n4358 & n4365 ) ;
  assign n4367 = ( n4358 & n4365 ) | ( n4358 & ~n4366 ) | ( n4365 & ~n4366 ) ;
  assign n4368 = ( n4357 & ~n4366 ) | ( n4357 & n4367 ) | ( ~n4366 & n4367 ) ;
  assign n4369 = ( x892 & x893 ) | ( x892 & x894 ) | ( x893 & x894 ) ;
  assign n4370 = ( x889 & x890 ) | ( x889 & x891 ) | ( x890 & x891 ) ;
  assign n4371 = ( x889 & ~x890 ) | ( x889 & x891 ) | ( ~x890 & x891 ) ;
  assign n4372 = ( ~x889 & x890 ) | ( ~x889 & n4371 ) | ( x890 & n4371 ) ;
  assign n4373 = ( ~x891 & n4371 ) | ( ~x891 & n4372 ) | ( n4371 & n4372 ) ;
  assign n4374 = ( x892 & ~x893 ) | ( x892 & x894 ) | ( ~x893 & x894 ) ;
  assign n4375 = ( ~x892 & x893 ) | ( ~x892 & n4374 ) | ( x893 & n4374 ) ;
  assign n4376 = ( ~x894 & n4374 ) | ( ~x894 & n4375 ) | ( n4374 & n4375 ) ;
  assign n4377 = n4373 & n4376 ;
  assign n4378 = ( n4369 & n4370 ) | ( n4369 & n4377 ) | ( n4370 & n4377 ) ;
  assign n4379 = ( n4370 & n4377 ) | ( n4370 & ~n4378 ) | ( n4377 & ~n4378 ) ;
  assign n4380 = ( n4369 & ~n4378 ) | ( n4369 & n4379 ) | ( ~n4378 & n4379 ) ;
  assign n4381 = n4366 & n4368 ;
  assign n4382 = n4361 & ~n4364 ;
  assign n4383 = ~n4361 & n4364 ;
  assign n4384 = n4382 | n4383 ;
  assign n4385 = n4373 & ~n4376 ;
  assign n4386 = ~n4373 & n4376 ;
  assign n4387 = n4385 | n4386 ;
  assign n4388 = n4384 & n4387 ;
  assign n4389 = ~n4381 & n4388 ;
  assign n4390 = ( n4368 & n4380 ) | ( n4368 & n4389 ) | ( n4380 & n4389 ) ;
  assign n4391 = ~n4366 & n4378 ;
  assign n4392 = n4366 & ~n4378 ;
  assign n4393 = n4391 | n4392 ;
  assign n4394 = n4390 & n4393 ;
  assign n4395 = n4390 | n4393 ;
  assign n4396 = ~n4394 & n4395 ;
  assign n4397 = n4356 | n4396 ;
  assign n4398 = ( n4321 & n4333 ) | ( n4321 & ~n4344 ) | ( n4333 & ~n4344 ) ;
  assign n4399 = n4321 & ~n4348 ;
  assign n4400 = ( n4333 & ~n4398 ) | ( n4333 & n4399 ) | ( ~n4398 & n4399 ) ;
  assign n4401 = ( n4345 & n4398 ) | ( n4345 & ~n4400 ) | ( n4398 & ~n4400 ) ;
  assign n4402 = n4384 & ~n4387 ;
  assign n4403 = ~n4384 & n4387 ;
  assign n4404 = n4402 | n4403 ;
  assign n4405 = n4338 & ~n4341 ;
  assign n4406 = ~n4338 & n4341 ;
  assign n4407 = n4405 | n4406 ;
  assign n4408 = n4404 & n4407 ;
  assign n4409 = n4380 | n4389 ;
  assign n4410 = ~n4390 & n4409 ;
  assign n4411 = n4380 & n4388 ;
  assign n4412 = ( n4368 & ~n4409 ) | ( n4368 & n4411 ) | ( ~n4409 & n4411 ) ;
  assign n4413 = n4410 | n4412 ;
  assign n4414 = n4408 | n4413 ;
  assign n4415 = ( n4408 & n4410 ) | ( n4408 & n4412 ) | ( n4410 & n4412 ) ;
  assign n4416 = ( n4401 & n4414 ) | ( n4401 & n4415 ) | ( n4414 & n4415 ) ;
  assign n4417 = n4397 & n4416 ;
  assign n4418 = n4356 & n4396 ;
  assign n4419 = ( n4366 & n4378 ) | ( n4366 & n4390 ) | ( n4378 & n4390 ) ;
  assign n4420 = ( n4319 & n4331 ) | ( n4319 & n4354 ) | ( n4331 & n4354 ) ;
  assign n4421 = ~n4419 & n4420 ;
  assign n4422 = n4419 & ~n4420 ;
  assign n4423 = n4421 | n4422 ;
  assign n4424 = n4418 | n4423 ;
  assign n4425 = n4417 | n4424 ;
  assign n4426 = n4417 | n4418 ;
  assign n4427 = n4423 & n4426 ;
  assign n4428 = n4425 & ~n4427 ;
  assign n4464 = ( x856 & x857 ) | ( x856 & x858 ) | ( x857 & x858 ) ;
  assign n4465 = ( x853 & x854 ) | ( x853 & x855 ) | ( x854 & x855 ) ;
  assign n4466 = ( x853 & ~x854 ) | ( x853 & x855 ) | ( ~x854 & x855 ) ;
  assign n4467 = ( ~x853 & x854 ) | ( ~x853 & n4466 ) | ( x854 & n4466 ) ;
  assign n4468 = ( ~x855 & n4466 ) | ( ~x855 & n4467 ) | ( n4466 & n4467 ) ;
  assign n4469 = ( x856 & ~x857 ) | ( x856 & x858 ) | ( ~x857 & x858 ) ;
  assign n4470 = ( ~x856 & x857 ) | ( ~x856 & n4469 ) | ( x857 & n4469 ) ;
  assign n4471 = ( ~x858 & n4469 ) | ( ~x858 & n4470 ) | ( n4469 & n4470 ) ;
  assign n4472 = n4468 & n4471 ;
  assign n4473 = ( n4464 & n4465 ) | ( n4464 & n4472 ) | ( n4465 & n4472 ) ;
  assign n4487 = ( n4465 & n4472 ) | ( n4465 & ~n4473 ) | ( n4472 & ~n4473 ) ;
  assign n4488 = ( n4464 & ~n4473 ) | ( n4464 & n4487 ) | ( ~n4473 & n4487 ) ;
  assign n4474 = ( x850 & x851 ) | ( x850 & x852 ) | ( x851 & x852 ) ;
  assign n4475 = ( x847 & x848 ) | ( x847 & x849 ) | ( x848 & x849 ) ;
  assign n4476 = ( x847 & ~x848 ) | ( x847 & x849 ) | ( ~x848 & x849 ) ;
  assign n4477 = ( ~x847 & x848 ) | ( ~x847 & n4476 ) | ( x848 & n4476 ) ;
  assign n4478 = ( ~x849 & n4476 ) | ( ~x849 & n4477 ) | ( n4476 & n4477 ) ;
  assign n4479 = ( x850 & ~x851 ) | ( x850 & x852 ) | ( ~x851 & x852 ) ;
  assign n4480 = ( ~x850 & x851 ) | ( ~x850 & n4479 ) | ( x851 & n4479 ) ;
  assign n4481 = ( ~x852 & n4479 ) | ( ~x852 & n4480 ) | ( n4479 & n4480 ) ;
  assign n4482 = n4478 & n4481 ;
  assign n4483 = ( n4474 & n4475 ) | ( n4474 & n4482 ) | ( n4475 & n4482 ) ;
  assign n4484 = ( n4475 & n4482 ) | ( n4475 & ~n4483 ) | ( n4482 & ~n4483 ) ;
  assign n4485 = ( n4474 & ~n4483 ) | ( n4474 & n4484 ) | ( ~n4483 & n4484 ) ;
  assign n4486 = n4483 & n4485 ;
  assign n4489 = n4473 & n4488 ;
  assign n4490 = n4468 & ~n4471 ;
  assign n4491 = ~n4468 & n4471 ;
  assign n4492 = n4490 | n4491 ;
  assign n4493 = n4478 & ~n4481 ;
  assign n4494 = ~n4478 & n4481 ;
  assign n4495 = n4493 | n4494 ;
  assign n4496 = n4492 & n4495 ;
  assign n4497 = ~n4489 & n4496 ;
  assign n4500 = ~n4486 & n4497 ;
  assign n4501 = ~n4488 & n4500 ;
  assign n4508 = ( n4485 & n4488 ) | ( n4485 & ~n4500 ) | ( n4488 & ~n4500 ) ;
  assign n4498 = n4488 & n4497 ;
  assign n4499 = ~n4486 & n4498 ;
  assign n4509 = n4485 & ~n4499 ;
  assign n4510 = ( n4488 & ~n4508 ) | ( n4488 & n4509 ) | ( ~n4508 & n4509 ) ;
  assign n4511 = ( n4501 & n4508 ) | ( n4501 & ~n4510 ) | ( n4508 & ~n4510 ) ;
  assign n4431 = ( x859 & ~x860 ) | ( x859 & x861 ) | ( ~x860 & x861 ) ;
  assign n4432 = ( ~x859 & x860 ) | ( ~x859 & n4431 ) | ( x860 & n4431 ) ;
  assign n4433 = ( ~x861 & n4431 ) | ( ~x861 & n4432 ) | ( n4431 & n4432 ) ;
  assign n4434 = ( x862 & ~x863 ) | ( x862 & x864 ) | ( ~x863 & x864 ) ;
  assign n4435 = ( ~x862 & x863 ) | ( ~x862 & n4434 ) | ( x863 & n4434 ) ;
  assign n4436 = ( ~x864 & n4434 ) | ( ~x864 & n4435 ) | ( n4434 & n4435 ) ;
  assign n4454 = n4433 & ~n4436 ;
  assign n4455 = ~n4433 & n4436 ;
  assign n4456 = n4454 | n4455 ;
  assign n4441 = ( x865 & ~x866 ) | ( x865 & x867 ) | ( ~x866 & x867 ) ;
  assign n4442 = ( ~x865 & x866 ) | ( ~x865 & n4441 ) | ( x866 & n4441 ) ;
  assign n4443 = ( ~x867 & n4441 ) | ( ~x867 & n4442 ) | ( n4441 & n4442 ) ;
  assign n4444 = ( x868 & ~x869 ) | ( x868 & x870 ) | ( ~x869 & x870 ) ;
  assign n4445 = ( ~x868 & x869 ) | ( ~x868 & n4444 ) | ( x869 & n4444 ) ;
  assign n4446 = ( ~x870 & n4444 ) | ( ~x870 & n4445 ) | ( n4444 & n4445 ) ;
  assign n4457 = n4443 & ~n4446 ;
  assign n4458 = ~n4443 & n4446 ;
  assign n4459 = n4457 | n4458 ;
  assign n4512 = n4456 & ~n4459 ;
  assign n4513 = ~n4456 & n4459 ;
  assign n4514 = n4512 | n4513 ;
  assign n4515 = ~n4492 & n4495 ;
  assign n4516 = n4492 & ~n4495 ;
  assign n4517 = n4515 | n4516 ;
  assign n4518 = n4514 & n4517 ;
  assign n4429 = ( x862 & x863 ) | ( x862 & x864 ) | ( x863 & x864 ) ;
  assign n4430 = ( x859 & x860 ) | ( x859 & x861 ) | ( x860 & x861 ) ;
  assign n4437 = n4433 & n4436 ;
  assign n4438 = ( n4429 & n4430 ) | ( n4429 & n4437 ) | ( n4430 & n4437 ) ;
  assign n4449 = ( n4430 & n4437 ) | ( n4430 & ~n4438 ) | ( n4437 & ~n4438 ) ;
  assign n4450 = ( n4429 & ~n4438 ) | ( n4429 & n4449 ) | ( ~n4438 & n4449 ) ;
  assign n4439 = ( x868 & x869 ) | ( x868 & x870 ) | ( x869 & x870 ) ;
  assign n4440 = ( x865 & x866 ) | ( x865 & x867 ) | ( x866 & x867 ) ;
  assign n4447 = n4443 & n4446 ;
  assign n4448 = ( n4439 & n4440 ) | ( n4439 & n4447 ) | ( n4440 & n4447 ) ;
  assign n4451 = ( n4440 & n4447 ) | ( n4440 & ~n4448 ) | ( n4447 & ~n4448 ) ;
  assign n4452 = ( n4439 & ~n4448 ) | ( n4439 & n4451 ) | ( ~n4448 & n4451 ) ;
  assign n4460 = n4456 & n4459 ;
  assign n4519 = n4452 & n4460 ;
  assign n4453 = n4438 & n4450 ;
  assign n4461 = ~n4453 & n4460 ;
  assign n4520 = n4452 | n4461 ;
  assign n4521 = ( n4450 & n4519 ) | ( n4450 & ~n4520 ) | ( n4519 & ~n4520 ) ;
  assign n4462 = ( n4450 & n4452 ) | ( n4450 & n4461 ) | ( n4452 & n4461 ) ;
  assign n4522 = ~n4462 & n4520 ;
  assign n4523 = n4521 | n4522 ;
  assign n4524 = n4518 | n4523 ;
  assign n4525 = n4511 & n4524 ;
  assign n4526 = ( n4518 & n4521 ) | ( n4518 & n4522 ) | ( n4521 & n4522 ) ;
  assign n4527 = n4525 | n4526 ;
  assign n4502 = ( n4485 & n4488 ) | ( n4485 & n4501 ) | ( n4488 & n4501 ) ;
  assign n4528 = n4473 & ~n4483 ;
  assign n4529 = ~n4473 & n4483 ;
  assign n4530 = n4528 | n4529 ;
  assign n4531 = n4499 | n4530 ;
  assign n4532 = n4502 | n4531 ;
  assign n4503 = n4499 | n4502 ;
  assign n4533 = n4503 & n4530 ;
  assign n4534 = n4532 & ~n4533 ;
  assign n4535 = ~n4438 & n4448 ;
  assign n4536 = n4438 & ~n4448 ;
  assign n4537 = n4535 | n4536 ;
  assign n4538 = n4462 & n4537 ;
  assign n4539 = n4462 | n4537 ;
  assign n4540 = ~n4538 & n4539 ;
  assign n4541 = ( n4527 & n4534 ) | ( n4527 & n4540 ) | ( n4534 & n4540 ) ;
  assign n4463 = ( n4438 & n4448 ) | ( n4438 & n4462 ) | ( n4448 & n4462 ) ;
  assign n4504 = ( n4473 & n4483 ) | ( n4473 & n4503 ) | ( n4483 & n4503 ) ;
  assign n4505 = n4463 & n4504 ;
  assign n4506 = n4504 & ~n4505 ;
  assign n4507 = ( n4463 & ~n4505 ) | ( n4463 & n4506 ) | ( ~n4505 & n4506 ) ;
  assign n4542 = n4507 | n4541 ;
  assign n4543 = ~n4507 & n4542 ;
  assign n4544 = ( ~n4541 & n4542 ) | ( ~n4541 & n4543 ) | ( n4542 & n4543 ) ;
  assign n4545 = n4428 | n4544 ;
  assign n4546 = ( n4527 & ~n4534 ) | ( n4527 & n4540 ) | ( ~n4534 & n4540 ) ;
  assign n4547 = ( ~n4527 & n4534 ) | ( ~n4527 & n4546 ) | ( n4534 & n4546 ) ;
  assign n4548 = ( ~n4540 & n4546 ) | ( ~n4540 & n4547 ) | ( n4546 & n4547 ) ;
  assign n4549 = ( ~n4356 & n4396 ) | ( ~n4356 & n4416 ) | ( n4396 & n4416 ) ;
  assign n4550 = ( n4356 & ~n4416 ) | ( n4356 & n4549 ) | ( ~n4416 & n4549 ) ;
  assign n4551 = ( ~n4396 & n4549 ) | ( ~n4396 & n4550 ) | ( n4549 & n4550 ) ;
  assign n4552 = n4404 & ~n4407 ;
  assign n4553 = ~n4404 & n4407 ;
  assign n4554 = n4552 | n4553 ;
  assign n4555 = n4514 & ~n4517 ;
  assign n4556 = ~n4514 & n4517 ;
  assign n4557 = n4555 | n4556 ;
  assign n4558 = n4554 & n4557 ;
  assign n4559 = ~n4408 & n4414 ;
  assign n4560 = ( ~n4413 & n4414 ) | ( ~n4413 & n4559 ) | ( n4414 & n4559 ) ;
  assign n4561 = n4401 & ~n4560 ;
  assign n4562 = ~n4401 & n4560 ;
  assign n4563 = n4561 | n4562 ;
  assign n4564 = ( n4511 & n4518 ) | ( n4511 & ~n4523 ) | ( n4518 & ~n4523 ) ;
  assign n4565 = ( ~n4511 & n4523 ) | ( ~n4511 & n4564 ) | ( n4523 & n4564 ) ;
  assign n4566 = ( ~n4518 & n4564 ) | ( ~n4518 & n4565 ) | ( n4564 & n4565 ) ;
  assign n4567 = ( n4558 & n4563 ) | ( n4558 & n4566 ) | ( n4563 & n4566 ) ;
  assign n4568 = ( n4548 & n4551 ) | ( n4548 & n4567 ) | ( n4551 & n4567 ) ;
  assign n4569 = n4545 & n4568 ;
  assign n4570 = n4428 & n4544 ;
  assign n4571 = n4569 | n4570 ;
  assign n4572 = n4505 | n4507 ;
  assign n4573 = ( n4505 & n4541 ) | ( n4505 & n4572 ) | ( n4541 & n4572 ) ;
  assign n4574 = ( n4419 & n4420 ) | ( n4419 & n4426 ) | ( n4420 & n4426 ) ;
  assign n4575 = n4573 & n4574 ;
  assign n4576 = n4574 & ~n4575 ;
  assign n4577 = ( n4573 & ~n4575 ) | ( n4573 & n4576 ) | ( ~n4575 & n4576 ) ;
  assign n4578 = ( n4572 & n4574 ) | ( n4572 & n4577 ) | ( n4574 & n4577 ) ;
  assign n4579 = ( n4571 & n4575 ) | ( n4571 & n4578 ) | ( n4575 & n4578 ) ;
  assign n4580 = ( x910 & x911 ) | ( x910 & x912 ) | ( x911 & x912 ) ;
  assign n4581 = ( x907 & x908 ) | ( x907 & x909 ) | ( x908 & x909 ) ;
  assign n4582 = ( x907 & ~x908 ) | ( x907 & x909 ) | ( ~x908 & x909 ) ;
  assign n4583 = ( ~x907 & x908 ) | ( ~x907 & n4582 ) | ( x908 & n4582 ) ;
  assign n4584 = ( ~x909 & n4582 ) | ( ~x909 & n4583 ) | ( n4582 & n4583 ) ;
  assign n4585 = ( x910 & ~x911 ) | ( x910 & x912 ) | ( ~x911 & x912 ) ;
  assign n4586 = ( ~x910 & x911 ) | ( ~x910 & n4585 ) | ( x911 & n4585 ) ;
  assign n4587 = ( ~x912 & n4585 ) | ( ~x912 & n4586 ) | ( n4585 & n4586 ) ;
  assign n4588 = n4584 & n4587 ;
  assign n4589 = ( n4580 & n4581 ) | ( n4580 & n4588 ) | ( n4581 & n4588 ) ;
  assign n4590 = ( x916 & x917 ) | ( x916 & x918 ) | ( x917 & x918 ) ;
  assign n4591 = ( x913 & x914 ) | ( x913 & x915 ) | ( x914 & x915 ) ;
  assign n4592 = ( x913 & ~x914 ) | ( x913 & x915 ) | ( ~x914 & x915 ) ;
  assign n4593 = ( ~x913 & x914 ) | ( ~x913 & n4592 ) | ( x914 & n4592 ) ;
  assign n4594 = ( ~x915 & n4592 ) | ( ~x915 & n4593 ) | ( n4592 & n4593 ) ;
  assign n4595 = ( x916 & ~x917 ) | ( x916 & x918 ) | ( ~x917 & x918 ) ;
  assign n4596 = ( ~x916 & x917 ) | ( ~x916 & n4595 ) | ( x917 & n4595 ) ;
  assign n4597 = ( ~x918 & n4595 ) | ( ~x918 & n4596 ) | ( n4595 & n4596 ) ;
  assign n4598 = n4594 & n4597 ;
  assign n4599 = ( n4590 & n4591 ) | ( n4590 & n4598 ) | ( n4591 & n4598 ) ;
  assign n4600 = ( n4581 & n4588 ) | ( n4581 & ~n4589 ) | ( n4588 & ~n4589 ) ;
  assign n4601 = ( n4580 & ~n4589 ) | ( n4580 & n4600 ) | ( ~n4589 & n4600 ) ;
  assign n4602 = ( n4591 & n4598 ) | ( n4591 & ~n4599 ) | ( n4598 & ~n4599 ) ;
  assign n4603 = ( n4590 & ~n4599 ) | ( n4590 & n4602 ) | ( ~n4599 & n4602 ) ;
  assign n4604 = n4589 & n4601 ;
  assign n4605 = n4584 & ~n4587 ;
  assign n4606 = ~n4584 & n4587 ;
  assign n4607 = n4605 | n4606 ;
  assign n4608 = n4594 & ~n4597 ;
  assign n4609 = ~n4594 & n4597 ;
  assign n4610 = n4608 | n4609 ;
  assign n4611 = n4607 & n4610 ;
  assign n4612 = ~n4604 & n4611 ;
  assign n4613 = ( n4601 & n4603 ) | ( n4601 & n4612 ) | ( n4603 & n4612 ) ;
  assign n4614 = ( n4589 & n4599 ) | ( n4589 & n4613 ) | ( n4599 & n4613 ) ;
  assign n4615 = ( x904 & x905 ) | ( x904 & x906 ) | ( x905 & x906 ) ;
  assign n4616 = ( x901 & x902 ) | ( x901 & x903 ) | ( x902 & x903 ) ;
  assign n4617 = ( x901 & ~x902 ) | ( x901 & x903 ) | ( ~x902 & x903 ) ;
  assign n4618 = ( ~x901 & x902 ) | ( ~x901 & n4617 ) | ( x902 & n4617 ) ;
  assign n4619 = ( ~x903 & n4617 ) | ( ~x903 & n4618 ) | ( n4617 & n4618 ) ;
  assign n4620 = ( x904 & ~x905 ) | ( x904 & x906 ) | ( ~x905 & x906 ) ;
  assign n4621 = ( ~x904 & x905 ) | ( ~x904 & n4620 ) | ( x905 & n4620 ) ;
  assign n4622 = ( ~x906 & n4620 ) | ( ~x906 & n4621 ) | ( n4620 & n4621 ) ;
  assign n4623 = n4619 & n4622 ;
  assign n4624 = ( n4615 & n4616 ) | ( n4615 & n4623 ) | ( n4616 & n4623 ) ;
  assign n4625 = ( x898 & x899 ) | ( x898 & x900 ) | ( x899 & x900 ) ;
  assign n4626 = ( x895 & x896 ) | ( x895 & x897 ) | ( x896 & x897 ) ;
  assign n4627 = ( x895 & ~x896 ) | ( x895 & x897 ) | ( ~x896 & x897 ) ;
  assign n4628 = ( ~x895 & x896 ) | ( ~x895 & n4627 ) | ( x896 & n4627 ) ;
  assign n4629 = ( ~x897 & n4627 ) | ( ~x897 & n4628 ) | ( n4627 & n4628 ) ;
  assign n4630 = ( x898 & ~x899 ) | ( x898 & x900 ) | ( ~x899 & x900 ) ;
  assign n4631 = ( ~x898 & x899 ) | ( ~x898 & n4630 ) | ( x899 & n4630 ) ;
  assign n4632 = ( ~x900 & n4630 ) | ( ~x900 & n4631 ) | ( n4630 & n4631 ) ;
  assign n4633 = n4629 & n4632 ;
  assign n4634 = ( n4625 & n4626 ) | ( n4625 & n4633 ) | ( n4626 & n4633 ) ;
  assign n4635 = ( n4626 & n4633 ) | ( n4626 & ~n4634 ) | ( n4633 & ~n4634 ) ;
  assign n4636 = ( n4625 & ~n4634 ) | ( n4625 & n4635 ) | ( ~n4634 & n4635 ) ;
  assign n4637 = n4634 & n4636 ;
  assign n4638 = ( n4616 & n4623 ) | ( n4616 & ~n4624 ) | ( n4623 & ~n4624 ) ;
  assign n4639 = ( n4615 & ~n4624 ) | ( n4615 & n4638 ) | ( ~n4624 & n4638 ) ;
  assign n4640 = n4624 & n4639 ;
  assign n4641 = n4619 & ~n4622 ;
  assign n4642 = ~n4619 & n4622 ;
  assign n4643 = n4641 | n4642 ;
  assign n4644 = n4629 & ~n4632 ;
  assign n4645 = ~n4629 & n4632 ;
  assign n4646 = n4644 | n4645 ;
  assign n4647 = n4643 & n4646 ;
  assign n4648 = ~n4640 & n4647 ;
  assign n4649 = n4639 & n4648 ;
  assign n4650 = ~n4637 & n4649 ;
  assign n4651 = ~n4637 & n4648 ;
  assign n4652 = ~n4639 & n4651 ;
  assign n4653 = ( n4636 & n4639 ) | ( n4636 & n4652 ) | ( n4639 & n4652 ) ;
  assign n4654 = n4650 | n4653 ;
  assign n4655 = ( n4624 & n4634 ) | ( n4624 & n4654 ) | ( n4634 & n4654 ) ;
  assign n4656 = ( n4636 & n4639 ) | ( n4636 & ~n4651 ) | ( n4639 & ~n4651 ) ;
  assign n4657 = n4636 & ~n4650 ;
  assign n4658 = ( n4639 & ~n4656 ) | ( n4639 & n4657 ) | ( ~n4656 & n4657 ) ;
  assign n4659 = ( n4652 & n4656 ) | ( n4652 & ~n4658 ) | ( n4656 & ~n4658 ) ;
  assign n4660 = n4607 & ~n4610 ;
  assign n4661 = ~n4607 & n4610 ;
  assign n4662 = n4660 | n4661 ;
  assign n4663 = ~n4643 & n4646 ;
  assign n4664 = n4643 & ~n4646 ;
  assign n4665 = n4663 | n4664 ;
  assign n4666 = n4662 & n4665 ;
  assign n4667 = n4603 & n4611 ;
  assign n4668 = n4603 | n4612 ;
  assign n4669 = ( n4601 & n4667 ) | ( n4601 & ~n4668 ) | ( n4667 & ~n4668 ) ;
  assign n4670 = ~n4613 & n4668 ;
  assign n4671 = n4669 | n4670 ;
  assign n4672 = n4666 | n4671 ;
  assign n4673 = n4659 & n4672 ;
  assign n4674 = ( n4666 & n4669 ) | ( n4666 & n4670 ) | ( n4669 & n4670 ) ;
  assign n4675 = n4673 | n4674 ;
  assign n4676 = n4624 & ~n4634 ;
  assign n4677 = ~n4624 & n4634 ;
  assign n4678 = n4676 | n4677 ;
  assign n4679 = n4650 | n4678 ;
  assign n4680 = n4653 | n4679 ;
  assign n4681 = n4654 & n4678 ;
  assign n4682 = n4680 & ~n4681 ;
  assign n4683 = ~n4589 & n4599 ;
  assign n4684 = n4589 & ~n4599 ;
  assign n4685 = n4683 | n4684 ;
  assign n4686 = n4613 & n4685 ;
  assign n4687 = n4613 | n4685 ;
  assign n4688 = ~n4686 & n4687 ;
  assign n4689 = ( n4675 & n4682 ) | ( n4675 & n4688 ) | ( n4682 & n4688 ) ;
  assign n4690 = ( n4614 & n4655 ) | ( n4614 & n4689 ) | ( n4655 & n4689 ) ;
  assign n4691 = ( x934 & x935 ) | ( x934 & x936 ) | ( x935 & x936 ) ;
  assign n4692 = ( x931 & x932 ) | ( x931 & x933 ) | ( x932 & x933 ) ;
  assign n4693 = ( x931 & ~x932 ) | ( x931 & x933 ) | ( ~x932 & x933 ) ;
  assign n4694 = ( ~x931 & x932 ) | ( ~x931 & n4693 ) | ( x932 & n4693 ) ;
  assign n4695 = ( ~x933 & n4693 ) | ( ~x933 & n4694 ) | ( n4693 & n4694 ) ;
  assign n4696 = ( x934 & ~x935 ) | ( x934 & x936 ) | ( ~x935 & x936 ) ;
  assign n4697 = ( ~x934 & x935 ) | ( ~x934 & n4696 ) | ( x935 & n4696 ) ;
  assign n4698 = ( ~x936 & n4696 ) | ( ~x936 & n4697 ) | ( n4696 & n4697 ) ;
  assign n4699 = n4695 & n4698 ;
  assign n4700 = ( n4691 & n4692 ) | ( n4691 & n4699 ) | ( n4692 & n4699 ) ;
  assign n4701 = ( x940 & x941 ) | ( x940 & x942 ) | ( x941 & x942 ) ;
  assign n4702 = ( x937 & x938 ) | ( x937 & x939 ) | ( x938 & x939 ) ;
  assign n4703 = ( x937 & ~x938 ) | ( x937 & x939 ) | ( ~x938 & x939 ) ;
  assign n4704 = ( ~x937 & x938 ) | ( ~x937 & n4703 ) | ( x938 & n4703 ) ;
  assign n4705 = ( ~x939 & n4703 ) | ( ~x939 & n4704 ) | ( n4703 & n4704 ) ;
  assign n4706 = ( x940 & ~x941 ) | ( x940 & x942 ) | ( ~x941 & x942 ) ;
  assign n4707 = ( ~x940 & x941 ) | ( ~x940 & n4706 ) | ( x941 & n4706 ) ;
  assign n4708 = ( ~x942 & n4706 ) | ( ~x942 & n4707 ) | ( n4706 & n4707 ) ;
  assign n4709 = n4705 & n4708 ;
  assign n4710 = ( n4701 & n4702 ) | ( n4701 & n4709 ) | ( n4702 & n4709 ) ;
  assign n4711 = ( n4692 & n4699 ) | ( n4692 & ~n4700 ) | ( n4699 & ~n4700 ) ;
  assign n4712 = ( n4691 & ~n4700 ) | ( n4691 & n4711 ) | ( ~n4700 & n4711 ) ;
  assign n4713 = ( n4702 & n4709 ) | ( n4702 & ~n4710 ) | ( n4709 & ~n4710 ) ;
  assign n4714 = ( n4701 & ~n4710 ) | ( n4701 & n4713 ) | ( ~n4710 & n4713 ) ;
  assign n4715 = n4700 & n4712 ;
  assign n4716 = n4695 & ~n4698 ;
  assign n4717 = ~n4695 & n4698 ;
  assign n4718 = n4716 | n4717 ;
  assign n4719 = n4705 & ~n4708 ;
  assign n4720 = ~n4705 & n4708 ;
  assign n4721 = n4719 | n4720 ;
  assign n4722 = n4718 & n4721 ;
  assign n4723 = ~n4715 & n4722 ;
  assign n4724 = ( n4712 & n4714 ) | ( n4712 & n4723 ) | ( n4714 & n4723 ) ;
  assign n4725 = ( n4700 & n4710 ) | ( n4700 & n4724 ) | ( n4710 & n4724 ) ;
  assign n4726 = ( x922 & x923 ) | ( x922 & x924 ) | ( x923 & x924 ) ;
  assign n4727 = ( x919 & x920 ) | ( x919 & x921 ) | ( x920 & x921 ) ;
  assign n4728 = ( x919 & ~x920 ) | ( x919 & x921 ) | ( ~x920 & x921 ) ;
  assign n4729 = ( ~x919 & x920 ) | ( ~x919 & n4728 ) | ( x920 & n4728 ) ;
  assign n4730 = ( ~x921 & n4728 ) | ( ~x921 & n4729 ) | ( n4728 & n4729 ) ;
  assign n4731 = ( x922 & ~x923 ) | ( x922 & x924 ) | ( ~x923 & x924 ) ;
  assign n4732 = ( ~x922 & x923 ) | ( ~x922 & n4731 ) | ( x923 & n4731 ) ;
  assign n4733 = ( ~x924 & n4731 ) | ( ~x924 & n4732 ) | ( n4731 & n4732 ) ;
  assign n4734 = n4730 & n4733 ;
  assign n4735 = ( n4726 & n4727 ) | ( n4726 & n4734 ) | ( n4727 & n4734 ) ;
  assign n4736 = ( x928 & x929 ) | ( x928 & x930 ) | ( x929 & x930 ) ;
  assign n4737 = ( x925 & x926 ) | ( x925 & x927 ) | ( x926 & x927 ) ;
  assign n4738 = ( x925 & ~x926 ) | ( x925 & x927 ) | ( ~x926 & x927 ) ;
  assign n4739 = ( ~x925 & x926 ) | ( ~x925 & n4738 ) | ( x926 & n4738 ) ;
  assign n4740 = ( ~x927 & n4738 ) | ( ~x927 & n4739 ) | ( n4738 & n4739 ) ;
  assign n4741 = ( x928 & ~x929 ) | ( x928 & x930 ) | ( ~x929 & x930 ) ;
  assign n4742 = ( ~x928 & x929 ) | ( ~x928 & n4741 ) | ( x929 & n4741 ) ;
  assign n4743 = ( ~x930 & n4741 ) | ( ~x930 & n4742 ) | ( n4741 & n4742 ) ;
  assign n4744 = n4740 & n4743 ;
  assign n4745 = ( n4736 & n4737 ) | ( n4736 & n4744 ) | ( n4737 & n4744 ) ;
  assign n4746 = ( n4727 & n4734 ) | ( n4727 & ~n4735 ) | ( n4734 & ~n4735 ) ;
  assign n4747 = ( n4726 & ~n4735 ) | ( n4726 & n4746 ) | ( ~n4735 & n4746 ) ;
  assign n4748 = ( n4737 & n4744 ) | ( n4737 & ~n4745 ) | ( n4744 & ~n4745 ) ;
  assign n4749 = ( n4736 & ~n4745 ) | ( n4736 & n4748 ) | ( ~n4745 & n4748 ) ;
  assign n4750 = n4735 & n4747 ;
  assign n4751 = n4745 & n4749 ;
  assign n4752 = n4730 & ~n4733 ;
  assign n4753 = ~n4730 & n4733 ;
  assign n4754 = n4752 | n4753 ;
  assign n4755 = n4740 & ~n4743 ;
  assign n4756 = ~n4740 & n4743 ;
  assign n4757 = n4755 | n4756 ;
  assign n4758 = n4754 & n4757 ;
  assign n4759 = ~n4751 & n4758 ;
  assign n4760 = ~n4750 & n4759 ;
  assign n4761 = ~n4749 & n4760 ;
  assign n4762 = ( n4747 & n4749 ) | ( n4747 & n4761 ) | ( n4749 & n4761 ) ;
  assign n4763 = n4749 & n4759 ;
  assign n4764 = ~n4750 & n4763 ;
  assign n4765 = n4762 | n4764 ;
  assign n4766 = ( n4735 & n4745 ) | ( n4735 & n4765 ) | ( n4745 & n4765 ) ;
  assign n4767 = ~n4735 & n4745 ;
  assign n4768 = n4735 & ~n4745 ;
  assign n4769 = n4767 | n4768 ;
  assign n4770 = n4764 | n4769 ;
  assign n4771 = n4762 | n4770 ;
  assign n4772 = n4765 & n4769 ;
  assign n4773 = n4771 & ~n4772 ;
  assign n4774 = ~n4700 & n4710 ;
  assign n4775 = n4700 & ~n4710 ;
  assign n4776 = n4774 | n4775 ;
  assign n4777 = n4724 & n4776 ;
  assign n4778 = n4724 | n4776 ;
  assign n4779 = ~n4777 & n4778 ;
  assign n4780 = n4773 | n4779 ;
  assign n4781 = ( n4747 & n4749 ) | ( n4747 & ~n4760 ) | ( n4749 & ~n4760 ) ;
  assign n4782 = n4747 & ~n4764 ;
  assign n4783 = ( n4749 & ~n4781 ) | ( n4749 & n4782 ) | ( ~n4781 & n4782 ) ;
  assign n4784 = ( n4761 & n4781 ) | ( n4761 & ~n4783 ) | ( n4781 & ~n4783 ) ;
  assign n4785 = n4718 & ~n4721 ;
  assign n4786 = ~n4718 & n4721 ;
  assign n4787 = n4785 | n4786 ;
  assign n4788 = n4754 & ~n4757 ;
  assign n4789 = ~n4754 & n4757 ;
  assign n4790 = n4788 | n4789 ;
  assign n4791 = n4787 & n4790 ;
  assign n4792 = n4714 | n4723 ;
  assign n4793 = ~n4724 & n4792 ;
  assign n4794 = n4714 & n4722 ;
  assign n4795 = ( n4712 & ~n4792 ) | ( n4712 & n4794 ) | ( ~n4792 & n4794 ) ;
  assign n4796 = n4793 | n4795 ;
  assign n4797 = n4791 | n4796 ;
  assign n4798 = ( n4791 & n4793 ) | ( n4791 & n4795 ) | ( n4793 & n4795 ) ;
  assign n4799 = ( n4784 & n4797 ) | ( n4784 & n4798 ) | ( n4797 & n4798 ) ;
  assign n4800 = n4780 & n4799 ;
  assign n4801 = n4773 & n4779 ;
  assign n4802 = n4800 | n4801 ;
  assign n4803 = ( n4725 & n4766 ) | ( n4725 & n4802 ) | ( n4766 & n4802 ) ;
  assign n4804 = n4690 & n4803 ;
  assign n4805 = ~n4725 & n4766 ;
  assign n4806 = n4725 & ~n4766 ;
  assign n4807 = n4805 | n4806 ;
  assign n4808 = n4801 | n4807 ;
  assign n4809 = n4800 | n4808 ;
  assign n4810 = n4802 & n4807 ;
  assign n4811 = n4809 & ~n4810 ;
  assign n4812 = ~n4614 & n4655 ;
  assign n4813 = n4614 & ~n4655 ;
  assign n4814 = n4812 | n4813 ;
  assign n4815 = n4689 | n4814 ;
  assign n4816 = ~n4814 & n4815 ;
  assign n4817 = ( ~n4689 & n4815 ) | ( ~n4689 & n4816 ) | ( n4815 & n4816 ) ;
  assign n4818 = n4811 | n4817 ;
  assign n4819 = ( n4675 & ~n4682 ) | ( n4675 & n4688 ) | ( ~n4682 & n4688 ) ;
  assign n4820 = ( ~n4675 & n4682 ) | ( ~n4675 & n4819 ) | ( n4682 & n4819 ) ;
  assign n4821 = ( ~n4688 & n4819 ) | ( ~n4688 & n4820 ) | ( n4819 & n4820 ) ;
  assign n4822 = ( ~n4773 & n4779 ) | ( ~n4773 & n4799 ) | ( n4779 & n4799 ) ;
  assign n4823 = ( n4773 & ~n4799 ) | ( n4773 & n4822 ) | ( ~n4799 & n4822 ) ;
  assign n4824 = ( ~n4779 & n4822 ) | ( ~n4779 & n4823 ) | ( n4822 & n4823 ) ;
  assign n4825 = n4787 & ~n4790 ;
  assign n4826 = ~n4787 & n4790 ;
  assign n4827 = n4825 | n4826 ;
  assign n4828 = n4662 & ~n4665 ;
  assign n4829 = ~n4662 & n4665 ;
  assign n4830 = n4828 | n4829 ;
  assign n4831 = n4827 & n4830 ;
  assign n4832 = ~n4791 & n4797 ;
  assign n4833 = ( ~n4796 & n4797 ) | ( ~n4796 & n4832 ) | ( n4797 & n4832 ) ;
  assign n4834 = n4784 & ~n4833 ;
  assign n4835 = ~n4784 & n4833 ;
  assign n4836 = n4834 | n4835 ;
  assign n4837 = ( n4659 & n4666 ) | ( n4659 & ~n4671 ) | ( n4666 & ~n4671 ) ;
  assign n4838 = ( ~n4659 & n4671 ) | ( ~n4659 & n4837 ) | ( n4671 & n4837 ) ;
  assign n4839 = ( ~n4666 & n4837 ) | ( ~n4666 & n4838 ) | ( n4837 & n4838 ) ;
  assign n4840 = ( n4831 & n4836 ) | ( n4831 & n4839 ) | ( n4836 & n4839 ) ;
  assign n4841 = ( n4821 & n4824 ) | ( n4821 & n4840 ) | ( n4824 & n4840 ) ;
  assign n4842 = n4818 & n4841 ;
  assign n4843 = n4811 & n4817 ;
  assign n4844 = n4842 | n4843 ;
  assign n4845 = n4803 & ~n4804 ;
  assign n4846 = ( n4690 & ~n4804 ) | ( n4690 & n4845 ) | ( ~n4804 & n4845 ) ;
  assign n4847 = n4844 & n4846 ;
  assign n4848 = ( n4803 & n4844 ) | ( n4803 & n4847 ) | ( n4844 & n4847 ) ;
  assign n4849 = n4804 | n4848 ;
  assign n4850 = n4579 & n4849 ;
  assign n4851 = n4575 | n4804 ;
  assign n4852 = n4578 | n4851 ;
  assign n4853 = ( n4571 & n4851 ) | ( n4571 & n4852 ) | ( n4851 & n4852 ) ;
  assign n4854 = n4848 | n4853 ;
  assign n4855 = n4850 | n4854 ;
  assign n4856 = n4570 | n4577 ;
  assign n4857 = n4569 | n4856 ;
  assign n4858 = n4571 & n4577 ;
  assign n4859 = n4857 & ~n4858 ;
  assign n4860 = n4843 | n4846 ;
  assign n4861 = n4842 | n4860 ;
  assign n4862 = ~n4847 & n4861 ;
  assign n4863 = ( ~n4548 & n4551 ) | ( ~n4548 & n4567 ) | ( n4551 & n4567 ) ;
  assign n4864 = ( n4548 & ~n4567 ) | ( n4548 & n4863 ) | ( ~n4567 & n4863 ) ;
  assign n4865 = ( ~n4551 & n4863 ) | ( ~n4551 & n4864 ) | ( n4863 & n4864 ) ;
  assign n4866 = ( ~n4821 & n4824 ) | ( ~n4821 & n4840 ) | ( n4824 & n4840 ) ;
  assign n4867 = ( n4821 & ~n4840 ) | ( n4821 & n4866 ) | ( ~n4840 & n4866 ) ;
  assign n4868 = ( ~n4824 & n4866 ) | ( ~n4824 & n4867 ) | ( n4866 & n4867 ) ;
  assign n4869 = n4827 & ~n4830 ;
  assign n4870 = ~n4827 & n4830 ;
  assign n4871 = n4869 | n4870 ;
  assign n4872 = n4554 & ~n4557 ;
  assign n4873 = ~n4554 & n4557 ;
  assign n4874 = n4872 | n4873 ;
  assign n4875 = n4871 & n4874 ;
  assign n4876 = ( n4831 & ~n4836 ) | ( n4831 & n4839 ) | ( ~n4836 & n4839 ) ;
  assign n4877 = ( ~n4831 & n4836 ) | ( ~n4831 & n4876 ) | ( n4836 & n4876 ) ;
  assign n4878 = ( ~n4839 & n4876 ) | ( ~n4839 & n4877 ) | ( n4876 & n4877 ) ;
  assign n4879 = ( n4558 & ~n4563 ) | ( n4558 & n4566 ) | ( ~n4563 & n4566 ) ;
  assign n4880 = ( ~n4558 & n4563 ) | ( ~n4558 & n4879 ) | ( n4563 & n4879 ) ;
  assign n4881 = ( ~n4566 & n4879 ) | ( ~n4566 & n4880 ) | ( n4879 & n4880 ) ;
  assign n4882 = ( n4875 & n4878 ) | ( n4875 & n4881 ) | ( n4878 & n4881 ) ;
  assign n4883 = ( n4865 & n4868 ) | ( n4865 & n4882 ) | ( n4868 & n4882 ) ;
  assign n4884 = ( ~n4811 & n4817 ) | ( ~n4811 & n4841 ) | ( n4817 & n4841 ) ;
  assign n4885 = ( n4811 & ~n4841 ) | ( n4811 & n4884 ) | ( ~n4841 & n4884 ) ;
  assign n4886 = ( ~n4817 & n4884 ) | ( ~n4817 & n4885 ) | ( n4884 & n4885 ) ;
  assign n4887 = ( ~n4428 & n4544 ) | ( ~n4428 & n4568 ) | ( n4544 & n4568 ) ;
  assign n4888 = ( n4428 & ~n4568 ) | ( n4428 & n4887 ) | ( ~n4568 & n4887 ) ;
  assign n4889 = ( ~n4544 & n4887 ) | ( ~n4544 & n4888 ) | ( n4887 & n4888 ) ;
  assign n4890 = ( n4883 & n4886 ) | ( n4883 & n4889 ) | ( n4886 & n4889 ) ;
  assign n4891 = ( n4859 & n4862 ) | ( n4859 & n4890 ) | ( n4862 & n4890 ) ;
  assign n4892 = ( n4850 & n4855 ) | ( n4850 & n4891 ) | ( n4855 & n4891 ) ;
  assign n4893 = ~n4260 & n4308 ;
  assign n4894 = ~n4258 & n4893 ;
  assign n4895 = ( ~n4301 & n4893 ) | ( ~n4301 & n4894 ) | ( n4893 & n4894 ) ;
  assign n4896 = ( n4309 & n4892 ) | ( n4309 & n4895 ) | ( n4892 & n4895 ) ;
  assign n4897 = n4892 | n4895 ;
  assign n4898 = n4309 | n4897 ;
  assign n4899 = ~n4896 & n4898 ;
  assign n4900 = n4295 | n4298 ;
  assign n4901 = ~n4299 & n4900 ;
  assign n4902 = ( ~n4859 & n4862 ) | ( ~n4859 & n4890 ) | ( n4862 & n4890 ) ;
  assign n4903 = ( n4859 & ~n4890 ) | ( n4859 & n4902 ) | ( ~n4890 & n4902 ) ;
  assign n4904 = ( ~n4862 & n4902 ) | ( ~n4862 & n4903 ) | ( n4902 & n4903 ) ;
  assign n4905 = ( n4883 & ~n4886 ) | ( n4883 & n4889 ) | ( ~n4886 & n4889 ) ;
  assign n4906 = ( ~n4883 & n4886 ) | ( ~n4883 & n4905 ) | ( n4886 & n4905 ) ;
  assign n4907 = ( ~n4889 & n4905 ) | ( ~n4889 & n4906 ) | ( n4905 & n4906 ) ;
  assign n4908 = ( ~n4865 & n4868 ) | ( ~n4865 & n4882 ) | ( n4868 & n4882 ) ;
  assign n4909 = ( n4865 & ~n4882 ) | ( n4865 & n4908 ) | ( ~n4882 & n4908 ) ;
  assign n4910 = ( ~n4868 & n4908 ) | ( ~n4868 & n4909 ) | ( n4908 & n4909 ) ;
  assign n4911 = n4871 & ~n4874 ;
  assign n4912 = ~n4871 & n4874 ;
  assign n4913 = n4911 | n4912 ;
  assign n4914 = n4273 | n4276 ;
  assign n4915 = ~n4276 & n4914 ;
  assign n4916 = ( ~n4273 & n4914 ) | ( ~n4273 & n4915 ) | ( n4914 & n4915 ) ;
  assign n4917 = n4913 & n4916 ;
  assign n4918 = ( n4277 & ~n4283 ) | ( n4277 & n4286 ) | ( ~n4283 & n4286 ) ;
  assign n4919 = ( ~n4277 & n4283 ) | ( ~n4277 & n4918 ) | ( n4283 & n4918 ) ;
  assign n4920 = ( ~n4286 & n4918 ) | ( ~n4286 & n4919 ) | ( n4918 & n4919 ) ;
  assign n4921 = ( n4875 & n4881 ) | ( n4875 & ~n4882 ) | ( n4881 & ~n4882 ) ;
  assign n4922 = ( n4878 & ~n4882 ) | ( n4878 & n4921 ) | ( ~n4882 & n4921 ) ;
  assign n4923 = ( n4917 & n4920 ) | ( n4917 & n4922 ) | ( n4920 & n4922 ) ;
  assign n4924 = ( n4270 & n4287 ) | ( n4270 & ~n4290 ) | ( n4287 & ~n4290 ) ;
  assign n4925 = ( ~n4270 & n4290 ) | ( ~n4270 & n4924 ) | ( n4290 & n4924 ) ;
  assign n4926 = ( ~n4287 & n4924 ) | ( ~n4287 & n4925 ) | ( n4924 & n4925 ) ;
  assign n4927 = ( n4910 & n4923 ) | ( n4910 & n4926 ) | ( n4923 & n4926 ) ;
  assign n4928 = n4267 & ~n4294 ;
  assign n4929 = ( ~n4267 & n4294 ) | ( ~n4267 & n4928 ) | ( n4294 & n4928 ) ;
  assign n4930 = n4928 | n4929 ;
  assign n4931 = ( n4291 & n4907 ) | ( n4291 & ~n4930 ) | ( n4907 & ~n4930 ) ;
  assign n4932 = ( ~n4291 & n4930 ) | ( ~n4291 & n4931 ) | ( n4930 & n4931 ) ;
  assign n4933 = ( ~n4907 & n4931 ) | ( ~n4907 & n4932 ) | ( n4931 & n4932 ) ;
  assign n4934 = n4927 & n4933 ;
  assign n4935 = n4927 | n4933 ;
  assign n4936 = ~n4934 & n4935 ;
  assign n4937 = ( n4907 & n4927 ) | ( n4907 & ~n4936 ) | ( n4927 & ~n4936 ) ;
  assign n4938 = ( n4907 & n4927 ) | ( n4907 & n4937 ) | ( n4927 & n4937 ) ;
  assign n4939 = ( n4901 & n4904 ) | ( n4901 & n4938 ) | ( n4904 & n4938 ) ;
  assign n4940 = ( n4579 & n4849 ) | ( n4579 & ~n4891 ) | ( n4849 & ~n4891 ) ;
  assign n4941 = ( ~n4849 & n4891 ) | ( ~n4849 & n4940 ) | ( n4891 & n4940 ) ;
  assign n4942 = ( ~n4579 & n4940 ) | ( ~n4579 & n4941 ) | ( n4940 & n4941 ) ;
  assign n4943 = ( n3994 & ~n4257 ) | ( n3994 & n4301 ) | ( ~n4257 & n4301 ) ;
  assign n4944 = ( ~n3994 & n4257 ) | ( ~n3994 & n4943 ) | ( n4257 & n4943 ) ;
  assign n4945 = ( ~n4301 & n4943 ) | ( ~n4301 & n4944 ) | ( n4943 & n4944 ) ;
  assign n4946 = ( n4939 & n4942 ) | ( n4939 & n4945 ) | ( n4942 & n4945 ) ;
  assign n4947 = n4899 & n4946 ;
  assign n4948 = n4302 & n4308 ;
  assign n4949 = ( n4896 & n4947 ) | ( n4896 & n4948 ) | ( n4947 & n4948 ) ;
  assign n4950 = n3485 | n4949 ;
  assign n4951 = n3482 | n4950 ;
  assign n4952 = n3482 | n3485 ;
  assign n4953 = n4949 & n4952 ;
  assign n4954 = n4899 | n4946 ;
  assign n4955 = ~n4947 & n4954 ;
  assign n4956 = ( n3424 & ~n3447 ) | ( n3424 & n3463 ) | ( ~n3447 & n3463 ) ;
  assign n4957 = ( ~n3424 & n3447 ) | ( ~n3424 & n4956 ) | ( n3447 & n4956 ) ;
  assign n4958 = ( ~n3463 & n4956 ) | ( ~n3463 & n4957 ) | ( n4956 & n4957 ) ;
  assign n4959 = ( n2190 & ~n3388 ) | ( n2190 & n3423 ) | ( ~n3388 & n3423 ) ;
  assign n4960 = ( ~n2190 & n3388 ) | ( ~n2190 & n4959 ) | ( n3388 & n4959 ) ;
  assign n4961 = ( ~n3423 & n4959 ) | ( ~n3423 & n4960 ) | ( n4959 & n4960 ) ;
  assign n4962 = ( ~n3397 & n3400 ) | ( ~n3397 & n3414 ) | ( n3400 & n3414 ) ;
  assign n4963 = ( n3397 & ~n3414 ) | ( n3397 & n4962 ) | ( ~n3414 & n4962 ) ;
  assign n4964 = ( ~n3400 & n4962 ) | ( ~n3400 & n4963 ) | ( n4962 & n4963 ) ;
  assign n4965 = n3403 & ~n3406 ;
  assign n4966 = ~n3403 & n3406 ;
  assign n4967 = n4965 | n4966 ;
  assign n4968 = n4913 | n4916 ;
  assign n4969 = ~n4913 & n4968 ;
  assign n4970 = ( ~n4916 & n4968 ) | ( ~n4916 & n4969 ) | ( n4968 & n4969 ) ;
  assign n4971 = n4967 & n4970 ;
  assign n4972 = ~n3407 & n3410 ;
  assign n4973 = n3407 & ~n3410 ;
  assign n4974 = n4972 | n4973 ;
  assign n4975 = n3413 & ~n4974 ;
  assign n4976 = ~n3413 & n4974 ;
  assign n4977 = n4975 | n4976 ;
  assign n4978 = ( n4917 & n4922 ) | ( n4917 & ~n4923 ) | ( n4922 & ~n4923 ) ;
  assign n4979 = ( n4920 & ~n4923 ) | ( n4920 & n4978 ) | ( ~n4923 & n4978 ) ;
  assign n4980 = ( n4971 & n4977 ) | ( n4971 & n4979 ) | ( n4977 & n4979 ) ;
  assign n4981 = ( ~n4910 & n4923 ) | ( ~n4910 & n4926 ) | ( n4923 & n4926 ) ;
  assign n4982 = ( n4910 & ~n4926 ) | ( n4910 & n4981 ) | ( ~n4926 & n4981 ) ;
  assign n4983 = ( ~n4923 & n4981 ) | ( ~n4923 & n4982 ) | ( n4981 & n4982 ) ;
  assign n4984 = ( n4964 & n4980 ) | ( n4964 & n4983 ) | ( n4980 & n4983 ) ;
  assign n4985 = ( n3415 & ~n3418 ) | ( n3415 & n3421 ) | ( ~n3418 & n3421 ) ;
  assign n4986 = ( ~n3415 & n3418 ) | ( ~n3415 & n4985 ) | ( n3418 & n4985 ) ;
  assign n4987 = ( ~n3421 & n4985 ) | ( ~n3421 & n4986 ) | ( n4985 & n4986 ) ;
  assign n4988 = ( n4936 & n4984 ) | ( n4936 & n4987 ) | ( n4984 & n4987 ) ;
  assign n4989 = ( n3391 & ~n3394 ) | ( n3391 & n3422 ) | ( ~n3394 & n3422 ) ;
  assign n4990 = ( ~n3391 & n3394 ) | ( ~n3391 & n4989 ) | ( n3394 & n4989 ) ;
  assign n4991 = ( ~n3422 & n4989 ) | ( ~n3422 & n4990 ) | ( n4989 & n4990 ) ;
  assign n4992 = ( n4901 & n4938 ) | ( n4901 & ~n4939 ) | ( n4938 & ~n4939 ) ;
  assign n4993 = ( n4904 & ~n4939 ) | ( n4904 & n4992 ) | ( ~n4939 & n4992 ) ;
  assign n4994 = ( n4988 & n4991 ) | ( n4988 & n4993 ) | ( n4991 & n4993 ) ;
  assign n4995 = ( n4939 & n4942 ) | ( n4939 & ~n4945 ) | ( n4942 & ~n4945 ) ;
  assign n4996 = ( ~n4942 & n4945 ) | ( ~n4942 & n4995 ) | ( n4945 & n4995 ) ;
  assign n4997 = ( ~n4939 & n4995 ) | ( ~n4939 & n4996 ) | ( n4995 & n4996 ) ;
  assign n4998 = ( n4961 & n4994 ) | ( n4961 & n4997 ) | ( n4994 & n4997 ) ;
  assign n4999 = ( n4955 & n4958 ) | ( n4955 & n4998 ) | ( n4958 & n4998 ) ;
  assign n5000 = n4896 | n4948 ;
  assign n5001 = n4898 | n5000 ;
  assign n5002 = ( n4946 & n5000 ) | ( n4946 & n5001 ) | ( n5000 & n5001 ) ;
  assign n5003 = ~n4949 & n5002 ;
  assign n5004 = n3484 & ~n3485 ;
  assign n5005 = ( n3483 & ~n3485 ) | ( n3483 & n5004 ) | ( ~n3485 & n5004 ) ;
  assign n5006 = n3467 & n5005 ;
  assign n5007 = n3466 | n5005 ;
  assign n5008 = n3465 | n5007 ;
  assign n5009 = ~n5006 & n5008 ;
  assign n5010 = ( n4999 & n5003 ) | ( n4999 & n5009 ) | ( n5003 & n5009 ) ;
  assign n5011 = ( n4951 & n4953 ) | ( n4951 & n5010 ) | ( n4953 & n5010 ) ;
  assign n5012 = ( x490 & x491 ) | ( x490 & x492 ) | ( x491 & x492 ) ;
  assign n5013 = ( x487 & x488 ) | ( x487 & x489 ) | ( x488 & x489 ) ;
  assign n5014 = ( x487 & ~x488 ) | ( x487 & x489 ) | ( ~x488 & x489 ) ;
  assign n5015 = ( ~x487 & x488 ) | ( ~x487 & n5014 ) | ( x488 & n5014 ) ;
  assign n5016 = ( ~x489 & n5014 ) | ( ~x489 & n5015 ) | ( n5014 & n5015 ) ;
  assign n5017 = ( x490 & ~x491 ) | ( x490 & x492 ) | ( ~x491 & x492 ) ;
  assign n5018 = ( ~x490 & x491 ) | ( ~x490 & n5017 ) | ( x491 & n5017 ) ;
  assign n5019 = ( ~x492 & n5017 ) | ( ~x492 & n5018 ) | ( n5017 & n5018 ) ;
  assign n5020 = n5016 & n5019 ;
  assign n5021 = ( n5012 & n5013 ) | ( n5012 & n5020 ) | ( n5013 & n5020 ) ;
  assign n5022 = ( n5013 & n5020 ) | ( n5013 & ~n5021 ) | ( n5020 & ~n5021 ) ;
  assign n5023 = ( n5012 & ~n5021 ) | ( n5012 & n5022 ) | ( ~n5021 & n5022 ) ;
  assign n5024 = ( x496 & x497 ) | ( x496 & x498 ) | ( x497 & x498 ) ;
  assign n5025 = ( x493 & x494 ) | ( x493 & x495 ) | ( x494 & x495 ) ;
  assign n5026 = ( x493 & ~x494 ) | ( x493 & x495 ) | ( ~x494 & x495 ) ;
  assign n5027 = ( ~x493 & x494 ) | ( ~x493 & n5026 ) | ( x494 & n5026 ) ;
  assign n5028 = ( ~x495 & n5026 ) | ( ~x495 & n5027 ) | ( n5026 & n5027 ) ;
  assign n5029 = ( x496 & ~x497 ) | ( x496 & x498 ) | ( ~x497 & x498 ) ;
  assign n5030 = ( ~x496 & x497 ) | ( ~x496 & n5029 ) | ( x497 & n5029 ) ;
  assign n5031 = ( ~x498 & n5029 ) | ( ~x498 & n5030 ) | ( n5029 & n5030 ) ;
  assign n5032 = n5028 & n5031 ;
  assign n5033 = ( n5024 & n5025 ) | ( n5024 & n5032 ) | ( n5025 & n5032 ) ;
  assign n5034 = ( n5025 & n5032 ) | ( n5025 & ~n5033 ) | ( n5032 & ~n5033 ) ;
  assign n5035 = ( n5024 & ~n5033 ) | ( n5024 & n5034 ) | ( ~n5033 & n5034 ) ;
  assign n5036 = n5021 & n5023 ;
  assign n5037 = n5033 & n5035 ;
  assign n5038 = n5016 & ~n5019 ;
  assign n5039 = ~n5016 & n5019 ;
  assign n5040 = n5038 | n5039 ;
  assign n5041 = n5028 & ~n5031 ;
  assign n5042 = ~n5028 & n5031 ;
  assign n5043 = n5041 | n5042 ;
  assign n5044 = n5040 & n5043 ;
  assign n5045 = ~n5037 & n5044 ;
  assign n5046 = ~n5036 & n5045 ;
  assign n5047 = ~n5035 & n5046 ;
  assign n5048 = ( n5023 & n5035 ) | ( n5023 & n5047 ) | ( n5035 & n5047 ) ;
  assign n5049 = n5035 & n5045 ;
  assign n5050 = ~n5036 & n5049 ;
  assign n5051 = ~n5021 & n5033 ;
  assign n5052 = n5021 & ~n5033 ;
  assign n5053 = n5051 | n5052 ;
  assign n5054 = n5050 | n5053 ;
  assign n5055 = n5048 | n5054 ;
  assign n5056 = n5048 | n5050 ;
  assign n5057 = n5053 & n5056 ;
  assign n5058 = n5055 & ~n5057 ;
  assign n5059 = ( x502 & x503 ) | ( x502 & x504 ) | ( x503 & x504 ) ;
  assign n5060 = ( x499 & x500 ) | ( x499 & x501 ) | ( x500 & x501 ) ;
  assign n5061 = ( x499 & ~x500 ) | ( x499 & x501 ) | ( ~x500 & x501 ) ;
  assign n5062 = ( ~x499 & x500 ) | ( ~x499 & n5061 ) | ( x500 & n5061 ) ;
  assign n5063 = ( ~x501 & n5061 ) | ( ~x501 & n5062 ) | ( n5061 & n5062 ) ;
  assign n5064 = ( x502 & ~x503 ) | ( x502 & x504 ) | ( ~x503 & x504 ) ;
  assign n5065 = ( ~x502 & x503 ) | ( ~x502 & n5064 ) | ( x503 & n5064 ) ;
  assign n5066 = ( ~x504 & n5064 ) | ( ~x504 & n5065 ) | ( n5064 & n5065 ) ;
  assign n5067 = n5063 & n5066 ;
  assign n5068 = ( n5059 & n5060 ) | ( n5059 & n5067 ) | ( n5060 & n5067 ) ;
  assign n5069 = ( n5060 & n5067 ) | ( n5060 & ~n5068 ) | ( n5067 & ~n5068 ) ;
  assign n5070 = ( n5059 & ~n5068 ) | ( n5059 & n5069 ) | ( ~n5068 & n5069 ) ;
  assign n5071 = ( x508 & x509 ) | ( x508 & x510 ) | ( x509 & x510 ) ;
  assign n5072 = ( x505 & x506 ) | ( x505 & x507 ) | ( x506 & x507 ) ;
  assign n5073 = ( x505 & ~x506 ) | ( x505 & x507 ) | ( ~x506 & x507 ) ;
  assign n5074 = ( ~x505 & x506 ) | ( ~x505 & n5073 ) | ( x506 & n5073 ) ;
  assign n5075 = ( ~x507 & n5073 ) | ( ~x507 & n5074 ) | ( n5073 & n5074 ) ;
  assign n5076 = ( x508 & ~x509 ) | ( x508 & x510 ) | ( ~x509 & x510 ) ;
  assign n5077 = ( ~x508 & x509 ) | ( ~x508 & n5076 ) | ( x509 & n5076 ) ;
  assign n5078 = ( ~x510 & n5076 ) | ( ~x510 & n5077 ) | ( n5076 & n5077 ) ;
  assign n5079 = n5075 & n5078 ;
  assign n5080 = ( n5071 & n5072 ) | ( n5071 & n5079 ) | ( n5072 & n5079 ) ;
  assign n5081 = ( n5072 & n5079 ) | ( n5072 & ~n5080 ) | ( n5079 & ~n5080 ) ;
  assign n5082 = ( n5071 & ~n5080 ) | ( n5071 & n5081 ) | ( ~n5080 & n5081 ) ;
  assign n5083 = n5068 & n5070 ;
  assign n5084 = n5063 & ~n5066 ;
  assign n5085 = ~n5063 & n5066 ;
  assign n5086 = n5084 | n5085 ;
  assign n5087 = n5075 & ~n5078 ;
  assign n5088 = ~n5075 & n5078 ;
  assign n5089 = n5087 | n5088 ;
  assign n5090 = n5086 & n5089 ;
  assign n5091 = ~n5083 & n5090 ;
  assign n5092 = ( n5070 & n5082 ) | ( n5070 & n5091 ) | ( n5082 & n5091 ) ;
  assign n5093 = ~n5068 & n5080 ;
  assign n5094 = n5068 & ~n5080 ;
  assign n5095 = n5093 | n5094 ;
  assign n5096 = n5092 & n5095 ;
  assign n5097 = n5092 | n5095 ;
  assign n5098 = ~n5096 & n5097 ;
  assign n5099 = n5058 | n5098 ;
  assign n5100 = ( n5023 & n5035 ) | ( n5023 & ~n5046 ) | ( n5035 & ~n5046 ) ;
  assign n5101 = n5023 & ~n5050 ;
  assign n5102 = ( n5035 & ~n5100 ) | ( n5035 & n5101 ) | ( ~n5100 & n5101 ) ;
  assign n5103 = ( n5047 & n5100 ) | ( n5047 & ~n5102 ) | ( n5100 & ~n5102 ) ;
  assign n5104 = n5086 & ~n5089 ;
  assign n5105 = ~n5086 & n5089 ;
  assign n5106 = n5104 | n5105 ;
  assign n5107 = n5040 & ~n5043 ;
  assign n5108 = ~n5040 & n5043 ;
  assign n5109 = n5107 | n5108 ;
  assign n5110 = n5106 & n5109 ;
  assign n5111 = n5082 | n5091 ;
  assign n5112 = ~n5092 & n5111 ;
  assign n5113 = n5082 & n5090 ;
  assign n5114 = ( n5070 & ~n5111 ) | ( n5070 & n5113 ) | ( ~n5111 & n5113 ) ;
  assign n5115 = n5112 | n5114 ;
  assign n5116 = n5110 | n5115 ;
  assign n5117 = ( n5110 & n5112 ) | ( n5110 & n5114 ) | ( n5112 & n5114 ) ;
  assign n5118 = ( n5103 & n5116 ) | ( n5103 & n5117 ) | ( n5116 & n5117 ) ;
  assign n5119 = n5099 & n5118 ;
  assign n5120 = n5058 & n5098 ;
  assign n5121 = ( n5068 & n5080 ) | ( n5068 & n5092 ) | ( n5080 & n5092 ) ;
  assign n5122 = ( n5021 & n5033 ) | ( n5021 & n5056 ) | ( n5033 & n5056 ) ;
  assign n5123 = ~n5121 & n5122 ;
  assign n5124 = n5121 & ~n5122 ;
  assign n5125 = n5123 | n5124 ;
  assign n5126 = n5120 | n5125 ;
  assign n5127 = n5119 | n5126 ;
  assign n5128 = n5119 | n5120 ;
  assign n5129 = n5125 & n5128 ;
  assign n5130 = n5127 & ~n5129 ;
  assign n5166 = ( x472 & x473 ) | ( x472 & x474 ) | ( x473 & x474 ) ;
  assign n5167 = ( x469 & x470 ) | ( x469 & x471 ) | ( x470 & x471 ) ;
  assign n5168 = ( x469 & ~x470 ) | ( x469 & x471 ) | ( ~x470 & x471 ) ;
  assign n5169 = ( ~x469 & x470 ) | ( ~x469 & n5168 ) | ( x470 & n5168 ) ;
  assign n5170 = ( ~x471 & n5168 ) | ( ~x471 & n5169 ) | ( n5168 & n5169 ) ;
  assign n5171 = ( x472 & ~x473 ) | ( x472 & x474 ) | ( ~x473 & x474 ) ;
  assign n5172 = ( ~x472 & x473 ) | ( ~x472 & n5171 ) | ( x473 & n5171 ) ;
  assign n5173 = ( ~x474 & n5171 ) | ( ~x474 & n5172 ) | ( n5171 & n5172 ) ;
  assign n5174 = n5170 & n5173 ;
  assign n5175 = ( n5166 & n5167 ) | ( n5166 & n5174 ) | ( n5167 & n5174 ) ;
  assign n5189 = ( n5167 & n5174 ) | ( n5167 & ~n5175 ) | ( n5174 & ~n5175 ) ;
  assign n5190 = ( n5166 & ~n5175 ) | ( n5166 & n5189 ) | ( ~n5175 & n5189 ) ;
  assign n5176 = ( x466 & ~x467 ) | ( x466 & x468 ) | ( ~x467 & x468 ) ;
  assign n5177 = ( ~x466 & x467 ) | ( ~x466 & n5176 ) | ( x467 & n5176 ) ;
  assign n5178 = ( ~x468 & n5176 ) | ( ~x468 & n5177 ) | ( n5176 & n5177 ) ;
  assign n5179 = ( x463 & ~x464 ) | ( x463 & x465 ) | ( ~x464 & x465 ) ;
  assign n5180 = ( ~x463 & x464 ) | ( ~x463 & n5179 ) | ( x464 & n5179 ) ;
  assign n5181 = ( ~x465 & n5179 ) | ( ~x465 & n5180 ) | ( n5179 & n5180 ) ;
  assign n5182 = n5178 & n5181 ;
  assign n5183 = ( x466 & x467 ) | ( x466 & x468 ) | ( x467 & x468 ) ;
  assign n5184 = ( x463 & x464 ) | ( x463 & x465 ) | ( x464 & x465 ) ;
  assign n5185 = ( n5182 & n5183 ) | ( n5182 & n5184 ) | ( n5183 & n5184 ) ;
  assign n5186 = ( n5182 & n5184 ) | ( n5182 & ~n5185 ) | ( n5184 & ~n5185 ) ;
  assign n5187 = ( n5183 & ~n5185 ) | ( n5183 & n5186 ) | ( ~n5185 & n5186 ) ;
  assign n5188 = n5185 & n5187 ;
  assign n5191 = n5175 & n5190 ;
  assign n5192 = n5170 & ~n5173 ;
  assign n5193 = ~n5170 & n5173 ;
  assign n5194 = n5192 | n5193 ;
  assign n5195 = n5178 & ~n5181 ;
  assign n5196 = ~n5178 & n5181 ;
  assign n5197 = n5195 | n5196 ;
  assign n5198 = n5194 & n5197 ;
  assign n5199 = ~n5191 & n5198 ;
  assign n5202 = ~n5188 & n5199 ;
  assign n5203 = ~n5190 & n5202 ;
  assign n5210 = ( n5187 & n5190 ) | ( n5187 & ~n5202 ) | ( n5190 & ~n5202 ) ;
  assign n5200 = n5190 & n5199 ;
  assign n5201 = ~n5188 & n5200 ;
  assign n5211 = n5187 & ~n5201 ;
  assign n5212 = ( n5190 & ~n5210 ) | ( n5190 & n5211 ) | ( ~n5210 & n5211 ) ;
  assign n5213 = ( n5203 & n5210 ) | ( n5203 & ~n5212 ) | ( n5210 & ~n5212 ) ;
  assign n5214 = ~n5194 & n5197 ;
  assign n5215 = n5194 & ~n5197 ;
  assign n5216 = n5214 | n5215 ;
  assign n5133 = ( x475 & ~x476 ) | ( x475 & x477 ) | ( ~x476 & x477 ) ;
  assign n5134 = ( ~x475 & x476 ) | ( ~x475 & n5133 ) | ( x476 & n5133 ) ;
  assign n5135 = ( ~x477 & n5133 ) | ( ~x477 & n5134 ) | ( n5133 & n5134 ) ;
  assign n5136 = ( x478 & ~x479 ) | ( x478 & x480 ) | ( ~x479 & x480 ) ;
  assign n5137 = ( ~x478 & x479 ) | ( ~x478 & n5136 ) | ( x479 & n5136 ) ;
  assign n5138 = ( ~x480 & n5136 ) | ( ~x480 & n5137 ) | ( n5136 & n5137 ) ;
  assign n5156 = n5135 & ~n5138 ;
  assign n5157 = ~n5135 & n5138 ;
  assign n5158 = n5156 | n5157 ;
  assign n5143 = ( x481 & ~x482 ) | ( x481 & x483 ) | ( ~x482 & x483 ) ;
  assign n5144 = ( ~x481 & x482 ) | ( ~x481 & n5143 ) | ( x482 & n5143 ) ;
  assign n5145 = ( ~x483 & n5143 ) | ( ~x483 & n5144 ) | ( n5143 & n5144 ) ;
  assign n5146 = ( x484 & ~x485 ) | ( x484 & x486 ) | ( ~x485 & x486 ) ;
  assign n5147 = ( ~x484 & x485 ) | ( ~x484 & n5146 ) | ( x485 & n5146 ) ;
  assign n5148 = ( ~x486 & n5146 ) | ( ~x486 & n5147 ) | ( n5146 & n5147 ) ;
  assign n5159 = n5145 & ~n5148 ;
  assign n5160 = ~n5145 & n5148 ;
  assign n5161 = n5159 | n5160 ;
  assign n5217 = n5158 & ~n5161 ;
  assign n5218 = ~n5158 & n5161 ;
  assign n5219 = n5217 | n5218 ;
  assign n5220 = n5216 & n5219 ;
  assign n5131 = ( x478 & x479 ) | ( x478 & x480 ) | ( x479 & x480 ) ;
  assign n5132 = ( x475 & x476 ) | ( x475 & x477 ) | ( x476 & x477 ) ;
  assign n5139 = n5135 & n5138 ;
  assign n5140 = ( n5131 & n5132 ) | ( n5131 & n5139 ) | ( n5132 & n5139 ) ;
  assign n5151 = ( n5132 & n5139 ) | ( n5132 & ~n5140 ) | ( n5139 & ~n5140 ) ;
  assign n5152 = ( n5131 & ~n5140 ) | ( n5131 & n5151 ) | ( ~n5140 & n5151 ) ;
  assign n5141 = ( x484 & x485 ) | ( x484 & x486 ) | ( x485 & x486 ) ;
  assign n5142 = ( x481 & x482 ) | ( x481 & x483 ) | ( x482 & x483 ) ;
  assign n5149 = n5145 & n5148 ;
  assign n5150 = ( n5141 & n5142 ) | ( n5141 & n5149 ) | ( n5142 & n5149 ) ;
  assign n5153 = ( n5142 & n5149 ) | ( n5142 & ~n5150 ) | ( n5149 & ~n5150 ) ;
  assign n5154 = ( n5141 & ~n5150 ) | ( n5141 & n5153 ) | ( ~n5150 & n5153 ) ;
  assign n5162 = n5158 & n5161 ;
  assign n5221 = n5154 & n5162 ;
  assign n5155 = n5140 & n5152 ;
  assign n5163 = ~n5155 & n5162 ;
  assign n5222 = n5154 | n5163 ;
  assign n5223 = ( n5152 & n5221 ) | ( n5152 & ~n5222 ) | ( n5221 & ~n5222 ) ;
  assign n5164 = ( n5152 & n5154 ) | ( n5152 & n5163 ) | ( n5154 & n5163 ) ;
  assign n5224 = ~n5164 & n5222 ;
  assign n5225 = n5223 | n5224 ;
  assign n5226 = n5220 | n5225 ;
  assign n5227 = n5213 & n5226 ;
  assign n5228 = ( n5220 & n5223 ) | ( n5220 & n5224 ) | ( n5223 & n5224 ) ;
  assign n5229 = n5227 | n5228 ;
  assign n5204 = ( n5187 & n5190 ) | ( n5187 & n5203 ) | ( n5190 & n5203 ) ;
  assign n5230 = n5175 & ~n5185 ;
  assign n5231 = ~n5175 & n5185 ;
  assign n5232 = n5230 | n5231 ;
  assign n5233 = n5201 | n5232 ;
  assign n5234 = n5204 | n5233 ;
  assign n5205 = n5201 | n5204 ;
  assign n5235 = n5205 & n5232 ;
  assign n5236 = n5234 & ~n5235 ;
  assign n5237 = ~n5140 & n5150 ;
  assign n5238 = n5140 & ~n5150 ;
  assign n5239 = n5237 | n5238 ;
  assign n5240 = n5164 & n5239 ;
  assign n5241 = n5164 | n5239 ;
  assign n5242 = ~n5240 & n5241 ;
  assign n5243 = ( n5229 & n5236 ) | ( n5229 & n5242 ) | ( n5236 & n5242 ) ;
  assign n5165 = ( n5140 & n5150 ) | ( n5140 & n5164 ) | ( n5150 & n5164 ) ;
  assign n5206 = ( n5175 & n5185 ) | ( n5175 & n5205 ) | ( n5185 & n5205 ) ;
  assign n5207 = n5165 & n5206 ;
  assign n5208 = n5206 & ~n5207 ;
  assign n5209 = ( n5165 & ~n5207 ) | ( n5165 & n5208 ) | ( ~n5207 & n5208 ) ;
  assign n5244 = n5209 | n5243 ;
  assign n5245 = ~n5209 & n5244 ;
  assign n5246 = ( ~n5243 & n5244 ) | ( ~n5243 & n5245 ) | ( n5244 & n5245 ) ;
  assign n5247 = n5130 | n5246 ;
  assign n5248 = ( n5229 & ~n5236 ) | ( n5229 & n5242 ) | ( ~n5236 & n5242 ) ;
  assign n5249 = ( ~n5229 & n5236 ) | ( ~n5229 & n5248 ) | ( n5236 & n5248 ) ;
  assign n5250 = ( ~n5242 & n5248 ) | ( ~n5242 & n5249 ) | ( n5248 & n5249 ) ;
  assign n5251 = ( ~n5058 & n5098 ) | ( ~n5058 & n5118 ) | ( n5098 & n5118 ) ;
  assign n5252 = ( n5058 & ~n5118 ) | ( n5058 & n5251 ) | ( ~n5118 & n5251 ) ;
  assign n5253 = ( ~n5098 & n5251 ) | ( ~n5098 & n5252 ) | ( n5251 & n5252 ) ;
  assign n5254 = n5216 & ~n5219 ;
  assign n5255 = ~n5216 & n5219 ;
  assign n5256 = n5254 | n5255 ;
  assign n5257 = n5106 & ~n5109 ;
  assign n5258 = ~n5106 & n5109 ;
  assign n5259 = n5257 | n5258 ;
  assign n5260 = n5256 & n5259 ;
  assign n5261 = ~n5110 & n5116 ;
  assign n5262 = ( ~n5115 & n5116 ) | ( ~n5115 & n5261 ) | ( n5116 & n5261 ) ;
  assign n5263 = n5103 & ~n5262 ;
  assign n5264 = ~n5103 & n5262 ;
  assign n5265 = n5263 | n5264 ;
  assign n5266 = ( n5213 & n5220 ) | ( n5213 & ~n5225 ) | ( n5220 & ~n5225 ) ;
  assign n5267 = ( ~n5213 & n5225 ) | ( ~n5213 & n5266 ) | ( n5225 & n5266 ) ;
  assign n5268 = ( ~n5220 & n5266 ) | ( ~n5220 & n5267 ) | ( n5266 & n5267 ) ;
  assign n5269 = ( n5260 & n5265 ) | ( n5260 & n5268 ) | ( n5265 & n5268 ) ;
  assign n5270 = ( n5250 & n5253 ) | ( n5250 & n5269 ) | ( n5253 & n5269 ) ;
  assign n5271 = n5247 & n5270 ;
  assign n5272 = n5130 & n5246 ;
  assign n5273 = n5271 | n5272 ;
  assign n5274 = n5207 | n5209 ;
  assign n5275 = ( n5207 & n5243 ) | ( n5207 & n5274 ) | ( n5243 & n5274 ) ;
  assign n5276 = ( n5121 & n5122 ) | ( n5121 & n5128 ) | ( n5122 & n5128 ) ;
  assign n5277 = n5275 & n5276 ;
  assign n5278 = n5276 & ~n5277 ;
  assign n5279 = ( n5275 & ~n5277 ) | ( n5275 & n5278 ) | ( ~n5277 & n5278 ) ;
  assign n5280 = ( n5274 & n5276 ) | ( n5274 & n5279 ) | ( n5276 & n5279 ) ;
  assign n5281 = ( n5273 & n5277 ) | ( n5273 & n5280 ) | ( n5277 & n5280 ) ;
  assign n5282 = ( x526 & x527 ) | ( x526 & x528 ) | ( x527 & x528 ) ;
  assign n5283 = ( x523 & x524 ) | ( x523 & x525 ) | ( x524 & x525 ) ;
  assign n5284 = ( x523 & ~x524 ) | ( x523 & x525 ) | ( ~x524 & x525 ) ;
  assign n5285 = ( ~x523 & x524 ) | ( ~x523 & n5284 ) | ( x524 & n5284 ) ;
  assign n5286 = ( ~x525 & n5284 ) | ( ~x525 & n5285 ) | ( n5284 & n5285 ) ;
  assign n5287 = ( x526 & ~x527 ) | ( x526 & x528 ) | ( ~x527 & x528 ) ;
  assign n5288 = ( ~x526 & x527 ) | ( ~x526 & n5287 ) | ( x527 & n5287 ) ;
  assign n5289 = ( ~x528 & n5287 ) | ( ~x528 & n5288 ) | ( n5287 & n5288 ) ;
  assign n5290 = n5286 & n5289 ;
  assign n5291 = ( n5282 & n5283 ) | ( n5282 & n5290 ) | ( n5283 & n5290 ) ;
  assign n5292 = ( x532 & x533 ) | ( x532 & x534 ) | ( x533 & x534 ) ;
  assign n5293 = ( x529 & x530 ) | ( x529 & x531 ) | ( x530 & x531 ) ;
  assign n5294 = ( x529 & ~x530 ) | ( x529 & x531 ) | ( ~x530 & x531 ) ;
  assign n5295 = ( ~x529 & x530 ) | ( ~x529 & n5294 ) | ( x530 & n5294 ) ;
  assign n5296 = ( ~x531 & n5294 ) | ( ~x531 & n5295 ) | ( n5294 & n5295 ) ;
  assign n5297 = ( x532 & ~x533 ) | ( x532 & x534 ) | ( ~x533 & x534 ) ;
  assign n5298 = ( ~x532 & x533 ) | ( ~x532 & n5297 ) | ( x533 & n5297 ) ;
  assign n5299 = ( ~x534 & n5297 ) | ( ~x534 & n5298 ) | ( n5297 & n5298 ) ;
  assign n5300 = n5296 & n5299 ;
  assign n5301 = ( n5292 & n5293 ) | ( n5292 & n5300 ) | ( n5293 & n5300 ) ;
  assign n5302 = ( n5283 & n5290 ) | ( n5283 & ~n5291 ) | ( n5290 & ~n5291 ) ;
  assign n5303 = ( n5282 & ~n5291 ) | ( n5282 & n5302 ) | ( ~n5291 & n5302 ) ;
  assign n5304 = ( n5293 & n5300 ) | ( n5293 & ~n5301 ) | ( n5300 & ~n5301 ) ;
  assign n5305 = ( n5292 & ~n5301 ) | ( n5292 & n5304 ) | ( ~n5301 & n5304 ) ;
  assign n5306 = n5291 & n5303 ;
  assign n5307 = n5286 & ~n5289 ;
  assign n5308 = ~n5286 & n5289 ;
  assign n5309 = n5307 | n5308 ;
  assign n5310 = n5296 & ~n5299 ;
  assign n5311 = ~n5296 & n5299 ;
  assign n5312 = n5310 | n5311 ;
  assign n5313 = n5309 & n5312 ;
  assign n5314 = ~n5306 & n5313 ;
  assign n5315 = ( n5303 & n5305 ) | ( n5303 & n5314 ) | ( n5305 & n5314 ) ;
  assign n5316 = ( n5291 & n5301 ) | ( n5291 & n5315 ) | ( n5301 & n5315 ) ;
  assign n5317 = ( x520 & x521 ) | ( x520 & x522 ) | ( x521 & x522 ) ;
  assign n5318 = ( x517 & x518 ) | ( x517 & x519 ) | ( x518 & x519 ) ;
  assign n5319 = ( x517 & ~x518 ) | ( x517 & x519 ) | ( ~x518 & x519 ) ;
  assign n5320 = ( ~x517 & x518 ) | ( ~x517 & n5319 ) | ( x518 & n5319 ) ;
  assign n5321 = ( ~x519 & n5319 ) | ( ~x519 & n5320 ) | ( n5319 & n5320 ) ;
  assign n5322 = ( x520 & ~x521 ) | ( x520 & x522 ) | ( ~x521 & x522 ) ;
  assign n5323 = ( ~x520 & x521 ) | ( ~x520 & n5322 ) | ( x521 & n5322 ) ;
  assign n5324 = ( ~x522 & n5322 ) | ( ~x522 & n5323 ) | ( n5322 & n5323 ) ;
  assign n5325 = n5321 & n5324 ;
  assign n5326 = ( n5317 & n5318 ) | ( n5317 & n5325 ) | ( n5318 & n5325 ) ;
  assign n5327 = ( x514 & x515 ) | ( x514 & x516 ) | ( x515 & x516 ) ;
  assign n5328 = ( x511 & x512 ) | ( x511 & x513 ) | ( x512 & x513 ) ;
  assign n5329 = ( x511 & ~x512 ) | ( x511 & x513 ) | ( ~x512 & x513 ) ;
  assign n5330 = ( ~x511 & x512 ) | ( ~x511 & n5329 ) | ( x512 & n5329 ) ;
  assign n5331 = ( ~x513 & n5329 ) | ( ~x513 & n5330 ) | ( n5329 & n5330 ) ;
  assign n5332 = ( x514 & ~x515 ) | ( x514 & x516 ) | ( ~x515 & x516 ) ;
  assign n5333 = ( ~x514 & x515 ) | ( ~x514 & n5332 ) | ( x515 & n5332 ) ;
  assign n5334 = ( ~x516 & n5332 ) | ( ~x516 & n5333 ) | ( n5332 & n5333 ) ;
  assign n5335 = n5331 & n5334 ;
  assign n5336 = ( n5327 & n5328 ) | ( n5327 & n5335 ) | ( n5328 & n5335 ) ;
  assign n5337 = ( n5328 & n5335 ) | ( n5328 & ~n5336 ) | ( n5335 & ~n5336 ) ;
  assign n5338 = ( n5327 & ~n5336 ) | ( n5327 & n5337 ) | ( ~n5336 & n5337 ) ;
  assign n5339 = n5336 & n5338 ;
  assign n5340 = ( n5318 & n5325 ) | ( n5318 & ~n5326 ) | ( n5325 & ~n5326 ) ;
  assign n5341 = ( n5317 & ~n5326 ) | ( n5317 & n5340 ) | ( ~n5326 & n5340 ) ;
  assign n5342 = n5326 & n5341 ;
  assign n5343 = n5321 & ~n5324 ;
  assign n5344 = ~n5321 & n5324 ;
  assign n5345 = n5343 | n5344 ;
  assign n5346 = n5331 & ~n5334 ;
  assign n5347 = ~n5331 & n5334 ;
  assign n5348 = n5346 | n5347 ;
  assign n5349 = n5345 & n5348 ;
  assign n5350 = ~n5342 & n5349 ;
  assign n5351 = n5341 & n5350 ;
  assign n5352 = ~n5339 & n5351 ;
  assign n5353 = ~n5339 & n5350 ;
  assign n5354 = ~n5341 & n5353 ;
  assign n5355 = ( n5338 & n5341 ) | ( n5338 & n5354 ) | ( n5341 & n5354 ) ;
  assign n5356 = n5352 | n5355 ;
  assign n5357 = ( n5326 & n5336 ) | ( n5326 & n5356 ) | ( n5336 & n5356 ) ;
  assign n5358 = ( n5338 & n5341 ) | ( n5338 & ~n5353 ) | ( n5341 & ~n5353 ) ;
  assign n5359 = n5338 & ~n5352 ;
  assign n5360 = ( n5341 & ~n5358 ) | ( n5341 & n5359 ) | ( ~n5358 & n5359 ) ;
  assign n5361 = ( n5354 & n5358 ) | ( n5354 & ~n5360 ) | ( n5358 & ~n5360 ) ;
  assign n5362 = n5309 & ~n5312 ;
  assign n5363 = ~n5309 & n5312 ;
  assign n5364 = n5362 | n5363 ;
  assign n5365 = ~n5345 & n5348 ;
  assign n5366 = n5345 & ~n5348 ;
  assign n5367 = n5365 | n5366 ;
  assign n5368 = n5364 & n5367 ;
  assign n5369 = n5305 & n5313 ;
  assign n5370 = n5305 | n5314 ;
  assign n5371 = ( n5303 & n5369 ) | ( n5303 & ~n5370 ) | ( n5369 & ~n5370 ) ;
  assign n5372 = ~n5315 & n5370 ;
  assign n5373 = n5371 | n5372 ;
  assign n5374 = n5368 | n5373 ;
  assign n5375 = n5361 & n5374 ;
  assign n5376 = ( n5368 & n5371 ) | ( n5368 & n5372 ) | ( n5371 & n5372 ) ;
  assign n5377 = n5375 | n5376 ;
  assign n5378 = n5326 & ~n5336 ;
  assign n5379 = ~n5326 & n5336 ;
  assign n5380 = n5378 | n5379 ;
  assign n5381 = n5352 | n5380 ;
  assign n5382 = n5355 | n5381 ;
  assign n5383 = n5356 & n5380 ;
  assign n5384 = n5382 & ~n5383 ;
  assign n5385 = ~n5291 & n5301 ;
  assign n5386 = n5291 & ~n5301 ;
  assign n5387 = n5385 | n5386 ;
  assign n5388 = n5315 & n5387 ;
  assign n5389 = n5315 | n5387 ;
  assign n5390 = ~n5388 & n5389 ;
  assign n5391 = ( n5377 & n5384 ) | ( n5377 & n5390 ) | ( n5384 & n5390 ) ;
  assign n5392 = ( n5316 & n5357 ) | ( n5316 & n5391 ) | ( n5357 & n5391 ) ;
  assign n5393 = ( x550 & x551 ) | ( x550 & x552 ) | ( x551 & x552 ) ;
  assign n5394 = ( x547 & x548 ) | ( x547 & x549 ) | ( x548 & x549 ) ;
  assign n5395 = ( x547 & ~x548 ) | ( x547 & x549 ) | ( ~x548 & x549 ) ;
  assign n5396 = ( ~x547 & x548 ) | ( ~x547 & n5395 ) | ( x548 & n5395 ) ;
  assign n5397 = ( ~x549 & n5395 ) | ( ~x549 & n5396 ) | ( n5395 & n5396 ) ;
  assign n5398 = ( x550 & ~x551 ) | ( x550 & x552 ) | ( ~x551 & x552 ) ;
  assign n5399 = ( ~x550 & x551 ) | ( ~x550 & n5398 ) | ( x551 & n5398 ) ;
  assign n5400 = ( ~x552 & n5398 ) | ( ~x552 & n5399 ) | ( n5398 & n5399 ) ;
  assign n5401 = n5397 & n5400 ;
  assign n5402 = ( n5393 & n5394 ) | ( n5393 & n5401 ) | ( n5394 & n5401 ) ;
  assign n5403 = ( x556 & x557 ) | ( x556 & x558 ) | ( x557 & x558 ) ;
  assign n5404 = ( x553 & x554 ) | ( x553 & x555 ) | ( x554 & x555 ) ;
  assign n5405 = ( x553 & ~x554 ) | ( x553 & x555 ) | ( ~x554 & x555 ) ;
  assign n5406 = ( ~x553 & x554 ) | ( ~x553 & n5405 ) | ( x554 & n5405 ) ;
  assign n5407 = ( ~x555 & n5405 ) | ( ~x555 & n5406 ) | ( n5405 & n5406 ) ;
  assign n5408 = ( x556 & ~x557 ) | ( x556 & x558 ) | ( ~x557 & x558 ) ;
  assign n5409 = ( ~x556 & x557 ) | ( ~x556 & n5408 ) | ( x557 & n5408 ) ;
  assign n5410 = ( ~x558 & n5408 ) | ( ~x558 & n5409 ) | ( n5408 & n5409 ) ;
  assign n5411 = n5407 & n5410 ;
  assign n5412 = ( n5403 & n5404 ) | ( n5403 & n5411 ) | ( n5404 & n5411 ) ;
  assign n5413 = ( n5394 & n5401 ) | ( n5394 & ~n5402 ) | ( n5401 & ~n5402 ) ;
  assign n5414 = ( n5393 & ~n5402 ) | ( n5393 & n5413 ) | ( ~n5402 & n5413 ) ;
  assign n5415 = ( n5404 & n5411 ) | ( n5404 & ~n5412 ) | ( n5411 & ~n5412 ) ;
  assign n5416 = ( n5403 & ~n5412 ) | ( n5403 & n5415 ) | ( ~n5412 & n5415 ) ;
  assign n5417 = n5402 & n5414 ;
  assign n5418 = n5397 & ~n5400 ;
  assign n5419 = ~n5397 & n5400 ;
  assign n5420 = n5418 | n5419 ;
  assign n5421 = n5407 & ~n5410 ;
  assign n5422 = ~n5407 & n5410 ;
  assign n5423 = n5421 | n5422 ;
  assign n5424 = n5420 & n5423 ;
  assign n5425 = ~n5417 & n5424 ;
  assign n5426 = ( n5414 & n5416 ) | ( n5414 & n5425 ) | ( n5416 & n5425 ) ;
  assign n5427 = ( n5402 & n5412 ) | ( n5402 & n5426 ) | ( n5412 & n5426 ) ;
  assign n5428 = ( x538 & x539 ) | ( x538 & x540 ) | ( x539 & x540 ) ;
  assign n5429 = ( x535 & x536 ) | ( x535 & x537 ) | ( x536 & x537 ) ;
  assign n5430 = ( x535 & ~x536 ) | ( x535 & x537 ) | ( ~x536 & x537 ) ;
  assign n5431 = ( ~x535 & x536 ) | ( ~x535 & n5430 ) | ( x536 & n5430 ) ;
  assign n5432 = ( ~x537 & n5430 ) | ( ~x537 & n5431 ) | ( n5430 & n5431 ) ;
  assign n5433 = ( x538 & ~x539 ) | ( x538 & x540 ) | ( ~x539 & x540 ) ;
  assign n5434 = ( ~x538 & x539 ) | ( ~x538 & n5433 ) | ( x539 & n5433 ) ;
  assign n5435 = ( ~x540 & n5433 ) | ( ~x540 & n5434 ) | ( n5433 & n5434 ) ;
  assign n5436 = n5432 & n5435 ;
  assign n5437 = ( n5428 & n5429 ) | ( n5428 & n5436 ) | ( n5429 & n5436 ) ;
  assign n5438 = ( x544 & x545 ) | ( x544 & x546 ) | ( x545 & x546 ) ;
  assign n5439 = ( x541 & x542 ) | ( x541 & x543 ) | ( x542 & x543 ) ;
  assign n5440 = ( x541 & ~x542 ) | ( x541 & x543 ) | ( ~x542 & x543 ) ;
  assign n5441 = ( ~x541 & x542 ) | ( ~x541 & n5440 ) | ( x542 & n5440 ) ;
  assign n5442 = ( ~x543 & n5440 ) | ( ~x543 & n5441 ) | ( n5440 & n5441 ) ;
  assign n5443 = ( x544 & ~x545 ) | ( x544 & x546 ) | ( ~x545 & x546 ) ;
  assign n5444 = ( ~x544 & x545 ) | ( ~x544 & n5443 ) | ( x545 & n5443 ) ;
  assign n5445 = ( ~x546 & n5443 ) | ( ~x546 & n5444 ) | ( n5443 & n5444 ) ;
  assign n5446 = n5442 & n5445 ;
  assign n5447 = ( n5438 & n5439 ) | ( n5438 & n5446 ) | ( n5439 & n5446 ) ;
  assign n5448 = ( n5429 & n5436 ) | ( n5429 & ~n5437 ) | ( n5436 & ~n5437 ) ;
  assign n5449 = ( n5428 & ~n5437 ) | ( n5428 & n5448 ) | ( ~n5437 & n5448 ) ;
  assign n5450 = ( n5439 & n5446 ) | ( n5439 & ~n5447 ) | ( n5446 & ~n5447 ) ;
  assign n5451 = ( n5438 & ~n5447 ) | ( n5438 & n5450 ) | ( ~n5447 & n5450 ) ;
  assign n5452 = n5437 & n5449 ;
  assign n5453 = n5447 & n5451 ;
  assign n5454 = n5432 & ~n5435 ;
  assign n5455 = ~n5432 & n5435 ;
  assign n5456 = n5454 | n5455 ;
  assign n5457 = n5442 & ~n5445 ;
  assign n5458 = ~n5442 & n5445 ;
  assign n5459 = n5457 | n5458 ;
  assign n5460 = n5456 & n5459 ;
  assign n5461 = ~n5453 & n5460 ;
  assign n5462 = ~n5452 & n5461 ;
  assign n5463 = ~n5451 & n5462 ;
  assign n5464 = ( n5449 & n5451 ) | ( n5449 & n5463 ) | ( n5451 & n5463 ) ;
  assign n5465 = n5451 & n5461 ;
  assign n5466 = ~n5452 & n5465 ;
  assign n5467 = n5464 | n5466 ;
  assign n5468 = ( n5437 & n5447 ) | ( n5437 & n5467 ) | ( n5447 & n5467 ) ;
  assign n5469 = ~n5437 & n5447 ;
  assign n5470 = n5437 & ~n5447 ;
  assign n5471 = n5469 | n5470 ;
  assign n5472 = n5466 | n5471 ;
  assign n5473 = n5464 | n5472 ;
  assign n5474 = n5467 & n5471 ;
  assign n5475 = n5473 & ~n5474 ;
  assign n5476 = ~n5402 & n5412 ;
  assign n5477 = n5402 & ~n5412 ;
  assign n5478 = n5476 | n5477 ;
  assign n5479 = n5426 & n5478 ;
  assign n5480 = n5426 | n5478 ;
  assign n5481 = ~n5479 & n5480 ;
  assign n5482 = n5475 | n5481 ;
  assign n5483 = ( n5449 & n5451 ) | ( n5449 & ~n5462 ) | ( n5451 & ~n5462 ) ;
  assign n5484 = n5449 & ~n5466 ;
  assign n5485 = ( n5451 & ~n5483 ) | ( n5451 & n5484 ) | ( ~n5483 & n5484 ) ;
  assign n5486 = ( n5463 & n5483 ) | ( n5463 & ~n5485 ) | ( n5483 & ~n5485 ) ;
  assign n5487 = n5420 & ~n5423 ;
  assign n5488 = ~n5420 & n5423 ;
  assign n5489 = n5487 | n5488 ;
  assign n5490 = n5456 & ~n5459 ;
  assign n5491 = ~n5456 & n5459 ;
  assign n5492 = n5490 | n5491 ;
  assign n5493 = n5489 & n5492 ;
  assign n5494 = n5416 | n5425 ;
  assign n5495 = ~n5426 & n5494 ;
  assign n5496 = n5416 & n5424 ;
  assign n5497 = ( n5414 & ~n5494 ) | ( n5414 & n5496 ) | ( ~n5494 & n5496 ) ;
  assign n5498 = n5495 | n5497 ;
  assign n5499 = n5493 | n5498 ;
  assign n5500 = ( n5493 & n5495 ) | ( n5493 & n5497 ) | ( n5495 & n5497 ) ;
  assign n5501 = ( n5486 & n5499 ) | ( n5486 & n5500 ) | ( n5499 & n5500 ) ;
  assign n5502 = n5482 & n5501 ;
  assign n5503 = n5475 & n5481 ;
  assign n5504 = n5502 | n5503 ;
  assign n5505 = ( n5427 & n5468 ) | ( n5427 & n5504 ) | ( n5468 & n5504 ) ;
  assign n5506 = n5392 & n5505 ;
  assign n5507 = ~n5427 & n5468 ;
  assign n5508 = n5427 & ~n5468 ;
  assign n5509 = n5507 | n5508 ;
  assign n5510 = n5503 | n5509 ;
  assign n5511 = n5502 | n5510 ;
  assign n5512 = n5504 & n5509 ;
  assign n5513 = n5511 & ~n5512 ;
  assign n5514 = ~n5316 & n5357 ;
  assign n5515 = n5316 & ~n5357 ;
  assign n5516 = n5514 | n5515 ;
  assign n5517 = n5391 | n5516 ;
  assign n5518 = ~n5516 & n5517 ;
  assign n5519 = ( ~n5391 & n5517 ) | ( ~n5391 & n5518 ) | ( n5517 & n5518 ) ;
  assign n5520 = n5513 | n5519 ;
  assign n5521 = ( n5377 & ~n5384 ) | ( n5377 & n5390 ) | ( ~n5384 & n5390 ) ;
  assign n5522 = ( ~n5377 & n5384 ) | ( ~n5377 & n5521 ) | ( n5384 & n5521 ) ;
  assign n5523 = ( ~n5390 & n5521 ) | ( ~n5390 & n5522 ) | ( n5521 & n5522 ) ;
  assign n5524 = ( ~n5475 & n5481 ) | ( ~n5475 & n5501 ) | ( n5481 & n5501 ) ;
  assign n5525 = ( n5475 & ~n5501 ) | ( n5475 & n5524 ) | ( ~n5501 & n5524 ) ;
  assign n5526 = ( ~n5481 & n5524 ) | ( ~n5481 & n5525 ) | ( n5524 & n5525 ) ;
  assign n5527 = n5489 & ~n5492 ;
  assign n5528 = ~n5489 & n5492 ;
  assign n5529 = n5527 | n5528 ;
  assign n5530 = n5364 & ~n5367 ;
  assign n5531 = ~n5364 & n5367 ;
  assign n5532 = n5530 | n5531 ;
  assign n5533 = n5529 & n5532 ;
  assign n5534 = ~n5493 & n5499 ;
  assign n5535 = ( ~n5498 & n5499 ) | ( ~n5498 & n5534 ) | ( n5499 & n5534 ) ;
  assign n5536 = n5486 & ~n5535 ;
  assign n5537 = ~n5486 & n5535 ;
  assign n5538 = n5536 | n5537 ;
  assign n5539 = ( n5361 & n5368 ) | ( n5361 & ~n5373 ) | ( n5368 & ~n5373 ) ;
  assign n5540 = ( ~n5361 & n5373 ) | ( ~n5361 & n5539 ) | ( n5373 & n5539 ) ;
  assign n5541 = ( ~n5368 & n5539 ) | ( ~n5368 & n5540 ) | ( n5539 & n5540 ) ;
  assign n5542 = ( n5533 & n5538 ) | ( n5533 & n5541 ) | ( n5538 & n5541 ) ;
  assign n5543 = ( n5523 & n5526 ) | ( n5523 & n5542 ) | ( n5526 & n5542 ) ;
  assign n5544 = n5520 & n5543 ;
  assign n5545 = n5513 & n5519 ;
  assign n5546 = n5544 | n5545 ;
  assign n5547 = n5505 & ~n5506 ;
  assign n5548 = ( n5392 & ~n5506 ) | ( n5392 & n5547 ) | ( ~n5506 & n5547 ) ;
  assign n5549 = n5546 & n5548 ;
  assign n5550 = ( n5505 & n5546 ) | ( n5505 & n5549 ) | ( n5546 & n5549 ) ;
  assign n5551 = n5506 | n5550 ;
  assign n5552 = n5281 & n5551 ;
  assign n5553 = n5277 | n5506 ;
  assign n5554 = n5280 | n5553 ;
  assign n5555 = ( n5273 & n5553 ) | ( n5273 & n5554 ) | ( n5553 & n5554 ) ;
  assign n5556 = n5550 | n5555 ;
  assign n5557 = n5272 | n5279 ;
  assign n5558 = n5271 | n5557 ;
  assign n5559 = n5273 & n5279 ;
  assign n5560 = n5558 & ~n5559 ;
  assign n5561 = n5545 | n5548 ;
  assign n5562 = n5544 | n5561 ;
  assign n5563 = ~n5549 & n5562 ;
  assign n5564 = ( ~n5250 & n5253 ) | ( ~n5250 & n5269 ) | ( n5253 & n5269 ) ;
  assign n5565 = ( n5250 & ~n5269 ) | ( n5250 & n5564 ) | ( ~n5269 & n5564 ) ;
  assign n5566 = ( ~n5253 & n5564 ) | ( ~n5253 & n5565 ) | ( n5564 & n5565 ) ;
  assign n5567 = ( ~n5523 & n5526 ) | ( ~n5523 & n5542 ) | ( n5526 & n5542 ) ;
  assign n5568 = ( n5523 & ~n5542 ) | ( n5523 & n5567 ) | ( ~n5542 & n5567 ) ;
  assign n5569 = ( ~n5526 & n5567 ) | ( ~n5526 & n5568 ) | ( n5567 & n5568 ) ;
  assign n5570 = n5256 & ~n5259 ;
  assign n5571 = ~n5256 & n5259 ;
  assign n5572 = n5570 | n5571 ;
  assign n5573 = n5529 & ~n5532 ;
  assign n5574 = ~n5529 & n5532 ;
  assign n5575 = n5573 | n5574 ;
  assign n5576 = n5572 & n5575 ;
  assign n5577 = ( n5533 & ~n5538 ) | ( n5533 & n5541 ) | ( ~n5538 & n5541 ) ;
  assign n5578 = ( ~n5533 & n5538 ) | ( ~n5533 & n5577 ) | ( n5538 & n5577 ) ;
  assign n5579 = ( ~n5541 & n5577 ) | ( ~n5541 & n5578 ) | ( n5577 & n5578 ) ;
  assign n5580 = ( n5260 & ~n5265 ) | ( n5260 & n5268 ) | ( ~n5265 & n5268 ) ;
  assign n5581 = ( ~n5260 & n5265 ) | ( ~n5260 & n5580 ) | ( n5265 & n5580 ) ;
  assign n5582 = ( ~n5268 & n5580 ) | ( ~n5268 & n5581 ) | ( n5580 & n5581 ) ;
  assign n5583 = ( n5576 & n5579 ) | ( n5576 & n5582 ) | ( n5579 & n5582 ) ;
  assign n5584 = ( n5566 & n5569 ) | ( n5566 & n5583 ) | ( n5569 & n5583 ) ;
  assign n5585 = ( ~n5513 & n5519 ) | ( ~n5513 & n5543 ) | ( n5519 & n5543 ) ;
  assign n5586 = ( n5513 & ~n5543 ) | ( n5513 & n5585 ) | ( ~n5543 & n5585 ) ;
  assign n5587 = ( ~n5519 & n5585 ) | ( ~n5519 & n5586 ) | ( n5585 & n5586 ) ;
  assign n5588 = ( ~n5130 & n5246 ) | ( ~n5130 & n5270 ) | ( n5246 & n5270 ) ;
  assign n5589 = ( n5130 & ~n5270 ) | ( n5130 & n5588 ) | ( ~n5270 & n5588 ) ;
  assign n5590 = ( ~n5246 & n5588 ) | ( ~n5246 & n5589 ) | ( n5588 & n5589 ) ;
  assign n5591 = ( n5584 & n5587 ) | ( n5584 & n5590 ) | ( n5587 & n5590 ) ;
  assign n5592 = ( n5560 & n5563 ) | ( n5560 & n5591 ) | ( n5563 & n5591 ) ;
  assign n5593 = ( n5552 & n5556 ) | ( n5552 & n5592 ) | ( n5556 & n5592 ) ;
  assign n5594 = ( x586 & x587 ) | ( x586 & x588 ) | ( x587 & x588 ) ;
  assign n5595 = ( x583 & x584 ) | ( x583 & x585 ) | ( x584 & x585 ) ;
  assign n5596 = ( x583 & ~x584 ) | ( x583 & x585 ) | ( ~x584 & x585 ) ;
  assign n5597 = ( ~x583 & x584 ) | ( ~x583 & n5596 ) | ( x584 & n5596 ) ;
  assign n5598 = ( ~x585 & n5596 ) | ( ~x585 & n5597 ) | ( n5596 & n5597 ) ;
  assign n5599 = ( x586 & ~x587 ) | ( x586 & x588 ) | ( ~x587 & x588 ) ;
  assign n5600 = ( ~x586 & x587 ) | ( ~x586 & n5599 ) | ( x587 & n5599 ) ;
  assign n5601 = ( ~x588 & n5599 ) | ( ~x588 & n5600 ) | ( n5599 & n5600 ) ;
  assign n5602 = n5598 & n5601 ;
  assign n5603 = ( n5594 & n5595 ) | ( n5594 & n5602 ) | ( n5595 & n5602 ) ;
  assign n5604 = ( n5595 & n5602 ) | ( n5595 & ~n5603 ) | ( n5602 & ~n5603 ) ;
  assign n5605 = ( n5594 & ~n5603 ) | ( n5594 & n5604 ) | ( ~n5603 & n5604 ) ;
  assign n5606 = ( x592 & x593 ) | ( x592 & x594 ) | ( x593 & x594 ) ;
  assign n5607 = ( x589 & x590 ) | ( x589 & x591 ) | ( x590 & x591 ) ;
  assign n5608 = ( x589 & ~x590 ) | ( x589 & x591 ) | ( ~x590 & x591 ) ;
  assign n5609 = ( ~x589 & x590 ) | ( ~x589 & n5608 ) | ( x590 & n5608 ) ;
  assign n5610 = ( ~x591 & n5608 ) | ( ~x591 & n5609 ) | ( n5608 & n5609 ) ;
  assign n5611 = ( x592 & ~x593 ) | ( x592 & x594 ) | ( ~x593 & x594 ) ;
  assign n5612 = ( ~x592 & x593 ) | ( ~x592 & n5611 ) | ( x593 & n5611 ) ;
  assign n5613 = ( ~x594 & n5611 ) | ( ~x594 & n5612 ) | ( n5611 & n5612 ) ;
  assign n5614 = n5610 & n5613 ;
  assign n5615 = ( n5606 & n5607 ) | ( n5606 & n5614 ) | ( n5607 & n5614 ) ;
  assign n5616 = ( n5607 & n5614 ) | ( n5607 & ~n5615 ) | ( n5614 & ~n5615 ) ;
  assign n5617 = ( n5606 & ~n5615 ) | ( n5606 & n5616 ) | ( ~n5615 & n5616 ) ;
  assign n5618 = n5603 & n5605 ;
  assign n5619 = n5615 & n5617 ;
  assign n5620 = n5598 & ~n5601 ;
  assign n5621 = ~n5598 & n5601 ;
  assign n5622 = n5620 | n5621 ;
  assign n5623 = n5610 & ~n5613 ;
  assign n5624 = ~n5610 & n5613 ;
  assign n5625 = n5623 | n5624 ;
  assign n5626 = n5622 & n5625 ;
  assign n5627 = ~n5619 & n5626 ;
  assign n5628 = ~n5618 & n5627 ;
  assign n5629 = ~n5617 & n5628 ;
  assign n5630 = ( n5605 & n5617 ) | ( n5605 & n5629 ) | ( n5617 & n5629 ) ;
  assign n5631 = n5617 & n5627 ;
  assign n5632 = ~n5618 & n5631 ;
  assign n5633 = ~n5603 & n5615 ;
  assign n5634 = n5603 & ~n5615 ;
  assign n5635 = n5633 | n5634 ;
  assign n5636 = n5632 | n5635 ;
  assign n5637 = n5630 | n5636 ;
  assign n5638 = n5630 | n5632 ;
  assign n5639 = n5635 & n5638 ;
  assign n5640 = n5637 & ~n5639 ;
  assign n5641 = ( x598 & x599 ) | ( x598 & x600 ) | ( x599 & x600 ) ;
  assign n5642 = ( x595 & x596 ) | ( x595 & x597 ) | ( x596 & x597 ) ;
  assign n5643 = ( x595 & ~x596 ) | ( x595 & x597 ) | ( ~x596 & x597 ) ;
  assign n5644 = ( ~x595 & x596 ) | ( ~x595 & n5643 ) | ( x596 & n5643 ) ;
  assign n5645 = ( ~x597 & n5643 ) | ( ~x597 & n5644 ) | ( n5643 & n5644 ) ;
  assign n5646 = ( x598 & ~x599 ) | ( x598 & x600 ) | ( ~x599 & x600 ) ;
  assign n5647 = ( ~x598 & x599 ) | ( ~x598 & n5646 ) | ( x599 & n5646 ) ;
  assign n5648 = ( ~x600 & n5646 ) | ( ~x600 & n5647 ) | ( n5646 & n5647 ) ;
  assign n5649 = n5645 & n5648 ;
  assign n5650 = ( n5641 & n5642 ) | ( n5641 & n5649 ) | ( n5642 & n5649 ) ;
  assign n5651 = ( n5642 & n5649 ) | ( n5642 & ~n5650 ) | ( n5649 & ~n5650 ) ;
  assign n5652 = ( n5641 & ~n5650 ) | ( n5641 & n5651 ) | ( ~n5650 & n5651 ) ;
  assign n5653 = ( x604 & x605 ) | ( x604 & x606 ) | ( x605 & x606 ) ;
  assign n5654 = ( x601 & x602 ) | ( x601 & x603 ) | ( x602 & x603 ) ;
  assign n5655 = ( x601 & ~x602 ) | ( x601 & x603 ) | ( ~x602 & x603 ) ;
  assign n5656 = ( ~x601 & x602 ) | ( ~x601 & n5655 ) | ( x602 & n5655 ) ;
  assign n5657 = ( ~x603 & n5655 ) | ( ~x603 & n5656 ) | ( n5655 & n5656 ) ;
  assign n5658 = ( x604 & ~x605 ) | ( x604 & x606 ) | ( ~x605 & x606 ) ;
  assign n5659 = ( ~x604 & x605 ) | ( ~x604 & n5658 ) | ( x605 & n5658 ) ;
  assign n5660 = ( ~x606 & n5658 ) | ( ~x606 & n5659 ) | ( n5658 & n5659 ) ;
  assign n5661 = n5657 & n5660 ;
  assign n5662 = ( n5653 & n5654 ) | ( n5653 & n5661 ) | ( n5654 & n5661 ) ;
  assign n5663 = ( n5654 & n5661 ) | ( n5654 & ~n5662 ) | ( n5661 & ~n5662 ) ;
  assign n5664 = ( n5653 & ~n5662 ) | ( n5653 & n5663 ) | ( ~n5662 & n5663 ) ;
  assign n5665 = n5650 & n5652 ;
  assign n5666 = n5645 & ~n5648 ;
  assign n5667 = ~n5645 & n5648 ;
  assign n5668 = n5666 | n5667 ;
  assign n5669 = n5657 & ~n5660 ;
  assign n5670 = ~n5657 & n5660 ;
  assign n5671 = n5669 | n5670 ;
  assign n5672 = n5668 & n5671 ;
  assign n5673 = ~n5665 & n5672 ;
  assign n5674 = ( n5652 & n5664 ) | ( n5652 & n5673 ) | ( n5664 & n5673 ) ;
  assign n5675 = ~n5650 & n5662 ;
  assign n5676 = n5650 & ~n5662 ;
  assign n5677 = n5675 | n5676 ;
  assign n5678 = n5674 & n5677 ;
  assign n5679 = n5674 | n5677 ;
  assign n5680 = ~n5678 & n5679 ;
  assign n5681 = n5640 | n5680 ;
  assign n5682 = ( n5605 & n5617 ) | ( n5605 & ~n5628 ) | ( n5617 & ~n5628 ) ;
  assign n5683 = n5605 & ~n5632 ;
  assign n5684 = ( n5617 & ~n5682 ) | ( n5617 & n5683 ) | ( ~n5682 & n5683 ) ;
  assign n5685 = ( n5629 & n5682 ) | ( n5629 & ~n5684 ) | ( n5682 & ~n5684 ) ;
  assign n5686 = n5668 & ~n5671 ;
  assign n5687 = ~n5668 & n5671 ;
  assign n5688 = n5686 | n5687 ;
  assign n5689 = n5622 & ~n5625 ;
  assign n5690 = ~n5622 & n5625 ;
  assign n5691 = n5689 | n5690 ;
  assign n5692 = n5688 & n5691 ;
  assign n5693 = n5664 | n5673 ;
  assign n5694 = ~n5674 & n5693 ;
  assign n5695 = n5664 & n5672 ;
  assign n5696 = ( n5652 & ~n5693 ) | ( n5652 & n5695 ) | ( ~n5693 & n5695 ) ;
  assign n5697 = n5694 | n5696 ;
  assign n5698 = n5692 | n5697 ;
  assign n5699 = ( n5692 & n5694 ) | ( n5692 & n5696 ) | ( n5694 & n5696 ) ;
  assign n5700 = ( n5685 & n5698 ) | ( n5685 & n5699 ) | ( n5698 & n5699 ) ;
  assign n5701 = n5681 & n5700 ;
  assign n5702 = n5640 & n5680 ;
  assign n5703 = ( n5650 & n5662 ) | ( n5650 & n5674 ) | ( n5662 & n5674 ) ;
  assign n5704 = ( n5603 & n5615 ) | ( n5603 & n5638 ) | ( n5615 & n5638 ) ;
  assign n5705 = ~n5703 & n5704 ;
  assign n5706 = n5703 & ~n5704 ;
  assign n5707 = n5705 | n5706 ;
  assign n5708 = n5702 | n5707 ;
  assign n5709 = n5701 | n5708 ;
  assign n5710 = n5701 | n5702 ;
  assign n5711 = n5707 & n5710 ;
  assign n5712 = n5709 & ~n5711 ;
  assign n5748 = ( x568 & x569 ) | ( x568 & x570 ) | ( x569 & x570 ) ;
  assign n5749 = ( x565 & x566 ) | ( x565 & x567 ) | ( x566 & x567 ) ;
  assign n5750 = ( x565 & ~x566 ) | ( x565 & x567 ) | ( ~x566 & x567 ) ;
  assign n5751 = ( ~x565 & x566 ) | ( ~x565 & n5750 ) | ( x566 & n5750 ) ;
  assign n5752 = ( ~x567 & n5750 ) | ( ~x567 & n5751 ) | ( n5750 & n5751 ) ;
  assign n5753 = ( x568 & ~x569 ) | ( x568 & x570 ) | ( ~x569 & x570 ) ;
  assign n5754 = ( ~x568 & x569 ) | ( ~x568 & n5753 ) | ( x569 & n5753 ) ;
  assign n5755 = ( ~x570 & n5753 ) | ( ~x570 & n5754 ) | ( n5753 & n5754 ) ;
  assign n5756 = n5752 & n5755 ;
  assign n5757 = ( n5748 & n5749 ) | ( n5748 & n5756 ) | ( n5749 & n5756 ) ;
  assign n5771 = ( n5749 & n5756 ) | ( n5749 & ~n5757 ) | ( n5756 & ~n5757 ) ;
  assign n5772 = ( n5748 & ~n5757 ) | ( n5748 & n5771 ) | ( ~n5757 & n5771 ) ;
  assign n5758 = ( x562 & x563 ) | ( x562 & x564 ) | ( x563 & x564 ) ;
  assign n5759 = ( x559 & x560 ) | ( x559 & x561 ) | ( x560 & x561 ) ;
  assign n5760 = ( x559 & ~x560 ) | ( x559 & x561 ) | ( ~x560 & x561 ) ;
  assign n5761 = ( ~x559 & x560 ) | ( ~x559 & n5760 ) | ( x560 & n5760 ) ;
  assign n5762 = ( ~x561 & n5760 ) | ( ~x561 & n5761 ) | ( n5760 & n5761 ) ;
  assign n5763 = ( x562 & ~x563 ) | ( x562 & x564 ) | ( ~x563 & x564 ) ;
  assign n5764 = ( ~x562 & x563 ) | ( ~x562 & n5763 ) | ( x563 & n5763 ) ;
  assign n5765 = ( ~x564 & n5763 ) | ( ~x564 & n5764 ) | ( n5763 & n5764 ) ;
  assign n5766 = n5762 & n5765 ;
  assign n5767 = ( n5758 & n5759 ) | ( n5758 & n5766 ) | ( n5759 & n5766 ) ;
  assign n5768 = ( n5759 & n5766 ) | ( n5759 & ~n5767 ) | ( n5766 & ~n5767 ) ;
  assign n5769 = ( n5758 & ~n5767 ) | ( n5758 & n5768 ) | ( ~n5767 & n5768 ) ;
  assign n5770 = n5767 & n5769 ;
  assign n5773 = n5757 & n5772 ;
  assign n5774 = n5752 & ~n5755 ;
  assign n5775 = ~n5752 & n5755 ;
  assign n5776 = n5774 | n5775 ;
  assign n5777 = n5762 & ~n5765 ;
  assign n5778 = ~n5762 & n5765 ;
  assign n5779 = n5777 | n5778 ;
  assign n5780 = n5776 & n5779 ;
  assign n5781 = ~n5773 & n5780 ;
  assign n5784 = ~n5770 & n5781 ;
  assign n5785 = ~n5772 & n5784 ;
  assign n5792 = ( n5769 & n5772 ) | ( n5769 & ~n5784 ) | ( n5772 & ~n5784 ) ;
  assign n5782 = n5772 & n5781 ;
  assign n5783 = ~n5770 & n5782 ;
  assign n5793 = n5769 & ~n5783 ;
  assign n5794 = ( n5772 & ~n5792 ) | ( n5772 & n5793 ) | ( ~n5792 & n5793 ) ;
  assign n5795 = ( n5785 & n5792 ) | ( n5785 & ~n5794 ) | ( n5792 & ~n5794 ) ;
  assign n5715 = ( x571 & ~x572 ) | ( x571 & x573 ) | ( ~x572 & x573 ) ;
  assign n5716 = ( ~x571 & x572 ) | ( ~x571 & n5715 ) | ( x572 & n5715 ) ;
  assign n5717 = ( ~x573 & n5715 ) | ( ~x573 & n5716 ) | ( n5715 & n5716 ) ;
  assign n5718 = ( x574 & ~x575 ) | ( x574 & x576 ) | ( ~x575 & x576 ) ;
  assign n5719 = ( ~x574 & x575 ) | ( ~x574 & n5718 ) | ( x575 & n5718 ) ;
  assign n5720 = ( ~x576 & n5718 ) | ( ~x576 & n5719 ) | ( n5718 & n5719 ) ;
  assign n5738 = n5717 & ~n5720 ;
  assign n5739 = ~n5717 & n5720 ;
  assign n5740 = n5738 | n5739 ;
  assign n5725 = ( x577 & ~x578 ) | ( x577 & x579 ) | ( ~x578 & x579 ) ;
  assign n5726 = ( ~x577 & x578 ) | ( ~x577 & n5725 ) | ( x578 & n5725 ) ;
  assign n5727 = ( ~x579 & n5725 ) | ( ~x579 & n5726 ) | ( n5725 & n5726 ) ;
  assign n5728 = ( x580 & ~x581 ) | ( x580 & x582 ) | ( ~x581 & x582 ) ;
  assign n5729 = ( ~x580 & x581 ) | ( ~x580 & n5728 ) | ( x581 & n5728 ) ;
  assign n5730 = ( ~x582 & n5728 ) | ( ~x582 & n5729 ) | ( n5728 & n5729 ) ;
  assign n5741 = n5727 & ~n5730 ;
  assign n5742 = ~n5727 & n5730 ;
  assign n5743 = n5741 | n5742 ;
  assign n5796 = n5740 & ~n5743 ;
  assign n5797 = ~n5740 & n5743 ;
  assign n5798 = n5796 | n5797 ;
  assign n5799 = ~n5776 & n5779 ;
  assign n5800 = n5776 & ~n5779 ;
  assign n5801 = n5799 | n5800 ;
  assign n5802 = n5798 & n5801 ;
  assign n5713 = ( x574 & x575 ) | ( x574 & x576 ) | ( x575 & x576 ) ;
  assign n5714 = ( x571 & x572 ) | ( x571 & x573 ) | ( x572 & x573 ) ;
  assign n5721 = n5717 & n5720 ;
  assign n5722 = ( n5713 & n5714 ) | ( n5713 & n5721 ) | ( n5714 & n5721 ) ;
  assign n5733 = ( n5714 & n5721 ) | ( n5714 & ~n5722 ) | ( n5721 & ~n5722 ) ;
  assign n5734 = ( n5713 & ~n5722 ) | ( n5713 & n5733 ) | ( ~n5722 & n5733 ) ;
  assign n5723 = ( x580 & x581 ) | ( x580 & x582 ) | ( x581 & x582 ) ;
  assign n5724 = ( x577 & x578 ) | ( x577 & x579 ) | ( x578 & x579 ) ;
  assign n5731 = n5727 & n5730 ;
  assign n5732 = ( n5723 & n5724 ) | ( n5723 & n5731 ) | ( n5724 & n5731 ) ;
  assign n5735 = ( n5724 & n5731 ) | ( n5724 & ~n5732 ) | ( n5731 & ~n5732 ) ;
  assign n5736 = ( n5723 & ~n5732 ) | ( n5723 & n5735 ) | ( ~n5732 & n5735 ) ;
  assign n5744 = n5740 & n5743 ;
  assign n5803 = n5736 & n5744 ;
  assign n5737 = n5722 & n5734 ;
  assign n5745 = ~n5737 & n5744 ;
  assign n5804 = n5736 | n5745 ;
  assign n5805 = ( n5734 & n5803 ) | ( n5734 & ~n5804 ) | ( n5803 & ~n5804 ) ;
  assign n5746 = ( n5734 & n5736 ) | ( n5734 & n5745 ) | ( n5736 & n5745 ) ;
  assign n5806 = ~n5746 & n5804 ;
  assign n5807 = n5805 | n5806 ;
  assign n5808 = n5802 | n5807 ;
  assign n5809 = n5795 & n5808 ;
  assign n5810 = ( n5802 & n5805 ) | ( n5802 & n5806 ) | ( n5805 & n5806 ) ;
  assign n5811 = n5809 | n5810 ;
  assign n5786 = ( n5769 & n5772 ) | ( n5769 & n5785 ) | ( n5772 & n5785 ) ;
  assign n5812 = n5757 & ~n5767 ;
  assign n5813 = ~n5757 & n5767 ;
  assign n5814 = n5812 | n5813 ;
  assign n5815 = n5783 | n5814 ;
  assign n5816 = n5786 | n5815 ;
  assign n5787 = n5783 | n5786 ;
  assign n5817 = n5787 & n5814 ;
  assign n5818 = n5816 & ~n5817 ;
  assign n5819 = ~n5722 & n5732 ;
  assign n5820 = n5722 & ~n5732 ;
  assign n5821 = n5819 | n5820 ;
  assign n5822 = n5746 & n5821 ;
  assign n5823 = n5746 | n5821 ;
  assign n5824 = ~n5822 & n5823 ;
  assign n5825 = ( n5811 & n5818 ) | ( n5811 & n5824 ) | ( n5818 & n5824 ) ;
  assign n5747 = ( n5722 & n5732 ) | ( n5722 & n5746 ) | ( n5732 & n5746 ) ;
  assign n5788 = ( n5757 & n5767 ) | ( n5757 & n5787 ) | ( n5767 & n5787 ) ;
  assign n5789 = n5747 & n5788 ;
  assign n5790 = n5788 & ~n5789 ;
  assign n5791 = ( n5747 & ~n5789 ) | ( n5747 & n5790 ) | ( ~n5789 & n5790 ) ;
  assign n5826 = n5791 | n5825 ;
  assign n5827 = ~n5791 & n5826 ;
  assign n5828 = ( ~n5825 & n5826 ) | ( ~n5825 & n5827 ) | ( n5826 & n5827 ) ;
  assign n5829 = n5712 | n5828 ;
  assign n5830 = ( n5811 & ~n5818 ) | ( n5811 & n5824 ) | ( ~n5818 & n5824 ) ;
  assign n5831 = ( ~n5811 & n5818 ) | ( ~n5811 & n5830 ) | ( n5818 & n5830 ) ;
  assign n5832 = ( ~n5824 & n5830 ) | ( ~n5824 & n5831 ) | ( n5830 & n5831 ) ;
  assign n5833 = ( ~n5640 & n5680 ) | ( ~n5640 & n5700 ) | ( n5680 & n5700 ) ;
  assign n5834 = ( n5640 & ~n5700 ) | ( n5640 & n5833 ) | ( ~n5700 & n5833 ) ;
  assign n5835 = ( ~n5680 & n5833 ) | ( ~n5680 & n5834 ) | ( n5833 & n5834 ) ;
  assign n5836 = n5688 & ~n5691 ;
  assign n5837 = ~n5688 & n5691 ;
  assign n5838 = n5836 | n5837 ;
  assign n5839 = n5798 & ~n5801 ;
  assign n5840 = ~n5798 & n5801 ;
  assign n5841 = n5839 | n5840 ;
  assign n5842 = n5838 & n5841 ;
  assign n5843 = ~n5692 & n5698 ;
  assign n5844 = ( ~n5697 & n5698 ) | ( ~n5697 & n5843 ) | ( n5698 & n5843 ) ;
  assign n5845 = n5685 & ~n5844 ;
  assign n5846 = ~n5685 & n5844 ;
  assign n5847 = n5845 | n5846 ;
  assign n5848 = ( n5795 & n5802 ) | ( n5795 & ~n5807 ) | ( n5802 & ~n5807 ) ;
  assign n5849 = ( ~n5795 & n5807 ) | ( ~n5795 & n5848 ) | ( n5807 & n5848 ) ;
  assign n5850 = ( ~n5802 & n5848 ) | ( ~n5802 & n5849 ) | ( n5848 & n5849 ) ;
  assign n5851 = ( n5842 & n5847 ) | ( n5842 & n5850 ) | ( n5847 & n5850 ) ;
  assign n5852 = ( n5832 & n5835 ) | ( n5832 & n5851 ) | ( n5835 & n5851 ) ;
  assign n5853 = n5829 & n5852 ;
  assign n5854 = n5712 & n5828 ;
  assign n5855 = n5853 | n5854 ;
  assign n5856 = n5789 | n5791 ;
  assign n5857 = ( n5789 & n5825 ) | ( n5789 & n5856 ) | ( n5825 & n5856 ) ;
  assign n5858 = ( n5703 & n5704 ) | ( n5703 & n5710 ) | ( n5704 & n5710 ) ;
  assign n5859 = n5857 & n5858 ;
  assign n5860 = n5858 & ~n5859 ;
  assign n5861 = ( n5857 & ~n5859 ) | ( n5857 & n5860 ) | ( ~n5859 & n5860 ) ;
  assign n5862 = ( n5856 & n5858 ) | ( n5856 & n5861 ) | ( n5858 & n5861 ) ;
  assign n5863 = ( n5855 & n5859 ) | ( n5855 & n5862 ) | ( n5859 & n5862 ) ;
  assign n5864 = ( x622 & x623 ) | ( x622 & x624 ) | ( x623 & x624 ) ;
  assign n5865 = ( x619 & x620 ) | ( x619 & x621 ) | ( x620 & x621 ) ;
  assign n5866 = ( x619 & ~x620 ) | ( x619 & x621 ) | ( ~x620 & x621 ) ;
  assign n5867 = ( ~x619 & x620 ) | ( ~x619 & n5866 ) | ( x620 & n5866 ) ;
  assign n5868 = ( ~x621 & n5866 ) | ( ~x621 & n5867 ) | ( n5866 & n5867 ) ;
  assign n5869 = ( x622 & ~x623 ) | ( x622 & x624 ) | ( ~x623 & x624 ) ;
  assign n5870 = ( ~x622 & x623 ) | ( ~x622 & n5869 ) | ( x623 & n5869 ) ;
  assign n5871 = ( ~x624 & n5869 ) | ( ~x624 & n5870 ) | ( n5869 & n5870 ) ;
  assign n5872 = n5868 & n5871 ;
  assign n5873 = ( n5864 & n5865 ) | ( n5864 & n5872 ) | ( n5865 & n5872 ) ;
  assign n5874 = ( x628 & x629 ) | ( x628 & x630 ) | ( x629 & x630 ) ;
  assign n5875 = ( x625 & x626 ) | ( x625 & x627 ) | ( x626 & x627 ) ;
  assign n5876 = ( x625 & ~x626 ) | ( x625 & x627 ) | ( ~x626 & x627 ) ;
  assign n5877 = ( ~x625 & x626 ) | ( ~x625 & n5876 ) | ( x626 & n5876 ) ;
  assign n5878 = ( ~x627 & n5876 ) | ( ~x627 & n5877 ) | ( n5876 & n5877 ) ;
  assign n5879 = ( x628 & ~x629 ) | ( x628 & x630 ) | ( ~x629 & x630 ) ;
  assign n5880 = ( ~x628 & x629 ) | ( ~x628 & n5879 ) | ( x629 & n5879 ) ;
  assign n5881 = ( ~x630 & n5879 ) | ( ~x630 & n5880 ) | ( n5879 & n5880 ) ;
  assign n5882 = n5878 & n5881 ;
  assign n5883 = ( n5874 & n5875 ) | ( n5874 & n5882 ) | ( n5875 & n5882 ) ;
  assign n5884 = ( n5865 & n5872 ) | ( n5865 & ~n5873 ) | ( n5872 & ~n5873 ) ;
  assign n5885 = ( n5864 & ~n5873 ) | ( n5864 & n5884 ) | ( ~n5873 & n5884 ) ;
  assign n5886 = ( n5875 & n5882 ) | ( n5875 & ~n5883 ) | ( n5882 & ~n5883 ) ;
  assign n5887 = ( n5874 & ~n5883 ) | ( n5874 & n5886 ) | ( ~n5883 & n5886 ) ;
  assign n5888 = n5873 & n5885 ;
  assign n5889 = n5868 & ~n5871 ;
  assign n5890 = ~n5868 & n5871 ;
  assign n5891 = n5889 | n5890 ;
  assign n5892 = n5878 & ~n5881 ;
  assign n5893 = ~n5878 & n5881 ;
  assign n5894 = n5892 | n5893 ;
  assign n5895 = n5891 & n5894 ;
  assign n5896 = ~n5888 & n5895 ;
  assign n5897 = ( n5885 & n5887 ) | ( n5885 & n5896 ) | ( n5887 & n5896 ) ;
  assign n5898 = ( n5873 & n5883 ) | ( n5873 & n5897 ) | ( n5883 & n5897 ) ;
  assign n5899 = ( x616 & x617 ) | ( x616 & x618 ) | ( x617 & x618 ) ;
  assign n5900 = ( x613 & x614 ) | ( x613 & x615 ) | ( x614 & x615 ) ;
  assign n5901 = ( x613 & ~x614 ) | ( x613 & x615 ) | ( ~x614 & x615 ) ;
  assign n5902 = ( ~x613 & x614 ) | ( ~x613 & n5901 ) | ( x614 & n5901 ) ;
  assign n5903 = ( ~x615 & n5901 ) | ( ~x615 & n5902 ) | ( n5901 & n5902 ) ;
  assign n5904 = ( x616 & ~x617 ) | ( x616 & x618 ) | ( ~x617 & x618 ) ;
  assign n5905 = ( ~x616 & x617 ) | ( ~x616 & n5904 ) | ( x617 & n5904 ) ;
  assign n5906 = ( ~x618 & n5904 ) | ( ~x618 & n5905 ) | ( n5904 & n5905 ) ;
  assign n5907 = n5903 & n5906 ;
  assign n5908 = ( n5899 & n5900 ) | ( n5899 & n5907 ) | ( n5900 & n5907 ) ;
  assign n5909 = ( x610 & x611 ) | ( x610 & x612 ) | ( x611 & x612 ) ;
  assign n5910 = ( x607 & x608 ) | ( x607 & x609 ) | ( x608 & x609 ) ;
  assign n5911 = ( x607 & ~x608 ) | ( x607 & x609 ) | ( ~x608 & x609 ) ;
  assign n5912 = ( ~x607 & x608 ) | ( ~x607 & n5911 ) | ( x608 & n5911 ) ;
  assign n5913 = ( ~x609 & n5911 ) | ( ~x609 & n5912 ) | ( n5911 & n5912 ) ;
  assign n5914 = ( x610 & ~x611 ) | ( x610 & x612 ) | ( ~x611 & x612 ) ;
  assign n5915 = ( ~x610 & x611 ) | ( ~x610 & n5914 ) | ( x611 & n5914 ) ;
  assign n5916 = ( ~x612 & n5914 ) | ( ~x612 & n5915 ) | ( n5914 & n5915 ) ;
  assign n5917 = n5913 & n5916 ;
  assign n5918 = ( n5909 & n5910 ) | ( n5909 & n5917 ) | ( n5910 & n5917 ) ;
  assign n5919 = ( n5910 & n5917 ) | ( n5910 & ~n5918 ) | ( n5917 & ~n5918 ) ;
  assign n5920 = ( n5909 & ~n5918 ) | ( n5909 & n5919 ) | ( ~n5918 & n5919 ) ;
  assign n5921 = n5918 & n5920 ;
  assign n5922 = ( n5900 & n5907 ) | ( n5900 & ~n5908 ) | ( n5907 & ~n5908 ) ;
  assign n5923 = ( n5899 & ~n5908 ) | ( n5899 & n5922 ) | ( ~n5908 & n5922 ) ;
  assign n5924 = n5908 & n5923 ;
  assign n5925 = n5903 & ~n5906 ;
  assign n5926 = ~n5903 & n5906 ;
  assign n5927 = n5925 | n5926 ;
  assign n5928 = n5913 & ~n5916 ;
  assign n5929 = ~n5913 & n5916 ;
  assign n5930 = n5928 | n5929 ;
  assign n5931 = n5927 & n5930 ;
  assign n5932 = ~n5924 & n5931 ;
  assign n5933 = n5923 & n5932 ;
  assign n5934 = ~n5921 & n5933 ;
  assign n5935 = ~n5921 & n5932 ;
  assign n5936 = ~n5923 & n5935 ;
  assign n5937 = ( n5920 & n5923 ) | ( n5920 & n5936 ) | ( n5923 & n5936 ) ;
  assign n5938 = n5934 | n5937 ;
  assign n5939 = ( n5908 & n5918 ) | ( n5908 & n5938 ) | ( n5918 & n5938 ) ;
  assign n5940 = ( n5920 & n5923 ) | ( n5920 & ~n5935 ) | ( n5923 & ~n5935 ) ;
  assign n5941 = n5920 & ~n5934 ;
  assign n5942 = ( n5923 & ~n5940 ) | ( n5923 & n5941 ) | ( ~n5940 & n5941 ) ;
  assign n5943 = ( n5936 & n5940 ) | ( n5936 & ~n5942 ) | ( n5940 & ~n5942 ) ;
  assign n5944 = n5891 & ~n5894 ;
  assign n5945 = ~n5891 & n5894 ;
  assign n5946 = n5944 | n5945 ;
  assign n5947 = ~n5927 & n5930 ;
  assign n5948 = n5927 & ~n5930 ;
  assign n5949 = n5947 | n5948 ;
  assign n5950 = n5946 & n5949 ;
  assign n5951 = n5887 & n5895 ;
  assign n5952 = n5887 | n5896 ;
  assign n5953 = ( n5885 & n5951 ) | ( n5885 & ~n5952 ) | ( n5951 & ~n5952 ) ;
  assign n5954 = ~n5897 & n5952 ;
  assign n5955 = n5953 | n5954 ;
  assign n5956 = n5950 | n5955 ;
  assign n5957 = n5943 & n5956 ;
  assign n5958 = ( n5950 & n5953 ) | ( n5950 & n5954 ) | ( n5953 & n5954 ) ;
  assign n5959 = n5957 | n5958 ;
  assign n5960 = n5908 & ~n5918 ;
  assign n5961 = ~n5908 & n5918 ;
  assign n5962 = n5960 | n5961 ;
  assign n5963 = n5934 | n5962 ;
  assign n5964 = n5937 | n5963 ;
  assign n5965 = n5938 & n5962 ;
  assign n5966 = n5964 & ~n5965 ;
  assign n5967 = ~n5873 & n5883 ;
  assign n5968 = n5873 & ~n5883 ;
  assign n5969 = n5967 | n5968 ;
  assign n5970 = n5897 & n5969 ;
  assign n5971 = n5897 | n5969 ;
  assign n5972 = ~n5970 & n5971 ;
  assign n5973 = ( n5959 & n5966 ) | ( n5959 & n5972 ) | ( n5966 & n5972 ) ;
  assign n5974 = ( n5898 & n5939 ) | ( n5898 & n5973 ) | ( n5939 & n5973 ) ;
  assign n5975 = ( x646 & x647 ) | ( x646 & x648 ) | ( x647 & x648 ) ;
  assign n5976 = ( x643 & x644 ) | ( x643 & x645 ) | ( x644 & x645 ) ;
  assign n5977 = ( x643 & ~x644 ) | ( x643 & x645 ) | ( ~x644 & x645 ) ;
  assign n5978 = ( ~x643 & x644 ) | ( ~x643 & n5977 ) | ( x644 & n5977 ) ;
  assign n5979 = ( ~x645 & n5977 ) | ( ~x645 & n5978 ) | ( n5977 & n5978 ) ;
  assign n5980 = ( x646 & ~x647 ) | ( x646 & x648 ) | ( ~x647 & x648 ) ;
  assign n5981 = ( ~x646 & x647 ) | ( ~x646 & n5980 ) | ( x647 & n5980 ) ;
  assign n5982 = ( ~x648 & n5980 ) | ( ~x648 & n5981 ) | ( n5980 & n5981 ) ;
  assign n5983 = n5979 & n5982 ;
  assign n5984 = ( n5975 & n5976 ) | ( n5975 & n5983 ) | ( n5976 & n5983 ) ;
  assign n5985 = ( x652 & x653 ) | ( x652 & x654 ) | ( x653 & x654 ) ;
  assign n5986 = ( x649 & x650 ) | ( x649 & x651 ) | ( x650 & x651 ) ;
  assign n5987 = ( x649 & ~x650 ) | ( x649 & x651 ) | ( ~x650 & x651 ) ;
  assign n5988 = ( ~x649 & x650 ) | ( ~x649 & n5987 ) | ( x650 & n5987 ) ;
  assign n5989 = ( ~x651 & n5987 ) | ( ~x651 & n5988 ) | ( n5987 & n5988 ) ;
  assign n5990 = ( x652 & ~x653 ) | ( x652 & x654 ) | ( ~x653 & x654 ) ;
  assign n5991 = ( ~x652 & x653 ) | ( ~x652 & n5990 ) | ( x653 & n5990 ) ;
  assign n5992 = ( ~x654 & n5990 ) | ( ~x654 & n5991 ) | ( n5990 & n5991 ) ;
  assign n5993 = n5989 & n5992 ;
  assign n5994 = ( n5985 & n5986 ) | ( n5985 & n5993 ) | ( n5986 & n5993 ) ;
  assign n5995 = ( n5976 & n5983 ) | ( n5976 & ~n5984 ) | ( n5983 & ~n5984 ) ;
  assign n5996 = ( n5975 & ~n5984 ) | ( n5975 & n5995 ) | ( ~n5984 & n5995 ) ;
  assign n5997 = ( n5986 & n5993 ) | ( n5986 & ~n5994 ) | ( n5993 & ~n5994 ) ;
  assign n5998 = ( n5985 & ~n5994 ) | ( n5985 & n5997 ) | ( ~n5994 & n5997 ) ;
  assign n5999 = n5984 & n5996 ;
  assign n6000 = n5979 & ~n5982 ;
  assign n6001 = ~n5979 & n5982 ;
  assign n6002 = n6000 | n6001 ;
  assign n6003 = n5989 & ~n5992 ;
  assign n6004 = ~n5989 & n5992 ;
  assign n6005 = n6003 | n6004 ;
  assign n6006 = n6002 & n6005 ;
  assign n6007 = ~n5999 & n6006 ;
  assign n6008 = ( n5996 & n5998 ) | ( n5996 & n6007 ) | ( n5998 & n6007 ) ;
  assign n6009 = ( n5984 & n5994 ) | ( n5984 & n6008 ) | ( n5994 & n6008 ) ;
  assign n6010 = ( x634 & x635 ) | ( x634 & x636 ) | ( x635 & x636 ) ;
  assign n6011 = ( x631 & x632 ) | ( x631 & x633 ) | ( x632 & x633 ) ;
  assign n6012 = ( x631 & ~x632 ) | ( x631 & x633 ) | ( ~x632 & x633 ) ;
  assign n6013 = ( ~x631 & x632 ) | ( ~x631 & n6012 ) | ( x632 & n6012 ) ;
  assign n6014 = ( ~x633 & n6012 ) | ( ~x633 & n6013 ) | ( n6012 & n6013 ) ;
  assign n6015 = ( x634 & ~x635 ) | ( x634 & x636 ) | ( ~x635 & x636 ) ;
  assign n6016 = ( ~x634 & x635 ) | ( ~x634 & n6015 ) | ( x635 & n6015 ) ;
  assign n6017 = ( ~x636 & n6015 ) | ( ~x636 & n6016 ) | ( n6015 & n6016 ) ;
  assign n6018 = n6014 & n6017 ;
  assign n6019 = ( n6010 & n6011 ) | ( n6010 & n6018 ) | ( n6011 & n6018 ) ;
  assign n6020 = ( x640 & x641 ) | ( x640 & x642 ) | ( x641 & x642 ) ;
  assign n6021 = ( x637 & x638 ) | ( x637 & x639 ) | ( x638 & x639 ) ;
  assign n6022 = ( x637 & ~x638 ) | ( x637 & x639 ) | ( ~x638 & x639 ) ;
  assign n6023 = ( ~x637 & x638 ) | ( ~x637 & n6022 ) | ( x638 & n6022 ) ;
  assign n6024 = ( ~x639 & n6022 ) | ( ~x639 & n6023 ) | ( n6022 & n6023 ) ;
  assign n6025 = ( x640 & ~x641 ) | ( x640 & x642 ) | ( ~x641 & x642 ) ;
  assign n6026 = ( ~x640 & x641 ) | ( ~x640 & n6025 ) | ( x641 & n6025 ) ;
  assign n6027 = ( ~x642 & n6025 ) | ( ~x642 & n6026 ) | ( n6025 & n6026 ) ;
  assign n6028 = n6024 & n6027 ;
  assign n6029 = ( n6020 & n6021 ) | ( n6020 & n6028 ) | ( n6021 & n6028 ) ;
  assign n6030 = ( n6011 & n6018 ) | ( n6011 & ~n6019 ) | ( n6018 & ~n6019 ) ;
  assign n6031 = ( n6010 & ~n6019 ) | ( n6010 & n6030 ) | ( ~n6019 & n6030 ) ;
  assign n6032 = ( n6021 & n6028 ) | ( n6021 & ~n6029 ) | ( n6028 & ~n6029 ) ;
  assign n6033 = ( n6020 & ~n6029 ) | ( n6020 & n6032 ) | ( ~n6029 & n6032 ) ;
  assign n6034 = n6019 & n6031 ;
  assign n6035 = n6029 & n6033 ;
  assign n6036 = n6014 & ~n6017 ;
  assign n6037 = ~n6014 & n6017 ;
  assign n6038 = n6036 | n6037 ;
  assign n6039 = n6024 & ~n6027 ;
  assign n6040 = ~n6024 & n6027 ;
  assign n6041 = n6039 | n6040 ;
  assign n6042 = n6038 & n6041 ;
  assign n6043 = ~n6035 & n6042 ;
  assign n6044 = ~n6034 & n6043 ;
  assign n6045 = ~n6033 & n6044 ;
  assign n6046 = ( n6031 & n6033 ) | ( n6031 & n6045 ) | ( n6033 & n6045 ) ;
  assign n6047 = n6033 & n6043 ;
  assign n6048 = ~n6034 & n6047 ;
  assign n6049 = n6046 | n6048 ;
  assign n6050 = ( n6019 & n6029 ) | ( n6019 & n6049 ) | ( n6029 & n6049 ) ;
  assign n6051 = ~n6019 & n6029 ;
  assign n6052 = n6019 & ~n6029 ;
  assign n6053 = n6051 | n6052 ;
  assign n6054 = n6048 | n6053 ;
  assign n6055 = n6046 | n6054 ;
  assign n6056 = n6049 & n6053 ;
  assign n6057 = n6055 & ~n6056 ;
  assign n6058 = ~n5984 & n5994 ;
  assign n6059 = n5984 & ~n5994 ;
  assign n6060 = n6058 | n6059 ;
  assign n6061 = n6008 & n6060 ;
  assign n6062 = n6008 | n6060 ;
  assign n6063 = ~n6061 & n6062 ;
  assign n6064 = n6057 | n6063 ;
  assign n6065 = ( n6031 & n6033 ) | ( n6031 & ~n6044 ) | ( n6033 & ~n6044 ) ;
  assign n6066 = n6031 & ~n6048 ;
  assign n6067 = ( n6033 & ~n6065 ) | ( n6033 & n6066 ) | ( ~n6065 & n6066 ) ;
  assign n6068 = ( n6045 & n6065 ) | ( n6045 & ~n6067 ) | ( n6065 & ~n6067 ) ;
  assign n6069 = n6002 & ~n6005 ;
  assign n6070 = ~n6002 & n6005 ;
  assign n6071 = n6069 | n6070 ;
  assign n6072 = n6038 & ~n6041 ;
  assign n6073 = ~n6038 & n6041 ;
  assign n6074 = n6072 | n6073 ;
  assign n6075 = n6071 & n6074 ;
  assign n6076 = n5998 | n6007 ;
  assign n6077 = ~n6008 & n6076 ;
  assign n6078 = n5998 & n6006 ;
  assign n6079 = ( n5996 & ~n6076 ) | ( n5996 & n6078 ) | ( ~n6076 & n6078 ) ;
  assign n6080 = n6077 | n6079 ;
  assign n6081 = n6075 | n6080 ;
  assign n6082 = ( n6075 & n6077 ) | ( n6075 & n6079 ) | ( n6077 & n6079 ) ;
  assign n6083 = ( n6068 & n6081 ) | ( n6068 & n6082 ) | ( n6081 & n6082 ) ;
  assign n6084 = n6064 & n6083 ;
  assign n6085 = n6057 & n6063 ;
  assign n6086 = n6084 | n6085 ;
  assign n6087 = ( n6009 & n6050 ) | ( n6009 & n6086 ) | ( n6050 & n6086 ) ;
  assign n6088 = n5974 & n6087 ;
  assign n6089 = ~n6009 & n6050 ;
  assign n6090 = n6009 & ~n6050 ;
  assign n6091 = n6089 | n6090 ;
  assign n6092 = n6085 | n6091 ;
  assign n6093 = n6084 | n6092 ;
  assign n6094 = n6086 & n6091 ;
  assign n6095 = n6093 & ~n6094 ;
  assign n6096 = ~n5898 & n5939 ;
  assign n6097 = n5898 & ~n5939 ;
  assign n6098 = n6096 | n6097 ;
  assign n6099 = n5973 | n6098 ;
  assign n6100 = ~n6098 & n6099 ;
  assign n6101 = ( ~n5973 & n6099 ) | ( ~n5973 & n6100 ) | ( n6099 & n6100 ) ;
  assign n6102 = n6095 | n6101 ;
  assign n6103 = ( n5959 & ~n5966 ) | ( n5959 & n5972 ) | ( ~n5966 & n5972 ) ;
  assign n6104 = ( ~n5959 & n5966 ) | ( ~n5959 & n6103 ) | ( n5966 & n6103 ) ;
  assign n6105 = ( ~n5972 & n6103 ) | ( ~n5972 & n6104 ) | ( n6103 & n6104 ) ;
  assign n6106 = ( ~n6057 & n6063 ) | ( ~n6057 & n6083 ) | ( n6063 & n6083 ) ;
  assign n6107 = ( n6057 & ~n6083 ) | ( n6057 & n6106 ) | ( ~n6083 & n6106 ) ;
  assign n6108 = ( ~n6063 & n6106 ) | ( ~n6063 & n6107 ) | ( n6106 & n6107 ) ;
  assign n6109 = n6071 & ~n6074 ;
  assign n6110 = ~n6071 & n6074 ;
  assign n6111 = n6109 | n6110 ;
  assign n6112 = n5946 & ~n5949 ;
  assign n6113 = ~n5946 & n5949 ;
  assign n6114 = n6112 | n6113 ;
  assign n6115 = n6111 & n6114 ;
  assign n6116 = ~n6075 & n6081 ;
  assign n6117 = ( ~n6080 & n6081 ) | ( ~n6080 & n6116 ) | ( n6081 & n6116 ) ;
  assign n6118 = n6068 & ~n6117 ;
  assign n6119 = ~n6068 & n6117 ;
  assign n6120 = n6118 | n6119 ;
  assign n6121 = ( n5943 & n5950 ) | ( n5943 & ~n5955 ) | ( n5950 & ~n5955 ) ;
  assign n6122 = ( ~n5943 & n5955 ) | ( ~n5943 & n6121 ) | ( n5955 & n6121 ) ;
  assign n6123 = ( ~n5950 & n6121 ) | ( ~n5950 & n6122 ) | ( n6121 & n6122 ) ;
  assign n6124 = ( n6115 & n6120 ) | ( n6115 & n6123 ) | ( n6120 & n6123 ) ;
  assign n6125 = ( n6105 & n6108 ) | ( n6105 & n6124 ) | ( n6108 & n6124 ) ;
  assign n6126 = n6102 & n6125 ;
  assign n6127 = n6095 & n6101 ;
  assign n6128 = n6126 | n6127 ;
  assign n6129 = n6087 & ~n6088 ;
  assign n6130 = ( n5974 & ~n6088 ) | ( n5974 & n6129 ) | ( ~n6088 & n6129 ) ;
  assign n6131 = n6128 & n6130 ;
  assign n6132 = ( n6087 & n6128 ) | ( n6087 & n6131 ) | ( n6128 & n6131 ) ;
  assign n6133 = n6088 | n6132 ;
  assign n6134 = n5863 & n6133 ;
  assign n6135 = n5859 | n6088 ;
  assign n6136 = n5862 | n6135 ;
  assign n6137 = ( n5855 & n6135 ) | ( n5855 & n6136 ) | ( n6135 & n6136 ) ;
  assign n6138 = n6132 | n6137 ;
  assign n6139 = n5854 | n5861 ;
  assign n6140 = n5853 | n6139 ;
  assign n6141 = n5855 & n5861 ;
  assign n6142 = n6140 & ~n6141 ;
  assign n6143 = n6127 | n6130 ;
  assign n6144 = n6126 | n6143 ;
  assign n6145 = ~n6131 & n6144 ;
  assign n6146 = n6142 | n6145 ;
  assign n6147 = ( ~n5832 & n5835 ) | ( ~n5832 & n5851 ) | ( n5835 & n5851 ) ;
  assign n6148 = ( n5832 & ~n5851 ) | ( n5832 & n6147 ) | ( ~n5851 & n6147 ) ;
  assign n6149 = ( ~n5835 & n6147 ) | ( ~n5835 & n6148 ) | ( n6147 & n6148 ) ;
  assign n6150 = ( ~n6105 & n6108 ) | ( ~n6105 & n6124 ) | ( n6108 & n6124 ) ;
  assign n6151 = ( n6105 & ~n6124 ) | ( n6105 & n6150 ) | ( ~n6124 & n6150 ) ;
  assign n6152 = ( ~n6108 & n6150 ) | ( ~n6108 & n6151 ) | ( n6150 & n6151 ) ;
  assign n6153 = n6111 & ~n6114 ;
  assign n6154 = ~n6111 & n6114 ;
  assign n6155 = n6153 | n6154 ;
  assign n6156 = n5838 & ~n5841 ;
  assign n6157 = ~n5838 & n5841 ;
  assign n6158 = n6156 | n6157 ;
  assign n6159 = n6155 & n6158 ;
  assign n6160 = ( n6115 & ~n6120 ) | ( n6115 & n6123 ) | ( ~n6120 & n6123 ) ;
  assign n6161 = ( ~n6115 & n6120 ) | ( ~n6115 & n6160 ) | ( n6120 & n6160 ) ;
  assign n6162 = ( ~n6123 & n6160 ) | ( ~n6123 & n6161 ) | ( n6160 & n6161 ) ;
  assign n6163 = ( n5842 & ~n5847 ) | ( n5842 & n5850 ) | ( ~n5847 & n5850 ) ;
  assign n6164 = ( ~n5842 & n5847 ) | ( ~n5842 & n6163 ) | ( n5847 & n6163 ) ;
  assign n6165 = ( ~n5850 & n6163 ) | ( ~n5850 & n6164 ) | ( n6163 & n6164 ) ;
  assign n6166 = ( n6159 & n6162 ) | ( n6159 & n6165 ) | ( n6162 & n6165 ) ;
  assign n6167 = ( n6149 & n6152 ) | ( n6149 & n6166 ) | ( n6152 & n6166 ) ;
  assign n6168 = ( ~n6095 & n6101 ) | ( ~n6095 & n6125 ) | ( n6101 & n6125 ) ;
  assign n6169 = ( n6095 & ~n6125 ) | ( n6095 & n6168 ) | ( ~n6125 & n6168 ) ;
  assign n6170 = ( ~n6101 & n6168 ) | ( ~n6101 & n6169 ) | ( n6168 & n6169 ) ;
  assign n6171 = ( ~n5712 & n5828 ) | ( ~n5712 & n5852 ) | ( n5828 & n5852 ) ;
  assign n6172 = ( n5712 & ~n5852 ) | ( n5712 & n6171 ) | ( ~n5852 & n6171 ) ;
  assign n6173 = ( ~n5828 & n6171 ) | ( ~n5828 & n6172 ) | ( n6171 & n6172 ) ;
  assign n6174 = ( n6167 & n6170 ) | ( n6167 & n6173 ) | ( n6170 & n6173 ) ;
  assign n6175 = n6146 & n6174 ;
  assign n6176 = n6142 & n6145 ;
  assign n6177 = n6175 | n6176 ;
  assign n6178 = n6138 & n6177 ;
  assign n6179 = n6134 | n6178 ;
  assign n6180 = n5593 & n6179 ;
  assign n6181 = n5552 | n6134 ;
  assign n6182 = n5556 | n6181 ;
  assign n6183 = ( n5592 & n6181 ) | ( n5592 & n6182 ) | ( n6181 & n6182 ) ;
  assign n6184 = n6178 | n6183 ;
  assign n6185 = n6133 & ~n6134 ;
  assign n6186 = ( n5863 & ~n6134 ) | ( n5863 & n6185 ) | ( ~n6134 & n6185 ) ;
  assign n6187 = n6176 | n6186 ;
  assign n6188 = n6175 | n6187 ;
  assign n6189 = n6177 & n6186 ;
  assign n6190 = n6188 & ~n6189 ;
  assign n6191 = ( n5281 & n5551 ) | ( n5281 & ~n5592 ) | ( n5551 & ~n5592 ) ;
  assign n6192 = ( ~n5551 & n5592 ) | ( ~n5551 & n6191 ) | ( n5592 & n6191 ) ;
  assign n6193 = ( ~n5281 & n6191 ) | ( ~n5281 & n6192 ) | ( n6191 & n6192 ) ;
  assign n6194 = n6190 | n6193 ;
  assign n6195 = ( ~n5560 & n5563 ) | ( ~n5560 & n5591 ) | ( n5563 & n5591 ) ;
  assign n6196 = ( n5560 & ~n5591 ) | ( n5560 & n6195 ) | ( ~n5591 & n6195 ) ;
  assign n6197 = ( ~n5563 & n6195 ) | ( ~n5563 & n6196 ) | ( n6195 & n6196 ) ;
  assign n6198 = ( ~n6142 & n6145 ) | ( ~n6142 & n6174 ) | ( n6145 & n6174 ) ;
  assign n6199 = ( n6142 & ~n6174 ) | ( n6142 & n6198 ) | ( ~n6174 & n6198 ) ;
  assign n6200 = ( ~n6145 & n6198 ) | ( ~n6145 & n6199 ) | ( n6198 & n6199 ) ;
  assign n6201 = ( ~n5566 & n5569 ) | ( ~n5566 & n5583 ) | ( n5569 & n5583 ) ;
  assign n6202 = ( n5566 & ~n5583 ) | ( n5566 & n6201 ) | ( ~n5583 & n6201 ) ;
  assign n6203 = ( ~n5569 & n6201 ) | ( ~n5569 & n6202 ) | ( n6201 & n6202 ) ;
  assign n6204 = ( ~n6149 & n6152 ) | ( ~n6149 & n6166 ) | ( n6152 & n6166 ) ;
  assign n6205 = ( n6149 & ~n6166 ) | ( n6149 & n6204 ) | ( ~n6166 & n6204 ) ;
  assign n6206 = ( ~n6152 & n6204 ) | ( ~n6152 & n6205 ) | ( n6204 & n6205 ) ;
  assign n6207 = n5572 & ~n5575 ;
  assign n6208 = ~n5572 & n5575 ;
  assign n6209 = n6207 | n6208 ;
  assign n6210 = n6155 & ~n6158 ;
  assign n6211 = ~n6155 & n6158 ;
  assign n6212 = n6210 | n6211 ;
  assign n6213 = n6209 & n6212 ;
  assign n6214 = ~n6159 & n6162 ;
  assign n6215 = n6159 & ~n6162 ;
  assign n6216 = n6214 | n6215 ;
  assign n6217 = n6165 & ~n6216 ;
  assign n6218 = ~n6165 & n6216 ;
  assign n6219 = n6217 | n6218 ;
  assign n6220 = ( n5576 & n5582 ) | ( n5576 & ~n5583 ) | ( n5582 & ~n5583 ) ;
  assign n6221 = ( n5579 & ~n5583 ) | ( n5579 & n6220 ) | ( ~n5583 & n6220 ) ;
  assign n6222 = ( n6213 & n6219 ) | ( n6213 & n6221 ) | ( n6219 & n6221 ) ;
  assign n6223 = ( n6203 & n6206 ) | ( n6203 & n6222 ) | ( n6206 & n6222 ) ;
  assign n6224 = ( n6167 & ~n6170 ) | ( n6167 & n6173 ) | ( ~n6170 & n6173 ) ;
  assign n6225 = ( ~n6167 & n6170 ) | ( ~n6167 & n6224 ) | ( n6170 & n6224 ) ;
  assign n6226 = ( ~n6173 & n6224 ) | ( ~n6173 & n6225 ) | ( n6224 & n6225 ) ;
  assign n6227 = ( n5584 & ~n5587 ) | ( n5584 & n5590 ) | ( ~n5587 & n5590 ) ;
  assign n6228 = ( ~n5584 & n5587 ) | ( ~n5584 & n6227 ) | ( n5587 & n6227 ) ;
  assign n6229 = ( ~n5590 & n6227 ) | ( ~n5590 & n6228 ) | ( n6227 & n6228 ) ;
  assign n6230 = ( n6223 & n6226 ) | ( n6223 & n6229 ) | ( n6226 & n6229 ) ;
  assign n6231 = ( n6197 & n6200 ) | ( n6197 & n6230 ) | ( n6200 & n6230 ) ;
  assign n6232 = n6194 & n6231 ;
  assign n6233 = n6190 & n6193 ;
  assign n6234 = n6232 | n6233 ;
  assign n6235 = ( n6180 & n6184 ) | ( n6180 & n6234 ) | ( n6184 & n6234 ) ;
  assign n6236 = ( x682 & x683 ) | ( x682 & x684 ) | ( x683 & x684 ) ;
  assign n6237 = ( x679 & x680 ) | ( x679 & x681 ) | ( x680 & x681 ) ;
  assign n6238 = ( x679 & ~x680 ) | ( x679 & x681 ) | ( ~x680 & x681 ) ;
  assign n6239 = ( ~x679 & x680 ) | ( ~x679 & n6238 ) | ( x680 & n6238 ) ;
  assign n6240 = ( ~x681 & n6238 ) | ( ~x681 & n6239 ) | ( n6238 & n6239 ) ;
  assign n6241 = ( x682 & ~x683 ) | ( x682 & x684 ) | ( ~x683 & x684 ) ;
  assign n6242 = ( ~x682 & x683 ) | ( ~x682 & n6241 ) | ( x683 & n6241 ) ;
  assign n6243 = ( ~x684 & n6241 ) | ( ~x684 & n6242 ) | ( n6241 & n6242 ) ;
  assign n6244 = n6240 & n6243 ;
  assign n6245 = ( n6236 & n6237 ) | ( n6236 & n6244 ) | ( n6237 & n6244 ) ;
  assign n6246 = ( n6237 & n6244 ) | ( n6237 & ~n6245 ) | ( n6244 & ~n6245 ) ;
  assign n6247 = ( n6236 & ~n6245 ) | ( n6236 & n6246 ) | ( ~n6245 & n6246 ) ;
  assign n6248 = ( x688 & x689 ) | ( x688 & x690 ) | ( x689 & x690 ) ;
  assign n6249 = ( x685 & x686 ) | ( x685 & x687 ) | ( x686 & x687 ) ;
  assign n6250 = ( x685 & ~x686 ) | ( x685 & x687 ) | ( ~x686 & x687 ) ;
  assign n6251 = ( ~x685 & x686 ) | ( ~x685 & n6250 ) | ( x686 & n6250 ) ;
  assign n6252 = ( ~x687 & n6250 ) | ( ~x687 & n6251 ) | ( n6250 & n6251 ) ;
  assign n6253 = ( x688 & ~x689 ) | ( x688 & x690 ) | ( ~x689 & x690 ) ;
  assign n6254 = ( ~x688 & x689 ) | ( ~x688 & n6253 ) | ( x689 & n6253 ) ;
  assign n6255 = ( ~x690 & n6253 ) | ( ~x690 & n6254 ) | ( n6253 & n6254 ) ;
  assign n6256 = n6252 & n6255 ;
  assign n6257 = ( n6248 & n6249 ) | ( n6248 & n6256 ) | ( n6249 & n6256 ) ;
  assign n6258 = ( n6249 & n6256 ) | ( n6249 & ~n6257 ) | ( n6256 & ~n6257 ) ;
  assign n6259 = ( n6248 & ~n6257 ) | ( n6248 & n6258 ) | ( ~n6257 & n6258 ) ;
  assign n6260 = n6245 & n6247 ;
  assign n6261 = n6257 & n6259 ;
  assign n6262 = n6240 & ~n6243 ;
  assign n6263 = ~n6240 & n6243 ;
  assign n6264 = n6262 | n6263 ;
  assign n6265 = n6252 & ~n6255 ;
  assign n6266 = ~n6252 & n6255 ;
  assign n6267 = n6265 | n6266 ;
  assign n6268 = n6264 & n6267 ;
  assign n6269 = ~n6261 & n6268 ;
  assign n6270 = ~n6260 & n6269 ;
  assign n6271 = ~n6259 & n6270 ;
  assign n6272 = ( n6247 & n6259 ) | ( n6247 & n6271 ) | ( n6259 & n6271 ) ;
  assign n6273 = n6259 & n6269 ;
  assign n6274 = ~n6260 & n6273 ;
  assign n6275 = ~n6245 & n6257 ;
  assign n6276 = n6245 & ~n6257 ;
  assign n6277 = n6275 | n6276 ;
  assign n6278 = n6274 | n6277 ;
  assign n6279 = n6272 | n6278 ;
  assign n6280 = n6272 | n6274 ;
  assign n6281 = n6277 & n6280 ;
  assign n6282 = n6279 & ~n6281 ;
  assign n6283 = ( x694 & x695 ) | ( x694 & x696 ) | ( x695 & x696 ) ;
  assign n6284 = ( x691 & x692 ) | ( x691 & x693 ) | ( x692 & x693 ) ;
  assign n6285 = ( x691 & ~x692 ) | ( x691 & x693 ) | ( ~x692 & x693 ) ;
  assign n6286 = ( ~x691 & x692 ) | ( ~x691 & n6285 ) | ( x692 & n6285 ) ;
  assign n6287 = ( ~x693 & n6285 ) | ( ~x693 & n6286 ) | ( n6285 & n6286 ) ;
  assign n6288 = ( x694 & ~x695 ) | ( x694 & x696 ) | ( ~x695 & x696 ) ;
  assign n6289 = ( ~x694 & x695 ) | ( ~x694 & n6288 ) | ( x695 & n6288 ) ;
  assign n6290 = ( ~x696 & n6288 ) | ( ~x696 & n6289 ) | ( n6288 & n6289 ) ;
  assign n6291 = n6287 & n6290 ;
  assign n6292 = ( n6283 & n6284 ) | ( n6283 & n6291 ) | ( n6284 & n6291 ) ;
  assign n6293 = ( n6284 & n6291 ) | ( n6284 & ~n6292 ) | ( n6291 & ~n6292 ) ;
  assign n6294 = ( n6283 & ~n6292 ) | ( n6283 & n6293 ) | ( ~n6292 & n6293 ) ;
  assign n6295 = ( x700 & x701 ) | ( x700 & x702 ) | ( x701 & x702 ) ;
  assign n6296 = ( x697 & x698 ) | ( x697 & x699 ) | ( x698 & x699 ) ;
  assign n6297 = ( x697 & ~x698 ) | ( x697 & x699 ) | ( ~x698 & x699 ) ;
  assign n6298 = ( ~x697 & x698 ) | ( ~x697 & n6297 ) | ( x698 & n6297 ) ;
  assign n6299 = ( ~x699 & n6297 ) | ( ~x699 & n6298 ) | ( n6297 & n6298 ) ;
  assign n6300 = ( x700 & ~x701 ) | ( x700 & x702 ) | ( ~x701 & x702 ) ;
  assign n6301 = ( ~x700 & x701 ) | ( ~x700 & n6300 ) | ( x701 & n6300 ) ;
  assign n6302 = ( ~x702 & n6300 ) | ( ~x702 & n6301 ) | ( n6300 & n6301 ) ;
  assign n6303 = n6299 & n6302 ;
  assign n6304 = ( n6295 & n6296 ) | ( n6295 & n6303 ) | ( n6296 & n6303 ) ;
  assign n6305 = ( n6296 & n6303 ) | ( n6296 & ~n6304 ) | ( n6303 & ~n6304 ) ;
  assign n6306 = ( n6295 & ~n6304 ) | ( n6295 & n6305 ) | ( ~n6304 & n6305 ) ;
  assign n6307 = n6292 & n6294 ;
  assign n6308 = n6287 & ~n6290 ;
  assign n6309 = ~n6287 & n6290 ;
  assign n6310 = n6308 | n6309 ;
  assign n6311 = n6299 & ~n6302 ;
  assign n6312 = ~n6299 & n6302 ;
  assign n6313 = n6311 | n6312 ;
  assign n6314 = n6310 & n6313 ;
  assign n6315 = ~n6307 & n6314 ;
  assign n6316 = ( n6294 & n6306 ) | ( n6294 & n6315 ) | ( n6306 & n6315 ) ;
  assign n6317 = ~n6292 & n6304 ;
  assign n6318 = n6292 & ~n6304 ;
  assign n6319 = n6317 | n6318 ;
  assign n6320 = n6316 & n6319 ;
  assign n6321 = n6316 | n6319 ;
  assign n6322 = ~n6320 & n6321 ;
  assign n6323 = n6282 | n6322 ;
  assign n6324 = ( n6247 & n6259 ) | ( n6247 & ~n6270 ) | ( n6259 & ~n6270 ) ;
  assign n6325 = n6247 & ~n6274 ;
  assign n6326 = ( n6259 & ~n6324 ) | ( n6259 & n6325 ) | ( ~n6324 & n6325 ) ;
  assign n6327 = ( n6271 & n6324 ) | ( n6271 & ~n6326 ) | ( n6324 & ~n6326 ) ;
  assign n6328 = n6310 & ~n6313 ;
  assign n6329 = ~n6310 & n6313 ;
  assign n6330 = n6328 | n6329 ;
  assign n6331 = n6264 & ~n6267 ;
  assign n6332 = ~n6264 & n6267 ;
  assign n6333 = n6331 | n6332 ;
  assign n6334 = n6330 & n6333 ;
  assign n6335 = n6306 | n6315 ;
  assign n6336 = ~n6316 & n6335 ;
  assign n6337 = n6306 & n6314 ;
  assign n6338 = ( n6294 & ~n6335 ) | ( n6294 & n6337 ) | ( ~n6335 & n6337 ) ;
  assign n6339 = n6336 | n6338 ;
  assign n6340 = n6334 | n6339 ;
  assign n6341 = ( n6334 & n6336 ) | ( n6334 & n6338 ) | ( n6336 & n6338 ) ;
  assign n6342 = ( n6327 & n6340 ) | ( n6327 & n6341 ) | ( n6340 & n6341 ) ;
  assign n6343 = n6323 & n6342 ;
  assign n6344 = n6282 & n6322 ;
  assign n6345 = ( n6292 & n6304 ) | ( n6292 & n6316 ) | ( n6304 & n6316 ) ;
  assign n6346 = ( n6245 & n6257 ) | ( n6245 & n6280 ) | ( n6257 & n6280 ) ;
  assign n6347 = ~n6345 & n6346 ;
  assign n6348 = n6345 & ~n6346 ;
  assign n6349 = n6347 | n6348 ;
  assign n6350 = n6344 | n6349 ;
  assign n6351 = n6343 | n6350 ;
  assign n6352 = n6343 | n6344 ;
  assign n6353 = n6349 & n6352 ;
  assign n6354 = n6351 & ~n6353 ;
  assign n6390 = ( x664 & x665 ) | ( x664 & x666 ) | ( x665 & x666 ) ;
  assign n6391 = ( x661 & x662 ) | ( x661 & x663 ) | ( x662 & x663 ) ;
  assign n6392 = ( x661 & ~x662 ) | ( x661 & x663 ) | ( ~x662 & x663 ) ;
  assign n6393 = ( ~x661 & x662 ) | ( ~x661 & n6392 ) | ( x662 & n6392 ) ;
  assign n6394 = ( ~x663 & n6392 ) | ( ~x663 & n6393 ) | ( n6392 & n6393 ) ;
  assign n6395 = ( x664 & ~x665 ) | ( x664 & x666 ) | ( ~x665 & x666 ) ;
  assign n6396 = ( ~x664 & x665 ) | ( ~x664 & n6395 ) | ( x665 & n6395 ) ;
  assign n6397 = ( ~x666 & n6395 ) | ( ~x666 & n6396 ) | ( n6395 & n6396 ) ;
  assign n6398 = n6394 & n6397 ;
  assign n6399 = ( n6390 & n6391 ) | ( n6390 & n6398 ) | ( n6391 & n6398 ) ;
  assign n6413 = ( n6391 & n6398 ) | ( n6391 & ~n6399 ) | ( n6398 & ~n6399 ) ;
  assign n6414 = ( n6390 & ~n6399 ) | ( n6390 & n6413 ) | ( ~n6399 & n6413 ) ;
  assign n6400 = ( x658 & x659 ) | ( x658 & x660 ) | ( x659 & x660 ) ;
  assign n6401 = ( x655 & x656 ) | ( x655 & x657 ) | ( x656 & x657 ) ;
  assign n6402 = ( x655 & ~x656 ) | ( x655 & x657 ) | ( ~x656 & x657 ) ;
  assign n6403 = ( ~x655 & x656 ) | ( ~x655 & n6402 ) | ( x656 & n6402 ) ;
  assign n6404 = ( ~x657 & n6402 ) | ( ~x657 & n6403 ) | ( n6402 & n6403 ) ;
  assign n6405 = ( x658 & ~x659 ) | ( x658 & x660 ) | ( ~x659 & x660 ) ;
  assign n6406 = ( ~x658 & x659 ) | ( ~x658 & n6405 ) | ( x659 & n6405 ) ;
  assign n6407 = ( ~x660 & n6405 ) | ( ~x660 & n6406 ) | ( n6405 & n6406 ) ;
  assign n6408 = n6404 & n6407 ;
  assign n6409 = ( n6400 & n6401 ) | ( n6400 & n6408 ) | ( n6401 & n6408 ) ;
  assign n6410 = ( n6401 & n6408 ) | ( n6401 & ~n6409 ) | ( n6408 & ~n6409 ) ;
  assign n6411 = ( n6400 & ~n6409 ) | ( n6400 & n6410 ) | ( ~n6409 & n6410 ) ;
  assign n6412 = n6409 & n6411 ;
  assign n6415 = n6399 & n6414 ;
  assign n6416 = n6394 & ~n6397 ;
  assign n6417 = ~n6394 & n6397 ;
  assign n6418 = n6416 | n6417 ;
  assign n6419 = n6404 & ~n6407 ;
  assign n6420 = ~n6404 & n6407 ;
  assign n6421 = n6419 | n6420 ;
  assign n6422 = n6418 & n6421 ;
  assign n6423 = ~n6415 & n6422 ;
  assign n6426 = ~n6412 & n6423 ;
  assign n6427 = ~n6414 & n6426 ;
  assign n6434 = ( n6411 & n6414 ) | ( n6411 & ~n6426 ) | ( n6414 & ~n6426 ) ;
  assign n6424 = n6414 & n6423 ;
  assign n6425 = ~n6412 & n6424 ;
  assign n6435 = n6411 & ~n6425 ;
  assign n6436 = ( n6414 & ~n6434 ) | ( n6414 & n6435 ) | ( ~n6434 & n6435 ) ;
  assign n6437 = ( n6427 & n6434 ) | ( n6427 & ~n6436 ) | ( n6434 & ~n6436 ) ;
  assign n6357 = ( x667 & ~x668 ) | ( x667 & x669 ) | ( ~x668 & x669 ) ;
  assign n6358 = ( ~x667 & x668 ) | ( ~x667 & n6357 ) | ( x668 & n6357 ) ;
  assign n6359 = ( ~x669 & n6357 ) | ( ~x669 & n6358 ) | ( n6357 & n6358 ) ;
  assign n6360 = ( x670 & ~x671 ) | ( x670 & x672 ) | ( ~x671 & x672 ) ;
  assign n6361 = ( ~x670 & x671 ) | ( ~x670 & n6360 ) | ( x671 & n6360 ) ;
  assign n6362 = ( ~x672 & n6360 ) | ( ~x672 & n6361 ) | ( n6360 & n6361 ) ;
  assign n6380 = n6359 & ~n6362 ;
  assign n6381 = ~n6359 & n6362 ;
  assign n6382 = n6380 | n6381 ;
  assign n6367 = ( x673 & ~x674 ) | ( x673 & x675 ) | ( ~x674 & x675 ) ;
  assign n6368 = ( ~x673 & x674 ) | ( ~x673 & n6367 ) | ( x674 & n6367 ) ;
  assign n6369 = ( ~x675 & n6367 ) | ( ~x675 & n6368 ) | ( n6367 & n6368 ) ;
  assign n6370 = ( x676 & ~x677 ) | ( x676 & x678 ) | ( ~x677 & x678 ) ;
  assign n6371 = ( ~x676 & x677 ) | ( ~x676 & n6370 ) | ( x677 & n6370 ) ;
  assign n6372 = ( ~x678 & n6370 ) | ( ~x678 & n6371 ) | ( n6370 & n6371 ) ;
  assign n6383 = n6369 & ~n6372 ;
  assign n6384 = ~n6369 & n6372 ;
  assign n6385 = n6383 | n6384 ;
  assign n6438 = n6382 & ~n6385 ;
  assign n6439 = ~n6382 & n6385 ;
  assign n6440 = n6438 | n6439 ;
  assign n6441 = ~n6418 & n6421 ;
  assign n6442 = n6418 & ~n6421 ;
  assign n6443 = n6441 | n6442 ;
  assign n6444 = n6440 & n6443 ;
  assign n6355 = ( x670 & x671 ) | ( x670 & x672 ) | ( x671 & x672 ) ;
  assign n6356 = ( x667 & x668 ) | ( x667 & x669 ) | ( x668 & x669 ) ;
  assign n6363 = n6359 & n6362 ;
  assign n6364 = ( n6355 & n6356 ) | ( n6355 & n6363 ) | ( n6356 & n6363 ) ;
  assign n6375 = ( n6356 & n6363 ) | ( n6356 & ~n6364 ) | ( n6363 & ~n6364 ) ;
  assign n6376 = ( n6355 & ~n6364 ) | ( n6355 & n6375 ) | ( ~n6364 & n6375 ) ;
  assign n6365 = ( x676 & x677 ) | ( x676 & x678 ) | ( x677 & x678 ) ;
  assign n6366 = ( x673 & x674 ) | ( x673 & x675 ) | ( x674 & x675 ) ;
  assign n6373 = n6369 & n6372 ;
  assign n6374 = ( n6365 & n6366 ) | ( n6365 & n6373 ) | ( n6366 & n6373 ) ;
  assign n6377 = ( n6366 & n6373 ) | ( n6366 & ~n6374 ) | ( n6373 & ~n6374 ) ;
  assign n6378 = ( n6365 & ~n6374 ) | ( n6365 & n6377 ) | ( ~n6374 & n6377 ) ;
  assign n6386 = n6382 & n6385 ;
  assign n6445 = n6378 & n6386 ;
  assign n6379 = n6364 & n6376 ;
  assign n6387 = ~n6379 & n6386 ;
  assign n6446 = n6378 | n6387 ;
  assign n6447 = ( n6376 & n6445 ) | ( n6376 & ~n6446 ) | ( n6445 & ~n6446 ) ;
  assign n6388 = ( n6376 & n6378 ) | ( n6376 & n6387 ) | ( n6378 & n6387 ) ;
  assign n6448 = ~n6388 & n6446 ;
  assign n6449 = n6447 | n6448 ;
  assign n6450 = n6444 | n6449 ;
  assign n6451 = n6437 & n6450 ;
  assign n6452 = ( n6444 & n6447 ) | ( n6444 & n6448 ) | ( n6447 & n6448 ) ;
  assign n6453 = n6451 | n6452 ;
  assign n6428 = ( n6411 & n6414 ) | ( n6411 & n6427 ) | ( n6414 & n6427 ) ;
  assign n6454 = n6399 & ~n6409 ;
  assign n6455 = ~n6399 & n6409 ;
  assign n6456 = n6454 | n6455 ;
  assign n6457 = n6425 | n6456 ;
  assign n6458 = n6428 | n6457 ;
  assign n6429 = n6425 | n6428 ;
  assign n6459 = n6429 & n6456 ;
  assign n6460 = n6458 & ~n6459 ;
  assign n6461 = ~n6364 & n6374 ;
  assign n6462 = n6364 & ~n6374 ;
  assign n6463 = n6461 | n6462 ;
  assign n6464 = n6388 & n6463 ;
  assign n6465 = n6388 | n6463 ;
  assign n6466 = ~n6464 & n6465 ;
  assign n6467 = ( n6453 & n6460 ) | ( n6453 & n6466 ) | ( n6460 & n6466 ) ;
  assign n6389 = ( n6364 & n6374 ) | ( n6364 & n6388 ) | ( n6374 & n6388 ) ;
  assign n6430 = ( n6399 & n6409 ) | ( n6399 & n6429 ) | ( n6409 & n6429 ) ;
  assign n6431 = n6389 & n6430 ;
  assign n6432 = n6430 & ~n6431 ;
  assign n6433 = ( n6389 & ~n6431 ) | ( n6389 & n6432 ) | ( ~n6431 & n6432 ) ;
  assign n6468 = n6433 | n6467 ;
  assign n6469 = ~n6433 & n6468 ;
  assign n6470 = ( ~n6467 & n6468 ) | ( ~n6467 & n6469 ) | ( n6468 & n6469 ) ;
  assign n6471 = n6354 | n6470 ;
  assign n6472 = ( n6453 & ~n6460 ) | ( n6453 & n6466 ) | ( ~n6460 & n6466 ) ;
  assign n6473 = ( ~n6453 & n6460 ) | ( ~n6453 & n6472 ) | ( n6460 & n6472 ) ;
  assign n6474 = ( ~n6466 & n6472 ) | ( ~n6466 & n6473 ) | ( n6472 & n6473 ) ;
  assign n6475 = ( ~n6282 & n6322 ) | ( ~n6282 & n6342 ) | ( n6322 & n6342 ) ;
  assign n6476 = ( n6282 & ~n6342 ) | ( n6282 & n6475 ) | ( ~n6342 & n6475 ) ;
  assign n6477 = ( ~n6322 & n6475 ) | ( ~n6322 & n6476 ) | ( n6475 & n6476 ) ;
  assign n6478 = n6330 & ~n6333 ;
  assign n6479 = ~n6330 & n6333 ;
  assign n6480 = n6478 | n6479 ;
  assign n6481 = n6440 & ~n6443 ;
  assign n6482 = ~n6440 & n6443 ;
  assign n6483 = n6481 | n6482 ;
  assign n6484 = n6480 & n6483 ;
  assign n6485 = ~n6334 & n6340 ;
  assign n6486 = ( ~n6339 & n6340 ) | ( ~n6339 & n6485 ) | ( n6340 & n6485 ) ;
  assign n6487 = n6327 & ~n6486 ;
  assign n6488 = ~n6327 & n6486 ;
  assign n6489 = n6487 | n6488 ;
  assign n6490 = ( n6437 & n6444 ) | ( n6437 & ~n6449 ) | ( n6444 & ~n6449 ) ;
  assign n6491 = ( ~n6437 & n6449 ) | ( ~n6437 & n6490 ) | ( n6449 & n6490 ) ;
  assign n6492 = ( ~n6444 & n6490 ) | ( ~n6444 & n6491 ) | ( n6490 & n6491 ) ;
  assign n6493 = ( n6484 & n6489 ) | ( n6484 & n6492 ) | ( n6489 & n6492 ) ;
  assign n6494 = ( n6474 & n6477 ) | ( n6474 & n6493 ) | ( n6477 & n6493 ) ;
  assign n6495 = n6471 & n6494 ;
  assign n6496 = n6354 & n6470 ;
  assign n6497 = n6495 | n6496 ;
  assign n6498 = n6431 | n6433 ;
  assign n6499 = ( n6431 & n6467 ) | ( n6431 & n6498 ) | ( n6467 & n6498 ) ;
  assign n6500 = ( n6345 & n6346 ) | ( n6345 & n6352 ) | ( n6346 & n6352 ) ;
  assign n6501 = n6499 & n6500 ;
  assign n6502 = n6500 & ~n6501 ;
  assign n6503 = ( n6499 & ~n6501 ) | ( n6499 & n6502 ) | ( ~n6501 & n6502 ) ;
  assign n6504 = ( n6498 & n6500 ) | ( n6498 & n6503 ) | ( n6500 & n6503 ) ;
  assign n6505 = ( n6497 & n6501 ) | ( n6497 & n6504 ) | ( n6501 & n6504 ) ;
  assign n6506 = ( x724 & x725 ) | ( x724 & x726 ) | ( x725 & x726 ) ;
  assign n6507 = ( x721 & x722 ) | ( x721 & x723 ) | ( x722 & x723 ) ;
  assign n6508 = ( x721 & ~x722 ) | ( x721 & x723 ) | ( ~x722 & x723 ) ;
  assign n6509 = ( ~x721 & x722 ) | ( ~x721 & n6508 ) | ( x722 & n6508 ) ;
  assign n6510 = ( ~x723 & n6508 ) | ( ~x723 & n6509 ) | ( n6508 & n6509 ) ;
  assign n6511 = ( x724 & ~x725 ) | ( x724 & x726 ) | ( ~x725 & x726 ) ;
  assign n6512 = ( ~x724 & x725 ) | ( ~x724 & n6511 ) | ( x725 & n6511 ) ;
  assign n6513 = ( ~x726 & n6511 ) | ( ~x726 & n6512 ) | ( n6511 & n6512 ) ;
  assign n6514 = n6510 & n6513 ;
  assign n6515 = ( n6506 & n6507 ) | ( n6506 & n6514 ) | ( n6507 & n6514 ) ;
  assign n6516 = ( x715 & ~x716 ) | ( x715 & x717 ) | ( ~x716 & x717 ) ;
  assign n6517 = ( ~x715 & x716 ) | ( ~x715 & n6516 ) | ( x716 & n6516 ) ;
  assign n6518 = ( ~x717 & n6516 ) | ( ~x717 & n6517 ) | ( n6516 & n6517 ) ;
  assign n6519 = ( x718 & ~x719 ) | ( x718 & x720 ) | ( ~x719 & x720 ) ;
  assign n6520 = ( ~x718 & x719 ) | ( ~x718 & n6519 ) | ( x719 & n6519 ) ;
  assign n6521 = ( ~x720 & n6519 ) | ( ~x720 & n6520 ) | ( n6519 & n6520 ) ;
  assign n6522 = n6518 & n6521 ;
  assign n6523 = ( x718 & x719 ) | ( x718 & x720 ) | ( x719 & x720 ) ;
  assign n6524 = ( x715 & x716 ) | ( x715 & x717 ) | ( x716 & x717 ) ;
  assign n6525 = ( n6522 & n6523 ) | ( n6522 & n6524 ) | ( n6523 & n6524 ) ;
  assign n6526 = ( n6507 & n6514 ) | ( n6507 & ~n6515 ) | ( n6514 & ~n6515 ) ;
  assign n6527 = ( n6506 & ~n6515 ) | ( n6506 & n6526 ) | ( ~n6515 & n6526 ) ;
  assign n6528 = ( n6522 & n6524 ) | ( n6522 & ~n6525 ) | ( n6524 & ~n6525 ) ;
  assign n6529 = ( n6523 & ~n6525 ) | ( n6523 & n6528 ) | ( ~n6525 & n6528 ) ;
  assign n6530 = n6525 & n6529 ;
  assign n6531 = n6510 & ~n6513 ;
  assign n6532 = ~n6510 & n6513 ;
  assign n6533 = n6531 | n6532 ;
  assign n6534 = n6518 & ~n6521 ;
  assign n6535 = ~n6518 & n6521 ;
  assign n6536 = n6534 | n6535 ;
  assign n6537 = n6533 & n6536 ;
  assign n6538 = ~n6530 & n6537 ;
  assign n6539 = ( n6527 & n6529 ) | ( n6527 & n6538 ) | ( n6529 & n6538 ) ;
  assign n6540 = ( n6515 & n6525 ) | ( n6515 & n6539 ) | ( n6525 & n6539 ) ;
  assign n6541 = ( x712 & x713 ) | ( x712 & x714 ) | ( x713 & x714 ) ;
  assign n6542 = ( x709 & x710 ) | ( x709 & x711 ) | ( x710 & x711 ) ;
  assign n6543 = ( x709 & ~x710 ) | ( x709 & x711 ) | ( ~x710 & x711 ) ;
  assign n6544 = ( ~x709 & x710 ) | ( ~x709 & n6543 ) | ( x710 & n6543 ) ;
  assign n6545 = ( ~x711 & n6543 ) | ( ~x711 & n6544 ) | ( n6543 & n6544 ) ;
  assign n6546 = ( x712 & ~x713 ) | ( x712 & x714 ) | ( ~x713 & x714 ) ;
  assign n6547 = ( ~x712 & x713 ) | ( ~x712 & n6546 ) | ( x713 & n6546 ) ;
  assign n6548 = ( ~x714 & n6546 ) | ( ~x714 & n6547 ) | ( n6546 & n6547 ) ;
  assign n6549 = n6545 & n6548 ;
  assign n6550 = ( n6541 & n6542 ) | ( n6541 & n6549 ) | ( n6542 & n6549 ) ;
  assign n6551 = ( x706 & x707 ) | ( x706 & x708 ) | ( x707 & x708 ) ;
  assign n6552 = ( x703 & x704 ) | ( x703 & x705 ) | ( x704 & x705 ) ;
  assign n6553 = ( x703 & ~x704 ) | ( x703 & x705 ) | ( ~x704 & x705 ) ;
  assign n6554 = ( ~x703 & x704 ) | ( ~x703 & n6553 ) | ( x704 & n6553 ) ;
  assign n6555 = ( ~x705 & n6553 ) | ( ~x705 & n6554 ) | ( n6553 & n6554 ) ;
  assign n6556 = ( x706 & ~x707 ) | ( x706 & x708 ) | ( ~x707 & x708 ) ;
  assign n6557 = ( ~x706 & x707 ) | ( ~x706 & n6556 ) | ( x707 & n6556 ) ;
  assign n6558 = ( ~x708 & n6556 ) | ( ~x708 & n6557 ) | ( n6556 & n6557 ) ;
  assign n6559 = n6555 & n6558 ;
  assign n6560 = ( n6551 & n6552 ) | ( n6551 & n6559 ) | ( n6552 & n6559 ) ;
  assign n6561 = ( n6552 & n6559 ) | ( n6552 & ~n6560 ) | ( n6559 & ~n6560 ) ;
  assign n6562 = ( n6551 & ~n6560 ) | ( n6551 & n6561 ) | ( ~n6560 & n6561 ) ;
  assign n6563 = n6560 & n6562 ;
  assign n6564 = ( n6542 & n6549 ) | ( n6542 & ~n6550 ) | ( n6549 & ~n6550 ) ;
  assign n6565 = ( n6541 & ~n6550 ) | ( n6541 & n6564 ) | ( ~n6550 & n6564 ) ;
  assign n6566 = n6550 & n6565 ;
  assign n6567 = n6545 & ~n6548 ;
  assign n6568 = ~n6545 & n6548 ;
  assign n6569 = n6567 | n6568 ;
  assign n6570 = n6555 & ~n6558 ;
  assign n6571 = ~n6555 & n6558 ;
  assign n6572 = n6570 | n6571 ;
  assign n6573 = n6569 & n6572 ;
  assign n6574 = ~n6566 & n6573 ;
  assign n6575 = n6565 & n6574 ;
  assign n6576 = ~n6563 & n6575 ;
  assign n6577 = ~n6563 & n6574 ;
  assign n6578 = ~n6565 & n6577 ;
  assign n6579 = ( n6562 & n6565 ) | ( n6562 & n6578 ) | ( n6565 & n6578 ) ;
  assign n6580 = n6576 | n6579 ;
  assign n6581 = ( n6550 & n6560 ) | ( n6550 & n6580 ) | ( n6560 & n6580 ) ;
  assign n6582 = ( n6562 & n6565 ) | ( n6562 & ~n6577 ) | ( n6565 & ~n6577 ) ;
  assign n6583 = n6562 & ~n6576 ;
  assign n6584 = ( n6565 & ~n6582 ) | ( n6565 & n6583 ) | ( ~n6582 & n6583 ) ;
  assign n6585 = ( n6578 & n6582 ) | ( n6578 & ~n6584 ) | ( n6582 & ~n6584 ) ;
  assign n6586 = ~n6533 & n6536 ;
  assign n6587 = n6533 & ~n6536 ;
  assign n6588 = n6586 | n6587 ;
  assign n6589 = ~n6569 & n6572 ;
  assign n6590 = n6569 & ~n6572 ;
  assign n6591 = n6589 | n6590 ;
  assign n6592 = n6588 & n6591 ;
  assign n6593 = n6527 & n6537 ;
  assign n6594 = n6527 | n6538 ;
  assign n6595 = ( n6529 & n6593 ) | ( n6529 & ~n6594 ) | ( n6593 & ~n6594 ) ;
  assign n6596 = ~n6539 & n6594 ;
  assign n6597 = n6595 | n6596 ;
  assign n6598 = n6592 | n6597 ;
  assign n6599 = n6585 & n6598 ;
  assign n6600 = ( n6592 & n6595 ) | ( n6592 & n6596 ) | ( n6595 & n6596 ) ;
  assign n6601 = n6599 | n6600 ;
  assign n6602 = n6550 & ~n6560 ;
  assign n6603 = ~n6550 & n6560 ;
  assign n6604 = n6602 | n6603 ;
  assign n6605 = n6576 | n6604 ;
  assign n6606 = n6579 | n6605 ;
  assign n6607 = n6580 & n6604 ;
  assign n6608 = n6606 & ~n6607 ;
  assign n6609 = ( n6515 & n6525 ) | ( n6515 & ~n6539 ) | ( n6525 & ~n6539 ) ;
  assign n6610 = ( n6515 & ~n6525 ) | ( n6515 & n6539 ) | ( ~n6525 & n6539 ) ;
  assign n6611 = ( ~n6515 & n6609 ) | ( ~n6515 & n6610 ) | ( n6609 & n6610 ) ;
  assign n6612 = ( n6601 & n6608 ) | ( n6601 & n6611 ) | ( n6608 & n6611 ) ;
  assign n6613 = ( n6540 & n6581 ) | ( n6540 & n6612 ) | ( n6581 & n6612 ) ;
  assign n6614 = ( x748 & x749 ) | ( x748 & x750 ) | ( x749 & x750 ) ;
  assign n6615 = ( x745 & x746 ) | ( x745 & x747 ) | ( x746 & x747 ) ;
  assign n6616 = ( x745 & ~x746 ) | ( x745 & x747 ) | ( ~x746 & x747 ) ;
  assign n6617 = ( ~x745 & x746 ) | ( ~x745 & n6616 ) | ( x746 & n6616 ) ;
  assign n6618 = ( ~x747 & n6616 ) | ( ~x747 & n6617 ) | ( n6616 & n6617 ) ;
  assign n6619 = ( x748 & ~x749 ) | ( x748 & x750 ) | ( ~x749 & x750 ) ;
  assign n6620 = ( ~x748 & x749 ) | ( ~x748 & n6619 ) | ( x749 & n6619 ) ;
  assign n6621 = ( ~x750 & n6619 ) | ( ~x750 & n6620 ) | ( n6619 & n6620 ) ;
  assign n6622 = n6618 & n6621 ;
  assign n6623 = ( n6614 & n6615 ) | ( n6614 & n6622 ) | ( n6615 & n6622 ) ;
  assign n6624 = ( x739 & ~x740 ) | ( x739 & x741 ) | ( ~x740 & x741 ) ;
  assign n6625 = ( ~x739 & x740 ) | ( ~x739 & n6624 ) | ( x740 & n6624 ) ;
  assign n6626 = ( ~x741 & n6624 ) | ( ~x741 & n6625 ) | ( n6624 & n6625 ) ;
  assign n6627 = ( x742 & ~x743 ) | ( x742 & x744 ) | ( ~x743 & x744 ) ;
  assign n6628 = ( ~x742 & x743 ) | ( ~x742 & n6627 ) | ( x743 & n6627 ) ;
  assign n6629 = ( ~x744 & n6627 ) | ( ~x744 & n6628 ) | ( n6627 & n6628 ) ;
  assign n6630 = n6626 & n6629 ;
  assign n6631 = ( x742 & x743 ) | ( x742 & x744 ) | ( x743 & x744 ) ;
  assign n6632 = ( x739 & x740 ) | ( x739 & x741 ) | ( x740 & x741 ) ;
  assign n6633 = ( n6630 & n6631 ) | ( n6630 & n6632 ) | ( n6631 & n6632 ) ;
  assign n6634 = ( n6615 & n6622 ) | ( n6615 & ~n6623 ) | ( n6622 & ~n6623 ) ;
  assign n6635 = ( n6614 & ~n6623 ) | ( n6614 & n6634 ) | ( ~n6623 & n6634 ) ;
  assign n6636 = ( n6630 & n6632 ) | ( n6630 & ~n6633 ) | ( n6632 & ~n6633 ) ;
  assign n6637 = ( n6631 & ~n6633 ) | ( n6631 & n6636 ) | ( ~n6633 & n6636 ) ;
  assign n6638 = n6633 & n6637 ;
  assign n6639 = n6626 & ~n6629 ;
  assign n6640 = ~n6626 & n6629 ;
  assign n6641 = n6639 | n6640 ;
  assign n6642 = n6618 & ~n6621 ;
  assign n6643 = ~n6618 & n6621 ;
  assign n6644 = n6642 | n6643 ;
  assign n6645 = ~n6622 & n6644 ;
  assign n6646 = n6641 & n6645 ;
  assign n6647 = ~n6638 & n6646 ;
  assign n6648 = ( n6635 & n6637 ) | ( n6635 & n6647 ) | ( n6637 & n6647 ) ;
  assign n6649 = ( n6623 & n6633 ) | ( n6623 & n6648 ) | ( n6633 & n6648 ) ;
  assign n6650 = ( x727 & ~x728 ) | ( x727 & x729 ) | ( ~x728 & x729 ) ;
  assign n6651 = ( ~x727 & x728 ) | ( ~x727 & n6650 ) | ( x728 & n6650 ) ;
  assign n6652 = ( ~x729 & n6650 ) | ( ~x729 & n6651 ) | ( n6650 & n6651 ) ;
  assign n6653 = ( x730 & ~x731 ) | ( x730 & x732 ) | ( ~x731 & x732 ) ;
  assign n6654 = ( ~x730 & x731 ) | ( ~x730 & n6653 ) | ( x731 & n6653 ) ;
  assign n6655 = ( ~x732 & n6653 ) | ( ~x732 & n6654 ) | ( n6653 & n6654 ) ;
  assign n6656 = n6652 & n6655 ;
  assign n6657 = ( x730 & x731 ) | ( x730 & x732 ) | ( x731 & x732 ) ;
  assign n6658 = ( x727 & x728 ) | ( x727 & x729 ) | ( x728 & x729 ) ;
  assign n6659 = ( n6656 & n6657 ) | ( n6656 & n6658 ) | ( n6657 & n6658 ) ;
  assign n6660 = ( x736 & x737 ) | ( x736 & x738 ) | ( x737 & x738 ) ;
  assign n6661 = ( x733 & x734 ) | ( x733 & x735 ) | ( x734 & x735 ) ;
  assign n6662 = ( x733 & ~x734 ) | ( x733 & x735 ) | ( ~x734 & x735 ) ;
  assign n6663 = ( ~x733 & x734 ) | ( ~x733 & n6662 ) | ( x734 & n6662 ) ;
  assign n6664 = ( ~x735 & n6662 ) | ( ~x735 & n6663 ) | ( n6662 & n6663 ) ;
  assign n6665 = ( x736 & ~x737 ) | ( x736 & x738 ) | ( ~x737 & x738 ) ;
  assign n6666 = ( ~x736 & x737 ) | ( ~x736 & n6665 ) | ( x737 & n6665 ) ;
  assign n6667 = ( ~x738 & n6665 ) | ( ~x738 & n6666 ) | ( n6665 & n6666 ) ;
  assign n6668 = n6664 & n6667 ;
  assign n6669 = ( n6660 & n6661 ) | ( n6660 & n6668 ) | ( n6661 & n6668 ) ;
  assign n6670 = ( n6656 & n6658 ) | ( n6656 & ~n6659 ) | ( n6658 & ~n6659 ) ;
  assign n6671 = ( n6657 & ~n6659 ) | ( n6657 & n6670 ) | ( ~n6659 & n6670 ) ;
  assign n6672 = ( n6661 & n6668 ) | ( n6661 & ~n6669 ) | ( n6668 & ~n6669 ) ;
  assign n6673 = ( n6660 & ~n6669 ) | ( n6660 & n6672 ) | ( ~n6669 & n6672 ) ;
  assign n6674 = n6659 & n6671 ;
  assign n6675 = n6669 & n6673 ;
  assign n6676 = n6652 & ~n6655 ;
  assign n6677 = ~n6652 & n6655 ;
  assign n6678 = n6676 | n6677 ;
  assign n6679 = n6664 & ~n6667 ;
  assign n6680 = ~n6664 & n6667 ;
  assign n6681 = n6679 | n6680 ;
  assign n6682 = n6678 & n6681 ;
  assign n6683 = ~n6675 & n6682 ;
  assign n6684 = ~n6674 & n6683 ;
  assign n6685 = ~n6673 & n6684 ;
  assign n6686 = ( n6671 & n6673 ) | ( n6671 & n6685 ) | ( n6673 & n6685 ) ;
  assign n6687 = n6673 & n6683 ;
  assign n6688 = ~n6674 & n6687 ;
  assign n6689 = n6686 | n6688 ;
  assign n6690 = ( n6659 & n6669 ) | ( n6659 & n6689 ) | ( n6669 & n6689 ) ;
  assign n6691 = ~n6659 & n6669 ;
  assign n6692 = n6659 & ~n6669 ;
  assign n6693 = n6691 | n6692 ;
  assign n6694 = n6688 | n6693 ;
  assign n6695 = n6686 | n6694 ;
  assign n6696 = n6689 & n6693 ;
  assign n6697 = n6695 & ~n6696 ;
  assign n6698 = ( n6623 & n6633 ) | ( n6623 & ~n6648 ) | ( n6633 & ~n6648 ) ;
  assign n6699 = ( n6623 & ~n6633 ) | ( n6623 & n6648 ) | ( ~n6633 & n6648 ) ;
  assign n6700 = ( ~n6623 & n6698 ) | ( ~n6623 & n6699 ) | ( n6698 & n6699 ) ;
  assign n6701 = n6697 | n6700 ;
  assign n6702 = ( n6671 & n6673 ) | ( n6671 & ~n6684 ) | ( n6673 & ~n6684 ) ;
  assign n6703 = n6671 & ~n6688 ;
  assign n6704 = ( n6673 & ~n6702 ) | ( n6673 & n6703 ) | ( ~n6702 & n6703 ) ;
  assign n6705 = ( n6685 & n6702 ) | ( n6685 & ~n6704 ) | ( n6702 & ~n6704 ) ;
  assign n6706 = n6641 & ~n6645 ;
  assign n6707 = ~n6641 & n6645 ;
  assign n6708 = n6706 | n6707 ;
  assign n6709 = n6678 & ~n6681 ;
  assign n6710 = ~n6678 & n6681 ;
  assign n6711 = n6709 | n6710 ;
  assign n6712 = n6708 & n6711 ;
  assign n6713 = n6635 | n6647 ;
  assign n6714 = ~n6648 & n6713 ;
  assign n6715 = n6635 & n6646 ;
  assign n6716 = ( n6637 & ~n6713 ) | ( n6637 & n6715 ) | ( ~n6713 & n6715 ) ;
  assign n6717 = n6714 | n6716 ;
  assign n6718 = n6712 | n6717 ;
  assign n6719 = ( n6712 & n6714 ) | ( n6712 & n6716 ) | ( n6714 & n6716 ) ;
  assign n6720 = ( n6705 & n6718 ) | ( n6705 & n6719 ) | ( n6718 & n6719 ) ;
  assign n6721 = n6701 & n6720 ;
  assign n6722 = n6697 & n6700 ;
  assign n6723 = n6721 | n6722 ;
  assign n6724 = ( n6649 & n6690 ) | ( n6649 & n6723 ) | ( n6690 & n6723 ) ;
  assign n6725 = n6613 & n6724 ;
  assign n6726 = ~n6649 & n6690 ;
  assign n6727 = n6649 & ~n6690 ;
  assign n6728 = n6726 | n6727 ;
  assign n6729 = n6722 | n6728 ;
  assign n6730 = n6721 | n6729 ;
  assign n6731 = n6723 & n6728 ;
  assign n6732 = n6730 & ~n6731 ;
  assign n6733 = ~n6540 & n6581 ;
  assign n6734 = n6540 & ~n6581 ;
  assign n6735 = n6733 | n6734 ;
  assign n6736 = n6612 | n6735 ;
  assign n6737 = ~n6735 & n6736 ;
  assign n6738 = ( ~n6612 & n6736 ) | ( ~n6612 & n6737 ) | ( n6736 & n6737 ) ;
  assign n6739 = n6732 | n6738 ;
  assign n6740 = ( n6601 & ~n6608 ) | ( n6601 & n6611 ) | ( ~n6608 & n6611 ) ;
  assign n6741 = ( ~n6601 & n6608 ) | ( ~n6601 & n6740 ) | ( n6608 & n6740 ) ;
  assign n6742 = ( ~n6611 & n6740 ) | ( ~n6611 & n6741 ) | ( n6740 & n6741 ) ;
  assign n6743 = ( ~n6697 & n6700 ) | ( ~n6697 & n6720 ) | ( n6700 & n6720 ) ;
  assign n6744 = ( n6697 & ~n6720 ) | ( n6697 & n6743 ) | ( ~n6720 & n6743 ) ;
  assign n6745 = ( ~n6700 & n6743 ) | ( ~n6700 & n6744 ) | ( n6743 & n6744 ) ;
  assign n6746 = n6708 & ~n6711 ;
  assign n6747 = ~n6708 & n6711 ;
  assign n6748 = n6746 | n6747 ;
  assign n6749 = n6588 & ~n6591 ;
  assign n6750 = ~n6588 & n6591 ;
  assign n6751 = n6749 | n6750 ;
  assign n6752 = n6748 & n6751 ;
  assign n6753 = ~n6712 & n6718 ;
  assign n6754 = ( ~n6717 & n6718 ) | ( ~n6717 & n6753 ) | ( n6718 & n6753 ) ;
  assign n6755 = n6705 & ~n6754 ;
  assign n6756 = ~n6705 & n6754 ;
  assign n6757 = n6755 | n6756 ;
  assign n6758 = ( n6585 & n6592 ) | ( n6585 & ~n6597 ) | ( n6592 & ~n6597 ) ;
  assign n6759 = ( ~n6585 & n6597 ) | ( ~n6585 & n6758 ) | ( n6597 & n6758 ) ;
  assign n6760 = ( ~n6592 & n6758 ) | ( ~n6592 & n6759 ) | ( n6758 & n6759 ) ;
  assign n6761 = ( n6752 & n6757 ) | ( n6752 & n6760 ) | ( n6757 & n6760 ) ;
  assign n6762 = ( n6742 & n6745 ) | ( n6742 & n6761 ) | ( n6745 & n6761 ) ;
  assign n6763 = n6739 & n6762 ;
  assign n6764 = n6732 & n6738 ;
  assign n6765 = n6763 | n6764 ;
  assign n6766 = n6724 & ~n6725 ;
  assign n6767 = ( n6613 & ~n6725 ) | ( n6613 & n6766 ) | ( ~n6725 & n6766 ) ;
  assign n6768 = n6765 & n6767 ;
  assign n6769 = ( n6724 & n6765 ) | ( n6724 & n6768 ) | ( n6765 & n6768 ) ;
  assign n6770 = n6725 | n6769 ;
  assign n6771 = n6505 & n6770 ;
  assign n6772 = n6501 | n6725 ;
  assign n6773 = n6504 | n6772 ;
  assign n6774 = ( n6497 & n6772 ) | ( n6497 & n6773 ) | ( n6772 & n6773 ) ;
  assign n6775 = n6769 | n6774 ;
  assign n6776 = n6496 | n6503 ;
  assign n6777 = n6495 | n6776 ;
  assign n6778 = n6497 & n6503 ;
  assign n6779 = n6777 & ~n6778 ;
  assign n6780 = n6764 | n6767 ;
  assign n6781 = n6763 | n6780 ;
  assign n6782 = ~n6768 & n6781 ;
  assign n6783 = ( ~n6474 & n6477 ) | ( ~n6474 & n6493 ) | ( n6477 & n6493 ) ;
  assign n6784 = ( n6474 & ~n6493 ) | ( n6474 & n6783 ) | ( ~n6493 & n6783 ) ;
  assign n6785 = ( ~n6477 & n6783 ) | ( ~n6477 & n6784 ) | ( n6783 & n6784 ) ;
  assign n6786 = ( ~n6742 & n6745 ) | ( ~n6742 & n6761 ) | ( n6745 & n6761 ) ;
  assign n6787 = ( n6742 & ~n6761 ) | ( n6742 & n6786 ) | ( ~n6761 & n6786 ) ;
  assign n6788 = ( ~n6745 & n6786 ) | ( ~n6745 & n6787 ) | ( n6786 & n6787 ) ;
  assign n6789 = n6748 & ~n6751 ;
  assign n6790 = ~n6748 & n6751 ;
  assign n6791 = n6789 | n6790 ;
  assign n6792 = n6480 & ~n6483 ;
  assign n6793 = ~n6480 & n6483 ;
  assign n6794 = n6792 | n6793 ;
  assign n6795 = n6791 & n6794 ;
  assign n6796 = ( n6752 & ~n6757 ) | ( n6752 & n6760 ) | ( ~n6757 & n6760 ) ;
  assign n6797 = ( ~n6752 & n6757 ) | ( ~n6752 & n6796 ) | ( n6757 & n6796 ) ;
  assign n6798 = ( ~n6760 & n6796 ) | ( ~n6760 & n6797 ) | ( n6796 & n6797 ) ;
  assign n6799 = ( n6484 & ~n6489 ) | ( n6484 & n6492 ) | ( ~n6489 & n6492 ) ;
  assign n6800 = ( ~n6484 & n6489 ) | ( ~n6484 & n6799 ) | ( n6489 & n6799 ) ;
  assign n6801 = ( ~n6492 & n6799 ) | ( ~n6492 & n6800 ) | ( n6799 & n6800 ) ;
  assign n6802 = ( n6795 & n6798 ) | ( n6795 & n6801 ) | ( n6798 & n6801 ) ;
  assign n6803 = ( n6785 & n6788 ) | ( n6785 & n6802 ) | ( n6788 & n6802 ) ;
  assign n6804 = ( ~n6732 & n6738 ) | ( ~n6732 & n6762 ) | ( n6738 & n6762 ) ;
  assign n6805 = ( n6732 & ~n6762 ) | ( n6732 & n6804 ) | ( ~n6762 & n6804 ) ;
  assign n6806 = ( ~n6738 & n6804 ) | ( ~n6738 & n6805 ) | ( n6804 & n6805 ) ;
  assign n6807 = ( ~n6354 & n6470 ) | ( ~n6354 & n6494 ) | ( n6470 & n6494 ) ;
  assign n6808 = ( n6354 & ~n6494 ) | ( n6354 & n6807 ) | ( ~n6494 & n6807 ) ;
  assign n6809 = ( ~n6470 & n6807 ) | ( ~n6470 & n6808 ) | ( n6807 & n6808 ) ;
  assign n6810 = ( n6803 & n6806 ) | ( n6803 & n6809 ) | ( n6806 & n6809 ) ;
  assign n6811 = ( n6779 & n6782 ) | ( n6779 & n6810 ) | ( n6782 & n6810 ) ;
  assign n6812 = ( n6771 & n6775 ) | ( n6771 & n6811 ) | ( n6775 & n6811 ) ;
  assign n6813 = ( x778 & x779 ) | ( x778 & x780 ) | ( x779 & x780 ) ;
  assign n6814 = ( x775 & ~x776 ) | ( x775 & x777 ) | ( ~x776 & x777 ) ;
  assign n6815 = ( ~x775 & x776 ) | ( ~x775 & n6814 ) | ( x776 & n6814 ) ;
  assign n6816 = ( ~x777 & n6814 ) | ( ~x777 & n6815 ) | ( n6814 & n6815 ) ;
  assign n6817 = ( x778 & ~x779 ) | ( x778 & x780 ) | ( ~x779 & x780 ) ;
  assign n6818 = ( ~x778 & x779 ) | ( ~x778 & n6817 ) | ( x779 & n6817 ) ;
  assign n6819 = ( ~x780 & n6817 ) | ( ~x780 & n6818 ) | ( n6817 & n6818 ) ;
  assign n6820 = n6816 & n6819 ;
  assign n6821 = ( x775 & x776 ) | ( x775 & x777 ) | ( x776 & x777 ) ;
  assign n6822 = ( n6813 & n6820 ) | ( n6813 & n6821 ) | ( n6820 & n6821 ) ;
  assign n6823 = ( n6820 & n6821 ) | ( n6820 & ~n6822 ) | ( n6821 & ~n6822 ) ;
  assign n6824 = ( n6813 & ~n6822 ) | ( n6813 & n6823 ) | ( ~n6822 & n6823 ) ;
  assign n6825 = ( x784 & x785 ) | ( x784 & x786 ) | ( x785 & x786 ) ;
  assign n6826 = ( x781 & x782 ) | ( x781 & x783 ) | ( x782 & x783 ) ;
  assign n6827 = ( x781 & ~x782 ) | ( x781 & x783 ) | ( ~x782 & x783 ) ;
  assign n6828 = ( ~x781 & x782 ) | ( ~x781 & n6827 ) | ( x782 & n6827 ) ;
  assign n6829 = ( ~x783 & n6827 ) | ( ~x783 & n6828 ) | ( n6827 & n6828 ) ;
  assign n6830 = ( x784 & ~x785 ) | ( x784 & x786 ) | ( ~x785 & x786 ) ;
  assign n6831 = ( ~x784 & x785 ) | ( ~x784 & n6830 ) | ( x785 & n6830 ) ;
  assign n6832 = ( ~x786 & n6830 ) | ( ~x786 & n6831 ) | ( n6830 & n6831 ) ;
  assign n6833 = n6829 & n6832 ;
  assign n6834 = ( n6825 & n6826 ) | ( n6825 & n6833 ) | ( n6826 & n6833 ) ;
  assign n6835 = ( n6826 & n6833 ) | ( n6826 & ~n6834 ) | ( n6833 & ~n6834 ) ;
  assign n6836 = ( n6825 & ~n6834 ) | ( n6825 & n6835 ) | ( ~n6834 & n6835 ) ;
  assign n6837 = n6822 & n6824 ;
  assign n6838 = n6834 & n6836 ;
  assign n6839 = n6816 & ~n6819 ;
  assign n6840 = ~n6816 & n6819 ;
  assign n6841 = n6839 | n6840 ;
  assign n6842 = n6829 & ~n6832 ;
  assign n6843 = ~n6829 & n6832 ;
  assign n6844 = n6842 | n6843 ;
  assign n6845 = n6841 & n6844 ;
  assign n6846 = ~n6838 & n6845 ;
  assign n6847 = ~n6837 & n6846 ;
  assign n6848 = ~n6836 & n6847 ;
  assign n6849 = ( n6824 & n6836 ) | ( n6824 & n6848 ) | ( n6836 & n6848 ) ;
  assign n6850 = n6836 & n6846 ;
  assign n6851 = ~n6837 & n6850 ;
  assign n6852 = ~n6822 & n6834 ;
  assign n6853 = n6822 & ~n6834 ;
  assign n6854 = n6852 | n6853 ;
  assign n6855 = n6851 | n6854 ;
  assign n6856 = n6849 | n6855 ;
  assign n6857 = n6849 | n6851 ;
  assign n6858 = n6854 & n6857 ;
  assign n6859 = n6856 & ~n6858 ;
  assign n6860 = ( x796 & x797 ) | ( x796 & x798 ) | ( x797 & x798 ) ;
  assign n6861 = ( x793 & x794 ) | ( x793 & x795 ) | ( x794 & x795 ) ;
  assign n6862 = ( x793 & ~x794 ) | ( x793 & x795 ) | ( ~x794 & x795 ) ;
  assign n6863 = ( ~x793 & x794 ) | ( ~x793 & n6862 ) | ( x794 & n6862 ) ;
  assign n6864 = ( ~x795 & n6862 ) | ( ~x795 & n6863 ) | ( n6862 & n6863 ) ;
  assign n6865 = ( x796 & ~x797 ) | ( x796 & x798 ) | ( ~x797 & x798 ) ;
  assign n6866 = ( ~x796 & x797 ) | ( ~x796 & n6865 ) | ( x797 & n6865 ) ;
  assign n6867 = ( ~x798 & n6865 ) | ( ~x798 & n6866 ) | ( n6865 & n6866 ) ;
  assign n6868 = n6864 & n6867 ;
  assign n6869 = ( n6860 & n6861 ) | ( n6860 & n6868 ) | ( n6861 & n6868 ) ;
  assign n6870 = ( x787 & ~x788 ) | ( x787 & x789 ) | ( ~x788 & x789 ) ;
  assign n6871 = ( ~x787 & x788 ) | ( ~x787 & n6870 ) | ( x788 & n6870 ) ;
  assign n6872 = ( ~x789 & n6870 ) | ( ~x789 & n6871 ) | ( n6870 & n6871 ) ;
  assign n6873 = ( x790 & ~x791 ) | ( x790 & x792 ) | ( ~x791 & x792 ) ;
  assign n6874 = ( ~x790 & x791 ) | ( ~x790 & n6873 ) | ( x791 & n6873 ) ;
  assign n6875 = ( ~x792 & n6873 ) | ( ~x792 & n6874 ) | ( n6873 & n6874 ) ;
  assign n6876 = n6872 & n6875 ;
  assign n6877 = ( x790 & x791 ) | ( x790 & x792 ) | ( x791 & x792 ) ;
  assign n6878 = ( x787 & x788 ) | ( x787 & x789 ) | ( x788 & x789 ) ;
  assign n6879 = ( n6876 & n6877 ) | ( n6876 & n6878 ) | ( n6877 & n6878 ) ;
  assign n6880 = ( n6861 & n6868 ) | ( n6861 & ~n6869 ) | ( n6868 & ~n6869 ) ;
  assign n6881 = ( n6860 & ~n6869 ) | ( n6860 & n6880 ) | ( ~n6869 & n6880 ) ;
  assign n6882 = ( n6876 & n6878 ) | ( n6876 & ~n6879 ) | ( n6878 & ~n6879 ) ;
  assign n6883 = ( n6877 & ~n6879 ) | ( n6877 & n6882 ) | ( ~n6879 & n6882 ) ;
  assign n6884 = n6879 & n6883 ;
  assign n6885 = n6872 & ~n6875 ;
  assign n6886 = ~n6872 & n6875 ;
  assign n6887 = n6885 | n6886 ;
  assign n6888 = n6864 & ~n6867 ;
  assign n6889 = ~n6864 & n6867 ;
  assign n6890 = n6888 | n6889 ;
  assign n6891 = ~n6868 & n6890 ;
  assign n6892 = n6887 & n6891 ;
  assign n6893 = ~n6884 & n6892 ;
  assign n6894 = ( n6881 & n6883 ) | ( n6881 & n6893 ) | ( n6883 & n6893 ) ;
  assign n6895 = ( n6869 & n6879 ) | ( n6869 & ~n6894 ) | ( n6879 & ~n6894 ) ;
  assign n6896 = ( n6869 & ~n6879 ) | ( n6869 & n6894 ) | ( ~n6879 & n6894 ) ;
  assign n6897 = ( ~n6869 & n6895 ) | ( ~n6869 & n6896 ) | ( n6895 & n6896 ) ;
  assign n6898 = n6859 | n6897 ;
  assign n6899 = ( n6824 & n6836 ) | ( n6824 & ~n6847 ) | ( n6836 & ~n6847 ) ;
  assign n6900 = n6824 & ~n6851 ;
  assign n6901 = ( n6836 & ~n6899 ) | ( n6836 & n6900 ) | ( ~n6899 & n6900 ) ;
  assign n6902 = ( n6848 & n6899 ) | ( n6848 & ~n6901 ) | ( n6899 & ~n6901 ) ;
  assign n6903 = n6887 & ~n6891 ;
  assign n6904 = ~n6887 & n6891 ;
  assign n6905 = n6903 | n6904 ;
  assign n6906 = n6841 & ~n6844 ;
  assign n6907 = ~n6841 & n6844 ;
  assign n6908 = n6906 | n6907 ;
  assign n6909 = n6905 & n6908 ;
  assign n6910 = n6881 | n6893 ;
  assign n6911 = ~n6894 & n6910 ;
  assign n6912 = n6881 & n6892 ;
  assign n6913 = ( n6883 & ~n6910 ) | ( n6883 & n6912 ) | ( ~n6910 & n6912 ) ;
  assign n6914 = n6911 | n6913 ;
  assign n6915 = n6909 | n6914 ;
  assign n6916 = ( n6909 & n6911 ) | ( n6909 & n6913 ) | ( n6911 & n6913 ) ;
  assign n6917 = ( n6902 & n6915 ) | ( n6902 & n6916 ) | ( n6915 & n6916 ) ;
  assign n6918 = n6898 & n6917 ;
  assign n6919 = n6859 & n6897 ;
  assign n6920 = ( n6869 & n6879 ) | ( n6869 & n6894 ) | ( n6879 & n6894 ) ;
  assign n6921 = ( n6822 & n6834 ) | ( n6822 & n6857 ) | ( n6834 & n6857 ) ;
  assign n6922 = ~n6920 & n6921 ;
  assign n6923 = n6920 & ~n6921 ;
  assign n6924 = n6922 | n6923 ;
  assign n6925 = n6919 | n6924 ;
  assign n6926 = n6918 | n6925 ;
  assign n6927 = n6918 | n6919 ;
  assign n6928 = n6924 & n6927 ;
  assign n6929 = n6926 & ~n6928 ;
  assign n6965 = ( x760 & x761 ) | ( x760 & x762 ) | ( x761 & x762 ) ;
  assign n6966 = ( x757 & x758 ) | ( x757 & x759 ) | ( x758 & x759 ) ;
  assign n6967 = ( x757 & ~x758 ) | ( x757 & x759 ) | ( ~x758 & x759 ) ;
  assign n6968 = ( ~x757 & x758 ) | ( ~x757 & n6967 ) | ( x758 & n6967 ) ;
  assign n6969 = ( ~x759 & n6967 ) | ( ~x759 & n6968 ) | ( n6967 & n6968 ) ;
  assign n6970 = ( x760 & ~x761 ) | ( x760 & x762 ) | ( ~x761 & x762 ) ;
  assign n6971 = ( ~x760 & x761 ) | ( ~x760 & n6970 ) | ( x761 & n6970 ) ;
  assign n6972 = ( ~x762 & n6970 ) | ( ~x762 & n6971 ) | ( n6970 & n6971 ) ;
  assign n6973 = n6969 & n6972 ;
  assign n6974 = ( n6965 & n6966 ) | ( n6965 & n6973 ) | ( n6966 & n6973 ) ;
  assign n6988 = ( n6966 & n6973 ) | ( n6966 & ~n6974 ) | ( n6973 & ~n6974 ) ;
  assign n6989 = ( n6965 & ~n6974 ) | ( n6965 & n6988 ) | ( ~n6974 & n6988 ) ;
  assign n6975 = ( x754 & x755 ) | ( x754 & x756 ) | ( x755 & x756 ) ;
  assign n6976 = ( x751 & x752 ) | ( x751 & x753 ) | ( x752 & x753 ) ;
  assign n6977 = ( x751 & ~x752 ) | ( x751 & x753 ) | ( ~x752 & x753 ) ;
  assign n6978 = ( ~x751 & x752 ) | ( ~x751 & n6977 ) | ( x752 & n6977 ) ;
  assign n6979 = ( ~x753 & n6977 ) | ( ~x753 & n6978 ) | ( n6977 & n6978 ) ;
  assign n6980 = ( x754 & ~x755 ) | ( x754 & x756 ) | ( ~x755 & x756 ) ;
  assign n6981 = ( ~x754 & x755 ) | ( ~x754 & n6980 ) | ( x755 & n6980 ) ;
  assign n6982 = ( ~x756 & n6980 ) | ( ~x756 & n6981 ) | ( n6980 & n6981 ) ;
  assign n6983 = n6979 & n6982 ;
  assign n6984 = ( n6975 & n6976 ) | ( n6975 & n6983 ) | ( n6976 & n6983 ) ;
  assign n6985 = ( n6976 & n6983 ) | ( n6976 & ~n6984 ) | ( n6983 & ~n6984 ) ;
  assign n6986 = ( n6975 & ~n6984 ) | ( n6975 & n6985 ) | ( ~n6984 & n6985 ) ;
  assign n6987 = n6984 & n6986 ;
  assign n6990 = n6974 & n6989 ;
  assign n6991 = n6969 & ~n6972 ;
  assign n6992 = ~n6969 & n6972 ;
  assign n6993 = n6991 | n6992 ;
  assign n6994 = n6979 & ~n6982 ;
  assign n6995 = ~n6979 & n6982 ;
  assign n6996 = n6994 | n6995 ;
  assign n6997 = n6993 & n6996 ;
  assign n6998 = ~n6990 & n6997 ;
  assign n7001 = ~n6987 & n6998 ;
  assign n7002 = ~n6989 & n7001 ;
  assign n7009 = ( n6986 & n6989 ) | ( n6986 & ~n7001 ) | ( n6989 & ~n7001 ) ;
  assign n6999 = n6989 & n6998 ;
  assign n7000 = ~n6987 & n6999 ;
  assign n7010 = n6986 & ~n7000 ;
  assign n7011 = ( n6989 & ~n7009 ) | ( n6989 & n7010 ) | ( ~n7009 & n7010 ) ;
  assign n7012 = ( n7002 & n7009 ) | ( n7002 & ~n7011 ) | ( n7009 & ~n7011 ) ;
  assign n6932 = ( x763 & ~x764 ) | ( x763 & x765 ) | ( ~x764 & x765 ) ;
  assign n6933 = ( ~x763 & x764 ) | ( ~x763 & n6932 ) | ( x764 & n6932 ) ;
  assign n6934 = ( ~x765 & n6932 ) | ( ~x765 & n6933 ) | ( n6932 & n6933 ) ;
  assign n6935 = ( x766 & ~x767 ) | ( x766 & x768 ) | ( ~x767 & x768 ) ;
  assign n6936 = ( ~x766 & x767 ) | ( ~x766 & n6935 ) | ( x767 & n6935 ) ;
  assign n6937 = ( ~x768 & n6935 ) | ( ~x768 & n6936 ) | ( n6935 & n6936 ) ;
  assign n6955 = n6934 & ~n6937 ;
  assign n6956 = ~n6934 & n6937 ;
  assign n6957 = n6955 | n6956 ;
  assign n6942 = ( x769 & ~x770 ) | ( x769 & x771 ) | ( ~x770 & x771 ) ;
  assign n6943 = ( ~x769 & x770 ) | ( ~x769 & n6942 ) | ( x770 & n6942 ) ;
  assign n6944 = ( ~x771 & n6942 ) | ( ~x771 & n6943 ) | ( n6942 & n6943 ) ;
  assign n6945 = ( x772 & ~x773 ) | ( x772 & x774 ) | ( ~x773 & x774 ) ;
  assign n6946 = ( ~x772 & x773 ) | ( ~x772 & n6945 ) | ( x773 & n6945 ) ;
  assign n6947 = ( ~x774 & n6945 ) | ( ~x774 & n6946 ) | ( n6945 & n6946 ) ;
  assign n6958 = n6944 & ~n6947 ;
  assign n6959 = ~n6944 & n6947 ;
  assign n6960 = n6958 | n6959 ;
  assign n7013 = n6957 & ~n6960 ;
  assign n7014 = ~n6957 & n6960 ;
  assign n7015 = n7013 | n7014 ;
  assign n7016 = ~n6993 & n6996 ;
  assign n7017 = n6993 & ~n6996 ;
  assign n7018 = n7016 | n7017 ;
  assign n7019 = n7015 & n7018 ;
  assign n6930 = ( x766 & x767 ) | ( x766 & x768 ) | ( x767 & x768 ) ;
  assign n6931 = ( x763 & x764 ) | ( x763 & x765 ) | ( x764 & x765 ) ;
  assign n6938 = n6934 & n6937 ;
  assign n6939 = ( n6930 & n6931 ) | ( n6930 & n6938 ) | ( n6931 & n6938 ) ;
  assign n6950 = ( n6931 & n6938 ) | ( n6931 & ~n6939 ) | ( n6938 & ~n6939 ) ;
  assign n6951 = ( n6930 & ~n6939 ) | ( n6930 & n6950 ) | ( ~n6939 & n6950 ) ;
  assign n6940 = ( x772 & x773 ) | ( x772 & x774 ) | ( x773 & x774 ) ;
  assign n6941 = ( x769 & x770 ) | ( x769 & x771 ) | ( x770 & x771 ) ;
  assign n6948 = n6944 & n6947 ;
  assign n6949 = ( n6940 & n6941 ) | ( n6940 & n6948 ) | ( n6941 & n6948 ) ;
  assign n6952 = ( n6941 & n6948 ) | ( n6941 & ~n6949 ) | ( n6948 & ~n6949 ) ;
  assign n6953 = ( n6940 & ~n6949 ) | ( n6940 & n6952 ) | ( ~n6949 & n6952 ) ;
  assign n6961 = n6957 & n6960 ;
  assign n7020 = n6953 & n6961 ;
  assign n6954 = n6939 & n6951 ;
  assign n6962 = ~n6954 & n6961 ;
  assign n7021 = n6953 | n6962 ;
  assign n7022 = ( n6951 & n7020 ) | ( n6951 & ~n7021 ) | ( n7020 & ~n7021 ) ;
  assign n6963 = ( n6951 & n6953 ) | ( n6951 & n6962 ) | ( n6953 & n6962 ) ;
  assign n7023 = ~n6963 & n7021 ;
  assign n7024 = n7022 | n7023 ;
  assign n7025 = n7019 | n7024 ;
  assign n7026 = n7012 & n7025 ;
  assign n7027 = ( n7019 & n7022 ) | ( n7019 & n7023 ) | ( n7022 & n7023 ) ;
  assign n7028 = n7026 | n7027 ;
  assign n7003 = ( n6986 & n6989 ) | ( n6986 & n7002 ) | ( n6989 & n7002 ) ;
  assign n7029 = n6974 & ~n6984 ;
  assign n7030 = ~n6974 & n6984 ;
  assign n7031 = n7029 | n7030 ;
  assign n7032 = n7000 | n7031 ;
  assign n7033 = n7003 | n7032 ;
  assign n7004 = n7000 | n7003 ;
  assign n7034 = n7004 & n7031 ;
  assign n7035 = n7033 & ~n7034 ;
  assign n7036 = ~n6939 & n6949 ;
  assign n7037 = n6939 & ~n6949 ;
  assign n7038 = n7036 | n7037 ;
  assign n7039 = n6963 & n7038 ;
  assign n7040 = n6963 | n7038 ;
  assign n7041 = ~n7039 & n7040 ;
  assign n7042 = ( n7028 & n7035 ) | ( n7028 & n7041 ) | ( n7035 & n7041 ) ;
  assign n6964 = ( n6939 & n6949 ) | ( n6939 & n6963 ) | ( n6949 & n6963 ) ;
  assign n7005 = ( n6974 & n6984 ) | ( n6974 & n7004 ) | ( n6984 & n7004 ) ;
  assign n7006 = n6964 & n7005 ;
  assign n7007 = n7005 & ~n7006 ;
  assign n7008 = ( n6964 & ~n7006 ) | ( n6964 & n7007 ) | ( ~n7006 & n7007 ) ;
  assign n7043 = n7008 | n7042 ;
  assign n7044 = ~n7008 & n7043 ;
  assign n7045 = ( ~n7042 & n7043 ) | ( ~n7042 & n7044 ) | ( n7043 & n7044 ) ;
  assign n7046 = n6929 | n7045 ;
  assign n7047 = ( n7028 & ~n7035 ) | ( n7028 & n7041 ) | ( ~n7035 & n7041 ) ;
  assign n7048 = ( ~n7028 & n7035 ) | ( ~n7028 & n7047 ) | ( n7035 & n7047 ) ;
  assign n7049 = ( ~n7041 & n7047 ) | ( ~n7041 & n7048 ) | ( n7047 & n7048 ) ;
  assign n7050 = ( ~n6859 & n6897 ) | ( ~n6859 & n6917 ) | ( n6897 & n6917 ) ;
  assign n7051 = ( n6859 & ~n6917 ) | ( n6859 & n7050 ) | ( ~n6917 & n7050 ) ;
  assign n7052 = ( ~n6897 & n7050 ) | ( ~n6897 & n7051 ) | ( n7050 & n7051 ) ;
  assign n7053 = n6905 & ~n6908 ;
  assign n7054 = ~n6905 & n6908 ;
  assign n7055 = n7053 | n7054 ;
  assign n7056 = n7015 & ~n7018 ;
  assign n7057 = ~n7015 & n7018 ;
  assign n7058 = n7056 | n7057 ;
  assign n7059 = n7055 & n7058 ;
  assign n7060 = ~n6909 & n6915 ;
  assign n7061 = ( ~n6914 & n6915 ) | ( ~n6914 & n7060 ) | ( n6915 & n7060 ) ;
  assign n7062 = n6902 & ~n7061 ;
  assign n7063 = ~n6902 & n7061 ;
  assign n7064 = n7062 | n7063 ;
  assign n7065 = ( n7012 & n7019 ) | ( n7012 & ~n7024 ) | ( n7019 & ~n7024 ) ;
  assign n7066 = ( ~n7012 & n7024 ) | ( ~n7012 & n7065 ) | ( n7024 & n7065 ) ;
  assign n7067 = ( ~n7019 & n7065 ) | ( ~n7019 & n7066 ) | ( n7065 & n7066 ) ;
  assign n7068 = ( n7059 & n7064 ) | ( n7059 & n7067 ) | ( n7064 & n7067 ) ;
  assign n7069 = ( n7049 & n7052 ) | ( n7049 & n7068 ) | ( n7052 & n7068 ) ;
  assign n7070 = n7046 & n7069 ;
  assign n7071 = n6929 & n7045 ;
  assign n7072 = n7070 | n7071 ;
  assign n7073 = n7006 | n7008 ;
  assign n7074 = ( n7006 & n7042 ) | ( n7006 & n7073 ) | ( n7042 & n7073 ) ;
  assign n7075 = ( n6920 & n6921 ) | ( n6920 & n6927 ) | ( n6921 & n6927 ) ;
  assign n7076 = n7074 & n7075 ;
  assign n7077 = n7075 & ~n7076 ;
  assign n7078 = ( n7074 & ~n7076 ) | ( n7074 & n7077 ) | ( ~n7076 & n7077 ) ;
  assign n7079 = ( n7073 & n7075 ) | ( n7073 & n7078 ) | ( n7075 & n7078 ) ;
  assign n7080 = ( n7072 & n7076 ) | ( n7072 & n7079 ) | ( n7076 & n7079 ) ;
  assign n7081 = ( x820 & x821 ) | ( x820 & x822 ) | ( x821 & x822 ) ;
  assign n7082 = ( x817 & x818 ) | ( x817 & x819 ) | ( x818 & x819 ) ;
  assign n7083 = ( x817 & ~x818 ) | ( x817 & x819 ) | ( ~x818 & x819 ) ;
  assign n7084 = ( ~x817 & x818 ) | ( ~x817 & n7083 ) | ( x818 & n7083 ) ;
  assign n7085 = ( ~x819 & n7083 ) | ( ~x819 & n7084 ) | ( n7083 & n7084 ) ;
  assign n7086 = ( x820 & ~x821 ) | ( x820 & x822 ) | ( ~x821 & x822 ) ;
  assign n7087 = ( ~x820 & x821 ) | ( ~x820 & n7086 ) | ( x821 & n7086 ) ;
  assign n7088 = ( ~x822 & n7086 ) | ( ~x822 & n7087 ) | ( n7086 & n7087 ) ;
  assign n7089 = n7085 & n7088 ;
  assign n7090 = ( n7081 & n7082 ) | ( n7081 & n7089 ) | ( n7082 & n7089 ) ;
  assign n7091 = ( x811 & ~x812 ) | ( x811 & x813 ) | ( ~x812 & x813 ) ;
  assign n7092 = ( ~x811 & x812 ) | ( ~x811 & n7091 ) | ( x812 & n7091 ) ;
  assign n7093 = ( ~x813 & n7091 ) | ( ~x813 & n7092 ) | ( n7091 & n7092 ) ;
  assign n7094 = ( x814 & ~x815 ) | ( x814 & x816 ) | ( ~x815 & x816 ) ;
  assign n7095 = ( ~x814 & x815 ) | ( ~x814 & n7094 ) | ( x815 & n7094 ) ;
  assign n7096 = ( ~x816 & n7094 ) | ( ~x816 & n7095 ) | ( n7094 & n7095 ) ;
  assign n7097 = n7093 & n7096 ;
  assign n7098 = ( x814 & x815 ) | ( x814 & x816 ) | ( x815 & x816 ) ;
  assign n7099 = ( x811 & x812 ) | ( x811 & x813 ) | ( x812 & x813 ) ;
  assign n7100 = ( n7097 & n7098 ) | ( n7097 & n7099 ) | ( n7098 & n7099 ) ;
  assign n7101 = ( n7082 & n7089 ) | ( n7082 & ~n7090 ) | ( n7089 & ~n7090 ) ;
  assign n7102 = ( n7081 & ~n7090 ) | ( n7081 & n7101 ) | ( ~n7090 & n7101 ) ;
  assign n7103 = ( n7097 & n7099 ) | ( n7097 & ~n7100 ) | ( n7099 & ~n7100 ) ;
  assign n7104 = ( n7098 & ~n7100 ) | ( n7098 & n7103 ) | ( ~n7100 & n7103 ) ;
  assign n7105 = n7100 & n7104 ;
  assign n7106 = n7085 & ~n7088 ;
  assign n7107 = ~n7085 & n7088 ;
  assign n7108 = n7106 | n7107 ;
  assign n7109 = n7093 & ~n7096 ;
  assign n7110 = ~n7093 & n7096 ;
  assign n7111 = n7109 | n7110 ;
  assign n7112 = n7108 & n7111 ;
  assign n7113 = ~n7105 & n7112 ;
  assign n7114 = ( n7102 & n7104 ) | ( n7102 & n7113 ) | ( n7104 & n7113 ) ;
  assign n7115 = ( n7090 & n7100 ) | ( n7090 & n7114 ) | ( n7100 & n7114 ) ;
  assign n7116 = ( x808 & x809 ) | ( x808 & x810 ) | ( x809 & x810 ) ;
  assign n7117 = ( x805 & x806 ) | ( x805 & x807 ) | ( x806 & x807 ) ;
  assign n7118 = ( x805 & ~x806 ) | ( x805 & x807 ) | ( ~x806 & x807 ) ;
  assign n7119 = ( ~x805 & x806 ) | ( ~x805 & n7118 ) | ( x806 & n7118 ) ;
  assign n7120 = ( ~x807 & n7118 ) | ( ~x807 & n7119 ) | ( n7118 & n7119 ) ;
  assign n7121 = ( x808 & ~x809 ) | ( x808 & x810 ) | ( ~x809 & x810 ) ;
  assign n7122 = ( ~x808 & x809 ) | ( ~x808 & n7121 ) | ( x809 & n7121 ) ;
  assign n7123 = ( ~x810 & n7121 ) | ( ~x810 & n7122 ) | ( n7121 & n7122 ) ;
  assign n7124 = n7120 & n7123 ;
  assign n7125 = ( n7116 & n7117 ) | ( n7116 & n7124 ) | ( n7117 & n7124 ) ;
  assign n7126 = ( x802 & x803 ) | ( x802 & x804 ) | ( x803 & x804 ) ;
  assign n7127 = ( x799 & x800 ) | ( x799 & x801 ) | ( x800 & x801 ) ;
  assign n7128 = ( x799 & ~x800 ) | ( x799 & x801 ) | ( ~x800 & x801 ) ;
  assign n7129 = ( ~x799 & x800 ) | ( ~x799 & n7128 ) | ( x800 & n7128 ) ;
  assign n7130 = ( ~x801 & n7128 ) | ( ~x801 & n7129 ) | ( n7128 & n7129 ) ;
  assign n7131 = ( x802 & ~x803 ) | ( x802 & x804 ) | ( ~x803 & x804 ) ;
  assign n7132 = ( ~x802 & x803 ) | ( ~x802 & n7131 ) | ( x803 & n7131 ) ;
  assign n7133 = ( ~x804 & n7131 ) | ( ~x804 & n7132 ) | ( n7131 & n7132 ) ;
  assign n7134 = n7130 & n7133 ;
  assign n7135 = ( n7126 & n7127 ) | ( n7126 & n7134 ) | ( n7127 & n7134 ) ;
  assign n7136 = ( n7127 & n7134 ) | ( n7127 & ~n7135 ) | ( n7134 & ~n7135 ) ;
  assign n7137 = ( n7126 & ~n7135 ) | ( n7126 & n7136 ) | ( ~n7135 & n7136 ) ;
  assign n7138 = n7135 & n7137 ;
  assign n7139 = ( n7117 & n7124 ) | ( n7117 & ~n7125 ) | ( n7124 & ~n7125 ) ;
  assign n7140 = ( n7116 & ~n7125 ) | ( n7116 & n7139 ) | ( ~n7125 & n7139 ) ;
  assign n7141 = n7125 & n7140 ;
  assign n7142 = n7120 & ~n7123 ;
  assign n7143 = ~n7120 & n7123 ;
  assign n7144 = n7142 | n7143 ;
  assign n7145 = n7130 & ~n7133 ;
  assign n7146 = ~n7130 & n7133 ;
  assign n7147 = n7145 | n7146 ;
  assign n7148 = n7144 & n7147 ;
  assign n7149 = ~n7141 & n7148 ;
  assign n7150 = n7140 & n7149 ;
  assign n7151 = ~n7138 & n7150 ;
  assign n7152 = ~n7138 & n7149 ;
  assign n7153 = ~n7140 & n7152 ;
  assign n7154 = ( n7137 & n7140 ) | ( n7137 & n7153 ) | ( n7140 & n7153 ) ;
  assign n7155 = n7151 | n7154 ;
  assign n7156 = ( n7125 & n7135 ) | ( n7125 & n7155 ) | ( n7135 & n7155 ) ;
  assign n7157 = ( n7137 & n7140 ) | ( n7137 & ~n7152 ) | ( n7140 & ~n7152 ) ;
  assign n7158 = n7137 & ~n7151 ;
  assign n7159 = ( n7140 & ~n7157 ) | ( n7140 & n7158 ) | ( ~n7157 & n7158 ) ;
  assign n7160 = ( n7153 & n7157 ) | ( n7153 & ~n7159 ) | ( n7157 & ~n7159 ) ;
  assign n7161 = ~n7108 & n7111 ;
  assign n7162 = n7108 & ~n7111 ;
  assign n7163 = n7161 | n7162 ;
  assign n7164 = ~n7144 & n7147 ;
  assign n7165 = n7144 & ~n7147 ;
  assign n7166 = n7164 | n7165 ;
  assign n7167 = n7163 & n7166 ;
  assign n7168 = n7102 & n7112 ;
  assign n7169 = n7102 | n7113 ;
  assign n7170 = ( n7104 & n7168 ) | ( n7104 & ~n7169 ) | ( n7168 & ~n7169 ) ;
  assign n7171 = ~n7114 & n7169 ;
  assign n7172 = n7170 | n7171 ;
  assign n7173 = n7167 | n7172 ;
  assign n7174 = n7160 & n7173 ;
  assign n7175 = ( n7167 & n7170 ) | ( n7167 & n7171 ) | ( n7170 & n7171 ) ;
  assign n7176 = n7174 | n7175 ;
  assign n7177 = n7125 & ~n7135 ;
  assign n7178 = ~n7125 & n7135 ;
  assign n7179 = n7177 | n7178 ;
  assign n7180 = n7151 | n7179 ;
  assign n7181 = n7154 | n7180 ;
  assign n7182 = n7155 & n7179 ;
  assign n7183 = n7181 & ~n7182 ;
  assign n7184 = ( n7090 & n7100 ) | ( n7090 & ~n7114 ) | ( n7100 & ~n7114 ) ;
  assign n7185 = ( n7090 & ~n7100 ) | ( n7090 & n7114 ) | ( ~n7100 & n7114 ) ;
  assign n7186 = ( ~n7090 & n7184 ) | ( ~n7090 & n7185 ) | ( n7184 & n7185 ) ;
  assign n7187 = ( n7176 & n7183 ) | ( n7176 & n7186 ) | ( n7183 & n7186 ) ;
  assign n7188 = ( n7115 & n7156 ) | ( n7115 & n7187 ) | ( n7156 & n7187 ) ;
  assign n7189 = ( x844 & x845 ) | ( x844 & x846 ) | ( x845 & x846 ) ;
  assign n7190 = ( x841 & x842 ) | ( x841 & x843 ) | ( x842 & x843 ) ;
  assign n7191 = ( x841 & ~x842 ) | ( x841 & x843 ) | ( ~x842 & x843 ) ;
  assign n7192 = ( ~x841 & x842 ) | ( ~x841 & n7191 ) | ( x842 & n7191 ) ;
  assign n7193 = ( ~x843 & n7191 ) | ( ~x843 & n7192 ) | ( n7191 & n7192 ) ;
  assign n7194 = ( x844 & ~x845 ) | ( x844 & x846 ) | ( ~x845 & x846 ) ;
  assign n7195 = ( ~x844 & x845 ) | ( ~x844 & n7194 ) | ( x845 & n7194 ) ;
  assign n7196 = ( ~x846 & n7194 ) | ( ~x846 & n7195 ) | ( n7194 & n7195 ) ;
  assign n7197 = n7193 & n7196 ;
  assign n7198 = ( n7189 & n7190 ) | ( n7189 & n7197 ) | ( n7190 & n7197 ) ;
  assign n7199 = ( x835 & ~x836 ) | ( x835 & x837 ) | ( ~x836 & x837 ) ;
  assign n7200 = ( ~x835 & x836 ) | ( ~x835 & n7199 ) | ( x836 & n7199 ) ;
  assign n7201 = ( ~x837 & n7199 ) | ( ~x837 & n7200 ) | ( n7199 & n7200 ) ;
  assign n7202 = ( x838 & ~x839 ) | ( x838 & x840 ) | ( ~x839 & x840 ) ;
  assign n7203 = ( ~x838 & x839 ) | ( ~x838 & n7202 ) | ( x839 & n7202 ) ;
  assign n7204 = ( ~x840 & n7202 ) | ( ~x840 & n7203 ) | ( n7202 & n7203 ) ;
  assign n7205 = n7201 & n7204 ;
  assign n7206 = ( x838 & x839 ) | ( x838 & x840 ) | ( x839 & x840 ) ;
  assign n7207 = ( x835 & x836 ) | ( x835 & x837 ) | ( x836 & x837 ) ;
  assign n7208 = ( n7205 & n7206 ) | ( n7205 & n7207 ) | ( n7206 & n7207 ) ;
  assign n7209 = ( n7190 & n7197 ) | ( n7190 & ~n7198 ) | ( n7197 & ~n7198 ) ;
  assign n7210 = ( n7189 & ~n7198 ) | ( n7189 & n7209 ) | ( ~n7198 & n7209 ) ;
  assign n7211 = ( n7205 & n7207 ) | ( n7205 & ~n7208 ) | ( n7207 & ~n7208 ) ;
  assign n7212 = ( n7206 & ~n7208 ) | ( n7206 & n7211 ) | ( ~n7208 & n7211 ) ;
  assign n7213 = n7208 & n7212 ;
  assign n7214 = n7201 & ~n7204 ;
  assign n7215 = ~n7201 & n7204 ;
  assign n7216 = n7214 | n7215 ;
  assign n7217 = n7193 & ~n7196 ;
  assign n7218 = ~n7193 & n7196 ;
  assign n7219 = n7217 | n7218 ;
  assign n7220 = ~n7197 & n7219 ;
  assign n7221 = n7216 & n7220 ;
  assign n7222 = ~n7213 & n7221 ;
  assign n7223 = ( n7210 & n7212 ) | ( n7210 & n7222 ) | ( n7212 & n7222 ) ;
  assign n7224 = ( n7198 & n7208 ) | ( n7198 & n7223 ) | ( n7208 & n7223 ) ;
  assign n7225 = ( x823 & ~x824 ) | ( x823 & x825 ) | ( ~x824 & x825 ) ;
  assign n7226 = ( ~x823 & x824 ) | ( ~x823 & n7225 ) | ( x824 & n7225 ) ;
  assign n7227 = ( ~x825 & n7225 ) | ( ~x825 & n7226 ) | ( n7225 & n7226 ) ;
  assign n7228 = ( x826 & ~x827 ) | ( x826 & x828 ) | ( ~x827 & x828 ) ;
  assign n7229 = ( ~x826 & x827 ) | ( ~x826 & n7228 ) | ( x827 & n7228 ) ;
  assign n7230 = ( ~x828 & n7228 ) | ( ~x828 & n7229 ) | ( n7228 & n7229 ) ;
  assign n7231 = n7227 & n7230 ;
  assign n7232 = ( x826 & x827 ) | ( x826 & x828 ) | ( x827 & x828 ) ;
  assign n7233 = ( x823 & x824 ) | ( x823 & x825 ) | ( x824 & x825 ) ;
  assign n7234 = ( n7231 & n7232 ) | ( n7231 & n7233 ) | ( n7232 & n7233 ) ;
  assign n7235 = ( x832 & x833 ) | ( x832 & x834 ) | ( x833 & x834 ) ;
  assign n7236 = ( x829 & x830 ) | ( x829 & x831 ) | ( x830 & x831 ) ;
  assign n7237 = ( x829 & ~x830 ) | ( x829 & x831 ) | ( ~x830 & x831 ) ;
  assign n7238 = ( ~x829 & x830 ) | ( ~x829 & n7237 ) | ( x830 & n7237 ) ;
  assign n7239 = ( ~x831 & n7237 ) | ( ~x831 & n7238 ) | ( n7237 & n7238 ) ;
  assign n7240 = ( x832 & ~x833 ) | ( x832 & x834 ) | ( ~x833 & x834 ) ;
  assign n7241 = ( ~x832 & x833 ) | ( ~x832 & n7240 ) | ( x833 & n7240 ) ;
  assign n7242 = ( ~x834 & n7240 ) | ( ~x834 & n7241 ) | ( n7240 & n7241 ) ;
  assign n7243 = n7239 & n7242 ;
  assign n7244 = ( n7235 & n7236 ) | ( n7235 & n7243 ) | ( n7236 & n7243 ) ;
  assign n7245 = ( n7231 & n7233 ) | ( n7231 & ~n7234 ) | ( n7233 & ~n7234 ) ;
  assign n7246 = ( n7232 & ~n7234 ) | ( n7232 & n7245 ) | ( ~n7234 & n7245 ) ;
  assign n7247 = ( n7236 & n7243 ) | ( n7236 & ~n7244 ) | ( n7243 & ~n7244 ) ;
  assign n7248 = ( n7235 & ~n7244 ) | ( n7235 & n7247 ) | ( ~n7244 & n7247 ) ;
  assign n7249 = n7234 & n7246 ;
  assign n7250 = n7244 & n7248 ;
  assign n7251 = n7227 & ~n7230 ;
  assign n7252 = ~n7227 & n7230 ;
  assign n7253 = n7251 | n7252 ;
  assign n7254 = n7239 & ~n7242 ;
  assign n7255 = ~n7239 & n7242 ;
  assign n7256 = n7254 | n7255 ;
  assign n7257 = n7253 & n7256 ;
  assign n7258 = ~n7250 & n7257 ;
  assign n7259 = ~n7249 & n7258 ;
  assign n7260 = ~n7248 & n7259 ;
  assign n7261 = ( n7246 & n7248 ) | ( n7246 & n7260 ) | ( n7248 & n7260 ) ;
  assign n7262 = n7248 & n7258 ;
  assign n7263 = ~n7249 & n7262 ;
  assign n7264 = n7261 | n7263 ;
  assign n7265 = ( n7234 & n7244 ) | ( n7234 & n7264 ) | ( n7244 & n7264 ) ;
  assign n7266 = ~n7234 & n7244 ;
  assign n7267 = n7234 & ~n7244 ;
  assign n7268 = n7266 | n7267 ;
  assign n7269 = n7263 | n7268 ;
  assign n7270 = n7261 | n7269 ;
  assign n7271 = n7264 & n7268 ;
  assign n7272 = n7270 & ~n7271 ;
  assign n7273 = ( n7198 & n7208 ) | ( n7198 & ~n7223 ) | ( n7208 & ~n7223 ) ;
  assign n7274 = ( n7198 & ~n7208 ) | ( n7198 & n7223 ) | ( ~n7208 & n7223 ) ;
  assign n7275 = ( ~n7198 & n7273 ) | ( ~n7198 & n7274 ) | ( n7273 & n7274 ) ;
  assign n7276 = n7272 | n7275 ;
  assign n7277 = ( n7246 & n7248 ) | ( n7246 & ~n7259 ) | ( n7248 & ~n7259 ) ;
  assign n7278 = n7246 & ~n7263 ;
  assign n7279 = ( n7248 & ~n7277 ) | ( n7248 & n7278 ) | ( ~n7277 & n7278 ) ;
  assign n7280 = ( n7260 & n7277 ) | ( n7260 & ~n7279 ) | ( n7277 & ~n7279 ) ;
  assign n7281 = n7216 & ~n7220 ;
  assign n7282 = ~n7216 & n7220 ;
  assign n7283 = n7281 | n7282 ;
  assign n7284 = n7253 & ~n7256 ;
  assign n7285 = ~n7253 & n7256 ;
  assign n7286 = n7284 | n7285 ;
  assign n7287 = n7283 & n7286 ;
  assign n7288 = n7210 | n7222 ;
  assign n7289 = ~n7223 & n7288 ;
  assign n7290 = n7210 & n7221 ;
  assign n7291 = ( n7212 & ~n7288 ) | ( n7212 & n7290 ) | ( ~n7288 & n7290 ) ;
  assign n7292 = n7289 | n7291 ;
  assign n7293 = n7287 | n7292 ;
  assign n7294 = ( n7287 & n7289 ) | ( n7287 & n7291 ) | ( n7289 & n7291 ) ;
  assign n7295 = ( n7280 & n7293 ) | ( n7280 & n7294 ) | ( n7293 & n7294 ) ;
  assign n7296 = n7276 & n7295 ;
  assign n7297 = n7272 & n7275 ;
  assign n7298 = n7296 | n7297 ;
  assign n7299 = ( n7224 & n7265 ) | ( n7224 & n7298 ) | ( n7265 & n7298 ) ;
  assign n7300 = n7188 & n7299 ;
  assign n7301 = ~n7224 & n7265 ;
  assign n7302 = n7224 & ~n7265 ;
  assign n7303 = n7301 | n7302 ;
  assign n7304 = n7297 | n7303 ;
  assign n7305 = n7296 | n7304 ;
  assign n7306 = n7298 & n7303 ;
  assign n7307 = n7305 & ~n7306 ;
  assign n7308 = ~n7115 & n7156 ;
  assign n7309 = n7115 & ~n7156 ;
  assign n7310 = n7308 | n7309 ;
  assign n7311 = n7187 | n7310 ;
  assign n7312 = ~n7310 & n7311 ;
  assign n7313 = ( ~n7187 & n7311 ) | ( ~n7187 & n7312 ) | ( n7311 & n7312 ) ;
  assign n7314 = n7307 | n7313 ;
  assign n7315 = ( n7176 & ~n7183 ) | ( n7176 & n7186 ) | ( ~n7183 & n7186 ) ;
  assign n7316 = ( ~n7176 & n7183 ) | ( ~n7176 & n7315 ) | ( n7183 & n7315 ) ;
  assign n7317 = ( ~n7186 & n7315 ) | ( ~n7186 & n7316 ) | ( n7315 & n7316 ) ;
  assign n7318 = ( ~n7272 & n7275 ) | ( ~n7272 & n7295 ) | ( n7275 & n7295 ) ;
  assign n7319 = ( n7272 & ~n7295 ) | ( n7272 & n7318 ) | ( ~n7295 & n7318 ) ;
  assign n7320 = ( ~n7275 & n7318 ) | ( ~n7275 & n7319 ) | ( n7318 & n7319 ) ;
  assign n7321 = n7283 & ~n7286 ;
  assign n7322 = ~n7283 & n7286 ;
  assign n7323 = n7321 | n7322 ;
  assign n7324 = n7163 & ~n7166 ;
  assign n7325 = ~n7163 & n7166 ;
  assign n7326 = n7324 | n7325 ;
  assign n7327 = n7323 & n7326 ;
  assign n7328 = ~n7287 & n7293 ;
  assign n7329 = ( ~n7292 & n7293 ) | ( ~n7292 & n7328 ) | ( n7293 & n7328 ) ;
  assign n7330 = n7280 & ~n7329 ;
  assign n7331 = ~n7280 & n7329 ;
  assign n7332 = n7330 | n7331 ;
  assign n7333 = ( n7160 & n7167 ) | ( n7160 & ~n7172 ) | ( n7167 & ~n7172 ) ;
  assign n7334 = ( ~n7160 & n7172 ) | ( ~n7160 & n7333 ) | ( n7172 & n7333 ) ;
  assign n7335 = ( ~n7167 & n7333 ) | ( ~n7167 & n7334 ) | ( n7333 & n7334 ) ;
  assign n7336 = ( n7327 & n7332 ) | ( n7327 & n7335 ) | ( n7332 & n7335 ) ;
  assign n7337 = ( n7317 & n7320 ) | ( n7317 & n7336 ) | ( n7320 & n7336 ) ;
  assign n7338 = n7314 & n7337 ;
  assign n7339 = n7307 & n7313 ;
  assign n7340 = n7338 | n7339 ;
  assign n7341 = n7299 & ~n7300 ;
  assign n7342 = ( n7188 & ~n7300 ) | ( n7188 & n7341 ) | ( ~n7300 & n7341 ) ;
  assign n7343 = n7340 & n7342 ;
  assign n7344 = ( n7299 & n7340 ) | ( n7299 & n7343 ) | ( n7340 & n7343 ) ;
  assign n7345 = n7300 | n7344 ;
  assign n7346 = n7080 & n7345 ;
  assign n7347 = n7076 | n7300 ;
  assign n7348 = n7079 | n7347 ;
  assign n7349 = ( n7072 & n7347 ) | ( n7072 & n7348 ) | ( n7347 & n7348 ) ;
  assign n7350 = n7344 | n7349 ;
  assign n7351 = n7071 | n7078 ;
  assign n7352 = n7070 | n7351 ;
  assign n7353 = n7072 & n7078 ;
  assign n7354 = n7352 & ~n7353 ;
  assign n7355 = n7339 | n7342 ;
  assign n7356 = n7338 | n7355 ;
  assign n7357 = ~n7343 & n7356 ;
  assign n7358 = n7354 | n7357 ;
  assign n7359 = ( ~n7049 & n7052 ) | ( ~n7049 & n7068 ) | ( n7052 & n7068 ) ;
  assign n7360 = ( n7049 & ~n7068 ) | ( n7049 & n7359 ) | ( ~n7068 & n7359 ) ;
  assign n7361 = ( ~n7052 & n7359 ) | ( ~n7052 & n7360 ) | ( n7359 & n7360 ) ;
  assign n7362 = ( ~n7317 & n7320 ) | ( ~n7317 & n7336 ) | ( n7320 & n7336 ) ;
  assign n7363 = ( n7317 & ~n7336 ) | ( n7317 & n7362 ) | ( ~n7336 & n7362 ) ;
  assign n7364 = ( ~n7320 & n7362 ) | ( ~n7320 & n7363 ) | ( n7362 & n7363 ) ;
  assign n7365 = n7323 & ~n7326 ;
  assign n7366 = ~n7323 & n7326 ;
  assign n7367 = n7365 | n7366 ;
  assign n7368 = n7055 & ~n7058 ;
  assign n7369 = ~n7055 & n7058 ;
  assign n7370 = n7368 | n7369 ;
  assign n7371 = n7367 & n7370 ;
  assign n7372 = ( n7327 & ~n7332 ) | ( n7327 & n7335 ) | ( ~n7332 & n7335 ) ;
  assign n7373 = ( ~n7327 & n7332 ) | ( ~n7327 & n7372 ) | ( n7332 & n7372 ) ;
  assign n7374 = ( ~n7335 & n7372 ) | ( ~n7335 & n7373 ) | ( n7372 & n7373 ) ;
  assign n7375 = ( n7059 & ~n7064 ) | ( n7059 & n7067 ) | ( ~n7064 & n7067 ) ;
  assign n7376 = ( ~n7059 & n7064 ) | ( ~n7059 & n7375 ) | ( n7064 & n7375 ) ;
  assign n7377 = ( ~n7067 & n7375 ) | ( ~n7067 & n7376 ) | ( n7375 & n7376 ) ;
  assign n7378 = ( n7371 & n7374 ) | ( n7371 & n7377 ) | ( n7374 & n7377 ) ;
  assign n7379 = ( n7361 & n7364 ) | ( n7361 & n7378 ) | ( n7364 & n7378 ) ;
  assign n7380 = ( ~n7307 & n7313 ) | ( ~n7307 & n7337 ) | ( n7313 & n7337 ) ;
  assign n7381 = ( n7307 & ~n7337 ) | ( n7307 & n7380 ) | ( ~n7337 & n7380 ) ;
  assign n7382 = ( ~n7313 & n7380 ) | ( ~n7313 & n7381 ) | ( n7380 & n7381 ) ;
  assign n7383 = ( ~n6929 & n7045 ) | ( ~n6929 & n7069 ) | ( n7045 & n7069 ) ;
  assign n7384 = ( n6929 & ~n7069 ) | ( n6929 & n7383 ) | ( ~n7069 & n7383 ) ;
  assign n7385 = ( ~n7045 & n7383 ) | ( ~n7045 & n7384 ) | ( n7383 & n7384 ) ;
  assign n7386 = ( n7379 & n7382 ) | ( n7379 & n7385 ) | ( n7382 & n7385 ) ;
  assign n7387 = n7358 & n7386 ;
  assign n7388 = n7354 & n7357 ;
  assign n7389 = n7387 | n7388 ;
  assign n7390 = n7350 & n7389 ;
  assign n7391 = n7346 | n7390 ;
  assign n7392 = n6812 & n7391 ;
  assign n7393 = n6771 | n7346 ;
  assign n7394 = n6775 | n7393 ;
  assign n7395 = ( n6811 & n7393 ) | ( n6811 & n7394 ) | ( n7393 & n7394 ) ;
  assign n7396 = n7390 | n7395 ;
  assign n7397 = n7345 & ~n7346 ;
  assign n7398 = ( n7080 & ~n7346 ) | ( n7080 & n7397 ) | ( ~n7346 & n7397 ) ;
  assign n7399 = n7388 | n7398 ;
  assign n7400 = n7387 | n7399 ;
  assign n7401 = n7389 & n7398 ;
  assign n7402 = n7400 & ~n7401 ;
  assign n7403 = ( n6505 & n6770 ) | ( n6505 & ~n6811 ) | ( n6770 & ~n6811 ) ;
  assign n7404 = ( ~n6770 & n6811 ) | ( ~n6770 & n7403 ) | ( n6811 & n7403 ) ;
  assign n7405 = ( ~n6505 & n7403 ) | ( ~n6505 & n7404 ) | ( n7403 & n7404 ) ;
  assign n7406 = ( ~n6779 & n6782 ) | ( ~n6779 & n6810 ) | ( n6782 & n6810 ) ;
  assign n7407 = ( n6779 & ~n6810 ) | ( n6779 & n7406 ) | ( ~n6810 & n7406 ) ;
  assign n7408 = ( ~n6782 & n7406 ) | ( ~n6782 & n7407 ) | ( n7406 & n7407 ) ;
  assign n7409 = ( ~n7354 & n7357 ) | ( ~n7354 & n7386 ) | ( n7357 & n7386 ) ;
  assign n7410 = ( n7354 & ~n7386 ) | ( n7354 & n7409 ) | ( ~n7386 & n7409 ) ;
  assign n7411 = ( ~n7357 & n7409 ) | ( ~n7357 & n7410 ) | ( n7409 & n7410 ) ;
  assign n7412 = ( ~n6785 & n6788 ) | ( ~n6785 & n6802 ) | ( n6788 & n6802 ) ;
  assign n7413 = ( n6785 & ~n6802 ) | ( n6785 & n7412 ) | ( ~n6802 & n7412 ) ;
  assign n7414 = ( ~n6788 & n7412 ) | ( ~n6788 & n7413 ) | ( n7412 & n7413 ) ;
  assign n7415 = ( ~n7361 & n7364 ) | ( ~n7361 & n7378 ) | ( n7364 & n7378 ) ;
  assign n7416 = ( n7361 & ~n7378 ) | ( n7361 & n7415 ) | ( ~n7378 & n7415 ) ;
  assign n7417 = ( ~n7364 & n7415 ) | ( ~n7364 & n7416 ) | ( n7415 & n7416 ) ;
  assign n7418 = n7367 & ~n7370 ;
  assign n7419 = ~n7367 & n7370 ;
  assign n7420 = n7418 | n7419 ;
  assign n7421 = n6791 & ~n6794 ;
  assign n7422 = ~n6791 & n6794 ;
  assign n7423 = n7421 | n7422 ;
  assign n7424 = n7420 & n7423 ;
  assign n7425 = ~n7371 & n7374 ;
  assign n7426 = n7371 & ~n7374 ;
  assign n7427 = n7425 | n7426 ;
  assign n7428 = n7377 & ~n7427 ;
  assign n7429 = ~n7377 & n7427 ;
  assign n7430 = n7428 | n7429 ;
  assign n7431 = ( n6795 & n6801 ) | ( n6795 & ~n6802 ) | ( n6801 & ~n6802 ) ;
  assign n7432 = ( n6798 & ~n6802 ) | ( n6798 & n7431 ) | ( ~n6802 & n7431 ) ;
  assign n7433 = ( n7424 & n7430 ) | ( n7424 & n7432 ) | ( n7430 & n7432 ) ;
  assign n7434 = ( n7414 & n7417 ) | ( n7414 & n7433 ) | ( n7417 & n7433 ) ;
  assign n7435 = ( n7379 & ~n7382 ) | ( n7379 & n7385 ) | ( ~n7382 & n7385 ) ;
  assign n7436 = ( ~n7379 & n7382 ) | ( ~n7379 & n7435 ) | ( n7382 & n7435 ) ;
  assign n7437 = ( ~n7385 & n7435 ) | ( ~n7385 & n7436 ) | ( n7435 & n7436 ) ;
  assign n7438 = ( n6803 & ~n6806 ) | ( n6803 & n6809 ) | ( ~n6806 & n6809 ) ;
  assign n7439 = ( ~n6803 & n6806 ) | ( ~n6803 & n7438 ) | ( n6806 & n7438 ) ;
  assign n7440 = ( ~n6809 & n7438 ) | ( ~n6809 & n7439 ) | ( n7438 & n7439 ) ;
  assign n7441 = ( n7434 & n7437 ) | ( n7434 & n7440 ) | ( n7437 & n7440 ) ;
  assign n7442 = ( n7408 & n7411 ) | ( n7408 & n7441 ) | ( n7411 & n7441 ) ;
  assign n7443 = ( n7402 & n7405 ) | ( n7402 & n7442 ) | ( n7405 & n7442 ) ;
  assign n7444 = n7396 & n7443 ;
  assign n7445 = n7392 | n7444 ;
  assign n7446 = n6179 & ~n6180 ;
  assign n7447 = ( n5593 & ~n6180 ) | ( n5593 & n7446 ) | ( ~n6180 & n7446 ) ;
  assign n7448 = n6233 | n7447 ;
  assign n7449 = n6232 | n7448 ;
  assign n7450 = n6234 & n7447 ;
  assign n7451 = n7449 & ~n7450 ;
  assign n7452 = ( n6812 & n7391 ) | ( n6812 & ~n7443 ) | ( n7391 & ~n7443 ) ;
  assign n7453 = ( ~n7391 & n7443 ) | ( ~n7391 & n7452 ) | ( n7443 & n7452 ) ;
  assign n7454 = ( ~n6812 & n7452 ) | ( ~n6812 & n7453 ) | ( n7452 & n7453 ) ;
  assign n7455 = ( ~n7402 & n7405 ) | ( ~n7402 & n7442 ) | ( n7405 & n7442 ) ;
  assign n7456 = ( n7402 & ~n7442 ) | ( n7402 & n7455 ) | ( ~n7442 & n7455 ) ;
  assign n7457 = ( ~n7405 & n7455 ) | ( ~n7405 & n7456 ) | ( n7455 & n7456 ) ;
  assign n7458 = ( ~n6190 & n6193 ) | ( ~n6190 & n6231 ) | ( n6193 & n6231 ) ;
  assign n7459 = ( n6190 & ~n6231 ) | ( n6190 & n7458 ) | ( ~n6231 & n7458 ) ;
  assign n7460 = ( ~n6193 & n7458 ) | ( ~n6193 & n7459 ) | ( n7458 & n7459 ) ;
  assign n7461 = ( n6197 & ~n6200 ) | ( n6197 & n6230 ) | ( ~n6200 & n6230 ) ;
  assign n7462 = ( ~n6197 & n6200 ) | ( ~n6197 & n7461 ) | ( n6200 & n7461 ) ;
  assign n7463 = ( ~n6230 & n7461 ) | ( ~n6230 & n7462 ) | ( n7461 & n7462 ) ;
  assign n7464 = ( n7408 & ~n7411 ) | ( n7408 & n7441 ) | ( ~n7411 & n7441 ) ;
  assign n7465 = ( ~n7408 & n7411 ) | ( ~n7408 & n7464 ) | ( n7411 & n7464 ) ;
  assign n7466 = ( ~n7441 & n7464 ) | ( ~n7441 & n7465 ) | ( n7464 & n7465 ) ;
  assign n7467 = ( ~n6203 & n6206 ) | ( ~n6203 & n6222 ) | ( n6206 & n6222 ) ;
  assign n7468 = ( n6203 & ~n6222 ) | ( n6203 & n7467 ) | ( ~n6222 & n7467 ) ;
  assign n7469 = ( ~n6206 & n7467 ) | ( ~n6206 & n7468 ) | ( n7467 & n7468 ) ;
  assign n7470 = ( ~n7414 & n7417 ) | ( ~n7414 & n7433 ) | ( n7417 & n7433 ) ;
  assign n7471 = ( n7414 & ~n7433 ) | ( n7414 & n7470 ) | ( ~n7433 & n7470 ) ;
  assign n7472 = ( ~n7417 & n7470 ) | ( ~n7417 & n7471 ) | ( n7470 & n7471 ) ;
  assign n7473 = n6209 & ~n6212 ;
  assign n7474 = ~n6209 & n6212 ;
  assign n7475 = n7473 | n7474 ;
  assign n7476 = n7420 & ~n7423 ;
  assign n7477 = ~n7420 & n7423 ;
  assign n7478 = n7476 | n7477 ;
  assign n7479 = n7475 & n7478 ;
  assign n7480 = ( n7424 & ~n7430 ) | ( n7424 & n7432 ) | ( ~n7430 & n7432 ) ;
  assign n7481 = ( ~n7424 & n7430 ) | ( ~n7424 & n7480 ) | ( n7430 & n7480 ) ;
  assign n7482 = ( ~n7432 & n7480 ) | ( ~n7432 & n7481 ) | ( n7480 & n7481 ) ;
  assign n7483 = ( n6213 & ~n6219 ) | ( n6213 & n6221 ) | ( ~n6219 & n6221 ) ;
  assign n7484 = ( ~n6213 & n6219 ) | ( ~n6213 & n7483 ) | ( n6219 & n7483 ) ;
  assign n7485 = ( ~n6221 & n7483 ) | ( ~n6221 & n7484 ) | ( n7483 & n7484 ) ;
  assign n7486 = ( n7479 & n7482 ) | ( n7479 & n7485 ) | ( n7482 & n7485 ) ;
  assign n7487 = ( n7469 & n7472 ) | ( n7469 & n7486 ) | ( n7472 & n7486 ) ;
  assign n7488 = ( n7434 & ~n7437 ) | ( n7434 & n7440 ) | ( ~n7437 & n7440 ) ;
  assign n7489 = ( ~n7434 & n7437 ) | ( ~n7434 & n7488 ) | ( n7437 & n7488 ) ;
  assign n7490 = ( ~n7440 & n7488 ) | ( ~n7440 & n7489 ) | ( n7488 & n7489 ) ;
  assign n7491 = ( n6223 & ~n6226 ) | ( n6223 & n6229 ) | ( ~n6226 & n6229 ) ;
  assign n7492 = ( ~n6223 & n6226 ) | ( ~n6223 & n7491 ) | ( n6226 & n7491 ) ;
  assign n7493 = ( ~n6229 & n7491 ) | ( ~n6229 & n7492 ) | ( n7491 & n7492 ) ;
  assign n7494 = ( n7487 & n7490 ) | ( n7487 & n7493 ) | ( n7490 & n7493 ) ;
  assign n7495 = ( n7463 & n7466 ) | ( n7463 & n7494 ) | ( n7466 & n7494 ) ;
  assign n7496 = ( n7457 & n7460 ) | ( n7457 & n7495 ) | ( n7460 & n7495 ) ;
  assign n7497 = ( n7451 & n7454 ) | ( n7451 & n7496 ) | ( n7454 & n7496 ) ;
  assign n7498 = ( n6235 & n7445 ) | ( n6235 & ~n7497 ) | ( n7445 & ~n7497 ) ;
  assign n7499 = ( ~n7445 & n7497 ) | ( ~n7445 & n7498 ) | ( n7497 & n7498 ) ;
  assign n7500 = ( ~n6235 & n7498 ) | ( ~n6235 & n7499 ) | ( n7498 & n7499 ) ;
  assign n7501 = n5003 & n5008 ;
  assign n7502 = ~n5006 & n7501 ;
  assign n7503 = n5003 | n5009 ;
  assign n7504 = ~n7502 & n7503 ;
  assign n7505 = n4999 | n7504 ;
  assign n7506 = n4999 & n7504 ;
  assign n7507 = n7505 & ~n7506 ;
  assign n7508 = ( ~n7451 & n7454 ) | ( ~n7451 & n7496 ) | ( n7454 & n7496 ) ;
  assign n7509 = ( n7451 & ~n7496 ) | ( n7451 & n7508 ) | ( ~n7496 & n7508 ) ;
  assign n7510 = ( ~n7454 & n7508 ) | ( ~n7454 & n7509 ) | ( n7508 & n7509 ) ;
  assign n7511 = ~n4955 & n4958 ;
  assign n7512 = n4955 & ~n4958 ;
  assign n7513 = n7511 | n7512 ;
  assign n7514 = n4998 | n7513 ;
  assign n7515 = n4998 & n7513 ;
  assign n7516 = n7514 & ~n7515 ;
  assign n7517 = ( n7457 & ~n7460 ) | ( n7457 & n7495 ) | ( ~n7460 & n7495 ) ;
  assign n7518 = ( ~n7457 & n7460 ) | ( ~n7457 & n7517 ) | ( n7460 & n7517 ) ;
  assign n7519 = ( ~n7495 & n7517 ) | ( ~n7495 & n7518 ) | ( n7517 & n7518 ) ;
  assign n7520 = ( ~n4961 & n4994 ) | ( ~n4961 & n4997 ) | ( n4994 & n4997 ) ;
  assign n7521 = ( n4961 & ~n4997 ) | ( n4961 & n7520 ) | ( ~n4997 & n7520 ) ;
  assign n7522 = ( ~n4994 & n7520 ) | ( ~n4994 & n7521 ) | ( n7520 & n7521 ) ;
  assign n7523 = ( n7463 & ~n7466 ) | ( n7463 & n7494 ) | ( ~n7466 & n7494 ) ;
  assign n7524 = ( ~n7463 & n7466 ) | ( ~n7463 & n7523 ) | ( n7466 & n7523 ) ;
  assign n7525 = ( ~n7494 & n7523 ) | ( ~n7494 & n7524 ) | ( n7523 & n7524 ) ;
  assign n7526 = n4991 & ~n4993 ;
  assign n7527 = ~n4991 & n4993 ;
  assign n7528 = n7526 | n7527 ;
  assign n7529 = n4988 | n7528 ;
  assign n7530 = n4988 & n7528 ;
  assign n7531 = n7529 & ~n7530 ;
  assign n7532 = ( n7487 & ~n7490 ) | ( n7487 & n7493 ) | ( ~n7490 & n7493 ) ;
  assign n7533 = ( ~n7487 & n7490 ) | ( ~n7487 & n7532 ) | ( n7490 & n7532 ) ;
  assign n7534 = ( ~n7493 & n7532 ) | ( ~n7493 & n7533 ) | ( n7532 & n7533 ) ;
  assign n7535 = n4964 & ~n4983 ;
  assign n7536 = ~n4964 & n4983 ;
  assign n7537 = n7535 | n7536 ;
  assign n7538 = n4980 | n7537 ;
  assign n7539 = ( ~n7469 & n7472 ) | ( ~n7469 & n7486 ) | ( n7472 & n7486 ) ;
  assign n7540 = ( n7469 & ~n7486 ) | ( n7469 & n7539 ) | ( ~n7486 & n7539 ) ;
  assign n7541 = ( ~n7472 & n7539 ) | ( ~n7472 & n7540 ) | ( n7539 & n7540 ) ;
  assign n7542 = ( n4980 & n7537 ) | ( n4980 & ~n7541 ) | ( n7537 & ~n7541 ) ;
  assign n7543 = n7475 & ~n7478 ;
  assign n7544 = ~n7475 & n7478 ;
  assign n7545 = n7543 | n7544 ;
  assign n7546 = n4967 & ~n4971 ;
  assign n7547 = ( n4970 & ~n4971 ) | ( n4970 & n7546 ) | ( ~n4971 & n7546 ) ;
  assign n7548 = n7545 & n7547 ;
  assign n7549 = n4971 & n4977 ;
  assign n7550 = ( n4979 & ~n4980 ) | ( n4979 & n7549 ) | ( ~n4980 & n7549 ) ;
  assign n7551 = ( n4971 & n4977 ) | ( n4971 & ~n4979 ) | ( n4977 & ~n4979 ) ;
  assign n7552 = ~n7549 & n7551 ;
  assign n7553 = n7550 | n7552 ;
  assign n7554 = ( n7479 & n7485 ) | ( n7479 & ~n7486 ) | ( n7485 & ~n7486 ) ;
  assign n7555 = ( n7482 & ~n7486 ) | ( n7482 & n7554 ) | ( ~n7486 & n7554 ) ;
  assign n7556 = ( n7548 & n7553 ) | ( n7548 & n7555 ) | ( n7553 & n7555 ) ;
  assign n7557 = n4980 & n7537 ;
  assign n7558 = ( ~n7538 & n7541 ) | ( ~n7538 & n7557 ) | ( n7541 & n7557 ) ;
  assign n7559 = n7542 & ~n7557 ;
  assign n7560 = ( n7556 & n7558 ) | ( n7556 & n7559 ) | ( n7558 & n7559 ) ;
  assign n7561 = ( n7538 & ~n7542 ) | ( n7538 & n7560 ) | ( ~n7542 & n7560 ) ;
  assign n7562 = n4936 & n4987 ;
  assign n7563 = n4987 & ~n7562 ;
  assign n7564 = ( n4936 & ~n7562 ) | ( n4936 & n7563 ) | ( ~n7562 & n7563 ) ;
  assign n7565 = ( n4984 & n7534 ) | ( n4984 & ~n7564 ) | ( n7534 & ~n7564 ) ;
  assign n7566 = ( ~n4984 & n7564 ) | ( ~n4984 & n7565 ) | ( n7564 & n7565 ) ;
  assign n7567 = ( ~n7534 & n7565 ) | ( ~n7534 & n7566 ) | ( n7565 & n7566 ) ;
  assign n7568 = n7561 & n7567 ;
  assign n7569 = n7561 | n7567 ;
  assign n7570 = ~n7568 & n7569 ;
  assign n7571 = ( n7534 & n7561 ) | ( n7534 & ~n7570 ) | ( n7561 & ~n7570 ) ;
  assign n7572 = ( n7534 & n7561 ) | ( n7534 & n7571 ) | ( n7561 & n7571 ) ;
  assign n7573 = ( n7525 & n7531 ) | ( n7525 & n7572 ) | ( n7531 & n7572 ) ;
  assign n7574 = ( n7519 & n7522 ) | ( n7519 & n7573 ) | ( n7522 & n7573 ) ;
  assign n7575 = ( n7510 & n7516 ) | ( n7510 & n7574 ) | ( n7516 & n7574 ) ;
  assign n7576 = ( n7500 & n7507 ) | ( n7500 & n7575 ) | ( n7507 & n7575 ) ;
  assign n7577 = n6235 & n7445 ;
  assign n7578 = n6180 | n7392 ;
  assign n7579 = n6184 | n7578 ;
  assign n7580 = ( n6234 & n7578 ) | ( n6234 & n7579 ) | ( n7578 & n7579 ) ;
  assign n7581 = n7444 | n7580 ;
  assign n7582 = n7577 | n7581 ;
  assign n7583 = ( n7497 & n7577 ) | ( n7497 & n7582 ) | ( n7577 & n7582 ) ;
  assign n7584 = n4951 & ~n4953 ;
  assign n7585 = n5010 & n7584 ;
  assign n7586 = ( n4951 & ~n4953 ) | ( n4951 & n5010 ) | ( ~n4953 & n5010 ) ;
  assign n7587 = ~n7585 & n7586 ;
  assign n7588 = n7583 & ~n7587 ;
  assign n7589 = ( ~n7583 & n7587 ) | ( ~n7583 & n7588 ) | ( n7587 & n7588 ) ;
  assign n7590 = n7588 | n7589 ;
  assign n7591 = n7576 & n7590 ;
  assign n7592 = n7500 & ~n7506 ;
  assign n7593 = n7505 & n7592 ;
  assign n7594 = n7590 | n7593 ;
  assign n7595 = n7576 | n7594 ;
  assign n7596 = ~n7591 & n7595 ;
  assign n7597 = n7583 & n7587 ;
  assign n7598 = ( n7576 & ~n7596 ) | ( n7576 & n7597 ) | ( ~n7596 & n7597 ) ;
  assign n7599 = n5011 & n7598 ;
  assign n7600 = ( x1000 & n7545 ) | ( x1000 & ~n7547 ) | ( n7545 & ~n7547 ) ;
  assign n7601 = ( ~n7545 & n7547 ) | ( ~n7545 & n7600 ) | ( n7547 & n7600 ) ;
  assign n7602 = ( ~x1000 & n7600 ) | ( ~x1000 & n7601 ) | ( n7600 & n7601 ) ;
  assign n7603 = x1000 & ~n7602 ;
  assign n7604 = ~n7560 & n7603 ;
  assign n7605 = n7548 & n7553 ;
  assign n7606 = n7548 | n7553 ;
  assign n7607 = ~n7605 & n7606 ;
  assign n7608 = ~n7555 & n7607 ;
  assign n7609 = n7555 & ~n7607 ;
  assign n7610 = n7556 | n7559 ;
  assign n7611 = n7558 | n7610 ;
  assign n7612 = ( n7608 & n7609 ) | ( n7608 & n7611 ) | ( n7609 & n7611 ) ;
  assign n7613 = n7604 & n7612 ;
  assign n7614 = ~n7568 & n7613 ;
  assign n7615 = n7569 & n7614 ;
  assign n7616 = ( n7525 & n7531 ) | ( n7525 & ~n7572 ) | ( n7531 & ~n7572 ) ;
  assign n7617 = ( ~n7531 & n7572 ) | ( ~n7531 & n7616 ) | ( n7572 & n7616 ) ;
  assign n7618 = ( ~n7525 & n7616 ) | ( ~n7525 & n7617 ) | ( n7616 & n7617 ) ;
  assign n7619 = n7615 & n7618 ;
  assign n7620 = ( n7522 & n7573 ) | ( n7522 & ~n7574 ) | ( n7573 & ~n7574 ) ;
  assign n7621 = ( n7519 & ~n7574 ) | ( n7519 & n7620 ) | ( ~n7574 & n7620 ) ;
  assign n7622 = n7619 & n7621 ;
  assign n7623 = ( n7516 & n7574 ) | ( n7516 & ~n7575 ) | ( n7574 & ~n7575 ) ;
  assign n7624 = ( n7510 & ~n7575 ) | ( n7510 & n7623 ) | ( ~n7575 & n7623 ) ;
  assign n7625 = n7622 & n7624 ;
  assign n7626 = ( n7507 & n7575 ) | ( n7507 & ~n7576 ) | ( n7575 & ~n7576 ) ;
  assign n7627 = ( n7500 & ~n7576 ) | ( n7500 & n7626 ) | ( ~n7576 & n7626 ) ;
  assign n7628 = n7625 & n7627 ;
  assign n7629 = n7596 & n7628 ;
  assign n7630 = ~n5011 & n7598 ;
  assign n7631 = ( n5011 & ~n7598 ) | ( n5011 & n7630 ) | ( ~n7598 & n7630 ) ;
  assign n7632 = ~n7597 & n7631 ;
  assign n7633 = n7630 | n7632 ;
  assign n7634 = n7629 & n7633 ;
  assign n7635 = n7629 | n7633 ;
  assign n7636 = n7615 | n7618 ;
  assign n7637 = ~n7619 & n7636 ;
  assign n7638 = n7570 | n7613 ;
  assign n7639 = ~n7615 & n7638 ;
  assign n7640 = ( n7603 & n7608 ) | ( n7603 & n7609 ) | ( n7608 & n7609 ) ;
  assign n7644 = ( n7603 & n7608 ) | ( n7603 & ~n7640 ) | ( n7608 & ~n7640 ) ;
  assign n7645 = ( n7609 & ~n7640 ) | ( n7609 & n7644 ) | ( ~n7640 & n7644 ) ;
  assign n7641 = ( ~n7560 & n7611 ) | ( ~n7560 & n7640 ) | ( n7611 & n7640 ) ;
  assign n7642 = ~n7613 & n7641 ;
  assign n7648 = ( n7615 & n7639 ) | ( n7615 & n7642 ) | ( n7639 & n7642 ) ;
  assign n7649 = ( n7639 & n7645 ) | ( n7639 & n7648 ) | ( n7645 & n7648 ) ;
  assign n7643 = ~n7639 & n7642 ;
  assign n7646 = ( n7602 & n7643 ) | ( n7602 & n7645 ) | ( n7643 & n7645 ) ;
  assign n7647 = n7643 & n7646 ;
  assign n7650 = ( n7639 & n7647 ) | ( n7639 & ~n7649 ) | ( n7647 & ~n7649 ) ;
  assign n7651 = ( n7637 & n7649 ) | ( n7637 & n7650 ) | ( n7649 & n7650 ) ;
  assign n7652 = n7625 | n7627 ;
  assign n7653 = ~n7628 & n7652 ;
  assign n7654 = n7619 | n7621 ;
  assign n7655 = ~n7622 & n7654 ;
  assign n7656 = n7637 | n7649 ;
  assign n7657 = n7655 & n7656 ;
  assign n7658 = n7622 | n7624 ;
  assign n7659 = ~n7625 & n7658 ;
  assign n7660 = n7657 & n7659 ;
  assign n7661 = n7653 & n7660 ;
  assign n7662 = n7596 & n7661 ;
  assign n7663 = n7651 & n7662 ;
  assign n7664 = ( ~n7629 & n7633 ) | ( ~n7629 & n7663 ) | ( n7633 & n7663 ) ;
  assign n7665 = ( ~n7633 & n7635 ) | ( ~n7633 & n7664 ) | ( n7635 & n7664 ) ;
  assign n7666 = ( ~n7599 & n7634 ) | ( ~n7599 & n7665 ) | ( n7634 & n7665 ) ;
  assign n7667 = n7599 | n7666 ;
  assign y0 = n7667 ;
endmodule
