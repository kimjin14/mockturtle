module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 ;
  wire n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , n3931 , n3932 , n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , n3940 , n3941 , n3942 , n3943 , n3944 , n3945 , n3946 , n3947 , n3948 , n3949 , n3950 , n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , n3970 , n3971 , n3972 , n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , n3980 , n3981 , n3982 , n3983 , n3984 , n3985 , n3986 , n3987 , n3988 , n3989 , n3990 , n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , n4000 , n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , n4009 , n4010 , n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , n4019 , n4020 , n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , n4029 , n4030 , n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , n4039 , n4040 , n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4049 , n4050 , n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , n4059 , n4060 , n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , n4070 , n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , n4079 , n4080 , n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , n4089 , n4090 , n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , n4097 , n4098 , n4099 , n4100 , n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , n4109 , n4110 , n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , n4119 , n4120 , n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , n4129 , n4130 , n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , n4139 , n4140 , n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , n4150 , n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , n4159 , n4160 , n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , n4169 , n4170 , n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , n4179 , n4180 , n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , n4189 , n4190 , n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , n4197 , n4198 , n4199 , n4200 , n4201 , n4202 , n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , n4209 , n4210 , n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , n4217 , n4218 , n4219 , n4220 , n4221 , n4222 , n4223 , n4224 , n4225 , n4226 , n4227 , n4228 , n4229 , n4230 , n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , n4237 , n4238 , n4239 , n4240 , n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , n4247 , n4248 , n4249 , n4250 , n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , n4259 , n4260 , n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , n4269 , n4270 , n4271 , n4272 , n4273 , n4274 , n4275 , n4276 , n4277 , n4278 , n4279 , n4280 , n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , n4289 , n4290 , n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , n4299 , n4300 , n4301 , n4302 , n4303 , n4304 , n4305 , n4306 , n4307 , n4308 , n4309 , n4310 , n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , n4319 , n4320 , n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , n4329 , n4330 , n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , n4340 , n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , n4349 , n4350 , n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , n4360 , n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , n4370 , n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , n4380 , n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , n4390 , n4391 , n4392 , n4393 , n4394 , n4395 , n4396 , n4397 , n4398 , n4399 , n4400 , n4401 , n4402 , n4403 , n4404 , n4405 , n4406 , n4407 , n4408 , n4409 , n4410 , n4411 , n4412 , n4413 , n4414 , n4415 , n4416 , n4417 , n4418 , n4419 , n4420 , n4421 , n4422 , n4423 , n4424 , n4425 , n4426 , n4427 , n4428 , n4429 , n4430 , n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , n4437 , n4438 , n4439 , n4440 , n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , n4449 , n4450 , n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , n4459 , n4460 , n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , n4469 , n4470 , n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , n4479 , n4480 , n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , n4487 , n4488 , n4489 , n4490 , n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , n4497 , n4498 , n4499 , n4500 , n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , n4509 , n4510 , n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , n4519 , n4520 , n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , n4529 , n4530 , n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , n4537 , n4538 , n4539 , n4540 , n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , n4547 , n4548 , n4549 , n4550 , n4551 , n4552 , n4553 , n4554 , n4555 , n4556 , n4557 , n4558 , n4559 , n4560 , n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , n4567 , n4568 , n4569 , n4570 , n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , n4579 , n4580 , n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , n4589 , n4590 , n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , n4597 , n4598 , n4599 , n4600 , n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , n4607 , n4608 , n4609 , n4610 , n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , n4617 , n4618 , n4619 , n4620 , n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , n4627 , n4628 , n4629 , n4630 , n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , n4637 , n4638 , n4639 , n4640 , n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , n4647 , n4648 , n4649 , n4650 , n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , n4657 , n4658 , n4659 , n4660 , n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , n4669 , n4670 , n4671 , n4672 , n4673 , n4674 , n4675 , n4676 , n4677 , n4678 , n4679 , n4680 , n4681 , n4682 , n4683 , n4684 , n4685 , n4686 , n4687 , n4688 , n4689 , n4690 , n4691 , n4692 , n4693 , n4694 , n4695 , n4696 , n4697 , n4698 , n4699 , n4700 , n4701 , n4702 , n4703 , n4704 , n4705 , n4706 , n4707 , n4708 , n4709 , n4710 , n4711 , n4712 , n4713 , n4714 , n4715 , n4716 , n4717 , n4718 , n4719 , n4720 , n4721 , n4722 , n4723 , n4724 , n4725 , n4726 , n4727 , n4728 , n4729 , n4730 , n4731 , n4732 , n4733 , n4734 , n4735 , n4736 , n4737 , n4738 , n4739 , n4740 , n4741 , n4742 , n4743 , n4744 , n4745 , n4746 , n4747 , n4748 , n4749 , n4750 , n4751 , n4752 , n4753 , n4754 , n4755 , n4756 , n4757 , n4758 , n4759 , n4760 , n4761 , n4762 , n4763 , n4764 , n4765 , n4766 , n4767 , n4768 , n4769 , n4770 , n4771 , n4772 , n4773 , n4774 , n4775 , n4776 , n4777 , n4778 , n4779 , n4780 , n4781 , n4782 , n4783 , n4784 , n4785 , n4786 , n4787 , n4788 , n4789 , n4790 , n4791 , n4792 , n4793 , n4794 , n4795 , n4796 , n4797 , n4798 , n4799 , n4800 , n4801 , n4802 , n4803 , n4804 , n4805 , n4806 , n4807 , n4808 , n4809 , n4810 , n4811 , n4812 , n4813 , n4814 , n4815 , n4816 , n4817 , n4818 , n4819 , n4820 , n4821 , n4822 , n4823 , n4824 , n4825 , n4826 , n4827 , n4828 , n4829 , n4830 , n4831 , n4832 , n4833 , n4834 , n4835 , n4836 , n4837 , n4838 , n4839 , n4840 , n4841 , n4842 , n4843 , n4844 , n4845 , n4846 , n4847 , n4848 , n4849 , n4850 , n4851 , n4852 , n4853 , n4854 , n4855 , n4856 , n4857 , n4858 , n4859 , n4860 , n4861 , n4862 , n4863 , n4864 , n4865 , n4866 , n4867 , n4868 , n4869 , n4870 , n4871 , n4872 , n4873 , n4874 , n4875 , n4876 , n4877 , n4878 , n4879 , n4880 , n4881 , n4882 , n4883 , n4884 , n4885 , n4886 , n4887 , n4888 , n4889 , n4890 , n4891 , n4892 , n4893 , n4894 , n4895 , n4896 , n4897 , n4898 , n4899 , n4900 , n4901 , n4902 , n4903 , n4904 , n4905 , n4906 , n4907 , n4908 , n4909 , n4910 , n4911 , n4912 , n4913 , n4914 , n4915 , n4916 , n4917 , n4918 , n4919 , n4920 , n4921 , n4922 , n4923 , n4924 , n4925 , n4926 , n4927 , n4928 , n4929 , n4930 , n4931 , n4932 , n4933 , n4934 , n4935 , n4936 , n4937 , n4938 , n4939 , n4940 , n4941 , n4942 , n4943 , n4944 , n4945 , n4946 , n4947 , n4948 , n4949 , n4950 , n4951 , n4952 , n4953 , n4954 , n4955 , n4956 , n4957 , n4958 , n4959 , n4960 , n4961 , n4962 , n4963 , n4964 , n4965 , n4966 , n4967 , n4968 , n4969 , n4970 , n4971 , n4972 , n4973 , n4974 , n4975 , n4976 , n4977 , n4978 , n4979 , n4980 , n4981 , n4982 , n4983 , n4984 , n4985 , n4986 , n4987 , n4988 , n4989 , n4990 , n4991 , n4992 , n4993 , n4994 , n4995 , n4996 , n4997 , n4998 , n4999 , n5000 , n5001 , n5002 , n5003 , n5004 , n5005 , n5006 , n5007 , n5008 , n5009 , n5010 , n5011 , n5012 , n5013 , n5014 , n5015 , n5016 , n5017 , n5018 , n5019 , n5020 , n5021 , n5022 , n5023 , n5024 , n5025 , n5026 , n5027 , n5028 , n5029 , n5030 , n5031 , n5032 , n5033 , n5034 , n5035 , n5036 , n5037 , n5038 , n5039 , n5040 , n5041 , n5042 , n5043 , n5044 , n5045 , n5046 , n5047 , n5048 , n5049 , n5050 , n5051 , n5052 , n5053 , n5054 , n5055 , n5056 , n5057 , n5058 , n5059 , n5060 , n5061 , n5062 , n5063 , n5064 , n5065 , n5066 , n5067 , n5068 , n5069 , n5070 , n5071 , n5072 , n5073 , n5074 , n5075 , n5076 , n5077 , n5078 , n5079 , n5080 , n5081 , n5082 , n5083 , n5084 , n5085 , n5086 , n5087 , n5088 , n5089 , n5090 , n5091 , n5092 , n5093 , n5094 , n5095 , n5096 , n5097 , n5098 , n5099 , n5100 , n5101 , n5102 , n5103 , n5104 , n5105 , n5106 , n5107 , n5108 , n5109 , n5110 , n5111 , n5112 , n5113 , n5114 , n5115 , n5116 , n5117 , n5118 , n5119 , n5120 , n5121 , n5122 , n5123 , n5124 , n5125 , n5126 , n5127 , n5128 , n5129 , n5130 , n5131 , n5132 , n5133 , n5134 , n5135 , n5136 , n5137 , n5138 , n5139 , n5140 , n5141 , n5142 , n5143 , n5144 , n5145 , n5146 , n5147 , n5148 , n5149 , n5150 , n5151 , n5152 , n5153 , n5154 , n5155 , n5156 , n5157 , n5158 , n5159 , n5160 , n5161 , n5162 , n5163 , n5164 , n5165 , n5166 , n5167 , n5168 , n5169 , n5170 , n5171 , n5172 , n5173 , n5174 , n5175 , n5176 , n5177 , n5178 , n5179 , n5180 , n5181 , n5182 , n5183 , n5184 , n5185 , n5186 , n5187 , n5188 , n5189 , n5190 , n5191 , n5192 , n5193 , n5194 , n5195 , n5196 , n5197 , n5198 , n5199 , n5200 , n5201 , n5202 , n5203 , n5204 , n5205 , n5206 , n5207 , n5208 , n5209 , n5210 , n5211 , n5212 , n5213 , n5214 , n5215 , n5216 , n5217 , n5218 , n5219 , n5220 , n5221 , n5222 , n5223 , n5224 , n5225 , n5226 , n5227 , n5228 , n5229 , n5230 , n5231 , n5232 , n5233 , n5234 , n5235 , n5236 , n5237 , n5238 , n5239 , n5240 , n5241 , n5242 , n5243 , n5244 , n5245 , n5246 , n5247 , n5248 , n5249 , n5250 , n5251 , n5252 , n5253 , n5254 , n5255 , n5256 , n5257 , n5258 , n5259 , n5260 , n5261 , n5262 , n5263 , n5264 , n5265 , n5266 , n5267 , n5268 , n5269 , n5270 , n5271 , n5272 , n5273 , n5274 , n5275 , n5276 , n5277 , n5278 , n5279 , n5280 , n5281 , n5282 , n5283 , n5284 , n5285 , n5286 , n5287 , n5288 , n5289 , n5290 , n5291 , n5292 , n5293 , n5294 , n5295 , n5296 , n5297 , n5298 , n5299 , n5300 , n5301 , n5302 , n5303 , n5304 , n5305 , n5306 , n5307 , n5308 , n5309 , n5310 , n5311 , n5312 , n5313 , n5314 , n5315 , n5316 , n5317 , n5318 , n5319 , n5320 , n5321 , n5322 , n5323 , n5324 , n5325 , n5326 , n5327 , n5328 , n5329 , n5330 , n5331 , n5332 , n5333 , n5334 , n5335 , n5336 , n5337 , n5338 , n5339 , n5340 , n5341 , n5342 , n5343 , n5344 , n5345 , n5346 , n5347 , n5348 , n5349 , n5350 , n5351 , n5352 , n5353 , n5354 , n5355 , n5356 , n5357 , n5358 , n5359 , n5360 , n5361 , n5362 , n5363 , n5364 , n5365 , n5366 , n5367 , n5368 , n5369 , n5370 , n5371 , n5372 , n5373 , n5374 , n5375 , n5376 , n5377 , n5378 , n5379 , n5380 , n5381 , n5382 , n5383 , n5384 , n5385 , n5386 , n5387 , n5388 , n5389 , n5390 , n5391 , n5392 , n5393 , n5394 , n5395 , n5396 , n5397 , n5398 , n5399 , n5400 , n5401 , n5402 , n5403 , n5404 , n5405 , n5406 , n5407 , n5408 , n5409 , n5410 , n5411 , n5412 , n5413 , n5414 , n5415 , n5416 , n5417 , n5418 , n5419 , n5420 , n5421 , n5422 , n5423 , n5424 , n5425 , n5426 , n5427 , n5428 , n5429 , n5430 , n5431 , n5432 , n5433 , n5434 , n5435 , n5436 , n5437 , n5438 , n5439 , n5440 , n5441 , n5442 , n5443 , n5444 , n5445 , n5446 , n5447 , n5448 , n5449 , n5450 , n5451 , n5452 , n5453 , n5454 , n5455 , n5456 , n5457 , n5458 , n5459 , n5460 , n5461 , n5462 , n5463 , n5464 , n5465 , n5466 , n5467 , n5468 , n5469 , n5470 , n5471 , n5472 , n5473 , n5474 , n5475 , n5476 , n5477 , n5478 , n5479 , n5480 , n5481 , n5482 , n5483 , n5484 , n5485 , n5486 , n5487 , n5488 , n5489 , n5490 , n5491 , n5492 , n5493 , n5494 , n5495 , n5496 , n5497 , n5498 , n5499 , n5500 , n5501 , n5502 , n5503 , n5504 , n5505 , n5506 , n5507 , n5508 , n5509 , n5510 , n5511 , n5512 , n5513 , n5514 , n5515 , n5516 , n5517 , n5518 , n5519 , n5520 , n5521 , n5522 , n5523 , n5524 , n5525 , n5526 , n5527 , n5528 , n5529 , n5530 , n5531 , n5532 , n5533 , n5534 , n5535 , n5536 , n5537 , n5538 , n5539 , n5540 , n5541 , n5542 , n5543 , n5544 , n5545 , n5546 , n5547 , n5548 , n5549 , n5550 , n5551 , n5552 , n5553 , n5554 , n5555 , n5556 , n5557 , n5558 , n5559 , n5560 , n5561 , n5562 , n5563 , n5564 , n5565 , n5566 , n5567 , n5568 , n5569 , n5570 , n5571 , n5572 , n5573 , n5574 , n5575 , n5576 , n5577 , n5578 , n5579 , n5580 , n5581 , n5582 , n5583 , n5584 , n5585 , n5586 , n5587 , n5588 , n5589 , n5590 , n5591 , n5592 , n5593 , n5594 , n5595 , n5596 , n5597 , n5598 , n5599 , n5600 , n5601 , n5602 , n5603 , n5604 , n5605 , n5606 , n5607 , n5608 , n5609 , n5610 , n5611 , n5612 , n5613 , n5614 , n5615 , n5616 , n5617 , n5618 , n5619 , n5620 , n5621 , n5622 , n5623 , n5624 , n5625 , n5626 , n5627 , n5628 , n5629 , n5630 , n5631 , n5632 , n5633 , n5634 , n5635 , n5636 , n5637 , n5638 , n5639 , n5640 , n5641 , n5642 , n5643 , n5644 , n5645 , n5646 , n5647 , n5648 , n5649 , n5650 , n5651 , n5652 , n5653 , n5654 , n5655 , n5656 , n5657 , n5658 , n5659 , n5660 , n5661 , n5662 , n5663 , n5664 , n5665 , n5666 , n5667 , n5668 , n5669 , n5670 , n5671 , n5672 , n5673 , n5674 , n5675 , n5676 , n5677 , n5678 , n5679 , n5680 , n5681 , n5682 , n5683 , n5684 , n5685 , n5686 , n5687 , n5688 , n5689 , n5690 , n5691 , n5692 , n5693 , n5694 , n5695 , n5696 , n5697 , n5698 , n5699 , n5700 , n5701 , n5702 , n5703 , n5704 , n5705 , n5706 , n5707 , n5708 , n5709 , n5710 , n5711 , n5712 , n5713 , n5714 , n5715 , n5716 , n5717 , n5718 , n5719 , n5720 , n5721 , n5722 , n5723 , n5724 , n5725 , n5726 , n5727 , n5728 , n5729 , n5730 , n5731 , n5732 , n5733 , n5734 , n5735 , n5736 , n5737 , n5738 , n5739 , n5740 , n5741 , n5742 , n5743 , n5744 , n5745 , n5746 , n5747 , n5748 , n5749 , n5750 , n5751 , n5752 , n5753 , n5754 , n5755 , n5756 , n5757 , n5758 , n5759 , n5760 , n5761 , n5762 , n5763 , n5764 , n5765 , n5766 , n5767 , n5768 , n5769 , n5770 , n5771 , n5772 , n5773 , n5774 , n5775 , n5776 , n5777 , n5778 , n5779 , n5780 , n5781 , n5782 , n5783 , n5784 , n5785 , n5786 , n5787 , n5788 , n5789 , n5790 , n5791 , n5792 , n5793 , n5794 , n5795 , n5796 , n5797 , n5798 , n5799 , n5800 , n5801 , n5802 , n5803 , n5804 , n5805 , n5806 , n5807 , n5808 , n5809 , n5810 , n5811 , n5812 , n5813 , n5814 , n5815 , n5816 , n5817 , n5818 , n5819 , n5820 , n5821 , n5822 , n5823 , n5824 , n5825 , n5826 , n5827 , n5828 , n5829 , n5830 , n5831 , n5832 , n5833 , n5834 , n5835 , n5836 , n5837 , n5838 , n5839 , n5840 , n5841 , n5842 , n5843 , n5844 , n5845 , n5846 , n5847 , n5848 , n5849 , n5850 , n5851 , n5852 , n5853 , n5854 , n5855 , n5856 , n5857 , n5858 , n5859 , n5860 , n5861 , n5862 , n5863 , n5864 , n5865 , n5866 , n5867 , n5868 , n5869 , n5870 , n5871 , n5872 , n5873 , n5874 , n5875 , n5876 , n5877 , n5878 , n5879 , n5880 , n5881 , n5882 , n5883 , n5884 , n5885 , n5886 , n5887 , n5888 , n5889 , n5890 , n5891 , n5892 , n5893 , n5894 , n5895 , n5896 , n5897 , n5898 , n5899 , n5900 , n5901 , n5902 , n5903 , n5904 , n5905 , n5906 , n5907 , n5908 , n5909 , n5910 , n5911 , n5912 , n5913 , n5914 , n5915 , n5916 , n5917 , n5918 , n5919 , n5920 , n5921 , n5922 , n5923 , n5924 , n5925 , n5926 , n5927 , n5928 , n5929 , n5930 , n5931 , n5932 , n5933 , n5934 , n5935 , n5936 , n5937 , n5938 , n5939 , n5940 , n5941 , n5942 , n5943 , n5944 , n5945 , n5946 , n5947 , n5948 , n5949 , n5950 , n5951 , n5952 , n5953 , n5954 , n5955 , n5956 , n5957 , n5958 , n5959 , n5960 , n5961 , n5962 , n5963 , n5964 , n5965 , n5966 , n5967 , n5968 , n5969 , n5970 , n5971 , n5972 , n5973 , n5974 , n5975 , n5976 , n5977 , n5978 , n5979 , n5980 , n5981 , n5982 , n5983 , n5984 , n5985 , n5986 , n5987 , n5988 , n5989 , n5990 , n5991 , n5992 , n5993 , n5994 , n5995 , n5996 , n5997 , n5998 , n5999 , n6000 , n6001 , n6002 , n6003 , n6004 , n6005 , n6006 , n6007 , n6008 , n6009 , n6010 , n6011 , n6012 , n6013 , n6014 , n6015 , n6016 , n6017 , n6018 , n6019 , n6020 , n6021 , n6022 , n6023 , n6024 , n6025 , n6026 , n6027 , n6028 , n6029 , n6030 , n6031 , n6032 , n6033 , n6034 , n6035 , n6036 , n6037 , n6038 , n6039 , n6040 , n6041 , n6042 , n6043 , n6044 , n6045 , n6046 , n6047 , n6048 , n6049 , n6050 , n6051 , n6052 , n6053 , n6054 , n6055 , n6056 , n6057 , n6058 , n6059 , n6060 , n6061 , n6062 , n6063 , n6064 , n6065 , n6066 , n6067 , n6068 , n6069 , n6070 , n6071 , n6072 , n6073 , n6074 , n6075 , n6076 , n6077 , n6078 , n6079 , n6080 , n6081 , n6082 , n6083 , n6084 , n6085 , n6086 , n6087 , n6088 , n6089 , n6090 , n6091 , n6092 , n6093 , n6094 , n6095 , n6096 , n6097 , n6098 , n6099 , n6100 , n6101 , n6102 , n6103 , n6104 , n6105 , n6106 , n6107 , n6108 , n6109 , n6110 , n6111 , n6112 , n6113 , n6114 , n6115 , n6116 , n6117 , n6118 , n6119 , n6120 , n6121 , n6122 , n6123 , n6124 , n6125 , n6126 , n6127 , n6128 , n6129 , n6130 , n6131 , n6132 , n6133 , n6134 , n6135 , n6136 , n6137 , n6138 , n6139 , n6140 , n6141 , n6142 , n6143 , n6144 , n6145 , n6146 , n6147 , n6148 , n6149 , n6150 , n6151 , n6152 , n6153 , n6154 , n6155 , n6156 , n6157 , n6158 , n6159 , n6160 , n6161 , n6162 , n6163 , n6164 , n6165 , n6166 , n6167 , n6168 , n6169 , n6170 , n6171 , n6172 , n6173 , n6174 , n6175 , n6176 , n6177 , n6178 , n6179 , n6180 , n6181 , n6182 , n6183 , n6184 , n6185 , n6186 , n6187 , n6188 , n6189 , n6190 , n6191 , n6192 , n6193 , n6194 , n6195 , n6196 , n6197 , n6198 , n6199 , n6200 , n6201 , n6202 , n6203 , n6204 , n6205 , n6206 , n6207 , n6208 , n6209 , n6210 , n6211 , n6212 , n6213 , n6214 , n6215 , n6216 , n6217 , n6218 , n6219 , n6220 , n6221 , n6222 , n6223 , n6224 , n6225 , n6226 , n6227 , n6228 , n6229 , n6230 , n6231 , n6232 , n6233 , n6234 , n6235 , n6236 , n6237 , n6238 , n6239 , n6240 , n6241 , n6242 , n6243 , n6244 , n6245 , n6246 , n6247 , n6248 , n6249 , n6250 , n6251 , n6252 , n6253 , n6254 , n6255 , n6256 , n6257 , n6258 , n6259 , n6260 , n6261 , n6262 , n6263 , n6264 , n6265 , n6266 , n6267 , n6268 , n6269 , n6270 , n6271 , n6272 , n6273 , n6274 , n6275 , n6276 , n6277 , n6278 , n6279 , n6280 , n6281 , n6282 , n6283 , n6284 , n6285 , n6286 , n6287 , n6288 , n6289 , n6290 , n6291 , n6292 , n6293 , n6294 , n6295 , n6296 , n6297 , n6298 , n6299 , n6300 , n6301 , n6302 , n6303 , n6304 , n6305 , n6306 , n6307 , n6308 , n6309 , n6310 , n6311 , n6312 , n6313 , n6314 , n6315 , n6316 , n6317 , n6318 , n6319 , n6320 , n6321 , n6322 , n6323 , n6324 , n6325 , n6326 , n6327 , n6328 , n6329 , n6330 , n6331 , n6332 , n6333 , n6334 , n6335 , n6336 , n6337 , n6338 , n6339 , n6340 , n6341 , n6342 , n6343 , n6344 , n6345 , n6346 , n6347 , n6348 , n6349 , n6350 , n6351 , n6352 , n6353 , n6354 , n6355 , n6356 , n6357 , n6358 , n6359 , n6360 , n6361 , n6362 , n6363 , n6364 , n6365 , n6366 , n6367 , n6368 , n6369 , n6370 , n6371 , n6372 , n6373 , n6374 , n6375 , n6376 , n6377 , n6378 , n6379 , n6380 , n6381 , n6382 , n6383 , n6384 , n6385 , n6386 , n6387 , n6388 , n6389 , n6390 , n6391 , n6392 , n6393 , n6394 , n6395 , n6396 , n6397 , n6398 , n6399 , n6400 , n6401 , n6402 , n6403 , n6404 , n6405 , n6406 , n6407 , n6408 , n6409 , n6410 , n6411 , n6412 , n6413 , n6414 , n6415 , n6416 , n6417 , n6418 , n6419 , n6420 , n6421 , n6422 , n6423 , n6424 , n6425 , n6426 , n6427 , n6428 , n6429 , n6430 , n6431 , n6432 , n6433 , n6434 , n6435 , n6436 , n6437 , n6438 , n6439 , n6440 , n6441 , n6442 , n6443 , n6444 , n6445 , n6446 , n6447 , n6448 , n6449 , n6450 , n6451 , n6452 , n6453 , n6454 , n6455 , n6456 , n6457 , n6458 , n6459 , n6460 , n6461 , n6462 , n6463 , n6464 , n6465 , n6466 , n6467 , n6468 , n6469 , n6470 , n6471 , n6472 , n6473 , n6474 , n6475 , n6476 , n6477 , n6478 , n6479 , n6480 , n6481 , n6482 , n6483 , n6484 , n6485 , n6486 , n6487 , n6488 , n6489 , n6490 , n6491 , n6492 , n6493 , n6494 , n6495 , n6496 , n6497 , n6498 , n6499 , n6500 , n6501 , n6502 , n6503 , n6504 , n6505 , n6506 , n6507 , n6508 , n6509 , n6510 , n6511 , n6512 , n6513 , n6514 , n6515 , n6516 , n6517 , n6518 , n6519 , n6520 , n6521 , n6522 , n6523 , n6524 , n6525 , n6526 , n6527 , n6528 , n6529 , n6530 , n6531 , n6532 , n6533 , n6534 , n6535 , n6536 , n6537 , n6538 , n6539 , n6540 , n6541 , n6542 , n6543 , n6544 , n6545 , n6546 , n6547 , n6548 , n6549 , n6550 , n6551 , n6552 , n6553 , n6554 , n6555 , n6556 , n6557 , n6558 , n6559 , n6560 , n6561 , n6562 , n6563 , n6564 , n6565 , n6566 , n6567 , n6568 , n6569 , n6570 , n6571 , n6572 , n6573 , n6574 , n6575 , n6576 , n6577 , n6578 , n6579 , n6580 , n6581 , n6582 , n6583 , n6584 , n6585 , n6586 , n6587 , n6588 , n6589 , n6590 , n6591 , n6592 , n6593 , n6594 , n6595 , n6596 , n6597 , n6598 , n6599 , n6600 , n6601 , n6602 , n6603 , n6604 , n6605 , n6606 , n6607 , n6608 , n6609 , n6610 , n6611 , n6612 , n6613 , n6614 , n6615 , n6616 , n6617 , n6618 , n6619 , n6620 , n6621 , n6622 , n6623 , n6624 , n6625 , n6626 , n6627 , n6628 , n6629 , n6630 , n6631 , n6632 , n6633 , n6634 , n6635 , n6636 , n6637 , n6638 , n6639 , n6640 , n6641 , n6642 , n6643 , n6644 , n6645 , n6646 , n6647 , n6648 , n6649 , n6650 , n6651 , n6652 , n6653 , n6654 , n6655 , n6656 , n6657 , n6658 , n6659 , n6660 , n6661 , n6662 , n6663 , n6664 , n6665 , n6666 , n6667 , n6668 , n6669 , n6670 , n6671 , n6672 , n6673 , n6674 , n6675 , n6676 , n6677 , n6678 , n6679 , n6680 , n6681 , n6682 , n6683 , n6684 , n6685 , n6686 , n6687 , n6688 , n6689 , n6690 , n6691 , n6692 , n6693 , n6694 , n6695 , n6696 , n6697 , n6698 , n6699 , n6700 , n6701 , n6702 , n6703 , n6704 , n6705 , n6706 , n6707 , n6708 , n6709 , n6710 , n6711 , n6712 , n6713 , n6714 , n6715 , n6716 , n6717 , n6718 , n6719 , n6720 , n6721 , n6722 , n6723 , n6724 , n6725 , n6726 , n6727 , n6728 , n6729 , n6730 , n6731 , n6732 , n6733 , n6734 , n6735 , n6736 , n6737 , n6738 , n6739 , n6740 , n6741 , n6742 , n6743 , n6744 , n6745 , n6746 , n6747 , n6748 , n6749 , n6750 , n6751 , n6752 , n6753 , n6754 , n6755 , n6756 , n6757 , n6758 , n6759 , n6760 , n6761 , n6762 , n6763 , n6764 , n6765 , n6766 , n6767 , n6768 , n6769 , n6770 , n6771 , n6772 , n6773 , n6774 , n6775 , n6776 , n6777 , n6778 , n6779 , n6780 , n6781 , n6782 , n6783 , n6784 , n6785 , n6786 , n6787 , n6788 , n6789 , n6790 , n6791 , n6792 , n6793 , n6794 , n6795 , n6796 , n6797 , n6798 , n6799 , n6800 , n6801 , n6802 , n6803 , n6804 , n6805 , n6806 , n6807 , n6808 , n6809 , n6810 , n6811 , n6812 , n6813 , n6814 , n6815 , n6816 , n6817 , n6818 , n6819 , n6820 , n6821 , n6822 , n6823 , n6824 , n6825 , n6826 , n6827 , n6828 , n6829 , n6830 , n6831 , n6832 , n6833 , n6834 , n6835 , n6836 , n6837 , n6838 , n6839 , n6840 , n6841 , n6842 , n6843 , n6844 , n6845 , n6846 , n6847 , n6848 , n6849 , n6850 , n6851 , n6852 , n6853 , n6854 , n6855 , n6856 , n6857 , n6858 , n6859 , n6860 , n6861 , n6862 , n6863 , n6864 , n6865 , n6866 , n6867 , n6868 , n6869 , n6870 , n6871 , n6872 , n6873 , n6874 , n6875 , n6876 , n6877 , n6878 , n6879 , n6880 , n6881 , n6882 , n6883 , n6884 , n6885 , n6886 , n6887 , n6888 , n6889 , n6890 , n6891 , n6892 , n6893 , n6894 , n6895 , n6896 , n6897 , n6898 , n6899 , n6900 , n6901 , n6902 , n6903 , n6904 , n6905 , n6906 , n6907 , n6908 , n6909 , n6910 , n6911 , n6912 , n6913 , n6914 , n6915 , n6916 , n6917 , n6918 , n6919 , n6920 , n6921 , n6922 , n6923 , n6924 , n6925 , n6926 , n6927 , n6928 , n6929 , n6930 , n6931 , n6932 , n6933 , n6934 , n6935 , n6936 , n6937 , n6938 , n6939 , n6940 , n6941 , n6942 , n6943 , n6944 , n6945 , n6946 , n6947 , n6948 , n6949 , n6950 , n6951 , n6952 , n6953 , n6954 , n6955 , n6956 , n6957 , n6958 , n6959 , n6960 , n6961 , n6962 , n6963 , n6964 , n6965 , n6966 , n6967 , n6968 , n6969 , n6970 , n6971 , n6972 , n6973 , n6974 , n6975 , n6976 , n6977 , n6978 , n6979 , n6980 , n6981 , n6982 , n6983 , n6984 , n6985 , n6986 , n6987 , n6988 , n6989 , n6990 , n6991 , n6992 , n6993 , n6994 , n6995 , n6996 , n6997 , n6998 , n6999 , n7000 , n7001 , n7002 , n7003 , n7004 , n7005 , n7006 , n7007 , n7008 , n7009 , n7010 , n7011 , n7012 , n7013 , n7014 , n7015 , n7016 , n7017 , n7018 , n7019 , n7020 , n7021 , n7022 , n7023 , n7024 , n7025 , n7026 , n7027 , n7028 , n7029 , n7030 , n7031 , n7032 , n7033 , n7034 , n7035 , n7036 , n7037 , n7038 , n7039 , n7040 , n7041 , n7042 , n7043 , n7044 , n7045 , n7046 , n7047 , n7048 , n7049 , n7050 , n7051 , n7052 , n7053 , n7054 , n7055 , n7056 , n7057 , n7058 , n7059 , n7060 , n7061 , n7062 , n7063 , n7064 , n7065 , n7066 , n7067 , n7068 , n7069 , n7070 , n7071 , n7072 , n7073 , n7074 , n7075 , n7076 , n7077 , n7078 , n7079 , n7080 , n7081 , n7082 , n7083 , n7084 , n7085 , n7086 , n7087 , n7088 , n7089 , n7090 , n7091 , n7092 , n7093 , n7094 , n7095 , n7096 , n7097 , n7098 , n7099 , n7100 , n7101 , n7102 , n7103 , n7104 , n7105 , n7106 , n7107 , n7108 , n7109 , n7110 , n7111 , n7112 , n7113 , n7114 , n7115 , n7116 , n7117 , n7118 , n7119 , n7120 , n7121 , n7122 , n7123 , n7124 , n7125 , n7126 , n7127 , n7128 , n7129 , n7130 , n7131 , n7132 , n7133 , n7134 , n7135 , n7136 , n7137 , n7138 , n7139 , n7140 , n7141 , n7142 , n7143 , n7144 , n7145 , n7146 , n7147 , n7148 , n7149 , n7150 , n7151 , n7152 , n7153 , n7154 , n7155 , n7156 , n7157 , n7158 , n7159 , n7160 , n7161 , n7162 , n7163 , n7164 , n7165 , n7166 , n7167 , n7168 , n7169 , n7170 , n7171 , n7172 , n7173 , n7174 , n7175 , n7176 , n7177 , n7178 , n7179 , n7180 , n7181 , n7182 , n7183 , n7184 , n7185 , n7186 , n7187 , n7188 , n7189 , n7190 , n7191 , n7192 , n7193 , n7194 , n7195 , n7196 , n7197 , n7198 , n7199 , n7200 , n7201 , n7202 , n7203 , n7204 , n7205 , n7206 , n7207 , n7208 , n7209 , n7210 , n7211 , n7212 , n7213 , n7214 , n7215 , n7216 , n7217 , n7218 , n7219 , n7220 , n7221 , n7222 , n7223 , n7224 , n7225 , n7226 , n7227 , n7228 , n7229 , n7230 , n7231 , n7232 , n7233 , n7234 , n7235 , n7236 , n7237 , n7238 , n7239 , n7240 , n7241 , n7242 , n7243 , n7244 , n7245 , n7246 , n7247 , n7248 , n7249 , n7250 , n7251 , n7252 , n7253 , n7254 , n7255 , n7256 , n7257 , n7258 , n7259 , n7260 , n7261 , n7262 , n7263 , n7264 , n7265 , n7266 , n7267 , n7268 , n7269 , n7270 , n7271 , n7272 , n7273 , n7274 , n7275 , n7276 , n7277 , n7278 , n7279 , n7280 , n7281 , n7282 , n7283 , n7284 , n7285 , n7286 , n7287 , n7288 , n7289 , n7290 , n7291 , n7292 , n7293 , n7294 , n7295 , n7296 , n7297 , n7298 , n7299 , n7300 , n7301 , n7302 , n7303 , n7304 , n7305 , n7306 , n7307 , n7308 , n7309 , n7310 , n7311 , n7312 , n7313 , n7314 , n7315 , n7316 , n7317 , n7318 , n7319 , n7320 , n7321 , n7322 , n7323 , n7324 , n7325 , n7326 , n7327 , n7328 , n7329 , n7330 , n7331 , n7332 , n7333 , n7334 , n7335 , n7336 , n7337 , n7338 , n7339 , n7340 , n7341 , n7342 , n7343 , n7344 , n7345 , n7346 , n7347 , n7348 , n7349 , n7350 , n7351 , n7352 , n7353 , n7354 , n7355 , n7356 , n7357 , n7358 , n7359 , n7360 , n7361 , n7362 , n7363 , n7364 , n7365 , n7366 , n7367 , n7368 , n7369 , n7370 , n7371 , n7372 , n7373 , n7374 , n7375 , n7376 , n7377 , n7378 , n7379 , n7380 , n7381 , n7382 , n7383 , n7384 , n7385 , n7386 , n7387 , n7388 , n7389 , n7390 , n7391 , n7392 , n7393 , n7394 , n7395 , n7396 , n7397 , n7398 , n7399 , n7400 , n7401 , n7402 , n7403 , n7404 , n7405 , n7406 , n7407 , n7408 , n7409 , n7410 , n7411 , n7412 , n7413 , n7414 , n7415 , n7416 , n7417 , n7418 , n7419 , n7420 , n7421 , n7422 , n7423 , n7424 , n7425 , n7426 , n7427 , n7428 , n7429 , n7430 , n7431 , n7432 , n7433 , n7434 , n7435 , n7436 , n7437 , n7438 , n7439 , n7440 , n7441 , n7442 , n7443 , n7444 , n7445 , n7446 , n7447 , n7448 , n7449 , n7450 , n7451 , n7452 , n7453 , n7454 , n7455 , n7456 , n7457 , n7458 , n7459 , n7460 , n7461 , n7462 , n7463 , n7464 , n7465 , n7466 , n7467 , n7468 , n7469 , n7470 , n7471 , n7472 , n7473 , n7474 , n7475 , n7476 , n7477 , n7478 , n7479 , n7480 , n7481 , n7482 , n7483 , n7484 , n7485 , n7486 , n7487 , n7488 , n7489 , n7490 , n7491 , n7492 , n7493 , n7494 , n7495 , n7496 , n7497 , n7498 , n7499 , n7500 , n7501 , n7502 , n7503 , n7504 , n7505 , n7506 , n7507 , n7508 , n7509 , n7510 , n7511 , n7512 , n7513 , n7514 , n7515 , n7516 , n7517 , n7518 , n7519 , n7520 , n7521 , n7522 , n7523 , n7524 , n7525 , n7526 , n7527 , n7528 , n7529 , n7530 , n7531 , n7532 , n7533 , n7534 , n7535 , n7536 , n7537 , n7538 , n7539 , n7540 , n7541 , n7542 , n7543 , n7544 , n7545 , n7546 , n7547 , n7548 , n7549 , n7550 , n7551 , n7552 , n7553 , n7554 , n7555 , n7556 , n7557 , n7558 , n7559 , n7560 , n7561 , n7562 , n7563 , n7564 , n7565 , n7566 , n7567 , n7568 , n7569 , n7570 , n7571 , n7572 , n7573 , n7574 , n7575 , n7576 , n7577 , n7578 , n7579 , n7580 , n7581 , n7582 , n7583 , n7584 , n7585 , n7586 , n7587 , n7588 , n7589 , n7590 , n7591 , n7592 , n7593 , n7594 , n7595 , n7596 , n7597 , n7598 , n7599 , n7600 , n7601 , n7602 , n7603 , n7604 , n7605 , n7606 , n7607 , n7608 , n7609 , n7610 , n7611 , n7612 , n7613 , n7614 , n7615 , n7616 , n7617 , n7618 , n7619 , n7620 , n7621 , n7622 , n7623 , n7624 , n7625 , n7626 , n7627 , n7628 , n7629 , n7630 , n7631 , n7632 , n7633 , n7634 , n7635 , n7636 , n7637 , n7638 , n7639 , n7640 , n7641 , n7642 , n7643 , n7644 , n7645 , n7646 , n7647 , n7648 , n7649 , n7650 , n7651 , n7652 , n7653 , n7654 , n7655 , n7656 , n7657 , n7658 , n7659 , n7660 , n7661 , n7662 , n7663 , n7664 , n7665 , n7666 , n7667 , n7668 , n7669 , n7670 , n7671 , n7672 , n7673 , n7674 , n7675 , n7676 , n7677 , n7678 , n7679 , n7680 , n7681 , n7682 , n7683 , n7684 , n7685 , n7686 , n7687 , n7688 , n7689 , n7690 , n7691 , n7692 , n7693 , n7694 , n7695 , n7696 , n7697 , n7698 , n7699 , n7700 , n7701 , n7702 , n7703 , n7704 , n7705 , n7706 , n7707 , n7708 , n7709 , n7710 , n7711 , n7712 , n7713 , n7714 , n7715 , n7716 , n7717 , n7718 , n7719 , n7720 , n7721 , n7722 , n7723 , n7724 , n7725 , n7726 , n7727 , n7728 , n7729 , n7730 , n7731 , n7732 , n7733 , n7734 , n7735 , n7736 , n7737 , n7738 , n7739 , n7740 , n7741 , n7742 , n7743 , n7744 , n7745 , n7746 , n7747 , n7748 , n7749 , n7750 , n7751 , n7752 , n7753 , n7754 , n7755 , n7756 , n7757 , n7758 , n7759 , n7760 , n7761 , n7762 , n7763 , n7764 , n7765 , n7766 , n7767 , n7768 , n7769 , n7770 , n7771 , n7772 , n7773 , n7774 , n7775 , n7776 , n7777 , n7778 , n7779 , n7780 , n7781 , n7782 , n7783 , n7784 , n7785 , n7786 , n7787 , n7788 , n7789 , n7790 , n7791 , n7792 , n7793 , n7794 , n7795 , n7796 , n7797 , n7798 , n7799 , n7800 , n7801 , n7802 , n7803 , n7804 , n7805 , n7806 , n7807 , n7808 , n7809 , n7810 , n7811 , n7812 , n7813 , n7814 , n7815 , n7816 , n7817 , n7818 , n7819 , n7820 , n7821 , n7822 , n7823 , n7824 , n7825 , n7826 , n7827 , n7828 , n7829 , n7830 , n7831 , n7832 , n7833 , n7834 , n7835 , n7836 , n7837 , n7838 , n7839 , n7840 , n7841 , n7842 , n7843 , n7844 , n7845 , n7846 , n7847 , n7848 , n7849 , n7850 , n7851 , n7852 , n7853 , n7854 , n7855 , n7856 , n7857 , n7858 , n7859 , n7860 , n7861 , n7862 , n7863 , n7864 , n7865 , n7866 , n7867 , n7868 , n7869 , n7870 , n7871 , n7872 , n7873 , n7874 , n7875 , n7876 , n7877 , n7878 , n7879 , n7880 , n7881 , n7882 , n7883 , n7884 , n7885 , n7886 , n7887 , n7888 , n7889 , n7890 , n7891 , n7892 , n7893 , n7894 , n7895 , n7896 , n7897 , n7898 , n7899 , n7900 , n7901 , n7902 , n7903 , n7904 , n7905 , n7906 , n7907 , n7908 , n7909 , n7910 , n7911 , n7912 , n7913 , n7914 , n7915 , n7916 , n7917 , n7918 , n7919 , n7920 , n7921 , n7922 , n7923 , n7924 , n7925 , n7926 , n7927 , n7928 , n7929 , n7930 , n7931 , n7932 , n7933 , n7934 , n7935 , n7936 , n7937 , n7938 , n7939 , n7940 , n7941 , n7942 , n7943 , n7944 , n7945 , n7946 , n7947 , n7948 , n7949 , n7950 , n7951 , n7952 , n7953 , n7954 , n7955 , n7956 , n7957 , n7958 , n7959 , n7960 , n7961 , n7962 , n7963 , n7964 , n7965 , n7966 , n7967 , n7968 , n7969 , n7970 , n7971 , n7972 , n7973 , n7974 , n7975 , n7976 , n7977 , n7978 , n7979 , n7980 , n7981 , n7982 , n7983 , n7984 , n7985 , n7986 , n7987 , n7988 , n7989 , n7990 , n7991 , n7992 , n7993 , n7994 , n7995 , n7996 , n7997 , n7998 , n7999 , n8000 , n8001 , n8002 , n8003 , n8004 , n8005 , n8006 , n8007 , n8008 , n8009 , n8010 , n8011 , n8012 , n8013 , n8014 , n8015 , n8016 , n8017 , n8018 , n8019 , n8020 , n8021 , n8022 , n8023 , n8024 , n8025 , n8026 , n8027 , n8028 , n8029 , n8030 , n8031 , n8032 , n8033 , n8034 , n8035 , n8036 , n8037 , n8038 , n8039 , n8040 , n8041 , n8042 , n8043 , n8044 , n8045 , n8046 , n8047 , n8048 , n8049 , n8050 , n8051 , n8052 , n8053 , n8054 , n8055 , n8056 , n8057 , n8058 , n8059 , n8060 , n8061 , n8062 , n8063 , n8064 , n8065 , n8066 , n8067 , n8068 , n8069 , n8070 , n8071 , n8072 , n8073 , n8074 , n8075 , n8076 , n8077 , n8078 , n8079 , n8080 , n8081 , n8082 , n8083 , n8084 , n8085 , n8086 , n8087 , n8088 , n8089 , n8090 , n8091 , n8092 , n8093 , n8094 , n8095 , n8096 , n8097 , n8098 , n8099 , n8100 , n8101 , n8102 , n8103 , n8104 , n8105 , n8106 , n8107 , n8108 , n8109 , n8110 , n8111 , n8112 , n8113 , n8114 , n8115 , n8116 , n8117 , n8118 , n8119 , n8120 , n8121 , n8122 , n8123 , n8124 , n8125 , n8126 , n8127 , n8128 , n8129 , n8130 , n8131 , n8132 , n8133 , n8134 ;
  assign n25 = x1 | x2 ;
  assign n26 = x0 | x3 ;
  assign n27 = n25 | n26 ;
  assign n28 = x4 | x5 ;
  assign n29 = x6 | n28 ;
  assign n30 = n27 | n29 ;
  assign n31 = x7 | x8 ;
  assign n32 = x9 | x10 ;
  assign n33 = n31 | n32 ;
  assign n34 = n30 | n33 ;
  assign n35 = x16 & ~x22 ;
  assign n36 = x17 & ~n35 ;
  assign n37 = x17 & x22 ;
  assign n38 = x11 | x12 ;
  assign n39 = x13 | x14 ;
  assign n40 = n38 | n39 ;
  assign n41 = x15 | n40 ;
  assign n42 = ( n36 & n37 ) | ( n36 & ~n41 ) | ( n37 & ~n41 ) ;
  assign n43 = n36 & n37 ;
  assign n44 = ( ~n34 & n42 ) | ( ~n34 & n43 ) | ( n42 & n43 ) ;
  assign n45 = ~x17 & n35 ;
  assign n46 = x17 | x22 ;
  assign n47 = ( n41 & n45 ) | ( n41 & ~n46 ) | ( n45 & ~n46 ) ;
  assign n48 = ~n45 & n46 ;
  assign n49 = ( n34 & n47 ) | ( n34 & ~n48 ) | ( n47 & ~n48 ) ;
  assign n50 = n44 | n49 ;
  assign n51 = ( ~x22 & n34 ) | ( ~x22 & n41 ) | ( n34 & n41 ) ;
  assign n52 = ( x15 & ~x16 ) | ( x15 & x22 ) | ( ~x16 & x22 ) ;
  assign n53 = ( ~n35 & n40 ) | ( ~n35 & n52 ) | ( n40 & n52 ) ;
  assign n54 = ( ~x16 & n34 ) | ( ~x16 & n53 ) | ( n34 & n53 ) ;
  assign n55 = n51 & ~n54 ;
  assign n56 = ~x22 & n53 ;
  assign n57 = x16 | x22 ;
  assign n58 = ( n34 & n56 ) | ( n34 & ~n57 ) | ( n56 & ~n57 ) ;
  assign n59 = ( x16 & ~n55 ) | ( x16 & n58 ) | ( ~n55 & n58 ) ;
  assign n60 = n50 & n59 ;
  assign n61 = x16 | x17 ;
  assign n62 = x18 & ~x22 ;
  assign n63 = ( ~x22 & n61 ) | ( ~x22 & n62 ) | ( n61 & n62 ) ;
  assign n64 = x19 & ~n63 ;
  assign n65 = x19 & x22 ;
  assign n66 = ( ~n41 & n64 ) | ( ~n41 & n65 ) | ( n64 & n65 ) ;
  assign n67 = x19 & n65 ;
  assign n68 = ~n63 & n67 ;
  assign n69 = ( ~n34 & n66 ) | ( ~n34 & n68 ) | ( n66 & n68 ) ;
  assign n70 = ~x19 & n63 ;
  assign n71 = x19 | x22 ;
  assign n72 = ( n41 & n70 ) | ( n41 & ~n71 ) | ( n70 & ~n71 ) ;
  assign n73 = x19 & n71 ;
  assign n74 = ( ~n63 & n71 ) | ( ~n63 & n73 ) | ( n71 & n73 ) ;
  assign n75 = ( n34 & n72 ) | ( n34 & ~n74 ) | ( n72 & ~n74 ) ;
  assign n76 = n69 | n75 ;
  assign n77 = x18 & x22 ;
  assign n78 = x15 | n61 ;
  assign n79 = n40 | n78 ;
  assign n80 = x18 & n33 ;
  assign n81 = ( x18 & n30 ) | ( x18 & n80 ) | ( n30 & n80 ) ;
  assign n82 = ( x18 & n79 ) | ( x18 & n81 ) | ( n79 & n81 ) ;
  assign n83 = ( ~x22 & n41 ) | ( ~x22 & n63 ) | ( n41 & n63 ) ;
  assign n84 = ( ~x22 & n34 ) | ( ~x22 & n83 ) | ( n34 & n83 ) ;
  assign n85 = ~n82 & n84 ;
  assign n86 = n77 | n85 ;
  assign n87 = n76 | n86 ;
  assign n88 = n60 & ~n87 ;
  assign n89 = x18 | x19 ;
  assign n90 = n61 | n89 ;
  assign n91 = n33 | n90 ;
  assign n92 = n30 | n91 ;
  assign n93 = n41 & ~n92 ;
  assign n94 = ( x20 & ~n92 ) | ( x20 & n93 ) | ( ~n92 & n93 ) ;
  assign n95 = ( x20 & n93 ) | ( x20 & ~n94 ) | ( n93 & ~n94 ) ;
  assign n96 = x20 & x22 ;
  assign n97 = x22 & ~n96 ;
  assign n98 = ( n92 & n96 ) | ( n92 & ~n97 ) | ( n96 & ~n97 ) ;
  assign n99 = ( n92 & ~n96 ) | ( n92 & n97 ) | ( ~n96 & n97 ) ;
  assign n100 = ( x20 & n96 ) | ( x20 & ~n97 ) | ( n96 & ~n97 ) ;
  assign n101 = ( n93 & ~n99 ) | ( n93 & n100 ) | ( ~n99 & n100 ) ;
  assign n102 = ( ~n95 & n98 ) | ( ~n95 & n101 ) | ( n98 & n101 ) ;
  assign n103 = x21 & x22 ;
  assign n104 = x20 | x21 ;
  assign n105 = n90 | n104 ;
  assign n106 = n41 | n105 ;
  assign n107 = n34 | n106 ;
  assign n108 = x20 & x21 ;
  assign n109 = ( x21 & n90 ) | ( x21 & n108 ) | ( n90 & n108 ) ;
  assign n110 = ( x21 & n41 ) | ( x21 & n109 ) | ( n41 & n109 ) ;
  assign n111 = ( x21 & n34 ) | ( x21 & n110 ) | ( n34 & n110 ) ;
  assign n112 = n107 & ~n111 ;
  assign n113 = x22 & ~n103 ;
  assign n114 = ( n103 & n112 ) | ( n103 & ~n113 ) | ( n112 & ~n113 ) ;
  assign n115 = ( ~x22 & n33 ) | ( ~x22 & n40 ) | ( n33 & n40 ) ;
  assign n116 = x22 & ~n40 ;
  assign n117 = ( n30 & n115 ) | ( n30 & ~n116 ) | ( n115 & ~n116 ) ;
  assign n118 = ( ~x15 & x22 ) | ( ~x15 & n117 ) | ( x22 & n117 ) ;
  assign n119 = n117 & ~n118 ;
  assign n120 = x15 | x22 ;
  assign n121 = n117 & ~n120 ;
  assign n122 = ( x15 & ~n119 ) | ( x15 & n121 ) | ( ~n119 & n121 ) ;
  assign n123 = ~n114 & n122 ;
  assign n124 = ~n102 & n123 ;
  assign n125 = n88 & n124 ;
  assign n126 = ~n50 & n59 ;
  assign n127 = n76 & n86 ;
  assign n128 = n126 & n127 ;
  assign n129 = n114 | n122 ;
  assign n130 = n102 | n129 ;
  assign n131 = n128 & ~n130 ;
  assign n132 = n60 & n127 ;
  assign n133 = n102 & n123 ;
  assign n134 = n132 & n133 ;
  assign n135 = n131 | n134 ;
  assign n136 = n50 | n59 ;
  assign n137 = ~n76 & n86 ;
  assign n138 = ~n136 & n137 ;
  assign n139 = n124 & n138 ;
  assign n140 = n126 & n137 ;
  assign n141 = n124 & n140 ;
  assign n142 = n114 & ~n122 ;
  assign n143 = ~n102 & n142 ;
  assign n144 = n138 & n143 ;
  assign n145 = n141 | n144 ;
  assign n146 = n139 | n145 ;
  assign n147 = n135 | n146 ;
  assign n148 = n60 & n137 ;
  assign n149 = n102 & n142 ;
  assign n150 = n148 & n149 ;
  assign n151 = n76 & ~n86 ;
  assign n152 = ~n136 & n151 ;
  assign n153 = n114 & n122 ;
  assign n154 = n102 & n153 ;
  assign n155 = n152 & n154 ;
  assign n156 = n150 | n155 ;
  assign n157 = n50 & ~n59 ;
  assign n158 = n151 & n157 ;
  assign n159 = n143 & n158 ;
  assign n160 = n137 & n157 ;
  assign n161 = n143 & n160 ;
  assign n162 = n159 | n161 ;
  assign n163 = n156 | n162 ;
  assign n164 = n127 & ~n136 ;
  assign n165 = n143 & n164 ;
  assign n166 = n102 & ~n129 ;
  assign n167 = n140 & n166 ;
  assign n168 = n165 | n167 ;
  assign n169 = n163 | n168 ;
  assign n170 = n147 | n169 ;
  assign n171 = n127 & n157 ;
  assign n172 = n166 & n171 ;
  assign n173 = n133 & n152 ;
  assign n174 = n124 & n160 ;
  assign n175 = n173 | n174 ;
  assign n176 = n143 & n152 ;
  assign n177 = n88 & n149 ;
  assign n178 = n176 | n177 ;
  assign n179 = n175 | n178 ;
  assign n180 = n172 | n179 ;
  assign n181 = n170 | n180 ;
  assign n182 = n133 & n160 ;
  assign n183 = n138 & n154 ;
  assign n184 = n87 | n136 ;
  assign n185 = n154 & ~n184 ;
  assign n186 = n183 | n185 ;
  assign n187 = n182 | n186 ;
  assign n188 = ~n102 & n153 ;
  assign n189 = n128 & n188 ;
  assign n190 = ~n87 & n157 ;
  assign n191 = n188 & n190 ;
  assign n192 = ~n87 & n126 ;
  assign n193 = n143 & n192 ;
  assign n194 = n191 | n193 ;
  assign n195 = n189 | n194 ;
  assign n196 = n187 | n195 ;
  assign n197 = n148 & n154 ;
  assign n198 = n148 & n188 ;
  assign n199 = n197 | n198 ;
  assign n200 = n88 & n166 ;
  assign n201 = n60 & n151 ;
  assign n202 = n133 & n201 ;
  assign n203 = n200 | n202 ;
  assign n204 = n199 | n203 ;
  assign n205 = n124 & n132 ;
  assign n206 = ~n130 & n201 ;
  assign n207 = n205 | n206 ;
  assign n208 = n204 | n207 ;
  assign n209 = n196 | n208 ;
  assign n210 = ~n130 & n148 ;
  assign n211 = n126 & n151 ;
  assign n212 = ~n130 & n211 ;
  assign n213 = n210 | n212 ;
  assign n214 = n209 | n213 ;
  assign n215 = n181 | n214 ;
  assign n216 = n149 & n152 ;
  assign n217 = n133 & n192 ;
  assign n218 = n216 | n217 ;
  assign n219 = n166 & n211 ;
  assign n220 = n160 & n166 ;
  assign n221 = n219 | n220 ;
  assign n222 = n218 | n221 ;
  assign n223 = n124 & n171 ;
  assign n224 = ~n130 & n152 ;
  assign n225 = n223 | n224 ;
  assign n226 = n222 | n225 ;
  assign n227 = n133 & ~n184 ;
  assign n228 = n138 & n188 ;
  assign n229 = n140 & n188 ;
  assign n230 = n228 | n229 ;
  assign n231 = n227 | n230 ;
  assign n232 = n188 & n211 ;
  assign n233 = n188 & n201 ;
  assign n234 = n232 | n233 ;
  assign n235 = n158 & n166 ;
  assign n236 = n124 & n192 ;
  assign n237 = n235 | n236 ;
  assign n238 = n234 | n237 ;
  assign n239 = n231 | n238 ;
  assign n240 = n226 | n239 ;
  assign n241 = n149 & n211 ;
  assign n242 = n133 & n148 ;
  assign n243 = n241 | n242 ;
  assign n244 = n133 & n164 ;
  assign n245 = n133 & n190 ;
  assign n246 = n244 | n245 ;
  assign n247 = n243 | n246 ;
  assign n248 = n124 & n190 ;
  assign n249 = ~n130 & n171 ;
  assign n250 = n248 | n249 ;
  assign n251 = n247 | n250 ;
  assign n252 = n240 | n251 ;
  assign n253 = n149 & ~n184 ;
  assign n254 = n149 & n192 ;
  assign n255 = n253 | n254 ;
  assign n256 = n88 & n154 ;
  assign n257 = n138 & n166 ;
  assign n258 = n256 | n257 ;
  assign n259 = n255 | n258 ;
  assign n260 = ~n130 & n158 ;
  assign n261 = n128 & n166 ;
  assign n262 = ~n130 & n164 ;
  assign n263 = n261 | n262 ;
  assign n264 = n260 | n263 ;
  assign n265 = n259 | n264 ;
  assign n266 = n171 & n188 ;
  assign n267 = n143 & n171 ;
  assign n268 = n266 | n267 ;
  assign n269 = n138 & n149 ;
  assign n270 = n124 & ~n184 ;
  assign n271 = n269 | n270 ;
  assign n272 = n268 | n271 ;
  assign n273 = n265 | n272 ;
  assign n274 = n252 | n273 ;
  assign n275 = n215 | n274 ;
  assign n276 = n125 | n275 ;
  assign n277 = n124 & n148 ;
  assign n278 = n154 & n190 ;
  assign n279 = n183 | n278 ;
  assign n280 = n166 & ~n184 ;
  assign n281 = n223 | n280 ;
  assign n282 = n279 | n281 ;
  assign n283 = n154 & n201 ;
  assign n284 = n140 & n143 ;
  assign n285 = n161 | n284 ;
  assign n286 = n283 | n285 ;
  assign n287 = n282 | n286 ;
  assign n288 = n277 | n287 ;
  assign n289 = n149 & n201 ;
  assign n290 = n149 & n158 ;
  assign n291 = n289 | n290 ;
  assign n292 = n154 & n171 ;
  assign n293 = n154 & n192 ;
  assign n294 = n292 | n293 ;
  assign n295 = n291 | n294 ;
  assign n296 = n235 | n242 ;
  assign n297 = n269 | n296 ;
  assign n298 = n295 | n297 ;
  assign n299 = n149 & n171 ;
  assign n300 = n177 | n299 ;
  assign n301 = n148 & n166 ;
  assign n302 = n229 | n301 ;
  assign n303 = n300 | n302 ;
  assign n304 = n132 & n154 ;
  assign n305 = ~n130 & n140 ;
  assign n306 = n304 | n305 ;
  assign n307 = n303 | n306 ;
  assign n308 = n298 | n307 ;
  assign n309 = n288 | n308 ;
  assign n310 = n88 & ~n130 ;
  assign n311 = n188 & n192 ;
  assign n312 = n310 | n311 ;
  assign n313 = n141 | n191 ;
  assign n314 = n312 | n313 ;
  assign n315 = ~n130 & n192 ;
  assign n316 = n133 & n171 ;
  assign n317 = n167 | n316 ;
  assign n318 = n315 | n317 ;
  assign n319 = n314 | n318 ;
  assign n320 = n152 & n188 ;
  assign n321 = n128 & n149 ;
  assign n322 = n320 | n321 ;
  assign n323 = n244 | n260 ;
  assign n324 = n224 | n245 ;
  assign n325 = n323 | n324 ;
  assign n326 = n322 | n325 ;
  assign n327 = n319 | n326 ;
  assign n328 = n309 | n327 ;
  assign n329 = n261 | n267 ;
  assign n330 = n124 & n128 ;
  assign n331 = n125 | n330 ;
  assign n332 = n329 | n331 ;
  assign n333 = n133 & n138 ;
  assign n334 = n132 & n149 ;
  assign n335 = n333 | n334 ;
  assign n336 = n227 | n335 ;
  assign n337 = n332 | n336 ;
  assign n338 = n166 & n190 ;
  assign n339 = n124 & n201 ;
  assign n340 = n236 | n339 ;
  assign n341 = n338 | n340 ;
  assign n342 = n337 | n341 ;
  assign n343 = n128 & n154 ;
  assign n344 = n164 & n166 ;
  assign n345 = n343 | n344 ;
  assign n346 = n262 | n345 ;
  assign n347 = n149 & n164 ;
  assign n348 = n154 & n211 ;
  assign n349 = n347 | n348 ;
  assign n350 = n134 | n349 ;
  assign n351 = n346 | n350 ;
  assign n352 = n143 & n190 ;
  assign n353 = n154 & n158 ;
  assign n354 = n149 & n190 ;
  assign n355 = n353 | n354 ;
  assign n356 = n352 | n355 ;
  assign n357 = n164 & n188 ;
  assign n358 = n133 & n211 ;
  assign n359 = n357 | n358 ;
  assign n360 = n132 & n166 ;
  assign n361 = n124 & n211 ;
  assign n362 = n360 | n361 ;
  assign n363 = n359 | n362 ;
  assign n364 = n356 | n363 ;
  assign n365 = n351 | n364 ;
  assign n366 = n154 & n164 ;
  assign n367 = n232 | n366 ;
  assign n368 = n143 & n211 ;
  assign n369 = n189 | n368 ;
  assign n370 = n367 | n369 ;
  assign n371 = n159 | n256 ;
  assign n372 = n128 & n143 ;
  assign n373 = n266 | n372 ;
  assign n374 = n371 | n373 ;
  assign n375 = n200 | n249 ;
  assign n376 = n374 | n375 ;
  assign n377 = n370 | n376 ;
  assign n378 = n365 | n377 ;
  assign n379 = n342 | n378 ;
  assign n380 = n328 | n379 ;
  assign n381 = n276 | n380 ;
  assign n382 = n276 & ~n380 ;
  assign n383 = ( ~n276 & n381 ) | ( ~n276 & n382 ) | ( n381 & n382 ) ;
  assign n384 = n88 & n188 ;
  assign n385 = n134 | n384 ;
  assign n386 = n262 | n385 ;
  assign n387 = n154 & n160 ;
  assign n388 = n233 | n387 ;
  assign n389 = n216 | n228 ;
  assign n390 = n388 | n389 ;
  assign n391 = n386 | n390 ;
  assign n392 = n277 | n292 ;
  assign n393 = n291 | n392 ;
  assign n394 = n172 | n321 ;
  assign n395 = n317 | n394 ;
  assign n396 = n393 | n395 ;
  assign n397 = n149 & n160 ;
  assign n398 = n241 | n397 ;
  assign n399 = n150 | n197 ;
  assign n400 = n398 | n399 ;
  assign n401 = n396 | n400 ;
  assign n402 = n266 | n348 ;
  assign n403 = n155 | n174 ;
  assign n404 = n402 | n403 ;
  assign n405 = n257 | n404 ;
  assign n406 = n401 | n405 ;
  assign n407 = n124 & n158 ;
  assign n408 = n152 & n166 ;
  assign n409 = n219 | n408 ;
  assign n410 = n335 | n409 ;
  assign n411 = n407 | n410 ;
  assign n412 = n88 & n143 ;
  assign n413 = n165 | n412 ;
  assign n414 = n128 & n133 ;
  assign n415 = n284 | n414 ;
  assign n416 = n413 | n415 ;
  assign n417 = n173 | n360 ;
  assign n418 = n280 | n417 ;
  assign n419 = n310 | n357 ;
  assign n420 = n418 | n419 ;
  assign n421 = n416 | n420 ;
  assign n422 = n411 | n421 ;
  assign n423 = n406 | n422 ;
  assign n424 = n391 | n423 ;
  assign n425 = ~n130 & n132 ;
  assign n426 = ~n130 & n160 ;
  assign n427 = n248 | n426 ;
  assign n428 = n140 & n154 ;
  assign n429 = n140 & n149 ;
  assign n430 = n428 | n429 ;
  assign n431 = n427 | n430 ;
  assign n432 = n425 | n431 ;
  assign n433 = n189 | n372 ;
  assign n434 = n339 | n433 ;
  assign n435 = n88 & n133 ;
  assign n436 = n205 | n435 ;
  assign n437 = n125 | n436 ;
  assign n438 = n283 | n304 ;
  assign n439 = n353 | n438 ;
  assign n440 = n437 | n439 ;
  assign n441 = n434 | n440 ;
  assign n442 = n432 | n441 ;
  assign n443 = n158 & n188 ;
  assign n444 = n267 | n443 ;
  assign n445 = n224 | n229 ;
  assign n446 = n444 | n445 ;
  assign n447 = n210 | n235 ;
  assign n448 = n446 | n447 ;
  assign n449 = n144 | n347 ;
  assign n450 = n343 | n366 ;
  assign n451 = n449 | n450 ;
  assign n452 = n143 & n201 ;
  assign n453 = n227 | n452 ;
  assign n454 = n358 | n453 ;
  assign n455 = n451 | n454 ;
  assign n456 = ~n130 & n190 ;
  assign n457 = n161 | n456 ;
  assign n458 = n206 | n299 ;
  assign n459 = n457 | n458 ;
  assign n460 = n455 | n459 ;
  assign n461 = n448 | n460 ;
  assign n462 = n442 | n461 ;
  assign n463 = n424 | n462 ;
  assign n464 = n381 & ~n463 ;
  assign n465 = n383 & ~n464 ;
  assign n466 = ( ~x22 & n30 ) | ( ~x22 & n31 ) | ( n30 & n31 ) ;
  assign n467 = ( ~x9 & x22 ) | ( ~x9 & n31 ) | ( x22 & n31 ) ;
  assign n468 = ( ~x9 & n30 ) | ( ~x9 & n467 ) | ( n30 & n467 ) ;
  assign n469 = n466 & ~n468 ;
  assign n470 = x9 | x22 ;
  assign n471 = n31 & ~n470 ;
  assign n472 = ( n30 & ~n470 ) | ( n30 & n471 ) | ( ~n470 & n471 ) ;
  assign n473 = ( x9 & ~n469 ) | ( x9 & n472 ) | ( ~n469 & n472 ) ;
  assign n474 = n276 & n380 ;
  assign n475 = ( x7 & ~x22 ) | ( x7 & n30 ) | ( ~x22 & n30 ) ;
  assign n476 = ( x7 & x8 ) | ( x7 & x22 ) | ( x8 & x22 ) ;
  assign n477 = ( x8 & n30 ) | ( x8 & n476 ) | ( n30 & n476 ) ;
  assign n478 = n475 & ~n477 ;
  assign n479 = ~x22 & n476 ;
  assign n480 = x8 & ~x22 ;
  assign n481 = ( n30 & n479 ) | ( n30 & n480 ) | ( n479 & n480 ) ;
  assign n482 = ( x8 & n478 ) | ( x8 & ~n481 ) | ( n478 & ~n481 ) ;
  assign n483 = n463 | n482 ;
  assign n484 = ( ~n474 & n482 ) | ( ~n474 & n483 ) | ( n482 & n483 ) ;
  assign n485 = n383 | n484 ;
  assign n486 = n463 & n482 ;
  assign n487 = ( ~n381 & n482 ) | ( ~n381 & n486 ) | ( n482 & n486 ) ;
  assign n488 = ~n383 & n487 ;
  assign n489 = n485 & ~n488 ;
  assign n490 = ( n465 & n473 ) | ( n465 & ~n489 ) | ( n473 & ~n489 ) ;
  assign n491 = n463 & ~n474 ;
  assign n492 = n383 & ~n491 ;
  assign n493 = ( n473 & n489 ) | ( n473 & ~n492 ) | ( n489 & ~n492 ) ;
  assign n494 = ~n490 & n493 ;
  assign n495 = n166 & n192 ;
  assign n496 = n333 | n495 ;
  assign n497 = n228 | n388 ;
  assign n498 = n496 | n497 ;
  assign n499 = n183 | n292 ;
  assign n500 = n224 | n499 ;
  assign n501 = n166 & n201 ;
  assign n502 = n304 | n501 ;
  assign n503 = n223 | n502 ;
  assign n504 = n500 | n503 ;
  assign n505 = n498 | n504 ;
  assign n506 = n165 | n185 ;
  assign n507 = ( n144 & n443 ) | ( n144 & ~n506 ) | ( n443 & ~n506 ) ;
  assign n508 = n506 | n507 ;
  assign n509 = n130 | n184 ;
  assign n510 = ~n232 & n509 ;
  assign n511 = n124 & n164 ;
  assign n512 = n236 | n266 ;
  assign n513 = n511 | n512 ;
  assign n514 = n510 & ~n513 ;
  assign n515 = ~n508 & n514 ;
  assign n516 = ~n505 & n515 ;
  assign n517 = n176 | n197 ;
  assign n518 = n320 | n517 ;
  assign n519 = n235 | n310 ;
  assign n520 = n425 | n519 ;
  assign n521 = ( n353 & ~n518 ) | ( n353 & n520 ) | ( ~n518 & n520 ) ;
  assign n522 = n518 | n521 ;
  assign n523 = n219 | n343 ;
  assign n524 = n143 & n148 ;
  assign n525 = n241 | n524 ;
  assign n526 = n523 | n525 ;
  assign n527 = n437 | n526 ;
  assign n528 = n124 & n152 ;
  assign n529 = n352 | n528 ;
  assign n530 = n212 | n360 ;
  assign n531 = n529 | n530 ;
  assign n532 = n256 | n368 ;
  assign n533 = n167 | n532 ;
  assign n534 = n531 | n533 ;
  assign n535 = n527 | n534 ;
  assign n536 = n522 | n535 ;
  assign n537 = n516 & ~n536 ;
  assign n538 = n160 & n188 ;
  assign n539 = n278 | n299 ;
  assign n540 = n538 | n539 ;
  assign n541 = n198 | n428 ;
  assign n542 = n200 | n408 ;
  assign n543 = n541 | n542 ;
  assign n544 = n540 | n543 ;
  assign n545 = n132 & n143 ;
  assign n546 = n134 | n545 ;
  assign n547 = n544 | n546 ;
  assign n548 = ~n184 & n188 ;
  assign n549 = n261 | n548 ;
  assign n550 = n394 | n549 ;
  assign n551 = n210 | n248 ;
  assign n552 = n339 | n551 ;
  assign n553 = n550 | n552 ;
  assign n554 = n262 | n452 ;
  assign n555 = n159 | n254 ;
  assign n556 = n554 | n555 ;
  assign n557 = n182 | n344 ;
  assign n558 = n270 | n557 ;
  assign n559 = n556 | n558 ;
  assign n560 = n553 | n559 ;
  assign n561 = n547 | n560 ;
  assign n562 = n289 | n334 ;
  assign n563 = n242 | n357 ;
  assign n564 = n562 | n563 ;
  assign n565 = n217 | n277 ;
  assign n566 = n191 | n565 ;
  assign n567 = n564 | n566 ;
  assign n568 = n561 | n567 ;
  assign n569 = n537 & ~n568 ;
  assign n570 = n132 & n188 ;
  assign n571 = n315 | n570 ;
  assign n572 = n456 | n571 ;
  assign n573 = n569 & ~n572 ;
  assign n574 = n176 | n266 ;
  assign n575 = n260 | n574 ;
  assign n576 = n205 | n407 ;
  assign n577 = n321 | n576 ;
  assign n578 = n575 | n577 ;
  assign n579 = n524 | n548 ;
  assign n580 = n200 | n579 ;
  assign n581 = n578 | n580 ;
  assign n582 = n182 | n501 ;
  assign n583 = n228 | n452 ;
  assign n584 = n582 | n583 ;
  assign n585 = n210 | n224 ;
  assign n586 = n206 | n585 ;
  assign n587 = n584 | n586 ;
  assign n588 = n398 | n587 ;
  assign n589 = n581 | n588 ;
  assign n590 = n254 | n269 ;
  assign n591 = n155 | n304 ;
  assign n592 = n590 | n591 ;
  assign n593 = n372 | n592 ;
  assign n594 = n193 | n570 ;
  assign n595 = n299 | n347 ;
  assign n596 = n334 | n414 ;
  assign n597 = n595 | n596 ;
  assign n598 = n594 | n597 ;
  assign n599 = n593 | n598 ;
  assign n600 = n343 | n354 ;
  assign n601 = n531 | n600 ;
  assign n602 = n227 | n387 ;
  assign n603 = n329 | n602 ;
  assign n604 = n216 | n361 ;
  assign n605 = n366 | n604 ;
  assign n606 = n603 | n605 ;
  assign n607 = n601 | n606 ;
  assign n608 = n599 | n607 ;
  assign n609 = n589 | n608 ;
  assign n610 = n159 | n165 ;
  assign n611 = n435 | n610 ;
  assign n612 = n358 | n384 ;
  assign n613 = n202 | n292 ;
  assign n614 = n612 | n613 ;
  assign n615 = n611 | n614 ;
  assign n616 = n257 | n301 ;
  assign n617 = n615 | n616 ;
  assign n618 = n288 | n617 ;
  assign n619 = n219 | n368 ;
  assign n620 = n618 | n619 ;
  assign n621 = n609 | n620 ;
  assign n622 = n425 | n621 ;
  assign n623 = n573 & ~n622 ;
  assign n624 = n622 | n623 ;
  assign n625 = ( ~n573 & n623 ) | ( ~n573 & n624 ) | ( n623 & n624 ) ;
  assign n626 = ~n573 & n622 ;
  assign n627 = n276 & ~n626 ;
  assign n628 = n625 | n627 ;
  assign n629 = ( ~x22 & n30 ) | ( ~x22 & n33 ) | ( n30 & n33 ) ;
  assign n630 = ( ~x11 & x22 ) | ( ~x11 & n33 ) | ( x22 & n33 ) ;
  assign n631 = ( ~x11 & n30 ) | ( ~x11 & n630 ) | ( n30 & n630 ) ;
  assign n632 = n629 & ~n631 ;
  assign n633 = ~x22 & n631 ;
  assign n634 = ( x11 & ~n632 ) | ( x11 & n633 ) | ( ~n632 & n633 ) ;
  assign n635 = x10 & x22 ;
  assign n636 = x10 & ~n635 ;
  assign n637 = ( x9 & n31 ) | ( x9 & n636 ) | ( n31 & n636 ) ;
  assign n638 = n636 & n637 ;
  assign n639 = ( n30 & n636 ) | ( n30 & n638 ) | ( n636 & n638 ) ;
  assign n640 = ~x22 & n33 ;
  assign n641 = ( ~x22 & n30 ) | ( ~x22 & n640 ) | ( n30 & n640 ) ;
  assign n642 = ( n635 & ~n639 ) | ( n635 & n641 ) | ( ~n639 & n641 ) ;
  assign n643 = n276 | n642 ;
  assign n644 = ( ~n626 & n642 ) | ( ~n626 & n643 ) | ( n642 & n643 ) ;
  assign n645 = n625 & ~n644 ;
  assign n646 = n276 & n642 ;
  assign n647 = ( n623 & n642 ) | ( n623 & n646 ) | ( n642 & n646 ) ;
  assign n648 = n625 & n647 ;
  assign n649 = n645 | n648 ;
  assign n650 = ( n628 & n634 ) | ( n628 & ~n649 ) | ( n634 & ~n649 ) ;
  assign n651 = n276 | n623 ;
  assign n652 = ~n625 & n651 ;
  assign n653 = ( n634 & n649 ) | ( n634 & n652 ) | ( n649 & n652 ) ;
  assign n654 = n650 & ~n653 ;
  assign n655 = ~n494 & n654 ;
  assign n656 = n494 & ~n654 ;
  assign n657 = n655 | n656 ;
  assign n658 = ~x22 & n30 ;
  assign n659 = x7 & ~x22 ;
  assign n660 = n30 & n659 ;
  assign n661 = x7 & ~n659 ;
  assign n662 = ( x7 & ~n30 ) | ( x7 & n661 ) | ( ~n30 & n661 ) ;
  assign n663 = ( n658 & ~n660 ) | ( n658 & n662 ) | ( ~n660 & n662 ) ;
  assign n664 = n139 | n249 ;
  assign n665 = n398 | n664 ;
  assign n666 = n348 | n387 ;
  assign n667 = n227 | n666 ;
  assign n668 = n665 | n667 ;
  assign n669 = n173 | n220 ;
  assign n670 = n426 | n669 ;
  assign n671 = n668 | n670 ;
  assign n672 = n216 | n254 ;
  assign n673 = n408 | n672 ;
  assign n674 = n185 | n429 ;
  assign n675 = n197 | n358 ;
  assign n676 = n674 | n675 ;
  assign n677 = n412 | n511 ;
  assign n678 = n224 | n677 ;
  assign n679 = n676 | n678 ;
  assign n680 = n673 | n679 ;
  assign n681 = n671 | n680 ;
  assign n682 = n309 | n681 ;
  assign n683 = n321 | n594 ;
  assign n684 = n356 | n683 ;
  assign n685 = n205 | n428 ;
  assign n686 = n174 | n256 ;
  assign n687 = n685 | n686 ;
  assign n688 = n684 | n687 ;
  assign n689 = n143 & ~n184 ;
  assign n690 = n131 | n689 ;
  assign n691 = n156 | n330 ;
  assign n692 = n311 | n449 ;
  assign n693 = n691 | n692 ;
  assign n694 = n690 | n693 ;
  assign n695 = n688 | n694 ;
  assign n696 = n253 | n545 ;
  assign n697 = n523 | n696 ;
  assign n698 = n334 | n366 ;
  assign n699 = n191 | n698 ;
  assign n700 = n697 | n699 ;
  assign n701 = ~n130 & n138 ;
  assign n702 = n141 | n701 ;
  assign n703 = n228 | n548 ;
  assign n704 = n702 | n703 ;
  assign n705 = n182 | n704 ;
  assign n706 = n700 | n705 ;
  assign n707 = n695 | n706 ;
  assign n708 = n682 | n707 ;
  assign n709 = n133 & n140 ;
  assign n710 = n384 | n709 ;
  assign n711 = n210 | n425 ;
  assign n712 = n710 | n711 ;
  assign n713 = n708 | n712 ;
  assign n714 = n463 | n713 ;
  assign n715 = ~n713 & n714 ;
  assign n716 = ( ~n463 & n714 ) | ( ~n463 & n715 ) | ( n714 & n715 ) ;
  assign n717 = n193 | n412 ;
  assign n718 = n133 & n158 ;
  assign n719 = n134 | n718 ;
  assign n720 = n717 | n719 ;
  assign n721 = n172 | n720 ;
  assign n722 = n191 | n311 ;
  assign n723 = n352 | n384 ;
  assign n724 = n161 | n360 ;
  assign n725 = n723 | n724 ;
  assign n726 = n722 | n725 ;
  assign n727 = n721 | n726 ;
  assign n728 = n244 | n414 ;
  assign n729 = n261 | n728 ;
  assign n730 = n202 | n501 ;
  assign n731 = n316 | n730 ;
  assign n732 = n729 | n731 ;
  assign n733 = n689 | n732 ;
  assign n734 = n727 | n733 ;
  assign n735 = n344 | n548 ;
  assign n736 = n734 | n735 ;
  assign n737 = n330 | n511 ;
  assign n738 = n281 | n737 ;
  assign n739 = n231 | n738 ;
  assign n740 = n144 | n284 ;
  assign n741 = n249 | n425 ;
  assign n742 = n740 | n741 ;
  assign n743 = n739 | n742 ;
  assign n744 = n212 | n260 ;
  assign n745 = n361 | n744 ;
  assign n746 = n131 | n205 ;
  assign n747 = n206 | n262 ;
  assign n748 = n746 | n747 ;
  assign n749 = n407 | n528 ;
  assign n750 = n339 | n749 ;
  assign n751 = n748 | n750 ;
  assign n752 = n745 | n751 ;
  assign n753 = n743 | n752 ;
  assign n754 = n736 | n753 ;
  assign n755 = n714 & ~n754 ;
  assign n756 = n716 & ~n755 ;
  assign n757 = n463 & n713 ;
  assign n758 = ( ~x22 & n27 ) | ( ~x22 & n28 ) | ( n27 & n28 ) ;
  assign n759 = ( ~x6 & x22 ) | ( ~x6 & n28 ) | ( x22 & n28 ) ;
  assign n760 = ( ~x6 & n27 ) | ( ~x6 & n759 ) | ( n27 & n759 ) ;
  assign n761 = n758 & ~n760 ;
  assign n762 = ~x22 & n760 ;
  assign n763 = ( x6 & ~n761 ) | ( x6 & n762 ) | ( ~n761 & n762 ) ;
  assign n764 = n754 | n763 ;
  assign n765 = ( ~n757 & n763 ) | ( ~n757 & n764 ) | ( n763 & n764 ) ;
  assign n766 = n716 | n765 ;
  assign n767 = n754 & n763 ;
  assign n768 = ( ~n714 & n763 ) | ( ~n714 & n767 ) | ( n763 & n767 ) ;
  assign n769 = ~n716 & n768 ;
  assign n770 = n766 & ~n769 ;
  assign n771 = ( n663 & n756 ) | ( n663 & ~n770 ) | ( n756 & ~n770 ) ;
  assign n772 = n754 & ~n757 ;
  assign n773 = n716 & ~n772 ;
  assign n774 = ( n663 & n770 ) | ( n663 & ~n773 ) | ( n770 & ~n773 ) ;
  assign n775 = ~n771 & n774 ;
  assign n776 = n657 & n775 ;
  assign n777 = n657 & ~n776 ;
  assign n778 = ~n657 & n775 ;
  assign n779 = n777 | n778 ;
  assign n780 = n361 | n701 ;
  assign n781 = n320 | n397 ;
  assign n782 = n780 | n781 ;
  assign n783 = n279 | n782 ;
  assign n784 = n432 | n783 ;
  assign n785 = n510 & ~n784 ;
  assign n786 = n159 | n443 ;
  assign n787 = n223 | n333 ;
  assign n788 = n786 | n787 ;
  assign n789 = n718 | n730 ;
  assign n790 = n788 | n789 ;
  assign n791 = n343 | n528 ;
  assign n792 = n723 | n791 ;
  assign n793 = n242 | n506 ;
  assign n794 = n792 | n793 ;
  assign n795 = n270 | n338 ;
  assign n796 = n794 | n795 ;
  assign n797 = n790 | n796 ;
  assign n798 = n785 & ~n797 ;
  assign n799 = n449 | n557 ;
  assign n800 = n197 | n313 ;
  assign n801 = n799 | n800 ;
  assign n802 = n228 | n368 ;
  assign n803 = n173 | n244 ;
  assign n804 = n802 | n803 ;
  assign n805 = n339 | n804 ;
  assign n806 = n801 | n805 ;
  assign n807 = n798 & ~n806 ;
  assign n808 = n334 | n524 ;
  assign n809 = n134 | n407 ;
  assign n810 = n808 | n809 ;
  assign n811 = ( n317 & ~n593 ) | ( n317 & n810 ) | ( ~n593 & n810 ) ;
  assign n812 = n593 | n811 ;
  assign n813 = n245 | n266 ;
  assign n814 = n210 | n261 ;
  assign n815 = n813 | n814 ;
  assign n816 = n267 | n548 ;
  assign n817 = n456 | n816 ;
  assign n818 = n366 | n412 ;
  assign n819 = n131 | n219 ;
  assign n820 = n818 | n819 ;
  assign n821 = n817 | n820 ;
  assign n822 = n161 | n217 ;
  assign n823 = n495 | n822 ;
  assign n824 = n177 | n823 ;
  assign n825 = n821 | n824 ;
  assign n826 = n815 | n825 ;
  assign n827 = n812 | n826 ;
  assign n828 = n807 & ~n827 ;
  assign n829 = n294 | n416 ;
  assign n830 = n159 | n387 ;
  assign n831 = n200 | n830 ;
  assign n832 = n574 | n831 ;
  assign n833 = n829 | n832 ;
  assign n834 = n185 | n216 ;
  assign n835 = n690 | n834 ;
  assign n836 = n372 | n835 ;
  assign n837 = n833 | n836 ;
  assign n838 = ~n384 & n509 ;
  assign n839 = n227 | n548 ;
  assign n840 = n838 & ~n839 ;
  assign n841 = n219 | n280 ;
  assign n842 = n235 | n841 ;
  assign n843 = n840 & ~n842 ;
  assign n844 = n425 | n435 ;
  assign n845 = n277 | n511 ;
  assign n846 = n664 | n845 ;
  assign n847 = n844 | n846 ;
  assign n848 = n843 & ~n847 ;
  assign n849 = ~n837 & n848 ;
  assign n850 = n428 | n452 ;
  assign n851 = n312 | n850 ;
  assign n852 = n191 | n232 ;
  assign n853 = n134 | n852 ;
  assign n854 = n851 | n853 ;
  assign n855 = n210 | n360 ;
  assign n856 = n456 | n855 ;
  assign n857 = n854 | n856 ;
  assign n858 = n177 | n357 ;
  assign n859 = n291 | n858 ;
  assign n860 = n256 | n353 ;
  assign n861 = n189 | n860 ;
  assign n862 = n859 | n861 ;
  assign n863 = n347 | n862 ;
  assign n864 = n857 | n863 ;
  assign n865 = n333 | n429 ;
  assign n866 = n315 | n709 ;
  assign n867 = n865 | n866 ;
  assign n868 = x13 & x14 ;
  assign n869 = ( x14 & n38 ) | ( x14 & n868 ) | ( n38 & n868 ) ;
  assign n870 = ( x14 & n33 ) | ( x14 & n869 ) | ( n33 & n869 ) ;
  assign n871 = ( x14 & n30 ) | ( x14 & n870 ) | ( n30 & n870 ) ;
  assign n872 = n40 & ~n871 ;
  assign n873 = x14 & x22 ;
  assign n874 = x22 & ~n873 ;
  assign n875 = ( n871 & ~n873 ) | ( n871 & n874 ) | ( ~n873 & n874 ) ;
  assign n876 = ( n33 & n873 ) | ( n33 & ~n874 ) | ( n873 & ~n874 ) ;
  assign n877 = ~n873 & n874 ;
  assign n878 = ( n30 & n876 ) | ( n30 & ~n877 ) | ( n876 & ~n877 ) ;
  assign n879 = ( n872 & ~n875 ) | ( n872 & n878 ) | ( ~n875 & n878 ) ;
  assign n880 = ~n702 & n879 ;
  assign n881 = ~n867 & n880 ;
  assign n882 = ~n864 & n881 ;
  assign n883 = n849 & n882 ;
  assign n884 = n150 | n269 ;
  assign n885 = n368 | n387 ;
  assign n886 = n884 | n885 ;
  assign n887 = n518 | n886 ;
  assign n888 = n183 | n232 ;
  assign n889 = n887 | n888 ;
  assign n890 = n253 | n570 ;
  assign n891 = n165 | n372 ;
  assign n892 = n890 | n891 ;
  assign n893 = n862 | n892 ;
  assign n894 = n889 | n893 ;
  assign n895 = n254 | n321 ;
  assign n896 = n299 | n343 ;
  assign n897 = n895 | n896 ;
  assign n898 = n185 | n348 ;
  assign n899 = n897 | n898 ;
  assign n900 = n894 | n899 ;
  assign n901 = x0 & ~x22 ;
  assign n902 = ( ~x22 & n25 ) | ( ~x22 & n901 ) | ( n25 & n901 ) ;
  assign n903 = x3 & ~n902 ;
  assign n904 = ~x3 & n902 ;
  assign n905 = n903 | n904 ;
  assign n906 = n216 | n452 ;
  assign n907 = n524 | n538 ;
  assign n908 = n906 | n907 ;
  assign n909 = n398 | n541 ;
  assign n910 = n908 | n909 ;
  assign n911 = n155 | n429 ;
  assign n912 = n786 | n911 ;
  assign n913 = n233 | n912 ;
  assign n914 = n910 | n913 ;
  assign n915 = n283 | n347 ;
  assign n916 = n366 | n545 ;
  assign n917 = n915 | n916 ;
  assign n918 = n268 | n294 ;
  assign n919 = n917 | n918 ;
  assign n920 = n354 | n919 ;
  assign n921 = n914 | n920 ;
  assign n922 = n278 | n334 ;
  assign n923 = n304 & n905 ;
  assign n924 = ( n905 & n922 ) | ( n905 & n923 ) | ( n922 & n923 ) ;
  assign n925 = ( n905 & n921 ) | ( n905 & n924 ) | ( n921 & n924 ) ;
  assign n926 = ( n900 & n905 ) | ( n900 & n925 ) | ( n905 & n925 ) ;
  assign n927 = ~n883 & n926 ;
  assign n928 = ~n828 & n927 ;
  assign n929 = n883 & ~n926 ;
  assign n930 = ( n828 & ~n926 ) | ( n828 & n929 ) | ( ~n926 & n929 ) ;
  assign n931 = n928 | n930 ;
  assign n932 = x13 & x22 ;
  assign n933 = ( x13 & ~n38 ) | ( x13 & n932 ) | ( ~n38 & n932 ) ;
  assign n934 = ( ~n33 & n932 ) | ( ~n33 & n933 ) | ( n932 & n933 ) ;
  assign n935 = n932 & n933 ;
  assign n936 = ( ~n30 & n934 ) | ( ~n30 & n935 ) | ( n934 & n935 ) ;
  assign n937 = x13 | x22 ;
  assign n938 = n38 & ~n937 ;
  assign n939 = ( n33 & ~n937 ) | ( n33 & n938 ) | ( ~n937 & n938 ) ;
  assign n940 = n937 & ~n938 ;
  assign n941 = ( n30 & n939 ) | ( n30 & ~n940 ) | ( n939 & ~n940 ) ;
  assign n942 = n936 | n941 ;
  assign n943 = n434 | n575 ;
  assign n944 = n509 & ~n943 ;
  assign n945 = n554 | n696 ;
  assign n946 = n185 | n293 ;
  assign n947 = n161 | n946 ;
  assign n948 = n945 | n947 ;
  assign n949 = n210 | n368 ;
  assign n950 = n236 | n949 ;
  assign n951 = n948 | n950 ;
  assign n952 = n944 & ~n951 ;
  assign n953 = n233 | n320 ;
  assign n954 = n230 | n953 ;
  assign n955 = n270 | n315 ;
  assign n956 = n954 | n955 ;
  assign n957 = n952 & ~n956 ;
  assign n958 = n269 | n429 ;
  assign n959 = n172 | n344 ;
  assign n960 = n958 | n959 ;
  assign n961 = n135 | n960 ;
  assign n962 = n296 | n729 ;
  assign n963 = n961 | n962 ;
  assign n964 = n139 | n277 ;
  assign n965 = n257 | n338 ;
  assign n966 = n710 | n965 ;
  assign n967 = n280 | n301 ;
  assign n968 = n398 | n967 ;
  assign n969 = n966 | n968 ;
  assign n970 = n964 | n969 ;
  assign n971 = n963 | n970 ;
  assign n972 = n957 & ~n971 ;
  assign n973 = n256 | n289 ;
  assign n974 = n495 | n973 ;
  assign n975 = n500 | n691 ;
  assign n976 = n541 | n975 ;
  assign n977 = n790 | n976 ;
  assign n978 = n290 | n334 ;
  assign n979 = n358 | n689 ;
  assign n980 = n978 | n979 ;
  assign n981 = n200 | n305 ;
  assign n982 = n980 | n981 ;
  assign n983 = n722 | n780 ;
  assign n984 = n367 | n387 ;
  assign n985 = n983 | n984 ;
  assign n986 = n299 | n304 ;
  assign n987 = n985 | n986 ;
  assign n988 = n982 | n987 ;
  assign n989 = n977 | n988 ;
  assign n990 = n974 | n989 ;
  assign n991 = n972 & ~n990 ;
  assign n992 = n828 & n991 ;
  assign n993 = n573 & ~n992 ;
  assign n994 = n828 & ~n992 ;
  assign n995 = ( n991 & ~n992 ) | ( n991 & n994 ) | ( ~n992 & n994 ) ;
  assign n996 = ~n993 & n995 ;
  assign n997 = x12 & x22 ;
  assign n998 = n33 | n38 ;
  assign n999 = ( ~x22 & n658 ) | ( ~x22 & n998 ) | ( n658 & n998 ) ;
  assign n1000 = x11 | n33 ;
  assign n1001 = x12 & n30 ;
  assign n1002 = ( x12 & n1000 ) | ( x12 & n1001 ) | ( n1000 & n1001 ) ;
  assign n1003 = n999 & ~n1002 ;
  assign n1004 = n997 | n1003 ;
  assign n1005 = n828 | n991 ;
  assign n1006 = n573 & ~n1004 ;
  assign n1007 = ( n1004 & n1005 ) | ( n1004 & ~n1006 ) | ( n1005 & ~n1006 ) ;
  assign n1008 = n995 | n1007 ;
  assign n1009 = ~n573 & n1004 ;
  assign n1010 = ( n992 & n1004 ) | ( n992 & n1009 ) | ( n1004 & n1009 ) ;
  assign n1011 = ~n995 & n1010 ;
  assign n1012 = n1008 & ~n1011 ;
  assign n1013 = ( n942 & n996 ) | ( n942 & ~n1012 ) | ( n996 & ~n1012 ) ;
  assign n1014 = ~n573 & n1005 ;
  assign n1015 = n995 & ~n1014 ;
  assign n1016 = ( n942 & n1012 ) | ( n942 & ~n1015 ) | ( n1012 & ~n1015 ) ;
  assign n1017 = ~n1013 & n1016 ;
  assign n1018 = ~n931 & n1017 ;
  assign n1019 = n931 & ~n1017 ;
  assign n1020 = n1018 | n1019 ;
  assign n1021 = n301 | n709 ;
  assign n1022 = n220 | n1021 ;
  assign n1023 = n182 | n296 ;
  assign n1024 = n1022 | n1023 ;
  assign n1025 = n173 | n358 ;
  assign n1026 = n409 | n1025 ;
  assign n1027 = n735 | n1026 ;
  assign n1028 = n1024 | n1027 ;
  assign n1029 = n734 | n1028 ;
  assign n1030 = n217 | n338 ;
  assign n1031 = n496 | n1030 ;
  assign n1032 = n200 | n435 ;
  assign n1033 = n245 | n1032 ;
  assign n1034 = n1031 | n1033 ;
  assign n1035 = n230 | n740 ;
  assign n1036 = n257 | n1035 ;
  assign n1037 = n1034 | n1036 ;
  assign n1038 = n167 | n1037 ;
  assign n1039 = n1029 | n1038 ;
  assign n1040 = n754 | n1039 ;
  assign n1041 = ~n754 & n1040 ;
  assign n1042 = ( ~n1039 & n1040 ) | ( ~n1039 & n1041 ) | ( n1040 & n1041 ) ;
  assign n1043 = n304 | n922 ;
  assign n1044 = n921 | n1043 ;
  assign n1045 = n900 | n1044 ;
  assign n1046 = n905 & n1045 ;
  assign n1047 = ( n905 & ~n1040 ) | ( n905 & n1046 ) | ( ~n1040 & n1046 ) ;
  assign n1048 = n1042 & n1047 ;
  assign n1049 = n754 & n1039 ;
  assign n1050 = n905 | n1045 ;
  assign n1051 = ( n905 & ~n1049 ) | ( n905 & n1050 ) | ( ~n1049 & n1050 ) ;
  assign n1052 = n1045 & ~n1049 ;
  assign n1053 = n1051 & n1052 ;
  assign n1054 = ( n1042 & n1051 ) | ( n1042 & n1053 ) | ( n1051 & n1053 ) ;
  assign n1055 = ~n1048 & n1054 ;
  assign n1056 = n702 | n867 ;
  assign n1057 = n864 | n1056 ;
  assign n1058 = n849 & ~n1057 ;
  assign n1059 = n815 & ~n942 ;
  assign n1060 = ( n825 & ~n942 ) | ( n825 & n1059 ) | ( ~n942 & n1059 ) ;
  assign n1061 = ( n812 & ~n942 ) | ( n812 & n1060 ) | ( ~n942 & n1060 ) ;
  assign n1062 = ( n807 & n942 ) | ( n807 & ~n1061 ) | ( n942 & ~n1061 ) ;
  assign n1063 = n1058 & n1062 ;
  assign n1064 = n879 | n1058 ;
  assign n1065 = n828 & ~n1064 ;
  assign n1066 = n1063 | n1065 ;
  assign n1067 = n879 & ~n1058 ;
  assign n1068 = ~n828 & n1067 ;
  assign n1069 = n1052 & ~n1068 ;
  assign n1070 = ~n1066 & n1069 ;
  assign n1071 = n1055 & n1070 ;
  assign n1072 = n1052 & n1055 ;
  assign n1073 = ~n1052 & n1068 ;
  assign n1074 = ( ~n1055 & n1068 ) | ( ~n1055 & n1073 ) | ( n1068 & n1073 ) ;
  assign n1075 = ( n1066 & ~n1072 ) | ( n1066 & n1074 ) | ( ~n1072 & n1074 ) ;
  assign n1076 = n1071 | n1075 ;
  assign n1077 = n573 & ~n634 ;
  assign n1078 = ( n634 & n1005 ) | ( n634 & ~n1077 ) | ( n1005 & ~n1077 ) ;
  assign n1079 = n995 | n1078 ;
  assign n1080 = ~n573 & n634 ;
  assign n1081 = ( n634 & n992 ) | ( n634 & n1080 ) | ( n992 & n1080 ) ;
  assign n1082 = ~n995 & n1081 ;
  assign n1083 = n1079 & ~n1082 ;
  assign n1084 = ( n1004 & ~n1015 ) | ( n1004 & n1083 ) | ( ~n1015 & n1083 ) ;
  assign n1085 = ( n996 & n1004 ) | ( n996 & ~n1083 ) | ( n1004 & ~n1083 ) ;
  assign n1086 = n1084 & ~n1085 ;
  assign n1087 = n1040 & ~n1045 ;
  assign n1088 = n1042 & ~n1087 ;
  assign n1089 = ~x22 & n27 ;
  assign n1090 = x4 & ~x22 ;
  assign n1091 = n27 & n1090 ;
  assign n1092 = x4 & ~n1090 ;
  assign n1093 = ( x4 & ~n27 ) | ( x4 & n1092 ) | ( ~n27 & n1092 ) ;
  assign n1094 = ( n1089 & ~n1091 ) | ( n1089 & n1093 ) | ( ~n1091 & n1093 ) ;
  assign n1095 = n1042 | n1051 ;
  assign n1096 = ~n1042 & n1047 ;
  assign n1097 = n1095 & ~n1096 ;
  assign n1098 = ( n1088 & n1094 ) | ( n1088 & ~n1097 ) | ( n1094 & ~n1097 ) ;
  assign n1099 = n1042 & ~n1052 ;
  assign n1100 = ( n1094 & n1097 ) | ( n1094 & ~n1099 ) | ( n1097 & ~n1099 ) ;
  assign n1101 = ~n1098 & n1100 ;
  assign n1102 = ( ~n1076 & n1086 ) | ( ~n1076 & n1101 ) | ( n1086 & n1101 ) ;
  assign n1103 = ~n1020 & n1102 ;
  assign n1104 = n1020 & ~n1102 ;
  assign n1105 = n1103 | n1104 ;
  assign n1106 = n779 & ~n1105 ;
  assign n1107 = n779 & ~n1106 ;
  assign n1108 = n779 | n1105 ;
  assign n1109 = ~n1107 & n1108 ;
  assign n1110 = ( ~x22 & n27 ) | ( ~x22 & n1090 ) | ( n27 & n1090 ) ;
  assign n1111 = ~x5 & n1090 ;
  assign n1112 = x5 | x22 ;
  assign n1113 = ( n27 & n1111 ) | ( n27 & ~n1112 ) | ( n1111 & ~n1112 ) ;
  assign n1114 = x5 | n1113 ;
  assign n1115 = ( ~n1110 & n1113 ) | ( ~n1110 & n1114 ) | ( n1113 & n1114 ) ;
  assign n1116 = n1045 | n1094 ;
  assign n1117 = ( ~n1049 & n1094 ) | ( ~n1049 & n1116 ) | ( n1094 & n1116 ) ;
  assign n1118 = n1042 | n1117 ;
  assign n1119 = n1045 & n1094 ;
  assign n1120 = ( ~n1040 & n1094 ) | ( ~n1040 & n1119 ) | ( n1094 & n1119 ) ;
  assign n1121 = ~n1042 & n1120 ;
  assign n1122 = n1118 & ~n1121 ;
  assign n1123 = ( n1088 & n1115 ) | ( n1088 & ~n1122 ) | ( n1115 & ~n1122 ) ;
  assign n1124 = ( ~n1099 & n1115 ) | ( ~n1099 & n1122 ) | ( n1115 & n1122 ) ;
  assign n1125 = ~n1123 & n1124 ;
  assign n1126 = n1071 & n1125 ;
  assign n1127 = n1071 | n1125 ;
  assign n1128 = ~n1126 & n1127 ;
  assign n1129 = n463 | n663 ;
  assign n1130 = ( ~n474 & n663 ) | ( ~n474 & n1129 ) | ( n663 & n1129 ) ;
  assign n1131 = n383 | n1130 ;
  assign n1132 = n463 & n663 ;
  assign n1133 = ( ~n381 & n663 ) | ( ~n381 & n1132 ) | ( n663 & n1132 ) ;
  assign n1134 = ~n383 & n1133 ;
  assign n1135 = n1131 & ~n1134 ;
  assign n1136 = ( n482 & ~n492 ) | ( n482 & n1135 ) | ( ~n492 & n1135 ) ;
  assign n1137 = ( n465 & n482 ) | ( n465 & ~n1135 ) | ( n482 & ~n1135 ) ;
  assign n1138 = n1136 & ~n1137 ;
  assign n1139 = n754 | n1115 ;
  assign n1140 = ( ~n757 & n1115 ) | ( ~n757 & n1139 ) | ( n1115 & n1139 ) ;
  assign n1141 = n716 | n1140 ;
  assign n1142 = n754 & n1115 ;
  assign n1143 = ( ~n714 & n1115 ) | ( ~n714 & n1142 ) | ( n1115 & n1142 ) ;
  assign n1144 = ~n716 & n1143 ;
  assign n1145 = n1141 & ~n1144 ;
  assign n1146 = ( n763 & ~n773 ) | ( n763 & n1145 ) | ( ~n773 & n1145 ) ;
  assign n1147 = ( n756 & n763 ) | ( n756 & ~n1145 ) | ( n763 & ~n1145 ) ;
  assign n1148 = n1146 & ~n1147 ;
  assign n1149 = n276 | n473 ;
  assign n1150 = ( n473 & ~n626 ) | ( n473 & n1149 ) | ( ~n626 & n1149 ) ;
  assign n1151 = n625 & ~n1150 ;
  assign n1152 = n276 & n473 ;
  assign n1153 = ( n473 & n623 ) | ( n473 & n1152 ) | ( n623 & n1152 ) ;
  assign n1154 = n625 & n1153 ;
  assign n1155 = n1151 | n1154 ;
  assign n1156 = ( n628 & n642 ) | ( n628 & ~n1155 ) | ( n642 & ~n1155 ) ;
  assign n1157 = ( n642 & n652 ) | ( n642 & n1155 ) | ( n652 & n1155 ) ;
  assign n1158 = n1156 & ~n1157 ;
  assign n1159 = ( n1138 & n1148 ) | ( n1138 & n1158 ) | ( n1148 & n1158 ) ;
  assign n1160 = n1128 & n1159 ;
  assign n1161 = n1128 | n1159 ;
  assign n1162 = ~n1160 & n1161 ;
  assign n1163 = n754 & n905 ;
  assign n1164 = ( ~n714 & n905 ) | ( ~n714 & n1163 ) | ( n905 & n1163 ) ;
  assign n1165 = n716 & n1164 ;
  assign n1166 = n753 | n905 ;
  assign n1167 = n736 | n1166 ;
  assign n1168 = ( ~n757 & n905 ) | ( ~n757 & n1167 ) | ( n905 & n1167 ) ;
  assign n1169 = n772 & n1168 ;
  assign n1170 = ( n716 & n1168 ) | ( n716 & n1169 ) | ( n1168 & n1169 ) ;
  assign n1171 = ~n1165 & n1170 ;
  assign n1172 = ~n634 & n815 ;
  assign n1173 = ( ~n634 & n825 ) | ( ~n634 & n1172 ) | ( n825 & n1172 ) ;
  assign n1174 = ( ~n634 & n812 ) | ( ~n634 & n1173 ) | ( n812 & n1173 ) ;
  assign n1175 = ( n634 & n807 ) | ( n634 & ~n1174 ) | ( n807 & ~n1174 ) ;
  assign n1176 = n1058 & n1175 ;
  assign n1177 = ( n828 & n1004 ) | ( n828 & ~n1058 ) | ( n1004 & ~n1058 ) ;
  assign n1178 = ~n827 & n1004 ;
  assign n1179 = n807 & n1178 ;
  assign n1180 = ( n1176 & n1177 ) | ( n1176 & ~n1179 ) | ( n1177 & ~n1179 ) ;
  assign n1181 = n772 & ~n1180 ;
  assign n1182 = n1171 & n1181 ;
  assign n1183 = n276 | n482 ;
  assign n1184 = ( n482 & ~n626 ) | ( n482 & n1183 ) | ( ~n626 & n1183 ) ;
  assign n1185 = n625 & ~n1184 ;
  assign n1186 = n276 & n482 ;
  assign n1187 = ( n482 & n623 ) | ( n482 & n1186 ) | ( n623 & n1186 ) ;
  assign n1188 = n625 & n1187 ;
  assign n1189 = n1185 | n1188 ;
  assign n1190 = ( n473 & n628 ) | ( n473 & ~n1189 ) | ( n628 & ~n1189 ) ;
  assign n1191 = ( n473 & n652 ) | ( n473 & n1189 ) | ( n652 & n1189 ) ;
  assign n1192 = n1190 & ~n1191 ;
  assign n1193 = n463 | n763 ;
  assign n1194 = ( ~n474 & n763 ) | ( ~n474 & n1193 ) | ( n763 & n1193 ) ;
  assign n1195 = n383 | n1194 ;
  assign n1196 = n463 & n763 ;
  assign n1197 = ( ~n381 & n763 ) | ( ~n381 & n1196 ) | ( n763 & n1196 ) ;
  assign n1198 = ~n383 & n1197 ;
  assign n1199 = n1195 & ~n1198 ;
  assign n1200 = ( ~n492 & n663 ) | ( ~n492 & n1199 ) | ( n663 & n1199 ) ;
  assign n1201 = ( n465 & n663 ) | ( n465 & ~n1199 ) | ( n663 & ~n1199 ) ;
  assign n1202 = n1200 & ~n1201 ;
  assign n1203 = ( n1182 & n1192 ) | ( n1182 & n1202 ) | ( n1192 & n1202 ) ;
  assign n1204 = n815 & ~n1004 ;
  assign n1205 = ( n825 & ~n1004 ) | ( n825 & n1204 ) | ( ~n1004 & n1204 ) ;
  assign n1206 = ( n812 & ~n1004 ) | ( n812 & n1205 ) | ( ~n1004 & n1205 ) ;
  assign n1207 = ( n807 & n1004 ) | ( n807 & ~n1206 ) | ( n1004 & ~n1206 ) ;
  assign n1208 = n1058 & n1207 ;
  assign n1209 = ( n828 & n942 ) | ( n828 & ~n1058 ) | ( n942 & ~n1058 ) ;
  assign n1210 = ~n827 & n942 ;
  assign n1211 = n807 & n1210 ;
  assign n1212 = ( n1208 & n1209 ) | ( n1208 & ~n1211 ) | ( n1209 & ~n1211 ) ;
  assign n1213 = n573 & ~n642 ;
  assign n1214 = ( n642 & n1005 ) | ( n642 & ~n1213 ) | ( n1005 & ~n1213 ) ;
  assign n1215 = n995 | n1214 ;
  assign n1216 = ~n573 & n642 ;
  assign n1217 = ( n642 & n992 ) | ( n642 & n1216 ) | ( n992 & n1216 ) ;
  assign n1218 = ~n995 & n1217 ;
  assign n1219 = n1215 & ~n1218 ;
  assign n1220 = ( n634 & ~n1015 ) | ( n634 & n1219 ) | ( ~n1015 & n1219 ) ;
  assign n1221 = ( n634 & n996 ) | ( n634 & ~n1219 ) | ( n996 & ~n1219 ) ;
  assign n1222 = n1220 & ~n1221 ;
  assign n1223 = n754 | n1094 ;
  assign n1224 = ( ~n757 & n1094 ) | ( ~n757 & n1223 ) | ( n1094 & n1223 ) ;
  assign n1225 = n716 | n1224 ;
  assign n1226 = n754 & n1094 ;
  assign n1227 = ( ~n714 & n1094 ) | ( ~n714 & n1226 ) | ( n1094 & n1226 ) ;
  assign n1228 = ~n716 & n1227 ;
  assign n1229 = n1225 & ~n1228 ;
  assign n1230 = ( ~n773 & n1115 ) | ( ~n773 & n1229 ) | ( n1115 & n1229 ) ;
  assign n1231 = ( n756 & n1115 ) | ( n756 & ~n1229 ) | ( n1115 & ~n1229 ) ;
  assign n1232 = n1230 & ~n1231 ;
  assign n1233 = ( ~n1212 & n1222 ) | ( ~n1212 & n1232 ) | ( n1222 & n1232 ) ;
  assign n1234 = n1203 & n1233 ;
  assign n1235 = n1138 & ~n1148 ;
  assign n1236 = ~n1138 & n1148 ;
  assign n1237 = n1235 | n1236 ;
  assign n1238 = n1158 & n1237 ;
  assign n1239 = n1237 & ~n1238 ;
  assign n1240 = n1158 & ~n1237 ;
  assign n1241 = n1239 | n1240 ;
  assign n1242 = n1203 & ~n1234 ;
  assign n1243 = n1233 & ~n1234 ;
  assign n1244 = n1242 | n1243 ;
  assign n1245 = n1234 | n1244 ;
  assign n1246 = ( n1234 & n1241 ) | ( n1234 & n1245 ) | ( n1241 & n1245 ) ;
  assign n1247 = n1162 & n1246 ;
  assign n1248 = n1162 | n1246 ;
  assign n1249 = ~n1247 & n1248 ;
  assign n1250 = ~n1109 & n1249 ;
  assign n1251 = n1109 & ~n1249 ;
  assign n1252 = n1250 | n1251 ;
  assign n1253 = n1241 & ~n1244 ;
  assign n1254 = ~n1241 & n1244 ;
  assign n1255 = n1253 | n1254 ;
  assign n1256 = n1086 | n1101 ;
  assign n1257 = ~n1102 & n1256 ;
  assign n1258 = n1086 & n1101 ;
  assign n1259 = n1256 & ~n1258 ;
  assign n1260 = n1076 | n1259 ;
  assign n1261 = ~n1257 & n1260 ;
  assign n1262 = n1052 | n1055 ;
  assign n1263 = ~n1072 & n1262 ;
  assign n1264 = ~n473 & n573 ;
  assign n1265 = ( n473 & n1005 ) | ( n473 & ~n1264 ) | ( n1005 & ~n1264 ) ;
  assign n1266 = n995 | n1265 ;
  assign n1267 = n473 & ~n573 ;
  assign n1268 = ( n473 & n992 ) | ( n473 & n1267 ) | ( n992 & n1267 ) ;
  assign n1269 = ~n995 & n1268 ;
  assign n1270 = n1266 & ~n1269 ;
  assign n1271 = ( n642 & ~n1015 ) | ( n642 & n1270 ) | ( ~n1015 & n1270 ) ;
  assign n1272 = ( n642 & n996 ) | ( n642 & ~n1270 ) | ( n996 & ~n1270 ) ;
  assign n1273 = n1271 & ~n1272 ;
  assign n1274 = n463 | n1115 ;
  assign n1275 = ( ~n474 & n1115 ) | ( ~n474 & n1274 ) | ( n1115 & n1274 ) ;
  assign n1276 = n383 | n1275 ;
  assign n1277 = n463 & n1115 ;
  assign n1278 = ( ~n381 & n1115 ) | ( ~n381 & n1277 ) | ( n1115 & n1277 ) ;
  assign n1279 = ~n383 & n1278 ;
  assign n1280 = n1276 & ~n1279 ;
  assign n1281 = ( ~n492 & n763 ) | ( ~n492 & n1280 ) | ( n763 & n1280 ) ;
  assign n1282 = ( n465 & n763 ) | ( n465 & ~n1280 ) | ( n763 & ~n1280 ) ;
  assign n1283 = n1281 & ~n1282 ;
  assign n1284 = n276 | n663 ;
  assign n1285 = ( ~n626 & n663 ) | ( ~n626 & n1284 ) | ( n663 & n1284 ) ;
  assign n1286 = n625 & ~n1285 ;
  assign n1287 = n276 & n663 ;
  assign n1288 = ( n623 & n663 ) | ( n623 & n1287 ) | ( n663 & n1287 ) ;
  assign n1289 = n625 & n1288 ;
  assign n1290 = n1286 | n1289 ;
  assign n1291 = ( n482 & n628 ) | ( n482 & ~n1290 ) | ( n628 & ~n1290 ) ;
  assign n1292 = ( n482 & n652 ) | ( n482 & n1290 ) | ( n652 & n1290 ) ;
  assign n1293 = n1291 & ~n1292 ;
  assign n1294 = ( n1273 & n1283 ) | ( n1273 & n1293 ) | ( n1283 & n1293 ) ;
  assign n1295 = n1263 & n1294 ;
  assign n1296 = n1192 & ~n1202 ;
  assign n1297 = ~n1192 & n1202 ;
  assign n1298 = n1296 | n1297 ;
  assign n1299 = n1182 & n1298 ;
  assign n1300 = n1182 | n1298 ;
  assign n1301 = ~n1299 & n1300 ;
  assign n1302 = n1294 & ~n1295 ;
  assign n1303 = n1263 & ~n1294 ;
  assign n1304 = n1302 | n1303 ;
  assign n1305 = n1301 & n1304 ;
  assign n1306 = n1295 | n1305 ;
  assign n1307 = ( n1255 & ~n1261 ) | ( n1255 & n1306 ) | ( ~n1261 & n1306 ) ;
  assign n1308 = ~n1252 & n1307 ;
  assign n1309 = n1252 & ~n1307 ;
  assign n1310 = n1308 | n1309 ;
  assign n1311 = ~n1257 & n1295 ;
  assign n1312 = n1260 & n1311 ;
  assign n1313 = ( n1261 & n1305 ) | ( n1261 & n1312 ) | ( n1305 & n1312 ) ;
  assign n1314 = n1257 & ~n1295 ;
  assign n1315 = ( n1260 & n1295 ) | ( n1260 & ~n1314 ) | ( n1295 & ~n1314 ) ;
  assign n1316 = n1305 | n1315 ;
  assign n1317 = ~n1313 & n1316 ;
  assign n1318 = n1255 & n1317 ;
  assign n1669 = n1273 & ~n1283 ;
  assign n1670 = ~n1273 & n1283 ;
  assign n1671 = n1669 | n1670 ;
  assign n1672 = n1293 & n1671 ;
  assign n1673 = n1293 | n1671 ;
  assign n1674 = ~n1672 & n1673 ;
  assign n1319 = n463 | n1094 ;
  assign n1320 = ( ~n474 & n1094 ) | ( ~n474 & n1319 ) | ( n1094 & n1319 ) ;
  assign n1321 = n383 | n1320 ;
  assign n1322 = n463 & n1094 ;
  assign n1323 = ( ~n381 & n1094 ) | ( ~n381 & n1322 ) | ( n1094 & n1322 ) ;
  assign n1324 = ~n383 & n1323 ;
  assign n1325 = n1321 & ~n1324 ;
  assign n1326 = ( ~n492 & n1115 ) | ( ~n492 & n1325 ) | ( n1115 & n1325 ) ;
  assign n1327 = ( n465 & n1115 ) | ( n465 & ~n1325 ) | ( n1115 & ~n1325 ) ;
  assign n1328 = n1326 & ~n1327 ;
  assign n1329 = n462 | n905 ;
  assign n1330 = n424 | n1329 ;
  assign n1331 = ( ~n474 & n905 ) | ( ~n474 & n1330 ) | ( n905 & n1330 ) ;
  assign n1332 = n491 & n1331 ;
  assign n1333 = ( n383 & n1331 ) | ( n383 & n1332 ) | ( n1331 & n1332 ) ;
  assign n1334 = ~n473 & n815 ;
  assign n1335 = ( ~n473 & n825 ) | ( ~n473 & n1334 ) | ( n825 & n1334 ) ;
  assign n1336 = ( ~n473 & n812 ) | ( ~n473 & n1335 ) | ( n812 & n1335 ) ;
  assign n1337 = ( n473 & n807 ) | ( n473 & ~n1336 ) | ( n807 & ~n1336 ) ;
  assign n1338 = n1058 & n1337 ;
  assign n1339 = ( n642 & n828 ) | ( n642 & n1058 ) | ( n828 & n1058 ) ;
  assign n1340 = ~n642 & n827 ;
  assign n1341 = ( n642 & n807 ) | ( n642 & ~n1340 ) | ( n807 & ~n1340 ) ;
  assign n1342 = ( n1338 & ~n1339 ) | ( n1338 & n1341 ) | ( ~n1339 & n1341 ) ;
  assign n1343 = n491 & ~n1342 ;
  assign n1344 = n463 & n905 ;
  assign n1345 = ( ~n381 & n905 ) | ( ~n381 & n1344 ) | ( n905 & n1344 ) ;
  assign n1346 = n383 & n1345 ;
  assign n1347 = n1343 & ~n1346 ;
  assign n1348 = n1333 & n1347 ;
  assign n1352 = n714 & n905 ;
  assign n1353 = ~n462 & n905 ;
  assign n1354 = ~n424 & n1353 ;
  assign n1355 = ( n715 & n1352 ) | ( n715 & n1354 ) | ( n1352 & n1354 ) ;
  assign n1675 = ( n1328 & n1348 ) | ( n1328 & n1355 ) | ( n1348 & n1355 ) ;
  assign n1676 = n1674 & n1675 ;
  assign n1677 = n1674 | n1675 ;
  assign n1678 = ~n1676 & n1677 ;
  assign n1359 = n276 | n763 ;
  assign n1360 = ( ~n626 & n763 ) | ( ~n626 & n1359 ) | ( n763 & n1359 ) ;
  assign n1361 = n625 & ~n1360 ;
  assign n1362 = n276 & n763 ;
  assign n1363 = ( n623 & n763 ) | ( n623 & n1362 ) | ( n763 & n1362 ) ;
  assign n1364 = n625 & n1363 ;
  assign n1365 = n1361 | n1364 ;
  assign n1366 = ( n652 & n663 ) | ( n652 & n1365 ) | ( n663 & n1365 ) ;
  assign n1367 = ( n628 & n663 ) | ( n628 & ~n1365 ) | ( n663 & ~n1365 ) ;
  assign n1368 = ~n1366 & n1367 ;
  assign n1369 = ~n642 & n815 ;
  assign n1370 = ( ~n642 & n825 ) | ( ~n642 & n1369 ) | ( n825 & n1369 ) ;
  assign n1371 = ( ~n642 & n812 ) | ( ~n642 & n1370 ) | ( n812 & n1370 ) ;
  assign n1372 = ( n642 & n807 ) | ( n642 & ~n1371 ) | ( n807 & ~n1371 ) ;
  assign n1373 = n1058 & n1372 ;
  assign n1374 = ( n634 & n828 ) | ( n634 & ~n1058 ) | ( n828 & ~n1058 ) ;
  assign n1375 = n634 & ~n827 ;
  assign n1376 = n807 & n1375 ;
  assign n1377 = ( n1373 & n1374 ) | ( n1373 & ~n1376 ) | ( n1374 & ~n1376 ) ;
  assign n1378 = ~n482 & n573 ;
  assign n1379 = ( n482 & n1005 ) | ( n482 & ~n1378 ) | ( n1005 & ~n1378 ) ;
  assign n1380 = n995 | n1379 ;
  assign n1381 = n482 & ~n573 ;
  assign n1382 = ( n482 & n992 ) | ( n482 & n1381 ) | ( n992 & n1381 ) ;
  assign n1383 = ~n995 & n1382 ;
  assign n1384 = n1380 & ~n1383 ;
  assign n1385 = ( n473 & ~n1015 ) | ( n473 & n1384 ) | ( ~n1015 & n1384 ) ;
  assign n1386 = ( n473 & n996 ) | ( n473 & ~n1384 ) | ( n996 & ~n1384 ) ;
  assign n1387 = n1385 & ~n1386 ;
  assign n1679 = ( n1368 & ~n1377 ) | ( n1368 & n1387 ) | ( ~n1377 & n1387 ) ;
  assign n1680 = ~n772 & n1180 ;
  assign n1681 = ( ~n1171 & n1180 ) | ( ~n1171 & n1680 ) | ( n1180 & n1680 ) ;
  assign n1682 = n1182 | n1681 ;
  assign n1683 = n754 | n905 ;
  assign n1684 = ( ~n757 & n905 ) | ( ~n757 & n1683 ) | ( n905 & n1683 ) ;
  assign n1685 = n716 | n1684 ;
  assign n1686 = ~n716 & n1164 ;
  assign n1687 = n1685 & ~n1686 ;
  assign n1688 = ( ~n773 & n1094 ) | ( ~n773 & n1687 ) | ( n1094 & n1687 ) ;
  assign n1689 = ( n756 & n1094 ) | ( n756 & ~n1687 ) | ( n1094 & ~n1687 ) ;
  assign n1690 = n1688 & ~n1689 ;
  assign n1691 = n1682 & n1690 ;
  assign n1692 = n1682 | n1690 ;
  assign n1693 = ~n1691 & n1692 ;
  assign n1694 = ~n1679 & n1693 ;
  assign n1695 = n1679 & ~n1693 ;
  assign n1696 = n1694 | n1695 ;
  assign n1697 = ~n1676 & n1696 ;
  assign n1698 = ( n1676 & n1678 ) | ( n1676 & ~n1697 ) | ( n1678 & ~n1697 ) ;
  assign n1349 = ~n1328 & n1348 ;
  assign n1350 = n1328 & ~n1348 ;
  assign n1351 = n1349 | n1350 ;
  assign n1356 = n1351 & n1355 ;
  assign n1357 = n1351 | n1355 ;
  assign n1358 = ~n1356 & n1357 ;
  assign n1388 = n1377 | n1387 ;
  assign n1389 = n1377 & n1387 ;
  assign n1390 = n1388 & ~n1389 ;
  assign n1391 = n1368 & ~n1390 ;
  assign n1392 = ~n1368 & n1390 ;
  assign n1393 = n1391 | n1392 ;
  assign n1394 = n573 & ~n663 ;
  assign n1395 = ( n663 & n1005 ) | ( n663 & ~n1394 ) | ( n1005 & ~n1394 ) ;
  assign n1396 = n995 | n1395 ;
  assign n1397 = ~n573 & n663 ;
  assign n1398 = ( n663 & n992 ) | ( n663 & n1397 ) | ( n992 & n1397 ) ;
  assign n1399 = ~n995 & n1398 ;
  assign n1400 = n1396 & ~n1399 ;
  assign n1401 = ( n482 & ~n1015 ) | ( n482 & n1400 ) | ( ~n1015 & n1400 ) ;
  assign n1402 = ( n482 & n996 ) | ( n482 & ~n1400 ) | ( n996 & ~n1400 ) ;
  assign n1403 = n1401 & ~n1402 ;
  assign n1404 = n276 | n1115 ;
  assign n1405 = ( ~n626 & n1115 ) | ( ~n626 & n1404 ) | ( n1115 & n1404 ) ;
  assign n1406 = n625 & ~n1405 ;
  assign n1407 = n276 & n1115 ;
  assign n1408 = ( n623 & n1115 ) | ( n623 & n1407 ) | ( n1115 & n1407 ) ;
  assign n1409 = n625 & n1408 ;
  assign n1410 = n1406 | n1409 ;
  assign n1411 = ( n652 & n763 ) | ( n652 & n1410 ) | ( n763 & n1410 ) ;
  assign n1412 = ( n628 & n763 ) | ( n628 & ~n1410 ) | ( n763 & ~n1410 ) ;
  assign n1413 = ~n1411 & n1412 ;
  assign n1414 = n463 | n905 ;
  assign n1415 = ( ~n474 & n905 ) | ( ~n474 & n1414 ) | ( n905 & n1414 ) ;
  assign n1416 = n383 | n1415 ;
  assign n1417 = ~n383 & n1345 ;
  assign n1418 = n1416 & ~n1417 ;
  assign n1419 = ( ~n492 & n1094 ) | ( ~n492 & n1418 ) | ( n1094 & n1418 ) ;
  assign n1420 = ( n465 & n1094 ) | ( n465 & ~n1418 ) | ( n1094 & ~n1418 ) ;
  assign n1421 = n1419 & ~n1420 ;
  assign n1422 = ( n1403 & n1413 ) | ( n1403 & n1421 ) | ( n1413 & n1421 ) ;
  assign n1423 = ~n1393 & n1422 ;
  assign n1424 = n1393 | n1423 ;
  assign n1425 = n1358 & n1422 ;
  assign n1426 = n1393 & n1425 ;
  assign n1427 = ( n1358 & ~n1424 ) | ( n1358 & n1426 ) | ( ~n1424 & n1426 ) ;
  assign n1428 = n1358 | n1422 ;
  assign n1429 = ( n1358 & n1393 ) | ( n1358 & n1428 ) | ( n1393 & n1428 ) ;
  assign n1430 = n1424 & ~n1429 ;
  assign n1431 = n1427 | n1430 ;
  assign n1432 = ~n491 & n1342 ;
  assign n1433 = ( n1342 & n1346 ) | ( n1342 & n1432 ) | ( n1346 & n1432 ) ;
  assign n1434 = n1342 | n1432 ;
  assign n1435 = ( ~n1333 & n1433 ) | ( ~n1333 & n1434 ) | ( n1433 & n1434 ) ;
  assign n1436 = n1348 | n1435 ;
  assign n1437 = ~n482 & n815 ;
  assign n1438 = ( ~n482 & n825 ) | ( ~n482 & n1437 ) | ( n825 & n1437 ) ;
  assign n1439 = ( ~n482 & n812 ) | ( ~n482 & n1438 ) | ( n812 & n1438 ) ;
  assign n1440 = ( n482 & n807 ) | ( n482 & ~n1439 ) | ( n807 & ~n1439 ) ;
  assign n1441 = n1058 & n1440 ;
  assign n1442 = ( n473 & n828 ) | ( n473 & n1058 ) | ( n828 & n1058 ) ;
  assign n1443 = ~n473 & n827 ;
  assign n1444 = ( n473 & n807 ) | ( n473 & ~n1443 ) | ( n807 & ~n1443 ) ;
  assign n1445 = ( n1441 & ~n1442 ) | ( n1441 & n1444 ) | ( ~n1442 & n1444 ) ;
  assign n1446 = n573 & ~n763 ;
  assign n1447 = ( n763 & n1005 ) | ( n763 & ~n1446 ) | ( n1005 & ~n1446 ) ;
  assign n1448 = n995 | n1447 ;
  assign n1449 = ~n573 & n763 ;
  assign n1450 = ( n763 & n992 ) | ( n763 & n1449 ) | ( n992 & n1449 ) ;
  assign n1451 = ~n995 & n1450 ;
  assign n1452 = n1448 & ~n1451 ;
  assign n1453 = ( n663 & ~n1015 ) | ( n663 & n1452 ) | ( ~n1015 & n1452 ) ;
  assign n1454 = ( n663 & n996 ) | ( n663 & ~n1452 ) | ( n996 & ~n1452 ) ;
  assign n1455 = n1453 & ~n1454 ;
  assign n1456 = n276 | n1094 ;
  assign n1457 = ( ~n626 & n1094 ) | ( ~n626 & n1456 ) | ( n1094 & n1456 ) ;
  assign n1458 = n625 & ~n1457 ;
  assign n1459 = n276 & n1094 ;
  assign n1460 = ( n623 & n1094 ) | ( n623 & n1459 ) | ( n1094 & n1459 ) ;
  assign n1461 = n625 & n1460 ;
  assign n1462 = n1458 | n1461 ;
  assign n1463 = ( n652 & n1115 ) | ( n652 & n1462 ) | ( n1115 & n1462 ) ;
  assign n1464 = ( n628 & n1115 ) | ( n628 & ~n1462 ) | ( n1115 & ~n1462 ) ;
  assign n1465 = ~n1463 & n1464 ;
  assign n1466 = ( ~n1445 & n1455 ) | ( ~n1445 & n1465 ) | ( n1455 & n1465 ) ;
  assign n1467 = ~n1436 & n1466 ;
  assign n1468 = n1403 & ~n1413 ;
  assign n1469 = ~n1403 & n1413 ;
  assign n1470 = n1468 | n1469 ;
  assign n1471 = n1421 & n1470 ;
  assign n1472 = n1470 & ~n1471 ;
  assign n1473 = n1436 & ~n1466 ;
  assign n1474 = n1467 | n1473 ;
  assign n1475 = n1421 & ~n1470 ;
  assign n1476 = ~n1474 & n1475 ;
  assign n1477 = ( n1472 & ~n1474 ) | ( n1472 & n1476 ) | ( ~n1474 & n1476 ) ;
  assign n1478 = n1467 | n1477 ;
  assign n1479 = n276 & n905 ;
  assign n1480 = ( n623 & n905 ) | ( n623 & n1479 ) | ( n905 & n1479 ) ;
  assign n1481 = ~n625 & n1480 ;
  assign n1482 = n125 | n905 ;
  assign n1483 = n275 | n1482 ;
  assign n1484 = ( ~n626 & n905 ) | ( ~n626 & n1483 ) | ( n905 & n1483 ) ;
  assign n1485 = n627 & n1484 ;
  assign n1486 = ( ~n625 & n1484 ) | ( ~n625 & n1485 ) | ( n1484 & n1485 ) ;
  assign n1487 = ~n1481 & n1486 ;
  assign n1488 = ~n663 & n815 ;
  assign n1489 = ( ~n663 & n825 ) | ( ~n663 & n1488 ) | ( n825 & n1488 ) ;
  assign n1490 = ( ~n663 & n812 ) | ( ~n663 & n1489 ) | ( n812 & n1489 ) ;
  assign n1491 = ( n663 & n807 ) | ( n663 & ~n1490 ) | ( n807 & ~n1490 ) ;
  assign n1492 = n1058 & n1491 ;
  assign n1493 = ( n482 & n828 ) | ( n482 & n1058 ) | ( n828 & n1058 ) ;
  assign n1494 = ~n482 & n827 ;
  assign n1495 = ( n482 & n807 ) | ( n482 & ~n1494 ) | ( n807 & ~n1494 ) ;
  assign n1496 = ( n1492 & ~n1493 ) | ( n1492 & n1495 ) | ( ~n1493 & n1495 ) ;
  assign n1497 = n627 & ~n1496 ;
  assign n1498 = n1487 & n1497 ;
  assign n1499 = ~n627 & n1496 ;
  assign n1500 = ( ~n1487 & n1496 ) | ( ~n1487 & n1499 ) | ( n1496 & n1499 ) ;
  assign n1501 = n1498 | n1500 ;
  assign n1502 = n573 & ~n1115 ;
  assign n1503 = ( n1005 & n1115 ) | ( n1005 & ~n1502 ) | ( n1115 & ~n1502 ) ;
  assign n1504 = n995 | n1503 ;
  assign n1505 = ~n573 & n1115 ;
  assign n1506 = ( n992 & n1115 ) | ( n992 & n1505 ) | ( n1115 & n1505 ) ;
  assign n1507 = ~n995 & n1506 ;
  assign n1508 = n1504 & ~n1507 ;
  assign n1509 = ( n763 & ~n1015 ) | ( n763 & n1508 ) | ( ~n1015 & n1508 ) ;
  assign n1510 = ( n763 & n996 ) | ( n763 & ~n1508 ) | ( n996 & ~n1508 ) ;
  assign n1511 = n1509 & ~n1510 ;
  assign n1512 = n276 | n905 ;
  assign n1513 = ( ~n626 & n905 ) | ( ~n626 & n1512 ) | ( n905 & n1512 ) ;
  assign n1514 = n625 & ~n1513 ;
  assign n1515 = n625 & n1480 ;
  assign n1516 = n1514 | n1515 ;
  assign n1517 = ( n628 & n1094 ) | ( n628 & ~n1516 ) | ( n1094 & ~n1516 ) ;
  assign n1518 = ( n652 & n1094 ) | ( n652 & n1516 ) | ( n1094 & n1516 ) ;
  assign n1519 = n1517 & ~n1518 ;
  assign n1520 = ( ~n1501 & n1511 ) | ( ~n1501 & n1519 ) | ( n1511 & n1519 ) ;
  assign n1521 = n1333 & ~n1346 ;
  assign n1522 = ( n491 & n1498 ) | ( n491 & ~n1521 ) | ( n1498 & ~n1521 ) ;
  assign n1523 = ( ~n491 & n1498 ) | ( ~n491 & n1521 ) | ( n1498 & n1521 ) ;
  assign n1524 = ( ~n1498 & n1522 ) | ( ~n1498 & n1523 ) | ( n1522 & n1523 ) ;
  assign n1525 = n1520 & n1524 ;
  assign n1526 = ~n491 & n1346 ;
  assign n1527 = ( n491 & n1333 ) | ( n491 & ~n1526 ) | ( n1333 & ~n1526 ) ;
  assign n1528 = n491 & ~n1346 ;
  assign n1529 = n1333 & n1528 ;
  assign n1530 = n1527 & ~n1529 ;
  assign n1531 = n1498 & n1530 ;
  assign n1532 = n1525 | n1531 ;
  assign n1533 = n1524 & ~n1525 ;
  assign n1534 = n1520 & ~n1524 ;
  assign n1535 = n1533 | n1534 ;
  assign n1536 = n1511 | n1519 ;
  assign n1537 = ~n1520 & n1536 ;
  assign n1538 = n1511 & n1519 ;
  assign n1539 = n1536 & ~n1538 ;
  assign n1540 = n1501 | n1539 ;
  assign n1541 = ~n1537 & n1540 ;
  assign n1566 = n573 & ~n905 ;
  assign n1567 = ( n905 & n1005 ) | ( n905 & ~n1566 ) | ( n1005 & ~n1566 ) ;
  assign n1568 = n995 | n1567 ;
  assign n1542 = ~n573 & n905 ;
  assign n1543 = ( n905 & n992 ) | ( n905 & n1542 ) | ( n992 & n1542 ) ;
  assign n1544 = n995 & n1543 ;
  assign n1545 = n456 | n905 ;
  assign n1546 = n571 | n1545 ;
  assign n1547 = n569 & ~n1546 ;
  assign n1548 = ( n905 & n1005 ) | ( n905 & ~n1547 ) | ( n1005 & ~n1547 ) ;
  assign n1549 = n1014 & n1548 ;
  assign n1550 = ( n995 & n1548 ) | ( n995 & n1549 ) | ( n1548 & n1549 ) ;
  assign n1551 = ~n1544 & n1550 ;
  assign n1552 = n815 & ~n1115 ;
  assign n1553 = ( n825 & ~n1115 ) | ( n825 & n1552 ) | ( ~n1115 & n1552 ) ;
  assign n1554 = ( n812 & ~n1115 ) | ( n812 & n1553 ) | ( ~n1115 & n1553 ) ;
  assign n1555 = ( n807 & n1115 ) | ( n807 & ~n1554 ) | ( n1115 & ~n1554 ) ;
  assign n1556 = n1058 & n1555 ;
  assign n1557 = ( n763 & n828 ) | ( n763 & n1058 ) | ( n828 & n1058 ) ;
  assign n1558 = ~n763 & n827 ;
  assign n1559 = ( n763 & n807 ) | ( n763 & ~n1558 ) | ( n807 & ~n1558 ) ;
  assign n1560 = ( n1556 & ~n1557 ) | ( n1556 & n1559 ) | ( ~n1557 & n1559 ) ;
  assign n1561 = n1014 & ~n1560 ;
  assign n1562 = n1551 & n1561 ;
  assign n1563 = ~n1014 & n1560 ;
  assign n1564 = ( ~n1551 & n1560 ) | ( ~n1551 & n1563 ) | ( n1560 & n1563 ) ;
  assign n1565 = n1562 | n1564 ;
  assign n1569 = ~n1565 & n1568 ;
  assign n1570 = n1014 & n1551 ;
  assign n1571 = ( n1014 & n1551 ) | ( n1014 & ~n1570 ) | ( n1551 & ~n1570 ) ;
  assign n1572 = n702 & n1094 ;
  assign n1573 = ( n867 & n1094 ) | ( n867 & n1572 ) | ( n1094 & n1572 ) ;
  assign n1574 = ( n849 & n864 ) | ( n849 & n1573 ) | ( n864 & n1573 ) ;
  assign n1575 = ( ~n849 & n1094 ) | ( ~n849 & n1574 ) | ( n1094 & n1574 ) ;
  assign n1576 = n806 & ~n905 ;
  assign n1577 = ( n798 & n905 ) | ( n798 & ~n1576 ) | ( n905 & ~n1576 ) ;
  assign n1578 = ( ~n827 & n905 ) | ( ~n827 & n1577 ) | ( n905 & n1577 ) ;
  assign n1579 = n1575 | n1578 ;
  assign n1580 = n1058 | n1094 ;
  assign n1581 = ( n828 & n1094 ) | ( n828 & n1580 ) | ( n1094 & n1580 ) ;
  assign n1582 = ~n1575 & n1581 ;
  assign n1583 = ( n828 & n1058 ) | ( n828 & n1115 ) | ( n1058 & n1115 ) ;
  assign n1584 = n827 & ~n1115 ;
  assign n1585 = ( n807 & n1115 ) | ( n807 & ~n1584 ) | ( n1115 & ~n1584 ) ;
  assign n1586 = ( n1582 & ~n1583 ) | ( n1582 & n1585 ) | ( ~n1583 & n1585 ) ;
  assign n1587 = ( n1014 & n1579 ) | ( n1014 & n1586 ) | ( n1579 & n1586 ) ;
  assign n1588 = n1579 & n1586 ;
  assign n1589 = ( n1551 & n1587 ) | ( n1551 & n1588 ) | ( n1587 & n1588 ) ;
  assign n1590 = ~n1579 & n1583 ;
  assign n1591 = n1579 | n1585 ;
  assign n1592 = ( n1582 & ~n1590 ) | ( n1582 & n1591 ) | ( ~n1590 & n1591 ) ;
  assign n1593 = ( ~n1571 & n1589 ) | ( ~n1571 & n1592 ) | ( n1589 & n1592 ) ;
  assign n1594 = ( n1568 & n1569 ) | ( n1568 & ~n1593 ) | ( n1569 & ~n1593 ) ;
  assign n1595 = ~n995 & n1543 ;
  assign n1596 = ( n996 & n1094 ) | ( n996 & n1595 ) | ( n1094 & n1595 ) ;
  assign n1597 = ( n1015 & ~n1094 ) | ( n1015 & n1595 ) | ( ~n1094 & n1595 ) ;
  assign n1598 = n1596 | n1597 ;
  assign n1599 = n1594 & ~n1598 ;
  assign n1600 = ~n623 & n905 ;
  assign n1601 = ~n572 & n905 ;
  assign n1602 = n569 & n1601 ;
  assign n1603 = ( ~n624 & n1600 ) | ( ~n624 & n1602 ) | ( n1600 & n1602 ) ;
  assign n1604 = ~n1565 & n1603 ;
  assign n1605 = ~n1593 & n1604 ;
  assign n1606 = ( n1599 & n1603 ) | ( n1599 & n1605 ) | ( n1603 & n1605 ) ;
  assign n1607 = ~n1541 & n1606 ;
  assign n1608 = ~n763 & n815 ;
  assign n1609 = ( ~n763 & n825 ) | ( ~n763 & n1608 ) | ( n825 & n1608 ) ;
  assign n1610 = ( ~n763 & n812 ) | ( ~n763 & n1609 ) | ( n812 & n1609 ) ;
  assign n1611 = ( n763 & n807 ) | ( n763 & ~n1610 ) | ( n807 & ~n1610 ) ;
  assign n1612 = n1058 & n1611 ;
  assign n1613 = ( n663 & n828 ) | ( n663 & n1058 ) | ( n828 & n1058 ) ;
  assign n1614 = ~n663 & n827 ;
  assign n1615 = ( n663 & n807 ) | ( n663 & ~n1614 ) | ( n807 & ~n1614 ) ;
  assign n1616 = ( n1612 & ~n1613 ) | ( n1612 & n1615 ) | ( ~n1613 & n1615 ) ;
  assign n1617 = n573 & ~n1094 ;
  assign n1618 = ( n1005 & n1094 ) | ( n1005 & ~n1617 ) | ( n1094 & ~n1617 ) ;
  assign n1619 = n995 | n1618 ;
  assign n1620 = ~n573 & n1094 ;
  assign n1621 = ( n992 & n1094 ) | ( n992 & n1620 ) | ( n1094 & n1620 ) ;
  assign n1622 = ~n995 & n1621 ;
  assign n1623 = n1619 & ~n1622 ;
  assign n1624 = ( ~n1015 & n1115 ) | ( ~n1015 & n1623 ) | ( n1115 & n1623 ) ;
  assign n1625 = ( n996 & n1115 ) | ( n996 & ~n1623 ) | ( n1115 & ~n1623 ) ;
  assign n1626 = n1624 & ~n1625 ;
  assign n1627 = n1616 | n1626 ;
  assign n1628 = n1616 & n1626 ;
  assign n1629 = n1627 & ~n1628 ;
  assign n1630 = n1562 & n1629 ;
  assign n1631 = n1565 & ~n1603 ;
  assign n1632 = ( n1593 & ~n1603 ) | ( n1593 & n1631 ) | ( ~n1603 & n1631 ) ;
  assign n1633 = ~n1599 & n1632 ;
  assign n1634 = ( n1562 & n1629 ) | ( n1562 & ~n1630 ) | ( n1629 & ~n1630 ) ;
  assign n1635 = ( ~n1630 & n1633 ) | ( ~n1630 & n1634 ) | ( n1633 & n1634 ) ;
  assign n1636 = ( n1541 & ~n1607 ) | ( n1541 & n1635 ) | ( ~n1607 & n1635 ) ;
  assign n1637 = n1535 & ~n1636 ;
  assign n1638 = n1541 & ~n1606 ;
  assign n1639 = n1635 & n1638 ;
  assign n1640 = ( n1562 & ~n1616 ) | ( n1562 & n1626 ) | ( ~n1616 & n1626 ) ;
  assign n1641 = ~n1639 & n1640 ;
  assign n1642 = ( n1535 & n1637 ) | ( n1535 & n1641 ) | ( n1637 & n1641 ) ;
  assign n1643 = n1532 & n1642 ;
  assign n1644 = n1445 | n1455 ;
  assign n1645 = n1445 & n1455 ;
  assign n1646 = n1644 & ~n1645 ;
  assign n1647 = n1465 & n1646 ;
  assign n1648 = ~n1535 & n1636 ;
  assign n1649 = ~n1641 & n1648 ;
  assign n1650 = ( n1465 & n1646 ) | ( n1465 & ~n1647 ) | ( n1646 & ~n1647 ) ;
  assign n1651 = ( ~n1647 & n1649 ) | ( ~n1647 & n1650 ) | ( n1649 & n1650 ) ;
  assign n1652 = ( n1532 & n1643 ) | ( n1532 & ~n1651 ) | ( n1643 & ~n1651 ) ;
  assign n1653 = n1478 | n1652 ;
  assign n1654 = n1532 | n1642 ;
  assign n1655 = n1651 & ~n1654 ;
  assign n1656 = n1472 | n1475 ;
  assign n1657 = ~n1477 & n1656 ;
  assign n1658 = n1474 | n1477 ;
  assign n1659 = ( n1655 & ~n1657 ) | ( n1655 & n1658 ) | ( ~n1657 & n1658 ) ;
  assign n1660 = ~n1653 & n1659 ;
  assign n1661 = n1431 | n1660 ;
  assign n1664 = n1423 | n1426 ;
  assign n1665 = n1358 | n1423 ;
  assign n1666 = ( ~n1424 & n1664 ) | ( ~n1424 & n1665 ) | ( n1664 & n1665 ) ;
  assign n1662 = n1478 & n1652 ;
  assign n1663 = ( n1478 & ~n1659 ) | ( n1478 & n1662 ) | ( ~n1659 & n1662 ) ;
  assign n1667 = n1663 & n1666 ;
  assign n1668 = ( ~n1661 & n1666 ) | ( ~n1661 & n1667 ) | ( n1666 & n1667 ) ;
  assign n1699 = n1668 & n1698 ;
  assign n1700 = n1678 | n1696 ;
  assign n1701 = n1663 | n1666 ;
  assign n1702 = n1661 & ~n1701 ;
  assign n1703 = ( n1678 & n1696 ) | ( n1678 & ~n1700 ) | ( n1696 & ~n1700 ) ;
  assign n1704 = ( n1700 & n1702 ) | ( n1700 & ~n1703 ) | ( n1702 & ~n1703 ) ;
  assign n1705 = ( n1698 & n1699 ) | ( n1698 & ~n1704 ) | ( n1699 & ~n1704 ) ;
  assign n1706 = ( n1679 & ~n1682 ) | ( n1679 & n1690 ) | ( ~n1682 & n1690 ) ;
  assign n1707 = n1212 | n1222 ;
  assign n1708 = n1212 & n1222 ;
  assign n1709 = n1707 & ~n1708 ;
  assign n1710 = n1232 & ~n1709 ;
  assign n1711 = n1709 | n1710 ;
  assign n1712 = n1232 & n1709 ;
  assign n1713 = n1706 & n1712 ;
  assign n1714 = ( n1706 & ~n1711 ) | ( n1706 & n1713 ) | ( ~n1711 & n1713 ) ;
  assign n1715 = n1706 & ~n1714 ;
  assign n1716 = n1711 & ~n1712 ;
  assign n1717 = n1714 | n1716 ;
  assign n1718 = ~n1715 & n1717 ;
  assign n1719 = n1301 | n1304 ;
  assign n1720 = ~n1305 & n1719 ;
  assign n1721 = n1714 | n1720 ;
  assign n1722 = ( n1714 & ~n1718 ) | ( n1714 & n1721 ) | ( ~n1718 & n1721 ) ;
  assign n1723 = n1705 | n1722 ;
  assign n1724 = n1668 | n1698 ;
  assign n1725 = n1704 & ~n1724 ;
  assign n1726 = ~n1718 & n1720 ;
  assign n1727 = n1718 | n1726 ;
  assign n1728 = n1718 & n1720 ;
  assign n1729 = ( n1725 & n1727 ) | ( n1725 & ~n1728 ) | ( n1727 & ~n1728 ) ;
  assign n1730 = ~n1723 & n1729 ;
  assign n1731 = ( n1255 & n1317 ) | ( n1255 & ~n1318 ) | ( n1317 & ~n1318 ) ;
  assign n1732 = ( ~n1318 & n1730 ) | ( ~n1318 & n1731 ) | ( n1730 & n1731 ) ;
  assign n1733 = n1705 & n1722 ;
  assign n1734 = ( n1722 & ~n1729 ) | ( n1722 & n1733 ) | ( ~n1729 & n1733 ) ;
  assign n1735 = ~n1310 & n1734 ;
  assign n1736 = ( n1310 & n1732 ) | ( n1310 & ~n1735 ) | ( n1732 & ~n1735 ) ;
  assign n1737 = n276 | n1004 ;
  assign n1738 = ( ~n626 & n1004 ) | ( ~n626 & n1737 ) | ( n1004 & n1737 ) ;
  assign n1739 = n625 & ~n1738 ;
  assign n1740 = n276 & n1004 ;
  assign n1741 = ( n623 & n1004 ) | ( n623 & n1740 ) | ( n1004 & n1740 ) ;
  assign n1742 = n625 & n1741 ;
  assign n1743 = n1739 | n1742 ;
  assign n1744 = ( n628 & n942 ) | ( n628 & ~n1743 ) | ( n942 & ~n1743 ) ;
  assign n1745 = ( n652 & n942 ) | ( n652 & n1743 ) | ( n942 & n1743 ) ;
  assign n1746 = n1744 & ~n1745 ;
  assign n1747 = n463 | n642 ;
  assign n1748 = ( ~n474 & n642 ) | ( ~n474 & n1747 ) | ( n642 & n1747 ) ;
  assign n1749 = n383 | n1748 ;
  assign n1750 = n463 & n642 ;
  assign n1751 = ( ~n381 & n642 ) | ( ~n381 & n1750 ) | ( n642 & n1750 ) ;
  assign n1752 = ~n383 & n1751 ;
  assign n1753 = n1749 & ~n1752 ;
  assign n1754 = ( ~n492 & n634 ) | ( ~n492 & n1753 ) | ( n634 & n1753 ) ;
  assign n1755 = ( n465 & n634 ) | ( n465 & ~n1753 ) | ( n634 & ~n1753 ) ;
  assign n1756 = n1754 & ~n1755 ;
  assign n1757 = n1746 & ~n1756 ;
  assign n1758 = ~n1746 & n1756 ;
  assign n1759 = n1757 | n1758 ;
  assign n1760 = n482 | n754 ;
  assign n1761 = ( n482 & ~n757 ) | ( n482 & n1760 ) | ( ~n757 & n1760 ) ;
  assign n1762 = n716 | n1761 ;
  assign n1763 = n482 & n754 ;
  assign n1764 = ( n482 & ~n714 ) | ( n482 & n1763 ) | ( ~n714 & n1763 ) ;
  assign n1765 = ~n716 & n1764 ;
  assign n1766 = n1762 & ~n1765 ;
  assign n1767 = ( n473 & ~n773 ) | ( n473 & n1766 ) | ( ~n773 & n1766 ) ;
  assign n1768 = ( n473 & n756 ) | ( n473 & ~n1766 ) | ( n756 & ~n1766 ) ;
  assign n1769 = n1767 & ~n1768 ;
  assign n1770 = n1759 & n1769 ;
  assign n1771 = n1759 & ~n1770 ;
  assign n1772 = ~n573 & n879 ;
  assign n1773 = ( n879 & n992 ) | ( n879 & n1772 ) | ( n992 & n1772 ) ;
  assign n1774 = ~n995 & n1773 ;
  assign n1775 = n456 | n879 ;
  assign n1776 = n571 | n1775 ;
  assign n1777 = n569 & ~n1776 ;
  assign n1778 = ( n879 & n1005 ) | ( n879 & ~n1777 ) | ( n1005 & ~n1777 ) ;
  assign n1779 = n1014 & n1778 ;
  assign n1780 = ( ~n995 & n1778 ) | ( ~n995 & n1779 ) | ( n1778 & n1779 ) ;
  assign n1781 = ~n1774 & n1780 ;
  assign n1782 = n304 & n1115 ;
  assign n1783 = ( n922 & n1115 ) | ( n922 & n1782 ) | ( n1115 & n1782 ) ;
  assign n1784 = ( ~n900 & n921 ) | ( ~n900 & n1783 ) | ( n921 & n1783 ) ;
  assign n1785 = ( n900 & n1115 ) | ( n900 & n1784 ) | ( n1115 & n1784 ) ;
  assign n1786 = ~n828 & n1785 ;
  assign n1787 = n828 & ~n1785 ;
  assign n1788 = n1786 | n1787 ;
  assign n1789 = n1781 & ~n1788 ;
  assign n1790 = n1781 | n1788 ;
  assign n1791 = ( ~n1781 & n1789 ) | ( ~n1781 & n1790 ) | ( n1789 & n1790 ) ;
  assign n1792 = n1769 & ~n1791 ;
  assign n1793 = ~n1759 & n1792 ;
  assign n1794 = ( n1771 & ~n1791 ) | ( n1771 & n1793 ) | ( ~n1791 & n1793 ) ;
  assign n1795 = ~n1769 & n1791 ;
  assign n1796 = ( n1759 & n1791 ) | ( n1759 & n1795 ) | ( n1791 & n1795 ) ;
  assign n1797 = ~n1771 & n1796 ;
  assign n1798 = n1794 | n1797 ;
  assign n1806 = n573 | n828 ;
  assign n1807 = n1005 & ~n1806 ;
  assign n1799 = n573 & n828 ;
  assign n1800 = ( n828 & ~n1005 ) | ( n828 & n1799 ) | ( ~n1005 & n1799 ) ;
  assign n1801 = n304 & n763 ;
  assign n1802 = ( n763 & n922 ) | ( n763 & n1801 ) | ( n922 & n1801 ) ;
  assign n1803 = ( ~n900 & n921 ) | ( ~n900 & n1802 ) | ( n921 & n1802 ) ;
  assign n1804 = ( n763 & n900 ) | ( n763 & n1803 ) | ( n900 & n1803 ) ;
  assign n1805 = ~n1800 & n1804 ;
  assign n1808 = ~n1800 & n1807 ;
  assign n1809 = ( n1800 & n1805 ) | ( n1800 & ~n1808 ) | ( n1805 & ~n1808 ) ;
  assign n1810 = n1807 | n1809 ;
  assign n1811 = n1804 & n1807 ;
  assign n1812 = ( n1804 & ~n1805 ) | ( n1804 & n1811 ) | ( ~n1805 & n1811 ) ;
  assign n1813 = n1810 & ~n1812 ;
  assign n1814 = n463 | n634 ;
  assign n1815 = ( ~n474 & n634 ) | ( ~n474 & n1814 ) | ( n634 & n1814 ) ;
  assign n1816 = n383 | n1815 ;
  assign n1817 = n463 & n634 ;
  assign n1818 = ( ~n381 & n634 ) | ( ~n381 & n1817 ) | ( n634 & n1817 ) ;
  assign n1819 = ~n383 & n1818 ;
  assign n1820 = n1816 & ~n1819 ;
  assign n1821 = ( ~n492 & n1004 ) | ( ~n492 & n1820 ) | ( n1004 & n1820 ) ;
  assign n1822 = ( n465 & n1004 ) | ( n465 & ~n1820 ) | ( n1004 & ~n1820 ) ;
  assign n1823 = n1821 & ~n1822 ;
  assign n1824 = ~n1813 & n1823 ;
  assign n1825 = n1813 & ~n1823 ;
  assign n1826 = n1824 | n1825 ;
  assign n1827 = ~n1786 & n1788 ;
  assign n1828 = ( n1781 & n1786 ) | ( n1781 & ~n1827 ) | ( n1786 & ~n1827 ) ;
  assign n1829 = ~n1826 & n1828 ;
  assign n1830 = n1826 & ~n1828 ;
  assign n1831 = n1829 | n1830 ;
  assign n1832 = n1045 | n1115 ;
  assign n1833 = ( ~n1049 & n1115 ) | ( ~n1049 & n1832 ) | ( n1115 & n1832 ) ;
  assign n1834 = n1042 | n1833 ;
  assign n1835 = n1045 & n1115 ;
  assign n1836 = ( ~n1040 & n1115 ) | ( ~n1040 & n1835 ) | ( n1115 & n1835 ) ;
  assign n1837 = ~n1042 & n1836 ;
  assign n1838 = n1834 & ~n1837 ;
  assign n1839 = ( n763 & ~n1099 ) | ( n763 & n1838 ) | ( ~n1099 & n1838 ) ;
  assign n1840 = ( n763 & n1088 ) | ( n763 & ~n1838 ) | ( n1088 & ~n1838 ) ;
  assign n1841 = n1839 & ~n1840 ;
  assign n1842 = ( n928 & ~n931 ) | ( n928 & n1841 ) | ( ~n931 & n1841 ) ;
  assign n1843 = n928 & n1841 ;
  assign n1844 = ( n1017 & n1842 ) | ( n1017 & n1843 ) | ( n1842 & n1843 ) ;
  assign n1845 = ~n928 & n931 ;
  assign n1846 = ~n1841 & n1845 ;
  assign n1847 = n928 | n1841 ;
  assign n1848 = ( n1017 & ~n1846 ) | ( n1017 & n1847 ) | ( ~n1846 & n1847 ) ;
  assign n1849 = ~n1844 & n1848 ;
  assign n1850 = ( n494 & n654 ) | ( n494 & n775 ) | ( n654 & n775 ) ;
  assign n1851 = n1844 | n1850 ;
  assign n1852 = ( n1844 & n1849 ) | ( n1844 & n1851 ) | ( n1849 & n1851 ) ;
  assign n1853 = ~n1793 & n1852 ;
  assign n1854 = n1791 & n1852 ;
  assign n1855 = ( ~n1771 & n1853 ) | ( ~n1771 & n1854 ) | ( n1853 & n1854 ) ;
  assign n1856 = ( n1794 & ~n1831 ) | ( n1794 & n1855 ) | ( ~n1831 & n1855 ) ;
  assign n1857 = n1794 & ~n1831 ;
  assign n1858 = ( ~n1798 & n1856 ) | ( ~n1798 & n1857 ) | ( n1856 & n1857 ) ;
  assign n1859 = ~n1793 & n1831 ;
  assign n1860 = n1791 & n1831 ;
  assign n1861 = ( ~n1771 & n1859 ) | ( ~n1771 & n1860 ) | ( n1859 & n1860 ) ;
  assign n1862 = ~n1852 & n1861 ;
  assign n1863 = ( n1798 & n1861 ) | ( n1798 & n1862 ) | ( n1861 & n1862 ) ;
  assign n1864 = n1858 | n1863 ;
  assign n1865 = n276 | n942 ;
  assign n1866 = ( ~n626 & n942 ) | ( ~n626 & n1865 ) | ( n942 & n1865 ) ;
  assign n1867 = n625 & ~n1866 ;
  assign n1868 = n276 & n942 ;
  assign n1869 = ( n623 & n942 ) | ( n623 & n1868 ) | ( n942 & n1868 ) ;
  assign n1870 = n625 & n1869 ;
  assign n1871 = n1867 | n1870 ;
  assign n1872 = ( n628 & n879 ) | ( n628 & ~n1871 ) | ( n879 & ~n1871 ) ;
  assign n1873 = ( n652 & n879 ) | ( n652 & n1871 ) | ( n879 & n1871 ) ;
  assign n1874 = n1872 & ~n1873 ;
  assign n1875 = n473 | n754 ;
  assign n1876 = ( n473 & ~n757 ) | ( n473 & n1875 ) | ( ~n757 & n1875 ) ;
  assign n1877 = n716 | n1876 ;
  assign n1878 = n473 & n754 ;
  assign n1879 = ( n473 & ~n714 ) | ( n473 & n1878 ) | ( ~n714 & n1878 ) ;
  assign n1880 = ~n716 & n1879 ;
  assign n1881 = n1877 & ~n1880 ;
  assign n1882 = ( n642 & ~n773 ) | ( n642 & n1881 ) | ( ~n773 & n1881 ) ;
  assign n1883 = ( n642 & n756 ) | ( n642 & ~n1881 ) | ( n756 & ~n1881 ) ;
  assign n1884 = n1882 & ~n1883 ;
  assign n1885 = n663 | n1045 ;
  assign n1886 = ( n663 & ~n1049 ) | ( n663 & n1885 ) | ( ~n1049 & n1885 ) ;
  assign n1887 = n1042 | n1886 ;
  assign n1888 = n663 & n1045 ;
  assign n1889 = ( n663 & ~n1040 ) | ( n663 & n1888 ) | ( ~n1040 & n1888 ) ;
  assign n1890 = ~n1042 & n1889 ;
  assign n1891 = n1887 & ~n1890 ;
  assign n1892 = ( n482 & ~n1099 ) | ( n482 & n1891 ) | ( ~n1099 & n1891 ) ;
  assign n1893 = ( n482 & n1088 ) | ( n482 & ~n1891 ) | ( n1088 & ~n1891 ) ;
  assign n1894 = n1892 & ~n1893 ;
  assign n1895 = n1884 & ~n1894 ;
  assign n1896 = ~n1884 & n1894 ;
  assign n1897 = n1895 | n1896 ;
  assign n1898 = n1874 & n1897 ;
  assign n1899 = n1874 | n1897 ;
  assign n1900 = ~n1898 & n1899 ;
  assign n1901 = ( n1746 & n1756 ) | ( n1746 & n1769 ) | ( n1756 & n1769 ) ;
  assign n1902 = n1900 | n1901 ;
  assign n1903 = n1900 & n1901 ;
  assign n1904 = n1902 & ~n1903 ;
  assign n1905 = n573 & ~n942 ;
  assign n1906 = ( n942 & n1005 ) | ( n942 & ~n1905 ) | ( n1005 & ~n1905 ) ;
  assign n1907 = n995 | n1906 ;
  assign n1908 = ~n573 & n942 ;
  assign n1909 = ( n942 & n992 ) | ( n942 & n1908 ) | ( n992 & n1908 ) ;
  assign n1910 = ~n995 & n1909 ;
  assign n1911 = n1907 & ~n1910 ;
  assign n1912 = ( n879 & ~n1015 ) | ( n879 & n1911 ) | ( ~n1015 & n1911 ) ;
  assign n1913 = ( n879 & n996 ) | ( n879 & ~n1911 ) | ( n996 & ~n1911 ) ;
  assign n1914 = n1912 & ~n1913 ;
  assign n1915 = n763 | n1045 ;
  assign n1916 = ( n763 & ~n1049 ) | ( n763 & n1915 ) | ( ~n1049 & n1915 ) ;
  assign n1917 = n1042 | n1916 ;
  assign n1918 = n763 & n1045 ;
  assign n1919 = ( n763 & ~n1040 ) | ( n763 & n1918 ) | ( ~n1040 & n1918 ) ;
  assign n1920 = ~n1042 & n1919 ;
  assign n1921 = n1917 & ~n1920 ;
  assign n1922 = ( n663 & ~n1099 ) | ( n663 & n1921 ) | ( ~n1099 & n1921 ) ;
  assign n1923 = ( n663 & n1088 ) | ( n663 & ~n1921 ) | ( n1088 & ~n1921 ) ;
  assign n1924 = n1922 & ~n1923 ;
  assign n1925 = n304 & n1094 ;
  assign n1926 = ( n922 & n1094 ) | ( n922 & n1925 ) | ( n1094 & n1925 ) ;
  assign n1927 = ( ~n900 & n921 ) | ( ~n900 & n1926 ) | ( n921 & n1926 ) ;
  assign n1928 = ( n900 & n1094 ) | ( n900 & n1927 ) | ( n1094 & n1927 ) ;
  assign n1929 = ~n828 & n1928 ;
  assign n1930 = n828 & ~n1928 ;
  assign n1931 = n1929 | n1930 ;
  assign n1932 = ~n1929 & n1931 ;
  assign n1933 = n1924 & ~n1932 ;
  assign n1934 = n1924 & n1929 ;
  assign n1935 = ( n1914 & n1933 ) | ( n1914 & n1934 ) | ( n1933 & n1934 ) ;
  assign n1936 = ~n1924 & n1932 ;
  assign n1937 = n1924 | n1929 ;
  assign n1938 = ( n1914 & ~n1936 ) | ( n1914 & n1937 ) | ( ~n1936 & n1937 ) ;
  assign n1939 = ~n1935 & n1938 ;
  assign n1940 = n463 | n473 ;
  assign n1941 = ( n473 & ~n474 ) | ( n473 & n1940 ) | ( ~n474 & n1940 ) ;
  assign n1942 = n383 | n1941 ;
  assign n1943 = n463 & n473 ;
  assign n1944 = ( ~n381 & n473 ) | ( ~n381 & n1943 ) | ( n473 & n1943 ) ;
  assign n1945 = ~n383 & n1944 ;
  assign n1946 = n1942 & ~n1945 ;
  assign n1947 = ( ~n492 & n642 ) | ( ~n492 & n1946 ) | ( n642 & n1946 ) ;
  assign n1948 = ( n465 & n642 ) | ( n465 & ~n1946 ) | ( n642 & ~n1946 ) ;
  assign n1949 = n1947 & ~n1948 ;
  assign n1950 = n276 | n634 ;
  assign n1951 = ( ~n626 & n634 ) | ( ~n626 & n1950 ) | ( n634 & n1950 ) ;
  assign n1952 = n625 & ~n1951 ;
  assign n1953 = n276 & n634 ;
  assign n1954 = ( n623 & n634 ) | ( n623 & n1953 ) | ( n634 & n1953 ) ;
  assign n1955 = n625 & n1954 ;
  assign n1956 = n1952 | n1955 ;
  assign n1957 = ( n628 & n1004 ) | ( n628 & ~n1956 ) | ( n1004 & ~n1956 ) ;
  assign n1958 = ( n652 & n1004 ) | ( n652 & n1956 ) | ( n1004 & n1956 ) ;
  assign n1959 = n1957 & ~n1958 ;
  assign n1960 = n663 | n754 ;
  assign n1961 = ( n663 & ~n757 ) | ( n663 & n1960 ) | ( ~n757 & n1960 ) ;
  assign n1962 = n716 | n1961 ;
  assign n1963 = n663 & n754 ;
  assign n1964 = ( n663 & ~n714 ) | ( n663 & n1963 ) | ( ~n714 & n1963 ) ;
  assign n1965 = ~n716 & n1964 ;
  assign n1966 = n1962 & ~n1965 ;
  assign n1967 = ( n482 & ~n773 ) | ( n482 & n1966 ) | ( ~n773 & n1966 ) ;
  assign n1968 = ( n482 & n756 ) | ( n482 & ~n1966 ) | ( n756 & ~n1966 ) ;
  assign n1969 = n1967 & ~n1968 ;
  assign n1970 = ( n1949 & n1959 ) | ( n1949 & n1969 ) | ( n1959 & n1969 ) ;
  assign n1971 = n1935 | n1970 ;
  assign n1972 = ( n1935 & n1939 ) | ( n1935 & n1971 ) | ( n1939 & n1971 ) ;
  assign n1973 = n1904 & n1972 ;
  assign n1974 = n1904 | n1972 ;
  assign n1975 = ~n1973 & n1974 ;
  assign n1976 = ~n1864 & n1975 ;
  assign n1977 = n1864 & ~n1975 ;
  assign n1978 = n1976 | n1977 ;
  assign n1979 = n1798 & n1852 ;
  assign n1980 = n1798 | n1852 ;
  assign n1981 = ~n1979 & n1980 ;
  assign n1982 = n1939 & n1970 ;
  assign n1983 = n1939 | n1970 ;
  assign n1984 = ~n1982 & n1983 ;
  assign n1985 = ~n1949 & n1959 ;
  assign n1986 = n1949 & ~n1959 ;
  assign n1987 = n1985 | n1986 ;
  assign n1988 = n1969 & n1987 ;
  assign n1989 = n1987 & ~n1988 ;
  assign n1990 = n1914 | n1931 ;
  assign n1991 = n1914 & n1931 ;
  assign n1992 = n1990 & ~n1991 ;
  assign n1993 = n1969 & ~n1987 ;
  assign n1994 = n1126 | n1160 ;
  assign n1995 = ( ~n1992 & n1993 ) | ( ~n1992 & n1994 ) | ( n1993 & n1994 ) ;
  assign n1996 = n1992 & ~n1994 ;
  assign n1997 = ( n1989 & n1995 ) | ( n1989 & ~n1996 ) | ( n1995 & ~n1996 ) ;
  assign n1998 = n1984 & n1997 ;
  assign n1999 = n1984 | n1997 ;
  assign n2000 = ~n1998 & n1999 ;
  assign n2001 = n1998 | n2000 ;
  assign n2002 = ( ~n1981 & n1998 ) | ( ~n1981 & n2001 ) | ( n1998 & n2001 ) ;
  assign n2003 = ~n1978 & n2002 ;
  assign n2004 = n1978 & ~n2002 ;
  assign n2005 = n2003 | n2004 ;
  assign n2006 = ~n1981 & n2000 ;
  assign n2007 = n1981 & ~n2000 ;
  assign n2008 = n2006 | n2007 ;
  assign n2009 = n1849 & n1850 ;
  assign n2010 = n1849 | n1850 ;
  assign n2011 = ~n2009 & n2010 ;
  assign n2014 = ( n1103 & ~n1105 ) | ( n1103 & n2011 ) | ( ~n1105 & n2011 ) ;
  assign n2015 = n1103 & n2011 ;
  assign n2016 = ( n779 & n2014 ) | ( n779 & n2015 ) | ( n2014 & n2015 ) ;
  assign n2012 = n1103 | n2011 ;
  assign n2013 = n1106 | n2012 ;
  assign n2017 = n2013 & ~n2016 ;
  assign n2018 = n1989 | n1993 ;
  assign n2019 = n1992 | n1994 ;
  assign n2020 = n1992 & n1994 ;
  assign n2021 = n2019 & ~n2020 ;
  assign n2022 = n2018 & ~n2021 ;
  assign n2023 = ~n2018 & n2021 ;
  assign n2024 = n2022 | n2023 ;
  assign n2025 = ~n2016 & n2024 ;
  assign n2026 = ( n2016 & n2017 ) | ( n2016 & ~n2025 ) | ( n2017 & ~n2025 ) ;
  assign n2027 = ~n2008 & n2026 ;
  assign n2028 = n2008 & ~n2026 ;
  assign n2029 = n2027 | n2028 ;
  assign n2030 = n2017 & ~n2024 ;
  assign n2031 = ~n2017 & n2024 ;
  assign n2032 = n2030 | n2031 ;
  assign n2033 = n1247 | n1250 ;
  assign n2034 = ~n2032 & n2033 ;
  assign n2035 = n2032 & ~n2033 ;
  assign n2036 = n2034 | n2035 ;
  assign n2037 = ~n2034 & n2036 ;
  assign n2038 = n2029 | n2037 ;
  assign n2039 = ~n2005 & n2027 ;
  assign n2040 = ( n2005 & n2038 ) | ( n2005 & ~n2039 ) | ( n2038 & ~n2039 ) ;
  assign n2041 = n276 & n879 ;
  assign n2042 = ( n623 & n879 ) | ( n623 & n2041 ) | ( n879 & n2041 ) ;
  assign n2043 = n625 & n2042 ;
  assign n2044 = n125 | n879 ;
  assign n2045 = n275 | n2044 ;
  assign n2046 = ( ~n626 & n879 ) | ( ~n626 & n2045 ) | ( n879 & n2045 ) ;
  assign n2047 = n627 & n2046 ;
  assign n2048 = ( n625 & n2046 ) | ( n625 & n2047 ) | ( n2046 & n2047 ) ;
  assign n2049 = ~n2043 & n2048 ;
  assign n2050 = n304 & n663 ;
  assign n2051 = ( n663 & n922 ) | ( n663 & n2050 ) | ( n922 & n2050 ) ;
  assign n2052 = ( ~n900 & n921 ) | ( ~n900 & n2051 ) | ( n921 & n2051 ) ;
  assign n2053 = ( n663 & n900 ) | ( n663 & n2052 ) | ( n900 & n2052 ) ;
  assign n2054 = n2049 & ~n2053 ;
  assign n2055 = ~n2049 & n2053 ;
  assign n2056 = n2054 | n2055 ;
  assign n2057 = n463 | n1004 ;
  assign n2058 = ( ~n474 & n1004 ) | ( ~n474 & n2057 ) | ( n1004 & n2057 ) ;
  assign n2059 = n383 | n2058 ;
  assign n2060 = n463 & n1004 ;
  assign n2061 = ( ~n381 & n1004 ) | ( ~n381 & n2060 ) | ( n1004 & n2060 ) ;
  assign n2062 = ~n383 & n2061 ;
  assign n2063 = n2059 & ~n2062 ;
  assign n2064 = ( ~n492 & n942 ) | ( ~n492 & n2063 ) | ( n942 & n2063 ) ;
  assign n2065 = ( n465 & n942 ) | ( n465 & ~n2063 ) | ( n942 & ~n2063 ) ;
  assign n2066 = n2064 & ~n2065 ;
  assign n2067 = ~n2056 & n2066 ;
  assign n2068 = n2056 & ~n2066 ;
  assign n2069 = n2067 | n2068 ;
  assign n2070 = ( n1874 & n1884 ) | ( n1874 & n1894 ) | ( n1884 & n1894 ) ;
  assign n2071 = ~n2069 & n2070 ;
  assign n2072 = n2069 | n2071 ;
  assign n2073 = n2069 & n2070 ;
  assign n2074 = n2072 & ~n2073 ;
  assign n2075 = n642 | n754 ;
  assign n2076 = ( n642 & ~n757 ) | ( n642 & n2075 ) | ( ~n757 & n2075 ) ;
  assign n2077 = n716 | n2076 ;
  assign n2078 = n642 & n754 ;
  assign n2079 = ( n642 & ~n714 ) | ( n642 & n2078 ) | ( ~n714 & n2078 ) ;
  assign n2080 = ~n716 & n2079 ;
  assign n2081 = n2077 & ~n2080 ;
  assign n2082 = ( n634 & ~n773 ) | ( n634 & n2081 ) | ( ~n773 & n2081 ) ;
  assign n2083 = ( n634 & n756 ) | ( n634 & ~n2081 ) | ( n756 & ~n2081 ) ;
  assign n2084 = n2082 & ~n2083 ;
  assign n2085 = n482 | n1045 ;
  assign n2086 = ( n482 & ~n1049 ) | ( n482 & n2085 ) | ( ~n1049 & n2085 ) ;
  assign n2087 = n1042 | n2086 ;
  assign n2088 = n482 & n1045 ;
  assign n2089 = ( n482 & ~n1040 ) | ( n482 & n2088 ) | ( ~n1040 & n2088 ) ;
  assign n2090 = ~n1042 & n2089 ;
  assign n2091 = n2087 & ~n2090 ;
  assign n2092 = ( n473 & ~n1099 ) | ( n473 & n2091 ) | ( ~n1099 & n2091 ) ;
  assign n2093 = ( n473 & n1088 ) | ( n473 & ~n2091 ) | ( n1088 & ~n2091 ) ;
  assign n2094 = n2092 & ~n2093 ;
  assign n2095 = n2084 & n2094 ;
  assign n2096 = n2084 | n2094 ;
  assign n2097 = ~n2095 & n2096 ;
  assign n2098 = n1809 & n2097 ;
  assign n2099 = n1809 | n2097 ;
  assign n2100 = ~n2098 & n2099 ;
  assign n2101 = n2071 | n2100 ;
  assign n2102 = ( n2071 & ~n2074 ) | ( n2071 & n2101 ) | ( ~n2074 & n2101 ) ;
  assign n2103 = n463 | n942 ;
  assign n2104 = ( ~n474 & n942 ) | ( ~n474 & n2103 ) | ( n942 & n2103 ) ;
  assign n2105 = n383 | n2104 ;
  assign n2106 = n463 & n942 ;
  assign n2107 = ( ~n381 & n942 ) | ( ~n381 & n2106 ) | ( n942 & n2106 ) ;
  assign n2108 = ~n383 & n2107 ;
  assign n2109 = n2105 & ~n2108 ;
  assign n2110 = ( ~n492 & n879 ) | ( ~n492 & n2109 ) | ( n879 & n2109 ) ;
  assign n2111 = ( n465 & n879 ) | ( n465 & ~n2109 ) | ( n879 & ~n2109 ) ;
  assign n2112 = n2110 & ~n2111 ;
  assign n2113 = n634 | n754 ;
  assign n2114 = ( n634 & ~n757 ) | ( n634 & n2113 ) | ( ~n757 & n2113 ) ;
  assign n2115 = n716 | n2114 ;
  assign n2116 = n634 & n754 ;
  assign n2117 = ( n634 & ~n714 ) | ( n634 & n2116 ) | ( ~n714 & n2116 ) ;
  assign n2118 = ~n716 & n2117 ;
  assign n2119 = n2115 & ~n2118 ;
  assign n2120 = ( ~n773 & n1004 ) | ( ~n773 & n2119 ) | ( n1004 & n2119 ) ;
  assign n2121 = ( n756 & n1004 ) | ( n756 & ~n2119 ) | ( n1004 & ~n2119 ) ;
  assign n2122 = n2120 & ~n2121 ;
  assign n2123 = n2112 & ~n2122 ;
  assign n2124 = ~n2112 & n2122 ;
  assign n2125 = n2123 | n2124 ;
  assign n2126 = n473 | n1045 ;
  assign n2127 = ( n473 & ~n1049 ) | ( n473 & n2126 ) | ( ~n1049 & n2126 ) ;
  assign n2128 = n1042 | n2127 ;
  assign n2129 = n473 & n1045 ;
  assign n2130 = ( n473 & ~n1040 ) | ( n473 & n2129 ) | ( ~n1040 & n2129 ) ;
  assign n2131 = ~n1042 & n2130 ;
  assign n2132 = n2128 & ~n2131 ;
  assign n2133 = ( n642 & ~n1099 ) | ( n642 & n2132 ) | ( ~n1099 & n2132 ) ;
  assign n2134 = ( n642 & n1088 ) | ( n642 & ~n2132 ) | ( n1088 & ~n2132 ) ;
  assign n2135 = n2133 & ~n2134 ;
  assign n2136 = n2125 & n2135 ;
  assign n2137 = n2125 & ~n2136 ;
  assign n2138 = ~n2125 & n2135 ;
  assign n2139 = n2137 | n2138 ;
  assign n2140 = n2102 & n2139 ;
  assign n2141 = n2102 | n2139 ;
  assign n2142 = ~n2140 & n2141 ;
  assign n2143 = n276 & ~n2053 ;
  assign n2144 = ~n626 & n2143 ;
  assign n2145 = ~n276 & n2053 ;
  assign n2146 = ( n626 & n2053 ) | ( n626 & n2145 ) | ( n2053 & n2145 ) ;
  assign n2147 = n2144 | n2146 ;
  assign n2148 = n2088 & n2147 ;
  assign n2149 = n2088 | n2147 ;
  assign n2150 = ~n2148 & n2149 ;
  assign n2151 = ( n1809 & n2084 ) | ( n1809 & n2094 ) | ( n2084 & n2094 ) ;
  assign n2152 = n2054 | n2066 ;
  assign n2153 = ( n2054 & ~n2056 ) | ( n2054 & n2152 ) | ( ~n2056 & n2152 ) ;
  assign n2154 = ( n2150 & n2151 ) | ( n2150 & ~n2153 ) | ( n2151 & ~n2153 ) ;
  assign n2155 = ( ~n2151 & n2153 ) | ( ~n2151 & n2154 ) | ( n2153 & n2154 ) ;
  assign n2156 = ( ~n2150 & n2154 ) | ( ~n2150 & n2155 ) | ( n2154 & n2155 ) ;
  assign n2157 = ~n2139 & n2156 ;
  assign n2158 = ( ~n2102 & n2156 ) | ( ~n2102 & n2157 ) | ( n2156 & n2157 ) ;
  assign n2159 = ( n2140 & n2142 ) | ( n2140 & ~n2158 ) | ( n2142 & ~n2158 ) ;
  assign n2160 = n2054 & ~n2150 ;
  assign n2161 = ( n2067 & ~n2150 ) | ( n2067 & n2160 ) | ( ~n2150 & n2160 ) ;
  assign n2162 = ~n2151 & n2161 ;
  assign n2163 = n2151 & ~n2153 ;
  assign n2164 = ( ~n2150 & n2162 ) | ( ~n2150 & n2163 ) | ( n2162 & n2163 ) ;
  assign n2165 = n462 | n879 ;
  assign n2166 = n424 | n2165 ;
  assign n2167 = ( ~n474 & n879 ) | ( ~n474 & n2166 ) | ( n879 & n2166 ) ;
  assign n2168 = n491 & n2167 ;
  assign n2169 = ( ~n383 & n2167 ) | ( ~n383 & n2168 ) | ( n2167 & n2168 ) ;
  assign n2170 = n304 & n473 ;
  assign n2171 = ( n473 & n922 ) | ( n473 & n2170 ) | ( n922 & n2170 ) ;
  assign n2172 = ( ~n900 & n921 ) | ( ~n900 & n2171 ) | ( n921 & n2171 ) ;
  assign n2173 = ( n473 & n900 ) | ( n473 & n2172 ) | ( n900 & n2172 ) ;
  assign n2174 = n463 & n879 ;
  assign n2175 = ( ~n381 & n879 ) | ( ~n381 & n2174 ) | ( n879 & n2174 ) ;
  assign n2176 = ~n383 & n2175 ;
  assign n2177 = n2173 | n2176 ;
  assign n2178 = n2169 & ~n2177 ;
  assign n2179 = n2173 & n2176 ;
  assign n2180 = ( ~n2169 & n2173 ) | ( ~n2169 & n2179 ) | ( n2173 & n2179 ) ;
  assign n2181 = n2178 | n2180 ;
  assign n2182 = n754 | n1004 ;
  assign n2183 = ( ~n757 & n1004 ) | ( ~n757 & n2182 ) | ( n1004 & n2182 ) ;
  assign n2184 = n716 | n2183 ;
  assign n2185 = n754 & n1004 ;
  assign n2186 = ( ~n714 & n1004 ) | ( ~n714 & n2185 ) | ( n1004 & n2185 ) ;
  assign n2187 = ~n716 & n2186 ;
  assign n2188 = n2184 & ~n2187 ;
  assign n2189 = ( ~n773 & n942 ) | ( ~n773 & n2188 ) | ( n942 & n2188 ) ;
  assign n2190 = ( n756 & n942 ) | ( n756 & ~n2188 ) | ( n942 & ~n2188 ) ;
  assign n2191 = n2189 & ~n2190 ;
  assign n2192 = ~n2181 & n2191 ;
  assign n2193 = n2181 & ~n2191 ;
  assign n2194 = n2192 | n2193 ;
  assign n2195 = n2151 & n2153 ;
  assign n2196 = ~n2194 & n2195 ;
  assign n2197 = ( n2164 & ~n2194 ) | ( n2164 & n2196 ) | ( ~n2194 & n2196 ) ;
  assign n2198 = n2194 & ~n2195 ;
  assign n2199 = ~n2164 & n2198 ;
  assign n2200 = n2197 | n2199 ;
  assign n2201 = ( n2112 & n2122 ) | ( n2112 & n2135 ) | ( n2122 & n2135 ) ;
  assign n2202 = n642 | n1045 ;
  assign n2203 = ( n642 & ~n1049 ) | ( n642 & n2202 ) | ( ~n1049 & n2202 ) ;
  assign n2204 = n1042 | n2203 ;
  assign n2205 = n642 & n1045 ;
  assign n2206 = ( n642 & ~n1040 ) | ( n642 & n2205 ) | ( ~n1040 & n2205 ) ;
  assign n2207 = ~n1042 & n2206 ;
  assign n2208 = n2204 & ~n2207 ;
  assign n2209 = ( n634 & ~n1099 ) | ( n634 & n2208 ) | ( ~n1099 & n2208 ) ;
  assign n2210 = ( n634 & n1088 ) | ( n634 & ~n2208 ) | ( n1088 & ~n2208 ) ;
  assign n2211 = n2209 & ~n2210 ;
  assign n2212 = n2088 | n2146 ;
  assign n2213 = ( n2146 & ~n2147 ) | ( n2146 & n2212 ) | ( ~n2147 & n2212 ) ;
  assign n2214 = ( n2135 & n2211 ) | ( n2135 & ~n2213 ) | ( n2211 & ~n2213 ) ;
  assign n2215 = ( n2112 & n2211 ) | ( n2112 & ~n2213 ) | ( n2211 & ~n2213 ) ;
  assign n2216 = ( n2122 & n2214 ) | ( n2122 & n2215 ) | ( n2214 & n2215 ) ;
  assign n2217 = ( n2135 & ~n2211 ) | ( n2135 & n2213 ) | ( ~n2211 & n2213 ) ;
  assign n2218 = ( n2112 & ~n2211 ) | ( n2112 & n2213 ) | ( ~n2211 & n2213 ) ;
  assign n2219 = ( n2122 & n2217 ) | ( n2122 & n2218 ) | ( n2217 & n2218 ) ;
  assign n2220 = ( ~n2201 & n2216 ) | ( ~n2201 & n2219 ) | ( n2216 & n2219 ) ;
  assign n2221 = n2200 | n2220 ;
  assign n2222 = n2200 & ~n2220 ;
  assign n2223 = ( ~n2200 & n2221 ) | ( ~n2200 & n2222 ) | ( n2221 & n2222 ) ;
  assign n2224 = n2159 & n2223 ;
  assign n2225 = n2159 | n2223 ;
  assign n2226 = ~n2224 & n2225 ;
  assign n2227 = n2142 & n2156 ;
  assign n2228 = n2142 | n2156 ;
  assign n2229 = ~n2227 & n2228 ;
  assign n2230 = n1901 | n1972 ;
  assign n2231 = ( n1900 & n1972 ) | ( n1900 & n2230 ) | ( n1972 & n2230 ) ;
  assign n2233 = n1824 | n1828 ;
  assign n2234 = ( n1824 & ~n1826 ) | ( n1824 & n2233 ) | ( ~n1826 & n2233 ) ;
  assign n2235 = n2231 & n2234 ;
  assign n2236 = n1903 & n2234 ;
  assign n2237 = ( n1904 & n2235 ) | ( n1904 & n2236 ) | ( n2235 & n2236 ) ;
  assign n2232 = ( n1903 & n1904 ) | ( n1903 & n2231 ) | ( n1904 & n2231 ) ;
  assign n2238 = n2232 & ~n2237 ;
  assign n2239 = n2074 & n2100 ;
  assign n2240 = n2074 | n2100 ;
  assign n2241 = ~n2239 & n2240 ;
  assign n2242 = ~n2231 & n2234 ;
  assign n2243 = ~n1903 & n2234 ;
  assign n2244 = ( ~n1904 & n2242 ) | ( ~n1904 & n2243 ) | ( n2242 & n2243 ) ;
  assign n2245 = ~n2241 & n2244 ;
  assign n2246 = ( n2238 & ~n2241 ) | ( n2238 & n2245 ) | ( ~n2241 & n2245 ) ;
  assign n2247 = n2237 | n2246 ;
  assign n2248 = ~n2229 & n2247 ;
  assign n2249 = ~n2226 & n2248 ;
  assign n2250 = n2229 & ~n2247 ;
  assign n2251 = n2248 | n2250 ;
  assign n2252 = n2238 | n2244 ;
  assign n2253 = ~n2246 & n2252 ;
  assign n2254 = n1858 | n1975 ;
  assign n2255 = ( n1858 & ~n1864 ) | ( n1858 & n2254 ) | ( ~n1864 & n2254 ) ;
  assign n2256 = n2241 | n2244 ;
  assign n2257 = n2238 | n2256 ;
  assign n2258 = n2255 & ~n2257 ;
  assign n2259 = ( n2253 & n2255 ) | ( n2253 & n2258 ) | ( n2255 & n2258 ) ;
  assign n2260 = ~n2251 & n2259 ;
  assign n2261 = ( ~n2241 & n2252 ) | ( ~n2241 & n2255 ) | ( n2252 & n2255 ) ;
  assign n2262 = ( n2241 & ~n2252 ) | ( n2241 & n2255 ) | ( ~n2252 & n2255 ) ;
  assign n2263 = ( ~n2255 & n2261 ) | ( ~n2255 & n2262 ) | ( n2261 & n2262 ) ;
  assign n2264 = ( n2251 & ~n2260 ) | ( n2251 & n2263 ) | ( ~n2260 & n2263 ) ;
  assign n2265 = ( n2226 & ~n2249 ) | ( n2226 & n2264 ) | ( ~n2249 & n2264 ) ;
  assign n2266 = n2003 & ~n2263 ;
  assign n2267 = ( ~n2251 & n2260 ) | ( ~n2251 & n2266 ) | ( n2260 & n2266 ) ;
  assign n2268 = ( ~n2226 & n2249 ) | ( ~n2226 & n2267 ) | ( n2249 & n2267 ) ;
  assign n2269 = ( n2040 & n2265 ) | ( n2040 & ~n2268 ) | ( n2265 & ~n2268 ) ;
  assign n2270 = n1308 | n2034 ;
  assign n2271 = ( n2034 & ~n2036 ) | ( n2034 & n2270 ) | ( ~n2036 & n2270 ) ;
  assign n2272 = ~n2027 & n2029 ;
  assign n2273 = ( n2027 & n2271 ) | ( n2027 & ~n2272 ) | ( n2271 & ~n2272 ) ;
  assign n2274 = ( ~n2251 & n2260 ) | ( ~n2251 & n2273 ) | ( n2260 & n2273 ) ;
  assign n2275 = ~n2003 & n2005 ;
  assign n2276 = n2263 | n2275 ;
  assign n2277 = ( n2226 & ~n2249 ) | ( n2226 & n2276 ) | ( ~n2249 & n2276 ) ;
  assign n2278 = ( n2268 & n2274 ) | ( n2268 & ~n2277 ) | ( n2274 & ~n2277 ) ;
  assign n2279 = ( n1736 & n2269 ) | ( n1736 & ~n2278 ) | ( n2269 & ~n2278 ) ;
  assign n2280 = n2226 & ~n2248 ;
  assign n2281 = ~n2267 & n2280 ;
  assign n2282 = n2276 & n2280 ;
  assign n2283 = ( ~n2274 & n2281 ) | ( ~n2274 & n2282 ) | ( n2281 & n2282 ) ;
  assign n2284 = n2264 & n2280 ;
  assign n2285 = ( n2040 & n2281 ) | ( n2040 & n2284 ) | ( n2281 & n2284 ) ;
  assign n2286 = ( n1736 & n2283 ) | ( n1736 & n2285 ) | ( n2283 & n2285 ) ;
  assign n2287 = n2279 & ~n2286 ;
  assign n2288 = n564 | n565 ;
  assign n2289 = n561 | n2288 ;
  assign n2290 = n155 | n229 ;
  assign n2291 = n141 | n316 ;
  assign n2292 = n2290 | n2291 ;
  assign n2293 = n249 | n305 ;
  assign n2294 = n407 | n2293 ;
  assign n2295 = ( ~n2288 & n2292 ) | ( ~n2288 & n2294 ) | ( n2292 & n2294 ) ;
  assign n2296 = n2292 & n2294 ;
  assign n2297 = ( ~n561 & n2295 ) | ( ~n561 & n2296 ) | ( n2295 & n2296 ) ;
  assign n2298 = n2289 | n2297 ;
  assign n2299 = n508 | n513 ;
  assign n2300 = n398 | n780 ;
  assign n2301 = n690 | n2300 ;
  assign n2302 = n260 | n353 ;
  assign n2303 = n216 | n311 ;
  assign n2304 = n2302 | n2303 ;
  assign n2305 = n202 | n2304 ;
  assign n2306 = n2301 | n2305 ;
  assign n2307 = n2299 | n2306 ;
  assign n2308 = n269 | n354 ;
  assign n2309 = n256 | n293 ;
  assign n2310 = n2308 | n2309 ;
  assign n2311 = n173 | n728 ;
  assign n2312 = n2310 | n2311 ;
  assign n2313 = n212 | n2312 ;
  assign n2314 = n150 | n283 ;
  assign n2315 = n227 | n232 ;
  assign n2316 = n2314 | n2315 ;
  assign n2317 = n301 | n435 ;
  assign n2318 = n235 | n2317 ;
  assign n2319 = n2316 | n2318 ;
  assign n2320 = n206 | n360 ;
  assign n2321 = n2319 | n2320 ;
  assign n2322 = n2313 | n2321 ;
  assign n2323 = n2307 | n2322 ;
  assign n2324 = n2298 | n2323 ;
  assign n2325 = ~n2287 & n2324 ;
  assign n2326 = n2287 | n2325 ;
  assign n2327 = n2287 & n2324 ;
  assign n2328 = n2326 & ~n2327 ;
  assign n2329 = ( n2040 & n2264 ) | ( n2040 & ~n2267 ) | ( n2264 & ~n2267 ) ;
  assign n2330 = ( n2267 & n2274 ) | ( n2267 & ~n2276 ) | ( n2274 & ~n2276 ) ;
  assign n2331 = ( n1736 & n2329 ) | ( n1736 & ~n2330 ) | ( n2329 & ~n2330 ) ;
  assign n2332 = ( n2266 & n2273 ) | ( n2266 & ~n2276 ) | ( n2273 & ~n2276 ) ;
  assign n2333 = n2251 & ~n2259 ;
  assign n2334 = ~n2332 & n2333 ;
  assign n2335 = ( n2039 & ~n2263 ) | ( n2039 & n2266 ) | ( ~n2263 & n2266 ) ;
  assign n2336 = ( n2005 & n2263 ) | ( n2005 & ~n2266 ) | ( n2263 & ~n2266 ) ;
  assign n2337 = ( n2038 & ~n2335 ) | ( n2038 & n2336 ) | ( ~n2335 & n2336 ) ;
  assign n2338 = n2333 & n2337 ;
  assign n2339 = ( n1736 & n2334 ) | ( n1736 & n2338 ) | ( n2334 & n2338 ) ;
  assign n2340 = n2331 & ~n2339 ;
  assign n2341 = n525 | n557 ;
  assign n2342 = n146 | n2341 ;
  assign n2343 = n358 | n408 ;
  assign n2344 = n305 | n407 ;
  assign n2345 = n2343 | n2344 ;
  assign n2346 = n2342 | n2345 ;
  assign n2347 = n161 | n249 ;
  assign n2348 = n248 | n2347 ;
  assign n2349 = n150 | n316 ;
  assign n2350 = n294 | n2349 ;
  assign n2351 = n2348 | n2350 ;
  assign n2352 = n677 | n788 ;
  assign n2353 = n2351 | n2352 ;
  assign n2354 = n541 | n2353 ;
  assign n2355 = n2346 | n2354 ;
  assign n2356 = n361 | n603 ;
  assign n2357 = n601 | n2356 ;
  assign n2358 = n599 | n2357 ;
  assign n2359 = n236 | n270 ;
  assign n2360 = n220 | n689 ;
  assign n2361 = n1021 | n2360 ;
  assign n2362 = n2359 | n2361 ;
  assign n2363 = n229 | n289 ;
  assign n2364 = n217 | n2363 ;
  assign n2365 = n2362 | n2364 ;
  assign n2366 = n522 | n2365 ;
  assign n2367 = n2358 | n2366 ;
  assign n2368 = n2355 | n2367 ;
  assign n2369 = ~n2340 & n2368 ;
  assign n2370 = n2340 & ~n2368 ;
  assign n2371 = n2369 | n2370 ;
  assign n2372 = ~n2369 & n2371 ;
  assign n2373 = n2328 | n2372 ;
  assign n2374 = n2159 & ~n2223 ;
  assign n2375 = n754 & n879 ;
  assign n2376 = ( ~n714 & n879 ) | ( ~n714 & n2375 ) | ( n879 & n2375 ) ;
  assign n2377 = ~n716 & n2376 ;
  assign n2378 = n753 | n879 ;
  assign n2379 = n736 | n2378 ;
  assign n2380 = ( ~n757 & n879 ) | ( ~n757 & n2379 ) | ( n879 & n2379 ) ;
  assign n2381 = n772 & n2380 ;
  assign n2382 = ( ~n716 & n2380 ) | ( ~n716 & n2381 ) | ( n2380 & n2381 ) ;
  assign n2383 = ~n2377 & n2382 ;
  assign n2384 = n304 & n634 ;
  assign n2385 = ( n634 & n922 ) | ( n634 & n2384 ) | ( n922 & n2384 ) ;
  assign n2386 = ( ~n900 & n921 ) | ( ~n900 & n2385 ) | ( n921 & n2385 ) ;
  assign n2387 = ( n634 & n900 ) | ( n634 & n2386 ) | ( n900 & n2386 ) ;
  assign n2388 = n2383 & ~n2387 ;
  assign n2389 = ~n2383 & n2387 ;
  assign n2390 = n2388 | n2389 ;
  assign n2391 = n1004 | n1045 ;
  assign n2392 = ( n1004 & ~n1049 ) | ( n1004 & n2391 ) | ( ~n1049 & n2391 ) ;
  assign n2393 = n1042 | n2392 ;
  assign n2394 = n1004 & n1045 ;
  assign n2395 = ( n1004 & ~n1040 ) | ( n1004 & n2394 ) | ( ~n1040 & n2394 ) ;
  assign n2396 = ~n1042 & n2395 ;
  assign n2397 = n2393 & ~n2396 ;
  assign n2398 = ( n942 & ~n1099 ) | ( n942 & n2397 ) | ( ~n1099 & n2397 ) ;
  assign n2399 = ( n942 & n1088 ) | ( n942 & ~n2397 ) | ( n1088 & ~n2397 ) ;
  assign n2400 = n2398 & ~n2399 ;
  assign n2401 = ~n2390 & n2400 ;
  assign n2402 = n2390 & ~n2400 ;
  assign n2403 = n2401 | n2402 ;
  assign n2404 = n754 | n942 ;
  assign n2405 = ( ~n757 & n942 ) | ( ~n757 & n2404 ) | ( n942 & n2404 ) ;
  assign n2406 = n716 | n2405 ;
  assign n2407 = n754 & n942 ;
  assign n2408 = ( ~n714 & n942 ) | ( ~n714 & n2407 ) | ( n942 & n2407 ) ;
  assign n2409 = ~n716 & n2408 ;
  assign n2410 = n2406 & ~n2409 ;
  assign n2411 = ( ~n773 & n879 ) | ( ~n773 & n2410 ) | ( n879 & n2410 ) ;
  assign n2412 = ( n756 & n879 ) | ( n756 & ~n2410 ) | ( n879 & ~n2410 ) ;
  assign n2413 = n2411 & ~n2412 ;
  assign n2414 = n634 | n1045 ;
  assign n2415 = ( n634 & ~n1049 ) | ( n634 & n2414 ) | ( ~n1049 & n2414 ) ;
  assign n2416 = n1042 | n2415 ;
  assign n2417 = n634 & n1045 ;
  assign n2418 = ( n634 & ~n1040 ) | ( n634 & n2417 ) | ( ~n1040 & n2417 ) ;
  assign n2419 = ~n1042 & n2418 ;
  assign n2420 = n2416 & ~n2419 ;
  assign n2421 = ( n1004 & ~n1099 ) | ( n1004 & n2420 ) | ( ~n1099 & n2420 ) ;
  assign n2422 = ( n1004 & n1088 ) | ( n1004 & ~n2420 ) | ( n1088 & ~n2420 ) ;
  assign n2423 = n2421 & ~n2422 ;
  assign n2424 = n2413 & n2423 ;
  assign n2425 = n2413 | n2423 ;
  assign n2426 = ~n2424 & n2425 ;
  assign n2427 = ~n2178 & n2181 ;
  assign n2428 = ( n2178 & n2191 ) | ( n2178 & ~n2427 ) | ( n2191 & ~n2427 ) ;
  assign n2429 = n2426 & n2428 ;
  assign n2432 = ~n463 & n2173 ;
  assign n2433 = ( n474 & n2173 ) | ( n474 & n2432 ) | ( n2173 & n2432 ) ;
  assign n2430 = n463 & ~n2173 ;
  assign n2431 = ~n474 & n2430 ;
  assign n2434 = n2431 | n2433 ;
  assign n2435 = n304 & n642 ;
  assign n2436 = ( n642 & n922 ) | ( n642 & n2435 ) | ( n922 & n2435 ) ;
  assign n2437 = ( ~n900 & n921 ) | ( ~n900 & n2436 ) | ( n921 & n2436 ) ;
  assign n2438 = ( n642 & n900 ) | ( n642 & n2437 ) | ( n900 & n2437 ) ;
  assign n2439 = n2433 | n2438 ;
  assign n2440 = ( n2433 & ~n2434 ) | ( n2433 & n2439 ) | ( ~n2434 & n2439 ) ;
  assign n2441 = n2423 & n2440 ;
  assign n2442 = n2413 & n2441 ;
  assign n2443 = ( n2428 & n2440 ) | ( n2428 & n2442 ) | ( n2440 & n2442 ) ;
  assign n2444 = n2440 & n2442 ;
  assign n2445 = ( n2426 & n2443 ) | ( n2426 & n2444 ) | ( n2443 & n2444 ) ;
  assign n2446 = ( n2424 & n2429 ) | ( n2424 & ~n2445 ) | ( n2429 & ~n2445 ) ;
  assign n2447 = n2440 & ~n2442 ;
  assign n2448 = ~n2403 & n2447 ;
  assign n2449 = ~n2429 & n2448 ;
  assign n2450 = ( ~n2403 & n2446 ) | ( ~n2403 & n2449 ) | ( n2446 & n2449 ) ;
  assign n2451 = n2403 & ~n2447 ;
  assign n2452 = ( n2403 & n2429 ) | ( n2403 & n2451 ) | ( n2429 & n2451 ) ;
  assign n2453 = ~n2446 & n2452 ;
  assign n2454 = n2450 | n2453 ;
  assign n2455 = n2211 & n2213 ;
  assign n2456 = n2211 & ~n2455 ;
  assign n2457 = ~n2211 & n2213 ;
  assign n2458 = n2455 | n2457 ;
  assign n2459 = n2456 | n2458 ;
  assign n2460 = ~n2434 & n2438 ;
  assign n2461 = n2434 & ~n2438 ;
  assign n2462 = n2460 | n2461 ;
  assign n2463 = n2135 & ~n2462 ;
  assign n2464 = n2112 & ~n2462 ;
  assign n2465 = ( n2122 & n2463 ) | ( n2122 & n2464 ) | ( n2463 & n2464 ) ;
  assign n2466 = n2213 & ~n2462 ;
  assign n2467 = n2211 & n2466 ;
  assign n2468 = ( n2459 & n2465 ) | ( n2459 & n2467 ) | ( n2465 & n2467 ) ;
  assign n2469 = ~n2135 & n2462 ;
  assign n2470 = ~n2112 & n2462 ;
  assign n2471 = ( ~n2122 & n2469 ) | ( ~n2122 & n2470 ) | ( n2469 & n2470 ) ;
  assign n2472 = ~n2213 & n2462 ;
  assign n2473 = ( ~n2211 & n2462 ) | ( ~n2211 & n2472 ) | ( n2462 & n2472 ) ;
  assign n2474 = ( ~n2459 & n2471 ) | ( ~n2459 & n2473 ) | ( n2471 & n2473 ) ;
  assign n2475 = n2468 | n2474 ;
  assign n2476 = n2426 | n2428 ;
  assign n2477 = ~n2429 & n2476 ;
  assign n2478 = ~n2475 & n2477 ;
  assign n2479 = n2468 | n2478 ;
  assign n2480 = n2454 & n2479 ;
  assign n2481 = n2454 | n2479 ;
  assign n2482 = ~n2480 & n2481 ;
  assign n2483 = n2475 & ~n2477 ;
  assign n2484 = n2478 | n2483 ;
  assign n2485 = n2196 | n2220 ;
  assign n2486 = n2194 & ~n2220 ;
  assign n2487 = ( n2164 & n2485 ) | ( n2164 & ~n2486 ) | ( n2485 & ~n2486 ) ;
  assign n2488 = ( n2197 & ~n2200 ) | ( n2197 & n2487 ) | ( ~n2200 & n2487 ) ;
  assign n2489 = ~n2484 & n2488 ;
  assign n2490 = ~n2482 & n2489 ;
  assign n2491 = n2484 & ~n2488 ;
  assign n2492 = n2489 | n2491 ;
  assign n2493 = ( n2482 & ~n2490 ) | ( n2482 & n2492 ) | ( ~n2490 & n2492 ) ;
  assign n2494 = ( n2374 & n2490 ) | ( n2374 & ~n2493 ) | ( n2490 & ~n2493 ) ;
  assign n2495 = ~n2490 & n2493 ;
  assign n2496 = ( n2226 & ~n2494 ) | ( n2226 & n2495 ) | ( ~n2494 & n2495 ) ;
  assign n2497 = n2374 & ~n2492 ;
  assign n2498 = ( n2226 & n2492 ) | ( n2226 & ~n2497 ) | ( n2492 & ~n2497 ) ;
  assign n2499 = ( ~n2482 & n2490 ) | ( ~n2482 & n2497 ) | ( n2490 & n2497 ) ;
  assign n2500 = ( n2248 & ~n2482 ) | ( n2248 & n2490 ) | ( ~n2482 & n2490 ) ;
  assign n2501 = ( ~n2498 & n2499 ) | ( ~n2498 & n2500 ) | ( n2499 & n2500 ) ;
  assign n2502 = ( n2264 & n2496 ) | ( n2264 & ~n2501 ) | ( n2496 & ~n2501 ) ;
  assign n2503 = ( n2267 & ~n2496 ) | ( n2267 & n2501 ) | ( ~n2496 & n2501 ) ;
  assign n2504 = ( n2040 & n2502 ) | ( n2040 & ~n2503 ) | ( n2502 & ~n2503 ) ;
  assign n2505 = ( n2276 & n2496 ) | ( n2276 & ~n2501 ) | ( n2496 & ~n2501 ) ;
  assign n2506 = ( n2274 & n2503 ) | ( n2274 & ~n2505 ) | ( n2503 & ~n2505 ) ;
  assign n2507 = ( n1736 & n2504 ) | ( n1736 & ~n2506 ) | ( n2504 & ~n2506 ) ;
  assign n2508 = ~n2489 & n2492 ;
  assign n2509 = ( n2374 & n2489 ) | ( n2374 & ~n2508 ) | ( n2489 & ~n2508 ) ;
  assign n2510 = ( n2226 & n2508 ) | ( n2226 & ~n2509 ) | ( n2508 & ~n2509 ) ;
  assign n2511 = n2482 & n2510 ;
  assign n2512 = n2482 & ~n2489 ;
  assign n2513 = ~n2497 & n2512 ;
  assign n2514 = ~n2248 & n2512 ;
  assign n2515 = ( n2498 & n2513 ) | ( n2498 & n2514 ) | ( n2513 & n2514 ) ;
  assign n2516 = ( n2264 & n2511 ) | ( n2264 & n2515 ) | ( n2511 & n2515 ) ;
  assign n2517 = ( ~n2267 & n2511 ) | ( ~n2267 & n2515 ) | ( n2511 & n2515 ) ;
  assign n2518 = ( n2040 & n2516 ) | ( n2040 & n2517 ) | ( n2516 & n2517 ) ;
  assign n2519 = ( n2276 & n2511 ) | ( n2276 & n2515 ) | ( n2511 & n2515 ) ;
  assign n2520 = ( ~n2274 & n2517 ) | ( ~n2274 & n2519 ) | ( n2517 & n2519 ) ;
  assign n2521 = ( n1736 & n2518 ) | ( n1736 & n2520 ) | ( n2518 & n2520 ) ;
  assign n2522 = n2507 & ~n2521 ;
  assign n2523 = n411 | n676 ;
  assign n2524 = n193 | n202 ;
  assign n2525 = n549 | n2524 ;
  assign n2526 = n167 | n344 ;
  assign n2527 = n248 | n2526 ;
  assign n2528 = n2525 | n2527 ;
  assign n2529 = n283 | n2528 ;
  assign n2530 = n2523 | n2529 ;
  assign n2531 = n232 | n372 ;
  assign n2532 = n236 | n2531 ;
  assign n2533 = n2530 | n2532 ;
  assign n2534 = n182 | n198 ;
  assign n2535 = n212 | n2534 ;
  assign n2536 = n737 | n2535 ;
  assign n2537 = n220 | n347 ;
  assign n2538 = n205 | n2537 ;
  assign n2539 = n392 | n2538 ;
  assign n2540 = n2536 | n2539 ;
  assign n2541 = n391 | n690 ;
  assign n2542 = n2540 | n2541 ;
  assign n2543 = n2533 | n2542 ;
  assign n2544 = n172 | n709 ;
  assign n2545 = n574 | n2544 ;
  assign n2546 = n284 | n354 ;
  assign n2547 = n570 | n2546 ;
  assign n2548 = n2545 | n2547 ;
  assign n2549 = n223 | n435 ;
  assign n2550 = n313 | n2549 ;
  assign n2551 = n696 | n2550 ;
  assign n2552 = n2548 | n2551 ;
  assign n2553 = n235 | n446 ;
  assign n2554 = n348 | n528 ;
  assign n2555 = n256 | n2554 ;
  assign n2556 = n2553 | n2555 ;
  assign n2557 = n2552 | n2556 ;
  assign n2558 = n304 | n428 ;
  assign n2559 = n189 | n245 ;
  assign n2560 = n2558 | n2559 ;
  assign n2561 = n320 | n426 ;
  assign n2562 = n278 | n2561 ;
  assign n2563 = n2560 | n2562 ;
  assign n2564 = n2557 | n2563 ;
  assign n2565 = n2543 | n2564 ;
  assign n2566 = ~n2522 & n2565 ;
  assign n2567 = n2522 & ~n2565 ;
  assign n2568 = n2566 | n2567 ;
  assign n2569 = ( n2248 & n2497 ) | ( n2248 & ~n2498 ) | ( n2497 & ~n2498 ) ;
  assign n2570 = ( n2264 & n2498 ) | ( n2264 & ~n2569 ) | ( n2498 & ~n2569 ) ;
  assign n2571 = ( n2267 & ~n2498 ) | ( n2267 & n2569 ) | ( ~n2498 & n2569 ) ;
  assign n2572 = ( n2040 & n2570 ) | ( n2040 & ~n2571 ) | ( n2570 & ~n2571 ) ;
  assign n2573 = ( n2276 & n2498 ) | ( n2276 & ~n2569 ) | ( n2498 & ~n2569 ) ;
  assign n2574 = ( n2274 & n2571 ) | ( n2274 & ~n2573 ) | ( n2571 & ~n2573 ) ;
  assign n2575 = ( n1736 & n2572 ) | ( n1736 & ~n2574 ) | ( n2572 & ~n2574 ) ;
  assign n2576 = ~n2374 & n2492 ;
  assign n2577 = n2226 & n2576 ;
  assign n2578 = ( ~n2248 & n2576 ) | ( ~n2248 & n2577 ) | ( n2576 & n2577 ) ;
  assign n2579 = ( n2264 & n2577 ) | ( n2264 & n2578 ) | ( n2577 & n2578 ) ;
  assign n2580 = ( ~n2267 & n2577 ) | ( ~n2267 & n2578 ) | ( n2577 & n2578 ) ;
  assign n2581 = ( n2040 & n2579 ) | ( n2040 & n2580 ) | ( n2579 & n2580 ) ;
  assign n2582 = ( n2276 & n2577 ) | ( n2276 & n2578 ) | ( n2577 & n2578 ) ;
  assign n2583 = ( ~n2274 & n2580 ) | ( ~n2274 & n2582 ) | ( n2580 & n2582 ) ;
  assign n2584 = ( n1736 & n2581 ) | ( n1736 & n2583 ) | ( n2581 & n2583 ) ;
  assign n2585 = n2575 & ~n2584 ;
  assign n2586 = n289 | n339 ;
  assign n2587 = n2560 | n2586 ;
  assign n2588 = n2557 | n2587 ;
  assign n2589 = n368 | n397 ;
  assign n2590 = n311 | n2589 ;
  assign n2591 = n363 | n2590 ;
  assign n2592 = n167 | n301 ;
  assign n2593 = n456 | n2592 ;
  assign n2594 = n2591 | n2593 ;
  assign n2595 = n202 | n210 ;
  assign n2596 = n125 | n2595 ;
  assign n2597 = ( n139 & ~n831 ) | ( n139 & n2596 ) | ( ~n831 & n2596 ) ;
  assign n2598 = n510 & ~n831 ;
  assign n2599 = ~n2597 & n2598 ;
  assign n2600 = ~n2594 & n2599 ;
  assign n2601 = n906 | n2538 ;
  assign n2602 = n241 | n261 ;
  assign n2603 = n728 | n2602 ;
  assign n2604 = n2601 | n2603 ;
  assign n2605 = n343 | n412 ;
  assign n2606 = n233 | n384 ;
  assign n2607 = n2605 | n2606 ;
  assign n2608 = n198 | n2607 ;
  assign n2609 = n257 | n495 ;
  assign n2610 = n300 | n2609 ;
  assign n2611 = n425 | n701 ;
  assign n2612 = n590 | n2611 ;
  assign n2613 = n2610 | n2612 ;
  assign n2614 = n2608 | n2613 ;
  assign n2615 = n2604 | n2614 ;
  assign n2616 = n2600 & ~n2615 ;
  assign n2617 = ~n2588 & n2616 ;
  assign n2618 = n2585 | n2617 ;
  assign n2619 = n2325 & n2618 ;
  assign n2620 = n2585 & n2617 ;
  assign n2621 = n2618 & n2620 ;
  assign n2622 = ( n2618 & ~n2619 ) | ( n2618 & n2621 ) | ( ~n2619 & n2621 ) ;
  assign n2623 = n2568 | n2622 ;
  assign n2624 = n2618 & ~n2620 ;
  assign n2625 = n2618 & ~n2624 ;
  assign n2626 = n2568 | n2625 ;
  assign n2627 = ( n2373 & n2623 ) | ( n2373 & n2626 ) | ( n2623 & n2626 ) ;
  assign n2628 = ( n1736 & ~n2332 ) | ( n1736 & n2337 ) | ( ~n2332 & n2337 ) ;
  assign n2629 = n2263 & n2275 ;
  assign n2630 = ~n2003 & n2263 ;
  assign n2631 = ( ~n2273 & n2629 ) | ( ~n2273 & n2630 ) | ( n2629 & n2630 ) ;
  assign n2632 = ~n2039 & n2630 ;
  assign n2633 = n2005 & n2630 ;
  assign n2634 = ( n2038 & n2632 ) | ( n2038 & n2633 ) | ( n2632 & n2633 ) ;
  assign n2635 = ( n1736 & n2631 ) | ( n1736 & n2634 ) | ( n2631 & n2634 ) ;
  assign n2636 = n2628 & ~n2635 ;
  assign n2637 = n966 | n967 ;
  assign n2638 = n352 | n425 ;
  assign n2639 = n2302 | n2638 ;
  assign n2640 = n664 | n2639 ;
  assign n2641 = n2637 | n2640 ;
  assign n2642 = n235 | n452 ;
  assign n2643 = n446 | n2642 ;
  assign n2644 = n2641 | n2643 ;
  assign n2645 = n266 | n316 ;
  assign n2646 = n361 | n2645 ;
  assign n2647 = n159 | n392 ;
  assign n2648 = n2646 | n2647 ;
  assign n2649 = n730 | n2648 ;
  assign n2650 = n2644 | n2649 ;
  assign n2651 = n414 | n570 ;
  assign n2652 = n426 | n2651 ;
  assign n2653 = n125 | n293 ;
  assign n2654 = n2652 | n2653 ;
  assign n2655 = n553 | n2654 ;
  assign n2656 = n177 | n524 ;
  assign n2657 = n285 | n2656 ;
  assign n2658 = n219 | n228 ;
  assign n2659 = n2657 | n2658 ;
  assign n2660 = n2655 | n2659 ;
  assign n2661 = n372 | n545 ;
  assign n2662 = n398 | n2661 ;
  assign n2663 = n198 | n718 ;
  assign n2664 = n456 | n2663 ;
  assign n2665 = n2662 | n2664 ;
  assign n2666 = n223 | n334 ;
  assign n2667 = n175 | n2666 ;
  assign n2668 = n428 | n2667 ;
  assign n2669 = n2665 | n2668 ;
  assign n2670 = n2660 | n2669 ;
  assign n2671 = n2650 | n2670 ;
  assign n2672 = n233 | n304 ;
  assign n2673 = n131 | n360 ;
  assign n2674 = n2672 | n2673 ;
  assign n2675 = n2671 | n2674 ;
  assign n2676 = ~n2636 & n2675 ;
  assign n2677 = ~n2369 & n2676 ;
  assign n2678 = ~n2369 & n2370 ;
  assign n2679 = ( n2369 & n2677 ) | ( n2369 & ~n2678 ) | ( n2677 & ~n2678 ) ;
  assign n2680 = ~n2328 & n2679 ;
  assign n2681 = ( n2623 & n2626 ) | ( n2623 & ~n2680 ) | ( n2626 & ~n2680 ) ;
  assign n2682 = n2636 & ~n2675 ;
  assign n2683 = n2676 | n2682 ;
  assign n2684 = ~n2005 & n2273 ;
  assign n2685 = ( n1736 & n2040 ) | ( n1736 & ~n2684 ) | ( n2040 & ~n2684 ) ;
  assign n2686 = n2005 & ~n2273 ;
  assign n2687 = n2005 & ~n2027 ;
  assign n2688 = n2038 & n2687 ;
  assign n2689 = ( n1736 & n2686 ) | ( n1736 & n2688 ) | ( n2686 & n2688 ) ;
  assign n2690 = n2685 & ~n2689 ;
  assign n2691 = n315 | n435 ;
  assign n2692 = n426 | n511 ;
  assign n2693 = n2691 | n2692 ;
  assign n2694 = n339 | n2693 ;
  assign n2695 = n439 | n2535 ;
  assign n2696 = n549 | n886 ;
  assign n2697 = n2695 | n2696 ;
  assign n2698 = n384 | n408 ;
  assign n2699 = n305 | n361 ;
  assign n2700 = n2698 | n2699 ;
  assign n2701 = n2697 | n2700 ;
  assign n2702 = n740 | n890 ;
  assign n2703 = n173 | n333 ;
  assign n2704 = n718 | n2703 ;
  assign n2705 = n2702 | n2704 ;
  assign n2706 = n419 | n425 ;
  assign n2707 = n2705 | n2706 ;
  assign n2708 = n2701 | n2707 ;
  assign n2709 = n155 | n317 ;
  assign n2710 = n597 | n2709 ;
  assign n2711 = n256 | n267 ;
  assign n2712 = n320 | n2711 ;
  assign n2713 = n2710 | n2712 ;
  assign n2714 = n252 | n2713 ;
  assign n2715 = n2708 | n2714 ;
  assign n2716 = n2694 | n2715 ;
  assign n2717 = ~n2690 & n2716 ;
  assign n2718 = n2690 & ~n2716 ;
  assign n2719 = n2717 | n2718 ;
  assign n2720 = ~n2717 & n2719 ;
  assign n2721 = n425 | n2705 ;
  assign n2722 = n369 | n906 ;
  assign n2723 = n224 | n242 ;
  assign n2724 = n510 & ~n2723 ;
  assign n2725 = ~n2722 & n2724 ;
  assign n2726 = ~n2721 & n2725 ;
  assign n2727 = n547 | n593 ;
  assign n2728 = n2726 & ~n2727 ;
  assign n2729 = n174 | n402 ;
  assign n2730 = n400 | n2729 ;
  assign n2731 = n396 | n2730 ;
  assign n2732 = n2728 & ~n2731 ;
  assign n2733 = n456 | n701 ;
  assign n2734 = n344 | n495 ;
  assign n2735 = n2733 | n2734 ;
  assign n2736 = n330 | n2735 ;
  assign n2737 = n339 | n414 ;
  assign n2738 = n576 | n2737 ;
  assign n2739 = n2596 | n2738 ;
  assign n2740 = n2736 | n2739 ;
  assign n2741 = n131 | n965 ;
  assign n2742 = n531 | n2741 ;
  assign n2743 = n664 | n2359 ;
  assign n2744 = n2361 | n2743 ;
  assign n2745 = n2742 | n2744 ;
  assign n2746 = n2740 | n2745 ;
  assign n2747 = n185 | n354 ;
  assign n2748 = n176 | n384 ;
  assign n2749 = n2747 | n2748 ;
  assign n2750 = n248 | n361 ;
  assign n2751 = n2749 | n2750 ;
  assign n2752 = n2746 | n2751 ;
  assign n2753 = n2732 & ~n2752 ;
  assign n2754 = ( n1736 & n2037 ) | ( n1736 & ~n2271 ) | ( n2037 & ~n2271 ) ;
  assign n2755 = n2029 & ~n2271 ;
  assign n2756 = n2029 & n2037 ;
  assign n2757 = ( n1736 & n2755 ) | ( n1736 & n2756 ) | ( n2755 & n2756 ) ;
  assign n2758 = n2029 & ~n2037 ;
  assign n2759 = n2029 & n2271 ;
  assign n2760 = ( ~n1736 & n2758 ) | ( ~n1736 & n2759 ) | ( n2758 & n2759 ) ;
  assign n2761 = ( n2754 & ~n2757 ) | ( n2754 & n2760 ) | ( ~n2757 & n2760 ) ;
  assign n2762 = n2753 | n2761 ;
  assign n2763 = n2753 & n2761 ;
  assign n2764 = n2762 & ~n2763 ;
  assign n2765 = n1308 & ~n2036 ;
  assign n2766 = ( n1736 & n2036 ) | ( n1736 & ~n2765 ) | ( n2036 & ~n2765 ) ;
  assign n2767 = ~n1308 & n2036 ;
  assign n2768 = n1736 & n2767 ;
  assign n2769 = n2766 & ~n2768 ;
  assign n2770 = n594 | n2737 ;
  assign n2771 = n281 | n2770 ;
  assign n2772 = n2346 | n2771 ;
  assign n2773 = n343 | n545 ;
  assign n2774 = n352 | n709 ;
  assign n2775 = n2773 | n2774 ;
  assign n2776 = n174 | n2775 ;
  assign n2777 = n283 | n289 ;
  assign n2778 = n781 | n2777 ;
  assign n2779 = n360 | n426 ;
  assign n2780 = n2778 | n2779 ;
  assign n2781 = n2776 | n2780 ;
  assign n2782 = n311 | n412 ;
  assign n2783 = n210 | n257 ;
  assign n2784 = n2782 | n2783 ;
  assign n2785 = n277 | n2784 ;
  assign n2786 = n2781 | n2785 ;
  assign n2787 = n2772 | n2786 ;
  assign n2788 = n216 | n429 ;
  assign n2789 = n348 | n2788 ;
  assign n2790 = n332 | n2789 ;
  assign n2791 = n232 | n718 ;
  assign n2792 = n212 | n301 ;
  assign n2793 = n2791 | n2792 ;
  assign n2794 = n443 | n2793 ;
  assign n2795 = n2790 | n2794 ;
  assign n2796 = n2787 | n2795 ;
  assign n2797 = n270 | n556 ;
  assign n2798 = n195 | n820 ;
  assign n2799 = n2797 | n2798 ;
  assign n2800 = n664 | n2799 ;
  assign n2801 = n2701 | n2800 ;
  assign n2802 = n238 | n2801 ;
  assign n2803 = n427 | n2545 ;
  assign n2804 = n231 | n823 ;
  assign n2805 = n2803 | n2804 ;
  assign n2806 = n244 | n253 ;
  assign n2807 = n674 | n2806 ;
  assign n2808 = n280 | n2807 ;
  assign n2809 = n597 | n2808 ;
  assign n2810 = n2805 | n2809 ;
  assign n2811 = n338 | n443 ;
  assign n2812 = n501 | n701 ;
  assign n2813 = n2811 | n2812 ;
  assign n2814 = n277 | n372 ;
  assign n2815 = n175 | n2814 ;
  assign n2816 = n2813 | n2815 ;
  assign n2817 = n2810 | n2816 ;
  assign n2818 = n2802 | n2817 ;
  assign n2819 = n1310 & ~n1734 ;
  assign n2820 = n1732 & n2819 ;
  assign n2821 = n1736 & ~n2820 ;
  assign n2822 = ~n2818 & n2821 ;
  assign n2823 = ( n2769 & ~n2796 ) | ( n2769 & n2822 ) | ( ~n2796 & n2822 ) ;
  assign n2824 = n2762 & n2823 ;
  assign n2825 = ( n2762 & ~n2764 ) | ( n2762 & n2824 ) | ( ~n2764 & n2824 ) ;
  assign n2826 = ( ~n2717 & n2720 ) | ( ~n2717 & n2825 ) | ( n2720 & n2825 ) ;
  assign n2827 = n2683 | n2826 ;
  assign n2828 = ( n2627 & n2681 ) | ( n2627 & n2827 ) | ( n2681 & n2827 ) ;
  assign n2829 = n2226 & ~n2374 ;
  assign n2830 = n942 | n1045 ;
  assign n2831 = ( n942 & ~n1049 ) | ( n942 & n2830 ) | ( ~n1049 & n2830 ) ;
  assign n2832 = n1042 | n2831 ;
  assign n2833 = n942 & n1045 ;
  assign n2834 = ( n942 & ~n1040 ) | ( n942 & n2833 ) | ( ~n1040 & n2833 ) ;
  assign n2835 = ~n1042 & n2834 ;
  assign n2836 = n2832 & ~n2835 ;
  assign n2837 = ( n879 & ~n1099 ) | ( n879 & n2836 ) | ( ~n1099 & n2836 ) ;
  assign n2838 = ( n879 & n1088 ) | ( n879 & ~n2836 ) | ( n1088 & ~n2836 ) ;
  assign n2839 = n2837 & ~n2838 ;
  assign n2840 = n2388 | n2400 ;
  assign n2841 = ( n2388 & ~n2390 ) | ( n2388 & n2840 ) | ( ~n2390 & n2840 ) ;
  assign n2842 = n2839 & n2841 ;
  assign n2843 = n2839 | n2841 ;
  assign n2844 = ~n2842 & n2843 ;
  assign n2845 = ~n754 & n2387 ;
  assign n2846 = ( n757 & n2387 ) | ( n757 & n2845 ) | ( n2387 & n2845 ) ;
  assign n2847 = n754 & ~n2387 ;
  assign n2848 = ~n757 & n2847 ;
  assign n2849 = n2846 | n2848 ;
  assign n2850 = n304 & n1004 ;
  assign n2851 = ( n922 & n1004 ) | ( n922 & n2850 ) | ( n1004 & n2850 ) ;
  assign n2852 = ( ~n900 & n921 ) | ( ~n900 & n2851 ) | ( n921 & n2851 ) ;
  assign n2853 = ( n900 & n1004 ) | ( n900 & n2852 ) | ( n1004 & n2852 ) ;
  assign n2854 = ~n2849 & n2853 ;
  assign n2855 = n2849 & ~n2853 ;
  assign n2856 = n2854 | n2855 ;
  assign n2857 = n2844 & ~n2856 ;
  assign n2858 = ~n2844 & n2856 ;
  assign n2859 = n2857 | n2858 ;
  assign n2860 = n2445 & ~n2859 ;
  assign n2861 = ( n2450 & ~n2859 ) | ( n2450 & n2860 ) | ( ~n2859 & n2860 ) ;
  assign n2862 = ~n2445 & n2859 ;
  assign n2863 = ~n2450 & n2862 ;
  assign n2864 = n2861 | n2863 ;
  assign n2865 = ~n2454 & n2479 ;
  assign n2866 = n2493 & ~n2865 ;
  assign n2867 = n2864 | n2866 ;
  assign n2868 = n2490 | n2865 ;
  assign n2869 = ~n2864 & n2868 ;
  assign n2870 = ( n2829 & n2867 ) | ( n2829 & ~n2869 ) | ( n2867 & ~n2869 ) ;
  assign n2871 = ~n2864 & n2865 ;
  assign n2872 = ( n2482 & n2864 ) | ( n2482 & ~n2871 ) | ( n2864 & ~n2871 ) ;
  assign n2873 = ( n2489 & n2871 ) | ( n2489 & ~n2872 ) | ( n2871 & ~n2872 ) ;
  assign n2874 = ~n2871 & n2872 ;
  assign n2875 = ( n2497 & n2873 ) | ( n2497 & ~n2874 ) | ( n2873 & ~n2874 ) ;
  assign n2876 = ( n2248 & n2873 ) | ( n2248 & ~n2874 ) | ( n2873 & ~n2874 ) ;
  assign n2877 = ( ~n2498 & n2875 ) | ( ~n2498 & n2876 ) | ( n2875 & n2876 ) ;
  assign n2878 = ( n2264 & n2870 ) | ( n2264 & ~n2877 ) | ( n2870 & ~n2877 ) ;
  assign n2879 = ( n2267 & ~n2870 ) | ( n2267 & n2877 ) | ( ~n2870 & n2877 ) ;
  assign n2880 = ( n2040 & n2878 ) | ( n2040 & ~n2879 ) | ( n2878 & ~n2879 ) ;
  assign n2881 = ( n2276 & n2870 ) | ( n2276 & ~n2877 ) | ( n2870 & ~n2877 ) ;
  assign n2882 = ( n2274 & n2879 ) | ( n2274 & ~n2881 ) | ( n2879 & ~n2881 ) ;
  assign n2883 = ( n1736 & n2880 ) | ( n1736 & ~n2882 ) | ( n2880 & ~n2882 ) ;
  assign n2884 = n2864 & n2866 ;
  assign n2885 = n2864 & ~n2868 ;
  assign n2886 = ( n2829 & n2884 ) | ( n2829 & n2885 ) | ( n2884 & n2885 ) ;
  assign n2887 = ( n2454 & ~n2479 ) | ( n2454 & n2484 ) | ( ~n2479 & n2484 ) ;
  assign n2888 = ( n2488 & n2865 ) | ( n2488 & ~n2887 ) | ( n2865 & ~n2887 ) ;
  assign n2889 = n2864 & ~n2888 ;
  assign n2890 = n2454 & ~n2479 ;
  assign n2891 = n2864 & n2890 ;
  assign n2892 = ( ~n2497 & n2889 ) | ( ~n2497 & n2891 ) | ( n2889 & n2891 ) ;
  assign n2893 = ( ~n2248 & n2889 ) | ( ~n2248 & n2891 ) | ( n2889 & n2891 ) ;
  assign n2894 = ( n2498 & n2892 ) | ( n2498 & n2893 ) | ( n2892 & n2893 ) ;
  assign n2895 = ( n2264 & n2886 ) | ( n2264 & n2894 ) | ( n2886 & n2894 ) ;
  assign n2896 = ( ~n2267 & n2886 ) | ( ~n2267 & n2894 ) | ( n2886 & n2894 ) ;
  assign n2897 = ( n2040 & n2895 ) | ( n2040 & n2896 ) | ( n2895 & n2896 ) ;
  assign n2898 = ( n2276 & n2886 ) | ( n2276 & n2894 ) | ( n2886 & n2894 ) ;
  assign n2899 = ( ~n2274 & n2896 ) | ( ~n2274 & n2898 ) | ( n2896 & n2898 ) ;
  assign n2900 = ( n1736 & n2897 ) | ( n1736 & n2899 ) | ( n2897 & n2899 ) ;
  assign n2901 = n2883 & ~n2900 ;
  assign n2902 = n346 | n394 ;
  assign n2903 = n281 | n540 ;
  assign n2904 = n2902 | n2903 ;
  assign n2905 = n238 | n696 ;
  assign n2906 = n2904 | n2905 ;
  assign n2907 = n617 | n671 ;
  assign n2908 = n2906 | n2907 ;
  assign n2909 = n821 | n823 ;
  assign n2910 = n244 | n311 ;
  assign n2911 = n206 | n338 ;
  assign n2912 = n2910 | n2911 ;
  assign n2913 = n125 | n2912 ;
  assign n2914 = n2909 | n2913 ;
  assign n2915 = n812 | n2914 ;
  assign n2916 = n2908 | n2915 ;
  assign n2917 = n2901 & ~n2916 ;
  assign n2918 = ~n2901 & n2916 ;
  assign n2919 = n2566 & ~n2918 ;
  assign n2920 = n2917 & ~n2918 ;
  assign n2921 = ( n2918 & n2919 ) | ( n2918 & ~n2920 ) | ( n2919 & ~n2920 ) ;
  assign n2922 = n2917 | n2921 ;
  assign n2923 = n2828 & ~n2922 ;
  assign n2924 = ~n2566 & n2828 ;
  assign n2925 = n2566 & n2918 ;
  assign n2926 = ( ~n2828 & n2918 ) | ( ~n2828 & n2925 ) | ( n2918 & n2925 ) ;
  assign n2927 = ( n2917 & ~n2924 ) | ( n2917 & n2926 ) | ( ~n2924 & n2926 ) ;
  assign n2928 = n2923 | n2927 ;
  assign n2929 = n2917 | n2918 ;
  assign n2930 = ~n2918 & n2929 ;
  assign n2931 = ( n2828 & ~n2921 ) | ( n2828 & n2930 ) | ( ~n2921 & n2930 ) ;
  assign n2932 = n175 | n277 ;
  assign n2933 = n2810 | n2932 ;
  assign n2934 = n291 | n322 ;
  assign n2935 = n907 | n2934 ;
  assign n2936 = n208 | n2935 ;
  assign n2937 = n2594 | n2936 ;
  assign n2938 = n193 | n284 ;
  assign n2939 = n305 | n338 ;
  assign n2940 = n2938 | n2939 ;
  assign n2941 = n135 | n511 ;
  assign n2942 = n2940 | n2941 ;
  assign n2943 = n310 | n501 ;
  assign n2944 = n236 | n2943 ;
  assign n2945 = n165 | n267 ;
  assign n2946 = n233 | n245 ;
  assign n2947 = n2945 | n2946 ;
  assign n2948 = n2944 | n2947 ;
  assign n2949 = n2942 | n2948 ;
  assign n2950 = n2937 | n2949 ;
  assign n2951 = n2933 | n2950 ;
  assign n2952 = n256 | n354 ;
  assign n2953 = n2554 | n2952 ;
  assign n2954 = n144 | n155 ;
  assign n2955 = n242 | n2954 ;
  assign n2956 = n2953 | n2955 ;
  assign n2957 = n139 | n425 ;
  assign n2958 = n2956 | n2957 ;
  assign n2959 = n2951 | n2958 ;
  assign n2960 = n2861 | n2871 ;
  assign n2961 = n2872 & ~n2960 ;
  assign n2962 = n2489 | n2861 ;
  assign n2963 = ( ~n2872 & n2960 ) | ( ~n2872 & n2962 ) | ( n2960 & n2962 ) ;
  assign n2964 = ( n2497 & ~n2961 ) | ( n2497 & n2963 ) | ( ~n2961 & n2963 ) ;
  assign n2965 = ( n2248 & ~n2961 ) | ( n2248 & n2963 ) | ( ~n2961 & n2963 ) ;
  assign n2966 = ( ~n2498 & n2964 ) | ( ~n2498 & n2965 ) | ( n2964 & n2965 ) ;
  assign n2967 = ~n2861 & n2864 ;
  assign n2968 = ( ~n2861 & n2866 ) | ( ~n2861 & n2967 ) | ( n2866 & n2967 ) ;
  assign n2969 = ( n2861 & n2868 ) | ( n2861 & ~n2967 ) | ( n2868 & ~n2967 ) ;
  assign n2970 = ( n2829 & n2968 ) | ( n2829 & ~n2969 ) | ( n2968 & ~n2969 ) ;
  assign n2971 = ( n2267 & n2966 ) | ( n2267 & ~n2970 ) | ( n2966 & ~n2970 ) ;
  assign n2972 = ( n2276 & ~n2966 ) | ( n2276 & n2970 ) | ( ~n2966 & n2970 ) ;
  assign n2973 = ( n2274 & n2971 ) | ( n2274 & ~n2972 ) | ( n2971 & ~n2972 ) ;
  assign n2974 = ( n2264 & ~n2966 ) | ( n2264 & n2970 ) | ( ~n2966 & n2970 ) ;
  assign n2975 = ( n2040 & ~n2971 ) | ( n2040 & n2974 ) | ( ~n2971 & n2974 ) ;
  assign n2976 = ( n1736 & ~n2973 ) | ( n1736 & n2975 ) | ( ~n2973 & n2975 ) ;
  assign n2977 = ~n2839 & n2856 ;
  assign n2978 = ( ~n2841 & n2856 ) | ( ~n2841 & n2977 ) | ( n2856 & n2977 ) ;
  assign n2979 = ( n2842 & n2844 ) | ( n2842 & ~n2978 ) | ( n2844 & ~n2978 ) ;
  assign n2980 = n879 & n1045 ;
  assign n2981 = ( n879 & ~n1040 ) | ( n879 & n2980 ) | ( ~n1040 & n2980 ) ;
  assign n2982 = ~n1042 & n2981 ;
  assign n2983 = n879 | n1045 ;
  assign n2984 = ( n879 & ~n1049 ) | ( n879 & n2983 ) | ( ~n1049 & n2983 ) ;
  assign n2985 = n1052 & n2984 ;
  assign n2986 = ( ~n1042 & n2984 ) | ( ~n1042 & n2985 ) | ( n2984 & n2985 ) ;
  assign n2987 = ~n2982 & n2986 ;
  assign n2988 = n304 & n942 ;
  assign n2989 = ( n922 & n942 ) | ( n922 & n2988 ) | ( n942 & n2988 ) ;
  assign n2990 = ( ~n900 & n921 ) | ( ~n900 & n2989 ) | ( n921 & n2989 ) ;
  assign n2991 = ( n900 & n942 ) | ( n900 & n2990 ) | ( n942 & n2990 ) ;
  assign n2992 = ~n2987 & n2991 ;
  assign n2993 = ( ~n754 & n2387 ) | ( ~n754 & n2853 ) | ( n2387 & n2853 ) ;
  assign n2994 = n2387 | n2853 ;
  assign n2995 = ( n757 & n2993 ) | ( n757 & n2994 ) | ( n2993 & n2994 ) ;
  assign n2996 = n2991 & n2995 ;
  assign n2997 = ( ~n2987 & n2995 ) | ( ~n2987 & n2996 ) | ( n2995 & n2996 ) ;
  assign n2998 = ( n2987 & ~n2991 ) | ( n2987 & n2997 ) | ( ~n2991 & n2997 ) ;
  assign n2999 = n2992 | n2998 ;
  assign n3000 = ~n2987 & n2996 ;
  assign n3001 = ( n2995 & ~n2997 ) | ( n2995 & n3000 ) | ( ~n2997 & n3000 ) ;
  assign n3002 = n2999 & ~n3001 ;
  assign n3003 = n2978 & n3002 ;
  assign n3004 = ~n2842 & n3002 ;
  assign n3005 = ( ~n2844 & n3003 ) | ( ~n2844 & n3004 ) | ( n3003 & n3004 ) ;
  assign n3006 = n3002 & ~n3005 ;
  assign n3007 = ( n2979 & n3005 ) | ( n2979 & ~n3006 ) | ( n3005 & ~n3006 ) ;
  assign n3008 = n2975 & ~n3007 ;
  assign n3009 = n2973 | n3007 ;
  assign n3010 = ( n1736 & n3008 ) | ( n1736 & ~n3009 ) | ( n3008 & ~n3009 ) ;
  assign n3011 = n2973 & ~n3007 ;
  assign n3012 = n2975 | n3007 ;
  assign n3013 = ( n1736 & ~n3011 ) | ( n1736 & n3012 ) | ( ~n3011 & n3012 ) ;
  assign n3014 = ( ~n2976 & n3010 ) | ( ~n2976 & n3013 ) | ( n3010 & n3013 ) ;
  assign n3015 = n2959 & ~n3014 ;
  assign n3016 = ~n2959 & n3014 ;
  assign n3017 = n3015 | n3016 ;
  assign n3018 = n2921 | n3017 ;
  assign n3019 = n2930 & ~n3017 ;
  assign n3020 = ( n2828 & ~n3018 ) | ( n2828 & n3019 ) | ( ~n3018 & n3019 ) ;
  assign n3021 = n2930 | n3017 ;
  assign n3022 = n2921 & ~n3017 ;
  assign n3023 = ( n2828 & n3021 ) | ( n2828 & ~n3022 ) | ( n3021 & ~n3022 ) ;
  assign n3024 = ( ~n2931 & n3020 ) | ( ~n2931 & n3023 ) | ( n3020 & n3023 ) ;
  assign n3025 = n2928 & n3024 ;
  assign n3026 = n2928 | n3024 ;
  assign n3027 = ~n3025 & n3026 ;
  assign n3028 = n2568 & n2622 ;
  assign n3029 = n2568 & n2625 ;
  assign n3030 = ( n2373 & n3028 ) | ( n2373 & n3029 ) | ( n3028 & n3029 ) ;
  assign n3031 = ( ~n2680 & n3028 ) | ( ~n2680 & n3029 ) | ( n3028 & n3029 ) ;
  assign n3032 = ( n2827 & n3030 ) | ( n2827 & n3031 ) | ( n3030 & n3031 ) ;
  assign n3033 = n2828 & ~n3032 ;
  assign n3036 = n2923 & n3033 ;
  assign n3037 = ( n2927 & n3033 ) | ( n2927 & n3036 ) | ( n3033 & n3036 ) ;
  assign n3034 = n2923 | n3033 ;
  assign n3035 = n2927 | n3034 ;
  assign n3038 = n3035 & ~n3037 ;
  assign n3039 = n3037 | n3038 ;
  assign n3040 = n3027 & n3039 ;
  assign n3041 = n3025 | n3040 ;
  assign n3042 = ( n2372 & ~n2679 ) | ( n2372 & n2683 ) | ( ~n2679 & n2683 ) ;
  assign n3043 = ~n2372 & n2679 ;
  assign n3044 = ( n2826 & n3042 ) | ( n2826 & ~n3043 ) | ( n3042 & ~n3043 ) ;
  assign n3045 = n2328 & ~n3044 ;
  assign n3046 = n2328 | n2680 ;
  assign n3047 = ~n2328 & n2373 ;
  assign n3048 = ( n2827 & ~n3046 ) | ( n2827 & n3047 ) | ( ~n3046 & n3047 ) ;
  assign n3049 = n3045 | n3048 ;
  assign n3050 = n2370 | n2679 ;
  assign n3051 = n2827 & ~n3050 ;
  assign n3052 = ~n2676 & n2683 ;
  assign n3053 = ( ~n2676 & n2826 ) | ( ~n2676 & n3052 ) | ( n2826 & n3052 ) ;
  assign n3054 = n2370 & n2676 ;
  assign n3055 = ( n2370 & ~n2683 ) | ( n2370 & n3054 ) | ( ~n2683 & n3054 ) ;
  assign n3056 = ( ~n2826 & n3054 ) | ( ~n2826 & n3055 ) | ( n3054 & n3055 ) ;
  assign n3057 = ( n2369 & ~n3053 ) | ( n2369 & n3056 ) | ( ~n3053 & n3056 ) ;
  assign n3058 = n3051 | n3057 ;
  assign n3059 = n3049 & n3058 ;
  assign n3060 = n3049 | n3058 ;
  assign n3061 = ~n3059 & n3060 ;
  assign n3062 = n2683 & n2826 ;
  assign n3063 = n2827 & ~n3062 ;
  assign n3064 = n3051 | n3063 ;
  assign n3065 = n3057 | n3064 ;
  assign n3066 = n3058 & n3063 ;
  assign n3067 = n3065 & ~n3066 ;
  assign n3068 = n2719 | n2825 ;
  assign n3069 = n2719 & n2825 ;
  assign n3070 = n3068 & ~n3069 ;
  assign n3071 = ~n2763 & n2825 ;
  assign n3072 = n2764 | n2823 ;
  assign n3073 = ~n3071 & n3072 ;
  assign n3074 = n3070 & ~n3073 ;
  assign n3075 = ~n3070 & n3073 ;
  assign n3076 = n3074 | n3075 ;
  assign n3077 = n2769 & ~n2796 ;
  assign n3078 = n2823 & ~n3077 ;
  assign n3079 = ~n2769 & n2796 ;
  assign n3080 = n2822 | n3079 ;
  assign n3081 = ~n2822 & n3077 ;
  assign n3082 = ( ~n2822 & n3080 ) | ( ~n2822 & n3081 ) | ( n3080 & n3081 ) ;
  assign n3083 = n3078 | n3082 ;
  assign n3084 = n2818 & ~n2821 ;
  assign n3085 = n2822 | n3084 ;
  assign n3086 = n3078 & n3085 ;
  assign n3087 = ( n3082 & n3085 ) | ( n3082 & n3086 ) | ( n3085 & n3086 ) ;
  assign n3088 = ( ~n3073 & n3083 ) | ( ~n3073 & n3087 ) | ( n3083 & n3087 ) ;
  assign n3089 = ~n3076 & n3088 ;
  assign n3090 = n3063 & n3070 ;
  assign n3091 = n3063 | n3070 ;
  assign n3092 = ~n3090 & n3091 ;
  assign n3093 = n3074 & n3092 ;
  assign n3094 = ( n3089 & n3092 ) | ( n3089 & n3093 ) | ( n3092 & n3093 ) ;
  assign n3095 = n3067 & n3090 ;
  assign n3096 = ( n3067 & n3094 ) | ( n3067 & n3095 ) | ( n3094 & n3095 ) ;
  assign n3097 = n3061 & n3066 ;
  assign n3098 = ( n3061 & n3096 ) | ( n3061 & n3097 ) | ( n3096 & n3097 ) ;
  assign n3099 = n2619 & ~n2620 ;
  assign n3100 = ( ~n2373 & n2624 ) | ( ~n2373 & n3099 ) | ( n2624 & n3099 ) ;
  assign n3101 = ( n2624 & n2680 ) | ( n2624 & n3099 ) | ( n2680 & n3099 ) ;
  assign n3102 = ( ~n2827 & n3100 ) | ( ~n2827 & n3101 ) | ( n3100 & n3101 ) ;
  assign n3103 = n2325 | n2680 ;
  assign n3104 = ~n2325 & n2373 ;
  assign n3105 = ( n2827 & ~n3103 ) | ( n2827 & n3104 ) | ( ~n3103 & n3104 ) ;
  assign n3106 = n3102 | n3105 ;
  assign n3107 = ~n2620 & n2622 ;
  assign n3108 = ~n2680 & n3107 ;
  assign n3109 = n2373 & n3107 ;
  assign n3110 = ( n2827 & n3108 ) | ( n2827 & n3109 ) | ( n3108 & n3109 ) ;
  assign n3111 = n3106 & ~n3110 ;
  assign n3112 = n3049 & ~n3111 ;
  assign n3113 = ~n3049 & n3111 ;
  assign n3114 = n3112 | n3113 ;
  assign n3115 = n3059 & ~n3114 ;
  assign n3116 = n3033 & ~n3111 ;
  assign n3117 = ~n3033 & n3111 ;
  assign n3118 = n3116 | n3117 ;
  assign n3119 = ~n3116 & n3118 ;
  assign n3120 = n3112 | n3116 ;
  assign n3121 = ( n3116 & ~n3118 ) | ( n3116 & n3120 ) | ( ~n3118 & n3120 ) ;
  assign n3122 = ( n3115 & ~n3119 ) | ( n3115 & n3121 ) | ( ~n3119 & n3121 ) ;
  assign n3123 = ( n3114 & n3119 ) | ( n3114 & ~n3121 ) | ( n3119 & ~n3121 ) ;
  assign n3124 = ( n3098 & n3122 ) | ( n3098 & ~n3123 ) | ( n3122 & ~n3123 ) ;
  assign n3125 = n3025 | n3037 ;
  assign n3126 = ( n3025 & n3027 ) | ( n3025 & n3125 ) | ( n3027 & n3125 ) ;
  assign n3127 = ( n3041 & n3124 ) | ( n3041 & n3126 ) | ( n3124 & n3126 ) ;
  assign n3128 = ~n3015 & n3017 ;
  assign n3129 = ( n2930 & ~n3015 ) | ( n2930 & n3128 ) | ( ~n3015 & n3128 ) ;
  assign n3130 = n2978 | n3002 ;
  assign n3131 = n2842 & ~n3002 ;
  assign n3132 = ( n2844 & ~n3130 ) | ( n2844 & n3131 ) | ( ~n3130 & n3131 ) ;
  assign n3133 = ~n2998 & n3132 ;
  assign n3134 = ( n2998 & n3007 ) | ( n2998 & ~n3133 ) | ( n3007 & ~n3133 ) ;
  assign n3135 = ( n2970 & ~n3133 ) | ( n2970 & n3134 ) | ( ~n3133 & n3134 ) ;
  assign n3136 = ( n2966 & n3133 ) | ( n2966 & ~n3134 ) | ( n3133 & ~n3134 ) ;
  assign n3137 = ( n2267 & ~n3135 ) | ( n2267 & n3136 ) | ( ~n3135 & n3136 ) ;
  assign n3138 = ( n2276 & n3135 ) | ( n2276 & ~n3136 ) | ( n3135 & ~n3136 ) ;
  assign n3139 = ( n2274 & n3137 ) | ( n2274 & ~n3138 ) | ( n3137 & ~n3138 ) ;
  assign n3140 = ( n2264 & n3135 ) | ( n2264 & ~n3136 ) | ( n3135 & ~n3136 ) ;
  assign n3141 = ( n2040 & ~n3137 ) | ( n2040 & n3140 ) | ( ~n3137 & n3140 ) ;
  assign n3142 = ( n1736 & ~n3139 ) | ( n1736 & n3141 ) | ( ~n3139 & n3141 ) ;
  assign n3143 = n2998 & ~n3132 ;
  assign n3144 = n3007 & n3143 ;
  assign n3145 = ( n2970 & n3143 ) | ( n2970 & n3144 ) | ( n3143 & n3144 ) ;
  assign n3146 = ( ~n2966 & n3143 ) | ( ~n2966 & n3144 ) | ( n3143 & n3144 ) ;
  assign n3147 = ( ~n2267 & n3145 ) | ( ~n2267 & n3146 ) | ( n3145 & n3146 ) ;
  assign n3148 = ( n2276 & n3145 ) | ( n2276 & n3146 ) | ( n3145 & n3146 ) ;
  assign n3149 = ( ~n2274 & n3147 ) | ( ~n2274 & n3148 ) | ( n3147 & n3148 ) ;
  assign n3150 = ( n2264 & n3145 ) | ( n2264 & n3146 ) | ( n3145 & n3146 ) ;
  assign n3151 = ( n2040 & n3147 ) | ( n2040 & n3150 ) | ( n3147 & n3150 ) ;
  assign n3152 = ( n1736 & n3149 ) | ( n1736 & n3151 ) | ( n3149 & n3151 ) ;
  assign n3153 = n3142 & ~n3152 ;
  assign n3154 = ( n754 & n1029 ) | ( n754 & n1038 ) | ( n1029 & n1038 ) ;
  assign n3155 = n879 & ~n942 ;
  assign n3156 = ~n879 & n942 ;
  assign n3157 = n3155 | n3156 ;
  assign n3158 = ( n754 & ~n3154 ) | ( n754 & n3157 ) | ( ~n3154 & n3157 ) ;
  assign n3159 = n3154 & n3158 ;
  assign n3160 = n1045 & ~n3157 ;
  assign n3161 = n753 & ~n3157 ;
  assign n3162 = ( n736 & ~n3157 ) | ( n736 & n3161 ) | ( ~n3157 & n3161 ) ;
  assign n3163 = n1045 & ~n3162 ;
  assign n3164 = ( n1045 & ~n3154 ) | ( n1045 & n3163 ) | ( ~n3154 & n3163 ) ;
  assign n3165 = ( n3159 & n3160 ) | ( n3159 & n3164 ) | ( n3160 & n3164 ) ;
  assign n3166 = n3153 & n3165 ;
  assign n3167 = n3153 | n3165 ;
  assign n3168 = ~n3166 & n3167 ;
  assign n3194 = n210 | n426 ;
  assign n3195 = n361 | n3194 ;
  assign n3196 = n177 | n283 ;
  assign n3197 = n452 | n3196 ;
  assign n3198 = n134 | n269 ;
  assign n3199 = n349 | n3198 ;
  assign n3200 = n3197 | n3199 ;
  assign n3201 = n260 | n3200 ;
  assign n3202 = n737 | n823 ;
  assign n3203 = n2346 | n3202 ;
  assign n3204 = n3201 | n3203 ;
  assign n3205 = n372 | n844 ;
  assign n3206 = n835 | n3205 ;
  assign n3207 = n833 | n3206 ;
  assign n3208 = n174 | n685 ;
  assign n3209 = n317 | n3208 ;
  assign n3210 = n684 | n3209 ;
  assign n3211 = n368 | n502 ;
  assign n3212 = n3210 | n3211 ;
  assign n3213 = n3207 | n3212 ;
  assign n3214 = n3204 | n3213 ;
  assign n3215 = n3195 | n3214 ;
  assign n3169 = n724 | n2648 ;
  assign n3170 = n2644 | n3169 ;
  assign n3171 = n177 | n216 ;
  assign n3172 = n320 | n366 ;
  assign n3173 = n3171 | n3172 ;
  assign n3174 = n495 | n3173 ;
  assign n3175 = n176 | n315 ;
  assign n3176 = n270 | n290 ;
  assign n3177 = n3175 | n3176 ;
  assign n3178 = n677 | n3177 ;
  assign n3179 = n3174 | n3178 ;
  assign n3180 = n524 | n570 ;
  assign n3181 = n2546 | n3180 ;
  assign n3182 = n206 | n305 ;
  assign n3183 = n510 & ~n3182 ;
  assign n3184 = ~n3181 & n3183 ;
  assign n3185 = ~n3179 & n3184 ;
  assign n3186 = ~n3170 & n3185 ;
  assign n3187 = n547 | n806 ;
  assign n3188 = n348 | n429 ;
  assign n3189 = n3187 | n3188 ;
  assign n3190 = n3186 & ~n3189 ;
  assign n3216 = n3190 & ~n3215 ;
  assign n3217 = ( n3168 & ~n3215 ) | ( n3168 & n3216 ) | ( ~n3215 & n3216 ) ;
  assign n3191 = n3168 | n3190 ;
  assign n3192 = n3168 & n3190 ;
  assign n3193 = n3191 & ~n3192 ;
  assign n3218 = ~n3193 & n3217 ;
  assign n3219 = ( n3129 & n3217 ) | ( n3129 & n3218 ) | ( n3217 & n3218 ) ;
  assign n3220 = ( n2921 & n3015 ) | ( n2921 & ~n3128 ) | ( n3015 & ~n3128 ) ;
  assign n3221 = ( n3217 & n3218 ) | ( n3217 & ~n3220 ) | ( n3218 & ~n3220 ) ;
  assign n3222 = ( n2828 & n3219 ) | ( n2828 & n3221 ) | ( n3219 & n3221 ) ;
  assign n3223 = n548 | n709 ;
  assign n3224 = n330 | n3223 ;
  assign n3225 = n392 | n2652 ;
  assign n3226 = n226 | n3225 ;
  assign n3227 = n213 | n3226 ;
  assign n3228 = n181 | n3227 ;
  assign n3229 = n343 | n387 ;
  assign n3230 = n283 | n3229 ;
  assign n3231 = n429 | n538 ;
  assign n3232 = n245 | n290 ;
  assign n3233 = n3231 | n3232 ;
  assign n3234 = n3230 | n3233 ;
  assign n3235 = n357 | n3234 ;
  assign n3236 = n293 | n334 ;
  assign n3237 = n228 | n443 ;
  assign n3238 = n3236 | n3237 ;
  assign n3239 = n501 | n3238 ;
  assign n3240 = n191 | n305 ;
  assign n3241 = n322 | n3240 ;
  assign n3242 = n2555 | n3241 ;
  assign n3243 = n3239 | n3242 ;
  assign n3244 = n253 | n267 ;
  assign n3245 = n352 | n689 ;
  assign n3246 = n3244 | n3245 ;
  assign n3247 = n202 | n3246 ;
  assign n3248 = n408 | n495 ;
  assign n3249 = n249 | n338 ;
  assign n3250 = n3248 | n3249 ;
  assign n3251 = n511 | n3250 ;
  assign n3252 = n3247 | n3251 ;
  assign n3253 = n3243 | n3252 ;
  assign n3254 = n3235 | n3253 ;
  assign n3255 = n3228 | n3254 ;
  assign n3256 = n3224 | n3255 ;
  assign n3257 = n3222 | n3256 ;
  assign n3258 = n3222 & n3256 ;
  assign n3259 = n3257 & ~n3258 ;
  assign n3260 = ~n3190 & n3215 ;
  assign n3261 = ~n3168 & n3260 ;
  assign n3262 = ( n3193 & n3215 ) | ( n3193 & n3261 ) | ( n3215 & n3261 ) ;
  assign n3263 = ( ~n3129 & n3261 ) | ( ~n3129 & n3262 ) | ( n3261 & n3262 ) ;
  assign n3264 = ( n3220 & n3261 ) | ( n3220 & n3262 ) | ( n3261 & n3262 ) ;
  assign n3265 = ( ~n2828 & n3263 ) | ( ~n2828 & n3264 ) | ( n3263 & n3264 ) ;
  assign n3266 = n3222 | n3265 ;
  assign n3267 = n3259 & n3266 ;
  assign n3268 = n3259 | n3266 ;
  assign n3269 = ~n3267 & n3268 ;
  assign n3270 = n3267 | n3269 ;
  assign n3271 = n134 | n315 ;
  assign n3272 = n125 | n3271 ;
  assign n3273 = ~n312 & n509 ;
  assign n3274 = ~n746 & n3273 ;
  assign n3275 = ~n2528 & n3274 ;
  assign n3276 = ~n743 & n3275 ;
  assign n3277 = n242 | n244 ;
  assign n3278 = n582 | n3277 ;
  assign n3279 = n2359 | n2733 ;
  assign n3280 = n2361 | n3279 ;
  assign n3281 = n3278 | n3280 ;
  assign n3282 = n3276 & ~n3281 ;
  assign n3283 = ~n900 & n3282 ;
  assign n3284 = ~n3272 & n3283 ;
  assign n3285 = ~n3256 & n3284 ;
  assign n3286 = n3222 & n3285 ;
  assign n3287 = n3256 & ~n3284 ;
  assign n3288 = ( n3222 & n3284 ) | ( n3222 & ~n3287 ) | ( n3284 & ~n3287 ) ;
  assign n3289 = ~n3286 & n3288 ;
  assign n3290 = n3259 & ~n3289 ;
  assign n3291 = ~n3259 & n3289 ;
  assign n3292 = n3290 | n3291 ;
  assign n3293 = n3270 & ~n3292 ;
  assign n3294 = n3267 & ~n3292 ;
  assign n3295 = n3129 & n3193 ;
  assign n3296 = n3193 & ~n3220 ;
  assign n3297 = ( n2828 & n3295 ) | ( n2828 & n3296 ) | ( n3295 & n3296 ) ;
  assign n3298 = ~n3193 & n3220 ;
  assign n3299 = n3129 | n3193 ;
  assign n3300 = ( n2828 & ~n3298 ) | ( n2828 & n3299 ) | ( ~n3298 & n3299 ) ;
  assign n3301 = ~n3297 & n3300 ;
  assign n3302 = n3266 & ~n3301 ;
  assign n3303 = n3024 & ~n3301 ;
  assign n3304 = ~n3024 & n3301 ;
  assign n3305 = n3303 | n3304 ;
  assign n3306 = ~n3303 & n3305 ;
  assign n3307 = ~n3266 & n3301 ;
  assign n3308 = n3302 | n3307 ;
  assign n3309 = ~n3302 & n3308 ;
  assign n3310 = ( ~n3302 & n3306 ) | ( ~n3302 & n3309 ) | ( n3306 & n3309 ) ;
  assign n3311 = ( n3293 & n3294 ) | ( n3293 & ~n3310 ) | ( n3294 & ~n3310 ) ;
  assign n3312 = n3302 | n3303 ;
  assign n3313 = ( n3302 & ~n3308 ) | ( n3302 & n3312 ) | ( ~n3308 & n3312 ) ;
  assign n3314 = ( n3293 & n3294 ) | ( n3293 & n3313 ) | ( n3294 & n3313 ) ;
  assign n3315 = ( n3127 & n3311 ) | ( n3127 & n3314 ) | ( n3311 & n3314 ) ;
  assign n3316 = ~n3270 & n3292 ;
  assign n3317 = ~n3267 & n3292 ;
  assign n3318 = ( n3310 & n3316 ) | ( n3310 & n3317 ) | ( n3316 & n3317 ) ;
  assign n3319 = ( ~n3313 & n3316 ) | ( ~n3313 & n3317 ) | ( n3316 & n3317 ) ;
  assign n3320 = ( ~n3127 & n3318 ) | ( ~n3127 & n3319 ) | ( n3318 & n3319 ) ;
  assign n3321 = n3315 | n3320 ;
  assign n3322 = x2 & x22 ;
  assign n3323 = x0 | x1 ;
  assign n3324 = x2 & n3323 ;
  assign n3325 = n902 & ~n3324 ;
  assign n3326 = n3322 | n3325 ;
  assign n3327 = x1 & ~n901 ;
  assign n3328 = ~x1 & n901 ;
  assign n3329 = n3327 | n3328 ;
  assign n3330 = n3326 & ~n3329 ;
  assign n3331 = ~n3326 & n3329 ;
  assign n3332 = n3330 | n3331 ;
  assign n3333 = ~n3323 & n3332 ;
  assign n3334 = n3266 & n3333 ;
  assign n3335 = ~x0 & n3329 ;
  assign n3336 = n3259 & n3335 ;
  assign n3337 = n3334 | n3336 ;
  assign n3338 = x0 & ~n3332 ;
  assign n3339 = ~n3289 & n3338 ;
  assign n3340 = x0 & n3332 ;
  assign n3341 = n3338 | n3340 ;
  assign n3342 = ( ~n3289 & n3340 ) | ( ~n3289 & n3341 ) | ( n3340 & n3341 ) ;
  assign n3343 = n3339 & n3342 ;
  assign n3344 = n3337 | n3343 ;
  assign n3345 = n3326 | n3344 ;
  assign n3346 = n3326 | n3341 ;
  assign n3347 = n3326 | n3340 ;
  assign n3348 = ( ~n3289 & n3346 ) | ( ~n3289 & n3347 ) | ( n3346 & n3347 ) ;
  assign n3349 = n3337 | n3348 ;
  assign n3350 = ( ~n3321 & n3345 ) | ( ~n3321 & n3349 ) | ( n3345 & n3349 ) ;
  assign n3351 = n3326 & n3344 ;
  assign n3352 = n3326 & n3341 ;
  assign n3353 = n3326 & n3340 ;
  assign n3354 = ( ~n3289 & n3352 ) | ( ~n3289 & n3353 ) | ( n3352 & n3353 ) ;
  assign n3355 = ( n3326 & n3337 ) | ( n3326 & n3354 ) | ( n3337 & n3354 ) ;
  assign n3356 = ( ~n3321 & n3351 ) | ( ~n3321 & n3355 ) | ( n3351 & n3355 ) ;
  assign n3357 = n3350 & ~n3356 ;
  assign n3358 = n3127 & ~n3305 ;
  assign n3359 = ~n3127 & n3305 ;
  assign n3360 = n3358 | n3359 ;
  assign n3361 = ~n905 & n3326 ;
  assign n3362 = n905 & ~n3326 ;
  assign n3363 = n3361 | n3362 ;
  assign n3364 = ~n905 & n1094 ;
  assign n3365 = n905 & ~n1094 ;
  assign n3366 = n3364 | n3365 ;
  assign n3367 = ~n3363 & n3366 ;
  assign n3368 = n3024 & n3367 ;
  assign n3369 = n1094 & ~n1115 ;
  assign n3370 = ~n1094 & n1115 ;
  assign n3371 = n3369 | n3370 ;
  assign n3372 = n3363 | n3366 ;
  assign n3373 = n3371 & ~n3372 ;
  assign n3374 = n2916 & n3373 ;
  assign n3375 = ( ~n2901 & n3373 ) | ( ~n2901 & n3374 ) | ( n3373 & n3374 ) ;
  assign n3376 = ~n2921 & n3375 ;
  assign n3377 = n2828 & n3376 ;
  assign n3378 = ( n2927 & n3373 ) | ( n2927 & n3377 ) | ( n3373 & n3377 ) ;
  assign n3379 = n3368 | n3378 ;
  assign n3380 = n3363 & ~n3371 ;
  assign n3381 = n3296 & n3380 ;
  assign n3382 = n3295 & n3380 ;
  assign n3383 = ( n2828 & n3381 ) | ( n2828 & n3382 ) | ( n3381 & n3382 ) ;
  assign n3384 = ( ~n3300 & n3380 ) | ( ~n3300 & n3383 ) | ( n3380 & n3383 ) ;
  assign n3385 = n1115 & n3384 ;
  assign n3386 = ( n1115 & n3379 ) | ( n1115 & n3385 ) | ( n3379 & n3385 ) ;
  assign n3387 = n3363 & n3371 ;
  assign n3388 = n1115 & n3387 ;
  assign n3389 = ( n1115 & n3384 ) | ( n1115 & n3388 ) | ( n3384 & n3388 ) ;
  assign n3390 = ( n1115 & n3379 ) | ( n1115 & n3389 ) | ( n3379 & n3389 ) ;
  assign n3391 = ( ~n3360 & n3386 ) | ( ~n3360 & n3390 ) | ( n3386 & n3390 ) ;
  assign n3392 = n1115 | n3384 ;
  assign n3393 = n3379 | n3392 ;
  assign n3394 = n1115 | n3387 ;
  assign n3395 = n3384 | n3394 ;
  assign n3396 = n3379 | n3395 ;
  assign n3397 = ( ~n3360 & n3393 ) | ( ~n3360 & n3396 ) | ( n3393 & n3396 ) ;
  assign n3398 = ~n3391 & n3397 ;
  assign n3399 = n3067 | n3090 ;
  assign n3400 = n3094 | n3399 ;
  assign n3401 = ~n3096 & n3400 ;
  assign n3402 = ~n473 & n482 ;
  assign n3403 = n473 & ~n482 ;
  assign n3404 = n3402 | n3403 ;
  assign n3405 = ~n634 & n642 ;
  assign n3406 = n634 & ~n642 ;
  assign n3407 = n3405 | n3406 ;
  assign n3408 = ~n473 & n642 ;
  assign n3409 = n473 & ~n642 ;
  assign n3410 = n3408 | n3409 ;
  assign n3411 = n3407 & ~n3410 ;
  assign n3412 = ~n3404 & n3411 ;
  assign n3413 = n3070 & n3412 ;
  assign n3414 = ~n3404 & n3410 ;
  assign n3415 = n3063 & n3414 ;
  assign n3416 = n3413 | n3415 ;
  assign n3417 = n3404 & ~n3407 ;
  assign n3418 = n2368 & n3417 ;
  assign n3419 = ( ~n2340 & n3417 ) | ( ~n2340 & n3418 ) | ( n3417 & n3418 ) ;
  assign n3420 = ~n2679 & n3419 ;
  assign n3421 = n2827 & n3420 ;
  assign n3422 = ( n3057 & n3417 ) | ( n3057 & n3421 ) | ( n3417 & n3421 ) ;
  assign n3423 = n3404 & n3407 ;
  assign n3424 = n634 & n3423 ;
  assign n3425 = ( n634 & n3422 ) | ( n634 & n3424 ) | ( n3422 & n3424 ) ;
  assign n3426 = n634 | n3424 ;
  assign n3427 = ( n3416 & n3425 ) | ( n3416 & n3426 ) | ( n3425 & n3426 ) ;
  assign n3428 = n634 & n3422 ;
  assign n3429 = ( n634 & n3416 ) | ( n634 & n3428 ) | ( n3416 & n3428 ) ;
  assign n3430 = ( n3401 & n3427 ) | ( n3401 & n3429 ) | ( n3427 & n3429 ) ;
  assign n3431 = n634 | n3423 ;
  assign n3432 = n3422 | n3431 ;
  assign n3433 = n3416 | n3432 ;
  assign n3434 = n634 | n3422 ;
  assign n3435 = n3416 | n3434 ;
  assign n3436 = ( n3401 & n3433 ) | ( n3401 & n3435 ) | ( n3433 & n3435 ) ;
  assign n3437 = ~n3430 & n3436 ;
  assign n3438 = ~n634 & n1004 ;
  assign n3439 = n634 & ~n1004 ;
  assign n3440 = n3438 | n3439 ;
  assign n3441 = ~n942 & n997 ;
  assign n3442 = ( ~n942 & n1003 ) | ( ~n942 & n3441 ) | ( n1003 & n3441 ) ;
  assign n3443 = n942 & ~n997 ;
  assign n3444 = ~n1003 & n3443 ;
  assign n3445 = n3442 | n3444 ;
  assign n3446 = ~n3440 & n3445 ;
  assign n3447 = n3085 & n3446 ;
  assign n3448 = ~n3157 & n3440 ;
  assign n3449 = n3078 & n3448 ;
  assign n3450 = ( n3082 & n3448 ) | ( n3082 & n3449 ) | ( n3448 & n3449 ) ;
  assign n3451 = n3447 | n3450 ;
  assign n3452 = n3157 & n3440 ;
  assign n3453 = ~n3078 & n3085 ;
  assign n3454 = ~n3082 & n3453 ;
  assign n3455 = n3078 & ~n3085 ;
  assign n3456 = ( n3082 & ~n3085 ) | ( n3082 & n3455 ) | ( ~n3085 & n3455 ) ;
  assign n3457 = n3454 | n3456 ;
  assign n3458 = n3452 & n3457 ;
  assign n3459 = n3451 | n3458 ;
  assign n3460 = n879 & n3446 ;
  assign n3461 = n3085 & n3460 ;
  assign n3462 = ( n879 & n3450 ) | ( n879 & n3461 ) | ( n3450 & n3461 ) ;
  assign n3463 = ( n879 & n3458 ) | ( n879 & n3462 ) | ( n3458 & n3462 ) ;
  assign n3464 = n3459 & ~n3463 ;
  assign n3465 = n879 & ~n3440 ;
  assign n3466 = ( n879 & ~n3085 ) | ( n879 & n3465 ) | ( ~n3085 & n3465 ) ;
  assign n3467 = n879 & ~n3460 ;
  assign n3468 = ( n879 & ~n3085 ) | ( n879 & n3467 ) | ( ~n3085 & n3467 ) ;
  assign n3469 = n3466 & n3468 ;
  assign n3470 = ~n3450 & n3469 ;
  assign n3471 = ~n3458 & n3470 ;
  assign n3472 = ( n3464 & n3466 ) | ( n3464 & n3471 ) | ( n3466 & n3471 ) ;
  assign n3473 = n3073 & ~n3456 ;
  assign n3474 = ~n3073 & n3456 ;
  assign n3475 = n3473 | n3474 ;
  assign n3482 = ~n2823 & n3448 ;
  assign n3483 = ~n2764 & n3482 ;
  assign n3484 = ( n3071 & n3448 ) | ( n3071 & n3483 ) | ( n3448 & n3483 ) ;
  assign n3476 = n3157 & ~n3445 ;
  assign n3477 = ~n3440 & n3476 ;
  assign n3478 = n3085 & n3477 ;
  assign n3479 = n3078 & n3446 ;
  assign n3480 = ( n3082 & n3446 ) | ( n3082 & n3479 ) | ( n3446 & n3479 ) ;
  assign n3481 = n3478 | n3480 ;
  assign n3485 = n3481 | n3484 ;
  assign n3487 = n3452 | n3477 ;
  assign n3488 = ( n3085 & n3452 ) | ( n3085 & n3487 ) | ( n3452 & n3487 ) ;
  assign n3489 = n3480 | n3488 ;
  assign n3490 = ( n3484 & n3485 ) | ( n3484 & n3489 ) | ( n3485 & n3489 ) ;
  assign n3491 = n3484 | n3489 ;
  assign n3492 = ( ~n3475 & n3490 ) | ( ~n3475 & n3491 ) | ( n3490 & n3491 ) ;
  assign n3486 = n3475 & ~n3485 ;
  assign n3493 = ( ~n879 & n3486 ) | ( ~n879 & n3492 ) | ( n3486 & n3492 ) ;
  assign n3494 = n3492 & ~n3493 ;
  assign n3495 = ~n3486 & n3493 ;
  assign n3496 = ( n879 & ~n3494 ) | ( n879 & n3495 ) | ( ~n3494 & n3495 ) ;
  assign n3497 = n3472 & n3496 ;
  assign n3498 = n3472 | n3496 ;
  assign n3499 = ~n3497 & n3498 ;
  assign n3500 = n3437 & n3499 ;
  assign n3501 = n3437 | n3499 ;
  assign n3502 = ~n3500 & n3501 ;
  assign n3503 = n3466 | n3468 ;
  assign n3504 = ( ~n3450 & n3466 ) | ( ~n3450 & n3503 ) | ( n3466 & n3503 ) ;
  assign n3505 = ( ~n3458 & n3466 ) | ( ~n3458 & n3504 ) | ( n3466 & n3504 ) ;
  assign n3506 = n3464 | n3505 ;
  assign n3507 = ~n3472 & n3506 ;
  assign n3508 = n3074 | n3088 ;
  assign n3509 = ( n3074 & ~n3076 ) | ( n3074 & n3508 ) | ( ~n3076 & n3508 ) ;
  assign n3510 = n3092 | n3509 ;
  assign n3511 = n3063 & n3417 ;
  assign n3512 = n3070 & n3414 ;
  assign n3513 = ~n2823 & n3412 ;
  assign n3514 = ~n2764 & n3513 ;
  assign n3515 = n3423 | n3514 ;
  assign n3516 = n3412 | n3423 ;
  assign n3517 = ( n3071 & n3515 ) | ( n3071 & n3516 ) | ( n3515 & n3516 ) ;
  assign n3518 = n3512 | n3517 ;
  assign n3519 = n3511 | n3518 ;
  assign n3520 = n634 | n3519 ;
  assign n3521 = n3511 | n3512 ;
  assign n3522 = ( n3071 & n3412 ) | ( n3071 & n3514 ) | ( n3412 & n3514 ) ;
  assign n3523 = n3517 & n3522 ;
  assign n3524 = n634 | n3523 ;
  assign n3525 = n3521 | n3524 ;
  assign n3526 = ( n3510 & n3520 ) | ( n3510 & n3525 ) | ( n3520 & n3525 ) ;
  assign n3527 = n3520 & n3525 ;
  assign n3528 = ( ~n3094 & n3526 ) | ( ~n3094 & n3527 ) | ( n3526 & n3527 ) ;
  assign n3529 = n634 & n3519 ;
  assign n3530 = n634 & n3523 ;
  assign n3531 = ( n634 & n3521 ) | ( n634 & n3530 ) | ( n3521 & n3530 ) ;
  assign n3532 = ( n3510 & n3529 ) | ( n3510 & n3531 ) | ( n3529 & n3531 ) ;
  assign n3533 = n3529 & n3531 ;
  assign n3534 = ( ~n3094 & n3532 ) | ( ~n3094 & n3533 ) | ( n3532 & n3533 ) ;
  assign n3535 = n3528 & ~n3534 ;
  assign n3536 = n3507 & n3535 ;
  assign n3541 = ~n2823 & n3417 ;
  assign n3542 = ~n2764 & n3541 ;
  assign n3543 = ( n3071 & n3417 ) | ( n3071 & n3542 ) | ( n3417 & n3542 ) ;
  assign n3537 = n3085 & n3412 ;
  assign n3538 = n3078 & n3414 ;
  assign n3539 = ( n3082 & n3414 ) | ( n3082 & n3538 ) | ( n3414 & n3538 ) ;
  assign n3540 = n3537 | n3539 ;
  assign n3544 = n3540 | n3543 ;
  assign n3546 = ( n3085 & n3423 ) | ( n3085 & n3516 ) | ( n3423 & n3516 ) ;
  assign n3547 = n3539 | n3546 ;
  assign n3548 = ( n3543 & n3544 ) | ( n3543 & n3547 ) | ( n3544 & n3547 ) ;
  assign n3549 = n3543 | n3547 ;
  assign n3550 = ( ~n3475 & n3548 ) | ( ~n3475 & n3549 ) | ( n3548 & n3549 ) ;
  assign n3545 = n3475 & ~n3544 ;
  assign n3551 = ( ~n634 & n3545 ) | ( ~n634 & n3550 ) | ( n3545 & n3550 ) ;
  assign n3552 = n3550 & ~n3551 ;
  assign n3553 = ~n3545 & n3551 ;
  assign n3554 = ( n634 & ~n3552 ) | ( n634 & n3553 ) | ( ~n3552 & n3553 ) ;
  assign n3556 = n3414 | n3423 ;
  assign n3557 = ( n3085 & n3423 ) | ( n3085 & n3556 ) | ( n3423 & n3556 ) ;
  assign n3559 = n3078 & n3417 ;
  assign n3560 = ( n3082 & n3417 ) | ( n3082 & n3559 ) | ( n3417 & n3559 ) ;
  assign n3561 = ~n3557 & n3560 ;
  assign n3555 = n3085 & n3414 ;
  assign n3562 = ~n3555 & n3560 ;
  assign n3563 = ( ~n3457 & n3561 ) | ( ~n3457 & n3562 ) | ( n3561 & n3562 ) ;
  assign n3558 = ( n3457 & n3555 ) | ( n3457 & n3557 ) | ( n3555 & n3557 ) ;
  assign n3564 = ( n634 & ~n3558 ) | ( n634 & n3563 ) | ( ~n3558 & n3563 ) ;
  assign n3565 = ( n634 & n3563 ) | ( n634 & ~n3564 ) | ( n3563 & ~n3564 ) ;
  assign n3566 = n3085 & n3440 ;
  assign n3567 = n634 & ~n3404 ;
  assign n3568 = ( n634 & ~n3085 ) | ( n634 & n3567 ) | ( ~n3085 & n3567 ) ;
  assign n3569 = n3566 & n3568 ;
  assign n3570 = n3564 & n3569 ;
  assign n3571 = n3557 & n3569 ;
  assign n3572 = n3555 & n3569 ;
  assign n3573 = ( n3457 & n3571 ) | ( n3457 & n3572 ) | ( n3571 & n3572 ) ;
  assign n3574 = ( ~n3565 & n3570 ) | ( ~n3565 & n3573 ) | ( n3570 & n3573 ) ;
  assign n3575 = n3554 & n3574 ;
  assign n3576 = n3564 & n3568 ;
  assign n3577 = n3557 & n3568 ;
  assign n3578 = n3555 & n3568 ;
  assign n3579 = ( n3457 & n3577 ) | ( n3457 & n3578 ) | ( n3577 & n3578 ) ;
  assign n3580 = ( ~n3565 & n3576 ) | ( ~n3565 & n3579 ) | ( n3576 & n3579 ) ;
  assign n3581 = n3554 & n3580 ;
  assign n3582 = ~n3575 & n3581 ;
  assign n3583 = n3076 | n3089 ;
  assign n3584 = n3078 & n3412 ;
  assign n3585 = ( n3082 & n3412 ) | ( n3082 & n3584 ) | ( n3412 & n3584 ) ;
  assign n3586 = n3417 | n3585 ;
  assign n3587 = ( n3070 & n3585 ) | ( n3070 & n3586 ) | ( n3585 & n3586 ) ;
  assign n3588 = ~n2823 & n3414 ;
  assign n3589 = ~n2764 & n3588 ;
  assign n3590 = ( n3071 & n3414 ) | ( n3071 & n3589 ) | ( n3414 & n3589 ) ;
  assign n3591 = n3587 | n3590 ;
  assign n3592 = n3088 & n3424 ;
  assign n3593 = n3076 & n3592 ;
  assign n3594 = ( n634 & n3591 ) | ( n634 & n3593 ) | ( n3591 & n3593 ) ;
  assign n3595 = ( n634 & n3424 ) | ( n634 & n3591 ) | ( n3424 & n3591 ) ;
  assign n3596 = ( ~n3583 & n3594 ) | ( ~n3583 & n3595 ) | ( n3594 & n3595 ) ;
  assign n3597 = ( n634 & n3088 ) | ( n634 & n3431 ) | ( n3088 & n3431 ) ;
  assign n3598 = n634 & n3431 ;
  assign n3599 = ( n3076 & n3597 ) | ( n3076 & n3598 ) | ( n3597 & n3598 ) ;
  assign n3600 = n3591 | n3599 ;
  assign n3601 = n3431 | n3591 ;
  assign n3602 = ( ~n3583 & n3600 ) | ( ~n3583 & n3601 ) | ( n3600 & n3601 ) ;
  assign n3603 = ~n3596 & n3602 ;
  assign n3604 = n3566 & ~n3574 ;
  assign n3605 = ( ~n3554 & n3566 ) | ( ~n3554 & n3604 ) | ( n3566 & n3604 ) ;
  assign n3606 = n3603 & n3605 ;
  assign n3607 = ( n3582 & n3603 ) | ( n3582 & n3606 ) | ( n3603 & n3606 ) ;
  assign n3608 = n3575 | n3607 ;
  assign n3609 = n3507 | n3535 ;
  assign n3610 = ~n3536 & n3609 ;
  assign n3611 = n3536 | n3610 ;
  assign n3612 = ( n3536 & n3608 ) | ( n3536 & n3611 ) | ( n3608 & n3611 ) ;
  assign n3613 = n3502 & n3612 ;
  assign n3614 = n3502 | n3612 ;
  assign n3615 = ~n3613 & n3614 ;
  assign n3616 = n3112 & ~n3118 ;
  assign n3617 = ( n3115 & ~n3118 ) | ( n3115 & n3616 ) | ( ~n3118 & n3616 ) ;
  assign n3618 = ( n3114 & n3118 ) | ( n3114 & ~n3616 ) | ( n3118 & ~n3616 ) ;
  assign n3619 = ( n3098 & n3617 ) | ( n3098 & ~n3618 ) | ( n3617 & ~n3618 ) ;
  assign n3620 = ~n3112 & n3118 ;
  assign n3621 = ~n3115 & n3620 ;
  assign n3622 = n3114 & n3620 ;
  assign n3623 = ( ~n3098 & n3621 ) | ( ~n3098 & n3622 ) | ( n3621 & n3622 ) ;
  assign n3624 = n3619 | n3623 ;
  assign n3625 = n482 & ~n663 ;
  assign n3626 = ~n482 & n663 ;
  assign n3627 = n3625 | n3626 ;
  assign n3628 = n763 & ~n1115 ;
  assign n3629 = ~n763 & n1115 ;
  assign n3630 = n3628 | n3629 ;
  assign n3631 = ~n663 & n763 ;
  assign n3632 = n663 & ~n763 ;
  assign n3633 = n3631 | n3632 ;
  assign n3634 = n3630 | n3633 ;
  assign n3635 = n3627 & ~n3634 ;
  assign n3636 = n3049 & n3635 ;
  assign n3637 = ~n3630 & n3633 ;
  assign n3638 = n3110 & n3637 ;
  assign n3639 = ( ~n3106 & n3637 ) | ( ~n3106 & n3638 ) | ( n3637 & n3638 ) ;
  assign n3640 = n3636 | n3639 ;
  assign n3641 = ~n3627 & n3630 ;
  assign n3642 = n3033 & n3641 ;
  assign n3643 = n3627 & n3630 ;
  assign n3644 = n3641 | n3643 ;
  assign n3645 = ( n3033 & n3643 ) | ( n3033 & n3644 ) | ( n3643 & n3644 ) ;
  assign n3646 = n3642 & n3645 ;
  assign n3647 = n3640 | n3646 ;
  assign n3648 = n482 | n3647 ;
  assign n3649 = n482 | n3644 ;
  assign n3650 = n482 | n3643 ;
  assign n3651 = ( n3033 & n3649 ) | ( n3033 & n3650 ) | ( n3649 & n3650 ) ;
  assign n3652 = n3640 | n3651 ;
  assign n3653 = ( ~n3624 & n3648 ) | ( ~n3624 & n3652 ) | ( n3648 & n3652 ) ;
  assign n3654 = n482 & n3647 ;
  assign n3655 = n482 & n3630 ;
  assign n3656 = n3627 & n3655 ;
  assign n3657 = n482 & n3644 ;
  assign n3658 = ( n3033 & n3656 ) | ( n3033 & n3657 ) | ( n3656 & n3657 ) ;
  assign n3659 = ( n482 & n3640 ) | ( n482 & n3658 ) | ( n3640 & n3658 ) ;
  assign n3660 = ( ~n3624 & n3654 ) | ( ~n3624 & n3659 ) | ( n3654 & n3659 ) ;
  assign n3661 = n3653 & ~n3660 ;
  assign n3662 = n3615 & n3661 ;
  assign n3663 = n3615 & ~n3662 ;
  assign n3664 = ~n3615 & n3661 ;
  assign n3665 = n3663 | n3664 ;
  assign n3666 = n2368 & n3635 ;
  assign n3667 = ( ~n2340 & n3635 ) | ( ~n2340 & n3666 ) | ( n3635 & n3666 ) ;
  assign n3668 = ~n2679 & n3667 ;
  assign n3669 = n2827 & n3668 ;
  assign n3670 = ( n3057 & n3635 ) | ( n3057 & n3669 ) | ( n3635 & n3669 ) ;
  assign n3671 = n3049 & n3637 ;
  assign n3672 = n3670 | n3671 ;
  assign n3673 = n3110 & n3641 ;
  assign n3674 = ( ~n3106 & n3641 ) | ( ~n3106 & n3673 ) | ( n3641 & n3673 ) ;
  assign n3675 = n3672 | n3674 ;
  assign n3676 = ( n3098 & ~n3114 ) | ( n3098 & n3115 ) | ( ~n3114 & n3115 ) ;
  assign n3677 = ~n3059 & n3114 ;
  assign n3678 = ~n3098 & n3677 ;
  assign n3679 = n3676 | n3678 ;
  assign n3680 = n3643 | n3674 ;
  assign n3681 = n3672 | n3680 ;
  assign n3682 = ( n3675 & ~n3679 ) | ( n3675 & n3681 ) | ( ~n3679 & n3681 ) ;
  assign n3683 = n482 & n3681 ;
  assign n3684 = n482 & n3674 ;
  assign n3685 = ( n482 & n3672 ) | ( n482 & n3684 ) | ( n3672 & n3684 ) ;
  assign n3686 = ( ~n3679 & n3683 ) | ( ~n3679 & n3685 ) | ( n3683 & n3685 ) ;
  assign n3687 = n3682 & ~n3686 ;
  assign n3688 = n482 & ~n3685 ;
  assign n3689 = n482 & ~n3681 ;
  assign n3690 = ( n3679 & n3688 ) | ( n3679 & n3689 ) | ( n3688 & n3689 ) ;
  assign n3691 = n3687 | n3690 ;
  assign n3692 = n3608 & n3610 ;
  assign n3693 = n3608 | n3610 ;
  assign n3694 = ~n3692 & n3693 ;
  assign n3695 = n3691 & n3694 ;
  assign n3696 = n3691 & ~n3695 ;
  assign n3697 = ( n3694 & ~n3695 ) | ( n3694 & n3696 ) | ( ~n3695 & n3696 ) ;
  assign n3698 = n3554 | n3580 ;
  assign n3699 = ~n3581 & n3698 ;
  assign n3700 = n3070 & n3635 ;
  assign n3701 = n3063 & n3637 ;
  assign n3702 = n3700 | n3701 ;
  assign n3703 = n2368 & n3641 ;
  assign n3704 = ( ~n2340 & n3641 ) | ( ~n2340 & n3703 ) | ( n3641 & n3703 ) ;
  assign n3705 = ~n2679 & n3704 ;
  assign n3706 = n2827 & n3705 ;
  assign n3707 = ( n3057 & n3641 ) | ( n3057 & n3706 ) | ( n3641 & n3706 ) ;
  assign n3708 = n3702 | n3707 ;
  assign n3709 = n3643 | n3707 ;
  assign n3710 = n3702 | n3709 ;
  assign n3711 = ( n3401 & n3708 ) | ( n3401 & n3710 ) | ( n3708 & n3710 ) ;
  assign n3712 = ( n482 & n3656 ) | ( n482 & n3707 ) | ( n3656 & n3707 ) ;
  assign n3713 = n482 | n3656 ;
  assign n3714 = ( n3702 & n3712 ) | ( n3702 & n3713 ) | ( n3712 & n3713 ) ;
  assign n3715 = n482 & n3707 ;
  assign n3716 = ( n482 & n3702 ) | ( n482 & n3715 ) | ( n3702 & n3715 ) ;
  assign n3717 = ( n3401 & n3714 ) | ( n3401 & n3716 ) | ( n3714 & n3716 ) ;
  assign n3718 = n3711 & ~n3717 ;
  assign n3719 = n482 & ~n3656 ;
  assign n3720 = ~n3707 & n3719 ;
  assign n3721 = ~n3702 & n3720 ;
  assign n3722 = n482 & ~n3707 ;
  assign n3723 = ~n3702 & n3722 ;
  assign n3724 = ( ~n3401 & n3721 ) | ( ~n3401 & n3723 ) | ( n3721 & n3723 ) ;
  assign n3725 = n3699 & n3724 ;
  assign n3726 = ( n3699 & n3718 ) | ( n3699 & n3725 ) | ( n3718 & n3725 ) ;
  assign n3727 = n3699 | n3724 ;
  assign n3728 = n3718 | n3727 ;
  assign n3729 = ~n3726 & n3728 ;
  assign n3730 = n3726 | n3729 ;
  assign n3731 = n3564 | n3568 ;
  assign n3732 = n3557 | n3568 ;
  assign n3733 = n3555 | n3568 ;
  assign n3734 = ( n3457 & n3732 ) | ( n3457 & n3733 ) | ( n3732 & n3733 ) ;
  assign n3735 = ( ~n3565 & n3731 ) | ( ~n3565 & n3734 ) | ( n3731 & n3734 ) ;
  assign n3736 = ~n3580 & n3735 ;
  assign n3737 = n3063 & n3641 ;
  assign n3738 = n3070 & n3637 ;
  assign n3739 = ~n2823 & n3635 ;
  assign n3740 = ~n2764 & n3739 ;
  assign n3741 = n3643 | n3740 ;
  assign n3742 = n3635 | n3643 ;
  assign n3743 = ( n3071 & n3741 ) | ( n3071 & n3742 ) | ( n3741 & n3742 ) ;
  assign n3744 = n3738 | n3743 ;
  assign n3745 = n3737 | n3744 ;
  assign n3746 = n482 | n3745 ;
  assign n3747 = n3737 | n3738 ;
  assign n3748 = ( n3071 & n3635 ) | ( n3071 & n3740 ) | ( n3635 & n3740 ) ;
  assign n3749 = n3743 & n3748 ;
  assign n3750 = n482 | n3749 ;
  assign n3751 = n3747 | n3750 ;
  assign n3752 = ( n3510 & n3746 ) | ( n3510 & n3751 ) | ( n3746 & n3751 ) ;
  assign n3753 = n3746 & n3751 ;
  assign n3754 = ( ~n3094 & n3752 ) | ( ~n3094 & n3753 ) | ( n3752 & n3753 ) ;
  assign n3755 = n482 & n3745 ;
  assign n3756 = n482 & n3749 ;
  assign n3757 = ( n482 & n3747 ) | ( n482 & n3756 ) | ( n3747 & n3756 ) ;
  assign n3758 = ( n3510 & n3755 ) | ( n3510 & n3757 ) | ( n3755 & n3757 ) ;
  assign n3759 = n3755 & n3757 ;
  assign n3760 = ( ~n3094 & n3758 ) | ( ~n3094 & n3759 ) | ( n3758 & n3759 ) ;
  assign n3761 = n3754 & ~n3760 ;
  assign n3762 = n3736 & n3761 ;
  assign n3767 = ~n2823 & n3641 ;
  assign n3768 = ~n2764 & n3767 ;
  assign n3769 = ( n3071 & n3641 ) | ( n3071 & n3768 ) | ( n3641 & n3768 ) ;
  assign n3763 = n3085 & n3635 ;
  assign n3764 = n3078 & n3637 ;
  assign n3765 = ( n3082 & n3637 ) | ( n3082 & n3764 ) | ( n3637 & n3764 ) ;
  assign n3766 = n3763 | n3765 ;
  assign n3770 = n3766 | n3769 ;
  assign n3772 = ( n3085 & n3643 ) | ( n3085 & n3742 ) | ( n3643 & n3742 ) ;
  assign n3773 = n3765 | n3772 ;
  assign n3774 = ( n3769 & n3770 ) | ( n3769 & n3773 ) | ( n3770 & n3773 ) ;
  assign n3775 = n3769 | n3773 ;
  assign n3776 = ( ~n3475 & n3774 ) | ( ~n3475 & n3775 ) | ( n3774 & n3775 ) ;
  assign n3771 = n3475 & ~n3770 ;
  assign n3777 = ( ~n482 & n3771 ) | ( ~n482 & n3776 ) | ( n3771 & n3776 ) ;
  assign n3778 = n3776 & ~n3777 ;
  assign n3779 = ~n3771 & n3777 ;
  assign n3780 = ( n482 & ~n3778 ) | ( n482 & n3779 ) | ( ~n3778 & n3779 ) ;
  assign n3781 = n3085 & n3637 ;
  assign n3782 = n3078 & n3641 ;
  assign n3783 = ( n3082 & n3641 ) | ( n3082 & n3782 ) | ( n3641 & n3782 ) ;
  assign n3784 = n3781 | n3783 ;
  assign n3785 = n3457 & n3643 ;
  assign n3786 = n3784 | n3785 ;
  assign n3787 = n482 & n3637 ;
  assign n3788 = n3085 & n3787 ;
  assign n3789 = ( n482 & n3783 ) | ( n482 & n3788 ) | ( n3783 & n3788 ) ;
  assign n3790 = ( n482 & n3785 ) | ( n482 & n3789 ) | ( n3785 & n3789 ) ;
  assign n3791 = n3786 & ~n3790 ;
  assign n3792 = n3085 & n3404 ;
  assign n3793 = n482 & ~n3630 ;
  assign n3794 = ( n482 & ~n3085 ) | ( n482 & n3793 ) | ( ~n3085 & n3793 ) ;
  assign n3795 = n3792 & n3794 ;
  assign n3796 = n482 & ~n3787 ;
  assign n3797 = ( n482 & ~n3085 ) | ( n482 & n3796 ) | ( ~n3085 & n3796 ) ;
  assign n3798 = n3794 & n3797 ;
  assign n3799 = ~n3783 & n3798 ;
  assign n3800 = n3792 & n3799 ;
  assign n3801 = ~n3785 & n3800 ;
  assign n3802 = ( n3791 & n3795 ) | ( n3791 & n3801 ) | ( n3795 & n3801 ) ;
  assign n3803 = n3780 & n3802 ;
  assign n3804 = ~n3785 & n3799 ;
  assign n3805 = ( n3791 & n3794 ) | ( n3791 & n3804 ) | ( n3794 & n3804 ) ;
  assign n3806 = n3780 & n3805 ;
  assign n3807 = ~n3803 & n3806 ;
  assign n3808 = n3792 & ~n3804 ;
  assign n3809 = n3792 & ~n3794 ;
  assign n3810 = ( ~n3791 & n3808 ) | ( ~n3791 & n3809 ) | ( n3808 & n3809 ) ;
  assign n3811 = ( ~n3780 & n3792 ) | ( ~n3780 & n3810 ) | ( n3792 & n3810 ) ;
  assign n3812 = n3807 | n3811 ;
  assign n3813 = n3078 & n3635 ;
  assign n3814 = ( n3082 & n3635 ) | ( n3082 & n3813 ) | ( n3635 & n3813 ) ;
  assign n3815 = n3641 | n3814 ;
  assign n3816 = ( n3070 & n3814 ) | ( n3070 & n3815 ) | ( n3814 & n3815 ) ;
  assign n3817 = ~n2823 & n3637 ;
  assign n3818 = ~n2764 & n3817 ;
  assign n3819 = ( n3071 & n3637 ) | ( n3071 & n3818 ) | ( n3637 & n3818 ) ;
  assign n3820 = n3816 | n3819 ;
  assign n3821 = n3076 & n3088 ;
  assign n3822 = n3643 | n3818 ;
  assign n3823 = n3637 | n3643 ;
  assign n3824 = ( n3071 & n3822 ) | ( n3071 & n3823 ) | ( n3822 & n3823 ) ;
  assign n3825 = n3816 | n3824 ;
  assign n3826 = ( n3820 & n3821 ) | ( n3820 & n3825 ) | ( n3821 & n3825 ) ;
  assign n3827 = n3820 | n3825 ;
  assign n3828 = ( ~n3583 & n3826 ) | ( ~n3583 & n3827 ) | ( n3826 & n3827 ) ;
  assign n3829 = n3088 & n3656 ;
  assign n3830 = n3076 & n3829 ;
  assign n3831 = ( n482 & n3820 ) | ( n482 & n3830 ) | ( n3820 & n3830 ) ;
  assign n3832 = ( n482 & n3656 ) | ( n482 & n3820 ) | ( n3656 & n3820 ) ;
  assign n3833 = ( ~n3583 & n3831 ) | ( ~n3583 & n3832 ) | ( n3831 & n3832 ) ;
  assign n3834 = n3828 & ~n3833 ;
  assign n3835 = ( n482 & ~n3088 ) | ( n482 & n3719 ) | ( ~n3088 & n3719 ) ;
  assign n3836 = n482 | n3719 ;
  assign n3837 = ( ~n3076 & n3835 ) | ( ~n3076 & n3836 ) | ( n3835 & n3836 ) ;
  assign n3838 = ~n3820 & n3837 ;
  assign n3839 = n3719 & ~n3820 ;
  assign n3840 = ( n3583 & n3838 ) | ( n3583 & n3839 ) | ( n3838 & n3839 ) ;
  assign n3841 = n3834 | n3840 ;
  assign n3842 = n3803 | n3841 ;
  assign n3843 = ( n3803 & n3812 ) | ( n3803 & n3842 ) | ( n3812 & n3842 ) ;
  assign n3844 = n3736 | n3761 ;
  assign n3845 = ~n3762 & n3844 ;
  assign n3846 = n3762 | n3845 ;
  assign n3847 = ( n3762 & n3843 ) | ( n3762 & n3846 ) | ( n3843 & n3846 ) ;
  assign n3848 = ( n3726 & n3730 ) | ( n3726 & n3847 ) | ( n3730 & n3847 ) ;
  assign n3849 = n3603 & ~n3605 ;
  assign n3850 = ~n3582 & n3849 ;
  assign n3851 = ~n3603 & n3605 ;
  assign n3852 = ( n3582 & ~n3603 ) | ( n3582 & n3851 ) | ( ~n3603 & n3851 ) ;
  assign n3853 = n3850 | n3852 ;
  assign n3854 = n3061 | n3066 ;
  assign n3855 = n3096 | n3854 ;
  assign n3856 = ~n3098 & n3855 ;
  assign n3857 = n3063 & n3635 ;
  assign n3858 = n2368 & n3637 ;
  assign n3859 = ( ~n2340 & n3637 ) | ( ~n2340 & n3858 ) | ( n3637 & n3858 ) ;
  assign n3860 = ~n2679 & n3859 ;
  assign n3861 = n2827 & n3860 ;
  assign n3862 = ( n3057 & n3637 ) | ( n3057 & n3861 ) | ( n3637 & n3861 ) ;
  assign n3863 = n3857 | n3862 ;
  assign n3864 = n3049 & n3641 ;
  assign n3865 = n3863 | n3864 ;
  assign n3866 = n3643 | n3865 ;
  assign n3867 = n3865 & n3866 ;
  assign n3868 = ( n3856 & n3866 ) | ( n3856 & n3867 ) | ( n3866 & n3867 ) ;
  assign n3869 = n482 & n3865 ;
  assign n3870 = n3866 & n3869 ;
  assign n3871 = ( n482 & n3656 ) | ( n482 & n3865 ) | ( n3656 & n3865 ) ;
  assign n3872 = ( n3856 & n3870 ) | ( n3856 & n3871 ) | ( n3870 & n3871 ) ;
  assign n3873 = n482 & ~n3870 ;
  assign n3874 = n3719 & ~n3865 ;
  assign n3875 = ( ~n3856 & n3873 ) | ( ~n3856 & n3874 ) | ( n3873 & n3874 ) ;
  assign n3876 = ( n3868 & ~n3872 ) | ( n3868 & n3875 ) | ( ~n3872 & n3875 ) ;
  assign n3877 = n3853 & n3876 ;
  assign n3878 = n3853 | n3876 ;
  assign n3879 = ~n3877 & n3878 ;
  assign n3880 = n3877 | n3879 ;
  assign n3881 = ( n3848 & n3877 ) | ( n3848 & n3880 ) | ( n3877 & n3880 ) ;
  assign n3882 = n3695 | n3881 ;
  assign n3883 = ( n3695 & n3697 ) | ( n3695 & n3882 ) | ( n3697 & n3882 ) ;
  assign n3884 = ( n3398 & ~n3665 ) | ( n3398 & n3883 ) | ( ~n3665 & n3883 ) ;
  assign n3885 = ( n3665 & ~n3883 ) | ( n3665 & n3884 ) | ( ~n3883 & n3884 ) ;
  assign n3886 = ( ~n3398 & n3884 ) | ( ~n3398 & n3885 ) | ( n3884 & n3885 ) ;
  assign n3887 = ~n3697 & n3881 ;
  assign n3888 = n3697 & ~n3881 ;
  assign n3889 = n3887 | n3888 ;
  assign n3890 = ( n3037 & n3039 ) | ( n3037 & n3124 ) | ( n3039 & n3124 ) ;
  assign n3891 = n3027 & n3037 ;
  assign n3892 = ( n3040 & n3124 ) | ( n3040 & n3891 ) | ( n3124 & n3891 ) ;
  assign n3893 = n3027 & ~n3891 ;
  assign n3894 = n3027 & ~n3040 ;
  assign n3895 = ( ~n3124 & n3893 ) | ( ~n3124 & n3894 ) | ( n3893 & n3894 ) ;
  assign n3896 = ( n3890 & ~n3892 ) | ( n3890 & n3895 ) | ( ~n3892 & n3895 ) ;
  assign n3897 = n3033 & n3373 ;
  assign n3898 = n2916 & n3367 ;
  assign n3899 = ( ~n2901 & n3367 ) | ( ~n2901 & n3898 ) | ( n3367 & n3898 ) ;
  assign n3900 = ~n2921 & n3899 ;
  assign n3901 = n2828 & n3900 ;
  assign n3902 = ( n2927 & n3367 ) | ( n2927 & n3901 ) | ( n3367 & n3901 ) ;
  assign n3903 = n3897 | n3902 ;
  assign n3904 = n3024 & n3380 ;
  assign n3905 = n3380 | n3387 ;
  assign n3906 = ( n3024 & n3387 ) | ( n3024 & n3905 ) | ( n3387 & n3905 ) ;
  assign n3907 = n3904 & n3906 ;
  assign n3908 = n3903 | n3907 ;
  assign n3909 = n1115 | n3908 ;
  assign n3910 = n1115 | n3905 ;
  assign n3911 = ( n3024 & n3394 ) | ( n3024 & n3910 ) | ( n3394 & n3910 ) ;
  assign n3912 = n3903 | n3911 ;
  assign n3913 = ( n3896 & n3909 ) | ( n3896 & n3912 ) | ( n3909 & n3912 ) ;
  assign n3914 = n1115 & n3908 ;
  assign n3915 = n1115 & n3905 ;
  assign n3916 = ( n3024 & n3388 ) | ( n3024 & n3915 ) | ( n3388 & n3915 ) ;
  assign n3917 = ( n1115 & n3903 ) | ( n1115 & n3916 ) | ( n3903 & n3916 ) ;
  assign n3918 = ( n3896 & n3914 ) | ( n3896 & n3917 ) | ( n3914 & n3917 ) ;
  assign n3919 = n3913 & ~n3918 ;
  assign n3920 = n3889 & n3919 ;
  assign n3921 = n3889 | n3919 ;
  assign n3922 = ~n3920 & n3921 ;
  assign n3923 = n3848 & n3879 ;
  assign n3924 = n3848 & ~n3923 ;
  assign n3925 = ~n3848 & n3879 ;
  assign n3926 = n3924 | n3925 ;
  assign n3927 = n3049 & n3373 ;
  assign n3928 = n3110 & n3367 ;
  assign n3929 = ( ~n3106 & n3367 ) | ( ~n3106 & n3928 ) | ( n3367 & n3928 ) ;
  assign n3930 = n3927 | n3929 ;
  assign n3931 = n3033 & n3380 ;
  assign n3932 = ( n3033 & n3387 ) | ( n3033 & n3905 ) | ( n3387 & n3905 ) ;
  assign n3933 = n3931 & n3932 ;
  assign n3934 = n3930 | n3933 ;
  assign n3935 = n1115 | n3934 ;
  assign n3936 = ( n3033 & n3394 ) | ( n3033 & n3910 ) | ( n3394 & n3910 ) ;
  assign n3937 = n3930 | n3936 ;
  assign n3938 = ( ~n3624 & n3935 ) | ( ~n3624 & n3937 ) | ( n3935 & n3937 ) ;
  assign n3939 = n1115 & n3934 ;
  assign n3940 = ( n3033 & n3388 ) | ( n3033 & n3915 ) | ( n3388 & n3915 ) ;
  assign n3941 = ( n1115 & n3930 ) | ( n1115 & n3940 ) | ( n3930 & n3940 ) ;
  assign n3942 = ( ~n3624 & n3939 ) | ( ~n3624 & n3941 ) | ( n3939 & n3941 ) ;
  assign n3943 = n3938 & ~n3942 ;
  assign n3944 = ~n3729 & n3847 ;
  assign n3945 = n3729 & ~n3847 ;
  assign n3946 = n3944 | n3945 ;
  assign n3947 = n3943 & n3946 ;
  assign n3948 = n3946 & ~n3947 ;
  assign n3949 = ( n3943 & ~n3947 ) | ( n3943 & n3948 ) | ( ~n3947 & n3948 ) ;
  assign n3950 = n3038 & n3124 ;
  assign n3951 = n3038 | n3124 ;
  assign n3952 = ~n3950 & n3951 ;
  assign n3953 = n3033 & n3367 ;
  assign n3954 = n3110 & n3373 ;
  assign n3955 = ( ~n3106 & n3373 ) | ( ~n3106 & n3954 ) | ( n3373 & n3954 ) ;
  assign n3956 = n3953 | n3955 ;
  assign n3957 = n2916 & n3380 ;
  assign n3958 = ( ~n2901 & n3380 ) | ( ~n2901 & n3957 ) | ( n3380 & n3957 ) ;
  assign n3959 = ~n2921 & n3958 ;
  assign n3960 = n2828 & n3959 ;
  assign n3961 = ( n2927 & n3380 ) | ( n2927 & n3960 ) | ( n3380 & n3960 ) ;
  assign n3962 = n3956 | n3961 ;
  assign n3963 = ( n3387 & n3952 ) | ( n3387 & n3962 ) | ( n3952 & n3962 ) ;
  assign n3964 = ( n1115 & n3387 ) | ( n1115 & ~n3962 ) | ( n3387 & ~n3962 ) ;
  assign n3965 = ( n1115 & n3952 ) | ( n1115 & n3964 ) | ( n3952 & n3964 ) ;
  assign n3966 = ~n3963 & n3965 ;
  assign n3967 = n3962 | n3964 ;
  assign n3968 = n1115 | n3962 ;
  assign n3969 = ( n3952 & n3967 ) | ( n3952 & n3968 ) | ( n3967 & n3968 ) ;
  assign n3970 = ( ~n1115 & n3966 ) | ( ~n1115 & n3969 ) | ( n3966 & n3969 ) ;
  assign n3971 = ( n3926 & n3949 ) | ( n3926 & n3970 ) | ( n3949 & n3970 ) ;
  assign n3972 = n2368 & n3373 ;
  assign n3973 = ( ~n2340 & n3373 ) | ( ~n2340 & n3972 ) | ( n3373 & n3972 ) ;
  assign n3974 = ~n2679 & n3973 ;
  assign n3975 = n2827 & n3974 ;
  assign n3976 = ( n3057 & n3373 ) | ( n3057 & n3975 ) | ( n3373 & n3975 ) ;
  assign n3977 = n3049 & n3367 ;
  assign n3978 = n3976 | n3977 ;
  assign n3979 = n3110 & n3380 ;
  assign n3980 = ( ~n3106 & n3380 ) | ( ~n3106 & n3979 ) | ( n3380 & n3979 ) ;
  assign n3981 = n3387 | n3980 ;
  assign n3982 = n3978 | n3981 ;
  assign n3983 = n1115 & n3982 ;
  assign n3984 = n1115 & n3980 ;
  assign n3985 = ( n1115 & n3978 ) | ( n1115 & n3984 ) | ( n3978 & n3984 ) ;
  assign n3986 = ( ~n3679 & n3983 ) | ( ~n3679 & n3985 ) | ( n3983 & n3985 ) ;
  assign n3987 = n1115 | n3982 ;
  assign n3988 = n1115 | n3980 ;
  assign n3989 = n3978 | n3988 ;
  assign n3990 = ( ~n3679 & n3987 ) | ( ~n3679 & n3989 ) | ( n3987 & n3989 ) ;
  assign n3991 = ~n3986 & n3990 ;
  assign n3992 = n3843 & n3845 ;
  assign n3993 = n3843 | n3845 ;
  assign n3994 = ~n3992 & n3993 ;
  assign n3995 = n3991 & n3994 ;
  assign n3996 = n3991 | n3994 ;
  assign n3997 = ~n3995 & n3996 ;
  assign n3998 = n3995 | n3997 ;
  assign n3999 = ~n3811 & n3841 ;
  assign n4000 = ~n3807 & n3999 ;
  assign n4001 = n3811 & ~n3841 ;
  assign n4002 = ( n3807 & ~n3841 ) | ( n3807 & n4001 ) | ( ~n3841 & n4001 ) ;
  assign n4003 = n4000 | n4002 ;
  assign n4004 = n3063 & n3373 ;
  assign n4005 = n2368 & n3367 ;
  assign n4006 = ( ~n2340 & n3367 ) | ( ~n2340 & n4005 ) | ( n3367 & n4005 ) ;
  assign n4007 = ~n2679 & n4006 ;
  assign n4008 = n2827 & n4007 ;
  assign n4009 = ( n3057 & n3367 ) | ( n3057 & n4008 ) | ( n3367 & n4008 ) ;
  assign n4010 = n4004 | n4009 ;
  assign n4011 = n3049 & n3380 ;
  assign n4012 = n4010 | n4011 ;
  assign n4013 = n3387 | n4012 ;
  assign n4014 = n4012 & n4013 ;
  assign n4015 = ( n3856 & n4013 ) | ( n3856 & n4014 ) | ( n4013 & n4014 ) ;
  assign n4016 = n1115 & n4012 ;
  assign n4017 = n4013 & n4016 ;
  assign n4018 = ( n1115 & n3388 ) | ( n1115 & n4012 ) | ( n3388 & n4012 ) ;
  assign n4019 = ( n3856 & n4017 ) | ( n3856 & n4018 ) | ( n4017 & n4018 ) ;
  assign n4020 = n1115 & ~n4017 ;
  assign n4021 = n1115 & ~n3388 ;
  assign n4022 = ~n4012 & n4021 ;
  assign n4023 = ( ~n3856 & n4020 ) | ( ~n3856 & n4022 ) | ( n4020 & n4022 ) ;
  assign n4024 = ( n4015 & ~n4019 ) | ( n4015 & n4023 ) | ( ~n4019 & n4023 ) ;
  assign n4025 = n4003 & n4024 ;
  assign n4026 = n3070 & n3373 ;
  assign n4027 = n3063 & n3367 ;
  assign n4028 = n4026 | n4027 ;
  assign n4029 = n2368 & n3380 ;
  assign n4030 = ( ~n2340 & n3380 ) | ( ~n2340 & n4029 ) | ( n3380 & n4029 ) ;
  assign n4031 = ~n2679 & n4030 ;
  assign n4032 = n2827 & n4031 ;
  assign n4033 = ( n3057 & n3380 ) | ( n3057 & n4032 ) | ( n3380 & n4032 ) ;
  assign n4034 = n1115 & n3363 ;
  assign n4035 = n3371 & n4034 ;
  assign n4036 = ( n1115 & n4033 ) | ( n1115 & n4035 ) | ( n4033 & n4035 ) ;
  assign n4037 = n1115 | n4035 ;
  assign n4038 = ( n4028 & n4036 ) | ( n4028 & n4037 ) | ( n4036 & n4037 ) ;
  assign n4039 = n1115 & n4033 ;
  assign n4040 = ( n1115 & n4028 ) | ( n1115 & n4039 ) | ( n4028 & n4039 ) ;
  assign n4041 = ( n3401 & n4038 ) | ( n3401 & n4040 ) | ( n4038 & n4040 ) ;
  assign n4042 = n1115 | n3363 ;
  assign n4043 = ( n1115 & n3371 ) | ( n1115 & n4042 ) | ( n3371 & n4042 ) ;
  assign n4044 = n4033 | n4043 ;
  assign n4045 = n4028 | n4044 ;
  assign n4046 = n1115 | n4033 ;
  assign n4047 = n4028 | n4046 ;
  assign n4048 = ( n3401 & n4045 ) | ( n3401 & n4047 ) | ( n4045 & n4047 ) ;
  assign n4049 = ~n4041 & n4048 ;
  assign n4050 = n3780 | n3805 ;
  assign n4051 = ~n3806 & n4050 ;
  assign n4052 = n4049 & n4051 ;
  assign n4053 = n4049 | n4051 ;
  assign n4054 = ~n4052 & n4053 ;
  assign n4055 = n3794 | n3797 ;
  assign n4056 = ( ~n3783 & n3794 ) | ( ~n3783 & n4055 ) | ( n3794 & n4055 ) ;
  assign n4057 = ( ~n3785 & n3794 ) | ( ~n3785 & n4056 ) | ( n3794 & n4056 ) ;
  assign n4058 = n3791 | n4057 ;
  assign n4059 = ~n3805 & n4058 ;
  assign n4060 = n3063 & n3380 ;
  assign n4061 = n3070 & n3367 ;
  assign n4062 = ~n2823 & n3373 ;
  assign n4063 = ~n2764 & n4062 ;
  assign n4064 = n3387 | n4063 ;
  assign n4065 = n3373 | n3387 ;
  assign n4066 = ( n3071 & n4064 ) | ( n3071 & n4065 ) | ( n4064 & n4065 ) ;
  assign n4067 = n4061 | n4066 ;
  assign n4068 = n4060 | n4067 ;
  assign n4069 = n1115 | n4068 ;
  assign n4070 = n4060 | n4061 ;
  assign n4071 = ( n3071 & n3373 ) | ( n3071 & n4063 ) | ( n3373 & n4063 ) ;
  assign n4072 = n4066 & n4071 ;
  assign n4073 = n1115 | n4072 ;
  assign n4074 = n4070 | n4073 ;
  assign n4075 = ( n3510 & n4069 ) | ( n3510 & n4074 ) | ( n4069 & n4074 ) ;
  assign n4076 = n4069 & n4074 ;
  assign n4077 = ( ~n3094 & n4075 ) | ( ~n3094 & n4076 ) | ( n4075 & n4076 ) ;
  assign n4078 = n1115 & n4068 ;
  assign n4079 = n1115 & n4072 ;
  assign n4080 = ( n1115 & n4070 ) | ( n1115 & n4079 ) | ( n4070 & n4079 ) ;
  assign n4081 = ( n3510 & n4078 ) | ( n3510 & n4080 ) | ( n4078 & n4080 ) ;
  assign n4082 = n4078 & n4080 ;
  assign n4083 = ( ~n3094 & n4081 ) | ( ~n3094 & n4082 ) | ( n4081 & n4082 ) ;
  assign n4084 = n4077 & ~n4083 ;
  assign n4085 = n4059 & n4084 ;
  assign n4090 = ~n2823 & n3380 ;
  assign n4091 = ~n2764 & n4090 ;
  assign n4092 = ( n3071 & n3380 ) | ( n3071 & n4091 ) | ( n3380 & n4091 ) ;
  assign n4086 = n3085 & n3373 ;
  assign n4087 = n3078 & n3367 ;
  assign n4088 = ( n3082 & n3367 ) | ( n3082 & n4087 ) | ( n3367 & n4087 ) ;
  assign n4089 = n4086 | n4088 ;
  assign n4093 = n4089 | n4092 ;
  assign n4095 = ( n3085 & n3387 ) | ( n3085 & n4065 ) | ( n3387 & n4065 ) ;
  assign n4096 = n4088 | n4095 ;
  assign n4097 = ( n4092 & n4093 ) | ( n4092 & n4096 ) | ( n4093 & n4096 ) ;
  assign n4098 = n4092 | n4096 ;
  assign n4099 = ( ~n3475 & n4097 ) | ( ~n3475 & n4098 ) | ( n4097 & n4098 ) ;
  assign n4094 = n3475 & ~n4093 ;
  assign n4100 = ( ~n1115 & n4094 ) | ( ~n1115 & n4099 ) | ( n4094 & n4099 ) ;
  assign n4101 = n4099 & ~n4100 ;
  assign n4102 = ~n4094 & n4100 ;
  assign n4103 = ( n1115 & ~n4101 ) | ( n1115 & n4102 ) | ( ~n4101 & n4102 ) ;
  assign n4105 = n3367 | n3387 ;
  assign n4106 = ( n3085 & n3387 ) | ( n3085 & n4105 ) | ( n3387 & n4105 ) ;
  assign n4108 = n3078 & n3380 ;
  assign n4109 = ( n3082 & n3380 ) | ( n3082 & n4108 ) | ( n3380 & n4108 ) ;
  assign n4110 = ~n4106 & n4109 ;
  assign n4104 = n3085 & n3367 ;
  assign n4111 = ~n4104 & n4109 ;
  assign n4112 = ( ~n3457 & n4110 ) | ( ~n3457 & n4111 ) | ( n4110 & n4111 ) ;
  assign n4107 = ( n3457 & n4104 ) | ( n3457 & n4106 ) | ( n4104 & n4106 ) ;
  assign n4113 = ( n1115 & ~n4107 ) | ( n1115 & n4112 ) | ( ~n4107 & n4112 ) ;
  assign n4114 = ( n1115 & n4112 ) | ( n1115 & ~n4113 ) | ( n4112 & ~n4113 ) ;
  assign n4115 = n3085 & n3630 ;
  assign n4116 = n1115 & ~n3363 ;
  assign n4117 = ( n1115 & ~n3085 ) | ( n1115 & n4116 ) | ( ~n3085 & n4116 ) ;
  assign n4118 = n4115 & n4117 ;
  assign n4119 = n4113 & n4118 ;
  assign n4120 = n4106 & n4118 ;
  assign n4121 = n4104 & n4118 ;
  assign n4122 = ( n3457 & n4120 ) | ( n3457 & n4121 ) | ( n4120 & n4121 ) ;
  assign n4123 = ( ~n4114 & n4119 ) | ( ~n4114 & n4122 ) | ( n4119 & n4122 ) ;
  assign n4124 = n4103 & n4123 ;
  assign n4125 = n4113 & n4117 ;
  assign n4126 = n4106 & n4117 ;
  assign n4127 = n4104 & n4117 ;
  assign n4128 = ( n3457 & n4126 ) | ( n3457 & n4127 ) | ( n4126 & n4127 ) ;
  assign n4129 = ( ~n4114 & n4125 ) | ( ~n4114 & n4128 ) | ( n4125 & n4128 ) ;
  assign n4130 = n4103 & n4129 ;
  assign n4131 = ~n4124 & n4130 ;
  assign n4132 = n3078 & n3373 ;
  assign n4133 = ( n3082 & n3373 ) | ( n3082 & n4132 ) | ( n3373 & n4132 ) ;
  assign n4134 = n3380 | n4133 ;
  assign n4135 = ( n3070 & n4133 ) | ( n3070 & n4134 ) | ( n4133 & n4134 ) ;
  assign n4136 = ~n2823 & n3367 ;
  assign n4137 = ~n2764 & n4136 ;
  assign n4138 = ( n3071 & n3367 ) | ( n3071 & n4137 ) | ( n3367 & n4137 ) ;
  assign n4139 = n4135 | n4138 ;
  assign n4140 = n3088 & n4035 ;
  assign n4141 = n3076 & n4140 ;
  assign n4142 = ( n1115 & n4139 ) | ( n1115 & n4141 ) | ( n4139 & n4141 ) ;
  assign n4143 = ( n1115 & n4035 ) | ( n1115 & n4139 ) | ( n4035 & n4139 ) ;
  assign n4144 = ( ~n3583 & n4142 ) | ( ~n3583 & n4143 ) | ( n4142 & n4143 ) ;
  assign n4145 = ( n1115 & n3088 ) | ( n1115 & n4043 ) | ( n3088 & n4043 ) ;
  assign n4146 = n1115 & n4043 ;
  assign n4147 = ( n3076 & n4145 ) | ( n3076 & n4146 ) | ( n4145 & n4146 ) ;
  assign n4148 = n4139 | n4147 ;
  assign n4149 = n1115 | n4043 ;
  assign n4150 = n4139 | n4149 ;
  assign n4151 = ( ~n3583 & n4148 ) | ( ~n3583 & n4150 ) | ( n4148 & n4150 ) ;
  assign n4152 = ~n4144 & n4151 ;
  assign n4153 = n4115 & ~n4123 ;
  assign n4154 = ( ~n4103 & n4115 ) | ( ~n4103 & n4153 ) | ( n4115 & n4153 ) ;
  assign n4155 = n4152 & n4154 ;
  assign n4156 = ( n4131 & n4152 ) | ( n4131 & n4155 ) | ( n4152 & n4155 ) ;
  assign n4157 = n4124 | n4156 ;
  assign n4158 = n4059 | n4084 ;
  assign n4159 = ~n4085 & n4158 ;
  assign n4160 = n4085 | n4159 ;
  assign n4161 = ( n4085 & n4157 ) | ( n4085 & n4160 ) | ( n4157 & n4160 ) ;
  assign n4162 = n4054 & n4161 ;
  assign n4163 = n4052 | n4162 ;
  assign n4164 = n4003 | n4024 ;
  assign n4165 = ~n4025 & n4164 ;
  assign n4166 = n4025 | n4165 ;
  assign n4167 = ( n4025 & n4163 ) | ( n4025 & n4166 ) | ( n4163 & n4166 ) ;
  assign n4168 = n3947 | n4167 ;
  assign n4169 = n3947 | n3995 ;
  assign n4170 = ( n3998 & n4168 ) | ( n3998 & n4169 ) | ( n4168 & n4169 ) ;
  assign n4171 = ( n3925 & n3947 ) | ( n3925 & n3970 ) | ( n3947 & n3970 ) ;
  assign n4172 = n3947 | n3970 ;
  assign n4173 = ( n3924 & n4171 ) | ( n3924 & n4172 ) | ( n4171 & n4172 ) ;
  assign n4174 = ( n3971 & n4170 ) | ( n3971 & n4173 ) | ( n4170 & n4173 ) ;
  assign n4175 = n3920 | n4174 ;
  assign n4176 = ( n3920 & n3922 ) | ( n3920 & n4175 ) | ( n3922 & n4175 ) ;
  assign n4177 = n3886 & n4176 ;
  assign n4178 = n3886 | n4176 ;
  assign n4179 = ~n4177 & n4178 ;
  assign n4180 = n3357 & n4179 ;
  assign n4181 = n4179 & ~n4180 ;
  assign n4182 = ( n3357 & ~n4180 ) | ( n3357 & n4181 ) | ( ~n4180 & n4181 ) ;
  assign n4183 = ( n3127 & n3303 ) | ( n3127 & ~n3306 ) | ( n3303 & ~n3306 ) ;
  assign n4184 = n3306 & n3308 ;
  assign n4185 = ~n3303 & n3308 ;
  assign n4186 = ( ~n3127 & n4184 ) | ( ~n3127 & n4185 ) | ( n4184 & n4185 ) ;
  assign n4187 = n3308 & ~n4185 ;
  assign n4188 = ~n3306 & n3308 ;
  assign n4189 = ( n3127 & n4187 ) | ( n3127 & n4188 ) | ( n4187 & n4188 ) ;
  assign n4190 = ( n4183 & n4186 ) | ( n4183 & ~n4189 ) | ( n4186 & ~n4189 ) ;
  assign n4191 = n3024 & n3333 ;
  assign n4192 = n3296 & n3335 ;
  assign n4193 = n3295 & n3335 ;
  assign n4194 = ( n2828 & n4192 ) | ( n2828 & n4193 ) | ( n4192 & n4193 ) ;
  assign n4195 = ( ~n3300 & n3335 ) | ( ~n3300 & n4194 ) | ( n3335 & n4194 ) ;
  assign n4196 = n4191 | n4195 ;
  assign n4197 = x0 & n3322 ;
  assign n4198 = ( x0 & n3325 ) | ( x0 & n4197 ) | ( n3325 & n4197 ) ;
  assign n4199 = ~n3332 & n4198 ;
  assign n4200 = n3266 & n4199 ;
  assign n4201 = ( n3326 & n4196 ) | ( n3326 & n4200 ) | ( n4196 & n4200 ) ;
  assign n4202 = ( n3266 & n3352 ) | ( n3266 & n3353 ) | ( n3352 & n3353 ) ;
  assign n4203 = ( n3326 & n4196 ) | ( n3326 & n4202 ) | ( n4196 & n4202 ) ;
  assign n4204 = ( ~n4190 & n4201 ) | ( ~n4190 & n4203 ) | ( n4201 & n4203 ) ;
  assign n4205 = x0 | n3322 ;
  assign n4206 = n3325 | n4205 ;
  assign n4207 = ( n3326 & ~n3332 ) | ( n3326 & n4206 ) | ( ~n3332 & n4206 ) ;
  assign n4208 = ( n3266 & n3326 ) | ( n3266 & n4207 ) | ( n3326 & n4207 ) ;
  assign n4209 = n4196 | n4208 ;
  assign n4210 = ( n3266 & n3346 ) | ( n3266 & n3347 ) | ( n3346 & n3347 ) ;
  assign n4211 = n4196 | n4210 ;
  assign n4212 = ( ~n4190 & n4209 ) | ( ~n4190 & n4211 ) | ( n4209 & n4211 ) ;
  assign n4213 = ~n4204 & n4212 ;
  assign n4214 = n3024 & n3335 ;
  assign n4215 = n2916 & n3333 ;
  assign n4216 = ( ~n2901 & n3333 ) | ( ~n2901 & n4215 ) | ( n3333 & n4215 ) ;
  assign n4217 = ~n2921 & n4216 ;
  assign n4218 = n2828 & n4217 ;
  assign n4219 = ( n2927 & n3333 ) | ( n2927 & n4218 ) | ( n3333 & n4218 ) ;
  assign n4220 = n4214 | n4219 ;
  assign n4221 = n3296 & n3338 ;
  assign n4222 = n3295 & n3338 ;
  assign n4223 = ( n2828 & n4221 ) | ( n2828 & n4222 ) | ( n4221 & n4222 ) ;
  assign n4224 = ( ~n3300 & n3338 ) | ( ~n3300 & n4223 ) | ( n3338 & n4223 ) ;
  assign n4225 = ~n3326 & n4224 ;
  assign n4226 = ( ~n3326 & n4220 ) | ( ~n3326 & n4225 ) | ( n4220 & n4225 ) ;
  assign n4227 = ~n3326 & n3340 ;
  assign n4228 = ( ~n3326 & n4224 ) | ( ~n3326 & n4227 ) | ( n4224 & n4227 ) ;
  assign n4229 = ( ~n3326 & n4220 ) | ( ~n3326 & n4228 ) | ( n4220 & n4228 ) ;
  assign n4230 = ( ~n3360 & n4226 ) | ( ~n3360 & n4229 ) | ( n4226 & n4229 ) ;
  assign n4231 = n3326 & ~n4224 ;
  assign n4232 = ~n4220 & n4231 ;
  assign n4233 = n3326 & ~n3340 ;
  assign n4234 = ~n4224 & n4233 ;
  assign n4235 = ~n4220 & n4234 ;
  assign n4236 = ( n3360 & n4232 ) | ( n3360 & n4235 ) | ( n4232 & n4235 ) ;
  assign n4237 = n4230 | n4236 ;
  assign n4238 = ( n3995 & n3998 ) | ( n3995 & n4167 ) | ( n3998 & n4167 ) ;
  assign n4239 = n3949 & n4238 ;
  assign n4240 = n3949 | n4238 ;
  assign n4241 = ~n4239 & n4240 ;
  assign n4242 = n2368 & n3333 ;
  assign n4243 = ( ~n2340 & n3333 ) | ( ~n2340 & n4242 ) | ( n3333 & n4242 ) ;
  assign n4244 = ~n2679 & n4243 ;
  assign n4245 = n2827 & n4244 ;
  assign n4246 = ( n3057 & n3333 ) | ( n3057 & n4245 ) | ( n3333 & n4245 ) ;
  assign n4247 = n3049 & n3335 ;
  assign n4248 = n4246 | n4247 ;
  assign n4249 = n3110 & n3338 ;
  assign n4250 = ( ~n3106 & n3338 ) | ( ~n3106 & n4249 ) | ( n3338 & n4249 ) ;
  assign n4251 = n4248 | n4250 ;
  assign n4252 = n3340 | n4250 ;
  assign n4253 = n4248 | n4252 ;
  assign n4254 = ( ~n3679 & n4251 ) | ( ~n3679 & n4253 ) | ( n4251 & n4253 ) ;
  assign n4255 = n3326 & n4253 ;
  assign n4256 = n3326 & n4250 ;
  assign n4257 = ( n3326 & n4248 ) | ( n3326 & n4256 ) | ( n4248 & n4256 ) ;
  assign n4258 = ( ~n3679 & n4255 ) | ( ~n3679 & n4257 ) | ( n4255 & n4257 ) ;
  assign n4259 = n4254 & ~n4258 ;
  assign n4260 = n3326 & ~n4257 ;
  assign n4261 = n3326 & ~n4253 ;
  assign n4262 = ( n3679 & n4260 ) | ( n3679 & n4261 ) | ( n4260 & n4261 ) ;
  assign n4263 = n4259 | n4262 ;
  assign n4264 = n4152 & ~n4154 ;
  assign n4265 = ~n4131 & n4264 ;
  assign n4266 = ~n4152 & n4154 ;
  assign n4267 = ( n4131 & ~n4152 ) | ( n4131 & n4266 ) | ( ~n4152 & n4266 ) ;
  assign n4268 = n4265 | n4267 ;
  assign n4269 = n3070 & n3333 ;
  assign n4270 = n3063 & n3335 ;
  assign n4271 = n4269 | n4270 ;
  assign n4272 = n2368 & n3338 ;
  assign n4273 = ( ~n2340 & n3338 ) | ( ~n2340 & n4272 ) | ( n3338 & n4272 ) ;
  assign n4274 = ~n2679 & n4273 ;
  assign n4275 = n2827 & n4274 ;
  assign n4276 = ( n3057 & n3338 ) | ( n3057 & n4275 ) | ( n3338 & n4275 ) ;
  assign n4277 = n4271 | n4276 ;
  assign n4278 = n3340 | n4276 ;
  assign n4279 = n4271 | n4278 ;
  assign n4280 = ( n3401 & n4277 ) | ( n3401 & n4279 ) | ( n4277 & n4279 ) ;
  assign n4281 = n3332 & n4198 ;
  assign n4282 = n3326 | n4281 ;
  assign n4283 = ( n3326 & n4276 ) | ( n3326 & n4281 ) | ( n4276 & n4281 ) ;
  assign n4284 = ( n4271 & n4282 ) | ( n4271 & n4283 ) | ( n4282 & n4283 ) ;
  assign n4285 = n3326 & n4276 ;
  assign n4286 = ( n3326 & n4271 ) | ( n3326 & n4285 ) | ( n4271 & n4285 ) ;
  assign n4287 = ( n3401 & n4284 ) | ( n3401 & n4286 ) | ( n4284 & n4286 ) ;
  assign n4288 = n4280 & ~n4287 ;
  assign n4289 = n3326 & ~n4198 ;
  assign n4290 = ( n3326 & ~n3332 ) | ( n3326 & n4289 ) | ( ~n3332 & n4289 ) ;
  assign n4291 = ~n4276 & n4290 ;
  assign n4292 = ~n4271 & n4291 ;
  assign n4293 = n3326 & ~n4276 ;
  assign n4294 = ~n4271 & n4293 ;
  assign n4295 = ( ~n3401 & n4292 ) | ( ~n3401 & n4294 ) | ( n4292 & n4294 ) ;
  assign n4296 = n4288 | n4295 ;
  assign n4297 = n3510 & n4281 ;
  assign n4298 = ~n3094 & n4297 ;
  assign n4299 = ( n3326 & n3332 ) | ( n3326 & n4206 ) | ( n3332 & n4206 ) ;
  assign n4300 = n3063 & n3338 ;
  assign n4301 = n3070 & n3335 ;
  assign n4302 = ~n2823 & n3333 ;
  assign n4303 = ~n2764 & n4302 ;
  assign n4304 = ( n3071 & n3333 ) | ( n3071 & n4303 ) | ( n3333 & n4303 ) ;
  assign n4305 = ( ~n4299 & n4301 ) | ( ~n4299 & n4304 ) | ( n4301 & n4304 ) ;
  assign n4306 = n4299 & ~n4303 ;
  assign n4307 = ~n3333 & n4299 ;
  assign n4308 = ( ~n3071 & n4306 ) | ( ~n3071 & n4307 ) | ( n4306 & n4307 ) ;
  assign n4309 = ( n4300 & n4305 ) | ( n4300 & ~n4308 ) | ( n4305 & ~n4308 ) ;
  assign n4310 = n4299 | n4309 ;
  assign n4311 = n3326 | n4303 ;
  assign n4312 = n3326 | n3333 ;
  assign n4313 = ( n3071 & n4311 ) | ( n3071 & n4312 ) | ( n4311 & n4312 ) ;
  assign n4314 = n4301 | n4313 ;
  assign n4315 = n4300 | n4314 ;
  assign n4316 = ( n3510 & n4310 ) | ( n3510 & n4315 ) | ( n4310 & n4315 ) ;
  assign n4317 = n4310 & n4315 ;
  assign n4318 = ( ~n3094 & n4316 ) | ( ~n3094 & n4317 ) | ( n4316 & n4317 ) ;
  assign n4319 = ~n4298 & n4318 ;
  assign n4320 = n3078 & n3333 ;
  assign n4321 = ( n3082 & n3333 ) | ( n3082 & n4320 ) | ( n3333 & n4320 ) ;
  assign n4322 = n3338 | n4321 ;
  assign n4323 = ( n3070 & n4321 ) | ( n3070 & n4322 ) | ( n4321 & n4322 ) ;
  assign n4324 = ~n2823 & n3335 ;
  assign n4325 = ~n2764 & n4324 ;
  assign n4326 = ( n3071 & n3335 ) | ( n3071 & n4325 ) | ( n3335 & n4325 ) ;
  assign n4327 = n4323 | n4326 ;
  assign n4328 = n3088 & n4281 ;
  assign n4329 = n3076 & n4328 ;
  assign n4330 = ( n3326 & n4327 ) | ( n3326 & n4329 ) | ( n4327 & n4329 ) ;
  assign n4331 = ( n3326 & n4281 ) | ( n3326 & n4327 ) | ( n4281 & n4327 ) ;
  assign n4332 = ( ~n3583 & n4330 ) | ( ~n3583 & n4331 ) | ( n4330 & n4331 ) ;
  assign n4333 = ( n3088 & n3326 ) | ( n3088 & n4299 ) | ( n3326 & n4299 ) ;
  assign n4334 = n3326 & n4299 ;
  assign n4335 = ( n3076 & n4333 ) | ( n3076 & n4334 ) | ( n4333 & n4334 ) ;
  assign n4336 = n4327 | n4335 ;
  assign n4337 = n3326 | n4206 ;
  assign n4338 = ( n3326 & n3332 ) | ( n3326 & n4337 ) | ( n3332 & n4337 ) ;
  assign n4339 = n4327 | n4338 ;
  assign n4340 = ( ~n3583 & n4336 ) | ( ~n3583 & n4339 ) | ( n4336 & n4339 ) ;
  assign n4341 = ~n4332 & n4340 ;
  assign n4342 = n4113 | n4117 ;
  assign n4343 = n4106 | n4117 ;
  assign n4344 = n4104 | n4117 ;
  assign n4345 = ( n3457 & n4343 ) | ( n3457 & n4344 ) | ( n4343 & n4344 ) ;
  assign n4346 = ( ~n4114 & n4342 ) | ( ~n4114 & n4345 ) | ( n4342 & n4345 ) ;
  assign n4347 = ~n4129 & n4346 ;
  assign n4348 = n3085 & n3363 ;
  assign n4349 = ~n3475 & n4281 ;
  assign n4350 = n3457 & n4281 ;
  assign n4351 = n3326 & ~n3335 ;
  assign n4352 = ( ~n3085 & n3326 ) | ( ~n3085 & n4351 ) | ( n3326 & n4351 ) ;
  assign n4353 = n3078 & n3338 ;
  assign n4354 = ( n3082 & n3338 ) | ( n3082 & n4353 ) | ( n3338 & n4353 ) ;
  assign n4355 = n4352 & ~n4354 ;
  assign n4356 = ~n4350 & n4355 ;
  assign n4357 = n3322 & ~n3323 ;
  assign n4358 = ( ~n3323 & n3325 ) | ( ~n3323 & n4357 ) | ( n3325 & n4357 ) ;
  assign n4359 = n3332 & n4358 ;
  assign n4360 = n3085 & n4359 ;
  assign n4361 = n3078 & n3335 ;
  assign n4362 = ( n3082 & n3335 ) | ( n3082 & n4361 ) | ( n3335 & n4361 ) ;
  assign n4363 = ( n3326 & n4360 ) | ( n3326 & n4362 ) | ( n4360 & n4362 ) ;
  assign n4364 = ~n2823 & n3338 ;
  assign n4365 = ~n2764 & n4364 ;
  assign n4366 = ( n3071 & n3338 ) | ( n3071 & n4365 ) | ( n3338 & n4365 ) ;
  assign n4367 = ( n3326 & n4363 ) | ( n3326 & n4366 ) | ( n4363 & n4366 ) ;
  assign n4368 = n4356 & ~n4367 ;
  assign n4369 = ~n4349 & n4368 ;
  assign n4370 = x0 & n3085 ;
  assign n4371 = ~n4348 & n4370 ;
  assign n4372 = ( n4348 & n4369 ) | ( n4348 & ~n4371 ) | ( n4369 & ~n4371 ) ;
  assign n4373 = n4347 | n4372 ;
  assign n4374 = n4348 & ~n4370 ;
  assign n4375 = n4369 & n4374 ;
  assign n4376 = n4347 | n4375 ;
  assign n4377 = ( n4341 & n4373 ) | ( n4341 & n4376 ) | ( n4373 & n4376 ) ;
  assign n4378 = n4319 & n4377 ;
  assign n4379 = n4347 & n4372 ;
  assign n4380 = n4347 & n4375 ;
  assign n4381 = ( n4341 & n4379 ) | ( n4341 & n4380 ) | ( n4379 & n4380 ) ;
  assign n4382 = ~n2823 & n4359 ;
  assign n4383 = ~n2764 & n4382 ;
  assign n4384 = ( n3071 & n4359 ) | ( n3071 & n4383 ) | ( n4359 & n4383 ) ;
  assign n4385 = ( n3326 & n4301 ) | ( n3326 & n4384 ) | ( n4301 & n4384 ) ;
  assign n4386 = n3326 | n4383 ;
  assign n4387 = n3326 | n4359 ;
  assign n4388 = ( n3071 & n4386 ) | ( n3071 & n4387 ) | ( n4386 & n4387 ) ;
  assign n4389 = ( n4300 & n4385 ) | ( n4300 & n4388 ) | ( n4385 & n4388 ) ;
  assign n4390 = ~n4380 & n4389 ;
  assign n4391 = ~n4379 & n4389 ;
  assign n4392 = ( ~n4341 & n4390 ) | ( ~n4341 & n4391 ) | ( n4390 & n4391 ) ;
  assign n4393 = ( n4378 & n4381 ) | ( n4378 & ~n4392 ) | ( n4381 & ~n4392 ) ;
  assign n4394 = n4296 & n4393 ;
  assign n4395 = n4268 & n4394 ;
  assign n4396 = ~n4130 & n4295 ;
  assign n4397 = ( ~n4130 & n4288 ) | ( ~n4130 & n4396 ) | ( n4288 & n4396 ) ;
  assign n4398 = n4103 | n4129 ;
  assign n4399 = n4393 & n4398 ;
  assign n4400 = ~n4130 & n4398 ;
  assign n4401 = ( n4397 & n4399 ) | ( n4397 & n4400 ) | ( n4399 & n4400 ) ;
  assign n4402 = ( n4268 & n4395 ) | ( n4268 & n4401 ) | ( n4395 & n4401 ) ;
  assign n4403 = n4263 & n4402 ;
  assign n4404 = n4054 | n4161 ;
  assign n4405 = ~n4162 & n4404 ;
  assign n4406 = n4268 | n4394 ;
  assign n4407 = n3856 & n4281 ;
  assign n4408 = n3063 & n3333 ;
  assign n4409 = n2368 & n3335 ;
  assign n4410 = ( ~n2340 & n3335 ) | ( ~n2340 & n4409 ) | ( n3335 & n4409 ) ;
  assign n4411 = ~n2679 & n4410 ;
  assign n4412 = n2827 & n4411 ;
  assign n4413 = ( n3057 & n3335 ) | ( n3057 & n4412 ) | ( n3335 & n4412 ) ;
  assign n4414 = n4408 | n4413 ;
  assign n4415 = ( n3049 & n3326 ) | ( n3049 & n4207 ) | ( n3326 & n4207 ) ;
  assign n4416 = n4414 | n4415 ;
  assign n4417 = n3049 & n3338 ;
  assign n4418 = ( ~n4299 & n4414 ) | ( ~n4299 & n4417 ) | ( n4414 & n4417 ) ;
  assign n4419 = n4299 | n4418 ;
  assign n4420 = ( n3856 & n4416 ) | ( n3856 & n4419 ) | ( n4416 & n4419 ) ;
  assign n4421 = ~n4407 & n4420 ;
  assign n4422 = n3049 & n4199 ;
  assign n4423 = ( n3326 & n4414 ) | ( n3326 & n4422 ) | ( n4414 & n4422 ) ;
  assign n4424 = n4421 & ~n4423 ;
  assign n4425 = n4401 & n4424 ;
  assign n4426 = ( n4406 & n4424 ) | ( n4406 & n4425 ) | ( n4424 & n4425 ) ;
  assign n4427 = n4405 | n4426 ;
  assign n4428 = n4263 | n4405 ;
  assign n4429 = ( n4403 & n4427 ) | ( n4403 & n4428 ) | ( n4427 & n4428 ) ;
  assign n4430 = n4263 | n4402 ;
  assign n4431 = ~n4157 & n4159 ;
  assign n4432 = ( n4157 & ~n4159 ) | ( n4157 & n4431 ) | ( ~n4159 & n4431 ) ;
  assign n4433 = ( n4426 & n4431 ) | ( n4426 & n4432 ) | ( n4431 & n4432 ) ;
  assign n4434 = n4431 | n4432 ;
  assign n4435 = ( n4430 & n4433 ) | ( n4430 & n4434 ) | ( n4433 & n4434 ) ;
  assign n4436 = n4429 | n4435 ;
  assign n4437 = n3049 & n3333 ;
  assign n4438 = n3110 & n3335 ;
  assign n4439 = ( ~n3106 & n3335 ) | ( ~n3106 & n4438 ) | ( n3335 & n4438 ) ;
  assign n4440 = n4437 | n4439 ;
  assign n4441 = n3033 & n4199 ;
  assign n4442 = ( n3326 & n4440 ) | ( n3326 & n4441 ) | ( n4440 & n4441 ) ;
  assign n4443 = ~n3624 & n4281 ;
  assign n4444 = ( n3033 & n3326 ) | ( n3033 & n4207 ) | ( n3326 & n4207 ) ;
  assign n4445 = n4440 | n4444 ;
  assign n4446 = n3338 | n4299 ;
  assign n4447 = ( n3033 & n4299 ) | ( n3033 & n4446 ) | ( n4299 & n4446 ) ;
  assign n4448 = n4440 | n4447 ;
  assign n4449 = ( ~n3624 & n4445 ) | ( ~n3624 & n4448 ) | ( n4445 & n4448 ) ;
  assign n4450 = ~n4443 & n4449 ;
  assign n4451 = ~n4442 & n4450 ;
  assign n4452 = n4436 & n4451 ;
  assign n4453 = n4163 & ~n4165 ;
  assign n4454 = ~n4163 & n4165 ;
  assign n4455 = n4453 | n4454 ;
  assign n4456 = n4405 & n4426 ;
  assign n4457 = n4263 & n4405 ;
  assign n4458 = ( n4403 & n4456 ) | ( n4403 & n4457 ) | ( n4456 & n4457 ) ;
  assign n4459 = ( n4405 & n4435 ) | ( n4405 & n4458 ) | ( n4435 & n4458 ) ;
  assign n4460 = n4455 | n4459 ;
  assign n4461 = n4452 | n4460 ;
  assign n4462 = n3033 & n3335 ;
  assign n4463 = n3110 & n3333 ;
  assign n4464 = ( ~n3106 & n3333 ) | ( ~n3106 & n4463 ) | ( n3333 & n4463 ) ;
  assign n4465 = n4462 | n4464 ;
  assign n4466 = n2916 & n3338 ;
  assign n4467 = ( ~n2901 & n3338 ) | ( ~n2901 & n4466 ) | ( n3338 & n4466 ) ;
  assign n4468 = ~n2921 & n4467 ;
  assign n4469 = n2828 & n4468 ;
  assign n4470 = ( n2927 & n3338 ) | ( n2927 & n4469 ) | ( n3338 & n4469 ) ;
  assign n4471 = n4465 | n4470 ;
  assign n4472 = n3326 & n4471 ;
  assign n4473 = n3952 & n4281 ;
  assign n4474 = n4299 | n4471 ;
  assign n4475 = n3326 | n4471 ;
  assign n4476 = ( n3952 & n4474 ) | ( n3952 & n4475 ) | ( n4474 & n4475 ) ;
  assign n4477 = ~n4473 & n4476 ;
  assign n4478 = ~n4472 & n4477 ;
  assign n4479 = n4461 & n4478 ;
  assign n4480 = n3997 & n4167 ;
  assign n4481 = n3997 | n4167 ;
  assign n4482 = ~n4480 & n4481 ;
  assign n4483 = n4455 & n4459 ;
  assign n4484 = ( n4452 & n4455 ) | ( n4452 & n4483 ) | ( n4455 & n4483 ) ;
  assign n4485 = n4482 | n4484 ;
  assign n4486 = n4479 | n4485 ;
  assign n4487 = n3033 & n3333 ;
  assign n4488 = n2916 & n3335 ;
  assign n4489 = ( ~n2901 & n3335 ) | ( ~n2901 & n4488 ) | ( n3335 & n4488 ) ;
  assign n4490 = ~n2921 & n4489 ;
  assign n4491 = n2828 & n4490 ;
  assign n4492 = ( n2927 & n3335 ) | ( n2927 & n4491 ) | ( n3335 & n4491 ) ;
  assign n4493 = n4487 | n4492 ;
  assign n4494 = n3024 & n4199 ;
  assign n4495 = ( n3326 & n4493 ) | ( n3326 & n4494 ) | ( n4493 & n4494 ) ;
  assign n4496 = n3896 & n4281 ;
  assign n4497 = ( n3024 & n3326 ) | ( n3024 & n4207 ) | ( n3326 & n4207 ) ;
  assign n4498 = n4493 | n4497 ;
  assign n4499 = ( n3024 & n4299 ) | ( n3024 & n4446 ) | ( n4299 & n4446 ) ;
  assign n4500 = n4493 | n4499 ;
  assign n4501 = ( n3896 & n4498 ) | ( n3896 & n4500 ) | ( n4498 & n4500 ) ;
  assign n4502 = ~n4496 & n4501 ;
  assign n4503 = ~n4495 & n4502 ;
  assign n4504 = n4486 & n4503 ;
  assign n4505 = n4482 & n4484 ;
  assign n4506 = ( n4479 & n4482 ) | ( n4479 & n4505 ) | ( n4482 & n4505 ) ;
  assign n4507 = n4241 & n4506 ;
  assign n4508 = ( n4241 & n4504 ) | ( n4241 & n4507 ) | ( n4504 & n4507 ) ;
  assign n4509 = n4237 | n4508 ;
  assign n4510 = n3925 & n3970 ;
  assign n4511 = ( n3924 & n3970 ) | ( n3924 & n4510 ) | ( n3970 & n4510 ) ;
  assign n4512 = n3926 & ~n4511 ;
  assign n4513 = ~n3925 & n3970 ;
  assign n4514 = ~n3924 & n4513 ;
  assign n4515 = n4512 | n4514 ;
  assign n4516 = ( n3947 & n3949 ) | ( n3947 & n4170 ) | ( n3949 & n4170 ) ;
  assign n4517 = n4515 | n4516 ;
  assign n4518 = n4515 & ~n4516 ;
  assign n4519 = ( ~n4515 & n4517 ) | ( ~n4515 & n4518 ) | ( n4517 & n4518 ) ;
  assign n4520 = n4241 | n4506 ;
  assign n4521 = n4504 | n4520 ;
  assign n4522 = n4519 | n4521 ;
  assign n4523 = ( n4509 & n4519 ) | ( n4509 & n4522 ) | ( n4519 & n4522 ) ;
  assign n4524 = n4213 & n4523 ;
  assign n4525 = ( n3127 & ~n3310 ) | ( n3127 & n3313 ) | ( ~n3310 & n3313 ) ;
  assign n4526 = n3269 | n3310 ;
  assign n4527 = ~n3269 & n3313 ;
  assign n4528 = ( n3127 & ~n4526 ) | ( n3127 & n4527 ) | ( ~n4526 & n4527 ) ;
  assign n4529 = n3269 | n4527 ;
  assign n4530 = ~n3269 & n3310 ;
  assign n4531 = ( n3127 & n4529 ) | ( n3127 & ~n4530 ) | ( n4529 & ~n4530 ) ;
  assign n4532 = ( ~n4525 & n4528 ) | ( ~n4525 & n4531 ) | ( n4528 & n4531 ) ;
  assign n4533 = n3259 & n3338 ;
  assign n4534 = n3266 & n3335 ;
  assign n4535 = n3296 & n3333 ;
  assign n4536 = n3295 & n3333 ;
  assign n4537 = ( n2828 & n4535 ) | ( n2828 & n4536 ) | ( n4535 & n4536 ) ;
  assign n4538 = ( ~n3300 & n3333 ) | ( ~n3300 & n4537 ) | ( n3333 & n4537 ) ;
  assign n4539 = n4534 | n4538 ;
  assign n4540 = n4533 | n4539 ;
  assign n4541 = ( n3340 & n4532 ) | ( n3340 & n4540 ) | ( n4532 & n4540 ) ;
  assign n4542 = ( n3326 & n3340 ) | ( n3326 & ~n4540 ) | ( n3340 & ~n4540 ) ;
  assign n4543 = ( n3326 & n4532 ) | ( n3326 & n4542 ) | ( n4532 & n4542 ) ;
  assign n4544 = ~n4541 & n4543 ;
  assign n4545 = n4540 | n4542 ;
  assign n4546 = n3326 | n4540 ;
  assign n4547 = ( n4532 & n4545 ) | ( n4532 & n4546 ) | ( n4545 & n4546 ) ;
  assign n4548 = ( ~n3326 & n4544 ) | ( ~n3326 & n4547 ) | ( n4544 & n4547 ) ;
  assign n4549 = n4519 & n4521 ;
  assign n4550 = n4509 & n4549 ;
  assign n4551 = n4548 & n4550 ;
  assign n4552 = ( n4524 & n4548 ) | ( n4524 & n4551 ) | ( n4548 & n4551 ) ;
  assign n4553 = n4182 & n4552 ;
  assign n4554 = ~n3922 & n4174 ;
  assign n4555 = n4548 | n4550 ;
  assign n4556 = n4524 | n4555 ;
  assign n4557 = ( n3922 & ~n4174 ) | ( n3922 & n4554 ) | ( ~n4174 & n4554 ) ;
  assign n4558 = ( n4554 & n4556 ) | ( n4554 & n4557 ) | ( n4556 & n4557 ) ;
  assign n4559 = ( n4182 & n4553 ) | ( n4182 & n4558 ) | ( n4553 & n4558 ) ;
  assign n4560 = n3259 & n3380 ;
  assign n4561 = n3266 & n3367 ;
  assign n4562 = n3296 & n3373 ;
  assign n4563 = n3295 & n3373 ;
  assign n4564 = ( n2828 & n4562 ) | ( n2828 & n4563 ) | ( n4562 & n4563 ) ;
  assign n4565 = ( ~n3300 & n3373 ) | ( ~n3300 & n4564 ) | ( n3373 & n4564 ) ;
  assign n4566 = n4561 | n4565 ;
  assign n4567 = n4560 | n4566 ;
  assign n4568 = ( n1115 & n4035 ) | ( n1115 & n4567 ) | ( n4035 & n4567 ) ;
  assign n4569 = n1115 & n4567 ;
  assign n4570 = ( n4532 & n4568 ) | ( n4532 & n4569 ) | ( n4568 & n4569 ) ;
  assign n4571 = n4043 | n4567 ;
  assign n4572 = n1115 | n4567 ;
  assign n4573 = ( n4532 & n4571 ) | ( n4532 & n4572 ) | ( n4571 & n4572 ) ;
  assign n4574 = ~n4570 & n4573 ;
  assign n4575 = n2368 & n3412 ;
  assign n4576 = ( ~n2340 & n3412 ) | ( ~n2340 & n4575 ) | ( n3412 & n4575 ) ;
  assign n4577 = ~n2679 & n4576 ;
  assign n4578 = n2827 & n4577 ;
  assign n4579 = ( n3057 & n3412 ) | ( n3057 & n4578 ) | ( n3412 & n4578 ) ;
  assign n4580 = n3049 & n3414 ;
  assign n4581 = n4579 | n4580 ;
  assign n4582 = n3110 & n3417 ;
  assign n4583 = ( ~n3106 & n3417 ) | ( ~n3106 & n4582 ) | ( n3417 & n4582 ) ;
  assign n4584 = n3423 | n4583 ;
  assign n4585 = n4581 | n4584 ;
  assign n4586 = n634 & n4585 ;
  assign n4587 = n634 & n4583 ;
  assign n4588 = ( n634 & n4581 ) | ( n634 & n4587 ) | ( n4581 & n4587 ) ;
  assign n4589 = ( ~n3679 & n4586 ) | ( ~n3679 & n4588 ) | ( n4586 & n4588 ) ;
  assign n4590 = n634 | n4585 ;
  assign n4591 = n634 | n4583 ;
  assign n4592 = n4581 | n4591 ;
  assign n4593 = ( ~n3679 & n4590 ) | ( ~n3679 & n4592 ) | ( n4590 & n4592 ) ;
  assign n4594 = ~n4589 & n4593 ;
  assign n4595 = n879 & n3085 ;
  assign n4596 = n3466 & n4595 ;
  assign n4597 = n3470 & n4595 ;
  assign n4598 = ~n3458 & n4597 ;
  assign n4599 = ( n3464 & n4596 ) | ( n3464 & n4598 ) | ( n4596 & n4598 ) ;
  assign n4600 = n3496 & n4599 ;
  assign n4601 = n3471 | n4595 ;
  assign n4602 = n3466 | n4595 ;
  assign n4603 = ( n3464 & n4601 ) | ( n3464 & n4602 ) | ( n4601 & n4602 ) ;
  assign n4604 = ( n3496 & n4595 ) | ( n3496 & n4603 ) | ( n4595 & n4603 ) ;
  assign n4605 = ~n4600 & n4604 ;
  assign n4606 = n3078 & n3477 ;
  assign n4607 = ( n3082 & n3477 ) | ( n3082 & n4606 ) | ( n3477 & n4606 ) ;
  assign n4608 = n3448 | n4607 ;
  assign n4609 = ( n3070 & n4607 ) | ( n3070 & n4608 ) | ( n4607 & n4608 ) ;
  assign n4610 = ~n2823 & n3446 ;
  assign n4611 = ~n2764 & n4610 ;
  assign n4612 = ( n3071 & n3446 ) | ( n3071 & n4611 ) | ( n3446 & n4611 ) ;
  assign n4613 = n4609 | n4612 ;
  assign n4614 = ( n3452 & n3821 ) | ( n3452 & n4613 ) | ( n3821 & n4613 ) ;
  assign n4615 = n3452 | n4612 ;
  assign n4616 = n4609 | n4615 ;
  assign n4617 = ( ~n3583 & n4614 ) | ( ~n3583 & n4616 ) | ( n4614 & n4616 ) ;
  assign n4618 = ( n879 & n4613 ) | ( n879 & ~n4617 ) | ( n4613 & ~n4617 ) ;
  assign n4619 = n4617 | n4618 ;
  assign n4620 = n879 & ~n4612 ;
  assign n4621 = ~n4609 & n4620 ;
  assign n4622 = ~n4617 & n4621 ;
  assign n4623 = ( ~n879 & n4619 ) | ( ~n879 & n4622 ) | ( n4619 & n4622 ) ;
  assign n4624 = n4605 & n4623 ;
  assign n4625 = n4600 | n4624 ;
  assign n4626 = n3063 & n3448 ;
  assign n4627 = n3070 & n3446 ;
  assign n4628 = ~n2823 & n3477 ;
  assign n4629 = ~n2764 & n4628 ;
  assign n4630 = n3452 | n4629 ;
  assign n4631 = ( n3071 & n3487 ) | ( n3071 & n4630 ) | ( n3487 & n4630 ) ;
  assign n4632 = n4627 | n4631 ;
  assign n4633 = n4626 | n4632 ;
  assign n4634 = n879 & n4633 ;
  assign n4635 = n879 & n4629 ;
  assign n4636 = n879 & n3477 ;
  assign n4637 = ( n3071 & n4635 ) | ( n3071 & n4636 ) | ( n4635 & n4636 ) ;
  assign n4638 = ( n879 & n4627 ) | ( n879 & n4637 ) | ( n4627 & n4637 ) ;
  assign n4639 = n879 | n4637 ;
  assign n4640 = ( n4626 & n4638 ) | ( n4626 & n4639 ) | ( n4638 & n4639 ) ;
  assign n4641 = ( n3510 & n4634 ) | ( n3510 & n4640 ) | ( n4634 & n4640 ) ;
  assign n4642 = n4634 & n4640 ;
  assign n4643 = ( ~n3094 & n4641 ) | ( ~n3094 & n4642 ) | ( n4641 & n4642 ) ;
  assign n4644 = n879 | n4633 ;
  assign n4645 = n879 | n4629 ;
  assign n4646 = n879 | n3477 ;
  assign n4647 = ( n3071 & n4645 ) | ( n3071 & n4646 ) | ( n4645 & n4646 ) ;
  assign n4648 = n4627 | n4647 ;
  assign n4649 = n4626 | n4648 ;
  assign n4650 = ( n3510 & n4644 ) | ( n3510 & n4649 ) | ( n4644 & n4649 ) ;
  assign n4651 = n4644 & n4649 ;
  assign n4652 = ( ~n3094 & n4650 ) | ( ~n3094 & n4651 ) | ( n4650 & n4651 ) ;
  assign n4653 = ~n4643 & n4652 ;
  assign n4654 = n879 & n3078 ;
  assign n4655 = ( n879 & n3082 ) | ( n879 & n4654 ) | ( n3082 & n4654 ) ;
  assign n4656 = ~n879 & n4655 ;
  assign n4657 = ( ~n4633 & n4655 ) | ( ~n4633 & n4656 ) | ( n4655 & n4656 ) ;
  assign n4658 = ~n4640 & n4655 ;
  assign n4659 = ( ~n3510 & n4657 ) | ( ~n3510 & n4658 ) | ( n4657 & n4658 ) ;
  assign n4660 = n4657 | n4658 ;
  assign n4661 = ( n3094 & n4659 ) | ( n3094 & n4660 ) | ( n4659 & n4660 ) ;
  assign n4662 = n4655 & ~n4661 ;
  assign n4663 = n4661 & ~n4662 ;
  assign n4664 = ( n4653 & n4662 ) | ( n4653 & ~n4663 ) | ( n4662 & ~n4663 ) ;
  assign n4665 = n4625 & n4664 ;
  assign n4666 = n4625 & ~n4665 ;
  assign n4667 = ~n4625 & n4664 ;
  assign n4669 = n4594 & n4667 ;
  assign n4670 = ( n4594 & n4666 ) | ( n4594 & n4669 ) | ( n4666 & n4669 ) ;
  assign n4668 = n4666 | n4667 ;
  assign n4671 = n4668 & ~n4670 ;
  assign n4672 = ( n4594 & ~n4670 ) | ( n4594 & n4671 ) | ( ~n4670 & n4671 ) ;
  assign n4673 = n4605 & ~n4623 ;
  assign n4674 = ~n4605 & n4623 ;
  assign n4675 = n4673 | n4674 ;
  assign n4676 = n3063 & n3412 ;
  assign n4677 = n2368 & n3414 ;
  assign n4678 = ( ~n2340 & n3414 ) | ( ~n2340 & n4677 ) | ( n3414 & n4677 ) ;
  assign n4679 = ~n2679 & n4678 ;
  assign n4680 = n2827 & n4679 ;
  assign n4681 = ( n3057 & n3414 ) | ( n3057 & n4680 ) | ( n3414 & n4680 ) ;
  assign n4682 = n4676 | n4681 ;
  assign n4683 = n3417 | n3423 ;
  assign n4684 = ( n3049 & n3423 ) | ( n3049 & n4683 ) | ( n3423 & n4683 ) ;
  assign n4685 = n4682 | n4684 ;
  assign n4686 = n634 & n4685 ;
  assign n4687 = n634 & n3417 ;
  assign n4688 = n3049 & n4687 ;
  assign n4689 = ( n634 & n4682 ) | ( n634 & n4688 ) | ( n4682 & n4688 ) ;
  assign n4690 = ( n3856 & n4686 ) | ( n3856 & n4689 ) | ( n4686 & n4689 ) ;
  assign n4691 = n634 | n4685 ;
  assign n4692 = n634 | n3417 ;
  assign n4693 = ( n634 & n3049 ) | ( n634 & n4692 ) | ( n3049 & n4692 ) ;
  assign n4694 = n4682 | n4693 ;
  assign n4695 = ( n3856 & n4691 ) | ( n3856 & n4694 ) | ( n4691 & n4694 ) ;
  assign n4696 = ~n4690 & n4695 ;
  assign n4697 = n4675 & n4696 ;
  assign n4698 = n4675 & ~n4697 ;
  assign n4699 = n3500 | n3613 ;
  assign n4700 = ~n4675 & n4696 ;
  assign n4701 = n3500 & n4700 ;
  assign n4702 = ( n3613 & n4700 ) | ( n3613 & n4701 ) | ( n4700 & n4701 ) ;
  assign n4703 = ( n4698 & n4699 ) | ( n4698 & n4702 ) | ( n4699 & n4702 ) ;
  assign n4704 = n4697 | n4703 ;
  assign n4705 = ~n4672 & n4704 ;
  assign n4706 = n4672 & ~n4704 ;
  assign n4707 = n4705 | n4706 ;
  assign n4708 = n3033 & n3635 ;
  assign n4709 = n2916 & n3637 ;
  assign n4710 = ( ~n2901 & n3637 ) | ( ~n2901 & n4709 ) | ( n3637 & n4709 ) ;
  assign n4711 = ~n2921 & n4710 ;
  assign n4712 = n2828 & n4711 ;
  assign n4713 = ( n2927 & n3637 ) | ( n2927 & n4712 ) | ( n3637 & n4712 ) ;
  assign n4714 = n4708 | n4713 ;
  assign n4715 = n3024 & n3641 ;
  assign n4716 = ( n3024 & n3643 ) | ( n3024 & n3644 ) | ( n3643 & n3644 ) ;
  assign n4717 = n4715 & n4716 ;
  assign n4718 = n4714 | n4717 ;
  assign n4719 = n482 | n4718 ;
  assign n4720 = ( n3024 & n3649 ) | ( n3024 & n3650 ) | ( n3649 & n3650 ) ;
  assign n4721 = n4714 | n4720 ;
  assign n4722 = ( n3896 & n4719 ) | ( n3896 & n4721 ) | ( n4719 & n4721 ) ;
  assign n4723 = n482 & n4718 ;
  assign n4724 = ( n3024 & n3656 ) | ( n3024 & n3657 ) | ( n3656 & n3657 ) ;
  assign n4725 = ( n482 & n4714 ) | ( n482 & n4724 ) | ( n4714 & n4724 ) ;
  assign n4726 = ( n3896 & n4723 ) | ( n3896 & n4725 ) | ( n4723 & n4725 ) ;
  assign n4727 = n4722 & ~n4726 ;
  assign n4728 = n4707 & n4727 ;
  assign n4729 = n4707 | n4727 ;
  assign n4730 = ~n4728 & n4729 ;
  assign n4731 = n3500 | n4700 ;
  assign n4732 = n3613 | n4731 ;
  assign n4733 = n4698 | n4732 ;
  assign n4734 = ~n4703 & n4733 ;
  assign n4735 = n3033 & n3637 ;
  assign n4736 = n3110 & n3635 ;
  assign n4737 = ( ~n3106 & n3635 ) | ( ~n3106 & n4736 ) | ( n3635 & n4736 ) ;
  assign n4738 = n4735 | n4737 ;
  assign n4739 = n2916 & n3641 ;
  assign n4740 = ( ~n2901 & n3641 ) | ( ~n2901 & n4739 ) | ( n3641 & n4739 ) ;
  assign n4741 = ~n2921 & n4740 ;
  assign n4742 = n2828 & n4741 ;
  assign n4743 = ( n2927 & n3641 ) | ( n2927 & n4742 ) | ( n3641 & n4742 ) ;
  assign n4744 = n4738 | n4743 ;
  assign n4745 = n3643 | n4744 ;
  assign n4746 = n482 & n4744 ;
  assign n4747 = n4745 & n4746 ;
  assign n4748 = ( n482 & n3656 ) | ( n482 & n4744 ) | ( n3656 & n4744 ) ;
  assign n4749 = ( n3952 & n4747 ) | ( n3952 & n4748 ) | ( n4747 & n4748 ) ;
  assign n4750 = n482 | n4744 ;
  assign n4751 = n3650 | n4744 ;
  assign n4752 = ( n3952 & n4750 ) | ( n3952 & n4751 ) | ( n4750 & n4751 ) ;
  assign n4753 = ~n4749 & n4752 ;
  assign n4754 = n4734 & n4753 ;
  assign n4755 = n4734 & ~n4754 ;
  assign n4756 = ( n4753 & ~n4754 ) | ( n4753 & n4755 ) | ( ~n4754 & n4755 ) ;
  assign n4757 = ( n3615 & n3661 ) | ( n3615 & n3883 ) | ( n3661 & n3883 ) ;
  assign n4758 = n4754 | n4757 ;
  assign n4759 = ( n4754 & n4756 ) | ( n4754 & n4758 ) | ( n4756 & n4758 ) ;
  assign n4760 = n4730 & n4759 ;
  assign n4761 = n4730 | n4759 ;
  assign n4762 = ~n4760 & n4761 ;
  assign n4763 = n4574 & n4762 ;
  assign n4764 = n4574 | n4762 ;
  assign n4765 = ~n4763 & n4764 ;
  assign n4766 = n3024 & n3373 ;
  assign n4767 = n3296 & n3367 ;
  assign n4768 = n3295 & n3367 ;
  assign n4769 = ( n2828 & n4767 ) | ( n2828 & n4768 ) | ( n4767 & n4768 ) ;
  assign n4770 = ( ~n3300 & n3367 ) | ( ~n3300 & n4769 ) | ( n3367 & n4769 ) ;
  assign n4771 = n4766 | n4770 ;
  assign n4772 = ~n3371 & n4034 ;
  assign n4773 = n3266 & n4772 ;
  assign n4774 = ( n1115 & n4771 ) | ( n1115 & n4773 ) | ( n4771 & n4773 ) ;
  assign n4775 = ( n3266 & n3388 ) | ( n3266 & n3915 ) | ( n3388 & n3915 ) ;
  assign n4776 = ( n1115 & n4771 ) | ( n1115 & n4775 ) | ( n4771 & n4775 ) ;
  assign n4777 = ( ~n4190 & n4774 ) | ( ~n4190 & n4776 ) | ( n4774 & n4776 ) ;
  assign n4778 = ( n1115 & ~n3371 ) | ( n1115 & n4042 ) | ( ~n3371 & n4042 ) ;
  assign n4779 = ( n1115 & n3266 ) | ( n1115 & n4778 ) | ( n3266 & n4778 ) ;
  assign n4780 = n4771 | n4779 ;
  assign n4781 = ( n3266 & n3394 ) | ( n3266 & n3910 ) | ( n3394 & n3910 ) ;
  assign n4782 = n4771 | n4781 ;
  assign n4783 = ( ~n4190 & n4780 ) | ( ~n4190 & n4782 ) | ( n4780 & n4782 ) ;
  assign n4784 = ~n4777 & n4783 ;
  assign n4785 = n4756 & n4757 ;
  assign n4786 = n4756 & ~n4785 ;
  assign n4787 = n4757 & n4784 ;
  assign n4788 = ~n4756 & n4787 ;
  assign n4789 = ( n4784 & n4786 ) | ( n4784 & n4788 ) | ( n4786 & n4788 ) ;
  assign n4790 = ~n4756 & n4757 ;
  assign n4791 = n4786 | n4790 ;
  assign n4792 = ~n4789 & n4791 ;
  assign n4793 = n3665 & n3883 ;
  assign n4794 = n3883 & ~n4793 ;
  assign n4795 = n3398 & n3664 ;
  assign n4796 = ( n3398 & n3663 ) | ( n3398 & n4795 ) | ( n3663 & n4795 ) ;
  assign n4797 = ~n3883 & n4796 ;
  assign n4798 = ( n3398 & n4794 ) | ( n3398 & n4797 ) | ( n4794 & n4797 ) ;
  assign n4799 = n3886 | n4798 ;
  assign n4800 = ( n4176 & n4798 ) | ( n4176 & n4799 ) | ( n4798 & n4799 ) ;
  assign n4801 = ~n4757 & n4784 ;
  assign n4802 = ( n4756 & n4784 ) | ( n4756 & n4801 ) | ( n4784 & n4801 ) ;
  assign n4803 = ~n4786 & n4802 ;
  assign n4804 = n4800 & n4803 ;
  assign n4805 = ( n4792 & n4800 ) | ( n4792 & n4804 ) | ( n4800 & n4804 ) ;
  assign n4806 = n4789 | n4805 ;
  assign n4807 = n4765 & n4806 ;
  assign n4808 = n4765 | n4806 ;
  assign n4809 = ~n4807 & n4808 ;
  assign n4810 = n257 | n1034 ;
  assign n4811 = n742 | n746 ;
  assign n4812 = n739 | n4811 ;
  assign n4813 = n4810 | n4812 ;
  assign n4814 = n724 | n891 ;
  assign n4815 = n960 | n4814 ;
  assign n4816 = n862 | n4815 ;
  assign n4817 = n268 | n907 ;
  assign n4818 = n917 | n4817 ;
  assign n4819 = n541 | n4818 ;
  assign n4820 = n4816 | n4819 ;
  assign n4821 = n4813 | n4820 ;
  assign n4822 = n183 | n348 ;
  assign n4823 = n397 | n4822 ;
  assign n4824 = n732 | n4823 ;
  assign n4825 = n4821 | n4824 ;
  assign n4826 = n3285 & n4825 ;
  assign n4827 = n3222 & n4826 ;
  assign n4828 = ~n3285 & n4825 ;
  assign n4829 = ( ~n3222 & n4825 ) | ( ~n3222 & n4828 ) | ( n4825 & n4828 ) ;
  assign n4830 = ( n3286 & ~n4827 ) | ( n3286 & n4829 ) | ( ~n4827 & n4829 ) ;
  assign n4831 = ~n3289 & n4830 ;
  assign n4832 = n3289 & ~n4830 ;
  assign n4833 = n4831 | n4832 ;
  assign n4834 = ~n4831 & n4833 ;
  assign n4835 = ~n3290 & n3292 ;
  assign n4836 = ( n3270 & n3290 ) | ( n3270 & ~n4835 ) | ( n3290 & ~n4835 ) ;
  assign n4837 = n3267 | n3290 ;
  assign n4838 = ( n3290 & ~n3292 ) | ( n3290 & n4837 ) | ( ~n3292 & n4837 ) ;
  assign n4839 = ( ~n3310 & n4836 ) | ( ~n3310 & n4838 ) | ( n4836 & n4838 ) ;
  assign n4840 = ( n3313 & n4836 ) | ( n3313 & n4838 ) | ( n4836 & n4838 ) ;
  assign n4841 = ( n3127 & n4839 ) | ( n3127 & n4840 ) | ( n4839 & n4840 ) ;
  assign n4842 = ( n4831 & ~n4834 ) | ( n4831 & n4841 ) | ( ~n4834 & n4841 ) ;
  assign n4843 = n1024 | n1026 ;
  assign n4844 = n161 | n257 ;
  assign n4845 = n167 | n4844 ;
  assign n4846 = n1034 | n4845 ;
  assign n4847 = n4843 | n4846 ;
  assign n4848 = n4812 | n4847 ;
  assign n4849 = n889 | n914 ;
  assign n4850 = n177 | n4849 ;
  assign n4851 = n4848 | n4850 ;
  assign n4852 = n256 | n718 ;
  assign n4853 = n4851 | n4852 ;
  assign n4854 = ( n3286 & n4827 ) | ( n3286 & n4853 ) | ( n4827 & n4853 ) ;
  assign n4855 = ( n4827 & n4853 ) | ( n4827 & ~n4854 ) | ( n4853 & ~n4854 ) ;
  assign n4856 = ~n4830 & n4854 ;
  assign n4857 = n3286 | n4830 ;
  assign n4858 = ( n4855 & ~n4856 ) | ( n4855 & n4857 ) | ( ~n4856 & n4857 ) ;
  assign n4859 = n4830 & ~n4854 ;
  assign n4860 = n3286 & n4830 ;
  assign n4861 = ( n4855 & n4859 ) | ( n4855 & n4860 ) | ( n4859 & n4860 ) ;
  assign n4862 = n4858 & ~n4861 ;
  assign n4863 = n4834 | n4862 ;
  assign n4864 = n4831 & ~n4862 ;
  assign n4865 = ( n4841 & ~n4863 ) | ( n4841 & n4864 ) | ( ~n4863 & n4864 ) ;
  assign n4866 = n4862 | n4864 ;
  assign n4867 = ~n4862 & n4863 ;
  assign n4868 = ( n4841 & n4866 ) | ( n4841 & ~n4867 ) | ( n4866 & ~n4867 ) ;
  assign n4869 = ( ~n4842 & n4865 ) | ( ~n4842 & n4868 ) | ( n4865 & n4868 ) ;
  assign n4870 = ~n3289 & n3333 ;
  assign n4871 = n3335 & n4830 ;
  assign n4872 = n4870 | n4871 ;
  assign n4873 = ( n3340 & n3341 ) | ( n3340 & ~n4854 ) | ( n3341 & ~n4854 ) ;
  assign n4874 = ( n3285 & n3340 ) | ( n3285 & n3341 ) | ( n3340 & n3341 ) ;
  assign n4875 = n3340 & n3341 ;
  assign n4876 = ( n3222 & n4874 ) | ( n3222 & n4875 ) | ( n4874 & n4875 ) ;
  assign n4877 = ( n4855 & n4873 ) | ( n4855 & n4876 ) | ( n4873 & n4876 ) ;
  assign n4878 = n4872 | n4877 ;
  assign n4879 = n3326 | n4878 ;
  assign n4880 = n3338 & ~n4854 ;
  assign n4881 = n3285 & n3338 ;
  assign n4882 = n3222 & n4881 ;
  assign n4883 = ( n4855 & n4880 ) | ( n4855 & n4882 ) | ( n4880 & n4882 ) ;
  assign n4884 = n4877 & n4883 ;
  assign n4885 = n3326 | n4872 ;
  assign n4886 = n4884 | n4885 ;
  assign n4887 = ( n4869 & n4879 ) | ( n4869 & n4886 ) | ( n4879 & n4886 ) ;
  assign n4888 = n3326 & n4878 ;
  assign n4889 = n3326 & n4872 ;
  assign n4890 = ( n3326 & n4884 ) | ( n3326 & n4889 ) | ( n4884 & n4889 ) ;
  assign n4891 = ( n4869 & n4888 ) | ( n4869 & n4890 ) | ( n4888 & n4890 ) ;
  assign n4892 = n4887 & ~n4891 ;
  assign n4893 = n4809 & n4892 ;
  assign n4894 = n4809 | n4892 ;
  assign n4895 = ~n4893 & n4894 ;
  assign n4896 = n4800 | n4803 ;
  assign n4897 = n4792 | n4896 ;
  assign n4898 = ~n4805 & n4897 ;
  assign n4899 = ~n4833 & n4841 ;
  assign n4900 = n4833 & ~n4841 ;
  assign n4901 = n4899 | n4900 ;
  assign n4902 = n3259 & n3333 ;
  assign n4903 = ~n3289 & n3335 ;
  assign n4904 = n4902 | n4903 ;
  assign n4905 = n3338 & n4830 ;
  assign n4906 = ( n3340 & n3341 ) | ( n3340 & n4830 ) | ( n3341 & n4830 ) ;
  assign n4907 = n4905 & n4906 ;
  assign n4908 = n4904 | n4907 ;
  assign n4909 = n3326 | n4908 ;
  assign n4910 = ( n3346 & n3347 ) | ( n3346 & n4830 ) | ( n3347 & n4830 ) ;
  assign n4911 = n4904 | n4910 ;
  assign n4912 = ( ~n4901 & n4909 ) | ( ~n4901 & n4911 ) | ( n4909 & n4911 ) ;
  assign n4913 = n3326 & n4908 ;
  assign n4914 = ( n3352 & n3353 ) | ( n3352 & n4830 ) | ( n3353 & n4830 ) ;
  assign n4915 = ( n3326 & n4904 ) | ( n3326 & n4914 ) | ( n4904 & n4914 ) ;
  assign n4916 = ( ~n4901 & n4913 ) | ( ~n4901 & n4915 ) | ( n4913 & n4915 ) ;
  assign n4917 = n4912 & ~n4916 ;
  assign n4918 = n4898 | n4917 ;
  assign n4919 = n4895 | n4918 ;
  assign n4920 = ( n4180 & n4898 ) | ( n4180 & n4917 ) | ( n4898 & n4917 ) ;
  assign n4921 = n4895 | n4920 ;
  assign n4922 = ( n4559 & n4919 ) | ( n4559 & n4921 ) | ( n4919 & n4921 ) ;
  assign n4923 = n4895 & n4918 ;
  assign n4924 = n4895 & n4920 ;
  assign n4925 = ( n4559 & n4923 ) | ( n4559 & n4924 ) | ( n4923 & n4924 ) ;
  assign n4926 = n4922 & ~n4925 ;
  assign n4927 = n206 | n455 ;
  assign n4928 = n501 | n858 ;
  assign n4929 = n3238 | n4928 ;
  assign n4930 = n233 | n4929 ;
  assign n4931 = n4927 | n4930 ;
  assign n4932 = n261 | n2731 ;
  assign n4933 = n4931 | n4932 ;
  assign n4936 = n387 | n428 ;
  assign n4937 = n165 | n256 ;
  assign n4938 = n4936 | n4937 ;
  assign n4939 = n139 | n235 ;
  assign n4940 = n229 | n4939 ;
  assign n4941 = n4938 | n4940 ;
  assign n4934 = n185 | n689 ;
  assign n4935 = n134 | n141 ;
  assign n4942 = ( n4934 & n4935 ) | ( n4934 & ~n4941 ) | ( n4935 & ~n4941 ) ;
  assign n4943 = n4941 | n4942 ;
  assign n4944 = n245 | n3231 ;
  assign n4945 = n594 | n3175 ;
  assign n4946 = n4944 | n4945 ;
  assign n4947 = n155 | n283 ;
  assign n4948 = n189 | n267 ;
  assign n4949 = n4947 | n4948 ;
  assign n4950 = n361 | n718 ;
  assign n4951 = n4949 | n4950 ;
  assign n4952 = n125 | n248 ;
  assign n4953 = n2549 | n4952 ;
  assign n4954 = n254 | n4953 ;
  assign n4955 = n4951 | n4954 ;
  assign n4956 = n4946 | n4955 ;
  assign n4957 = n4943 | n4956 ;
  assign n4958 = n4933 | n4957 ;
  assign n4959 = n299 | n353 ;
  assign n4960 = n232 | n333 ;
  assign n4961 = n4959 | n4960 ;
  assign n4962 = n344 | n408 ;
  assign n4963 = n249 | n4962 ;
  assign n4964 = n4961 | n4963 ;
  assign n4965 = n4958 | n4964 ;
  assign n4966 = n4926 & n4965 ;
  assign n4967 = n4926 & ~n4966 ;
  assign n4968 = n4898 & n4917 ;
  assign n4969 = n4898 & ~n4968 ;
  assign n4970 = n3357 | n4917 ;
  assign n4971 = ( n4179 & n4917 ) | ( n4179 & n4970 ) | ( n4917 & n4970 ) ;
  assign n4972 = ( n4180 & ~n4898 ) | ( n4180 & n4971 ) | ( ~n4898 & n4971 ) ;
  assign n4973 = n4969 | n4972 ;
  assign n4974 = n4559 | n4973 ;
  assign n4975 = ~n4898 & n4917 ;
  assign n4976 = n4969 | n4975 ;
  assign n4977 = n4180 & n4975 ;
  assign n4978 = ( n4180 & n4969 ) | ( n4180 & n4977 ) | ( n4969 & n4977 ) ;
  assign n4979 = ( n4559 & n4976 ) | ( n4559 & n4978 ) | ( n4976 & n4978 ) ;
  assign n4980 = n4974 & ~n4979 ;
  assign n4981 = n4182 | n4552 ;
  assign n4982 = n4558 | n4981 ;
  assign n4983 = ~n4559 & n4982 ;
  assign n4984 = n260 | n319 ;
  assign n4985 = n197 | n495 ;
  assign n4986 = n3173 | n4985 ;
  assign n4987 = n4984 | n4986 ;
  assign n4988 = n723 | n2737 ;
  assign n4989 = n677 | n2723 ;
  assign n4990 = n4988 | n4989 ;
  assign n4991 = n292 | n4990 ;
  assign n4992 = n4987 | n4991 ;
  assign n4993 = n206 | n2319 ;
  assign n4994 = n330 | n841 ;
  assign n4995 = n321 | n907 ;
  assign n4996 = n2596 | n4995 ;
  assign n4997 = n4994 | n4996 ;
  assign n4998 = n4993 | n4997 ;
  assign n4999 = n223 | n253 ;
  assign n5000 = n278 | n290 ;
  assign n5001 = n4999 | n5000 ;
  assign n5002 = n2665 | n5001 ;
  assign n5003 = n4998 | n5002 ;
  assign n5004 = n4992 | n5003 ;
  assign n5005 = ( n182 & n452 ) | ( n182 & ~n4937 ) | ( n452 & ~n4937 ) ;
  assign n5006 = n4937 | n5005 ;
  assign n5007 = n5004 | n5006 ;
  assign n5008 = n4983 & n5007 ;
  assign n5009 = n173 | n372 ;
  assign n5010 = n332 | n5009 ;
  assign n5011 = n2780 | n5010 ;
  assign n5012 = n220 | n408 ;
  assign n5013 = n340 | n5012 ;
  assign n5014 = n277 | n369 ;
  assign n5015 = n5013 | n5014 ;
  assign n5016 = n241 | n290 ;
  assign n5017 = n198 | n357 ;
  assign n5018 = n5016 | n5017 ;
  assign n5019 = n257 | n266 ;
  assign n5020 = n172 | n249 ;
  assign n5021 = n5019 | n5020 ;
  assign n5022 = n5018 | n5021 ;
  assign n5023 = n5015 | n5022 ;
  assign n5024 = n5011 | n5023 ;
  assign n5025 = n304 | n985 ;
  assign n5026 = n229 | n296 ;
  assign n5027 = n2639 | n5026 ;
  assign n5028 = n217 | n570 ;
  assign n5029 = n212 | n456 ;
  assign n5030 = n5028 | n5029 ;
  assign n5031 = n139 | n205 ;
  assign n5032 = n5030 | n5031 ;
  assign n5033 = n5027 | n5032 ;
  assign n5034 = n5025 | n5033 ;
  assign n5035 = n5024 | n5034 ;
  assign n5036 = n193 | n197 ;
  assign n5037 = n590 | n5036 ;
  assign n5038 = n316 | n579 ;
  assign n5039 = n5037 | n5038 ;
  assign n5040 = n262 | n495 ;
  assign n5041 = n244 | n511 ;
  assign n5042 = n5040 | n5041 ;
  assign n5043 = n5039 | n5042 ;
  assign n5044 = n5035 | n5043 ;
  assign n5045 = ( n4980 & n5008 ) | ( n4980 & n5044 ) | ( n5008 & n5044 ) ;
  assign n5046 = ~n4926 & n4965 ;
  assign n5047 = n5045 & n5046 ;
  assign n5048 = ( n4967 & n5045 ) | ( n4967 & n5047 ) | ( n5045 & n5047 ) ;
  assign n5049 = n4966 | n5048 ;
  assign n5050 = n4825 | n4853 ;
  assign n5051 = n3285 & ~n5050 ;
  assign n5052 = n3222 & n5051 ;
  assign n5053 = n174 | n361 ;
  assign n5054 = n419 | n4952 ;
  assign n5055 = n159 | n232 ;
  assign n5056 = n198 | n5055 ;
  assign n5057 = n5054 | n5056 ;
  assign n5058 = n212 | n538 ;
  assign n5059 = n407 | n5058 ;
  assign n5060 = n5057 | n5059 ;
  assign n5061 = n3181 | n3182 ;
  assign n5062 = n224 | n528 ;
  assign n5063 = n444 | n5062 ;
  assign n5064 = n964 | n5063 ;
  assign n5065 = n5061 | n5064 ;
  assign n5066 = n5060 | n5065 ;
  assign n5067 = n254 | n278 ;
  assign n5068 = n2733 | n5067 ;
  assign n5069 = n144 | n165 ;
  assign n5070 = n426 | n5069 ;
  assign n5071 = n5068 | n5070 ;
  assign n5072 = n141 | n5071 ;
  assign n5073 = n5066 | n5072 ;
  assign n5074 = n957 & ~n5073 ;
  assign n5075 = ~n5053 & n5074 ;
  assign n5076 = n5051 & ~n5075 ;
  assign n5077 = n3222 & n5076 ;
  assign n5078 = n5051 | n5075 ;
  assign n5079 = ( n3222 & n5075 ) | ( n3222 & n5078 ) | ( n5075 & n5078 ) ;
  assign n5080 = ( ~n5052 & n5077 ) | ( ~n5052 & n5079 ) | ( n5077 & n5079 ) ;
  assign n5081 = n4854 & n5080 ;
  assign n5082 = ~n3286 & n5080 ;
  assign n5083 = ( ~n4855 & n5081 ) | ( ~n4855 & n5082 ) | ( n5081 & n5082 ) ;
  assign n5084 = n4854 | n5080 ;
  assign n5085 = n3286 & ~n5080 ;
  assign n5086 = ( n4855 & ~n5084 ) | ( n4855 & n5085 ) | ( ~n5084 & n5085 ) ;
  assign n5087 = n5083 | n5086 ;
  assign n5088 = n4831 | n4861 ;
  assign n5089 = ( n4861 & n4862 ) | ( n4861 & n5088 ) | ( n4862 & n5088 ) ;
  assign n5090 = ~n5087 & n5089 ;
  assign n5091 = ~n4834 & n4862 ;
  assign n5092 = n4861 & ~n5087 ;
  assign n5093 = ( ~n5087 & n5091 ) | ( ~n5087 & n5092 ) | ( n5091 & n5092 ) ;
  assign n5094 = ( n4841 & n5090 ) | ( n4841 & n5093 ) | ( n5090 & n5093 ) ;
  assign n5095 = n5087 & ~n5089 ;
  assign n5096 = ~n4861 & n5087 ;
  assign n5097 = ~n5091 & n5096 ;
  assign n5098 = ( ~n4841 & n5095 ) | ( ~n4841 & n5097 ) | ( n5095 & n5097 ) ;
  assign n5099 = n5094 | n5098 ;
  assign n5100 = n3335 & ~n4854 ;
  assign n5101 = n3285 & n3335 ;
  assign n5102 = n3222 & n5101 ;
  assign n5103 = ( n4855 & n5100 ) | ( n4855 & n5102 ) | ( n5100 & n5102 ) ;
  assign n5104 = n3338 & ~n5080 ;
  assign n5105 = n3333 & n4830 ;
  assign n5106 = n5104 | n5105 ;
  assign n5107 = n5103 | n5106 ;
  assign n5108 = n3340 | n5107 ;
  assign n5109 = ( ~n5099 & n5107 ) | ( ~n5099 & n5108 ) | ( n5107 & n5108 ) ;
  assign n5110 = n3326 & n5107 ;
  assign n5111 = ( n3326 & n4281 ) | ( n3326 & n5107 ) | ( n4281 & n5107 ) ;
  assign n5112 = ( ~n5099 & n5110 ) | ( ~n5099 & n5111 ) | ( n5110 & n5111 ) ;
  assign n5113 = n5109 & ~n5112 ;
  assign n5114 = n3326 & ~n5107 ;
  assign n5115 = n4233 & ~n5107 ;
  assign n5116 = ( n5099 & n5114 ) | ( n5099 & n5115 ) | ( n5114 & n5115 ) ;
  assign n5117 = n5113 | n5116 ;
  assign n5118 = n3266 & n3373 ;
  assign n5119 = n3259 & n3367 ;
  assign n5120 = n5118 | n5119 ;
  assign n5121 = ~n3289 & n3380 ;
  assign n5122 = ( ~n3289 & n3387 ) | ( ~n3289 & n3905 ) | ( n3387 & n3905 ) ;
  assign n5123 = n5121 & n5122 ;
  assign n5124 = n5120 | n5123 ;
  assign n5125 = n1115 | n5124 ;
  assign n5126 = ( ~n3289 & n3394 ) | ( ~n3289 & n3910 ) | ( n3394 & n3910 ) ;
  assign n5127 = n5120 | n5126 ;
  assign n5128 = ( ~n3321 & n5125 ) | ( ~n3321 & n5127 ) | ( n5125 & n5127 ) ;
  assign n5129 = n1115 & n5124 ;
  assign n5130 = ( ~n3289 & n3388 ) | ( ~n3289 & n3915 ) | ( n3388 & n3915 ) ;
  assign n5131 = ( n1115 & n5120 ) | ( n1115 & n5130 ) | ( n5120 & n5130 ) ;
  assign n5132 = ( ~n3321 & n5129 ) | ( ~n3321 & n5131 ) | ( n5129 & n5131 ) ;
  assign n5133 = n5128 & ~n5132 ;
  assign n5134 = n3024 & n3637 ;
  assign n5135 = n2916 & n3635 ;
  assign n5136 = ( ~n2901 & n3635 ) | ( ~n2901 & n5135 ) | ( n3635 & n5135 ) ;
  assign n5137 = ~n2921 & n5136 ;
  assign n5138 = n2828 & n5137 ;
  assign n5139 = ( n2927 & n3635 ) | ( n2927 & n5138 ) | ( n3635 & n5138 ) ;
  assign n5140 = n5134 | n5139 ;
  assign n5141 = n3296 & n3641 ;
  assign n5142 = n3295 & n3641 ;
  assign n5143 = ( n2828 & n5141 ) | ( n2828 & n5142 ) | ( n5141 & n5142 ) ;
  assign n5144 = ( ~n3300 & n3641 ) | ( ~n3300 & n5143 ) | ( n3641 & n5143 ) ;
  assign n5145 = n5140 | n5144 ;
  assign n5146 = n3643 | n5144 ;
  assign n5147 = n5140 | n5146 ;
  assign n5148 = ( ~n3360 & n5145 ) | ( ~n3360 & n5147 ) | ( n5145 & n5147 ) ;
  assign n5149 = ( n482 & n3656 ) | ( n482 & n5144 ) | ( n3656 & n5144 ) ;
  assign n5150 = ( n482 & n5140 ) | ( n482 & n5149 ) | ( n5140 & n5149 ) ;
  assign n5151 = n482 & n5144 ;
  assign n5152 = ( n482 & n5140 ) | ( n482 & n5151 ) | ( n5140 & n5151 ) ;
  assign n5153 = ( ~n3360 & n5150 ) | ( ~n3360 & n5152 ) | ( n5150 & n5152 ) ;
  assign n5154 = n5148 & ~n5153 ;
  assign n5155 = n482 & ~n5151 ;
  assign n5156 = ~n5140 & n5155 ;
  assign n5157 = n482 & ~n5146 ;
  assign n5158 = ~n5140 & n5157 ;
  assign n5159 = ( n3360 & n5156 ) | ( n3360 & n5158 ) | ( n5156 & n5158 ) ;
  assign n5160 = n5154 | n5159 ;
  assign n5184 = n4661 | n4662 ;
  assign n5185 = n4653 | n4661 ;
  assign n5186 = ( ~n4663 & n5184 ) | ( ~n4663 & n5185 ) | ( n5184 & n5185 ) ;
  assign n5187 = ( n4625 & n4661 ) | ( n4625 & n5186 ) | ( n4661 & n5186 ) ;
  assign n5171 = n879 & n2823 ;
  assign n5172 = ( n879 & n2764 ) | ( n879 & n5171 ) | ( n2764 & n5171 ) ;
  assign n5173 = ~n3071 & n5172 ;
  assign n5161 = n3070 & n3477 ;
  assign n5162 = n3063 & n3446 ;
  assign n5163 = n5161 | n5162 ;
  assign n5164 = n2368 & n3448 ;
  assign n5165 = ( ~n2340 & n3448 ) | ( ~n2340 & n5164 ) | ( n3448 & n5164 ) ;
  assign n5166 = ~n2679 & n5165 ;
  assign n5167 = n2827 & n5166 ;
  assign n5168 = ( n3057 & n3448 ) | ( n3057 & n5167 ) | ( n3448 & n5167 ) ;
  assign n5169 = n5163 | n5168 ;
  assign n5170 = ( n3401 & n3452 ) | ( n3401 & n5169 ) | ( n3452 & n5169 ) ;
  assign n5174 = ( n3452 & ~n5168 ) | ( n3452 & n5173 ) | ( ~n5168 & n5173 ) ;
  assign n5175 = n3452 & n5173 ;
  assign n5176 = ( ~n5163 & n5174 ) | ( ~n5163 & n5175 ) | ( n5174 & n5175 ) ;
  assign n5177 = ( n3401 & n5173 ) | ( n3401 & n5176 ) | ( n5173 & n5176 ) ;
  assign n5178 = ~n5170 & n5177 ;
  assign n5179 = n5169 | n5176 ;
  assign n5180 = n5168 | n5173 ;
  assign n5181 = n5163 | n5180 ;
  assign n5182 = ( n3401 & n5179 ) | ( n3401 & n5181 ) | ( n5179 & n5181 ) ;
  assign n5183 = ( ~n5173 & n5178 ) | ( ~n5173 & n5182 ) | ( n5178 & n5182 ) ;
  assign n5188 = n5183 | n5187 ;
  assign n5189 = ~n5183 & n5187 ;
  assign n5190 = ( ~n5187 & n5188 ) | ( ~n5187 & n5189 ) | ( n5188 & n5189 ) ;
  assign n5191 = n3049 & n3412 ;
  assign n5192 = n3110 & n3414 ;
  assign n5193 = ( ~n3106 & n3414 ) | ( ~n3106 & n5192 ) | ( n3414 & n5192 ) ;
  assign n5194 = n5191 | n5193 ;
  assign n5195 = n3033 & n3417 ;
  assign n5196 = ( n3033 & n3423 ) | ( n3033 & n4683 ) | ( n3423 & n4683 ) ;
  assign n5197 = n5195 & n5196 ;
  assign n5198 = n5194 | n5197 ;
  assign n5199 = n634 | n5198 ;
  assign n5200 = n634 | n4683 ;
  assign n5201 = ( n3033 & n3431 ) | ( n3033 & n5200 ) | ( n3431 & n5200 ) ;
  assign n5202 = n5194 | n5201 ;
  assign n5203 = ( ~n3624 & n5199 ) | ( ~n3624 & n5202 ) | ( n5199 & n5202 ) ;
  assign n5204 = n634 & n5198 ;
  assign n5205 = n634 & n4683 ;
  assign n5206 = ( n3033 & n3424 ) | ( n3033 & n5205 ) | ( n3424 & n5205 ) ;
  assign n5207 = ( n634 & n5194 ) | ( n634 & n5206 ) | ( n5194 & n5206 ) ;
  assign n5208 = ( ~n3624 & n5204 ) | ( ~n3624 & n5207 ) | ( n5204 & n5207 ) ;
  assign n5209 = n5203 & ~n5208 ;
  assign n5210 = n5190 & n5209 ;
  assign n5211 = n5190 & ~n5210 ;
  assign n5212 = ~n5190 & n5209 ;
  assign n5213 = n5211 | n5212 ;
  assign n5214 = n4670 | n4697 ;
  assign n5215 = n4703 | n5214 ;
  assign n5216 = ( n4670 & n4672 ) | ( n4670 & n5215 ) | ( n4672 & n5215 ) ;
  assign n5217 = ( n5160 & n5213 ) | ( n5160 & ~n5216 ) | ( n5213 & ~n5216 ) ;
  assign n5218 = ( ~n5213 & n5216 ) | ( ~n5213 & n5217 ) | ( n5216 & n5217 ) ;
  assign n5219 = ( ~n5160 & n5217 ) | ( ~n5160 & n5218 ) | ( n5217 & n5218 ) ;
  assign n5220 = n4728 | n5219 ;
  assign n5221 = n4760 | n5220 ;
  assign n5222 = n4728 & n5219 ;
  assign n5223 = ( n4760 & n5219 ) | ( n4760 & n5222 ) | ( n5219 & n5222 ) ;
  assign n5224 = n5221 & ~n5223 ;
  assign n5225 = n5133 & n5224 ;
  assign n5226 = n5224 & ~n5225 ;
  assign n5227 = ( n5133 & ~n5225 ) | ( n5133 & n5226 ) | ( ~n5225 & n5226 ) ;
  assign n5228 = n4763 | n4765 ;
  assign n5229 = ( n4763 & n4806 ) | ( n4763 & n5228 ) | ( n4806 & n5228 ) ;
  assign n5230 = n5227 & n5229 ;
  assign n5231 = n5227 & ~n5230 ;
  assign n5232 = ~n5227 & n5229 ;
  assign n5233 = n5117 & n5232 ;
  assign n5234 = ( n5117 & n5231 ) | ( n5117 & n5233 ) | ( n5231 & n5233 ) ;
  assign n5235 = n5117 | n5232 ;
  assign n5236 = n5231 | n5235 ;
  assign n5237 = ~n5234 & n5236 ;
  assign n5238 = n4893 | n5237 ;
  assign n5239 = n4925 | n5238 ;
  assign n5240 = n4893 & n5237 ;
  assign n5241 = ( n4925 & n5237 ) | ( n4925 & n5240 ) | ( n5237 & n5240 ) ;
  assign n5242 = n5239 & ~n5241 ;
  assign n5243 = n303 | n305 ;
  assign n5244 = n298 | n5243 ;
  assign n5245 = n288 | n5244 ;
  assign n5246 = n4944 | n5245 ;
  assign n5247 = n182 | n700 ;
  assign n5248 = n369 | n4952 ;
  assign n5249 = n817 | n5248 ;
  assign n5250 = n200 | n360 ;
  assign n5251 = n830 | n5250 ;
  assign n5252 = n5249 | n5251 ;
  assign n5253 = n5247 | n5252 ;
  assign n5254 = n2307 | n5253 ;
  assign n5255 = n5246 | n5254 ;
  assign n5256 = n167 | n570 ;
  assign n5257 = n270 | n5256 ;
  assign n5258 = n5255 | n5257 ;
  assign n5259 = n5242 | n5258 ;
  assign n5260 = n5242 & n5258 ;
  assign n5261 = n5259 & ~n5260 ;
  assign n5262 = n5049 & n5261 ;
  assign n5263 = n5049 | n5261 ;
  assign n5264 = ~n5262 & n5263 ;
  assign n5265 = n5045 | n5046 ;
  assign n5266 = n4967 | n5265 ;
  assign n5267 = ~n5048 & n5266 ;
  assign n5268 = n5264 & n5267 ;
  assign n5269 = n5264 & ~n5268 ;
  assign n5270 = ~n5264 & n5267 ;
  assign n5271 = n5269 | n5270 ;
  assign n5272 = n5234 | n5241 ;
  assign n5273 = n3335 & ~n5080 ;
  assign n5274 = n3333 & ~n4854 ;
  assign n5275 = n3285 & n3333 ;
  assign n5276 = n3222 & n5275 ;
  assign n5277 = ( n4855 & n5274 ) | ( n4855 & n5276 ) | ( n5274 & n5276 ) ;
  assign n5278 = n5273 | n5277 ;
  assign n5279 = n843 & ~n845 ;
  assign n5280 = n245 | n323 ;
  assign n5281 = n427 | n542 ;
  assign n5282 = n5280 | n5281 ;
  assign n5283 = n319 | n5282 ;
  assign n5284 = n5279 & ~n5283 ;
  assign n5285 = n2549 | n2723 ;
  assign n5286 = n175 | n5285 ;
  assign n5287 = n721 | n5286 ;
  assign n5288 = n333 | n358 ;
  assign n5289 = n206 | n261 ;
  assign n5290 = n5288 | n5289 ;
  assign n5291 = n5287 | n5290 ;
  assign n5292 = n5284 & ~n5291 ;
  assign n5293 = ~n582 & n5292 ;
  assign n5294 = n217 | n262 ;
  assign n5295 = n305 | n425 ;
  assign n5296 = n5294 | n5295 ;
  assign n5297 = n361 | n5296 ;
  assign n5298 = n2746 | n5297 ;
  assign n5299 = n5293 & ~n5298 ;
  assign n5301 = ~n5051 & n5075 ;
  assign n5302 = n3222 & n5301 ;
  assign n5300 = n3222 & n5075 ;
  assign n5303 = ( n5299 & n5300 ) | ( n5299 & n5302 ) | ( n5300 & n5302 ) ;
  assign n5304 = ( n5299 & n5302 ) | ( n5299 & ~n5303 ) | ( n5302 & ~n5303 ) ;
  assign n5305 = n3338 & n5303 ;
  assign n5306 = n3338 & ~n5075 ;
  assign n5307 = ( ~n3222 & n3338 ) | ( ~n3222 & n5306 ) | ( n3338 & n5306 ) ;
  assign n5308 = ( ~n5304 & n5305 ) | ( ~n5304 & n5307 ) | ( n5305 & n5307 ) ;
  assign n5309 = n5278 | n5308 ;
  assign n5310 = n5080 & ~n5303 ;
  assign n5311 = n5080 & n5300 ;
  assign n5312 = ( n5304 & n5310 ) | ( n5304 & n5311 ) | ( n5310 & n5311 ) ;
  assign n5313 = ~n5080 & n5303 ;
  assign n5314 = n5080 | n5300 ;
  assign n5315 = ( n5304 & ~n5313 ) | ( n5304 & n5314 ) | ( ~n5313 & n5314 ) ;
  assign n5316 = ~n5312 & n5315 ;
  assign n5317 = n5086 & n5316 ;
  assign n5318 = ( n5093 & n5316 ) | ( n5093 & n5317 ) | ( n5316 & n5317 ) ;
  assign n5319 = ( n5090 & n5316 ) | ( n5090 & n5317 ) | ( n5316 & n5317 ) ;
  assign n5320 = ( n4841 & n5318 ) | ( n4841 & n5319 ) | ( n5318 & n5319 ) ;
  assign n5321 = n5086 | n5316 ;
  assign n5322 = n5093 | n5321 ;
  assign n5323 = n5090 | n5321 ;
  assign n5324 = ( n4841 & n5322 ) | ( n4841 & n5323 ) | ( n5322 & n5323 ) ;
  assign n5325 = ~n5320 & n5324 ;
  assign n5326 = n3340 | n5308 ;
  assign n5327 = n5278 | n5326 ;
  assign n5328 = ( n5309 & n5325 ) | ( n5309 & n5327 ) | ( n5325 & n5327 ) ;
  assign n5329 = n3326 & n5327 ;
  assign n5330 = n3326 & n5308 ;
  assign n5331 = ( n3326 & n5278 ) | ( n3326 & n5330 ) | ( n5278 & n5330 ) ;
  assign n5332 = ( n5325 & n5329 ) | ( n5325 & n5331 ) | ( n5329 & n5331 ) ;
  assign n5333 = n5328 & ~n5332 ;
  assign n5334 = n3326 & ~n5331 ;
  assign n5335 = n3326 & ~n5327 ;
  assign n5336 = ( ~n5325 & n5334 ) | ( ~n5325 & n5335 ) | ( n5334 & n5335 ) ;
  assign n5337 = n5333 | n5336 ;
  assign n5338 = n5225 | n5229 ;
  assign n5339 = ( n5225 & n5227 ) | ( n5225 & n5338 ) | ( n5227 & n5338 ) ;
  assign n5340 = n3259 & n3373 ;
  assign n5341 = ~n3289 & n3367 ;
  assign n5342 = n5340 | n5341 ;
  assign n5343 = n3380 & n4830 ;
  assign n5344 = ( n3387 & n3905 ) | ( n3387 & n4830 ) | ( n3905 & n4830 ) ;
  assign n5345 = n5343 & n5344 ;
  assign n5346 = n5342 | n5345 ;
  assign n5347 = n1115 | n5346 ;
  assign n5348 = ( n3394 & n3910 ) | ( n3394 & n4830 ) | ( n3910 & n4830 ) ;
  assign n5349 = n5342 | n5348 ;
  assign n5350 = ( ~n4901 & n5347 ) | ( ~n4901 & n5349 ) | ( n5347 & n5349 ) ;
  assign n5351 = n1115 & n5346 ;
  assign n5352 = ( n3388 & n3915 ) | ( n3388 & n4830 ) | ( n3915 & n4830 ) ;
  assign n5353 = ( n1115 & n5342 ) | ( n1115 & n5352 ) | ( n5342 & n5352 ) ;
  assign n5354 = ( ~n4901 & n5351 ) | ( ~n4901 & n5353 ) | ( n5351 & n5353 ) ;
  assign n5355 = n5350 & ~n5354 ;
  assign n5356 = ( n5190 & n5209 ) | ( n5190 & n5216 ) | ( n5209 & n5216 ) ;
  assign n5357 = n879 & ~n3070 ;
  assign n5358 = n3063 & n3477 ;
  assign n5359 = n2368 & n3446 ;
  assign n5360 = ( ~n2340 & n3446 ) | ( ~n2340 & n5359 ) | ( n3446 & n5359 ) ;
  assign n5361 = ~n2679 & n5360 ;
  assign n5362 = n2827 & n5361 ;
  assign n5363 = ( n3057 & n3446 ) | ( n3057 & n5362 ) | ( n3446 & n5362 ) ;
  assign n5364 = n5358 | n5363 ;
  assign n5365 = n3448 | n3452 ;
  assign n5366 = ( n3049 & n3452 ) | ( n3049 & n5365 ) | ( n3452 & n5365 ) ;
  assign n5367 = n5364 | n5366 ;
  assign n5368 = n5357 & n5367 ;
  assign n5369 = n879 & n3448 ;
  assign n5370 = ~n3070 & n5369 ;
  assign n5371 = n3049 & n5370 ;
  assign n5372 = ( n5357 & n5364 ) | ( n5357 & n5371 ) | ( n5364 & n5371 ) ;
  assign n5373 = ( n3856 & n5368 ) | ( n3856 & n5372 ) | ( n5368 & n5372 ) ;
  assign n5374 = n5357 | n5367 ;
  assign n5375 = n879 | n3448 ;
  assign n5376 = ( ~n3070 & n3448 ) | ( ~n3070 & n5375 ) | ( n3448 & n5375 ) ;
  assign n5377 = ( n3049 & n5357 ) | ( n3049 & n5376 ) | ( n5357 & n5376 ) ;
  assign n5378 = n5364 | n5377 ;
  assign n5379 = ( n3856 & n5374 ) | ( n3856 & n5378 ) | ( n5374 & n5378 ) ;
  assign n5380 = ~n5373 & n5379 ;
  assign n5381 = n879 & ~n2823 ;
  assign n5382 = ~n2764 & n5381 ;
  assign n5383 = ( n879 & n3071 ) | ( n879 & n5382 ) | ( n3071 & n5382 ) ;
  assign n5384 = ~n5168 & n5383 ;
  assign n5385 = ~n5163 & n5384 ;
  assign n5386 = ~n3452 & n5385 ;
  assign n5387 = ( ~n3401 & n5385 ) | ( ~n3401 & n5386 ) | ( n5385 & n5386 ) ;
  assign n5388 = n4661 & n5179 ;
  assign n5389 = n4661 & n5181 ;
  assign n5390 = ( n3401 & n5388 ) | ( n3401 & n5389 ) | ( n5388 & n5389 ) ;
  assign n5391 = n5387 | n5390 ;
  assign n5392 = n4661 & ~n5173 ;
  assign n5393 = n5387 | n5392 ;
  assign n5394 = ( n5178 & n5391 ) | ( n5178 & n5393 ) | ( n5391 & n5393 ) ;
  assign n5395 = n5380 & n5394 ;
  assign n5396 = n5182 | n5387 ;
  assign n5397 = n5173 & ~n5386 ;
  assign n5398 = n5173 & ~n5385 ;
  assign n5399 = ( n3401 & n5397 ) | ( n3401 & n5398 ) | ( n5397 & n5398 ) ;
  assign n5400 = ( n5178 & n5396 ) | ( n5178 & ~n5399 ) | ( n5396 & ~n5399 ) ;
  assign n5401 = n5380 & n5400 ;
  assign n5402 = ( n4665 & n5395 ) | ( n4665 & n5401 ) | ( n5395 & n5401 ) ;
  assign n5403 = n5380 | n5394 ;
  assign n5404 = n5380 | n5400 ;
  assign n5405 = ( n4665 & n5403 ) | ( n4665 & n5404 ) | ( n5403 & n5404 ) ;
  assign n5406 = ~n5402 & n5405 ;
  assign n5407 = n3033 & n3414 ;
  assign n5408 = n3110 & n3412 ;
  assign n5409 = ( ~n3106 & n3412 ) | ( ~n3106 & n5408 ) | ( n3412 & n5408 ) ;
  assign n5410 = n5407 | n5409 ;
  assign n5411 = n2916 & n3417 ;
  assign n5412 = ( ~n2901 & n3417 ) | ( ~n2901 & n5411 ) | ( n3417 & n5411 ) ;
  assign n5413 = ~n2921 & n5412 ;
  assign n5414 = n2828 & n5413 ;
  assign n5415 = ( n2927 & n3417 ) | ( n2927 & n5414 ) | ( n3417 & n5414 ) ;
  assign n5416 = n5410 | n5415 ;
  assign n5417 = ( n3423 & n3952 ) | ( n3423 & n5416 ) | ( n3952 & n5416 ) ;
  assign n5418 = ( n634 & n3423 ) | ( n634 & ~n5416 ) | ( n3423 & ~n5416 ) ;
  assign n5419 = ( n634 & n3952 ) | ( n634 & n5418 ) | ( n3952 & n5418 ) ;
  assign n5420 = ~n5417 & n5419 ;
  assign n5421 = n5416 | n5418 ;
  assign n5422 = n634 | n5416 ;
  assign n5423 = ( n3952 & n5421 ) | ( n3952 & n5422 ) | ( n5421 & n5422 ) ;
  assign n5424 = ( ~n634 & n5420 ) | ( ~n634 & n5423 ) | ( n5420 & n5423 ) ;
  assign n5425 = n5406 & n5424 ;
  assign n5426 = n5406 & ~n5425 ;
  assign n5427 = ~n5406 & n5424 ;
  assign n5428 = n5426 | n5427 ;
  assign n5429 = n5356 & n5428 ;
  assign n5430 = n5356 & ~n5429 ;
  assign n5431 = n3266 & n3641 ;
  assign n5432 = n3024 & n3635 ;
  assign n5433 = n3296 & n3637 ;
  assign n5434 = n3295 & n3637 ;
  assign n5435 = ( n2828 & n5433 ) | ( n2828 & n5434 ) | ( n5433 & n5434 ) ;
  assign n5436 = ( ~n3300 & n3637 ) | ( ~n3300 & n5435 ) | ( n3637 & n5435 ) ;
  assign n5437 = n5432 | n5436 ;
  assign n5438 = n5431 | n5437 ;
  assign n5439 = ( n3266 & n3643 ) | ( n3266 & n3644 ) | ( n3643 & n3644 ) ;
  assign n5440 = n5437 | n5439 ;
  assign n5441 = ( ~n4190 & n5438 ) | ( ~n4190 & n5440 ) | ( n5438 & n5440 ) ;
  assign n5442 = n482 & n3641 ;
  assign n5443 = n3266 & n5442 ;
  assign n5444 = ( n482 & n5437 ) | ( n482 & n5443 ) | ( n5437 & n5443 ) ;
  assign n5445 = n482 & n5439 ;
  assign n5446 = ( n482 & n5437 ) | ( n482 & n5445 ) | ( n5437 & n5445 ) ;
  assign n5447 = ( ~n4190 & n5444 ) | ( ~n4190 & n5446 ) | ( n5444 & n5446 ) ;
  assign n5448 = n5441 & ~n5447 ;
  assign n5449 = n482 & ~n5443 ;
  assign n5450 = ~n5437 & n5449 ;
  assign n5451 = n482 & ~n5439 ;
  assign n5452 = ~n5437 & n5451 ;
  assign n5453 = ( n4190 & n5450 ) | ( n4190 & n5452 ) | ( n5450 & n5452 ) ;
  assign n5454 = n5448 | n5453 ;
  assign n5455 = n5427 & n5454 ;
  assign n5456 = ( n5426 & n5454 ) | ( n5426 & n5455 ) | ( n5454 & n5455 ) ;
  assign n5457 = n5454 & ~n5456 ;
  assign n5458 = ( n5356 & n5454 ) | ( n5356 & n5457 ) | ( n5454 & n5457 ) ;
  assign n5459 = ~n5430 & n5458 ;
  assign n5460 = ~n5356 & n5456 ;
  assign n5461 = ( n5356 & n5428 ) | ( n5356 & ~n5460 ) | ( n5428 & ~n5460 ) ;
  assign n5462 = ( n5356 & n5428 ) | ( n5356 & ~n5454 ) | ( n5428 & ~n5454 ) ;
  assign n5463 = ( ~n5430 & n5461 ) | ( ~n5430 & n5462 ) | ( n5461 & n5462 ) ;
  assign n5464 = ~n5429 & n5463 ;
  assign n5465 = n5459 | n5464 ;
  assign n5466 = n5213 & n5216 ;
  assign n5467 = n5216 & ~n5466 ;
  assign n5468 = n5160 & n5212 ;
  assign n5469 = ( n5160 & n5211 ) | ( n5160 & n5468 ) | ( n5211 & n5468 ) ;
  assign n5470 = ~n5216 & n5469 ;
  assign n5471 = ( n5160 & n5467 ) | ( n5160 & n5470 ) | ( n5467 & n5470 ) ;
  assign n5472 = n5223 | n5471 ;
  assign n5473 = n5465 | n5472 ;
  assign n5474 = n5465 & n5472 ;
  assign n5475 = n5473 & ~n5474 ;
  assign n5476 = n5355 & n5475 ;
  assign n5477 = n5475 & ~n5476 ;
  assign n5478 = ( n5355 & ~n5476 ) | ( n5355 & n5477 ) | ( ~n5476 & n5477 ) ;
  assign n5479 = n5339 & ~n5478 ;
  assign n5480 = ~n5339 & n5478 ;
  assign n5481 = n5479 | n5480 ;
  assign n5482 = n5337 & n5481 ;
  assign n5483 = n5337 | n5481 ;
  assign n5484 = ~n5482 & n5483 ;
  assign n5485 = n5272 | n5484 ;
  assign n5486 = n5272 & n5484 ;
  assign n5487 = n5485 & ~n5486 ;
  assign n5488 = n4941 | n4955 ;
  assign n5489 = n425 | n2610 ;
  assign n5490 = n696 | n2349 ;
  assign n5491 = n701 | n5490 ;
  assign n5492 = n5489 | n5491 ;
  assign n5493 = n2604 | n5492 ;
  assign n5494 = n5488 | n5493 ;
  assign n5495 = n183 | n397 ;
  assign n5496 = n866 | n5495 ;
  assign n5497 = n175 | n5496 ;
  assign n5498 = n3241 | n4944 ;
  assign n5499 = n5497 | n5498 ;
  assign n5500 = n292 | n366 ;
  assign n5501 = n228 | n524 ;
  assign n5502 = n212 | n333 ;
  assign n5503 = n5501 | n5502 ;
  assign n5504 = n5500 | n5503 ;
  assign n5505 = n5499 | n5504 ;
  assign n5506 = n5494 | n5505 ;
  assign n5507 = n5487 | n5506 ;
  assign n5508 = n5487 & n5506 ;
  assign n5509 = n5507 & ~n5508 ;
  assign n5510 = n5260 | n5261 ;
  assign n5511 = ( n5049 & n5260 ) | ( n5049 & n5510 ) | ( n5260 & n5510 ) ;
  assign n5512 = n5509 & n5511 ;
  assign n5513 = n5509 | n5511 ;
  assign n5514 = ~n5512 & n5513 ;
  assign n5515 = n5268 & n5514 ;
  assign n5516 = n5268 | n5514 ;
  assign n5517 = ~n5515 & n5516 ;
  assign n5518 = x22 & ~x23 ;
  assign n5519 = ~x22 & x23 ;
  assign n5520 = n5518 | n5519 ;
  assign n5521 = n5271 & n5520 ;
  assign n5522 = ~n5517 & n5521 ;
  assign n5523 = n5517 & ~n5521 ;
  assign n5524 = n5522 | n5523 ;
  assign n5525 = n5508 | n5512 ;
  assign n5526 = n3333 & ~n5080 ;
  assign n5527 = n3335 & n5303 ;
  assign n5528 = n3335 & ~n5075 ;
  assign n5529 = ( ~n3222 & n3335 ) | ( ~n3222 & n5528 ) | ( n3335 & n5528 ) ;
  assign n5530 = ( ~n5304 & n5527 ) | ( ~n5304 & n5529 ) | ( n5527 & n5529 ) ;
  assign n5531 = n5526 | n5530 ;
  assign n5532 = ( n5300 & ~n5303 ) | ( n5300 & n5304 ) | ( ~n5303 & n5304 ) ;
  assign n5533 = n5080 & ~n5086 ;
  assign n5534 = ( n5080 & ~n5316 ) | ( n5080 & n5533 ) | ( ~n5316 & n5533 ) ;
  assign n5535 = n5532 | n5534 ;
  assign n5536 = ( n5315 & ~n5316 ) | ( n5315 & n5532 ) | ( ~n5316 & n5532 ) ;
  assign n5537 = ( ~n5093 & n5535 ) | ( ~n5093 & n5536 ) | ( n5535 & n5536 ) ;
  assign n5538 = ( ~n5090 & n5535 ) | ( ~n5090 & n5536 ) | ( n5535 & n5536 ) ;
  assign n5539 = ( ~n4841 & n5537 ) | ( ~n4841 & n5538 ) | ( n5537 & n5538 ) ;
  assign n5540 = ~n5316 & n5532 ;
  assign n5541 = ~n5086 & n5532 ;
  assign n5542 = ( ~n5316 & n5532 ) | ( ~n5316 & n5541 ) | ( n5532 & n5541 ) ;
  assign n5543 = ( ~n5093 & n5540 ) | ( ~n5093 & n5542 ) | ( n5540 & n5542 ) ;
  assign n5544 = ( ~n5090 & n5540 ) | ( ~n5090 & n5542 ) | ( n5540 & n5542 ) ;
  assign n5545 = ( ~n4841 & n5543 ) | ( ~n4841 & n5544 ) | ( n5543 & n5544 ) ;
  assign n5546 = n5539 & ~n5545 ;
  assign n5547 = n3333 | n3340 ;
  assign n5548 = ( n3340 & ~n5080 ) | ( n3340 & n5547 ) | ( ~n5080 & n5547 ) ;
  assign n5549 = n5530 | n5548 ;
  assign n5550 = ( n5531 & n5546 ) | ( n5531 & n5549 ) | ( n5546 & n5549 ) ;
  assign n5551 = ( n3326 & n4281 ) | ( n3326 & n5526 ) | ( n4281 & n5526 ) ;
  assign n5552 = ( n4282 & n5530 ) | ( n4282 & n5551 ) | ( n5530 & n5551 ) ;
  assign n5553 = n3326 & n5526 ;
  assign n5554 = ( n3326 & n5530 ) | ( n3326 & n5553 ) | ( n5530 & n5553 ) ;
  assign n5555 = ( n5546 & n5552 ) | ( n5546 & n5554 ) | ( n5552 & n5554 ) ;
  assign n5556 = n5550 & ~n5555 ;
  assign n5557 = n4290 & ~n5526 ;
  assign n5558 = ~n5530 & n5557 ;
  assign n5559 = n3326 & ~n5526 ;
  assign n5560 = ~n5530 & n5559 ;
  assign n5561 = ( ~n5546 & n5558 ) | ( ~n5546 & n5560 ) | ( n5558 & n5560 ) ;
  assign n5562 = n5556 | n5561 ;
  assign n5563 = n5227 | n5476 ;
  assign n5564 = n5225 | n5355 ;
  assign n5565 = ( n5225 & n5475 ) | ( n5225 & n5564 ) | ( n5475 & n5564 ) ;
  assign n5566 = ( n5338 & n5563 ) | ( n5338 & n5565 ) | ( n5563 & n5565 ) ;
  assign n5567 = ( n5476 & n5478 ) | ( n5476 & n5566 ) | ( n5478 & n5566 ) ;
  assign n5568 = ~n3289 & n3373 ;
  assign n5569 = n3367 & n4830 ;
  assign n5570 = n5568 | n5569 ;
  assign n5571 = ( n3387 & n3905 ) | ( n3387 & ~n4854 ) | ( n3905 & ~n4854 ) ;
  assign n5572 = ( n3285 & n3387 ) | ( n3285 & n3905 ) | ( n3387 & n3905 ) ;
  assign n5573 = n3387 & n3905 ;
  assign n5574 = ( n3222 & n5572 ) | ( n3222 & n5573 ) | ( n5572 & n5573 ) ;
  assign n5575 = ( n4855 & n5571 ) | ( n4855 & n5574 ) | ( n5571 & n5574 ) ;
  assign n5576 = n5570 | n5575 ;
  assign n5577 = n1115 | n5576 ;
  assign n5578 = n3380 & ~n4854 ;
  assign n5579 = n3285 & n3380 ;
  assign n5580 = n3222 & n5579 ;
  assign n5581 = ( n4855 & n5578 ) | ( n4855 & n5580 ) | ( n5578 & n5580 ) ;
  assign n5582 = n5575 & n5581 ;
  assign n5583 = n1115 | n5570 ;
  assign n5584 = n5582 | n5583 ;
  assign n5585 = ( n4869 & n5577 ) | ( n4869 & n5584 ) | ( n5577 & n5584 ) ;
  assign n5586 = n1115 & n5576 ;
  assign n5587 = n1115 & n5570 ;
  assign n5588 = ( n1115 & n5582 ) | ( n1115 & n5587 ) | ( n5582 & n5587 ) ;
  assign n5589 = ( n4869 & n5586 ) | ( n4869 & n5588 ) | ( n5586 & n5588 ) ;
  assign n5590 = n5585 & ~n5589 ;
  assign n5591 = ( n5430 & n5454 ) | ( n5430 & n5460 ) | ( n5454 & n5460 ) ;
  assign n5592 = n5459 | n5591 ;
  assign n5593 = n5464 | n5592 ;
  assign n5594 = ( n5472 & n5591 ) | ( n5472 & n5593 ) | ( n5591 & n5593 ) ;
  assign n5595 = n879 & ~n3063 ;
  assign n5596 = n2368 & n3477 ;
  assign n5597 = ( ~n2340 & n3477 ) | ( ~n2340 & n5596 ) | ( n3477 & n5596 ) ;
  assign n5598 = ~n2679 & n5597 ;
  assign n5599 = n2827 & n5598 ;
  assign n5600 = ( n3057 & n3477 ) | ( n3057 & n5599 ) | ( n3477 & n5599 ) ;
  assign n5601 = n3049 & n3446 ;
  assign n5602 = n5600 | n5601 ;
  assign n5603 = n3110 & n3448 ;
  assign n5604 = ( ~n3106 & n3448 ) | ( ~n3106 & n5603 ) | ( n3448 & n5603 ) ;
  assign n5605 = n3452 | n5604 ;
  assign n5606 = n5602 | n5605 ;
  assign n5607 = n5595 & n5606 ;
  assign n5608 = n5595 & n5604 ;
  assign n5609 = ( n5595 & n5602 ) | ( n5595 & n5608 ) | ( n5602 & n5608 ) ;
  assign n5610 = ( ~n3679 & n5607 ) | ( ~n3679 & n5609 ) | ( n5607 & n5609 ) ;
  assign n5611 = n5595 | n5606 ;
  assign n5612 = n5595 | n5604 ;
  assign n5613 = n5602 | n5612 ;
  assign n5614 = ( ~n3679 & n5611 ) | ( ~n3679 & n5613 ) | ( n5611 & n5613 ) ;
  assign n5615 = ~n5610 & n5614 ;
  assign n5616 = n3033 & n3412 ;
  assign n5617 = n2916 & n3414 ;
  assign n5618 = ( ~n2901 & n3414 ) | ( ~n2901 & n5617 ) | ( n3414 & n5617 ) ;
  assign n5619 = ~n2921 & n5618 ;
  assign n5620 = n2828 & n5619 ;
  assign n5621 = ( n2927 & n3414 ) | ( n2927 & n5620 ) | ( n3414 & n5620 ) ;
  assign n5622 = n5616 | n5621 ;
  assign n5623 = n3024 & n3417 ;
  assign n5624 = ( n3024 & n3423 ) | ( n3024 & n4683 ) | ( n3423 & n4683 ) ;
  assign n5625 = n5623 & n5624 ;
  assign n5626 = n5622 | n5625 ;
  assign n5627 = n634 | n5626 ;
  assign n5628 = ( n3024 & n3431 ) | ( n3024 & n5200 ) | ( n3431 & n5200 ) ;
  assign n5629 = n5622 | n5628 ;
  assign n5630 = ( n3896 & n5627 ) | ( n3896 & n5629 ) | ( n5627 & n5629 ) ;
  assign n5631 = n634 & n5626 ;
  assign n5632 = ( n3024 & n3424 ) | ( n3024 & n5205 ) | ( n3424 & n5205 ) ;
  assign n5633 = ( n634 & n5622 ) | ( n634 & n5632 ) | ( n5622 & n5632 ) ;
  assign n5634 = ( n3896 & n5631 ) | ( n3896 & n5633 ) | ( n5631 & n5633 ) ;
  assign n5635 = n5630 & ~n5634 ;
  assign n5636 = ( n4665 & n5394 ) | ( n4665 & n5400 ) | ( n5394 & n5400 ) ;
  assign n5637 = n879 & n3070 ;
  assign n5638 = ~n5367 & n5637 ;
  assign n5639 = n3049 & n3448 ;
  assign n5640 = ( n5364 & n5637 ) | ( n5364 & n5639 ) | ( n5637 & n5639 ) ;
  assign n5641 = n5637 & ~n5640 ;
  assign n5642 = ( ~n3856 & n5638 ) | ( ~n3856 & n5641 ) | ( n5638 & n5641 ) ;
  assign n5643 = n5380 | n5642 ;
  assign n5644 = ( n5636 & n5642 ) | ( n5636 & n5643 ) | ( n5642 & n5643 ) ;
  assign n5645 = ( n5615 & n5635 ) | ( n5615 & ~n5644 ) | ( n5635 & ~n5644 ) ;
  assign n5646 = ( ~n5635 & n5644 ) | ( ~n5635 & n5645 ) | ( n5644 & n5645 ) ;
  assign n5647 = ( ~n5615 & n5645 ) | ( ~n5615 & n5646 ) | ( n5645 & n5646 ) ;
  assign n5648 = n5425 | n5427 ;
  assign n5649 = n5426 | n5648 ;
  assign n5650 = ~n5647 & n5649 ;
  assign n5651 = n5425 & ~n5647 ;
  assign n5652 = ( n5356 & n5650 ) | ( n5356 & n5651 ) | ( n5650 & n5651 ) ;
  assign n5653 = n5647 & ~n5649 ;
  assign n5654 = ~n5425 & n5647 ;
  assign n5655 = ( ~n5356 & n5653 ) | ( ~n5356 & n5654 ) | ( n5653 & n5654 ) ;
  assign n5656 = n5652 | n5655 ;
  assign n5657 = n3259 & n3641 ;
  assign n5658 = n3266 & n3637 ;
  assign n5659 = n3296 & n3635 ;
  assign n5660 = n3295 & n3635 ;
  assign n5661 = ( n2828 & n5659 ) | ( n2828 & n5660 ) | ( n5659 & n5660 ) ;
  assign n5662 = ( ~n3300 & n3635 ) | ( ~n3300 & n5661 ) | ( n3635 & n5661 ) ;
  assign n5663 = n5658 | n5662 ;
  assign n5664 = n5657 | n5663 ;
  assign n5665 = ( n3643 & n4532 ) | ( n3643 & n5664 ) | ( n4532 & n5664 ) ;
  assign n5666 = ( n482 & n3643 ) | ( n482 & ~n5664 ) | ( n3643 & ~n5664 ) ;
  assign n5667 = ( n482 & n4532 ) | ( n482 & n5666 ) | ( n4532 & n5666 ) ;
  assign n5668 = ~n5665 & n5667 ;
  assign n5669 = n5664 | n5666 ;
  assign n5670 = n482 | n5664 ;
  assign n5671 = ( n4532 & n5669 ) | ( n4532 & n5670 ) | ( n5669 & n5670 ) ;
  assign n5672 = ( ~n482 & n5668 ) | ( ~n482 & n5671 ) | ( n5668 & n5671 ) ;
  assign n5673 = n5656 & n5672 ;
  assign n5674 = n5656 | n5672 ;
  assign n5675 = ~n5673 & n5674 ;
  assign n5676 = n5594 & n5675 ;
  assign n5677 = ~n5594 & n5675 ;
  assign n5678 = ( n5594 & ~n5676 ) | ( n5594 & n5677 ) | ( ~n5676 & n5677 ) ;
  assign n5679 = n5590 & n5678 ;
  assign n5680 = n5678 & ~n5679 ;
  assign n5681 = ( n5590 & ~n5679 ) | ( n5590 & n5680 ) | ( ~n5679 & n5680 ) ;
  assign n5682 = ( n5562 & ~n5567 ) | ( n5562 & n5681 ) | ( ~n5567 & n5681 ) ;
  assign n5683 = ( n5567 & ~n5681 ) | ( n5567 & n5682 ) | ( ~n5681 & n5682 ) ;
  assign n5684 = ( ~n5562 & n5682 ) | ( ~n5562 & n5683 ) | ( n5682 & n5683 ) ;
  assign n5685 = n5482 | n5484 ;
  assign n5686 = ( n5272 & n5482 ) | ( n5272 & n5685 ) | ( n5482 & n5685 ) ;
  assign n5687 = ~n5684 & n5686 ;
  assign n5688 = n5684 & ~n5686 ;
  assign n5689 = n5687 | n5688 ;
  assign n5690 = n200 | n374 ;
  assign n5691 = n365 | n5690 ;
  assign n5692 = n269 | n299 ;
  assign n5693 = n3176 | n5692 ;
  assign n5694 = n155 | n172 ;
  assign n5695 = n174 | n5694 ;
  assign n5696 = n5693 | n5695 ;
  assign n5697 = n249 | n890 ;
  assign n5698 = n673 | n5697 ;
  assign n5699 = n5696 | n5698 ;
  assign n5700 = n5691 | n5699 ;
  assign n5701 = n198 | n311 ;
  assign n5702 = n173 | n242 ;
  assign n5703 = n5701 | n5702 ;
  assign n5704 = n220 | n316 ;
  assign n5705 = n305 | n5704 ;
  assign n5706 = n5703 | n5705 ;
  assign n5707 = n4998 | n5706 ;
  assign n5708 = n5700 | n5707 ;
  assign n5709 = n5689 & n5708 ;
  assign n5710 = n5689 | n5708 ;
  assign n5711 = ~n5709 & n5710 ;
  assign n5712 = n5525 & n5711 ;
  assign n5713 = n5525 & ~n5712 ;
  assign n5714 = n5515 & ~n5712 ;
  assign n5715 = n5515 & n5711 ;
  assign n5716 = ( n5713 & n5714 ) | ( n5713 & n5715 ) | ( n5714 & n5715 ) ;
  assign n5717 = ~n5515 & n5712 ;
  assign n5718 = n5515 | n5711 ;
  assign n5719 = ( n5713 & ~n5717 ) | ( n5713 & n5718 ) | ( ~n5717 & n5718 ) ;
  assign n5720 = ~n5716 & n5719 ;
  assign n5721 = n5271 | n5517 ;
  assign n5722 = n5520 & n5721 ;
  assign n5723 = ~n5720 & n5722 ;
  assign n5724 = n5720 & ~n5722 ;
  assign n5725 = n5723 | n5724 ;
  assign n5726 = n5720 | n5721 ;
  assign n5727 = n5520 & n5726 ;
  assign n5728 = n3340 & ~n5315 ;
  assign n5729 = n3340 & n5303 ;
  assign n5730 = n3340 & ~n5075 ;
  assign n5731 = ( ~n3222 & n3340 ) | ( ~n3222 & n5730 ) | ( n3340 & n5730 ) ;
  assign n5732 = ( ~n5304 & n5729 ) | ( ~n5304 & n5731 ) | ( n5729 & n5731 ) ;
  assign n5733 = ( n5316 & n5728 ) | ( n5316 & n5732 ) | ( n5728 & n5732 ) ;
  assign n5734 = n3333 & n5303 ;
  assign n5735 = n3333 & ~n5075 ;
  assign n5736 = ( ~n3222 & n3333 ) | ( ~n3222 & n5735 ) | ( n3333 & n5735 ) ;
  assign n5737 = ( ~n5304 & n5734 ) | ( ~n5304 & n5736 ) | ( n5734 & n5736 ) ;
  assign n5738 = n5733 | n5737 ;
  assign n5739 = n5732 | n5737 ;
  assign n5740 = ( ~n5534 & n5737 ) | ( ~n5534 & n5739 ) | ( n5737 & n5739 ) ;
  assign n5741 = ( n5093 & n5738 ) | ( n5093 & n5740 ) | ( n5738 & n5740 ) ;
  assign n5742 = ( n5090 & n5738 ) | ( n5090 & n5740 ) | ( n5738 & n5740 ) ;
  assign n5743 = ( n4841 & n5741 ) | ( n4841 & n5742 ) | ( n5741 & n5742 ) ;
  assign n5744 = n3326 & ~n5743 ;
  assign n5745 = ~n3326 & n5743 ;
  assign n5746 = n5744 | n5745 ;
  assign n5747 = n3367 & ~n4854 ;
  assign n5748 = n3285 & n3367 ;
  assign n5749 = n3222 & n5748 ;
  assign n5750 = ( n4855 & n5747 ) | ( n4855 & n5749 ) | ( n5747 & n5749 ) ;
  assign n5751 = n3373 & n4830 ;
  assign n5752 = ( n3387 & n3905 ) | ( n3387 & ~n5080 ) | ( n3905 & ~n5080 ) ;
  assign n5753 = n5751 | n5752 ;
  assign n5754 = n5750 | n5753 ;
  assign n5755 = n1115 | n5754 ;
  assign n5756 = n5750 | n5751 ;
  assign n5757 = n3380 & ~n5080 ;
  assign n5758 = n5752 & n5757 ;
  assign n5759 = n1115 | n5758 ;
  assign n5760 = n5756 | n5759 ;
  assign n5761 = ( ~n5099 & n5755 ) | ( ~n5099 & n5760 ) | ( n5755 & n5760 ) ;
  assign n5762 = n1115 & n5754 ;
  assign n5763 = n1115 & n5758 ;
  assign n5764 = ( n1115 & n5756 ) | ( n1115 & n5763 ) | ( n5756 & n5763 ) ;
  assign n5765 = ( ~n5099 & n5762 ) | ( ~n5099 & n5764 ) | ( n5762 & n5764 ) ;
  assign n5766 = n5761 & ~n5765 ;
  assign n5767 = n5673 | n5675 ;
  assign n5768 = ( n5594 & n5673 ) | ( n5594 & n5767 ) | ( n5673 & n5767 ) ;
  assign n5769 = ( n5356 & n5425 ) | ( n5356 & n5649 ) | ( n5425 & n5649 ) ;
  assign n5770 = n3024 & n3414 ;
  assign n5771 = n2916 & n3412 ;
  assign n5772 = ( ~n2901 & n3412 ) | ( ~n2901 & n5771 ) | ( n3412 & n5771 ) ;
  assign n5773 = ~n2921 & n5772 ;
  assign n5774 = n2828 & n5773 ;
  assign n5775 = ( n2927 & n3412 ) | ( n2927 & n5774 ) | ( n3412 & n5774 ) ;
  assign n5776 = n5770 | n5775 ;
  assign n5777 = n3296 & n3417 ;
  assign n5778 = n3295 & n3417 ;
  assign n5779 = ( n2828 & n5777 ) | ( n2828 & n5778 ) | ( n5777 & n5778 ) ;
  assign n5780 = ( ~n3300 & n3417 ) | ( ~n3300 & n5779 ) | ( n3417 & n5779 ) ;
  assign n5782 = n3423 | n5780 ;
  assign n5783 = n5776 | n5782 ;
  assign n5781 = n5776 | n5780 ;
  assign n5784 = n5781 & n5783 ;
  assign n5785 = ( ~n3360 & n5783 ) | ( ~n3360 & n5784 ) | ( n5783 & n5784 ) ;
  assign n5786 = ~n634 & n5784 ;
  assign n5787 = ~n634 & n5782 ;
  assign n5788 = ( ~n634 & n5776 ) | ( ~n634 & n5787 ) | ( n5776 & n5787 ) ;
  assign n5789 = ( ~n3360 & n5786 ) | ( ~n3360 & n5788 ) | ( n5786 & n5788 ) ;
  assign n5790 = n634 | n5788 ;
  assign n5791 = n634 | n5784 ;
  assign n5792 = ( ~n3360 & n5790 ) | ( ~n3360 & n5791 ) | ( n5790 & n5791 ) ;
  assign n5793 = ( ~n5785 & n5789 ) | ( ~n5785 & n5792 ) | ( n5789 & n5792 ) ;
  assign n5794 = n879 & n2370 ;
  assign n5795 = ( n879 & n2679 ) | ( n879 & n5794 ) | ( n2679 & n5794 ) ;
  assign n5796 = ( n879 & ~n2827 ) | ( n879 & n5795 ) | ( ~n2827 & n5795 ) ;
  assign n5797 = ~n3057 & n5796 ;
  assign n5798 = n3049 & n3477 ;
  assign n5799 = n3110 & n3446 ;
  assign n5800 = ( ~n3106 & n3446 ) | ( ~n3106 & n5799 ) | ( n3446 & n5799 ) ;
  assign n5801 = n5798 | n5800 ;
  assign n5802 = n3033 & n3448 ;
  assign n5803 = n5797 & n5802 ;
  assign n5804 = ( n5797 & n5801 ) | ( n5797 & n5803 ) | ( n5801 & n5803 ) ;
  assign n5805 = ( n3033 & n3452 ) | ( n3033 & n5365 ) | ( n3452 & n5365 ) ;
  assign n5806 = n5797 & n5805 ;
  assign n5807 = ( n5797 & n5801 ) | ( n5797 & n5806 ) | ( n5801 & n5806 ) ;
  assign n5808 = ( ~n3624 & n5804 ) | ( ~n3624 & n5807 ) | ( n5804 & n5807 ) ;
  assign n5809 = n5797 | n5802 ;
  assign n5810 = n5801 | n5809 ;
  assign n5811 = n5797 | n5805 ;
  assign n5812 = n5801 | n5811 ;
  assign n5813 = ( ~n3624 & n5810 ) | ( ~n3624 & n5812 ) | ( n5810 & n5812 ) ;
  assign n5814 = ~n5808 & n5813 ;
  assign n5815 = n879 & n3063 ;
  assign n5816 = ~n5606 & n5815 ;
  assign n5817 = ~n5604 & n5815 ;
  assign n5818 = ~n5602 & n5817 ;
  assign n5819 = ( n3679 & n5816 ) | ( n3679 & n5818 ) | ( n5816 & n5818 ) ;
  assign n5820 = n5642 | n5819 ;
  assign n5821 = ( n5615 & n5819 ) | ( n5615 & n5820 ) | ( n5819 & n5820 ) ;
  assign n5822 = n5814 & ~n5821 ;
  assign n5823 = n5615 | n5819 ;
  assign n5824 = n5814 & ~n5823 ;
  assign n5825 = ( ~n5402 & n5822 ) | ( ~n5402 & n5824 ) | ( n5822 & n5824 ) ;
  assign n5826 = n5793 & n5825 ;
  assign n5827 = ~n5814 & n5821 ;
  assign n5828 = ~n5814 & n5823 ;
  assign n5829 = ( n5402 & n5827 ) | ( n5402 & n5828 ) | ( n5827 & n5828 ) ;
  assign n5830 = ( n5793 & n5826 ) | ( n5793 & n5829 ) | ( n5826 & n5829 ) ;
  assign n5831 = n5793 | n5825 ;
  assign n5832 = n5829 | n5831 ;
  assign n5833 = ~n5830 & n5832 ;
  assign n5834 = n5615 & n5642 ;
  assign n5835 = ( n5402 & n5615 ) | ( n5402 & n5834 ) | ( n5615 & n5834 ) ;
  assign n5836 = n5644 & ~n5835 ;
  assign n5837 = n5615 & ~n5834 ;
  assign n5838 = ~n5402 & n5635 ;
  assign n5839 = n5837 & n5838 ;
  assign n5840 = ( n5635 & n5836 ) | ( n5635 & n5839 ) | ( n5836 & n5839 ) ;
  assign n5841 = n5647 | n5840 ;
  assign n5842 = n5833 & n5841 ;
  assign n5843 = n5833 & n5840 ;
  assign n5844 = ( n5769 & n5842 ) | ( n5769 & n5843 ) | ( n5842 & n5843 ) ;
  assign n5845 = n5833 | n5841 ;
  assign n5846 = n5833 | n5840 ;
  assign n5847 = ( n5769 & n5845 ) | ( n5769 & n5846 ) | ( n5845 & n5846 ) ;
  assign n5848 = ~n5844 & n5847 ;
  assign n5849 = ~n3289 & n3641 ;
  assign n5850 = n3266 & n3635 ;
  assign n5851 = n3259 & n3637 ;
  assign n5852 = n5850 | n5851 ;
  assign n5853 = n5849 | n5852 ;
  assign n5854 = ( ~n3289 & n3643 ) | ( ~n3289 & n3644 ) | ( n3643 & n3644 ) ;
  assign n5855 = n5852 | n5854 ;
  assign n5856 = ( ~n3321 & n5853 ) | ( ~n3321 & n5855 ) | ( n5853 & n5855 ) ;
  assign n5857 = ~n3289 & n5442 ;
  assign n5858 = ( n482 & n5852 ) | ( n482 & n5857 ) | ( n5852 & n5857 ) ;
  assign n5859 = n482 & n5854 ;
  assign n5860 = ( n482 & n5852 ) | ( n482 & n5859 ) | ( n5852 & n5859 ) ;
  assign n5861 = ( ~n3321 & n5858 ) | ( ~n3321 & n5860 ) | ( n5858 & n5860 ) ;
  assign n5862 = n5856 & ~n5861 ;
  assign n5863 = n482 & ~n5857 ;
  assign n5864 = ~n5852 & n5863 ;
  assign n5865 = n482 & ~n5854 ;
  assign n5866 = ~n5852 & n5865 ;
  assign n5867 = ( n3321 & n5864 ) | ( n3321 & n5866 ) | ( n5864 & n5866 ) ;
  assign n5868 = n5862 | n5867 ;
  assign n5869 = n5848 & n5868 ;
  assign n5870 = n5848 & ~n5869 ;
  assign n5871 = ~n5848 & n5868 ;
  assign n5872 = n5870 | n5871 ;
  assign n5873 = n5768 & n5872 ;
  assign n5874 = ~n5768 & n5872 ;
  assign n5875 = ( n5768 & ~n5873 ) | ( n5768 & n5874 ) | ( ~n5873 & n5874 ) ;
  assign n5876 = n5766 & n5875 ;
  assign n5877 = n5766 | n5875 ;
  assign n5878 = ~n5876 & n5877 ;
  assign n5879 = n5746 & n5878 ;
  assign n5880 = n5746 | n5878 ;
  assign n5881 = ~n5879 & n5880 ;
  assign n5882 = n5567 & n5681 ;
  assign n5883 = n5679 | n5882 ;
  assign n5884 = n5881 & n5883 ;
  assign n5885 = n5881 | n5883 ;
  assign n5886 = ~n5884 & n5885 ;
  assign n5887 = n5567 & ~n5882 ;
  assign n5888 = ~n5567 & n5681 ;
  assign n5889 = n5562 & n5888 ;
  assign n5890 = ( n5562 & n5887 ) | ( n5562 & n5889 ) | ( n5887 & n5889 ) ;
  assign n5891 = ( n5684 & n5686 ) | ( n5684 & n5890 ) | ( n5686 & n5890 ) ;
  assign n5892 = ( n5684 & n5886 ) | ( n5684 & ~n5890 ) | ( n5886 & ~n5890 ) ;
  assign n5893 = ( n5686 & n5886 ) | ( n5686 & n5892 ) | ( n5886 & n5892 ) ;
  assign n5894 = ~n5891 & n5893 ;
  assign n5895 = n5890 | n5893 ;
  assign n5896 = ( ~n5886 & n5894 ) | ( ~n5886 & n5895 ) | ( n5894 & n5895 ) ;
  assign n5897 = n248 | n315 ;
  assign n5898 = n265 | n270 ;
  assign n5899 = n277 | n2349 ;
  assign n5900 = n5013 | n5899 ;
  assign n5901 = n503 | n907 ;
  assign n5902 = n5900 | n5901 ;
  assign n5903 = n2594 | n5902 ;
  assign n5904 = n5898 | n5903 ;
  assign n5905 = n235 | n278 ;
  assign n5906 = n366 | n5905 ;
  assign n5907 = n446 | n5906 ;
  assign n5908 = n344 | n352 ;
  assign n5909 = n5907 | n5908 ;
  assign n5910 = n3207 | n5909 ;
  assign n5911 = n5904 | n5910 ;
  assign n5912 = n5897 | n5911 ;
  assign n5913 = n5896 & n5912 ;
  assign n5914 = n5896 & ~n5913 ;
  assign n5915 = ~n5896 & n5912 ;
  assign n5916 = n5914 | n5915 ;
  assign n5917 = n5709 | n5711 ;
  assign n5918 = ( n5525 & n5709 ) | ( n5525 & n5917 ) | ( n5709 & n5917 ) ;
  assign n5919 = n5916 & n5918 ;
  assign n5920 = n5916 | n5918 ;
  assign n5921 = ~n5919 & n5920 ;
  assign n5922 = n5716 & n5921 ;
  assign n5923 = n5716 & ~n5922 ;
  assign n5924 = ( n5921 & ~n5922 ) | ( n5921 & n5923 ) | ( ~n5922 & n5923 ) ;
  assign n5925 = n5727 & n5924 ;
  assign n5926 = n5727 | n5924 ;
  assign n5927 = ~n5925 & n5926 ;
  assign n5928 = n5886 & n5890 ;
  assign n5929 = n5830 | n5844 ;
  assign n5930 = n3033 & n3446 ;
  assign n5931 = n3110 & n3477 ;
  assign n5932 = ( ~n3106 & n3477 ) | ( ~n3106 & n5931 ) | ( n3477 & n5931 ) ;
  assign n5933 = n5930 | n5932 ;
  assign n5934 = n2916 & n3448 ;
  assign n5935 = ( ~n2901 & n3448 ) | ( ~n2901 & n5934 ) | ( n3448 & n5934 ) ;
  assign n5936 = ~n2921 & n5935 ;
  assign n5937 = n2828 & n5936 ;
  assign n5938 = ( n2927 & n3448 ) | ( n2927 & n5937 ) | ( n3448 & n5937 ) ;
  assign n5939 = n5933 | n5938 ;
  assign n5940 = n3452 | n5939 ;
  assign n5941 = ( n3952 & n5939 ) | ( n3952 & n5940 ) | ( n5939 & n5940 ) ;
  assign n5942 = n879 & n3157 ;
  assign n5943 = n3440 & n5942 ;
  assign n5944 = ( n879 & n5939 ) | ( n879 & n5943 ) | ( n5939 & n5943 ) ;
  assign n5945 = n879 & n5939 ;
  assign n5946 = ( n3952 & n5944 ) | ( n3952 & n5945 ) | ( n5944 & n5945 ) ;
  assign n5947 = n5941 & ~n5946 ;
  assign n5948 = ~n874 & n3322 ;
  assign n5949 = ( ~n874 & n3325 ) | ( ~n874 & n5948 ) | ( n3325 & n5948 ) ;
  assign n5950 = n873 & n3322 ;
  assign n5951 = ( n873 & n3325 ) | ( n873 & n5950 ) | ( n3325 & n5950 ) ;
  assign n5952 = ( ~n871 & n5949 ) | ( ~n871 & n5951 ) | ( n5949 & n5951 ) ;
  assign n5953 = ( n34 & n5949 ) | ( n34 & n5951 ) | ( n5949 & n5951 ) ;
  assign n5954 = ( n872 & n5952 ) | ( n872 & n5953 ) | ( n5952 & n5953 ) ;
  assign n5955 = n3049 & n5954 ;
  assign n5956 = n879 & n3049 ;
  assign n5957 = ~n5955 & n5956 ;
  assign n5958 = n3326 & ~n5954 ;
  assign n5959 = ( ~n3049 & n3326 ) | ( ~n3049 & n5958 ) | ( n3326 & n5958 ) ;
  assign n5960 = n5957 | n5959 ;
  assign n5961 = n879 & ~n5939 ;
  assign n5962 = n5960 & n5961 ;
  assign n5963 = n879 & ~n5943 ;
  assign n5964 = ~n5939 & n5963 ;
  assign n5965 = n5960 & n5964 ;
  assign n5966 = ( ~n3952 & n5962 ) | ( ~n3952 & n5965 ) | ( n5962 & n5965 ) ;
  assign n5967 = ( n5947 & n5960 ) | ( n5947 & n5966 ) | ( n5960 & n5966 ) ;
  assign n5968 = n5960 | n5961 ;
  assign n5969 = n5960 | n5964 ;
  assign n5970 = ( ~n3952 & n5968 ) | ( ~n3952 & n5969 ) | ( n5968 & n5969 ) ;
  assign n5971 = n5947 | n5970 ;
  assign n5972 = ~n5967 & n5971 ;
  assign n5973 = n879 & ~n2370 ;
  assign n5974 = ~n2679 & n5973 ;
  assign n5975 = n2827 & n5974 ;
  assign n5976 = ( n879 & n3057 ) | ( n879 & n5975 ) | ( n3057 & n5975 ) ;
  assign n5977 = ~n5802 & n5976 ;
  assign n5978 = ~n5801 & n5977 ;
  assign n5979 = ~n5805 & n5976 ;
  assign n5980 = ~n5801 & n5979 ;
  assign n5981 = ( n3624 & n5978 ) | ( n3624 & n5980 ) | ( n5978 & n5980 ) ;
  assign n5982 = n5814 & n5821 ;
  assign n5983 = n5814 & n5823 ;
  assign n5984 = ( n5402 & n5982 ) | ( n5402 & n5983 ) | ( n5982 & n5983 ) ;
  assign n5985 = n5981 | n5984 ;
  assign n5986 = ~n5972 & n5985 ;
  assign n5987 = n5972 & ~n5985 ;
  assign n5988 = n5986 | n5987 ;
  assign n5989 = n3024 & n3412 ;
  assign n5990 = n3296 & n3414 ;
  assign n5991 = n3295 & n3414 ;
  assign n5992 = ( n2828 & n5990 ) | ( n2828 & n5991 ) | ( n5990 & n5991 ) ;
  assign n5993 = ( ~n3300 & n3414 ) | ( ~n3300 & n5992 ) | ( n3414 & n5992 ) ;
  assign n5994 = n5989 | n5993 ;
  assign n5995 = n3266 & n4687 ;
  assign n5996 = ( n634 & n5994 ) | ( n634 & n5995 ) | ( n5994 & n5995 ) ;
  assign n5997 = ( n3266 & n3424 ) | ( n3266 & n5205 ) | ( n3424 & n5205 ) ;
  assign n5998 = ( n634 & n5994 ) | ( n634 & n5997 ) | ( n5994 & n5997 ) ;
  assign n5999 = ( ~n4190 & n5996 ) | ( ~n4190 & n5998 ) | ( n5996 & n5998 ) ;
  assign n6000 = ( n634 & n3266 ) | ( n634 & n4692 ) | ( n3266 & n4692 ) ;
  assign n6001 = n5994 | n6000 ;
  assign n6002 = ( n3266 & n3431 ) | ( n3266 & n5200 ) | ( n3431 & n5200 ) ;
  assign n6003 = n5994 | n6002 ;
  assign n6004 = ( ~n4190 & n6001 ) | ( ~n4190 & n6003 ) | ( n6001 & n6003 ) ;
  assign n6005 = ~n5999 & n6004 ;
  assign n6006 = ~n5988 & n6005 ;
  assign n6007 = n5988 & ~n6005 ;
  assign n6008 = n6006 | n6007 ;
  assign n6009 = n5929 & ~n6008 ;
  assign n6010 = ~n5929 & n6008 ;
  assign n6011 = n6009 | n6010 ;
  assign n6012 = n3641 & n4830 ;
  assign n6013 = n3259 & n3635 ;
  assign n6014 = ~n3289 & n3637 ;
  assign n6015 = n6013 | n6014 ;
  assign n6016 = n6012 | n6015 ;
  assign n6017 = ( n3643 & n3644 ) | ( n3643 & n4830 ) | ( n3644 & n4830 ) ;
  assign n6018 = n6015 | n6017 ;
  assign n6019 = ( ~n4901 & n6016 ) | ( ~n4901 & n6018 ) | ( n6016 & n6018 ) ;
  assign n6020 = n4830 & n5442 ;
  assign n6021 = ( n482 & n6015 ) | ( n482 & n6020 ) | ( n6015 & n6020 ) ;
  assign n6022 = n482 & n6017 ;
  assign n6023 = ( n482 & n6015 ) | ( n482 & n6022 ) | ( n6015 & n6022 ) ;
  assign n6024 = ( ~n4901 & n6021 ) | ( ~n4901 & n6023 ) | ( n6021 & n6023 ) ;
  assign n6025 = n6019 & ~n6024 ;
  assign n6026 = n482 & ~n6020 ;
  assign n6027 = ~n6015 & n6026 ;
  assign n6028 = n482 & ~n6017 ;
  assign n6029 = ~n6015 & n6028 ;
  assign n6030 = ( n4901 & n6027 ) | ( n4901 & n6029 ) | ( n6027 & n6029 ) ;
  assign n6031 = n6025 | n6030 ;
  assign n6032 = n6011 & n6031 ;
  assign n6033 = n6011 | n6031 ;
  assign n6034 = ~n6032 & n6033 ;
  assign n6035 = n5869 | n5871 ;
  assign n6036 = n5870 | n6035 ;
  assign n6037 = ( n5768 & n5869 ) | ( n5768 & n6036 ) | ( n5869 & n6036 ) ;
  assign n6038 = n6034 & n6037 ;
  assign n6039 = n6034 | n6037 ;
  assign n6040 = ~n6038 & n6039 ;
  assign n6041 = n3367 & ~n5080 ;
  assign n6042 = n3373 & ~n4854 ;
  assign n6043 = n3285 & n3373 ;
  assign n6044 = n3222 & n6043 ;
  assign n6045 = ( n4855 & n6042 ) | ( n4855 & n6044 ) | ( n6042 & n6044 ) ;
  assign n6046 = n6041 | n6045 ;
  assign n6047 = n3380 & n5303 ;
  assign n6048 = n3380 & ~n5075 ;
  assign n6049 = ( ~n3222 & n3380 ) | ( ~n3222 & n6048 ) | ( n3380 & n6048 ) ;
  assign n6050 = ( ~n5304 & n6047 ) | ( ~n5304 & n6049 ) | ( n6047 & n6049 ) ;
  assign n6051 = n3387 | n6050 ;
  assign n6052 = n6046 | n6051 ;
  assign n6053 = n1115 & n6052 ;
  assign n6054 = n1115 & n6050 ;
  assign n6055 = ( n1115 & n6046 ) | ( n1115 & n6054 ) | ( n6046 & n6054 ) ;
  assign n6056 = ( n5325 & n6053 ) | ( n5325 & n6055 ) | ( n6053 & n6055 ) ;
  assign n6057 = n1115 | n6052 ;
  assign n6058 = n1115 | n6050 ;
  assign n6059 = n6046 | n6058 ;
  assign n6060 = ( n5325 & n6057 ) | ( n5325 & n6059 ) | ( n6057 & n6059 ) ;
  assign n6061 = ~n6056 & n6060 ;
  assign n6062 = n6040 & n6061 ;
  assign n6063 = n6040 | n6061 ;
  assign n6064 = ~n6062 & n6063 ;
  assign n6065 = ( n5746 & n5766 ) | ( n5746 & n5875 ) | ( n5766 & n5875 ) ;
  assign n6066 = n6064 | n6065 ;
  assign n6067 = n6064 & n6065 ;
  assign n6068 = n6066 & ~n6067 ;
  assign n6069 = n5884 & n6068 ;
  assign n6070 = ( n5928 & n6068 ) | ( n5928 & n6069 ) | ( n6068 & n6069 ) ;
  assign n6071 = ( n5886 & n6068 ) | ( n5886 & n6069 ) | ( n6068 & n6069 ) ;
  assign n6072 = n5684 & n5686 ;
  assign n6073 = ( n6070 & n6071 ) | ( n6070 & n6072 ) | ( n6071 & n6072 ) ;
  assign n6074 = n5884 | n6068 ;
  assign n6075 = n5928 | n6074 ;
  assign n6076 = n5886 | n6074 ;
  assign n6077 = ( n6072 & n6075 ) | ( n6072 & n6076 ) | ( n6075 & n6076 ) ;
  assign n6078 = ~n6073 & n6077 ;
  assign n6079 = n496 | n3176 ;
  assign n6080 = n313 | n6079 ;
  assign n6081 = n581 | n6080 ;
  assign n6082 = n2786 | n6081 ;
  assign n6083 = n690 | n2733 ;
  assign n6084 = n293 | n347 ;
  assign n6085 = n310 | n6084 ;
  assign n6086 = n6083 | n6085 ;
  assign n6087 = n251 | n6086 ;
  assign n6088 = n240 | n6087 ;
  assign n6089 = n6082 | n6088 ;
  assign n6090 = n6078 | n6089 ;
  assign n6091 = n6078 & n6089 ;
  assign n6092 = n6090 & ~n6091 ;
  assign n6093 = ( n5913 & n5916 ) | ( n5913 & n5918 ) | ( n5916 & n5918 ) ;
  assign n6094 = ( ~n5913 & n6092 ) | ( ~n5913 & n6093 ) | ( n6092 & n6093 ) ;
  assign n6095 = ~n6093 & n6094 ;
  assign n6096 = n5913 | n6092 ;
  assign n6097 = n6093 | n6096 ;
  assign n6098 = ( ~n6092 & n6095 ) | ( ~n6092 & n6097 ) | ( n6095 & n6097 ) ;
  assign n6099 = n5922 | n6098 ;
  assign n6100 = n5922 & n6098 ;
  assign n6101 = n6099 & ~n6100 ;
  assign n6102 = n5726 | n5924 ;
  assign n6103 = n5520 & n6102 ;
  assign n6104 = ~n6101 & n6103 ;
  assign n6105 = n6101 & ~n6103 ;
  assign n6106 = n6104 | n6105 ;
  assign n6107 = n3367 & n5303 ;
  assign n6108 = n3367 & ~n5075 ;
  assign n6109 = ( ~n3222 & n3367 ) | ( ~n3222 & n6108 ) | ( n3367 & n6108 ) ;
  assign n6110 = ( ~n5304 & n6107 ) | ( ~n5304 & n6109 ) | ( n6107 & n6109 ) ;
  assign n6111 = n3373 & ~n5080 ;
  assign n6112 = ( n1115 & n4035 ) | ( n1115 & n6111 ) | ( n4035 & n6111 ) ;
  assign n6113 = ( n4037 & n6110 ) | ( n4037 & n6112 ) | ( n6110 & n6112 ) ;
  assign n6114 = n1115 & n6111 ;
  assign n6115 = ( n1115 & n6110 ) | ( n1115 & n6114 ) | ( n6110 & n6114 ) ;
  assign n6116 = ( n5546 & n6113 ) | ( n5546 & n6115 ) | ( n6113 & n6115 ) ;
  assign n6117 = n4043 | n6111 ;
  assign n6118 = n6110 | n6117 ;
  assign n6119 = n1115 | n6111 ;
  assign n6120 = n6110 | n6119 ;
  assign n6121 = ( n5546 & n6118 ) | ( n5546 & n6120 ) | ( n6118 & n6120 ) ;
  assign n6122 = ~n6116 & n6121 ;
  assign n6123 = ~n3289 & n3635 ;
  assign n6124 = n3637 & n4830 ;
  assign n6125 = n6123 | n6124 ;
  assign n6126 = n3641 & ~n4854 ;
  assign n6127 = n3285 & n3641 ;
  assign n6128 = n3222 & n6127 ;
  assign n6129 = ( n4855 & n6126 ) | ( n4855 & n6128 ) | ( n6126 & n6128 ) ;
  assign n6130 = n6125 | n6129 ;
  assign n6131 = n3643 | n6130 ;
  assign n6132 = ( n4869 & n6130 ) | ( n4869 & n6131 ) | ( n6130 & n6131 ) ;
  assign n6133 = n482 & n6130 ;
  assign n6134 = ( n482 & n3656 ) | ( n482 & n6130 ) | ( n3656 & n6130 ) ;
  assign n6135 = ( n4869 & n6133 ) | ( n4869 & n6134 ) | ( n6133 & n6134 ) ;
  assign n6136 = n6132 & ~n6135 ;
  assign n6137 = n482 & ~n6130 ;
  assign n6138 = n482 & ~n3643 ;
  assign n6139 = ~n6130 & n6138 ;
  assign n6140 = ( ~n4869 & n6137 ) | ( ~n4869 & n6139 ) | ( n6137 & n6139 ) ;
  assign n6141 = n6136 | n6140 ;
  assign n6195 = n3259 & n3417 ;
  assign n6196 = n3266 & n3414 ;
  assign n6197 = n3296 & n3412 ;
  assign n6198 = n3295 & n3412 ;
  assign n6199 = ( n2828 & n6197 ) | ( n2828 & n6198 ) | ( n6197 & n6198 ) ;
  assign n6200 = ( ~n3300 & n3412 ) | ( ~n3300 & n6199 ) | ( n3412 & n6199 ) ;
  assign n6201 = n6196 | n6200 ;
  assign n6202 = n6195 | n6201 ;
  assign n6203 = ( n634 & n3424 ) | ( n634 & n6202 ) | ( n3424 & n6202 ) ;
  assign n6204 = n634 & n6202 ;
  assign n6205 = ( n4532 & n6203 ) | ( n4532 & n6204 ) | ( n6203 & n6204 ) ;
  assign n6206 = n3431 | n6202 ;
  assign n6207 = n634 | n6202 ;
  assign n6208 = ( n4532 & n6206 ) | ( n4532 & n6207 ) | ( n6206 & n6207 ) ;
  assign n6209 = ~n6205 & n6208 ;
  assign n6142 = n3110 & n5954 ;
  assign n6143 = ( ~n3106 & n5954 ) | ( ~n3106 & n6142 ) | ( n5954 & n6142 ) ;
  assign n6144 = n3326 & ~n6143 ;
  assign n6145 = n3111 | n6143 ;
  assign n6146 = n879 & ~n6145 ;
  assign n6147 = n6144 | n6146 ;
  assign n6148 = n5955 & n6144 ;
  assign n6149 = ( n5955 & n6146 ) | ( n5955 & n6148 ) | ( n6146 & n6148 ) ;
  assign n6150 = ( n5960 & n6147 ) | ( n5960 & n6149 ) | ( n6147 & n6149 ) ;
  assign n6151 = ( n5965 & n6147 ) | ( n5965 & n6149 ) | ( n6147 & n6149 ) ;
  assign n6152 = ( n5962 & n6147 ) | ( n5962 & n6149 ) | ( n6147 & n6149 ) ;
  assign n6153 = ( ~n3952 & n6151 ) | ( ~n3952 & n6152 ) | ( n6151 & n6152 ) ;
  assign n6154 = ( n5947 & n6150 ) | ( n5947 & n6153 ) | ( n6150 & n6153 ) ;
  assign n6155 = n5955 | n5965 ;
  assign n6156 = n5955 | n5962 ;
  assign n6157 = ( ~n3952 & n6155 ) | ( ~n3952 & n6156 ) | ( n6155 & n6156 ) ;
  assign n6158 = n5955 | n5959 ;
  assign n6159 = n5957 | n6158 ;
  assign n6160 = ( n5947 & n6157 ) | ( n5947 & n6159 ) | ( n6157 & n6159 ) ;
  assign n6161 = ~n6154 & n6160 ;
  assign n6162 = n6147 & ~n6149 ;
  assign n6163 = ~n5960 & n6162 ;
  assign n6164 = ~n5965 & n6162 ;
  assign n6165 = ~n5962 & n6162 ;
  assign n6166 = ( n3952 & n6164 ) | ( n3952 & n6165 ) | ( n6164 & n6165 ) ;
  assign n6167 = ( ~n5947 & n6163 ) | ( ~n5947 & n6166 ) | ( n6163 & n6166 ) ;
  assign n6168 = n6161 | n6167 ;
  assign n6169 = n3033 & n3477 ;
  assign n6170 = n2916 & n3446 ;
  assign n6171 = ( ~n2901 & n3446 ) | ( ~n2901 & n6170 ) | ( n3446 & n6170 ) ;
  assign n6172 = ~n2921 & n6171 ;
  assign n6173 = n2828 & n6172 ;
  assign n6174 = ( n2927 & n3446 ) | ( n2927 & n6173 ) | ( n3446 & n6173 ) ;
  assign n6175 = n6169 | n6174 ;
  assign n6176 = n3024 & n3448 ;
  assign n6177 = ( n3024 & n3452 ) | ( n3024 & n5365 ) | ( n3452 & n5365 ) ;
  assign n6178 = n6176 & n6177 ;
  assign n6179 = n6175 | n6178 ;
  assign n6180 = n879 | n6179 ;
  assign n6181 = n879 | n5365 ;
  assign n6182 = n879 | n3452 ;
  assign n6183 = ( n3024 & n6181 ) | ( n3024 & n6182 ) | ( n6181 & n6182 ) ;
  assign n6184 = n6175 | n6183 ;
  assign n6185 = ( n3896 & n6180 ) | ( n3896 & n6184 ) | ( n6180 & n6184 ) ;
  assign n6186 = n879 & n6179 ;
  assign n6187 = n879 & n5365 ;
  assign n6188 = ( n3024 & n5943 ) | ( n3024 & n6187 ) | ( n5943 & n6187 ) ;
  assign n6189 = ( n879 & n6175 ) | ( n879 & n6188 ) | ( n6175 & n6188 ) ;
  assign n6190 = ( n3896 & n6186 ) | ( n3896 & n6189 ) | ( n6186 & n6189 ) ;
  assign n6191 = n6185 & ~n6190 ;
  assign n6192 = n6167 & n6191 ;
  assign n6193 = ( n6161 & n6191 ) | ( n6161 & n6192 ) | ( n6191 & n6192 ) ;
  assign n6194 = n6168 & ~n6193 ;
  assign n6213 = n6191 & ~n6193 ;
  assign n6214 = n6194 | n6213 ;
  assign n6215 = n6209 & n6214 ;
  assign n6210 = n6191 | n6209 ;
  assign n6211 = ( ~n6193 & n6209 ) | ( ~n6193 & n6210 ) | ( n6209 & n6210 ) ;
  assign n6212 = n6194 | n6211 ;
  assign n6217 = ( n5972 & n5985 ) | ( n5972 & n6005 ) | ( n5985 & n6005 ) ;
  assign n6218 = ( n6141 & n6212 ) | ( n6141 & ~n6217 ) | ( n6212 & ~n6217 ) ;
  assign n6219 = n6141 & ~n6217 ;
  assign n6220 = ( ~n6215 & n6218 ) | ( ~n6215 & n6219 ) | ( n6218 & n6219 ) ;
  assign n6216 = n6212 & ~n6215 ;
  assign n6221 = ( ~n6216 & n6217 ) | ( ~n6216 & n6220 ) | ( n6217 & n6220 ) ;
  assign n6222 = ( ~n6141 & n6220 ) | ( ~n6141 & n6221 ) | ( n6220 & n6221 ) ;
  assign n6223 = ( n5929 & n6008 ) | ( n5929 & n6031 ) | ( n6008 & n6031 ) ;
  assign n6224 = ( n6122 & n6222 ) | ( n6122 & ~n6223 ) | ( n6222 & ~n6223 ) ;
  assign n6225 = ( ~n6222 & n6223 ) | ( ~n6222 & n6224 ) | ( n6223 & n6224 ) ;
  assign n6226 = ( ~n6122 & n6224 ) | ( ~n6122 & n6225 ) | ( n6224 & n6225 ) ;
  assign n6227 = n6034 | n6061 ;
  assign n6228 = ( n6037 & n6061 ) | ( n6037 & n6227 ) | ( n6061 & n6227 ) ;
  assign n6229 = n6226 & n6228 ;
  assign n6230 = n6038 & n6226 ;
  assign n6231 = ( n6040 & n6229 ) | ( n6040 & n6230 ) | ( n6229 & n6230 ) ;
  assign n6232 = n6226 | n6228 ;
  assign n6233 = n6038 | n6226 ;
  assign n6234 = ( n6040 & n6232 ) | ( n6040 & n6233 ) | ( n6232 & n6233 ) ;
  assign n6235 = ~n6231 & n6234 ;
  assign n6236 = n6067 & n6235 ;
  assign n6237 = ( n6073 & n6235 ) | ( n6073 & n6236 ) | ( n6235 & n6236 ) ;
  assign n6238 = n6067 | n6235 ;
  assign n6239 = n6073 | n6238 ;
  assign n6240 = ~n6237 & n6239 ;
  assign n6241 = n407 | n2292 ;
  assign n6242 = n257 | n278 ;
  assign n6243 = n131 | n6242 ;
  assign n6244 = n367 | n858 ;
  assign n6245 = n6243 | n6244 ;
  assign n6246 = n6241 | n6245 ;
  assign n6247 = n541 | n6246 ;
  assign n6248 = n5291 | n6247 ;
  assign n6249 = n347 | n2302 ;
  assign n6250 = n5496 | n6249 ;
  assign n6251 = n368 | n372 ;
  assign n6252 = n125 | n6251 ;
  assign n6253 = n6250 | n6252 ;
  assign n6254 = n3253 | n6253 ;
  assign n6255 = n6248 | n6254 ;
  assign n6256 = n6240 | n6255 ;
  assign n6257 = n6240 & n6255 ;
  assign n6258 = n6256 & ~n6257 ;
  assign n6259 = n5913 | n6091 ;
  assign n6260 = ( n6091 & n6092 ) | ( n6091 & n6259 ) | ( n6092 & n6259 ) ;
  assign n6261 = n6258 & n6260 ;
  assign n6262 = n6091 | n6092 ;
  assign n6263 = n6258 & n6262 ;
  assign n6264 = ( n5919 & n6261 ) | ( n5919 & n6263 ) | ( n6261 & n6263 ) ;
  assign n6265 = n6258 | n6260 ;
  assign n6266 = n6258 | n6262 ;
  assign n6267 = ( n5919 & n6265 ) | ( n5919 & n6266 ) | ( n6265 & n6266 ) ;
  assign n6268 = ~n6264 & n6267 ;
  assign n6269 = n5922 | n6268 ;
  assign n6270 = ( n6098 & n6268 ) | ( n6098 & n6269 ) | ( n6268 & n6269 ) ;
  assign n6271 = n5922 & n6268 ;
  assign n6272 = n6098 & n6271 ;
  assign n6273 = n6270 & ~n6272 ;
  assign n6274 = n6101 | n6102 ;
  assign n6275 = n5520 & n6274 ;
  assign n6276 = ~n6273 & n6275 ;
  assign n6277 = n6273 & ~n6275 ;
  assign n6278 = n6276 | n6277 ;
  assign n6279 = ( n5919 & n6260 ) | ( n5919 & n6262 ) | ( n6260 & n6262 ) ;
  assign n6280 = n6212 & n6217 ;
  assign n6281 = n5972 & n6209 ;
  assign n6282 = n6005 & n6209 ;
  assign n6283 = ( n5985 & n6281 ) | ( n5985 & n6282 ) | ( n6281 & n6282 ) ;
  assign n6284 = n6214 & n6283 ;
  assign n6285 = ( n6217 & ~n6280 ) | ( n6217 & n6284 ) | ( ~n6280 & n6284 ) ;
  assign n6286 = ~n6215 & n6280 ;
  assign n6287 = n6216 & ~n6286 ;
  assign n6288 = n6285 | n6287 ;
  assign n6289 = n3387 & ~n5315 ;
  assign n6290 = n3387 & n5303 ;
  assign n6291 = n3387 & ~n5075 ;
  assign n6292 = ( ~n3222 & n3387 ) | ( ~n3222 & n6291 ) | ( n3387 & n6291 ) ;
  assign n6293 = ( ~n5304 & n6290 ) | ( ~n5304 & n6292 ) | ( n6290 & n6292 ) ;
  assign n6294 = ( n5316 & n6289 ) | ( n5316 & n6293 ) | ( n6289 & n6293 ) ;
  assign n6295 = n3373 & n5303 ;
  assign n6296 = n3373 & ~n5075 ;
  assign n6297 = ( ~n3222 & n3373 ) | ( ~n3222 & n6296 ) | ( n3373 & n6296 ) ;
  assign n6298 = ( ~n5304 & n6295 ) | ( ~n5304 & n6297 ) | ( n6295 & n6297 ) ;
  assign n6299 = n6294 | n6298 ;
  assign n6300 = n6293 | n6298 ;
  assign n6301 = ( ~n5534 & n6298 ) | ( ~n5534 & n6300 ) | ( n6298 & n6300 ) ;
  assign n6302 = ( n5093 & n6299 ) | ( n5093 & n6301 ) | ( n6299 & n6301 ) ;
  assign n6303 = ( n5090 & n6299 ) | ( n5090 & n6301 ) | ( n6299 & n6301 ) ;
  assign n6304 = ( n4841 & n6302 ) | ( n4841 & n6303 ) | ( n6302 & n6303 ) ;
  assign n6305 = ~n1115 & n6304 ;
  assign n6306 = n1115 & ~n6304 ;
  assign n6307 = n6305 | n6306 ;
  assign n6308 = ~n6209 & n6307 ;
  assign n6309 = ( ~n6214 & n6307 ) | ( ~n6214 & n6308 ) | ( n6307 & n6308 ) ;
  assign n6310 = n6280 & n6309 ;
  assign n6311 = n6140 & n6307 ;
  assign n6312 = ( n6136 & n6307 ) | ( n6136 & n6311 ) | ( n6307 & n6311 ) ;
  assign n6313 = ( n6286 & n6307 ) | ( n6286 & n6312 ) | ( n6307 & n6312 ) ;
  assign n6314 = ( n6288 & n6310 ) | ( n6288 & n6313 ) | ( n6310 & n6313 ) ;
  assign n6315 = n6286 | n6307 ;
  assign n6316 = n6140 | n6307 ;
  assign n6317 = n6136 | n6316 ;
  assign n6318 = n6286 | n6317 ;
  assign n6319 = ( n6288 & n6315 ) | ( n6288 & n6318 ) | ( n6315 & n6318 ) ;
  assign n6320 = ~n6314 & n6319 ;
  assign n6419 = n6193 | n6209 ;
  assign n6420 = ( n6193 & n6214 ) | ( n6193 & n6419 ) | ( n6214 & n6419 ) ;
  assign n6321 = n6143 | n6149 ;
  assign n6322 = n6143 | n6144 ;
  assign n6323 = n6146 | n6322 ;
  assign n6324 = ( n5960 & n6321 ) | ( n5960 & n6323 ) | ( n6321 & n6323 ) ;
  assign n6325 = ( n5965 & n6321 ) | ( n5965 & n6323 ) | ( n6321 & n6323 ) ;
  assign n6326 = ( n5962 & n6321 ) | ( n5962 & n6323 ) | ( n6321 & n6323 ) ;
  assign n6327 = ( ~n3952 & n6325 ) | ( ~n3952 & n6326 ) | ( n6325 & n6326 ) ;
  assign n6328 = ( n5947 & n6324 ) | ( n5947 & n6327 ) | ( n6324 & n6327 ) ;
  assign n6329 = ( ~n3033 & n3326 ) | ( ~n3033 & n5958 ) | ( n3326 & n5958 ) ;
  assign n6330 = n3033 & n5954 ;
  assign n6331 = n879 & n3033 ;
  assign n6332 = ~n6330 & n6331 ;
  assign n6333 = n6329 | n6332 ;
  assign n6334 = n6323 & n6333 ;
  assign n6335 = n6143 & n6329 ;
  assign n6336 = ( n6143 & n6332 ) | ( n6143 & n6335 ) | ( n6332 & n6335 ) ;
  assign n6337 = ( n6149 & n6333 ) | ( n6149 & n6336 ) | ( n6333 & n6336 ) ;
  assign n6338 = ( n5960 & n6334 ) | ( n5960 & n6337 ) | ( n6334 & n6337 ) ;
  assign n6339 = ( n5965 & n6334 ) | ( n5965 & n6337 ) | ( n6334 & n6337 ) ;
  assign n6340 = ( n5962 & n6334 ) | ( n5962 & n6337 ) | ( n6334 & n6337 ) ;
  assign n6341 = ( ~n3952 & n6339 ) | ( ~n3952 & n6340 ) | ( n6339 & n6340 ) ;
  assign n6342 = ( n5947 & n6338 ) | ( n5947 & n6341 ) | ( n6338 & n6341 ) ;
  assign n6343 = n6328 & ~n6342 ;
  assign n6344 = ~n6323 & n6333 ;
  assign n6345 = n6333 & ~n6336 ;
  assign n6346 = ~n6149 & n6345 ;
  assign n6347 = ( ~n5960 & n6344 ) | ( ~n5960 & n6346 ) | ( n6344 & n6346 ) ;
  assign n6348 = ( ~n5965 & n6344 ) | ( ~n5965 & n6346 ) | ( n6344 & n6346 ) ;
  assign n6349 = ( ~n5962 & n6344 ) | ( ~n5962 & n6346 ) | ( n6344 & n6346 ) ;
  assign n6350 = ( n3952 & n6348 ) | ( n3952 & n6349 ) | ( n6348 & n6349 ) ;
  assign n6351 = ( ~n5947 & n6347 ) | ( ~n5947 & n6350 ) | ( n6347 & n6350 ) ;
  assign n6352 = n6343 | n6351 ;
  assign n6353 = n3024 & n3446 ;
  assign n6354 = n2916 & n3477 ;
  assign n6355 = ( ~n2901 & n3477 ) | ( ~n2901 & n6354 ) | ( n3477 & n6354 ) ;
  assign n6356 = ~n2921 & n6355 ;
  assign n6357 = n2828 & n6356 ;
  assign n6358 = ( n2927 & n3477 ) | ( n2927 & n6357 ) | ( n3477 & n6357 ) ;
  assign n6359 = n6353 | n6358 ;
  assign n6360 = n3296 & n3448 ;
  assign n6361 = n3295 & n3448 ;
  assign n6362 = ( n2828 & n6360 ) | ( n2828 & n6361 ) | ( n6360 & n6361 ) ;
  assign n6363 = ( ~n3300 & n3448 ) | ( ~n3300 & n6362 ) | ( n3448 & n6362 ) ;
  assign n6365 = n3452 | n6363 ;
  assign n6366 = n6359 | n6365 ;
  assign n6364 = n6359 | n6363 ;
  assign n6367 = n6364 & n6366 ;
  assign n6368 = ( ~n3360 & n6366 ) | ( ~n3360 & n6367 ) | ( n6366 & n6367 ) ;
  assign n6369 = ~n879 & n6367 ;
  assign n6370 = ~n879 & n6365 ;
  assign n6371 = ( ~n879 & n6359 ) | ( ~n879 & n6370 ) | ( n6359 & n6370 ) ;
  assign n6372 = ( ~n3360 & n6369 ) | ( ~n3360 & n6371 ) | ( n6369 & n6371 ) ;
  assign n6373 = n879 | n6371 ;
  assign n6374 = n879 | n6367 ;
  assign n6375 = ( ~n3360 & n6373 ) | ( ~n3360 & n6374 ) | ( n6373 & n6374 ) ;
  assign n6376 = ( ~n6368 & n6372 ) | ( ~n6368 & n6375 ) | ( n6372 & n6375 ) ;
  assign n6377 = n6351 & n6376 ;
  assign n6378 = ( n6343 & n6376 ) | ( n6343 & n6377 ) | ( n6376 & n6377 ) ;
  assign n6379 = n6352 & ~n6378 ;
  assign n6380 = n6376 & ~n6378 ;
  assign n6381 = n6379 | n6380 ;
  assign n6382 = n3266 & n3412 ;
  assign n6383 = n3259 & n3414 ;
  assign n6384 = n6382 | n6383 ;
  assign n6385 = ~n3289 & n4687 ;
  assign n6386 = ( n634 & n6384 ) | ( n634 & n6385 ) | ( n6384 & n6385 ) ;
  assign n6387 = ( ~n3289 & n3424 ) | ( ~n3289 & n5205 ) | ( n3424 & n5205 ) ;
  assign n6388 = ( n634 & n6384 ) | ( n634 & n6387 ) | ( n6384 & n6387 ) ;
  assign n6389 = ( ~n3321 & n6386 ) | ( ~n3321 & n6388 ) | ( n6386 & n6388 ) ;
  assign n6390 = ( n634 & ~n3289 ) | ( n634 & n4692 ) | ( ~n3289 & n4692 ) ;
  assign n6391 = n6384 | n6390 ;
  assign n6392 = ( ~n3289 & n3431 ) | ( ~n3289 & n5200 ) | ( n3431 & n5200 ) ;
  assign n6393 = n6384 | n6392 ;
  assign n6394 = ( ~n3321 & n6391 ) | ( ~n3321 & n6393 ) | ( n6391 & n6393 ) ;
  assign n6395 = ~n6389 & n6394 ;
  assign n6396 = n6381 & n6395 ;
  assign n6397 = n6376 | n6395 ;
  assign n6398 = ( ~n6378 & n6395 ) | ( ~n6378 & n6397 ) | ( n6395 & n6397 ) ;
  assign n6399 = n6379 | n6398 ;
  assign n6400 = ~n6396 & n6399 ;
  assign n6401 = n3637 & ~n4854 ;
  assign n6402 = n3285 & n3637 ;
  assign n6403 = n3222 & n6402 ;
  assign n6404 = ( n4855 & n6401 ) | ( n4855 & n6403 ) | ( n6401 & n6403 ) ;
  assign n6405 = n3641 & ~n5080 ;
  assign n6406 = n3635 & n4830 ;
  assign n6407 = n6405 | n6406 ;
  assign n6408 = n6404 | n6407 ;
  assign n6409 = n3643 | n6408 ;
  assign n6410 = ( ~n5099 & n6408 ) | ( ~n5099 & n6409 ) | ( n6408 & n6409 ) ;
  assign n6411 = n482 & n6408 ;
  assign n6412 = ( n482 & n3656 ) | ( n482 & n6408 ) | ( n3656 & n6408 ) ;
  assign n6413 = ( ~n5099 & n6411 ) | ( ~n5099 & n6412 ) | ( n6411 & n6412 ) ;
  assign n6414 = n6410 & ~n6413 ;
  assign n6415 = n482 & ~n6408 ;
  assign n6416 = n6138 & ~n6408 ;
  assign n6417 = ( n5099 & n6415 ) | ( n5099 & n6416 ) | ( n6415 & n6416 ) ;
  assign n6418 = n6414 | n6417 ;
  assign n6421 = ( n6400 & n6418 ) | ( n6400 & n6420 ) | ( n6418 & n6420 ) ;
  assign n6422 = ( n6400 & n6418 ) | ( n6400 & ~n6421 ) | ( n6418 & ~n6421 ) ;
  assign n6423 = ( n6420 & ~n6421 ) | ( n6420 & n6422 ) | ( ~n6421 & n6422 ) ;
  assign n6424 = n6320 & n6423 ;
  assign n6425 = n6320 | n6423 ;
  assign n6426 = ~n6424 & n6425 ;
  assign n6427 = n6222 & n6223 ;
  assign n6428 = n6223 & ~n6427 ;
  assign n6429 = n6222 & ~n6223 ;
  assign n6430 = n6122 | n6220 ;
  assign n6431 = ~n6122 & n6141 ;
  assign n6432 = ( n6221 & n6430 ) | ( n6221 & ~n6431 ) | ( n6430 & ~n6431 ) ;
  assign n6433 = ( n6122 & n6223 ) | ( n6122 & n6432 ) | ( n6223 & n6432 ) ;
  assign n6434 = ( n6427 & n6429 ) | ( n6427 & n6433 ) | ( n6429 & n6433 ) ;
  assign n6435 = n6427 | n6433 ;
  assign n6436 = ( n6428 & n6434 ) | ( n6428 & n6435 ) | ( n6434 & n6435 ) ;
  assign n6437 = n6426 & n6436 ;
  assign n6438 = n6426 | n6436 ;
  assign n6439 = ~n6437 & n6438 ;
  assign n6440 = ( n6038 & n6040 ) | ( n6038 & n6228 ) | ( n6040 & n6228 ) ;
  assign n6441 = n6226 & n6439 ;
  assign n6442 = n6440 & n6441 ;
  assign n6443 = ( n6235 & n6439 ) | ( n6235 & n6442 ) | ( n6439 & n6442 ) ;
  assign n6444 = n6439 & n6442 ;
  assign n6445 = ( n6067 & n6443 ) | ( n6067 & n6444 ) | ( n6443 & n6444 ) ;
  assign n6446 = ( n6073 & n6443 ) | ( n6073 & n6445 ) | ( n6443 & n6445 ) ;
  assign n6447 = n6226 | n6439 ;
  assign n6448 = ( n6439 & n6440 ) | ( n6439 & n6447 ) | ( n6440 & n6447 ) ;
  assign n6449 = n6235 | n6448 ;
  assign n6450 = ( n6067 & n6448 ) | ( n6067 & n6449 ) | ( n6448 & n6449 ) ;
  assign n6451 = ( n6073 & n6449 ) | ( n6073 & n6450 ) | ( n6449 & n6450 ) ;
  assign n6452 = ~n6446 & n6451 ;
  assign n6453 = n542 | n781 ;
  assign n6454 = n418 | n6453 ;
  assign n6455 = n2736 | n6454 ;
  assign n6456 = n392 | n2349 ;
  assign n6457 = n582 | n2302 ;
  assign n6458 = n6456 | n6457 ;
  assign n6459 = n301 | n6458 ;
  assign n6460 = n6455 | n6459 ;
  assign n6461 = n216 | n6460 ;
  assign n6462 = n174 | n576 ;
  assign n6463 = n2775 | n6462 ;
  assign n6464 = n4822 | n6463 ;
  assign n6465 = n4955 | n6464 ;
  assign n6466 = n4943 | n6465 ;
  assign n6467 = n6461 | n6466 ;
  assign n6468 = n227 | n290 ;
  assign n6469 = n202 | n358 ;
  assign n6470 = n6468 | n6469 ;
  assign n6471 = n167 | n6470 ;
  assign n6472 = n6467 | n6471 ;
  assign n6473 = n6452 | n6472 ;
  assign n6474 = n6452 & n6472 ;
  assign n6475 = n6473 & ~n6474 ;
  assign n6476 = n6257 | n6258 ;
  assign n6477 = n6475 & n6476 ;
  assign n6478 = n6257 & n6475 ;
  assign n6479 = ( n6279 & n6477 ) | ( n6279 & n6478 ) | ( n6477 & n6478 ) ;
  assign n6480 = n6475 | n6476 ;
  assign n6481 = n6257 | n6475 ;
  assign n6482 = ( n6279 & n6480 ) | ( n6279 & n6481 ) | ( n6480 & n6481 ) ;
  assign n6483 = ~n6479 & n6482 ;
  assign n6484 = n6268 & n6483 ;
  assign n6485 = n6100 & n6484 ;
  assign n6486 = n6272 | n6483 ;
  assign n6487 = ~n6485 & n6486 ;
  assign n6488 = ( n5520 & n6273 ) | ( n5520 & n6275 ) | ( n6273 & n6275 ) ;
  assign n6489 = ~n6487 & n6488 ;
  assign n6490 = n6487 & ~n6488 ;
  assign n6491 = n6489 | n6490 ;
  assign n6492 = n6474 | n6479 ;
  assign n6641 = n6314 | n6423 ;
  assign n6642 = ( n6314 & n6320 ) | ( n6314 & n6641 ) | ( n6320 & n6641 ) ;
  assign n6493 = n6400 & n6420 ;
  assign n6494 = n6400 & ~n6493 ;
  assign n6495 = n6418 & n6419 ;
  assign n6496 = n6193 & n6418 ;
  assign n6497 = ( n6214 & n6495 ) | ( n6214 & n6496 ) | ( n6495 & n6496 ) ;
  assign n6498 = ~n6400 & n6497 ;
  assign n6499 = n3637 & ~n5080 ;
  assign n6500 = n3635 & ~n4854 ;
  assign n6501 = n3285 & n3635 ;
  assign n6502 = n3222 & n6501 ;
  assign n6503 = ( n4855 & n6500 ) | ( n4855 & n6502 ) | ( n6500 & n6502 ) ;
  assign n6504 = n6499 | n6503 ;
  assign n6505 = n3641 & n5303 ;
  assign n6506 = n3641 & ~n5075 ;
  assign n6507 = ( ~n3222 & n3641 ) | ( ~n3222 & n6506 ) | ( n3641 & n6506 ) ;
  assign n6508 = ( ~n5304 & n6505 ) | ( ~n5304 & n6507 ) | ( n6505 & n6507 ) ;
  assign n6509 = ( n3643 & n3644 ) | ( n3643 & n5303 ) | ( n3644 & n5303 ) ;
  assign n6510 = ( n3643 & n3644 ) | ( n3643 & ~n5075 ) | ( n3644 & ~n5075 ) ;
  assign n6511 = n3643 | n3644 ;
  assign n6512 = ( ~n3222 & n6510 ) | ( ~n3222 & n6511 ) | ( n6510 & n6511 ) ;
  assign n6513 = ( ~n5304 & n6509 ) | ( ~n5304 & n6512 ) | ( n6509 & n6512 ) ;
  assign n6514 = n6508 & n6513 ;
  assign n6515 = n6504 | n6514 ;
  assign n6516 = n482 | n6515 ;
  assign n6517 = n482 | n6513 ;
  assign n6518 = n6504 | n6517 ;
  assign n6519 = ( n5325 & n6516 ) | ( n5325 & n6518 ) | ( n6516 & n6518 ) ;
  assign n6520 = n482 & n6515 ;
  assign n6521 = n482 & n6513 ;
  assign n6522 = ( n482 & n6504 ) | ( n482 & n6521 ) | ( n6504 & n6521 ) ;
  assign n6523 = ( n5325 & n6520 ) | ( n5325 & n6522 ) | ( n6520 & n6522 ) ;
  assign n6524 = n6519 & ~n6523 ;
  assign n6525 = n6193 & n6524 ;
  assign n6526 = n6209 & n6524 ;
  assign n6527 = ( n6193 & n6524 ) | ( n6193 & n6526 ) | ( n6524 & n6526 ) ;
  assign n6528 = ( n6214 & n6525 ) | ( n6214 & n6527 ) | ( n6525 & n6527 ) ;
  assign n6529 = n6400 & n6528 ;
  assign n6530 = ( n6498 & n6524 ) | ( n6498 & n6529 ) | ( n6524 & n6529 ) ;
  assign n6531 = n6418 & n6524 ;
  assign n6532 = ( n6418 & n6524 ) | ( n6418 & n6527 ) | ( n6524 & n6527 ) ;
  assign n6533 = ( n6418 & n6524 ) | ( n6418 & n6525 ) | ( n6524 & n6525 ) ;
  assign n6534 = ( n6214 & n6532 ) | ( n6214 & n6533 ) | ( n6532 & n6533 ) ;
  assign n6535 = ( n6400 & n6531 ) | ( n6400 & n6534 ) | ( n6531 & n6534 ) ;
  assign n6536 = ( n6494 & n6530 ) | ( n6494 & n6535 ) | ( n6530 & n6535 ) ;
  assign n6537 = n6419 | n6524 ;
  assign n6538 = n6193 | n6524 ;
  assign n6539 = ( n6214 & n6537 ) | ( n6214 & n6538 ) | ( n6537 & n6538 ) ;
  assign n6540 = ( n6400 & n6524 ) | ( n6400 & n6539 ) | ( n6524 & n6539 ) ;
  assign n6541 = n6498 | n6540 ;
  assign n6542 = n6418 | n6539 ;
  assign n6543 = n6418 | n6524 ;
  assign n6544 = ( n6400 & n6542 ) | ( n6400 & n6543 ) | ( n6542 & n6543 ) ;
  assign n6545 = ( n6494 & n6541 ) | ( n6494 & n6544 ) | ( n6541 & n6544 ) ;
  assign n6546 = ~n6536 & n6545 ;
  assign n6547 = n3266 & n3448 ;
  assign n6548 = n3024 & n3477 ;
  assign n6549 = n3296 & n3446 ;
  assign n6550 = n3295 & n3446 ;
  assign n6551 = ( n2828 & n6549 ) | ( n2828 & n6550 ) | ( n6549 & n6550 ) ;
  assign n6552 = ( ~n3300 & n3446 ) | ( ~n3300 & n6551 ) | ( n3446 & n6551 ) ;
  assign n6553 = n6548 | n6552 ;
  assign n6554 = n6547 | n6553 ;
  assign n6555 = ( n3266 & n3452 ) | ( n3266 & n5365 ) | ( n3452 & n5365 ) ;
  assign n6556 = n6553 | n6555 ;
  assign n6557 = ( ~n4190 & n6554 ) | ( ~n4190 & n6556 ) | ( n6554 & n6556 ) ;
  assign n6558 = n3266 & n5369 ;
  assign n6559 = ( n879 & n6553 ) | ( n879 & n6558 ) | ( n6553 & n6558 ) ;
  assign n6560 = n879 & n6555 ;
  assign n6561 = ( n879 & n6553 ) | ( n879 & n6560 ) | ( n6553 & n6560 ) ;
  assign n6562 = ( ~n4190 & n6559 ) | ( ~n4190 & n6561 ) | ( n6559 & n6561 ) ;
  assign n6563 = n6557 & ~n6562 ;
  assign n6564 = n879 & ~n6558 ;
  assign n6565 = ~n6553 & n6564 ;
  assign n6566 = n879 & ~n6555 ;
  assign n6567 = ~n6553 & n6566 ;
  assign n6568 = ( n4190 & n6565 ) | ( n4190 & n6567 ) | ( n6565 & n6567 ) ;
  assign n6569 = n6563 | n6568 ;
  assign n6570 = n879 & ~n2917 ;
  assign n6571 = ~n2921 & n6570 ;
  assign n6572 = n2828 & n6571 ;
  assign n6573 = ( n879 & n2927 ) | ( n879 & n6572 ) | ( n2927 & n6572 ) ;
  assign n6574 = n1115 | n3326 ;
  assign n6575 = n1115 & n3326 ;
  assign n6576 = n6574 & ~n6575 ;
  assign n6577 = n879 & n6576 ;
  assign n6578 = n6571 & n6576 ;
  assign n6579 = n2828 & n6578 ;
  assign n6580 = ( n2927 & n6577 ) | ( n2927 & n6579 ) | ( n6577 & n6579 ) ;
  assign n6581 = n6576 & ~n6579 ;
  assign n6582 = n6576 & ~n6577 ;
  assign n6583 = ( ~n2927 & n6581 ) | ( ~n2927 & n6582 ) | ( n6581 & n6582 ) ;
  assign n6584 = ( n6573 & ~n6580 ) | ( n6573 & n6583 ) | ( ~n6580 & n6583 ) ;
  assign n6585 = n6567 & n6584 ;
  assign n6586 = n6565 & n6584 ;
  assign n6587 = ( n4190 & n6585 ) | ( n4190 & n6586 ) | ( n6585 & n6586 ) ;
  assign n6588 = ( n6563 & n6584 ) | ( n6563 & n6587 ) | ( n6584 & n6587 ) ;
  assign n6589 = n6569 & ~n6588 ;
  assign n6590 = ~n6565 & n6584 ;
  assign n6591 = ~n6567 & n6584 ;
  assign n6592 = ( ~n4190 & n6590 ) | ( ~n4190 & n6591 ) | ( n6590 & n6591 ) ;
  assign n6593 = ~n6563 & n6592 ;
  assign n6594 = n6589 | n6593 ;
  assign n6595 = n6329 | n6330 ;
  assign n6596 = n6332 | n6595 ;
  assign n6597 = ( n6323 & n6330 ) | ( n6323 & n6596 ) | ( n6330 & n6596 ) ;
  assign n6598 = n6330 | n6336 ;
  assign n6599 = ( n6149 & n6596 ) | ( n6149 & n6598 ) | ( n6596 & n6598 ) ;
  assign n6600 = ( n5960 & n6597 ) | ( n5960 & n6599 ) | ( n6597 & n6599 ) ;
  assign n6601 = ( n5965 & n6597 ) | ( n5965 & n6599 ) | ( n6597 & n6599 ) ;
  assign n6602 = ( n5962 & n6597 ) | ( n5962 & n6599 ) | ( n6597 & n6599 ) ;
  assign n6603 = ( ~n3952 & n6601 ) | ( ~n3952 & n6602 ) | ( n6601 & n6602 ) ;
  assign n6604 = ( n5947 & n6600 ) | ( n5947 & n6603 ) | ( n6600 & n6603 ) ;
  assign n6605 = n6593 | n6604 ;
  assign n6606 = n6589 | n6605 ;
  assign n6607 = ~n6604 & n6606 ;
  assign n6608 = ( ~n6594 & n6606 ) | ( ~n6594 & n6607 ) | ( n6606 & n6607 ) ;
  assign n6609 = n3259 & n3412 ;
  assign n6610 = ~n3289 & n3414 ;
  assign n6611 = n6609 | n6610 ;
  assign n6612 = n3417 & n4830 ;
  assign n6613 = ( n3423 & n4683 ) | ( n3423 & n4830 ) | ( n4683 & n4830 ) ;
  assign n6614 = n6612 & n6613 ;
  assign n6615 = n6611 | n6614 ;
  assign n6616 = n634 | n6615 ;
  assign n6617 = ( n3431 & n4830 ) | ( n3431 & n5200 ) | ( n4830 & n5200 ) ;
  assign n6618 = n6611 | n6617 ;
  assign n6619 = ( ~n4901 & n6616 ) | ( ~n4901 & n6618 ) | ( n6616 & n6618 ) ;
  assign n6620 = n634 & n6615 ;
  assign n6621 = ( n3424 & n4830 ) | ( n3424 & n5205 ) | ( n4830 & n5205 ) ;
  assign n6622 = ( n634 & n6611 ) | ( n634 & n6621 ) | ( n6611 & n6621 ) ;
  assign n6623 = ( ~n4901 & n6620 ) | ( ~n4901 & n6622 ) | ( n6620 & n6622 ) ;
  assign n6624 = n6619 & ~n6623 ;
  assign n6625 = n6606 & n6624 ;
  assign n6626 = ~n6593 & n6624 ;
  assign n6627 = ~n6589 & n6626 ;
  assign n6628 = ( n6607 & n6625 ) | ( n6607 & n6627 ) | ( n6625 & n6627 ) ;
  assign n6629 = n6608 & ~n6628 ;
  assign n6630 = n6378 | n6395 ;
  assign n6631 = ( n6378 & n6381 ) | ( n6378 & n6630 ) | ( n6381 & n6630 ) ;
  assign n6632 = ~n6606 & n6624 ;
  assign n6633 = n6593 & n6624 ;
  assign n6634 = ( n6589 & n6624 ) | ( n6589 & n6633 ) | ( n6624 & n6633 ) ;
  assign n6635 = ( ~n6607 & n6632 ) | ( ~n6607 & n6634 ) | ( n6632 & n6634 ) ;
  assign n6636 = n6631 & n6635 ;
  assign n6637 = ( n6629 & n6631 ) | ( n6629 & n6636 ) | ( n6631 & n6636 ) ;
  assign n6638 = n6631 | n6635 ;
  assign n6639 = n6629 | n6638 ;
  assign n6640 = ~n6637 & n6639 ;
  assign n6643 = ( n6546 & ~n6640 ) | ( n6546 & n6642 ) | ( ~n6640 & n6642 ) ;
  assign n6644 = ( ~n6546 & n6640 ) | ( ~n6546 & n6642 ) | ( n6640 & n6642 ) ;
  assign n6645 = ( ~n6642 & n6643 ) | ( ~n6642 & n6644 ) | ( n6643 & n6644 ) ;
  assign n6646 = n6437 & n6645 ;
  assign n6647 = ( n6442 & n6645 ) | ( n6442 & n6646 ) | ( n6645 & n6646 ) ;
  assign n6648 = ( n6439 & n6645 ) | ( n6439 & n6646 ) | ( n6645 & n6646 ) ;
  assign n6649 = ( n6236 & n6647 ) | ( n6236 & n6648 ) | ( n6647 & n6648 ) ;
  assign n6650 = ( n6235 & n6647 ) | ( n6235 & n6648 ) | ( n6647 & n6648 ) ;
  assign n6651 = ( n6073 & n6649 ) | ( n6073 & n6650 ) | ( n6649 & n6650 ) ;
  assign n6652 = n6437 | n6645 ;
  assign n6653 = n6442 | n6652 ;
  assign n6654 = n6439 | n6652 ;
  assign n6655 = ( n6236 & n6653 ) | ( n6236 & n6654 ) | ( n6653 & n6654 ) ;
  assign n6656 = ( n6235 & n6653 ) | ( n6235 & n6654 ) | ( n6653 & n6654 ) ;
  assign n6657 = ( n6073 & n6655 ) | ( n6073 & n6656 ) | ( n6655 & n6656 ) ;
  assign n6658 = ~n6651 & n6657 ;
  assign n6659 = n299 | n6460 ;
  assign n6660 = n139 | n525 ;
  assign n6661 = n6243 | n6660 ;
  assign n6662 = n312 | n6661 ;
  assign n6663 = ( ~n2588 & n6659 ) | ( ~n2588 & n6662 ) | ( n6659 & n6662 ) ;
  assign n6664 = n197 | n293 ;
  assign n6665 = n165 | n6664 ;
  assign n6666 = n206 | n822 ;
  assign n6667 = n6665 | n6666 ;
  assign n6668 = n212 | n6667 ;
  assign n6669 = n2587 | n6668 ;
  assign n6670 = n2557 | n6669 ;
  assign n6671 = n6663 | n6670 ;
  assign n6672 = n6658 & n6671 ;
  assign n6673 = n6658 | n6671 ;
  assign n6674 = ~n6672 & n6673 ;
  assign n6675 = n6474 | n6674 ;
  assign n6676 = n6479 | n6675 ;
  assign n6677 = ~n6674 & n6675 ;
  assign n6678 = ( n6479 & ~n6674 ) | ( n6479 & n6677 ) | ( ~n6674 & n6677 ) ;
  assign n6679 = ( ~n6492 & n6676 ) | ( ~n6492 & n6678 ) | ( n6676 & n6678 ) ;
  assign n6680 = n6485 & n6679 ;
  assign n6681 = n6485 | n6679 ;
  assign n6682 = ~n6680 & n6681 ;
  assign n6683 = n6273 | n6487 ;
  assign n6684 = n6274 | n6683 ;
  assign n6685 = n5520 & n6684 ;
  assign n6686 = ~n6682 & n6685 ;
  assign n6687 = n6682 & ~n6685 ;
  assign n6688 = n6686 | n6687 ;
  assign n6689 = n206 | n584 ;
  assign n6690 = n202 | n612 ;
  assign n6691 = n2348 | n6690 ;
  assign n6692 = n6689 | n6691 ;
  assign n6693 = n5010 | n6692 ;
  assign n6694 = n5034 | n6693 ;
  assign n6695 = n279 | n280 ;
  assign n6696 = n2807 | n6695 ;
  assign n6697 = n2729 | n6696 ;
  assign n6698 = n401 | n6697 ;
  assign n6699 = n256 | n428 ;
  assign n6700 = n189 | n233 ;
  assign n6701 = n6699 | n6700 ;
  assign n6702 = n141 | n735 ;
  assign n6703 = n6701 | n6702 ;
  assign n6704 = n6698 | n6703 ;
  assign n6705 = n6694 | n6704 ;
  assign n6706 = n176 | n269 ;
  assign n6707 = n538 | n709 ;
  assign n6708 = n6706 | n6707 ;
  assign n6709 = n718 | n2344 ;
  assign n6710 = n6708 | n6709 ;
  assign n6711 = n6705 | n6710 ;
  assign n6712 = n6546 & n6640 ;
  assign n6713 = n6546 & ~n6712 ;
  assign n6714 = ~n6546 & n6640 ;
  assign n6715 = n6642 & n6714 ;
  assign n6716 = ( n6642 & n6713 ) | ( n6642 & n6715 ) | ( n6713 & n6715 ) ;
  assign n6717 = n6645 | n6716 ;
  assign n6718 = n6437 | n6439 ;
  assign n6719 = ( n6716 & n6717 ) | ( n6716 & n6718 ) | ( n6717 & n6718 ) ;
  assign n6720 = ( n6437 & n6716 ) | ( n6437 & n6717 ) | ( n6716 & n6717 ) ;
  assign n6721 = n6716 | n6717 ;
  assign n6722 = ( n6442 & n6720 ) | ( n6442 & n6721 ) | ( n6720 & n6721 ) ;
  assign n6723 = ( n6236 & n6719 ) | ( n6236 & n6722 ) | ( n6719 & n6722 ) ;
  assign n6724 = n6235 | n6716 ;
  assign n6725 = n6648 | n6716 ;
  assign n6726 = ( n6647 & n6724 ) | ( n6647 & n6725 ) | ( n6724 & n6725 ) ;
  assign n6727 = ( n6073 & n6723 ) | ( n6073 & n6726 ) | ( n6723 & n6726 ) ;
  assign n6728 = n3635 & ~n5080 ;
  assign n6729 = n3637 & n5303 ;
  assign n6730 = n3637 & ~n5075 ;
  assign n6731 = ( ~n3222 & n3637 ) | ( ~n3222 & n6730 ) | ( n3637 & n6730 ) ;
  assign n6732 = ( ~n5304 & n6729 ) | ( ~n5304 & n6731 ) | ( n6729 & n6731 ) ;
  assign n6733 = n6728 | n6732 ;
  assign n6734 = ( n3643 & n3742 ) | ( n3643 & ~n5080 ) | ( n3742 & ~n5080 ) ;
  assign n6735 = n6732 | n6734 ;
  assign n6736 = ( n5546 & n6733 ) | ( n5546 & n6735 ) | ( n6733 & n6735 ) ;
  assign n6737 = ( n482 & n3656 ) | ( n482 & n6728 ) | ( n3656 & n6728 ) ;
  assign n6738 = ( n3713 & n6732 ) | ( n3713 & n6737 ) | ( n6732 & n6737 ) ;
  assign n6739 = n482 & n6728 ;
  assign n6740 = ( n482 & n6732 ) | ( n482 & n6739 ) | ( n6732 & n6739 ) ;
  assign n6741 = ( n5546 & n6738 ) | ( n5546 & n6740 ) | ( n6738 & n6740 ) ;
  assign n6742 = n6736 & ~n6741 ;
  assign n6743 = n3719 & ~n6728 ;
  assign n6744 = ~n6732 & n6743 ;
  assign n6745 = n482 & ~n6728 ;
  assign n6746 = ~n6732 & n6745 ;
  assign n6747 = ( ~n5546 & n6744 ) | ( ~n5546 & n6746 ) | ( n6744 & n6746 ) ;
  assign n6748 = n6742 | n6747 ;
  assign n6749 = n6628 | n6637 ;
  assign n6750 = n6588 | n6604 ;
  assign n6751 = ( n6588 & n6594 ) | ( n6588 & n6750 ) | ( n6594 & n6750 ) ;
  assign n6752 = n6574 & ~n6576 ;
  assign n6753 = ( ~n6570 & n6574 ) | ( ~n6570 & n6752 ) | ( n6574 & n6752 ) ;
  assign n6754 = ( n2921 & n6574 ) | ( n2921 & n6753 ) | ( n6574 & n6753 ) ;
  assign n6755 = ( ~n2828 & n6574 ) | ( ~n2828 & n6754 ) | ( n6574 & n6754 ) ;
  assign n6756 = ~n879 & n6574 ;
  assign n6757 = ( n6574 & ~n6576 ) | ( n6574 & n6756 ) | ( ~n6576 & n6756 ) ;
  assign n6758 = ( ~n2927 & n6755 ) | ( ~n2927 & n6757 ) | ( n6755 & n6757 ) ;
  assign n6759 = n879 & n3024 ;
  assign n6760 = n6758 | n6759 ;
  assign n6761 = ~n6758 & n6760 ;
  assign n6762 = n6758 & ~n6759 ;
  assign n6763 = n6761 | n6762 ;
  assign n6764 = n3259 & n3448 ;
  assign n6765 = n3266 & n3446 ;
  assign n6766 = n3296 & n3477 ;
  assign n6767 = n3295 & n3477 ;
  assign n6768 = ( n2828 & n6766 ) | ( n2828 & n6767 ) | ( n6766 & n6767 ) ;
  assign n6769 = ( ~n3300 & n3477 ) | ( ~n3300 & n6768 ) | ( n3477 & n6768 ) ;
  assign n6770 = n6765 | n6769 ;
  assign n6771 = n6764 | n6770 ;
  assign n6772 = n3452 | n6771 ;
  assign n6773 = n879 & n6771 ;
  assign n6774 = n6772 & n6773 ;
  assign n6775 = ( n879 & n5943 ) | ( n879 & n6771 ) | ( n5943 & n6771 ) ;
  assign n6776 = ( n4532 & n6774 ) | ( n4532 & n6775 ) | ( n6774 & n6775 ) ;
  assign n6777 = n879 | n6771 ;
  assign n6778 = n6182 | n6771 ;
  assign n6779 = ( n4532 & n6777 ) | ( n4532 & n6778 ) | ( n6777 & n6778 ) ;
  assign n6780 = ~n6776 & n6779 ;
  assign n6781 = n6763 & n6780 ;
  assign n6782 = n6763 | n6780 ;
  assign n6783 = ~n6781 & n6782 ;
  assign n6784 = n6750 & n6783 ;
  assign n6785 = n6588 & n6783 ;
  assign n6786 = ( n6594 & n6784 ) | ( n6594 & n6785 ) | ( n6784 & n6785 ) ;
  assign n6787 = n6751 & ~n6786 ;
  assign n6788 = ~n3289 & n3412 ;
  assign n6789 = n3414 & n4830 ;
  assign n6790 = n6788 | n6789 ;
  assign n6791 = n3417 & ~n4854 ;
  assign n6792 = n3285 & n3417 ;
  assign n6793 = n3222 & n6792 ;
  assign n6794 = ( n4855 & n6791 ) | ( n4855 & n6793 ) | ( n6791 & n6793 ) ;
  assign n6795 = n634 & n6794 ;
  assign n6796 = ( n634 & n6790 ) | ( n634 & n6795 ) | ( n6790 & n6795 ) ;
  assign n6797 = n3423 | n6794 ;
  assign n6798 = n634 & n6790 ;
  assign n6799 = ( n634 & n6797 ) | ( n634 & n6798 ) | ( n6797 & n6798 ) ;
  assign n6800 = ( n4869 & n6796 ) | ( n4869 & n6799 ) | ( n6796 & n6799 ) ;
  assign n6801 = n634 | n6794 ;
  assign n6802 = n6790 | n6801 ;
  assign n6803 = n634 | n6790 ;
  assign n6804 = n6797 | n6803 ;
  assign n6805 = ( n4869 & n6802 ) | ( n4869 & n6804 ) | ( n6802 & n6804 ) ;
  assign n6806 = ~n6800 & n6805 ;
  assign n6807 = n6783 | n6806 ;
  assign n6808 = ( ~n6751 & n6806 ) | ( ~n6751 & n6807 ) | ( n6806 & n6807 ) ;
  assign n6809 = n6787 | n6808 ;
  assign n6810 = ~n6750 & n6783 ;
  assign n6811 = ~n6588 & n6783 ;
  assign n6812 = ( ~n6594 & n6810 ) | ( ~n6594 & n6811 ) | ( n6810 & n6811 ) ;
  assign n6813 = n6806 & n6812 ;
  assign n6814 = ( n6787 & n6806 ) | ( n6787 & n6813 ) | ( n6806 & n6813 ) ;
  assign n6815 = n6809 & ~n6814 ;
  assign n6816 = n6749 & n6815 ;
  assign n6817 = n6749 | n6815 ;
  assign n6818 = ~n6816 & n6817 ;
  assign n6819 = n6748 & n6818 ;
  assign n6820 = n6748 | n6818 ;
  assign n6821 = ~n6819 & n6820 ;
  assign n6822 = n6536 | n6640 ;
  assign n6823 = ( n6536 & n6546 ) | ( n6536 & n6822 ) | ( n6546 & n6822 ) ;
  assign n6824 = n6821 & n6823 ;
  assign n6825 = n6821 | n6823 ;
  assign n6826 = ~n6824 & n6825 ;
  assign n6827 = n6726 & n6826 ;
  assign n6828 = n6722 & n6826 ;
  assign n6829 = n6719 & n6826 ;
  assign n6830 = ( n6236 & n6828 ) | ( n6236 & n6829 ) | ( n6828 & n6829 ) ;
  assign n6831 = ( n6073 & n6827 ) | ( n6073 & n6830 ) | ( n6827 & n6830 ) ;
  assign n6832 = n6826 & ~n6830 ;
  assign n6833 = ~n6726 & n6826 ;
  assign n6834 = ( ~n6073 & n6832 ) | ( ~n6073 & n6833 ) | ( n6832 & n6833 ) ;
  assign n6835 = ( n6727 & ~n6831 ) | ( n6727 & n6834 ) | ( ~n6831 & n6834 ) ;
  assign n6836 = n6711 | n6835 ;
  assign n6837 = n6711 & n6835 ;
  assign n6838 = n6836 & ~n6837 ;
  assign n6839 = n6474 | n6672 ;
  assign n6840 = ( n6672 & n6674 ) | ( n6672 & n6839 ) | ( n6674 & n6839 ) ;
  assign n6841 = n6838 & n6840 ;
  assign n6842 = n6672 | n6674 ;
  assign n6843 = n6838 & n6842 ;
  assign n6844 = ( n6479 & n6841 ) | ( n6479 & n6843 ) | ( n6841 & n6843 ) ;
  assign n6845 = n6838 | n6840 ;
  assign n6846 = n6838 | n6842 ;
  assign n6847 = ( n6479 & n6845 ) | ( n6479 & n6846 ) | ( n6845 & n6846 ) ;
  assign n6848 = ~n6844 & n6847 ;
  assign n6849 = n6679 & n6848 ;
  assign n6850 = n6485 & n6849 ;
  assign n6851 = n6679 | n6848 ;
  assign n6852 = ( n6485 & n6848 ) | ( n6485 & n6851 ) | ( n6848 & n6851 ) ;
  assign n6853 = ~n6850 & n6852 ;
  assign n6854 = n6682 | n6684 ;
  assign n6855 = n5520 & n6854 ;
  assign n6856 = ~n6853 & n6855 ;
  assign n6857 = n6853 & ~n6855 ;
  assign n6858 = n6856 | n6857 ;
  assign n6859 = n3643 & ~n5315 ;
  assign n6860 = n3643 & n5303 ;
  assign n6861 = n3643 & ~n5075 ;
  assign n6862 = ( ~n3222 & n3643 ) | ( ~n3222 & n6861 ) | ( n3643 & n6861 ) ;
  assign n6863 = ( ~n5304 & n6860 ) | ( ~n5304 & n6862 ) | ( n6860 & n6862 ) ;
  assign n6864 = ( n5316 & n6859 ) | ( n5316 & n6863 ) | ( n6859 & n6863 ) ;
  assign n6865 = n3635 & n5303 ;
  assign n6866 = n3635 & ~n5075 ;
  assign n6867 = ( ~n3222 & n3635 ) | ( ~n3222 & n6866 ) | ( n3635 & n6866 ) ;
  assign n6868 = ( ~n5304 & n6865 ) | ( ~n5304 & n6867 ) | ( n6865 & n6867 ) ;
  assign n6869 = n6864 | n6868 ;
  assign n6870 = n6863 | n6868 ;
  assign n6871 = ( ~n5534 & n6868 ) | ( ~n5534 & n6870 ) | ( n6868 & n6870 ) ;
  assign n6872 = ( n5093 & n6869 ) | ( n5093 & n6871 ) | ( n6869 & n6871 ) ;
  assign n6873 = ( n5090 & n6869 ) | ( n5090 & n6871 ) | ( n6869 & n6871 ) ;
  assign n6874 = ( n4841 & n6872 ) | ( n4841 & n6873 ) | ( n6872 & n6873 ) ;
  assign n6875 = n482 & ~n6874 ;
  assign n6876 = ~n482 & n6874 ;
  assign n6877 = n6875 | n6876 ;
  assign n6878 = n6786 & n6877 ;
  assign n6879 = ( n6814 & n6877 ) | ( n6814 & n6878 ) | ( n6877 & n6878 ) ;
  assign n6880 = n6786 | n6877 ;
  assign n6881 = n6814 | n6880 ;
  assign n6882 = ~n6879 & n6881 ;
  assign n6883 = ~n3289 & n3448 ;
  assign n6884 = n3266 & n3477 ;
  assign n6885 = n3259 & n3446 ;
  assign n6886 = n6884 | n6885 ;
  assign n6887 = n6883 | n6886 ;
  assign n6888 = ( ~n3289 & n3452 ) | ( ~n3289 & n5365 ) | ( n3452 & n5365 ) ;
  assign n6889 = n6886 | n6888 ;
  assign n6890 = ( ~n3321 & n6887 ) | ( ~n3321 & n6889 ) | ( n6887 & n6889 ) ;
  assign n6891 = ~n3289 & n5369 ;
  assign n6892 = ( n879 & n6886 ) | ( n879 & n6891 ) | ( n6886 & n6891 ) ;
  assign n6893 = n879 & n6888 ;
  assign n6894 = ( n879 & n6886 ) | ( n879 & n6893 ) | ( n6886 & n6893 ) ;
  assign n6895 = ( ~n3321 & n6892 ) | ( ~n3321 & n6894 ) | ( n6892 & n6894 ) ;
  assign n6896 = n6890 & ~n6895 ;
  assign n6897 = n879 & ~n6891 ;
  assign n6898 = ~n6886 & n6897 ;
  assign n6899 = n879 & ~n6888 ;
  assign n6900 = ~n6886 & n6899 ;
  assign n6901 = ( n3321 & n6898 ) | ( n3321 & n6900 ) | ( n6898 & n6900 ) ;
  assign n6902 = n6896 | n6901 ;
  assign n6903 = n879 & ~n3305 ;
  assign n6904 = n6900 & ~n6903 ;
  assign n6905 = n6898 & ~n6903 ;
  assign n6906 = ( n3321 & n6904 ) | ( n3321 & n6905 ) | ( n6904 & n6905 ) ;
  assign n6907 = ( n6896 & ~n6903 ) | ( n6896 & n6906 ) | ( ~n6903 & n6906 ) ;
  assign n6908 = n6902 & ~n6907 ;
  assign n6909 = n6898 | n6903 ;
  assign n6910 = n6900 | n6903 ;
  assign n6911 = ( n3321 & n6909 ) | ( n3321 & n6910 ) | ( n6909 & n6910 ) ;
  assign n6912 = n6896 | n6911 ;
  assign n6913 = ( n6758 & n6759 ) | ( n6758 & ~n6780 ) | ( n6759 & ~n6780 ) ;
  assign n6914 = n6912 & ~n6913 ;
  assign n6915 = ~n6908 & n6914 ;
  assign n6916 = ~n6912 & n6913 ;
  assign n6917 = ( n6908 & n6913 ) | ( n6908 & n6916 ) | ( n6913 & n6916 ) ;
  assign n6918 = n6915 | n6917 ;
  assign n6919 = n3414 & ~n4854 ;
  assign n6920 = n3285 & n3414 ;
  assign n6921 = n3222 & n6920 ;
  assign n6922 = ( n4855 & n6919 ) | ( n4855 & n6921 ) | ( n6919 & n6921 ) ;
  assign n6923 = n3412 & n4830 ;
  assign n6924 = ( n3423 & n4683 ) | ( n3423 & ~n5080 ) | ( n4683 & ~n5080 ) ;
  assign n6925 = n6923 | n6924 ;
  assign n6926 = n6922 | n6925 ;
  assign n6927 = n634 & n6926 ;
  assign n6928 = n4687 & ~n5080 ;
  assign n6929 = ( n634 & n6923 ) | ( n634 & n6928 ) | ( n6923 & n6928 ) ;
  assign n6930 = n634 | n4687 ;
  assign n6931 = ( n634 & ~n5080 ) | ( n634 & n6930 ) | ( ~n5080 & n6930 ) ;
  assign n6932 = ( n6922 & n6929 ) | ( n6922 & n6931 ) | ( n6929 & n6931 ) ;
  assign n6933 = ( ~n5099 & n6927 ) | ( ~n5099 & n6932 ) | ( n6927 & n6932 ) ;
  assign n6934 = n634 | n6926 ;
  assign n6935 = ( n634 & n4692 ) | ( n634 & ~n5080 ) | ( n4692 & ~n5080 ) ;
  assign n6936 = n6923 | n6935 ;
  assign n6937 = n6922 | n6936 ;
  assign n6938 = ( ~n5099 & n6934 ) | ( ~n5099 & n6937 ) | ( n6934 & n6937 ) ;
  assign n6939 = ~n6933 & n6938 ;
  assign n6940 = ~n6918 & n6939 ;
  assign n6941 = n6918 & ~n6939 ;
  assign n6942 = n6940 | n6941 ;
  assign n6943 = n6882 & ~n6942 ;
  assign n6944 = n6882 | n6942 ;
  assign n6945 = ( ~n6882 & n6943 ) | ( ~n6882 & n6944 ) | ( n6943 & n6944 ) ;
  assign n6946 = ( n6748 & n6749 ) | ( n6748 & n6815 ) | ( n6749 & n6815 ) ;
  assign n6947 = ~n6945 & n6946 ;
  assign n6948 = n6945 & ~n6946 ;
  assign n6949 = n6947 | n6948 ;
  assign n6950 = n6824 & n6949 ;
  assign n6951 = ( n6826 & n6949 ) | ( n6826 & n6950 ) | ( n6949 & n6950 ) ;
  assign n6952 = ( n6722 & n6950 ) | ( n6722 & n6951 ) | ( n6950 & n6951 ) ;
  assign n6953 = ( n6719 & n6950 ) | ( n6719 & n6951 ) | ( n6950 & n6951 ) ;
  assign n6954 = ( n6236 & n6952 ) | ( n6236 & n6953 ) | ( n6952 & n6953 ) ;
  assign n6955 = ( n6716 & n6950 ) | ( n6716 & n6951 ) | ( n6950 & n6951 ) ;
  assign n6956 = n6950 | n6951 ;
  assign n6957 = ( n6235 & n6955 ) | ( n6235 & n6956 ) | ( n6955 & n6956 ) ;
  assign n6958 = ( n6648 & n6955 ) | ( n6648 & n6956 ) | ( n6955 & n6956 ) ;
  assign n6959 = ( n6647 & n6957 ) | ( n6647 & n6958 ) | ( n6957 & n6958 ) ;
  assign n6960 = ( n6073 & n6954 ) | ( n6073 & n6959 ) | ( n6954 & n6959 ) ;
  assign n6961 = n6824 | n6949 ;
  assign n6962 = n6826 | n6961 ;
  assign n6963 = ( n6722 & n6961 ) | ( n6722 & n6962 ) | ( n6961 & n6962 ) ;
  assign n6964 = ( n6719 & n6961 ) | ( n6719 & n6962 ) | ( n6961 & n6962 ) ;
  assign n6965 = ( n6236 & n6963 ) | ( n6236 & n6964 ) | ( n6963 & n6964 ) ;
  assign n6966 = ( n6716 & n6961 ) | ( n6716 & n6962 ) | ( n6961 & n6962 ) ;
  assign n6967 = n6961 | n6962 ;
  assign n6968 = ( n6235 & n6966 ) | ( n6235 & n6967 ) | ( n6966 & n6967 ) ;
  assign n6969 = ( n6648 & n6966 ) | ( n6648 & n6967 ) | ( n6966 & n6967 ) ;
  assign n6970 = ( n6647 & n6968 ) | ( n6647 & n6969 ) | ( n6968 & n6969 ) ;
  assign n6971 = ( n6073 & n6965 ) | ( n6073 & n6970 ) | ( n6965 & n6970 ) ;
  assign n6972 = ~n6960 & n6971 ;
  assign n6973 = n361 | n2746 ;
  assign n6974 = n261 | n3241 ;
  assign n6975 = n168 | n312 ;
  assign n6976 = n163 | n6975 ;
  assign n6977 = n6974 | n6976 ;
  assign n6978 = n4822 | n6977 ;
  assign n6979 = n4931 | n6978 ;
  assign n6980 = n6973 | n6979 ;
  assign n6981 = n216 | n524 ;
  assign n6982 = n189 | n266 ;
  assign n6983 = n6981 | n6982 ;
  assign n6984 = n280 | n435 ;
  assign n6985 = n235 | n6984 ;
  assign n6986 = n6983 | n6985 ;
  assign n6987 = n6980 | n6986 ;
  assign n6988 = n6972 | n6987 ;
  assign n6989 = n6972 & n6987 ;
  assign n6990 = n6988 & ~n6989 ;
  assign n6991 = n6837 & n6990 ;
  assign n6992 = ( n6843 & n6990 ) | ( n6843 & n6991 ) | ( n6990 & n6991 ) ;
  assign n6993 = ( n6841 & n6990 ) | ( n6841 & n6991 ) | ( n6990 & n6991 ) ;
  assign n6994 = ( n6479 & n6992 ) | ( n6479 & n6993 ) | ( n6992 & n6993 ) ;
  assign n6995 = n6837 | n6990 ;
  assign n6996 = n6843 | n6995 ;
  assign n6997 = n6841 | n6995 ;
  assign n6998 = ( n6479 & n6996 ) | ( n6479 & n6997 ) | ( n6996 & n6997 ) ;
  assign n6999 = ~n6994 & n6998 ;
  assign n7000 = n6850 | n6999 ;
  assign n7001 = n6850 & n6999 ;
  assign n7002 = n7000 & ~n7001 ;
  assign n7003 = n6682 | n6853 ;
  assign n7004 = n6684 | n7003 ;
  assign n7005 = n5520 & n7004 ;
  assign n7006 = ~n7002 & n7005 ;
  assign n7007 = n7002 & ~n7005 ;
  assign n7008 = n7006 | n7007 ;
  assign n7035 = ( n6912 & n6913 ) | ( n6912 & ~n6939 ) | ( n6913 & ~n6939 ) ;
  assign n7036 = n6913 & ~n6939 ;
  assign n7037 = ( ~n6908 & n7035 ) | ( ~n6908 & n7036 ) | ( n7035 & n7036 ) ;
  assign n7009 = n3414 & ~n5080 ;
  assign n7010 = n3412 & ~n4854 ;
  assign n7011 = n3285 & n3412 ;
  assign n7012 = n3222 & n7011 ;
  assign n7013 = ( n4855 & n7010 ) | ( n4855 & n7012 ) | ( n7010 & n7012 ) ;
  assign n7014 = n7009 | n7013 ;
  assign n7015 = n3417 & n5303 ;
  assign n7016 = n3417 & ~n5075 ;
  assign n7017 = ( ~n3222 & n3417 ) | ( ~n3222 & n7016 ) | ( n3417 & n7016 ) ;
  assign n7018 = ( ~n5304 & n7015 ) | ( ~n5304 & n7017 ) | ( n7015 & n7017 ) ;
  assign n7019 = ( n3423 & n4683 ) | ( n3423 & n5303 ) | ( n4683 & n5303 ) ;
  assign n7020 = ( n3423 & n4683 ) | ( n3423 & ~n5075 ) | ( n4683 & ~n5075 ) ;
  assign n7021 = n3423 | n4683 ;
  assign n7022 = ( ~n3222 & n7020 ) | ( ~n3222 & n7021 ) | ( n7020 & n7021 ) ;
  assign n7023 = ( ~n5304 & n7019 ) | ( ~n5304 & n7022 ) | ( n7019 & n7022 ) ;
  assign n7024 = n7018 & n7023 ;
  assign n7025 = n7014 | n7024 ;
  assign n7026 = n634 | n7025 ;
  assign n7027 = n634 | n7023 ;
  assign n7028 = n7014 | n7027 ;
  assign n7029 = ( n5325 & n7026 ) | ( n5325 & n7028 ) | ( n7026 & n7028 ) ;
  assign n7030 = n634 & n7025 ;
  assign n7031 = n634 & n7023 ;
  assign n7032 = ( n634 & n7014 ) | ( n634 & n7031 ) | ( n7014 & n7031 ) ;
  assign n7033 = ( n5325 & n7030 ) | ( n5325 & n7032 ) | ( n7030 & n7032 ) ;
  assign n7034 = n7029 & ~n7033 ;
  assign n7038 = n7034 & ~n7037 ;
  assign n7039 = n7037 | n7038 ;
  assign n7040 = n7034 & n7037 ;
  assign n7041 = n3448 & n4830 ;
  assign n7042 = n3259 & n3477 ;
  assign n7043 = ~n3289 & n3446 ;
  assign n7044 = n7042 | n7043 ;
  assign n7045 = n7041 | n7044 ;
  assign n7046 = ( n3452 & n4830 ) | ( n3452 & n5365 ) | ( n4830 & n5365 ) ;
  assign n7047 = n7044 | n7046 ;
  assign n7048 = ( ~n4901 & n7045 ) | ( ~n4901 & n7047 ) | ( n7045 & n7047 ) ;
  assign n7049 = n4830 & n5369 ;
  assign n7050 = ( n879 & n7044 ) | ( n879 & n7049 ) | ( n7044 & n7049 ) ;
  assign n7051 = n879 & n7046 ;
  assign n7052 = ( n879 & n7044 ) | ( n879 & n7051 ) | ( n7044 & n7051 ) ;
  assign n7053 = ( ~n4901 & n7050 ) | ( ~n4901 & n7052 ) | ( n7050 & n7052 ) ;
  assign n7054 = n7048 & ~n7053 ;
  assign n7055 = n879 & ~n7049 ;
  assign n7056 = ~n7044 & n7055 ;
  assign n7057 = n879 & ~n7046 ;
  assign n7058 = ~n7044 & n7057 ;
  assign n7059 = ( n4901 & n7056 ) | ( n4901 & n7058 ) | ( n7056 & n7058 ) ;
  assign n7060 = n7054 | n7059 ;
  assign n7061 = n482 & ~n879 ;
  assign n7062 = ( n482 & ~n3266 ) | ( n482 & n7061 ) | ( ~n3266 & n7061 ) ;
  assign n7063 = ~n482 & n879 ;
  assign n7064 = n3266 & n7063 ;
  assign n7065 = n6759 & ~n7064 ;
  assign n7066 = n7062 & ~n7064 ;
  assign n7067 = ( n7064 & n7065 ) | ( n7064 & ~n7066 ) | ( n7065 & ~n7066 ) ;
  assign n7068 = n7062 | n7067 ;
  assign n7069 = n6759 & n7062 ;
  assign n7070 = ( n6759 & ~n7065 ) | ( n6759 & n7069 ) | ( ~n7065 & n7069 ) ;
  assign n7071 = n7068 & ~n7070 ;
  assign n7072 = n879 & ~n3024 ;
  assign n7073 = ~n3301 & n7072 ;
  assign n7074 = n7070 & n7073 ;
  assign n7075 = ( ~n7068 & n7073 ) | ( ~n7068 & n7074 ) | ( n7073 & n7074 ) ;
  assign n7076 = ( n6903 & n7071 ) | ( n6903 & ~n7075 ) | ( n7071 & ~n7075 ) ;
  assign n7077 = ( n6905 & ~n7071 ) | ( n6905 & n7075 ) | ( ~n7071 & n7075 ) ;
  assign n7078 = ( n6904 & ~n7071 ) | ( n6904 & n7075 ) | ( ~n7071 & n7075 ) ;
  assign n7079 = ( n3321 & n7077 ) | ( n3321 & n7078 ) | ( n7077 & n7078 ) ;
  assign n7080 = ( n6896 & ~n7076 ) | ( n6896 & n7079 ) | ( ~n7076 & n7079 ) ;
  assign n7081 = n6903 & ~n7073 ;
  assign n7082 = n6905 | n7073 ;
  assign n7083 = n6904 | n7073 ;
  assign n7084 = ( n3321 & n7082 ) | ( n3321 & n7083 ) | ( n7082 & n7083 ) ;
  assign n7085 = ( n6896 & ~n7081 ) | ( n6896 & n7084 ) | ( ~n7081 & n7084 ) ;
  assign n7086 = ~n7080 & n7085 ;
  assign n7087 = n7071 | n7075 ;
  assign n7088 = n6903 & ~n7087 ;
  assign n7089 = n6905 | n7087 ;
  assign n7090 = n6904 | n7087 ;
  assign n7091 = ( n3321 & n7089 ) | ( n3321 & n7090 ) | ( n7089 & n7090 ) ;
  assign n7092 = ( n6896 & ~n7088 ) | ( n6896 & n7091 ) | ( ~n7088 & n7091 ) ;
  assign n7093 = n7060 & ~n7092 ;
  assign n7094 = ( n7060 & n7086 ) | ( n7060 & n7093 ) | ( n7086 & n7093 ) ;
  assign n7095 = ~n7086 & n7092 ;
  assign n7096 = n7060 | n7095 ;
  assign n7097 = ( ~n7060 & n7094 ) | ( ~n7060 & n7096 ) | ( n7094 & n7096 ) ;
  assign n7098 = ~n7040 & n7097 ;
  assign n7099 = n7039 & n7098 ;
  assign n7100 = n7040 & ~n7097 ;
  assign n7101 = ( n7039 & n7097 ) | ( n7039 & ~n7100 ) | ( n7097 & ~n7100 ) ;
  assign n7102 = ~n7099 & n7101 ;
  assign n7103 = n6879 | n6942 ;
  assign n7104 = ( n6879 & n6882 ) | ( n6879 & n7103 ) | ( n6882 & n7103 ) ;
  assign n7105 = n7102 & n7104 ;
  assign n7106 = n7102 | n7104 ;
  assign n7107 = ~n7105 & n7106 ;
  assign n7108 = n6945 & n6946 ;
  assign n7109 = n7107 & n7108 ;
  assign n7110 = ( n6951 & n7107 ) | ( n6951 & n7109 ) | ( n7107 & n7109 ) ;
  assign n7111 = ( n6949 & n7107 ) | ( n6949 & n7109 ) | ( n7107 & n7109 ) ;
  assign n7112 = n7107 & n7109 ;
  assign n7113 = ( n6824 & n7111 ) | ( n6824 & n7112 ) | ( n7111 & n7112 ) ;
  assign n7114 = ( n6722 & n7110 ) | ( n6722 & n7113 ) | ( n7110 & n7113 ) ;
  assign n7115 = ( n6719 & n7110 ) | ( n6719 & n7113 ) | ( n7110 & n7113 ) ;
  assign n7116 = ( n6236 & n7114 ) | ( n6236 & n7115 ) | ( n7114 & n7115 ) ;
  assign n7117 = ( n6716 & n7109 ) | ( n6716 & n7113 ) | ( n7109 & n7113 ) ;
  assign n7118 = ( n6716 & n7107 ) | ( n6716 & n7113 ) | ( n7107 & n7113 ) ;
  assign n7119 = ( n6951 & n7117 ) | ( n6951 & n7118 ) | ( n7117 & n7118 ) ;
  assign n7120 = n7109 | n7113 ;
  assign n7121 = n7107 | n7113 ;
  assign n7122 = ( n6951 & n7120 ) | ( n6951 & n7121 ) | ( n7120 & n7121 ) ;
  assign n7123 = ( n6235 & n7119 ) | ( n6235 & n7122 ) | ( n7119 & n7122 ) ;
  assign n7124 = ( n6648 & n7119 ) | ( n6648 & n7122 ) | ( n7119 & n7122 ) ;
  assign n7125 = ( n6647 & n7123 ) | ( n6647 & n7124 ) | ( n7123 & n7124 ) ;
  assign n7126 = ( n6073 & n7116 ) | ( n6073 & n7125 ) | ( n7116 & n7125 ) ;
  assign n7127 = n7107 | n7108 ;
  assign n7128 = n6951 | n7127 ;
  assign n7129 = n6949 | n7127 ;
  assign n7130 = ( n6824 & n7127 ) | ( n6824 & n7129 ) | ( n7127 & n7129 ) ;
  assign n7131 = ( n6722 & n7128 ) | ( n6722 & n7130 ) | ( n7128 & n7130 ) ;
  assign n7132 = ( n6719 & n7128 ) | ( n6719 & n7130 ) | ( n7128 & n7130 ) ;
  assign n7133 = ( n6236 & n7131 ) | ( n6236 & n7132 ) | ( n7131 & n7132 ) ;
  assign n7134 = ( n6716 & n7127 ) | ( n6716 & n7130 ) | ( n7127 & n7130 ) ;
  assign n7135 = n6716 | n7130 ;
  assign n7136 = ( n6951 & n7134 ) | ( n6951 & n7135 ) | ( n7134 & n7135 ) ;
  assign n7137 = n7127 | n7130 ;
  assign n7138 = n6951 | n7137 ;
  assign n7139 = ( n6235 & n7136 ) | ( n6235 & n7138 ) | ( n7136 & n7138 ) ;
  assign n7140 = ( n6648 & n7136 ) | ( n6648 & n7138 ) | ( n7136 & n7138 ) ;
  assign n7141 = ( n6647 & n7139 ) | ( n6647 & n7140 ) | ( n7139 & n7140 ) ;
  assign n7142 = ( n6073 & n7133 ) | ( n6073 & n7141 ) | ( n7133 & n7141 ) ;
  assign n7143 = ~n7126 & n7142 ;
  assign n7144 = n311 | n3175 ;
  assign n7145 = n231 | n7144 ;
  assign n7146 = n296 | n7145 ;
  assign n7147 = n688 | n7146 ;
  assign n7148 = n4944 | n5023 ;
  assign n7149 = n7147 | n7148 ;
  assign n7150 = n823 | n4822 ;
  assign n7151 = n821 | n7150 ;
  assign n7152 = n812 | n7151 ;
  assign n7153 = n7149 | n7152 ;
  assign n7154 = n452 | n545 ;
  assign n7155 = n582 | n7154 ;
  assign n7156 = n200 | n443 ;
  assign n7157 = n7155 | n7156 ;
  assign n7158 = n7153 | n7157 ;
  assign n7159 = n7143 | n7158 ;
  assign n7160 = n7143 & n7158 ;
  assign n7161 = n7159 & ~n7160 ;
  assign n7162 = n6837 | n6989 ;
  assign n7163 = ( n6989 & n6990 ) | ( n6989 & n7162 ) | ( n6990 & n7162 ) ;
  assign n7164 = n7161 & n7163 ;
  assign n7165 = n6989 | n6990 ;
  assign n7166 = n7161 & n7165 ;
  assign n7167 = ( n6843 & n7164 ) | ( n6843 & n7166 ) | ( n7164 & n7166 ) ;
  assign n7168 = ( n6841 & n7164 ) | ( n6841 & n7166 ) | ( n7164 & n7166 ) ;
  assign n7169 = ( n6479 & n7167 ) | ( n6479 & n7168 ) | ( n7167 & n7168 ) ;
  assign n7170 = n7161 | n7163 ;
  assign n7171 = n7161 | n7165 ;
  assign n7172 = ( n6843 & n7170 ) | ( n6843 & n7171 ) | ( n7170 & n7171 ) ;
  assign n7173 = ( n6841 & n7170 ) | ( n6841 & n7171 ) | ( n7170 & n7171 ) ;
  assign n7174 = ( n6479 & n7172 ) | ( n6479 & n7173 ) | ( n7172 & n7173 ) ;
  assign n7175 = ~n7169 & n7174 ;
  assign n7176 = n6999 & n7175 ;
  assign n7177 = n6850 & n7176 ;
  assign n7178 = n6999 | n7175 ;
  assign n7179 = ( n6850 & n7175 ) | ( n6850 & n7178 ) | ( n7175 & n7178 ) ;
  assign n7180 = ~n7177 & n7179 ;
  assign n7181 = n7002 | n7004 ;
  assign n7182 = n5520 & n7181 ;
  assign n7183 = ~n7180 & n7182 ;
  assign n7184 = n7180 & ~n7182 ;
  assign n7185 = n7183 | n7184 ;
  assign n7186 = n7002 | n7180 ;
  assign n7187 = n7004 | n7186 ;
  assign n7188 = n5520 & n7187 ;
  assign n7189 = n7160 | n7169 ;
  assign n7190 = n200 | n1031 ;
  assign n7191 = n554 | n575 ;
  assign n7192 = n7190 | n7191 ;
  assign n7193 = n5060 | n7192 ;
  assign n7194 = n704 | n732 ;
  assign n7195 = n7193 | n7194 ;
  assign n7196 = n682 | n7195 ;
  assign n7197 = n320 | n7196 ;
  assign n7198 = n879 & n3259 ;
  assign n7199 = n7067 & n7198 ;
  assign n7200 = n7067 | n7198 ;
  assign n7201 = ~n7199 & n7200 ;
  assign n7202 = ~n3289 & n3477 ;
  assign n7203 = n3446 & n4830 ;
  assign n7204 = n7202 | n7203 ;
  assign n7205 = ( n3452 & ~n4854 ) | ( n3452 & n5365 ) | ( ~n4854 & n5365 ) ;
  assign n7206 = ( n3285 & n3452 ) | ( n3285 & n5365 ) | ( n3452 & n5365 ) ;
  assign n7207 = n3452 & n5365 ;
  assign n7208 = ( n3222 & n7206 ) | ( n3222 & n7207 ) | ( n7206 & n7207 ) ;
  assign n7209 = ( n4855 & n7205 ) | ( n4855 & n7208 ) | ( n7205 & n7208 ) ;
  assign n7210 = n7204 | n7209 ;
  assign n7211 = n879 | n7210 ;
  assign n7212 = n3448 & ~n4854 ;
  assign n7213 = n3285 & n3448 ;
  assign n7214 = n3222 & n7213 ;
  assign n7215 = ( n4855 & n7212 ) | ( n4855 & n7214 ) | ( n7212 & n7214 ) ;
  assign n7216 = n7209 & n7215 ;
  assign n7217 = n879 | n7204 ;
  assign n7218 = n7216 | n7217 ;
  assign n7219 = ( n4869 & n7211 ) | ( n4869 & n7218 ) | ( n7211 & n7218 ) ;
  assign n7220 = n879 & n7210 ;
  assign n7221 = n879 & n7204 ;
  assign n7222 = ( n879 & n7216 ) | ( n879 & n7221 ) | ( n7216 & n7221 ) ;
  assign n7223 = ( n4869 & n7220 ) | ( n4869 & n7222 ) | ( n7220 & n7222 ) ;
  assign n7224 = n7219 & ~n7223 ;
  assign n7225 = ~n7201 & n7224 ;
  assign n7226 = n7201 & ~n7224 ;
  assign n7227 = n7225 | n7226 ;
  assign n7228 = n7080 & ~n7227 ;
  assign n7229 = ( n7094 & ~n7227 ) | ( n7094 & n7228 ) | ( ~n7227 & n7228 ) ;
  assign n7230 = n7080 | n7086 ;
  assign n7231 = n7060 | n7080 ;
  assign n7232 = ( n7093 & n7230 ) | ( n7093 & n7231 ) | ( n7230 & n7231 ) ;
  assign n7233 = ~n7229 & n7232 ;
  assign n7234 = n7227 | n7229 ;
  assign n7235 = ~n7233 & n7234 ;
  assign n7236 = n3414 & n5303 ;
  assign n7237 = n3414 & ~n5075 ;
  assign n7238 = ( ~n3222 & n3414 ) | ( ~n3222 & n7237 ) | ( n3414 & n7237 ) ;
  assign n7239 = ( ~n5304 & n7236 ) | ( ~n5304 & n7238 ) | ( n7236 & n7238 ) ;
  assign n7240 = n3412 & ~n5080 ;
  assign n7241 = ( n634 & n3424 ) | ( n634 & n7240 ) | ( n3424 & n7240 ) ;
  assign n7242 = ( n3426 & n7239 ) | ( n3426 & n7241 ) | ( n7239 & n7241 ) ;
  assign n7243 = n634 & n7240 ;
  assign n7244 = ( n634 & n7239 ) | ( n634 & n7243 ) | ( n7239 & n7243 ) ;
  assign n7245 = ( n5546 & n7242 ) | ( n5546 & n7244 ) | ( n7242 & n7244 ) ;
  assign n7246 = n3431 | n7240 ;
  assign n7247 = n7239 | n7246 ;
  assign n7248 = n634 | n7240 ;
  assign n7249 = n7239 | n7248 ;
  assign n7250 = ( n5546 & n7247 ) | ( n5546 & n7249 ) | ( n7247 & n7249 ) ;
  assign n7251 = ~n7245 & n7250 ;
  assign n7252 = ~n7235 & n7251 ;
  assign n7253 = n7227 & ~n7251 ;
  assign n7254 = ( n7229 & ~n7251 ) | ( n7229 & n7253 ) | ( ~n7251 & n7253 ) ;
  assign n7255 = ~n7233 & n7254 ;
  assign n7256 = ~n7038 & n7097 ;
  assign n7257 = ~n7038 & n7039 ;
  assign n7258 = ( ~n7100 & n7256 ) | ( ~n7100 & n7257 ) | ( n7256 & n7257 ) ;
  assign n7259 = n7255 | n7258 ;
  assign n7260 = n7252 | n7259 ;
  assign n7261 = n7255 & n7258 ;
  assign n7262 = ( n7252 & n7258 ) | ( n7252 & n7261 ) | ( n7258 & n7261 ) ;
  assign n7263 = n7260 & ~n7262 ;
  assign n7264 = n7105 & n7263 ;
  assign n7265 = ( n7109 & n7263 ) | ( n7109 & n7264 ) | ( n7263 & n7264 ) ;
  assign n7266 = ( n7107 & n7263 ) | ( n7107 & n7264 ) | ( n7263 & n7264 ) ;
  assign n7267 = ( n6950 & n7265 ) | ( n6950 & n7266 ) | ( n7265 & n7266 ) ;
  assign n7268 = ( n6951 & n7265 ) | ( n6951 & n7266 ) | ( n7265 & n7266 ) ;
  assign n7269 = ( n6716 & n7267 ) | ( n6716 & n7268 ) | ( n7267 & n7268 ) ;
  assign n7270 = n7267 | n7268 ;
  assign n7271 = ( n6650 & n7269 ) | ( n6650 & n7270 ) | ( n7269 & n7270 ) ;
  assign n7272 = ( n6722 & n7267 ) | ( n6722 & n7268 ) | ( n7267 & n7268 ) ;
  assign n7273 = ( n6719 & n7267 ) | ( n6719 & n7268 ) | ( n7267 & n7268 ) ;
  assign n7274 = ( n6236 & n7272 ) | ( n6236 & n7273 ) | ( n7272 & n7273 ) ;
  assign n7275 = ( n6073 & n7271 ) | ( n6073 & n7274 ) | ( n7271 & n7274 ) ;
  assign n7276 = n7105 | n7263 ;
  assign n7277 = n7109 | n7276 ;
  assign n7278 = n7107 | n7276 ;
  assign n7279 = ( n6950 & n7277 ) | ( n6950 & n7278 ) | ( n7277 & n7278 ) ;
  assign n7280 = ( n6951 & n7277 ) | ( n6951 & n7278 ) | ( n7277 & n7278 ) ;
  assign n7281 = ( n6716 & n7279 ) | ( n6716 & n7280 ) | ( n7279 & n7280 ) ;
  assign n7282 = n7279 | n7280 ;
  assign n7283 = ( n6650 & n7281 ) | ( n6650 & n7282 ) | ( n7281 & n7282 ) ;
  assign n7284 = ( n6722 & n7279 ) | ( n6722 & n7280 ) | ( n7279 & n7280 ) ;
  assign n7285 = ( n6719 & n7279 ) | ( n6719 & n7280 ) | ( n7279 & n7280 ) ;
  assign n7286 = ( n6236 & n7284 ) | ( n6236 & n7285 ) | ( n7284 & n7285 ) ;
  assign n7287 = ( n6073 & n7283 ) | ( n6073 & n7286 ) | ( n7283 & n7286 ) ;
  assign n7288 = ~n7275 & n7287 ;
  assign n7289 = n7197 | n7288 ;
  assign n7290 = n7197 & n7288 ;
  assign n7291 = n7289 & ~n7290 ;
  assign n7292 = n7160 | n7291 ;
  assign n7293 = n7169 | n7292 ;
  assign n7294 = ~n7291 & n7292 ;
  assign n7295 = ( n7169 & ~n7291 ) | ( n7169 & n7294 ) | ( ~n7291 & n7294 ) ;
  assign n7296 = ( ~n7189 & n7293 ) | ( ~n7189 & n7295 ) | ( n7293 & n7295 ) ;
  assign n7297 = n7176 & ~n7296 ;
  assign n7298 = n6850 & n7297 ;
  assign n7299 = n7296 | n7298 ;
  assign n7300 = ( ~n7177 & n7298 ) | ( ~n7177 & n7299 ) | ( n7298 & n7299 ) ;
  assign n7301 = n7188 & ~n7300 ;
  assign n7302 = ~n7188 & n7300 ;
  assign n7303 = n7301 | n7302 ;
  assign n7304 = n7290 | n7291 ;
  assign n7305 = n7160 | n7290 ;
  assign n7306 = ( n7290 & n7291 ) | ( n7290 & n7305 ) | ( n7291 & n7305 ) ;
  assign n7307 = ( n7169 & n7304 ) | ( n7169 & n7306 ) | ( n7304 & n7306 ) ;
  assign n7308 = n3446 & ~n4854 ;
  assign n7309 = n3285 & n3446 ;
  assign n7310 = n3222 & n7309 ;
  assign n7311 = ( n4855 & n7308 ) | ( n4855 & n7310 ) | ( n7308 & n7310 ) ;
  assign n7312 = n3448 & ~n5080 ;
  assign n7313 = n3477 & n4830 ;
  assign n7314 = n7312 | n7313 ;
  assign n7315 = n7311 | n7314 ;
  assign n7316 = n3452 | n7315 ;
  assign n7317 = ( ~n5099 & n7315 ) | ( ~n5099 & n7316 ) | ( n7315 & n7316 ) ;
  assign n7318 = n879 & n7315 ;
  assign n7319 = ( n879 & n5943 ) | ( n879 & n7315 ) | ( n5943 & n7315 ) ;
  assign n7320 = ( ~n5099 & n7318 ) | ( ~n5099 & n7319 ) | ( n7318 & n7319 ) ;
  assign n7321 = n7317 & ~n7320 ;
  assign n7322 = n879 & ~n7315 ;
  assign n7323 = n879 & ~n3452 ;
  assign n7324 = ~n7315 & n7323 ;
  assign n7325 = ( n5099 & n7322 ) | ( n5099 & n7324 ) | ( n7322 & n7324 ) ;
  assign n7326 = n7321 | n7325 ;
  assign n7327 = n3423 & ~n5315 ;
  assign n7328 = n3423 & n5303 ;
  assign n7329 = n3423 & ~n5075 ;
  assign n7330 = ( ~n3222 & n3423 ) | ( ~n3222 & n7329 ) | ( n3423 & n7329 ) ;
  assign n7331 = ( ~n5304 & n7328 ) | ( ~n5304 & n7330 ) | ( n7328 & n7330 ) ;
  assign n7332 = ( n5316 & n7327 ) | ( n5316 & n7331 ) | ( n7327 & n7331 ) ;
  assign n7333 = n3412 & n5303 ;
  assign n7334 = n3412 & ~n5075 ;
  assign n7335 = ( ~n3222 & n3412 ) | ( ~n3222 & n7334 ) | ( n3412 & n7334 ) ;
  assign n7336 = ( ~n5304 & n7333 ) | ( ~n5304 & n7335 ) | ( n7333 & n7335 ) ;
  assign n7337 = n7332 | n7336 ;
  assign n7338 = n7331 | n7336 ;
  assign n7339 = ( ~n5534 & n7336 ) | ( ~n5534 & n7338 ) | ( n7336 & n7338 ) ;
  assign n7340 = ( n5093 & n7337 ) | ( n5093 & n7339 ) | ( n7337 & n7339 ) ;
  assign n7341 = ( n5090 & n7337 ) | ( n5090 & n7339 ) | ( n7337 & n7339 ) ;
  assign n7342 = ( n4841 & n7340 ) | ( n4841 & n7341 ) | ( n7340 & n7341 ) ;
  assign n7343 = n634 & n7342 ;
  assign n7344 = n634 | n7342 ;
  assign n7345 = ~n7343 & n7344 ;
  assign n7346 = n7325 & n7345 ;
  assign n7347 = ( n7321 & n7345 ) | ( n7321 & n7346 ) | ( n7345 & n7346 ) ;
  assign n7348 = n7326 & ~n7347 ;
  assign n7349 = ~n7325 & n7345 ;
  assign n7350 = ~n7321 & n7349 ;
  assign n7351 = n7348 | n7350 ;
  assign n7352 = n879 & ~n3289 ;
  assign n7353 = n7198 & ~n7352 ;
  assign n7354 = n7067 & ~n7198 ;
  assign n7355 = ~n7353 & n7354 ;
  assign n7356 = ( n7201 & n7353 ) | ( n7201 & ~n7355 ) | ( n7353 & ~n7355 ) ;
  assign n7357 = ~n7198 & n7352 ;
  assign n7358 = n7353 | n7357 ;
  assign n7359 = ~n7353 & n7357 ;
  assign n7360 = ~n7357 & n7359 ;
  assign n7361 = ( n7356 & ~n7358 ) | ( n7356 & n7360 ) | ( ~n7358 & n7360 ) ;
  assign n7362 = n7354 & ~n7358 ;
  assign n7363 = n7358 | n7362 ;
  assign n7364 = ( n7224 & ~n7361 ) | ( n7224 & n7363 ) | ( ~n7361 & n7363 ) ;
  assign n7365 = ( ~n7067 & n7198 ) | ( ~n7067 & n7352 ) | ( n7198 & n7352 ) ;
  assign n7366 = ( n7352 & n7357 ) | ( n7352 & ~n7365 ) | ( n7357 & ~n7365 ) ;
  assign n7367 = ( n7198 & n7357 ) | ( n7198 & ~n7365 ) | ( n7357 & ~n7365 ) ;
  assign n7368 = ( n7224 & n7366 ) | ( n7224 & n7367 ) | ( n7366 & n7367 ) ;
  assign n7369 = n7364 & ~n7368 ;
  assign n7370 = n7351 & n7369 ;
  assign n7371 = n7351 | n7369 ;
  assign n7372 = ~n7370 & n7371 ;
  assign n7373 = n7229 | n7251 ;
  assign n7374 = ~n7372 & n7373 ;
  assign n7375 = n7229 & ~n7372 ;
  assign n7376 = ( ~n7235 & n7374 ) | ( ~n7235 & n7375 ) | ( n7374 & n7375 ) ;
  assign n7377 = n7372 & ~n7373 ;
  assign n7378 = ~n7229 & n7372 ;
  assign n7379 = ( n7235 & n7377 ) | ( n7235 & n7378 ) | ( n7377 & n7378 ) ;
  assign n7380 = n7376 | n7379 ;
  assign n7381 = n7260 | n7380 ;
  assign n7382 = ( ~n7266 & n7380 ) | ( ~n7266 & n7381 ) | ( n7380 & n7381 ) ;
  assign n7383 = ( ~n7263 & n7380 ) | ( ~n7263 & n7381 ) | ( n7380 & n7381 ) ;
  assign n7384 = ( ~n7264 & n7380 ) | ( ~n7264 & n7381 ) | ( n7380 & n7381 ) ;
  assign n7385 = ( ~n7109 & n7383 ) | ( ~n7109 & n7384 ) | ( n7383 & n7384 ) ;
  assign n7386 = ( ~n6951 & n7382 ) | ( ~n6951 & n7385 ) | ( n7382 & n7385 ) ;
  assign n7387 = n7105 | n7107 ;
  assign n7388 = ( n7381 & n7383 ) | ( n7381 & ~n7387 ) | ( n7383 & ~n7387 ) ;
  assign n7389 = ( ~n7105 & n7381 ) | ( ~n7105 & n7383 ) | ( n7381 & n7383 ) ;
  assign n7390 = n7381 & n7383 ;
  assign n7391 = ( ~n7109 & n7389 ) | ( ~n7109 & n7390 ) | ( n7389 & n7390 ) ;
  assign n7392 = ( ~n6950 & n7388 ) | ( ~n6950 & n7391 ) | ( n7388 & n7391 ) ;
  assign n7393 = ( ~n6716 & n7386 ) | ( ~n6716 & n7392 ) | ( n7386 & n7392 ) ;
  assign n7394 = n7386 & n7392 ;
  assign n7395 = ( ~n6650 & n7393 ) | ( ~n6650 & n7394 ) | ( n7393 & n7394 ) ;
  assign n7396 = ( ~n6722 & n7386 ) | ( ~n6722 & n7392 ) | ( n7386 & n7392 ) ;
  assign n7397 = ( ~n6719 & n7386 ) | ( ~n6719 & n7392 ) | ( n7386 & n7392 ) ;
  assign n7398 = ( ~n6236 & n7396 ) | ( ~n6236 & n7397 ) | ( n7396 & n7397 ) ;
  assign n7399 = ( ~n6073 & n7395 ) | ( ~n6073 & n7398 ) | ( n7395 & n7398 ) ;
  assign n7400 = n7260 & n7380 ;
  assign n7401 = ~n7266 & n7400 ;
  assign n7402 = ~n7263 & n7400 ;
  assign n7403 = ~n7264 & n7400 ;
  assign n7404 = ( ~n7109 & n7402 ) | ( ~n7109 & n7403 ) | ( n7402 & n7403 ) ;
  assign n7405 = ( ~n6951 & n7401 ) | ( ~n6951 & n7404 ) | ( n7401 & n7404 ) ;
  assign n7406 = ( ~n7387 & n7400 ) | ( ~n7387 & n7402 ) | ( n7400 & n7402 ) ;
  assign n7407 = ( ~n7105 & n7400 ) | ( ~n7105 & n7402 ) | ( n7400 & n7402 ) ;
  assign n7408 = n7400 & n7402 ;
  assign n7409 = ( ~n7109 & n7407 ) | ( ~n7109 & n7408 ) | ( n7407 & n7408 ) ;
  assign n7410 = ( ~n6950 & n7406 ) | ( ~n6950 & n7409 ) | ( n7406 & n7409 ) ;
  assign n7411 = ( ~n6716 & n7405 ) | ( ~n6716 & n7410 ) | ( n7405 & n7410 ) ;
  assign n7412 = n7405 & n7410 ;
  assign n7413 = ( ~n6650 & n7411 ) | ( ~n6650 & n7412 ) | ( n7411 & n7412 ) ;
  assign n7414 = ( ~n6722 & n7405 ) | ( ~n6722 & n7410 ) | ( n7405 & n7410 ) ;
  assign n7415 = ( ~n6719 & n7405 ) | ( ~n6719 & n7410 ) | ( n7405 & n7410 ) ;
  assign n7416 = ( ~n6236 & n7414 ) | ( ~n6236 & n7415 ) | ( n7414 & n7415 ) ;
  assign n7417 = ( ~n6073 & n7413 ) | ( ~n6073 & n7416 ) | ( n7413 & n7416 ) ;
  assign n7418 = n7399 & ~n7417 ;
  assign n7419 = n144 | n357 ;
  assign n7420 = n435 | n538 ;
  assign n7421 = n7419 | n7420 ;
  assign n7422 = n495 | n2653 ;
  assign n7423 = n7421 | n7422 ;
  assign n7424 = n503 | n7423 ;
  assign n7425 = n5696 | n7424 ;
  assign n7426 = n2533 | n7425 ;
  assign n7427 = n2643 | n2646 ;
  assign n7428 = n2641 | n7427 ;
  assign n7429 = n141 | n348 ;
  assign n7430 = n241 | n7429 ;
  assign n7431 = n7428 | n7430 ;
  assign n7432 = n7426 | n7431 ;
  assign n7433 = n7418 | n7432 ;
  assign n7434 = n7418 & n7432 ;
  assign n7435 = n7433 & ~n7434 ;
  assign n7436 = n7306 & n7435 ;
  assign n7437 = n7304 & n7435 ;
  assign n7438 = ( n7169 & n7436 ) | ( n7169 & n7437 ) | ( n7436 & n7437 ) ;
  assign n7439 = ~n7304 & n7435 ;
  assign n7440 = ~n7306 & n7435 ;
  assign n7441 = ( ~n7169 & n7439 ) | ( ~n7169 & n7440 ) | ( n7439 & n7440 ) ;
  assign n7442 = ( n7307 & ~n7438 ) | ( n7307 & n7441 ) | ( ~n7438 & n7441 ) ;
  assign n7443 = n7296 & n7442 ;
  assign n7444 = n7177 & n7443 ;
  assign n7445 = n7296 | n7442 ;
  assign n7446 = ( n7177 & n7442 ) | ( n7177 & n7445 ) | ( n7442 & n7445 ) ;
  assign n7447 = ~n7444 & n7446 ;
  assign n7448 = n7187 | n7300 ;
  assign n7449 = n5520 & n7448 ;
  assign n7450 = ~n7447 & n7449 ;
  assign n7451 = n7447 & ~n7449 ;
  assign n7452 = n7450 | n7451 ;
  assign n7453 = n7434 | n7435 ;
  assign n7454 = ( n7306 & n7434 ) | ( n7306 & n7453 ) | ( n7434 & n7453 ) ;
  assign n7455 = ( n7304 & n7434 ) | ( n7304 & n7453 ) | ( n7434 & n7453 ) ;
  assign n7456 = ( n7169 & n7454 ) | ( n7169 & n7455 ) | ( n7454 & n7455 ) ;
  assign n7457 = ~n7347 & n7369 ;
  assign n7458 = ( n7347 & n7351 ) | ( n7347 & ~n7457 ) | ( n7351 & ~n7457 ) ;
  assign n7459 = n3446 & ~n5080 ;
  assign n7460 = n3477 & ~n4854 ;
  assign n7461 = n3285 & n3477 ;
  assign n7462 = n3222 & n7461 ;
  assign n7463 = ( n4855 & n7460 ) | ( n4855 & n7462 ) | ( n7460 & n7462 ) ;
  assign n7464 = n7459 | n7463 ;
  assign n7465 = n3448 & n5303 ;
  assign n7466 = n3448 & ~n5075 ;
  assign n7467 = ( ~n3222 & n3448 ) | ( ~n3222 & n7466 ) | ( n3448 & n7466 ) ;
  assign n7468 = ( ~n5304 & n7465 ) | ( ~n5304 & n7467 ) | ( n7465 & n7467 ) ;
  assign n7469 = n7464 | n7468 ;
  assign n7470 = n3452 | n7468 ;
  assign n7471 = n7464 | n7470 ;
  assign n7472 = ( n5325 & n7469 ) | ( n5325 & n7471 ) | ( n7469 & n7471 ) ;
  assign n7473 = n879 & n7471 ;
  assign n7474 = n879 & n7468 ;
  assign n7475 = ( n879 & n7464 ) | ( n879 & n7474 ) | ( n7464 & n7474 ) ;
  assign n7476 = ( n5325 & n7473 ) | ( n5325 & n7475 ) | ( n7473 & n7475 ) ;
  assign n7477 = n7472 & ~n7476 ;
  assign n7478 = n879 & ~n7475 ;
  assign n7479 = n879 & ~n7471 ;
  assign n7480 = ( ~n5325 & n7478 ) | ( ~n5325 & n7479 ) | ( n7478 & n7479 ) ;
  assign n7481 = n7477 | n7480 ;
  assign n7482 = ~n634 & n879 ;
  assign n7483 = ~n3289 & n7482 ;
  assign n7484 = n634 & ~n879 ;
  assign n7485 = ( n634 & n3289 ) | ( n634 & n7484 ) | ( n3289 & n7484 ) ;
  assign n7486 = n7483 | n7485 ;
  assign n7487 = n879 & n4830 ;
  assign n7488 = ~n7486 & n7487 ;
  assign n7489 = n7486 & ~n7487 ;
  assign n7490 = n7488 | n7489 ;
  assign n7491 = n7479 & ~n7490 ;
  assign n7492 = n7478 & ~n7490 ;
  assign n7493 = ( ~n5325 & n7491 ) | ( ~n5325 & n7492 ) | ( n7491 & n7492 ) ;
  assign n7494 = ( n7477 & ~n7490 ) | ( n7477 & n7493 ) | ( ~n7490 & n7493 ) ;
  assign n7495 = n7481 & ~n7494 ;
  assign n7496 = n7478 | n7490 ;
  assign n7497 = n7479 | n7490 ;
  assign n7498 = ( ~n5325 & n7496 ) | ( ~n5325 & n7497 ) | ( n7496 & n7497 ) ;
  assign n7499 = n7477 | n7498 ;
  assign n7500 = ~n7495 & n7499 ;
  assign n7501 = n7353 | n7362 ;
  assign n7502 = ( ~n7353 & n7356 ) | ( ~n7353 & n7359 ) | ( n7356 & n7359 ) ;
  assign n7503 = ( n7224 & n7501 ) | ( n7224 & ~n7502 ) | ( n7501 & ~n7502 ) ;
  assign n7504 = n7499 & n7503 ;
  assign n7505 = ~n7495 & n7504 ;
  assign n7506 = n7503 & ~n7505 ;
  assign n7507 = ( n7500 & ~n7505 ) | ( n7500 & n7506 ) | ( ~n7505 & n7506 ) ;
  assign n7508 = n7458 & ~n7507 ;
  assign n7509 = ~n7458 & n7507 ;
  assign n7510 = n7508 | n7509 ;
  assign n7511 = n7376 & ~n7510 ;
  assign n7512 = ( n7381 & n7510 ) | ( n7381 & ~n7511 ) | ( n7510 & ~n7511 ) ;
  assign n7513 = ( n7380 & n7510 ) | ( n7380 & ~n7511 ) | ( n7510 & ~n7511 ) ;
  assign n7514 = ( ~n7266 & n7512 ) | ( ~n7266 & n7513 ) | ( n7512 & n7513 ) ;
  assign n7515 = ( ~n7264 & n7512 ) | ( ~n7264 & n7513 ) | ( n7512 & n7513 ) ;
  assign n7516 = ( ~n7263 & n7512 ) | ( ~n7263 & n7513 ) | ( n7512 & n7513 ) ;
  assign n7517 = ( ~n7109 & n7515 ) | ( ~n7109 & n7516 ) | ( n7515 & n7516 ) ;
  assign n7518 = ( ~n6951 & n7514 ) | ( ~n6951 & n7517 ) | ( n7514 & n7517 ) ;
  assign n7519 = n7105 | n7109 ;
  assign n7520 = ( n7383 & n7510 ) | ( n7383 & ~n7511 ) | ( n7510 & ~n7511 ) ;
  assign n7521 = ( n7512 & ~n7519 ) | ( n7512 & n7520 ) | ( ~n7519 & n7520 ) ;
  assign n7522 = ( ~n7387 & n7512 ) | ( ~n7387 & n7520 ) | ( n7512 & n7520 ) ;
  assign n7523 = ( ~n6950 & n7521 ) | ( ~n6950 & n7522 ) | ( n7521 & n7522 ) ;
  assign n7524 = ( ~n6716 & n7518 ) | ( ~n6716 & n7523 ) | ( n7518 & n7523 ) ;
  assign n7525 = n7518 & n7523 ;
  assign n7526 = ( ~n6650 & n7524 ) | ( ~n6650 & n7525 ) | ( n7524 & n7525 ) ;
  assign n7527 = ( ~n6722 & n7518 ) | ( ~n6722 & n7523 ) | ( n7518 & n7523 ) ;
  assign n7528 = ( ~n6719 & n7518 ) | ( ~n6719 & n7523 ) | ( n7518 & n7523 ) ;
  assign n7529 = ( ~n6236 & n7527 ) | ( ~n6236 & n7528 ) | ( n7527 & n7528 ) ;
  assign n7530 = ( ~n6073 & n7526 ) | ( ~n6073 & n7529 ) | ( n7526 & n7529 ) ;
  assign n7531 = ~n7376 & n7510 ;
  assign n7532 = n7381 & n7531 ;
  assign n7533 = n7380 & n7531 ;
  assign n7534 = ( ~n7266 & n7532 ) | ( ~n7266 & n7533 ) | ( n7532 & n7533 ) ;
  assign n7535 = ( ~n7264 & n7532 ) | ( ~n7264 & n7533 ) | ( n7532 & n7533 ) ;
  assign n7536 = ( ~n7263 & n7532 ) | ( ~n7263 & n7533 ) | ( n7532 & n7533 ) ;
  assign n7537 = ( ~n7109 & n7535 ) | ( ~n7109 & n7536 ) | ( n7535 & n7536 ) ;
  assign n7538 = ( ~n6951 & n7534 ) | ( ~n6951 & n7537 ) | ( n7534 & n7537 ) ;
  assign n7539 = n7383 & n7531 ;
  assign n7540 = ( ~n7519 & n7532 ) | ( ~n7519 & n7539 ) | ( n7532 & n7539 ) ;
  assign n7541 = ( ~n7387 & n7532 ) | ( ~n7387 & n7539 ) | ( n7532 & n7539 ) ;
  assign n7542 = ( ~n6950 & n7540 ) | ( ~n6950 & n7541 ) | ( n7540 & n7541 ) ;
  assign n7543 = ( ~n6716 & n7538 ) | ( ~n6716 & n7542 ) | ( n7538 & n7542 ) ;
  assign n7544 = n7538 & n7542 ;
  assign n7545 = ( ~n6650 & n7543 ) | ( ~n6650 & n7544 ) | ( n7543 & n7544 ) ;
  assign n7546 = ( ~n6722 & n7538 ) | ( ~n6722 & n7542 ) | ( n7538 & n7542 ) ;
  assign n7547 = ( ~n6719 & n7538 ) | ( ~n6719 & n7542 ) | ( n7538 & n7542 ) ;
  assign n7548 = ( ~n6236 & n7546 ) | ( ~n6236 & n7547 ) | ( n7546 & n7547 ) ;
  assign n7549 = ( ~n6073 & n7545 ) | ( ~n6073 & n7548 ) | ( n7545 & n7548 ) ;
  assign n7550 = n7530 & ~n7549 ;
  assign n7551 = n293 | n304 ;
  assign n7552 = n384 | n570 ;
  assign n7553 = n7551 | n7552 ;
  assign n7554 = n333 | n392 ;
  assign n7555 = n7553 | n7554 ;
  assign n7556 = n5496 | n7555 ;
  assign n7557 = n806 | n7556 ;
  assign n7558 = n590 | n2949 ;
  assign n7559 = n7557 | n7558 ;
  assign n7560 = n334 | n4998 ;
  assign n7561 = n7559 | n7560 ;
  assign n7562 = n176 | n412 ;
  assign n7563 = n172 | n358 ;
  assign n7564 = n7562 | n7563 ;
  assign n7565 = n224 | n262 ;
  assign n7566 = n7564 | n7565 ;
  assign n7567 = n7561 | n7566 ;
  assign n7568 = n7550 & n7567 ;
  assign n7569 = n7550 | n7567 ;
  assign n7570 = ~n7568 & n7569 ;
  assign n7571 = n7455 & n7570 ;
  assign n7572 = n7454 & n7570 ;
  assign n7573 = ( n7169 & n7571 ) | ( n7169 & n7572 ) | ( n7571 & n7572 ) ;
  assign n7574 = ~n7454 & n7570 ;
  assign n7575 = ~n7455 & n7570 ;
  assign n7576 = ( ~n7169 & n7574 ) | ( ~n7169 & n7575 ) | ( n7574 & n7575 ) ;
  assign n7577 = ( n7456 & ~n7573 ) | ( n7456 & n7576 ) | ( ~n7573 & n7576 ) ;
  assign n7578 = n7443 & n7577 ;
  assign n7579 = n7177 & n7578 ;
  assign n7580 = n7443 | n7577 ;
  assign n7581 = ( n7177 & n7577 ) | ( n7177 & n7580 ) | ( n7577 & n7580 ) ;
  assign n7582 = ~n7579 & n7581 ;
  assign n7583 = n7300 | n7447 ;
  assign n7584 = n7187 | n7583 ;
  assign n7585 = n5520 & n7584 ;
  assign n7586 = ~n7582 & n7585 ;
  assign n7587 = n7582 & ~n7585 ;
  assign n7588 = n7586 | n7587 ;
  assign n7589 = n2653 | n2723 ;
  assign n7590 = n740 | n7589 ;
  assign n7591 = n617 | n7590 ;
  assign n7592 = n857 | n7591 ;
  assign n7593 = n2933 | n7592 ;
  assign n7594 = n150 | n343 ;
  assign n7595 = n353 | n7594 ;
  assign n7596 = ( ~n593 & n4822 ) | ( ~n593 & n7595 ) | ( n4822 & n7595 ) ;
  assign n7597 = n352 | n412 ;
  assign n7598 = n220 | n320 ;
  assign n7599 = n7597 | n7598 ;
  assign n7600 = n593 | n7599 ;
  assign n7601 = n7596 | n7600 ;
  assign n7602 = n7593 | n7601 ;
  assign n7603 = ~n7508 & n7523 ;
  assign n7604 = ~n7508 & n7517 ;
  assign n7605 = ~n7508 & n7514 ;
  assign n7606 = ( ~n6951 & n7604 ) | ( ~n6951 & n7605 ) | ( n7604 & n7605 ) ;
  assign n7607 = ( ~n6716 & n7603 ) | ( ~n6716 & n7606 ) | ( n7603 & n7606 ) ;
  assign n7608 = n7603 & n7606 ;
  assign n7609 = ( ~n6650 & n7607 ) | ( ~n6650 & n7608 ) | ( n7607 & n7608 ) ;
  assign n7610 = ( ~n6722 & n7603 ) | ( ~n6722 & n7606 ) | ( n7603 & n7606 ) ;
  assign n7611 = ( ~n6719 & n7603 ) | ( ~n6719 & n7606 ) | ( n7603 & n7606 ) ;
  assign n7612 = ( ~n6236 & n7610 ) | ( ~n6236 & n7611 ) | ( n7610 & n7611 ) ;
  assign n7613 = ( ~n6073 & n7609 ) | ( ~n6073 & n7612 ) | ( n7609 & n7612 ) ;
  assign n7614 = n7483 | n7487 ;
  assign n7615 = ( n7483 & ~n7486 ) | ( n7483 & n7614 ) | ( ~n7486 & n7614 ) ;
  assign n7616 = n879 & ~n4854 ;
  assign n7617 = n879 & n3285 ;
  assign n7618 = n3222 & n7617 ;
  assign n7619 = ( n4855 & n7616 ) | ( n4855 & n7618 ) | ( n7616 & n7618 ) ;
  assign n7620 = n7615 & ~n7619 ;
  assign n7621 = n7615 & ~n7620 ;
  assign n7622 = n7615 | n7619 ;
  assign n7623 = ~n7621 & n7622 ;
  assign n7624 = n3446 & n5303 ;
  assign n7625 = n3446 & ~n5075 ;
  assign n7626 = ( ~n3222 & n3446 ) | ( ~n3222 & n7625 ) | ( n3446 & n7625 ) ;
  assign n7627 = ( ~n5304 & n7624 ) | ( ~n5304 & n7626 ) | ( n7624 & n7626 ) ;
  assign n7628 = ( n3452 & n3487 ) | ( n3452 & ~n5080 ) | ( n3487 & ~n5080 ) ;
  assign n7629 = n7627 | n7628 ;
  assign n7630 = ( n879 & n4646 ) | ( n879 & ~n5080 ) | ( n4646 & ~n5080 ) ;
  assign n7631 = n7627 | n7630 ;
  assign n7632 = ( n879 & n7629 ) | ( n879 & n7631 ) | ( n7629 & n7631 ) ;
  assign n7633 = n879 | n3157 ;
  assign n7634 = ( n879 & n3440 ) | ( n879 & n7633 ) | ( n3440 & n7633 ) ;
  assign n7635 = n3477 | n7634 ;
  assign n7636 = ( ~n5080 & n7634 ) | ( ~n5080 & n7635 ) | ( n7634 & n7635 ) ;
  assign n7637 = n7627 | n7636 ;
  assign n7638 = ( n5546 & n7632 ) | ( n5546 & n7637 ) | ( n7632 & n7637 ) ;
  assign n7639 = n4636 & ~n5080 ;
  assign n7640 = ( n879 & n7627 ) | ( n879 & n7639 ) | ( n7627 & n7639 ) ;
  assign n7641 = n7629 & n7640 ;
  assign n7642 = n879 | n5943 ;
  assign n7643 = ( n879 & n3477 ) | ( n879 & n5943 ) | ( n3477 & n5943 ) ;
  assign n7644 = n879 & n5943 ;
  assign n7645 = ( ~n5080 & n7643 ) | ( ~n5080 & n7644 ) | ( n7643 & n7644 ) ;
  assign n7646 = ( n7627 & n7642 ) | ( n7627 & n7645 ) | ( n7642 & n7645 ) ;
  assign n7647 = ( n5546 & n7641 ) | ( n5546 & n7646 ) | ( n7641 & n7646 ) ;
  assign n7648 = n7638 & ~n7647 ;
  assign n7649 = ~n7623 & n7648 ;
  assign n7650 = n7623 & ~n7648 ;
  assign n7651 = n7649 | n7650 ;
  assign n7652 = n7494 | n7503 ;
  assign n7653 = ~n7651 & n7652 ;
  assign n7654 = n7494 & ~n7651 ;
  assign n7655 = ( ~n7500 & n7653 ) | ( ~n7500 & n7654 ) | ( n7653 & n7654 ) ;
  assign n7656 = n7651 & ~n7652 ;
  assign n7657 = ~n7494 & n7651 ;
  assign n7658 = ( n7500 & n7656 ) | ( n7500 & n7657 ) | ( n7656 & n7657 ) ;
  assign n7659 = n7655 | n7658 ;
  assign n7660 = n7612 & n7659 ;
  assign n7661 = n7608 & n7659 ;
  assign n7662 = n7607 & n7659 ;
  assign n7663 = ( ~n6650 & n7661 ) | ( ~n6650 & n7662 ) | ( n7661 & n7662 ) ;
  assign n7664 = ( ~n6073 & n7660 ) | ( ~n6073 & n7663 ) | ( n7660 & n7663 ) ;
  assign n7665 = n7659 & ~n7663 ;
  assign n7666 = ~n7612 & n7659 ;
  assign n7667 = ( n6073 & n7665 ) | ( n6073 & n7666 ) | ( n7665 & n7666 ) ;
  assign n7668 = ( n7613 & ~n7664 ) | ( n7613 & n7667 ) | ( ~n7664 & n7667 ) ;
  assign n7669 = n7602 | n7668 ;
  assign n7670 = n7602 & n7668 ;
  assign n7671 = n7669 & ~n7670 ;
  assign n7672 = n7568 | n7570 ;
  assign n7673 = n7671 & n7672 ;
  assign n7674 = n7568 & n7671 ;
  assign n7675 = ( n7455 & n7673 ) | ( n7455 & n7674 ) | ( n7673 & n7674 ) ;
  assign n7676 = ( n7454 & n7673 ) | ( n7454 & n7674 ) | ( n7673 & n7674 ) ;
  assign n7677 = ( n7169 & n7675 ) | ( n7169 & n7676 ) | ( n7675 & n7676 ) ;
  assign n7678 = n7671 | n7672 ;
  assign n7679 = n7568 | n7671 ;
  assign n7680 = ( n7455 & n7678 ) | ( n7455 & n7679 ) | ( n7678 & n7679 ) ;
  assign n7681 = ( n7454 & n7678 ) | ( n7454 & n7679 ) | ( n7678 & n7679 ) ;
  assign n7682 = ( n7169 & n7680 ) | ( n7169 & n7681 ) | ( n7680 & n7681 ) ;
  assign n7683 = ~n7677 & n7682 ;
  assign n7684 = n7579 | n7683 ;
  assign n7685 = n7579 & n7683 ;
  assign n7686 = n7684 & ~n7685 ;
  assign n7687 = n7582 | n7584 ;
  assign n7688 = n5520 & n7687 ;
  assign n7689 = ~n7686 & n7688 ;
  assign n7690 = n7686 & ~n7688 ;
  assign n7691 = n7689 | n7690 ;
  assign n7692 = n879 & ~n5087 ;
  assign n7693 = n3452 & ~n5315 ;
  assign n7694 = n3452 & n5303 ;
  assign n7695 = n3452 & ~n5075 ;
  assign n7696 = ( ~n3222 & n3452 ) | ( ~n3222 & n7695 ) | ( n3452 & n7695 ) ;
  assign n7697 = ( ~n5304 & n7694 ) | ( ~n5304 & n7696 ) | ( n7694 & n7696 ) ;
  assign n7698 = ( n5316 & n7693 ) | ( n5316 & n7697 ) | ( n7693 & n7697 ) ;
  assign n7699 = n3477 & n5303 ;
  assign n7700 = n3477 & ~n5075 ;
  assign n7701 = ( ~n3222 & n3477 ) | ( ~n3222 & n7700 ) | ( n3477 & n7700 ) ;
  assign n7702 = ( ~n5304 & n7699 ) | ( ~n5304 & n7701 ) | ( n7699 & n7701 ) ;
  assign n7703 = n7698 | n7702 ;
  assign n7704 = n7697 | n7702 ;
  assign n7705 = ( ~n5534 & n7702 ) | ( ~n5534 & n7704 ) | ( n7702 & n7704 ) ;
  assign n7706 = ( n5093 & n7703 ) | ( n5093 & n7705 ) | ( n7703 & n7705 ) ;
  assign n7707 = ( n5090 & n7703 ) | ( n5090 & n7705 ) | ( n7703 & n7705 ) ;
  assign n7708 = ( n4841 & n7706 ) | ( n4841 & n7707 ) | ( n7706 & n7707 ) ;
  assign n7709 = ( n879 & n7692 ) | ( n879 & ~n7708 ) | ( n7692 & ~n7708 ) ;
  assign n7710 = ( ~n879 & n7708 ) | ( ~n879 & n7709 ) | ( n7708 & n7709 ) ;
  assign n7711 = ( ~n7692 & n7709 ) | ( ~n7692 & n7710 ) | ( n7709 & n7710 ) ;
  assign n7712 = ( n7615 & ~n7619 ) | ( n7615 & n7648 ) | ( ~n7619 & n7648 ) ;
  assign n7713 = n7711 & ~n7712 ;
  assign n7714 = ~n7711 & n7712 ;
  assign n7715 = n7713 | n7714 ;
  assign n7716 = n7655 & ~n7715 ;
  assign n7717 = ( n7659 & n7715 ) | ( n7659 & ~n7716 ) | ( n7715 & ~n7716 ) ;
  assign n7718 = ( n7608 & ~n7716 ) | ( n7608 & n7717 ) | ( ~n7716 & n7717 ) ;
  assign n7719 = ( n7607 & ~n7716 ) | ( n7607 & n7717 ) | ( ~n7716 & n7717 ) ;
  assign n7720 = ( ~n6650 & n7718 ) | ( ~n6650 & n7719 ) | ( n7718 & n7719 ) ;
  assign n7721 = ( n7605 & ~n7716 ) | ( n7605 & n7717 ) | ( ~n7716 & n7717 ) ;
  assign n7722 = ( n7604 & ~n7716 ) | ( n7604 & n7717 ) | ( ~n7716 & n7717 ) ;
  assign n7723 = ( ~n6951 & n7721 ) | ( ~n6951 & n7722 ) | ( n7721 & n7722 ) ;
  assign n7724 = ( n7508 & n7716 ) | ( n7508 & ~n7717 ) | ( n7716 & ~n7717 ) ;
  assign n7725 = ~n7716 & n7717 ;
  assign n7726 = ( n7523 & ~n7724 ) | ( n7523 & n7725 ) | ( ~n7724 & n7725 ) ;
  assign n7727 = ( ~n6722 & n7723 ) | ( ~n6722 & n7726 ) | ( n7723 & n7726 ) ;
  assign n7728 = ( ~n6719 & n7723 ) | ( ~n6719 & n7726 ) | ( n7723 & n7726 ) ;
  assign n7729 = ( ~n6236 & n7727 ) | ( ~n6236 & n7728 ) | ( n7727 & n7728 ) ;
  assign n7730 = ( ~n6073 & n7720 ) | ( ~n6073 & n7729 ) | ( n7720 & n7729 ) ;
  assign n7731 = ~n7655 & n7715 ;
  assign n7732 = n7659 & n7731 ;
  assign n7733 = ( n7608 & n7731 ) | ( n7608 & n7732 ) | ( n7731 & n7732 ) ;
  assign n7734 = ( n7607 & n7731 ) | ( n7607 & n7732 ) | ( n7731 & n7732 ) ;
  assign n7735 = ( ~n6650 & n7733 ) | ( ~n6650 & n7734 ) | ( n7733 & n7734 ) ;
  assign n7736 = ( n7605 & n7731 ) | ( n7605 & n7732 ) | ( n7731 & n7732 ) ;
  assign n7737 = ( n7604 & n7731 ) | ( n7604 & n7732 ) | ( n7731 & n7732 ) ;
  assign n7738 = ( ~n6951 & n7736 ) | ( ~n6951 & n7737 ) | ( n7736 & n7737 ) ;
  assign n7739 = ( ~n7508 & n7731 ) | ( ~n7508 & n7732 ) | ( n7731 & n7732 ) ;
  assign n7740 = n7731 & n7732 ;
  assign n7741 = ( n7523 & n7739 ) | ( n7523 & n7740 ) | ( n7739 & n7740 ) ;
  assign n7742 = ( ~n6722 & n7738 ) | ( ~n6722 & n7741 ) | ( n7738 & n7741 ) ;
  assign n7743 = ( ~n6719 & n7738 ) | ( ~n6719 & n7741 ) | ( n7738 & n7741 ) ;
  assign n7744 = ( ~n6236 & n7742 ) | ( ~n6236 & n7743 ) | ( n7742 & n7743 ) ;
  assign n7745 = ( ~n6073 & n7735 ) | ( ~n6073 & n7744 ) | ( n7735 & n7744 ) ;
  assign n7746 = n7730 & ~n7745 ;
  assign n7747 = n495 | n7421 ;
  assign n7748 = n193 | n354 ;
  assign n7749 = n576 | n7748 ;
  assign n7750 = n677 | n7749 ;
  assign n7751 = n7747 | n7750 ;
  assign n7752 = n2660 | n7751 ;
  assign n7753 = n216 | n981 ;
  assign n7754 = n980 | n7753 ;
  assign n7755 = n987 | n7754 ;
  assign n7756 = n977 | n7755 ;
  assign n7757 = n7752 | n7756 ;
  assign n7758 = n220 | n236 ;
  assign n7759 = n229 | n280 ;
  assign n7760 = n267 | n353 ;
  assign n7761 = n795 | n7760 ;
  assign n7762 = n7759 | n7761 ;
  assign n7763 = n794 | n7762 ;
  assign n7764 = n7758 | n7763 ;
  assign n7765 = n7757 | n7764 ;
  assign n7766 = n7746 & n7765 ;
  assign n7767 = n7746 | n7765 ;
  assign n7768 = ~n7766 & n7767 ;
  assign n7769 = n7568 | n7670 ;
  assign n7770 = ( n7670 & n7671 ) | ( n7670 & n7769 ) | ( n7671 & n7769 ) ;
  assign n7771 = n7768 & n7770 ;
  assign n7772 = n7670 | n7671 ;
  assign n7773 = ( n7670 & n7672 ) | ( n7670 & n7772 ) | ( n7672 & n7772 ) ;
  assign n7774 = n7768 & n7773 ;
  assign n7775 = ( n7455 & n7771 ) | ( n7455 & n7774 ) | ( n7771 & n7774 ) ;
  assign n7776 = ( n7454 & n7771 ) | ( n7454 & n7774 ) | ( n7771 & n7774 ) ;
  assign n7777 = ( n7169 & n7775 ) | ( n7169 & n7776 ) | ( n7775 & n7776 ) ;
  assign n7778 = ( n7454 & n7770 ) | ( n7454 & n7773 ) | ( n7770 & n7773 ) ;
  assign n7779 = n7768 | n7778 ;
  assign n7780 = ( n7455 & n7770 ) | ( n7455 & n7773 ) | ( n7770 & n7773 ) ;
  assign n7781 = n7768 | n7780 ;
  assign n7782 = ( n7169 & n7779 ) | ( n7169 & n7781 ) | ( n7779 & n7781 ) ;
  assign n7783 = ~n7777 & n7782 ;
  assign n7784 = n7683 & n7783 ;
  assign n7785 = n7579 & n7784 ;
  assign n7786 = n7683 | n7783 ;
  assign n7787 = ( n7579 & n7783 ) | ( n7579 & n7786 ) | ( n7783 & n7786 ) ;
  assign n7788 = ~n7785 & n7787 ;
  assign n7789 = n7686 | n7687 ;
  assign n7790 = n5520 & n7789 ;
  assign n7791 = ~n7788 & n7790 ;
  assign n7792 = n7788 & ~n7790 ;
  assign n7793 = n7791 | n7792 ;
  assign n7794 = n7686 | n7788 ;
  assign n7795 = n7687 | n7794 ;
  assign n7796 = n5520 & n7795 ;
  assign n7797 = n879 & n7708 ;
  assign n7798 = n7708 & ~n7797 ;
  assign n7799 = n879 & ~n5080 ;
  assign n7800 = ~n7619 & n7799 ;
  assign n7801 = n7692 & ~n7800 ;
  assign n7802 = n879 & n5087 ;
  assign n7803 = n7800 | n7802 ;
  assign n7804 = ( ~n7708 & n7800 ) | ( ~n7708 & n7803 ) | ( n7800 & n7803 ) ;
  assign n7805 = ( n7798 & ~n7801 ) | ( n7798 & n7804 ) | ( ~n7801 & n7804 ) ;
  assign n7806 = n7711 | n7805 ;
  assign n7807 = n7712 & ~n7806 ;
  assign n7808 = ( n7717 & n7805 ) | ( n7717 & ~n7807 ) | ( n7805 & ~n7807 ) ;
  assign n7809 = ( n7715 & n7805 ) | ( n7715 & ~n7807 ) | ( n7805 & ~n7807 ) ;
  assign n7810 = ~n7805 & n7807 ;
  assign n7811 = ( n7655 & ~n7809 ) | ( n7655 & n7810 ) | ( ~n7809 & n7810 ) ;
  assign n7812 = ( n7608 & n7808 ) | ( n7608 & ~n7811 ) | ( n7808 & ~n7811 ) ;
  assign n7813 = ( n7607 & n7808 ) | ( n7607 & ~n7811 ) | ( n7808 & ~n7811 ) ;
  assign n7814 = ( ~n6650 & n7812 ) | ( ~n6650 & n7813 ) | ( n7812 & n7813 ) ;
  assign n7815 = ( n7605 & n7808 ) | ( n7605 & ~n7811 ) | ( n7808 & ~n7811 ) ;
  assign n7816 = ( n7604 & n7808 ) | ( n7604 & ~n7811 ) | ( n7808 & ~n7811 ) ;
  assign n7817 = ( ~n6951 & n7815 ) | ( ~n6951 & n7816 ) | ( n7815 & n7816 ) ;
  assign n7818 = ( n7508 & ~n7808 ) | ( n7508 & n7811 ) | ( ~n7808 & n7811 ) ;
  assign n7819 = n7808 & ~n7811 ;
  assign n7820 = ( n7523 & ~n7818 ) | ( n7523 & n7819 ) | ( ~n7818 & n7819 ) ;
  assign n7821 = ( ~n6722 & n7817 ) | ( ~n6722 & n7820 ) | ( n7817 & n7820 ) ;
  assign n7822 = ( ~n6719 & n7817 ) | ( ~n6719 & n7820 ) | ( n7817 & n7820 ) ;
  assign n7823 = ( ~n6236 & n7821 ) | ( ~n6236 & n7822 ) | ( n7821 & n7822 ) ;
  assign n7824 = ( ~n6073 & n7814 ) | ( ~n6073 & n7823 ) | ( n7814 & n7823 ) ;
  assign n7825 = n7711 & n7805 ;
  assign n7826 = ( ~n7712 & n7805 ) | ( ~n7712 & n7825 ) | ( n7805 & n7825 ) ;
  assign n7827 = n7717 & n7826 ;
  assign n7828 = n7715 & n7826 ;
  assign n7829 = ( ~n7655 & n7826 ) | ( ~n7655 & n7828 ) | ( n7826 & n7828 ) ;
  assign n7830 = ( n7608 & n7827 ) | ( n7608 & n7829 ) | ( n7827 & n7829 ) ;
  assign n7831 = ( n7607 & n7827 ) | ( n7607 & n7829 ) | ( n7827 & n7829 ) ;
  assign n7832 = ( ~n6650 & n7830 ) | ( ~n6650 & n7831 ) | ( n7830 & n7831 ) ;
  assign n7833 = ( n7605 & n7827 ) | ( n7605 & n7829 ) | ( n7827 & n7829 ) ;
  assign n7834 = ( n7604 & n7827 ) | ( n7604 & n7829 ) | ( n7827 & n7829 ) ;
  assign n7835 = ( ~n6951 & n7833 ) | ( ~n6951 & n7834 ) | ( n7833 & n7834 ) ;
  assign n7836 = ( ~n7508 & n7827 ) | ( ~n7508 & n7829 ) | ( n7827 & n7829 ) ;
  assign n7837 = n7827 & n7829 ;
  assign n7838 = ( n7523 & n7836 ) | ( n7523 & n7837 ) | ( n7836 & n7837 ) ;
  assign n7839 = ( ~n6722 & n7835 ) | ( ~n6722 & n7838 ) | ( n7835 & n7838 ) ;
  assign n7840 = ( ~n6719 & n7835 ) | ( ~n6719 & n7838 ) | ( n7835 & n7838 ) ;
  assign n7841 = ( ~n6236 & n7839 ) | ( ~n6236 & n7840 ) | ( n7839 & n7840 ) ;
  assign n7842 = ( ~n6073 & n7832 ) | ( ~n6073 & n7841 ) | ( n7832 & n7841 ) ;
  assign n7843 = n7824 & ~n7842 ;
  assign n7844 = n879 & n7619 ;
  assign n7845 = n879 & ~n5303 ;
  assign n7846 = n879 & n5300 ;
  assign n7847 = ( n5304 & n7845 ) | ( n5304 & n7846 ) | ( n7845 & n7846 ) ;
  assign n7848 = ( n7843 & n7844 ) | ( n7843 & n7847 ) | ( n7844 & n7847 ) ;
  assign n7849 = ( ~n7843 & n7844 ) | ( ~n7843 & n7847 ) | ( n7844 & n7847 ) ;
  assign n7850 = ( n7843 & ~n7848 ) | ( n7843 & n7849 ) | ( ~n7848 & n7849 ) ;
  assign n7851 = n333 | n7553 ;
  assign n7852 = n523 | n2293 ;
  assign n7853 = n2538 | n7852 ;
  assign n7854 = n7851 | n7853 ;
  assign n7855 = n230 | n4950 ;
  assign n7856 = n4949 | n7855 ;
  assign n7857 = n7854 | n7856 ;
  assign n7858 = n202 | n330 ;
  assign n7859 = n429 | n7858 ;
  assign n7860 = n292 | n4985 ;
  assign n7861 = n3173 | n7860 ;
  assign n7862 = n7859 | n7861 ;
  assign n7863 = n4984 | n7862 ;
  assign n7864 = n7857 | n7863 ;
  assign n7865 = n2289 | n7864 ;
  assign n7866 = n7850 & n7865 ;
  assign n7867 = n7765 & n7865 ;
  assign n7868 = n7746 & n7867 ;
  assign n7869 = ( n7766 & n7850 ) | ( n7766 & n7868 ) | ( n7850 & n7868 ) ;
  assign n7870 = ~n7866 & n7869 ;
  assign n7871 = n7850 | n7865 ;
  assign n7872 = ~n7866 & n7871 ;
  assign n7873 = ( n7777 & n7870 ) | ( n7777 & n7872 ) | ( n7870 & n7872 ) ;
  assign n7874 = n7766 | n7872 ;
  assign n7875 = n7777 | n7874 ;
  assign n7876 = ~n7873 & n7875 ;
  assign n7877 = n7784 & ~n7876 ;
  assign n7878 = n7579 & n7877 ;
  assign n7879 = n7876 | n7877 ;
  assign n7880 = ( n7579 & n7876 ) | ( n7579 & n7879 ) | ( n7876 & n7879 ) ;
  assign n7881 = ( ~n7785 & n7878 ) | ( ~n7785 & n7880 ) | ( n7878 & n7880 ) ;
  assign n7882 = n7796 & ~n7881 ;
  assign n7883 = ~n7796 & n7881 ;
  assign n7884 = n7882 | n7883 ;
  assign n7885 = n7795 | n7881 ;
  assign n7886 = n5520 & n7885 ;
  assign n7887 = n442 | n460 ;
  assign n7888 = n317 | n393 ;
  assign n7889 = n187 | n549 ;
  assign n7890 = n7888 | n7889 ;
  assign n7891 = n3175 | n7890 ;
  assign n7892 = n3253 | n7891 ;
  assign n7893 = n7887 | n7892 ;
  assign n7894 = n241 | n538 ;
  assign n7895 = n590 | n7894 ;
  assign n7896 = n139 | n323 ;
  assign n7897 = n7895 | n7896 ;
  assign n7898 = n7893 | n7897 ;
  assign n7899 = n7865 & n7898 ;
  assign n7900 = n7850 & n7899 ;
  assign n7901 = ( n7870 & n7898 ) | ( n7870 & n7900 ) | ( n7898 & n7900 ) ;
  assign n7902 = ( n7872 & n7898 ) | ( n7872 & n7900 ) | ( n7898 & n7900 ) ;
  assign n7903 = ( n7777 & n7901 ) | ( n7777 & n7902 ) | ( n7901 & n7902 ) ;
  assign n7904 = n7865 | n7898 ;
  assign n7905 = ( n7850 & n7898 ) | ( n7850 & n7904 ) | ( n7898 & n7904 ) ;
  assign n7906 = n7872 | n7905 ;
  assign n7907 = n7870 | n7905 ;
  assign n7908 = ( n7777 & n7906 ) | ( n7777 & n7907 ) | ( n7906 & n7907 ) ;
  assign n7909 = ~n7903 & n7908 ;
  assign n7910 = n7784 & n7876 ;
  assign n7911 = ~n7909 & n7910 ;
  assign n7912 = n7579 & n7911 ;
  assign n7913 = n7909 | n7912 ;
  assign n7914 = n7579 & n7910 ;
  assign n7915 = ( n7912 & n7913 ) | ( n7912 & ~n7914 ) | ( n7913 & ~n7914 ) ;
  assign n7916 = n7886 & n7915 ;
  assign n7917 = n7886 | n7915 ;
  assign n7918 = ~n7916 & n7917 ;
  assign n7919 = n7881 | n7915 ;
  assign n7920 = n7795 | n7919 ;
  assign n7921 = n5520 & n7920 ;
  assign n7922 = n7876 & n7909 ;
  assign n7923 = n511 | n2940 ;
  assign n7924 = n673 | n7923 ;
  assign n7925 = n951 | n7924 ;
  assign n7926 = n406 | n7925 ;
  assign n7927 = n597 | n790 ;
  assign n7928 = n7926 | n7927 ;
  assign n7929 = n283 | n538 ;
  assign n7930 = n248 | n301 ;
  assign n7931 = n7929 | n7930 ;
  assign n7932 = n343 | n7931 ;
  assign n7933 = n5034 | n7932 ;
  assign n7934 = n7928 | n7933 ;
  assign n7935 = n7900 | n7934 ;
  assign n7936 = n7898 | n7934 ;
  assign n7937 = ( n7872 & n7935 ) | ( n7872 & n7936 ) | ( n7935 & n7936 ) ;
  assign n7938 = ( n7870 & n7935 ) | ( n7870 & n7936 ) | ( n7935 & n7936 ) ;
  assign n7939 = ( n7777 & n7937 ) | ( n7777 & n7938 ) | ( n7937 & n7938 ) ;
  assign n7940 = ~n7784 & n7922 ;
  assign n7941 = ( ~n7579 & n7922 ) | ( ~n7579 & n7940 ) | ( n7922 & n7940 ) ;
  assign n7942 = ( n7922 & ~n7939 ) | ( n7922 & n7941 ) | ( ~n7939 & n7941 ) ;
  assign n7943 = n7900 & n7934 ;
  assign n7944 = n7898 & n7934 ;
  assign n7945 = ( n7872 & n7943 ) | ( n7872 & n7944 ) | ( n7943 & n7944 ) ;
  assign n7946 = ( n7870 & n7943 ) | ( n7870 & n7944 ) | ( n7943 & n7944 ) ;
  assign n7947 = ( n7777 & n7945 ) | ( n7777 & n7946 ) | ( n7945 & n7946 ) ;
  assign n7948 = n7939 & ~n7947 ;
  assign n7949 = ( n7922 & ~n7941 ) | ( n7922 & n7948 ) | ( ~n7941 & n7948 ) ;
  assign n7950 = ( ~n7922 & n7942 ) | ( ~n7922 & n7949 ) | ( n7942 & n7949 ) ;
  assign n7951 = n7921 & ~n7950 ;
  assign n7952 = ~n7921 & n7950 ;
  assign n7953 = n7951 | n7952 ;
  assign n7954 = n7920 | n7950 ;
  assign n7955 = n5520 & n7954 ;
  assign n7983 = n7784 & n7922 ;
  assign n7984 = n7579 & n7983 ;
  assign n7956 = n664 | n7748 ;
  assign n7957 = n6243 | n7956 ;
  assign n7958 = n3201 | n7957 ;
  assign n7959 = n536 | n7958 ;
  assign n7960 = n7756 | n7959 ;
  assign n7961 = n289 | n321 ;
  assign n7962 = n397 | n429 ;
  assign n7963 = n7961 | n7962 ;
  assign n7964 = n173 | n548 ;
  assign n7965 = n245 | n7964 ;
  assign n7966 = n7963 | n7965 ;
  assign n7967 = n7960 | n7966 ;
  assign n7968 = n7934 | n7967 ;
  assign n7969 = ( n7898 & n7967 ) | ( n7898 & n7968 ) | ( n7967 & n7968 ) ;
  assign n7970 = ( n7899 & n7967 ) | ( n7899 & n7968 ) | ( n7967 & n7968 ) ;
  assign n7971 = n7967 & n7968 ;
  assign n7972 = ( n7850 & n7970 ) | ( n7850 & n7971 ) | ( n7970 & n7971 ) ;
  assign n7973 = ( n7872 & n7969 ) | ( n7872 & n7972 ) | ( n7969 & n7972 ) ;
  assign n7974 = ( n7870 & n7969 ) | ( n7870 & n7972 ) | ( n7969 & n7972 ) ;
  assign n7975 = ( n7777 & n7973 ) | ( n7777 & n7974 ) | ( n7973 & n7974 ) ;
  assign n7976 = n7934 & n7967 ;
  assign n7977 = n7900 & n7976 ;
  assign n7978 = n7898 & n7976 ;
  assign n7979 = ( n7872 & n7977 ) | ( n7872 & n7978 ) | ( n7977 & n7978 ) ;
  assign n7980 = ( n7870 & n7977 ) | ( n7870 & n7978 ) | ( n7977 & n7978 ) ;
  assign n7981 = ( n7777 & n7979 ) | ( n7777 & n7980 ) | ( n7979 & n7980 ) ;
  assign n7982 = n7975 & ~n7981 ;
  assign n7985 = ~n7939 & n7984 ;
  assign n7986 = ( n7982 & n7984 ) | ( n7982 & n7985 ) | ( n7984 & n7985 ) ;
  assign n7987 = ( n7982 & n7985 ) | ( n7982 & ~n7986 ) | ( n7985 & ~n7986 ) ;
  assign n7988 = ( n7984 & ~n7986 ) | ( n7984 & n7987 ) | ( ~n7986 & n7987 ) ;
  assign n7989 = n7955 & ~n7988 ;
  assign n7990 = ~n7955 & n7988 ;
  assign n7991 = n7989 | n7990 ;
  assign n7992 = n7922 & n7939 ;
  assign n7993 = n722 | n858 ;
  assign n7994 = n585 | n7993 ;
  assign n7995 = n4810 | n7994 ;
  assign n7996 = n608 | n7995 ;
  assign n7997 = n6704 | n7996 ;
  assign n7998 = n283 | n293 ;
  assign n7999 = n2302 | n7998 ;
  assign n8000 = n165 | n545 ;
  assign n8001 = n689 | n8000 ;
  assign n8002 = n7999 | n8001 ;
  assign n8003 = n134 | n426 ;
  assign n8004 = n8002 | n8003 ;
  assign n8005 = n7997 | n8004 ;
  assign n8006 = n7976 | n8005 ;
  assign n8007 = ( n7899 & n8005 ) | ( n7899 & n8006 ) | ( n8005 & n8006 ) ;
  assign n8008 = n8005 & n8006 ;
  assign n8009 = ( n7850 & n8007 ) | ( n7850 & n8008 ) | ( n8007 & n8008 ) ;
  assign n8010 = n7898 | n8005 ;
  assign n8011 = ( n7976 & n8005 ) | ( n7976 & n8010 ) | ( n8005 & n8010 ) ;
  assign n8012 = ( n7872 & n8009 ) | ( n7872 & n8011 ) | ( n8009 & n8011 ) ;
  assign n8013 = ( n7870 & n8009 ) | ( n7870 & n8011 ) | ( n8009 & n8011 ) ;
  assign n8014 = ( n7777 & n8012 ) | ( n7777 & n8013 ) | ( n8012 & n8013 ) ;
  assign n8015 = ( ~n7939 & n7982 ) | ( ~n7939 & n8014 ) | ( n7982 & n8014 ) ;
  assign n8016 = n7982 | n8014 ;
  assign n8017 = ( ~n7922 & n8015 ) | ( ~n7922 & n8016 ) | ( n8015 & n8016 ) ;
  assign n8018 = n7992 & n8017 ;
  assign n8019 = n7785 & n8018 ;
  assign n8020 = n7976 & n8005 ;
  assign n8021 = n7900 & n8020 ;
  assign n8022 = n7898 & n8020 ;
  assign n8023 = ( n7872 & n8021 ) | ( n7872 & n8022 ) | ( n8021 & n8022 ) ;
  assign n8024 = ( n7870 & n8021 ) | ( n7870 & n8022 ) | ( n8021 & n8022 ) ;
  assign n8025 = ( n7777 & n8023 ) | ( n7777 & n8024 ) | ( n8023 & n8024 ) ;
  assign n8026 = n8014 & ~n8025 ;
  assign n8027 = n7939 & n7982 ;
  assign n8028 = n8026 | n8027 ;
  assign n8029 = ( n7984 & n8026 ) | ( n7984 & n8028 ) | ( n8026 & n8028 ) ;
  assign n8030 = ~n8019 & n8029 ;
  assign n8031 = ~n7950 & n7986 ;
  assign n8032 = n7950 | n7984 ;
  assign n8033 = ( n7987 & ~n8031 ) | ( n7987 & n8032 ) | ( ~n8031 & n8032 ) ;
  assign n8034 = n7919 | n8033 ;
  assign n8035 = n7795 | n8034 ;
  assign n8036 = n5520 & n8035 ;
  assign n8037 = ~n8030 & n8036 ;
  assign n8038 = n8030 & ~n8036 ;
  assign n8039 = n8037 | n8038 ;
  assign n8040 = n900 | n921 ;
  assign n8041 = n339 | n748 ;
  assign n8042 = n743 | n8041 ;
  assign n8043 = n384 | n412 ;
  assign n8044 = n167 | n407 ;
  assign n8045 = n4844 | n8044 ;
  assign n8046 = n1043 | n8045 ;
  assign n8047 = n1034 | n8046 ;
  assign n8048 = n8043 | n8047 ;
  assign n8049 = n8042 | n8048 ;
  assign n8050 = n8040 | n8049 ;
  assign n8051 = n8005 | n8050 ;
  assign n8052 = ( n7976 & n8050 ) | ( n7976 & n8051 ) | ( n8050 & n8051 ) ;
  assign n8053 = ( n7898 & n8050 ) | ( n7898 & n8052 ) | ( n8050 & n8052 ) ;
  assign n8054 = ( n7899 & n8050 ) | ( n7899 & n8052 ) | ( n8050 & n8052 ) ;
  assign n8055 = n8050 & n8052 ;
  assign n8056 = ( n7850 & n8054 ) | ( n7850 & n8055 ) | ( n8054 & n8055 ) ;
  assign n8057 = ( n7872 & n8053 ) | ( n7872 & n8056 ) | ( n8053 & n8056 ) ;
  assign n8058 = ( n7870 & n8053 ) | ( n7870 & n8056 ) | ( n8053 & n8056 ) ;
  assign n8059 = ( n7777 & n8057 ) | ( n7777 & n8058 ) | ( n8057 & n8058 ) ;
  assign n8060 = n8005 & n8050 ;
  assign n8061 = n7976 & n8060 ;
  assign n8062 = n7900 & n8061 ;
  assign n8063 = n7898 & n8061 ;
  assign n8064 = ( n7872 & n8062 ) | ( n7872 & n8063 ) | ( n8062 & n8063 ) ;
  assign n8065 = ( n7870 & n8062 ) | ( n7870 & n8063 ) | ( n8062 & n8063 ) ;
  assign n8066 = ( n7777 & n8064 ) | ( n7777 & n8065 ) | ( n8064 & n8065 ) ;
  assign n8067 = n8059 & ~n8066 ;
  assign n8068 = n8019 | n8067 ;
  assign n8069 = n8019 & n8067 ;
  assign n8070 = n8068 & ~n8069 ;
  assign n8071 = n8030 | n8035 ;
  assign n8072 = n5520 & n8071 ;
  assign n8073 = ~n8070 & n8072 ;
  assign n8074 = n8070 & ~n8072 ;
  assign n8075 = n8073 | n8074 ;
  assign n8076 = n8030 | n8070 ;
  assign n8077 = n7795 | n8076 ;
  assign n8078 = n8034 | n8077 ;
  assign n8079 = n5520 & n8078 ;
  assign n8080 = n1028 | n1035 ;
  assign n8081 = n734 | n8080 ;
  assign n8082 = n1045 | n8081 ;
  assign n8083 = n8061 | n8082 ;
  assign n8084 = ( n7899 & n8082 ) | ( n7899 & n8083 ) | ( n8082 & n8083 ) ;
  assign n8085 = n8082 & n8083 ;
  assign n8086 = ( n7850 & n8084 ) | ( n7850 & n8085 ) | ( n8084 & n8085 ) ;
  assign n8087 = n7898 | n8082 ;
  assign n8088 = ( n8061 & n8082 ) | ( n8061 & n8087 ) | ( n8082 & n8087 ) ;
  assign n8089 = ( n7872 & n8086 ) | ( n7872 & n8088 ) | ( n8086 & n8088 ) ;
  assign n8090 = ( n7870 & n8086 ) | ( n7870 & n8088 ) | ( n8086 & n8088 ) ;
  assign n8091 = ( n7777 & n8089 ) | ( n7777 & n8090 ) | ( n8089 & n8090 ) ;
  assign n8092 = n8061 & n8082 ;
  assign n8093 = n7900 & n8092 ;
  assign n8094 = n7898 & n8092 ;
  assign n8095 = ( n7872 & n8093 ) | ( n7872 & n8094 ) | ( n8093 & n8094 ) ;
  assign n8096 = ( n7870 & n8093 ) | ( n7870 & n8094 ) | ( n8093 & n8094 ) ;
  assign n8097 = ( n7777 & n8095 ) | ( n7777 & n8096 ) | ( n8095 & n8096 ) ;
  assign n8098 = n8091 & ~n8097 ;
  assign n8099 = n8067 | n8098 ;
  assign n8100 = ( n8019 & n8098 ) | ( n8019 & n8099 ) | ( n8098 & n8099 ) ;
  assign n8101 = ~n8091 & n8099 ;
  assign n8102 = ~n8091 & n8098 ;
  assign n8103 = ( n8019 & n8101 ) | ( n8019 & n8102 ) | ( n8101 & n8102 ) ;
  assign n8104 = ( ~n8069 & n8100 ) | ( ~n8069 & n8103 ) | ( n8100 & n8103 ) ;
  assign n8105 = n8079 & ~n8104 ;
  assign n8106 = ~n8079 & n8104 ;
  assign n8107 = n8105 | n8106 ;
  assign n8108 = x22 | n107 ;
  assign n8109 = n5520 & n8104 ;
  assign n8110 = ( n5520 & n8078 ) | ( n5520 & n8109 ) | ( n8078 & n8109 ) ;
  assign n8111 = n8091 | n8097 ;
  assign n8112 = ( n8067 & n8097 ) | ( n8067 & n8111 ) | ( n8097 & n8111 ) ;
  assign n8113 = ( n8019 & n8097 ) | ( n8019 & n8112 ) | ( n8097 & n8112 ) ;
  assign n8114 = ( ~n8067 & n8091 ) | ( ~n8067 & n8097 ) | ( n8091 & n8097 ) ;
  assign n8115 = ( ~n8019 & n8111 ) | ( ~n8019 & n8114 ) | ( n8111 & n8114 ) ;
  assign n8116 = n8069 & n8115 ;
  assign n8117 = n8113 & ~n8116 ;
  assign n8118 = n8109 & n8117 ;
  assign n8119 = n5520 & n8117 ;
  assign n8120 = ( n8078 & n8118 ) | ( n8078 & n8119 ) | ( n8118 & n8119 ) ;
  assign n8121 = n8117 & ~n8119 ;
  assign n8122 = n8117 & ~n8118 ;
  assign n8123 = ( ~n8078 & n8121 ) | ( ~n8078 & n8122 ) | ( n8121 & n8122 ) ;
  assign n8124 = ( n8110 & ~n8120 ) | ( n8110 & n8123 ) | ( ~n8120 & n8123 ) ;
  assign n8125 = n8108 & ~n8124 ;
  assign n8126 = n8076 | n8104 ;
  assign n8127 = n8113 & ~n8126 ;
  assign n8128 = ~n8035 & n8127 ;
  assign n8129 = ~n8116 & n8126 ;
  assign n8130 = ( n8035 & ~n8116 ) | ( n8035 & n8129 ) | ( ~n8116 & n8129 ) ;
  assign n8131 = n8128 | n8130 ;
  assign n8132 = ~x22 & n5520 ;
  assign n8133 = ~n107 & n8132 ;
  assign n8134 = ( n5520 & n8131 ) | ( n5520 & n8133 ) | ( n8131 & n8133 ) ;
  assign y0 = n5271 ;
  assign y1 = n5524 ;
  assign y2 = n5725 ;
  assign y3 = n5927 ;
  assign y4 = n6106 ;
  assign y5 = n6278 ;
  assign y6 = n6491 ;
  assign y7 = n6688 ;
  assign y8 = n6858 ;
  assign y9 = n7008 ;
  assign y10 = n7185 ;
  assign y11 = n7303 ;
  assign y12 = n7452 ;
  assign y13 = n7588 ;
  assign y14 = n7691 ;
  assign y15 = n7793 ;
  assign y16 = n7884 ;
  assign y17 = n7918 ;
  assign y18 = n7953 ;
  assign y19 = n7991 ;
  assign y20 = n8039 ;
  assign y21 = n8075 ;
  assign y22 = n8107 ;
  assign y23 = ~n8125 ;
  assign y24 = n8134 ;
endmodule
