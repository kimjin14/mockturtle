module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 ;
  wire n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 ;
  assign n61 = x17 | x18 ;
  assign n62 = x19 & n61 ;
  assign n63 = x9 | x10 ;
  assign n64 = x11 | x12 ;
  assign n65 = ( x12 & n63 ) | ( x12 & n64 ) | ( n63 & n64 ) ;
  assign n66 = x13 & x14 ;
  assign n67 = x15 & n66 ;
  assign n68 = x14 & x15 ;
  assign n69 = ( n65 & n67 ) | ( n65 & n68 ) | ( n67 & n68 ) ;
  assign n70 = x16 & x17 ;
  assign n71 = x18 & x19 ;
  assign n72 = ( x19 & n70 ) | ( x19 & n71 ) | ( n70 & n71 ) ;
  assign n73 = ( n62 & n69 ) | ( n62 & n72 ) | ( n69 & n72 ) ;
  assign n74 = x20 | x21 ;
  assign n75 = x22 & x23 ;
  assign n76 = ( x23 & n74 ) | ( x23 & n75 ) | ( n74 & n75 ) ;
  assign n77 = x24 & n76 ;
  assign n78 = x25 | x26 ;
  assign n79 = x27 & x28 ;
  assign n80 = n78 & n79 ;
  assign n81 = x29 & n80 ;
  assign n82 = x26 & x27 ;
  assign n83 = x28 & x29 ;
  assign n84 = n82 & n83 ;
  assign n85 = ( n77 & n81 ) | ( n77 & n84 ) | ( n81 & n84 ) ;
  assign n86 = x21 | x22 ;
  assign n87 = x23 & x24 ;
  assign n88 = n86 & n87 ;
  assign n89 = ( n81 & n84 ) | ( n81 & n88 ) | ( n84 & n88 ) ;
  assign n90 = ( n73 & n85 ) | ( n73 & n89 ) | ( n85 & n89 ) ;
  assign n91 = x27 & n78 ;
  assign n92 = ( n77 & n82 ) | ( n77 & n91 ) | ( n82 & n91 ) ;
  assign n93 = ( n82 & n88 ) | ( n82 & n91 ) | ( n88 & n91 ) ;
  assign n94 = ( n73 & n92 ) | ( n73 & n93 ) | ( n92 & n93 ) ;
  assign n95 = x27 | n78 ;
  assign n96 = x26 | x27 ;
  assign n97 = ( n77 & n95 ) | ( n77 & n96 ) | ( n95 & n96 ) ;
  assign n98 = ( n88 & n95 ) | ( n88 & n96 ) | ( n95 & n96 ) ;
  assign n99 = ( n73 & n97 ) | ( n73 & n98 ) | ( n97 & n98 ) ;
  assign n100 = ~n94 & n99 ;
  assign n101 = x28 & ~n82 ;
  assign n102 = ~x27 & x28 ;
  assign n103 = ( x28 & ~n78 ) | ( x28 & n102 ) | ( ~n78 & n102 ) ;
  assign n104 = ( ~n77 & n101 ) | ( ~n77 & n103 ) | ( n101 & n103 ) ;
  assign n105 = ( ~n88 & n101 ) | ( ~n88 & n103 ) | ( n101 & n103 ) ;
  assign n106 = ( ~n73 & n104 ) | ( ~n73 & n105 ) | ( n104 & n105 ) ;
  assign n107 = ~x28 & n82 ;
  assign n108 = x27 & ~x28 ;
  assign n109 = n78 & n108 ;
  assign n110 = ( n77 & n107 ) | ( n77 & n109 ) | ( n107 & n109 ) ;
  assign n111 = ( n88 & n107 ) | ( n88 & n109 ) | ( n107 & n109 ) ;
  assign n112 = ( n73 & n110 ) | ( n73 & n111 ) | ( n110 & n111 ) ;
  assign n113 = n106 | n112 ;
  assign n114 = n100 | n113 ;
  assign n115 = ~x9 & n90 ;
  assign n116 = ( n90 & n114 ) | ( n90 & n115 ) | ( n114 & n115 ) ;
  assign n117 = x1 | x2 ;
  assign n118 = x3 | x4 ;
  assign n119 = n117 | n118 ;
  assign n120 = x5 | x6 ;
  assign n121 = x7 | n120 ;
  assign n122 = n119 | n121 ;
  assign n123 = x9 & x10 ;
  assign n124 = n63 & ~n123 ;
  assign n125 = ~x8 & n124 ;
  assign n126 = ~n122 & n125 ;
  assign n127 = x11 & n63 ;
  assign n128 = x11 | n63 ;
  assign n129 = ~n127 & n128 ;
  assign n130 = x11 & x12 ;
  assign n131 = n63 & n130 ;
  assign n132 = n65 & ~n131 ;
  assign n133 = ~n129 & n132 ;
  assign n134 = n126 & n133 ;
  assign n135 = x13 | n65 ;
  assign n136 = x13 & n65 ;
  assign n137 = n135 & ~n136 ;
  assign n138 = x13 | x14 ;
  assign n139 = n65 | n138 ;
  assign n140 = ~x14 & n138 ;
  assign n141 = ( ~x14 & n65 ) | ( ~x14 & n140 ) | ( n65 & n140 ) ;
  assign n142 = ( ~n135 & n139 ) | ( ~n135 & n141 ) | ( n139 & n141 ) ;
  assign n143 = n137 & ~n142 ;
  assign n144 = n134 & n143 ;
  assign n145 = x16 | n69 ;
  assign n146 = x16 & n69 ;
  assign n147 = n145 & ~n146 ;
  assign n148 = ( x14 & n65 ) | ( x14 & n66 ) | ( n65 & n66 ) ;
  assign n149 = x15 & ~n69 ;
  assign n150 = ( ~n69 & n148 ) | ( ~n69 & n149 ) | ( n148 & n149 ) ;
  assign n151 = n147 & ~n150 ;
  assign n152 = n144 & n151 ;
  assign n153 = x19 | n61 ;
  assign n154 = x18 | x19 ;
  assign n155 = n70 | n154 ;
  assign n156 = ( n69 & n153 ) | ( n69 & n155 ) | ( n153 & n155 ) ;
  assign n157 = ~n73 & n156 ;
  assign n158 = x18 | n70 ;
  assign n159 = ( n61 & n69 ) | ( n61 & n158 ) | ( n69 & n158 ) ;
  assign n160 = x18 & n70 ;
  assign n161 = x17 & x18 ;
  assign n162 = ( n69 & n160 ) | ( n69 & n161 ) | ( n160 & n161 ) ;
  assign n163 = n159 & ~n162 ;
  assign n164 = x16 | x17 ;
  assign n165 = n69 | n164 ;
  assign n166 = ~x17 & n164 ;
  assign n167 = ( ~x17 & n69 ) | ( ~x17 & n166 ) | ( n69 & n166 ) ;
  assign n168 = ( ~n145 & n165 ) | ( ~n145 & n167 ) | ( n165 & n167 ) ;
  assign n169 = n163 & ~n168 ;
  assign n170 = ~n157 & n169 ;
  assign n171 = n152 & n170 ;
  assign n172 = x20 & n72 ;
  assign n173 = x20 & n62 ;
  assign n174 = ( n69 & n172 ) | ( n69 & n173 ) | ( n172 & n173 ) ;
  assign n175 = x20 & ~n174 ;
  assign n176 = ( n73 & ~n174 ) | ( n73 & n175 ) | ( ~n174 & n175 ) ;
  assign n177 = x22 | n74 ;
  assign n178 = ( n72 & n86 ) | ( n72 & n177 ) | ( n86 & n177 ) ;
  assign n179 = ( n62 & n86 ) | ( n62 & n177 ) | ( n86 & n177 ) ;
  assign n180 = ( n69 & n178 ) | ( n69 & n179 ) | ( n178 & n179 ) ;
  assign n181 = x22 & n74 ;
  assign n182 = x21 & x22 ;
  assign n183 = ( n72 & n181 ) | ( n72 & n182 ) | ( n181 & n182 ) ;
  assign n184 = ( n62 & n181 ) | ( n62 & n182 ) | ( n181 & n182 ) ;
  assign n185 = ( n69 & n183 ) | ( n69 & n184 ) | ( n183 & n184 ) ;
  assign n186 = n180 & ~n185 ;
  assign n187 = ( x21 & n72 ) | ( x21 & n74 ) | ( n72 & n74 ) ;
  assign n188 = ( x21 & n62 ) | ( x21 & n74 ) | ( n62 & n74 ) ;
  assign n189 = ( n69 & n187 ) | ( n69 & n188 ) | ( n187 & n188 ) ;
  assign n190 = x20 & x21 ;
  assign n191 = n72 & n190 ;
  assign n192 = n62 & n190 ;
  assign n193 = ( n69 & n191 ) | ( n69 & n192 ) | ( n191 & n192 ) ;
  assign n194 = n189 & ~n193 ;
  assign n195 = n186 & n194 ;
  assign n196 = ~n176 & n195 ;
  assign n197 = n171 & n196 ;
  assign n198 = x23 & n86 ;
  assign n199 = ( n72 & n76 ) | ( n72 & n198 ) | ( n76 & n198 ) ;
  assign n200 = ( n62 & n76 ) | ( n62 & n198 ) | ( n76 & n198 ) ;
  assign n201 = ( n69 & n199 ) | ( n69 & n200 ) | ( n199 & n200 ) ;
  assign n202 = x23 | n86 ;
  assign n203 = x22 | x23 ;
  assign n204 = n74 | n203 ;
  assign n205 = ( n72 & n202 ) | ( n72 & n204 ) | ( n202 & n204 ) ;
  assign n206 = ( n62 & n202 ) | ( n62 & n204 ) | ( n202 & n204 ) ;
  assign n207 = ( n69 & n205 ) | ( n69 & n206 ) | ( n205 & n206 ) ;
  assign n208 = ~n201 & n207 ;
  assign n209 = x24 & ~n76 ;
  assign n210 = ~x23 & x24 ;
  assign n211 = ( x24 & ~n86 ) | ( x24 & n210 ) | ( ~n86 & n210 ) ;
  assign n212 = ( ~n73 & n209 ) | ( ~n73 & n211 ) | ( n209 & n211 ) ;
  assign n213 = ~x24 & n76 ;
  assign n214 = x23 & ~x24 ;
  assign n215 = n86 & n214 ;
  assign n216 = ( n73 & n213 ) | ( n73 & n215 ) | ( n213 & n215 ) ;
  assign n217 = n212 | n216 ;
  assign n218 = n208 | n217 ;
  assign n219 = ( x26 & n78 ) | ( x26 & n88 ) | ( n78 & n88 ) ;
  assign n220 = ( x24 & x26 ) | ( x24 & n78 ) | ( x26 & n78 ) ;
  assign n221 = x26 & n78 ;
  assign n222 = ( n76 & n220 ) | ( n76 & n221 ) | ( n220 & n221 ) ;
  assign n223 = ( n73 & n219 ) | ( n73 & n222 ) | ( n219 & n222 ) ;
  assign n224 = x25 & x26 ;
  assign n225 = n77 & n224 ;
  assign n226 = n88 & n224 ;
  assign n227 = ( n73 & n225 ) | ( n73 & n226 ) | ( n225 & n226 ) ;
  assign n228 = n223 & ~n227 ;
  assign n229 = ( n73 & n77 ) | ( n73 & n88 ) | ( n77 & n88 ) ;
  assign n230 = x25 & n77 ;
  assign n231 = x25 & n88 ;
  assign n232 = ( n73 & n230 ) | ( n73 & n231 ) | ( n230 & n231 ) ;
  assign n233 = x25 & ~n232 ;
  assign n234 = ( n229 & ~n232 ) | ( n229 & n233 ) | ( ~n232 & n233 ) ;
  assign n235 = n228 & ~n234 ;
  assign n236 = ~n218 & n235 ;
  assign n237 = ( n116 & n197 ) | ( n116 & n236 ) | ( n197 & n236 ) ;
  assign n238 = ( n90 & n116 ) | ( n90 & ~n237 ) | ( n116 & ~n237 ) ;
  assign n239 = ~x29 & n80 ;
  assign n240 = x28 & ~x29 ;
  assign n241 = n82 & n240 ;
  assign n242 = ( n77 & n239 ) | ( n77 & n241 ) | ( n239 & n241 ) ;
  assign n243 = ( n88 & n239 ) | ( n88 & n241 ) | ( n239 & n241 ) ;
  assign n244 = ( n73 & n242 ) | ( n73 & n243 ) | ( n242 & n243 ) ;
  assign n245 = x29 & ~n80 ;
  assign n246 = ~x28 & x29 ;
  assign n247 = ( x29 & ~n82 ) | ( x29 & n246 ) | ( ~n82 & n246 ) ;
  assign n248 = ( ~n77 & n245 ) | ( ~n77 & n247 ) | ( n245 & n247 ) ;
  assign n249 = ( ~n88 & n245 ) | ( ~n88 & n247 ) | ( n245 & n247 ) ;
  assign n250 = ( ~n73 & n248 ) | ( ~n73 & n249 ) | ( n248 & n249 ) ;
  assign n251 = n244 | n250 ;
  assign n252 = ~x9 & n251 ;
  assign n253 = n100 & n113 ;
  assign n254 = n252 & n253 ;
  assign n255 = n217 & ~n228 ;
  assign n256 = n234 & n255 ;
  assign n257 = n254 & n256 ;
  assign n258 = ~n163 & n168 ;
  assign n259 = ~n147 & n150 ;
  assign n260 = n258 & n259 ;
  assign n261 = ~n137 & n142 ;
  assign n262 = ~n132 & n261 ;
  assign n263 = n260 & n262 ;
  assign n264 = n176 & ~n194 ;
  assign n265 = ~n186 & n208 ;
  assign n266 = n157 & n265 ;
  assign n267 = n264 & n266 ;
  assign n268 = n263 & n267 ;
  assign n269 = n257 & n268 ;
  assign n270 = x0 | n90 ;
  assign n271 = x8 & ~n124 ;
  assign n272 = n129 & n271 ;
  assign n273 = x6 & x7 ;
  assign n274 = x4 & x5 ;
  assign n275 = n273 & n274 ;
  assign n276 = x3 & n275 ;
  assign n277 = x1 & x2 ;
  assign n278 = n276 & n277 ;
  assign n279 = n272 & n278 ;
  assign n280 = ( n90 & n270 ) | ( n90 & n279 ) | ( n270 & n279 ) ;
  assign n281 = ( n90 & n269 ) | ( n90 & n280 ) | ( n269 & n280 ) ;
  assign n282 = ~n238 & n281 ;
  assign n283 = x47 | x48 ;
  assign n284 = x49 & n283 ;
  assign n285 = x39 | x40 ;
  assign n286 = x41 | x42 ;
  assign n287 = ( x42 & n285 ) | ( x42 & n286 ) | ( n285 & n286 ) ;
  assign n288 = x43 & x44 ;
  assign n289 = x45 & n288 ;
  assign n290 = x44 & x45 ;
  assign n291 = ( n287 & n289 ) | ( n287 & n290 ) | ( n289 & n290 ) ;
  assign n292 = x46 & x47 ;
  assign n293 = x48 & x49 ;
  assign n294 = ( x49 & n292 ) | ( x49 & n293 ) | ( n292 & n293 ) ;
  assign n295 = ( n284 & n291 ) | ( n284 & n294 ) | ( n291 & n294 ) ;
  assign n296 = x50 | x51 ;
  assign n297 = x52 & x53 ;
  assign n298 = ( x53 & n296 ) | ( x53 & n297 ) | ( n296 & n297 ) ;
  assign n299 = x54 & n298 ;
  assign n300 = x55 | x56 ;
  assign n301 = x57 & x58 ;
  assign n302 = n300 & n301 ;
  assign n303 = x59 & n302 ;
  assign n304 = x56 & x57 ;
  assign n305 = x58 & x59 ;
  assign n306 = n304 & n305 ;
  assign n307 = ( n299 & n303 ) | ( n299 & n306 ) | ( n303 & n306 ) ;
  assign n308 = x51 | x52 ;
  assign n309 = x53 & x54 ;
  assign n310 = n308 & n309 ;
  assign n311 = ( n303 & n306 ) | ( n303 & n310 ) | ( n306 & n310 ) ;
  assign n312 = ( n295 & n307 ) | ( n295 & n311 ) | ( n307 & n311 ) ;
  assign n313 = x0 & ~n312 ;
  assign n314 = ~n116 & n313 ;
  assign n315 = ~n90 & n313 ;
  assign n316 = ( n237 & n314 ) | ( n237 & n315 ) | ( n314 & n315 ) ;
  assign n317 = x58 & ~n304 ;
  assign n318 = ~x57 & x58 ;
  assign n319 = ( x58 & ~n300 ) | ( x58 & n318 ) | ( ~n300 & n318 ) ;
  assign n320 = ( ~n299 & n317 ) | ( ~n299 & n319 ) | ( n317 & n319 ) ;
  assign n321 = ( ~n310 & n317 ) | ( ~n310 & n319 ) | ( n317 & n319 ) ;
  assign n322 = ( ~n295 & n320 ) | ( ~n295 & n321 ) | ( n320 & n321 ) ;
  assign n323 = ~x58 & n304 ;
  assign n324 = x57 & ~x58 ;
  assign n325 = n300 & n324 ;
  assign n326 = ( n299 & n323 ) | ( n299 & n325 ) | ( n323 & n325 ) ;
  assign n327 = ( n310 & n323 ) | ( n310 & n325 ) | ( n323 & n325 ) ;
  assign n328 = ( n295 & n326 ) | ( n295 & n327 ) | ( n326 & n327 ) ;
  assign n329 = n322 | n328 ;
  assign n330 = x57 & n300 ;
  assign n331 = ( n299 & n304 ) | ( n299 & n330 ) | ( n304 & n330 ) ;
  assign n332 = ( n304 & n310 ) | ( n304 & n330 ) | ( n310 & n330 ) ;
  assign n333 = ( n295 & n331 ) | ( n295 & n332 ) | ( n331 & n332 ) ;
  assign n334 = x57 | n300 ;
  assign n335 = x56 | x57 ;
  assign n336 = ( n299 & n334 ) | ( n299 & n335 ) | ( n334 & n335 ) ;
  assign n337 = ( n310 & n334 ) | ( n310 & n335 ) | ( n334 & n335 ) ;
  assign n338 = ( n295 & n336 ) | ( n295 & n337 ) | ( n336 & n337 ) ;
  assign n339 = ~n333 & n338 ;
  assign n340 = n329 | n339 ;
  assign n341 = ~x39 & n312 ;
  assign n342 = ( n312 & n340 ) | ( n312 & n341 ) | ( n340 & n341 ) ;
  assign n343 = x31 | x32 ;
  assign n344 = x33 | x34 ;
  assign n345 = n343 | n344 ;
  assign n346 = x35 | x36 ;
  assign n347 = x37 | n346 ;
  assign n348 = n345 | n347 ;
  assign n349 = x39 & x40 ;
  assign n350 = n285 & ~n349 ;
  assign n351 = ~x38 & n350 ;
  assign n352 = ~n348 & n351 ;
  assign n353 = x41 & n285 ;
  assign n354 = x41 | n285 ;
  assign n355 = ~n353 & n354 ;
  assign n356 = x41 & x42 ;
  assign n357 = n285 & n356 ;
  assign n358 = n287 & ~n357 ;
  assign n359 = ~n355 & n358 ;
  assign n360 = n352 & n359 ;
  assign n361 = x43 | n287 ;
  assign n362 = x43 & n287 ;
  assign n363 = n361 & ~n362 ;
  assign n364 = x43 | x44 ;
  assign n365 = n287 | n364 ;
  assign n366 = ~x44 & n364 ;
  assign n367 = ( ~x44 & n287 ) | ( ~x44 & n366 ) | ( n287 & n366 ) ;
  assign n368 = ( ~n361 & n365 ) | ( ~n361 & n367 ) | ( n365 & n367 ) ;
  assign n369 = n363 & ~n368 ;
  assign n370 = n360 & n369 ;
  assign n371 = x46 | n291 ;
  assign n372 = x46 & n291 ;
  assign n373 = n371 & ~n372 ;
  assign n374 = ( x44 & n287 ) | ( x44 & n288 ) | ( n287 & n288 ) ;
  assign n375 = x45 & ~n291 ;
  assign n376 = ( ~n291 & n374 ) | ( ~n291 & n375 ) | ( n374 & n375 ) ;
  assign n377 = n373 & ~n376 ;
  assign n378 = n370 & n377 ;
  assign n379 = x49 | n283 ;
  assign n380 = x48 | x49 ;
  assign n381 = n292 | n380 ;
  assign n382 = ( n291 & n379 ) | ( n291 & n381 ) | ( n379 & n381 ) ;
  assign n383 = ~n295 & n382 ;
  assign n384 = x48 | n292 ;
  assign n385 = ( n283 & n291 ) | ( n283 & n384 ) | ( n291 & n384 ) ;
  assign n386 = x48 & n292 ;
  assign n387 = x47 & x48 ;
  assign n388 = ( n291 & n386 ) | ( n291 & n387 ) | ( n386 & n387 ) ;
  assign n389 = n385 & ~n388 ;
  assign n390 = x46 | x47 ;
  assign n391 = n291 | n390 ;
  assign n392 = ~x47 & n390 ;
  assign n393 = ( ~x47 & n291 ) | ( ~x47 & n392 ) | ( n291 & n392 ) ;
  assign n394 = ( ~n371 & n391 ) | ( ~n371 & n393 ) | ( n391 & n393 ) ;
  assign n395 = n389 & ~n394 ;
  assign n396 = ~n383 & n395 ;
  assign n397 = n378 & n396 ;
  assign n398 = x50 & n294 ;
  assign n399 = x50 & n284 ;
  assign n400 = ( n291 & n398 ) | ( n291 & n399 ) | ( n398 & n399 ) ;
  assign n401 = x50 & ~n400 ;
  assign n402 = ( n295 & ~n400 ) | ( n295 & n401 ) | ( ~n400 & n401 ) ;
  assign n403 = ( x51 & n294 ) | ( x51 & n296 ) | ( n294 & n296 ) ;
  assign n404 = ( x51 & n284 ) | ( x51 & n296 ) | ( n284 & n296 ) ;
  assign n405 = ( n291 & n403 ) | ( n291 & n404 ) | ( n403 & n404 ) ;
  assign n406 = x50 & x51 ;
  assign n407 = n294 & n406 ;
  assign n408 = n284 & n406 ;
  assign n409 = ( n291 & n407 ) | ( n291 & n408 ) | ( n407 & n408 ) ;
  assign n410 = n405 & ~n409 ;
  assign n411 = x52 | n296 ;
  assign n412 = ( n294 & n308 ) | ( n294 & n411 ) | ( n308 & n411 ) ;
  assign n413 = ( n284 & n308 ) | ( n284 & n411 ) | ( n308 & n411 ) ;
  assign n414 = ( n291 & n412 ) | ( n291 & n413 ) | ( n412 & n413 ) ;
  assign n415 = x52 & n296 ;
  assign n416 = x51 & x52 ;
  assign n417 = ( n294 & n415 ) | ( n294 & n416 ) | ( n415 & n416 ) ;
  assign n418 = ( n284 & n415 ) | ( n284 & n416 ) | ( n415 & n416 ) ;
  assign n419 = ( n291 & n417 ) | ( n291 & n418 ) | ( n417 & n418 ) ;
  assign n420 = n414 & ~n419 ;
  assign n421 = n410 & n420 ;
  assign n422 = ~n402 & n421 ;
  assign n423 = n397 & n422 ;
  assign n424 = x53 & n308 ;
  assign n425 = ( n294 & n298 ) | ( n294 & n424 ) | ( n298 & n424 ) ;
  assign n426 = ( n284 & n298 ) | ( n284 & n424 ) | ( n298 & n424 ) ;
  assign n427 = ( n291 & n425 ) | ( n291 & n426 ) | ( n425 & n426 ) ;
  assign n428 = x53 | n308 ;
  assign n429 = x52 | x53 ;
  assign n430 = n296 | n429 ;
  assign n431 = ( n294 & n428 ) | ( n294 & n430 ) | ( n428 & n430 ) ;
  assign n432 = ( n284 & n428 ) | ( n284 & n430 ) | ( n428 & n430 ) ;
  assign n433 = ( n291 & n431 ) | ( n291 & n432 ) | ( n431 & n432 ) ;
  assign n434 = ~n427 & n433 ;
  assign n435 = x54 & ~n298 ;
  assign n436 = ~x53 & x54 ;
  assign n437 = ( x54 & ~n308 ) | ( x54 & n436 ) | ( ~n308 & n436 ) ;
  assign n438 = ( ~n295 & n435 ) | ( ~n295 & n437 ) | ( n435 & n437 ) ;
  assign n439 = ~x54 & n298 ;
  assign n440 = x53 & ~x54 ;
  assign n441 = n308 & n440 ;
  assign n442 = ( n295 & n439 ) | ( n295 & n441 ) | ( n439 & n441 ) ;
  assign n443 = n438 | n442 ;
  assign n444 = n434 | n443 ;
  assign n445 = ( x56 & n300 ) | ( x56 & n310 ) | ( n300 & n310 ) ;
  assign n446 = ( x54 & x56 ) | ( x54 & n300 ) | ( x56 & n300 ) ;
  assign n447 = x56 & n300 ;
  assign n448 = ( n298 & n446 ) | ( n298 & n447 ) | ( n446 & n447 ) ;
  assign n449 = ( n295 & n445 ) | ( n295 & n448 ) | ( n445 & n448 ) ;
  assign n450 = x55 & x56 ;
  assign n451 = n299 & n450 ;
  assign n452 = n310 & n450 ;
  assign n453 = ( n295 & n451 ) | ( n295 & n452 ) | ( n451 & n452 ) ;
  assign n454 = n449 & ~n453 ;
  assign n455 = ( n295 & n299 ) | ( n295 & n310 ) | ( n299 & n310 ) ;
  assign n456 = x55 & n299 ;
  assign n457 = x55 & n310 ;
  assign n458 = ( n295 & n456 ) | ( n295 & n457 ) | ( n456 & n457 ) ;
  assign n459 = x55 & ~n458 ;
  assign n460 = ( n455 & ~n458 ) | ( n455 & n459 ) | ( ~n458 & n459 ) ;
  assign n461 = n454 & ~n460 ;
  assign n462 = ~n444 & n461 ;
  assign n463 = ( n342 & n423 ) | ( n342 & n462 ) | ( n423 & n462 ) ;
  assign n464 = ( n312 & n342 ) | ( n312 & ~n463 ) | ( n342 & ~n463 ) ;
  assign n465 = x30 & ~x39 ;
  assign n466 = x59 & n465 ;
  assign n467 = n329 & n466 ;
  assign n468 = n339 & ~n454 ;
  assign n469 = n467 & n468 ;
  assign n470 = n434 & n443 ;
  assign n471 = n460 & n470 ;
  assign n472 = n469 & n471 ;
  assign n473 = n410 | n420 ;
  assign n474 = n402 & ~n473 ;
  assign n475 = n383 & ~n389 ;
  assign n476 = n474 & n475 ;
  assign n477 = ~n373 & n394 ;
  assign n478 = n368 & n376 ;
  assign n479 = n477 & n478 ;
  assign n480 = n358 | n363 ;
  assign n481 = n355 & ~n480 ;
  assign n482 = n479 & n481 ;
  assign n483 = n476 & n482 ;
  assign n484 = n472 & n483 ;
  assign n485 = x37 & x38 ;
  assign n486 = x36 & n485 ;
  assign n487 = ~n350 & n486 ;
  assign n488 = x34 & x35 ;
  assign n489 = x33 & n488 ;
  assign n490 = x32 & n489 ;
  assign n491 = n487 & n490 ;
  assign n492 = x31 & n491 ;
  assign n493 = n342 | n492 ;
  assign n494 = n312 | n492 ;
  assign n495 = ( ~n463 & n493 ) | ( ~n463 & n494 ) | ( n493 & n494 ) ;
  assign n496 = ( n464 & n484 ) | ( n464 & n495 ) | ( n484 & n495 ) ;
  assign n497 = x0 | x30 ;
  assign n498 = n312 & n497 ;
  assign n499 = n281 & n498 ;
  assign n500 = ( n281 & n496 ) | ( n281 & n499 ) | ( n496 & n499 ) ;
  assign n501 = ( n238 & ~n316 ) | ( n238 & n500 ) | ( ~n316 & n500 ) ;
  assign n502 = x0 & x30 ;
  assign n503 = n312 & n502 ;
  assign n504 = n464 | n503 ;
  assign n505 = n282 & n504 ;
  assign y0 = ~n282 ;
  assign y1 = ~n501 ;
  assign y2 = n505 ;
  assign y3 = 1'b0 ;
  assign y4 = 1'b0 ;
  assign y5 = 1'b0 ;
  assign y6 = 1'b0 ;
  assign y7 = 1'b0 ;
  assign y8 = 1'b0 ;
  assign y9 = 1'b0 ;
  assign y10 = 1'b0 ;
  assign y11 = 1'b0 ;
  assign y12 = 1'b0 ;
  assign y13 = 1'b0 ;
  assign y14 = 1'b0 ;
  assign y15 = 1'b0 ;
  assign y16 = 1'b0 ;
  assign y17 = 1'b0 ;
  assign y18 = 1'b0 ;
  assign y19 = 1'b0 ;
  assign y20 = 1'b0 ;
  assign y21 = 1'b0 ;
  assign y22 = 1'b0 ;
  assign y23 = 1'b0 ;
  assign y24 = 1'b0 ;
  assign y25 = 1'b0 ;
  assign y26 = 1'b0 ;
  assign y27 = 1'b0 ;
  assign y28 = 1'b0 ;
  assign y29 = 1'b0 ;
endmodule
