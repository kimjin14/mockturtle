module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 , x147 , x148 , x149 , x150 , x151 , x152 , x153 , x154 , x155 , x156 , x157 , x158 , x159 , x160 , x161 , x162 , x163 , x164 , x165 , x166 , x167 , x168 , x169 , x170 , x171 , x172 , x173 , x174 , x175 , x176 , x177 , x178 , x179 , x180 , x181 , x182 , x183 , x184 , x185 , x186 , x187 , x188 , x189 , x190 , x191 , x192 , x193 , x194 , x195 , x196 , x197 , x198 , x199 , x200 , x201 , x202 , x203 , x204 , x205 , x206 , x207 , x208 , x209 , x210 , x211 , x212 , x213 , x214 , x215 , x216 , x217 , x218 , x219 , x220 , x221 , x222 , x223 , x224 , x225 , x226 , x227 , x228 , x229 , x230 , x231 , x232 , x233 , x234 , x235 , x236 , x237 , x238 , x239 , x240 , x241 , x242 , x243 , x244 , x245 , x246 , x247 , x248 , x249 , x250 , x251 , x252 , x253 , x254 , x255 , x256 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 , y128 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 , x147 , x148 , x149 , x150 , x151 , x152 , x153 , x154 , x155 , x156 , x157 , x158 , x159 , x160 , x161 , x162 , x163 , x164 , x165 , x166 , x167 , x168 , x169 , x170 , x171 , x172 , x173 , x174 , x175 , x176 , x177 , x178 , x179 , x180 , x181 , x182 , x183 , x184 , x185 , x186 , x187 , x188 , x189 , x190 , x191 , x192 , x193 , x194 , x195 , x196 , x197 , x198 , x199 , x200 , x201 , x202 , x203 , x204 , x205 , x206 , x207 , x208 , x209 , x210 , x211 , x212 , x213 , x214 , x215 , x216 , x217 , x218 , x219 , x220 , x221 , x222 , x223 , x224 , x225 , x226 , x227 , x228 , x229 , x230 , x231 , x232 , x233 , x234 , x235 , x236 , x237 , x238 , x239 , x240 , x241 , x242 , x243 , x244 , x245 , x246 , x247 , x248 , x249 , x250 , x251 , x252 , x253 , x254 , x255 , x256 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 , y128 ;
  wire n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 ;
  assign n258 = ( x0 & ~x1 ) | ( x0 & x2 ) | ( ~x1 & x2 ) ;
  assign n259 = ( ~x0 & x1 ) | ( ~x0 & n258 ) | ( x1 & n258 ) ;
  assign n260 = ( ~x2 & n258 ) | ( ~x2 & n259 ) | ( n258 & n259 ) ;
  assign n261 = ( x0 & x1 ) | ( x0 & x2 ) | ( x1 & x2 ) ;
  assign n262 = ( x3 & ~x4 ) | ( x3 & n261 ) | ( ~x4 & n261 ) ;
  assign n263 = ( ~x3 & x4 ) | ( ~x3 & n262 ) | ( x4 & n262 ) ;
  assign n264 = ( ~n261 & n262 ) | ( ~n261 & n263 ) | ( n262 & n263 ) ;
  assign n265 = ( x3 & x4 ) | ( x3 & n261 ) | ( x4 & n261 ) ;
  assign n266 = ( x5 & ~x6 ) | ( x5 & n265 ) | ( ~x6 & n265 ) ;
  assign n267 = ( ~x5 & x6 ) | ( ~x5 & n266 ) | ( x6 & n266 ) ;
  assign n268 = ( ~n265 & n266 ) | ( ~n265 & n267 ) | ( n266 & n267 ) ;
  assign n269 = ( x5 & x6 ) | ( x5 & n265 ) | ( x6 & n265 ) ;
  assign n270 = ( x7 & ~x8 ) | ( x7 & n269 ) | ( ~x8 & n269 ) ;
  assign n271 = ( ~x7 & x8 ) | ( ~x7 & n270 ) | ( x8 & n270 ) ;
  assign n272 = ( ~n269 & n270 ) | ( ~n269 & n271 ) | ( n270 & n271 ) ;
  assign n273 = ( x7 & x8 ) | ( x7 & n269 ) | ( x8 & n269 ) ;
  assign n274 = ( x9 & ~x10 ) | ( x9 & n273 ) | ( ~x10 & n273 ) ;
  assign n275 = ( ~x9 & x10 ) | ( ~x9 & n274 ) | ( x10 & n274 ) ;
  assign n276 = ( ~n273 & n274 ) | ( ~n273 & n275 ) | ( n274 & n275 ) ;
  assign n277 = ( x9 & x10 ) | ( x9 & n273 ) | ( x10 & n273 ) ;
  assign n278 = ( x11 & ~x12 ) | ( x11 & n277 ) | ( ~x12 & n277 ) ;
  assign n279 = ( ~x11 & x12 ) | ( ~x11 & n278 ) | ( x12 & n278 ) ;
  assign n280 = ( ~n277 & n278 ) | ( ~n277 & n279 ) | ( n278 & n279 ) ;
  assign n281 = ( x11 & x12 ) | ( x11 & n277 ) | ( x12 & n277 ) ;
  assign n282 = ( x13 & ~x14 ) | ( x13 & n281 ) | ( ~x14 & n281 ) ;
  assign n283 = ( ~x13 & x14 ) | ( ~x13 & n282 ) | ( x14 & n282 ) ;
  assign n284 = ( ~n281 & n282 ) | ( ~n281 & n283 ) | ( n282 & n283 ) ;
  assign n285 = ( x13 & x14 ) | ( x13 & n281 ) | ( x14 & n281 ) ;
  assign n286 = ( x15 & ~x16 ) | ( x15 & n285 ) | ( ~x16 & n285 ) ;
  assign n287 = ( ~x15 & x16 ) | ( ~x15 & n286 ) | ( x16 & n286 ) ;
  assign n288 = ( ~n285 & n286 ) | ( ~n285 & n287 ) | ( n286 & n287 ) ;
  assign n289 = ( x15 & x16 ) | ( x15 & n285 ) | ( x16 & n285 ) ;
  assign n290 = ( x17 & ~x18 ) | ( x17 & n289 ) | ( ~x18 & n289 ) ;
  assign n291 = ( ~x17 & x18 ) | ( ~x17 & n290 ) | ( x18 & n290 ) ;
  assign n292 = ( ~n289 & n290 ) | ( ~n289 & n291 ) | ( n290 & n291 ) ;
  assign n293 = ( x17 & x18 ) | ( x17 & n289 ) | ( x18 & n289 ) ;
  assign n294 = ( x19 & ~x20 ) | ( x19 & n293 ) | ( ~x20 & n293 ) ;
  assign n295 = ( ~x19 & x20 ) | ( ~x19 & n294 ) | ( x20 & n294 ) ;
  assign n296 = ( ~n293 & n294 ) | ( ~n293 & n295 ) | ( n294 & n295 ) ;
  assign n297 = ( x19 & x20 ) | ( x19 & n293 ) | ( x20 & n293 ) ;
  assign n298 = ( x21 & ~x22 ) | ( x21 & n297 ) | ( ~x22 & n297 ) ;
  assign n299 = ( ~x21 & x22 ) | ( ~x21 & n298 ) | ( x22 & n298 ) ;
  assign n300 = ( ~n297 & n298 ) | ( ~n297 & n299 ) | ( n298 & n299 ) ;
  assign n301 = ( x21 & x22 ) | ( x21 & n297 ) | ( x22 & n297 ) ;
  assign n302 = ( x23 & ~x24 ) | ( x23 & n301 ) | ( ~x24 & n301 ) ;
  assign n303 = ( ~x23 & x24 ) | ( ~x23 & n302 ) | ( x24 & n302 ) ;
  assign n304 = ( ~n301 & n302 ) | ( ~n301 & n303 ) | ( n302 & n303 ) ;
  assign n305 = ( x23 & x24 ) | ( x23 & n301 ) | ( x24 & n301 ) ;
  assign n306 = ( x25 & ~x26 ) | ( x25 & n305 ) | ( ~x26 & n305 ) ;
  assign n307 = ( ~x25 & x26 ) | ( ~x25 & n306 ) | ( x26 & n306 ) ;
  assign n308 = ( ~n305 & n306 ) | ( ~n305 & n307 ) | ( n306 & n307 ) ;
  assign n309 = ( x25 & x26 ) | ( x25 & n305 ) | ( x26 & n305 ) ;
  assign n310 = ( x27 & ~x28 ) | ( x27 & n309 ) | ( ~x28 & n309 ) ;
  assign n311 = ( ~x27 & x28 ) | ( ~x27 & n310 ) | ( x28 & n310 ) ;
  assign n312 = ( ~n309 & n310 ) | ( ~n309 & n311 ) | ( n310 & n311 ) ;
  assign n313 = ( x27 & x28 ) | ( x27 & n309 ) | ( x28 & n309 ) ;
  assign n314 = ( x29 & ~x30 ) | ( x29 & n313 ) | ( ~x30 & n313 ) ;
  assign n315 = ( ~x29 & x30 ) | ( ~x29 & n314 ) | ( x30 & n314 ) ;
  assign n316 = ( ~n313 & n314 ) | ( ~n313 & n315 ) | ( n314 & n315 ) ;
  assign n317 = ( x29 & x30 ) | ( x29 & n313 ) | ( x30 & n313 ) ;
  assign n318 = ( x31 & ~x32 ) | ( x31 & n317 ) | ( ~x32 & n317 ) ;
  assign n319 = ( ~x31 & x32 ) | ( ~x31 & n318 ) | ( x32 & n318 ) ;
  assign n320 = ( ~n317 & n318 ) | ( ~n317 & n319 ) | ( n318 & n319 ) ;
  assign n321 = ( x31 & x32 ) | ( x31 & n317 ) | ( x32 & n317 ) ;
  assign n322 = ( x33 & ~x34 ) | ( x33 & n321 ) | ( ~x34 & n321 ) ;
  assign n323 = ( ~x33 & x34 ) | ( ~x33 & n322 ) | ( x34 & n322 ) ;
  assign n324 = ( ~n321 & n322 ) | ( ~n321 & n323 ) | ( n322 & n323 ) ;
  assign n325 = ( x33 & x34 ) | ( x33 & n321 ) | ( x34 & n321 ) ;
  assign n326 = ( x35 & ~x36 ) | ( x35 & n325 ) | ( ~x36 & n325 ) ;
  assign n327 = ( ~x35 & x36 ) | ( ~x35 & n326 ) | ( x36 & n326 ) ;
  assign n328 = ( ~n325 & n326 ) | ( ~n325 & n327 ) | ( n326 & n327 ) ;
  assign n329 = ( x35 & x36 ) | ( x35 & n325 ) | ( x36 & n325 ) ;
  assign n330 = ( x37 & ~x38 ) | ( x37 & n329 ) | ( ~x38 & n329 ) ;
  assign n331 = ( ~x37 & x38 ) | ( ~x37 & n330 ) | ( x38 & n330 ) ;
  assign n332 = ( ~n329 & n330 ) | ( ~n329 & n331 ) | ( n330 & n331 ) ;
  assign n333 = ( x37 & x38 ) | ( x37 & n329 ) | ( x38 & n329 ) ;
  assign n334 = ( x39 & ~x40 ) | ( x39 & n333 ) | ( ~x40 & n333 ) ;
  assign n335 = ( ~x39 & x40 ) | ( ~x39 & n334 ) | ( x40 & n334 ) ;
  assign n336 = ( ~n333 & n334 ) | ( ~n333 & n335 ) | ( n334 & n335 ) ;
  assign n337 = ( x39 & x40 ) | ( x39 & n333 ) | ( x40 & n333 ) ;
  assign n338 = ( x41 & ~x42 ) | ( x41 & n337 ) | ( ~x42 & n337 ) ;
  assign n339 = ( ~x41 & x42 ) | ( ~x41 & n338 ) | ( x42 & n338 ) ;
  assign n340 = ( ~n337 & n338 ) | ( ~n337 & n339 ) | ( n338 & n339 ) ;
  assign n341 = ( x41 & x42 ) | ( x41 & n337 ) | ( x42 & n337 ) ;
  assign n342 = ( x43 & ~x44 ) | ( x43 & n341 ) | ( ~x44 & n341 ) ;
  assign n343 = ( ~x43 & x44 ) | ( ~x43 & n342 ) | ( x44 & n342 ) ;
  assign n344 = ( ~n341 & n342 ) | ( ~n341 & n343 ) | ( n342 & n343 ) ;
  assign n345 = ( x43 & x44 ) | ( x43 & n341 ) | ( x44 & n341 ) ;
  assign n346 = ( x45 & ~x46 ) | ( x45 & n345 ) | ( ~x46 & n345 ) ;
  assign n347 = ( ~x45 & x46 ) | ( ~x45 & n346 ) | ( x46 & n346 ) ;
  assign n348 = ( ~n345 & n346 ) | ( ~n345 & n347 ) | ( n346 & n347 ) ;
  assign n349 = ( x45 & x46 ) | ( x45 & n345 ) | ( x46 & n345 ) ;
  assign n350 = ( x47 & ~x48 ) | ( x47 & n349 ) | ( ~x48 & n349 ) ;
  assign n351 = ( ~x47 & x48 ) | ( ~x47 & n350 ) | ( x48 & n350 ) ;
  assign n352 = ( ~n349 & n350 ) | ( ~n349 & n351 ) | ( n350 & n351 ) ;
  assign n353 = ( x47 & x48 ) | ( x47 & n349 ) | ( x48 & n349 ) ;
  assign n354 = ( x49 & ~x50 ) | ( x49 & n353 ) | ( ~x50 & n353 ) ;
  assign n355 = ( ~x49 & x50 ) | ( ~x49 & n354 ) | ( x50 & n354 ) ;
  assign n356 = ( ~n353 & n354 ) | ( ~n353 & n355 ) | ( n354 & n355 ) ;
  assign n357 = ( x49 & x50 ) | ( x49 & n353 ) | ( x50 & n353 ) ;
  assign n358 = ( x51 & ~x52 ) | ( x51 & n357 ) | ( ~x52 & n357 ) ;
  assign n359 = ( ~x51 & x52 ) | ( ~x51 & n358 ) | ( x52 & n358 ) ;
  assign n360 = ( ~n357 & n358 ) | ( ~n357 & n359 ) | ( n358 & n359 ) ;
  assign n361 = ( x51 & x52 ) | ( x51 & n357 ) | ( x52 & n357 ) ;
  assign n362 = ( x53 & ~x54 ) | ( x53 & n361 ) | ( ~x54 & n361 ) ;
  assign n363 = ( ~x53 & x54 ) | ( ~x53 & n362 ) | ( x54 & n362 ) ;
  assign n364 = ( ~n361 & n362 ) | ( ~n361 & n363 ) | ( n362 & n363 ) ;
  assign n365 = ( x53 & x54 ) | ( x53 & n361 ) | ( x54 & n361 ) ;
  assign n366 = ( x55 & ~x56 ) | ( x55 & n365 ) | ( ~x56 & n365 ) ;
  assign n367 = ( ~x55 & x56 ) | ( ~x55 & n366 ) | ( x56 & n366 ) ;
  assign n368 = ( ~n365 & n366 ) | ( ~n365 & n367 ) | ( n366 & n367 ) ;
  assign n369 = ( x55 & x56 ) | ( x55 & n365 ) | ( x56 & n365 ) ;
  assign n370 = ( x57 & ~x58 ) | ( x57 & n369 ) | ( ~x58 & n369 ) ;
  assign n371 = ( ~x57 & x58 ) | ( ~x57 & n370 ) | ( x58 & n370 ) ;
  assign n372 = ( ~n369 & n370 ) | ( ~n369 & n371 ) | ( n370 & n371 ) ;
  assign n373 = ( x57 & x58 ) | ( x57 & n369 ) | ( x58 & n369 ) ;
  assign n374 = ( x59 & ~x60 ) | ( x59 & n373 ) | ( ~x60 & n373 ) ;
  assign n375 = ( ~x59 & x60 ) | ( ~x59 & n374 ) | ( x60 & n374 ) ;
  assign n376 = ( ~n373 & n374 ) | ( ~n373 & n375 ) | ( n374 & n375 ) ;
  assign n377 = ( x59 & x60 ) | ( x59 & n373 ) | ( x60 & n373 ) ;
  assign n378 = ( x61 & ~x62 ) | ( x61 & n377 ) | ( ~x62 & n377 ) ;
  assign n379 = ( ~x61 & x62 ) | ( ~x61 & n378 ) | ( x62 & n378 ) ;
  assign n380 = ( ~n377 & n378 ) | ( ~n377 & n379 ) | ( n378 & n379 ) ;
  assign n381 = ( x61 & x62 ) | ( x61 & n377 ) | ( x62 & n377 ) ;
  assign n382 = ( x63 & ~x64 ) | ( x63 & n381 ) | ( ~x64 & n381 ) ;
  assign n383 = ( ~x63 & x64 ) | ( ~x63 & n382 ) | ( x64 & n382 ) ;
  assign n384 = ( ~n381 & n382 ) | ( ~n381 & n383 ) | ( n382 & n383 ) ;
  assign n385 = ( x63 & x64 ) | ( x63 & n381 ) | ( x64 & n381 ) ;
  assign n386 = ( x65 & ~x66 ) | ( x65 & n385 ) | ( ~x66 & n385 ) ;
  assign n387 = ( ~x65 & x66 ) | ( ~x65 & n386 ) | ( x66 & n386 ) ;
  assign n388 = ( ~n385 & n386 ) | ( ~n385 & n387 ) | ( n386 & n387 ) ;
  assign n389 = ( x65 & x66 ) | ( x65 & n385 ) | ( x66 & n385 ) ;
  assign n390 = ( x67 & ~x68 ) | ( x67 & n389 ) | ( ~x68 & n389 ) ;
  assign n391 = ( ~x67 & x68 ) | ( ~x67 & n390 ) | ( x68 & n390 ) ;
  assign n392 = ( ~n389 & n390 ) | ( ~n389 & n391 ) | ( n390 & n391 ) ;
  assign n393 = ( x67 & x68 ) | ( x67 & n389 ) | ( x68 & n389 ) ;
  assign n394 = ( x69 & ~x70 ) | ( x69 & n393 ) | ( ~x70 & n393 ) ;
  assign n395 = ( ~x69 & x70 ) | ( ~x69 & n394 ) | ( x70 & n394 ) ;
  assign n396 = ( ~n393 & n394 ) | ( ~n393 & n395 ) | ( n394 & n395 ) ;
  assign n397 = ( x69 & x70 ) | ( x69 & n393 ) | ( x70 & n393 ) ;
  assign n398 = ( x71 & ~x72 ) | ( x71 & n397 ) | ( ~x72 & n397 ) ;
  assign n399 = ( ~x71 & x72 ) | ( ~x71 & n398 ) | ( x72 & n398 ) ;
  assign n400 = ( ~n397 & n398 ) | ( ~n397 & n399 ) | ( n398 & n399 ) ;
  assign n401 = ( x71 & x72 ) | ( x71 & n397 ) | ( x72 & n397 ) ;
  assign n402 = ( x73 & ~x74 ) | ( x73 & n401 ) | ( ~x74 & n401 ) ;
  assign n403 = ( ~x73 & x74 ) | ( ~x73 & n402 ) | ( x74 & n402 ) ;
  assign n404 = ( ~n401 & n402 ) | ( ~n401 & n403 ) | ( n402 & n403 ) ;
  assign n405 = ( x73 & x74 ) | ( x73 & n401 ) | ( x74 & n401 ) ;
  assign n406 = ( x75 & ~x76 ) | ( x75 & n405 ) | ( ~x76 & n405 ) ;
  assign n407 = ( ~x75 & x76 ) | ( ~x75 & n406 ) | ( x76 & n406 ) ;
  assign n408 = ( ~n405 & n406 ) | ( ~n405 & n407 ) | ( n406 & n407 ) ;
  assign n409 = ( x75 & x76 ) | ( x75 & n405 ) | ( x76 & n405 ) ;
  assign n410 = ( x77 & ~x78 ) | ( x77 & n409 ) | ( ~x78 & n409 ) ;
  assign n411 = ( ~x77 & x78 ) | ( ~x77 & n410 ) | ( x78 & n410 ) ;
  assign n412 = ( ~n409 & n410 ) | ( ~n409 & n411 ) | ( n410 & n411 ) ;
  assign n413 = ( x77 & x78 ) | ( x77 & n409 ) | ( x78 & n409 ) ;
  assign n414 = ( x79 & ~x80 ) | ( x79 & n413 ) | ( ~x80 & n413 ) ;
  assign n415 = ( ~x79 & x80 ) | ( ~x79 & n414 ) | ( x80 & n414 ) ;
  assign n416 = ( ~n413 & n414 ) | ( ~n413 & n415 ) | ( n414 & n415 ) ;
  assign n417 = ( x79 & x80 ) | ( x79 & n413 ) | ( x80 & n413 ) ;
  assign n418 = ( x81 & ~x82 ) | ( x81 & n417 ) | ( ~x82 & n417 ) ;
  assign n419 = ( ~x81 & x82 ) | ( ~x81 & n418 ) | ( x82 & n418 ) ;
  assign n420 = ( ~n417 & n418 ) | ( ~n417 & n419 ) | ( n418 & n419 ) ;
  assign n421 = ( x81 & x82 ) | ( x81 & n417 ) | ( x82 & n417 ) ;
  assign n422 = ( x83 & ~x84 ) | ( x83 & n421 ) | ( ~x84 & n421 ) ;
  assign n423 = ( ~x83 & x84 ) | ( ~x83 & n422 ) | ( x84 & n422 ) ;
  assign n424 = ( ~n421 & n422 ) | ( ~n421 & n423 ) | ( n422 & n423 ) ;
  assign n425 = ( x83 & x84 ) | ( x83 & n421 ) | ( x84 & n421 ) ;
  assign n426 = ( x85 & ~x86 ) | ( x85 & n425 ) | ( ~x86 & n425 ) ;
  assign n427 = ( ~x85 & x86 ) | ( ~x85 & n426 ) | ( x86 & n426 ) ;
  assign n428 = ( ~n425 & n426 ) | ( ~n425 & n427 ) | ( n426 & n427 ) ;
  assign n429 = ( x85 & x86 ) | ( x85 & n425 ) | ( x86 & n425 ) ;
  assign n430 = ( x87 & ~x88 ) | ( x87 & n429 ) | ( ~x88 & n429 ) ;
  assign n431 = ( ~x87 & x88 ) | ( ~x87 & n430 ) | ( x88 & n430 ) ;
  assign n432 = ( ~n429 & n430 ) | ( ~n429 & n431 ) | ( n430 & n431 ) ;
  assign n433 = ( x87 & x88 ) | ( x87 & n429 ) | ( x88 & n429 ) ;
  assign n434 = ( x89 & ~x90 ) | ( x89 & n433 ) | ( ~x90 & n433 ) ;
  assign n435 = ( ~x89 & x90 ) | ( ~x89 & n434 ) | ( x90 & n434 ) ;
  assign n436 = ( ~n433 & n434 ) | ( ~n433 & n435 ) | ( n434 & n435 ) ;
  assign n437 = ( x89 & x90 ) | ( x89 & n433 ) | ( x90 & n433 ) ;
  assign n438 = ( x91 & ~x92 ) | ( x91 & n437 ) | ( ~x92 & n437 ) ;
  assign n439 = ( ~x91 & x92 ) | ( ~x91 & n438 ) | ( x92 & n438 ) ;
  assign n440 = ( ~n437 & n438 ) | ( ~n437 & n439 ) | ( n438 & n439 ) ;
  assign n441 = ( x91 & x92 ) | ( x91 & n437 ) | ( x92 & n437 ) ;
  assign n442 = ( x93 & ~x94 ) | ( x93 & n441 ) | ( ~x94 & n441 ) ;
  assign n443 = ( ~x93 & x94 ) | ( ~x93 & n442 ) | ( x94 & n442 ) ;
  assign n444 = ( ~n441 & n442 ) | ( ~n441 & n443 ) | ( n442 & n443 ) ;
  assign n445 = ( x93 & x94 ) | ( x93 & n441 ) | ( x94 & n441 ) ;
  assign n446 = ( x95 & ~x96 ) | ( x95 & n445 ) | ( ~x96 & n445 ) ;
  assign n447 = ( ~x95 & x96 ) | ( ~x95 & n446 ) | ( x96 & n446 ) ;
  assign n448 = ( ~n445 & n446 ) | ( ~n445 & n447 ) | ( n446 & n447 ) ;
  assign n449 = ( x95 & x96 ) | ( x95 & n445 ) | ( x96 & n445 ) ;
  assign n450 = ( x97 & ~x98 ) | ( x97 & n449 ) | ( ~x98 & n449 ) ;
  assign n451 = ( ~x97 & x98 ) | ( ~x97 & n450 ) | ( x98 & n450 ) ;
  assign n452 = ( ~n449 & n450 ) | ( ~n449 & n451 ) | ( n450 & n451 ) ;
  assign n453 = ( x97 & x98 ) | ( x97 & n449 ) | ( x98 & n449 ) ;
  assign n454 = ( x99 & ~x100 ) | ( x99 & n453 ) | ( ~x100 & n453 ) ;
  assign n455 = ( ~x99 & x100 ) | ( ~x99 & n454 ) | ( x100 & n454 ) ;
  assign n456 = ( ~n453 & n454 ) | ( ~n453 & n455 ) | ( n454 & n455 ) ;
  assign n457 = ( x99 & x100 ) | ( x99 & n453 ) | ( x100 & n453 ) ;
  assign n458 = ( x101 & ~x102 ) | ( x101 & n457 ) | ( ~x102 & n457 ) ;
  assign n459 = ( ~x101 & x102 ) | ( ~x101 & n458 ) | ( x102 & n458 ) ;
  assign n460 = ( ~n457 & n458 ) | ( ~n457 & n459 ) | ( n458 & n459 ) ;
  assign n461 = ( x101 & x102 ) | ( x101 & n457 ) | ( x102 & n457 ) ;
  assign n462 = ( x103 & ~x104 ) | ( x103 & n461 ) | ( ~x104 & n461 ) ;
  assign n463 = ( ~x103 & x104 ) | ( ~x103 & n462 ) | ( x104 & n462 ) ;
  assign n464 = ( ~n461 & n462 ) | ( ~n461 & n463 ) | ( n462 & n463 ) ;
  assign n465 = ( x103 & x104 ) | ( x103 & n461 ) | ( x104 & n461 ) ;
  assign n466 = ( x105 & ~x106 ) | ( x105 & n465 ) | ( ~x106 & n465 ) ;
  assign n467 = ( ~x105 & x106 ) | ( ~x105 & n466 ) | ( x106 & n466 ) ;
  assign n468 = ( ~n465 & n466 ) | ( ~n465 & n467 ) | ( n466 & n467 ) ;
  assign n469 = ( x105 & x106 ) | ( x105 & n465 ) | ( x106 & n465 ) ;
  assign n470 = ( x107 & ~x108 ) | ( x107 & n469 ) | ( ~x108 & n469 ) ;
  assign n471 = ( ~x107 & x108 ) | ( ~x107 & n470 ) | ( x108 & n470 ) ;
  assign n472 = ( ~n469 & n470 ) | ( ~n469 & n471 ) | ( n470 & n471 ) ;
  assign n473 = ( x107 & x108 ) | ( x107 & n469 ) | ( x108 & n469 ) ;
  assign n474 = ( x109 & ~x110 ) | ( x109 & n473 ) | ( ~x110 & n473 ) ;
  assign n475 = ( ~x109 & x110 ) | ( ~x109 & n474 ) | ( x110 & n474 ) ;
  assign n476 = ( ~n473 & n474 ) | ( ~n473 & n475 ) | ( n474 & n475 ) ;
  assign n477 = ( x109 & x110 ) | ( x109 & n473 ) | ( x110 & n473 ) ;
  assign n478 = ( x111 & ~x112 ) | ( x111 & n477 ) | ( ~x112 & n477 ) ;
  assign n479 = ( ~x111 & x112 ) | ( ~x111 & n478 ) | ( x112 & n478 ) ;
  assign n480 = ( ~n477 & n478 ) | ( ~n477 & n479 ) | ( n478 & n479 ) ;
  assign n481 = ( x111 & x112 ) | ( x111 & n477 ) | ( x112 & n477 ) ;
  assign n482 = ( x113 & ~x114 ) | ( x113 & n481 ) | ( ~x114 & n481 ) ;
  assign n483 = ( ~x113 & x114 ) | ( ~x113 & n482 ) | ( x114 & n482 ) ;
  assign n484 = ( ~n481 & n482 ) | ( ~n481 & n483 ) | ( n482 & n483 ) ;
  assign n485 = ( x113 & x114 ) | ( x113 & n481 ) | ( x114 & n481 ) ;
  assign n486 = ( x115 & ~x116 ) | ( x115 & n485 ) | ( ~x116 & n485 ) ;
  assign n487 = ( ~x115 & x116 ) | ( ~x115 & n486 ) | ( x116 & n486 ) ;
  assign n488 = ( ~n485 & n486 ) | ( ~n485 & n487 ) | ( n486 & n487 ) ;
  assign n489 = ( x115 & x116 ) | ( x115 & n485 ) | ( x116 & n485 ) ;
  assign n490 = ( x117 & ~x118 ) | ( x117 & n489 ) | ( ~x118 & n489 ) ;
  assign n491 = ( ~x117 & x118 ) | ( ~x117 & n490 ) | ( x118 & n490 ) ;
  assign n492 = ( ~n489 & n490 ) | ( ~n489 & n491 ) | ( n490 & n491 ) ;
  assign n493 = ( x117 & x118 ) | ( x117 & n489 ) | ( x118 & n489 ) ;
  assign n494 = ( x119 & ~x120 ) | ( x119 & n493 ) | ( ~x120 & n493 ) ;
  assign n495 = ( ~x119 & x120 ) | ( ~x119 & n494 ) | ( x120 & n494 ) ;
  assign n496 = ( ~n493 & n494 ) | ( ~n493 & n495 ) | ( n494 & n495 ) ;
  assign n497 = ( x119 & x120 ) | ( x119 & n493 ) | ( x120 & n493 ) ;
  assign n498 = ( x121 & ~x122 ) | ( x121 & n497 ) | ( ~x122 & n497 ) ;
  assign n499 = ( ~x121 & x122 ) | ( ~x121 & n498 ) | ( x122 & n498 ) ;
  assign n500 = ( ~n497 & n498 ) | ( ~n497 & n499 ) | ( n498 & n499 ) ;
  assign n501 = ( x121 & x122 ) | ( x121 & n497 ) | ( x122 & n497 ) ;
  assign n502 = ( x123 & ~x124 ) | ( x123 & n501 ) | ( ~x124 & n501 ) ;
  assign n503 = ( ~x123 & x124 ) | ( ~x123 & n502 ) | ( x124 & n502 ) ;
  assign n504 = ( ~n501 & n502 ) | ( ~n501 & n503 ) | ( n502 & n503 ) ;
  assign n505 = ( x123 & x124 ) | ( x123 & n501 ) | ( x124 & n501 ) ;
  assign n506 = ( x125 & ~x126 ) | ( x125 & n505 ) | ( ~x126 & n505 ) ;
  assign n507 = ( ~x125 & x126 ) | ( ~x125 & n506 ) | ( x126 & n506 ) ;
  assign n508 = ( ~n505 & n506 ) | ( ~n505 & n507 ) | ( n506 & n507 ) ;
  assign n509 = ( x125 & x126 ) | ( x125 & n505 ) | ( x126 & n505 ) ;
  assign n510 = ( x127 & ~x128 ) | ( x127 & n509 ) | ( ~x128 & n509 ) ;
  assign n511 = ( ~x127 & x128 ) | ( ~x127 & n510 ) | ( x128 & n510 ) ;
  assign n512 = ( ~n509 & n510 ) | ( ~n509 & n511 ) | ( n510 & n511 ) ;
  assign n513 = ( x127 & x128 ) | ( x127 & n509 ) | ( x128 & n509 ) ;
  assign n514 = ( x129 & ~x130 ) | ( x129 & n513 ) | ( ~x130 & n513 ) ;
  assign n515 = ( ~x129 & x130 ) | ( ~x129 & n514 ) | ( x130 & n514 ) ;
  assign n516 = ( ~n513 & n514 ) | ( ~n513 & n515 ) | ( n514 & n515 ) ;
  assign n517 = ( x129 & x130 ) | ( x129 & n513 ) | ( x130 & n513 ) ;
  assign n518 = ( x131 & ~x132 ) | ( x131 & n517 ) | ( ~x132 & n517 ) ;
  assign n519 = ( ~x131 & x132 ) | ( ~x131 & n518 ) | ( x132 & n518 ) ;
  assign n520 = ( ~n517 & n518 ) | ( ~n517 & n519 ) | ( n518 & n519 ) ;
  assign n521 = ( x131 & x132 ) | ( x131 & n517 ) | ( x132 & n517 ) ;
  assign n522 = ( x133 & ~x134 ) | ( x133 & n521 ) | ( ~x134 & n521 ) ;
  assign n523 = ( ~x133 & x134 ) | ( ~x133 & n522 ) | ( x134 & n522 ) ;
  assign n524 = ( ~n521 & n522 ) | ( ~n521 & n523 ) | ( n522 & n523 ) ;
  assign n525 = ( x133 & x134 ) | ( x133 & n521 ) | ( x134 & n521 ) ;
  assign n526 = ( x135 & ~x136 ) | ( x135 & n525 ) | ( ~x136 & n525 ) ;
  assign n527 = ( ~x135 & x136 ) | ( ~x135 & n526 ) | ( x136 & n526 ) ;
  assign n528 = ( ~n525 & n526 ) | ( ~n525 & n527 ) | ( n526 & n527 ) ;
  assign n529 = ( x135 & x136 ) | ( x135 & n525 ) | ( x136 & n525 ) ;
  assign n530 = ( x137 & ~x138 ) | ( x137 & n529 ) | ( ~x138 & n529 ) ;
  assign n531 = ( ~x137 & x138 ) | ( ~x137 & n530 ) | ( x138 & n530 ) ;
  assign n532 = ( ~n529 & n530 ) | ( ~n529 & n531 ) | ( n530 & n531 ) ;
  assign n533 = ( x137 & x138 ) | ( x137 & n529 ) | ( x138 & n529 ) ;
  assign n534 = ( x139 & ~x140 ) | ( x139 & n533 ) | ( ~x140 & n533 ) ;
  assign n535 = ( ~x139 & x140 ) | ( ~x139 & n534 ) | ( x140 & n534 ) ;
  assign n536 = ( ~n533 & n534 ) | ( ~n533 & n535 ) | ( n534 & n535 ) ;
  assign n537 = ( x139 & x140 ) | ( x139 & n533 ) | ( x140 & n533 ) ;
  assign n538 = ( x141 & ~x142 ) | ( x141 & n537 ) | ( ~x142 & n537 ) ;
  assign n539 = ( ~x141 & x142 ) | ( ~x141 & n538 ) | ( x142 & n538 ) ;
  assign n540 = ( ~n537 & n538 ) | ( ~n537 & n539 ) | ( n538 & n539 ) ;
  assign n541 = ( x141 & x142 ) | ( x141 & n537 ) | ( x142 & n537 ) ;
  assign n542 = ( x143 & ~x144 ) | ( x143 & n541 ) | ( ~x144 & n541 ) ;
  assign n543 = ( ~x143 & x144 ) | ( ~x143 & n542 ) | ( x144 & n542 ) ;
  assign n544 = ( ~n541 & n542 ) | ( ~n541 & n543 ) | ( n542 & n543 ) ;
  assign n545 = ( x143 & x144 ) | ( x143 & n541 ) | ( x144 & n541 ) ;
  assign n546 = ( x145 & ~x146 ) | ( x145 & n545 ) | ( ~x146 & n545 ) ;
  assign n547 = ( ~x145 & x146 ) | ( ~x145 & n546 ) | ( x146 & n546 ) ;
  assign n548 = ( ~n545 & n546 ) | ( ~n545 & n547 ) | ( n546 & n547 ) ;
  assign n549 = ( x145 & x146 ) | ( x145 & n545 ) | ( x146 & n545 ) ;
  assign n550 = ( x147 & ~x148 ) | ( x147 & n549 ) | ( ~x148 & n549 ) ;
  assign n551 = ( ~x147 & x148 ) | ( ~x147 & n550 ) | ( x148 & n550 ) ;
  assign n552 = ( ~n549 & n550 ) | ( ~n549 & n551 ) | ( n550 & n551 ) ;
  assign n553 = ( x147 & x148 ) | ( x147 & n549 ) | ( x148 & n549 ) ;
  assign n554 = ( x149 & ~x150 ) | ( x149 & n553 ) | ( ~x150 & n553 ) ;
  assign n555 = ( ~x149 & x150 ) | ( ~x149 & n554 ) | ( x150 & n554 ) ;
  assign n556 = ( ~n553 & n554 ) | ( ~n553 & n555 ) | ( n554 & n555 ) ;
  assign n557 = ( x149 & x150 ) | ( x149 & n553 ) | ( x150 & n553 ) ;
  assign n558 = ( x151 & ~x152 ) | ( x151 & n557 ) | ( ~x152 & n557 ) ;
  assign n559 = ( ~x151 & x152 ) | ( ~x151 & n558 ) | ( x152 & n558 ) ;
  assign n560 = ( ~n557 & n558 ) | ( ~n557 & n559 ) | ( n558 & n559 ) ;
  assign n561 = ( x151 & x152 ) | ( x151 & n557 ) | ( x152 & n557 ) ;
  assign n562 = ( x153 & ~x154 ) | ( x153 & n561 ) | ( ~x154 & n561 ) ;
  assign n563 = ( ~x153 & x154 ) | ( ~x153 & n562 ) | ( x154 & n562 ) ;
  assign n564 = ( ~n561 & n562 ) | ( ~n561 & n563 ) | ( n562 & n563 ) ;
  assign n565 = ( x153 & x154 ) | ( x153 & n561 ) | ( x154 & n561 ) ;
  assign n566 = ( x155 & ~x156 ) | ( x155 & n565 ) | ( ~x156 & n565 ) ;
  assign n567 = ( ~x155 & x156 ) | ( ~x155 & n566 ) | ( x156 & n566 ) ;
  assign n568 = ( ~n565 & n566 ) | ( ~n565 & n567 ) | ( n566 & n567 ) ;
  assign n569 = ( x155 & x156 ) | ( x155 & n565 ) | ( x156 & n565 ) ;
  assign n570 = ( x157 & ~x158 ) | ( x157 & n569 ) | ( ~x158 & n569 ) ;
  assign n571 = ( ~x157 & x158 ) | ( ~x157 & n570 ) | ( x158 & n570 ) ;
  assign n572 = ( ~n569 & n570 ) | ( ~n569 & n571 ) | ( n570 & n571 ) ;
  assign n573 = ( x157 & x158 ) | ( x157 & n569 ) | ( x158 & n569 ) ;
  assign n574 = ( x159 & ~x160 ) | ( x159 & n573 ) | ( ~x160 & n573 ) ;
  assign n575 = ( ~x159 & x160 ) | ( ~x159 & n574 ) | ( x160 & n574 ) ;
  assign n576 = ( ~n573 & n574 ) | ( ~n573 & n575 ) | ( n574 & n575 ) ;
  assign n577 = ( x159 & x160 ) | ( x159 & n573 ) | ( x160 & n573 ) ;
  assign n578 = ( x161 & ~x162 ) | ( x161 & n577 ) | ( ~x162 & n577 ) ;
  assign n579 = ( ~x161 & x162 ) | ( ~x161 & n578 ) | ( x162 & n578 ) ;
  assign n580 = ( ~n577 & n578 ) | ( ~n577 & n579 ) | ( n578 & n579 ) ;
  assign n581 = ( x161 & x162 ) | ( x161 & n577 ) | ( x162 & n577 ) ;
  assign n582 = ( x163 & ~x164 ) | ( x163 & n581 ) | ( ~x164 & n581 ) ;
  assign n583 = ( ~x163 & x164 ) | ( ~x163 & n582 ) | ( x164 & n582 ) ;
  assign n584 = ( ~n581 & n582 ) | ( ~n581 & n583 ) | ( n582 & n583 ) ;
  assign n585 = ( x163 & x164 ) | ( x163 & n581 ) | ( x164 & n581 ) ;
  assign n586 = ( x165 & ~x166 ) | ( x165 & n585 ) | ( ~x166 & n585 ) ;
  assign n587 = ( ~x165 & x166 ) | ( ~x165 & n586 ) | ( x166 & n586 ) ;
  assign n588 = ( ~n585 & n586 ) | ( ~n585 & n587 ) | ( n586 & n587 ) ;
  assign n589 = ( x165 & x166 ) | ( x165 & n585 ) | ( x166 & n585 ) ;
  assign n590 = ( x167 & ~x168 ) | ( x167 & n589 ) | ( ~x168 & n589 ) ;
  assign n591 = ( ~x167 & x168 ) | ( ~x167 & n590 ) | ( x168 & n590 ) ;
  assign n592 = ( ~n589 & n590 ) | ( ~n589 & n591 ) | ( n590 & n591 ) ;
  assign n593 = ( x167 & x168 ) | ( x167 & n589 ) | ( x168 & n589 ) ;
  assign n594 = ( x169 & ~x170 ) | ( x169 & n593 ) | ( ~x170 & n593 ) ;
  assign n595 = ( ~x169 & x170 ) | ( ~x169 & n594 ) | ( x170 & n594 ) ;
  assign n596 = ( ~n593 & n594 ) | ( ~n593 & n595 ) | ( n594 & n595 ) ;
  assign n597 = ( x169 & x170 ) | ( x169 & n593 ) | ( x170 & n593 ) ;
  assign n598 = ( x171 & ~x172 ) | ( x171 & n597 ) | ( ~x172 & n597 ) ;
  assign n599 = ( ~x171 & x172 ) | ( ~x171 & n598 ) | ( x172 & n598 ) ;
  assign n600 = ( ~n597 & n598 ) | ( ~n597 & n599 ) | ( n598 & n599 ) ;
  assign n601 = ( x171 & x172 ) | ( x171 & n597 ) | ( x172 & n597 ) ;
  assign n602 = ( x173 & ~x174 ) | ( x173 & n601 ) | ( ~x174 & n601 ) ;
  assign n603 = ( ~x173 & x174 ) | ( ~x173 & n602 ) | ( x174 & n602 ) ;
  assign n604 = ( ~n601 & n602 ) | ( ~n601 & n603 ) | ( n602 & n603 ) ;
  assign n605 = ( x173 & x174 ) | ( x173 & n601 ) | ( x174 & n601 ) ;
  assign n606 = ( x175 & ~x176 ) | ( x175 & n605 ) | ( ~x176 & n605 ) ;
  assign n607 = ( ~x175 & x176 ) | ( ~x175 & n606 ) | ( x176 & n606 ) ;
  assign n608 = ( ~n605 & n606 ) | ( ~n605 & n607 ) | ( n606 & n607 ) ;
  assign n609 = ( x175 & x176 ) | ( x175 & n605 ) | ( x176 & n605 ) ;
  assign n610 = ( x177 & ~x178 ) | ( x177 & n609 ) | ( ~x178 & n609 ) ;
  assign n611 = ( ~x177 & x178 ) | ( ~x177 & n610 ) | ( x178 & n610 ) ;
  assign n612 = ( ~n609 & n610 ) | ( ~n609 & n611 ) | ( n610 & n611 ) ;
  assign n613 = ( x177 & x178 ) | ( x177 & n609 ) | ( x178 & n609 ) ;
  assign n614 = ( x179 & ~x180 ) | ( x179 & n613 ) | ( ~x180 & n613 ) ;
  assign n615 = ( ~x179 & x180 ) | ( ~x179 & n614 ) | ( x180 & n614 ) ;
  assign n616 = ( ~n613 & n614 ) | ( ~n613 & n615 ) | ( n614 & n615 ) ;
  assign n617 = ( x179 & x180 ) | ( x179 & n613 ) | ( x180 & n613 ) ;
  assign n618 = ( x181 & ~x182 ) | ( x181 & n617 ) | ( ~x182 & n617 ) ;
  assign n619 = ( ~x181 & x182 ) | ( ~x181 & n618 ) | ( x182 & n618 ) ;
  assign n620 = ( ~n617 & n618 ) | ( ~n617 & n619 ) | ( n618 & n619 ) ;
  assign n621 = ( x181 & x182 ) | ( x181 & n617 ) | ( x182 & n617 ) ;
  assign n622 = ( x183 & ~x184 ) | ( x183 & n621 ) | ( ~x184 & n621 ) ;
  assign n623 = ( ~x183 & x184 ) | ( ~x183 & n622 ) | ( x184 & n622 ) ;
  assign n624 = ( ~n621 & n622 ) | ( ~n621 & n623 ) | ( n622 & n623 ) ;
  assign n625 = ( x183 & x184 ) | ( x183 & n621 ) | ( x184 & n621 ) ;
  assign n626 = ( x185 & ~x186 ) | ( x185 & n625 ) | ( ~x186 & n625 ) ;
  assign n627 = ( ~x185 & x186 ) | ( ~x185 & n626 ) | ( x186 & n626 ) ;
  assign n628 = ( ~n625 & n626 ) | ( ~n625 & n627 ) | ( n626 & n627 ) ;
  assign n629 = ( x185 & x186 ) | ( x185 & n625 ) | ( x186 & n625 ) ;
  assign n630 = ( x187 & ~x188 ) | ( x187 & n629 ) | ( ~x188 & n629 ) ;
  assign n631 = ( ~x187 & x188 ) | ( ~x187 & n630 ) | ( x188 & n630 ) ;
  assign n632 = ( ~n629 & n630 ) | ( ~n629 & n631 ) | ( n630 & n631 ) ;
  assign n633 = ( x187 & x188 ) | ( x187 & n629 ) | ( x188 & n629 ) ;
  assign n634 = ( x189 & ~x190 ) | ( x189 & n633 ) | ( ~x190 & n633 ) ;
  assign n635 = ( ~x189 & x190 ) | ( ~x189 & n634 ) | ( x190 & n634 ) ;
  assign n636 = ( ~n633 & n634 ) | ( ~n633 & n635 ) | ( n634 & n635 ) ;
  assign n637 = ( x189 & x190 ) | ( x189 & n633 ) | ( x190 & n633 ) ;
  assign n638 = ( x191 & ~x192 ) | ( x191 & n637 ) | ( ~x192 & n637 ) ;
  assign n639 = ( ~x191 & x192 ) | ( ~x191 & n638 ) | ( x192 & n638 ) ;
  assign n640 = ( ~n637 & n638 ) | ( ~n637 & n639 ) | ( n638 & n639 ) ;
  assign n641 = ( x191 & x192 ) | ( x191 & n637 ) | ( x192 & n637 ) ;
  assign n642 = ( x193 & ~x194 ) | ( x193 & n641 ) | ( ~x194 & n641 ) ;
  assign n643 = ( ~x193 & x194 ) | ( ~x193 & n642 ) | ( x194 & n642 ) ;
  assign n644 = ( ~n641 & n642 ) | ( ~n641 & n643 ) | ( n642 & n643 ) ;
  assign n645 = ( x193 & x194 ) | ( x193 & n641 ) | ( x194 & n641 ) ;
  assign n646 = ( x195 & ~x196 ) | ( x195 & n645 ) | ( ~x196 & n645 ) ;
  assign n647 = ( ~x195 & x196 ) | ( ~x195 & n646 ) | ( x196 & n646 ) ;
  assign n648 = ( ~n645 & n646 ) | ( ~n645 & n647 ) | ( n646 & n647 ) ;
  assign n649 = ( x195 & x196 ) | ( x195 & n645 ) | ( x196 & n645 ) ;
  assign n650 = ( x197 & ~x198 ) | ( x197 & n649 ) | ( ~x198 & n649 ) ;
  assign n651 = ( ~x197 & x198 ) | ( ~x197 & n650 ) | ( x198 & n650 ) ;
  assign n652 = ( ~n649 & n650 ) | ( ~n649 & n651 ) | ( n650 & n651 ) ;
  assign n653 = ( x197 & x198 ) | ( x197 & n649 ) | ( x198 & n649 ) ;
  assign n654 = ( x199 & ~x200 ) | ( x199 & n653 ) | ( ~x200 & n653 ) ;
  assign n655 = ( ~x199 & x200 ) | ( ~x199 & n654 ) | ( x200 & n654 ) ;
  assign n656 = ( ~n653 & n654 ) | ( ~n653 & n655 ) | ( n654 & n655 ) ;
  assign n657 = ( x199 & x200 ) | ( x199 & n653 ) | ( x200 & n653 ) ;
  assign n658 = ( x201 & ~x202 ) | ( x201 & n657 ) | ( ~x202 & n657 ) ;
  assign n659 = ( ~x201 & x202 ) | ( ~x201 & n658 ) | ( x202 & n658 ) ;
  assign n660 = ( ~n657 & n658 ) | ( ~n657 & n659 ) | ( n658 & n659 ) ;
  assign n661 = ( x201 & x202 ) | ( x201 & n657 ) | ( x202 & n657 ) ;
  assign n662 = ( x203 & ~x204 ) | ( x203 & n661 ) | ( ~x204 & n661 ) ;
  assign n663 = ( ~x203 & x204 ) | ( ~x203 & n662 ) | ( x204 & n662 ) ;
  assign n664 = ( ~n661 & n662 ) | ( ~n661 & n663 ) | ( n662 & n663 ) ;
  assign n665 = ( x203 & x204 ) | ( x203 & n661 ) | ( x204 & n661 ) ;
  assign n666 = ( x205 & ~x206 ) | ( x205 & n665 ) | ( ~x206 & n665 ) ;
  assign n667 = ( ~x205 & x206 ) | ( ~x205 & n666 ) | ( x206 & n666 ) ;
  assign n668 = ( ~n665 & n666 ) | ( ~n665 & n667 ) | ( n666 & n667 ) ;
  assign n669 = ( x205 & x206 ) | ( x205 & n665 ) | ( x206 & n665 ) ;
  assign n670 = ( x207 & ~x208 ) | ( x207 & n669 ) | ( ~x208 & n669 ) ;
  assign n671 = ( ~x207 & x208 ) | ( ~x207 & n670 ) | ( x208 & n670 ) ;
  assign n672 = ( ~n669 & n670 ) | ( ~n669 & n671 ) | ( n670 & n671 ) ;
  assign n673 = ( x207 & x208 ) | ( x207 & n669 ) | ( x208 & n669 ) ;
  assign n674 = ( x209 & ~x210 ) | ( x209 & n673 ) | ( ~x210 & n673 ) ;
  assign n675 = ( ~x209 & x210 ) | ( ~x209 & n674 ) | ( x210 & n674 ) ;
  assign n676 = ( ~n673 & n674 ) | ( ~n673 & n675 ) | ( n674 & n675 ) ;
  assign n677 = ( x209 & x210 ) | ( x209 & n673 ) | ( x210 & n673 ) ;
  assign n678 = ( x211 & ~x212 ) | ( x211 & n677 ) | ( ~x212 & n677 ) ;
  assign n679 = ( ~x211 & x212 ) | ( ~x211 & n678 ) | ( x212 & n678 ) ;
  assign n680 = ( ~n677 & n678 ) | ( ~n677 & n679 ) | ( n678 & n679 ) ;
  assign n681 = ( x211 & x212 ) | ( x211 & n677 ) | ( x212 & n677 ) ;
  assign n682 = ( x213 & ~x214 ) | ( x213 & n681 ) | ( ~x214 & n681 ) ;
  assign n683 = ( ~x213 & x214 ) | ( ~x213 & n682 ) | ( x214 & n682 ) ;
  assign n684 = ( ~n681 & n682 ) | ( ~n681 & n683 ) | ( n682 & n683 ) ;
  assign n685 = ( x213 & x214 ) | ( x213 & n681 ) | ( x214 & n681 ) ;
  assign n686 = ( x215 & ~x216 ) | ( x215 & n685 ) | ( ~x216 & n685 ) ;
  assign n687 = ( ~x215 & x216 ) | ( ~x215 & n686 ) | ( x216 & n686 ) ;
  assign n688 = ( ~n685 & n686 ) | ( ~n685 & n687 ) | ( n686 & n687 ) ;
  assign n689 = ( x215 & x216 ) | ( x215 & n685 ) | ( x216 & n685 ) ;
  assign n690 = ( x217 & ~x218 ) | ( x217 & n689 ) | ( ~x218 & n689 ) ;
  assign n691 = ( ~x217 & x218 ) | ( ~x217 & n690 ) | ( x218 & n690 ) ;
  assign n692 = ( ~n689 & n690 ) | ( ~n689 & n691 ) | ( n690 & n691 ) ;
  assign n693 = ( x217 & x218 ) | ( x217 & n689 ) | ( x218 & n689 ) ;
  assign n694 = ( x219 & ~x220 ) | ( x219 & n693 ) | ( ~x220 & n693 ) ;
  assign n695 = ( ~x219 & x220 ) | ( ~x219 & n694 ) | ( x220 & n694 ) ;
  assign n696 = ( ~n693 & n694 ) | ( ~n693 & n695 ) | ( n694 & n695 ) ;
  assign n697 = ( x219 & x220 ) | ( x219 & n693 ) | ( x220 & n693 ) ;
  assign n698 = ( x221 & ~x222 ) | ( x221 & n697 ) | ( ~x222 & n697 ) ;
  assign n699 = ( ~x221 & x222 ) | ( ~x221 & n698 ) | ( x222 & n698 ) ;
  assign n700 = ( ~n697 & n698 ) | ( ~n697 & n699 ) | ( n698 & n699 ) ;
  assign n701 = ( x221 & x222 ) | ( x221 & n697 ) | ( x222 & n697 ) ;
  assign n702 = ( x223 & ~x224 ) | ( x223 & n701 ) | ( ~x224 & n701 ) ;
  assign n703 = ( ~x223 & x224 ) | ( ~x223 & n702 ) | ( x224 & n702 ) ;
  assign n704 = ( ~n701 & n702 ) | ( ~n701 & n703 ) | ( n702 & n703 ) ;
  assign n705 = ( x223 & x224 ) | ( x223 & n701 ) | ( x224 & n701 ) ;
  assign n706 = ( x225 & ~x226 ) | ( x225 & n705 ) | ( ~x226 & n705 ) ;
  assign n707 = ( ~x225 & x226 ) | ( ~x225 & n706 ) | ( x226 & n706 ) ;
  assign n708 = ( ~n705 & n706 ) | ( ~n705 & n707 ) | ( n706 & n707 ) ;
  assign n709 = ( x225 & x226 ) | ( x225 & n705 ) | ( x226 & n705 ) ;
  assign n710 = ( x227 & ~x228 ) | ( x227 & n709 ) | ( ~x228 & n709 ) ;
  assign n711 = ( ~x227 & x228 ) | ( ~x227 & n710 ) | ( x228 & n710 ) ;
  assign n712 = ( ~n709 & n710 ) | ( ~n709 & n711 ) | ( n710 & n711 ) ;
  assign n713 = ( x227 & x228 ) | ( x227 & n709 ) | ( x228 & n709 ) ;
  assign n714 = ( x229 & ~x230 ) | ( x229 & n713 ) | ( ~x230 & n713 ) ;
  assign n715 = ( ~x229 & x230 ) | ( ~x229 & n714 ) | ( x230 & n714 ) ;
  assign n716 = ( ~n713 & n714 ) | ( ~n713 & n715 ) | ( n714 & n715 ) ;
  assign n717 = ( x229 & x230 ) | ( x229 & n713 ) | ( x230 & n713 ) ;
  assign n718 = ( x231 & ~x232 ) | ( x231 & n717 ) | ( ~x232 & n717 ) ;
  assign n719 = ( ~x231 & x232 ) | ( ~x231 & n718 ) | ( x232 & n718 ) ;
  assign n720 = ( ~n717 & n718 ) | ( ~n717 & n719 ) | ( n718 & n719 ) ;
  assign n721 = ( x231 & x232 ) | ( x231 & n717 ) | ( x232 & n717 ) ;
  assign n722 = ( x233 & ~x234 ) | ( x233 & n721 ) | ( ~x234 & n721 ) ;
  assign n723 = ( ~x233 & x234 ) | ( ~x233 & n722 ) | ( x234 & n722 ) ;
  assign n724 = ( ~n721 & n722 ) | ( ~n721 & n723 ) | ( n722 & n723 ) ;
  assign n725 = ( x233 & x234 ) | ( x233 & n721 ) | ( x234 & n721 ) ;
  assign n726 = ( x235 & ~x236 ) | ( x235 & n725 ) | ( ~x236 & n725 ) ;
  assign n727 = ( ~x235 & x236 ) | ( ~x235 & n726 ) | ( x236 & n726 ) ;
  assign n728 = ( ~n725 & n726 ) | ( ~n725 & n727 ) | ( n726 & n727 ) ;
  assign n729 = ( x235 & x236 ) | ( x235 & n725 ) | ( x236 & n725 ) ;
  assign n730 = ( x237 & ~x238 ) | ( x237 & n729 ) | ( ~x238 & n729 ) ;
  assign n731 = ( ~x237 & x238 ) | ( ~x237 & n730 ) | ( x238 & n730 ) ;
  assign n732 = ( ~n729 & n730 ) | ( ~n729 & n731 ) | ( n730 & n731 ) ;
  assign n733 = ( x237 & x238 ) | ( x237 & n729 ) | ( x238 & n729 ) ;
  assign n734 = ( x239 & ~x240 ) | ( x239 & n733 ) | ( ~x240 & n733 ) ;
  assign n735 = ( ~x239 & x240 ) | ( ~x239 & n734 ) | ( x240 & n734 ) ;
  assign n736 = ( ~n733 & n734 ) | ( ~n733 & n735 ) | ( n734 & n735 ) ;
  assign n737 = ( x239 & x240 ) | ( x239 & n733 ) | ( x240 & n733 ) ;
  assign n738 = ( x241 & ~x242 ) | ( x241 & n737 ) | ( ~x242 & n737 ) ;
  assign n739 = ( ~x241 & x242 ) | ( ~x241 & n738 ) | ( x242 & n738 ) ;
  assign n740 = ( ~n737 & n738 ) | ( ~n737 & n739 ) | ( n738 & n739 ) ;
  assign n741 = ( x241 & x242 ) | ( x241 & n737 ) | ( x242 & n737 ) ;
  assign n742 = ( x243 & ~x244 ) | ( x243 & n741 ) | ( ~x244 & n741 ) ;
  assign n743 = ( ~x243 & x244 ) | ( ~x243 & n742 ) | ( x244 & n742 ) ;
  assign n744 = ( ~n741 & n742 ) | ( ~n741 & n743 ) | ( n742 & n743 ) ;
  assign n745 = ( x243 & x244 ) | ( x243 & n741 ) | ( x244 & n741 ) ;
  assign n746 = ( x245 & ~x246 ) | ( x245 & n745 ) | ( ~x246 & n745 ) ;
  assign n747 = ( ~x245 & x246 ) | ( ~x245 & n746 ) | ( x246 & n746 ) ;
  assign n748 = ( ~n745 & n746 ) | ( ~n745 & n747 ) | ( n746 & n747 ) ;
  assign n749 = ( x245 & x246 ) | ( x245 & n745 ) | ( x246 & n745 ) ;
  assign n750 = ( x247 & ~x248 ) | ( x247 & n749 ) | ( ~x248 & n749 ) ;
  assign n751 = ( ~x247 & x248 ) | ( ~x247 & n750 ) | ( x248 & n750 ) ;
  assign n752 = ( ~n749 & n750 ) | ( ~n749 & n751 ) | ( n750 & n751 ) ;
  assign n753 = ( x247 & x248 ) | ( x247 & n749 ) | ( x248 & n749 ) ;
  assign n754 = ( x249 & ~x250 ) | ( x249 & n753 ) | ( ~x250 & n753 ) ;
  assign n755 = ( ~x249 & x250 ) | ( ~x249 & n754 ) | ( x250 & n754 ) ;
  assign n756 = ( ~n753 & n754 ) | ( ~n753 & n755 ) | ( n754 & n755 ) ;
  assign n757 = ( x249 & x250 ) | ( x249 & n753 ) | ( x250 & n753 ) ;
  assign n758 = ( x251 & ~x252 ) | ( x251 & n757 ) | ( ~x252 & n757 ) ;
  assign n759 = ( ~x251 & x252 ) | ( ~x251 & n758 ) | ( x252 & n758 ) ;
  assign n760 = ( ~n757 & n758 ) | ( ~n757 & n759 ) | ( n758 & n759 ) ;
  assign n761 = ( x251 & x252 ) | ( x251 & n757 ) | ( x252 & n757 ) ;
  assign n762 = ( x253 & ~x254 ) | ( x253 & n761 ) | ( ~x254 & n761 ) ;
  assign n763 = ( ~x253 & x254 ) | ( ~x253 & n762 ) | ( x254 & n762 ) ;
  assign n764 = ( ~n761 & n762 ) | ( ~n761 & n763 ) | ( n762 & n763 ) ;
  assign n765 = ( x253 & x254 ) | ( x253 & n761 ) | ( x254 & n761 ) ;
  assign n766 = ( x255 & ~x256 ) | ( x255 & n765 ) | ( ~x256 & n765 ) ;
  assign n767 = ( ~x255 & x256 ) | ( ~x255 & n766 ) | ( x256 & n766 ) ;
  assign n768 = ( ~n765 & n766 ) | ( ~n765 & n767 ) | ( n766 & n767 ) ;
  assign n769 = ( x255 & x256 ) | ( x255 & n765 ) | ( x256 & n765 ) ;
  assign y0 = n260 ;
  assign y1 = n264 ;
  assign y2 = n268 ;
  assign y3 = n272 ;
  assign y4 = n276 ;
  assign y5 = n280 ;
  assign y6 = n284 ;
  assign y7 = n288 ;
  assign y8 = n292 ;
  assign y9 = n296 ;
  assign y10 = n300 ;
  assign y11 = n304 ;
  assign y12 = n308 ;
  assign y13 = n312 ;
  assign y14 = n316 ;
  assign y15 = n320 ;
  assign y16 = n324 ;
  assign y17 = n328 ;
  assign y18 = n332 ;
  assign y19 = n336 ;
  assign y20 = n340 ;
  assign y21 = n344 ;
  assign y22 = n348 ;
  assign y23 = n352 ;
  assign y24 = n356 ;
  assign y25 = n360 ;
  assign y26 = n364 ;
  assign y27 = n368 ;
  assign y28 = n372 ;
  assign y29 = n376 ;
  assign y30 = n380 ;
  assign y31 = n384 ;
  assign y32 = n388 ;
  assign y33 = n392 ;
  assign y34 = n396 ;
  assign y35 = n400 ;
  assign y36 = n404 ;
  assign y37 = n408 ;
  assign y38 = n412 ;
  assign y39 = n416 ;
  assign y40 = n420 ;
  assign y41 = n424 ;
  assign y42 = n428 ;
  assign y43 = n432 ;
  assign y44 = n436 ;
  assign y45 = n440 ;
  assign y46 = n444 ;
  assign y47 = n448 ;
  assign y48 = n452 ;
  assign y49 = n456 ;
  assign y50 = n460 ;
  assign y51 = n464 ;
  assign y52 = n468 ;
  assign y53 = n472 ;
  assign y54 = n476 ;
  assign y55 = n480 ;
  assign y56 = n484 ;
  assign y57 = n488 ;
  assign y58 = n492 ;
  assign y59 = n496 ;
  assign y60 = n500 ;
  assign y61 = n504 ;
  assign y62 = n508 ;
  assign y63 = n512 ;
  assign y64 = n516 ;
  assign y65 = n520 ;
  assign y66 = n524 ;
  assign y67 = n528 ;
  assign y68 = n532 ;
  assign y69 = n536 ;
  assign y70 = n540 ;
  assign y71 = n544 ;
  assign y72 = n548 ;
  assign y73 = n552 ;
  assign y74 = n556 ;
  assign y75 = n560 ;
  assign y76 = n564 ;
  assign y77 = n568 ;
  assign y78 = n572 ;
  assign y79 = n576 ;
  assign y80 = n580 ;
  assign y81 = n584 ;
  assign y82 = n588 ;
  assign y83 = n592 ;
  assign y84 = n596 ;
  assign y85 = n600 ;
  assign y86 = n604 ;
  assign y87 = n608 ;
  assign y88 = n612 ;
  assign y89 = n616 ;
  assign y90 = n620 ;
  assign y91 = n624 ;
  assign y92 = n628 ;
  assign y93 = n632 ;
  assign y94 = n636 ;
  assign y95 = n640 ;
  assign y96 = n644 ;
  assign y97 = n648 ;
  assign y98 = n652 ;
  assign y99 = n656 ;
  assign y100 = n660 ;
  assign y101 = n664 ;
  assign y102 = n668 ;
  assign y103 = n672 ;
  assign y104 = n676 ;
  assign y105 = n680 ;
  assign y106 = n684 ;
  assign y107 = n688 ;
  assign y108 = n692 ;
  assign y109 = n696 ;
  assign y110 = n700 ;
  assign y111 = n704 ;
  assign y112 = n708 ;
  assign y113 = n712 ;
  assign y114 = n716 ;
  assign y115 = n720 ;
  assign y116 = n724 ;
  assign y117 = n728 ;
  assign y118 = n732 ;
  assign y119 = n736 ;
  assign y120 = n740 ;
  assign y121 = n744 ;
  assign y122 = n748 ;
  assign y123 = n752 ;
  assign y124 = n756 ;
  assign y125 = n760 ;
  assign y126 = n764 ;
  assign y127 = n768 ;
  assign y128 = n769 ;
endmodule
