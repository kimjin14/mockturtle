module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 ;
  wire n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 ;
  assign n8 = x3 & x4 ;
  assign n9 = ( x1 & x2 ) | ( x1 & x4 ) | ( x2 & x4 ) ;
  assign n10 = x1 | n8 ;
  assign n11 = ~x3 & x4 ;
  assign n12 = x3 | n11 ;
  assign n13 = ~n8 & n12 ;
  assign n14 = ~x0 & n12 ;
  assign n15 = ( n12 & n13 ) | ( n12 & n14 ) | ( n13 & n14 ) ;
  assign n16 = x0 & ~x1 ;
  assign n17 = x3 & ~n8 ;
  assign n18 = n16 & n17 ;
  assign n19 = ( n10 & ~n15 ) | ( n10 & n18 ) | ( ~n15 & n18 ) ;
  assign n20 = ( n8 & n9 ) | ( n8 & n19 ) | ( n9 & n19 ) ;
  assign n21 = x1 | x2 ;
  assign n22 = ( x0 & x3 ) | ( x0 & n12 ) | ( x3 & n12 ) ;
  assign n23 = x1 & n22 ;
  assign n24 = ( x1 & n19 ) | ( x1 & n23 ) | ( n19 & n23 ) ;
  assign n25 = n10 & ~n24 ;
  assign n26 = x2 | n25 ;
  assign n27 = x1 & ~x2 ;
  assign n28 = ( x2 & n15 ) | ( x2 & ~n27 ) | ( n15 & ~n27 ) ;
  assign n29 = ( ~x2 & n11 ) | ( ~x2 & n28 ) | ( n11 & n28 ) ;
  assign n30 = ( n21 & n26 ) | ( n21 & n29 ) | ( n26 & n29 ) ;
  assign n31 = ( ~x1 & x2 ) | ( ~x1 & n13 ) | ( x2 & n13 ) ;
  assign n32 = ( x2 & n8 ) | ( x2 & n31 ) | ( n8 & n31 ) ;
  assign n33 = n30 & ~n32 ;
  assign n34 = ~x0 & x3 ;
  assign n35 = ( x1 & n10 ) | ( x1 & n34 ) | ( n10 & n34 ) ;
  assign n36 = ( n17 & n25 ) | ( n17 & n35 ) | ( n25 & n35 ) ;
  assign n37 = ~x2 & n36 ;
  assign n38 = x2 & ~n11 ;
  assign n39 = ( x2 & n14 ) | ( x2 & n38 ) | ( n14 & n38 ) ;
  assign n40 = x4 & x5 ;
  assign n41 = n34 & n40 ;
  assign n42 = x3 & ~x6 ;
  assign n43 = ~n8 & n42 ;
  assign n44 = x0 & x1 ;
  assign n45 = ( x3 & x5 ) | ( x3 & n17 ) | ( x5 & n17 ) ;
  assign n46 = n44 & n45 ;
  assign n47 = ( x6 & n43 ) | ( x6 & n46 ) | ( n43 & n46 ) ;
  assign n48 = ( x2 & n21 ) | ( x2 & n47 ) | ( n21 & n47 ) ;
  assign n49 = ( n21 & n41 ) | ( n21 & n48 ) | ( n41 & n48 ) ;
  assign n50 = ~n39 & n49 ;
  assign n51 = ( x3 & x6 ) | ( x3 & n43 ) | ( x6 & n43 ) ;
  assign n52 = ( x1 & x2 ) | ( x1 & n51 ) | ( x2 & n51 ) ;
  assign n53 = ~n38 & n52 ;
  assign n54 = x2 & n8 ;
  assign n55 = x2 | n31 ;
  assign n56 = n23 | n55 ;
  assign n57 = n8 & ~n44 ;
  assign n58 = ( n30 & n56 ) | ( n30 & ~n57 ) | ( n56 & ~n57 ) ;
  assign n59 = ( ~x2 & n54 ) | ( ~x2 & n58 ) | ( n54 & n58 ) ;
  assign n60 = ( n19 & n28 ) | ( n19 & n37 ) | ( n28 & n37 ) ;
  assign n61 = n26 & ~n32 ;
  assign n62 = ( x1 & n54 ) | ( x1 & n61 ) | ( n54 & n61 ) ;
  assign n63 = ~n38 & n56 ;
  assign n64 = x0 | n14 ;
  assign n65 = x2 | n64 ;
  assign n66 = x1 | n65 ;
  assign n67 = ( x1 & ~x2 ) | ( x1 & n17 ) | ( ~x2 & n17 ) ;
  assign n68 = n9 & ~n67 ;
  assign n69 = ( ~x2 & n22 ) | ( ~x2 & n61 ) | ( n22 & n61 ) ;
  assign n70 = n68 | n69 ;
  assign n71 = x2 & ~n12 ;
  assign n72 = x0 & n71 ;
  assign n73 = x2 & ~n64 ;
  assign n74 = ~x0 & n17 ;
  assign n75 = x2 & n74 ;
  assign n76 = ~x1 & n75 ;
  assign n77 = ( x2 & n18 ) | ( x2 & n27 ) | ( n18 & n27 ) ;
  assign n78 = x0 & ~n11 ;
  assign n79 = ( x2 & n16 ) | ( x2 & n78 ) | ( n16 & n78 ) ;
  assign n80 = ( n36 & n76 ) | ( n36 & n79 ) | ( n76 & n79 ) ;
  assign n81 = x1 & n75 ;
  assign n82 = x2 | n18 ;
  assign n83 = n46 | n82 ;
  assign n84 = x2 & ~n57 ;
  assign n85 = n83 & ~n84 ;
  assign n86 = ( n18 & n46 ) | ( n18 & ~n47 ) | ( n46 & ~n47 ) ;
  assign n87 = ( x1 & n16 ) | ( x1 & n86 ) | ( n16 & n86 ) ;
  assign n88 = ~x2 & n87 ;
  assign n89 = ( n47 & n57 ) | ( n47 & n85 ) | ( n57 & n85 ) ;
  assign n90 = ( x0 & ~x1 ) | ( x0 & x2 ) | ( ~x1 & x2 ) ;
  assign n91 = ( x0 & ~x1 ) | ( x0 & n11 ) | ( ~x1 & n11 ) ;
  assign n92 = ~n90 & n91 ;
  assign n93 = n16 & ~n79 ;
  assign y0 = n20 ;
  assign y1 = n33 ;
  assign y2 = n37 ;
  assign y3 = n29 ;
  assign y4 = n50 ;
  assign y5 = n53 ;
  assign y6 = n59 ;
  assign y7 = n60 ;
  assign y8 = n62 ;
  assign y9 = n61 ;
  assign y10 = n63 ;
  assign y11 = ~n66 ;
  assign y12 = n70 ;
  assign y13 = n72 ;
  assign y14 = n73 ;
  assign y15 = n76 ;
  assign y16 = n77 ;
  assign y17 = n80 ;
  assign y18 = n81 ;
  assign y19 = n71 ;
  assign y20 = n85 ;
  assign y21 = n88 ;
  assign y22 = n89 ;
  assign y23 = ~1'b0 ;
  assign y24 = n92 ;
  assign y25 = n93 ;
endmodule
