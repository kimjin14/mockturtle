module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 , x147 , x148 , x149 , x150 , x151 , x152 , x153 , x154 , x155 , x156 , x157 , x158 , x159 , x160 , x161 , x162 , x163 , x164 , x165 , x166 , x167 , x168 , x169 , x170 , x171 , x172 , x173 , x174 , x175 , x176 , x177 , x178 , x179 , x180 , x181 , x182 , x183 , x184 , x185 , x186 , x187 , x188 , x189 , x190 , x191 , x192 , x193 , x194 , x195 , x196 , x197 , x198 , x199 , x200 , x201 , x202 , x203 , x204 , x205 , x206 , x207 , x208 , x209 , x210 , x211 , x212 , x213 , x214 , x215 , x216 , x217 , x218 , x219 , x220 , x221 , x222 , x223 , x224 , x225 , x226 , x227 , x228 , x229 , x230 , x231 , x232 , x233 , x234 , x235 , x236 , x237 , x238 , x239 , x240 , x241 , x242 , x243 , x244 , x245 , x246 , x247 , x248 , x249 , x250 , x251 , x252 , x253 , x254 , x255 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 , y128 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 , x147 , x148 , x149 , x150 , x151 , x152 , x153 , x154 , x155 , x156 , x157 , x158 , x159 , x160 , x161 , x162 , x163 , x164 , x165 , x166 , x167 , x168 , x169 , x170 , x171 , x172 , x173 , x174 , x175 , x176 , x177 , x178 , x179 , x180 , x181 , x182 , x183 , x184 , x185 , x186 , x187 , x188 , x189 , x190 , x191 , x192 , x193 , x194 , x195 , x196 , x197 , x198 , x199 , x200 , x201 , x202 , x203 , x204 , x205 , x206 , x207 , x208 , x209 , x210 , x211 , x212 , x213 , x214 , x215 , x216 , x217 , x218 , x219 , x220 , x221 , x222 , x223 , x224 , x225 , x226 , x227 , x228 , x229 , x230 , x231 , x232 , x233 , x234 , x235 , x236 , x237 , x238 , x239 , x240 , x241 , x242 , x243 , x244 , x245 , x246 , x247 , x248 , x249 , x250 , x251 , x252 , x253 , x254 , x255 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 , y128 ;
  wire n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 ;
  assign n257 = x0 & ~x128 ;
  assign n258 = ~x0 & x128 ;
  assign n259 = n257 | n258 ;
  assign n260 = x0 & x128 ;
  assign n261 = ( x1 & ~x129 ) | ( x1 & n260 ) | ( ~x129 & n260 ) ;
  assign n262 = ( ~x1 & x129 ) | ( ~x1 & n261 ) | ( x129 & n261 ) ;
  assign n263 = ( ~n260 & n261 ) | ( ~n260 & n262 ) | ( n261 & n262 ) ;
  assign n264 = x1 & x129 ;
  assign n265 = x1 | x129 ;
  assign n266 = n260 & n265 ;
  assign n267 = n264 | n266 ;
  assign n268 = ( x2 & ~x130 ) | ( x2 & n267 ) | ( ~x130 & n267 ) ;
  assign n269 = ( ~x2 & x130 ) | ( ~x2 & n268 ) | ( x130 & n268 ) ;
  assign n270 = ( ~n267 & n268 ) | ( ~n267 & n269 ) | ( n268 & n269 ) ;
  assign n271 = x3 | x131 ;
  assign n272 = x3 & x131 ;
  assign n273 = n271 | n272 ;
  assign n274 = x2 & x130 ;
  assign n275 = x2 | x130 ;
  assign n276 = n264 & n275 ;
  assign n277 = ( n266 & n275 ) | ( n266 & n276 ) | ( n275 & n276 ) ;
  assign n278 = n274 | n277 ;
  assign n279 = ( n272 & ~n273 ) | ( n272 & n278 ) | ( ~n273 & n278 ) ;
  assign n280 = ( n272 & n273 ) | ( n272 & n278 ) | ( n273 & n278 ) ;
  assign n281 = ( n273 & n279 ) | ( n273 & ~n280 ) | ( n279 & ~n280 ) ;
  assign n282 = ( x3 & x131 ) | ( x3 & n274 ) | ( x131 & n274 ) ;
  assign n283 = ( n271 & n277 ) | ( n271 & n282 ) | ( n277 & n282 ) ;
  assign n284 = ( x4 & ~x132 ) | ( x4 & n283 ) | ( ~x132 & n283 ) ;
  assign n285 = ( ~x4 & x132 ) | ( ~x4 & n284 ) | ( x132 & n284 ) ;
  assign n286 = ( ~n283 & n284 ) | ( ~n283 & n285 ) | ( n284 & n285 ) ;
  assign n287 = x4 & x132 ;
  assign n288 = x4 | x132 ;
  assign n289 = n287 | n288 ;
  assign n290 = ( n283 & n287 ) | ( n283 & n289 ) | ( n287 & n289 ) ;
  assign n291 = ( x5 & ~x133 ) | ( x5 & n290 ) | ( ~x133 & n290 ) ;
  assign n292 = ( ~x5 & x133 ) | ( ~x5 & n291 ) | ( x133 & n291 ) ;
  assign n293 = ( ~n290 & n291 ) | ( ~n290 & n292 ) | ( n291 & n292 ) ;
  assign n294 = x5 & x133 ;
  assign n295 = x5 | x133 ;
  assign n296 = n287 & n295 ;
  assign n297 = n294 | n296 ;
  assign n298 = n294 | n295 ;
  assign n299 = ( n289 & n294 ) | ( n289 & n298 ) | ( n294 & n298 ) ;
  assign n300 = ( n283 & n297 ) | ( n283 & n299 ) | ( n297 & n299 ) ;
  assign n301 = ( x6 & ~x134 ) | ( x6 & n300 ) | ( ~x134 & n300 ) ;
  assign n302 = ( ~x6 & x134 ) | ( ~x6 & n301 ) | ( x134 & n301 ) ;
  assign n303 = ( ~n300 & n301 ) | ( ~n300 & n302 ) | ( n301 & n302 ) ;
  assign n304 = x6 & x134 ;
  assign n305 = x6 | x134 ;
  assign n306 = n304 | n305 ;
  assign n307 = ( n300 & n304 ) | ( n300 & n306 ) | ( n304 & n306 ) ;
  assign n308 = ( x7 & ~x135 ) | ( x7 & n307 ) | ( ~x135 & n307 ) ;
  assign n309 = ( ~x7 & x135 ) | ( ~x7 & n308 ) | ( x135 & n308 ) ;
  assign n310 = ( ~n307 & n308 ) | ( ~n307 & n309 ) | ( n308 & n309 ) ;
  assign n311 = x7 & x135 ;
  assign n312 = x7 | x135 ;
  assign n313 = n304 & n312 ;
  assign n314 = n311 | n313 ;
  assign n315 = n311 | n312 ;
  assign n316 = ( n306 & n311 ) | ( n306 & n315 ) | ( n311 & n315 ) ;
  assign n317 = ( n300 & n314 ) | ( n300 & n316 ) | ( n314 & n316 ) ;
  assign n318 = ( x8 & ~x136 ) | ( x8 & n317 ) | ( ~x136 & n317 ) ;
  assign n319 = ( ~x8 & x136 ) | ( ~x8 & n318 ) | ( x136 & n318 ) ;
  assign n320 = ( ~n317 & n318 ) | ( ~n317 & n319 ) | ( n318 & n319 ) ;
  assign n321 = x9 | x137 ;
  assign n322 = x9 & x137 ;
  assign n323 = n321 | n322 ;
  assign n324 = x8 & x136 ;
  assign n325 = x8 | x136 ;
  assign n326 = n316 & n325 ;
  assign n327 = n311 & n325 ;
  assign n328 = ( n313 & n325 ) | ( n313 & n327 ) | ( n325 & n327 ) ;
  assign n329 = ( n300 & n326 ) | ( n300 & n328 ) | ( n326 & n328 ) ;
  assign n330 = n324 | n329 ;
  assign n331 = ( n322 & ~n323 ) | ( n322 & n330 ) | ( ~n323 & n330 ) ;
  assign n332 = ( n322 & n323 ) | ( n322 & n330 ) | ( n323 & n330 ) ;
  assign n333 = ( n323 & n331 ) | ( n323 & ~n332 ) | ( n331 & ~n332 ) ;
  assign n334 = ( x9 & x137 ) | ( x9 & n330 ) | ( x137 & n330 ) ;
  assign n335 = ( x10 & ~x138 ) | ( x10 & n334 ) | ( ~x138 & n334 ) ;
  assign n336 = ( ~x10 & x138 ) | ( ~x10 & n335 ) | ( x138 & n335 ) ;
  assign n337 = ( ~n334 & n335 ) | ( ~n334 & n336 ) | ( n335 & n336 ) ;
  assign n338 = x10 & x138 ;
  assign n339 = x10 | x138 ;
  assign n340 = n321 & n324 ;
  assign n341 = n322 & n339 ;
  assign n342 = ( n339 & n340 ) | ( n339 & n341 ) | ( n340 & n341 ) ;
  assign n343 = n338 | n342 ;
  assign n344 = n338 | n339 ;
  assign n345 = ( n323 & n338 ) | ( n323 & n344 ) | ( n338 & n344 ) ;
  assign n346 = ( n329 & n343 ) | ( n329 & n345 ) | ( n343 & n345 ) ;
  assign n347 = ( x11 & ~x139 ) | ( x11 & n346 ) | ( ~x139 & n346 ) ;
  assign n348 = ( ~x11 & x139 ) | ( ~x11 & n347 ) | ( x139 & n347 ) ;
  assign n349 = ( ~n346 & n347 ) | ( ~n346 & n348 ) | ( n347 & n348 ) ;
  assign n350 = x12 | x140 ;
  assign n351 = x12 & x140 ;
  assign n352 = n350 | n351 ;
  assign n353 = x11 & x139 ;
  assign n354 = x11 | x139 ;
  assign n355 = n345 & n354 ;
  assign n356 = n338 & n354 ;
  assign n357 = ( n342 & n354 ) | ( n342 & n356 ) | ( n354 & n356 ) ;
  assign n358 = ( n326 & n355 ) | ( n326 & n357 ) | ( n355 & n357 ) ;
  assign n359 = ( n328 & n355 ) | ( n328 & n357 ) | ( n355 & n357 ) ;
  assign n360 = ( n300 & n358 ) | ( n300 & n359 ) | ( n358 & n359 ) ;
  assign n361 = n353 | n360 ;
  assign n362 = ( n351 & ~n352 ) | ( n351 & n361 ) | ( ~n352 & n361 ) ;
  assign n363 = ( n351 & n352 ) | ( n351 & n361 ) | ( n352 & n361 ) ;
  assign n364 = ( n352 & n362 ) | ( n352 & ~n363 ) | ( n362 & ~n363 ) ;
  assign n365 = ( x12 & x140 ) | ( x12 & n361 ) | ( x140 & n361 ) ;
  assign n366 = ( x13 & ~x141 ) | ( x13 & n365 ) | ( ~x141 & n365 ) ;
  assign n367 = ( ~x13 & x141 ) | ( ~x13 & n366 ) | ( x141 & n366 ) ;
  assign n368 = ( ~n365 & n366 ) | ( ~n365 & n367 ) | ( n366 & n367 ) ;
  assign n369 = x14 | x142 ;
  assign n370 = x14 & x142 ;
  assign n371 = n369 & ~n370 ;
  assign n372 = x13 & x141 ;
  assign n373 = x13 | x141 ;
  assign n374 = n350 & n353 ;
  assign n375 = n351 & n373 ;
  assign n376 = ( n373 & n374 ) | ( n373 & n375 ) | ( n374 & n375 ) ;
  assign n377 = n372 | n376 ;
  assign n378 = n372 | n373 ;
  assign n379 = ( n352 & n372 ) | ( n352 & n378 ) | ( n372 & n378 ) ;
  assign n380 = ( n360 & n377 ) | ( n360 & n379 ) | ( n377 & n379 ) ;
  assign n381 = n371 | n380 ;
  assign n382 = n371 & n380 ;
  assign n383 = n381 & ~n382 ;
  assign n384 = n369 | n370 ;
  assign n385 = ( n370 & n379 ) | ( n370 & n384 ) | ( n379 & n384 ) ;
  assign n386 = ( x14 & x142 ) | ( x14 & n372 ) | ( x142 & n372 ) ;
  assign n387 = ( n369 & n376 ) | ( n369 & n386 ) | ( n376 & n386 ) ;
  assign n388 = ( n360 & n385 ) | ( n360 & n387 ) | ( n385 & n387 ) ;
  assign n389 = ( x15 & ~x143 ) | ( x15 & n388 ) | ( ~x143 & n388 ) ;
  assign n390 = ( ~x15 & x143 ) | ( ~x15 & n389 ) | ( x143 & n389 ) ;
  assign n391 = ( ~n388 & n389 ) | ( ~n388 & n390 ) | ( n389 & n390 ) ;
  assign n392 = x15 & x143 ;
  assign n393 = x15 | x143 ;
  assign n394 = n392 | n393 ;
  assign n395 = ( n388 & n392 ) | ( n388 & n394 ) | ( n392 & n394 ) ;
  assign n396 = ( x16 & ~x144 ) | ( x16 & n395 ) | ( ~x144 & n395 ) ;
  assign n397 = ( ~x16 & x144 ) | ( ~x16 & n396 ) | ( x144 & n396 ) ;
  assign n398 = ( ~n395 & n396 ) | ( ~n395 & n397 ) | ( n396 & n397 ) ;
  assign n399 = x16 & x144 ;
  assign n400 = x16 | x144 ;
  assign n401 = n392 & n400 ;
  assign n402 = n399 | n401 ;
  assign n403 = n399 | n400 ;
  assign n404 = ( n394 & n399 ) | ( n394 & n403 ) | ( n399 & n403 ) ;
  assign n405 = ( n388 & n402 ) | ( n388 & n404 ) | ( n402 & n404 ) ;
  assign n406 = ( x17 & ~x145 ) | ( x17 & n405 ) | ( ~x145 & n405 ) ;
  assign n407 = ( ~x17 & x145 ) | ( ~x17 & n406 ) | ( x145 & n406 ) ;
  assign n408 = ( ~n405 & n406 ) | ( ~n405 & n407 ) | ( n406 & n407 ) ;
  assign n409 = x17 & x145 ;
  assign n410 = x17 | x145 ;
  assign n411 = n399 & n410 ;
  assign n412 = ( n401 & n410 ) | ( n401 & n411 ) | ( n410 & n411 ) ;
  assign n413 = n409 | n412 ;
  assign n414 = n409 | n410 ;
  assign n415 = ( n404 & n409 ) | ( n404 & n414 ) | ( n409 & n414 ) ;
  assign n416 = ( n388 & n413 ) | ( n388 & n415 ) | ( n413 & n415 ) ;
  assign n417 = ( x18 & ~x146 ) | ( x18 & n416 ) | ( ~x146 & n416 ) ;
  assign n418 = ( ~x18 & x146 ) | ( ~x18 & n417 ) | ( x146 & n417 ) ;
  assign n419 = ( ~n416 & n417 ) | ( ~n416 & n418 ) | ( n417 & n418 ) ;
  assign n420 = x18 & x146 ;
  assign n421 = x18 | x146 ;
  assign n422 = n409 & n421 ;
  assign n423 = n414 & n421 ;
  assign n424 = ( n404 & n422 ) | ( n404 & n423 ) | ( n422 & n423 ) ;
  assign n425 = n420 | n424 ;
  assign n426 = n420 | n422 ;
  assign n427 = n420 | n421 ;
  assign n428 = ( n412 & n426 ) | ( n412 & n427 ) | ( n426 & n427 ) ;
  assign n429 = ( n385 & n425 ) | ( n385 & n428 ) | ( n425 & n428 ) ;
  assign n430 = ( n387 & n425 ) | ( n387 & n428 ) | ( n425 & n428 ) ;
  assign n431 = ( n360 & n429 ) | ( n360 & n430 ) | ( n429 & n430 ) ;
  assign n432 = ( x19 & ~x147 ) | ( x19 & n431 ) | ( ~x147 & n431 ) ;
  assign n433 = ( ~x19 & x147 ) | ( ~x19 & n432 ) | ( x147 & n432 ) ;
  assign n434 = ( ~n431 & n432 ) | ( ~n431 & n433 ) | ( n432 & n433 ) ;
  assign n435 = x19 & x147 ;
  assign n436 = x19 | x147 ;
  assign n437 = n435 | n436 ;
  assign n438 = ( n431 & n435 ) | ( n431 & n437 ) | ( n435 & n437 ) ;
  assign n439 = ( x20 & ~x148 ) | ( x20 & n438 ) | ( ~x148 & n438 ) ;
  assign n440 = ( ~x20 & x148 ) | ( ~x20 & n439 ) | ( x148 & n439 ) ;
  assign n441 = ( ~n438 & n439 ) | ( ~n438 & n440 ) | ( n439 & n440 ) ;
  assign n442 = x20 & x148 ;
  assign n443 = x20 | x148 ;
  assign n444 = n435 & n443 ;
  assign n445 = n442 | n444 ;
  assign n446 = n442 | n443 ;
  assign n447 = ( n437 & n442 ) | ( n437 & n446 ) | ( n442 & n446 ) ;
  assign n448 = ( n431 & n445 ) | ( n431 & n447 ) | ( n445 & n447 ) ;
  assign n449 = ( x21 & ~x149 ) | ( x21 & n448 ) | ( ~x149 & n448 ) ;
  assign n450 = ( ~x21 & x149 ) | ( ~x21 & n449 ) | ( x149 & n449 ) ;
  assign n451 = ( ~n448 & n449 ) | ( ~n448 & n450 ) | ( n449 & n450 ) ;
  assign n452 = x21 & x149 ;
  assign n453 = x21 | x149 ;
  assign n454 = n442 & n453 ;
  assign n455 = ( n444 & n453 ) | ( n444 & n454 ) | ( n453 & n454 ) ;
  assign n456 = n452 | n455 ;
  assign n457 = n452 | n453 ;
  assign n458 = ( n447 & n452 ) | ( n447 & n457 ) | ( n452 & n457 ) ;
  assign n459 = ( n431 & n456 ) | ( n431 & n458 ) | ( n456 & n458 ) ;
  assign n460 = ( x22 & ~x150 ) | ( x22 & n459 ) | ( ~x150 & n459 ) ;
  assign n461 = ( ~x22 & x150 ) | ( ~x22 & n460 ) | ( x150 & n460 ) ;
  assign n462 = ( ~n459 & n460 ) | ( ~n459 & n461 ) | ( n460 & n461 ) ;
  assign n463 = x22 & x150 ;
  assign n464 = x22 | x150 ;
  assign n465 = n452 & n464 ;
  assign n466 = n457 & n464 ;
  assign n467 = ( n447 & n465 ) | ( n447 & n466 ) | ( n465 & n466 ) ;
  assign n468 = n463 | n467 ;
  assign n469 = n463 | n465 ;
  assign n470 = n463 | n464 ;
  assign n471 = ( n455 & n469 ) | ( n455 & n470 ) | ( n469 & n470 ) ;
  assign n472 = ( n431 & n468 ) | ( n431 & n471 ) | ( n468 & n471 ) ;
  assign n473 = ( x23 & ~x151 ) | ( x23 & n472 ) | ( ~x151 & n472 ) ;
  assign n474 = ( ~x23 & x151 ) | ( ~x23 & n473 ) | ( x151 & n473 ) ;
  assign n475 = ( ~n472 & n473 ) | ( ~n472 & n474 ) | ( n473 & n474 ) ;
  assign n476 = x24 | x152 ;
  assign n477 = x24 & x152 ;
  assign n478 = n476 | n477 ;
  assign n479 = x23 & x151 ;
  assign n480 = x23 | x151 ;
  assign n481 = n471 & n480 ;
  assign n482 = n463 & n480 ;
  assign n483 = ( n467 & n480 ) | ( n467 & n482 ) | ( n480 & n482 ) ;
  assign n484 = ( n431 & n481 ) | ( n431 & n483 ) | ( n481 & n483 ) ;
  assign n485 = n479 | n484 ;
  assign n486 = ( n477 & ~n478 ) | ( n477 & n485 ) | ( ~n478 & n485 ) ;
  assign n487 = ( n477 & n478 ) | ( n477 & n485 ) | ( n478 & n485 ) ;
  assign n488 = ( n478 & n486 ) | ( n478 & ~n487 ) | ( n486 & ~n487 ) ;
  assign n489 = ( x24 & x152 ) | ( x24 & n485 ) | ( x152 & n485 ) ;
  assign n490 = ( x25 & ~x153 ) | ( x25 & n489 ) | ( ~x153 & n489 ) ;
  assign n491 = ( ~x25 & x153 ) | ( ~x25 & n490 ) | ( x153 & n490 ) ;
  assign n492 = ( ~n489 & n490 ) | ( ~n489 & n491 ) | ( n490 & n491 ) ;
  assign n493 = x26 | x154 ;
  assign n494 = x26 & x154 ;
  assign n495 = n493 & ~n494 ;
  assign n496 = x25 & x153 ;
  assign n497 = x25 | x153 ;
  assign n498 = n476 & n479 ;
  assign n499 = n477 & n497 ;
  assign n500 = ( n497 & n498 ) | ( n497 & n499 ) | ( n498 & n499 ) ;
  assign n501 = n496 | n500 ;
  assign n502 = n496 | n497 ;
  assign n503 = ( n478 & n496 ) | ( n478 & n502 ) | ( n496 & n502 ) ;
  assign n504 = ( n484 & n501 ) | ( n484 & n503 ) | ( n501 & n503 ) ;
  assign n505 = n495 | n504 ;
  assign n506 = n495 & n504 ;
  assign n507 = n505 & ~n506 ;
  assign n508 = n493 | n494 ;
  assign n509 = ( n494 & n503 ) | ( n494 & n508 ) | ( n503 & n508 ) ;
  assign n510 = ( x26 & x154 ) | ( x26 & n496 ) | ( x154 & n496 ) ;
  assign n511 = ( n493 & n500 ) | ( n493 & n510 ) | ( n500 & n510 ) ;
  assign n512 = ( n484 & n509 ) | ( n484 & n511 ) | ( n509 & n511 ) ;
  assign n513 = ( x27 & ~x155 ) | ( x27 & n512 ) | ( ~x155 & n512 ) ;
  assign n514 = ( ~x27 & x155 ) | ( ~x27 & n513 ) | ( x155 & n513 ) ;
  assign n515 = ( ~n512 & n513 ) | ( ~n512 & n514 ) | ( n513 & n514 ) ;
  assign n516 = x27 & x155 ;
  assign n517 = x27 | x155 ;
  assign n518 = n508 & n517 ;
  assign n519 = n494 & n517 ;
  assign n520 = ( n503 & n518 ) | ( n503 & n519 ) | ( n518 & n519 ) ;
  assign n521 = n516 | n520 ;
  assign n522 = n516 | n517 ;
  assign n523 = ( n510 & n516 ) | ( n510 & n522 ) | ( n516 & n522 ) ;
  assign n524 = ( n493 & n516 ) | ( n493 & n522 ) | ( n516 & n522 ) ;
  assign n525 = ( n500 & n523 ) | ( n500 & n524 ) | ( n523 & n524 ) ;
  assign n526 = ( n484 & n521 ) | ( n484 & n525 ) | ( n521 & n525 ) ;
  assign n527 = ( x28 & ~x156 ) | ( x28 & n526 ) | ( ~x156 & n526 ) ;
  assign n528 = ( ~x28 & x156 ) | ( ~x28 & n527 ) | ( x156 & n527 ) ;
  assign n529 = ( ~n526 & n527 ) | ( ~n526 & n528 ) | ( n527 & n528 ) ;
  assign n530 = x29 | x157 ;
  assign n531 = x29 & x157 ;
  assign n532 = n530 | n531 ;
  assign n533 = x28 & x156 ;
  assign n534 = x28 | x156 ;
  assign n535 = n516 & n534 ;
  assign n536 = ( n520 & n534 ) | ( n520 & n535 ) | ( n534 & n535 ) ;
  assign n537 = n525 & n534 ;
  assign n538 = ( n483 & n536 ) | ( n483 & n537 ) | ( n536 & n537 ) ;
  assign n539 = ( n481 & n536 ) | ( n481 & n537 ) | ( n536 & n537 ) ;
  assign n540 = ( n431 & n538 ) | ( n431 & n539 ) | ( n538 & n539 ) ;
  assign n541 = n533 | n540 ;
  assign n542 = ( n531 & ~n532 ) | ( n531 & n541 ) | ( ~n532 & n541 ) ;
  assign n543 = ( n531 & n532 ) | ( n531 & n541 ) | ( n532 & n541 ) ;
  assign n544 = ( n532 & n542 ) | ( n532 & ~n543 ) | ( n542 & ~n543 ) ;
  assign n545 = ( x29 & x157 ) | ( x29 & n541 ) | ( x157 & n541 ) ;
  assign n546 = ( x30 & ~x158 ) | ( x30 & n545 ) | ( ~x158 & n545 ) ;
  assign n547 = ( ~x30 & x158 ) | ( ~x30 & n546 ) | ( x158 & n546 ) ;
  assign n548 = ( ~n545 & n546 ) | ( ~n545 & n547 ) | ( n546 & n547 ) ;
  assign n549 = x31 | x159 ;
  assign n550 = x31 & x159 ;
  assign n551 = n549 & ~n550 ;
  assign n552 = x30 & x158 ;
  assign n553 = x30 | x158 ;
  assign n554 = n530 & n533 ;
  assign n555 = n531 & n553 ;
  assign n556 = ( n553 & n554 ) | ( n553 & n555 ) | ( n554 & n555 ) ;
  assign n557 = n552 | n556 ;
  assign n558 = n552 | n553 ;
  assign n559 = ( n532 & n552 ) | ( n532 & n558 ) | ( n552 & n558 ) ;
  assign n560 = ( n540 & n557 ) | ( n540 & n559 ) | ( n557 & n559 ) ;
  assign n561 = n551 | n560 ;
  assign n562 = n551 & n560 ;
  assign n563 = n561 & ~n562 ;
  assign n564 = n549 | n550 ;
  assign n565 = ( n550 & n559 ) | ( n550 & n564 ) | ( n559 & n564 ) ;
  assign n566 = ( x31 & x159 ) | ( x31 & n552 ) | ( x159 & n552 ) ;
  assign n567 = ( n549 & n556 ) | ( n549 & n566 ) | ( n556 & n566 ) ;
  assign n568 = ( n540 & n565 ) | ( n540 & n567 ) | ( n565 & n567 ) ;
  assign n569 = ( x32 & ~x160 ) | ( x32 & n568 ) | ( ~x160 & n568 ) ;
  assign n570 = ( ~x32 & x160 ) | ( ~x32 & n569 ) | ( x160 & n569 ) ;
  assign n571 = ( ~n568 & n569 ) | ( ~n568 & n570 ) | ( n569 & n570 ) ;
  assign n572 = x32 & x160 ;
  assign n573 = x32 | x160 ;
  assign n574 = n564 & n573 ;
  assign n575 = n550 & n573 ;
  assign n576 = ( n559 & n574 ) | ( n559 & n575 ) | ( n574 & n575 ) ;
  assign n577 = n572 | n576 ;
  assign n578 = n572 | n573 ;
  assign n579 = ( n567 & n572 ) | ( n567 & n578 ) | ( n572 & n578 ) ;
  assign n580 = ( n540 & n577 ) | ( n540 & n579 ) | ( n577 & n579 ) ;
  assign n581 = ( x33 & ~x161 ) | ( x33 & n580 ) | ( ~x161 & n580 ) ;
  assign n582 = ( ~x33 & x161 ) | ( ~x33 & n581 ) | ( x161 & n581 ) ;
  assign n583 = ( ~n580 & n581 ) | ( ~n580 & n582 ) | ( n581 & n582 ) ;
  assign n584 = x33 & x161 ;
  assign n585 = x33 | x161 ;
  assign n586 = n572 & n585 ;
  assign n587 = n584 | n586 ;
  assign n588 = n584 | n585 ;
  assign n589 = ( n578 & n584 ) | ( n578 & n588 ) | ( n584 & n588 ) ;
  assign n590 = ( n567 & n587 ) | ( n567 & n589 ) | ( n587 & n589 ) ;
  assign n591 = ( n576 & n587 ) | ( n576 & n588 ) | ( n587 & n588 ) ;
  assign n592 = ( n539 & n590 ) | ( n539 & n591 ) | ( n590 & n591 ) ;
  assign n593 = ( n538 & n590 ) | ( n538 & n591 ) | ( n590 & n591 ) ;
  assign n594 = ( n431 & n592 ) | ( n431 & n593 ) | ( n592 & n593 ) ;
  assign n595 = ( x34 & ~x162 ) | ( x34 & n594 ) | ( ~x162 & n594 ) ;
  assign n596 = ( ~x34 & x162 ) | ( ~x34 & n595 ) | ( x162 & n595 ) ;
  assign n597 = ( ~n594 & n595 ) | ( ~n594 & n596 ) | ( n595 & n596 ) ;
  assign n598 = x34 & x162 ;
  assign n599 = x34 | x162 ;
  assign n600 = n598 | n599 ;
  assign n601 = ( n594 & n598 ) | ( n594 & n600 ) | ( n598 & n600 ) ;
  assign n602 = ( x35 & ~x163 ) | ( x35 & n601 ) | ( ~x163 & n601 ) ;
  assign n603 = ( ~x35 & x163 ) | ( ~x35 & n602 ) | ( x163 & n602 ) ;
  assign n604 = ( ~n601 & n602 ) | ( ~n601 & n603 ) | ( n602 & n603 ) ;
  assign n605 = x35 & x163 ;
  assign n606 = x35 | x163 ;
  assign n607 = n598 & n606 ;
  assign n608 = n605 | n607 ;
  assign n609 = n605 | n606 ;
  assign n610 = ( n600 & n605 ) | ( n600 & n609 ) | ( n605 & n609 ) ;
  assign n611 = ( n594 & n608 ) | ( n594 & n610 ) | ( n608 & n610 ) ;
  assign n612 = ( x36 & ~x164 ) | ( x36 & n611 ) | ( ~x164 & n611 ) ;
  assign n613 = ( ~x36 & x164 ) | ( ~x36 & n612 ) | ( x164 & n612 ) ;
  assign n614 = ( ~n611 & n612 ) | ( ~n611 & n613 ) | ( n612 & n613 ) ;
  assign n615 = x36 & x164 ;
  assign n616 = x36 | x164 ;
  assign n617 = n605 & n616 ;
  assign n618 = ( n607 & n616 ) | ( n607 & n617 ) | ( n616 & n617 ) ;
  assign n619 = n615 | n618 ;
  assign n620 = n615 | n616 ;
  assign n621 = ( n610 & n615 ) | ( n610 & n620 ) | ( n615 & n620 ) ;
  assign n622 = ( n594 & n619 ) | ( n594 & n621 ) | ( n619 & n621 ) ;
  assign n623 = ( x37 & ~x165 ) | ( x37 & n622 ) | ( ~x165 & n622 ) ;
  assign n624 = ( ~x37 & x165 ) | ( ~x37 & n623 ) | ( x165 & n623 ) ;
  assign n625 = ( ~n622 & n623 ) | ( ~n622 & n624 ) | ( n623 & n624 ) ;
  assign n626 = x37 & x165 ;
  assign n627 = x37 | x165 ;
  assign n628 = n615 & n627 ;
  assign n629 = n620 & n627 ;
  assign n630 = ( n610 & n628 ) | ( n610 & n629 ) | ( n628 & n629 ) ;
  assign n631 = n626 | n630 ;
  assign n632 = n626 | n628 ;
  assign n633 = n626 | n627 ;
  assign n634 = ( n618 & n632 ) | ( n618 & n633 ) | ( n632 & n633 ) ;
  assign n635 = ( n594 & n631 ) | ( n594 & n634 ) | ( n631 & n634 ) ;
  assign n636 = ( x38 & ~x166 ) | ( x38 & n635 ) | ( ~x166 & n635 ) ;
  assign n637 = ( ~x38 & x166 ) | ( ~x38 & n636 ) | ( x166 & n636 ) ;
  assign n638 = ( ~n635 & n636 ) | ( ~n635 & n637 ) | ( n636 & n637 ) ;
  assign n639 = x38 & x166 ;
  assign n640 = x38 | x166 ;
  assign n641 = n626 & n640 ;
  assign n642 = n639 | n641 ;
  assign n643 = n639 | n640 ;
  assign n644 = ( n630 & n642 ) | ( n630 & n643 ) | ( n642 & n643 ) ;
  assign n645 = ( n634 & n639 ) | ( n634 & n643 ) | ( n639 & n643 ) ;
  assign n646 = ( n594 & n644 ) | ( n594 & n645 ) | ( n644 & n645 ) ;
  assign n647 = ( x39 & ~x167 ) | ( x39 & n646 ) | ( ~x167 & n646 ) ;
  assign n648 = ( ~x39 & x167 ) | ( ~x39 & n647 ) | ( x167 & n647 ) ;
  assign n649 = ( ~n646 & n647 ) | ( ~n646 & n648 ) | ( n647 & n648 ) ;
  assign n650 = x39 & x167 ;
  assign n651 = x39 | x167 ;
  assign n652 = n643 & n651 ;
  assign n653 = n642 & n651 ;
  assign n654 = ( n630 & n652 ) | ( n630 & n653 ) | ( n652 & n653 ) ;
  assign n655 = n650 | n654 ;
  assign n656 = n650 | n652 ;
  assign n657 = n639 & n651 ;
  assign n658 = n650 | n657 ;
  assign n659 = ( n634 & n656 ) | ( n634 & n658 ) | ( n656 & n658 ) ;
  assign n660 = ( n594 & n655 ) | ( n594 & n659 ) | ( n655 & n659 ) ;
  assign n661 = ( x40 & ~x168 ) | ( x40 & n660 ) | ( ~x168 & n660 ) ;
  assign n662 = ( ~x40 & x168 ) | ( ~x40 & n661 ) | ( x168 & n661 ) ;
  assign n663 = ( ~n660 & n661 ) | ( ~n660 & n662 ) | ( n661 & n662 ) ;
  assign n664 = x40 & x168 ;
  assign n665 = x40 | x168 ;
  assign n666 = n664 | n665 ;
  assign n667 = ( n660 & n664 ) | ( n660 & n666 ) | ( n664 & n666 ) ;
  assign n668 = ( x41 & ~x169 ) | ( x41 & n667 ) | ( ~x169 & n667 ) ;
  assign n669 = ( ~x41 & x169 ) | ( ~x41 & n668 ) | ( x169 & n668 ) ;
  assign n670 = ( ~n667 & n668 ) | ( ~n667 & n669 ) | ( n668 & n669 ) ;
  assign n671 = x41 & x169 ;
  assign n672 = x41 | x169 ;
  assign n673 = n664 & n672 ;
  assign n674 = n671 | n673 ;
  assign n675 = n671 | n672 ;
  assign n676 = ( n666 & n671 ) | ( n666 & n675 ) | ( n671 & n675 ) ;
  assign n677 = ( n660 & n674 ) | ( n660 & n676 ) | ( n674 & n676 ) ;
  assign n678 = ( x42 & ~x170 ) | ( x42 & n677 ) | ( ~x170 & n677 ) ;
  assign n679 = ( ~x42 & x170 ) | ( ~x42 & n678 ) | ( x170 & n678 ) ;
  assign n680 = ( ~n677 & n678 ) | ( ~n677 & n679 ) | ( n678 & n679 ) ;
  assign n681 = x42 & x170 ;
  assign n682 = x42 | x170 ;
  assign n683 = n671 & n682 ;
  assign n684 = ( n673 & n682 ) | ( n673 & n683 ) | ( n682 & n683 ) ;
  assign n685 = n681 | n684 ;
  assign n686 = n681 | n682 ;
  assign n687 = ( n676 & n681 ) | ( n676 & n686 ) | ( n681 & n686 ) ;
  assign n688 = ( n660 & n685 ) | ( n660 & n687 ) | ( n685 & n687 ) ;
  assign n689 = ( x43 & ~x171 ) | ( x43 & n688 ) | ( ~x171 & n688 ) ;
  assign n690 = ( ~x43 & x171 ) | ( ~x43 & n689 ) | ( x171 & n689 ) ;
  assign n691 = ( ~n688 & n689 ) | ( ~n688 & n690 ) | ( n689 & n690 ) ;
  assign n692 = x43 & x171 ;
  assign n693 = x43 | x171 ;
  assign n694 = n681 & n693 ;
  assign n695 = n686 & n693 ;
  assign n696 = ( n676 & n694 ) | ( n676 & n695 ) | ( n694 & n695 ) ;
  assign n697 = n692 | n696 ;
  assign n698 = n692 | n694 ;
  assign n699 = n692 | n693 ;
  assign n700 = ( n684 & n698 ) | ( n684 & n699 ) | ( n698 & n699 ) ;
  assign n701 = ( n660 & n697 ) | ( n660 & n700 ) | ( n697 & n700 ) ;
  assign n702 = ( x44 & ~x172 ) | ( x44 & n701 ) | ( ~x172 & n701 ) ;
  assign n703 = ( ~x44 & x172 ) | ( ~x44 & n702 ) | ( x172 & n702 ) ;
  assign n704 = ( ~n701 & n702 ) | ( ~n701 & n703 ) | ( n702 & n703 ) ;
  assign n705 = x44 & x172 ;
  assign n706 = x44 | x172 ;
  assign n707 = n692 & n706 ;
  assign n708 = n705 | n707 ;
  assign n709 = n705 | n706 ;
  assign n710 = ( n696 & n708 ) | ( n696 & n709 ) | ( n708 & n709 ) ;
  assign n711 = ( n700 & n705 ) | ( n700 & n709 ) | ( n705 & n709 ) ;
  assign n712 = ( n660 & n710 ) | ( n660 & n711 ) | ( n710 & n711 ) ;
  assign n713 = ( x45 & ~x173 ) | ( x45 & n712 ) | ( ~x173 & n712 ) ;
  assign n714 = ( ~x45 & x173 ) | ( ~x45 & n713 ) | ( x173 & n713 ) ;
  assign n715 = ( ~n712 & n713 ) | ( ~n712 & n714 ) | ( n713 & n714 ) ;
  assign n716 = x45 & x173 ;
  assign n717 = x45 | x173 ;
  assign n718 = n709 & n717 ;
  assign n719 = n708 & n717 ;
  assign n720 = ( n696 & n718 ) | ( n696 & n719 ) | ( n718 & n719 ) ;
  assign n721 = n716 | n720 ;
  assign n722 = n716 | n718 ;
  assign n723 = n705 & n717 ;
  assign n724 = n716 | n723 ;
  assign n725 = ( n700 & n722 ) | ( n700 & n724 ) | ( n722 & n724 ) ;
  assign n726 = ( n660 & n721 ) | ( n660 & n725 ) | ( n721 & n725 ) ;
  assign n727 = ( x46 & ~x174 ) | ( x46 & n726 ) | ( ~x174 & n726 ) ;
  assign n728 = ( ~x46 & x174 ) | ( ~x46 & n727 ) | ( x174 & n727 ) ;
  assign n729 = ( ~n726 & n727 ) | ( ~n726 & n728 ) | ( n727 & n728 ) ;
  assign n730 = x47 | x175 ;
  assign n731 = x47 & x175 ;
  assign n732 = n730 | n731 ;
  assign n733 = x46 & x174 ;
  assign n734 = x46 | x174 ;
  assign n735 = n725 & n734 ;
  assign n736 = n716 & n734 ;
  assign n737 = ( n720 & n734 ) | ( n720 & n736 ) | ( n734 & n736 ) ;
  assign n738 = ( n655 & n735 ) | ( n655 & n737 ) | ( n735 & n737 ) ;
  assign n739 = ( n659 & n735 ) | ( n659 & n737 ) | ( n735 & n737 ) ;
  assign n740 = ( n594 & n738 ) | ( n594 & n739 ) | ( n738 & n739 ) ;
  assign n741 = n733 | n740 ;
  assign n742 = ( n731 & ~n732 ) | ( n731 & n741 ) | ( ~n732 & n741 ) ;
  assign n743 = ( n731 & n732 ) | ( n731 & n741 ) | ( n732 & n741 ) ;
  assign n744 = ( n732 & n742 ) | ( n732 & ~n743 ) | ( n742 & ~n743 ) ;
  assign n745 = ( x47 & x175 ) | ( x47 & n741 ) | ( x175 & n741 ) ;
  assign n746 = ( x48 & ~x176 ) | ( x48 & n745 ) | ( ~x176 & n745 ) ;
  assign n747 = ( ~x48 & x176 ) | ( ~x48 & n746 ) | ( x176 & n746 ) ;
  assign n748 = ( ~n745 & n746 ) | ( ~n745 & n747 ) | ( n746 & n747 ) ;
  assign n749 = x49 | x177 ;
  assign n750 = x49 & x177 ;
  assign n751 = n749 & ~n750 ;
  assign n752 = x48 & x176 ;
  assign n753 = x48 | x176 ;
  assign n754 = n730 & n733 ;
  assign n755 = n731 & n753 ;
  assign n756 = ( n753 & n754 ) | ( n753 & n755 ) | ( n754 & n755 ) ;
  assign n757 = n752 | n756 ;
  assign n758 = n752 | n753 ;
  assign n759 = ( n732 & n752 ) | ( n732 & n758 ) | ( n752 & n758 ) ;
  assign n760 = ( n740 & n757 ) | ( n740 & n759 ) | ( n757 & n759 ) ;
  assign n761 = n751 | n760 ;
  assign n762 = n751 & n760 ;
  assign n763 = n761 & ~n762 ;
  assign n764 = n749 | n750 ;
  assign n765 = ( n750 & n759 ) | ( n750 & n764 ) | ( n759 & n764 ) ;
  assign n766 = ( x49 & x177 ) | ( x49 & n752 ) | ( x177 & n752 ) ;
  assign n767 = ( n749 & n756 ) | ( n749 & n766 ) | ( n756 & n766 ) ;
  assign n768 = ( n740 & n765 ) | ( n740 & n767 ) | ( n765 & n767 ) ;
  assign n769 = ( x50 & ~x178 ) | ( x50 & n768 ) | ( ~x178 & n768 ) ;
  assign n770 = ( ~x50 & x178 ) | ( ~x50 & n769 ) | ( x178 & n769 ) ;
  assign n771 = ( ~n768 & n769 ) | ( ~n768 & n770 ) | ( n769 & n770 ) ;
  assign n772 = x50 & x178 ;
  assign n773 = x50 | x178 ;
  assign n774 = n764 & n773 ;
  assign n775 = n750 & n773 ;
  assign n776 = ( n759 & n774 ) | ( n759 & n775 ) | ( n774 & n775 ) ;
  assign n777 = n772 | n776 ;
  assign n778 = n772 | n773 ;
  assign n779 = ( n767 & n772 ) | ( n767 & n778 ) | ( n772 & n778 ) ;
  assign n780 = ( n740 & n777 ) | ( n740 & n779 ) | ( n777 & n779 ) ;
  assign n781 = ( x51 & ~x179 ) | ( x51 & n780 ) | ( ~x179 & n780 ) ;
  assign n782 = ( ~x51 & x179 ) | ( ~x51 & n781 ) | ( x179 & n781 ) ;
  assign n783 = ( ~n780 & n781 ) | ( ~n780 & n782 ) | ( n781 & n782 ) ;
  assign n784 = x51 & x179 ;
  assign n785 = x51 | x179 ;
  assign n786 = n772 & n785 ;
  assign n787 = n784 | n786 ;
  assign n788 = n784 | n785 ;
  assign n789 = ( n778 & n784 ) | ( n778 & n788 ) | ( n784 & n788 ) ;
  assign n790 = ( n767 & n787 ) | ( n767 & n789 ) | ( n787 & n789 ) ;
  assign n791 = ( n776 & n787 ) | ( n776 & n788 ) | ( n787 & n788 ) ;
  assign n792 = ( n740 & n790 ) | ( n740 & n791 ) | ( n790 & n791 ) ;
  assign n793 = ( x52 & ~x180 ) | ( x52 & n792 ) | ( ~x180 & n792 ) ;
  assign n794 = ( ~x52 & x180 ) | ( ~x52 & n793 ) | ( x180 & n793 ) ;
  assign n795 = ( ~n792 & n793 ) | ( ~n792 & n794 ) | ( n793 & n794 ) ;
  assign n796 = x52 & x180 ;
  assign n797 = x52 | x180 ;
  assign n798 = n787 & n797 ;
  assign n799 = n788 & n797 ;
  assign n800 = ( n776 & n798 ) | ( n776 & n799 ) | ( n798 & n799 ) ;
  assign n801 = n796 | n800 ;
  assign n802 = n796 | n797 ;
  assign n803 = ( n789 & n796 ) | ( n789 & n802 ) | ( n796 & n802 ) ;
  assign n804 = ( n787 & n796 ) | ( n787 & n802 ) | ( n796 & n802 ) ;
  assign n805 = ( n767 & n803 ) | ( n767 & n804 ) | ( n803 & n804 ) ;
  assign n806 = ( n740 & n801 ) | ( n740 & n805 ) | ( n801 & n805 ) ;
  assign n807 = ( x53 & ~x181 ) | ( x53 & n806 ) | ( ~x181 & n806 ) ;
  assign n808 = ( ~x53 & x181 ) | ( ~x53 & n807 ) | ( x181 & n807 ) ;
  assign n809 = ( ~n806 & n807 ) | ( ~n806 & n808 ) | ( n807 & n808 ) ;
  assign n810 = x54 | x182 ;
  assign n811 = x54 & x182 ;
  assign n812 = n810 | n811 ;
  assign n813 = x53 & x181 ;
  assign n814 = x53 | x181 ;
  assign n815 = n796 & n814 ;
  assign n816 = ( n800 & n814 ) | ( n800 & n815 ) | ( n814 & n815 ) ;
  assign n817 = n805 & n814 ;
  assign n818 = ( n739 & n816 ) | ( n739 & n817 ) | ( n816 & n817 ) ;
  assign n819 = ( n738 & n816 ) | ( n738 & n817 ) | ( n816 & n817 ) ;
  assign n820 = ( n594 & n818 ) | ( n594 & n819 ) | ( n818 & n819 ) ;
  assign n821 = n813 | n820 ;
  assign n822 = ( n811 & ~n812 ) | ( n811 & n821 ) | ( ~n812 & n821 ) ;
  assign n823 = ( n811 & n812 ) | ( n811 & n821 ) | ( n812 & n821 ) ;
  assign n824 = ( n812 & n822 ) | ( n812 & ~n823 ) | ( n822 & ~n823 ) ;
  assign n825 = ( x54 & x182 ) | ( x54 & n821 ) | ( x182 & n821 ) ;
  assign n826 = ( x55 & ~x183 ) | ( x55 & n825 ) | ( ~x183 & n825 ) ;
  assign n827 = ( ~x55 & x183 ) | ( ~x55 & n826 ) | ( x183 & n826 ) ;
  assign n828 = ( ~n825 & n826 ) | ( ~n825 & n827 ) | ( n826 & n827 ) ;
  assign n829 = x56 | x184 ;
  assign n830 = x56 & x184 ;
  assign n831 = n829 & ~n830 ;
  assign n832 = x55 & x183 ;
  assign n833 = x55 | x183 ;
  assign n834 = n810 & n813 ;
  assign n835 = n811 & n833 ;
  assign n836 = ( n833 & n834 ) | ( n833 & n835 ) | ( n834 & n835 ) ;
  assign n837 = n832 | n836 ;
  assign n838 = n832 | n833 ;
  assign n839 = ( n812 & n832 ) | ( n812 & n838 ) | ( n832 & n838 ) ;
  assign n840 = ( n820 & n837 ) | ( n820 & n839 ) | ( n837 & n839 ) ;
  assign n841 = n831 | n840 ;
  assign n842 = n831 & n840 ;
  assign n843 = n841 & ~n842 ;
  assign n844 = n829 | n830 ;
  assign n845 = ( n830 & n839 ) | ( n830 & n844 ) | ( n839 & n844 ) ;
  assign n846 = ( x56 & x184 ) | ( x56 & n832 ) | ( x184 & n832 ) ;
  assign n847 = ( n829 & n836 ) | ( n829 & n846 ) | ( n836 & n846 ) ;
  assign n848 = ( n820 & n845 ) | ( n820 & n847 ) | ( n845 & n847 ) ;
  assign n849 = ( x57 & ~x185 ) | ( x57 & n848 ) | ( ~x185 & n848 ) ;
  assign n850 = ( ~x57 & x185 ) | ( ~x57 & n849 ) | ( x185 & n849 ) ;
  assign n851 = ( ~n848 & n849 ) | ( ~n848 & n850 ) | ( n849 & n850 ) ;
  assign n852 = x57 & x185 ;
  assign n853 = x57 | x185 ;
  assign n854 = n844 & n853 ;
  assign n855 = n830 & n853 ;
  assign n856 = ( n839 & n854 ) | ( n839 & n855 ) | ( n854 & n855 ) ;
  assign n857 = n852 | n856 ;
  assign n858 = n852 | n853 ;
  assign n859 = ( n847 & n852 ) | ( n847 & n858 ) | ( n852 & n858 ) ;
  assign n860 = ( n820 & n857 ) | ( n820 & n859 ) | ( n857 & n859 ) ;
  assign n861 = ( x58 & ~x186 ) | ( x58 & n860 ) | ( ~x186 & n860 ) ;
  assign n862 = ( ~x58 & x186 ) | ( ~x58 & n861 ) | ( x186 & n861 ) ;
  assign n863 = ( ~n860 & n861 ) | ( ~n860 & n862 ) | ( n861 & n862 ) ;
  assign n864 = x58 & x186 ;
  assign n865 = x58 | x186 ;
  assign n866 = n852 & n865 ;
  assign n867 = n864 | n866 ;
  assign n868 = n864 | n865 ;
  assign n869 = ( n858 & n864 ) | ( n858 & n868 ) | ( n864 & n868 ) ;
  assign n870 = ( n847 & n867 ) | ( n847 & n869 ) | ( n867 & n869 ) ;
  assign n871 = ( n856 & n867 ) | ( n856 & n868 ) | ( n867 & n868 ) ;
  assign n872 = ( n820 & n870 ) | ( n820 & n871 ) | ( n870 & n871 ) ;
  assign n873 = ( x59 & ~x187 ) | ( x59 & n872 ) | ( ~x187 & n872 ) ;
  assign n874 = ( ~x59 & x187 ) | ( ~x59 & n873 ) | ( x187 & n873 ) ;
  assign n875 = ( ~n872 & n873 ) | ( ~n872 & n874 ) | ( n873 & n874 ) ;
  assign n876 = x59 & x187 ;
  assign n877 = x59 | x187 ;
  assign n878 = n867 & n877 ;
  assign n879 = n868 & n877 ;
  assign n880 = ( n856 & n878 ) | ( n856 & n879 ) | ( n878 & n879 ) ;
  assign n881 = n876 | n880 ;
  assign n882 = n876 | n877 ;
  assign n883 = ( n870 & n876 ) | ( n870 & n882 ) | ( n876 & n882 ) ;
  assign n884 = ( n820 & n881 ) | ( n820 & n883 ) | ( n881 & n883 ) ;
  assign n885 = ( x60 & ~x188 ) | ( x60 & n884 ) | ( ~x188 & n884 ) ;
  assign n886 = ( ~x60 & x188 ) | ( ~x60 & n885 ) | ( x188 & n885 ) ;
  assign n887 = ( ~n884 & n885 ) | ( ~n884 & n886 ) | ( n885 & n886 ) ;
  assign n888 = x60 & x188 ;
  assign n889 = x60 | x188 ;
  assign n890 = n876 & n889 ;
  assign n891 = n888 | n890 ;
  assign n892 = n888 | n889 ;
  assign n893 = ( n880 & n891 ) | ( n880 & n892 ) | ( n891 & n892 ) ;
  assign n894 = ( n882 & n888 ) | ( n882 & n892 ) | ( n888 & n892 ) ;
  assign n895 = ( n869 & n891 ) | ( n869 & n894 ) | ( n891 & n894 ) ;
  assign n896 = ( n867 & n891 ) | ( n867 & n894 ) | ( n891 & n894 ) ;
  assign n897 = ( n847 & n895 ) | ( n847 & n896 ) | ( n895 & n896 ) ;
  assign n898 = ( n820 & n893 ) | ( n820 & n897 ) | ( n893 & n897 ) ;
  assign n899 = ( x61 & ~x189 ) | ( x61 & n898 ) | ( ~x189 & n898 ) ;
  assign n900 = ( ~x61 & x189 ) | ( ~x61 & n899 ) | ( x189 & n899 ) ;
  assign n901 = ( ~n898 & n899 ) | ( ~n898 & n900 ) | ( n899 & n900 ) ;
  assign n902 = x61 & x189 ;
  assign n903 = x61 | x189 ;
  assign n904 = n902 | n903 ;
  assign n905 = ( n898 & n902 ) | ( n898 & n904 ) | ( n902 & n904 ) ;
  assign n906 = ( x62 & ~x190 ) | ( x62 & n905 ) | ( ~x190 & n905 ) ;
  assign n907 = ( ~x62 & x190 ) | ( ~x62 & n906 ) | ( x190 & n906 ) ;
  assign n908 = ( ~n905 & n906 ) | ( ~n905 & n907 ) | ( n906 & n907 ) ;
  assign n909 = x62 & x190 ;
  assign n910 = x62 | x190 ;
  assign n911 = n902 & n910 ;
  assign n912 = n909 | n911 ;
  assign n913 = n909 | n910 ;
  assign n914 = ( n904 & n909 ) | ( n904 & n913 ) | ( n909 & n913 ) ;
  assign n915 = ( n898 & n912 ) | ( n898 & n914 ) | ( n912 & n914 ) ;
  assign n916 = ( x63 & ~x191 ) | ( x63 & n915 ) | ( ~x191 & n915 ) ;
  assign n917 = ( ~x63 & x191 ) | ( ~x63 & n916 ) | ( x191 & n916 ) ;
  assign n918 = ( ~n915 & n916 ) | ( ~n915 & n917 ) | ( n916 & n917 ) ;
  assign n919 = x63 & x191 ;
  assign n920 = x63 | x191 ;
  assign n921 = n909 & n920 ;
  assign n922 = ( n911 & n920 ) | ( n911 & n921 ) | ( n920 & n921 ) ;
  assign n923 = n919 | n922 ;
  assign n924 = n919 | n920 ;
  assign n925 = ( n914 & n919 ) | ( n914 & n924 ) | ( n919 & n924 ) ;
  assign n926 = ( n898 & n923 ) | ( n898 & n925 ) | ( n923 & n925 ) ;
  assign n927 = ( x64 & ~x192 ) | ( x64 & n926 ) | ( ~x192 & n926 ) ;
  assign n928 = ( ~x64 & x192 ) | ( ~x64 & n927 ) | ( x192 & n927 ) ;
  assign n929 = ( ~n926 & n927 ) | ( ~n926 & n928 ) | ( n927 & n928 ) ;
  assign n930 = x64 & x192 ;
  assign n931 = x64 | x192 ;
  assign n932 = n919 & n931 ;
  assign n933 = n924 & n931 ;
  assign n934 = ( n914 & n932 ) | ( n914 & n933 ) | ( n932 & n933 ) ;
  assign n935 = n930 | n934 ;
  assign n936 = n930 | n932 ;
  assign n937 = n930 | n931 ;
  assign n938 = ( n922 & n936 ) | ( n922 & n937 ) | ( n936 & n937 ) ;
  assign n939 = ( n898 & n935 ) | ( n898 & n938 ) | ( n935 & n938 ) ;
  assign n940 = ( x65 & ~x193 ) | ( x65 & n939 ) | ( ~x193 & n939 ) ;
  assign n941 = ( ~x65 & x193 ) | ( ~x65 & n940 ) | ( x193 & n940 ) ;
  assign n942 = ( ~n939 & n940 ) | ( ~n939 & n941 ) | ( n940 & n941 ) ;
  assign n943 = x65 & x193 ;
  assign n944 = x65 | x193 ;
  assign n945 = n930 & n944 ;
  assign n946 = n943 | n945 ;
  assign n947 = n943 | n944 ;
  assign n948 = ( n934 & n946 ) | ( n934 & n947 ) | ( n946 & n947 ) ;
  assign n949 = ( n938 & n943 ) | ( n938 & n947 ) | ( n943 & n947 ) ;
  assign n950 = ( n898 & n948 ) | ( n898 & n949 ) | ( n948 & n949 ) ;
  assign n951 = ( x66 & ~x194 ) | ( x66 & n950 ) | ( ~x194 & n950 ) ;
  assign n952 = ( ~x66 & x194 ) | ( ~x66 & n951 ) | ( x194 & n951 ) ;
  assign n953 = ( ~n950 & n951 ) | ( ~n950 & n952 ) | ( n951 & n952 ) ;
  assign n954 = x66 & x194 ;
  assign n955 = x66 | x194 ;
  assign n956 = n947 & n955 ;
  assign n957 = n946 & n955 ;
  assign n958 = ( n934 & n956 ) | ( n934 & n957 ) | ( n956 & n957 ) ;
  assign n959 = n954 | n958 ;
  assign n960 = n954 | n956 ;
  assign n961 = n943 & n955 ;
  assign n962 = n954 | n961 ;
  assign n963 = ( n938 & n960 ) | ( n938 & n962 ) | ( n960 & n962 ) ;
  assign n964 = ( n898 & n959 ) | ( n898 & n963 ) | ( n959 & n963 ) ;
  assign n965 = ( x67 & ~x195 ) | ( x67 & n964 ) | ( ~x195 & n964 ) ;
  assign n966 = ( ~x67 & x195 ) | ( ~x67 & n965 ) | ( x195 & n965 ) ;
  assign n967 = ( ~n964 & n965 ) | ( ~n964 & n966 ) | ( n965 & n966 ) ;
  assign n968 = x67 & x195 ;
  assign n969 = x67 | x195 ;
  assign n970 = n954 & n969 ;
  assign n971 = n968 | n970 ;
  assign n972 = n968 | n969 ;
  assign n973 = ( n958 & n971 ) | ( n958 & n972 ) | ( n971 & n972 ) ;
  assign n974 = ( n963 & n968 ) | ( n963 & n972 ) | ( n968 & n972 ) ;
  assign n975 = ( n898 & n973 ) | ( n898 & n974 ) | ( n973 & n974 ) ;
  assign n976 = ( x68 & ~x196 ) | ( x68 & n975 ) | ( ~x196 & n975 ) ;
  assign n977 = ( ~x68 & x196 ) | ( ~x68 & n976 ) | ( x196 & n976 ) ;
  assign n978 = ( ~n975 & n976 ) | ( ~n975 & n977 ) | ( n976 & n977 ) ;
  assign n979 = x68 & x196 ;
  assign n980 = x68 | x196 ;
  assign n981 = n968 & n980 ;
  assign n982 = ( n970 & n980 ) | ( n970 & n981 ) | ( n980 & n981 ) ;
  assign n983 = n979 | n982 ;
  assign n984 = n979 | n980 ;
  assign n985 = ( n972 & n979 ) | ( n972 & n984 ) | ( n979 & n984 ) ;
  assign n986 = ( n958 & n983 ) | ( n958 & n985 ) | ( n983 & n985 ) ;
  assign n987 = n979 | n981 ;
  assign n988 = ( n963 & n985 ) | ( n963 & n987 ) | ( n985 & n987 ) ;
  assign n989 = ( n893 & n986 ) | ( n893 & n988 ) | ( n986 & n988 ) ;
  assign n990 = ( n897 & n986 ) | ( n897 & n988 ) | ( n986 & n988 ) ;
  assign n991 = ( n820 & n989 ) | ( n820 & n990 ) | ( n989 & n990 ) ;
  assign n992 = ( x69 & ~x197 ) | ( x69 & n991 ) | ( ~x197 & n991 ) ;
  assign n993 = ( ~x69 & x197 ) | ( ~x69 & n992 ) | ( x197 & n992 ) ;
  assign n994 = ( ~n991 & n992 ) | ( ~n991 & n993 ) | ( n992 & n993 ) ;
  assign n995 = x69 & x197 ;
  assign n996 = x69 | x197 ;
  assign n997 = n995 | n996 ;
  assign n998 = ( n991 & n995 ) | ( n991 & n997 ) | ( n995 & n997 ) ;
  assign n999 = ( x70 & ~x198 ) | ( x70 & n998 ) | ( ~x198 & n998 ) ;
  assign n1000 = ( ~x70 & x198 ) | ( ~x70 & n999 ) | ( x198 & n999 ) ;
  assign n1001 = ( ~n998 & n999 ) | ( ~n998 & n1000 ) | ( n999 & n1000 ) ;
  assign n1002 = x70 & x198 ;
  assign n1003 = x70 | x198 ;
  assign n1004 = n995 & n1003 ;
  assign n1005 = n1002 | n1004 ;
  assign n1006 = n1002 | n1003 ;
  assign n1007 = ( n997 & n1002 ) | ( n997 & n1006 ) | ( n1002 & n1006 ) ;
  assign n1008 = ( n991 & n1005 ) | ( n991 & n1007 ) | ( n1005 & n1007 ) ;
  assign n1009 = ( x71 & ~x199 ) | ( x71 & n1008 ) | ( ~x199 & n1008 ) ;
  assign n1010 = ( ~x71 & x199 ) | ( ~x71 & n1009 ) | ( x199 & n1009 ) ;
  assign n1011 = ( ~n1008 & n1009 ) | ( ~n1008 & n1010 ) | ( n1009 & n1010 ) ;
  assign n1012 = x71 & x199 ;
  assign n1013 = x71 | x199 ;
  assign n1014 = n1002 & n1013 ;
  assign n1015 = ( n1004 & n1013 ) | ( n1004 & n1014 ) | ( n1013 & n1014 ) ;
  assign n1016 = n1012 | n1015 ;
  assign n1017 = n1012 | n1013 ;
  assign n1018 = ( n1007 & n1012 ) | ( n1007 & n1017 ) | ( n1012 & n1017 ) ;
  assign n1019 = ( n991 & n1016 ) | ( n991 & n1018 ) | ( n1016 & n1018 ) ;
  assign n1020 = ( x72 & ~x200 ) | ( x72 & n1019 ) | ( ~x200 & n1019 ) ;
  assign n1021 = ( ~x72 & x200 ) | ( ~x72 & n1020 ) | ( x200 & n1020 ) ;
  assign n1022 = ( ~n1019 & n1020 ) | ( ~n1019 & n1021 ) | ( n1020 & n1021 ) ;
  assign n1023 = x72 & x200 ;
  assign n1024 = x72 | x200 ;
  assign n1025 = n1012 & n1024 ;
  assign n1026 = n1017 & n1024 ;
  assign n1027 = ( n1007 & n1025 ) | ( n1007 & n1026 ) | ( n1025 & n1026 ) ;
  assign n1028 = n1023 | n1027 ;
  assign n1029 = n1023 | n1025 ;
  assign n1030 = n1023 | n1024 ;
  assign n1031 = ( n1015 & n1029 ) | ( n1015 & n1030 ) | ( n1029 & n1030 ) ;
  assign n1032 = ( n991 & n1028 ) | ( n991 & n1031 ) | ( n1028 & n1031 ) ;
  assign n1033 = ( x73 & ~x201 ) | ( x73 & n1032 ) | ( ~x201 & n1032 ) ;
  assign n1034 = ( ~x73 & x201 ) | ( ~x73 & n1033 ) | ( x201 & n1033 ) ;
  assign n1035 = ( ~n1032 & n1033 ) | ( ~n1032 & n1034 ) | ( n1033 & n1034 ) ;
  assign n1036 = x73 & x201 ;
  assign n1037 = x73 | x201 ;
  assign n1038 = n1023 & n1037 ;
  assign n1039 = n1036 | n1038 ;
  assign n1040 = n1036 | n1037 ;
  assign n1041 = ( n1027 & n1039 ) | ( n1027 & n1040 ) | ( n1039 & n1040 ) ;
  assign n1042 = ( n1031 & n1036 ) | ( n1031 & n1040 ) | ( n1036 & n1040 ) ;
  assign n1043 = ( n991 & n1041 ) | ( n991 & n1042 ) | ( n1041 & n1042 ) ;
  assign n1044 = ( x74 & ~x202 ) | ( x74 & n1043 ) | ( ~x202 & n1043 ) ;
  assign n1045 = ( ~x74 & x202 ) | ( ~x74 & n1044 ) | ( x202 & n1044 ) ;
  assign n1046 = ( ~n1043 & n1044 ) | ( ~n1043 & n1045 ) | ( n1044 & n1045 ) ;
  assign n1047 = x74 & x202 ;
  assign n1048 = x74 | x202 ;
  assign n1049 = n1040 & n1048 ;
  assign n1050 = n1039 & n1048 ;
  assign n1051 = ( n1027 & n1049 ) | ( n1027 & n1050 ) | ( n1049 & n1050 ) ;
  assign n1052 = n1047 | n1051 ;
  assign n1053 = n1047 | n1049 ;
  assign n1054 = n1036 & n1048 ;
  assign n1055 = n1047 | n1054 ;
  assign n1056 = ( n1031 & n1053 ) | ( n1031 & n1055 ) | ( n1053 & n1055 ) ;
  assign n1057 = ( n991 & n1052 ) | ( n991 & n1056 ) | ( n1052 & n1056 ) ;
  assign n1058 = ( x75 & ~x203 ) | ( x75 & n1057 ) | ( ~x203 & n1057 ) ;
  assign n1059 = ( ~x75 & x203 ) | ( ~x75 & n1058 ) | ( x203 & n1058 ) ;
  assign n1060 = ( ~n1057 & n1058 ) | ( ~n1057 & n1059 ) | ( n1058 & n1059 ) ;
  assign n1061 = x75 & x203 ;
  assign n1062 = x75 | x203 ;
  assign n1063 = n1047 & n1062 ;
  assign n1064 = n1061 | n1063 ;
  assign n1065 = n1061 | n1062 ;
  assign n1066 = ( n1051 & n1064 ) | ( n1051 & n1065 ) | ( n1064 & n1065 ) ;
  assign n1067 = ( n1056 & n1061 ) | ( n1056 & n1065 ) | ( n1061 & n1065 ) ;
  assign n1068 = ( n991 & n1066 ) | ( n991 & n1067 ) | ( n1066 & n1067 ) ;
  assign n1069 = ( x76 & ~x204 ) | ( x76 & n1068 ) | ( ~x204 & n1068 ) ;
  assign n1070 = ( ~x76 & x204 ) | ( ~x76 & n1069 ) | ( x204 & n1069 ) ;
  assign n1071 = ( ~n1068 & n1069 ) | ( ~n1068 & n1070 ) | ( n1069 & n1070 ) ;
  assign n1072 = x76 & x204 ;
  assign n1073 = x76 | x204 ;
  assign n1074 = n1061 & n1073 ;
  assign n1075 = ( n1063 & n1073 ) | ( n1063 & n1074 ) | ( n1073 & n1074 ) ;
  assign n1076 = n1072 | n1075 ;
  assign n1077 = n1072 | n1073 ;
  assign n1078 = ( n1065 & n1072 ) | ( n1065 & n1077 ) | ( n1072 & n1077 ) ;
  assign n1079 = ( n1051 & n1076 ) | ( n1051 & n1078 ) | ( n1076 & n1078 ) ;
  assign n1080 = n1072 | n1074 ;
  assign n1081 = ( n1056 & n1078 ) | ( n1056 & n1080 ) | ( n1078 & n1080 ) ;
  assign n1082 = ( n991 & n1079 ) | ( n991 & n1081 ) | ( n1079 & n1081 ) ;
  assign n1083 = ( x77 & ~x205 ) | ( x77 & n1082 ) | ( ~x205 & n1082 ) ;
  assign n1084 = ( ~x77 & x205 ) | ( ~x77 & n1083 ) | ( x205 & n1083 ) ;
  assign n1085 = ( ~n1082 & n1083 ) | ( ~n1082 & n1084 ) | ( n1083 & n1084 ) ;
  assign n1086 = x78 | x206 ;
  assign n1087 = x78 & x206 ;
  assign n1088 = n1086 | n1087 ;
  assign n1089 = x77 & x205 ;
  assign n1090 = x77 | x205 ;
  assign n1091 = n1076 & n1090 ;
  assign n1092 = n1078 & n1090 ;
  assign n1093 = ( n1051 & n1091 ) | ( n1051 & n1092 ) | ( n1091 & n1092 ) ;
  assign n1094 = n1080 & n1090 ;
  assign n1095 = ( n1056 & n1092 ) | ( n1056 & n1094 ) | ( n1092 & n1094 ) ;
  assign n1096 = ( n990 & n1093 ) | ( n990 & n1095 ) | ( n1093 & n1095 ) ;
  assign n1097 = ( n989 & n1093 ) | ( n989 & n1095 ) | ( n1093 & n1095 ) ;
  assign n1098 = ( n820 & n1096 ) | ( n820 & n1097 ) | ( n1096 & n1097 ) ;
  assign n1099 = n1089 | n1098 ;
  assign n1100 = ( n1087 & ~n1088 ) | ( n1087 & n1099 ) | ( ~n1088 & n1099 ) ;
  assign n1101 = ( n1087 & n1088 ) | ( n1087 & n1099 ) | ( n1088 & n1099 ) ;
  assign n1102 = ( n1088 & n1100 ) | ( n1088 & ~n1101 ) | ( n1100 & ~n1101 ) ;
  assign n1103 = ( x78 & x206 ) | ( x78 & n1099 ) | ( x206 & n1099 ) ;
  assign n1104 = ( x79 & ~x207 ) | ( x79 & n1103 ) | ( ~x207 & n1103 ) ;
  assign n1105 = ( ~x79 & x207 ) | ( ~x79 & n1104 ) | ( x207 & n1104 ) ;
  assign n1106 = ( ~n1103 & n1104 ) | ( ~n1103 & n1105 ) | ( n1104 & n1105 ) ;
  assign n1107 = x80 | x208 ;
  assign n1108 = x80 & x208 ;
  assign n1109 = n1107 & ~n1108 ;
  assign n1110 = x79 & x207 ;
  assign n1111 = x79 | x207 ;
  assign n1112 = n1086 & n1089 ;
  assign n1113 = n1087 & n1111 ;
  assign n1114 = ( n1111 & n1112 ) | ( n1111 & n1113 ) | ( n1112 & n1113 ) ;
  assign n1115 = n1110 | n1114 ;
  assign n1116 = n1110 | n1111 ;
  assign n1117 = ( n1088 & n1110 ) | ( n1088 & n1116 ) | ( n1110 & n1116 ) ;
  assign n1118 = ( n1098 & n1115 ) | ( n1098 & n1117 ) | ( n1115 & n1117 ) ;
  assign n1119 = n1109 | n1118 ;
  assign n1120 = n1109 & n1118 ;
  assign n1121 = n1119 & ~n1120 ;
  assign n1122 = n1107 | n1108 ;
  assign n1123 = ( n1108 & n1117 ) | ( n1108 & n1122 ) | ( n1117 & n1122 ) ;
  assign n1124 = ( x80 & x208 ) | ( x80 & n1110 ) | ( x208 & n1110 ) ;
  assign n1125 = ( n1107 & n1114 ) | ( n1107 & n1124 ) | ( n1114 & n1124 ) ;
  assign n1126 = ( n1098 & n1123 ) | ( n1098 & n1125 ) | ( n1123 & n1125 ) ;
  assign n1127 = ( x81 & ~x209 ) | ( x81 & n1126 ) | ( ~x209 & n1126 ) ;
  assign n1128 = ( ~x81 & x209 ) | ( ~x81 & n1127 ) | ( x209 & n1127 ) ;
  assign n1129 = ( ~n1126 & n1127 ) | ( ~n1126 & n1128 ) | ( n1127 & n1128 ) ;
  assign n1130 = x81 & x209 ;
  assign n1131 = x81 | x209 ;
  assign n1132 = n1122 & n1131 ;
  assign n1133 = n1108 & n1131 ;
  assign n1134 = ( n1117 & n1132 ) | ( n1117 & n1133 ) | ( n1132 & n1133 ) ;
  assign n1135 = n1130 | n1134 ;
  assign n1136 = n1130 | n1131 ;
  assign n1137 = ( n1125 & n1130 ) | ( n1125 & n1136 ) | ( n1130 & n1136 ) ;
  assign n1138 = ( n1098 & n1135 ) | ( n1098 & n1137 ) | ( n1135 & n1137 ) ;
  assign n1139 = ( x82 & ~x210 ) | ( x82 & n1138 ) | ( ~x210 & n1138 ) ;
  assign n1140 = ( ~x82 & x210 ) | ( ~x82 & n1139 ) | ( x210 & n1139 ) ;
  assign n1141 = ( ~n1138 & n1139 ) | ( ~n1138 & n1140 ) | ( n1139 & n1140 ) ;
  assign n1142 = x82 & x210 ;
  assign n1143 = x82 | x210 ;
  assign n1144 = n1130 & n1143 ;
  assign n1145 = n1142 | n1144 ;
  assign n1146 = n1142 | n1143 ;
  assign n1147 = ( n1136 & n1142 ) | ( n1136 & n1146 ) | ( n1142 & n1146 ) ;
  assign n1148 = ( n1125 & n1145 ) | ( n1125 & n1147 ) | ( n1145 & n1147 ) ;
  assign n1149 = ( n1134 & n1145 ) | ( n1134 & n1146 ) | ( n1145 & n1146 ) ;
  assign n1150 = ( n1098 & n1148 ) | ( n1098 & n1149 ) | ( n1148 & n1149 ) ;
  assign n1151 = ( x83 & ~x211 ) | ( x83 & n1150 ) | ( ~x211 & n1150 ) ;
  assign n1152 = ( ~x83 & x211 ) | ( ~x83 & n1151 ) | ( x211 & n1151 ) ;
  assign n1153 = ( ~n1150 & n1151 ) | ( ~n1150 & n1152 ) | ( n1151 & n1152 ) ;
  assign n1154 = x83 & x211 ;
  assign n1155 = x83 | x211 ;
  assign n1156 = n1145 & n1155 ;
  assign n1157 = n1146 & n1155 ;
  assign n1158 = ( n1134 & n1156 ) | ( n1134 & n1157 ) | ( n1156 & n1157 ) ;
  assign n1159 = n1154 | n1158 ;
  assign n1160 = n1154 | n1155 ;
  assign n1161 = ( n1148 & n1154 ) | ( n1148 & n1160 ) | ( n1154 & n1160 ) ;
  assign n1162 = ( n1098 & n1159 ) | ( n1098 & n1161 ) | ( n1159 & n1161 ) ;
  assign n1163 = ( x84 & ~x212 ) | ( x84 & n1162 ) | ( ~x212 & n1162 ) ;
  assign n1164 = ( ~x84 & x212 ) | ( ~x84 & n1163 ) | ( x212 & n1163 ) ;
  assign n1165 = ( ~n1162 & n1163 ) | ( ~n1162 & n1164 ) | ( n1163 & n1164 ) ;
  assign n1166 = x84 & x212 ;
  assign n1167 = x84 | x212 ;
  assign n1168 = n1154 & n1167 ;
  assign n1169 = n1166 | n1168 ;
  assign n1170 = n1166 | n1167 ;
  assign n1171 = ( n1158 & n1169 ) | ( n1158 & n1170 ) | ( n1169 & n1170 ) ;
  assign n1172 = ( n1160 & n1166 ) | ( n1160 & n1170 ) | ( n1166 & n1170 ) ;
  assign n1173 = ( n1147 & n1169 ) | ( n1147 & n1172 ) | ( n1169 & n1172 ) ;
  assign n1174 = ( n1145 & n1169 ) | ( n1145 & n1172 ) | ( n1169 & n1172 ) ;
  assign n1175 = ( n1125 & n1173 ) | ( n1125 & n1174 ) | ( n1173 & n1174 ) ;
  assign n1176 = ( n1098 & n1171 ) | ( n1098 & n1175 ) | ( n1171 & n1175 ) ;
  assign n1177 = ( x85 & ~x213 ) | ( x85 & n1176 ) | ( ~x213 & n1176 ) ;
  assign n1178 = ( ~x85 & x213 ) | ( ~x85 & n1177 ) | ( x213 & n1177 ) ;
  assign n1179 = ( ~n1176 & n1177 ) | ( ~n1176 & n1178 ) | ( n1177 & n1178 ) ;
  assign n1180 = x85 & x213 ;
  assign n1181 = x85 | x213 ;
  assign n1182 = n1166 & n1181 ;
  assign n1183 = ( n1168 & n1181 ) | ( n1168 & n1182 ) | ( n1181 & n1182 ) ;
  assign n1184 = n1180 | n1183 ;
  assign n1185 = n1170 & n1181 ;
  assign n1186 = n1180 | n1185 ;
  assign n1187 = ( n1158 & n1184 ) | ( n1158 & n1186 ) | ( n1184 & n1186 ) ;
  assign n1188 = n1180 | n1181 ;
  assign n1189 = ( n1175 & n1180 ) | ( n1175 & n1188 ) | ( n1180 & n1188 ) ;
  assign n1190 = ( n1098 & n1187 ) | ( n1098 & n1189 ) | ( n1187 & n1189 ) ;
  assign n1191 = ( x86 & ~x214 ) | ( x86 & n1190 ) | ( ~x214 & n1190 ) ;
  assign n1192 = ( ~x86 & x214 ) | ( ~x86 & n1191 ) | ( x214 & n1191 ) ;
  assign n1193 = ( ~n1190 & n1191 ) | ( ~n1190 & n1192 ) | ( n1191 & n1192 ) ;
  assign n1194 = x87 | x215 ;
  assign n1195 = x87 & x215 ;
  assign n1196 = n1194 | n1195 ;
  assign n1197 = x86 & x214 ;
  assign n1198 = x86 | x214 ;
  assign n1199 = n1186 & n1198 ;
  assign n1200 = n1184 & n1198 ;
  assign n1201 = ( n1158 & n1199 ) | ( n1158 & n1200 ) | ( n1199 & n1200 ) ;
  assign n1202 = n1188 & n1198 ;
  assign n1203 = n1180 & n1198 ;
  assign n1204 = ( n1175 & n1202 ) | ( n1175 & n1203 ) | ( n1202 & n1203 ) ;
  assign n1205 = ( n1095 & n1201 ) | ( n1095 & n1204 ) | ( n1201 & n1204 ) ;
  assign n1206 = ( n1093 & n1201 ) | ( n1093 & n1204 ) | ( n1201 & n1204 ) ;
  assign n1207 = ( n989 & n1205 ) | ( n989 & n1206 ) | ( n1205 & n1206 ) ;
  assign n1208 = ( n990 & n1205 ) | ( n990 & n1206 ) | ( n1205 & n1206 ) ;
  assign n1209 = ( n820 & n1207 ) | ( n820 & n1208 ) | ( n1207 & n1208 ) ;
  assign n1210 = n1197 | n1209 ;
  assign n1211 = ( n1195 & ~n1196 ) | ( n1195 & n1210 ) | ( ~n1196 & n1210 ) ;
  assign n1212 = ( n1195 & n1196 ) | ( n1195 & n1210 ) | ( n1196 & n1210 ) ;
  assign n1213 = ( n1196 & n1211 ) | ( n1196 & ~n1212 ) | ( n1211 & ~n1212 ) ;
  assign n1214 = ( x87 & x215 ) | ( x87 & n1210 ) | ( x215 & n1210 ) ;
  assign n1215 = ( x88 & ~x216 ) | ( x88 & n1214 ) | ( ~x216 & n1214 ) ;
  assign n1216 = ( ~x88 & x216 ) | ( ~x88 & n1215 ) | ( x216 & n1215 ) ;
  assign n1217 = ( ~n1214 & n1215 ) | ( ~n1214 & n1216 ) | ( n1215 & n1216 ) ;
  assign n1218 = x89 | x217 ;
  assign n1219 = x89 & x217 ;
  assign n1220 = n1218 & ~n1219 ;
  assign n1221 = x88 & x216 ;
  assign n1222 = x88 | x216 ;
  assign n1223 = n1194 & n1197 ;
  assign n1224 = n1195 & n1222 ;
  assign n1225 = ( n1222 & n1223 ) | ( n1222 & n1224 ) | ( n1223 & n1224 ) ;
  assign n1226 = n1221 | n1225 ;
  assign n1227 = n1221 | n1222 ;
  assign n1228 = ( n1196 & n1221 ) | ( n1196 & n1227 ) | ( n1221 & n1227 ) ;
  assign n1229 = ( n1209 & n1226 ) | ( n1209 & n1228 ) | ( n1226 & n1228 ) ;
  assign n1230 = n1220 | n1229 ;
  assign n1231 = n1220 & n1229 ;
  assign n1232 = n1230 & ~n1231 ;
  assign n1233 = n1218 | n1219 ;
  assign n1234 = ( n1219 & n1228 ) | ( n1219 & n1233 ) | ( n1228 & n1233 ) ;
  assign n1235 = ( x89 & x217 ) | ( x89 & n1221 ) | ( x217 & n1221 ) ;
  assign n1236 = ( n1218 & n1225 ) | ( n1218 & n1235 ) | ( n1225 & n1235 ) ;
  assign n1237 = ( n1209 & n1234 ) | ( n1209 & n1236 ) | ( n1234 & n1236 ) ;
  assign n1238 = ( x90 & ~x218 ) | ( x90 & n1237 ) | ( ~x218 & n1237 ) ;
  assign n1239 = ( ~x90 & x218 ) | ( ~x90 & n1238 ) | ( x218 & n1238 ) ;
  assign n1240 = ( ~n1237 & n1238 ) | ( ~n1237 & n1239 ) | ( n1238 & n1239 ) ;
  assign n1241 = x90 & x218 ;
  assign n1242 = x90 | x218 ;
  assign n1243 = n1233 & n1242 ;
  assign n1244 = n1219 & n1242 ;
  assign n1245 = ( n1228 & n1243 ) | ( n1228 & n1244 ) | ( n1243 & n1244 ) ;
  assign n1246 = n1241 | n1245 ;
  assign n1247 = n1241 | n1242 ;
  assign n1248 = ( n1236 & n1241 ) | ( n1236 & n1247 ) | ( n1241 & n1247 ) ;
  assign n1249 = ( n1209 & n1246 ) | ( n1209 & n1248 ) | ( n1246 & n1248 ) ;
  assign n1250 = ( x91 & ~x219 ) | ( x91 & n1249 ) | ( ~x219 & n1249 ) ;
  assign n1251 = ( ~x91 & x219 ) | ( ~x91 & n1250 ) | ( x219 & n1250 ) ;
  assign n1252 = ( ~n1249 & n1250 ) | ( ~n1249 & n1251 ) | ( n1250 & n1251 ) ;
  assign n1253 = x91 & x219 ;
  assign n1254 = x91 | x219 ;
  assign n1255 = n1241 & n1254 ;
  assign n1256 = n1253 | n1255 ;
  assign n1257 = n1253 | n1254 ;
  assign n1258 = ( n1247 & n1253 ) | ( n1247 & n1257 ) | ( n1253 & n1257 ) ;
  assign n1259 = ( n1236 & n1256 ) | ( n1236 & n1258 ) | ( n1256 & n1258 ) ;
  assign n1260 = ( n1245 & n1256 ) | ( n1245 & n1257 ) | ( n1256 & n1257 ) ;
  assign n1261 = ( n1209 & n1259 ) | ( n1209 & n1260 ) | ( n1259 & n1260 ) ;
  assign n1262 = ( x92 & ~x220 ) | ( x92 & n1261 ) | ( ~x220 & n1261 ) ;
  assign n1263 = ( ~x92 & x220 ) | ( ~x92 & n1262 ) | ( x220 & n1262 ) ;
  assign n1264 = ( ~n1261 & n1262 ) | ( ~n1261 & n1263 ) | ( n1262 & n1263 ) ;
  assign n1265 = x92 & x220 ;
  assign n1266 = x92 | x220 ;
  assign n1267 = n1256 & n1266 ;
  assign n1268 = n1257 & n1266 ;
  assign n1269 = ( n1245 & n1267 ) | ( n1245 & n1268 ) | ( n1267 & n1268 ) ;
  assign n1270 = n1265 | n1269 ;
  assign n1271 = n1265 | n1266 ;
  assign n1272 = ( n1259 & n1265 ) | ( n1259 & n1271 ) | ( n1265 & n1271 ) ;
  assign n1273 = ( n1209 & n1270 ) | ( n1209 & n1272 ) | ( n1270 & n1272 ) ;
  assign n1274 = ( x93 & ~x221 ) | ( x93 & n1273 ) | ( ~x221 & n1273 ) ;
  assign n1275 = ( ~x93 & x221 ) | ( ~x93 & n1274 ) | ( x221 & n1274 ) ;
  assign n1276 = ( ~n1273 & n1274 ) | ( ~n1273 & n1275 ) | ( n1274 & n1275 ) ;
  assign n1277 = x93 & x221 ;
  assign n1278 = x93 | x221 ;
  assign n1279 = n1265 & n1278 ;
  assign n1280 = n1277 | n1279 ;
  assign n1281 = n1277 | n1278 ;
  assign n1282 = ( n1269 & n1280 ) | ( n1269 & n1281 ) | ( n1280 & n1281 ) ;
  assign n1283 = ( n1271 & n1277 ) | ( n1271 & n1281 ) | ( n1277 & n1281 ) ;
  assign n1284 = ( n1258 & n1280 ) | ( n1258 & n1283 ) | ( n1280 & n1283 ) ;
  assign n1285 = ( n1256 & n1280 ) | ( n1256 & n1283 ) | ( n1280 & n1283 ) ;
  assign n1286 = ( n1236 & n1284 ) | ( n1236 & n1285 ) | ( n1284 & n1285 ) ;
  assign n1287 = ( n1209 & n1282 ) | ( n1209 & n1286 ) | ( n1282 & n1286 ) ;
  assign n1288 = ( x94 & ~x222 ) | ( x94 & n1287 ) | ( ~x222 & n1287 ) ;
  assign n1289 = ( ~x94 & x222 ) | ( ~x94 & n1288 ) | ( x222 & n1288 ) ;
  assign n1290 = ( ~n1287 & n1288 ) | ( ~n1287 & n1289 ) | ( n1288 & n1289 ) ;
  assign n1291 = x95 | x223 ;
  assign n1292 = x95 & x223 ;
  assign n1293 = n1291 & ~n1292 ;
  assign n1294 = x94 & x222 ;
  assign n1295 = x94 | x222 ;
  assign n1296 = n1294 | n1295 ;
  assign n1297 = ( n1286 & n1294 ) | ( n1286 & n1296 ) | ( n1294 & n1296 ) ;
  assign n1298 = n1277 & n1295 ;
  assign n1299 = ( n1279 & n1295 ) | ( n1279 & n1298 ) | ( n1295 & n1298 ) ;
  assign n1300 = n1294 | n1299 ;
  assign n1301 = n1281 & n1295 ;
  assign n1302 = n1294 | n1301 ;
  assign n1303 = ( n1269 & n1300 ) | ( n1269 & n1302 ) | ( n1300 & n1302 ) ;
  assign n1304 = ( n1209 & n1297 ) | ( n1209 & n1303 ) | ( n1297 & n1303 ) ;
  assign n1305 = n1293 | n1304 ;
  assign n1306 = n1293 & n1304 ;
  assign n1307 = n1305 & ~n1306 ;
  assign n1308 = ( x95 & x223 ) | ( x95 & n1296 ) | ( x223 & n1296 ) ;
  assign n1309 = ( x95 & x223 ) | ( x95 & n1294 ) | ( x223 & n1294 ) ;
  assign n1310 = ( n1286 & n1308 ) | ( n1286 & n1309 ) | ( n1308 & n1309 ) ;
  assign n1311 = n1291 | n1292 ;
  assign n1312 = ( n1292 & n1302 ) | ( n1292 & n1311 ) | ( n1302 & n1311 ) ;
  assign n1313 = ( n1292 & n1300 ) | ( n1292 & n1311 ) | ( n1300 & n1311 ) ;
  assign n1314 = ( n1269 & n1312 ) | ( n1269 & n1313 ) | ( n1312 & n1313 ) ;
  assign n1315 = ( n1209 & n1310 ) | ( n1209 & n1314 ) | ( n1310 & n1314 ) ;
  assign n1316 = ( x96 & ~x224 ) | ( x96 & n1315 ) | ( ~x224 & n1315 ) ;
  assign n1317 = ( ~x96 & x224 ) | ( ~x96 & n1316 ) | ( x224 & n1316 ) ;
  assign n1318 = ( ~n1315 & n1316 ) | ( ~n1315 & n1317 ) | ( n1316 & n1317 ) ;
  assign n1319 = x96 & x224 ;
  assign n1320 = x96 | x224 ;
  assign n1321 = n1319 | n1320 ;
  assign n1322 = ( n1315 & n1319 ) | ( n1315 & n1321 ) | ( n1319 & n1321 ) ;
  assign n1323 = ( x97 & ~x225 ) | ( x97 & n1322 ) | ( ~x225 & n1322 ) ;
  assign n1324 = ( ~x97 & x225 ) | ( ~x97 & n1323 ) | ( x225 & n1323 ) ;
  assign n1325 = ( ~n1322 & n1323 ) | ( ~n1322 & n1324 ) | ( n1323 & n1324 ) ;
  assign n1326 = x97 & x225 ;
  assign n1327 = x97 | x225 ;
  assign n1328 = n1319 & n1327 ;
  assign n1329 = n1326 | n1328 ;
  assign n1330 = n1326 | n1327 ;
  assign n1331 = ( n1321 & n1326 ) | ( n1321 & n1330 ) | ( n1326 & n1330 ) ;
  assign n1332 = ( n1315 & n1329 ) | ( n1315 & n1331 ) | ( n1329 & n1331 ) ;
  assign n1333 = ( x98 & ~x226 ) | ( x98 & n1332 ) | ( ~x226 & n1332 ) ;
  assign n1334 = ( ~x98 & x226 ) | ( ~x98 & n1333 ) | ( x226 & n1333 ) ;
  assign n1335 = ( ~n1332 & n1333 ) | ( ~n1332 & n1334 ) | ( n1333 & n1334 ) ;
  assign n1336 = x98 & x226 ;
  assign n1337 = x98 | x226 ;
  assign n1338 = n1326 & n1337 ;
  assign n1339 = ( n1328 & n1337 ) | ( n1328 & n1338 ) | ( n1337 & n1338 ) ;
  assign n1340 = n1336 | n1339 ;
  assign n1341 = n1336 | n1337 ;
  assign n1342 = ( n1331 & n1336 ) | ( n1331 & n1341 ) | ( n1336 & n1341 ) ;
  assign n1343 = ( n1315 & n1340 ) | ( n1315 & n1342 ) | ( n1340 & n1342 ) ;
  assign n1344 = ( x99 & ~x227 ) | ( x99 & n1343 ) | ( ~x227 & n1343 ) ;
  assign n1345 = ( ~x99 & x227 ) | ( ~x99 & n1344 ) | ( x227 & n1344 ) ;
  assign n1346 = ( ~n1343 & n1344 ) | ( ~n1343 & n1345 ) | ( n1344 & n1345 ) ;
  assign n1347 = x99 & x227 ;
  assign n1348 = x99 | x227 ;
  assign n1349 = n1336 & n1348 ;
  assign n1350 = n1341 & n1348 ;
  assign n1351 = ( n1331 & n1349 ) | ( n1331 & n1350 ) | ( n1349 & n1350 ) ;
  assign n1352 = n1347 | n1351 ;
  assign n1353 = n1347 | n1349 ;
  assign n1354 = n1347 | n1348 ;
  assign n1355 = ( n1339 & n1353 ) | ( n1339 & n1354 ) | ( n1353 & n1354 ) ;
  assign n1356 = ( n1315 & n1352 ) | ( n1315 & n1355 ) | ( n1352 & n1355 ) ;
  assign n1357 = ( x100 & ~x228 ) | ( x100 & n1356 ) | ( ~x228 & n1356 ) ;
  assign n1358 = ( ~x100 & x228 ) | ( ~x100 & n1357 ) | ( x228 & n1357 ) ;
  assign n1359 = ( ~n1356 & n1357 ) | ( ~n1356 & n1358 ) | ( n1357 & n1358 ) ;
  assign n1360 = x100 & x228 ;
  assign n1361 = x100 | x228 ;
  assign n1362 = n1347 & n1361 ;
  assign n1363 = n1360 | n1362 ;
  assign n1364 = n1360 | n1361 ;
  assign n1365 = ( n1351 & n1363 ) | ( n1351 & n1364 ) | ( n1363 & n1364 ) ;
  assign n1366 = ( n1355 & n1360 ) | ( n1355 & n1364 ) | ( n1360 & n1364 ) ;
  assign n1367 = ( n1315 & n1365 ) | ( n1315 & n1366 ) | ( n1365 & n1366 ) ;
  assign n1368 = ( x101 & ~x229 ) | ( x101 & n1367 ) | ( ~x229 & n1367 ) ;
  assign n1369 = ( ~x101 & x229 ) | ( ~x101 & n1368 ) | ( x229 & n1368 ) ;
  assign n1370 = ( ~n1367 & n1368 ) | ( ~n1367 & n1369 ) | ( n1368 & n1369 ) ;
  assign n1371 = x101 & x229 ;
  assign n1372 = x101 | x229 ;
  assign n1373 = n1364 & n1372 ;
  assign n1374 = n1363 & n1372 ;
  assign n1375 = ( n1351 & n1373 ) | ( n1351 & n1374 ) | ( n1373 & n1374 ) ;
  assign n1376 = n1371 | n1375 ;
  assign n1377 = n1371 | n1373 ;
  assign n1378 = n1360 & n1372 ;
  assign n1379 = n1371 | n1378 ;
  assign n1380 = ( n1355 & n1377 ) | ( n1355 & n1379 ) | ( n1377 & n1379 ) ;
  assign n1381 = ( n1315 & n1376 ) | ( n1315 & n1380 ) | ( n1376 & n1380 ) ;
  assign n1382 = ( x102 & ~x230 ) | ( x102 & n1381 ) | ( ~x230 & n1381 ) ;
  assign n1383 = ( ~x102 & x230 ) | ( ~x102 & n1382 ) | ( x230 & n1382 ) ;
  assign n1384 = ( ~n1381 & n1382 ) | ( ~n1381 & n1383 ) | ( n1382 & n1383 ) ;
  assign n1385 = x102 & x230 ;
  assign n1386 = x102 | x230 ;
  assign n1387 = n1371 & n1386 ;
  assign n1388 = n1385 | n1387 ;
  assign n1389 = n1385 | n1386 ;
  assign n1390 = ( n1375 & n1388 ) | ( n1375 & n1389 ) | ( n1388 & n1389 ) ;
  assign n1391 = ( n1380 & n1385 ) | ( n1380 & n1389 ) | ( n1385 & n1389 ) ;
  assign n1392 = ( n1315 & n1390 ) | ( n1315 & n1391 ) | ( n1390 & n1391 ) ;
  assign n1393 = ( x103 & ~x231 ) | ( x103 & n1392 ) | ( ~x231 & n1392 ) ;
  assign n1394 = ( ~x103 & x231 ) | ( ~x103 & n1393 ) | ( x231 & n1393 ) ;
  assign n1395 = ( ~n1392 & n1393 ) | ( ~n1392 & n1394 ) | ( n1393 & n1394 ) ;
  assign n1396 = x103 & x231 ;
  assign n1397 = x103 | x231 ;
  assign n1398 = n1385 & n1397 ;
  assign n1399 = ( n1387 & n1397 ) | ( n1387 & n1398 ) | ( n1397 & n1398 ) ;
  assign n1400 = n1396 | n1399 ;
  assign n1401 = n1396 | n1397 ;
  assign n1402 = ( n1389 & n1396 ) | ( n1389 & n1401 ) | ( n1396 & n1401 ) ;
  assign n1403 = ( n1375 & n1400 ) | ( n1375 & n1402 ) | ( n1400 & n1402 ) ;
  assign n1404 = n1396 | n1398 ;
  assign n1405 = ( n1380 & n1402 ) | ( n1380 & n1404 ) | ( n1402 & n1404 ) ;
  assign n1406 = ( n1315 & n1403 ) | ( n1315 & n1405 ) | ( n1403 & n1405 ) ;
  assign n1407 = ( x104 & ~x232 ) | ( x104 & n1406 ) | ( ~x232 & n1406 ) ;
  assign n1408 = ( ~x104 & x232 ) | ( ~x104 & n1407 ) | ( x232 & n1407 ) ;
  assign n1409 = ( ~n1406 & n1407 ) | ( ~n1406 & n1408 ) | ( n1407 & n1408 ) ;
  assign n1410 = x104 & x232 ;
  assign n1411 = x104 | x232 ;
  assign n1412 = n1402 & n1411 ;
  assign n1413 = n1404 & n1411 ;
  assign n1414 = ( n1380 & n1412 ) | ( n1380 & n1413 ) | ( n1412 & n1413 ) ;
  assign n1415 = n1410 | n1414 ;
  assign n1416 = n1410 | n1411 ;
  assign n1417 = ( n1403 & n1410 ) | ( n1403 & n1416 ) | ( n1410 & n1416 ) ;
  assign n1418 = ( n1315 & n1415 ) | ( n1315 & n1417 ) | ( n1415 & n1417 ) ;
  assign n1419 = ( x105 & ~x233 ) | ( x105 & n1418 ) | ( ~x233 & n1418 ) ;
  assign n1420 = ( ~x105 & x233 ) | ( ~x105 & n1419 ) | ( x233 & n1419 ) ;
  assign n1421 = ( ~n1418 & n1419 ) | ( ~n1418 & n1420 ) | ( n1419 & n1420 ) ;
  assign n1422 = x105 & x233 ;
  assign n1423 = x105 | x233 ;
  assign n1424 = n1410 & n1423 ;
  assign n1425 = n1422 | n1424 ;
  assign n1426 = n1422 | n1423 ;
  assign n1427 = ( n1416 & n1422 ) | ( n1416 & n1426 ) | ( n1422 & n1426 ) ;
  assign n1428 = ( n1400 & n1425 ) | ( n1400 & n1427 ) | ( n1425 & n1427 ) ;
  assign n1429 = ( n1402 & n1425 ) | ( n1402 & n1427 ) | ( n1425 & n1427 ) ;
  assign n1430 = ( n1375 & n1428 ) | ( n1375 & n1429 ) | ( n1428 & n1429 ) ;
  assign n1431 = ( n1413 & n1425 ) | ( n1413 & n1426 ) | ( n1425 & n1426 ) ;
  assign n1432 = ( n1412 & n1425 ) | ( n1412 & n1426 ) | ( n1425 & n1426 ) ;
  assign n1433 = ( n1380 & n1431 ) | ( n1380 & n1432 ) | ( n1431 & n1432 ) ;
  assign n1434 = ( n1314 & n1430 ) | ( n1314 & n1433 ) | ( n1430 & n1433 ) ;
  assign n1435 = ( n1310 & n1430 ) | ( n1310 & n1433 ) | ( n1430 & n1433 ) ;
  assign n1436 = ( n1209 & n1434 ) | ( n1209 & n1435 ) | ( n1434 & n1435 ) ;
  assign n1437 = ( x106 & ~x234 ) | ( x106 & n1436 ) | ( ~x234 & n1436 ) ;
  assign n1438 = ( ~x106 & x234 ) | ( ~x106 & n1437 ) | ( x234 & n1437 ) ;
  assign n1439 = ( ~n1436 & n1437 ) | ( ~n1436 & n1438 ) | ( n1437 & n1438 ) ;
  assign n1440 = x106 & x234 ;
  assign n1441 = x106 | x234 ;
  assign n1442 = n1440 | n1441 ;
  assign n1443 = ( n1436 & n1440 ) | ( n1436 & n1442 ) | ( n1440 & n1442 ) ;
  assign n1444 = ( x107 & ~x235 ) | ( x107 & n1443 ) | ( ~x235 & n1443 ) ;
  assign n1445 = ( ~x107 & x235 ) | ( ~x107 & n1444 ) | ( x235 & n1444 ) ;
  assign n1446 = ( ~n1443 & n1444 ) | ( ~n1443 & n1445 ) | ( n1444 & n1445 ) ;
  assign n1447 = x107 & x235 ;
  assign n1448 = x107 | x235 ;
  assign n1449 = n1440 & n1448 ;
  assign n1450 = n1447 | n1449 ;
  assign n1451 = n1447 | n1448 ;
  assign n1452 = ( n1442 & n1447 ) | ( n1442 & n1451 ) | ( n1447 & n1451 ) ;
  assign n1453 = ( n1436 & n1450 ) | ( n1436 & n1452 ) | ( n1450 & n1452 ) ;
  assign n1454 = ( x108 & ~x236 ) | ( x108 & n1453 ) | ( ~x236 & n1453 ) ;
  assign n1455 = ( ~x108 & x236 ) | ( ~x108 & n1454 ) | ( x236 & n1454 ) ;
  assign n1456 = ( ~n1453 & n1454 ) | ( ~n1453 & n1455 ) | ( n1454 & n1455 ) ;
  assign n1457 = x108 & x236 ;
  assign n1458 = x108 | x236 ;
  assign n1459 = n1447 & n1458 ;
  assign n1460 = ( n1449 & n1458 ) | ( n1449 & n1459 ) | ( n1458 & n1459 ) ;
  assign n1461 = n1457 | n1460 ;
  assign n1462 = n1457 | n1458 ;
  assign n1463 = ( n1452 & n1457 ) | ( n1452 & n1462 ) | ( n1457 & n1462 ) ;
  assign n1464 = ( n1436 & n1461 ) | ( n1436 & n1463 ) | ( n1461 & n1463 ) ;
  assign n1465 = ( x109 & ~x237 ) | ( x109 & n1464 ) | ( ~x237 & n1464 ) ;
  assign n1466 = ( ~x109 & x237 ) | ( ~x109 & n1465 ) | ( x237 & n1465 ) ;
  assign n1467 = ( ~n1464 & n1465 ) | ( ~n1464 & n1466 ) | ( n1465 & n1466 ) ;
  assign n1468 = x109 & x237 ;
  assign n1469 = x109 | x237 ;
  assign n1470 = n1457 & n1469 ;
  assign n1471 = n1462 & n1469 ;
  assign n1472 = ( n1452 & n1470 ) | ( n1452 & n1471 ) | ( n1470 & n1471 ) ;
  assign n1473 = n1468 | n1472 ;
  assign n1474 = n1468 | n1470 ;
  assign n1475 = n1468 | n1469 ;
  assign n1476 = ( n1460 & n1474 ) | ( n1460 & n1475 ) | ( n1474 & n1475 ) ;
  assign n1477 = ( n1436 & n1473 ) | ( n1436 & n1476 ) | ( n1473 & n1476 ) ;
  assign n1478 = ( x110 & ~x238 ) | ( x110 & n1477 ) | ( ~x238 & n1477 ) ;
  assign n1479 = ( ~x110 & x238 ) | ( ~x110 & n1478 ) | ( x238 & n1478 ) ;
  assign n1480 = ( ~n1477 & n1478 ) | ( ~n1477 & n1479 ) | ( n1478 & n1479 ) ;
  assign n1481 = x110 & x238 ;
  assign n1482 = x110 | x238 ;
  assign n1483 = n1468 & n1482 ;
  assign n1484 = n1481 | n1483 ;
  assign n1485 = n1481 | n1482 ;
  assign n1486 = ( n1472 & n1484 ) | ( n1472 & n1485 ) | ( n1484 & n1485 ) ;
  assign n1487 = ( n1476 & n1481 ) | ( n1476 & n1485 ) | ( n1481 & n1485 ) ;
  assign n1488 = ( n1436 & n1486 ) | ( n1436 & n1487 ) | ( n1486 & n1487 ) ;
  assign n1489 = ( x111 & ~x239 ) | ( x111 & n1488 ) | ( ~x239 & n1488 ) ;
  assign n1490 = ( ~x111 & x239 ) | ( ~x111 & n1489 ) | ( x239 & n1489 ) ;
  assign n1491 = ( ~n1488 & n1489 ) | ( ~n1488 & n1490 ) | ( n1489 & n1490 ) ;
  assign n1492 = x111 & x239 ;
  assign n1493 = x111 | x239 ;
  assign n1494 = n1485 & n1493 ;
  assign n1495 = n1484 & n1493 ;
  assign n1496 = ( n1472 & n1494 ) | ( n1472 & n1495 ) | ( n1494 & n1495 ) ;
  assign n1497 = n1492 | n1496 ;
  assign n1498 = n1492 | n1494 ;
  assign n1499 = n1481 & n1493 ;
  assign n1500 = n1492 | n1499 ;
  assign n1501 = ( n1476 & n1498 ) | ( n1476 & n1500 ) | ( n1498 & n1500 ) ;
  assign n1502 = ( n1436 & n1497 ) | ( n1436 & n1501 ) | ( n1497 & n1501 ) ;
  assign n1503 = ( x112 & ~x240 ) | ( x112 & n1502 ) | ( ~x240 & n1502 ) ;
  assign n1504 = ( ~x112 & x240 ) | ( ~x112 & n1503 ) | ( x240 & n1503 ) ;
  assign n1505 = ( ~n1502 & n1503 ) | ( ~n1502 & n1504 ) | ( n1503 & n1504 ) ;
  assign n1506 = x112 & x240 ;
  assign n1507 = x112 | x240 ;
  assign n1508 = n1492 & n1507 ;
  assign n1509 = n1506 | n1508 ;
  assign n1510 = n1506 | n1507 ;
  assign n1511 = ( n1496 & n1509 ) | ( n1496 & n1510 ) | ( n1509 & n1510 ) ;
  assign n1512 = ( n1501 & n1506 ) | ( n1501 & n1510 ) | ( n1506 & n1510 ) ;
  assign n1513 = ( n1436 & n1511 ) | ( n1436 & n1512 ) | ( n1511 & n1512 ) ;
  assign n1514 = ( x113 & ~x241 ) | ( x113 & n1513 ) | ( ~x241 & n1513 ) ;
  assign n1515 = ( ~x113 & x241 ) | ( ~x113 & n1514 ) | ( x241 & n1514 ) ;
  assign n1516 = ( ~n1513 & n1514 ) | ( ~n1513 & n1515 ) | ( n1514 & n1515 ) ;
  assign n1517 = x113 & x241 ;
  assign n1518 = x113 | x241 ;
  assign n1519 = n1506 & n1518 ;
  assign n1520 = ( n1508 & n1518 ) | ( n1508 & n1519 ) | ( n1518 & n1519 ) ;
  assign n1521 = n1517 | n1520 ;
  assign n1522 = n1517 | n1518 ;
  assign n1523 = ( n1510 & n1517 ) | ( n1510 & n1522 ) | ( n1517 & n1522 ) ;
  assign n1524 = ( n1496 & n1521 ) | ( n1496 & n1523 ) | ( n1521 & n1523 ) ;
  assign n1525 = n1517 | n1519 ;
  assign n1526 = ( n1501 & n1523 ) | ( n1501 & n1525 ) | ( n1523 & n1525 ) ;
  assign n1527 = ( n1436 & n1524 ) | ( n1436 & n1526 ) | ( n1524 & n1526 ) ;
  assign n1528 = ( x114 & ~x242 ) | ( x114 & n1527 ) | ( ~x242 & n1527 ) ;
  assign n1529 = ( ~x114 & x242 ) | ( ~x114 & n1528 ) | ( x242 & n1528 ) ;
  assign n1530 = ( ~n1527 & n1528 ) | ( ~n1527 & n1529 ) | ( n1528 & n1529 ) ;
  assign n1531 = x114 & x242 ;
  assign n1532 = x114 | x242 ;
  assign n1533 = n1523 & n1532 ;
  assign n1534 = n1525 & n1532 ;
  assign n1535 = ( n1501 & n1533 ) | ( n1501 & n1534 ) | ( n1533 & n1534 ) ;
  assign n1536 = n1531 | n1535 ;
  assign n1537 = n1531 | n1532 ;
  assign n1538 = ( n1524 & n1531 ) | ( n1524 & n1537 ) | ( n1531 & n1537 ) ;
  assign n1539 = ( n1436 & n1536 ) | ( n1436 & n1538 ) | ( n1536 & n1538 ) ;
  assign n1540 = ( x115 & ~x243 ) | ( x115 & n1539 ) | ( ~x243 & n1539 ) ;
  assign n1541 = ( ~x115 & x243 ) | ( ~x115 & n1540 ) | ( x243 & n1540 ) ;
  assign n1542 = ( ~n1539 & n1540 ) | ( ~n1539 & n1541 ) | ( n1540 & n1541 ) ;
  assign n1543 = x115 & x243 ;
  assign n1544 = x115 | x243 ;
  assign n1545 = n1531 & n1544 ;
  assign n1546 = n1543 | n1545 ;
  assign n1547 = n1543 | n1544 ;
  assign n1548 = ( n1535 & n1546 ) | ( n1535 & n1547 ) | ( n1546 & n1547 ) ;
  assign n1549 = ( n1537 & n1543 ) | ( n1537 & n1547 ) | ( n1543 & n1547 ) ;
  assign n1550 = ( n1521 & n1546 ) | ( n1521 & n1549 ) | ( n1546 & n1549 ) ;
  assign n1551 = ( n1523 & n1546 ) | ( n1523 & n1549 ) | ( n1546 & n1549 ) ;
  assign n1552 = ( n1496 & n1550 ) | ( n1496 & n1551 ) | ( n1550 & n1551 ) ;
  assign n1553 = ( n1436 & n1548 ) | ( n1436 & n1552 ) | ( n1548 & n1552 ) ;
  assign n1554 = ( x116 & ~x244 ) | ( x116 & n1553 ) | ( ~x244 & n1553 ) ;
  assign n1555 = ( ~x116 & x244 ) | ( ~x116 & n1554 ) | ( x244 & n1554 ) ;
  assign n1556 = ( ~n1553 & n1554 ) | ( ~n1553 & n1555 ) | ( n1554 & n1555 ) ;
  assign n1557 = x117 | x245 ;
  assign n1558 = x117 & x245 ;
  assign n1559 = n1557 | n1558 ;
  assign n1560 = x116 & x244 ;
  assign n1561 = x116 | x244 ;
  assign n1562 = n1552 & n1561 ;
  assign n1563 = n1547 & n1561 ;
  assign n1564 = n1543 & n1561 ;
  assign n1565 = ( n1545 & n1561 ) | ( n1545 & n1564 ) | ( n1561 & n1564 ) ;
  assign n1566 = ( n1534 & n1563 ) | ( n1534 & n1565 ) | ( n1563 & n1565 ) ;
  assign n1567 = ( n1533 & n1563 ) | ( n1533 & n1565 ) | ( n1563 & n1565 ) ;
  assign n1568 = ( n1501 & n1566 ) | ( n1501 & n1567 ) | ( n1566 & n1567 ) ;
  assign n1569 = ( n1435 & n1562 ) | ( n1435 & n1568 ) | ( n1562 & n1568 ) ;
  assign n1570 = ( n1434 & n1562 ) | ( n1434 & n1568 ) | ( n1562 & n1568 ) ;
  assign n1571 = ( n1208 & n1569 ) | ( n1208 & n1570 ) | ( n1569 & n1570 ) ;
  assign n1572 = ( n1207 & n1569 ) | ( n1207 & n1570 ) | ( n1569 & n1570 ) ;
  assign n1573 = ( n820 & n1571 ) | ( n820 & n1572 ) | ( n1571 & n1572 ) ;
  assign n1574 = n1560 | n1573 ;
  assign n1575 = ( n1558 & ~n1559 ) | ( n1558 & n1574 ) | ( ~n1559 & n1574 ) ;
  assign n1576 = ( n1558 & n1559 ) | ( n1558 & n1574 ) | ( n1559 & n1574 ) ;
  assign n1577 = ( n1559 & n1575 ) | ( n1559 & ~n1576 ) | ( n1575 & ~n1576 ) ;
  assign n1578 = ( x117 & x245 ) | ( x117 & n1560 ) | ( x245 & n1560 ) ;
  assign n1579 = ( n1557 & n1573 ) | ( n1557 & n1578 ) | ( n1573 & n1578 ) ;
  assign n1580 = ( x118 & ~x246 ) | ( x118 & n1578 ) | ( ~x246 & n1578 ) ;
  assign n1581 = ( x118 & ~x246 ) | ( x118 & n1557 ) | ( ~x246 & n1557 ) ;
  assign n1582 = ( n1573 & n1580 ) | ( n1573 & n1581 ) | ( n1580 & n1581 ) ;
  assign n1583 = ( ~x118 & x246 ) | ( ~x118 & n1580 ) | ( x246 & n1580 ) ;
  assign n1584 = ( ~x118 & x246 ) | ( ~x118 & n1581 ) | ( x246 & n1581 ) ;
  assign n1585 = ( n1573 & n1583 ) | ( n1573 & n1584 ) | ( n1583 & n1584 ) ;
  assign n1586 = ( ~n1579 & n1582 ) | ( ~n1579 & n1585 ) | ( n1582 & n1585 ) ;
  assign n1587 = x119 | x247 ;
  assign n1588 = x119 & x247 ;
  assign n1589 = n1587 & ~n1588 ;
  assign n1590 = x118 & x246 ;
  assign n1591 = x118 | x246 ;
  assign n1592 = n1557 & n1560 ;
  assign n1593 = n1558 | n1592 ;
  assign n1594 = n1591 & n1593 ;
  assign n1595 = n1590 | n1594 ;
  assign n1596 = n1590 | n1591 ;
  assign n1597 = ( n1559 & n1590 ) | ( n1559 & n1596 ) | ( n1590 & n1596 ) ;
  assign n1598 = ( n1573 & n1595 ) | ( n1573 & n1597 ) | ( n1595 & n1597 ) ;
  assign n1599 = n1589 | n1598 ;
  assign n1600 = n1589 & n1598 ;
  assign n1601 = n1599 & ~n1600 ;
  assign n1602 = n1587 | n1588 ;
  assign n1603 = ( n1588 & n1597 ) | ( n1588 & n1602 ) | ( n1597 & n1602 ) ;
  assign n1604 = ( x119 & x247 ) | ( x119 & n1595 ) | ( x247 & n1595 ) ;
  assign n1605 = ( n1573 & n1603 ) | ( n1573 & n1604 ) | ( n1603 & n1604 ) ;
  assign n1606 = ( x120 & ~x248 ) | ( x120 & n1605 ) | ( ~x248 & n1605 ) ;
  assign n1607 = ( ~x120 & x248 ) | ( ~x120 & n1606 ) | ( x248 & n1606 ) ;
  assign n1608 = ( ~n1605 & n1606 ) | ( ~n1605 & n1607 ) | ( n1606 & n1607 ) ;
  assign n1609 = x120 & x248 ;
  assign n1610 = x120 | x248 ;
  assign n1611 = n1603 & n1610 ;
  assign n1612 = n1609 | n1611 ;
  assign n1613 = n1609 | n1610 ;
  assign n1614 = ( n1604 & n1609 ) | ( n1604 & n1613 ) | ( n1609 & n1613 ) ;
  assign n1615 = ( n1573 & n1612 ) | ( n1573 & n1614 ) | ( n1612 & n1614 ) ;
  assign n1616 = ( x121 & ~x249 ) | ( x121 & n1615 ) | ( ~x249 & n1615 ) ;
  assign n1617 = ( ~x121 & x249 ) | ( ~x121 & n1616 ) | ( x249 & n1616 ) ;
  assign n1618 = ( ~n1615 & n1616 ) | ( ~n1615 & n1617 ) | ( n1616 & n1617 ) ;
  assign n1619 = x121 & x249 ;
  assign n1620 = x121 | x249 ;
  assign n1621 = n1613 & n1620 ;
  assign n1622 = n1619 | n1621 ;
  assign n1623 = n1609 & n1620 ;
  assign n1624 = n1619 | n1623 ;
  assign n1625 = ( n1604 & n1622 ) | ( n1604 & n1624 ) | ( n1622 & n1624 ) ;
  assign n1626 = n1619 | n1620 ;
  assign n1627 = ( n1611 & n1624 ) | ( n1611 & n1626 ) | ( n1624 & n1626 ) ;
  assign n1628 = ( n1573 & n1625 ) | ( n1573 & n1627 ) | ( n1625 & n1627 ) ;
  assign n1629 = ( x122 & ~x250 ) | ( x122 & n1628 ) | ( ~x250 & n1628 ) ;
  assign n1630 = ( ~x122 & x250 ) | ( ~x122 & n1629 ) | ( x250 & n1629 ) ;
  assign n1631 = ( ~n1628 & n1629 ) | ( ~n1628 & n1630 ) | ( n1629 & n1630 ) ;
  assign n1632 = x122 & x250 ;
  assign n1633 = x122 | x250 ;
  assign n1634 = n1627 & n1633 ;
  assign n1635 = n1632 | n1634 ;
  assign n1636 = n1632 | n1633 ;
  assign n1637 = ( n1625 & n1632 ) | ( n1625 & n1636 ) | ( n1632 & n1636 ) ;
  assign n1638 = ( n1573 & n1635 ) | ( n1573 & n1637 ) | ( n1635 & n1637 ) ;
  assign n1639 = ( x123 & ~x251 ) | ( x123 & n1638 ) | ( ~x251 & n1638 ) ;
  assign n1640 = ( ~x123 & x251 ) | ( ~x123 & n1639 ) | ( x251 & n1639 ) ;
  assign n1641 = ( ~n1638 & n1639 ) | ( ~n1638 & n1640 ) | ( n1639 & n1640 ) ;
  assign n1642 = x123 & x251 ;
  assign n1643 = x123 | x251 ;
  assign n1644 = n1636 & n1643 ;
  assign n1645 = n1642 | n1644 ;
  assign n1646 = n1632 & n1643 ;
  assign n1647 = n1642 | n1646 ;
  assign n1648 = ( n1625 & n1645 ) | ( n1625 & n1647 ) | ( n1645 & n1647 ) ;
  assign n1649 = n1642 | n1643 ;
  assign n1650 = ( n1634 & n1647 ) | ( n1634 & n1649 ) | ( n1647 & n1649 ) ;
  assign n1651 = ( n1573 & n1648 ) | ( n1573 & n1650 ) | ( n1648 & n1650 ) ;
  assign n1652 = ( x124 & ~x252 ) | ( x124 & n1651 ) | ( ~x252 & n1651 ) ;
  assign n1653 = ( ~x124 & x252 ) | ( ~x124 & n1652 ) | ( x252 & n1652 ) ;
  assign n1654 = ( ~n1651 & n1652 ) | ( ~n1651 & n1653 ) | ( n1652 & n1653 ) ;
  assign n1655 = x124 & x252 ;
  assign n1656 = x124 | x252 ;
  assign n1657 = n1648 & n1656 ;
  assign n1658 = n1655 | n1657 ;
  assign n1659 = n1647 & n1656 ;
  assign n1660 = n1649 & n1656 ;
  assign n1661 = ( n1634 & n1659 ) | ( n1634 & n1660 ) | ( n1659 & n1660 ) ;
  assign n1662 = n1655 | n1661 ;
  assign n1663 = ( n1573 & n1658 ) | ( n1573 & n1662 ) | ( n1658 & n1662 ) ;
  assign n1664 = ( x125 & ~x253 ) | ( x125 & n1663 ) | ( ~x253 & n1663 ) ;
  assign n1665 = ( ~x125 & x253 ) | ( ~x125 & n1664 ) | ( x253 & n1664 ) ;
  assign n1666 = ( ~n1663 & n1664 ) | ( ~n1663 & n1665 ) | ( n1664 & n1665 ) ;
  assign n1667 = x125 & x253 ;
  assign n1668 = x125 | x253 ;
  assign n1669 = n1655 & n1668 ;
  assign n1670 = n1667 | n1669 ;
  assign n1671 = n1667 | n1668 ;
  assign n1672 = ( n1657 & n1670 ) | ( n1657 & n1671 ) | ( n1670 & n1671 ) ;
  assign n1673 = ( n1662 & n1667 ) | ( n1662 & n1671 ) | ( n1667 & n1671 ) ;
  assign n1674 = ( n1573 & n1672 ) | ( n1573 & n1673 ) | ( n1672 & n1673 ) ;
  assign n1675 = ( x126 & ~x254 ) | ( x126 & n1674 ) | ( ~x254 & n1674 ) ;
  assign n1676 = ( ~x126 & x254 ) | ( ~x126 & n1675 ) | ( x254 & n1675 ) ;
  assign n1677 = ( ~n1674 & n1675 ) | ( ~n1674 & n1676 ) | ( n1675 & n1676 ) ;
  assign n1678 = x126 & x254 ;
  assign n1679 = x126 | x254 ;
  assign n1680 = n1670 & n1679 ;
  assign n1681 = n1678 | n1680 ;
  assign n1682 = n1671 & n1679 ;
  assign n1683 = n1678 | n1682 ;
  assign n1684 = ( n1657 & n1681 ) | ( n1657 & n1683 ) | ( n1681 & n1683 ) ;
  assign n1685 = n1667 & n1679 ;
  assign n1686 = n1678 | n1685 ;
  assign n1687 = ( n1662 & n1683 ) | ( n1662 & n1686 ) | ( n1683 & n1686 ) ;
  assign n1688 = ( n1573 & n1684 ) | ( n1573 & n1687 ) | ( n1684 & n1687 ) ;
  assign n1689 = x127 | x255 ;
  assign n1690 = x127 & x255 ;
  assign n1691 = n1689 & ~n1690 ;
  assign n1692 = n1688 & n1691 ;
  assign n1693 = n1691 & ~n1692 ;
  assign n1694 = ( n1688 & ~n1692 ) | ( n1688 & n1693 ) | ( ~n1692 & n1693 ) ;
  assign n1695 = ( n1570 & n1684 ) | ( n1570 & n1687 ) | ( n1684 & n1687 ) ;
  assign n1696 = ( n1569 & n1684 ) | ( n1569 & n1687 ) | ( n1684 & n1687 ) ;
  assign n1697 = ( n1209 & n1695 ) | ( n1209 & n1696 ) | ( n1695 & n1696 ) ;
  assign n1698 = ( x127 & x255 ) | ( x127 & n1697 ) | ( x255 & n1697 ) ;
  assign y0 = n259 ;
  assign y1 = n263 ;
  assign y2 = n270 ;
  assign y3 = n281 ;
  assign y4 = n286 ;
  assign y5 = n293 ;
  assign y6 = n303 ;
  assign y7 = n310 ;
  assign y8 = n320 ;
  assign y9 = n333 ;
  assign y10 = n337 ;
  assign y11 = n349 ;
  assign y12 = n364 ;
  assign y13 = n368 ;
  assign y14 = n383 ;
  assign y15 = n391 ;
  assign y16 = n398 ;
  assign y17 = n408 ;
  assign y18 = n419 ;
  assign y19 = n434 ;
  assign y20 = n441 ;
  assign y21 = n451 ;
  assign y22 = n462 ;
  assign y23 = n475 ;
  assign y24 = n488 ;
  assign y25 = n492 ;
  assign y26 = n507 ;
  assign y27 = n515 ;
  assign y28 = n529 ;
  assign y29 = n544 ;
  assign y30 = n548 ;
  assign y31 = n563 ;
  assign y32 = n571 ;
  assign y33 = n583 ;
  assign y34 = n597 ;
  assign y35 = n604 ;
  assign y36 = n614 ;
  assign y37 = n625 ;
  assign y38 = n638 ;
  assign y39 = n649 ;
  assign y40 = n663 ;
  assign y41 = n670 ;
  assign y42 = n680 ;
  assign y43 = n691 ;
  assign y44 = n704 ;
  assign y45 = n715 ;
  assign y46 = n729 ;
  assign y47 = n744 ;
  assign y48 = n748 ;
  assign y49 = n763 ;
  assign y50 = n771 ;
  assign y51 = n783 ;
  assign y52 = n795 ;
  assign y53 = n809 ;
  assign y54 = n824 ;
  assign y55 = n828 ;
  assign y56 = n843 ;
  assign y57 = n851 ;
  assign y58 = n863 ;
  assign y59 = n875 ;
  assign y60 = n887 ;
  assign y61 = n901 ;
  assign y62 = n908 ;
  assign y63 = n918 ;
  assign y64 = n929 ;
  assign y65 = n942 ;
  assign y66 = n953 ;
  assign y67 = n967 ;
  assign y68 = n978 ;
  assign y69 = n994 ;
  assign y70 = n1001 ;
  assign y71 = n1011 ;
  assign y72 = n1022 ;
  assign y73 = n1035 ;
  assign y74 = n1046 ;
  assign y75 = n1060 ;
  assign y76 = n1071 ;
  assign y77 = n1085 ;
  assign y78 = n1102 ;
  assign y79 = n1106 ;
  assign y80 = n1121 ;
  assign y81 = n1129 ;
  assign y82 = n1141 ;
  assign y83 = n1153 ;
  assign y84 = n1165 ;
  assign y85 = n1179 ;
  assign y86 = n1193 ;
  assign y87 = n1213 ;
  assign y88 = n1217 ;
  assign y89 = n1232 ;
  assign y90 = n1240 ;
  assign y91 = n1252 ;
  assign y92 = n1264 ;
  assign y93 = n1276 ;
  assign y94 = n1290 ;
  assign y95 = n1307 ;
  assign y96 = n1318 ;
  assign y97 = n1325 ;
  assign y98 = n1335 ;
  assign y99 = n1346 ;
  assign y100 = n1359 ;
  assign y101 = n1370 ;
  assign y102 = n1384 ;
  assign y103 = n1395 ;
  assign y104 = n1409 ;
  assign y105 = n1421 ;
  assign y106 = n1439 ;
  assign y107 = n1446 ;
  assign y108 = n1456 ;
  assign y109 = n1467 ;
  assign y110 = n1480 ;
  assign y111 = n1491 ;
  assign y112 = n1505 ;
  assign y113 = n1516 ;
  assign y114 = n1530 ;
  assign y115 = n1542 ;
  assign y116 = n1556 ;
  assign y117 = n1577 ;
  assign y118 = n1586 ;
  assign y119 = n1601 ;
  assign y120 = n1608 ;
  assign y121 = n1618 ;
  assign y122 = n1631 ;
  assign y123 = n1641 ;
  assign y124 = n1654 ;
  assign y125 = n1666 ;
  assign y126 = n1677 ;
  assign y127 = n1694 ;
  assign y128 = n1698 ;
endmodule
