module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 , x147 , x148 , x149 , x150 , x151 , x152 , x153 , x154 , x155 , x156 , x157 , x158 , x159 , x160 , x161 , x162 , x163 , x164 , x165 , x166 , x167 , x168 , x169 , x170 , x171 , x172 , x173 , x174 , x175 , x176 , x177 , x178 , x179 , x180 , x181 , x182 , x183 , x184 , x185 , x186 , x187 , x188 , x189 , x190 , x191 , x192 , x193 , x194 , x195 , x196 , x197 , x198 , x199 , x200 , x201 , x202 , x203 , x204 , x205 , x206 , x207 , x208 , x209 , x210 , x211 , x212 , x213 , x214 , x215 , x216 , x217 , x218 , x219 , x220 , x221 , x222 , x223 , x224 , x225 , x226 , x227 , x228 , x229 , x230 , x231 , x232 , x233 , x234 , x235 , x236 , x237 , x238 , x239 , x240 , x241 , x242 , x243 , x244 , x245 , x246 , x247 , x248 , x249 , x250 , x251 , x252 , x253 , x254 , x255 , x256 , x257 , x258 , x259 , x260 , x261 , x262 , x263 , x264 , x265 , x266 , x267 , x268 , x269 , x270 , x271 , x272 , x273 , x274 , x275 , x276 , x277 , x278 , x279 , x280 , x281 , x282 , x283 , x284 , x285 , x286 , x287 , x288 , x289 , x290 , x291 , x292 , x293 , x294 , x295 , x296 , x297 , x298 , x299 , x300 , x301 , x302 , x303 , x304 , x305 , x306 , x307 , x308 , x309 , x310 , x311 , x312 , x313 , x314 , x315 , x316 , x317 , x318 , x319 , x320 , x321 , x322 , x323 , x324 , x325 , x326 , x327 , x328 , x329 , x330 , x331 , x332 , x333 , x334 , x335 , x336 , x337 , x338 , x339 , x340 , x341 , x342 , x343 , x344 , x345 , x346 , x347 , x348 , x349 , x350 , x351 , x352 , x353 , x354 , x355 , x356 , x357 , x358 , x359 , x360 , x361 , x362 , x363 , x364 , x365 , x366 , x367 , x368 , x369 , x370 , x371 , x372 , x373 , x374 , x375 , x376 , x377 , x378 , x379 , x380 , x381 , x382 , x383 , x384 , x385 , x386 , x387 , x388 , x389 , x390 , x391 , x392 , x393 , x394 , x395 , x396 , x397 , x398 , x399 , x400 , x401 , x402 , x403 , x404 , x405 , x406 , x407 , x408 , x409 , x410 , x411 , x412 , x413 , x414 , x415 , x416 , x417 , x418 , x419 , x420 , x421 , x422 , x423 , x424 , x425 , x426 , x427 , x428 , x429 , x430 , x431 , x432 , x433 , x434 , x435 , x436 , x437 , x438 , x439 , x440 , x441 , x442 , x443 , x444 , x445 , x446 , x447 , x448 , x449 , x450 , x451 , x452 , x453 , x454 , x455 , x456 , x457 , x458 , x459 , x460 , x461 , x462 , x463 , x464 , x465 , x466 , x467 , x468 , x469 , x470 , x471 , x472 , x473 , x474 , x475 , x476 , x477 , x478 , x479 , x480 , x481 , x482 , x483 , x484 , x485 , x486 , x487 , x488 , x489 , x490 , x491 , x492 , x493 , x494 , x495 , x496 , x497 , x498 , x499 , x500 , x501 , x502 , x503 , x504 , x505 , x506 , x507 , x508 , x509 , x510 , x511 , x512 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 , y128 , y129 , y130 , y131 , y132 , y133 , y134 , y135 , y136 , y137 , y138 , y139 , y140 , y141 , y142 , y143 , y144 , y145 , y146 , y147 , y148 , y149 , y150 , y151 , y152 , y153 , y154 , y155 , y156 , y157 , y158 , y159 , y160 , y161 , y162 , y163 , y164 , y165 , y166 , y167 , y168 , y169 , y170 , y171 , y172 , y173 , y174 , y175 , y176 , y177 , y178 , y179 , y180 , y181 , y182 , y183 , y184 , y185 , y186 , y187 , y188 , y189 , y190 , y191 , y192 , y193 , y194 , y195 , y196 , y197 , y198 , y199 , y200 , y201 , y202 , y203 , y204 , y205 , y206 , y207 , y208 , y209 , y210 , y211 , y212 , y213 , y214 , y215 , y216 , y217 , y218 , y219 , y220 , y221 , y222 , y223 , y224 , y225 , y226 , y227 , y228 , y229 , y230 , y231 , y232 , y233 , y234 , y235 , y236 , y237 , y238 , y239 , y240 , y241 , y242 , y243 , y244 , y245 , y246 , y247 , y248 , y249 , y250 , y251 , y252 , y253 , y254 , y255 , y256 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 , x147 , x148 , x149 , x150 , x151 , x152 , x153 , x154 , x155 , x156 , x157 , x158 , x159 , x160 , x161 , x162 , x163 , x164 , x165 , x166 , x167 , x168 , x169 , x170 , x171 , x172 , x173 , x174 , x175 , x176 , x177 , x178 , x179 , x180 , x181 , x182 , x183 , x184 , x185 , x186 , x187 , x188 , x189 , x190 , x191 , x192 , x193 , x194 , x195 , x196 , x197 , x198 , x199 , x200 , x201 , x202 , x203 , x204 , x205 , x206 , x207 , x208 , x209 , x210 , x211 , x212 , x213 , x214 , x215 , x216 , x217 , x218 , x219 , x220 , x221 , x222 , x223 , x224 , x225 , x226 , x227 , x228 , x229 , x230 , x231 , x232 , x233 , x234 , x235 , x236 , x237 , x238 , x239 , x240 , x241 , x242 , x243 , x244 , x245 , x246 , x247 , x248 , x249 , x250 , x251 , x252 , x253 , x254 , x255 , x256 , x257 , x258 , x259 , x260 , x261 , x262 , x263 , x264 , x265 , x266 , x267 , x268 , x269 , x270 , x271 , x272 , x273 , x274 , x275 , x276 , x277 , x278 , x279 , x280 , x281 , x282 , x283 , x284 , x285 , x286 , x287 , x288 , x289 , x290 , x291 , x292 , x293 , x294 , x295 , x296 , x297 , x298 , x299 , x300 , x301 , x302 , x303 , x304 , x305 , x306 , x307 , x308 , x309 , x310 , x311 , x312 , x313 , x314 , x315 , x316 , x317 , x318 , x319 , x320 , x321 , x322 , x323 , x324 , x325 , x326 , x327 , x328 , x329 , x330 , x331 , x332 , x333 , x334 , x335 , x336 , x337 , x338 , x339 , x340 , x341 , x342 , x343 , x344 , x345 , x346 , x347 , x348 , x349 , x350 , x351 , x352 , x353 , x354 , x355 , x356 , x357 , x358 , x359 , x360 , x361 , x362 , x363 , x364 , x365 , x366 , x367 , x368 , x369 , x370 , x371 , x372 , x373 , x374 , x375 , x376 , x377 , x378 , x379 , x380 , x381 , x382 , x383 , x384 , x385 , x386 , x387 , x388 , x389 , x390 , x391 , x392 , x393 , x394 , x395 , x396 , x397 , x398 , x399 , x400 , x401 , x402 , x403 , x404 , x405 , x406 , x407 , x408 , x409 , x410 , x411 , x412 , x413 , x414 , x415 , x416 , x417 , x418 , x419 , x420 , x421 , x422 , x423 , x424 , x425 , x426 , x427 , x428 , x429 , x430 , x431 , x432 , x433 , x434 , x435 , x436 , x437 , x438 , x439 , x440 , x441 , x442 , x443 , x444 , x445 , x446 , x447 , x448 , x449 , x450 , x451 , x452 , x453 , x454 , x455 , x456 , x457 , x458 , x459 , x460 , x461 , x462 , x463 , x464 , x465 , x466 , x467 , x468 , x469 , x470 , x471 , x472 , x473 , x474 , x475 , x476 , x477 , x478 , x479 , x480 , x481 , x482 , x483 , x484 , x485 , x486 , x487 , x488 , x489 , x490 , x491 , x492 , x493 , x494 , x495 , x496 , x497 , x498 , x499 , x500 , x501 , x502 , x503 , x504 , x505 , x506 , x507 , x508 , x509 , x510 , x511 , x512 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 , y128 , y129 , y130 , y131 , y132 , y133 , y134 , y135 , y136 , y137 , y138 , y139 , y140 , y141 , y142 , y143 , y144 , y145 , y146 , y147 , y148 , y149 , y150 , y151 , y152 , y153 , y154 , y155 , y156 , y157 , y158 , y159 , y160 , y161 , y162 , y163 , y164 , y165 , y166 , y167 , y168 , y169 , y170 , y171 , y172 , y173 , y174 , y175 , y176 , y177 , y178 , y179 , y180 , y181 , y182 , y183 , y184 , y185 , y186 , y187 , y188 , y189 , y190 , y191 , y192 , y193 , y194 , y195 , y196 , y197 , y198 , y199 , y200 , y201 , y202 , y203 , y204 , y205 , y206 , y207 , y208 , y209 , y210 , y211 , y212 , y213 , y214 , y215 , y216 , y217 , y218 , y219 , y220 , y221 , y222 , y223 , y224 , y225 , y226 , y227 , y228 , y229 , y230 , y231 , y232 , y233 , y234 , y235 , y236 , y237 , y238 , y239 , y240 , y241 , y242 , y243 , y244 , y245 , y246 , y247 , y248 , y249 , y250 , y251 , y252 , y253 , y254 , y255 , y256 ;
  wire n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 ;
  assign n514 = ( x0 & ~x1 ) | ( x0 & x2 ) | ( ~x1 & x2 ) ;
  assign n515 = ( ~x0 & x1 ) | ( ~x0 & n514 ) | ( x1 & n514 ) ;
  assign n516 = ( ~x2 & n514 ) | ( ~x2 & n515 ) | ( n514 & n515 ) ;
  assign n517 = ( x0 & x1 ) | ( x0 & x2 ) | ( x1 & x2 ) ;
  assign n518 = ( x3 & ~x4 ) | ( x3 & n517 ) | ( ~x4 & n517 ) ;
  assign n519 = ( ~x3 & x4 ) | ( ~x3 & n518 ) | ( x4 & n518 ) ;
  assign n520 = ( ~n517 & n518 ) | ( ~n517 & n519 ) | ( n518 & n519 ) ;
  assign n521 = ( x3 & x4 ) | ( x3 & n517 ) | ( x4 & n517 ) ;
  assign n522 = ( x5 & ~x6 ) | ( x5 & n521 ) | ( ~x6 & n521 ) ;
  assign n523 = ( ~x5 & x6 ) | ( ~x5 & n522 ) | ( x6 & n522 ) ;
  assign n524 = ( ~n521 & n522 ) | ( ~n521 & n523 ) | ( n522 & n523 ) ;
  assign n525 = ( x5 & x6 ) | ( x5 & n521 ) | ( x6 & n521 ) ;
  assign n526 = ( x7 & ~x8 ) | ( x7 & n525 ) | ( ~x8 & n525 ) ;
  assign n527 = ( ~x7 & x8 ) | ( ~x7 & n526 ) | ( x8 & n526 ) ;
  assign n528 = ( ~n525 & n526 ) | ( ~n525 & n527 ) | ( n526 & n527 ) ;
  assign n529 = ( x7 & x8 ) | ( x7 & n525 ) | ( x8 & n525 ) ;
  assign n530 = ( x9 & ~x10 ) | ( x9 & n529 ) | ( ~x10 & n529 ) ;
  assign n531 = ( ~x9 & x10 ) | ( ~x9 & n530 ) | ( x10 & n530 ) ;
  assign n532 = ( ~n529 & n530 ) | ( ~n529 & n531 ) | ( n530 & n531 ) ;
  assign n533 = ( x9 & x10 ) | ( x9 & n529 ) | ( x10 & n529 ) ;
  assign n534 = ( x11 & ~x12 ) | ( x11 & n533 ) | ( ~x12 & n533 ) ;
  assign n535 = ( ~x11 & x12 ) | ( ~x11 & n534 ) | ( x12 & n534 ) ;
  assign n536 = ( ~n533 & n534 ) | ( ~n533 & n535 ) | ( n534 & n535 ) ;
  assign n537 = ( x11 & x12 ) | ( x11 & n533 ) | ( x12 & n533 ) ;
  assign n538 = ( x13 & ~x14 ) | ( x13 & n537 ) | ( ~x14 & n537 ) ;
  assign n539 = ( ~x13 & x14 ) | ( ~x13 & n538 ) | ( x14 & n538 ) ;
  assign n540 = ( ~n537 & n538 ) | ( ~n537 & n539 ) | ( n538 & n539 ) ;
  assign n541 = ( x13 & x14 ) | ( x13 & n537 ) | ( x14 & n537 ) ;
  assign n542 = ( x15 & ~x16 ) | ( x15 & n541 ) | ( ~x16 & n541 ) ;
  assign n543 = ( ~x15 & x16 ) | ( ~x15 & n542 ) | ( x16 & n542 ) ;
  assign n544 = ( ~n541 & n542 ) | ( ~n541 & n543 ) | ( n542 & n543 ) ;
  assign n545 = ( x15 & x16 ) | ( x15 & n541 ) | ( x16 & n541 ) ;
  assign n546 = ( x17 & ~x18 ) | ( x17 & n545 ) | ( ~x18 & n545 ) ;
  assign n547 = ( ~x17 & x18 ) | ( ~x17 & n546 ) | ( x18 & n546 ) ;
  assign n548 = ( ~n545 & n546 ) | ( ~n545 & n547 ) | ( n546 & n547 ) ;
  assign n549 = ( x17 & x18 ) | ( x17 & n545 ) | ( x18 & n545 ) ;
  assign n550 = ( x19 & ~x20 ) | ( x19 & n549 ) | ( ~x20 & n549 ) ;
  assign n551 = ( ~x19 & x20 ) | ( ~x19 & n550 ) | ( x20 & n550 ) ;
  assign n552 = ( ~n549 & n550 ) | ( ~n549 & n551 ) | ( n550 & n551 ) ;
  assign n553 = ( x19 & x20 ) | ( x19 & n549 ) | ( x20 & n549 ) ;
  assign n554 = ( x21 & ~x22 ) | ( x21 & n553 ) | ( ~x22 & n553 ) ;
  assign n555 = ( ~x21 & x22 ) | ( ~x21 & n554 ) | ( x22 & n554 ) ;
  assign n556 = ( ~n553 & n554 ) | ( ~n553 & n555 ) | ( n554 & n555 ) ;
  assign n557 = ( x21 & x22 ) | ( x21 & n553 ) | ( x22 & n553 ) ;
  assign n558 = ( x23 & ~x24 ) | ( x23 & n557 ) | ( ~x24 & n557 ) ;
  assign n559 = ( ~x23 & x24 ) | ( ~x23 & n558 ) | ( x24 & n558 ) ;
  assign n560 = ( ~n557 & n558 ) | ( ~n557 & n559 ) | ( n558 & n559 ) ;
  assign n561 = ( x23 & x24 ) | ( x23 & n557 ) | ( x24 & n557 ) ;
  assign n562 = ( x25 & ~x26 ) | ( x25 & n561 ) | ( ~x26 & n561 ) ;
  assign n563 = ( ~x25 & x26 ) | ( ~x25 & n562 ) | ( x26 & n562 ) ;
  assign n564 = ( ~n561 & n562 ) | ( ~n561 & n563 ) | ( n562 & n563 ) ;
  assign n565 = ( x25 & x26 ) | ( x25 & n561 ) | ( x26 & n561 ) ;
  assign n566 = ( x27 & ~x28 ) | ( x27 & n565 ) | ( ~x28 & n565 ) ;
  assign n567 = ( ~x27 & x28 ) | ( ~x27 & n566 ) | ( x28 & n566 ) ;
  assign n568 = ( ~n565 & n566 ) | ( ~n565 & n567 ) | ( n566 & n567 ) ;
  assign n569 = ( x27 & x28 ) | ( x27 & n565 ) | ( x28 & n565 ) ;
  assign n570 = ( x29 & ~x30 ) | ( x29 & n569 ) | ( ~x30 & n569 ) ;
  assign n571 = ( ~x29 & x30 ) | ( ~x29 & n570 ) | ( x30 & n570 ) ;
  assign n572 = ( ~n569 & n570 ) | ( ~n569 & n571 ) | ( n570 & n571 ) ;
  assign n573 = ( x29 & x30 ) | ( x29 & n569 ) | ( x30 & n569 ) ;
  assign n574 = ( x31 & ~x32 ) | ( x31 & n573 ) | ( ~x32 & n573 ) ;
  assign n575 = ( ~x31 & x32 ) | ( ~x31 & n574 ) | ( x32 & n574 ) ;
  assign n576 = ( ~n573 & n574 ) | ( ~n573 & n575 ) | ( n574 & n575 ) ;
  assign n577 = ( x31 & x32 ) | ( x31 & n573 ) | ( x32 & n573 ) ;
  assign n578 = ( x33 & ~x34 ) | ( x33 & n577 ) | ( ~x34 & n577 ) ;
  assign n579 = ( ~x33 & x34 ) | ( ~x33 & n578 ) | ( x34 & n578 ) ;
  assign n580 = ( ~n577 & n578 ) | ( ~n577 & n579 ) | ( n578 & n579 ) ;
  assign n581 = ( x33 & x34 ) | ( x33 & n577 ) | ( x34 & n577 ) ;
  assign n582 = ( x35 & ~x36 ) | ( x35 & n581 ) | ( ~x36 & n581 ) ;
  assign n583 = ( ~x35 & x36 ) | ( ~x35 & n582 ) | ( x36 & n582 ) ;
  assign n584 = ( ~n581 & n582 ) | ( ~n581 & n583 ) | ( n582 & n583 ) ;
  assign n585 = ( x35 & x36 ) | ( x35 & n581 ) | ( x36 & n581 ) ;
  assign n586 = ( x37 & ~x38 ) | ( x37 & n585 ) | ( ~x38 & n585 ) ;
  assign n587 = ( ~x37 & x38 ) | ( ~x37 & n586 ) | ( x38 & n586 ) ;
  assign n588 = ( ~n585 & n586 ) | ( ~n585 & n587 ) | ( n586 & n587 ) ;
  assign n589 = ( x37 & x38 ) | ( x37 & n585 ) | ( x38 & n585 ) ;
  assign n590 = ( x39 & ~x40 ) | ( x39 & n589 ) | ( ~x40 & n589 ) ;
  assign n591 = ( ~x39 & x40 ) | ( ~x39 & n590 ) | ( x40 & n590 ) ;
  assign n592 = ( ~n589 & n590 ) | ( ~n589 & n591 ) | ( n590 & n591 ) ;
  assign n593 = ( x39 & x40 ) | ( x39 & n589 ) | ( x40 & n589 ) ;
  assign n594 = ( x41 & ~x42 ) | ( x41 & n593 ) | ( ~x42 & n593 ) ;
  assign n595 = ( ~x41 & x42 ) | ( ~x41 & n594 ) | ( x42 & n594 ) ;
  assign n596 = ( ~n593 & n594 ) | ( ~n593 & n595 ) | ( n594 & n595 ) ;
  assign n597 = ( x41 & x42 ) | ( x41 & n593 ) | ( x42 & n593 ) ;
  assign n598 = ( x43 & ~x44 ) | ( x43 & n597 ) | ( ~x44 & n597 ) ;
  assign n599 = ( ~x43 & x44 ) | ( ~x43 & n598 ) | ( x44 & n598 ) ;
  assign n600 = ( ~n597 & n598 ) | ( ~n597 & n599 ) | ( n598 & n599 ) ;
  assign n601 = ( x43 & x44 ) | ( x43 & n597 ) | ( x44 & n597 ) ;
  assign n602 = ( x45 & ~x46 ) | ( x45 & n601 ) | ( ~x46 & n601 ) ;
  assign n603 = ( ~x45 & x46 ) | ( ~x45 & n602 ) | ( x46 & n602 ) ;
  assign n604 = ( ~n601 & n602 ) | ( ~n601 & n603 ) | ( n602 & n603 ) ;
  assign n605 = ( x45 & x46 ) | ( x45 & n601 ) | ( x46 & n601 ) ;
  assign n606 = ( x47 & ~x48 ) | ( x47 & n605 ) | ( ~x48 & n605 ) ;
  assign n607 = ( ~x47 & x48 ) | ( ~x47 & n606 ) | ( x48 & n606 ) ;
  assign n608 = ( ~n605 & n606 ) | ( ~n605 & n607 ) | ( n606 & n607 ) ;
  assign n609 = ( x47 & x48 ) | ( x47 & n605 ) | ( x48 & n605 ) ;
  assign n610 = ( x49 & ~x50 ) | ( x49 & n609 ) | ( ~x50 & n609 ) ;
  assign n611 = ( ~x49 & x50 ) | ( ~x49 & n610 ) | ( x50 & n610 ) ;
  assign n612 = ( ~n609 & n610 ) | ( ~n609 & n611 ) | ( n610 & n611 ) ;
  assign n613 = ( x49 & x50 ) | ( x49 & n609 ) | ( x50 & n609 ) ;
  assign n614 = ( x51 & ~x52 ) | ( x51 & n613 ) | ( ~x52 & n613 ) ;
  assign n615 = ( ~x51 & x52 ) | ( ~x51 & n614 ) | ( x52 & n614 ) ;
  assign n616 = ( ~n613 & n614 ) | ( ~n613 & n615 ) | ( n614 & n615 ) ;
  assign n617 = ( x51 & x52 ) | ( x51 & n613 ) | ( x52 & n613 ) ;
  assign n618 = ( x53 & ~x54 ) | ( x53 & n617 ) | ( ~x54 & n617 ) ;
  assign n619 = ( ~x53 & x54 ) | ( ~x53 & n618 ) | ( x54 & n618 ) ;
  assign n620 = ( ~n617 & n618 ) | ( ~n617 & n619 ) | ( n618 & n619 ) ;
  assign n621 = ( x53 & x54 ) | ( x53 & n617 ) | ( x54 & n617 ) ;
  assign n622 = ( x55 & ~x56 ) | ( x55 & n621 ) | ( ~x56 & n621 ) ;
  assign n623 = ( ~x55 & x56 ) | ( ~x55 & n622 ) | ( x56 & n622 ) ;
  assign n624 = ( ~n621 & n622 ) | ( ~n621 & n623 ) | ( n622 & n623 ) ;
  assign n625 = ( x55 & x56 ) | ( x55 & n621 ) | ( x56 & n621 ) ;
  assign n626 = ( x57 & ~x58 ) | ( x57 & n625 ) | ( ~x58 & n625 ) ;
  assign n627 = ( ~x57 & x58 ) | ( ~x57 & n626 ) | ( x58 & n626 ) ;
  assign n628 = ( ~n625 & n626 ) | ( ~n625 & n627 ) | ( n626 & n627 ) ;
  assign n629 = ( x57 & x58 ) | ( x57 & n625 ) | ( x58 & n625 ) ;
  assign n630 = ( x59 & ~x60 ) | ( x59 & n629 ) | ( ~x60 & n629 ) ;
  assign n631 = ( ~x59 & x60 ) | ( ~x59 & n630 ) | ( x60 & n630 ) ;
  assign n632 = ( ~n629 & n630 ) | ( ~n629 & n631 ) | ( n630 & n631 ) ;
  assign n633 = ( x59 & x60 ) | ( x59 & n629 ) | ( x60 & n629 ) ;
  assign n634 = ( x61 & ~x62 ) | ( x61 & n633 ) | ( ~x62 & n633 ) ;
  assign n635 = ( ~x61 & x62 ) | ( ~x61 & n634 ) | ( x62 & n634 ) ;
  assign n636 = ( ~n633 & n634 ) | ( ~n633 & n635 ) | ( n634 & n635 ) ;
  assign n637 = ( x61 & x62 ) | ( x61 & n633 ) | ( x62 & n633 ) ;
  assign n638 = ( x63 & ~x64 ) | ( x63 & n637 ) | ( ~x64 & n637 ) ;
  assign n639 = ( ~x63 & x64 ) | ( ~x63 & n638 ) | ( x64 & n638 ) ;
  assign n640 = ( ~n637 & n638 ) | ( ~n637 & n639 ) | ( n638 & n639 ) ;
  assign n641 = ( x63 & x64 ) | ( x63 & n637 ) | ( x64 & n637 ) ;
  assign n642 = ( x65 & ~x66 ) | ( x65 & n641 ) | ( ~x66 & n641 ) ;
  assign n643 = ( ~x65 & x66 ) | ( ~x65 & n642 ) | ( x66 & n642 ) ;
  assign n644 = ( ~n641 & n642 ) | ( ~n641 & n643 ) | ( n642 & n643 ) ;
  assign n645 = ( x65 & x66 ) | ( x65 & n641 ) | ( x66 & n641 ) ;
  assign n646 = ( x67 & ~x68 ) | ( x67 & n645 ) | ( ~x68 & n645 ) ;
  assign n647 = ( ~x67 & x68 ) | ( ~x67 & n646 ) | ( x68 & n646 ) ;
  assign n648 = ( ~n645 & n646 ) | ( ~n645 & n647 ) | ( n646 & n647 ) ;
  assign n649 = ( x67 & x68 ) | ( x67 & n645 ) | ( x68 & n645 ) ;
  assign n650 = ( x69 & ~x70 ) | ( x69 & n649 ) | ( ~x70 & n649 ) ;
  assign n651 = ( ~x69 & x70 ) | ( ~x69 & n650 ) | ( x70 & n650 ) ;
  assign n652 = ( ~n649 & n650 ) | ( ~n649 & n651 ) | ( n650 & n651 ) ;
  assign n653 = ( x69 & x70 ) | ( x69 & n649 ) | ( x70 & n649 ) ;
  assign n654 = ( x71 & ~x72 ) | ( x71 & n653 ) | ( ~x72 & n653 ) ;
  assign n655 = ( ~x71 & x72 ) | ( ~x71 & n654 ) | ( x72 & n654 ) ;
  assign n656 = ( ~n653 & n654 ) | ( ~n653 & n655 ) | ( n654 & n655 ) ;
  assign n657 = ( x71 & x72 ) | ( x71 & n653 ) | ( x72 & n653 ) ;
  assign n658 = ( x73 & ~x74 ) | ( x73 & n657 ) | ( ~x74 & n657 ) ;
  assign n659 = ( ~x73 & x74 ) | ( ~x73 & n658 ) | ( x74 & n658 ) ;
  assign n660 = ( ~n657 & n658 ) | ( ~n657 & n659 ) | ( n658 & n659 ) ;
  assign n661 = ( x73 & x74 ) | ( x73 & n657 ) | ( x74 & n657 ) ;
  assign n662 = ( x75 & ~x76 ) | ( x75 & n661 ) | ( ~x76 & n661 ) ;
  assign n663 = ( ~x75 & x76 ) | ( ~x75 & n662 ) | ( x76 & n662 ) ;
  assign n664 = ( ~n661 & n662 ) | ( ~n661 & n663 ) | ( n662 & n663 ) ;
  assign n665 = ( x75 & x76 ) | ( x75 & n661 ) | ( x76 & n661 ) ;
  assign n666 = ( x77 & ~x78 ) | ( x77 & n665 ) | ( ~x78 & n665 ) ;
  assign n667 = ( ~x77 & x78 ) | ( ~x77 & n666 ) | ( x78 & n666 ) ;
  assign n668 = ( ~n665 & n666 ) | ( ~n665 & n667 ) | ( n666 & n667 ) ;
  assign n669 = ( x77 & x78 ) | ( x77 & n665 ) | ( x78 & n665 ) ;
  assign n670 = ( x79 & ~x80 ) | ( x79 & n669 ) | ( ~x80 & n669 ) ;
  assign n671 = ( ~x79 & x80 ) | ( ~x79 & n670 ) | ( x80 & n670 ) ;
  assign n672 = ( ~n669 & n670 ) | ( ~n669 & n671 ) | ( n670 & n671 ) ;
  assign n673 = ( x79 & x80 ) | ( x79 & n669 ) | ( x80 & n669 ) ;
  assign n674 = ( x81 & ~x82 ) | ( x81 & n673 ) | ( ~x82 & n673 ) ;
  assign n675 = ( ~x81 & x82 ) | ( ~x81 & n674 ) | ( x82 & n674 ) ;
  assign n676 = ( ~n673 & n674 ) | ( ~n673 & n675 ) | ( n674 & n675 ) ;
  assign n677 = ( x81 & x82 ) | ( x81 & n673 ) | ( x82 & n673 ) ;
  assign n678 = ( x83 & ~x84 ) | ( x83 & n677 ) | ( ~x84 & n677 ) ;
  assign n679 = ( ~x83 & x84 ) | ( ~x83 & n678 ) | ( x84 & n678 ) ;
  assign n680 = ( ~n677 & n678 ) | ( ~n677 & n679 ) | ( n678 & n679 ) ;
  assign n681 = ( x83 & x84 ) | ( x83 & n677 ) | ( x84 & n677 ) ;
  assign n682 = ( x85 & ~x86 ) | ( x85 & n681 ) | ( ~x86 & n681 ) ;
  assign n683 = ( ~x85 & x86 ) | ( ~x85 & n682 ) | ( x86 & n682 ) ;
  assign n684 = ( ~n681 & n682 ) | ( ~n681 & n683 ) | ( n682 & n683 ) ;
  assign n685 = ( x85 & x86 ) | ( x85 & n681 ) | ( x86 & n681 ) ;
  assign n686 = ( x87 & ~x88 ) | ( x87 & n685 ) | ( ~x88 & n685 ) ;
  assign n687 = ( ~x87 & x88 ) | ( ~x87 & n686 ) | ( x88 & n686 ) ;
  assign n688 = ( ~n685 & n686 ) | ( ~n685 & n687 ) | ( n686 & n687 ) ;
  assign n689 = ( x87 & x88 ) | ( x87 & n685 ) | ( x88 & n685 ) ;
  assign n690 = ( x89 & ~x90 ) | ( x89 & n689 ) | ( ~x90 & n689 ) ;
  assign n691 = ( ~x89 & x90 ) | ( ~x89 & n690 ) | ( x90 & n690 ) ;
  assign n692 = ( ~n689 & n690 ) | ( ~n689 & n691 ) | ( n690 & n691 ) ;
  assign n693 = ( x89 & x90 ) | ( x89 & n689 ) | ( x90 & n689 ) ;
  assign n694 = ( x91 & ~x92 ) | ( x91 & n693 ) | ( ~x92 & n693 ) ;
  assign n695 = ( ~x91 & x92 ) | ( ~x91 & n694 ) | ( x92 & n694 ) ;
  assign n696 = ( ~n693 & n694 ) | ( ~n693 & n695 ) | ( n694 & n695 ) ;
  assign n697 = ( x91 & x92 ) | ( x91 & n693 ) | ( x92 & n693 ) ;
  assign n698 = ( x93 & ~x94 ) | ( x93 & n697 ) | ( ~x94 & n697 ) ;
  assign n699 = ( ~x93 & x94 ) | ( ~x93 & n698 ) | ( x94 & n698 ) ;
  assign n700 = ( ~n697 & n698 ) | ( ~n697 & n699 ) | ( n698 & n699 ) ;
  assign n701 = ( x93 & x94 ) | ( x93 & n697 ) | ( x94 & n697 ) ;
  assign n702 = ( x95 & ~x96 ) | ( x95 & n701 ) | ( ~x96 & n701 ) ;
  assign n703 = ( ~x95 & x96 ) | ( ~x95 & n702 ) | ( x96 & n702 ) ;
  assign n704 = ( ~n701 & n702 ) | ( ~n701 & n703 ) | ( n702 & n703 ) ;
  assign n705 = ( x95 & x96 ) | ( x95 & n701 ) | ( x96 & n701 ) ;
  assign n706 = ( x97 & ~x98 ) | ( x97 & n705 ) | ( ~x98 & n705 ) ;
  assign n707 = ( ~x97 & x98 ) | ( ~x97 & n706 ) | ( x98 & n706 ) ;
  assign n708 = ( ~n705 & n706 ) | ( ~n705 & n707 ) | ( n706 & n707 ) ;
  assign n709 = ( x97 & x98 ) | ( x97 & n705 ) | ( x98 & n705 ) ;
  assign n710 = ( x99 & ~x100 ) | ( x99 & n709 ) | ( ~x100 & n709 ) ;
  assign n711 = ( ~x99 & x100 ) | ( ~x99 & n710 ) | ( x100 & n710 ) ;
  assign n712 = ( ~n709 & n710 ) | ( ~n709 & n711 ) | ( n710 & n711 ) ;
  assign n713 = ( x99 & x100 ) | ( x99 & n709 ) | ( x100 & n709 ) ;
  assign n714 = ( x101 & ~x102 ) | ( x101 & n713 ) | ( ~x102 & n713 ) ;
  assign n715 = ( ~x101 & x102 ) | ( ~x101 & n714 ) | ( x102 & n714 ) ;
  assign n716 = ( ~n713 & n714 ) | ( ~n713 & n715 ) | ( n714 & n715 ) ;
  assign n717 = ( x101 & x102 ) | ( x101 & n713 ) | ( x102 & n713 ) ;
  assign n718 = ( x103 & ~x104 ) | ( x103 & n717 ) | ( ~x104 & n717 ) ;
  assign n719 = ( ~x103 & x104 ) | ( ~x103 & n718 ) | ( x104 & n718 ) ;
  assign n720 = ( ~n717 & n718 ) | ( ~n717 & n719 ) | ( n718 & n719 ) ;
  assign n721 = ( x103 & x104 ) | ( x103 & n717 ) | ( x104 & n717 ) ;
  assign n722 = ( x105 & ~x106 ) | ( x105 & n721 ) | ( ~x106 & n721 ) ;
  assign n723 = ( ~x105 & x106 ) | ( ~x105 & n722 ) | ( x106 & n722 ) ;
  assign n724 = ( ~n721 & n722 ) | ( ~n721 & n723 ) | ( n722 & n723 ) ;
  assign n725 = ( x105 & x106 ) | ( x105 & n721 ) | ( x106 & n721 ) ;
  assign n726 = ( x107 & ~x108 ) | ( x107 & n725 ) | ( ~x108 & n725 ) ;
  assign n727 = ( ~x107 & x108 ) | ( ~x107 & n726 ) | ( x108 & n726 ) ;
  assign n728 = ( ~n725 & n726 ) | ( ~n725 & n727 ) | ( n726 & n727 ) ;
  assign n729 = ( x107 & x108 ) | ( x107 & n725 ) | ( x108 & n725 ) ;
  assign n730 = ( x109 & ~x110 ) | ( x109 & n729 ) | ( ~x110 & n729 ) ;
  assign n731 = ( ~x109 & x110 ) | ( ~x109 & n730 ) | ( x110 & n730 ) ;
  assign n732 = ( ~n729 & n730 ) | ( ~n729 & n731 ) | ( n730 & n731 ) ;
  assign n733 = ( x109 & x110 ) | ( x109 & n729 ) | ( x110 & n729 ) ;
  assign n734 = ( x111 & ~x112 ) | ( x111 & n733 ) | ( ~x112 & n733 ) ;
  assign n735 = ( ~x111 & x112 ) | ( ~x111 & n734 ) | ( x112 & n734 ) ;
  assign n736 = ( ~n733 & n734 ) | ( ~n733 & n735 ) | ( n734 & n735 ) ;
  assign n737 = ( x111 & x112 ) | ( x111 & n733 ) | ( x112 & n733 ) ;
  assign n738 = ( x113 & ~x114 ) | ( x113 & n737 ) | ( ~x114 & n737 ) ;
  assign n739 = ( ~x113 & x114 ) | ( ~x113 & n738 ) | ( x114 & n738 ) ;
  assign n740 = ( ~n737 & n738 ) | ( ~n737 & n739 ) | ( n738 & n739 ) ;
  assign n741 = ( x113 & x114 ) | ( x113 & n737 ) | ( x114 & n737 ) ;
  assign n742 = ( x115 & ~x116 ) | ( x115 & n741 ) | ( ~x116 & n741 ) ;
  assign n743 = ( ~x115 & x116 ) | ( ~x115 & n742 ) | ( x116 & n742 ) ;
  assign n744 = ( ~n741 & n742 ) | ( ~n741 & n743 ) | ( n742 & n743 ) ;
  assign n745 = ( x115 & x116 ) | ( x115 & n741 ) | ( x116 & n741 ) ;
  assign n746 = ( x117 & ~x118 ) | ( x117 & n745 ) | ( ~x118 & n745 ) ;
  assign n747 = ( ~x117 & x118 ) | ( ~x117 & n746 ) | ( x118 & n746 ) ;
  assign n748 = ( ~n745 & n746 ) | ( ~n745 & n747 ) | ( n746 & n747 ) ;
  assign n749 = ( x117 & x118 ) | ( x117 & n745 ) | ( x118 & n745 ) ;
  assign n750 = ( x119 & ~x120 ) | ( x119 & n749 ) | ( ~x120 & n749 ) ;
  assign n751 = ( ~x119 & x120 ) | ( ~x119 & n750 ) | ( x120 & n750 ) ;
  assign n752 = ( ~n749 & n750 ) | ( ~n749 & n751 ) | ( n750 & n751 ) ;
  assign n753 = ( x119 & x120 ) | ( x119 & n749 ) | ( x120 & n749 ) ;
  assign n754 = ( x121 & ~x122 ) | ( x121 & n753 ) | ( ~x122 & n753 ) ;
  assign n755 = ( ~x121 & x122 ) | ( ~x121 & n754 ) | ( x122 & n754 ) ;
  assign n756 = ( ~n753 & n754 ) | ( ~n753 & n755 ) | ( n754 & n755 ) ;
  assign n757 = ( x121 & x122 ) | ( x121 & n753 ) | ( x122 & n753 ) ;
  assign n758 = ( x123 & ~x124 ) | ( x123 & n757 ) | ( ~x124 & n757 ) ;
  assign n759 = ( ~x123 & x124 ) | ( ~x123 & n758 ) | ( x124 & n758 ) ;
  assign n760 = ( ~n757 & n758 ) | ( ~n757 & n759 ) | ( n758 & n759 ) ;
  assign n761 = ( x123 & x124 ) | ( x123 & n757 ) | ( x124 & n757 ) ;
  assign n762 = ( x125 & ~x126 ) | ( x125 & n761 ) | ( ~x126 & n761 ) ;
  assign n763 = ( ~x125 & x126 ) | ( ~x125 & n762 ) | ( x126 & n762 ) ;
  assign n764 = ( ~n761 & n762 ) | ( ~n761 & n763 ) | ( n762 & n763 ) ;
  assign n765 = ( x125 & x126 ) | ( x125 & n761 ) | ( x126 & n761 ) ;
  assign n766 = ( x127 & ~x128 ) | ( x127 & n765 ) | ( ~x128 & n765 ) ;
  assign n767 = ( ~x127 & x128 ) | ( ~x127 & n766 ) | ( x128 & n766 ) ;
  assign n768 = ( ~n765 & n766 ) | ( ~n765 & n767 ) | ( n766 & n767 ) ;
  assign n769 = ( x127 & x128 ) | ( x127 & n765 ) | ( x128 & n765 ) ;
  assign n770 = ( x129 & ~x130 ) | ( x129 & n769 ) | ( ~x130 & n769 ) ;
  assign n771 = ( ~x129 & x130 ) | ( ~x129 & n770 ) | ( x130 & n770 ) ;
  assign n772 = ( ~n769 & n770 ) | ( ~n769 & n771 ) | ( n770 & n771 ) ;
  assign n773 = ( x129 & x130 ) | ( x129 & n769 ) | ( x130 & n769 ) ;
  assign n774 = ( x131 & ~x132 ) | ( x131 & n773 ) | ( ~x132 & n773 ) ;
  assign n775 = ( ~x131 & x132 ) | ( ~x131 & n774 ) | ( x132 & n774 ) ;
  assign n776 = ( ~n773 & n774 ) | ( ~n773 & n775 ) | ( n774 & n775 ) ;
  assign n777 = ( x131 & x132 ) | ( x131 & n773 ) | ( x132 & n773 ) ;
  assign n778 = ( x133 & ~x134 ) | ( x133 & n777 ) | ( ~x134 & n777 ) ;
  assign n779 = ( ~x133 & x134 ) | ( ~x133 & n778 ) | ( x134 & n778 ) ;
  assign n780 = ( ~n777 & n778 ) | ( ~n777 & n779 ) | ( n778 & n779 ) ;
  assign n781 = ( x133 & x134 ) | ( x133 & n777 ) | ( x134 & n777 ) ;
  assign n782 = ( x135 & ~x136 ) | ( x135 & n781 ) | ( ~x136 & n781 ) ;
  assign n783 = ( ~x135 & x136 ) | ( ~x135 & n782 ) | ( x136 & n782 ) ;
  assign n784 = ( ~n781 & n782 ) | ( ~n781 & n783 ) | ( n782 & n783 ) ;
  assign n785 = ( x135 & x136 ) | ( x135 & n781 ) | ( x136 & n781 ) ;
  assign n786 = ( x137 & ~x138 ) | ( x137 & n785 ) | ( ~x138 & n785 ) ;
  assign n787 = ( ~x137 & x138 ) | ( ~x137 & n786 ) | ( x138 & n786 ) ;
  assign n788 = ( ~n785 & n786 ) | ( ~n785 & n787 ) | ( n786 & n787 ) ;
  assign n789 = ( x137 & x138 ) | ( x137 & n785 ) | ( x138 & n785 ) ;
  assign n790 = ( x139 & ~x140 ) | ( x139 & n789 ) | ( ~x140 & n789 ) ;
  assign n791 = ( ~x139 & x140 ) | ( ~x139 & n790 ) | ( x140 & n790 ) ;
  assign n792 = ( ~n789 & n790 ) | ( ~n789 & n791 ) | ( n790 & n791 ) ;
  assign n793 = ( x139 & x140 ) | ( x139 & n789 ) | ( x140 & n789 ) ;
  assign n794 = ( x141 & ~x142 ) | ( x141 & n793 ) | ( ~x142 & n793 ) ;
  assign n795 = ( ~x141 & x142 ) | ( ~x141 & n794 ) | ( x142 & n794 ) ;
  assign n796 = ( ~n793 & n794 ) | ( ~n793 & n795 ) | ( n794 & n795 ) ;
  assign n797 = ( x141 & x142 ) | ( x141 & n793 ) | ( x142 & n793 ) ;
  assign n798 = ( x143 & ~x144 ) | ( x143 & n797 ) | ( ~x144 & n797 ) ;
  assign n799 = ( ~x143 & x144 ) | ( ~x143 & n798 ) | ( x144 & n798 ) ;
  assign n800 = ( ~n797 & n798 ) | ( ~n797 & n799 ) | ( n798 & n799 ) ;
  assign n801 = ( x143 & x144 ) | ( x143 & n797 ) | ( x144 & n797 ) ;
  assign n802 = ( x145 & ~x146 ) | ( x145 & n801 ) | ( ~x146 & n801 ) ;
  assign n803 = ( ~x145 & x146 ) | ( ~x145 & n802 ) | ( x146 & n802 ) ;
  assign n804 = ( ~n801 & n802 ) | ( ~n801 & n803 ) | ( n802 & n803 ) ;
  assign n805 = ( x145 & x146 ) | ( x145 & n801 ) | ( x146 & n801 ) ;
  assign n806 = ( x147 & ~x148 ) | ( x147 & n805 ) | ( ~x148 & n805 ) ;
  assign n807 = ( ~x147 & x148 ) | ( ~x147 & n806 ) | ( x148 & n806 ) ;
  assign n808 = ( ~n805 & n806 ) | ( ~n805 & n807 ) | ( n806 & n807 ) ;
  assign n809 = ( x147 & x148 ) | ( x147 & n805 ) | ( x148 & n805 ) ;
  assign n810 = ( x149 & ~x150 ) | ( x149 & n809 ) | ( ~x150 & n809 ) ;
  assign n811 = ( ~x149 & x150 ) | ( ~x149 & n810 ) | ( x150 & n810 ) ;
  assign n812 = ( ~n809 & n810 ) | ( ~n809 & n811 ) | ( n810 & n811 ) ;
  assign n813 = ( x149 & x150 ) | ( x149 & n809 ) | ( x150 & n809 ) ;
  assign n814 = ( x151 & ~x152 ) | ( x151 & n813 ) | ( ~x152 & n813 ) ;
  assign n815 = ( ~x151 & x152 ) | ( ~x151 & n814 ) | ( x152 & n814 ) ;
  assign n816 = ( ~n813 & n814 ) | ( ~n813 & n815 ) | ( n814 & n815 ) ;
  assign n817 = ( x151 & x152 ) | ( x151 & n813 ) | ( x152 & n813 ) ;
  assign n818 = ( x153 & ~x154 ) | ( x153 & n817 ) | ( ~x154 & n817 ) ;
  assign n819 = ( ~x153 & x154 ) | ( ~x153 & n818 ) | ( x154 & n818 ) ;
  assign n820 = ( ~n817 & n818 ) | ( ~n817 & n819 ) | ( n818 & n819 ) ;
  assign n821 = ( x153 & x154 ) | ( x153 & n817 ) | ( x154 & n817 ) ;
  assign n822 = ( x155 & ~x156 ) | ( x155 & n821 ) | ( ~x156 & n821 ) ;
  assign n823 = ( ~x155 & x156 ) | ( ~x155 & n822 ) | ( x156 & n822 ) ;
  assign n824 = ( ~n821 & n822 ) | ( ~n821 & n823 ) | ( n822 & n823 ) ;
  assign n825 = ( x155 & x156 ) | ( x155 & n821 ) | ( x156 & n821 ) ;
  assign n826 = ( x157 & ~x158 ) | ( x157 & n825 ) | ( ~x158 & n825 ) ;
  assign n827 = ( ~x157 & x158 ) | ( ~x157 & n826 ) | ( x158 & n826 ) ;
  assign n828 = ( ~n825 & n826 ) | ( ~n825 & n827 ) | ( n826 & n827 ) ;
  assign n829 = ( x157 & x158 ) | ( x157 & n825 ) | ( x158 & n825 ) ;
  assign n830 = ( x159 & ~x160 ) | ( x159 & n829 ) | ( ~x160 & n829 ) ;
  assign n831 = ( ~x159 & x160 ) | ( ~x159 & n830 ) | ( x160 & n830 ) ;
  assign n832 = ( ~n829 & n830 ) | ( ~n829 & n831 ) | ( n830 & n831 ) ;
  assign n833 = ( x159 & x160 ) | ( x159 & n829 ) | ( x160 & n829 ) ;
  assign n834 = ( x161 & ~x162 ) | ( x161 & n833 ) | ( ~x162 & n833 ) ;
  assign n835 = ( ~x161 & x162 ) | ( ~x161 & n834 ) | ( x162 & n834 ) ;
  assign n836 = ( ~n833 & n834 ) | ( ~n833 & n835 ) | ( n834 & n835 ) ;
  assign n837 = ( x161 & x162 ) | ( x161 & n833 ) | ( x162 & n833 ) ;
  assign n838 = ( x163 & ~x164 ) | ( x163 & n837 ) | ( ~x164 & n837 ) ;
  assign n839 = ( ~x163 & x164 ) | ( ~x163 & n838 ) | ( x164 & n838 ) ;
  assign n840 = ( ~n837 & n838 ) | ( ~n837 & n839 ) | ( n838 & n839 ) ;
  assign n841 = ( x163 & x164 ) | ( x163 & n837 ) | ( x164 & n837 ) ;
  assign n842 = ( x165 & ~x166 ) | ( x165 & n841 ) | ( ~x166 & n841 ) ;
  assign n843 = ( ~x165 & x166 ) | ( ~x165 & n842 ) | ( x166 & n842 ) ;
  assign n844 = ( ~n841 & n842 ) | ( ~n841 & n843 ) | ( n842 & n843 ) ;
  assign n845 = ( x165 & x166 ) | ( x165 & n841 ) | ( x166 & n841 ) ;
  assign n846 = ( x167 & ~x168 ) | ( x167 & n845 ) | ( ~x168 & n845 ) ;
  assign n847 = ( ~x167 & x168 ) | ( ~x167 & n846 ) | ( x168 & n846 ) ;
  assign n848 = ( ~n845 & n846 ) | ( ~n845 & n847 ) | ( n846 & n847 ) ;
  assign n849 = ( x167 & x168 ) | ( x167 & n845 ) | ( x168 & n845 ) ;
  assign n850 = ( x169 & ~x170 ) | ( x169 & n849 ) | ( ~x170 & n849 ) ;
  assign n851 = ( ~x169 & x170 ) | ( ~x169 & n850 ) | ( x170 & n850 ) ;
  assign n852 = ( ~n849 & n850 ) | ( ~n849 & n851 ) | ( n850 & n851 ) ;
  assign n853 = ( x169 & x170 ) | ( x169 & n849 ) | ( x170 & n849 ) ;
  assign n854 = ( x171 & ~x172 ) | ( x171 & n853 ) | ( ~x172 & n853 ) ;
  assign n855 = ( ~x171 & x172 ) | ( ~x171 & n854 ) | ( x172 & n854 ) ;
  assign n856 = ( ~n853 & n854 ) | ( ~n853 & n855 ) | ( n854 & n855 ) ;
  assign n857 = ( x171 & x172 ) | ( x171 & n853 ) | ( x172 & n853 ) ;
  assign n858 = ( x173 & ~x174 ) | ( x173 & n857 ) | ( ~x174 & n857 ) ;
  assign n859 = ( ~x173 & x174 ) | ( ~x173 & n858 ) | ( x174 & n858 ) ;
  assign n860 = ( ~n857 & n858 ) | ( ~n857 & n859 ) | ( n858 & n859 ) ;
  assign n861 = ( x173 & x174 ) | ( x173 & n857 ) | ( x174 & n857 ) ;
  assign n862 = ( x175 & ~x176 ) | ( x175 & n861 ) | ( ~x176 & n861 ) ;
  assign n863 = ( ~x175 & x176 ) | ( ~x175 & n862 ) | ( x176 & n862 ) ;
  assign n864 = ( ~n861 & n862 ) | ( ~n861 & n863 ) | ( n862 & n863 ) ;
  assign n865 = ( x175 & x176 ) | ( x175 & n861 ) | ( x176 & n861 ) ;
  assign n866 = ( x177 & ~x178 ) | ( x177 & n865 ) | ( ~x178 & n865 ) ;
  assign n867 = ( ~x177 & x178 ) | ( ~x177 & n866 ) | ( x178 & n866 ) ;
  assign n868 = ( ~n865 & n866 ) | ( ~n865 & n867 ) | ( n866 & n867 ) ;
  assign n869 = ( x177 & x178 ) | ( x177 & n865 ) | ( x178 & n865 ) ;
  assign n870 = ( x179 & ~x180 ) | ( x179 & n869 ) | ( ~x180 & n869 ) ;
  assign n871 = ( ~x179 & x180 ) | ( ~x179 & n870 ) | ( x180 & n870 ) ;
  assign n872 = ( ~n869 & n870 ) | ( ~n869 & n871 ) | ( n870 & n871 ) ;
  assign n873 = ( x179 & x180 ) | ( x179 & n869 ) | ( x180 & n869 ) ;
  assign n874 = ( x181 & ~x182 ) | ( x181 & n873 ) | ( ~x182 & n873 ) ;
  assign n875 = ( ~x181 & x182 ) | ( ~x181 & n874 ) | ( x182 & n874 ) ;
  assign n876 = ( ~n873 & n874 ) | ( ~n873 & n875 ) | ( n874 & n875 ) ;
  assign n877 = ( x181 & x182 ) | ( x181 & n873 ) | ( x182 & n873 ) ;
  assign n878 = ( x183 & ~x184 ) | ( x183 & n877 ) | ( ~x184 & n877 ) ;
  assign n879 = ( ~x183 & x184 ) | ( ~x183 & n878 ) | ( x184 & n878 ) ;
  assign n880 = ( ~n877 & n878 ) | ( ~n877 & n879 ) | ( n878 & n879 ) ;
  assign n881 = ( x183 & x184 ) | ( x183 & n877 ) | ( x184 & n877 ) ;
  assign n882 = ( x185 & ~x186 ) | ( x185 & n881 ) | ( ~x186 & n881 ) ;
  assign n883 = ( ~x185 & x186 ) | ( ~x185 & n882 ) | ( x186 & n882 ) ;
  assign n884 = ( ~n881 & n882 ) | ( ~n881 & n883 ) | ( n882 & n883 ) ;
  assign n885 = ( x185 & x186 ) | ( x185 & n881 ) | ( x186 & n881 ) ;
  assign n886 = ( x187 & ~x188 ) | ( x187 & n885 ) | ( ~x188 & n885 ) ;
  assign n887 = ( ~x187 & x188 ) | ( ~x187 & n886 ) | ( x188 & n886 ) ;
  assign n888 = ( ~n885 & n886 ) | ( ~n885 & n887 ) | ( n886 & n887 ) ;
  assign n889 = ( x187 & x188 ) | ( x187 & n885 ) | ( x188 & n885 ) ;
  assign n890 = ( x189 & ~x190 ) | ( x189 & n889 ) | ( ~x190 & n889 ) ;
  assign n891 = ( ~x189 & x190 ) | ( ~x189 & n890 ) | ( x190 & n890 ) ;
  assign n892 = ( ~n889 & n890 ) | ( ~n889 & n891 ) | ( n890 & n891 ) ;
  assign n893 = ( x189 & x190 ) | ( x189 & n889 ) | ( x190 & n889 ) ;
  assign n894 = ( x191 & ~x192 ) | ( x191 & n893 ) | ( ~x192 & n893 ) ;
  assign n895 = ( ~x191 & x192 ) | ( ~x191 & n894 ) | ( x192 & n894 ) ;
  assign n896 = ( ~n893 & n894 ) | ( ~n893 & n895 ) | ( n894 & n895 ) ;
  assign n897 = ( x191 & x192 ) | ( x191 & n893 ) | ( x192 & n893 ) ;
  assign n898 = ( x193 & ~x194 ) | ( x193 & n897 ) | ( ~x194 & n897 ) ;
  assign n899 = ( ~x193 & x194 ) | ( ~x193 & n898 ) | ( x194 & n898 ) ;
  assign n900 = ( ~n897 & n898 ) | ( ~n897 & n899 ) | ( n898 & n899 ) ;
  assign n901 = ( x193 & x194 ) | ( x193 & n897 ) | ( x194 & n897 ) ;
  assign n902 = ( x195 & ~x196 ) | ( x195 & n901 ) | ( ~x196 & n901 ) ;
  assign n903 = ( ~x195 & x196 ) | ( ~x195 & n902 ) | ( x196 & n902 ) ;
  assign n904 = ( ~n901 & n902 ) | ( ~n901 & n903 ) | ( n902 & n903 ) ;
  assign n905 = ( x195 & x196 ) | ( x195 & n901 ) | ( x196 & n901 ) ;
  assign n906 = ( x197 & ~x198 ) | ( x197 & n905 ) | ( ~x198 & n905 ) ;
  assign n907 = ( ~x197 & x198 ) | ( ~x197 & n906 ) | ( x198 & n906 ) ;
  assign n908 = ( ~n905 & n906 ) | ( ~n905 & n907 ) | ( n906 & n907 ) ;
  assign n909 = ( x197 & x198 ) | ( x197 & n905 ) | ( x198 & n905 ) ;
  assign n910 = ( x199 & ~x200 ) | ( x199 & n909 ) | ( ~x200 & n909 ) ;
  assign n911 = ( ~x199 & x200 ) | ( ~x199 & n910 ) | ( x200 & n910 ) ;
  assign n912 = ( ~n909 & n910 ) | ( ~n909 & n911 ) | ( n910 & n911 ) ;
  assign n913 = ( x199 & x200 ) | ( x199 & n909 ) | ( x200 & n909 ) ;
  assign n914 = ( x201 & ~x202 ) | ( x201 & n913 ) | ( ~x202 & n913 ) ;
  assign n915 = ( ~x201 & x202 ) | ( ~x201 & n914 ) | ( x202 & n914 ) ;
  assign n916 = ( ~n913 & n914 ) | ( ~n913 & n915 ) | ( n914 & n915 ) ;
  assign n917 = ( x201 & x202 ) | ( x201 & n913 ) | ( x202 & n913 ) ;
  assign n918 = ( x203 & ~x204 ) | ( x203 & n917 ) | ( ~x204 & n917 ) ;
  assign n919 = ( ~x203 & x204 ) | ( ~x203 & n918 ) | ( x204 & n918 ) ;
  assign n920 = ( ~n917 & n918 ) | ( ~n917 & n919 ) | ( n918 & n919 ) ;
  assign n921 = ( x203 & x204 ) | ( x203 & n917 ) | ( x204 & n917 ) ;
  assign n922 = ( x205 & ~x206 ) | ( x205 & n921 ) | ( ~x206 & n921 ) ;
  assign n923 = ( ~x205 & x206 ) | ( ~x205 & n922 ) | ( x206 & n922 ) ;
  assign n924 = ( ~n921 & n922 ) | ( ~n921 & n923 ) | ( n922 & n923 ) ;
  assign n925 = ( x205 & x206 ) | ( x205 & n921 ) | ( x206 & n921 ) ;
  assign n926 = ( x207 & ~x208 ) | ( x207 & n925 ) | ( ~x208 & n925 ) ;
  assign n927 = ( ~x207 & x208 ) | ( ~x207 & n926 ) | ( x208 & n926 ) ;
  assign n928 = ( ~n925 & n926 ) | ( ~n925 & n927 ) | ( n926 & n927 ) ;
  assign n929 = ( x207 & x208 ) | ( x207 & n925 ) | ( x208 & n925 ) ;
  assign n930 = ( x209 & ~x210 ) | ( x209 & n929 ) | ( ~x210 & n929 ) ;
  assign n931 = ( ~x209 & x210 ) | ( ~x209 & n930 ) | ( x210 & n930 ) ;
  assign n932 = ( ~n929 & n930 ) | ( ~n929 & n931 ) | ( n930 & n931 ) ;
  assign n933 = ( x209 & x210 ) | ( x209 & n929 ) | ( x210 & n929 ) ;
  assign n934 = ( x211 & ~x212 ) | ( x211 & n933 ) | ( ~x212 & n933 ) ;
  assign n935 = ( ~x211 & x212 ) | ( ~x211 & n934 ) | ( x212 & n934 ) ;
  assign n936 = ( ~n933 & n934 ) | ( ~n933 & n935 ) | ( n934 & n935 ) ;
  assign n937 = ( x211 & x212 ) | ( x211 & n933 ) | ( x212 & n933 ) ;
  assign n938 = ( x213 & ~x214 ) | ( x213 & n937 ) | ( ~x214 & n937 ) ;
  assign n939 = ( ~x213 & x214 ) | ( ~x213 & n938 ) | ( x214 & n938 ) ;
  assign n940 = ( ~n937 & n938 ) | ( ~n937 & n939 ) | ( n938 & n939 ) ;
  assign n941 = ( x213 & x214 ) | ( x213 & n937 ) | ( x214 & n937 ) ;
  assign n942 = ( x215 & ~x216 ) | ( x215 & n941 ) | ( ~x216 & n941 ) ;
  assign n943 = ( ~x215 & x216 ) | ( ~x215 & n942 ) | ( x216 & n942 ) ;
  assign n944 = ( ~n941 & n942 ) | ( ~n941 & n943 ) | ( n942 & n943 ) ;
  assign n945 = ( x215 & x216 ) | ( x215 & n941 ) | ( x216 & n941 ) ;
  assign n946 = ( x217 & ~x218 ) | ( x217 & n945 ) | ( ~x218 & n945 ) ;
  assign n947 = ( ~x217 & x218 ) | ( ~x217 & n946 ) | ( x218 & n946 ) ;
  assign n948 = ( ~n945 & n946 ) | ( ~n945 & n947 ) | ( n946 & n947 ) ;
  assign n949 = ( x217 & x218 ) | ( x217 & n945 ) | ( x218 & n945 ) ;
  assign n950 = ( x219 & ~x220 ) | ( x219 & n949 ) | ( ~x220 & n949 ) ;
  assign n951 = ( ~x219 & x220 ) | ( ~x219 & n950 ) | ( x220 & n950 ) ;
  assign n952 = ( ~n949 & n950 ) | ( ~n949 & n951 ) | ( n950 & n951 ) ;
  assign n953 = ( x219 & x220 ) | ( x219 & n949 ) | ( x220 & n949 ) ;
  assign n954 = ( x221 & ~x222 ) | ( x221 & n953 ) | ( ~x222 & n953 ) ;
  assign n955 = ( ~x221 & x222 ) | ( ~x221 & n954 ) | ( x222 & n954 ) ;
  assign n956 = ( ~n953 & n954 ) | ( ~n953 & n955 ) | ( n954 & n955 ) ;
  assign n957 = ( x221 & x222 ) | ( x221 & n953 ) | ( x222 & n953 ) ;
  assign n958 = ( x223 & ~x224 ) | ( x223 & n957 ) | ( ~x224 & n957 ) ;
  assign n959 = ( ~x223 & x224 ) | ( ~x223 & n958 ) | ( x224 & n958 ) ;
  assign n960 = ( ~n957 & n958 ) | ( ~n957 & n959 ) | ( n958 & n959 ) ;
  assign n961 = ( x223 & x224 ) | ( x223 & n957 ) | ( x224 & n957 ) ;
  assign n962 = ( x225 & ~x226 ) | ( x225 & n961 ) | ( ~x226 & n961 ) ;
  assign n963 = ( ~x225 & x226 ) | ( ~x225 & n962 ) | ( x226 & n962 ) ;
  assign n964 = ( ~n961 & n962 ) | ( ~n961 & n963 ) | ( n962 & n963 ) ;
  assign n965 = ( x225 & x226 ) | ( x225 & n961 ) | ( x226 & n961 ) ;
  assign n966 = ( x227 & ~x228 ) | ( x227 & n965 ) | ( ~x228 & n965 ) ;
  assign n967 = ( ~x227 & x228 ) | ( ~x227 & n966 ) | ( x228 & n966 ) ;
  assign n968 = ( ~n965 & n966 ) | ( ~n965 & n967 ) | ( n966 & n967 ) ;
  assign n969 = ( x227 & x228 ) | ( x227 & n965 ) | ( x228 & n965 ) ;
  assign n970 = ( x229 & ~x230 ) | ( x229 & n969 ) | ( ~x230 & n969 ) ;
  assign n971 = ( ~x229 & x230 ) | ( ~x229 & n970 ) | ( x230 & n970 ) ;
  assign n972 = ( ~n969 & n970 ) | ( ~n969 & n971 ) | ( n970 & n971 ) ;
  assign n973 = ( x229 & x230 ) | ( x229 & n969 ) | ( x230 & n969 ) ;
  assign n974 = ( x231 & ~x232 ) | ( x231 & n973 ) | ( ~x232 & n973 ) ;
  assign n975 = ( ~x231 & x232 ) | ( ~x231 & n974 ) | ( x232 & n974 ) ;
  assign n976 = ( ~n973 & n974 ) | ( ~n973 & n975 ) | ( n974 & n975 ) ;
  assign n977 = ( x231 & x232 ) | ( x231 & n973 ) | ( x232 & n973 ) ;
  assign n978 = ( x233 & ~x234 ) | ( x233 & n977 ) | ( ~x234 & n977 ) ;
  assign n979 = ( ~x233 & x234 ) | ( ~x233 & n978 ) | ( x234 & n978 ) ;
  assign n980 = ( ~n977 & n978 ) | ( ~n977 & n979 ) | ( n978 & n979 ) ;
  assign n981 = ( x233 & x234 ) | ( x233 & n977 ) | ( x234 & n977 ) ;
  assign n982 = ( x235 & ~x236 ) | ( x235 & n981 ) | ( ~x236 & n981 ) ;
  assign n983 = ( ~x235 & x236 ) | ( ~x235 & n982 ) | ( x236 & n982 ) ;
  assign n984 = ( ~n981 & n982 ) | ( ~n981 & n983 ) | ( n982 & n983 ) ;
  assign n985 = ( x235 & x236 ) | ( x235 & n981 ) | ( x236 & n981 ) ;
  assign n986 = ( x237 & ~x238 ) | ( x237 & n985 ) | ( ~x238 & n985 ) ;
  assign n987 = ( ~x237 & x238 ) | ( ~x237 & n986 ) | ( x238 & n986 ) ;
  assign n988 = ( ~n985 & n986 ) | ( ~n985 & n987 ) | ( n986 & n987 ) ;
  assign n989 = ( x237 & x238 ) | ( x237 & n985 ) | ( x238 & n985 ) ;
  assign n990 = ( x239 & ~x240 ) | ( x239 & n989 ) | ( ~x240 & n989 ) ;
  assign n991 = ( ~x239 & x240 ) | ( ~x239 & n990 ) | ( x240 & n990 ) ;
  assign n992 = ( ~n989 & n990 ) | ( ~n989 & n991 ) | ( n990 & n991 ) ;
  assign n993 = ( x239 & x240 ) | ( x239 & n989 ) | ( x240 & n989 ) ;
  assign n994 = ( x241 & ~x242 ) | ( x241 & n993 ) | ( ~x242 & n993 ) ;
  assign n995 = ( ~x241 & x242 ) | ( ~x241 & n994 ) | ( x242 & n994 ) ;
  assign n996 = ( ~n993 & n994 ) | ( ~n993 & n995 ) | ( n994 & n995 ) ;
  assign n997 = ( x241 & x242 ) | ( x241 & n993 ) | ( x242 & n993 ) ;
  assign n998 = ( x243 & ~x244 ) | ( x243 & n997 ) | ( ~x244 & n997 ) ;
  assign n999 = ( ~x243 & x244 ) | ( ~x243 & n998 ) | ( x244 & n998 ) ;
  assign n1000 = ( ~n997 & n998 ) | ( ~n997 & n999 ) | ( n998 & n999 ) ;
  assign n1001 = ( x243 & x244 ) | ( x243 & n997 ) | ( x244 & n997 ) ;
  assign n1002 = ( x245 & ~x246 ) | ( x245 & n1001 ) | ( ~x246 & n1001 ) ;
  assign n1003 = ( ~x245 & x246 ) | ( ~x245 & n1002 ) | ( x246 & n1002 ) ;
  assign n1004 = ( ~n1001 & n1002 ) | ( ~n1001 & n1003 ) | ( n1002 & n1003 ) ;
  assign n1005 = ( x245 & x246 ) | ( x245 & n1001 ) | ( x246 & n1001 ) ;
  assign n1006 = ( x247 & ~x248 ) | ( x247 & n1005 ) | ( ~x248 & n1005 ) ;
  assign n1007 = ( ~x247 & x248 ) | ( ~x247 & n1006 ) | ( x248 & n1006 ) ;
  assign n1008 = ( ~n1005 & n1006 ) | ( ~n1005 & n1007 ) | ( n1006 & n1007 ) ;
  assign n1009 = ( x247 & x248 ) | ( x247 & n1005 ) | ( x248 & n1005 ) ;
  assign n1010 = ( x249 & ~x250 ) | ( x249 & n1009 ) | ( ~x250 & n1009 ) ;
  assign n1011 = ( ~x249 & x250 ) | ( ~x249 & n1010 ) | ( x250 & n1010 ) ;
  assign n1012 = ( ~n1009 & n1010 ) | ( ~n1009 & n1011 ) | ( n1010 & n1011 ) ;
  assign n1013 = ( x249 & x250 ) | ( x249 & n1009 ) | ( x250 & n1009 ) ;
  assign n1014 = ( x251 & ~x252 ) | ( x251 & n1013 ) | ( ~x252 & n1013 ) ;
  assign n1015 = ( ~x251 & x252 ) | ( ~x251 & n1014 ) | ( x252 & n1014 ) ;
  assign n1016 = ( ~n1013 & n1014 ) | ( ~n1013 & n1015 ) | ( n1014 & n1015 ) ;
  assign n1017 = ( x251 & x252 ) | ( x251 & n1013 ) | ( x252 & n1013 ) ;
  assign n1018 = ( x253 & ~x254 ) | ( x253 & n1017 ) | ( ~x254 & n1017 ) ;
  assign n1019 = ( ~x253 & x254 ) | ( ~x253 & n1018 ) | ( x254 & n1018 ) ;
  assign n1020 = ( ~n1017 & n1018 ) | ( ~n1017 & n1019 ) | ( n1018 & n1019 ) ;
  assign n1021 = ( x253 & x254 ) | ( x253 & n1017 ) | ( x254 & n1017 ) ;
  assign n1022 = ( x255 & ~x256 ) | ( x255 & n1021 ) | ( ~x256 & n1021 ) ;
  assign n1023 = ( ~x255 & x256 ) | ( ~x255 & n1022 ) | ( x256 & n1022 ) ;
  assign n1024 = ( ~n1021 & n1022 ) | ( ~n1021 & n1023 ) | ( n1022 & n1023 ) ;
  assign n1025 = ( x255 & x256 ) | ( x255 & n1021 ) | ( x256 & n1021 ) ;
  assign n1026 = ( x257 & ~x258 ) | ( x257 & n1025 ) | ( ~x258 & n1025 ) ;
  assign n1027 = ( ~x257 & x258 ) | ( ~x257 & n1026 ) | ( x258 & n1026 ) ;
  assign n1028 = ( ~n1025 & n1026 ) | ( ~n1025 & n1027 ) | ( n1026 & n1027 ) ;
  assign n1029 = ( x257 & x258 ) | ( x257 & n1025 ) | ( x258 & n1025 ) ;
  assign n1030 = ( x259 & ~x260 ) | ( x259 & n1029 ) | ( ~x260 & n1029 ) ;
  assign n1031 = ( ~x259 & x260 ) | ( ~x259 & n1030 ) | ( x260 & n1030 ) ;
  assign n1032 = ( ~n1029 & n1030 ) | ( ~n1029 & n1031 ) | ( n1030 & n1031 ) ;
  assign n1033 = ( x259 & x260 ) | ( x259 & n1029 ) | ( x260 & n1029 ) ;
  assign n1034 = ( x261 & ~x262 ) | ( x261 & n1033 ) | ( ~x262 & n1033 ) ;
  assign n1035 = ( ~x261 & x262 ) | ( ~x261 & n1034 ) | ( x262 & n1034 ) ;
  assign n1036 = ( ~n1033 & n1034 ) | ( ~n1033 & n1035 ) | ( n1034 & n1035 ) ;
  assign n1037 = ( x261 & x262 ) | ( x261 & n1033 ) | ( x262 & n1033 ) ;
  assign n1038 = ( x263 & ~x264 ) | ( x263 & n1037 ) | ( ~x264 & n1037 ) ;
  assign n1039 = ( ~x263 & x264 ) | ( ~x263 & n1038 ) | ( x264 & n1038 ) ;
  assign n1040 = ( ~n1037 & n1038 ) | ( ~n1037 & n1039 ) | ( n1038 & n1039 ) ;
  assign n1041 = ( x263 & x264 ) | ( x263 & n1037 ) | ( x264 & n1037 ) ;
  assign n1042 = ( x265 & ~x266 ) | ( x265 & n1041 ) | ( ~x266 & n1041 ) ;
  assign n1043 = ( ~x265 & x266 ) | ( ~x265 & n1042 ) | ( x266 & n1042 ) ;
  assign n1044 = ( ~n1041 & n1042 ) | ( ~n1041 & n1043 ) | ( n1042 & n1043 ) ;
  assign n1045 = ( x265 & x266 ) | ( x265 & n1041 ) | ( x266 & n1041 ) ;
  assign n1046 = ( x267 & ~x268 ) | ( x267 & n1045 ) | ( ~x268 & n1045 ) ;
  assign n1047 = ( ~x267 & x268 ) | ( ~x267 & n1046 ) | ( x268 & n1046 ) ;
  assign n1048 = ( ~n1045 & n1046 ) | ( ~n1045 & n1047 ) | ( n1046 & n1047 ) ;
  assign n1049 = ( x267 & x268 ) | ( x267 & n1045 ) | ( x268 & n1045 ) ;
  assign n1050 = ( x269 & ~x270 ) | ( x269 & n1049 ) | ( ~x270 & n1049 ) ;
  assign n1051 = ( ~x269 & x270 ) | ( ~x269 & n1050 ) | ( x270 & n1050 ) ;
  assign n1052 = ( ~n1049 & n1050 ) | ( ~n1049 & n1051 ) | ( n1050 & n1051 ) ;
  assign n1053 = ( x269 & x270 ) | ( x269 & n1049 ) | ( x270 & n1049 ) ;
  assign n1054 = ( x271 & ~x272 ) | ( x271 & n1053 ) | ( ~x272 & n1053 ) ;
  assign n1055 = ( ~x271 & x272 ) | ( ~x271 & n1054 ) | ( x272 & n1054 ) ;
  assign n1056 = ( ~n1053 & n1054 ) | ( ~n1053 & n1055 ) | ( n1054 & n1055 ) ;
  assign n1057 = ( x271 & x272 ) | ( x271 & n1053 ) | ( x272 & n1053 ) ;
  assign n1058 = ( x273 & ~x274 ) | ( x273 & n1057 ) | ( ~x274 & n1057 ) ;
  assign n1059 = ( ~x273 & x274 ) | ( ~x273 & n1058 ) | ( x274 & n1058 ) ;
  assign n1060 = ( ~n1057 & n1058 ) | ( ~n1057 & n1059 ) | ( n1058 & n1059 ) ;
  assign n1061 = ( x273 & x274 ) | ( x273 & n1057 ) | ( x274 & n1057 ) ;
  assign n1062 = ( x275 & ~x276 ) | ( x275 & n1061 ) | ( ~x276 & n1061 ) ;
  assign n1063 = ( ~x275 & x276 ) | ( ~x275 & n1062 ) | ( x276 & n1062 ) ;
  assign n1064 = ( ~n1061 & n1062 ) | ( ~n1061 & n1063 ) | ( n1062 & n1063 ) ;
  assign n1065 = ( x275 & x276 ) | ( x275 & n1061 ) | ( x276 & n1061 ) ;
  assign n1066 = ( x277 & ~x278 ) | ( x277 & n1065 ) | ( ~x278 & n1065 ) ;
  assign n1067 = ( ~x277 & x278 ) | ( ~x277 & n1066 ) | ( x278 & n1066 ) ;
  assign n1068 = ( ~n1065 & n1066 ) | ( ~n1065 & n1067 ) | ( n1066 & n1067 ) ;
  assign n1069 = ( x277 & x278 ) | ( x277 & n1065 ) | ( x278 & n1065 ) ;
  assign n1070 = ( x279 & ~x280 ) | ( x279 & n1069 ) | ( ~x280 & n1069 ) ;
  assign n1071 = ( ~x279 & x280 ) | ( ~x279 & n1070 ) | ( x280 & n1070 ) ;
  assign n1072 = ( ~n1069 & n1070 ) | ( ~n1069 & n1071 ) | ( n1070 & n1071 ) ;
  assign n1073 = ( x279 & x280 ) | ( x279 & n1069 ) | ( x280 & n1069 ) ;
  assign n1074 = ( x281 & ~x282 ) | ( x281 & n1073 ) | ( ~x282 & n1073 ) ;
  assign n1075 = ( ~x281 & x282 ) | ( ~x281 & n1074 ) | ( x282 & n1074 ) ;
  assign n1076 = ( ~n1073 & n1074 ) | ( ~n1073 & n1075 ) | ( n1074 & n1075 ) ;
  assign n1077 = ( x281 & x282 ) | ( x281 & n1073 ) | ( x282 & n1073 ) ;
  assign n1078 = ( x283 & ~x284 ) | ( x283 & n1077 ) | ( ~x284 & n1077 ) ;
  assign n1079 = ( ~x283 & x284 ) | ( ~x283 & n1078 ) | ( x284 & n1078 ) ;
  assign n1080 = ( ~n1077 & n1078 ) | ( ~n1077 & n1079 ) | ( n1078 & n1079 ) ;
  assign n1081 = ( x283 & x284 ) | ( x283 & n1077 ) | ( x284 & n1077 ) ;
  assign n1082 = ( x285 & ~x286 ) | ( x285 & n1081 ) | ( ~x286 & n1081 ) ;
  assign n1083 = ( ~x285 & x286 ) | ( ~x285 & n1082 ) | ( x286 & n1082 ) ;
  assign n1084 = ( ~n1081 & n1082 ) | ( ~n1081 & n1083 ) | ( n1082 & n1083 ) ;
  assign n1085 = ( x285 & x286 ) | ( x285 & n1081 ) | ( x286 & n1081 ) ;
  assign n1086 = ( x287 & ~x288 ) | ( x287 & n1085 ) | ( ~x288 & n1085 ) ;
  assign n1087 = ( ~x287 & x288 ) | ( ~x287 & n1086 ) | ( x288 & n1086 ) ;
  assign n1088 = ( ~n1085 & n1086 ) | ( ~n1085 & n1087 ) | ( n1086 & n1087 ) ;
  assign n1089 = ( x287 & x288 ) | ( x287 & n1085 ) | ( x288 & n1085 ) ;
  assign n1090 = ( x289 & ~x290 ) | ( x289 & n1089 ) | ( ~x290 & n1089 ) ;
  assign n1091 = ( ~x289 & x290 ) | ( ~x289 & n1090 ) | ( x290 & n1090 ) ;
  assign n1092 = ( ~n1089 & n1090 ) | ( ~n1089 & n1091 ) | ( n1090 & n1091 ) ;
  assign n1093 = ( x289 & x290 ) | ( x289 & n1089 ) | ( x290 & n1089 ) ;
  assign n1094 = ( x291 & ~x292 ) | ( x291 & n1093 ) | ( ~x292 & n1093 ) ;
  assign n1095 = ( ~x291 & x292 ) | ( ~x291 & n1094 ) | ( x292 & n1094 ) ;
  assign n1096 = ( ~n1093 & n1094 ) | ( ~n1093 & n1095 ) | ( n1094 & n1095 ) ;
  assign n1097 = ( x291 & x292 ) | ( x291 & n1093 ) | ( x292 & n1093 ) ;
  assign n1098 = ( x293 & ~x294 ) | ( x293 & n1097 ) | ( ~x294 & n1097 ) ;
  assign n1099 = ( ~x293 & x294 ) | ( ~x293 & n1098 ) | ( x294 & n1098 ) ;
  assign n1100 = ( ~n1097 & n1098 ) | ( ~n1097 & n1099 ) | ( n1098 & n1099 ) ;
  assign n1101 = ( x293 & x294 ) | ( x293 & n1097 ) | ( x294 & n1097 ) ;
  assign n1102 = ( x295 & ~x296 ) | ( x295 & n1101 ) | ( ~x296 & n1101 ) ;
  assign n1103 = ( ~x295 & x296 ) | ( ~x295 & n1102 ) | ( x296 & n1102 ) ;
  assign n1104 = ( ~n1101 & n1102 ) | ( ~n1101 & n1103 ) | ( n1102 & n1103 ) ;
  assign n1105 = ( x295 & x296 ) | ( x295 & n1101 ) | ( x296 & n1101 ) ;
  assign n1106 = ( x297 & ~x298 ) | ( x297 & n1105 ) | ( ~x298 & n1105 ) ;
  assign n1107 = ( ~x297 & x298 ) | ( ~x297 & n1106 ) | ( x298 & n1106 ) ;
  assign n1108 = ( ~n1105 & n1106 ) | ( ~n1105 & n1107 ) | ( n1106 & n1107 ) ;
  assign n1109 = ( x297 & x298 ) | ( x297 & n1105 ) | ( x298 & n1105 ) ;
  assign n1110 = ( x299 & ~x300 ) | ( x299 & n1109 ) | ( ~x300 & n1109 ) ;
  assign n1111 = ( ~x299 & x300 ) | ( ~x299 & n1110 ) | ( x300 & n1110 ) ;
  assign n1112 = ( ~n1109 & n1110 ) | ( ~n1109 & n1111 ) | ( n1110 & n1111 ) ;
  assign n1113 = ( x299 & x300 ) | ( x299 & n1109 ) | ( x300 & n1109 ) ;
  assign n1114 = ( x301 & ~x302 ) | ( x301 & n1113 ) | ( ~x302 & n1113 ) ;
  assign n1115 = ( ~x301 & x302 ) | ( ~x301 & n1114 ) | ( x302 & n1114 ) ;
  assign n1116 = ( ~n1113 & n1114 ) | ( ~n1113 & n1115 ) | ( n1114 & n1115 ) ;
  assign n1117 = ( x301 & x302 ) | ( x301 & n1113 ) | ( x302 & n1113 ) ;
  assign n1118 = ( x303 & ~x304 ) | ( x303 & n1117 ) | ( ~x304 & n1117 ) ;
  assign n1119 = ( ~x303 & x304 ) | ( ~x303 & n1118 ) | ( x304 & n1118 ) ;
  assign n1120 = ( ~n1117 & n1118 ) | ( ~n1117 & n1119 ) | ( n1118 & n1119 ) ;
  assign n1121 = ( x303 & x304 ) | ( x303 & n1117 ) | ( x304 & n1117 ) ;
  assign n1122 = ( x305 & ~x306 ) | ( x305 & n1121 ) | ( ~x306 & n1121 ) ;
  assign n1123 = ( ~x305 & x306 ) | ( ~x305 & n1122 ) | ( x306 & n1122 ) ;
  assign n1124 = ( ~n1121 & n1122 ) | ( ~n1121 & n1123 ) | ( n1122 & n1123 ) ;
  assign n1125 = ( x305 & x306 ) | ( x305 & n1121 ) | ( x306 & n1121 ) ;
  assign n1126 = ( x307 & ~x308 ) | ( x307 & n1125 ) | ( ~x308 & n1125 ) ;
  assign n1127 = ( ~x307 & x308 ) | ( ~x307 & n1126 ) | ( x308 & n1126 ) ;
  assign n1128 = ( ~n1125 & n1126 ) | ( ~n1125 & n1127 ) | ( n1126 & n1127 ) ;
  assign n1129 = ( x307 & x308 ) | ( x307 & n1125 ) | ( x308 & n1125 ) ;
  assign n1130 = ( x309 & ~x310 ) | ( x309 & n1129 ) | ( ~x310 & n1129 ) ;
  assign n1131 = ( ~x309 & x310 ) | ( ~x309 & n1130 ) | ( x310 & n1130 ) ;
  assign n1132 = ( ~n1129 & n1130 ) | ( ~n1129 & n1131 ) | ( n1130 & n1131 ) ;
  assign n1133 = ( x309 & x310 ) | ( x309 & n1129 ) | ( x310 & n1129 ) ;
  assign n1134 = ( x311 & ~x312 ) | ( x311 & n1133 ) | ( ~x312 & n1133 ) ;
  assign n1135 = ( ~x311 & x312 ) | ( ~x311 & n1134 ) | ( x312 & n1134 ) ;
  assign n1136 = ( ~n1133 & n1134 ) | ( ~n1133 & n1135 ) | ( n1134 & n1135 ) ;
  assign n1137 = ( x311 & x312 ) | ( x311 & n1133 ) | ( x312 & n1133 ) ;
  assign n1138 = ( x313 & ~x314 ) | ( x313 & n1137 ) | ( ~x314 & n1137 ) ;
  assign n1139 = ( ~x313 & x314 ) | ( ~x313 & n1138 ) | ( x314 & n1138 ) ;
  assign n1140 = ( ~n1137 & n1138 ) | ( ~n1137 & n1139 ) | ( n1138 & n1139 ) ;
  assign n1141 = ( x313 & x314 ) | ( x313 & n1137 ) | ( x314 & n1137 ) ;
  assign n1142 = ( x315 & ~x316 ) | ( x315 & n1141 ) | ( ~x316 & n1141 ) ;
  assign n1143 = ( ~x315 & x316 ) | ( ~x315 & n1142 ) | ( x316 & n1142 ) ;
  assign n1144 = ( ~n1141 & n1142 ) | ( ~n1141 & n1143 ) | ( n1142 & n1143 ) ;
  assign n1145 = ( x315 & x316 ) | ( x315 & n1141 ) | ( x316 & n1141 ) ;
  assign n1146 = ( x317 & ~x318 ) | ( x317 & n1145 ) | ( ~x318 & n1145 ) ;
  assign n1147 = ( ~x317 & x318 ) | ( ~x317 & n1146 ) | ( x318 & n1146 ) ;
  assign n1148 = ( ~n1145 & n1146 ) | ( ~n1145 & n1147 ) | ( n1146 & n1147 ) ;
  assign n1149 = ( x317 & x318 ) | ( x317 & n1145 ) | ( x318 & n1145 ) ;
  assign n1150 = ( x319 & ~x320 ) | ( x319 & n1149 ) | ( ~x320 & n1149 ) ;
  assign n1151 = ( ~x319 & x320 ) | ( ~x319 & n1150 ) | ( x320 & n1150 ) ;
  assign n1152 = ( ~n1149 & n1150 ) | ( ~n1149 & n1151 ) | ( n1150 & n1151 ) ;
  assign n1153 = ( x319 & x320 ) | ( x319 & n1149 ) | ( x320 & n1149 ) ;
  assign n1154 = ( x321 & ~x322 ) | ( x321 & n1153 ) | ( ~x322 & n1153 ) ;
  assign n1155 = ( ~x321 & x322 ) | ( ~x321 & n1154 ) | ( x322 & n1154 ) ;
  assign n1156 = ( ~n1153 & n1154 ) | ( ~n1153 & n1155 ) | ( n1154 & n1155 ) ;
  assign n1157 = ( x321 & x322 ) | ( x321 & n1153 ) | ( x322 & n1153 ) ;
  assign n1158 = ( x323 & ~x324 ) | ( x323 & n1157 ) | ( ~x324 & n1157 ) ;
  assign n1159 = ( ~x323 & x324 ) | ( ~x323 & n1158 ) | ( x324 & n1158 ) ;
  assign n1160 = ( ~n1157 & n1158 ) | ( ~n1157 & n1159 ) | ( n1158 & n1159 ) ;
  assign n1161 = ( x323 & x324 ) | ( x323 & n1157 ) | ( x324 & n1157 ) ;
  assign n1162 = ( x325 & ~x326 ) | ( x325 & n1161 ) | ( ~x326 & n1161 ) ;
  assign n1163 = ( ~x325 & x326 ) | ( ~x325 & n1162 ) | ( x326 & n1162 ) ;
  assign n1164 = ( ~n1161 & n1162 ) | ( ~n1161 & n1163 ) | ( n1162 & n1163 ) ;
  assign n1165 = ( x325 & x326 ) | ( x325 & n1161 ) | ( x326 & n1161 ) ;
  assign n1166 = ( x327 & ~x328 ) | ( x327 & n1165 ) | ( ~x328 & n1165 ) ;
  assign n1167 = ( ~x327 & x328 ) | ( ~x327 & n1166 ) | ( x328 & n1166 ) ;
  assign n1168 = ( ~n1165 & n1166 ) | ( ~n1165 & n1167 ) | ( n1166 & n1167 ) ;
  assign n1169 = ( x327 & x328 ) | ( x327 & n1165 ) | ( x328 & n1165 ) ;
  assign n1170 = ( x329 & ~x330 ) | ( x329 & n1169 ) | ( ~x330 & n1169 ) ;
  assign n1171 = ( ~x329 & x330 ) | ( ~x329 & n1170 ) | ( x330 & n1170 ) ;
  assign n1172 = ( ~n1169 & n1170 ) | ( ~n1169 & n1171 ) | ( n1170 & n1171 ) ;
  assign n1173 = ( x329 & x330 ) | ( x329 & n1169 ) | ( x330 & n1169 ) ;
  assign n1174 = ( x331 & ~x332 ) | ( x331 & n1173 ) | ( ~x332 & n1173 ) ;
  assign n1175 = ( ~x331 & x332 ) | ( ~x331 & n1174 ) | ( x332 & n1174 ) ;
  assign n1176 = ( ~n1173 & n1174 ) | ( ~n1173 & n1175 ) | ( n1174 & n1175 ) ;
  assign n1177 = ( x331 & x332 ) | ( x331 & n1173 ) | ( x332 & n1173 ) ;
  assign n1178 = ( x333 & ~x334 ) | ( x333 & n1177 ) | ( ~x334 & n1177 ) ;
  assign n1179 = ( ~x333 & x334 ) | ( ~x333 & n1178 ) | ( x334 & n1178 ) ;
  assign n1180 = ( ~n1177 & n1178 ) | ( ~n1177 & n1179 ) | ( n1178 & n1179 ) ;
  assign n1181 = ( x333 & x334 ) | ( x333 & n1177 ) | ( x334 & n1177 ) ;
  assign n1182 = ( x335 & ~x336 ) | ( x335 & n1181 ) | ( ~x336 & n1181 ) ;
  assign n1183 = ( ~x335 & x336 ) | ( ~x335 & n1182 ) | ( x336 & n1182 ) ;
  assign n1184 = ( ~n1181 & n1182 ) | ( ~n1181 & n1183 ) | ( n1182 & n1183 ) ;
  assign n1185 = ( x335 & x336 ) | ( x335 & n1181 ) | ( x336 & n1181 ) ;
  assign n1186 = ( x337 & ~x338 ) | ( x337 & n1185 ) | ( ~x338 & n1185 ) ;
  assign n1187 = ( ~x337 & x338 ) | ( ~x337 & n1186 ) | ( x338 & n1186 ) ;
  assign n1188 = ( ~n1185 & n1186 ) | ( ~n1185 & n1187 ) | ( n1186 & n1187 ) ;
  assign n1189 = ( x337 & x338 ) | ( x337 & n1185 ) | ( x338 & n1185 ) ;
  assign n1190 = ( x339 & ~x340 ) | ( x339 & n1189 ) | ( ~x340 & n1189 ) ;
  assign n1191 = ( ~x339 & x340 ) | ( ~x339 & n1190 ) | ( x340 & n1190 ) ;
  assign n1192 = ( ~n1189 & n1190 ) | ( ~n1189 & n1191 ) | ( n1190 & n1191 ) ;
  assign n1193 = ( x339 & x340 ) | ( x339 & n1189 ) | ( x340 & n1189 ) ;
  assign n1194 = ( x341 & ~x342 ) | ( x341 & n1193 ) | ( ~x342 & n1193 ) ;
  assign n1195 = ( ~x341 & x342 ) | ( ~x341 & n1194 ) | ( x342 & n1194 ) ;
  assign n1196 = ( ~n1193 & n1194 ) | ( ~n1193 & n1195 ) | ( n1194 & n1195 ) ;
  assign n1197 = ( x341 & x342 ) | ( x341 & n1193 ) | ( x342 & n1193 ) ;
  assign n1198 = ( x343 & ~x344 ) | ( x343 & n1197 ) | ( ~x344 & n1197 ) ;
  assign n1199 = ( ~x343 & x344 ) | ( ~x343 & n1198 ) | ( x344 & n1198 ) ;
  assign n1200 = ( ~n1197 & n1198 ) | ( ~n1197 & n1199 ) | ( n1198 & n1199 ) ;
  assign n1201 = ( x343 & x344 ) | ( x343 & n1197 ) | ( x344 & n1197 ) ;
  assign n1202 = ( x345 & ~x346 ) | ( x345 & n1201 ) | ( ~x346 & n1201 ) ;
  assign n1203 = ( ~x345 & x346 ) | ( ~x345 & n1202 ) | ( x346 & n1202 ) ;
  assign n1204 = ( ~n1201 & n1202 ) | ( ~n1201 & n1203 ) | ( n1202 & n1203 ) ;
  assign n1205 = ( x345 & x346 ) | ( x345 & n1201 ) | ( x346 & n1201 ) ;
  assign n1206 = ( x347 & ~x348 ) | ( x347 & n1205 ) | ( ~x348 & n1205 ) ;
  assign n1207 = ( ~x347 & x348 ) | ( ~x347 & n1206 ) | ( x348 & n1206 ) ;
  assign n1208 = ( ~n1205 & n1206 ) | ( ~n1205 & n1207 ) | ( n1206 & n1207 ) ;
  assign n1209 = ( x347 & x348 ) | ( x347 & n1205 ) | ( x348 & n1205 ) ;
  assign n1210 = ( x349 & ~x350 ) | ( x349 & n1209 ) | ( ~x350 & n1209 ) ;
  assign n1211 = ( ~x349 & x350 ) | ( ~x349 & n1210 ) | ( x350 & n1210 ) ;
  assign n1212 = ( ~n1209 & n1210 ) | ( ~n1209 & n1211 ) | ( n1210 & n1211 ) ;
  assign n1213 = ( x349 & x350 ) | ( x349 & n1209 ) | ( x350 & n1209 ) ;
  assign n1214 = ( x351 & ~x352 ) | ( x351 & n1213 ) | ( ~x352 & n1213 ) ;
  assign n1215 = ( ~x351 & x352 ) | ( ~x351 & n1214 ) | ( x352 & n1214 ) ;
  assign n1216 = ( ~n1213 & n1214 ) | ( ~n1213 & n1215 ) | ( n1214 & n1215 ) ;
  assign n1217 = ( x351 & x352 ) | ( x351 & n1213 ) | ( x352 & n1213 ) ;
  assign n1218 = ( x353 & ~x354 ) | ( x353 & n1217 ) | ( ~x354 & n1217 ) ;
  assign n1219 = ( ~x353 & x354 ) | ( ~x353 & n1218 ) | ( x354 & n1218 ) ;
  assign n1220 = ( ~n1217 & n1218 ) | ( ~n1217 & n1219 ) | ( n1218 & n1219 ) ;
  assign n1221 = ( x353 & x354 ) | ( x353 & n1217 ) | ( x354 & n1217 ) ;
  assign n1222 = ( x355 & ~x356 ) | ( x355 & n1221 ) | ( ~x356 & n1221 ) ;
  assign n1223 = ( ~x355 & x356 ) | ( ~x355 & n1222 ) | ( x356 & n1222 ) ;
  assign n1224 = ( ~n1221 & n1222 ) | ( ~n1221 & n1223 ) | ( n1222 & n1223 ) ;
  assign n1225 = ( x355 & x356 ) | ( x355 & n1221 ) | ( x356 & n1221 ) ;
  assign n1226 = ( x357 & ~x358 ) | ( x357 & n1225 ) | ( ~x358 & n1225 ) ;
  assign n1227 = ( ~x357 & x358 ) | ( ~x357 & n1226 ) | ( x358 & n1226 ) ;
  assign n1228 = ( ~n1225 & n1226 ) | ( ~n1225 & n1227 ) | ( n1226 & n1227 ) ;
  assign n1229 = ( x357 & x358 ) | ( x357 & n1225 ) | ( x358 & n1225 ) ;
  assign n1230 = ( x359 & ~x360 ) | ( x359 & n1229 ) | ( ~x360 & n1229 ) ;
  assign n1231 = ( ~x359 & x360 ) | ( ~x359 & n1230 ) | ( x360 & n1230 ) ;
  assign n1232 = ( ~n1229 & n1230 ) | ( ~n1229 & n1231 ) | ( n1230 & n1231 ) ;
  assign n1233 = ( x359 & x360 ) | ( x359 & n1229 ) | ( x360 & n1229 ) ;
  assign n1234 = ( x361 & ~x362 ) | ( x361 & n1233 ) | ( ~x362 & n1233 ) ;
  assign n1235 = ( ~x361 & x362 ) | ( ~x361 & n1234 ) | ( x362 & n1234 ) ;
  assign n1236 = ( ~n1233 & n1234 ) | ( ~n1233 & n1235 ) | ( n1234 & n1235 ) ;
  assign n1237 = ( x361 & x362 ) | ( x361 & n1233 ) | ( x362 & n1233 ) ;
  assign n1238 = ( x363 & ~x364 ) | ( x363 & n1237 ) | ( ~x364 & n1237 ) ;
  assign n1239 = ( ~x363 & x364 ) | ( ~x363 & n1238 ) | ( x364 & n1238 ) ;
  assign n1240 = ( ~n1237 & n1238 ) | ( ~n1237 & n1239 ) | ( n1238 & n1239 ) ;
  assign n1241 = ( x363 & x364 ) | ( x363 & n1237 ) | ( x364 & n1237 ) ;
  assign n1242 = ( x365 & ~x366 ) | ( x365 & n1241 ) | ( ~x366 & n1241 ) ;
  assign n1243 = ( ~x365 & x366 ) | ( ~x365 & n1242 ) | ( x366 & n1242 ) ;
  assign n1244 = ( ~n1241 & n1242 ) | ( ~n1241 & n1243 ) | ( n1242 & n1243 ) ;
  assign n1245 = ( x365 & x366 ) | ( x365 & n1241 ) | ( x366 & n1241 ) ;
  assign n1246 = ( x367 & ~x368 ) | ( x367 & n1245 ) | ( ~x368 & n1245 ) ;
  assign n1247 = ( ~x367 & x368 ) | ( ~x367 & n1246 ) | ( x368 & n1246 ) ;
  assign n1248 = ( ~n1245 & n1246 ) | ( ~n1245 & n1247 ) | ( n1246 & n1247 ) ;
  assign n1249 = ( x367 & x368 ) | ( x367 & n1245 ) | ( x368 & n1245 ) ;
  assign n1250 = ( x369 & ~x370 ) | ( x369 & n1249 ) | ( ~x370 & n1249 ) ;
  assign n1251 = ( ~x369 & x370 ) | ( ~x369 & n1250 ) | ( x370 & n1250 ) ;
  assign n1252 = ( ~n1249 & n1250 ) | ( ~n1249 & n1251 ) | ( n1250 & n1251 ) ;
  assign n1253 = ( x369 & x370 ) | ( x369 & n1249 ) | ( x370 & n1249 ) ;
  assign n1254 = ( x371 & ~x372 ) | ( x371 & n1253 ) | ( ~x372 & n1253 ) ;
  assign n1255 = ( ~x371 & x372 ) | ( ~x371 & n1254 ) | ( x372 & n1254 ) ;
  assign n1256 = ( ~n1253 & n1254 ) | ( ~n1253 & n1255 ) | ( n1254 & n1255 ) ;
  assign n1257 = ( x371 & x372 ) | ( x371 & n1253 ) | ( x372 & n1253 ) ;
  assign n1258 = ( x373 & ~x374 ) | ( x373 & n1257 ) | ( ~x374 & n1257 ) ;
  assign n1259 = ( ~x373 & x374 ) | ( ~x373 & n1258 ) | ( x374 & n1258 ) ;
  assign n1260 = ( ~n1257 & n1258 ) | ( ~n1257 & n1259 ) | ( n1258 & n1259 ) ;
  assign n1261 = ( x373 & x374 ) | ( x373 & n1257 ) | ( x374 & n1257 ) ;
  assign n1262 = ( x375 & ~x376 ) | ( x375 & n1261 ) | ( ~x376 & n1261 ) ;
  assign n1263 = ( ~x375 & x376 ) | ( ~x375 & n1262 ) | ( x376 & n1262 ) ;
  assign n1264 = ( ~n1261 & n1262 ) | ( ~n1261 & n1263 ) | ( n1262 & n1263 ) ;
  assign n1265 = ( x375 & x376 ) | ( x375 & n1261 ) | ( x376 & n1261 ) ;
  assign n1266 = ( x377 & ~x378 ) | ( x377 & n1265 ) | ( ~x378 & n1265 ) ;
  assign n1267 = ( ~x377 & x378 ) | ( ~x377 & n1266 ) | ( x378 & n1266 ) ;
  assign n1268 = ( ~n1265 & n1266 ) | ( ~n1265 & n1267 ) | ( n1266 & n1267 ) ;
  assign n1269 = ( x377 & x378 ) | ( x377 & n1265 ) | ( x378 & n1265 ) ;
  assign n1270 = ( x379 & ~x380 ) | ( x379 & n1269 ) | ( ~x380 & n1269 ) ;
  assign n1271 = ( ~x379 & x380 ) | ( ~x379 & n1270 ) | ( x380 & n1270 ) ;
  assign n1272 = ( ~n1269 & n1270 ) | ( ~n1269 & n1271 ) | ( n1270 & n1271 ) ;
  assign n1273 = ( x379 & x380 ) | ( x379 & n1269 ) | ( x380 & n1269 ) ;
  assign n1274 = ( x381 & ~x382 ) | ( x381 & n1273 ) | ( ~x382 & n1273 ) ;
  assign n1275 = ( ~x381 & x382 ) | ( ~x381 & n1274 ) | ( x382 & n1274 ) ;
  assign n1276 = ( ~n1273 & n1274 ) | ( ~n1273 & n1275 ) | ( n1274 & n1275 ) ;
  assign n1277 = ( x381 & x382 ) | ( x381 & n1273 ) | ( x382 & n1273 ) ;
  assign n1278 = ( x383 & ~x384 ) | ( x383 & n1277 ) | ( ~x384 & n1277 ) ;
  assign n1279 = ( ~x383 & x384 ) | ( ~x383 & n1278 ) | ( x384 & n1278 ) ;
  assign n1280 = ( ~n1277 & n1278 ) | ( ~n1277 & n1279 ) | ( n1278 & n1279 ) ;
  assign n1281 = ( x383 & x384 ) | ( x383 & n1277 ) | ( x384 & n1277 ) ;
  assign n1282 = ( x385 & ~x386 ) | ( x385 & n1281 ) | ( ~x386 & n1281 ) ;
  assign n1283 = ( ~x385 & x386 ) | ( ~x385 & n1282 ) | ( x386 & n1282 ) ;
  assign n1284 = ( ~n1281 & n1282 ) | ( ~n1281 & n1283 ) | ( n1282 & n1283 ) ;
  assign n1285 = ( x385 & x386 ) | ( x385 & n1281 ) | ( x386 & n1281 ) ;
  assign n1286 = ( x387 & ~x388 ) | ( x387 & n1285 ) | ( ~x388 & n1285 ) ;
  assign n1287 = ( ~x387 & x388 ) | ( ~x387 & n1286 ) | ( x388 & n1286 ) ;
  assign n1288 = ( ~n1285 & n1286 ) | ( ~n1285 & n1287 ) | ( n1286 & n1287 ) ;
  assign n1289 = ( x387 & x388 ) | ( x387 & n1285 ) | ( x388 & n1285 ) ;
  assign n1290 = ( x389 & ~x390 ) | ( x389 & n1289 ) | ( ~x390 & n1289 ) ;
  assign n1291 = ( ~x389 & x390 ) | ( ~x389 & n1290 ) | ( x390 & n1290 ) ;
  assign n1292 = ( ~n1289 & n1290 ) | ( ~n1289 & n1291 ) | ( n1290 & n1291 ) ;
  assign n1293 = ( x389 & x390 ) | ( x389 & n1289 ) | ( x390 & n1289 ) ;
  assign n1294 = ( x391 & ~x392 ) | ( x391 & n1293 ) | ( ~x392 & n1293 ) ;
  assign n1295 = ( ~x391 & x392 ) | ( ~x391 & n1294 ) | ( x392 & n1294 ) ;
  assign n1296 = ( ~n1293 & n1294 ) | ( ~n1293 & n1295 ) | ( n1294 & n1295 ) ;
  assign n1297 = ( x391 & x392 ) | ( x391 & n1293 ) | ( x392 & n1293 ) ;
  assign n1298 = ( x393 & ~x394 ) | ( x393 & n1297 ) | ( ~x394 & n1297 ) ;
  assign n1299 = ( ~x393 & x394 ) | ( ~x393 & n1298 ) | ( x394 & n1298 ) ;
  assign n1300 = ( ~n1297 & n1298 ) | ( ~n1297 & n1299 ) | ( n1298 & n1299 ) ;
  assign n1301 = ( x393 & x394 ) | ( x393 & n1297 ) | ( x394 & n1297 ) ;
  assign n1302 = ( x395 & ~x396 ) | ( x395 & n1301 ) | ( ~x396 & n1301 ) ;
  assign n1303 = ( ~x395 & x396 ) | ( ~x395 & n1302 ) | ( x396 & n1302 ) ;
  assign n1304 = ( ~n1301 & n1302 ) | ( ~n1301 & n1303 ) | ( n1302 & n1303 ) ;
  assign n1305 = ( x395 & x396 ) | ( x395 & n1301 ) | ( x396 & n1301 ) ;
  assign n1306 = ( x397 & ~x398 ) | ( x397 & n1305 ) | ( ~x398 & n1305 ) ;
  assign n1307 = ( ~x397 & x398 ) | ( ~x397 & n1306 ) | ( x398 & n1306 ) ;
  assign n1308 = ( ~n1305 & n1306 ) | ( ~n1305 & n1307 ) | ( n1306 & n1307 ) ;
  assign n1309 = ( x397 & x398 ) | ( x397 & n1305 ) | ( x398 & n1305 ) ;
  assign n1310 = ( x399 & ~x400 ) | ( x399 & n1309 ) | ( ~x400 & n1309 ) ;
  assign n1311 = ( ~x399 & x400 ) | ( ~x399 & n1310 ) | ( x400 & n1310 ) ;
  assign n1312 = ( ~n1309 & n1310 ) | ( ~n1309 & n1311 ) | ( n1310 & n1311 ) ;
  assign n1313 = ( x399 & x400 ) | ( x399 & n1309 ) | ( x400 & n1309 ) ;
  assign n1314 = ( x401 & ~x402 ) | ( x401 & n1313 ) | ( ~x402 & n1313 ) ;
  assign n1315 = ( ~x401 & x402 ) | ( ~x401 & n1314 ) | ( x402 & n1314 ) ;
  assign n1316 = ( ~n1313 & n1314 ) | ( ~n1313 & n1315 ) | ( n1314 & n1315 ) ;
  assign n1317 = ( x401 & x402 ) | ( x401 & n1313 ) | ( x402 & n1313 ) ;
  assign n1318 = ( x403 & ~x404 ) | ( x403 & n1317 ) | ( ~x404 & n1317 ) ;
  assign n1319 = ( ~x403 & x404 ) | ( ~x403 & n1318 ) | ( x404 & n1318 ) ;
  assign n1320 = ( ~n1317 & n1318 ) | ( ~n1317 & n1319 ) | ( n1318 & n1319 ) ;
  assign n1321 = ( x403 & x404 ) | ( x403 & n1317 ) | ( x404 & n1317 ) ;
  assign n1322 = ( x405 & ~x406 ) | ( x405 & n1321 ) | ( ~x406 & n1321 ) ;
  assign n1323 = ( ~x405 & x406 ) | ( ~x405 & n1322 ) | ( x406 & n1322 ) ;
  assign n1324 = ( ~n1321 & n1322 ) | ( ~n1321 & n1323 ) | ( n1322 & n1323 ) ;
  assign n1325 = ( x405 & x406 ) | ( x405 & n1321 ) | ( x406 & n1321 ) ;
  assign n1326 = ( x407 & ~x408 ) | ( x407 & n1325 ) | ( ~x408 & n1325 ) ;
  assign n1327 = ( ~x407 & x408 ) | ( ~x407 & n1326 ) | ( x408 & n1326 ) ;
  assign n1328 = ( ~n1325 & n1326 ) | ( ~n1325 & n1327 ) | ( n1326 & n1327 ) ;
  assign n1329 = ( x407 & x408 ) | ( x407 & n1325 ) | ( x408 & n1325 ) ;
  assign n1330 = ( x409 & ~x410 ) | ( x409 & n1329 ) | ( ~x410 & n1329 ) ;
  assign n1331 = ( ~x409 & x410 ) | ( ~x409 & n1330 ) | ( x410 & n1330 ) ;
  assign n1332 = ( ~n1329 & n1330 ) | ( ~n1329 & n1331 ) | ( n1330 & n1331 ) ;
  assign n1333 = ( x409 & x410 ) | ( x409 & n1329 ) | ( x410 & n1329 ) ;
  assign n1334 = ( x411 & ~x412 ) | ( x411 & n1333 ) | ( ~x412 & n1333 ) ;
  assign n1335 = ( ~x411 & x412 ) | ( ~x411 & n1334 ) | ( x412 & n1334 ) ;
  assign n1336 = ( ~n1333 & n1334 ) | ( ~n1333 & n1335 ) | ( n1334 & n1335 ) ;
  assign n1337 = ( x411 & x412 ) | ( x411 & n1333 ) | ( x412 & n1333 ) ;
  assign n1338 = ( x413 & ~x414 ) | ( x413 & n1337 ) | ( ~x414 & n1337 ) ;
  assign n1339 = ( ~x413 & x414 ) | ( ~x413 & n1338 ) | ( x414 & n1338 ) ;
  assign n1340 = ( ~n1337 & n1338 ) | ( ~n1337 & n1339 ) | ( n1338 & n1339 ) ;
  assign n1341 = ( x413 & x414 ) | ( x413 & n1337 ) | ( x414 & n1337 ) ;
  assign n1342 = ( x415 & ~x416 ) | ( x415 & n1341 ) | ( ~x416 & n1341 ) ;
  assign n1343 = ( ~x415 & x416 ) | ( ~x415 & n1342 ) | ( x416 & n1342 ) ;
  assign n1344 = ( ~n1341 & n1342 ) | ( ~n1341 & n1343 ) | ( n1342 & n1343 ) ;
  assign n1345 = ( x415 & x416 ) | ( x415 & n1341 ) | ( x416 & n1341 ) ;
  assign n1346 = ( x417 & ~x418 ) | ( x417 & n1345 ) | ( ~x418 & n1345 ) ;
  assign n1347 = ( ~x417 & x418 ) | ( ~x417 & n1346 ) | ( x418 & n1346 ) ;
  assign n1348 = ( ~n1345 & n1346 ) | ( ~n1345 & n1347 ) | ( n1346 & n1347 ) ;
  assign n1349 = ( x417 & x418 ) | ( x417 & n1345 ) | ( x418 & n1345 ) ;
  assign n1350 = ( x419 & ~x420 ) | ( x419 & n1349 ) | ( ~x420 & n1349 ) ;
  assign n1351 = ( ~x419 & x420 ) | ( ~x419 & n1350 ) | ( x420 & n1350 ) ;
  assign n1352 = ( ~n1349 & n1350 ) | ( ~n1349 & n1351 ) | ( n1350 & n1351 ) ;
  assign n1353 = ( x419 & x420 ) | ( x419 & n1349 ) | ( x420 & n1349 ) ;
  assign n1354 = ( x421 & ~x422 ) | ( x421 & n1353 ) | ( ~x422 & n1353 ) ;
  assign n1355 = ( ~x421 & x422 ) | ( ~x421 & n1354 ) | ( x422 & n1354 ) ;
  assign n1356 = ( ~n1353 & n1354 ) | ( ~n1353 & n1355 ) | ( n1354 & n1355 ) ;
  assign n1357 = ( x421 & x422 ) | ( x421 & n1353 ) | ( x422 & n1353 ) ;
  assign n1358 = ( x423 & ~x424 ) | ( x423 & n1357 ) | ( ~x424 & n1357 ) ;
  assign n1359 = ( ~x423 & x424 ) | ( ~x423 & n1358 ) | ( x424 & n1358 ) ;
  assign n1360 = ( ~n1357 & n1358 ) | ( ~n1357 & n1359 ) | ( n1358 & n1359 ) ;
  assign n1361 = ( x423 & x424 ) | ( x423 & n1357 ) | ( x424 & n1357 ) ;
  assign n1362 = ( x425 & ~x426 ) | ( x425 & n1361 ) | ( ~x426 & n1361 ) ;
  assign n1363 = ( ~x425 & x426 ) | ( ~x425 & n1362 ) | ( x426 & n1362 ) ;
  assign n1364 = ( ~n1361 & n1362 ) | ( ~n1361 & n1363 ) | ( n1362 & n1363 ) ;
  assign n1365 = ( x425 & x426 ) | ( x425 & n1361 ) | ( x426 & n1361 ) ;
  assign n1366 = ( x427 & ~x428 ) | ( x427 & n1365 ) | ( ~x428 & n1365 ) ;
  assign n1367 = ( ~x427 & x428 ) | ( ~x427 & n1366 ) | ( x428 & n1366 ) ;
  assign n1368 = ( ~n1365 & n1366 ) | ( ~n1365 & n1367 ) | ( n1366 & n1367 ) ;
  assign n1369 = ( x427 & x428 ) | ( x427 & n1365 ) | ( x428 & n1365 ) ;
  assign n1370 = ( x429 & ~x430 ) | ( x429 & n1369 ) | ( ~x430 & n1369 ) ;
  assign n1371 = ( ~x429 & x430 ) | ( ~x429 & n1370 ) | ( x430 & n1370 ) ;
  assign n1372 = ( ~n1369 & n1370 ) | ( ~n1369 & n1371 ) | ( n1370 & n1371 ) ;
  assign n1373 = ( x429 & x430 ) | ( x429 & n1369 ) | ( x430 & n1369 ) ;
  assign n1374 = ( x431 & ~x432 ) | ( x431 & n1373 ) | ( ~x432 & n1373 ) ;
  assign n1375 = ( ~x431 & x432 ) | ( ~x431 & n1374 ) | ( x432 & n1374 ) ;
  assign n1376 = ( ~n1373 & n1374 ) | ( ~n1373 & n1375 ) | ( n1374 & n1375 ) ;
  assign n1377 = ( x431 & x432 ) | ( x431 & n1373 ) | ( x432 & n1373 ) ;
  assign n1378 = ( x433 & ~x434 ) | ( x433 & n1377 ) | ( ~x434 & n1377 ) ;
  assign n1379 = ( ~x433 & x434 ) | ( ~x433 & n1378 ) | ( x434 & n1378 ) ;
  assign n1380 = ( ~n1377 & n1378 ) | ( ~n1377 & n1379 ) | ( n1378 & n1379 ) ;
  assign n1381 = ( x433 & x434 ) | ( x433 & n1377 ) | ( x434 & n1377 ) ;
  assign n1382 = ( x435 & ~x436 ) | ( x435 & n1381 ) | ( ~x436 & n1381 ) ;
  assign n1383 = ( ~x435 & x436 ) | ( ~x435 & n1382 ) | ( x436 & n1382 ) ;
  assign n1384 = ( ~n1381 & n1382 ) | ( ~n1381 & n1383 ) | ( n1382 & n1383 ) ;
  assign n1385 = ( x435 & x436 ) | ( x435 & n1381 ) | ( x436 & n1381 ) ;
  assign n1386 = ( x437 & ~x438 ) | ( x437 & n1385 ) | ( ~x438 & n1385 ) ;
  assign n1387 = ( ~x437 & x438 ) | ( ~x437 & n1386 ) | ( x438 & n1386 ) ;
  assign n1388 = ( ~n1385 & n1386 ) | ( ~n1385 & n1387 ) | ( n1386 & n1387 ) ;
  assign n1389 = ( x437 & x438 ) | ( x437 & n1385 ) | ( x438 & n1385 ) ;
  assign n1390 = ( x439 & ~x440 ) | ( x439 & n1389 ) | ( ~x440 & n1389 ) ;
  assign n1391 = ( ~x439 & x440 ) | ( ~x439 & n1390 ) | ( x440 & n1390 ) ;
  assign n1392 = ( ~n1389 & n1390 ) | ( ~n1389 & n1391 ) | ( n1390 & n1391 ) ;
  assign n1393 = ( x439 & x440 ) | ( x439 & n1389 ) | ( x440 & n1389 ) ;
  assign n1394 = ( x441 & ~x442 ) | ( x441 & n1393 ) | ( ~x442 & n1393 ) ;
  assign n1395 = ( ~x441 & x442 ) | ( ~x441 & n1394 ) | ( x442 & n1394 ) ;
  assign n1396 = ( ~n1393 & n1394 ) | ( ~n1393 & n1395 ) | ( n1394 & n1395 ) ;
  assign n1397 = ( x441 & x442 ) | ( x441 & n1393 ) | ( x442 & n1393 ) ;
  assign n1398 = ( x443 & ~x444 ) | ( x443 & n1397 ) | ( ~x444 & n1397 ) ;
  assign n1399 = ( ~x443 & x444 ) | ( ~x443 & n1398 ) | ( x444 & n1398 ) ;
  assign n1400 = ( ~n1397 & n1398 ) | ( ~n1397 & n1399 ) | ( n1398 & n1399 ) ;
  assign n1401 = ( x443 & x444 ) | ( x443 & n1397 ) | ( x444 & n1397 ) ;
  assign n1402 = ( x445 & ~x446 ) | ( x445 & n1401 ) | ( ~x446 & n1401 ) ;
  assign n1403 = ( ~x445 & x446 ) | ( ~x445 & n1402 ) | ( x446 & n1402 ) ;
  assign n1404 = ( ~n1401 & n1402 ) | ( ~n1401 & n1403 ) | ( n1402 & n1403 ) ;
  assign n1405 = ( x445 & x446 ) | ( x445 & n1401 ) | ( x446 & n1401 ) ;
  assign n1406 = ( x447 & ~x448 ) | ( x447 & n1405 ) | ( ~x448 & n1405 ) ;
  assign n1407 = ( ~x447 & x448 ) | ( ~x447 & n1406 ) | ( x448 & n1406 ) ;
  assign n1408 = ( ~n1405 & n1406 ) | ( ~n1405 & n1407 ) | ( n1406 & n1407 ) ;
  assign n1409 = ( x447 & x448 ) | ( x447 & n1405 ) | ( x448 & n1405 ) ;
  assign n1410 = ( x449 & ~x450 ) | ( x449 & n1409 ) | ( ~x450 & n1409 ) ;
  assign n1411 = ( ~x449 & x450 ) | ( ~x449 & n1410 ) | ( x450 & n1410 ) ;
  assign n1412 = ( ~n1409 & n1410 ) | ( ~n1409 & n1411 ) | ( n1410 & n1411 ) ;
  assign n1413 = ( x449 & x450 ) | ( x449 & n1409 ) | ( x450 & n1409 ) ;
  assign n1414 = ( x451 & ~x452 ) | ( x451 & n1413 ) | ( ~x452 & n1413 ) ;
  assign n1415 = ( ~x451 & x452 ) | ( ~x451 & n1414 ) | ( x452 & n1414 ) ;
  assign n1416 = ( ~n1413 & n1414 ) | ( ~n1413 & n1415 ) | ( n1414 & n1415 ) ;
  assign n1417 = ( x451 & x452 ) | ( x451 & n1413 ) | ( x452 & n1413 ) ;
  assign n1418 = ( x453 & ~x454 ) | ( x453 & n1417 ) | ( ~x454 & n1417 ) ;
  assign n1419 = ( ~x453 & x454 ) | ( ~x453 & n1418 ) | ( x454 & n1418 ) ;
  assign n1420 = ( ~n1417 & n1418 ) | ( ~n1417 & n1419 ) | ( n1418 & n1419 ) ;
  assign n1421 = ( x453 & x454 ) | ( x453 & n1417 ) | ( x454 & n1417 ) ;
  assign n1422 = ( x455 & ~x456 ) | ( x455 & n1421 ) | ( ~x456 & n1421 ) ;
  assign n1423 = ( ~x455 & x456 ) | ( ~x455 & n1422 ) | ( x456 & n1422 ) ;
  assign n1424 = ( ~n1421 & n1422 ) | ( ~n1421 & n1423 ) | ( n1422 & n1423 ) ;
  assign n1425 = ( x455 & x456 ) | ( x455 & n1421 ) | ( x456 & n1421 ) ;
  assign n1426 = ( x457 & ~x458 ) | ( x457 & n1425 ) | ( ~x458 & n1425 ) ;
  assign n1427 = ( ~x457 & x458 ) | ( ~x457 & n1426 ) | ( x458 & n1426 ) ;
  assign n1428 = ( ~n1425 & n1426 ) | ( ~n1425 & n1427 ) | ( n1426 & n1427 ) ;
  assign n1429 = ( x457 & x458 ) | ( x457 & n1425 ) | ( x458 & n1425 ) ;
  assign n1430 = ( x459 & ~x460 ) | ( x459 & n1429 ) | ( ~x460 & n1429 ) ;
  assign n1431 = ( ~x459 & x460 ) | ( ~x459 & n1430 ) | ( x460 & n1430 ) ;
  assign n1432 = ( ~n1429 & n1430 ) | ( ~n1429 & n1431 ) | ( n1430 & n1431 ) ;
  assign n1433 = ( x459 & x460 ) | ( x459 & n1429 ) | ( x460 & n1429 ) ;
  assign n1434 = ( x461 & ~x462 ) | ( x461 & n1433 ) | ( ~x462 & n1433 ) ;
  assign n1435 = ( ~x461 & x462 ) | ( ~x461 & n1434 ) | ( x462 & n1434 ) ;
  assign n1436 = ( ~n1433 & n1434 ) | ( ~n1433 & n1435 ) | ( n1434 & n1435 ) ;
  assign n1437 = ( x461 & x462 ) | ( x461 & n1433 ) | ( x462 & n1433 ) ;
  assign n1438 = ( x463 & ~x464 ) | ( x463 & n1437 ) | ( ~x464 & n1437 ) ;
  assign n1439 = ( ~x463 & x464 ) | ( ~x463 & n1438 ) | ( x464 & n1438 ) ;
  assign n1440 = ( ~n1437 & n1438 ) | ( ~n1437 & n1439 ) | ( n1438 & n1439 ) ;
  assign n1441 = ( x463 & x464 ) | ( x463 & n1437 ) | ( x464 & n1437 ) ;
  assign n1442 = ( x465 & ~x466 ) | ( x465 & n1441 ) | ( ~x466 & n1441 ) ;
  assign n1443 = ( ~x465 & x466 ) | ( ~x465 & n1442 ) | ( x466 & n1442 ) ;
  assign n1444 = ( ~n1441 & n1442 ) | ( ~n1441 & n1443 ) | ( n1442 & n1443 ) ;
  assign n1445 = ( x465 & x466 ) | ( x465 & n1441 ) | ( x466 & n1441 ) ;
  assign n1446 = ( x467 & ~x468 ) | ( x467 & n1445 ) | ( ~x468 & n1445 ) ;
  assign n1447 = ( ~x467 & x468 ) | ( ~x467 & n1446 ) | ( x468 & n1446 ) ;
  assign n1448 = ( ~n1445 & n1446 ) | ( ~n1445 & n1447 ) | ( n1446 & n1447 ) ;
  assign n1449 = ( x467 & x468 ) | ( x467 & n1445 ) | ( x468 & n1445 ) ;
  assign n1450 = ( x469 & ~x470 ) | ( x469 & n1449 ) | ( ~x470 & n1449 ) ;
  assign n1451 = ( ~x469 & x470 ) | ( ~x469 & n1450 ) | ( x470 & n1450 ) ;
  assign n1452 = ( ~n1449 & n1450 ) | ( ~n1449 & n1451 ) | ( n1450 & n1451 ) ;
  assign n1453 = ( x469 & x470 ) | ( x469 & n1449 ) | ( x470 & n1449 ) ;
  assign n1454 = ( x471 & ~x472 ) | ( x471 & n1453 ) | ( ~x472 & n1453 ) ;
  assign n1455 = ( ~x471 & x472 ) | ( ~x471 & n1454 ) | ( x472 & n1454 ) ;
  assign n1456 = ( ~n1453 & n1454 ) | ( ~n1453 & n1455 ) | ( n1454 & n1455 ) ;
  assign n1457 = ( x471 & x472 ) | ( x471 & n1453 ) | ( x472 & n1453 ) ;
  assign n1458 = ( x473 & ~x474 ) | ( x473 & n1457 ) | ( ~x474 & n1457 ) ;
  assign n1459 = ( ~x473 & x474 ) | ( ~x473 & n1458 ) | ( x474 & n1458 ) ;
  assign n1460 = ( ~n1457 & n1458 ) | ( ~n1457 & n1459 ) | ( n1458 & n1459 ) ;
  assign n1461 = ( x473 & x474 ) | ( x473 & n1457 ) | ( x474 & n1457 ) ;
  assign n1462 = ( x475 & ~x476 ) | ( x475 & n1461 ) | ( ~x476 & n1461 ) ;
  assign n1463 = ( ~x475 & x476 ) | ( ~x475 & n1462 ) | ( x476 & n1462 ) ;
  assign n1464 = ( ~n1461 & n1462 ) | ( ~n1461 & n1463 ) | ( n1462 & n1463 ) ;
  assign n1465 = ( x475 & x476 ) | ( x475 & n1461 ) | ( x476 & n1461 ) ;
  assign n1466 = ( x477 & ~x478 ) | ( x477 & n1465 ) | ( ~x478 & n1465 ) ;
  assign n1467 = ( ~x477 & x478 ) | ( ~x477 & n1466 ) | ( x478 & n1466 ) ;
  assign n1468 = ( ~n1465 & n1466 ) | ( ~n1465 & n1467 ) | ( n1466 & n1467 ) ;
  assign n1469 = ( x477 & x478 ) | ( x477 & n1465 ) | ( x478 & n1465 ) ;
  assign n1470 = ( x479 & ~x480 ) | ( x479 & n1469 ) | ( ~x480 & n1469 ) ;
  assign n1471 = ( ~x479 & x480 ) | ( ~x479 & n1470 ) | ( x480 & n1470 ) ;
  assign n1472 = ( ~n1469 & n1470 ) | ( ~n1469 & n1471 ) | ( n1470 & n1471 ) ;
  assign n1473 = ( x479 & x480 ) | ( x479 & n1469 ) | ( x480 & n1469 ) ;
  assign n1474 = ( x481 & ~x482 ) | ( x481 & n1473 ) | ( ~x482 & n1473 ) ;
  assign n1475 = ( ~x481 & x482 ) | ( ~x481 & n1474 ) | ( x482 & n1474 ) ;
  assign n1476 = ( ~n1473 & n1474 ) | ( ~n1473 & n1475 ) | ( n1474 & n1475 ) ;
  assign n1477 = ( x481 & x482 ) | ( x481 & n1473 ) | ( x482 & n1473 ) ;
  assign n1478 = ( x483 & ~x484 ) | ( x483 & n1477 ) | ( ~x484 & n1477 ) ;
  assign n1479 = ( ~x483 & x484 ) | ( ~x483 & n1478 ) | ( x484 & n1478 ) ;
  assign n1480 = ( ~n1477 & n1478 ) | ( ~n1477 & n1479 ) | ( n1478 & n1479 ) ;
  assign n1481 = ( x483 & x484 ) | ( x483 & n1477 ) | ( x484 & n1477 ) ;
  assign n1482 = ( x485 & ~x486 ) | ( x485 & n1481 ) | ( ~x486 & n1481 ) ;
  assign n1483 = ( ~x485 & x486 ) | ( ~x485 & n1482 ) | ( x486 & n1482 ) ;
  assign n1484 = ( ~n1481 & n1482 ) | ( ~n1481 & n1483 ) | ( n1482 & n1483 ) ;
  assign n1485 = ( x485 & x486 ) | ( x485 & n1481 ) | ( x486 & n1481 ) ;
  assign n1486 = ( x487 & ~x488 ) | ( x487 & n1485 ) | ( ~x488 & n1485 ) ;
  assign n1487 = ( ~x487 & x488 ) | ( ~x487 & n1486 ) | ( x488 & n1486 ) ;
  assign n1488 = ( ~n1485 & n1486 ) | ( ~n1485 & n1487 ) | ( n1486 & n1487 ) ;
  assign n1489 = ( x487 & x488 ) | ( x487 & n1485 ) | ( x488 & n1485 ) ;
  assign n1490 = ( x489 & ~x490 ) | ( x489 & n1489 ) | ( ~x490 & n1489 ) ;
  assign n1491 = ( ~x489 & x490 ) | ( ~x489 & n1490 ) | ( x490 & n1490 ) ;
  assign n1492 = ( ~n1489 & n1490 ) | ( ~n1489 & n1491 ) | ( n1490 & n1491 ) ;
  assign n1493 = ( x489 & x490 ) | ( x489 & n1489 ) | ( x490 & n1489 ) ;
  assign n1494 = ( x491 & ~x492 ) | ( x491 & n1493 ) | ( ~x492 & n1493 ) ;
  assign n1495 = ( ~x491 & x492 ) | ( ~x491 & n1494 ) | ( x492 & n1494 ) ;
  assign n1496 = ( ~n1493 & n1494 ) | ( ~n1493 & n1495 ) | ( n1494 & n1495 ) ;
  assign n1497 = ( x491 & x492 ) | ( x491 & n1493 ) | ( x492 & n1493 ) ;
  assign n1498 = ( x493 & ~x494 ) | ( x493 & n1497 ) | ( ~x494 & n1497 ) ;
  assign n1499 = ( ~x493 & x494 ) | ( ~x493 & n1498 ) | ( x494 & n1498 ) ;
  assign n1500 = ( ~n1497 & n1498 ) | ( ~n1497 & n1499 ) | ( n1498 & n1499 ) ;
  assign n1501 = ( x493 & x494 ) | ( x493 & n1497 ) | ( x494 & n1497 ) ;
  assign n1502 = ( x495 & ~x496 ) | ( x495 & n1501 ) | ( ~x496 & n1501 ) ;
  assign n1503 = ( ~x495 & x496 ) | ( ~x495 & n1502 ) | ( x496 & n1502 ) ;
  assign n1504 = ( ~n1501 & n1502 ) | ( ~n1501 & n1503 ) | ( n1502 & n1503 ) ;
  assign n1505 = ( x495 & x496 ) | ( x495 & n1501 ) | ( x496 & n1501 ) ;
  assign n1506 = ( x497 & ~x498 ) | ( x497 & n1505 ) | ( ~x498 & n1505 ) ;
  assign n1507 = ( ~x497 & x498 ) | ( ~x497 & n1506 ) | ( x498 & n1506 ) ;
  assign n1508 = ( ~n1505 & n1506 ) | ( ~n1505 & n1507 ) | ( n1506 & n1507 ) ;
  assign n1509 = ( x497 & x498 ) | ( x497 & n1505 ) | ( x498 & n1505 ) ;
  assign n1510 = ( x499 & ~x500 ) | ( x499 & n1509 ) | ( ~x500 & n1509 ) ;
  assign n1511 = ( ~x499 & x500 ) | ( ~x499 & n1510 ) | ( x500 & n1510 ) ;
  assign n1512 = ( ~n1509 & n1510 ) | ( ~n1509 & n1511 ) | ( n1510 & n1511 ) ;
  assign n1513 = ( x499 & x500 ) | ( x499 & n1509 ) | ( x500 & n1509 ) ;
  assign n1514 = ( x501 & ~x502 ) | ( x501 & n1513 ) | ( ~x502 & n1513 ) ;
  assign n1515 = ( ~x501 & x502 ) | ( ~x501 & n1514 ) | ( x502 & n1514 ) ;
  assign n1516 = ( ~n1513 & n1514 ) | ( ~n1513 & n1515 ) | ( n1514 & n1515 ) ;
  assign n1517 = ( x501 & x502 ) | ( x501 & n1513 ) | ( x502 & n1513 ) ;
  assign n1518 = ( x503 & ~x504 ) | ( x503 & n1517 ) | ( ~x504 & n1517 ) ;
  assign n1519 = ( ~x503 & x504 ) | ( ~x503 & n1518 ) | ( x504 & n1518 ) ;
  assign n1520 = ( ~n1517 & n1518 ) | ( ~n1517 & n1519 ) | ( n1518 & n1519 ) ;
  assign n1521 = ( x503 & x504 ) | ( x503 & n1517 ) | ( x504 & n1517 ) ;
  assign n1522 = ( x505 & ~x506 ) | ( x505 & n1521 ) | ( ~x506 & n1521 ) ;
  assign n1523 = ( ~x505 & x506 ) | ( ~x505 & n1522 ) | ( x506 & n1522 ) ;
  assign n1524 = ( ~n1521 & n1522 ) | ( ~n1521 & n1523 ) | ( n1522 & n1523 ) ;
  assign n1525 = ( x505 & x506 ) | ( x505 & n1521 ) | ( x506 & n1521 ) ;
  assign n1526 = ( x507 & ~x508 ) | ( x507 & n1525 ) | ( ~x508 & n1525 ) ;
  assign n1527 = ( ~x507 & x508 ) | ( ~x507 & n1526 ) | ( x508 & n1526 ) ;
  assign n1528 = ( ~n1525 & n1526 ) | ( ~n1525 & n1527 ) | ( n1526 & n1527 ) ;
  assign n1529 = ( x507 & x508 ) | ( x507 & n1525 ) | ( x508 & n1525 ) ;
  assign n1530 = ( x509 & ~x510 ) | ( x509 & n1529 ) | ( ~x510 & n1529 ) ;
  assign n1531 = ( ~x509 & x510 ) | ( ~x509 & n1530 ) | ( x510 & n1530 ) ;
  assign n1532 = ( ~n1529 & n1530 ) | ( ~n1529 & n1531 ) | ( n1530 & n1531 ) ;
  assign n1533 = ( x509 & x510 ) | ( x509 & n1529 ) | ( x510 & n1529 ) ;
  assign n1534 = ( x511 & ~x512 ) | ( x511 & n1533 ) | ( ~x512 & n1533 ) ;
  assign n1535 = ( ~x511 & x512 ) | ( ~x511 & n1534 ) | ( x512 & n1534 ) ;
  assign n1536 = ( ~n1533 & n1534 ) | ( ~n1533 & n1535 ) | ( n1534 & n1535 ) ;
  assign n1537 = ( x511 & x512 ) | ( x511 & n1533 ) | ( x512 & n1533 ) ;
  assign y0 = n516 ;
  assign y1 = n520 ;
  assign y2 = n524 ;
  assign y3 = n528 ;
  assign y4 = n532 ;
  assign y5 = n536 ;
  assign y6 = n540 ;
  assign y7 = n544 ;
  assign y8 = n548 ;
  assign y9 = n552 ;
  assign y10 = n556 ;
  assign y11 = n560 ;
  assign y12 = n564 ;
  assign y13 = n568 ;
  assign y14 = n572 ;
  assign y15 = n576 ;
  assign y16 = n580 ;
  assign y17 = n584 ;
  assign y18 = n588 ;
  assign y19 = n592 ;
  assign y20 = n596 ;
  assign y21 = n600 ;
  assign y22 = n604 ;
  assign y23 = n608 ;
  assign y24 = n612 ;
  assign y25 = n616 ;
  assign y26 = n620 ;
  assign y27 = n624 ;
  assign y28 = n628 ;
  assign y29 = n632 ;
  assign y30 = n636 ;
  assign y31 = n640 ;
  assign y32 = n644 ;
  assign y33 = n648 ;
  assign y34 = n652 ;
  assign y35 = n656 ;
  assign y36 = n660 ;
  assign y37 = n664 ;
  assign y38 = n668 ;
  assign y39 = n672 ;
  assign y40 = n676 ;
  assign y41 = n680 ;
  assign y42 = n684 ;
  assign y43 = n688 ;
  assign y44 = n692 ;
  assign y45 = n696 ;
  assign y46 = n700 ;
  assign y47 = n704 ;
  assign y48 = n708 ;
  assign y49 = n712 ;
  assign y50 = n716 ;
  assign y51 = n720 ;
  assign y52 = n724 ;
  assign y53 = n728 ;
  assign y54 = n732 ;
  assign y55 = n736 ;
  assign y56 = n740 ;
  assign y57 = n744 ;
  assign y58 = n748 ;
  assign y59 = n752 ;
  assign y60 = n756 ;
  assign y61 = n760 ;
  assign y62 = n764 ;
  assign y63 = n768 ;
  assign y64 = n772 ;
  assign y65 = n776 ;
  assign y66 = n780 ;
  assign y67 = n784 ;
  assign y68 = n788 ;
  assign y69 = n792 ;
  assign y70 = n796 ;
  assign y71 = n800 ;
  assign y72 = n804 ;
  assign y73 = n808 ;
  assign y74 = n812 ;
  assign y75 = n816 ;
  assign y76 = n820 ;
  assign y77 = n824 ;
  assign y78 = n828 ;
  assign y79 = n832 ;
  assign y80 = n836 ;
  assign y81 = n840 ;
  assign y82 = n844 ;
  assign y83 = n848 ;
  assign y84 = n852 ;
  assign y85 = n856 ;
  assign y86 = n860 ;
  assign y87 = n864 ;
  assign y88 = n868 ;
  assign y89 = n872 ;
  assign y90 = n876 ;
  assign y91 = n880 ;
  assign y92 = n884 ;
  assign y93 = n888 ;
  assign y94 = n892 ;
  assign y95 = n896 ;
  assign y96 = n900 ;
  assign y97 = n904 ;
  assign y98 = n908 ;
  assign y99 = n912 ;
  assign y100 = n916 ;
  assign y101 = n920 ;
  assign y102 = n924 ;
  assign y103 = n928 ;
  assign y104 = n932 ;
  assign y105 = n936 ;
  assign y106 = n940 ;
  assign y107 = n944 ;
  assign y108 = n948 ;
  assign y109 = n952 ;
  assign y110 = n956 ;
  assign y111 = n960 ;
  assign y112 = n964 ;
  assign y113 = n968 ;
  assign y114 = n972 ;
  assign y115 = n976 ;
  assign y116 = n980 ;
  assign y117 = n984 ;
  assign y118 = n988 ;
  assign y119 = n992 ;
  assign y120 = n996 ;
  assign y121 = n1000 ;
  assign y122 = n1004 ;
  assign y123 = n1008 ;
  assign y124 = n1012 ;
  assign y125 = n1016 ;
  assign y126 = n1020 ;
  assign y127 = n1024 ;
  assign y128 = n1028 ;
  assign y129 = n1032 ;
  assign y130 = n1036 ;
  assign y131 = n1040 ;
  assign y132 = n1044 ;
  assign y133 = n1048 ;
  assign y134 = n1052 ;
  assign y135 = n1056 ;
  assign y136 = n1060 ;
  assign y137 = n1064 ;
  assign y138 = n1068 ;
  assign y139 = n1072 ;
  assign y140 = n1076 ;
  assign y141 = n1080 ;
  assign y142 = n1084 ;
  assign y143 = n1088 ;
  assign y144 = n1092 ;
  assign y145 = n1096 ;
  assign y146 = n1100 ;
  assign y147 = n1104 ;
  assign y148 = n1108 ;
  assign y149 = n1112 ;
  assign y150 = n1116 ;
  assign y151 = n1120 ;
  assign y152 = n1124 ;
  assign y153 = n1128 ;
  assign y154 = n1132 ;
  assign y155 = n1136 ;
  assign y156 = n1140 ;
  assign y157 = n1144 ;
  assign y158 = n1148 ;
  assign y159 = n1152 ;
  assign y160 = n1156 ;
  assign y161 = n1160 ;
  assign y162 = n1164 ;
  assign y163 = n1168 ;
  assign y164 = n1172 ;
  assign y165 = n1176 ;
  assign y166 = n1180 ;
  assign y167 = n1184 ;
  assign y168 = n1188 ;
  assign y169 = n1192 ;
  assign y170 = n1196 ;
  assign y171 = n1200 ;
  assign y172 = n1204 ;
  assign y173 = n1208 ;
  assign y174 = n1212 ;
  assign y175 = n1216 ;
  assign y176 = n1220 ;
  assign y177 = n1224 ;
  assign y178 = n1228 ;
  assign y179 = n1232 ;
  assign y180 = n1236 ;
  assign y181 = n1240 ;
  assign y182 = n1244 ;
  assign y183 = n1248 ;
  assign y184 = n1252 ;
  assign y185 = n1256 ;
  assign y186 = n1260 ;
  assign y187 = n1264 ;
  assign y188 = n1268 ;
  assign y189 = n1272 ;
  assign y190 = n1276 ;
  assign y191 = n1280 ;
  assign y192 = n1284 ;
  assign y193 = n1288 ;
  assign y194 = n1292 ;
  assign y195 = n1296 ;
  assign y196 = n1300 ;
  assign y197 = n1304 ;
  assign y198 = n1308 ;
  assign y199 = n1312 ;
  assign y200 = n1316 ;
  assign y201 = n1320 ;
  assign y202 = n1324 ;
  assign y203 = n1328 ;
  assign y204 = n1332 ;
  assign y205 = n1336 ;
  assign y206 = n1340 ;
  assign y207 = n1344 ;
  assign y208 = n1348 ;
  assign y209 = n1352 ;
  assign y210 = n1356 ;
  assign y211 = n1360 ;
  assign y212 = n1364 ;
  assign y213 = n1368 ;
  assign y214 = n1372 ;
  assign y215 = n1376 ;
  assign y216 = n1380 ;
  assign y217 = n1384 ;
  assign y218 = n1388 ;
  assign y219 = n1392 ;
  assign y220 = n1396 ;
  assign y221 = n1400 ;
  assign y222 = n1404 ;
  assign y223 = n1408 ;
  assign y224 = n1412 ;
  assign y225 = n1416 ;
  assign y226 = n1420 ;
  assign y227 = n1424 ;
  assign y228 = n1428 ;
  assign y229 = n1432 ;
  assign y230 = n1436 ;
  assign y231 = n1440 ;
  assign y232 = n1444 ;
  assign y233 = n1448 ;
  assign y234 = n1452 ;
  assign y235 = n1456 ;
  assign y236 = n1460 ;
  assign y237 = n1464 ;
  assign y238 = n1468 ;
  assign y239 = n1472 ;
  assign y240 = n1476 ;
  assign y241 = n1480 ;
  assign y242 = n1484 ;
  assign y243 = n1488 ;
  assign y244 = n1492 ;
  assign y245 = n1496 ;
  assign y246 = n1500 ;
  assign y247 = n1504 ;
  assign y248 = n1508 ;
  assign y249 = n1512 ;
  assign y250 = n1516 ;
  assign y251 = n1520 ;
  assign y252 = n1524 ;
  assign y253 = n1528 ;
  assign y254 = n1532 ;
  assign y255 = n1536 ;
  assign y256 = n1537 ;
endmodule
