module top( cin , a0 , b0 , a1 , b1 , a2 , b2 , a3 , b3 , a4 , b4 , a5 , b5 , a6 , b6 , a7 , b7 , a8 , b8 , a9 , b9 , a10 , b10 , a11 , b11 , a12 , b12 , a13 , b13 , a14 , b14 , a15 , b15 , a16 , b16 , a17 , b17 , a18 , b18 , a19 , b19 , a20 , b20 , a21 , b21 , a22 , b22 , a23 , b23 , a24 , b24 , a25 , b25 , a26 , b26 , a27 , b27 , a28 , b28 , a29 , b29 , a30 , b30 , a31 , b31 , s0 , s1 , s2 , s3 , s4 , s5 , s6 , s7 , s8 , s9 , s10 , s11 , s12 , s13 , s14 , s15 , s16 , s17 , s18 , s19 , s20 , s21 , s22 , s23 , s24 , s25 , s26 , s27 , s28 , s29 , s30 , s31 , s32 );
  input cin , a0 , b0 , a1 , b1 , a2 , b2 , a3 , b3 , a4 , b4 , a5 , b5 , a6 , b6 , a7 , b7 , a8 , b8 , a9 , b9 , a10 , b10 , a11 , b11 , a12 , b12 , a13 , b13 , a14 , b14 , a15 , b15 , a16 , b16 , a17 , b17 , a18 , b18 , a19 , b19 , a20 , b20 , a21 , b21 , a22 , b22 , a23 , b23 , a24 , b24 , a25 , b25 , a26 , b26 , a27 , b27 , a28 , b28 , a29 , b29 , a30 , b30 , a31 , b31 ;
  output s0 , s1 , s2 , s3 , s4 , s5 , s6 , s7 , s8 , s9 , s10 , s11 , s12 , s13 , s14 , s15 , s16 , s17 , s18 , s19 , s20 , s21 , s22 , s23 , s24 , s25 , s26 , s27 , s28 , s29 , s30 , s31 , s32 ;
  wire n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 ;
  assign n66 = a0 & ~b0 ;
  assign n67 = ~a0 & b0 ;
  assign n68 = n66 | n67 ;
  assign n69 = ~cin & n68 ;
  assign n70 = cin & ~n68 ;
  assign n71 = n69 | n70 ;
  assign n72 = a0 & b0 ;
  assign n73 = cin & a0 ;
  assign n74 = n72 | n73 ;
  assign n75 = cin & b0 ;
  assign n76 = n74 | n75 ;
  assign n77 = a1 & ~b1 ;
  assign n78 = ~a1 & b1 ;
  assign n79 = n77 | n78 ;
  assign n80 = ~n76 & n79 ;
  assign n81 = n76 & ~n79 ;
  assign n82 = n80 | n81 ;
  assign n83 = a1 & b1 ;
  assign n84 = a1 & n76 ;
  assign n85 = n83 | n84 ;
  assign n86 = b1 & n76 ;
  assign n87 = n85 | n86 ;
  assign n88 = a2 & ~b2 ;
  assign n89 = ~a2 & b2 ;
  assign n90 = n88 | n89 ;
  assign n91 = ~n87 & n90 ;
  assign n92 = n87 & ~n90 ;
  assign n93 = n91 | n92 ;
  assign n94 = a2 & b2 ;
  assign n95 = a2 & n87 ;
  assign n96 = n94 | n95 ;
  assign n97 = b2 & n87 ;
  assign n98 = n96 | n97 ;
  assign n99 = a3 & ~b3 ;
  assign n100 = ~a3 & b3 ;
  assign n101 = n99 | n100 ;
  assign n102 = ~n98 & n101 ;
  assign n103 = n98 & ~n101 ;
  assign n104 = n102 | n103 ;
  assign n105 = a3 & b3 ;
  assign n106 = a3 & n98 ;
  assign n107 = n105 | n106 ;
  assign n108 = b3 & n98 ;
  assign n109 = n107 | n108 ;
  assign n110 = a4 & ~b4 ;
  assign n111 = ~a4 & b4 ;
  assign n112 = n110 | n111 ;
  assign n113 = ~n109 & n112 ;
  assign n114 = n109 & ~n112 ;
  assign n115 = n113 | n114 ;
  assign n116 = a4 & b4 ;
  assign n117 = a4 & n109 ;
  assign n118 = n116 | n117 ;
  assign n119 = b4 & n109 ;
  assign n120 = n118 | n119 ;
  assign n121 = a5 & ~b5 ;
  assign n122 = ~a5 & b5 ;
  assign n123 = n121 | n122 ;
  assign n124 = ~n120 & n123 ;
  assign n125 = n120 & ~n123 ;
  assign n126 = n124 | n125 ;
  assign n127 = a5 & b5 ;
  assign n128 = a5 & n120 ;
  assign n129 = n127 | n128 ;
  assign n130 = b5 & n120 ;
  assign n131 = n129 | n130 ;
  assign n132 = a6 & ~b6 ;
  assign n133 = ~a6 & b6 ;
  assign n134 = n132 | n133 ;
  assign n135 = ~n131 & n134 ;
  assign n136 = n131 & ~n134 ;
  assign n137 = n135 | n136 ;
  assign n138 = a6 & b6 ;
  assign n139 = a6 & n131 ;
  assign n140 = n138 | n139 ;
  assign n141 = b6 & n131 ;
  assign n142 = n140 | n141 ;
  assign n143 = a7 & ~b7 ;
  assign n144 = ~a7 & b7 ;
  assign n145 = n143 | n144 ;
  assign n146 = ~n142 & n145 ;
  assign n147 = n142 & ~n145 ;
  assign n148 = n146 | n147 ;
  assign n149 = a7 & b7 ;
  assign n150 = a7 & n142 ;
  assign n151 = n149 | n150 ;
  assign n152 = b7 & n142 ;
  assign n153 = n151 | n152 ;
  assign n154 = a8 & ~b8 ;
  assign n155 = ~a8 & b8 ;
  assign n156 = n154 | n155 ;
  assign n157 = ~n153 & n156 ;
  assign n158 = n153 & ~n156 ;
  assign n159 = n157 | n158 ;
  assign n160 = a8 & b8 ;
  assign n161 = a8 & n153 ;
  assign n162 = n160 | n161 ;
  assign n163 = b8 & n153 ;
  assign n164 = n162 | n163 ;
  assign n165 = a9 & ~b9 ;
  assign n166 = ~a9 & b9 ;
  assign n167 = n165 | n166 ;
  assign n168 = ~n164 & n167 ;
  assign n169 = n164 & ~n167 ;
  assign n170 = n168 | n169 ;
  assign n171 = a9 & b9 ;
  assign n172 = a9 & n164 ;
  assign n173 = n171 | n172 ;
  assign n174 = b9 & n164 ;
  assign n175 = n173 | n174 ;
  assign n176 = a10 & ~b10 ;
  assign n177 = ~a10 & b10 ;
  assign n178 = n176 | n177 ;
  assign n179 = ~n175 & n178 ;
  assign n180 = n175 & ~n178 ;
  assign n181 = n179 | n180 ;
  assign n182 = a10 & b10 ;
  assign n183 = a10 & n175 ;
  assign n184 = n182 | n183 ;
  assign n185 = b10 & n175 ;
  assign n186 = n184 | n185 ;
  assign n187 = a11 & ~b11 ;
  assign n188 = ~a11 & b11 ;
  assign n189 = n187 | n188 ;
  assign n190 = ~n186 & n189 ;
  assign n191 = n186 & ~n189 ;
  assign n192 = n190 | n191 ;
  assign n193 = a11 & b11 ;
  assign n194 = a11 & n186 ;
  assign n195 = n193 | n194 ;
  assign n196 = b11 & n186 ;
  assign n197 = n195 | n196 ;
  assign n198 = a12 & ~b12 ;
  assign n199 = ~a12 & b12 ;
  assign n200 = n198 | n199 ;
  assign n201 = ~n197 & n200 ;
  assign n202 = n197 & ~n200 ;
  assign n203 = n201 | n202 ;
  assign n204 = a12 & b12 ;
  assign n205 = a12 & n197 ;
  assign n206 = n204 | n205 ;
  assign n207 = b12 & n197 ;
  assign n208 = n206 | n207 ;
  assign n209 = a13 & ~b13 ;
  assign n210 = ~a13 & b13 ;
  assign n211 = n209 | n210 ;
  assign n212 = ~n208 & n211 ;
  assign n213 = n208 & ~n211 ;
  assign n214 = n212 | n213 ;
  assign n215 = a13 & b13 ;
  assign n216 = a13 & n208 ;
  assign n217 = n215 | n216 ;
  assign n218 = b13 & n208 ;
  assign n219 = n217 | n218 ;
  assign n220 = a14 & ~b14 ;
  assign n221 = ~a14 & b14 ;
  assign n222 = n220 | n221 ;
  assign n223 = ~n219 & n222 ;
  assign n224 = n219 & ~n222 ;
  assign n225 = n223 | n224 ;
  assign n226 = a14 & b14 ;
  assign n227 = a14 & n219 ;
  assign n228 = n226 | n227 ;
  assign n229 = b14 & n219 ;
  assign n230 = n228 | n229 ;
  assign n231 = a15 & ~b15 ;
  assign n232 = ~a15 & b15 ;
  assign n233 = n231 | n232 ;
  assign n234 = ~n230 & n233 ;
  assign n235 = n230 & ~n233 ;
  assign n236 = n234 | n235 ;
  assign n237 = a15 & b15 ;
  assign n238 = a15 & n230 ;
  assign n239 = n237 | n238 ;
  assign n240 = b15 & n230 ;
  assign n241 = n239 | n240 ;
  assign n242 = a16 & ~b16 ;
  assign n243 = ~a16 & b16 ;
  assign n244 = n242 | n243 ;
  assign n245 = ~n241 & n244 ;
  assign n246 = n241 & ~n244 ;
  assign n247 = n245 | n246 ;
  assign n248 = a16 & b16 ;
  assign n249 = a16 & n241 ;
  assign n250 = n248 | n249 ;
  assign n251 = b16 & n241 ;
  assign n252 = n250 | n251 ;
  assign n253 = a17 & ~b17 ;
  assign n254 = ~a17 & b17 ;
  assign n255 = n253 | n254 ;
  assign n256 = ~n252 & n255 ;
  assign n257 = n252 & ~n255 ;
  assign n258 = n256 | n257 ;
  assign n259 = a17 & b17 ;
  assign n260 = a17 & n252 ;
  assign n261 = n259 | n260 ;
  assign n262 = b17 & n252 ;
  assign n263 = n261 | n262 ;
  assign n264 = a18 & ~b18 ;
  assign n265 = ~a18 & b18 ;
  assign n266 = n264 | n265 ;
  assign n267 = ~n263 & n266 ;
  assign n268 = n263 & ~n266 ;
  assign n269 = n267 | n268 ;
  assign n270 = a18 & b18 ;
  assign n271 = a18 & n263 ;
  assign n272 = n270 | n271 ;
  assign n273 = b18 & n263 ;
  assign n274 = n272 | n273 ;
  assign n275 = a19 & ~b19 ;
  assign n276 = ~a19 & b19 ;
  assign n277 = n275 | n276 ;
  assign n278 = ~n274 & n277 ;
  assign n279 = n274 & ~n277 ;
  assign n280 = n278 | n279 ;
  assign n281 = a19 & b19 ;
  assign n282 = a19 & n274 ;
  assign n283 = n281 | n282 ;
  assign n284 = b19 & n274 ;
  assign n285 = n283 | n284 ;
  assign n286 = a20 & ~b20 ;
  assign n287 = ~a20 & b20 ;
  assign n288 = n286 | n287 ;
  assign n289 = ~n285 & n288 ;
  assign n290 = n285 & ~n288 ;
  assign n291 = n289 | n290 ;
  assign n292 = a20 & b20 ;
  assign n293 = a20 & n285 ;
  assign n294 = n292 | n293 ;
  assign n295 = b20 & n285 ;
  assign n296 = n294 | n295 ;
  assign n297 = a21 & ~b21 ;
  assign n298 = ~a21 & b21 ;
  assign n299 = n297 | n298 ;
  assign n300 = ~n296 & n299 ;
  assign n301 = n296 & ~n299 ;
  assign n302 = n300 | n301 ;
  assign n303 = a21 & b21 ;
  assign n304 = a21 & n296 ;
  assign n305 = n303 | n304 ;
  assign n306 = b21 & n296 ;
  assign n307 = n305 | n306 ;
  assign n308 = a22 & ~b22 ;
  assign n309 = ~a22 & b22 ;
  assign n310 = n308 | n309 ;
  assign n311 = ~n307 & n310 ;
  assign n312 = n307 & ~n310 ;
  assign n313 = n311 | n312 ;
  assign n314 = a22 & b22 ;
  assign n315 = a22 & n307 ;
  assign n316 = n314 | n315 ;
  assign n317 = b22 & n307 ;
  assign n318 = n316 | n317 ;
  assign n319 = a23 & ~b23 ;
  assign n320 = ~a23 & b23 ;
  assign n321 = n319 | n320 ;
  assign n322 = ~n318 & n321 ;
  assign n323 = n318 & ~n321 ;
  assign n324 = n322 | n323 ;
  assign n325 = a23 & b23 ;
  assign n326 = a23 & n318 ;
  assign n327 = n325 | n326 ;
  assign n328 = b23 & n318 ;
  assign n329 = n327 | n328 ;
  assign n330 = a24 & ~b24 ;
  assign n331 = ~a24 & b24 ;
  assign n332 = n330 | n331 ;
  assign n333 = ~n329 & n332 ;
  assign n334 = n329 & ~n332 ;
  assign n335 = n333 | n334 ;
  assign n336 = a24 & b24 ;
  assign n337 = a24 & n329 ;
  assign n338 = n336 | n337 ;
  assign n339 = b24 & n329 ;
  assign n340 = n338 | n339 ;
  assign n341 = a25 & ~b25 ;
  assign n342 = ~a25 & b25 ;
  assign n343 = n341 | n342 ;
  assign n344 = ~n340 & n343 ;
  assign n345 = n340 & ~n343 ;
  assign n346 = n344 | n345 ;
  assign n347 = a25 & b25 ;
  assign n348 = a25 & n340 ;
  assign n349 = n347 | n348 ;
  assign n350 = b25 & n340 ;
  assign n351 = n349 | n350 ;
  assign n352 = a26 & ~b26 ;
  assign n353 = ~a26 & b26 ;
  assign n354 = n352 | n353 ;
  assign n355 = ~n351 & n354 ;
  assign n356 = n351 & ~n354 ;
  assign n357 = n355 | n356 ;
  assign n358 = a26 & b26 ;
  assign n359 = a26 & n351 ;
  assign n360 = n358 | n359 ;
  assign n361 = b26 & n351 ;
  assign n362 = n360 | n361 ;
  assign n363 = a27 & ~b27 ;
  assign n364 = ~a27 & b27 ;
  assign n365 = n363 | n364 ;
  assign n366 = ~n362 & n365 ;
  assign n367 = n362 & ~n365 ;
  assign n368 = n366 | n367 ;
  assign n369 = a27 & b27 ;
  assign n370 = a27 & n362 ;
  assign n371 = n369 | n370 ;
  assign n372 = b27 & n362 ;
  assign n373 = n371 | n372 ;
  assign n374 = a28 & ~b28 ;
  assign n375 = ~a28 & b28 ;
  assign n376 = n374 | n375 ;
  assign n377 = ~n373 & n376 ;
  assign n378 = n373 & ~n376 ;
  assign n379 = n377 | n378 ;
  assign n380 = a28 & b28 ;
  assign n381 = a28 & n373 ;
  assign n382 = n380 | n381 ;
  assign n383 = b28 & n373 ;
  assign n384 = n382 | n383 ;
  assign n385 = a29 & ~b29 ;
  assign n386 = ~a29 & b29 ;
  assign n387 = n385 | n386 ;
  assign n388 = ~n384 & n387 ;
  assign n389 = n384 & ~n387 ;
  assign n390 = n388 | n389 ;
  assign n391 = a29 & b29 ;
  assign n392 = a29 & n384 ;
  assign n393 = n391 | n392 ;
  assign n394 = b29 & n384 ;
  assign n395 = n393 | n394 ;
  assign n396 = a30 & ~b30 ;
  assign n397 = ~a30 & b30 ;
  assign n398 = n396 | n397 ;
  assign n399 = ~n395 & n398 ;
  assign n400 = n395 & ~n398 ;
  assign n401 = n399 | n400 ;
  assign n402 = a30 & b30 ;
  assign n403 = a30 & n395 ;
  assign n404 = n402 | n403 ;
  assign n405 = b30 & n395 ;
  assign n406 = n404 | n405 ;
  assign n407 = a31 & ~b31 ;
  assign n408 = ~a31 & b31 ;
  assign n409 = n407 | n408 ;
  assign n410 = ~n406 & n409 ;
  assign n411 = n406 & ~n409 ;
  assign n412 = n410 | n411 ;
  assign n413 = a31 & b31 ;
  assign n414 = a31 & n406 ;
  assign n415 = n413 | n414 ;
  assign n416 = b31 & n406 ;
  assign n417 = n415 | n416 ;
  assign s0 = n71 ;
  assign s1 = n82 ;
  assign s2 = n93 ;
  assign s3 = n104 ;
  assign s4 = n115 ;
  assign s5 = n126 ;
  assign s6 = n137 ;
  assign s7 = n148 ;
  assign s8 = n159 ;
  assign s9 = n170 ;
  assign s10 = n181 ;
  assign s11 = n192 ;
  assign s12 = n203 ;
  assign s13 = n214 ;
  assign s14 = n225 ;
  assign s15 = n236 ;
  assign s16 = n247 ;
  assign s17 = n258 ;
  assign s18 = n269 ;
  assign s19 = n280 ;
  assign s20 = n291 ;
  assign s21 = n302 ;
  assign s22 = n313 ;
  assign s23 = n324 ;
  assign s24 = n335 ;
  assign s25 = n346 ;
  assign s26 = n357 ;
  assign s27 = n368 ;
  assign s28 = n379 ;
  assign s29 = n390 ;
  assign s30 = n401 ;
  assign s31 = n412 ;
  assign s32 = n417 ;
endmodule
