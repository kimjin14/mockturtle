module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 ;
  wire n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 ;
  assign n66 = ( x0 & ~x1 ) | ( x0 & x2 ) | ( ~x1 & x2 ) ;
  assign n67 = ( ~x0 & x1 ) | ( ~x0 & n66 ) | ( x1 & n66 ) ;
  assign n68 = ( ~x2 & n66 ) | ( ~x2 & n67 ) | ( n66 & n67 ) ;
  assign n69 = ( x0 & x1 ) | ( x0 & x2 ) | ( x1 & x2 ) ;
  assign n70 = ( x3 & ~x4 ) | ( x3 & n69 ) | ( ~x4 & n69 ) ;
  assign n71 = ( ~x3 & x4 ) | ( ~x3 & n70 ) | ( x4 & n70 ) ;
  assign n72 = ( ~n69 & n70 ) | ( ~n69 & n71 ) | ( n70 & n71 ) ;
  assign n73 = ( x3 & x4 ) | ( x3 & n69 ) | ( x4 & n69 ) ;
  assign n74 = ( x5 & ~x6 ) | ( x5 & n73 ) | ( ~x6 & n73 ) ;
  assign n75 = ( ~x5 & x6 ) | ( ~x5 & n74 ) | ( x6 & n74 ) ;
  assign n76 = ( ~n73 & n74 ) | ( ~n73 & n75 ) | ( n74 & n75 ) ;
  assign n77 = ( x4 & x5 ) | ( x4 & x6 ) | ( x5 & x6 ) ;
  assign n78 = ( x3 & x5 ) | ( x3 & x6 ) | ( x5 & x6 ) ;
  assign n79 = ( n69 & n77 ) | ( n69 & n78 ) | ( n77 & n78 ) ;
  assign n80 = ( x7 & ~x8 ) | ( x7 & n79 ) | ( ~x8 & n79 ) ;
  assign n81 = ( ~x7 & x8 ) | ( ~x7 & n80 ) | ( x8 & n80 ) ;
  assign n82 = ( ~n79 & n80 ) | ( ~n79 & n81 ) | ( n80 & n81 ) ;
  assign n83 = ( x7 & x8 ) | ( x7 & n79 ) | ( x8 & n79 ) ;
  assign n84 = ( x9 & ~x10 ) | ( x9 & n83 ) | ( ~x10 & n83 ) ;
  assign n85 = ( ~x9 & x10 ) | ( ~x9 & n84 ) | ( x10 & n84 ) ;
  assign n86 = ( ~n83 & n84 ) | ( ~n83 & n85 ) | ( n84 & n85 ) ;
  assign n87 = ( x8 & x9 ) | ( x8 & x10 ) | ( x9 & x10 ) ;
  assign n88 = ( x7 & x9 ) | ( x7 & x10 ) | ( x9 & x10 ) ;
  assign n89 = ( n79 & n87 ) | ( n79 & n88 ) | ( n87 & n88 ) ;
  assign n90 = ( x11 & ~x12 ) | ( x11 & n89 ) | ( ~x12 & n89 ) ;
  assign n91 = ( ~x11 & x12 ) | ( ~x11 & n90 ) | ( x12 & n90 ) ;
  assign n92 = ( ~n89 & n90 ) | ( ~n89 & n91 ) | ( n90 & n91 ) ;
  assign n93 = ( x11 & x12 ) | ( x11 & n88 ) | ( x12 & n88 ) ;
  assign n94 = ( x11 & x12 ) | ( x11 & n87 ) | ( x12 & n87 ) ;
  assign n95 = ( n79 & n93 ) | ( n79 & n94 ) | ( n93 & n94 ) ;
  assign n96 = ( x13 & ~x14 ) | ( x13 & n95 ) | ( ~x14 & n95 ) ;
  assign n97 = ( ~x13 & x14 ) | ( ~x13 & n96 ) | ( x14 & n96 ) ;
  assign n98 = ( ~n95 & n96 ) | ( ~n95 & n97 ) | ( n96 & n97 ) ;
  assign n99 = ( x13 & x14 ) | ( x13 & n95 ) | ( x14 & n95 ) ;
  assign n100 = ( x15 & ~x16 ) | ( x15 & n99 ) | ( ~x16 & n99 ) ;
  assign n101 = ( ~x15 & x16 ) | ( ~x15 & n100 ) | ( x16 & n100 ) ;
  assign n102 = ( ~n99 & n100 ) | ( ~n99 & n101 ) | ( n100 & n101 ) ;
  assign n103 = ( x14 & x15 ) | ( x14 & x16 ) | ( x15 & x16 ) ;
  assign n104 = ( x13 & x15 ) | ( x13 & x16 ) | ( x15 & x16 ) ;
  assign n105 = ( n95 & n103 ) | ( n95 & n104 ) | ( n103 & n104 ) ;
  assign n106 = ( x17 & ~x18 ) | ( x17 & n105 ) | ( ~x18 & n105 ) ;
  assign n107 = ( ~x17 & x18 ) | ( ~x17 & n106 ) | ( x18 & n106 ) ;
  assign n108 = ( ~n105 & n106 ) | ( ~n105 & n107 ) | ( n106 & n107 ) ;
  assign n109 = ( x17 & x18 ) | ( x17 & n104 ) | ( x18 & n104 ) ;
  assign n110 = ( x17 & x18 ) | ( x17 & n103 ) | ( x18 & n103 ) ;
  assign n111 = ( n95 & n109 ) | ( n95 & n110 ) | ( n109 & n110 ) ;
  assign n112 = ( x19 & ~x20 ) | ( x19 & n111 ) | ( ~x20 & n111 ) ;
  assign n113 = ( ~x19 & x20 ) | ( ~x19 & n112 ) | ( x20 & n112 ) ;
  assign n114 = ( ~n111 & n112 ) | ( ~n111 & n113 ) | ( n112 & n113 ) ;
  assign n115 = ( x19 & x20 ) | ( x19 & n110 ) | ( x20 & n110 ) ;
  assign n116 = ( x19 & x20 ) | ( x19 & n109 ) | ( x20 & n109 ) ;
  assign n117 = ( n95 & n115 ) | ( n95 & n116 ) | ( n115 & n116 ) ;
  assign n118 = ( x21 & ~x22 ) | ( x21 & n117 ) | ( ~x22 & n117 ) ;
  assign n119 = ( ~x21 & x22 ) | ( ~x21 & n118 ) | ( x22 & n118 ) ;
  assign n120 = ( ~n117 & n118 ) | ( ~n117 & n119 ) | ( n118 & n119 ) ;
  assign n121 = ( x21 & x22 ) | ( x21 & n117 ) | ( x22 & n117 ) ;
  assign n122 = ( x23 & ~x24 ) | ( x23 & n121 ) | ( ~x24 & n121 ) ;
  assign n123 = ( ~x23 & x24 ) | ( ~x23 & n122 ) | ( x24 & n122 ) ;
  assign n124 = ( ~n121 & n122 ) | ( ~n121 & n123 ) | ( n122 & n123 ) ;
  assign n125 = ( x22 & x23 ) | ( x22 & x24 ) | ( x23 & x24 ) ;
  assign n126 = ( x21 & x23 ) | ( x21 & x24 ) | ( x23 & x24 ) ;
  assign n127 = ( n117 & n125 ) | ( n117 & n126 ) | ( n125 & n126 ) ;
  assign n128 = ( x25 & ~x26 ) | ( x25 & n127 ) | ( ~x26 & n127 ) ;
  assign n129 = ( ~x25 & x26 ) | ( ~x25 & n128 ) | ( x26 & n128 ) ;
  assign n130 = ( ~n127 & n128 ) | ( ~n127 & n129 ) | ( n128 & n129 ) ;
  assign n131 = ( x25 & x26 ) | ( x25 & n126 ) | ( x26 & n126 ) ;
  assign n132 = ( x25 & x26 ) | ( x25 & n125 ) | ( x26 & n125 ) ;
  assign n133 = ( n117 & n131 ) | ( n117 & n132 ) | ( n131 & n132 ) ;
  assign n134 = ( x27 & ~x28 ) | ( x27 & n133 ) | ( ~x28 & n133 ) ;
  assign n135 = ( ~x27 & x28 ) | ( ~x27 & n134 ) | ( x28 & n134 ) ;
  assign n136 = ( ~n133 & n134 ) | ( ~n133 & n135 ) | ( n134 & n135 ) ;
  assign n137 = ( x27 & x28 ) | ( x27 & n132 ) | ( x28 & n132 ) ;
  assign n138 = ( x27 & x28 ) | ( x27 & n131 ) | ( x28 & n131 ) ;
  assign n139 = ( n117 & n137 ) | ( n117 & n138 ) | ( n137 & n138 ) ;
  assign n140 = ( x29 & ~x30 ) | ( x29 & n139 ) | ( ~x30 & n139 ) ;
  assign n141 = ( ~x29 & x30 ) | ( ~x29 & n140 ) | ( x30 & n140 ) ;
  assign n142 = ( ~n139 & n140 ) | ( ~n139 & n141 ) | ( n140 & n141 ) ;
  assign n143 = ( x29 & x30 ) | ( x29 & n138 ) | ( x30 & n138 ) ;
  assign n144 = ( x29 & x30 ) | ( x29 & n137 ) | ( x30 & n137 ) ;
  assign n145 = ( n117 & n143 ) | ( n117 & n144 ) | ( n143 & n144 ) ;
  assign n146 = ( x31 & ~x32 ) | ( x31 & n145 ) | ( ~x32 & n145 ) ;
  assign n147 = ( ~x31 & x32 ) | ( ~x31 & n146 ) | ( x32 & n146 ) ;
  assign n148 = ( ~n145 & n146 ) | ( ~n145 & n147 ) | ( n146 & n147 ) ;
  assign n149 = ( x31 & x32 ) | ( x31 & n145 ) | ( x32 & n145 ) ;
  assign n150 = ( x33 & ~x34 ) | ( x33 & n149 ) | ( ~x34 & n149 ) ;
  assign n151 = ( ~x33 & x34 ) | ( ~x33 & n150 ) | ( x34 & n150 ) ;
  assign n152 = ( ~n149 & n150 ) | ( ~n149 & n151 ) | ( n150 & n151 ) ;
  assign n153 = ( x32 & x33 ) | ( x32 & x34 ) | ( x33 & x34 ) ;
  assign n154 = ( x31 & x33 ) | ( x31 & x34 ) | ( x33 & x34 ) ;
  assign n155 = ( n145 & n153 ) | ( n145 & n154 ) | ( n153 & n154 ) ;
  assign n156 = ( x35 & ~x36 ) | ( x35 & n155 ) | ( ~x36 & n155 ) ;
  assign n157 = ( ~x35 & x36 ) | ( ~x35 & n156 ) | ( x36 & n156 ) ;
  assign n158 = ( ~n155 & n156 ) | ( ~n155 & n157 ) | ( n156 & n157 ) ;
  assign n159 = ( x35 & x36 ) | ( x35 & n154 ) | ( x36 & n154 ) ;
  assign n160 = ( x35 & x36 ) | ( x35 & n153 ) | ( x36 & n153 ) ;
  assign n161 = ( n145 & n159 ) | ( n145 & n160 ) | ( n159 & n160 ) ;
  assign n162 = ( x37 & ~x38 ) | ( x37 & n161 ) | ( ~x38 & n161 ) ;
  assign n163 = ( ~x37 & x38 ) | ( ~x37 & n162 ) | ( x38 & n162 ) ;
  assign n164 = ( ~n161 & n162 ) | ( ~n161 & n163 ) | ( n162 & n163 ) ;
  assign n165 = ( x37 & x38 ) | ( x37 & n160 ) | ( x38 & n160 ) ;
  assign n166 = ( x37 & x38 ) | ( x37 & n159 ) | ( x38 & n159 ) ;
  assign n167 = ( n145 & n165 ) | ( n145 & n166 ) | ( n165 & n166 ) ;
  assign n168 = ( x39 & ~x40 ) | ( x39 & n167 ) | ( ~x40 & n167 ) ;
  assign n169 = ( ~x39 & x40 ) | ( ~x39 & n168 ) | ( x40 & n168 ) ;
  assign n170 = ( ~n167 & n168 ) | ( ~n167 & n169 ) | ( n168 & n169 ) ;
  assign n171 = ( x39 & x40 ) | ( x39 & n166 ) | ( x40 & n166 ) ;
  assign n172 = ( x39 & x40 ) | ( x39 & n165 ) | ( x40 & n165 ) ;
  assign n173 = ( n145 & n171 ) | ( n145 & n172 ) | ( n171 & n172 ) ;
  assign n174 = ( x41 & ~x42 ) | ( x41 & n173 ) | ( ~x42 & n173 ) ;
  assign n175 = ( ~x41 & x42 ) | ( ~x41 & n174 ) | ( x42 & n174 ) ;
  assign n176 = ( ~n173 & n174 ) | ( ~n173 & n175 ) | ( n174 & n175 ) ;
  assign n177 = ( x41 & x42 ) | ( x41 & n172 ) | ( x42 & n172 ) ;
  assign n178 = ( x41 & x42 ) | ( x41 & n171 ) | ( x42 & n171 ) ;
  assign n179 = ( n145 & n177 ) | ( n145 & n178 ) | ( n177 & n178 ) ;
  assign n180 = ( x43 & ~x44 ) | ( x43 & n179 ) | ( ~x44 & n179 ) ;
  assign n181 = ( ~x43 & x44 ) | ( ~x43 & n180 ) | ( x44 & n180 ) ;
  assign n182 = ( ~n179 & n180 ) | ( ~n179 & n181 ) | ( n180 & n181 ) ;
  assign n183 = ( x43 & x44 ) | ( x43 & n179 ) | ( x44 & n179 ) ;
  assign n184 = ( x45 & ~x46 ) | ( x45 & n183 ) | ( ~x46 & n183 ) ;
  assign n185 = ( ~x45 & x46 ) | ( ~x45 & n184 ) | ( x46 & n184 ) ;
  assign n186 = ( ~n183 & n184 ) | ( ~n183 & n185 ) | ( n184 & n185 ) ;
  assign n187 = ( x44 & x45 ) | ( x44 & x46 ) | ( x45 & x46 ) ;
  assign n188 = ( x43 & x45 ) | ( x43 & x46 ) | ( x45 & x46 ) ;
  assign n189 = ( n179 & n187 ) | ( n179 & n188 ) | ( n187 & n188 ) ;
  assign n190 = ( x47 & ~x48 ) | ( x47 & n189 ) | ( ~x48 & n189 ) ;
  assign n191 = ( ~x47 & x48 ) | ( ~x47 & n190 ) | ( x48 & n190 ) ;
  assign n192 = ( ~n189 & n190 ) | ( ~n189 & n191 ) | ( n190 & n191 ) ;
  assign n193 = ( x47 & x48 ) | ( x47 & n188 ) | ( x48 & n188 ) ;
  assign n194 = ( x47 & x48 ) | ( x47 & n187 ) | ( x48 & n187 ) ;
  assign n195 = ( n179 & n193 ) | ( n179 & n194 ) | ( n193 & n194 ) ;
  assign n196 = ( x49 & ~x50 ) | ( x49 & n195 ) | ( ~x50 & n195 ) ;
  assign n197 = ( ~x49 & x50 ) | ( ~x49 & n196 ) | ( x50 & n196 ) ;
  assign n198 = ( ~n195 & n196 ) | ( ~n195 & n197 ) | ( n196 & n197 ) ;
  assign n199 = ( x49 & x50 ) | ( x49 & n194 ) | ( x50 & n194 ) ;
  assign n200 = ( x49 & x50 ) | ( x49 & n193 ) | ( x50 & n193 ) ;
  assign n201 = ( n179 & n199 ) | ( n179 & n200 ) | ( n199 & n200 ) ;
  assign n202 = ( x51 & ~x52 ) | ( x51 & n201 ) | ( ~x52 & n201 ) ;
  assign n203 = ( ~x51 & x52 ) | ( ~x51 & n202 ) | ( x52 & n202 ) ;
  assign n204 = ( ~n201 & n202 ) | ( ~n201 & n203 ) | ( n202 & n203 ) ;
  assign n205 = ( x51 & x52 ) | ( x51 & n200 ) | ( x52 & n200 ) ;
  assign n206 = ( x51 & x52 ) | ( x51 & n199 ) | ( x52 & n199 ) ;
  assign n207 = ( n179 & n205 ) | ( n179 & n206 ) | ( n205 & n206 ) ;
  assign n208 = ( x53 & ~x54 ) | ( x53 & n207 ) | ( ~x54 & n207 ) ;
  assign n209 = ( ~x53 & x54 ) | ( ~x53 & n208 ) | ( x54 & n208 ) ;
  assign n210 = ( ~n207 & n208 ) | ( ~n207 & n209 ) | ( n208 & n209 ) ;
  assign n211 = ( x53 & x54 ) | ( x53 & n206 ) | ( x54 & n206 ) ;
  assign n212 = ( x53 & x54 ) | ( x53 & n205 ) | ( x54 & n205 ) ;
  assign n213 = ( n179 & n211 ) | ( n179 & n212 ) | ( n211 & n212 ) ;
  assign n214 = ( x55 & ~x56 ) | ( x55 & n213 ) | ( ~x56 & n213 ) ;
  assign n215 = ( ~x55 & x56 ) | ( ~x55 & n214 ) | ( x56 & n214 ) ;
  assign n216 = ( ~n213 & n214 ) | ( ~n213 & n215 ) | ( n214 & n215 ) ;
  assign n217 = ( x55 & x56 ) | ( x55 & n212 ) | ( x56 & n212 ) ;
  assign n218 = ( x55 & x56 ) | ( x55 & n211 ) | ( x56 & n211 ) ;
  assign n219 = ( n179 & n217 ) | ( n179 & n218 ) | ( n217 & n218 ) ;
  assign n220 = ( x57 & ~x58 ) | ( x57 & n219 ) | ( ~x58 & n219 ) ;
  assign n221 = ( ~x57 & x58 ) | ( ~x57 & n220 ) | ( x58 & n220 ) ;
  assign n222 = ( ~n219 & n220 ) | ( ~n219 & n221 ) | ( n220 & n221 ) ;
  assign n223 = ( x57 & x58 ) | ( x57 & n219 ) | ( x58 & n219 ) ;
  assign n224 = ( x59 & ~x60 ) | ( x59 & n223 ) | ( ~x60 & n223 ) ;
  assign n225 = ( ~x59 & x60 ) | ( ~x59 & n224 ) | ( x60 & n224 ) ;
  assign n226 = ( ~n223 & n224 ) | ( ~n223 & n225 ) | ( n224 & n225 ) ;
  assign n227 = ( x58 & x59 ) | ( x58 & x60 ) | ( x59 & x60 ) ;
  assign n228 = ( x57 & x59 ) | ( x57 & x60 ) | ( x59 & x60 ) ;
  assign n229 = ( n219 & n227 ) | ( n219 & n228 ) | ( n227 & n228 ) ;
  assign n230 = ( x61 & ~x62 ) | ( x61 & n229 ) | ( ~x62 & n229 ) ;
  assign n231 = ( ~x61 & x62 ) | ( ~x61 & n230 ) | ( x62 & n230 ) ;
  assign n232 = ( ~n229 & n230 ) | ( ~n229 & n231 ) | ( n230 & n231 ) ;
  assign n233 = ( x61 & x62 ) | ( x61 & n228 ) | ( x62 & n228 ) ;
  assign n234 = ( x61 & x62 ) | ( x61 & n227 ) | ( x62 & n227 ) ;
  assign n235 = ( n219 & n233 ) | ( n219 & n234 ) | ( n233 & n234 ) ;
  assign n236 = ( x63 & ~x64 ) | ( x63 & n234 ) | ( ~x64 & n234 ) ;
  assign n237 = ( x63 & ~x64 ) | ( x63 & n233 ) | ( ~x64 & n233 ) ;
  assign n238 = ( n219 & n236 ) | ( n219 & n237 ) | ( n236 & n237 ) ;
  assign n239 = ( ~x63 & x64 ) | ( ~x63 & n237 ) | ( x64 & n237 ) ;
  assign n240 = ( ~x63 & x64 ) | ( ~x63 & n236 ) | ( x64 & n236 ) ;
  assign n241 = ( n219 & n239 ) | ( n219 & n240 ) | ( n239 & n240 ) ;
  assign n242 = ( ~n235 & n238 ) | ( ~n235 & n241 ) | ( n238 & n241 ) ;
  assign n243 = ( x63 & x64 ) | ( x63 & n235 ) | ( x64 & n235 ) ;
  assign y0 = n68 ;
  assign y1 = n72 ;
  assign y2 = n76 ;
  assign y3 = n82 ;
  assign y4 = n86 ;
  assign y5 = n92 ;
  assign y6 = n98 ;
  assign y7 = n102 ;
  assign y8 = n108 ;
  assign y9 = n114 ;
  assign y10 = n120 ;
  assign y11 = n124 ;
  assign y12 = n130 ;
  assign y13 = n136 ;
  assign y14 = n142 ;
  assign y15 = n148 ;
  assign y16 = n152 ;
  assign y17 = n158 ;
  assign y18 = n164 ;
  assign y19 = n170 ;
  assign y20 = n176 ;
  assign y21 = n182 ;
  assign y22 = n186 ;
  assign y23 = n192 ;
  assign y24 = n198 ;
  assign y25 = n204 ;
  assign y26 = n210 ;
  assign y27 = n216 ;
  assign y28 = n222 ;
  assign y29 = n226 ;
  assign y30 = n232 ;
  assign y31 = n242 ;
  assign y32 = n243 ;
endmodule
