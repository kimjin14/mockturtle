module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 , x147 , x148 , x149 , x150 , x151 , x152 , x153 , x154 , x155 , x156 , x157 , x158 , x159 , x160 , x161 , x162 , x163 , x164 , x165 , x166 , x167 , x168 , x169 , x170 , x171 , x172 , x173 , x174 , x175 , x176 , x177 , x178 , x179 , x180 , x181 , x182 , x183 , x184 , x185 , x186 , x187 , x188 , x189 , x190 , x191 , x192 , x193 , x194 , x195 , x196 , x197 , x198 , x199 , x200 , x201 , x202 , x203 , x204 , x205 , x206 , x207 , x208 , x209 , x210 , x211 , x212 , x213 , x214 , x215 , x216 , x217 , x218 , x219 , x220 , x221 , x222 , x223 , x224 , x225 , x226 , x227 , x228 , x229 , x230 , x231 , x232 , x233 , x234 , x235 , x236 , x237 , x238 , x239 , x240 , x241 , x242 , x243 , x244 , x245 , x246 , x247 , x248 , x249 , x250 , x251 , x252 , x253 , x254 , x255 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 , y128 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 , x147 , x148 , x149 , x150 , x151 , x152 , x153 , x154 , x155 , x156 , x157 , x158 , x159 , x160 , x161 , x162 , x163 , x164 , x165 , x166 , x167 , x168 , x169 , x170 , x171 , x172 , x173 , x174 , x175 , x176 , x177 , x178 , x179 , x180 , x181 , x182 , x183 , x184 , x185 , x186 , x187 , x188 , x189 , x190 , x191 , x192 , x193 , x194 , x195 , x196 , x197 , x198 , x199 , x200 , x201 , x202 , x203 , x204 , x205 , x206 , x207 , x208 , x209 , x210 , x211 , x212 , x213 , x214 , x215 , x216 , x217 , x218 , x219 , x220 , x221 , x222 , x223 , x224 , x225 , x226 , x227 , x228 , x229 , x230 , x231 , x232 , x233 , x234 , x235 , x236 , x237 , x238 , x239 , x240 , x241 , x242 , x243 , x244 , x245 , x246 , x247 , x248 , x249 , x250 , x251 , x252 , x253 , x254 , x255 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 , y128 ;
  wire n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , n3931 , n3932 , n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , n3940 , n3941 , n3942 , n3943 , n3944 , n3945 , n3946 , n3947 , n3948 , n3949 , n3950 , n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , n3970 , n3971 , n3972 , n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , n3980 , n3981 , n3982 , n3983 , n3984 , n3985 , n3986 , n3987 , n3988 , n3989 , n3990 , n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , n4000 , n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , n4009 , n4010 , n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , n4019 , n4020 , n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , n4029 , n4030 , n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , n4039 , n4040 , n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4049 , n4050 , n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , n4059 , n4060 , n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , n4070 , n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , n4079 , n4080 , n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , n4089 , n4090 , n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , n4097 , n4098 , n4099 , n4100 , n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , n4109 , n4110 , n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , n4119 , n4120 , n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , n4129 , n4130 , n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , n4139 , n4140 , n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , n4150 , n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , n4159 , n4160 , n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , n4169 , n4170 , n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , n4179 , n4180 , n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , n4189 , n4190 , n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , n4197 , n4198 , n4199 , n4200 , n4201 , n4202 , n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , n4209 , n4210 , n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , n4217 , n4218 , n4219 , n4220 , n4221 , n4222 , n4223 , n4224 , n4225 , n4226 , n4227 , n4228 , n4229 , n4230 , n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , n4237 , n4238 , n4239 , n4240 , n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , n4247 , n4248 , n4249 , n4250 , n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , n4259 , n4260 , n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , n4269 , n4270 , n4271 , n4272 , n4273 , n4274 , n4275 , n4276 , n4277 , n4278 , n4279 , n4280 , n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , n4289 , n4290 , n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , n4299 , n4300 , n4301 , n4302 , n4303 , n4304 , n4305 , n4306 , n4307 , n4308 , n4309 , n4310 , n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , n4319 , n4320 , n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , n4329 , n4330 , n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , n4340 , n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , n4349 , n4350 , n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , n4360 , n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , n4370 , n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , n4380 , n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , n4390 , n4391 , n4392 , n4393 , n4394 , n4395 , n4396 , n4397 , n4398 , n4399 , n4400 , n4401 , n4402 , n4403 , n4404 , n4405 , n4406 , n4407 , n4408 , n4409 , n4410 , n4411 , n4412 , n4413 , n4414 , n4415 , n4416 , n4417 , n4418 , n4419 , n4420 , n4421 , n4422 , n4423 , n4424 , n4425 , n4426 , n4427 , n4428 , n4429 , n4430 , n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , n4437 , n4438 , n4439 , n4440 , n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , n4449 , n4450 , n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , n4459 , n4460 , n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , n4469 , n4470 , n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , n4479 , n4480 , n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , n4487 , n4488 , n4489 , n4490 , n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , n4497 , n4498 , n4499 , n4500 , n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , n4509 , n4510 , n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , n4519 , n4520 , n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , n4529 , n4530 , n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , n4537 , n4538 , n4539 , n4540 , n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , n4547 , n4548 , n4549 , n4550 , n4551 , n4552 , n4553 , n4554 , n4555 , n4556 , n4557 , n4558 , n4559 , n4560 , n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , n4567 , n4568 , n4569 , n4570 , n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , n4579 , n4580 , n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , n4589 , n4590 , n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , n4597 , n4598 , n4599 , n4600 , n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , n4607 , n4608 , n4609 , n4610 , n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , n4617 , n4618 , n4619 , n4620 , n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , n4627 , n4628 , n4629 , n4630 , n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , n4637 , n4638 , n4639 , n4640 , n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , n4647 , n4648 , n4649 , n4650 , n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , n4657 , n4658 , n4659 , n4660 , n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , n4669 , n4670 , n4671 , n4672 , n4673 , n4674 , n4675 , n4676 , n4677 , n4678 , n4679 , n4680 , n4681 , n4682 , n4683 , n4684 , n4685 , n4686 , n4687 , n4688 , n4689 , n4690 , n4691 , n4692 , n4693 , n4694 , n4695 , n4696 , n4697 , n4698 , n4699 , n4700 , n4701 , n4702 , n4703 , n4704 , n4705 , n4706 , n4707 , n4708 , n4709 , n4710 , n4711 , n4712 , n4713 , n4714 , n4715 , n4716 , n4717 , n4718 , n4719 , n4720 , n4721 , n4722 , n4723 , n4724 , n4725 , n4726 , n4727 , n4728 , n4729 , n4730 , n4731 , n4732 , n4733 , n4734 , n4735 , n4736 , n4737 , n4738 , n4739 , n4740 , n4741 , n4742 , n4743 , n4744 , n4745 , n4746 , n4747 , n4748 , n4749 , n4750 , n4751 , n4752 , n4753 , n4754 , n4755 , n4756 , n4757 , n4758 , n4759 , n4760 , n4761 , n4762 , n4763 , n4764 , n4765 , n4766 , n4767 , n4768 , n4769 , n4770 , n4771 , n4772 , n4773 , n4774 , n4775 , n4776 , n4777 , n4778 , n4779 , n4780 , n4781 , n4782 , n4783 , n4784 , n4785 , n4786 , n4787 , n4788 , n4789 , n4790 , n4791 , n4792 , n4793 , n4794 , n4795 , n4796 , n4797 , n4798 , n4799 , n4800 , n4801 , n4802 , n4803 , n4804 , n4805 , n4806 , n4807 , n4808 , n4809 , n4810 , n4811 , n4812 , n4813 , n4814 , n4815 , n4816 , n4817 , n4818 , n4819 , n4820 , n4821 , n4822 , n4823 , n4824 , n4825 , n4826 , n4827 , n4828 , n4829 , n4830 , n4831 , n4832 , n4833 , n4834 , n4835 , n4836 , n4837 , n4838 , n4839 , n4840 , n4841 , n4842 , n4843 , n4844 , n4845 , n4846 , n4847 , n4848 , n4849 , n4850 , n4851 , n4852 , n4853 , n4854 , n4855 , n4856 , n4857 , n4858 , n4859 , n4860 , n4861 , n4862 , n4863 , n4864 , n4865 , n4866 , n4867 , n4868 , n4869 , n4870 , n4871 , n4872 , n4873 , n4874 , n4875 , n4876 , n4877 , n4878 , n4879 , n4880 , n4881 , n4882 , n4883 , n4884 , n4885 , n4886 , n4887 , n4888 , n4889 , n4890 , n4891 , n4892 , n4893 , n4894 , n4895 , n4896 , n4897 , n4898 , n4899 , n4900 , n4901 , n4902 , n4903 , n4904 , n4905 , n4906 , n4907 , n4908 , n4909 , n4910 , n4911 , n4912 , n4913 , n4914 , n4915 , n4916 , n4917 , n4918 , n4919 , n4920 , n4921 , n4922 , n4923 , n4924 , n4925 , n4926 , n4927 , n4928 , n4929 , n4930 , n4931 , n4932 , n4933 , n4934 , n4935 , n4936 , n4937 , n4938 , n4939 , n4940 , n4941 , n4942 , n4943 , n4944 , n4945 , n4946 , n4947 , n4948 , n4949 , n4950 , n4951 , n4952 , n4953 , n4954 , n4955 , n4956 , n4957 , n4958 , n4959 , n4960 , n4961 , n4962 , n4963 , n4964 , n4965 , n4966 , n4967 , n4968 , n4969 , n4970 , n4971 , n4972 , n4973 , n4974 , n4975 , n4976 , n4977 , n4978 , n4979 , n4980 , n4981 , n4982 , n4983 , n4984 , n4985 , n4986 , n4987 , n4988 , n4989 , n4990 , n4991 , n4992 , n4993 , n4994 , n4995 , n4996 , n4997 , n4998 , n4999 , n5000 , n5001 , n5002 , n5003 , n5004 , n5005 , n5006 , n5007 , n5008 , n5009 , n5010 , n5011 , n5012 , n5013 , n5014 , n5015 , n5016 , n5017 , n5018 , n5019 , n5020 , n5021 , n5022 , n5023 , n5024 , n5025 , n5026 , n5027 , n5028 , n5029 , n5030 , n5031 , n5032 , n5033 , n5034 , n5035 , n5036 , n5037 , n5038 , n5039 , n5040 , n5041 , n5042 , n5043 , n5044 , n5045 , n5046 , n5047 , n5048 , n5049 , n5050 , n5051 , n5052 , n5053 , n5054 , n5055 , n5056 , n5057 , n5058 , n5059 , n5060 , n5061 , n5062 , n5063 , n5064 , n5065 , n5066 , n5067 , n5068 , n5069 , n5070 , n5071 , n5072 , n5073 , n5074 , n5075 , n5076 , n5077 , n5078 , n5079 , n5080 , n5081 , n5082 , n5083 , n5084 , n5085 , n5086 , n5087 , n5088 , n5089 , n5090 , n5091 , n5092 , n5093 , n5094 , n5095 , n5096 , n5097 , n5098 , n5099 , n5100 , n5101 , n5102 , n5103 , n5104 , n5105 , n5106 , n5107 , n5108 , n5109 , n5110 , n5111 , n5112 , n5113 , n5114 , n5115 , n5116 , n5117 , n5118 , n5119 , n5120 , n5121 , n5122 , n5123 , n5124 , n5125 , n5126 , n5127 , n5128 , n5129 , n5130 , n5131 , n5132 , n5133 , n5134 , n5135 , n5136 , n5137 , n5138 , n5139 , n5140 , n5141 , n5142 , n5143 , n5144 , n5145 , n5146 , n5147 , n5148 , n5149 , n5150 , n5151 , n5152 , n5153 , n5154 , n5155 , n5156 , n5157 , n5158 , n5159 , n5160 , n5161 , n5162 , n5163 , n5164 , n5165 , n5166 , n5167 , n5168 , n5169 , n5170 , n5171 , n5172 , n5173 , n5174 , n5175 , n5176 , n5177 , n5178 , n5179 , n5180 , n5181 , n5182 , n5183 , n5184 , n5185 , n5186 , n5187 , n5188 , n5189 , n5190 , n5191 , n5192 , n5193 , n5194 , n5195 , n5196 , n5197 , n5198 , n5199 , n5200 , n5201 , n5202 , n5203 , n5204 , n5205 , n5206 , n5207 , n5208 , n5209 , n5210 , n5211 , n5212 , n5213 , n5214 , n5215 , n5216 , n5217 , n5218 , n5219 , n5220 , n5221 , n5222 , n5223 , n5224 , n5225 , n5226 , n5227 , n5228 , n5229 , n5230 , n5231 , n5232 , n5233 , n5234 , n5235 , n5236 , n5237 , n5238 , n5239 , n5240 , n5241 , n5242 , n5243 , n5244 , n5245 , n5246 , n5247 , n5248 , n5249 , n5250 , n5251 , n5252 , n5253 , n5254 , n5255 , n5256 , n5257 , n5258 , n5259 , n5260 , n5261 , n5262 , n5263 , n5264 , n5265 , n5266 , n5267 , n5268 , n5269 , n5270 , n5271 , n5272 , n5273 , n5274 , n5275 , n5276 , n5277 , n5278 , n5279 , n5280 , n5281 , n5282 , n5283 , n5284 , n5285 , n5286 , n5287 , n5288 , n5289 , n5290 , n5291 , n5292 , n5293 , n5294 , n5295 , n5296 , n5297 , n5298 , n5299 , n5300 , n5301 , n5302 , n5303 , n5304 , n5305 , n5306 , n5307 , n5308 , n5309 , n5310 , n5311 , n5312 , n5313 , n5314 , n5315 , n5316 , n5317 , n5318 , n5319 , n5320 , n5321 , n5322 , n5323 , n5324 , n5325 , n5326 , n5327 , n5328 , n5329 , n5330 , n5331 , n5332 , n5333 , n5334 , n5335 , n5336 , n5337 , n5338 , n5339 , n5340 , n5341 , n5342 , n5343 , n5344 , n5345 , n5346 , n5347 , n5348 , n5349 , n5350 , n5351 , n5352 , n5353 , n5354 , n5355 , n5356 , n5357 , n5358 , n5359 , n5360 , n5361 , n5362 , n5363 , n5364 , n5365 , n5366 , n5367 , n5368 , n5369 , n5370 , n5371 , n5372 , n5373 , n5374 , n5375 , n5376 , n5377 , n5378 , n5379 , n5380 , n5381 , n5382 , n5383 , n5384 , n5385 , n5386 , n5387 , n5388 , n5389 , n5390 , n5391 , n5392 , n5393 , n5394 , n5395 , n5396 , n5397 , n5398 , n5399 , n5400 , n5401 , n5402 , n5403 , n5404 , n5405 , n5406 , n5407 , n5408 , n5409 , n5410 , n5411 , n5412 , n5413 , n5414 , n5415 , n5416 , n5417 , n5418 , n5419 , n5420 , n5421 , n5422 , n5423 , n5424 , n5425 , n5426 , n5427 , n5428 , n5429 , n5430 , n5431 , n5432 , n5433 , n5434 , n5435 , n5436 , n5437 , n5438 , n5439 , n5440 , n5441 , n5442 , n5443 , n5444 , n5445 , n5446 , n5447 , n5448 , n5449 , n5450 , n5451 , n5452 , n5453 , n5454 , n5455 , n5456 , n5457 , n5458 , n5459 , n5460 , n5461 , n5462 , n5463 , n5464 , n5465 , n5466 , n5467 , n5468 , n5469 , n5470 , n5471 , n5472 , n5473 , n5474 , n5475 , n5476 , n5477 , n5478 , n5479 , n5480 , n5481 , n5482 , n5483 , n5484 , n5485 , n5486 , n5487 , n5488 , n5489 , n5490 , n5491 , n5492 , n5493 , n5494 , n5495 , n5496 , n5497 , n5498 , n5499 , n5500 , n5501 , n5502 , n5503 , n5504 , n5505 , n5506 , n5507 , n5508 , n5509 , n5510 , n5511 , n5512 , n5513 , n5514 , n5515 , n5516 , n5517 , n5518 , n5519 , n5520 , n5521 , n5522 , n5523 , n5524 , n5525 , n5526 , n5527 , n5528 , n5529 , n5530 , n5531 , n5532 , n5533 , n5534 , n5535 , n5536 , n5537 , n5538 , n5539 , n5540 , n5541 , n5542 , n5543 , n5544 , n5545 , n5546 , n5547 , n5548 , n5549 , n5550 , n5551 , n5552 , n5553 , n5554 , n5555 , n5556 , n5557 , n5558 , n5559 , n5560 , n5561 , n5562 , n5563 , n5564 , n5565 , n5566 , n5567 , n5568 , n5569 , n5570 , n5571 , n5572 , n5573 , n5574 , n5575 , n5576 , n5577 , n5578 , n5579 , n5580 , n5581 , n5582 , n5583 , n5584 , n5585 , n5586 , n5587 , n5588 , n5589 , n5590 , n5591 , n5592 , n5593 , n5594 , n5595 , n5596 , n5597 , n5598 , n5599 , n5600 , n5601 , n5602 , n5603 , n5604 , n5605 , n5606 , n5607 , n5608 , n5609 , n5610 , n5611 , n5612 , n5613 , n5614 , n5615 , n5616 , n5617 , n5618 , n5619 , n5620 , n5621 , n5622 , n5623 , n5624 , n5625 , n5626 , n5627 , n5628 , n5629 , n5630 , n5631 , n5632 , n5633 , n5634 , n5635 , n5636 , n5637 , n5638 , n5639 , n5640 , n5641 , n5642 , n5643 , n5644 , n5645 , n5646 , n5647 , n5648 , n5649 , n5650 , n5651 , n5652 , n5653 , n5654 , n5655 , n5656 , n5657 , n5658 , n5659 , n5660 , n5661 , n5662 , n5663 , n5664 , n5665 , n5666 , n5667 , n5668 , n5669 , n5670 , n5671 , n5672 , n5673 , n5674 , n5675 , n5676 , n5677 , n5678 , n5679 , n5680 , n5681 , n5682 , n5683 , n5684 , n5685 , n5686 , n5687 , n5688 , n5689 , n5690 , n5691 , n5692 , n5693 , n5694 , n5695 , n5696 , n5697 , n5698 , n5699 , n5700 , n5701 , n5702 , n5703 , n5704 , n5705 , n5706 , n5707 , n5708 , n5709 , n5710 , n5711 , n5712 , n5713 , n5714 , n5715 , n5716 , n5717 , n5718 , n5719 , n5720 , n5721 , n5722 , n5723 , n5724 , n5725 , n5726 , n5727 , n5728 , n5729 , n5730 , n5731 , n5732 , n5733 , n5734 , n5735 , n5736 , n5737 , n5738 , n5739 , n5740 , n5741 , n5742 , n5743 , n5744 , n5745 , n5746 , n5747 , n5748 , n5749 , n5750 , n5751 , n5752 , n5753 , n5754 , n5755 , n5756 , n5757 , n5758 , n5759 , n5760 , n5761 , n5762 , n5763 , n5764 , n5765 , n5766 , n5767 , n5768 , n5769 , n5770 , n5771 , n5772 , n5773 , n5774 , n5775 , n5776 , n5777 , n5778 , n5779 , n5780 , n5781 , n5782 , n5783 , n5784 , n5785 , n5786 , n5787 , n5788 , n5789 , n5790 , n5791 , n5792 , n5793 , n5794 , n5795 , n5796 , n5797 , n5798 , n5799 , n5800 , n5801 , n5802 , n5803 , n5804 , n5805 , n5806 , n5807 , n5808 , n5809 , n5810 , n5811 , n5812 , n5813 , n5814 , n5815 , n5816 , n5817 , n5818 , n5819 , n5820 , n5821 , n5822 , n5823 , n5824 , n5825 , n5826 , n5827 , n5828 , n5829 , n5830 , n5831 , n5832 , n5833 , n5834 , n5835 , n5836 , n5837 , n5838 , n5839 , n5840 , n5841 , n5842 , n5843 , n5844 , n5845 , n5846 , n5847 , n5848 , n5849 , n5850 , n5851 , n5852 , n5853 , n5854 , n5855 , n5856 , n5857 , n5858 , n5859 , n5860 , n5861 , n5862 , n5863 , n5864 , n5865 , n5866 , n5867 , n5868 , n5869 , n5870 , n5871 , n5872 , n5873 , n5874 , n5875 , n5876 , n5877 , n5878 , n5879 , n5880 , n5881 , n5882 , n5883 , n5884 , n5885 , n5886 , n5887 , n5888 , n5889 , n5890 , n5891 , n5892 , n5893 , n5894 , n5895 , n5896 , n5897 , n5898 , n5899 , n5900 , n5901 , n5902 , n5903 , n5904 , n5905 , n5906 , n5907 , n5908 , n5909 , n5910 , n5911 , n5912 , n5913 , n5914 , n5915 , n5916 , n5917 , n5918 , n5919 , n5920 , n5921 , n5922 , n5923 , n5924 , n5925 , n5926 , n5927 , n5928 , n5929 , n5930 , n5931 , n5932 , n5933 , n5934 , n5935 , n5936 , n5937 , n5938 , n5939 , n5940 , n5941 , n5942 , n5943 , n5944 , n5945 , n5946 , n5947 , n5948 , n5949 , n5950 , n5951 , n5952 , n5953 , n5954 , n5955 , n5956 , n5957 , n5958 , n5959 , n5960 , n5961 , n5962 , n5963 , n5964 , n5965 , n5966 , n5967 , n5968 , n5969 , n5970 , n5971 , n5972 , n5973 , n5974 , n5975 , n5976 , n5977 , n5978 , n5979 , n5980 , n5981 , n5982 , n5983 , n5984 , n5985 , n5986 , n5987 , n5988 , n5989 , n5990 , n5991 , n5992 , n5993 , n5994 , n5995 , n5996 , n5997 , n5998 , n5999 , n6000 , n6001 , n6002 , n6003 , n6004 , n6005 , n6006 , n6007 , n6008 , n6009 , n6010 , n6011 , n6012 , n6013 , n6014 , n6015 , n6016 , n6017 , n6018 , n6019 , n6020 , n6021 , n6022 , n6023 , n6024 , n6025 , n6026 , n6027 , n6028 , n6029 , n6030 , n6031 , n6032 , n6033 , n6034 , n6035 , n6036 , n6037 , n6038 , n6039 , n6040 , n6041 , n6042 , n6043 , n6044 , n6045 , n6046 , n6047 , n6048 , n6049 , n6050 , n6051 , n6052 , n6053 , n6054 , n6055 , n6056 , n6057 , n6058 , n6059 , n6060 , n6061 , n6062 , n6063 , n6064 , n6065 , n6066 , n6067 , n6068 , n6069 , n6070 , n6071 , n6072 , n6073 , n6074 , n6075 , n6076 , n6077 , n6078 , n6079 , n6080 , n6081 , n6082 , n6083 , n6084 , n6085 , n6086 , n6087 , n6088 , n6089 , n6090 , n6091 , n6092 , n6093 , n6094 , n6095 , n6096 , n6097 , n6098 , n6099 , n6100 , n6101 , n6102 , n6103 , n6104 , n6105 , n6106 , n6107 , n6108 , n6109 , n6110 , n6111 , n6112 , n6113 , n6114 , n6115 , n6116 , n6117 , n6118 , n6119 , n6120 , n6121 , n6122 , n6123 , n6124 , n6125 , n6126 , n6127 , n6128 , n6129 , n6130 , n6131 , n6132 , n6133 , n6134 , n6135 , n6136 , n6137 , n6138 , n6139 , n6140 , n6141 , n6142 , n6143 , n6144 , n6145 , n6146 , n6147 , n6148 , n6149 , n6150 , n6151 , n6152 , n6153 , n6154 , n6155 , n6156 , n6157 , n6158 , n6159 , n6160 , n6161 , n6162 , n6163 , n6164 , n6165 , n6166 , n6167 , n6168 , n6169 , n6170 , n6171 , n6172 , n6173 , n6174 , n6175 , n6176 , n6177 , n6178 , n6179 , n6180 , n6181 , n6182 , n6183 , n6184 , n6185 , n6186 , n6187 , n6188 , n6189 , n6190 , n6191 , n6192 , n6193 , n6194 , n6195 , n6196 , n6197 , n6198 , n6199 , n6200 , n6201 , n6202 , n6203 , n6204 , n6205 , n6206 , n6207 , n6208 , n6209 , n6210 , n6211 , n6212 , n6213 , n6214 , n6215 , n6216 , n6217 , n6218 , n6219 , n6220 , n6221 , n6222 , n6223 , n6224 , n6225 , n6226 , n6227 , n6228 , n6229 , n6230 , n6231 , n6232 , n6233 , n6234 , n6235 , n6236 , n6237 , n6238 , n6239 , n6240 , n6241 , n6242 , n6243 , n6244 , n6245 , n6246 , n6247 , n6248 , n6249 , n6250 , n6251 , n6252 , n6253 , n6254 , n6255 , n6256 , n6257 , n6258 , n6259 , n6260 , n6261 , n6262 , n6263 , n6264 , n6265 , n6266 , n6267 , n6268 , n6269 , n6270 , n6271 , n6272 , n6273 , n6274 , n6275 , n6276 , n6277 , n6278 , n6279 , n6280 , n6281 , n6282 , n6283 , n6284 , n6285 , n6286 , n6287 , n6288 , n6289 , n6290 , n6291 , n6292 , n6293 , n6294 , n6295 , n6296 , n6297 , n6298 , n6299 , n6300 , n6301 , n6302 , n6303 , n6304 , n6305 , n6306 , n6307 , n6308 , n6309 , n6310 , n6311 , n6312 , n6313 , n6314 , n6315 , n6316 , n6317 , n6318 , n6319 , n6320 , n6321 , n6322 , n6323 , n6324 , n6325 , n6326 , n6327 , n6328 , n6329 , n6330 , n6331 , n6332 , n6333 , n6334 , n6335 , n6336 , n6337 , n6338 , n6339 , n6340 , n6341 , n6342 , n6343 , n6344 , n6345 , n6346 , n6347 , n6348 , n6349 , n6350 , n6351 , n6352 , n6353 , n6354 , n6355 , n6356 , n6357 , n6358 , n6359 , n6360 , n6361 , n6362 , n6363 , n6364 , n6365 , n6366 , n6367 , n6368 , n6369 , n6370 , n6371 , n6372 , n6373 , n6374 , n6375 , n6376 , n6377 , n6378 , n6379 , n6380 , n6381 , n6382 , n6383 , n6384 , n6385 , n6386 , n6387 , n6388 , n6389 , n6390 , n6391 , n6392 , n6393 , n6394 , n6395 , n6396 , n6397 , n6398 , n6399 , n6400 , n6401 , n6402 , n6403 , n6404 , n6405 , n6406 , n6407 , n6408 , n6409 , n6410 , n6411 , n6412 , n6413 , n6414 , n6415 , n6416 , n6417 , n6418 , n6419 , n6420 , n6421 , n6422 , n6423 , n6424 , n6425 , n6426 , n6427 , n6428 , n6429 , n6430 , n6431 , n6432 , n6433 , n6434 , n6435 , n6436 , n6437 , n6438 , n6439 , n6440 , n6441 , n6442 , n6443 , n6444 ;
  assign n257 = ~x0 & x255 ;
  assign n258 = x128 & ~n257 ;
  assign n259 = x1 & ~x129 ;
  assign n260 = x2 | n259 ;
  assign n261 = x130 | x131 ;
  assign n262 = n260 & ~n261 ;
  assign n263 = ~x5 & x132 ;
  assign n264 = x133 | x134 ;
  assign n265 = n263 | n264 ;
  assign n266 = x3 & ~x131 ;
  assign n267 = x4 | x5 ;
  assign n268 = n266 | n267 ;
  assign n269 = ~n265 & n268 ;
  assign n270 = ( n262 & ~n265 ) | ( n262 & n269 ) | ( ~n265 & n269 ) ;
  assign n271 = ~x8 & x135 ;
  assign n272 = x136 | x137 ;
  assign n273 = n271 | n272 ;
  assign n274 = x6 & ~x134 ;
  assign n275 = x7 | x8 ;
  assign n276 = n274 | n275 ;
  assign n277 = ~n273 & n276 ;
  assign n278 = x9 & ~x137 ;
  assign n279 = x10 | x11 ;
  assign n280 = n278 | n279 ;
  assign n281 = n277 | n280 ;
  assign n282 = n273 & ~n280 ;
  assign n283 = ( n270 & n281 ) | ( n270 & ~n282 ) | ( n281 & ~n282 ) ;
  assign n284 = x15 & ~x143 ;
  assign n285 = x16 | x17 ;
  assign n286 = n284 | n285 ;
  assign n287 = ~x14 & x141 ;
  assign n288 = x142 | x143 ;
  assign n289 = n287 | n288 ;
  assign n290 = x12 & ~x140 ;
  assign n291 = x13 | x14 ;
  assign n292 = n290 | n291 ;
  assign n293 = ~n289 & n292 ;
  assign n294 = n286 | n293 ;
  assign n295 = ~x11 & x138 ;
  assign n296 = x139 | x140 ;
  assign n297 = n295 | n296 ;
  assign n298 = ~n292 & n297 ;
  assign n299 = ~n286 & n289 ;
  assign n300 = ( ~n286 & n298 ) | ( ~n286 & n299 ) | ( n298 & n299 ) ;
  assign n301 = ( n283 & n294 ) | ( n283 & ~n300 ) | ( n294 & ~n300 ) ;
  assign n302 = ~x23 & x150 ;
  assign n303 = x151 | x152 ;
  assign n304 = n302 | n303 ;
  assign n305 = ~x17 & x144 ;
  assign n306 = x145 | x146 ;
  assign n307 = n305 | n306 ;
  assign n308 = x18 & ~x146 ;
  assign n309 = x19 | x20 ;
  assign n310 = n308 | n309 ;
  assign n311 = n307 & ~n310 ;
  assign n312 = x21 & ~x149 ;
  assign n313 = x22 | x23 ;
  assign n314 = n312 | n313 ;
  assign n315 = ~x20 & x147 ;
  assign n316 = x148 | x149 ;
  assign n317 = n315 | n316 ;
  assign n318 = ~n314 & n317 ;
  assign n319 = ( n311 & ~n314 ) | ( n311 & n318 ) | ( ~n314 & n318 ) ;
  assign n320 = n304 | n319 ;
  assign n321 = n310 & ~n317 ;
  assign n322 = ~n304 & n314 ;
  assign n323 = ( ~n304 & n321 ) | ( ~n304 & n322 ) | ( n321 & n322 ) ;
  assign n324 = ( n301 & ~n320 ) | ( n301 & n323 ) | ( ~n320 & n323 ) ;
  assign n325 = ~x32 & x159 ;
  assign n326 = x160 | x161 ;
  assign n327 = n325 | n326 ;
  assign n328 = x30 & ~x158 ;
  assign n329 = x31 | x32 ;
  assign n330 = n328 | n329 ;
  assign n331 = ~x26 & x153 ;
  assign n332 = x154 | x155 ;
  assign n333 = n331 | n332 ;
  assign n334 = x27 & ~x155 ;
  assign n335 = x28 | x29 ;
  assign n336 = n334 | n335 ;
  assign n337 = n333 & ~n336 ;
  assign n338 = ~x29 & x156 ;
  assign n339 = x157 | x158 ;
  assign n340 = n338 | n339 ;
  assign n341 = ~n330 & n340 ;
  assign n342 = ( ~n330 & n337 ) | ( ~n330 & n341 ) | ( n337 & n341 ) ;
  assign n343 = n327 | n342 ;
  assign n344 = ~n327 & n330 ;
  assign n345 = x24 & ~x152 ;
  assign n346 = x25 | x26 ;
  assign n347 = n345 | n346 ;
  assign n348 = ~n333 & n347 ;
  assign n349 = n336 & ~n340 ;
  assign n350 = ( ~n340 & n348 ) | ( ~n340 & n349 ) | ( n348 & n349 ) ;
  assign n351 = ( ~n327 & n344 ) | ( ~n327 & n350 ) | ( n344 & n350 ) ;
  assign n352 = ( n324 & ~n343 ) | ( n324 & n351 ) | ( ~n343 & n351 ) ;
  assign n353 = x42 & ~x170 ;
  assign n354 = x43 | x44 ;
  assign n355 = n353 | n354 ;
  assign n356 = ~x41 & x168 ;
  assign n357 = x169 | x170 ;
  assign n358 = n356 | n357 ;
  assign n359 = ~n355 & n358 ;
  assign n360 = x39 & ~x167 ;
  assign n361 = x40 | x41 ;
  assign n362 = n360 | n361 ;
  assign n363 = ~x35 & x162 ;
  assign n364 = x163 | x164 ;
  assign n365 = n363 | n364 ;
  assign n366 = x36 & ~x164 ;
  assign n367 = x37 | x38 ;
  assign n368 = n366 | n367 ;
  assign n369 = n365 & ~n368 ;
  assign n370 = ~x38 & x165 ;
  assign n371 = x166 | x167 ;
  assign n372 = n370 | n371 ;
  assign n373 = ~n362 & n372 ;
  assign n374 = ( ~n362 & n369 ) | ( ~n362 & n373 ) | ( n369 & n373 ) ;
  assign n375 = ( ~n355 & n359 ) | ( ~n355 & n374 ) | ( n359 & n374 ) ;
  assign n376 = ~n358 & n362 ;
  assign n377 = n355 | n376 ;
  assign n378 = x33 & ~x161 ;
  assign n379 = x34 | x35 ;
  assign n380 = n378 | n379 ;
  assign n381 = ~n365 & n380 ;
  assign n382 = n368 & ~n372 ;
  assign n383 = ( ~n372 & n381 ) | ( ~n372 & n382 ) | ( n381 & n382 ) ;
  assign n384 = ( ~n359 & n377 ) | ( ~n359 & n383 ) | ( n377 & n383 ) ;
  assign n385 = ( n352 & ~n375 ) | ( n352 & n384 ) | ( ~n375 & n384 ) ;
  assign n386 = x54 & ~x182 ;
  assign n387 = x55 | x56 ;
  assign n388 = n386 | n387 ;
  assign n389 = ~x53 & x180 ;
  assign n390 = x181 | x182 ;
  assign n391 = n389 | n390 ;
  assign n392 = x51 & ~x179 ;
  assign n393 = x52 | x53 ;
  assign n394 = n392 | n393 ;
  assign n395 = ~n391 & n394 ;
  assign n396 = ~x44 & x171 ;
  assign n397 = x172 | x173 ;
  assign n398 = n396 | n397 ;
  assign n399 = x45 & ~x173 ;
  assign n400 = x46 | x47 ;
  assign n401 = n399 | n400 ;
  assign n402 = n398 & ~n401 ;
  assign n403 = x48 & ~x176 ;
  assign n404 = x49 | x50 ;
  assign n405 = n403 | n404 ;
  assign n406 = ~x47 & x174 ;
  assign n407 = x175 | x176 ;
  assign n408 = n406 | n407 ;
  assign n409 = ~n405 & n408 ;
  assign n410 = ( n402 & ~n405 ) | ( n402 & n409 ) | ( ~n405 & n409 ) ;
  assign n411 = ~x50 & x177 ;
  assign n412 = x178 | x179 ;
  assign n413 = n411 | n412 ;
  assign n414 = ~n394 & n413 ;
  assign n415 = n391 | n414 ;
  assign n416 = ( ~n395 & n410 ) | ( ~n395 & n415 ) | ( n410 & n415 ) ;
  assign n417 = ~n388 & n416 ;
  assign n418 = n388 | n395 ;
  assign n419 = ~n388 & n391 ;
  assign n420 = n401 & ~n408 ;
  assign n421 = n405 & ~n413 ;
  assign n422 = ( ~n413 & n420 ) | ( ~n413 & n421 ) | ( n420 & n421 ) ;
  assign n423 = ( n418 & ~n419 ) | ( n418 & n422 ) | ( ~n419 & n422 ) ;
  assign n424 = ( n385 & ~n417 ) | ( n385 & n423 ) | ( ~n417 & n423 ) ;
  assign n425 = ~x68 & x195 ;
  assign n426 = x196 | x197 ;
  assign n427 = n425 | n426 ;
  assign n428 = x66 & ~x194 ;
  assign n429 = x67 | x68 ;
  assign n430 = n428 | n429 ;
  assign n431 = ~x65 & x192 ;
  assign n432 = x193 | x194 ;
  assign n433 = n431 | n432 ;
  assign n434 = x63 & ~x191 ;
  assign n435 = x64 | x65 ;
  assign n436 = n434 | n435 ;
  assign n437 = ~n433 & n436 ;
  assign n438 = n430 | n437 ;
  assign n439 = ~n430 & n433 ;
  assign n440 = ~x62 & x189 ;
  assign n441 = x190 | x191 ;
  assign n442 = n440 | n441 ;
  assign n443 = ~x59 & x186 ;
  assign n444 = x187 | x188 ;
  assign n445 = n443 | n444 ;
  assign n446 = x57 & ~x185 ;
  assign n447 = x58 | x59 ;
  assign n448 = n446 | n447 ;
  assign n449 = ~n445 & n448 ;
  assign n450 = x60 & ~x188 ;
  assign n451 = x61 | x62 ;
  assign n452 = n450 | n451 ;
  assign n453 = ~n442 & n452 ;
  assign n454 = ( ~n442 & n449 ) | ( ~n442 & n453 ) | ( n449 & n453 ) ;
  assign n455 = ( n438 & ~n439 ) | ( n438 & n454 ) | ( ~n439 & n454 ) ;
  assign n456 = ~n427 & n455 ;
  assign n457 = ~n427 & n430 ;
  assign n458 = ~x56 & x183 ;
  assign n459 = x184 | x185 ;
  assign n460 = n458 | n459 ;
  assign n461 = ~n448 & n460 ;
  assign n462 = n445 & ~n452 ;
  assign n463 = ( ~n452 & n461 ) | ( ~n452 & n462 ) | ( n461 & n462 ) ;
  assign n464 = ~n436 & n442 ;
  assign n465 = n433 | n464 ;
  assign n466 = ( ~n437 & n463 ) | ( ~n437 & n465 ) | ( n463 & n465 ) ;
  assign n467 = ( n427 & ~n457 ) | ( n427 & n466 ) | ( ~n457 & n466 ) ;
  assign n468 = ( n424 & n456 ) | ( n424 & ~n467 ) | ( n456 & ~n467 ) ;
  assign n469 = ~x83 & x210 ;
  assign n470 = x211 | x212 ;
  assign n471 = n469 | n470 ;
  assign n472 = x81 & ~x209 ;
  assign n473 = x82 | x83 ;
  assign n474 = n472 | n473 ;
  assign n475 = ~n471 & n474 ;
  assign n476 = x78 & ~x206 ;
  assign n477 = x79 | x80 ;
  assign n478 = n476 | n477 ;
  assign n479 = ~x77 & x204 ;
  assign n480 = x205 | x206 ;
  assign n481 = n479 | n480 ;
  assign n482 = x75 & ~x203 ;
  assign n483 = x76 | x77 ;
  assign n484 = n482 | n483 ;
  assign n485 = ~n481 & n484 ;
  assign n486 = n478 | n485 ;
  assign n487 = ~n478 & n481 ;
  assign n488 = ~x74 & x201 ;
  assign n489 = x202 | x203 ;
  assign n490 = n488 | n489 ;
  assign n491 = ~x71 & x198 ;
  assign n492 = x199 | x200 ;
  assign n493 = n491 | n492 ;
  assign n494 = x69 & ~x197 ;
  assign n495 = x70 | x71 ;
  assign n496 = n494 | n495 ;
  assign n497 = ~n493 & n496 ;
  assign n498 = x72 & ~x200 ;
  assign n499 = x73 | x74 ;
  assign n500 = n498 | n499 ;
  assign n501 = ~n490 & n500 ;
  assign n502 = ( ~n490 & n497 ) | ( ~n490 & n501 ) | ( n497 & n501 ) ;
  assign n503 = ( n486 & ~n487 ) | ( n486 & n502 ) | ( ~n487 & n502 ) ;
  assign n504 = ~x80 & x207 ;
  assign n505 = x208 | x209 ;
  assign n506 = n504 | n505 ;
  assign n507 = ~n474 & n506 ;
  assign n508 = n471 | n507 ;
  assign n509 = ( n475 & n503 ) | ( n475 & ~n508 ) | ( n503 & ~n508 ) ;
  assign n510 = n487 | n506 ;
  assign n511 = n478 & ~n506 ;
  assign n512 = n493 & ~n500 ;
  assign n513 = ~n484 & n490 ;
  assign n514 = ( ~n484 & n512 ) | ( ~n484 & n513 ) | ( n512 & n513 ) ;
  assign n515 = ( n510 & ~n511 ) | ( n510 & n514 ) | ( ~n511 & n514 ) ;
  assign n516 = ( n471 & ~n475 ) | ( n471 & n515 ) | ( ~n475 & n515 ) ;
  assign n517 = ( n468 & n509 ) | ( n468 & ~n516 ) | ( n509 & ~n516 ) ;
  assign n518 = x99 & ~x227 ;
  assign n519 = x100 | x101 ;
  assign n520 = n518 | n519 ;
  assign n521 = ~x98 & x225 ;
  assign n522 = x226 | x227 ;
  assign n523 = n521 | n522 ;
  assign n524 = x96 & ~x224 ;
  assign n525 = x97 | x98 ;
  assign n526 = n524 | n525 ;
  assign n527 = ~n523 & n526 ;
  assign n528 = n520 | n527 ;
  assign n529 = x93 & ~x221 ;
  assign n530 = x94 | x95 ;
  assign n531 = n529 | n530 ;
  assign n532 = ~x92 & x219 ;
  assign n533 = x220 | x221 ;
  assign n534 = n532 | n533 ;
  assign n535 = x90 & ~x218 ;
  assign n536 = x91 | x92 ;
  assign n537 = n535 | n536 ;
  assign n538 = ~n534 & n537 ;
  assign n539 = n531 | n538 ;
  assign n540 = ~n531 & n534 ;
  assign n541 = ~x89 & x216 ;
  assign n542 = x217 | x218 ;
  assign n543 = n541 | n542 ;
  assign n544 = ~x86 & x213 ;
  assign n545 = x214 | x215 ;
  assign n546 = n544 | n545 ;
  assign n547 = x84 & ~x212 ;
  assign n548 = x85 | x86 ;
  assign n549 = n547 | n548 ;
  assign n550 = ~n546 & n549 ;
  assign n551 = x87 & ~x215 ;
  assign n552 = x88 | x89 ;
  assign n553 = n551 | n552 ;
  assign n554 = ~n543 & n553 ;
  assign n555 = ( ~n543 & n550 ) | ( ~n543 & n554 ) | ( n550 & n554 ) ;
  assign n556 = ( n539 & ~n540 ) | ( n539 & n555 ) | ( ~n540 & n555 ) ;
  assign n557 = ~x95 & x222 ;
  assign n558 = x223 | x224 ;
  assign n559 = n557 | n558 ;
  assign n560 = ~n526 & n559 ;
  assign n561 = n523 | n560 ;
  assign n562 = ~n520 & n561 ;
  assign n563 = ( n528 & n556 ) | ( n528 & ~n562 ) | ( n556 & ~n562 ) ;
  assign n564 = ~n520 & n523 ;
  assign n565 = n540 | n559 ;
  assign n566 = n531 & ~n559 ;
  assign n567 = n546 & ~n553 ;
  assign n568 = ~n537 & n543 ;
  assign n569 = ( ~n537 & n567 ) | ( ~n537 & n568 ) | ( n567 & n568 ) ;
  assign n570 = ( n565 & ~n566 ) | ( n565 & n569 ) | ( ~n566 & n569 ) ;
  assign n571 = ( ~n528 & n564 ) | ( ~n528 & n570 ) | ( n564 & n570 ) ;
  assign n572 = ( n517 & n563 ) | ( n517 & ~n571 ) | ( n563 & ~n571 ) ;
  assign n573 = ~x116 & x243 ;
  assign n574 = x244 | x245 ;
  assign n575 = n573 | n574 ;
  assign n576 = x114 & ~x242 ;
  assign n577 = x115 | x116 ;
  assign n578 = n576 | n577 ;
  assign n579 = ~x113 & x240 ;
  assign n580 = x241 | x242 ;
  assign n581 = n579 | n580 ;
  assign n582 = x111 & ~x239 ;
  assign n583 = x112 | x113 ;
  assign n584 = n582 | n583 ;
  assign n585 = ~n581 & n584 ;
  assign n586 = ~x110 & x237 ;
  assign n587 = x238 | x239 ;
  assign n588 = n586 | n587 ;
  assign n589 = ~x107 & x234 ;
  assign n590 = x235 | x236 ;
  assign n591 = n589 | n590 ;
  assign n592 = x108 & ~x236 ;
  assign n593 = x109 | x110 ;
  assign n594 = n592 | n593 ;
  assign n595 = n591 & ~n594 ;
  assign n596 = n588 | n595 ;
  assign n597 = ~n588 & n594 ;
  assign n598 = ~x101 & x228 ;
  assign n599 = x229 | x230 ;
  assign n600 = n598 | n599 ;
  assign n601 = x102 & ~x230 ;
  assign n602 = x103 | x104 ;
  assign n603 = n601 | n602 ;
  assign n604 = n600 & ~n603 ;
  assign n605 = x105 & ~x233 ;
  assign n606 = x106 | x107 ;
  assign n607 = n605 | n606 ;
  assign n608 = ~x104 & x231 ;
  assign n609 = x232 | x233 ;
  assign n610 = n608 | n609 ;
  assign n611 = ~n607 & n610 ;
  assign n612 = ( n604 & ~n607 ) | ( n604 & n611 ) | ( ~n607 & n611 ) ;
  assign n613 = ( n596 & ~n597 ) | ( n596 & n612 ) | ( ~n597 & n612 ) ;
  assign n614 = ( n581 & ~n585 ) | ( n581 & n613 ) | ( ~n585 & n613 ) ;
  assign n615 = ~n578 & n614 ;
  assign n616 = n575 | n615 ;
  assign n617 = x117 & ~x245 ;
  assign n618 = x118 | x119 ;
  assign n619 = n617 | n618 ;
  assign n620 = n616 & ~n619 ;
  assign n621 = ~n575 & n578 ;
  assign n622 = n584 | n597 ;
  assign n623 = ~n584 & n588 ;
  assign n624 = n603 & ~n610 ;
  assign n625 = ~n591 & n607 ;
  assign n626 = ( ~n591 & n624 ) | ( ~n591 & n625 ) | ( n624 & n625 ) ;
  assign n627 = ( n622 & ~n623 ) | ( n622 & n626 ) | ( ~n623 & n626 ) ;
  assign n628 = ~n578 & n581 ;
  assign n629 = n575 | n628 ;
  assign n630 = ( n621 & n627 ) | ( n621 & ~n629 ) | ( n627 & ~n629 ) ;
  assign n631 = n619 | n630 ;
  assign n632 = ( n572 & ~n620 ) | ( n572 & n631 ) | ( ~n620 & n631 ) ;
  assign n633 = x126 & ~x254 ;
  assign n634 = x0 | x127 ;
  assign n635 = n633 | n634 ;
  assign n636 = ~x125 & x252 ;
  assign n637 = x253 | x254 ;
  assign n638 = n636 | n637 ;
  assign n639 = ~x122 & x249 ;
  assign n640 = x250 | x251 ;
  assign n641 = n639 | n640 ;
  assign n642 = x120 & ~x248 ;
  assign n643 = x121 | x122 ;
  assign n644 = n642 | n643 ;
  assign n645 = ~n641 & n644 ;
  assign n646 = x123 & ~x251 ;
  assign n647 = x124 | x125 ;
  assign n648 = n646 | n647 ;
  assign n649 = ~n638 & n648 ;
  assign n650 = ( ~n638 & n645 ) | ( ~n638 & n649 ) | ( n645 & n649 ) ;
  assign n651 = n635 | n650 ;
  assign n652 = ~n635 & n638 ;
  assign n653 = ~x119 & x246 ;
  assign n654 = x247 | x248 ;
  assign n655 = n653 | n654 ;
  assign n656 = ~n644 & n655 ;
  assign n657 = n641 & ~n648 ;
  assign n658 = ( ~n648 & n656 ) | ( ~n648 & n657 ) | ( n656 & n657 ) ;
  assign n659 = ( ~n635 & n652 ) | ( ~n635 & n658 ) | ( n652 & n658 ) ;
  assign n660 = ( n632 & n651 ) | ( n632 & ~n659 ) | ( n651 & ~n659 ) ;
  assign n661 = n258 & n660 ;
  assign n662 = ~x1 & x128 ;
  assign n663 = x129 & ~n662 ;
  assign n664 = x2 & ~x130 ;
  assign n665 = x3 | n664 ;
  assign n666 = x131 | x132 ;
  assign n667 = n665 & ~n666 ;
  assign n668 = ~x6 & x133 ;
  assign n669 = x134 | x135 ;
  assign n670 = n668 | n669 ;
  assign n671 = x4 & ~x132 ;
  assign n672 = x5 | x6 ;
  assign n673 = n671 | n672 ;
  assign n674 = ~n670 & n673 ;
  assign n675 = ( n667 & ~n670 ) | ( n667 & n674 ) | ( ~n670 & n674 ) ;
  assign n676 = ~x9 & x136 ;
  assign n677 = x137 | x138 ;
  assign n678 = n676 | n677 ;
  assign n679 = x7 & ~x135 ;
  assign n680 = x8 | x9 ;
  assign n681 = n679 | n680 ;
  assign n682 = ~n678 & n681 ;
  assign n683 = x10 & ~x138 ;
  assign n684 = x11 | x12 ;
  assign n685 = n683 | n684 ;
  assign n686 = n682 | n685 ;
  assign n687 = n678 & ~n685 ;
  assign n688 = ( n675 & n686 ) | ( n675 & ~n687 ) | ( n686 & ~n687 ) ;
  assign n689 = x16 & ~x144 ;
  assign n690 = x17 | x18 ;
  assign n691 = n689 | n690 ;
  assign n692 = ~x15 & x142 ;
  assign n693 = x143 | x144 ;
  assign n694 = n692 | n693 ;
  assign n695 = x13 & ~x141 ;
  assign n696 = x14 | x15 ;
  assign n697 = n695 | n696 ;
  assign n698 = ~n694 & n697 ;
  assign n699 = n691 | n698 ;
  assign n700 = ~x12 & x139 ;
  assign n701 = x140 | x141 ;
  assign n702 = n700 | n701 ;
  assign n703 = ~n697 & n702 ;
  assign n704 = ~n691 & n694 ;
  assign n705 = ( ~n691 & n703 ) | ( ~n691 & n704 ) | ( n703 & n704 ) ;
  assign n706 = ( n688 & n699 ) | ( n688 & ~n705 ) | ( n699 & ~n705 ) ;
  assign n707 = ~x24 & x151 ;
  assign n708 = x152 | x153 ;
  assign n709 = n707 | n708 ;
  assign n710 = ~x18 & x145 ;
  assign n711 = x146 | x147 ;
  assign n712 = n710 | n711 ;
  assign n713 = x19 & ~x147 ;
  assign n714 = x20 | x21 ;
  assign n715 = n713 | n714 ;
  assign n716 = n712 & ~n715 ;
  assign n717 = x22 & ~x150 ;
  assign n718 = x23 | x24 ;
  assign n719 = n717 | n718 ;
  assign n720 = ~x21 & x148 ;
  assign n721 = x149 | x150 ;
  assign n722 = n720 | n721 ;
  assign n723 = ~n719 & n722 ;
  assign n724 = ( n716 & ~n719 ) | ( n716 & n723 ) | ( ~n719 & n723 ) ;
  assign n725 = n709 | n724 ;
  assign n726 = n715 & ~n722 ;
  assign n727 = ~n709 & n719 ;
  assign n728 = ( ~n709 & n726 ) | ( ~n709 & n727 ) | ( n726 & n727 ) ;
  assign n729 = ( n706 & ~n725 ) | ( n706 & n728 ) | ( ~n725 & n728 ) ;
  assign n730 = ~x33 & x160 ;
  assign n731 = x161 | x162 ;
  assign n732 = n730 | n731 ;
  assign n733 = x31 & ~x159 ;
  assign n734 = x32 | x33 ;
  assign n735 = n733 | n734 ;
  assign n736 = ~x27 & x154 ;
  assign n737 = x155 | x156 ;
  assign n738 = n736 | n737 ;
  assign n739 = x28 & ~x156 ;
  assign n740 = x29 | x30 ;
  assign n741 = n739 | n740 ;
  assign n742 = n738 & ~n741 ;
  assign n743 = ~x30 & x157 ;
  assign n744 = x158 | x159 ;
  assign n745 = n743 | n744 ;
  assign n746 = ~n735 & n745 ;
  assign n747 = ( ~n735 & n742 ) | ( ~n735 & n746 ) | ( n742 & n746 ) ;
  assign n748 = n732 | n747 ;
  assign n749 = ~n732 & n735 ;
  assign n750 = x25 & ~x153 ;
  assign n751 = x26 | x27 ;
  assign n752 = n750 | n751 ;
  assign n753 = ~n738 & n752 ;
  assign n754 = n741 & ~n745 ;
  assign n755 = ( ~n745 & n753 ) | ( ~n745 & n754 ) | ( n753 & n754 ) ;
  assign n756 = ( ~n732 & n749 ) | ( ~n732 & n755 ) | ( n749 & n755 ) ;
  assign n757 = ( n729 & ~n748 ) | ( n729 & n756 ) | ( ~n748 & n756 ) ;
  assign n758 = x43 & ~x171 ;
  assign n759 = x44 | x45 ;
  assign n760 = n758 | n759 ;
  assign n761 = ~x42 & x169 ;
  assign n762 = x170 | x171 ;
  assign n763 = n761 | n762 ;
  assign n764 = ~n760 & n763 ;
  assign n765 = x40 & ~x168 ;
  assign n766 = x41 | x42 ;
  assign n767 = n765 | n766 ;
  assign n768 = ~x36 & x163 ;
  assign n769 = x164 | x165 ;
  assign n770 = n768 | n769 ;
  assign n771 = x37 & ~x165 ;
  assign n772 = x38 | x39 ;
  assign n773 = n771 | n772 ;
  assign n774 = n770 & ~n773 ;
  assign n775 = ~x39 & x166 ;
  assign n776 = x167 | x168 ;
  assign n777 = n775 | n776 ;
  assign n778 = ~n767 & n777 ;
  assign n779 = ( ~n767 & n774 ) | ( ~n767 & n778 ) | ( n774 & n778 ) ;
  assign n780 = ( ~n760 & n764 ) | ( ~n760 & n779 ) | ( n764 & n779 ) ;
  assign n781 = ~n763 & n767 ;
  assign n782 = n760 | n781 ;
  assign n783 = x34 & ~x162 ;
  assign n784 = x35 | x36 ;
  assign n785 = n783 | n784 ;
  assign n786 = ~n770 & n785 ;
  assign n787 = n773 & ~n777 ;
  assign n788 = ( ~n777 & n786 ) | ( ~n777 & n787 ) | ( n786 & n787 ) ;
  assign n789 = ( ~n764 & n782 ) | ( ~n764 & n788 ) | ( n782 & n788 ) ;
  assign n790 = ( n757 & ~n780 ) | ( n757 & n789 ) | ( ~n780 & n789 ) ;
  assign n791 = x55 & ~x183 ;
  assign n792 = x56 | x57 ;
  assign n793 = n791 | n792 ;
  assign n794 = ~x54 & x181 ;
  assign n795 = x182 | x183 ;
  assign n796 = n794 | n795 ;
  assign n797 = x52 & ~x180 ;
  assign n798 = x53 | x54 ;
  assign n799 = n797 | n798 ;
  assign n800 = ~n796 & n799 ;
  assign n801 = ~x45 & x172 ;
  assign n802 = x173 | x174 ;
  assign n803 = n801 | n802 ;
  assign n804 = x46 & ~x174 ;
  assign n805 = x47 | x48 ;
  assign n806 = n804 | n805 ;
  assign n807 = n803 & ~n806 ;
  assign n808 = x49 & ~x177 ;
  assign n809 = x50 | x51 ;
  assign n810 = n808 | n809 ;
  assign n811 = ~x48 & x175 ;
  assign n812 = x176 | x177 ;
  assign n813 = n811 | n812 ;
  assign n814 = ~n810 & n813 ;
  assign n815 = ( n807 & ~n810 ) | ( n807 & n814 ) | ( ~n810 & n814 ) ;
  assign n816 = ~x51 & x178 ;
  assign n817 = x179 | x180 ;
  assign n818 = n816 | n817 ;
  assign n819 = ~n799 & n818 ;
  assign n820 = n796 | n819 ;
  assign n821 = ( ~n800 & n815 ) | ( ~n800 & n820 ) | ( n815 & n820 ) ;
  assign n822 = ~n793 & n821 ;
  assign n823 = n793 | n800 ;
  assign n824 = ~n793 & n796 ;
  assign n825 = n806 & ~n813 ;
  assign n826 = n810 & ~n818 ;
  assign n827 = ( ~n818 & n825 ) | ( ~n818 & n826 ) | ( n825 & n826 ) ;
  assign n828 = ( n823 & ~n824 ) | ( n823 & n827 ) | ( ~n824 & n827 ) ;
  assign n829 = ( n790 & ~n822 ) | ( n790 & n828 ) | ( ~n822 & n828 ) ;
  assign n830 = ~x69 & x196 ;
  assign n831 = x197 | x198 ;
  assign n832 = n830 | n831 ;
  assign n833 = x67 & ~x195 ;
  assign n834 = x68 | x69 ;
  assign n835 = n833 | n834 ;
  assign n836 = ~x66 & x193 ;
  assign n837 = x194 | x195 ;
  assign n838 = n836 | n837 ;
  assign n839 = x64 & ~x192 ;
  assign n840 = x65 | x66 ;
  assign n841 = n839 | n840 ;
  assign n842 = ~n838 & n841 ;
  assign n843 = n835 | n842 ;
  assign n844 = ~n835 & n838 ;
  assign n845 = ~x63 & x190 ;
  assign n846 = x191 | x192 ;
  assign n847 = n845 | n846 ;
  assign n848 = ~x60 & x187 ;
  assign n849 = x188 | x189 ;
  assign n850 = n848 | n849 ;
  assign n851 = x58 & ~x186 ;
  assign n852 = x59 | x60 ;
  assign n853 = n851 | n852 ;
  assign n854 = ~n850 & n853 ;
  assign n855 = x61 & ~x189 ;
  assign n856 = x62 | x63 ;
  assign n857 = n855 | n856 ;
  assign n858 = ~n847 & n857 ;
  assign n859 = ( ~n847 & n854 ) | ( ~n847 & n858 ) | ( n854 & n858 ) ;
  assign n860 = ( n843 & ~n844 ) | ( n843 & n859 ) | ( ~n844 & n859 ) ;
  assign n861 = ~n832 & n860 ;
  assign n862 = ~n832 & n835 ;
  assign n863 = ~x57 & x184 ;
  assign n864 = x185 | x186 ;
  assign n865 = n863 | n864 ;
  assign n866 = ~n853 & n865 ;
  assign n867 = n850 & ~n857 ;
  assign n868 = ( ~n857 & n866 ) | ( ~n857 & n867 ) | ( n866 & n867 ) ;
  assign n869 = ~n841 & n847 ;
  assign n870 = n838 | n869 ;
  assign n871 = ( ~n842 & n868 ) | ( ~n842 & n870 ) | ( n868 & n870 ) ;
  assign n872 = ( n832 & ~n862 ) | ( n832 & n871 ) | ( ~n862 & n871 ) ;
  assign n873 = ( n829 & n861 ) | ( n829 & ~n872 ) | ( n861 & ~n872 ) ;
  assign n874 = ~x84 & x211 ;
  assign n875 = x212 | x213 ;
  assign n876 = n874 | n875 ;
  assign n877 = x82 & ~x210 ;
  assign n878 = x83 | x84 ;
  assign n879 = n877 | n878 ;
  assign n880 = ~n876 & n879 ;
  assign n881 = x79 & ~x207 ;
  assign n882 = x80 | x81 ;
  assign n883 = n881 | n882 ;
  assign n884 = ~x78 & x205 ;
  assign n885 = x206 | x207 ;
  assign n886 = n884 | n885 ;
  assign n887 = x76 & ~x204 ;
  assign n888 = x77 | x78 ;
  assign n889 = n887 | n888 ;
  assign n890 = ~n886 & n889 ;
  assign n891 = n883 | n890 ;
  assign n892 = ~n883 & n886 ;
  assign n893 = ~x75 & x202 ;
  assign n894 = x203 | x204 ;
  assign n895 = n893 | n894 ;
  assign n896 = ~x72 & x199 ;
  assign n897 = x200 | x201 ;
  assign n898 = n896 | n897 ;
  assign n899 = x70 & ~x198 ;
  assign n900 = x71 | x72 ;
  assign n901 = n899 | n900 ;
  assign n902 = ~n898 & n901 ;
  assign n903 = x73 & ~x201 ;
  assign n904 = x74 | x75 ;
  assign n905 = n903 | n904 ;
  assign n906 = ~n895 & n905 ;
  assign n907 = ( ~n895 & n902 ) | ( ~n895 & n906 ) | ( n902 & n906 ) ;
  assign n908 = ( n891 & ~n892 ) | ( n891 & n907 ) | ( ~n892 & n907 ) ;
  assign n909 = ~x81 & x208 ;
  assign n910 = x209 | x210 ;
  assign n911 = n909 | n910 ;
  assign n912 = ~n879 & n911 ;
  assign n913 = n876 | n912 ;
  assign n914 = ( n880 & n908 ) | ( n880 & ~n913 ) | ( n908 & ~n913 ) ;
  assign n915 = n892 | n911 ;
  assign n916 = n883 & ~n911 ;
  assign n917 = n898 & ~n905 ;
  assign n918 = ~n889 & n895 ;
  assign n919 = ( ~n889 & n917 ) | ( ~n889 & n918 ) | ( n917 & n918 ) ;
  assign n920 = ( n915 & ~n916 ) | ( n915 & n919 ) | ( ~n916 & n919 ) ;
  assign n921 = ( n876 & ~n880 ) | ( n876 & n920 ) | ( ~n880 & n920 ) ;
  assign n922 = ( n873 & n914 ) | ( n873 & ~n921 ) | ( n914 & ~n921 ) ;
  assign n923 = x100 & ~x228 ;
  assign n924 = x101 | x102 ;
  assign n925 = n923 | n924 ;
  assign n926 = ~x99 & x226 ;
  assign n927 = x227 | x228 ;
  assign n928 = n926 | n927 ;
  assign n929 = x97 & ~x225 ;
  assign n930 = x98 | x99 ;
  assign n931 = n929 | n930 ;
  assign n932 = ~n928 & n931 ;
  assign n933 = n925 | n932 ;
  assign n934 = x94 & ~x222 ;
  assign n935 = x95 | x96 ;
  assign n936 = n934 | n935 ;
  assign n937 = ~x93 & x220 ;
  assign n938 = x221 | x222 ;
  assign n939 = n937 | n938 ;
  assign n940 = x91 & ~x219 ;
  assign n941 = x92 | x93 ;
  assign n942 = n940 | n941 ;
  assign n943 = ~n939 & n942 ;
  assign n944 = n936 | n943 ;
  assign n945 = ~n936 & n939 ;
  assign n946 = ~x90 & x217 ;
  assign n947 = x218 | x219 ;
  assign n948 = n946 | n947 ;
  assign n949 = ~x87 & x214 ;
  assign n950 = x215 | x216 ;
  assign n951 = n949 | n950 ;
  assign n952 = x85 & ~x213 ;
  assign n953 = x86 | x87 ;
  assign n954 = n952 | n953 ;
  assign n955 = ~n951 & n954 ;
  assign n956 = x88 & ~x216 ;
  assign n957 = x89 | x90 ;
  assign n958 = n956 | n957 ;
  assign n959 = ~n948 & n958 ;
  assign n960 = ( ~n948 & n955 ) | ( ~n948 & n959 ) | ( n955 & n959 ) ;
  assign n961 = ( n944 & ~n945 ) | ( n944 & n960 ) | ( ~n945 & n960 ) ;
  assign n962 = ~x96 & x223 ;
  assign n963 = x224 | x225 ;
  assign n964 = n962 | n963 ;
  assign n965 = ~n931 & n964 ;
  assign n966 = n928 | n965 ;
  assign n967 = ~n925 & n966 ;
  assign n968 = ( n933 & n961 ) | ( n933 & ~n967 ) | ( n961 & ~n967 ) ;
  assign n969 = ~n925 & n928 ;
  assign n970 = n945 | n964 ;
  assign n971 = n936 & ~n964 ;
  assign n972 = n951 & ~n958 ;
  assign n973 = ~n942 & n948 ;
  assign n974 = ( ~n942 & n972 ) | ( ~n942 & n973 ) | ( n972 & n973 ) ;
  assign n975 = ( n970 & ~n971 ) | ( n970 & n974 ) | ( ~n971 & n974 ) ;
  assign n976 = ( ~n933 & n969 ) | ( ~n933 & n975 ) | ( n969 & n975 ) ;
  assign n977 = ( n922 & n968 ) | ( n922 & ~n976 ) | ( n968 & ~n976 ) ;
  assign n978 = ~x117 & x244 ;
  assign n979 = x245 | x246 ;
  assign n980 = n978 | n979 ;
  assign n981 = x115 & ~x243 ;
  assign n982 = x116 | x117 ;
  assign n983 = n981 | n982 ;
  assign n984 = ~x114 & x241 ;
  assign n985 = x242 | x243 ;
  assign n986 = n984 | n985 ;
  assign n987 = x112 & ~x240 ;
  assign n988 = x113 | x114 ;
  assign n989 = n987 | n988 ;
  assign n990 = ~n986 & n989 ;
  assign n991 = ~x111 & x238 ;
  assign n992 = x239 | x240 ;
  assign n993 = n991 | n992 ;
  assign n994 = ~x108 & x235 ;
  assign n995 = x236 | x237 ;
  assign n996 = n994 | n995 ;
  assign n997 = x109 & ~x237 ;
  assign n998 = x110 | x111 ;
  assign n999 = n997 | n998 ;
  assign n1000 = n996 & ~n999 ;
  assign n1001 = n993 | n1000 ;
  assign n1002 = ~n993 & n999 ;
  assign n1003 = ~x102 & x229 ;
  assign n1004 = x230 | x231 ;
  assign n1005 = n1003 | n1004 ;
  assign n1006 = x103 & ~x231 ;
  assign n1007 = x104 | x105 ;
  assign n1008 = n1006 | n1007 ;
  assign n1009 = n1005 & ~n1008 ;
  assign n1010 = x106 & ~x234 ;
  assign n1011 = x107 | x108 ;
  assign n1012 = n1010 | n1011 ;
  assign n1013 = ~x105 & x232 ;
  assign n1014 = x233 | x234 ;
  assign n1015 = n1013 | n1014 ;
  assign n1016 = ~n1012 & n1015 ;
  assign n1017 = ( n1009 & ~n1012 ) | ( n1009 & n1016 ) | ( ~n1012 & n1016 ) ;
  assign n1018 = ( n1001 & ~n1002 ) | ( n1001 & n1017 ) | ( ~n1002 & n1017 ) ;
  assign n1019 = ( n986 & ~n990 ) | ( n986 & n1018 ) | ( ~n990 & n1018 ) ;
  assign n1020 = ~n983 & n1019 ;
  assign n1021 = n980 | n1020 ;
  assign n1022 = x118 & ~x246 ;
  assign n1023 = x119 | x120 ;
  assign n1024 = n1022 | n1023 ;
  assign n1025 = n1021 & ~n1024 ;
  assign n1026 = ~n980 & n983 ;
  assign n1027 = n989 | n1002 ;
  assign n1028 = ~n989 & n993 ;
  assign n1029 = n1008 & ~n1015 ;
  assign n1030 = ~n996 & n1012 ;
  assign n1031 = ( ~n996 & n1029 ) | ( ~n996 & n1030 ) | ( n1029 & n1030 ) ;
  assign n1032 = ( n1027 & ~n1028 ) | ( n1027 & n1031 ) | ( ~n1028 & n1031 ) ;
  assign n1033 = ~n983 & n986 ;
  assign n1034 = n980 | n1033 ;
  assign n1035 = ( n1026 & n1032 ) | ( n1026 & ~n1034 ) | ( n1032 & ~n1034 ) ;
  assign n1036 = n1024 | n1035 ;
  assign n1037 = ( n977 & ~n1025 ) | ( n977 & n1036 ) | ( ~n1025 & n1036 ) ;
  assign n1038 = x127 & ~x255 ;
  assign n1039 = x0 | x1 ;
  assign n1040 = n1038 | n1039 ;
  assign n1041 = ~x126 & x253 ;
  assign n1042 = x254 | x255 ;
  assign n1043 = n1041 | n1042 ;
  assign n1044 = ~x123 & x250 ;
  assign n1045 = x251 | x252 ;
  assign n1046 = n1044 | n1045 ;
  assign n1047 = x121 & ~x249 ;
  assign n1048 = x122 | x123 ;
  assign n1049 = n1047 | n1048 ;
  assign n1050 = ~n1046 & n1049 ;
  assign n1051 = x124 & ~x252 ;
  assign n1052 = x125 | x126 ;
  assign n1053 = n1051 | n1052 ;
  assign n1054 = ~n1043 & n1053 ;
  assign n1055 = ( ~n1043 & n1050 ) | ( ~n1043 & n1054 ) | ( n1050 & n1054 ) ;
  assign n1056 = n1040 | n1055 ;
  assign n1057 = ~n1040 & n1043 ;
  assign n1058 = ~x120 & x247 ;
  assign n1059 = x248 | x249 ;
  assign n1060 = n1058 | n1059 ;
  assign n1061 = ~n1049 & n1060 ;
  assign n1062 = n1046 & ~n1053 ;
  assign n1063 = ( ~n1053 & n1061 ) | ( ~n1053 & n1062 ) | ( n1061 & n1062 ) ;
  assign n1064 = ( ~n1040 & n1057 ) | ( ~n1040 & n1063 ) | ( n1057 & n1063 ) ;
  assign n1065 = ( n1037 & n1056 ) | ( n1037 & ~n1064 ) | ( n1056 & ~n1064 ) ;
  assign n1066 = n663 & n1065 ;
  assign n1067 = ~x2 & x129 ;
  assign n1068 = x130 & ~n1067 ;
  assign n1069 = x4 | n266 ;
  assign n1070 = x132 | x133 ;
  assign n1071 = n1069 & ~n1070 ;
  assign n1072 = ~x7 & x134 ;
  assign n1073 = x135 | x136 ;
  assign n1074 = n1072 | n1073 ;
  assign n1075 = x5 & ~x133 ;
  assign n1076 = x6 | x7 ;
  assign n1077 = n1075 | n1076 ;
  assign n1078 = ~n1074 & n1077 ;
  assign n1079 = ( n1071 & ~n1074 ) | ( n1071 & n1078 ) | ( ~n1074 & n1078 ) ;
  assign n1080 = ~x10 & x137 ;
  assign n1081 = x138 | x139 ;
  assign n1082 = n1080 | n1081 ;
  assign n1083 = x8 & ~x136 ;
  assign n1084 = x9 | x10 ;
  assign n1085 = n1083 | n1084 ;
  assign n1086 = ~n1082 & n1085 ;
  assign n1087 = x11 & ~x139 ;
  assign n1088 = x12 | x13 ;
  assign n1089 = n1087 | n1088 ;
  assign n1090 = n1086 | n1089 ;
  assign n1091 = n1082 & ~n1089 ;
  assign n1092 = ( n1079 & n1090 ) | ( n1079 & ~n1091 ) | ( n1090 & ~n1091 ) ;
  assign n1093 = x17 & ~x145 ;
  assign n1094 = x18 | x19 ;
  assign n1095 = n1093 | n1094 ;
  assign n1096 = ~x16 & x143 ;
  assign n1097 = x144 | x145 ;
  assign n1098 = n1096 | n1097 ;
  assign n1099 = x14 & ~x142 ;
  assign n1100 = x15 | x16 ;
  assign n1101 = n1099 | n1100 ;
  assign n1102 = ~n1098 & n1101 ;
  assign n1103 = n1095 | n1102 ;
  assign n1104 = ~x13 & x140 ;
  assign n1105 = x141 | x142 ;
  assign n1106 = n1104 | n1105 ;
  assign n1107 = ~n1101 & n1106 ;
  assign n1108 = ~n1095 & n1098 ;
  assign n1109 = ( ~n1095 & n1107 ) | ( ~n1095 & n1108 ) | ( n1107 & n1108 ) ;
  assign n1110 = ( n1092 & n1103 ) | ( n1092 & ~n1109 ) | ( n1103 & ~n1109 ) ;
  assign n1111 = ~x25 & x152 ;
  assign n1112 = x153 | x154 ;
  assign n1113 = n1111 | n1112 ;
  assign n1114 = ~x19 & x146 ;
  assign n1115 = x147 | x148 ;
  assign n1116 = n1114 | n1115 ;
  assign n1117 = x20 & ~x148 ;
  assign n1118 = x21 | x22 ;
  assign n1119 = n1117 | n1118 ;
  assign n1120 = n1116 & ~n1119 ;
  assign n1121 = x23 & ~x151 ;
  assign n1122 = x24 | x25 ;
  assign n1123 = n1121 | n1122 ;
  assign n1124 = ~x22 & x149 ;
  assign n1125 = x150 | x151 ;
  assign n1126 = n1124 | n1125 ;
  assign n1127 = ~n1123 & n1126 ;
  assign n1128 = ( n1120 & ~n1123 ) | ( n1120 & n1127 ) | ( ~n1123 & n1127 ) ;
  assign n1129 = n1113 | n1128 ;
  assign n1130 = n1119 & ~n1126 ;
  assign n1131 = ~n1113 & n1123 ;
  assign n1132 = ( ~n1113 & n1130 ) | ( ~n1113 & n1131 ) | ( n1130 & n1131 ) ;
  assign n1133 = ( n1110 & ~n1129 ) | ( n1110 & n1132 ) | ( ~n1129 & n1132 ) ;
  assign n1134 = ~x34 & x161 ;
  assign n1135 = x162 | x163 ;
  assign n1136 = n1134 | n1135 ;
  assign n1137 = x32 & ~x160 ;
  assign n1138 = x33 | x34 ;
  assign n1139 = n1137 | n1138 ;
  assign n1140 = ~x28 & x155 ;
  assign n1141 = x156 | x157 ;
  assign n1142 = n1140 | n1141 ;
  assign n1143 = x29 & ~x157 ;
  assign n1144 = x30 | x31 ;
  assign n1145 = n1143 | n1144 ;
  assign n1146 = n1142 & ~n1145 ;
  assign n1147 = ~x31 & x158 ;
  assign n1148 = x159 | x160 ;
  assign n1149 = n1147 | n1148 ;
  assign n1150 = ~n1139 & n1149 ;
  assign n1151 = ( ~n1139 & n1146 ) | ( ~n1139 & n1150 ) | ( n1146 & n1150 ) ;
  assign n1152 = n1136 | n1151 ;
  assign n1153 = ~n1136 & n1139 ;
  assign n1154 = x26 & ~x154 ;
  assign n1155 = x27 | x28 ;
  assign n1156 = n1154 | n1155 ;
  assign n1157 = ~n1142 & n1156 ;
  assign n1158 = n1145 & ~n1149 ;
  assign n1159 = ( ~n1149 & n1157 ) | ( ~n1149 & n1158 ) | ( n1157 & n1158 ) ;
  assign n1160 = ( ~n1136 & n1153 ) | ( ~n1136 & n1159 ) | ( n1153 & n1159 ) ;
  assign n1161 = ( n1133 & ~n1152 ) | ( n1133 & n1160 ) | ( ~n1152 & n1160 ) ;
  assign n1162 = x44 & ~x172 ;
  assign n1163 = x45 | x46 ;
  assign n1164 = n1162 | n1163 ;
  assign n1165 = ~x43 & x170 ;
  assign n1166 = x171 | x172 ;
  assign n1167 = n1165 | n1166 ;
  assign n1168 = ~n1164 & n1167 ;
  assign n1169 = x41 & ~x169 ;
  assign n1170 = x42 | x43 ;
  assign n1171 = n1169 | n1170 ;
  assign n1172 = ~x37 & x164 ;
  assign n1173 = x165 | x166 ;
  assign n1174 = n1172 | n1173 ;
  assign n1175 = x38 & ~x166 ;
  assign n1176 = x39 | x40 ;
  assign n1177 = n1175 | n1176 ;
  assign n1178 = n1174 & ~n1177 ;
  assign n1179 = ~x40 & x167 ;
  assign n1180 = x168 | x169 ;
  assign n1181 = n1179 | n1180 ;
  assign n1182 = ~n1171 & n1181 ;
  assign n1183 = ( ~n1171 & n1178 ) | ( ~n1171 & n1182 ) | ( n1178 & n1182 ) ;
  assign n1184 = ( ~n1164 & n1168 ) | ( ~n1164 & n1183 ) | ( n1168 & n1183 ) ;
  assign n1185 = ~n1167 & n1171 ;
  assign n1186 = n1164 | n1185 ;
  assign n1187 = x35 & ~x163 ;
  assign n1188 = x36 | x37 ;
  assign n1189 = n1187 | n1188 ;
  assign n1190 = ~n1174 & n1189 ;
  assign n1191 = n1177 & ~n1181 ;
  assign n1192 = ( ~n1181 & n1190 ) | ( ~n1181 & n1191 ) | ( n1190 & n1191 ) ;
  assign n1193 = ( ~n1168 & n1186 ) | ( ~n1168 & n1192 ) | ( n1186 & n1192 ) ;
  assign n1194 = ( n1161 & ~n1184 ) | ( n1161 & n1193 ) | ( ~n1184 & n1193 ) ;
  assign n1195 = x56 & ~x184 ;
  assign n1196 = x57 | x58 ;
  assign n1197 = n1195 | n1196 ;
  assign n1198 = ~x55 & x182 ;
  assign n1199 = x183 | x184 ;
  assign n1200 = n1198 | n1199 ;
  assign n1201 = x53 & ~x181 ;
  assign n1202 = x54 | x55 ;
  assign n1203 = n1201 | n1202 ;
  assign n1204 = ~n1200 & n1203 ;
  assign n1205 = ~x46 & x173 ;
  assign n1206 = x174 | x175 ;
  assign n1207 = n1205 | n1206 ;
  assign n1208 = x47 & ~x175 ;
  assign n1209 = x48 | x49 ;
  assign n1210 = n1208 | n1209 ;
  assign n1211 = n1207 & ~n1210 ;
  assign n1212 = x50 & ~x178 ;
  assign n1213 = x51 | x52 ;
  assign n1214 = n1212 | n1213 ;
  assign n1215 = ~x49 & x176 ;
  assign n1216 = x177 | x178 ;
  assign n1217 = n1215 | n1216 ;
  assign n1218 = ~n1214 & n1217 ;
  assign n1219 = ( n1211 & ~n1214 ) | ( n1211 & n1218 ) | ( ~n1214 & n1218 ) ;
  assign n1220 = ~x52 & x179 ;
  assign n1221 = x180 | x181 ;
  assign n1222 = n1220 | n1221 ;
  assign n1223 = ~n1203 & n1222 ;
  assign n1224 = n1200 | n1223 ;
  assign n1225 = ( ~n1204 & n1219 ) | ( ~n1204 & n1224 ) | ( n1219 & n1224 ) ;
  assign n1226 = ~n1197 & n1225 ;
  assign n1227 = n1197 | n1204 ;
  assign n1228 = ~n1197 & n1200 ;
  assign n1229 = n1210 & ~n1217 ;
  assign n1230 = n1214 & ~n1222 ;
  assign n1231 = ( ~n1222 & n1229 ) | ( ~n1222 & n1230 ) | ( n1229 & n1230 ) ;
  assign n1232 = ( n1227 & ~n1228 ) | ( n1227 & n1231 ) | ( ~n1228 & n1231 ) ;
  assign n1233 = ( n1194 & ~n1226 ) | ( n1194 & n1232 ) | ( ~n1226 & n1232 ) ;
  assign n1234 = ~x70 & x197 ;
  assign n1235 = x198 | x199 ;
  assign n1236 = n1234 | n1235 ;
  assign n1237 = x68 & ~x196 ;
  assign n1238 = x69 | x70 ;
  assign n1239 = n1237 | n1238 ;
  assign n1240 = ~x67 & x194 ;
  assign n1241 = x195 | x196 ;
  assign n1242 = n1240 | n1241 ;
  assign n1243 = x65 & ~x193 ;
  assign n1244 = x66 | x67 ;
  assign n1245 = n1243 | n1244 ;
  assign n1246 = ~n1242 & n1245 ;
  assign n1247 = n1239 | n1246 ;
  assign n1248 = ~n1239 & n1242 ;
  assign n1249 = ~x64 & x191 ;
  assign n1250 = x192 | x193 ;
  assign n1251 = n1249 | n1250 ;
  assign n1252 = ~x61 & x188 ;
  assign n1253 = x189 | x190 ;
  assign n1254 = n1252 | n1253 ;
  assign n1255 = x59 & ~x187 ;
  assign n1256 = x60 | x61 ;
  assign n1257 = n1255 | n1256 ;
  assign n1258 = ~n1254 & n1257 ;
  assign n1259 = x62 & ~x190 ;
  assign n1260 = x63 | x64 ;
  assign n1261 = n1259 | n1260 ;
  assign n1262 = ~n1251 & n1261 ;
  assign n1263 = ( ~n1251 & n1258 ) | ( ~n1251 & n1262 ) | ( n1258 & n1262 ) ;
  assign n1264 = ( n1247 & ~n1248 ) | ( n1247 & n1263 ) | ( ~n1248 & n1263 ) ;
  assign n1265 = ~n1236 & n1264 ;
  assign n1266 = ~n1236 & n1239 ;
  assign n1267 = ~x58 & x185 ;
  assign n1268 = x186 | x187 ;
  assign n1269 = n1267 | n1268 ;
  assign n1270 = ~n1257 & n1269 ;
  assign n1271 = n1254 & ~n1261 ;
  assign n1272 = ( ~n1261 & n1270 ) | ( ~n1261 & n1271 ) | ( n1270 & n1271 ) ;
  assign n1273 = ~n1245 & n1251 ;
  assign n1274 = n1242 | n1273 ;
  assign n1275 = ( ~n1246 & n1272 ) | ( ~n1246 & n1274 ) | ( n1272 & n1274 ) ;
  assign n1276 = ( n1236 & ~n1266 ) | ( n1236 & n1275 ) | ( ~n1266 & n1275 ) ;
  assign n1277 = ( n1233 & n1265 ) | ( n1233 & ~n1276 ) | ( n1265 & ~n1276 ) ;
  assign n1278 = ~x85 & x212 ;
  assign n1279 = x213 | x214 ;
  assign n1280 = n1278 | n1279 ;
  assign n1281 = x83 & ~x211 ;
  assign n1282 = x84 | x85 ;
  assign n1283 = n1281 | n1282 ;
  assign n1284 = ~n1280 & n1283 ;
  assign n1285 = x80 & ~x208 ;
  assign n1286 = x81 | x82 ;
  assign n1287 = n1285 | n1286 ;
  assign n1288 = ~x79 & x206 ;
  assign n1289 = x207 | x208 ;
  assign n1290 = n1288 | n1289 ;
  assign n1291 = x77 & ~x205 ;
  assign n1292 = x78 | x79 ;
  assign n1293 = n1291 | n1292 ;
  assign n1294 = ~n1290 & n1293 ;
  assign n1295 = n1287 | n1294 ;
  assign n1296 = ~n1287 & n1290 ;
  assign n1297 = ~x76 & x203 ;
  assign n1298 = x204 | x205 ;
  assign n1299 = n1297 | n1298 ;
  assign n1300 = ~x73 & x200 ;
  assign n1301 = x201 | x202 ;
  assign n1302 = n1300 | n1301 ;
  assign n1303 = x71 & ~x199 ;
  assign n1304 = x72 | x73 ;
  assign n1305 = n1303 | n1304 ;
  assign n1306 = ~n1302 & n1305 ;
  assign n1307 = x74 & ~x202 ;
  assign n1308 = x75 | x76 ;
  assign n1309 = n1307 | n1308 ;
  assign n1310 = ~n1299 & n1309 ;
  assign n1311 = ( ~n1299 & n1306 ) | ( ~n1299 & n1310 ) | ( n1306 & n1310 ) ;
  assign n1312 = ( n1295 & ~n1296 ) | ( n1295 & n1311 ) | ( ~n1296 & n1311 ) ;
  assign n1313 = ~x82 & x209 ;
  assign n1314 = x210 | x211 ;
  assign n1315 = n1313 | n1314 ;
  assign n1316 = ~n1283 & n1315 ;
  assign n1317 = n1280 | n1316 ;
  assign n1318 = ( n1284 & n1312 ) | ( n1284 & ~n1317 ) | ( n1312 & ~n1317 ) ;
  assign n1319 = n1296 | n1315 ;
  assign n1320 = n1287 & ~n1315 ;
  assign n1321 = n1302 & ~n1309 ;
  assign n1322 = ~n1293 & n1299 ;
  assign n1323 = ( ~n1293 & n1321 ) | ( ~n1293 & n1322 ) | ( n1321 & n1322 ) ;
  assign n1324 = ( n1319 & ~n1320 ) | ( n1319 & n1323 ) | ( ~n1320 & n1323 ) ;
  assign n1325 = ( n1280 & ~n1284 ) | ( n1280 & n1324 ) | ( ~n1284 & n1324 ) ;
  assign n1326 = ( n1277 & n1318 ) | ( n1277 & ~n1325 ) | ( n1318 & ~n1325 ) ;
  assign n1327 = x101 & ~x229 ;
  assign n1328 = x102 | x103 ;
  assign n1329 = n1327 | n1328 ;
  assign n1330 = ~x100 & x227 ;
  assign n1331 = x228 | x229 ;
  assign n1332 = n1330 | n1331 ;
  assign n1333 = x98 & ~x226 ;
  assign n1334 = x99 | x100 ;
  assign n1335 = n1333 | n1334 ;
  assign n1336 = ~n1332 & n1335 ;
  assign n1337 = n1329 | n1336 ;
  assign n1338 = x95 & ~x223 ;
  assign n1339 = x96 | x97 ;
  assign n1340 = n1338 | n1339 ;
  assign n1341 = ~x94 & x221 ;
  assign n1342 = x222 | x223 ;
  assign n1343 = n1341 | n1342 ;
  assign n1344 = x92 & ~x220 ;
  assign n1345 = x93 | x94 ;
  assign n1346 = n1344 | n1345 ;
  assign n1347 = ~n1343 & n1346 ;
  assign n1348 = n1340 | n1347 ;
  assign n1349 = ~n1340 & n1343 ;
  assign n1350 = ~x91 & x218 ;
  assign n1351 = x219 | x220 ;
  assign n1352 = n1350 | n1351 ;
  assign n1353 = ~x88 & x215 ;
  assign n1354 = x216 | x217 ;
  assign n1355 = n1353 | n1354 ;
  assign n1356 = x86 & ~x214 ;
  assign n1357 = x87 | x88 ;
  assign n1358 = n1356 | n1357 ;
  assign n1359 = ~n1355 & n1358 ;
  assign n1360 = x89 & ~x217 ;
  assign n1361 = x90 | x91 ;
  assign n1362 = n1360 | n1361 ;
  assign n1363 = ~n1352 & n1362 ;
  assign n1364 = ( ~n1352 & n1359 ) | ( ~n1352 & n1363 ) | ( n1359 & n1363 ) ;
  assign n1365 = ( n1348 & ~n1349 ) | ( n1348 & n1364 ) | ( ~n1349 & n1364 ) ;
  assign n1366 = ~x97 & x224 ;
  assign n1367 = x225 | x226 ;
  assign n1368 = n1366 | n1367 ;
  assign n1369 = ~n1335 & n1368 ;
  assign n1370 = n1332 | n1369 ;
  assign n1371 = ~n1329 & n1370 ;
  assign n1372 = ( n1337 & n1365 ) | ( n1337 & ~n1371 ) | ( n1365 & ~n1371 ) ;
  assign n1373 = ~n1329 & n1332 ;
  assign n1374 = n1349 | n1368 ;
  assign n1375 = n1340 & ~n1368 ;
  assign n1376 = n1355 & ~n1362 ;
  assign n1377 = ~n1346 & n1352 ;
  assign n1378 = ( ~n1346 & n1376 ) | ( ~n1346 & n1377 ) | ( n1376 & n1377 ) ;
  assign n1379 = ( n1374 & ~n1375 ) | ( n1374 & n1378 ) | ( ~n1375 & n1378 ) ;
  assign n1380 = ( ~n1337 & n1373 ) | ( ~n1337 & n1379 ) | ( n1373 & n1379 ) ;
  assign n1381 = ( n1326 & n1372 ) | ( n1326 & ~n1380 ) | ( n1372 & ~n1380 ) ;
  assign n1382 = ~x118 & x245 ;
  assign n1383 = x246 | x247 ;
  assign n1384 = n1382 | n1383 ;
  assign n1385 = x116 & ~x244 ;
  assign n1386 = x117 | x118 ;
  assign n1387 = n1385 | n1386 ;
  assign n1388 = ~x115 & x242 ;
  assign n1389 = x243 | x244 ;
  assign n1390 = n1388 | n1389 ;
  assign n1391 = x113 & ~x241 ;
  assign n1392 = x114 | x115 ;
  assign n1393 = n1391 | n1392 ;
  assign n1394 = ~n1390 & n1393 ;
  assign n1395 = ~x112 & x239 ;
  assign n1396 = x240 | x241 ;
  assign n1397 = n1395 | n1396 ;
  assign n1398 = ~x109 & x236 ;
  assign n1399 = x237 | x238 ;
  assign n1400 = n1398 | n1399 ;
  assign n1401 = x110 & ~x238 ;
  assign n1402 = x111 | x112 ;
  assign n1403 = n1401 | n1402 ;
  assign n1404 = n1400 & ~n1403 ;
  assign n1405 = n1397 | n1404 ;
  assign n1406 = ~n1397 & n1403 ;
  assign n1407 = ~x103 & x230 ;
  assign n1408 = x231 | x232 ;
  assign n1409 = n1407 | n1408 ;
  assign n1410 = x104 & ~x232 ;
  assign n1411 = x105 | x106 ;
  assign n1412 = n1410 | n1411 ;
  assign n1413 = n1409 & ~n1412 ;
  assign n1414 = x107 & ~x235 ;
  assign n1415 = x108 | x109 ;
  assign n1416 = n1414 | n1415 ;
  assign n1417 = ~x106 & x233 ;
  assign n1418 = x234 | x235 ;
  assign n1419 = n1417 | n1418 ;
  assign n1420 = ~n1416 & n1419 ;
  assign n1421 = ( n1413 & ~n1416 ) | ( n1413 & n1420 ) | ( ~n1416 & n1420 ) ;
  assign n1422 = ( n1405 & ~n1406 ) | ( n1405 & n1421 ) | ( ~n1406 & n1421 ) ;
  assign n1423 = ( n1390 & ~n1394 ) | ( n1390 & n1422 ) | ( ~n1394 & n1422 ) ;
  assign n1424 = ~n1387 & n1423 ;
  assign n1425 = n1384 | n1424 ;
  assign n1426 = x119 & ~x247 ;
  assign n1427 = x120 | x121 ;
  assign n1428 = n1426 | n1427 ;
  assign n1429 = n1425 & ~n1428 ;
  assign n1430 = ~n1384 & n1387 ;
  assign n1431 = n1393 | n1406 ;
  assign n1432 = ~n1393 & n1397 ;
  assign n1433 = n1412 & ~n1419 ;
  assign n1434 = ~n1400 & n1416 ;
  assign n1435 = ( ~n1400 & n1433 ) | ( ~n1400 & n1434 ) | ( n1433 & n1434 ) ;
  assign n1436 = ( n1431 & ~n1432 ) | ( n1431 & n1435 ) | ( ~n1432 & n1435 ) ;
  assign n1437 = ~n1387 & n1390 ;
  assign n1438 = n1384 | n1437 ;
  assign n1439 = ( n1430 & n1436 ) | ( n1430 & ~n1438 ) | ( n1436 & ~n1438 ) ;
  assign n1440 = n1428 | n1439 ;
  assign n1441 = ( n1381 & ~n1429 ) | ( n1381 & n1440 ) | ( ~n1429 & n1440 ) ;
  assign n1442 = x0 & ~x128 ;
  assign n1443 = x1 | x2 ;
  assign n1444 = n1442 | n1443 ;
  assign n1445 = ~x127 & x254 ;
  assign n1446 = x128 | x255 ;
  assign n1447 = n1445 | n1446 ;
  assign n1448 = ~x124 & x251 ;
  assign n1449 = x252 | x253 ;
  assign n1450 = n1448 | n1449 ;
  assign n1451 = x122 & ~x250 ;
  assign n1452 = x123 | x124 ;
  assign n1453 = n1451 | n1452 ;
  assign n1454 = ~n1450 & n1453 ;
  assign n1455 = x125 & ~x253 ;
  assign n1456 = x126 | x127 ;
  assign n1457 = n1455 | n1456 ;
  assign n1458 = ~n1447 & n1457 ;
  assign n1459 = ( ~n1447 & n1454 ) | ( ~n1447 & n1458 ) | ( n1454 & n1458 ) ;
  assign n1460 = n1444 | n1459 ;
  assign n1461 = ~n1444 & n1447 ;
  assign n1462 = ~x121 & x248 ;
  assign n1463 = x249 | x250 ;
  assign n1464 = n1462 | n1463 ;
  assign n1465 = ~n1453 & n1464 ;
  assign n1466 = n1450 & ~n1457 ;
  assign n1467 = ( ~n1457 & n1465 ) | ( ~n1457 & n1466 ) | ( n1465 & n1466 ) ;
  assign n1468 = ( ~n1444 & n1461 ) | ( ~n1444 & n1467 ) | ( n1461 & n1467 ) ;
  assign n1469 = ( n1441 & n1460 ) | ( n1441 & ~n1468 ) | ( n1460 & ~n1468 ) ;
  assign n1470 = n1068 & n1469 ;
  assign n1471 = ~x3 & x130 ;
  assign n1472 = x131 & ~n1471 ;
  assign n1473 = x5 | n671 ;
  assign n1474 = ~n264 & n1473 ;
  assign n1475 = ( ~n273 & n277 ) | ( ~n273 & n1474 ) | ( n277 & n1474 ) ;
  assign n1476 = n280 & ~n297 ;
  assign n1477 = n292 | n1476 ;
  assign n1478 = ( ~n298 & n1475 ) | ( ~n298 & n1477 ) | ( n1475 & n1477 ) ;
  assign n1479 = n286 & ~n307 ;
  assign n1480 = n310 | n1479 ;
  assign n1481 = ( n299 & ~n310 ) | ( n299 & n311 ) | ( ~n310 & n311 ) ;
  assign n1482 = ( n1478 & n1480 ) | ( n1478 & ~n1481 ) | ( n1480 & ~n1481 ) ;
  assign n1483 = n304 & ~n347 ;
  assign n1484 = ( n318 & ~n347 ) | ( n318 & n1483 ) | ( ~n347 & n1483 ) ;
  assign n1485 = n333 | n1484 ;
  assign n1486 = ( n322 & ~n333 ) | ( n322 & n348 ) | ( ~n333 & n348 ) ;
  assign n1487 = ( n1482 & ~n1485 ) | ( n1482 & n1486 ) | ( ~n1485 & n1486 ) ;
  assign n1488 = n327 & ~n380 ;
  assign n1489 = ( n341 & ~n380 ) | ( n341 & n1488 ) | ( ~n380 & n1488 ) ;
  assign n1490 = n365 | n1489 ;
  assign n1491 = ( ~n327 & n344 ) | ( ~n327 & n349 ) | ( n344 & n349 ) ;
  assign n1492 = ( ~n365 & n381 ) | ( ~n365 & n1491 ) | ( n381 & n1491 ) ;
  assign n1493 = ( n1487 & ~n1490 ) | ( n1487 & n1492 ) | ( ~n1490 & n1492 ) ;
  assign n1494 = ( ~n355 & n359 ) | ( ~n355 & n373 ) | ( n359 & n373 ) ;
  assign n1495 = ( ~n401 & n402 ) | ( ~n401 & n1494 ) | ( n402 & n1494 ) ;
  assign n1496 = n355 & ~n398 ;
  assign n1497 = n401 | n1496 ;
  assign n1498 = ( ~n358 & n376 ) | ( ~n358 & n382 ) | ( n376 & n382 ) ;
  assign n1499 = ( ~n402 & n1497 ) | ( ~n402 & n1498 ) | ( n1497 & n1498 ) ;
  assign n1500 = ( n1493 & ~n1495 ) | ( n1493 & n1499 ) | ( ~n1495 & n1499 ) ;
  assign n1501 = n388 & ~n460 ;
  assign n1502 = ( ~n394 & n409 ) | ( ~n394 & n414 ) | ( n409 & n414 ) ;
  assign n1503 = n419 | n460 ;
  assign n1504 = ( ~n1501 & n1502 ) | ( ~n1501 & n1503 ) | ( n1502 & n1503 ) ;
  assign n1505 = ~n448 & n1504 ;
  assign n1506 = n448 | n1501 ;
  assign n1507 = ( ~n391 & n395 ) | ( ~n391 & n421 ) | ( n395 & n421 ) ;
  assign n1508 = ( ~n461 & n1506 ) | ( ~n461 & n1507 ) | ( n1506 & n1507 ) ;
  assign n1509 = ( n1500 & ~n1505 ) | ( n1500 & n1508 ) | ( ~n1505 & n1508 ) ;
  assign n1510 = n457 | n496 ;
  assign n1511 = n427 & ~n496 ;
  assign n1512 = ( ~n433 & n437 ) | ( ~n433 & n453 ) | ( n437 & n453 ) ;
  assign n1513 = ( n1510 & ~n1511 ) | ( n1510 & n1512 ) | ( ~n1511 & n1512 ) ;
  assign n1514 = ~n493 & n1513 ;
  assign n1515 = ( ~n436 & n462 ) | ( ~n436 & n464 ) | ( n462 & n464 ) ;
  assign n1516 = n427 | n439 ;
  assign n1517 = ( ~n457 & n1515 ) | ( ~n457 & n1516 ) | ( n1515 & n1516 ) ;
  assign n1518 = ( n493 & ~n497 ) | ( n493 & n1517 ) | ( ~n497 & n1517 ) ;
  assign n1519 = ( n1509 & n1514 ) | ( n1509 & ~n1518 ) | ( n1514 & ~n1518 ) ;
  assign n1520 = n474 | n511 ;
  assign n1521 = ( ~n481 & n485 ) | ( ~n481 & n501 ) | ( n485 & n501 ) ;
  assign n1522 = ( ~n507 & n1520 ) | ( ~n507 & n1521 ) | ( n1520 & n1521 ) ;
  assign n1523 = n471 & ~n549 ;
  assign n1524 = n546 | n1523 ;
  assign n1525 = ( n550 & n1522 ) | ( n550 & ~n1524 ) | ( n1522 & ~n1524 ) ;
  assign n1526 = ( ~n478 & n487 ) | ( ~n478 & n513 ) | ( n487 & n513 ) ;
  assign n1527 = ( ~n475 & n508 ) | ( ~n475 & n1526 ) | ( n508 & n1526 ) ;
  assign n1528 = ( n546 & ~n550 ) | ( n546 & n1527 ) | ( ~n550 & n1527 ) ;
  assign n1529 = ( n1519 & n1525 ) | ( n1519 & ~n1528 ) | ( n1525 & ~n1528 ) ;
  assign n1530 = n520 & ~n600 ;
  assign n1531 = n603 | n1530 ;
  assign n1532 = n526 | n566 ;
  assign n1533 = ( ~n534 & n538 ) | ( ~n534 & n554 ) | ( n538 & n554 ) ;
  assign n1534 = ( ~n560 & n1532 ) | ( ~n560 & n1533 ) | ( n1532 & n1533 ) ;
  assign n1535 = n564 | n600 ;
  assign n1536 = ~n603 & n1535 ;
  assign n1537 = ( n1531 & n1534 ) | ( n1531 & ~n1536 ) | ( n1534 & ~n1536 ) ;
  assign n1538 = ( ~n531 & n540 ) | ( ~n531 & n568 ) | ( n540 & n568 ) ;
  assign n1539 = ( ~n527 & n561 ) | ( ~n527 & n1538 ) | ( n561 & n1538 ) ;
  assign n1540 = ( n604 & ~n1531 ) | ( n604 & n1539 ) | ( ~n1531 & n1539 ) ;
  assign n1541 = ( n1529 & n1537 ) | ( n1529 & ~n1540 ) | ( n1537 & ~n1540 ) ;
  assign n1542 = n581 | n623 ;
  assign n1543 = ( ~n594 & n595 ) | ( ~n594 & n611 ) | ( n595 & n611 ) ;
  assign n1544 = ( ~n585 & n1542 ) | ( ~n585 & n1543 ) | ( n1542 & n1543 ) ;
  assign n1545 = ( n575 & ~n621 ) | ( n575 & n1544 ) | ( ~n621 & n1544 ) ;
  assign n1546 = ~n619 & n1545 ;
  assign n1547 = n655 | n1546 ;
  assign n1548 = ~n644 & n1547 ;
  assign n1549 = n575 & ~n619 ;
  assign n1550 = n655 | n1549 ;
  assign n1551 = n619 & ~n655 ;
  assign n1552 = n578 | n585 ;
  assign n1553 = ( ~n588 & n597 ) | ( ~n588 & n625 ) | ( n597 & n625 ) ;
  assign n1554 = ( ~n628 & n1552 ) | ( ~n628 & n1553 ) | ( n1552 & n1553 ) ;
  assign n1555 = ( ~n1550 & n1551 ) | ( ~n1550 & n1554 ) | ( n1551 & n1554 ) ;
  assign n1556 = n644 | n1555 ;
  assign n1557 = ( n1541 & ~n1548 ) | ( n1541 & n1556 ) | ( ~n1548 & n1556 ) ;
  assign n1558 = x2 | x3 ;
  assign n1559 = n259 | n1558 ;
  assign n1560 = x128 | x129 ;
  assign n1561 = n257 | n1560 ;
  assign n1562 = n635 & ~n1561 ;
  assign n1563 = ( n649 & ~n1561 ) | ( n649 & n1562 ) | ( ~n1561 & n1562 ) ;
  assign n1564 = n1559 | n1563 ;
  assign n1565 = ~n1559 & n1561 ;
  assign n1566 = ( ~n635 & n652 ) | ( ~n635 & n657 ) | ( n652 & n657 ) ;
  assign n1567 = ( ~n1559 & n1565 ) | ( ~n1559 & n1566 ) | ( n1565 & n1566 ) ;
  assign n1568 = ( n1557 & n1564 ) | ( n1557 & ~n1567 ) | ( n1564 & ~n1567 ) ;
  assign n1569 = n1472 & n1568 ;
  assign n1570 = ~x4 & x131 ;
  assign n1571 = x132 & ~n1570 ;
  assign n1572 = x6 | n1075 ;
  assign n1573 = ~n669 & n1572 ;
  assign n1574 = ( ~n678 & n682 ) | ( ~n678 & n1573 ) | ( n682 & n1573 ) ;
  assign n1575 = n685 & ~n702 ;
  assign n1576 = n697 | n1575 ;
  assign n1577 = ( ~n703 & n1574 ) | ( ~n703 & n1576 ) | ( n1574 & n1576 ) ;
  assign n1578 = n691 & ~n712 ;
  assign n1579 = n715 | n1578 ;
  assign n1580 = ( n704 & ~n715 ) | ( n704 & n716 ) | ( ~n715 & n716 ) ;
  assign n1581 = ( n1577 & n1579 ) | ( n1577 & ~n1580 ) | ( n1579 & ~n1580 ) ;
  assign n1582 = n709 & ~n752 ;
  assign n1583 = ( n723 & ~n752 ) | ( n723 & n1582 ) | ( ~n752 & n1582 ) ;
  assign n1584 = n738 | n1583 ;
  assign n1585 = ( n727 & ~n738 ) | ( n727 & n753 ) | ( ~n738 & n753 ) ;
  assign n1586 = ( n1581 & ~n1584 ) | ( n1581 & n1585 ) | ( ~n1584 & n1585 ) ;
  assign n1587 = n732 & ~n785 ;
  assign n1588 = ( n746 & ~n785 ) | ( n746 & n1587 ) | ( ~n785 & n1587 ) ;
  assign n1589 = n770 | n1588 ;
  assign n1590 = ( ~n732 & n749 ) | ( ~n732 & n754 ) | ( n749 & n754 ) ;
  assign n1591 = ( ~n770 & n786 ) | ( ~n770 & n1590 ) | ( n786 & n1590 ) ;
  assign n1592 = ( n1586 & ~n1589 ) | ( n1586 & n1591 ) | ( ~n1589 & n1591 ) ;
  assign n1593 = ( ~n760 & n764 ) | ( ~n760 & n778 ) | ( n764 & n778 ) ;
  assign n1594 = ( ~n806 & n807 ) | ( ~n806 & n1593 ) | ( n807 & n1593 ) ;
  assign n1595 = n760 & ~n803 ;
  assign n1596 = n806 | n1595 ;
  assign n1597 = ( ~n763 & n781 ) | ( ~n763 & n787 ) | ( n781 & n787 ) ;
  assign n1598 = ( ~n807 & n1596 ) | ( ~n807 & n1597 ) | ( n1596 & n1597 ) ;
  assign n1599 = ( n1592 & ~n1594 ) | ( n1592 & n1598 ) | ( ~n1594 & n1598 ) ;
  assign n1600 = n793 & ~n865 ;
  assign n1601 = ( ~n799 & n814 ) | ( ~n799 & n819 ) | ( n814 & n819 ) ;
  assign n1602 = n824 | n865 ;
  assign n1603 = ( ~n1600 & n1601 ) | ( ~n1600 & n1602 ) | ( n1601 & n1602 ) ;
  assign n1604 = ~n853 & n1603 ;
  assign n1605 = n853 | n1600 ;
  assign n1606 = ( ~n796 & n800 ) | ( ~n796 & n826 ) | ( n800 & n826 ) ;
  assign n1607 = ( ~n866 & n1605 ) | ( ~n866 & n1606 ) | ( n1605 & n1606 ) ;
  assign n1608 = ( n1599 & ~n1604 ) | ( n1599 & n1607 ) | ( ~n1604 & n1607 ) ;
  assign n1609 = n862 | n901 ;
  assign n1610 = n832 & ~n901 ;
  assign n1611 = ( ~n838 & n842 ) | ( ~n838 & n858 ) | ( n842 & n858 ) ;
  assign n1612 = ( n1609 & ~n1610 ) | ( n1609 & n1611 ) | ( ~n1610 & n1611 ) ;
  assign n1613 = ~n898 & n1612 ;
  assign n1614 = ( ~n841 & n867 ) | ( ~n841 & n869 ) | ( n867 & n869 ) ;
  assign n1615 = n832 | n844 ;
  assign n1616 = ( ~n862 & n1614 ) | ( ~n862 & n1615 ) | ( n1614 & n1615 ) ;
  assign n1617 = ( n898 & ~n902 ) | ( n898 & n1616 ) | ( ~n902 & n1616 ) ;
  assign n1618 = ( n1608 & n1613 ) | ( n1608 & ~n1617 ) | ( n1613 & ~n1617 ) ;
  assign n1619 = n879 | n916 ;
  assign n1620 = ( ~n886 & n890 ) | ( ~n886 & n906 ) | ( n890 & n906 ) ;
  assign n1621 = ( ~n912 & n1619 ) | ( ~n912 & n1620 ) | ( n1619 & n1620 ) ;
  assign n1622 = n876 & ~n954 ;
  assign n1623 = n951 | n1622 ;
  assign n1624 = ( n955 & n1621 ) | ( n955 & ~n1623 ) | ( n1621 & ~n1623 ) ;
  assign n1625 = ( ~n883 & n892 ) | ( ~n883 & n918 ) | ( n892 & n918 ) ;
  assign n1626 = ( ~n880 & n913 ) | ( ~n880 & n1625 ) | ( n913 & n1625 ) ;
  assign n1627 = ( n951 & ~n955 ) | ( n951 & n1626 ) | ( ~n955 & n1626 ) ;
  assign n1628 = ( n1618 & n1624 ) | ( n1618 & ~n1627 ) | ( n1624 & ~n1627 ) ;
  assign n1629 = n925 & ~n1005 ;
  assign n1630 = n1008 | n1629 ;
  assign n1631 = n931 | n971 ;
  assign n1632 = ( ~n939 & n943 ) | ( ~n939 & n959 ) | ( n943 & n959 ) ;
  assign n1633 = ( ~n965 & n1631 ) | ( ~n965 & n1632 ) | ( n1631 & n1632 ) ;
  assign n1634 = n969 | n1005 ;
  assign n1635 = ~n1008 & n1634 ;
  assign n1636 = ( n1630 & n1633 ) | ( n1630 & ~n1635 ) | ( n1633 & ~n1635 ) ;
  assign n1637 = ( ~n936 & n945 ) | ( ~n936 & n973 ) | ( n945 & n973 ) ;
  assign n1638 = ( ~n932 & n966 ) | ( ~n932 & n1637 ) | ( n966 & n1637 ) ;
  assign n1639 = ( n1009 & ~n1630 ) | ( n1009 & n1638 ) | ( ~n1630 & n1638 ) ;
  assign n1640 = ( n1628 & n1636 ) | ( n1628 & ~n1639 ) | ( n1636 & ~n1639 ) ;
  assign n1641 = n986 | n1028 ;
  assign n1642 = ( ~n999 & n1000 ) | ( ~n999 & n1016 ) | ( n1000 & n1016 ) ;
  assign n1643 = ( ~n990 & n1641 ) | ( ~n990 & n1642 ) | ( n1641 & n1642 ) ;
  assign n1644 = ( n980 & ~n1026 ) | ( n980 & n1643 ) | ( ~n1026 & n1643 ) ;
  assign n1645 = ~n1024 & n1644 ;
  assign n1646 = n1060 | n1645 ;
  assign n1647 = ~n1049 & n1646 ;
  assign n1648 = n980 & ~n1024 ;
  assign n1649 = n1060 | n1648 ;
  assign n1650 = n1024 & ~n1060 ;
  assign n1651 = n983 | n990 ;
  assign n1652 = ( ~n993 & n1002 ) | ( ~n993 & n1030 ) | ( n1002 & n1030 ) ;
  assign n1653 = ( ~n1033 & n1651 ) | ( ~n1033 & n1652 ) | ( n1651 & n1652 ) ;
  assign n1654 = ( ~n1649 & n1650 ) | ( ~n1649 & n1653 ) | ( n1650 & n1653 ) ;
  assign n1655 = n1049 | n1654 ;
  assign n1656 = ( n1640 & ~n1647 ) | ( n1640 & n1655 ) | ( ~n1647 & n1655 ) ;
  assign n1657 = x3 | x4 ;
  assign n1658 = n664 | n1657 ;
  assign n1659 = x129 | x130 ;
  assign n1660 = n662 | n1659 ;
  assign n1661 = n1040 & ~n1660 ;
  assign n1662 = ( n1054 & ~n1660 ) | ( n1054 & n1661 ) | ( ~n1660 & n1661 ) ;
  assign n1663 = n1658 | n1662 ;
  assign n1664 = ~n1658 & n1660 ;
  assign n1665 = ( ~n1040 & n1057 ) | ( ~n1040 & n1062 ) | ( n1057 & n1062 ) ;
  assign n1666 = ( ~n1658 & n1664 ) | ( ~n1658 & n1665 ) | ( n1664 & n1665 ) ;
  assign n1667 = ( n1656 & n1663 ) | ( n1656 & ~n1666 ) | ( n1663 & ~n1666 ) ;
  assign n1668 = n1571 & n1667 ;
  assign n1669 = x133 & ~n263 ;
  assign n1670 = x7 | n274 ;
  assign n1671 = ~n1073 & n1670 ;
  assign n1672 = ( ~n1082 & n1086 ) | ( ~n1082 & n1671 ) | ( n1086 & n1671 ) ;
  assign n1673 = n1089 & ~n1106 ;
  assign n1674 = n1101 | n1673 ;
  assign n1675 = ( ~n1107 & n1672 ) | ( ~n1107 & n1674 ) | ( n1672 & n1674 ) ;
  assign n1676 = n1095 & ~n1116 ;
  assign n1677 = n1119 | n1676 ;
  assign n1678 = ( n1108 & ~n1119 ) | ( n1108 & n1120 ) | ( ~n1119 & n1120 ) ;
  assign n1679 = ( n1675 & n1677 ) | ( n1675 & ~n1678 ) | ( n1677 & ~n1678 ) ;
  assign n1680 = n1113 & ~n1156 ;
  assign n1681 = ( n1127 & ~n1156 ) | ( n1127 & n1680 ) | ( ~n1156 & n1680 ) ;
  assign n1682 = n1142 | n1681 ;
  assign n1683 = ( n1131 & ~n1142 ) | ( n1131 & n1157 ) | ( ~n1142 & n1157 ) ;
  assign n1684 = ( n1679 & ~n1682 ) | ( n1679 & n1683 ) | ( ~n1682 & n1683 ) ;
  assign n1685 = n1136 & ~n1189 ;
  assign n1686 = ( n1150 & ~n1189 ) | ( n1150 & n1685 ) | ( ~n1189 & n1685 ) ;
  assign n1687 = n1174 | n1686 ;
  assign n1688 = ( ~n1136 & n1153 ) | ( ~n1136 & n1158 ) | ( n1153 & n1158 ) ;
  assign n1689 = ( ~n1174 & n1190 ) | ( ~n1174 & n1688 ) | ( n1190 & n1688 ) ;
  assign n1690 = ( n1684 & ~n1687 ) | ( n1684 & n1689 ) | ( ~n1687 & n1689 ) ;
  assign n1691 = ( ~n1164 & n1168 ) | ( ~n1164 & n1182 ) | ( n1168 & n1182 ) ;
  assign n1692 = ( ~n1210 & n1211 ) | ( ~n1210 & n1691 ) | ( n1211 & n1691 ) ;
  assign n1693 = n1164 & ~n1207 ;
  assign n1694 = n1210 | n1693 ;
  assign n1695 = ( ~n1167 & n1185 ) | ( ~n1167 & n1191 ) | ( n1185 & n1191 ) ;
  assign n1696 = ( ~n1211 & n1694 ) | ( ~n1211 & n1695 ) | ( n1694 & n1695 ) ;
  assign n1697 = ( n1690 & ~n1692 ) | ( n1690 & n1696 ) | ( ~n1692 & n1696 ) ;
  assign n1698 = n1197 & ~n1269 ;
  assign n1699 = ( ~n1203 & n1218 ) | ( ~n1203 & n1223 ) | ( n1218 & n1223 ) ;
  assign n1700 = n1228 | n1269 ;
  assign n1701 = ( ~n1698 & n1699 ) | ( ~n1698 & n1700 ) | ( n1699 & n1700 ) ;
  assign n1702 = ~n1257 & n1701 ;
  assign n1703 = n1257 | n1698 ;
  assign n1704 = ( ~n1200 & n1204 ) | ( ~n1200 & n1230 ) | ( n1204 & n1230 ) ;
  assign n1705 = ( ~n1270 & n1703 ) | ( ~n1270 & n1704 ) | ( n1703 & n1704 ) ;
  assign n1706 = ( n1697 & ~n1702 ) | ( n1697 & n1705 ) | ( ~n1702 & n1705 ) ;
  assign n1707 = n1266 | n1305 ;
  assign n1708 = n1236 & ~n1305 ;
  assign n1709 = ( ~n1242 & n1246 ) | ( ~n1242 & n1262 ) | ( n1246 & n1262 ) ;
  assign n1710 = ( n1707 & ~n1708 ) | ( n1707 & n1709 ) | ( ~n1708 & n1709 ) ;
  assign n1711 = ~n1302 & n1710 ;
  assign n1712 = ( ~n1245 & n1271 ) | ( ~n1245 & n1273 ) | ( n1271 & n1273 ) ;
  assign n1713 = n1236 | n1248 ;
  assign n1714 = ( ~n1266 & n1712 ) | ( ~n1266 & n1713 ) | ( n1712 & n1713 ) ;
  assign n1715 = ( n1302 & ~n1306 ) | ( n1302 & n1714 ) | ( ~n1306 & n1714 ) ;
  assign n1716 = ( n1706 & n1711 ) | ( n1706 & ~n1715 ) | ( n1711 & ~n1715 ) ;
  assign n1717 = n1283 | n1320 ;
  assign n1718 = ( ~n1290 & n1294 ) | ( ~n1290 & n1310 ) | ( n1294 & n1310 ) ;
  assign n1719 = ( ~n1316 & n1717 ) | ( ~n1316 & n1718 ) | ( n1717 & n1718 ) ;
  assign n1720 = n1280 & ~n1358 ;
  assign n1721 = n1355 | n1720 ;
  assign n1722 = ( n1359 & n1719 ) | ( n1359 & ~n1721 ) | ( n1719 & ~n1721 ) ;
  assign n1723 = ( ~n1287 & n1296 ) | ( ~n1287 & n1322 ) | ( n1296 & n1322 ) ;
  assign n1724 = ( ~n1284 & n1317 ) | ( ~n1284 & n1723 ) | ( n1317 & n1723 ) ;
  assign n1725 = ( n1355 & ~n1359 ) | ( n1355 & n1724 ) | ( ~n1359 & n1724 ) ;
  assign n1726 = ( n1716 & n1722 ) | ( n1716 & ~n1725 ) | ( n1722 & ~n1725 ) ;
  assign n1727 = n1329 & ~n1409 ;
  assign n1728 = n1412 | n1727 ;
  assign n1729 = n1335 | n1375 ;
  assign n1730 = ( ~n1343 & n1347 ) | ( ~n1343 & n1363 ) | ( n1347 & n1363 ) ;
  assign n1731 = ( ~n1369 & n1729 ) | ( ~n1369 & n1730 ) | ( n1729 & n1730 ) ;
  assign n1732 = n1373 | n1409 ;
  assign n1733 = ~n1412 & n1732 ;
  assign n1734 = ( n1728 & n1731 ) | ( n1728 & ~n1733 ) | ( n1731 & ~n1733 ) ;
  assign n1735 = ( ~n1340 & n1349 ) | ( ~n1340 & n1377 ) | ( n1349 & n1377 ) ;
  assign n1736 = ( ~n1336 & n1370 ) | ( ~n1336 & n1735 ) | ( n1370 & n1735 ) ;
  assign n1737 = ( n1413 & ~n1728 ) | ( n1413 & n1736 ) | ( ~n1728 & n1736 ) ;
  assign n1738 = ( n1726 & n1734 ) | ( n1726 & ~n1737 ) | ( n1734 & ~n1737 ) ;
  assign n1739 = n1390 | n1432 ;
  assign n1740 = ( ~n1403 & n1404 ) | ( ~n1403 & n1420 ) | ( n1404 & n1420 ) ;
  assign n1741 = ( ~n1394 & n1739 ) | ( ~n1394 & n1740 ) | ( n1739 & n1740 ) ;
  assign n1742 = ( n1384 & ~n1430 ) | ( n1384 & n1741 ) | ( ~n1430 & n1741 ) ;
  assign n1743 = ~n1428 & n1742 ;
  assign n1744 = n1464 | n1743 ;
  assign n1745 = ~n1453 & n1744 ;
  assign n1746 = n1384 & ~n1428 ;
  assign n1747 = n1464 | n1746 ;
  assign n1748 = n1428 & ~n1464 ;
  assign n1749 = n1387 | n1394 ;
  assign n1750 = ( ~n1397 & n1406 ) | ( ~n1397 & n1434 ) | ( n1406 & n1434 ) ;
  assign n1751 = ( ~n1437 & n1749 ) | ( ~n1437 & n1750 ) | ( n1749 & n1750 ) ;
  assign n1752 = ( ~n1747 & n1748 ) | ( ~n1747 & n1751 ) | ( n1748 & n1751 ) ;
  assign n1753 = n1453 | n1752 ;
  assign n1754 = ( n1738 & ~n1745 ) | ( n1738 & n1753 ) | ( ~n1745 & n1753 ) ;
  assign n1755 = n261 | n1067 ;
  assign n1756 = n1444 & ~n1755 ;
  assign n1757 = ( n1458 & ~n1755 ) | ( n1458 & n1756 ) | ( ~n1755 & n1756 ) ;
  assign n1758 = n268 | n1757 ;
  assign n1759 = ~n268 & n1755 ;
  assign n1760 = ( ~n1444 & n1461 ) | ( ~n1444 & n1466 ) | ( n1461 & n1466 ) ;
  assign n1761 = ( ~n268 & n1759 ) | ( ~n268 & n1760 ) | ( n1759 & n1760 ) ;
  assign n1762 = ( n1754 & n1758 ) | ( n1754 & ~n1761 ) | ( n1758 & ~n1761 ) ;
  assign n1763 = n1669 & n1762 ;
  assign n1764 = x134 & ~n668 ;
  assign n1765 = n314 | n321 ;
  assign n1766 = x8 | n679 ;
  assign n1767 = ~n272 & n1766 ;
  assign n1768 = ( ~n297 & n1476 ) | ( ~n297 & n1767 ) | ( n1476 & n1767 ) ;
  assign n1769 = ( n294 & ~n299 ) | ( n294 & n1768 ) | ( ~n299 & n1768 ) ;
  assign n1770 = ( ~n319 & n1765 ) | ( ~n319 & n1769 ) | ( n1765 & n1769 ) ;
  assign n1771 = ( ~n336 & n337 ) | ( ~n336 & n1483 ) | ( n337 & n1483 ) ;
  assign n1772 = n340 | n1771 ;
  assign n1773 = ( n350 & n1770 ) | ( n350 & ~n1772 ) | ( n1770 & ~n1772 ) ;
  assign n1774 = ( ~n368 & n369 ) | ( ~n368 & n1488 ) | ( n369 & n1488 ) ;
  assign n1775 = n372 | n1774 ;
  assign n1776 = ( n344 & ~n365 ) | ( n344 & n381 ) | ( ~n365 & n381 ) ;
  assign n1777 = ( ~n372 & n382 ) | ( ~n372 & n1776 ) | ( n382 & n1776 ) ;
  assign n1778 = ( n1773 & ~n1775 ) | ( n1773 & n1777 ) | ( ~n1775 & n1777 ) ;
  assign n1779 = ( n359 & ~n401 ) | ( n359 & n402 ) | ( ~n401 & n402 ) ;
  assign n1780 = ( ~n405 & n409 ) | ( ~n405 & n1779 ) | ( n409 & n1779 ) ;
  assign n1781 = n405 | n420 ;
  assign n1782 = ( n376 & ~n398 ) | ( n376 & n1496 ) | ( ~n398 & n1496 ) ;
  assign n1783 = ( ~n409 & n1781 ) | ( ~n409 & n1782 ) | ( n1781 & n1782 ) ;
  assign n1784 = ( n1778 & ~n1780 ) | ( n1778 & n1783 ) | ( ~n1780 & n1783 ) ;
  assign n1785 = ( ~n388 & n414 ) | ( ~n388 & n419 ) | ( n414 & n419 ) ;
  assign n1786 = n445 | n461 ;
  assign n1787 = ( ~n449 & n1785 ) | ( ~n449 & n1786 ) | ( n1785 & n1786 ) ;
  assign n1788 = ~n452 & n1787 ;
  assign n1789 = n449 | n452 ;
  assign n1790 = ( n395 & ~n460 ) | ( n395 & n1501 ) | ( ~n460 & n1501 ) ;
  assign n1791 = ( ~n462 & n1789 ) | ( ~n462 & n1790 ) | ( n1789 & n1790 ) ;
  assign n1792 = ( n1784 & ~n1788 ) | ( n1784 & n1791 ) | ( ~n1788 & n1791 ) ;
  assign n1793 = n497 | n500 ;
  assign n1794 = ( ~n427 & n437 ) | ( ~n427 & n457 ) | ( n437 & n457 ) ;
  assign n1795 = ( ~n512 & n1793 ) | ( ~n512 & n1794 ) | ( n1793 & n1794 ) ;
  assign n1796 = ~n490 & n1795 ;
  assign n1797 = ( ~n430 & n439 ) | ( ~n430 & n464 ) | ( n439 & n464 ) ;
  assign n1798 = n493 | n1511 ;
  assign n1799 = ( ~n497 & n1797 ) | ( ~n497 & n1798 ) | ( n1797 & n1798 ) ;
  assign n1800 = ( n490 & ~n501 ) | ( n490 & n1799 ) | ( ~n501 & n1799 ) ;
  assign n1801 = ( n1792 & n1796 ) | ( n1792 & ~n1800 ) | ( n1796 & ~n1800 ) ;
  assign n1802 = n543 | n567 ;
  assign n1803 = n475 | n549 ;
  assign n1804 = ( n485 & ~n506 ) | ( n485 & n511 ) | ( ~n506 & n511 ) ;
  assign n1805 = ( ~n1523 & n1803 ) | ( ~n1523 & n1804 ) | ( n1803 & n1804 ) ;
  assign n1806 = ( n554 & ~n1802 ) | ( n554 & n1805 ) | ( ~n1802 & n1805 ) ;
  assign n1807 = ( ~n474 & n487 ) | ( ~n474 & n507 ) | ( n487 & n507 ) ;
  assign n1808 = ( ~n550 & n1524 ) | ( ~n550 & n1807 ) | ( n1524 & n1807 ) ;
  assign n1809 = ( n543 & ~n554 ) | ( n543 & n1808 ) | ( ~n554 & n1808 ) ;
  assign n1810 = ( n1801 & n1806 ) | ( n1801 & ~n1809 ) | ( n1806 & ~n1809 ) ;
  assign n1811 = n607 | n624 ;
  assign n1812 = ( n538 & ~n559 ) | ( n538 & n566 ) | ( ~n559 & n566 ) ;
  assign n1813 = ( n528 & ~n564 ) | ( n528 & n1812 ) | ( ~n564 & n1812 ) ;
  assign n1814 = n604 | n610 ;
  assign n1815 = ~n607 & n1814 ;
  assign n1816 = ( n1811 & n1813 ) | ( n1811 & ~n1815 ) | ( n1813 & ~n1815 ) ;
  assign n1817 = ( ~n526 & n540 ) | ( ~n526 & n560 ) | ( n540 & n560 ) ;
  assign n1818 = ( ~n1530 & n1535 ) | ( ~n1530 & n1817 ) | ( n1535 & n1817 ) ;
  assign n1819 = ( n611 & ~n1811 ) | ( n611 & n1818 ) | ( ~n1811 & n1818 ) ;
  assign n1820 = ( n1810 & n1816 ) | ( n1810 & ~n1819 ) | ( n1816 & ~n1819 ) ;
  assign n1821 = ( ~n584 & n595 ) | ( ~n584 & n623 ) | ( n595 & n623 ) ;
  assign n1822 = ( ~n621 & n629 ) | ( ~n621 & n1821 ) | ( n629 & n1821 ) ;
  assign n1823 = ( n655 & ~n1551 ) | ( n655 & n1822 ) | ( ~n1551 & n1822 ) ;
  assign n1824 = ~n644 & n1823 ;
  assign n1825 = n641 | n1824 ;
  assign n1826 = ~n648 & n1825 ;
  assign n1827 = n645 | n648 ;
  assign n1828 = n619 | n621 ;
  assign n1829 = ( ~n581 & n585 ) | ( ~n581 & n597 ) | ( n585 & n597 ) ;
  assign n1830 = ( ~n1549 & n1828 ) | ( ~n1549 & n1829 ) | ( n1828 & n1829 ) ;
  assign n1831 = ( ~n658 & n1827 ) | ( ~n658 & n1830 ) | ( n1827 & n1830 ) ;
  assign n1832 = ( n1820 & ~n1826 ) | ( n1820 & n1831 ) | ( ~n1826 & n1831 ) ;
  assign n1833 = n666 | n1471 ;
  assign n1834 = n1559 & ~n1833 ;
  assign n1835 = ( n1562 & ~n1833 ) | ( n1562 & n1834 ) | ( ~n1833 & n1834 ) ;
  assign n1836 = n673 | n1835 ;
  assign n1837 = ~n673 & n1833 ;
  assign n1838 = ( n652 & ~n1559 ) | ( n652 & n1565 ) | ( ~n1559 & n1565 ) ;
  assign n1839 = ( ~n673 & n1837 ) | ( ~n673 & n1838 ) | ( n1837 & n1838 ) ;
  assign n1840 = ( n1832 & n1836 ) | ( n1832 & ~n1839 ) | ( n1836 & ~n1839 ) ;
  assign n1841 = n1764 & n1840 ;
  assign n1842 = x135 & ~n1072 ;
  assign n1843 = n719 | n726 ;
  assign n1844 = x9 | n1083 ;
  assign n1845 = ~n677 & n1844 ;
  assign n1846 = ( ~n702 & n1575 ) | ( ~n702 & n1845 ) | ( n1575 & n1845 ) ;
  assign n1847 = ( n699 & ~n704 ) | ( n699 & n1846 ) | ( ~n704 & n1846 ) ;
  assign n1848 = ( ~n724 & n1843 ) | ( ~n724 & n1847 ) | ( n1843 & n1847 ) ;
  assign n1849 = ( ~n741 & n742 ) | ( ~n741 & n1582 ) | ( n742 & n1582 ) ;
  assign n1850 = n745 | n1849 ;
  assign n1851 = ( n755 & n1848 ) | ( n755 & ~n1850 ) | ( n1848 & ~n1850 ) ;
  assign n1852 = ( ~n773 & n774 ) | ( ~n773 & n1587 ) | ( n774 & n1587 ) ;
  assign n1853 = n777 | n1852 ;
  assign n1854 = ( n749 & ~n770 ) | ( n749 & n786 ) | ( ~n770 & n786 ) ;
  assign n1855 = ( ~n777 & n787 ) | ( ~n777 & n1854 ) | ( n787 & n1854 ) ;
  assign n1856 = ( n1851 & ~n1853 ) | ( n1851 & n1855 ) | ( ~n1853 & n1855 ) ;
  assign n1857 = ( n764 & ~n806 ) | ( n764 & n807 ) | ( ~n806 & n807 ) ;
  assign n1858 = ( ~n810 & n814 ) | ( ~n810 & n1857 ) | ( n814 & n1857 ) ;
  assign n1859 = n810 | n825 ;
  assign n1860 = ( n781 & ~n803 ) | ( n781 & n1595 ) | ( ~n803 & n1595 ) ;
  assign n1861 = ( ~n814 & n1859 ) | ( ~n814 & n1860 ) | ( n1859 & n1860 ) ;
  assign n1862 = ( n1856 & ~n1858 ) | ( n1856 & n1861 ) | ( ~n1858 & n1861 ) ;
  assign n1863 = ( ~n793 & n819 ) | ( ~n793 & n824 ) | ( n819 & n824 ) ;
  assign n1864 = n850 | n866 ;
  assign n1865 = ( ~n854 & n1863 ) | ( ~n854 & n1864 ) | ( n1863 & n1864 ) ;
  assign n1866 = ~n857 & n1865 ;
  assign n1867 = n854 | n857 ;
  assign n1868 = ( n800 & ~n865 ) | ( n800 & n1600 ) | ( ~n865 & n1600 ) ;
  assign n1869 = ( ~n867 & n1867 ) | ( ~n867 & n1868 ) | ( n1867 & n1868 ) ;
  assign n1870 = ( n1862 & ~n1866 ) | ( n1862 & n1869 ) | ( ~n1866 & n1869 ) ;
  assign n1871 = n902 | n905 ;
  assign n1872 = ( ~n832 & n842 ) | ( ~n832 & n862 ) | ( n842 & n862 ) ;
  assign n1873 = ( ~n917 & n1871 ) | ( ~n917 & n1872 ) | ( n1871 & n1872 ) ;
  assign n1874 = ~n895 & n1873 ;
  assign n1875 = ( ~n835 & n844 ) | ( ~n835 & n869 ) | ( n844 & n869 ) ;
  assign n1876 = n898 | n1610 ;
  assign n1877 = ( ~n902 & n1875 ) | ( ~n902 & n1876 ) | ( n1875 & n1876 ) ;
  assign n1878 = ( n895 & ~n906 ) | ( n895 & n1877 ) | ( ~n906 & n1877 ) ;
  assign n1879 = ( n1870 & n1874 ) | ( n1870 & ~n1878 ) | ( n1874 & ~n1878 ) ;
  assign n1880 = n948 | n972 ;
  assign n1881 = n880 | n954 ;
  assign n1882 = ( n890 & ~n911 ) | ( n890 & n916 ) | ( ~n911 & n916 ) ;
  assign n1883 = ( ~n1622 & n1881 ) | ( ~n1622 & n1882 ) | ( n1881 & n1882 ) ;
  assign n1884 = ( n959 & ~n1880 ) | ( n959 & n1883 ) | ( ~n1880 & n1883 ) ;
  assign n1885 = ( ~n879 & n892 ) | ( ~n879 & n912 ) | ( n892 & n912 ) ;
  assign n1886 = ( ~n955 & n1623 ) | ( ~n955 & n1885 ) | ( n1623 & n1885 ) ;
  assign n1887 = ( n948 & ~n959 ) | ( n948 & n1886 ) | ( ~n959 & n1886 ) ;
  assign n1888 = ( n1879 & n1884 ) | ( n1879 & ~n1887 ) | ( n1884 & ~n1887 ) ;
  assign n1889 = n1012 | n1029 ;
  assign n1890 = ( n943 & ~n964 ) | ( n943 & n971 ) | ( ~n964 & n971 ) ;
  assign n1891 = ( n933 & ~n969 ) | ( n933 & n1890 ) | ( ~n969 & n1890 ) ;
  assign n1892 = n1009 | n1015 ;
  assign n1893 = ~n1012 & n1892 ;
  assign n1894 = ( n1889 & n1891 ) | ( n1889 & ~n1893 ) | ( n1891 & ~n1893 ) ;
  assign n1895 = ( ~n931 & n945 ) | ( ~n931 & n965 ) | ( n945 & n965 ) ;
  assign n1896 = ( ~n1629 & n1634 ) | ( ~n1629 & n1895 ) | ( n1634 & n1895 ) ;
  assign n1897 = ( n1016 & ~n1889 ) | ( n1016 & n1896 ) | ( ~n1889 & n1896 ) ;
  assign n1898 = ( n1888 & n1894 ) | ( n1888 & ~n1897 ) | ( n1894 & ~n1897 ) ;
  assign n1899 = ( ~n989 & n1000 ) | ( ~n989 & n1028 ) | ( n1000 & n1028 ) ;
  assign n1900 = ( ~n1026 & n1034 ) | ( ~n1026 & n1899 ) | ( n1034 & n1899 ) ;
  assign n1901 = ( n1060 & ~n1650 ) | ( n1060 & n1900 ) | ( ~n1650 & n1900 ) ;
  assign n1902 = ~n1049 & n1901 ;
  assign n1903 = n1046 | n1902 ;
  assign n1904 = ~n1053 & n1903 ;
  assign n1905 = n1050 | n1053 ;
  assign n1906 = n1024 | n1026 ;
  assign n1907 = ( ~n986 & n990 ) | ( ~n986 & n1002 ) | ( n990 & n1002 ) ;
  assign n1908 = ( ~n1648 & n1906 ) | ( ~n1648 & n1907 ) | ( n1906 & n1907 ) ;
  assign n1909 = ( ~n1063 & n1905 ) | ( ~n1063 & n1908 ) | ( n1905 & n1908 ) ;
  assign n1910 = ( n1898 & ~n1904 ) | ( n1898 & n1909 ) | ( ~n1904 & n1909 ) ;
  assign n1911 = n1070 | n1570 ;
  assign n1912 = n1658 & ~n1911 ;
  assign n1913 = ( n1661 & ~n1911 ) | ( n1661 & n1912 ) | ( ~n1911 & n1912 ) ;
  assign n1914 = n1077 | n1913 ;
  assign n1915 = ~n1077 & n1911 ;
  assign n1916 = ( n1057 & ~n1658 ) | ( n1057 & n1664 ) | ( ~n1658 & n1664 ) ;
  assign n1917 = ( ~n1077 & n1915 ) | ( ~n1077 & n1916 ) | ( n1915 & n1916 ) ;
  assign n1918 = ( n1910 & n1914 ) | ( n1910 & ~n1917 ) | ( n1914 & ~n1917 ) ;
  assign n1919 = n1842 & n1918 ;
  assign n1920 = x136 & ~n271 ;
  assign n1921 = n1123 | n1130 ;
  assign n1922 = x10 | n278 ;
  assign n1923 = ~n1081 & n1922 ;
  assign n1924 = ( ~n1106 & n1673 ) | ( ~n1106 & n1923 ) | ( n1673 & n1923 ) ;
  assign n1925 = ( n1103 & ~n1108 ) | ( n1103 & n1924 ) | ( ~n1108 & n1924 ) ;
  assign n1926 = ( ~n1128 & n1921 ) | ( ~n1128 & n1925 ) | ( n1921 & n1925 ) ;
  assign n1927 = ( ~n1145 & n1146 ) | ( ~n1145 & n1680 ) | ( n1146 & n1680 ) ;
  assign n1928 = n1149 | n1927 ;
  assign n1929 = ( n1159 & n1926 ) | ( n1159 & ~n1928 ) | ( n1926 & ~n1928 ) ;
  assign n1930 = ( ~n1177 & n1178 ) | ( ~n1177 & n1685 ) | ( n1178 & n1685 ) ;
  assign n1931 = n1181 | n1930 ;
  assign n1932 = ( n1153 & ~n1174 ) | ( n1153 & n1190 ) | ( ~n1174 & n1190 ) ;
  assign n1933 = ( ~n1181 & n1191 ) | ( ~n1181 & n1932 ) | ( n1191 & n1932 ) ;
  assign n1934 = ( n1929 & ~n1931 ) | ( n1929 & n1933 ) | ( ~n1931 & n1933 ) ;
  assign n1935 = ( n1168 & ~n1210 ) | ( n1168 & n1211 ) | ( ~n1210 & n1211 ) ;
  assign n1936 = ( ~n1214 & n1218 ) | ( ~n1214 & n1935 ) | ( n1218 & n1935 ) ;
  assign n1937 = n1214 | n1229 ;
  assign n1938 = ( n1185 & ~n1207 ) | ( n1185 & n1693 ) | ( ~n1207 & n1693 ) ;
  assign n1939 = ( ~n1218 & n1937 ) | ( ~n1218 & n1938 ) | ( n1937 & n1938 ) ;
  assign n1940 = ( n1934 & ~n1936 ) | ( n1934 & n1939 ) | ( ~n1936 & n1939 ) ;
  assign n1941 = ( ~n1197 & n1223 ) | ( ~n1197 & n1228 ) | ( n1223 & n1228 ) ;
  assign n1942 = n1254 | n1270 ;
  assign n1943 = ( ~n1258 & n1941 ) | ( ~n1258 & n1942 ) | ( n1941 & n1942 ) ;
  assign n1944 = ~n1261 & n1943 ;
  assign n1945 = n1258 | n1261 ;
  assign n1946 = ( n1204 & ~n1269 ) | ( n1204 & n1698 ) | ( ~n1269 & n1698 ) ;
  assign n1947 = ( ~n1271 & n1945 ) | ( ~n1271 & n1946 ) | ( n1945 & n1946 ) ;
  assign n1948 = ( n1940 & ~n1944 ) | ( n1940 & n1947 ) | ( ~n1944 & n1947 ) ;
  assign n1949 = n1306 | n1309 ;
  assign n1950 = ( ~n1236 & n1246 ) | ( ~n1236 & n1266 ) | ( n1246 & n1266 ) ;
  assign n1951 = ( ~n1321 & n1949 ) | ( ~n1321 & n1950 ) | ( n1949 & n1950 ) ;
  assign n1952 = ~n1299 & n1951 ;
  assign n1953 = ( ~n1239 & n1248 ) | ( ~n1239 & n1273 ) | ( n1248 & n1273 ) ;
  assign n1954 = n1302 | n1708 ;
  assign n1955 = ( ~n1306 & n1953 ) | ( ~n1306 & n1954 ) | ( n1953 & n1954 ) ;
  assign n1956 = ( n1299 & ~n1310 ) | ( n1299 & n1955 ) | ( ~n1310 & n1955 ) ;
  assign n1957 = ( n1948 & n1952 ) | ( n1948 & ~n1956 ) | ( n1952 & ~n1956 ) ;
  assign n1958 = n1352 | n1376 ;
  assign n1959 = n1284 | n1358 ;
  assign n1960 = ( n1294 & ~n1315 ) | ( n1294 & n1320 ) | ( ~n1315 & n1320 ) ;
  assign n1961 = ( ~n1720 & n1959 ) | ( ~n1720 & n1960 ) | ( n1959 & n1960 ) ;
  assign n1962 = ( n1363 & ~n1958 ) | ( n1363 & n1961 ) | ( ~n1958 & n1961 ) ;
  assign n1963 = ( ~n1283 & n1296 ) | ( ~n1283 & n1316 ) | ( n1296 & n1316 ) ;
  assign n1964 = ( ~n1359 & n1721 ) | ( ~n1359 & n1963 ) | ( n1721 & n1963 ) ;
  assign n1965 = ( n1352 & ~n1363 ) | ( n1352 & n1964 ) | ( ~n1363 & n1964 ) ;
  assign n1966 = ( n1957 & n1962 ) | ( n1957 & ~n1965 ) | ( n1962 & ~n1965 ) ;
  assign n1967 = n1416 | n1433 ;
  assign n1968 = ( n1347 & ~n1368 ) | ( n1347 & n1375 ) | ( ~n1368 & n1375 ) ;
  assign n1969 = ( n1337 & ~n1373 ) | ( n1337 & n1968 ) | ( ~n1373 & n1968 ) ;
  assign n1970 = n1413 | n1419 ;
  assign n1971 = ~n1416 & n1970 ;
  assign n1972 = ( n1967 & n1969 ) | ( n1967 & ~n1971 ) | ( n1969 & ~n1971 ) ;
  assign n1973 = ( ~n1335 & n1349 ) | ( ~n1335 & n1369 ) | ( n1349 & n1369 ) ;
  assign n1974 = ( ~n1727 & n1732 ) | ( ~n1727 & n1973 ) | ( n1732 & n1973 ) ;
  assign n1975 = ( n1420 & ~n1967 ) | ( n1420 & n1974 ) | ( ~n1967 & n1974 ) ;
  assign n1976 = ( n1966 & n1972 ) | ( n1966 & ~n1975 ) | ( n1972 & ~n1975 ) ;
  assign n1977 = ( ~n1393 & n1404 ) | ( ~n1393 & n1432 ) | ( n1404 & n1432 ) ;
  assign n1978 = ( ~n1430 & n1438 ) | ( ~n1430 & n1977 ) | ( n1438 & n1977 ) ;
  assign n1979 = ( n1464 & ~n1748 ) | ( n1464 & n1978 ) | ( ~n1748 & n1978 ) ;
  assign n1980 = ~n1453 & n1979 ;
  assign n1981 = n1450 | n1980 ;
  assign n1982 = ~n1457 & n1981 ;
  assign n1983 = n1454 | n1457 ;
  assign n1984 = n1428 | n1430 ;
  assign n1985 = ( ~n1390 & n1394 ) | ( ~n1390 & n1406 ) | ( n1394 & n1406 ) ;
  assign n1986 = ( ~n1746 & n1984 ) | ( ~n1746 & n1985 ) | ( n1984 & n1985 ) ;
  assign n1987 = ( ~n1467 & n1983 ) | ( ~n1467 & n1986 ) | ( n1983 & n1986 ) ;
  assign n1988 = ( n1976 & ~n1982 ) | ( n1976 & n1987 ) | ( ~n1982 & n1987 ) ;
  assign n1989 = ( ~n265 & n269 ) | ( ~n265 & n1756 ) | ( n269 & n1756 ) ;
  assign n1990 = n276 | n1989 ;
  assign n1991 = n265 & ~n276 ;
  assign n1992 = ( ~n268 & n1461 ) | ( ~n268 & n1759 ) | ( n1461 & n1759 ) ;
  assign n1993 = ( ~n276 & n1991 ) | ( ~n276 & n1992 ) | ( n1991 & n1992 ) ;
  assign n1994 = ( n1988 & n1990 ) | ( n1988 & ~n1993 ) | ( n1990 & ~n1993 ) ;
  assign n1995 = n1920 & n1994 ;
  assign n1996 = x137 & ~n676 ;
  assign n1997 = n358 | n374 ;
  assign n1998 = n322 | n347 ;
  assign n1999 = x11 | n683 ;
  assign n2000 = ~n296 & n1999 ;
  assign n2001 = ( ~n289 & n293 ) | ( ~n289 & n2000 ) | ( n293 & n2000 ) ;
  assign n2002 = ( ~n311 & n1480 ) | ( ~n311 & n2001 ) | ( n1480 & n2001 ) ;
  assign n2003 = ( ~n1484 & n1998 ) | ( ~n1484 & n2002 ) | ( n1998 & n2002 ) ;
  assign n2004 = ( ~n343 & n1491 ) | ( ~n343 & n2003 ) | ( n1491 & n2003 ) ;
  assign n2005 = ( ~n358 & n376 ) | ( ~n358 & n383 ) | ( n376 & n383 ) ;
  assign n2006 = ( ~n1997 & n2004 ) | ( ~n1997 & n2005 ) | ( n2004 & n2005 ) ;
  assign n2007 = ( ~n394 & n410 ) | ( ~n394 & n414 ) | ( n410 & n414 ) ;
  assign n2008 = n394 | n421 ;
  assign n2009 = ( ~n408 & n420 ) | ( ~n408 & n1496 ) | ( n420 & n1496 ) ;
  assign n2010 = ( ~n414 & n2008 ) | ( ~n414 & n2009 ) | ( n2008 & n2009 ) ;
  assign n2011 = ( n2006 & ~n2007 ) | ( n2006 & n2010 ) | ( ~n2007 & n2010 ) ;
  assign n2012 = ( n419 & ~n448 ) | ( n419 & n461 ) | ( ~n448 & n461 ) ;
  assign n2013 = n442 | n462 ;
  assign n2014 = ( ~n453 & n2012 ) | ( ~n453 & n2013 ) | ( n2012 & n2013 ) ;
  assign n2015 = ~n436 & n2014 ;
  assign n2016 = n436 | n453 ;
  assign n2017 = ( ~n445 & n449 ) | ( ~n445 & n1501 ) | ( n449 & n1501 ) ;
  assign n2018 = ( ~n464 & n2016 ) | ( ~n464 & n2017 ) | ( n2016 & n2017 ) ;
  assign n2019 = ( n2011 & ~n2015 ) | ( n2011 & n2018 ) | ( ~n2015 & n2018 ) ;
  assign n2020 = n484 | n501 ;
  assign n2021 = ( n457 & ~n493 ) | ( n457 & n497 ) | ( ~n493 & n497 ) ;
  assign n2022 = ( ~n513 & n2020 ) | ( ~n513 & n2021 ) | ( n2020 & n2021 ) ;
  assign n2023 = ~n481 & n2022 ;
  assign n2024 = ( n439 & ~n496 ) | ( n439 & n1511 ) | ( ~n496 & n1511 ) ;
  assign n2025 = n490 | n512 ;
  assign n2026 = ( ~n501 & n2024 ) | ( ~n501 & n2025 ) | ( n2024 & n2025 ) ;
  assign n2027 = ( n481 & ~n485 ) | ( n481 & n2026 ) | ( ~n485 & n2026 ) ;
  assign n2028 = ( n2019 & n2023 ) | ( n2019 & ~n2027 ) | ( n2023 & ~n2027 ) ;
  assign n2029 = ( n507 & ~n549 ) | ( n507 & n1523 ) | ( ~n549 & n1523 ) ;
  assign n2030 = ( ~n554 & n1802 ) | ( ~n554 & n2029 ) | ( n1802 & n2029 ) ;
  assign n2031 = ( n534 & ~n538 ) | ( n534 & n2030 ) | ( ~n538 & n2030 ) ;
  assign n2032 = n534 | n568 ;
  assign n2033 = n550 | n553 ;
  assign n2034 = ( ~n471 & n475 ) | ( ~n471 & n511 ) | ( n475 & n511 ) ;
  assign n2035 = ( ~n567 & n2033 ) | ( ~n567 & n2034 ) | ( n2033 & n2034 ) ;
  assign n2036 = ( n538 & ~n2032 ) | ( n538 & n2035 ) | ( ~n2032 & n2035 ) ;
  assign n2037 = ( n2028 & ~n2031 ) | ( n2028 & n2036 ) | ( ~n2031 & n2036 ) ;
  assign n2038 = n594 | n625 ;
  assign n2039 = ( ~n523 & n527 ) | ( ~n523 & n566 ) | ( n527 & n566 ) ;
  assign n2040 = ( ~n604 & n1531 ) | ( ~n604 & n2039 ) | ( n1531 & n2039 ) ;
  assign n2041 = n591 | n611 ;
  assign n2042 = ~n594 & n2041 ;
  assign n2043 = ( n2038 & n2040 ) | ( n2038 & ~n2042 ) | ( n2040 & ~n2042 ) ;
  assign n2044 = ( ~n520 & n560 ) | ( ~n520 & n564 ) | ( n560 & n564 ) ;
  assign n2045 = ( ~n624 & n1814 ) | ( ~n624 & n2044 ) | ( n1814 & n2044 ) ;
  assign n2046 = ( n595 & ~n2038 ) | ( n595 & n2045 ) | ( ~n2038 & n2045 ) ;
  assign n2047 = ( n2037 & n2043 ) | ( n2037 & ~n2046 ) | ( n2043 & ~n2046 ) ;
  assign n2048 = ( ~n578 & n623 ) | ( ~n578 & n628 ) | ( n623 & n628 ) ;
  assign n2049 = ( n1550 & ~n1551 ) | ( n1550 & n2048 ) | ( ~n1551 & n2048 ) ;
  assign n2050 = ( n657 & ~n1827 ) | ( n657 & n2049 ) | ( ~n1827 & n2049 ) ;
  assign n2051 = n638 | n2050 ;
  assign n2052 = ~n635 & n2051 ;
  assign n2053 = n635 | n649 ;
  assign n2054 = n644 | n1551 ;
  assign n2055 = ( ~n575 & n585 ) | ( ~n575 & n621 ) | ( n585 & n621 ) ;
  assign n2056 = ( ~n656 & n2054 ) | ( ~n656 & n2055 ) | ( n2054 & n2055 ) ;
  assign n2057 = ( ~n1566 & n2053 ) | ( ~n1566 & n2056 ) | ( n2053 & n2056 ) ;
  assign n2058 = ( n2047 & ~n2052 ) | ( n2047 & n2057 ) | ( ~n2052 & n2057 ) ;
  assign n2059 = ( ~n670 & n674 ) | ( ~n670 & n1834 ) | ( n674 & n1834 ) ;
  assign n2060 = n681 | n2059 ;
  assign n2061 = n670 & ~n681 ;
  assign n2062 = ( ~n673 & n1565 ) | ( ~n673 & n1837 ) | ( n1565 & n1837 ) ;
  assign n2063 = ( ~n681 & n2061 ) | ( ~n681 & n2062 ) | ( n2061 & n2062 ) ;
  assign n2064 = ( n2058 & n2060 ) | ( n2058 & ~n2063 ) | ( n2060 & ~n2063 ) ;
  assign n2065 = n1996 & n2064 ;
  assign n2066 = x138 & ~n1080 ;
  assign n2067 = n763 | n779 ;
  assign n2068 = n727 | n752 ;
  assign n2069 = x12 | n1087 ;
  assign n2070 = ~n701 & n2069 ;
  assign n2071 = ( ~n694 & n698 ) | ( ~n694 & n2070 ) | ( n698 & n2070 ) ;
  assign n2072 = ( ~n716 & n1579 ) | ( ~n716 & n2071 ) | ( n1579 & n2071 ) ;
  assign n2073 = ( ~n1583 & n2068 ) | ( ~n1583 & n2072 ) | ( n2068 & n2072 ) ;
  assign n2074 = ( ~n748 & n1590 ) | ( ~n748 & n2073 ) | ( n1590 & n2073 ) ;
  assign n2075 = ( ~n763 & n781 ) | ( ~n763 & n788 ) | ( n781 & n788 ) ;
  assign n2076 = ( ~n2067 & n2074 ) | ( ~n2067 & n2075 ) | ( n2074 & n2075 ) ;
  assign n2077 = ( ~n799 & n815 ) | ( ~n799 & n819 ) | ( n815 & n819 ) ;
  assign n2078 = n799 | n826 ;
  assign n2079 = ( ~n813 & n825 ) | ( ~n813 & n1595 ) | ( n825 & n1595 ) ;
  assign n2080 = ( ~n819 & n2078 ) | ( ~n819 & n2079 ) | ( n2078 & n2079 ) ;
  assign n2081 = ( n2076 & ~n2077 ) | ( n2076 & n2080 ) | ( ~n2077 & n2080 ) ;
  assign n2082 = ( n824 & ~n853 ) | ( n824 & n866 ) | ( ~n853 & n866 ) ;
  assign n2083 = n847 | n867 ;
  assign n2084 = ( ~n858 & n2082 ) | ( ~n858 & n2083 ) | ( n2082 & n2083 ) ;
  assign n2085 = ~n841 & n2084 ;
  assign n2086 = n841 | n858 ;
  assign n2087 = ( ~n850 & n854 ) | ( ~n850 & n1600 ) | ( n854 & n1600 ) ;
  assign n2088 = ( ~n869 & n2086 ) | ( ~n869 & n2087 ) | ( n2086 & n2087 ) ;
  assign n2089 = ( n2081 & ~n2085 ) | ( n2081 & n2088 ) | ( ~n2085 & n2088 ) ;
  assign n2090 = n889 | n906 ;
  assign n2091 = ( n862 & ~n898 ) | ( n862 & n902 ) | ( ~n898 & n902 ) ;
  assign n2092 = ( ~n918 & n2090 ) | ( ~n918 & n2091 ) | ( n2090 & n2091 ) ;
  assign n2093 = ~n886 & n2092 ;
  assign n2094 = ( n844 & ~n901 ) | ( n844 & n1610 ) | ( ~n901 & n1610 ) ;
  assign n2095 = n895 | n917 ;
  assign n2096 = ( ~n906 & n2094 ) | ( ~n906 & n2095 ) | ( n2094 & n2095 ) ;
  assign n2097 = ( n886 & ~n890 ) | ( n886 & n2096 ) | ( ~n890 & n2096 ) ;
  assign n2098 = ( n2089 & n2093 ) | ( n2089 & ~n2097 ) | ( n2093 & ~n2097 ) ;
  assign n2099 = ( n912 & ~n954 ) | ( n912 & n1622 ) | ( ~n954 & n1622 ) ;
  assign n2100 = ( ~n959 & n1880 ) | ( ~n959 & n2099 ) | ( n1880 & n2099 ) ;
  assign n2101 = ( n939 & ~n943 ) | ( n939 & n2100 ) | ( ~n943 & n2100 ) ;
  assign n2102 = n939 | n973 ;
  assign n2103 = n955 | n958 ;
  assign n2104 = ( ~n876 & n880 ) | ( ~n876 & n916 ) | ( n880 & n916 ) ;
  assign n2105 = ( ~n972 & n2103 ) | ( ~n972 & n2104 ) | ( n2103 & n2104 ) ;
  assign n2106 = ( n943 & ~n2102 ) | ( n943 & n2105 ) | ( ~n2102 & n2105 ) ;
  assign n2107 = ( n2098 & ~n2101 ) | ( n2098 & n2106 ) | ( ~n2101 & n2106 ) ;
  assign n2108 = n999 | n1030 ;
  assign n2109 = ( ~n928 & n932 ) | ( ~n928 & n971 ) | ( n932 & n971 ) ;
  assign n2110 = ( ~n1009 & n1630 ) | ( ~n1009 & n2109 ) | ( n1630 & n2109 ) ;
  assign n2111 = n996 | n1016 ;
  assign n2112 = ~n999 & n2111 ;
  assign n2113 = ( n2108 & n2110 ) | ( n2108 & ~n2112 ) | ( n2110 & ~n2112 ) ;
  assign n2114 = ( ~n925 & n965 ) | ( ~n925 & n969 ) | ( n965 & n969 ) ;
  assign n2115 = ( ~n1029 & n1892 ) | ( ~n1029 & n2114 ) | ( n1892 & n2114 ) ;
  assign n2116 = ( n1000 & ~n2108 ) | ( n1000 & n2115 ) | ( ~n2108 & n2115 ) ;
  assign n2117 = ( n2107 & n2113 ) | ( n2107 & ~n2116 ) | ( n2113 & ~n2116 ) ;
  assign n2118 = ( ~n983 & n1028 ) | ( ~n983 & n1033 ) | ( n1028 & n1033 ) ;
  assign n2119 = ( n1649 & ~n1650 ) | ( n1649 & n2118 ) | ( ~n1650 & n2118 ) ;
  assign n2120 = ( n1062 & ~n1905 ) | ( n1062 & n2119 ) | ( ~n1905 & n2119 ) ;
  assign n2121 = n1043 | n2120 ;
  assign n2122 = ~n1040 & n2121 ;
  assign n2123 = n1040 | n1054 ;
  assign n2124 = n1049 | n1650 ;
  assign n2125 = ( ~n980 & n990 ) | ( ~n980 & n1026 ) | ( n990 & n1026 ) ;
  assign n2126 = ( ~n1061 & n2124 ) | ( ~n1061 & n2125 ) | ( n2124 & n2125 ) ;
  assign n2127 = ( ~n1665 & n2123 ) | ( ~n1665 & n2126 ) | ( n2123 & n2126 ) ;
  assign n2128 = ( n2117 & ~n2122 ) | ( n2117 & n2127 ) | ( ~n2122 & n2127 ) ;
  assign n2129 = ( ~n1074 & n1078 ) | ( ~n1074 & n1912 ) | ( n1078 & n1912 ) ;
  assign n2130 = n1085 | n2129 ;
  assign n2131 = n1074 & ~n1085 ;
  assign n2132 = ( ~n1077 & n1664 ) | ( ~n1077 & n1915 ) | ( n1664 & n1915 ) ;
  assign n2133 = ( ~n1085 & n2131 ) | ( ~n1085 & n2132 ) | ( n2131 & n2132 ) ;
  assign n2134 = ( n2128 & n2130 ) | ( n2128 & ~n2133 ) | ( n2130 & ~n2133 ) ;
  assign n2135 = n2066 & n2134 ;
  assign n2136 = x139 & ~n295 ;
  assign n2137 = n1167 | n1183 ;
  assign n2138 = n1131 | n1156 ;
  assign n2139 = x13 | n290 ;
  assign n2140 = ~n1105 & n2139 ;
  assign n2141 = ( ~n1098 & n1102 ) | ( ~n1098 & n2140 ) | ( n1102 & n2140 ) ;
  assign n2142 = ( ~n1120 & n1677 ) | ( ~n1120 & n2141 ) | ( n1677 & n2141 ) ;
  assign n2143 = ( ~n1681 & n2138 ) | ( ~n1681 & n2142 ) | ( n2138 & n2142 ) ;
  assign n2144 = ( ~n1152 & n1688 ) | ( ~n1152 & n2143 ) | ( n1688 & n2143 ) ;
  assign n2145 = ( ~n1167 & n1185 ) | ( ~n1167 & n1192 ) | ( n1185 & n1192 ) ;
  assign n2146 = ( ~n2137 & n2144 ) | ( ~n2137 & n2145 ) | ( n2144 & n2145 ) ;
  assign n2147 = ( ~n1203 & n1219 ) | ( ~n1203 & n1223 ) | ( n1219 & n1223 ) ;
  assign n2148 = n1203 | n1230 ;
  assign n2149 = ( ~n1217 & n1229 ) | ( ~n1217 & n1693 ) | ( n1229 & n1693 ) ;
  assign n2150 = ( ~n1223 & n2148 ) | ( ~n1223 & n2149 ) | ( n2148 & n2149 ) ;
  assign n2151 = ( n2146 & ~n2147 ) | ( n2146 & n2150 ) | ( ~n2147 & n2150 ) ;
  assign n2152 = ( n1228 & ~n1257 ) | ( n1228 & n1270 ) | ( ~n1257 & n1270 ) ;
  assign n2153 = n1251 | n1271 ;
  assign n2154 = ( ~n1262 & n2152 ) | ( ~n1262 & n2153 ) | ( n2152 & n2153 ) ;
  assign n2155 = ~n1245 & n2154 ;
  assign n2156 = n1245 | n1262 ;
  assign n2157 = ( ~n1254 & n1258 ) | ( ~n1254 & n1698 ) | ( n1258 & n1698 ) ;
  assign n2158 = ( ~n1273 & n2156 ) | ( ~n1273 & n2157 ) | ( n2156 & n2157 ) ;
  assign n2159 = ( n2151 & ~n2155 ) | ( n2151 & n2158 ) | ( ~n2155 & n2158 ) ;
  assign n2160 = n1293 | n1310 ;
  assign n2161 = ( n1266 & ~n1302 ) | ( n1266 & n1306 ) | ( ~n1302 & n1306 ) ;
  assign n2162 = ( ~n1322 & n2160 ) | ( ~n1322 & n2161 ) | ( n2160 & n2161 ) ;
  assign n2163 = ~n1290 & n2162 ;
  assign n2164 = ( n1248 & ~n1305 ) | ( n1248 & n1708 ) | ( ~n1305 & n1708 ) ;
  assign n2165 = n1299 | n1321 ;
  assign n2166 = ( ~n1310 & n2164 ) | ( ~n1310 & n2165 ) | ( n2164 & n2165 ) ;
  assign n2167 = ( n1290 & ~n1294 ) | ( n1290 & n2166 ) | ( ~n1294 & n2166 ) ;
  assign n2168 = ( n2159 & n2163 ) | ( n2159 & ~n2167 ) | ( n2163 & ~n2167 ) ;
  assign n2169 = ( n1316 & ~n1358 ) | ( n1316 & n1720 ) | ( ~n1358 & n1720 ) ;
  assign n2170 = ( ~n1363 & n1958 ) | ( ~n1363 & n2169 ) | ( n1958 & n2169 ) ;
  assign n2171 = ( n1343 & ~n1347 ) | ( n1343 & n2170 ) | ( ~n1347 & n2170 ) ;
  assign n2172 = n1343 | n1377 ;
  assign n2173 = n1359 | n1362 ;
  assign n2174 = ( ~n1280 & n1284 ) | ( ~n1280 & n1320 ) | ( n1284 & n1320 ) ;
  assign n2175 = ( ~n1376 & n2173 ) | ( ~n1376 & n2174 ) | ( n2173 & n2174 ) ;
  assign n2176 = ( n1347 & ~n2172 ) | ( n1347 & n2175 ) | ( ~n2172 & n2175 ) ;
  assign n2177 = ( n2168 & ~n2171 ) | ( n2168 & n2176 ) | ( ~n2171 & n2176 ) ;
  assign n2178 = n1403 | n1434 ;
  assign n2179 = ( ~n1332 & n1336 ) | ( ~n1332 & n1375 ) | ( n1336 & n1375 ) ;
  assign n2180 = ( ~n1413 & n1728 ) | ( ~n1413 & n2179 ) | ( n1728 & n2179 ) ;
  assign n2181 = n1400 | n1420 ;
  assign n2182 = ~n1403 & n2181 ;
  assign n2183 = ( n2178 & n2180 ) | ( n2178 & ~n2182 ) | ( n2180 & ~n2182 ) ;
  assign n2184 = ( ~n1329 & n1369 ) | ( ~n1329 & n1373 ) | ( n1369 & n1373 ) ;
  assign n2185 = ( ~n1433 & n1970 ) | ( ~n1433 & n2184 ) | ( n1970 & n2184 ) ;
  assign n2186 = ( n1404 & ~n2178 ) | ( n1404 & n2185 ) | ( ~n2178 & n2185 ) ;
  assign n2187 = ( n2177 & n2183 ) | ( n2177 & ~n2186 ) | ( n2183 & ~n2186 ) ;
  assign n2188 = ( ~n1387 & n1432 ) | ( ~n1387 & n1437 ) | ( n1432 & n1437 ) ;
  assign n2189 = ( n1747 & ~n1748 ) | ( n1747 & n2188 ) | ( ~n1748 & n2188 ) ;
  assign n2190 = ( n1466 & ~n1983 ) | ( n1466 & n2189 ) | ( ~n1983 & n2189 ) ;
  assign n2191 = n1447 | n2190 ;
  assign n2192 = ~n1444 & n2191 ;
  assign n2193 = n1444 | n1458 ;
  assign n2194 = n1453 | n1748 ;
  assign n2195 = ( ~n1384 & n1394 ) | ( ~n1384 & n1430 ) | ( n1394 & n1430 ) ;
  assign n2196 = ( ~n1465 & n2194 ) | ( ~n1465 & n2195 ) | ( n2194 & n2195 ) ;
  assign n2197 = ( ~n1760 & n2193 ) | ( ~n1760 & n2196 ) | ( n2193 & n2196 ) ;
  assign n2198 = ( n2187 & ~n2192 ) | ( n2187 & n2197 ) | ( ~n2192 & n2197 ) ;
  assign n2199 = ( n269 & ~n273 ) | ( n269 & n277 ) | ( ~n273 & n277 ) ;
  assign n2200 = n280 | n2199 ;
  assign n2201 = ( ~n276 & n1759 ) | ( ~n276 & n1991 ) | ( n1759 & n1991 ) ;
  assign n2202 = ( ~n280 & n282 ) | ( ~n280 & n2201 ) | ( n282 & n2201 ) ;
  assign n2203 = ( n2198 & n2200 ) | ( n2198 & ~n2202 ) | ( n2200 & ~n2202 ) ;
  assign n2204 = n2136 & n2203 ;
  assign n2205 = x140 & ~n700 ;
  assign n2206 = n503 & ~n506 ;
  assign n2207 = ~n430 & n466 ;
  assign n2208 = n398 | n1494 ;
  assign n2209 = n336 | n348 ;
  assign n2210 = x14 | n695 ;
  assign n2211 = ~n288 & n2210 ;
  assign n2212 = ( ~n307 & n1479 ) | ( ~n307 & n2211 ) | ( n1479 & n2211 ) ;
  assign n2213 = ( ~n318 & n1765 ) | ( ~n318 & n2212 ) | ( n1765 & n2212 ) ;
  assign n2214 = ( ~n1771 & n2209 ) | ( ~n1771 & n2213 ) | ( n2209 & n2213 ) ;
  assign n2215 = ( ~n1490 & n1776 ) | ( ~n1490 & n2214 ) | ( n1776 & n2214 ) ;
  assign n2216 = ( ~n398 & n1496 ) | ( ~n398 & n1498 ) | ( n1496 & n1498 ) ;
  assign n2217 = ( ~n2208 & n2215 ) | ( ~n2208 & n2216 ) | ( n2215 & n2216 ) ;
  assign n2218 = ( ~n388 & n419 ) | ( ~n388 & n1502 ) | ( n419 & n1502 ) ;
  assign n2219 = ( n423 & n2217 ) | ( n423 & ~n2218 ) | ( n2217 & ~n2218 ) ;
  assign n2220 = ( n455 & ~n2207 ) | ( n455 & n2219 ) | ( ~n2207 & n2219 ) ;
  assign n2221 = n481 | n513 ;
  assign n2222 = ( ~n500 & n512 ) | ( ~n500 & n1511 ) | ( n512 & n1511 ) ;
  assign n2223 = ( ~n485 & n2221 ) | ( ~n485 & n2222 ) | ( n2221 & n2222 ) ;
  assign n2224 = ( n506 & ~n511 ) | ( n506 & n2223 ) | ( ~n511 & n2223 ) ;
  assign n2225 = ( n2206 & n2220 ) | ( n2206 & ~n2224 ) | ( n2220 & ~n2224 ) ;
  assign n2226 = ( ~n553 & n567 ) | ( ~n553 & n1523 ) | ( n567 & n1523 ) ;
  assign n2227 = ( ~n538 & n2032 ) | ( ~n538 & n2226 ) | ( n2032 & n2226 ) ;
  assign n2228 = ( n559 & ~n566 ) | ( n559 & n2227 ) | ( ~n566 & n2227 ) ;
  assign n2229 = n537 | n554 ;
  assign n2230 = ( n475 & ~n546 ) | ( n475 & n550 ) | ( ~n546 & n550 ) ;
  assign n2231 = ( ~n568 & n2229 ) | ( ~n568 & n2230 ) | ( n2229 & n2230 ) ;
  assign n2232 = ( ~n565 & n566 ) | ( ~n565 & n2231 ) | ( n566 & n2231 ) ;
  assign n2233 = ( n2225 & ~n2228 ) | ( n2225 & n2232 ) | ( ~n2228 & n2232 ) ;
  assign n2234 = ( n527 & ~n600 ) | ( n527 & n1530 ) | ( ~n600 & n1530 ) ;
  assign n2235 = ( ~n611 & n1811 ) | ( ~n611 & n2234 ) | ( n1811 & n2234 ) ;
  assign n2236 = ~n584 & n596 ;
  assign n2237 = ( n622 & n2235 ) | ( n622 & ~n2236 ) | ( n2235 & ~n2236 ) ;
  assign n2238 = ( n564 & ~n603 ) | ( n564 & n604 ) | ( ~n603 & n604 ) ;
  assign n2239 = ( ~n625 & n2041 ) | ( ~n625 & n2238 ) | ( n2041 & n2238 ) ;
  assign n2240 = ( ~n622 & n623 ) | ( ~n622 & n2239 ) | ( n623 & n2239 ) ;
  assign n2241 = ( n2233 & n2237 ) | ( n2233 & ~n2240 ) | ( n2237 & ~n2240 ) ;
  assign n2242 = n641 | n656 ;
  assign n2243 = ( ~n619 & n628 ) | ( ~n619 & n1549 ) | ( n628 & n1549 ) ;
  assign n2244 = ( ~n645 & n2242 ) | ( ~n645 & n2243 ) | ( n2242 & n2243 ) ;
  assign n2245 = ( n652 & ~n2053 ) | ( n652 & n2244 ) | ( ~n2053 & n2244 ) ;
  assign n2246 = n1561 | n2245 ;
  assign n2247 = ~n1559 & n2246 ;
  assign n2248 = n1559 | n1562 ;
  assign n2249 = ( n621 & ~n655 ) | ( n621 & n1551 ) | ( ~n655 & n1551 ) ;
  assign n2250 = ( ~n657 & n1827 ) | ( ~n657 & n2249 ) | ( n1827 & n2249 ) ;
  assign n2251 = n652 | n1561 ;
  assign n2252 = ~n1559 & n2251 ;
  assign n2253 = ( n2248 & n2250 ) | ( n2248 & ~n2252 ) | ( n2250 & ~n2252 ) ;
  assign n2254 = ( n2241 & ~n2247 ) | ( n2241 & n2253 ) | ( ~n2247 & n2253 ) ;
  assign n2255 = ( n674 & ~n678 ) | ( n674 & n682 ) | ( ~n678 & n682 ) ;
  assign n2256 = n685 | n2255 ;
  assign n2257 = ( ~n681 & n1837 ) | ( ~n681 & n2061 ) | ( n1837 & n2061 ) ;
  assign n2258 = ( ~n685 & n687 ) | ( ~n685 & n2257 ) | ( n687 & n2257 ) ;
  assign n2259 = ( n2254 & n2256 ) | ( n2254 & ~n2258 ) | ( n2256 & ~n2258 ) ;
  assign n2260 = n2205 & n2259 ;
  assign n2261 = x141 & ~n1104 ;
  assign n2262 = n908 & ~n911 ;
  assign n2263 = ~n835 & n871 ;
  assign n2264 = n803 | n1593 ;
  assign n2265 = n741 | n753 ;
  assign n2266 = x15 | n1099 ;
  assign n2267 = ~n693 & n2266 ;
  assign n2268 = ( ~n712 & n1578 ) | ( ~n712 & n2267 ) | ( n1578 & n2267 ) ;
  assign n2269 = ( ~n723 & n1843 ) | ( ~n723 & n2268 ) | ( n1843 & n2268 ) ;
  assign n2270 = ( ~n1849 & n2265 ) | ( ~n1849 & n2269 ) | ( n2265 & n2269 ) ;
  assign n2271 = ( ~n1589 & n1854 ) | ( ~n1589 & n2270 ) | ( n1854 & n2270 ) ;
  assign n2272 = ( ~n803 & n1595 ) | ( ~n803 & n1597 ) | ( n1595 & n1597 ) ;
  assign n2273 = ( ~n2264 & n2271 ) | ( ~n2264 & n2272 ) | ( n2271 & n2272 ) ;
  assign n2274 = ( ~n793 & n824 ) | ( ~n793 & n1601 ) | ( n824 & n1601 ) ;
  assign n2275 = ( n828 & n2273 ) | ( n828 & ~n2274 ) | ( n2273 & ~n2274 ) ;
  assign n2276 = ( n860 & ~n2263 ) | ( n860 & n2275 ) | ( ~n2263 & n2275 ) ;
  assign n2277 = n886 | n918 ;
  assign n2278 = ( ~n905 & n917 ) | ( ~n905 & n1610 ) | ( n917 & n1610 ) ;
  assign n2279 = ( ~n890 & n2277 ) | ( ~n890 & n2278 ) | ( n2277 & n2278 ) ;
  assign n2280 = ( n911 & ~n916 ) | ( n911 & n2279 ) | ( ~n916 & n2279 ) ;
  assign n2281 = ( n2262 & n2276 ) | ( n2262 & ~n2280 ) | ( n2276 & ~n2280 ) ;
  assign n2282 = ( ~n958 & n972 ) | ( ~n958 & n1622 ) | ( n972 & n1622 ) ;
  assign n2283 = ( ~n943 & n2102 ) | ( ~n943 & n2282 ) | ( n2102 & n2282 ) ;
  assign n2284 = ( n964 & ~n971 ) | ( n964 & n2283 ) | ( ~n971 & n2283 ) ;
  assign n2285 = n942 | n959 ;
  assign n2286 = ( n880 & ~n951 ) | ( n880 & n955 ) | ( ~n951 & n955 ) ;
  assign n2287 = ( ~n973 & n2285 ) | ( ~n973 & n2286 ) | ( n2285 & n2286 ) ;
  assign n2288 = ( ~n970 & n971 ) | ( ~n970 & n2287 ) | ( n971 & n2287 ) ;
  assign n2289 = ( n2281 & ~n2284 ) | ( n2281 & n2288 ) | ( ~n2284 & n2288 ) ;
  assign n2290 = ( n932 & ~n1005 ) | ( n932 & n1629 ) | ( ~n1005 & n1629 ) ;
  assign n2291 = ( ~n1016 & n1889 ) | ( ~n1016 & n2290 ) | ( n1889 & n2290 ) ;
  assign n2292 = ~n989 & n1001 ;
  assign n2293 = ( n1027 & n2291 ) | ( n1027 & ~n2292 ) | ( n2291 & ~n2292 ) ;
  assign n2294 = ( n969 & ~n1008 ) | ( n969 & n1009 ) | ( ~n1008 & n1009 ) ;
  assign n2295 = ( ~n1030 & n2111 ) | ( ~n1030 & n2294 ) | ( n2111 & n2294 ) ;
  assign n2296 = ( ~n1027 & n1028 ) | ( ~n1027 & n2295 ) | ( n1028 & n2295 ) ;
  assign n2297 = ( n2289 & n2293 ) | ( n2289 & ~n2296 ) | ( n2293 & ~n2296 ) ;
  assign n2298 = n1046 | n1061 ;
  assign n2299 = ( ~n1024 & n1033 ) | ( ~n1024 & n1648 ) | ( n1033 & n1648 ) ;
  assign n2300 = ( ~n1050 & n2298 ) | ( ~n1050 & n2299 ) | ( n2298 & n2299 ) ;
  assign n2301 = ( n1057 & ~n2123 ) | ( n1057 & n2300 ) | ( ~n2123 & n2300 ) ;
  assign n2302 = n1660 | n2301 ;
  assign n2303 = ~n1658 & n2302 ;
  assign n2304 = n1658 | n1661 ;
  assign n2305 = ( n1026 & ~n1060 ) | ( n1026 & n1650 ) | ( ~n1060 & n1650 ) ;
  assign n2306 = ( ~n1062 & n1905 ) | ( ~n1062 & n2305 ) | ( n1905 & n2305 ) ;
  assign n2307 = n1057 | n1660 ;
  assign n2308 = ~n1658 & n2307 ;
  assign n2309 = ( n2304 & n2306 ) | ( n2304 & ~n2308 ) | ( n2306 & ~n2308 ) ;
  assign n2310 = ( n2297 & ~n2303 ) | ( n2297 & n2309 ) | ( ~n2303 & n2309 ) ;
  assign n2311 = ( n1078 & ~n1082 ) | ( n1078 & n1086 ) | ( ~n1082 & n1086 ) ;
  assign n2312 = n1089 | n2311 ;
  assign n2313 = ( ~n1085 & n1915 ) | ( ~n1085 & n2131 ) | ( n1915 & n2131 ) ;
  assign n2314 = ( ~n1089 & n1091 ) | ( ~n1089 & n2313 ) | ( n1091 & n2313 ) ;
  assign n2315 = ( n2310 & n2312 ) | ( n2310 & ~n2314 ) | ( n2312 & ~n2314 ) ;
  assign n2316 = n2261 & n2315 ;
  assign n2317 = x142 & ~n287 ;
  assign n2318 = n1312 & ~n1315 ;
  assign n2319 = ~n1239 & n1275 ;
  assign n2320 = n1207 | n1691 ;
  assign n2321 = n1145 | n1157 ;
  assign n2322 = x16 | n284 ;
  assign n2323 = ~n1097 & n2322 ;
  assign n2324 = ( ~n1116 & n1676 ) | ( ~n1116 & n2323 ) | ( n1676 & n2323 ) ;
  assign n2325 = ( ~n1127 & n1921 ) | ( ~n1127 & n2324 ) | ( n1921 & n2324 ) ;
  assign n2326 = ( ~n1927 & n2321 ) | ( ~n1927 & n2325 ) | ( n2321 & n2325 ) ;
  assign n2327 = ( ~n1687 & n1932 ) | ( ~n1687 & n2326 ) | ( n1932 & n2326 ) ;
  assign n2328 = ( ~n1207 & n1693 ) | ( ~n1207 & n1695 ) | ( n1693 & n1695 ) ;
  assign n2329 = ( ~n2320 & n2327 ) | ( ~n2320 & n2328 ) | ( n2327 & n2328 ) ;
  assign n2330 = ( ~n1197 & n1228 ) | ( ~n1197 & n1699 ) | ( n1228 & n1699 ) ;
  assign n2331 = ( n1232 & n2329 ) | ( n1232 & ~n2330 ) | ( n2329 & ~n2330 ) ;
  assign n2332 = ( n1264 & ~n2319 ) | ( n1264 & n2331 ) | ( ~n2319 & n2331 ) ;
  assign n2333 = n1290 | n1322 ;
  assign n2334 = ( ~n1309 & n1321 ) | ( ~n1309 & n1708 ) | ( n1321 & n1708 ) ;
  assign n2335 = ( ~n1294 & n2333 ) | ( ~n1294 & n2334 ) | ( n2333 & n2334 ) ;
  assign n2336 = ( n1315 & ~n1320 ) | ( n1315 & n2335 ) | ( ~n1320 & n2335 ) ;
  assign n2337 = ( n2318 & n2332 ) | ( n2318 & ~n2336 ) | ( n2332 & ~n2336 ) ;
  assign n2338 = ( ~n1362 & n1376 ) | ( ~n1362 & n1720 ) | ( n1376 & n1720 ) ;
  assign n2339 = ( ~n1347 & n2172 ) | ( ~n1347 & n2338 ) | ( n2172 & n2338 ) ;
  assign n2340 = ( n1368 & ~n1375 ) | ( n1368 & n2339 ) | ( ~n1375 & n2339 ) ;
  assign n2341 = n1346 | n1363 ;
  assign n2342 = ( n1284 & ~n1355 ) | ( n1284 & n1359 ) | ( ~n1355 & n1359 ) ;
  assign n2343 = ( ~n1377 & n2341 ) | ( ~n1377 & n2342 ) | ( n2341 & n2342 ) ;
  assign n2344 = ( ~n1374 & n1375 ) | ( ~n1374 & n2343 ) | ( n1375 & n2343 ) ;
  assign n2345 = ( n2337 & ~n2340 ) | ( n2337 & n2344 ) | ( ~n2340 & n2344 ) ;
  assign n2346 = ( n1336 & ~n1409 ) | ( n1336 & n1727 ) | ( ~n1409 & n1727 ) ;
  assign n2347 = ( ~n1420 & n1967 ) | ( ~n1420 & n2346 ) | ( n1967 & n2346 ) ;
  assign n2348 = ~n1393 & n1405 ;
  assign n2349 = ( n1431 & n2347 ) | ( n1431 & ~n2348 ) | ( n2347 & ~n2348 ) ;
  assign n2350 = ( n1373 & ~n1412 ) | ( n1373 & n1413 ) | ( ~n1412 & n1413 ) ;
  assign n2351 = ( ~n1434 & n2181 ) | ( ~n1434 & n2350 ) | ( n2181 & n2350 ) ;
  assign n2352 = ( ~n1431 & n1432 ) | ( ~n1431 & n2351 ) | ( n1432 & n2351 ) ;
  assign n2353 = ( n2345 & n2349 ) | ( n2345 & ~n2352 ) | ( n2349 & ~n2352 ) ;
  assign n2354 = n1450 | n1465 ;
  assign n2355 = ( ~n1428 & n1437 ) | ( ~n1428 & n1746 ) | ( n1437 & n1746 ) ;
  assign n2356 = ( ~n1454 & n2354 ) | ( ~n1454 & n2355 ) | ( n2354 & n2355 ) ;
  assign n2357 = ( n1461 & ~n2193 ) | ( n1461 & n2356 ) | ( ~n2193 & n2356 ) ;
  assign n2358 = n1755 | n2357 ;
  assign n2359 = ~n268 & n2358 ;
  assign n2360 = n268 | n1756 ;
  assign n2361 = ( n1430 & ~n1464 ) | ( n1430 & n1748 ) | ( ~n1464 & n1748 ) ;
  assign n2362 = ( ~n1466 & n1983 ) | ( ~n1466 & n2361 ) | ( n1983 & n2361 ) ;
  assign n2363 = n1461 | n1755 ;
  assign n2364 = ~n268 & n2363 ;
  assign n2365 = ( n2360 & n2362 ) | ( n2360 & ~n2364 ) | ( n2362 & ~n2364 ) ;
  assign n2366 = ( n2353 & ~n2359 ) | ( n2353 & n2365 ) | ( ~n2359 & n2365 ) ;
  assign n2367 = ( n277 & ~n297 ) | ( n277 & n1476 ) | ( ~n297 & n1476 ) ;
  assign n2368 = n292 | n2367 ;
  assign n2369 = ( ~n280 & n282 ) | ( ~n280 & n1991 ) | ( n282 & n1991 ) ;
  assign n2370 = ( ~n292 & n298 ) | ( ~n292 & n2369 ) | ( n298 & n2369 ) ;
  assign n2371 = ( n2366 & n2368 ) | ( n2366 & ~n2370 ) | ( n2368 & ~n2370 ) ;
  assign n2372 = n2317 & n2371 ;
  assign n2373 = x143 & ~n692 ;
  assign n2374 = ~n471 & n1522 ;
  assign n2375 = ~n496 & n1517 ;
  assign n2376 = n408 | n1779 ;
  assign n2377 = n330 | n349 ;
  assign n2378 = x17 | n689 ;
  assign n2379 = ~n306 & n2378 ;
  assign n2380 = ( ~n317 & n321 ) | ( ~n317 & n2379 ) | ( n321 & n2379 ) ;
  assign n2381 = ( ~n1483 & n1998 ) | ( ~n1483 & n2380 ) | ( n1998 & n2380 ) ;
  assign n2382 = ( ~n342 & n2377 ) | ( ~n342 & n2381 ) | ( n2377 & n2381 ) ;
  assign n2383 = ( n383 & ~n1775 ) | ( n383 & n2382 ) | ( ~n1775 & n2382 ) ;
  assign n2384 = ( ~n408 & n420 ) | ( ~n408 & n1782 ) | ( n420 & n1782 ) ;
  assign n2385 = ( ~n2376 & n2383 ) | ( ~n2376 & n2384 ) | ( n2383 & n2384 ) ;
  assign n2386 = ( ~n448 & n461 ) | ( ~n448 & n1785 ) | ( n461 & n1785 ) ;
  assign n2387 = ( n1508 & n2385 ) | ( n1508 & ~n2386 ) | ( n2385 & ~n2386 ) ;
  assign n2388 = ( n1513 & ~n2375 ) | ( n1513 & n2387 ) | ( ~n2375 & n2387 ) ;
  assign n2389 = ( ~n516 & n2374 ) | ( ~n516 & n2388 ) | ( n2374 & n2388 ) ;
  assign n2390 = ( n523 & ~n527 ) | ( n523 & n570 ) | ( ~n527 & n570 ) ;
  assign n2391 = ( n527 & n556 ) | ( n527 & ~n561 ) | ( n556 & ~n561 ) ;
  assign n2392 = ( n2389 & ~n2390 ) | ( n2389 & n2391 ) | ( ~n2390 & n2391 ) ;
  assign n2393 = ( ~n610 & n624 ) | ( ~n610 & n1530 ) | ( n624 & n1530 ) ;
  assign n2394 = ( ~n595 & n2038 ) | ( ~n595 & n2393 ) | ( n2038 & n2393 ) ;
  assign n2395 = ~n578 & n1542 ;
  assign n2396 = ( n1552 & n2394 ) | ( n1552 & ~n2395 ) | ( n2394 & ~n2395 ) ;
  assign n2397 = ( ~n615 & n2392 ) | ( ~n615 & n2396 ) | ( n2392 & n2396 ) ;
  assign n2398 = n638 | n657 ;
  assign n2399 = ( ~n644 & n656 ) | ( ~n644 & n1549 ) | ( n656 & n1549 ) ;
  assign n2400 = ( ~n649 & n2398 ) | ( ~n649 & n2399 ) | ( n2398 & n2399 ) ;
  assign n2401 = ( n1565 & ~n2248 ) | ( n1565 & n2400 ) | ( ~n2248 & n2400 ) ;
  assign n2402 = n1833 | n2401 ;
  assign n2403 = ~n673 & n2402 ;
  assign n2404 = n673 | n1834 ;
  assign n2405 = ( ~n641 & n645 ) | ( ~n641 & n1551 ) | ( n645 & n1551 ) ;
  assign n2406 = ( ~n652 & n2053 ) | ( ~n652 & n2405 ) | ( n2053 & n2405 ) ;
  assign n2407 = n1565 | n1833 ;
  assign n2408 = ~n673 & n2407 ;
  assign n2409 = ( n2404 & n2406 ) | ( n2404 & ~n2408 ) | ( n2406 & ~n2408 ) ;
  assign n2410 = ( n2397 & ~n2403 ) | ( n2397 & n2409 ) | ( ~n2403 & n2409 ) ;
  assign n2411 = ( n682 & ~n702 ) | ( n682 & n1575 ) | ( ~n702 & n1575 ) ;
  assign n2412 = n697 | n2411 ;
  assign n2413 = ( ~n685 & n687 ) | ( ~n685 & n2061 ) | ( n687 & n2061 ) ;
  assign n2414 = ( ~n697 & n703 ) | ( ~n697 & n2413 ) | ( n703 & n2413 ) ;
  assign n2415 = ( n2410 & n2412 ) | ( n2410 & ~n2414 ) | ( n2412 & ~n2414 ) ;
  assign n2416 = n2373 & n2415 ;
  assign n2417 = x144 & ~n1096 ;
  assign n2418 = ~n876 & n1621 ;
  assign n2419 = ~n901 & n1616 ;
  assign n2420 = n813 | n1857 ;
  assign n2421 = n735 | n754 ;
  assign n2422 = x18 | n1093 ;
  assign n2423 = ~n711 & n2422 ;
  assign n2424 = ( ~n722 & n726 ) | ( ~n722 & n2423 ) | ( n726 & n2423 ) ;
  assign n2425 = ( ~n1582 & n2068 ) | ( ~n1582 & n2424 ) | ( n2068 & n2424 ) ;
  assign n2426 = ( ~n747 & n2421 ) | ( ~n747 & n2425 ) | ( n2421 & n2425 ) ;
  assign n2427 = ( n788 & ~n1853 ) | ( n788 & n2426 ) | ( ~n1853 & n2426 ) ;
  assign n2428 = ( ~n813 & n825 ) | ( ~n813 & n1860 ) | ( n825 & n1860 ) ;
  assign n2429 = ( ~n2420 & n2427 ) | ( ~n2420 & n2428 ) | ( n2427 & n2428 ) ;
  assign n2430 = ( ~n853 & n866 ) | ( ~n853 & n1863 ) | ( n866 & n1863 ) ;
  assign n2431 = ( n1607 & n2429 ) | ( n1607 & ~n2430 ) | ( n2429 & ~n2430 ) ;
  assign n2432 = ( n1612 & ~n2419 ) | ( n1612 & n2431 ) | ( ~n2419 & n2431 ) ;
  assign n2433 = ( ~n921 & n2418 ) | ( ~n921 & n2432 ) | ( n2418 & n2432 ) ;
  assign n2434 = ( n928 & ~n932 ) | ( n928 & n975 ) | ( ~n932 & n975 ) ;
  assign n2435 = ( n932 & n961 ) | ( n932 & ~n966 ) | ( n961 & ~n966 ) ;
  assign n2436 = ( n2433 & ~n2434 ) | ( n2433 & n2435 ) | ( ~n2434 & n2435 ) ;
  assign n2437 = ( ~n1015 & n1029 ) | ( ~n1015 & n1629 ) | ( n1029 & n1629 ) ;
  assign n2438 = ( ~n1000 & n2108 ) | ( ~n1000 & n2437 ) | ( n2108 & n2437 ) ;
  assign n2439 = ~n983 & n1641 ;
  assign n2440 = ( n1651 & n2438 ) | ( n1651 & ~n2439 ) | ( n2438 & ~n2439 ) ;
  assign n2441 = ( ~n1020 & n2436 ) | ( ~n1020 & n2440 ) | ( n2436 & n2440 ) ;
  assign n2442 = n1043 | n1062 ;
  assign n2443 = ( ~n1049 & n1061 ) | ( ~n1049 & n1648 ) | ( n1061 & n1648 ) ;
  assign n2444 = ( ~n1054 & n2442 ) | ( ~n1054 & n2443 ) | ( n2442 & n2443 ) ;
  assign n2445 = ( n1664 & ~n2304 ) | ( n1664 & n2444 ) | ( ~n2304 & n2444 ) ;
  assign n2446 = n1911 | n2445 ;
  assign n2447 = ~n1077 & n2446 ;
  assign n2448 = n1077 | n1912 ;
  assign n2449 = ( ~n1046 & n1050 ) | ( ~n1046 & n1650 ) | ( n1050 & n1650 ) ;
  assign n2450 = ( ~n1057 & n2123 ) | ( ~n1057 & n2449 ) | ( n2123 & n2449 ) ;
  assign n2451 = n1664 | n1911 ;
  assign n2452 = ~n1077 & n2451 ;
  assign n2453 = ( n2448 & n2450 ) | ( n2448 & ~n2452 ) | ( n2450 & ~n2452 ) ;
  assign n2454 = ( n2441 & ~n2447 ) | ( n2441 & n2453 ) | ( ~n2447 & n2453 ) ;
  assign n2455 = ( n1086 & ~n1106 ) | ( n1086 & n1673 ) | ( ~n1106 & n1673 ) ;
  assign n2456 = n1101 | n2455 ;
  assign n2457 = ( ~n1089 & n1091 ) | ( ~n1089 & n2131 ) | ( n1091 & n2131 ) ;
  assign n2458 = ( ~n1101 & n1107 ) | ( ~n1101 & n2457 ) | ( n1107 & n2457 ) ;
  assign n2459 = ( n2454 & n2456 ) | ( n2454 & ~n2458 ) | ( n2456 & ~n2458 ) ;
  assign n2460 = n2417 & n2459 ;
  assign n2461 = x145 & ~n305 ;
  assign n2462 = ~n1280 & n1719 ;
  assign n2463 = ~n1305 & n1714 ;
  assign n2464 = n1217 | n1935 ;
  assign n2465 = n1139 | n1158 ;
  assign n2466 = x19 | n308 ;
  assign n2467 = ~n1115 & n2466 ;
  assign n2468 = ( ~n1126 & n1130 ) | ( ~n1126 & n2467 ) | ( n1130 & n2467 ) ;
  assign n2469 = ( ~n1680 & n2138 ) | ( ~n1680 & n2468 ) | ( n2138 & n2468 ) ;
  assign n2470 = ( ~n1151 & n2465 ) | ( ~n1151 & n2469 ) | ( n2465 & n2469 ) ;
  assign n2471 = ( n1192 & ~n1931 ) | ( n1192 & n2470 ) | ( ~n1931 & n2470 ) ;
  assign n2472 = ( ~n1217 & n1229 ) | ( ~n1217 & n1938 ) | ( n1229 & n1938 ) ;
  assign n2473 = ( ~n2464 & n2471 ) | ( ~n2464 & n2472 ) | ( n2471 & n2472 ) ;
  assign n2474 = ( ~n1257 & n1270 ) | ( ~n1257 & n1941 ) | ( n1270 & n1941 ) ;
  assign n2475 = ( n1705 & n2473 ) | ( n1705 & ~n2474 ) | ( n2473 & ~n2474 ) ;
  assign n2476 = ( n1710 & ~n2463 ) | ( n1710 & n2475 ) | ( ~n2463 & n2475 ) ;
  assign n2477 = ( ~n1325 & n2462 ) | ( ~n1325 & n2476 ) | ( n2462 & n2476 ) ;
  assign n2478 = ( n1332 & ~n1336 ) | ( n1332 & n1379 ) | ( ~n1336 & n1379 ) ;
  assign n2479 = ( n1336 & n1365 ) | ( n1336 & ~n1370 ) | ( n1365 & ~n1370 ) ;
  assign n2480 = ( n2477 & ~n2478 ) | ( n2477 & n2479 ) | ( ~n2478 & n2479 ) ;
  assign n2481 = ( ~n1419 & n1433 ) | ( ~n1419 & n1727 ) | ( n1433 & n1727 ) ;
  assign n2482 = ( ~n1404 & n2178 ) | ( ~n1404 & n2481 ) | ( n2178 & n2481 ) ;
  assign n2483 = ~n1387 & n1739 ;
  assign n2484 = ( n1749 & n2482 ) | ( n1749 & ~n2483 ) | ( n2482 & ~n2483 ) ;
  assign n2485 = ( ~n1424 & n2480 ) | ( ~n1424 & n2484 ) | ( n2480 & n2484 ) ;
  assign n2486 = n1447 | n1466 ;
  assign n2487 = ( ~n1453 & n1465 ) | ( ~n1453 & n1746 ) | ( n1465 & n1746 ) ;
  assign n2488 = ( ~n1458 & n2486 ) | ( ~n1458 & n2487 ) | ( n2486 & n2487 ) ;
  assign n2489 = ( n1759 & ~n2360 ) | ( n1759 & n2488 ) | ( ~n2360 & n2488 ) ;
  assign n2490 = n265 | n2489 ;
  assign n2491 = ~n276 & n2490 ;
  assign n2492 = n269 | n276 ;
  assign n2493 = ( ~n1450 & n1454 ) | ( ~n1450 & n1748 ) | ( n1454 & n1748 ) ;
  assign n2494 = ( ~n1461 & n2193 ) | ( ~n1461 & n2493 ) | ( n2193 & n2493 ) ;
  assign n2495 = n265 | n1759 ;
  assign n2496 = ~n276 & n2495 ;
  assign n2497 = ( n2492 & n2494 ) | ( n2492 & ~n2496 ) | ( n2494 & ~n2496 ) ;
  assign n2498 = ( n2485 & ~n2491 ) | ( n2485 & n2497 ) | ( ~n2491 & n2497 ) ;
  assign n2499 = ( ~n289 & n293 ) | ( ~n289 & n1476 ) | ( n293 & n1476 ) ;
  assign n2500 = n286 | n2499 ;
  assign n2501 = ( n282 & ~n292 ) | ( n282 & n298 ) | ( ~n292 & n298 ) ;
  assign n2502 = ( ~n286 & n299 ) | ( ~n286 & n2501 ) | ( n299 & n2501 ) ;
  assign n2503 = ( n2498 & n2500 ) | ( n2498 & ~n2502 ) | ( n2500 & ~n2502 ) ;
  assign n2504 = n2461 & n2503 ;
  assign n2505 = x146 & ~n710 ;
  assign n2506 = ~n546 & n1805 ;
  assign n2507 = ~n500 & n1799 ;
  assign n2508 = n410 | n413 ;
  assign n2509 = n344 | n380 ;
  assign n2510 = x20 | n713 ;
  assign n2511 = ~n316 & n2510 ;
  assign n2512 = ( ~n304 & n322 ) | ( ~n304 & n2511 ) | ( n322 & n2511 ) ;
  assign n2513 = ( ~n337 & n2209 ) | ( ~n337 & n2512 ) | ( n2209 & n2512 ) ;
  assign n2514 = ( ~n1489 & n2509 ) | ( ~n1489 & n2513 ) | ( n2509 & n2513 ) ;
  assign n2515 = ( n1498 & ~n1997 ) | ( n1498 & n2514 ) | ( ~n1997 & n2514 ) ;
  assign n2516 = ( ~n413 & n421 ) | ( ~n413 & n2009 ) | ( n421 & n2009 ) ;
  assign n2517 = ( ~n2508 & n2515 ) | ( ~n2508 & n2516 ) | ( n2515 & n2516 ) ;
  assign n2518 = ( ~n452 & n462 ) | ( ~n452 & n2012 ) | ( n462 & n2012 ) ;
  assign n2519 = ( n1791 & n2517 ) | ( n1791 & ~n2518 ) | ( n2517 & ~n2518 ) ;
  assign n2520 = ( n1795 & ~n2507 ) | ( n1795 & n2519 ) | ( ~n2507 & n2519 ) ;
  assign n2521 = ( ~n1528 & n2506 ) | ( ~n1528 & n2520 ) | ( n2506 & n2520 ) ;
  assign n2522 = ( n600 & ~n1530 ) | ( n600 & n1539 ) | ( ~n1530 & n1539 ) ;
  assign n2523 = ( n1530 & n1534 ) | ( n1530 & ~n1535 ) | ( n1534 & ~n1535 ) ;
  assign n2524 = ( n2521 & ~n2522 ) | ( n2521 & n2523 ) | ( ~n2522 & n2523 ) ;
  assign n2525 = ( n631 & ~n1546 ) | ( n631 & n2524 ) | ( ~n1546 & n2524 ) ;
  assign n2526 = ( n658 & ~n1562 ) | ( n658 & n2251 ) | ( ~n1562 & n2251 ) ;
  assign n2527 = ( n1837 & ~n2404 ) | ( n1837 & n2526 ) | ( ~n2404 & n2526 ) ;
  assign n2528 = n670 | n2527 ;
  assign n2529 = ~n681 & n2528 ;
  assign n2530 = n674 | n681 ;
  assign n2531 = ( n650 & ~n1565 ) | ( n650 & n2248 ) | ( ~n1565 & n2248 ) ;
  assign n2532 = n670 | n1837 ;
  assign n2533 = ~n681 & n2532 ;
  assign n2534 = ( n2530 & n2531 ) | ( n2530 & ~n2533 ) | ( n2531 & ~n2533 ) ;
  assign n2535 = ( n2525 & ~n2529 ) | ( n2525 & n2534 ) | ( ~n2529 & n2534 ) ;
  assign n2536 = ( ~n694 & n698 ) | ( ~n694 & n1575 ) | ( n698 & n1575 ) ;
  assign n2537 = n691 | n2536 ;
  assign n2538 = ( n687 & ~n697 ) | ( n687 & n703 ) | ( ~n697 & n703 ) ;
  assign n2539 = ( ~n691 & n704 ) | ( ~n691 & n2538 ) | ( n704 & n2538 ) ;
  assign n2540 = ( n2535 & n2537 ) | ( n2535 & ~n2539 ) | ( n2537 & ~n2539 ) ;
  assign n2541 = n2505 & n2540 ;
  assign n2542 = x147 & ~n1114 ;
  assign n2543 = ~n951 & n1883 ;
  assign n2544 = ~n905 & n1877 ;
  assign n2545 = n815 | n818 ;
  assign n2546 = n749 | n785 ;
  assign n2547 = x21 | n1117 ;
  assign n2548 = ~n721 & n2547 ;
  assign n2549 = ( ~n709 & n727 ) | ( ~n709 & n2548 ) | ( n727 & n2548 ) ;
  assign n2550 = ( ~n742 & n2265 ) | ( ~n742 & n2549 ) | ( n2265 & n2549 ) ;
  assign n2551 = ( ~n1588 & n2546 ) | ( ~n1588 & n2550 ) | ( n2546 & n2550 ) ;
  assign n2552 = ( n1597 & ~n2067 ) | ( n1597 & n2551 ) | ( ~n2067 & n2551 ) ;
  assign n2553 = ( ~n818 & n826 ) | ( ~n818 & n2079 ) | ( n826 & n2079 ) ;
  assign n2554 = ( ~n2545 & n2552 ) | ( ~n2545 & n2553 ) | ( n2552 & n2553 ) ;
  assign n2555 = ( ~n857 & n867 ) | ( ~n857 & n2082 ) | ( n867 & n2082 ) ;
  assign n2556 = ( n1869 & n2554 ) | ( n1869 & ~n2555 ) | ( n2554 & ~n2555 ) ;
  assign n2557 = ( n1873 & ~n2544 ) | ( n1873 & n2556 ) | ( ~n2544 & n2556 ) ;
  assign n2558 = ( ~n1627 & n2543 ) | ( ~n1627 & n2557 ) | ( n2543 & n2557 ) ;
  assign n2559 = ( n1005 & ~n1629 ) | ( n1005 & n1638 ) | ( ~n1629 & n1638 ) ;
  assign n2560 = ( n1629 & n1633 ) | ( n1629 & ~n1634 ) | ( n1633 & ~n1634 ) ;
  assign n2561 = ( n2558 & ~n2559 ) | ( n2558 & n2560 ) | ( ~n2559 & n2560 ) ;
  assign n2562 = ( n1036 & ~n1645 ) | ( n1036 & n2561 ) | ( ~n1645 & n2561 ) ;
  assign n2563 = ( n1063 & ~n1661 ) | ( n1063 & n2307 ) | ( ~n1661 & n2307 ) ;
  assign n2564 = ( n1915 & ~n2448 ) | ( n1915 & n2563 ) | ( ~n2448 & n2563 ) ;
  assign n2565 = n1074 | n2564 ;
  assign n2566 = ~n1085 & n2565 ;
  assign n2567 = n1078 | n1085 ;
  assign n2568 = ( n1055 & ~n1664 ) | ( n1055 & n2304 ) | ( ~n1664 & n2304 ) ;
  assign n2569 = n1074 | n1915 ;
  assign n2570 = ~n1085 & n2569 ;
  assign n2571 = ( n2567 & n2568 ) | ( n2567 & ~n2570 ) | ( n2568 & ~n2570 ) ;
  assign n2572 = ( n2562 & ~n2566 ) | ( n2562 & n2571 ) | ( ~n2566 & n2571 ) ;
  assign n2573 = ( ~n1098 & n1102 ) | ( ~n1098 & n1673 ) | ( n1102 & n1673 ) ;
  assign n2574 = n1095 | n2573 ;
  assign n2575 = ( n1091 & ~n1101 ) | ( n1091 & n1107 ) | ( ~n1101 & n1107 ) ;
  assign n2576 = ( ~n1095 & n1108 ) | ( ~n1095 & n2575 ) | ( n1108 & n2575 ) ;
  assign n2577 = ( n2572 & n2574 ) | ( n2572 & ~n2576 ) | ( n2574 & ~n2576 ) ;
  assign n2578 = n2542 & n2577 ;
  assign n2579 = x148 & ~n315 ;
  assign n2580 = ~n1355 & n1961 ;
  assign n2581 = ~n1309 & n1955 ;
  assign n2582 = n1219 | n1222 ;
  assign n2583 = n1153 | n1189 ;
  assign n2584 = x22 | n312 ;
  assign n2585 = ~n1125 & n2584 ;
  assign n2586 = ( ~n1113 & n1131 ) | ( ~n1113 & n2585 ) | ( n1131 & n2585 ) ;
  assign n2587 = ( ~n1146 & n2321 ) | ( ~n1146 & n2586 ) | ( n2321 & n2586 ) ;
  assign n2588 = ( ~n1686 & n2583 ) | ( ~n1686 & n2587 ) | ( n2583 & n2587 ) ;
  assign n2589 = ( n1695 & ~n2137 ) | ( n1695 & n2588 ) | ( ~n2137 & n2588 ) ;
  assign n2590 = ( ~n1222 & n1230 ) | ( ~n1222 & n2149 ) | ( n1230 & n2149 ) ;
  assign n2591 = ( ~n2582 & n2589 ) | ( ~n2582 & n2590 ) | ( n2589 & n2590 ) ;
  assign n2592 = ( ~n1261 & n1271 ) | ( ~n1261 & n2152 ) | ( n1271 & n2152 ) ;
  assign n2593 = ( n1947 & n2591 ) | ( n1947 & ~n2592 ) | ( n2591 & ~n2592 ) ;
  assign n2594 = ( n1951 & ~n2581 ) | ( n1951 & n2593 ) | ( ~n2581 & n2593 ) ;
  assign n2595 = ( ~n1725 & n2580 ) | ( ~n1725 & n2594 ) | ( n2580 & n2594 ) ;
  assign n2596 = ( n1409 & ~n1727 ) | ( n1409 & n1736 ) | ( ~n1727 & n1736 ) ;
  assign n2597 = ( n1727 & n1731 ) | ( n1727 & ~n1732 ) | ( n1731 & ~n1732 ) ;
  assign n2598 = ( n2595 & ~n2596 ) | ( n2595 & n2597 ) | ( ~n2596 & n2597 ) ;
  assign n2599 = ( n1440 & ~n1743 ) | ( n1440 & n2598 ) | ( ~n1743 & n2598 ) ;
  assign n2600 = ( n1467 & ~n1756 ) | ( n1467 & n2363 ) | ( ~n1756 & n2363 ) ;
  assign n2601 = ( n1991 & ~n2492 ) | ( n1991 & n2600 ) | ( ~n2492 & n2600 ) ;
  assign n2602 = n273 | n2601 ;
  assign n2603 = ~n280 & n2602 ;
  assign n2604 = ( n1459 & ~n1759 ) | ( n1459 & n2360 ) | ( ~n1759 & n2360 ) ;
  assign n2605 = n273 | n1991 ;
  assign n2606 = ~n280 & n2605 ;
  assign n2607 = ( n281 & n2604 ) | ( n281 & ~n2606 ) | ( n2604 & ~n2606 ) ;
  assign n2608 = ( n2599 & ~n2603 ) | ( n2599 & n2607 ) | ( ~n2603 & n2607 ) ;
  assign n2609 = ( n293 & ~n307 ) | ( n293 & n1479 ) | ( ~n307 & n1479 ) ;
  assign n2610 = n310 | n2609 ;
  assign n2611 = ( n300 & ~n310 ) | ( n300 & n311 ) | ( ~n310 & n311 ) ;
  assign n2612 = ( n2608 & n2610 ) | ( n2608 & ~n2611 ) | ( n2610 & ~n2611 ) ;
  assign n2613 = n2579 & n2612 ;
  assign n2614 = x149 & ~n720 ;
  assign n2615 = ~n543 & n2035 ;
  assign n2616 = ~n484 & n2026 ;
  assign n2617 = n391 | n1502 ;
  assign n2618 = n368 | n381 ;
  assign n2619 = x23 | n717 ;
  assign n2620 = ~n303 & n2619 ;
  assign n2621 = ( ~n333 & n348 ) | ( ~n333 & n2620 ) | ( n348 & n2620 ) ;
  assign n2622 = ( ~n341 & n2377 ) | ( ~n341 & n2621 ) | ( n2377 & n2621 ) ;
  assign n2623 = ( ~n1774 & n2618 ) | ( ~n1774 & n2622 ) | ( n2618 & n2622 ) ;
  assign n2624 = ( n1782 & ~n2208 ) | ( n1782 & n2623 ) | ( ~n2208 & n2623 ) ;
  assign n2625 = ( ~n391 & n395 ) | ( ~n391 & n422 ) | ( n395 & n422 ) ;
  assign n2626 = ( ~n2617 & n2624 ) | ( ~n2617 & n2625 ) | ( n2624 & n2625 ) ;
  assign n2627 = ( ~n436 & n463 ) | ( ~n436 & n464 ) | ( n463 & n464 ) ;
  assign n2628 = ( n2018 & n2626 ) | ( n2018 & ~n2627 ) | ( n2626 & ~n2627 ) ;
  assign n2629 = ( n2022 & ~n2616 ) | ( n2022 & n2628 ) | ( ~n2616 & n2628 ) ;
  assign n2630 = ( ~n1809 & n2615 ) | ( ~n1809 & n2629 ) | ( n2615 & n2629 ) ;
  assign n2631 = ( n610 & ~n624 ) | ( n610 & n1818 ) | ( ~n624 & n1818 ) ;
  assign n2632 = ( n624 & n1813 ) | ( n624 & ~n1814 ) | ( n1813 & ~n1814 ) ;
  assign n2633 = ( n2630 & ~n2631 ) | ( n2630 & n2632 ) | ( ~n2631 & n2632 ) ;
  assign n2634 = ( n1556 & ~n1824 ) | ( n1556 & n2633 ) | ( ~n1824 & n2633 ) ;
  assign n2635 = ( n1566 & ~n1834 ) | ( n1566 & n2407 ) | ( ~n1834 & n2407 ) ;
  assign n2636 = ( n2061 & ~n2530 ) | ( n2061 & n2635 ) | ( ~n2530 & n2635 ) ;
  assign n2637 = n678 | n2636 ;
  assign n2638 = ~n685 & n2637 ;
  assign n2639 = ( n1563 & ~n1837 ) | ( n1563 & n2404 ) | ( ~n1837 & n2404 ) ;
  assign n2640 = n678 | n2061 ;
  assign n2641 = ~n685 & n2640 ;
  assign n2642 = ( n686 & n2639 ) | ( n686 & ~n2641 ) | ( n2639 & ~n2641 ) ;
  assign n2643 = ( n2634 & ~n2638 ) | ( n2634 & n2642 ) | ( ~n2638 & n2642 ) ;
  assign n2644 = ( n698 & ~n712 ) | ( n698 & n1578 ) | ( ~n712 & n1578 ) ;
  assign n2645 = n715 | n2644 ;
  assign n2646 = ( n705 & ~n715 ) | ( n705 & n716 ) | ( ~n715 & n716 ) ;
  assign n2647 = ( n2643 & n2645 ) | ( n2643 & ~n2646 ) | ( n2645 & ~n2646 ) ;
  assign n2648 = n2614 & n2647 ;
  assign n2649 = x150 & ~n1124 ;
  assign n2650 = ~n948 & n2105 ;
  assign n2651 = ~n889 & n2096 ;
  assign n2652 = n796 | n1601 ;
  assign n2653 = n773 | n786 ;
  assign n2654 = x24 | n1121 ;
  assign n2655 = ~n708 & n2654 ;
  assign n2656 = ( ~n738 & n753 ) | ( ~n738 & n2655 ) | ( n753 & n2655 ) ;
  assign n2657 = ( ~n746 & n2421 ) | ( ~n746 & n2656 ) | ( n2421 & n2656 ) ;
  assign n2658 = ( ~n1852 & n2653 ) | ( ~n1852 & n2657 ) | ( n2653 & n2657 ) ;
  assign n2659 = ( n1860 & ~n2264 ) | ( n1860 & n2658 ) | ( ~n2264 & n2658 ) ;
  assign n2660 = ( ~n796 & n800 ) | ( ~n796 & n827 ) | ( n800 & n827 ) ;
  assign n2661 = ( ~n2652 & n2659 ) | ( ~n2652 & n2660 ) | ( n2659 & n2660 ) ;
  assign n2662 = ( ~n841 & n868 ) | ( ~n841 & n869 ) | ( n868 & n869 ) ;
  assign n2663 = ( n2088 & n2661 ) | ( n2088 & ~n2662 ) | ( n2661 & ~n2662 ) ;
  assign n2664 = ( n2092 & ~n2651 ) | ( n2092 & n2663 ) | ( ~n2651 & n2663 ) ;
  assign n2665 = ( ~n1887 & n2650 ) | ( ~n1887 & n2664 ) | ( n2650 & n2664 ) ;
  assign n2666 = ( n1015 & ~n1029 ) | ( n1015 & n1896 ) | ( ~n1029 & n1896 ) ;
  assign n2667 = ( n1029 & n1891 ) | ( n1029 & ~n1892 ) | ( n1891 & ~n1892 ) ;
  assign n2668 = ( n2665 & ~n2666 ) | ( n2665 & n2667 ) | ( ~n2666 & n2667 ) ;
  assign n2669 = ( n1655 & ~n1902 ) | ( n1655 & n2668 ) | ( ~n1902 & n2668 ) ;
  assign n2670 = ( n1665 & ~n1912 ) | ( n1665 & n2451 ) | ( ~n1912 & n2451 ) ;
  assign n2671 = ( n2131 & ~n2567 ) | ( n2131 & n2670 ) | ( ~n2567 & n2670 ) ;
  assign n2672 = n1082 | n2671 ;
  assign n2673 = ~n1089 & n2672 ;
  assign n2674 = ( n1662 & ~n1915 ) | ( n1662 & n2448 ) | ( ~n1915 & n2448 ) ;
  assign n2675 = n1082 | n2131 ;
  assign n2676 = ~n1089 & n2675 ;
  assign n2677 = ( n1090 & n2674 ) | ( n1090 & ~n2676 ) | ( n2674 & ~n2676 ) ;
  assign n2678 = ( n2669 & ~n2673 ) | ( n2669 & n2677 ) | ( ~n2673 & n2677 ) ;
  assign n2679 = ( n1102 & ~n1116 ) | ( n1102 & n1676 ) | ( ~n1116 & n1676 ) ;
  assign n2680 = n1119 | n2679 ;
  assign n2681 = ( n1109 & ~n1119 ) | ( n1109 & n1120 ) | ( ~n1119 & n1120 ) ;
  assign n2682 = ( n2678 & n2680 ) | ( n2678 & ~n2681 ) | ( n2680 & ~n2681 ) ;
  assign n2683 = n2649 & n2682 ;
  assign n2684 = x151 & ~n302 ;
  assign n2685 = ~n1352 & n2175 ;
  assign n2686 = ~n1293 & n2166 ;
  assign n2687 = n1200 | n1699 ;
  assign n2688 = n1177 | n1190 ;
  assign n2689 = x25 | n345 ;
  assign n2690 = ~n1112 & n2689 ;
  assign n2691 = ( ~n1142 & n1157 ) | ( ~n1142 & n2690 ) | ( n1157 & n2690 ) ;
  assign n2692 = ( ~n1150 & n2465 ) | ( ~n1150 & n2691 ) | ( n2465 & n2691 ) ;
  assign n2693 = ( ~n1930 & n2688 ) | ( ~n1930 & n2692 ) | ( n2688 & n2692 ) ;
  assign n2694 = ( n1938 & ~n2320 ) | ( n1938 & n2693 ) | ( ~n2320 & n2693 ) ;
  assign n2695 = ( ~n1200 & n1204 ) | ( ~n1200 & n1231 ) | ( n1204 & n1231 ) ;
  assign n2696 = ( ~n2687 & n2694 ) | ( ~n2687 & n2695 ) | ( n2694 & n2695 ) ;
  assign n2697 = ( ~n1245 & n1272 ) | ( ~n1245 & n1273 ) | ( n1272 & n1273 ) ;
  assign n2698 = ( n2158 & n2696 ) | ( n2158 & ~n2697 ) | ( n2696 & ~n2697 ) ;
  assign n2699 = ( n2162 & ~n2686 ) | ( n2162 & n2698 ) | ( ~n2686 & n2698 ) ;
  assign n2700 = ( ~n1965 & n2685 ) | ( ~n1965 & n2699 ) | ( n2685 & n2699 ) ;
  assign n2701 = ( n1419 & ~n1433 ) | ( n1419 & n1974 ) | ( ~n1433 & n1974 ) ;
  assign n2702 = ( n1433 & n1969 ) | ( n1433 & ~n1970 ) | ( n1969 & ~n1970 ) ;
  assign n2703 = ( n2700 & ~n2701 ) | ( n2700 & n2702 ) | ( ~n2701 & n2702 ) ;
  assign n2704 = ( n1753 & ~n1980 ) | ( n1753 & n2703 ) | ( ~n1980 & n2703 ) ;
  assign n2705 = ( ~n269 & n1760 ) | ( ~n269 & n2495 ) | ( n1760 & n2495 ) ;
  assign n2706 = ( ~n281 & n282 ) | ( ~n281 & n2705 ) | ( n282 & n2705 ) ;
  assign n2707 = n297 | n2706 ;
  assign n2708 = ~n292 & n2707 ;
  assign n2709 = ( n1757 & ~n1991 ) | ( n1757 & n2492 ) | ( ~n1991 & n2492 ) ;
  assign n2710 = n282 | n297 ;
  assign n2711 = ~n292 & n2710 ;
  assign n2712 = ( n1477 & n2709 ) | ( n1477 & ~n2711 ) | ( n2709 & ~n2711 ) ;
  assign n2713 = ( n2704 & ~n2708 ) | ( n2704 & n2712 ) | ( ~n2708 & n2712 ) ;
  assign n2714 = ( ~n317 & n321 ) | ( ~n317 & n1479 ) | ( n321 & n1479 ) ;
  assign n2715 = n314 | n2714 ;
  assign n2716 = ( ~n314 & n318 ) | ( ~n314 & n1481 ) | ( n318 & n1481 ) ;
  assign n2717 = ( n2713 & n2715 ) | ( n2713 & ~n2716 ) | ( n2715 & ~n2716 ) ;
  assign n2718 = n2684 & n2717 ;
  assign n2719 = n362 | n382 ;
  assign n2720 = x26 | n750 ;
  assign n2721 = ~n332 & n2720 ;
  assign n2722 = ( ~n340 & n349 ) | ( ~n340 & n2721 ) | ( n349 & n2721 ) ;
  assign n2723 = ( ~n1488 & n2509 ) | ( ~n1488 & n2722 ) | ( n2509 & n2722 ) ;
  assign n2724 = ( ~n374 & n2719 ) | ( ~n374 & n2723 ) | ( n2719 & n2723 ) ;
  assign n2725 = n460 | n1785 ;
  assign n2726 = ( ~n460 & n1501 ) | ( ~n460 & n1507 ) | ( n1501 & n1507 ) ;
  assign n2727 = ( n2376 & n2725 ) | ( n2376 & ~n2726 ) | ( n2725 & ~n2726 ) ;
  assign n2728 = ( n2009 & ~n2725 ) | ( n2009 & n2726 ) | ( ~n2725 & n2726 ) ;
  assign n2729 = ( n2724 & ~n2727 ) | ( n2724 & n2728 ) | ( ~n2727 & n2728 ) ;
  assign n2730 = ~n478 & n2223 ;
  assign n2731 = ( ~n430 & n439 ) | ( ~n430 & n1515 ) | ( n439 & n1515 ) ;
  assign n2732 = ( ~n503 & n2730 ) | ( ~n503 & n2731 ) | ( n2730 & n2731 ) ;
  assign n2733 = ( n455 & n503 ) | ( n455 & ~n2730 ) | ( n503 & ~n2730 ) ;
  assign n2734 = ( n2729 & ~n2732 ) | ( n2729 & n2733 ) | ( ~n2732 & n2733 ) ;
  assign n2735 = ~n534 & n2231 ;
  assign n2736 = ( n625 & n2040 ) | ( n625 & ~n2041 ) | ( n2040 & ~n2041 ) ;
  assign n2737 = ( n591 & ~n625 ) | ( n591 & n2045 ) | ( ~n625 & n2045 ) ;
  assign n2738 = ( n2735 & n2736 ) | ( n2735 & ~n2737 ) | ( n2736 & ~n2737 ) ;
  assign n2739 = ( n1831 & ~n2050 ) | ( n1831 & n2738 ) | ( ~n2050 & n2738 ) ;
  assign n2740 = ( n2031 & ~n2736 ) | ( n2031 & n2737 ) | ( ~n2736 & n2737 ) ;
  assign n2741 = ( ~n1831 & n2050 ) | ( ~n1831 & n2740 ) | ( n2050 & n2740 ) ;
  assign n2742 = ( n2734 & n2739 ) | ( n2734 & ~n2741 ) | ( n2739 & ~n2741 ) ;
  assign n2743 = x152 & ~n707 ;
  assign n2744 = n687 | n702 ;
  assign n2745 = ( ~n674 & n1838 ) | ( ~n674 & n2532 ) | ( n1838 & n2532 ) ;
  assign n2746 = ( ~n2411 & n2744 ) | ( ~n2411 & n2745 ) | ( n2744 & n2745 ) ;
  assign n2747 = ~n697 & n2746 ;
  assign n2748 = ( ~n722 & n726 ) | ( ~n722 & n1578 ) | ( n726 & n1578 ) ;
  assign n2749 = n719 | n2748 ;
  assign n2750 = ( ~n719 & n723 ) | ( ~n719 & n1580 ) | ( n723 & n1580 ) ;
  assign n2751 = ( n2747 & ~n2749 ) | ( n2747 & n2750 ) | ( ~n2749 & n2750 ) ;
  assign n2752 = n2743 & ~n2751 ;
  assign n2753 = ( n1835 & ~n2061 ) | ( n1835 & n2530 ) | ( ~n2061 & n2530 ) ;
  assign n2754 = ( n1576 & ~n2538 ) | ( n1576 & n2753 ) | ( ~n2538 & n2753 ) ;
  assign n2755 = ( n2749 & ~n2750 ) | ( n2749 & n2754 ) | ( ~n2750 & n2754 ) ;
  assign n2756 = n2743 & n2755 ;
  assign n2757 = ( n2742 & n2752 ) | ( n2742 & n2756 ) | ( n2752 & n2756 ) ;
  assign n2758 = n767 | n787 ;
  assign n2759 = x27 | n1154 ;
  assign n2760 = ~n737 & n2759 ;
  assign n2761 = ( ~n745 & n754 ) | ( ~n745 & n2760 ) | ( n754 & n2760 ) ;
  assign n2762 = ( ~n1587 & n2546 ) | ( ~n1587 & n2761 ) | ( n2546 & n2761 ) ;
  assign n2763 = ( ~n779 & n2758 ) | ( ~n779 & n2762 ) | ( n2758 & n2762 ) ;
  assign n2764 = n865 | n1863 ;
  assign n2765 = ( ~n865 & n1600 ) | ( ~n865 & n1606 ) | ( n1600 & n1606 ) ;
  assign n2766 = ( n2420 & n2764 ) | ( n2420 & ~n2765 ) | ( n2764 & ~n2765 ) ;
  assign n2767 = ( n2079 & ~n2764 ) | ( n2079 & n2765 ) | ( ~n2764 & n2765 ) ;
  assign n2768 = ( n2763 & ~n2766 ) | ( n2763 & n2767 ) | ( ~n2766 & n2767 ) ;
  assign n2769 = ~n883 & n2279 ;
  assign n2770 = ( ~n835 & n844 ) | ( ~n835 & n1614 ) | ( n844 & n1614 ) ;
  assign n2771 = ( ~n908 & n2769 ) | ( ~n908 & n2770 ) | ( n2769 & n2770 ) ;
  assign n2772 = ( n860 & n908 ) | ( n860 & ~n2769 ) | ( n908 & ~n2769 ) ;
  assign n2773 = ( n2768 & ~n2771 ) | ( n2768 & n2772 ) | ( ~n2771 & n2772 ) ;
  assign n2774 = ~n939 & n2287 ;
  assign n2775 = ( n1030 & n2110 ) | ( n1030 & ~n2111 ) | ( n2110 & ~n2111 ) ;
  assign n2776 = ( n996 & ~n1030 ) | ( n996 & n2115 ) | ( ~n1030 & n2115 ) ;
  assign n2777 = ( n2774 & n2775 ) | ( n2774 & ~n2776 ) | ( n2775 & ~n2776 ) ;
  assign n2778 = ( n1909 & ~n2120 ) | ( n1909 & n2777 ) | ( ~n2120 & n2777 ) ;
  assign n2779 = ( n2101 & ~n2775 ) | ( n2101 & n2776 ) | ( ~n2775 & n2776 ) ;
  assign n2780 = ( ~n1909 & n2120 ) | ( ~n1909 & n2779 ) | ( n2120 & n2779 ) ;
  assign n2781 = ( n2773 & n2778 ) | ( n2773 & ~n2780 ) | ( n2778 & ~n2780 ) ;
  assign n2782 = x153 & ~n1111 ;
  assign n2783 = n1091 | n1106 ;
  assign n2784 = ( ~n1078 & n1916 ) | ( ~n1078 & n2569 ) | ( n1916 & n2569 ) ;
  assign n2785 = ( ~n2455 & n2783 ) | ( ~n2455 & n2784 ) | ( n2783 & n2784 ) ;
  assign n2786 = ~n1101 & n2785 ;
  assign n2787 = ( ~n1126 & n1130 ) | ( ~n1126 & n1676 ) | ( n1130 & n1676 ) ;
  assign n2788 = n1123 | n2787 ;
  assign n2789 = ( ~n1123 & n1127 ) | ( ~n1123 & n1678 ) | ( n1127 & n1678 ) ;
  assign n2790 = ( n2786 & ~n2788 ) | ( n2786 & n2789 ) | ( ~n2788 & n2789 ) ;
  assign n2791 = n2782 & ~n2790 ;
  assign n2792 = ( n1913 & ~n2131 ) | ( n1913 & n2567 ) | ( ~n2131 & n2567 ) ;
  assign n2793 = ( n1674 & ~n2575 ) | ( n1674 & n2792 ) | ( ~n2575 & n2792 ) ;
  assign n2794 = ( n2788 & ~n2789 ) | ( n2788 & n2793 ) | ( ~n2789 & n2793 ) ;
  assign n2795 = n2782 & n2794 ;
  assign n2796 = ( n2781 & n2791 ) | ( n2781 & n2795 ) | ( n2791 & n2795 ) ;
  assign n2797 = n1171 | n1191 ;
  assign n2798 = x28 | n334 ;
  assign n2799 = ~n1141 & n2798 ;
  assign n2800 = ( ~n1149 & n1158 ) | ( ~n1149 & n2799 ) | ( n1158 & n2799 ) ;
  assign n2801 = ( ~n1685 & n2583 ) | ( ~n1685 & n2800 ) | ( n2583 & n2800 ) ;
  assign n2802 = ( ~n1183 & n2797 ) | ( ~n1183 & n2801 ) | ( n2797 & n2801 ) ;
  assign n2803 = n1269 | n1941 ;
  assign n2804 = ( ~n1269 & n1698 ) | ( ~n1269 & n1704 ) | ( n1698 & n1704 ) ;
  assign n2805 = ( n2464 & n2803 ) | ( n2464 & ~n2804 ) | ( n2803 & ~n2804 ) ;
  assign n2806 = ( n2149 & ~n2803 ) | ( n2149 & n2804 ) | ( ~n2803 & n2804 ) ;
  assign n2807 = ( n2802 & ~n2805 ) | ( n2802 & n2806 ) | ( ~n2805 & n2806 ) ;
  assign n2808 = ~n1287 & n2335 ;
  assign n2809 = ( ~n1239 & n1248 ) | ( ~n1239 & n1712 ) | ( n1248 & n1712 ) ;
  assign n2810 = ( ~n1312 & n2808 ) | ( ~n1312 & n2809 ) | ( n2808 & n2809 ) ;
  assign n2811 = ( n1264 & n1312 ) | ( n1264 & ~n2808 ) | ( n1312 & ~n2808 ) ;
  assign n2812 = ( n2807 & ~n2810 ) | ( n2807 & n2811 ) | ( ~n2810 & n2811 ) ;
  assign n2813 = ~n1343 & n2343 ;
  assign n2814 = ( n1434 & n2180 ) | ( n1434 & ~n2181 ) | ( n2180 & ~n2181 ) ;
  assign n2815 = ( n1400 & ~n1434 ) | ( n1400 & n2185 ) | ( ~n1434 & n2185 ) ;
  assign n2816 = ( n2813 & n2814 ) | ( n2813 & ~n2815 ) | ( n2814 & ~n2815 ) ;
  assign n2817 = ( n1987 & ~n2190 ) | ( n1987 & n2816 ) | ( ~n2190 & n2816 ) ;
  assign n2818 = ( n2171 & ~n2814 ) | ( n2171 & n2815 ) | ( ~n2814 & n2815 ) ;
  assign n2819 = ( ~n1987 & n2190 ) | ( ~n1987 & n2818 ) | ( n2190 & n2818 ) ;
  assign n2820 = ( n2812 & n2817 ) | ( n2812 & ~n2819 ) | ( n2817 & ~n2819 ) ;
  assign n2821 = x154 & ~n331 ;
  assign n2822 = n289 | n298 ;
  assign n2823 = ( ~n277 & n1992 ) | ( ~n277 & n2605 ) | ( n1992 & n2605 ) ;
  assign n2824 = ( ~n2499 & n2822 ) | ( ~n2499 & n2823 ) | ( n2822 & n2823 ) ;
  assign n2825 = ~n286 & n2824 ;
  assign n2826 = n323 | n347 ;
  assign n2827 = ( n319 & ~n347 ) | ( n319 & n1483 ) | ( ~n347 & n1483 ) ;
  assign n2828 = ( n2825 & ~n2826 ) | ( n2825 & n2827 ) | ( ~n2826 & n2827 ) ;
  assign n2829 = n2821 & ~n2828 ;
  assign n2830 = ( n281 & ~n282 ) | ( n281 & n1989 ) | ( ~n282 & n1989 ) ;
  assign n2831 = ( n294 & ~n300 ) | ( n294 & n2830 ) | ( ~n300 & n2830 ) ;
  assign n2832 = ( n2826 & ~n2827 ) | ( n2826 & n2831 ) | ( ~n2827 & n2831 ) ;
  assign n2833 = n2821 & n2832 ;
  assign n2834 = ( n2820 & n2829 ) | ( n2820 & n2833 ) | ( n2829 & n2833 ) ;
  assign n2835 = x29 | n739 ;
  assign n2836 = ~n339 & n2835 ;
  assign n2837 = ( ~n327 & n344 ) | ( ~n327 & n2836 ) | ( n344 & n2836 ) ;
  assign n2838 = ( ~n369 & n2618 ) | ( ~n369 & n2837 ) | ( n2618 & n2837 ) ;
  assign n2839 = ( n377 & ~n1494 ) | ( n377 & n2838 ) | ( ~n1494 & n2838 ) ;
  assign n2840 = n445 | n2012 ;
  assign n2841 = ( ~n445 & n449 ) | ( ~n445 & n1790 ) | ( n449 & n1790 ) ;
  assign n2842 = ( n2508 & n2840 ) | ( n2508 & ~n2841 ) | ( n2840 & ~n2841 ) ;
  assign n2843 = ( n422 & ~n2840 ) | ( n422 & n2841 ) | ( ~n2840 & n2841 ) ;
  assign n2844 = ( n2839 & ~n2842 ) | ( n2839 & n2843 ) | ( ~n2842 & n2843 ) ;
  assign n2845 = ~n474 & n515 ;
  assign n2846 = ( ~n496 & n1511 ) | ( ~n496 & n1797 ) | ( n1511 & n1797 ) ;
  assign n2847 = ( ~n1522 & n2845 ) | ( ~n1522 & n2846 ) | ( n2845 & n2846 ) ;
  assign n2848 = ( n1513 & n1522 ) | ( n1513 & ~n2845 ) | ( n1522 & ~n2845 ) ;
  assign n2849 = ( n2844 & ~n2847 ) | ( n2844 & n2848 ) | ( ~n2847 & n2848 ) ;
  assign n2850 = n556 & ~n559 ;
  assign n2851 = ( ~n596 & n597 ) | ( ~n596 & n2235 ) | ( n597 & n2235 ) ;
  assign n2852 = ( n588 & ~n597 ) | ( n588 & n2239 ) | ( ~n597 & n2239 ) ;
  assign n2853 = ( n2850 & n2851 ) | ( n2850 & ~n2852 ) | ( n2851 & ~n2852 ) ;
  assign n2854 = ( n2057 & ~n2245 ) | ( n2057 & n2853 ) | ( ~n2245 & n2853 ) ;
  assign n2855 = ( n2228 & ~n2851 ) | ( n2228 & n2852 ) | ( ~n2851 & n2852 ) ;
  assign n2856 = ( ~n2057 & n2245 ) | ( ~n2057 & n2855 ) | ( n2245 & n2855 ) ;
  assign n2857 = ( n2849 & n2854 ) | ( n2849 & ~n2856 ) | ( n2854 & ~n2856 ) ;
  assign n2858 = x155 & ~n736 ;
  assign n2859 = n694 | n703 ;
  assign n2860 = ( ~n682 & n2062 ) | ( ~n682 & n2640 ) | ( n2062 & n2640 ) ;
  assign n2861 = ( ~n2536 & n2859 ) | ( ~n2536 & n2860 ) | ( n2859 & n2860 ) ;
  assign n2862 = ~n691 & n2861 ;
  assign n2863 = n728 | n752 ;
  assign n2864 = ( n724 & ~n752 ) | ( n724 & n1582 ) | ( ~n752 & n1582 ) ;
  assign n2865 = ( n2862 & ~n2863 ) | ( n2862 & n2864 ) | ( ~n2863 & n2864 ) ;
  assign n2866 = n2858 & ~n2865 ;
  assign n2867 = ( n686 & ~n687 ) | ( n686 & n2059 ) | ( ~n687 & n2059 ) ;
  assign n2868 = ( n699 & ~n705 ) | ( n699 & n2867 ) | ( ~n705 & n2867 ) ;
  assign n2869 = ( n2863 & ~n2864 ) | ( n2863 & n2868 ) | ( ~n2864 & n2868 ) ;
  assign n2870 = n2858 & n2869 ;
  assign n2871 = ( n2857 & n2866 ) | ( n2857 & n2870 ) | ( n2866 & n2870 ) ;
  assign n2872 = x30 | n1143 ;
  assign n2873 = ~n744 & n2872 ;
  assign n2874 = ( ~n732 & n749 ) | ( ~n732 & n2873 ) | ( n749 & n2873 ) ;
  assign n2875 = ( ~n774 & n2653 ) | ( ~n774 & n2874 ) | ( n2653 & n2874 ) ;
  assign n2876 = ( n782 & ~n1593 ) | ( n782 & n2875 ) | ( ~n1593 & n2875 ) ;
  assign n2877 = n850 | n2082 ;
  assign n2878 = ( ~n850 & n854 ) | ( ~n850 & n1868 ) | ( n854 & n1868 ) ;
  assign n2879 = ( n2545 & n2877 ) | ( n2545 & ~n2878 ) | ( n2877 & ~n2878 ) ;
  assign n2880 = ( n827 & ~n2877 ) | ( n827 & n2878 ) | ( ~n2877 & n2878 ) ;
  assign n2881 = ( n2876 & ~n2879 ) | ( n2876 & n2880 ) | ( ~n2879 & n2880 ) ;
  assign n2882 = ~n879 & n920 ;
  assign n2883 = ( ~n901 & n1610 ) | ( ~n901 & n1875 ) | ( n1610 & n1875 ) ;
  assign n2884 = ( ~n1621 & n2882 ) | ( ~n1621 & n2883 ) | ( n2882 & n2883 ) ;
  assign n2885 = ( n1612 & n1621 ) | ( n1612 & ~n2882 ) | ( n1621 & ~n2882 ) ;
  assign n2886 = ( n2881 & ~n2884 ) | ( n2881 & n2885 ) | ( ~n2884 & n2885 ) ;
  assign n2887 = n961 & ~n964 ;
  assign n2888 = ( ~n1001 & n1002 ) | ( ~n1001 & n2291 ) | ( n1002 & n2291 ) ;
  assign n2889 = ( n993 & ~n1002 ) | ( n993 & n2295 ) | ( ~n1002 & n2295 ) ;
  assign n2890 = ( n2887 & n2888 ) | ( n2887 & ~n2889 ) | ( n2888 & ~n2889 ) ;
  assign n2891 = ( n2127 & ~n2301 ) | ( n2127 & n2890 ) | ( ~n2301 & n2890 ) ;
  assign n2892 = ( n2284 & ~n2888 ) | ( n2284 & n2889 ) | ( ~n2888 & n2889 ) ;
  assign n2893 = ( ~n2127 & n2301 ) | ( ~n2127 & n2892 ) | ( n2301 & n2892 ) ;
  assign n2894 = ( n2886 & n2891 ) | ( n2886 & ~n2893 ) | ( n2891 & ~n2893 ) ;
  assign n2895 = x156 & ~n1140 ;
  assign n2896 = n1098 | n1107 ;
  assign n2897 = ( ~n1086 & n2132 ) | ( ~n1086 & n2675 ) | ( n2132 & n2675 ) ;
  assign n2898 = ( ~n2573 & n2896 ) | ( ~n2573 & n2897 ) | ( n2896 & n2897 ) ;
  assign n2899 = ~n1095 & n2898 ;
  assign n2900 = n1132 | n1156 ;
  assign n2901 = ( n1128 & ~n1156 ) | ( n1128 & n1680 ) | ( ~n1156 & n1680 ) ;
  assign n2902 = ( n2899 & ~n2900 ) | ( n2899 & n2901 ) | ( ~n2900 & n2901 ) ;
  assign n2903 = n2895 & ~n2902 ;
  assign n2904 = ( n1090 & ~n1091 ) | ( n1090 & n2129 ) | ( ~n1091 & n2129 ) ;
  assign n2905 = ( n1103 & ~n1109 ) | ( n1103 & n2904 ) | ( ~n1109 & n2904 ) ;
  assign n2906 = ( n2900 & ~n2901 ) | ( n2900 & n2905 ) | ( ~n2901 & n2905 ) ;
  assign n2907 = n2895 & n2906 ;
  assign n2908 = ( n2894 & n2903 ) | ( n2894 & n2907 ) | ( n2903 & n2907 ) ;
  assign n2909 = x31 | n328 ;
  assign n2910 = ~n1148 & n2909 ;
  assign n2911 = ( ~n1136 & n1153 ) | ( ~n1136 & n2910 ) | ( n1153 & n2910 ) ;
  assign n2912 = ( ~n1178 & n2688 ) | ( ~n1178 & n2911 ) | ( n2688 & n2911 ) ;
  assign n2913 = ( n1186 & ~n1691 ) | ( n1186 & n2912 ) | ( ~n1691 & n2912 ) ;
  assign n2914 = n1254 | n2152 ;
  assign n2915 = ( ~n1254 & n1258 ) | ( ~n1254 & n1946 ) | ( n1258 & n1946 ) ;
  assign n2916 = ( n2582 & n2914 ) | ( n2582 & ~n2915 ) | ( n2914 & ~n2915 ) ;
  assign n2917 = ( n1231 & ~n2914 ) | ( n1231 & n2915 ) | ( ~n2914 & n2915 ) ;
  assign n2918 = ( n2913 & ~n2916 ) | ( n2913 & n2917 ) | ( ~n2916 & n2917 ) ;
  assign n2919 = ~n1283 & n1324 ;
  assign n2920 = ( ~n1305 & n1708 ) | ( ~n1305 & n1953 ) | ( n1708 & n1953 ) ;
  assign n2921 = ( ~n1719 & n2919 ) | ( ~n1719 & n2920 ) | ( n2919 & n2920 ) ;
  assign n2922 = ( n1710 & n1719 ) | ( n1710 & ~n2919 ) | ( n1719 & ~n2919 ) ;
  assign n2923 = ( n2918 & ~n2921 ) | ( n2918 & n2922 ) | ( ~n2921 & n2922 ) ;
  assign n2924 = n1365 & ~n1368 ;
  assign n2925 = ( ~n1405 & n1406 ) | ( ~n1405 & n2347 ) | ( n1406 & n2347 ) ;
  assign n2926 = ( n1397 & ~n1406 ) | ( n1397 & n2351 ) | ( ~n1406 & n2351 ) ;
  assign n2927 = ( n2924 & n2925 ) | ( n2924 & ~n2926 ) | ( n2925 & ~n2926 ) ;
  assign n2928 = ( n2197 & ~n2357 ) | ( n2197 & n2927 ) | ( ~n2357 & n2927 ) ;
  assign n2929 = ( n2340 & ~n2925 ) | ( n2340 & n2926 ) | ( ~n2925 & n2926 ) ;
  assign n2930 = ( ~n2197 & n2357 ) | ( ~n2197 & n2929 ) | ( n2357 & n2929 ) ;
  assign n2931 = ( n2923 & n2928 ) | ( n2923 & ~n2930 ) | ( n2928 & ~n2930 ) ;
  assign n2932 = x157 & ~n338 ;
  assign n2933 = n299 | n307 ;
  assign n2934 = ( ~n1476 & n2201 ) | ( ~n1476 & n2710 ) | ( n2201 & n2710 ) ;
  assign n2935 = ( ~n2609 & n2933 ) | ( ~n2609 & n2934 ) | ( n2933 & n2934 ) ;
  assign n2936 = ~n310 & n2935 ;
  assign n2937 = n336 | n1486 ;
  assign n2938 = ( ~n336 & n337 ) | ( ~n336 & n1484 ) | ( n337 & n1484 ) ;
  assign n2939 = ( n2936 & ~n2937 ) | ( n2936 & n2938 ) | ( ~n2937 & n2938 ) ;
  assign n2940 = n2932 & ~n2939 ;
  assign n2941 = ( ~n298 & n1477 ) | ( ~n298 & n2199 ) | ( n1477 & n2199 ) ;
  assign n2942 = ( n1480 & ~n1481 ) | ( n1480 & n2941 ) | ( ~n1481 & n2941 ) ;
  assign n2943 = ( n2937 & ~n2938 ) | ( n2937 & n2942 ) | ( ~n2938 & n2942 ) ;
  assign n2944 = n2932 & n2943 ;
  assign n2945 = ( n2931 & n2940 ) | ( n2931 & n2944 ) | ( n2940 & n2944 ) ;
  assign n2946 = x32 | n733 ;
  assign n2947 = ~n326 & n2946 ;
  assign n2948 = ( ~n365 & n381 ) | ( ~n365 & n2947 ) | ( n381 & n2947 ) ;
  assign n2949 = ( ~n373 & n2719 ) | ( ~n373 & n2948 ) | ( n2719 & n2948 ) ;
  assign n2950 = ( n1497 & ~n1779 ) | ( n1497 & n2949 ) | ( ~n1779 & n2949 ) ;
  assign n2951 = n442 | n463 ;
  assign n2952 = ( ~n442 & n453 ) | ( ~n442 & n2017 ) | ( n453 & n2017 ) ;
  assign n2953 = ( n2617 & n2951 ) | ( n2617 & ~n2952 ) | ( n2951 & ~n2952 ) ;
  assign n2954 = ( n1507 & ~n2951 ) | ( n1507 & n2952 ) | ( ~n2951 & n2952 ) ;
  assign n2955 = ( n2950 & ~n2953 ) | ( n2950 & n2954 ) | ( ~n2953 & n2954 ) ;
  assign n2956 = ~n549 & n1527 ;
  assign n2957 = ( ~n500 & n512 ) | ( ~n500 & n2024 ) | ( n512 & n2024 ) ;
  assign n2958 = ( ~n1805 & n2956 ) | ( ~n1805 & n2957 ) | ( n2956 & n2957 ) ;
  assign n2959 = ( n1795 & n1805 ) | ( n1795 & ~n2956 ) | ( n1805 & ~n2956 ) ;
  assign n2960 = ( n2955 & ~n2958 ) | ( n2955 & n2959 ) | ( ~n2958 & n2959 ) ;
  assign n2961 = ~n523 & n1534 ;
  assign n2962 = ( n585 & ~n1542 ) | ( n585 & n2394 ) | ( ~n1542 & n2394 ) ;
  assign n2963 = ( ~n614 & n2961 ) | ( ~n614 & n2962 ) | ( n2961 & n2962 ) ;
  assign n2964 = ( n2253 & ~n2401 ) | ( n2253 & n2963 ) | ( ~n2401 & n2963 ) ;
  assign n2965 = ( n614 & n2390 ) | ( n614 & ~n2962 ) | ( n2390 & ~n2962 ) ;
  assign n2966 = ( ~n2253 & n2401 ) | ( ~n2253 & n2965 ) | ( n2401 & n2965 ) ;
  assign n2967 = ( n2960 & n2964 ) | ( n2960 & ~n2966 ) | ( n2964 & ~n2966 ) ;
  assign n2968 = x158 & ~n743 ;
  assign n2969 = ( ~n1575 & n2257 ) | ( ~n1575 & n2744 ) | ( n2257 & n2744 ) ;
  assign n2970 = n704 | n712 ;
  assign n2971 = ( ~n2644 & n2969 ) | ( ~n2644 & n2970 ) | ( n2969 & n2970 ) ;
  assign n2972 = ~n715 & n2971 ;
  assign n2973 = n741 | n1585 ;
  assign n2974 = ( ~n741 & n742 ) | ( ~n741 & n1583 ) | ( n742 & n1583 ) ;
  assign n2975 = ( n2972 & ~n2973 ) | ( n2972 & n2974 ) | ( ~n2973 & n2974 ) ;
  assign n2976 = n2968 & ~n2975 ;
  assign n2977 = ( ~n703 & n1576 ) | ( ~n703 & n2255 ) | ( n1576 & n2255 ) ;
  assign n2978 = ( n1579 & ~n1580 ) | ( n1579 & n2977 ) | ( ~n1580 & n2977 ) ;
  assign n2979 = ( n2973 & ~n2974 ) | ( n2973 & n2978 ) | ( ~n2974 & n2978 ) ;
  assign n2980 = n2968 & n2979 ;
  assign n2981 = ( n2967 & n2976 ) | ( n2967 & n2980 ) | ( n2976 & n2980 ) ;
  assign n2982 = x33 | n1137 ;
  assign n2983 = ~n731 & n2982 ;
  assign n2984 = ( ~n770 & n786 ) | ( ~n770 & n2983 ) | ( n786 & n2983 ) ;
  assign n2985 = ( ~n778 & n2758 ) | ( ~n778 & n2984 ) | ( n2758 & n2984 ) ;
  assign n2986 = ( n1596 & ~n1857 ) | ( n1596 & n2985 ) | ( ~n1857 & n2985 ) ;
  assign n2987 = n847 | n868 ;
  assign n2988 = ( ~n847 & n858 ) | ( ~n847 & n2087 ) | ( n858 & n2087 ) ;
  assign n2989 = ( n2652 & n2987 ) | ( n2652 & ~n2988 ) | ( n2987 & ~n2988 ) ;
  assign n2990 = ( n1606 & ~n2987 ) | ( n1606 & n2988 ) | ( ~n2987 & n2988 ) ;
  assign n2991 = ( n2986 & ~n2989 ) | ( n2986 & n2990 ) | ( ~n2989 & n2990 ) ;
  assign n2992 = ~n954 & n1626 ;
  assign n2993 = ( ~n905 & n917 ) | ( ~n905 & n2094 ) | ( n917 & n2094 ) ;
  assign n2994 = ( ~n1883 & n2992 ) | ( ~n1883 & n2993 ) | ( n2992 & n2993 ) ;
  assign n2995 = ( n1873 & n1883 ) | ( n1873 & ~n2992 ) | ( n1883 & ~n2992 ) ;
  assign n2996 = ( n2991 & ~n2994 ) | ( n2991 & n2995 ) | ( ~n2994 & n2995 ) ;
  assign n2997 = ~n928 & n1633 ;
  assign n2998 = ( n990 & ~n1641 ) | ( n990 & n2438 ) | ( ~n1641 & n2438 ) ;
  assign n2999 = ( ~n1019 & n2997 ) | ( ~n1019 & n2998 ) | ( n2997 & n2998 ) ;
  assign n3000 = ( n2309 & ~n2445 ) | ( n2309 & n2999 ) | ( ~n2445 & n2999 ) ;
  assign n3001 = ( n1019 & n2434 ) | ( n1019 & ~n2998 ) | ( n2434 & ~n2998 ) ;
  assign n3002 = ( ~n2309 & n2445 ) | ( ~n2309 & n3001 ) | ( n2445 & n3001 ) ;
  assign n3003 = ( n2996 & n3000 ) | ( n2996 & ~n3002 ) | ( n3000 & ~n3002 ) ;
  assign n3004 = x159 & ~n1147 ;
  assign n3005 = ( ~n1673 & n2313 ) | ( ~n1673 & n2783 ) | ( n2313 & n2783 ) ;
  assign n3006 = n1108 | n1116 ;
  assign n3007 = ( ~n2679 & n3005 ) | ( ~n2679 & n3006 ) | ( n3005 & n3006 ) ;
  assign n3008 = ~n1119 & n3007 ;
  assign n3009 = n1145 | n1683 ;
  assign n3010 = ( ~n1145 & n1146 ) | ( ~n1145 & n1681 ) | ( n1146 & n1681 ) ;
  assign n3011 = ( n3008 & ~n3009 ) | ( n3008 & n3010 ) | ( ~n3009 & n3010 ) ;
  assign n3012 = n3004 & ~n3011 ;
  assign n3013 = ( ~n1107 & n1674 ) | ( ~n1107 & n2311 ) | ( n1674 & n2311 ) ;
  assign n3014 = ( n1677 & ~n1678 ) | ( n1677 & n3013 ) | ( ~n1678 & n3013 ) ;
  assign n3015 = ( n3009 & ~n3010 ) | ( n3009 & n3014 ) | ( ~n3010 & n3014 ) ;
  assign n3016 = n3004 & n3015 ;
  assign n3017 = ( n3003 & n3012 ) | ( n3003 & n3016 ) | ( n3012 & n3016 ) ;
  assign n3018 = x34 | n378 ;
  assign n3019 = ~n1135 & n3018 ;
  assign n3020 = ( ~n1174 & n1190 ) | ( ~n1174 & n3019 ) | ( n1190 & n3019 ) ;
  assign n3021 = ( ~n1182 & n2797 ) | ( ~n1182 & n3020 ) | ( n2797 & n3020 ) ;
  assign n3022 = ( n1694 & ~n1935 ) | ( n1694 & n3021 ) | ( ~n1935 & n3021 ) ;
  assign n3023 = n1251 | n1272 ;
  assign n3024 = ( ~n1251 & n1262 ) | ( ~n1251 & n2157 ) | ( n1262 & n2157 ) ;
  assign n3025 = ( n2687 & n3023 ) | ( n2687 & ~n3024 ) | ( n3023 & ~n3024 ) ;
  assign n3026 = ( n1704 & ~n3023 ) | ( n1704 & n3024 ) | ( ~n3023 & n3024 ) ;
  assign n3027 = ( n3022 & ~n3025 ) | ( n3022 & n3026 ) | ( ~n3025 & n3026 ) ;
  assign n3028 = ~n1358 & n1724 ;
  assign n3029 = ( ~n1309 & n1321 ) | ( ~n1309 & n2164 ) | ( n1321 & n2164 ) ;
  assign n3030 = ( ~n1961 & n3028 ) | ( ~n1961 & n3029 ) | ( n3028 & n3029 ) ;
  assign n3031 = ( n1951 & n1961 ) | ( n1951 & ~n3028 ) | ( n1961 & ~n3028 ) ;
  assign n3032 = ( n3027 & ~n3030 ) | ( n3027 & n3031 ) | ( ~n3030 & n3031 ) ;
  assign n3033 = ~n1332 & n1731 ;
  assign n3034 = ( n1394 & ~n1739 ) | ( n1394 & n2482 ) | ( ~n1739 & n2482 ) ;
  assign n3035 = ( ~n1423 & n3033 ) | ( ~n1423 & n3034 ) | ( n3033 & n3034 ) ;
  assign n3036 = ( n2365 & ~n2489 ) | ( n2365 & n3035 ) | ( ~n2489 & n3035 ) ;
  assign n3037 = ( n1423 & n2478 ) | ( n1423 & ~n3034 ) | ( n2478 & ~n3034 ) ;
  assign n3038 = ( ~n2365 & n2489 ) | ( ~n2365 & n3037 ) | ( n2489 & n3037 ) ;
  assign n3039 = ( n3032 & n3036 ) | ( n3032 & ~n3038 ) | ( n3036 & ~n3038 ) ;
  assign n3040 = x160 & ~n325 ;
  assign n3041 = n330 | n350 ;
  assign n3042 = ( ~n293 & n2369 ) | ( ~n293 & n2822 ) | ( n2369 & n2822 ) ;
  assign n3043 = n311 | n317 ;
  assign n3044 = ( ~n2714 & n3042 ) | ( ~n2714 & n3043 ) | ( n3042 & n3043 ) ;
  assign n3045 = ~n314 & n3044 ;
  assign n3046 = ( ~n330 & n341 ) | ( ~n330 & n1771 ) | ( n341 & n1771 ) ;
  assign n3047 = ( ~n3041 & n3045 ) | ( ~n3041 & n3046 ) | ( n3045 & n3046 ) ;
  assign n3048 = n3040 & ~n3047 ;
  assign n3049 = ( n294 & ~n299 ) | ( n294 & n2367 ) | ( ~n299 & n2367 ) ;
  assign n3050 = ( ~n319 & n1765 ) | ( ~n319 & n3049 ) | ( n1765 & n3049 ) ;
  assign n3051 = ( n3041 & ~n3046 ) | ( n3041 & n3050 ) | ( ~n3046 & n3050 ) ;
  assign n3052 = n3040 & n3051 ;
  assign n3053 = ( n3039 & n3048 ) | ( n3039 & n3052 ) | ( n3048 & n3052 ) ;
  assign n3054 = x35 | n783 ;
  assign n3055 = ~n364 & n3054 ;
  assign n3056 = ( ~n372 & n382 ) | ( ~n372 & n3055 ) | ( n382 & n3055 ) ;
  assign n3057 = ( ~n359 & n377 ) | ( ~n359 & n3056 ) | ( n377 & n3056 ) ;
  assign n3058 = ( ~n410 & n1781 ) | ( ~n410 & n3057 ) | ( n1781 & n3057 ) ;
  assign n3059 = n433 | n1515 ;
  assign n3060 = ( ~n433 & n437 ) | ( ~n433 & n454 ) | ( n437 & n454 ) ;
  assign n3061 = ( n2725 & n3059 ) | ( n2725 & ~n3060 ) | ( n3059 & ~n3060 ) ;
  assign n3062 = ( n1790 & ~n3059 ) | ( n1790 & n3060 ) | ( ~n3059 & n3060 ) ;
  assign n3063 = ( n3058 & ~n3061 ) | ( n3058 & n3062 ) | ( ~n3061 & n3062 ) ;
  assign n3064 = ~n553 & n1808 ;
  assign n3065 = ( n2022 & n2035 ) | ( n2022 & ~n3064 ) | ( n2035 & ~n3064 ) ;
  assign n3066 = ( ~n484 & n513 ) | ( ~n484 & n2222 ) | ( n513 & n2222 ) ;
  assign n3067 = ( ~n2035 & n3064 ) | ( ~n2035 & n3066 ) | ( n3064 & n3066 ) ;
  assign n3068 = ( n3063 & n3065 ) | ( n3063 & ~n3067 ) | ( n3065 & ~n3067 ) ;
  assign n3069 = ~n600 & n1813 ;
  assign n3070 = ( n630 & ~n1545 ) | ( n630 & n3069 ) | ( ~n1545 & n3069 ) ;
  assign n3071 = ( n2409 & ~n2527 ) | ( n2409 & n3070 ) | ( ~n2527 & n3070 ) ;
  assign n3072 = ( ~n630 & n1545 ) | ( ~n630 & n2522 ) | ( n1545 & n2522 ) ;
  assign n3073 = ( ~n2409 & n2527 ) | ( ~n2409 & n3072 ) | ( n2527 & n3072 ) ;
  assign n3074 = ( n3068 & n3071 ) | ( n3068 & ~n3073 ) | ( n3071 & ~n3073 ) ;
  assign n3075 = x161 & ~n730 ;
  assign n3076 = n735 | n755 ;
  assign n3077 = ( ~n698 & n2413 ) | ( ~n698 & n2859 ) | ( n2413 & n2859 ) ;
  assign n3078 = ~n722 & n1579 ;
  assign n3079 = n716 | n722 ;
  assign n3080 = ( n3077 & ~n3078 ) | ( n3077 & n3079 ) | ( ~n3078 & n3079 ) ;
  assign n3081 = ~n719 & n3080 ;
  assign n3082 = ( ~n735 & n746 ) | ( ~n735 & n1849 ) | ( n746 & n1849 ) ;
  assign n3083 = ( ~n3076 & n3081 ) | ( ~n3076 & n3082 ) | ( n3081 & n3082 ) ;
  assign n3084 = n3075 & ~n3083 ;
  assign n3085 = ( n699 & ~n704 ) | ( n699 & n2411 ) | ( ~n704 & n2411 ) ;
  assign n3086 = ( ~n724 & n1843 ) | ( ~n724 & n3085 ) | ( n1843 & n3085 ) ;
  assign n3087 = ( n3076 & ~n3082 ) | ( n3076 & n3086 ) | ( ~n3082 & n3086 ) ;
  assign n3088 = n3075 & n3087 ;
  assign n3089 = ( n3074 & n3084 ) | ( n3074 & n3088 ) | ( n3084 & n3088 ) ;
  assign n3090 = x36 | n1187 ;
  assign n3091 = ~n769 & n3090 ;
  assign n3092 = ( ~n777 & n787 ) | ( ~n777 & n3091 ) | ( n787 & n3091 ) ;
  assign n3093 = ( ~n764 & n782 ) | ( ~n764 & n3092 ) | ( n782 & n3092 ) ;
  assign n3094 = ( ~n815 & n1859 ) | ( ~n815 & n3093 ) | ( n1859 & n3093 ) ;
  assign n3095 = n838 | n1614 ;
  assign n3096 = ( ~n838 & n842 ) | ( ~n838 & n859 ) | ( n842 & n859 ) ;
  assign n3097 = ( n2764 & n3095 ) | ( n2764 & ~n3096 ) | ( n3095 & ~n3096 ) ;
  assign n3098 = ( n1868 & ~n3095 ) | ( n1868 & n3096 ) | ( ~n3095 & n3096 ) ;
  assign n3099 = ( n3094 & ~n3097 ) | ( n3094 & n3098 ) | ( ~n3097 & n3098 ) ;
  assign n3100 = ~n958 & n1886 ;
  assign n3101 = ( n2092 & n2105 ) | ( n2092 & ~n3100 ) | ( n2105 & ~n3100 ) ;
  assign n3102 = ( ~n889 & n918 ) | ( ~n889 & n2278 ) | ( n918 & n2278 ) ;
  assign n3103 = ( ~n2105 & n3100 ) | ( ~n2105 & n3102 ) | ( n3100 & n3102 ) ;
  assign n3104 = ( n3099 & n3101 ) | ( n3099 & ~n3103 ) | ( n3101 & ~n3103 ) ;
  assign n3105 = ~n1005 & n1891 ;
  assign n3106 = ( n1035 & ~n1644 ) | ( n1035 & n3105 ) | ( ~n1644 & n3105 ) ;
  assign n3107 = ( n2453 & ~n2564 ) | ( n2453 & n3106 ) | ( ~n2564 & n3106 ) ;
  assign n3108 = ( ~n1035 & n1644 ) | ( ~n1035 & n2559 ) | ( n1644 & n2559 ) ;
  assign n3109 = ( ~n2453 & n2564 ) | ( ~n2453 & n3108 ) | ( n2564 & n3108 ) ;
  assign n3110 = ( n3104 & n3107 ) | ( n3104 & ~n3109 ) | ( n3107 & ~n3109 ) ;
  assign n3111 = x162 & ~n1134 ;
  assign n3112 = n1139 | n1159 ;
  assign n3113 = ( ~n1102 & n2457 ) | ( ~n1102 & n2896 ) | ( n2457 & n2896 ) ;
  assign n3114 = ~n1126 & n1677 ;
  assign n3115 = n1120 | n1126 ;
  assign n3116 = ( n3113 & ~n3114 ) | ( n3113 & n3115 ) | ( ~n3114 & n3115 ) ;
  assign n3117 = ~n1123 & n3116 ;
  assign n3118 = ( ~n1139 & n1150 ) | ( ~n1139 & n1927 ) | ( n1150 & n1927 ) ;
  assign n3119 = ( ~n3112 & n3117 ) | ( ~n3112 & n3118 ) | ( n3117 & n3118 ) ;
  assign n3120 = n3111 & ~n3119 ;
  assign n3121 = ( n1103 & ~n1108 ) | ( n1103 & n2455 ) | ( ~n1108 & n2455 ) ;
  assign n3122 = ( ~n1128 & n1921 ) | ( ~n1128 & n3121 ) | ( n1921 & n3121 ) ;
  assign n3123 = ( n3112 & ~n3118 ) | ( n3112 & n3122 ) | ( ~n3118 & n3122 ) ;
  assign n3124 = n3111 & n3123 ;
  assign n3125 = ( n3110 & n3120 ) | ( n3110 & n3124 ) | ( n3120 & n3124 ) ;
  assign n3126 = x37 | n366 ;
  assign n3127 = ~n1173 & n3126 ;
  assign n3128 = ( ~n1181 & n1191 ) | ( ~n1181 & n3127 ) | ( n1191 & n3127 ) ;
  assign n3129 = ( ~n1168 & n1186 ) | ( ~n1168 & n3128 ) | ( n1186 & n3128 ) ;
  assign n3130 = ( ~n1219 & n1937 ) | ( ~n1219 & n3129 ) | ( n1937 & n3129 ) ;
  assign n3131 = n1242 | n1712 ;
  assign n3132 = ( ~n1242 & n1246 ) | ( ~n1242 & n1263 ) | ( n1246 & n1263 ) ;
  assign n3133 = ( n2803 & n3131 ) | ( n2803 & ~n3132 ) | ( n3131 & ~n3132 ) ;
  assign n3134 = ( n1946 & ~n3131 ) | ( n1946 & n3132 ) | ( ~n3131 & n3132 ) ;
  assign n3135 = ( n3130 & ~n3133 ) | ( n3130 & n3134 ) | ( ~n3133 & n3134 ) ;
  assign n3136 = ~n1362 & n1964 ;
  assign n3137 = ( n2162 & n2175 ) | ( n2162 & ~n3136 ) | ( n2175 & ~n3136 ) ;
  assign n3138 = ( ~n1293 & n1322 ) | ( ~n1293 & n2334 ) | ( n1322 & n2334 ) ;
  assign n3139 = ( ~n2175 & n3136 ) | ( ~n2175 & n3138 ) | ( n3136 & n3138 ) ;
  assign n3140 = ( n3135 & n3137 ) | ( n3135 & ~n3139 ) | ( n3137 & ~n3139 ) ;
  assign n3141 = ~n1409 & n1969 ;
  assign n3142 = ( n1439 & ~n1742 ) | ( n1439 & n3141 ) | ( ~n1742 & n3141 ) ;
  assign n3143 = ( n2497 & ~n2601 ) | ( n2497 & n3142 ) | ( ~n2601 & n3142 ) ;
  assign n3144 = ( ~n1439 & n1742 ) | ( ~n1439 & n2596 ) | ( n1742 & n2596 ) ;
  assign n3145 = ( ~n2497 & n2601 ) | ( ~n2497 & n3144 ) | ( n2601 & n3144 ) ;
  assign n3146 = ( n3140 & n3143 ) | ( n3140 & ~n3145 ) | ( n3143 & ~n3145 ) ;
  assign n3147 = x163 & ~n363 ;
  assign n3148 = n380 | n1491 ;
  assign n3149 = ( ~n1479 & n2501 ) | ( ~n1479 & n2933 ) | ( n2501 & n2933 ) ;
  assign n3150 = ~n304 & n1765 ;
  assign n3151 = n304 | n318 ;
  assign n3152 = ( n3149 & ~n3150 ) | ( n3149 & n3151 ) | ( ~n3150 & n3151 ) ;
  assign n3153 = ~n347 & n3152 ;
  assign n3154 = ( n342 & ~n380 ) | ( n342 & n1488 ) | ( ~n380 & n1488 ) ;
  assign n3155 = ( ~n3148 & n3153 ) | ( ~n3148 & n3154 ) | ( n3153 & n3154 ) ;
  assign n3156 = n3147 & ~n3155 ;
  assign n3157 = ( ~n311 & n1480 ) | ( ~n311 & n2499 ) | ( n1480 & n2499 ) ;
  assign n3158 = ( ~n1484 & n1998 ) | ( ~n1484 & n3157 ) | ( n1998 & n3157 ) ;
  assign n3159 = ( n3148 & ~n3154 ) | ( n3148 & n3158 ) | ( ~n3154 & n3158 ) ;
  assign n3160 = n3147 & n3159 ;
  assign n3161 = ( n3146 & n3156 ) | ( n3146 & n3160 ) | ( n3156 & n3160 ) ;
  assign n3162 = x38 | n771 ;
  assign n3163 = ~n371 & n3162 ;
  assign n3164 = ( ~n358 & n376 ) | ( ~n358 & n3163 ) | ( n376 & n3163 ) ;
  assign n3165 = ( ~n402 & n1497 ) | ( ~n402 & n3164 ) | ( n1497 & n3164 ) ;
  assign n3166 = ( ~n1502 & n2008 ) | ( ~n1502 & n3165 ) | ( n2008 & n3165 ) ;
  assign n3167 = n427 | n1797 ;
  assign n3168 = ( ~n427 & n457 ) | ( ~n427 & n1512 ) | ( n457 & n1512 ) ;
  assign n3169 = ( n2840 & n3167 ) | ( n2840 & ~n3168 ) | ( n3167 & ~n3168 ) ;
  assign n3170 = ( n2017 & ~n3167 ) | ( n2017 & n3168 ) | ( ~n3167 & n3168 ) ;
  assign n3171 = ( n3166 & ~n3169 ) | ( n3166 & n3170 ) | ( ~n3169 & n3170 ) ;
  assign n3172 = ~n537 & n2030 ;
  assign n3173 = ( ~n478 & n487 ) | ( ~n478 & n514 ) | ( n487 & n514 ) ;
  assign n3174 = ( ~n2231 & n3172 ) | ( ~n2231 & n3173 ) | ( n3172 & n3173 ) ;
  assign n3175 = ( n503 & n2231 ) | ( n503 & ~n3172 ) | ( n2231 & ~n3172 ) ;
  assign n3176 = ( n3171 & ~n3174 ) | ( n3171 & n3175 ) | ( ~n3174 & n3175 ) ;
  assign n3177 = ~n610 & n2040 ;
  assign n3178 = ( n1555 & ~n1823 ) | ( n1555 & n3177 ) | ( ~n1823 & n3177 ) ;
  assign n3179 = ( n2534 & ~n2636 ) | ( n2534 & n3178 ) | ( ~n2636 & n3178 ) ;
  assign n3180 = ( ~n1555 & n1823 ) | ( ~n1555 & n2631 ) | ( n1823 & n2631 ) ;
  assign n3181 = ( ~n2534 & n2636 ) | ( ~n2534 & n3180 ) | ( n2636 & n3180 ) ;
  assign n3182 = ( n3176 & n3179 ) | ( n3176 & ~n3181 ) | ( n3179 & ~n3181 ) ;
  assign n3183 = x164 & ~n768 ;
  assign n3184 = n785 | n1590 ;
  assign n3185 = ( ~n1578 & n2538 ) | ( ~n1578 & n2970 ) | ( n2538 & n2970 ) ;
  assign n3186 = ~n709 & n1843 ;
  assign n3187 = n709 | n723 ;
  assign n3188 = ( n3185 & ~n3186 ) | ( n3185 & n3187 ) | ( ~n3186 & n3187 ) ;
  assign n3189 = ~n752 & n3188 ;
  assign n3190 = ( n747 & ~n785 ) | ( n747 & n1587 ) | ( ~n785 & n1587 ) ;
  assign n3191 = ( ~n3184 & n3189 ) | ( ~n3184 & n3190 ) | ( n3189 & n3190 ) ;
  assign n3192 = n3183 & ~n3191 ;
  assign n3193 = ( ~n716 & n1579 ) | ( ~n716 & n2536 ) | ( n1579 & n2536 ) ;
  assign n3194 = ( ~n1583 & n2068 ) | ( ~n1583 & n3193 ) | ( n2068 & n3193 ) ;
  assign n3195 = ( n3184 & ~n3190 ) | ( n3184 & n3194 ) | ( ~n3190 & n3194 ) ;
  assign n3196 = n3183 & n3195 ;
  assign n3197 = ( n3182 & n3192 ) | ( n3182 & n3196 ) | ( n3192 & n3196 ) ;
  assign n3198 = x39 | n1175 ;
  assign n3199 = ~n776 & n3198 ;
  assign n3200 = ( ~n763 & n781 ) | ( ~n763 & n3199 ) | ( n781 & n3199 ) ;
  assign n3201 = ( ~n807 & n1596 ) | ( ~n807 & n3200 ) | ( n1596 & n3200 ) ;
  assign n3202 = ( ~n1601 & n2078 ) | ( ~n1601 & n3201 ) | ( n2078 & n3201 ) ;
  assign n3203 = n832 | n1875 ;
  assign n3204 = ( ~n832 & n862 ) | ( ~n832 & n1611 ) | ( n862 & n1611 ) ;
  assign n3205 = ( n2877 & n3203 ) | ( n2877 & ~n3204 ) | ( n3203 & ~n3204 ) ;
  assign n3206 = ( n2087 & ~n3203 ) | ( n2087 & n3204 ) | ( ~n3203 & n3204 ) ;
  assign n3207 = ( n3202 & ~n3205 ) | ( n3202 & n3206 ) | ( ~n3205 & n3206 ) ;
  assign n3208 = ~n942 & n2100 ;
  assign n3209 = ( ~n883 & n892 ) | ( ~n883 & n919 ) | ( n892 & n919 ) ;
  assign n3210 = ( ~n2287 & n3208 ) | ( ~n2287 & n3209 ) | ( n3208 & n3209 ) ;
  assign n3211 = ( n908 & n2287 ) | ( n908 & ~n3208 ) | ( n2287 & ~n3208 ) ;
  assign n3212 = ( n3207 & ~n3210 ) | ( n3207 & n3211 ) | ( ~n3210 & n3211 ) ;
  assign n3213 = ~n1015 & n2110 ;
  assign n3214 = ( n1654 & ~n1901 ) | ( n1654 & n3213 ) | ( ~n1901 & n3213 ) ;
  assign n3215 = ( n2571 & ~n2671 ) | ( n2571 & n3214 ) | ( ~n2671 & n3214 ) ;
  assign n3216 = ( ~n1654 & n1901 ) | ( ~n1654 & n2666 ) | ( n1901 & n2666 ) ;
  assign n3217 = ( ~n2571 & n2671 ) | ( ~n2571 & n3216 ) | ( n2671 & n3216 ) ;
  assign n3218 = ( n3212 & n3215 ) | ( n3212 & ~n3217 ) | ( n3215 & ~n3217 ) ;
  assign n3219 = x165 & ~n1172 ;
  assign n3220 = n1189 | n1688 ;
  assign n3221 = ( ~n1676 & n2575 ) | ( ~n1676 & n3006 ) | ( n2575 & n3006 ) ;
  assign n3222 = ~n1113 & n1921 ;
  assign n3223 = n1113 | n1127 ;
  assign n3224 = ( n3221 & ~n3222 ) | ( n3221 & n3223 ) | ( ~n3222 & n3223 ) ;
  assign n3225 = ~n1156 & n3224 ;
  assign n3226 = ( n1151 & ~n1189 ) | ( n1151 & n1685 ) | ( ~n1189 & n1685 ) ;
  assign n3227 = ( ~n3220 & n3225 ) | ( ~n3220 & n3226 ) | ( n3225 & n3226 ) ;
  assign n3228 = n3219 & ~n3227 ;
  assign n3229 = ( ~n1120 & n1677 ) | ( ~n1120 & n2573 ) | ( n1677 & n2573 ) ;
  assign n3230 = ( ~n1681 & n2138 ) | ( ~n1681 & n3229 ) | ( n2138 & n3229 ) ;
  assign n3231 = ( n3220 & ~n3226 ) | ( n3220 & n3230 ) | ( ~n3226 & n3230 ) ;
  assign n3232 = n3219 & n3231 ;
  assign n3233 = ( n3218 & n3228 ) | ( n3218 & n3232 ) | ( n3228 & n3232 ) ;
  assign n3234 = x40 | n360 ;
  assign n3235 = ~n1180 & n3234 ;
  assign n3236 = ( ~n1167 & n1185 ) | ( ~n1167 & n3235 ) | ( n1185 & n3235 ) ;
  assign n3237 = ( ~n1211 & n1694 ) | ( ~n1211 & n3236 ) | ( n1694 & n3236 ) ;
  assign n3238 = ( ~n1699 & n2148 ) | ( ~n1699 & n3237 ) | ( n2148 & n3237 ) ;
  assign n3239 = n1236 | n1953 ;
  assign n3240 = ( ~n1236 & n1266 ) | ( ~n1236 & n1709 ) | ( n1266 & n1709 ) ;
  assign n3241 = ( n2914 & n3239 ) | ( n2914 & ~n3240 ) | ( n3239 & ~n3240 ) ;
  assign n3242 = ( n2157 & ~n3239 ) | ( n2157 & n3240 ) | ( ~n3239 & n3240 ) ;
  assign n3243 = ( n3238 & ~n3241 ) | ( n3238 & n3242 ) | ( ~n3241 & n3242 ) ;
  assign n3244 = ~n1346 & n2170 ;
  assign n3245 = ( ~n1287 & n1296 ) | ( ~n1287 & n1323 ) | ( n1296 & n1323 ) ;
  assign n3246 = ( ~n2343 & n3244 ) | ( ~n2343 & n3245 ) | ( n3244 & n3245 ) ;
  assign n3247 = ( n1312 & n2343 ) | ( n1312 & ~n3244 ) | ( n2343 & ~n3244 ) ;
  assign n3248 = ( n3243 & ~n3246 ) | ( n3243 & n3247 ) | ( ~n3246 & n3247 ) ;
  assign n3249 = ~n1419 & n2180 ;
  assign n3250 = ( n1752 & ~n1979 ) | ( n1752 & n3249 ) | ( ~n1979 & n3249 ) ;
  assign n3251 = ( n2607 & ~n2706 ) | ( n2607 & n3250 ) | ( ~n2706 & n3250 ) ;
  assign n3252 = ( ~n1752 & n1979 ) | ( ~n1752 & n2701 ) | ( n1979 & n2701 ) ;
  assign n3253 = ( ~n2607 & n2706 ) | ( ~n2607 & n3252 ) | ( n2706 & n3252 ) ;
  assign n3254 = ( n3248 & n3251 ) | ( n3248 & ~n3253 ) | ( n3251 & ~n3253 ) ;
  assign n3255 = x166 & ~n370 ;
  assign n3256 = n368 | n1776 ;
  assign n3257 = ( n300 & ~n321 ) | ( n300 & n3043 ) | ( ~n321 & n3043 ) ;
  assign n3258 = ~n333 & n1998 ;
  assign n3259 = n333 | n1483 ;
  assign n3260 = ( n3257 & ~n3258 ) | ( n3257 & n3259 ) | ( ~n3258 & n3259 ) ;
  assign n3261 = ~n336 & n3260 ;
  assign n3262 = ( ~n368 & n369 ) | ( ~n368 & n1489 ) | ( n369 & n1489 ) ;
  assign n3263 = ( ~n3256 & n3261 ) | ( ~n3256 & n3262 ) | ( n3261 & n3262 ) ;
  assign n3264 = n3255 & ~n3263 ;
  assign n3265 = ( ~n318 & n1765 ) | ( ~n318 & n2609 ) | ( n1765 & n2609 ) ;
  assign n3266 = ( ~n1771 & n2209 ) | ( ~n1771 & n3265 ) | ( n2209 & n3265 ) ;
  assign n3267 = ( n3256 & ~n3262 ) | ( n3256 & n3266 ) | ( ~n3262 & n3266 ) ;
  assign n3268 = n3255 & n3267 ;
  assign n3269 = ( n3254 & n3264 ) | ( n3254 & n3268 ) | ( n3264 & n3268 ) ;
  assign n3270 = x41 | n765 ;
  assign n3271 = ~n357 & n3270 ;
  assign n3272 = ( ~n398 & n1496 ) | ( ~n398 & n3271 ) | ( n1496 & n3271 ) ;
  assign n3273 = ( ~n409 & n1781 ) | ( ~n409 & n3272 ) | ( n1781 & n3272 ) ;
  assign n3274 = ( n418 & ~n1785 ) | ( n418 & n3273 ) | ( ~n1785 & n3273 ) ;
  assign n3275 = n493 | n2024 ;
  assign n3276 = ( ~n493 & n497 ) | ( ~n493 & n1794 ) | ( n497 & n1794 ) ;
  assign n3277 = ( n2951 & n3275 ) | ( n2951 & ~n3276 ) | ( n3275 & ~n3276 ) ;
  assign n3278 = ( n454 & ~n3275 ) | ( n454 & n3276 ) | ( ~n3275 & n3276 ) ;
  assign n3279 = ( n3274 & ~n3277 ) | ( n3274 & n3278 ) | ( ~n3277 & n3278 ) ;
  assign n3280 = ~n531 & n2227 ;
  assign n3281 = ( ~n474 & n507 ) | ( ~n474 & n1526 ) | ( n507 & n1526 ) ;
  assign n3282 = ( ~n556 & n3280 ) | ( ~n556 & n3281 ) | ( n3280 & n3281 ) ;
  assign n3283 = ( n556 & n1522 ) | ( n556 & ~n3280 ) | ( n1522 & ~n3280 ) ;
  assign n3284 = ( n3279 & ~n3282 ) | ( n3279 & n3283 ) | ( ~n3282 & n3283 ) ;
  assign n3285 = ( ~n686 & n687 ) | ( ~n686 & n2745 ) | ( n687 & n2745 ) ;
  assign n3286 = ~n591 & n2235 ;
  assign n3287 = ( n645 & n1830 ) | ( n645 & ~n2242 ) | ( n1830 & ~n2242 ) ;
  assign n3288 = ( n641 & ~n645 ) | ( n641 & n2049 ) | ( ~n645 & n2049 ) ;
  assign n3289 = ( n3286 & n3287 ) | ( n3286 & ~n3288 ) | ( n3287 & ~n3288 ) ;
  assign n3290 = ( n2642 & ~n3285 ) | ( n2642 & n3289 ) | ( ~n3285 & n3289 ) ;
  assign n3291 = ( n2737 & ~n3287 ) | ( n2737 & n3288 ) | ( ~n3287 & n3288 ) ;
  assign n3292 = ( ~n2642 & n3285 ) | ( ~n2642 & n3291 ) | ( n3285 & n3291 ) ;
  assign n3293 = ( n3284 & n3290 ) | ( n3284 & ~n3292 ) | ( n3290 & ~n3292 ) ;
  assign n3294 = x167 & ~n775 ;
  assign n3295 = n773 | n1854 ;
  assign n3296 = ( n705 & ~n726 ) | ( n705 & n3079 ) | ( ~n726 & n3079 ) ;
  assign n3297 = ~n738 & n2068 ;
  assign n3298 = n738 | n1582 ;
  assign n3299 = ( n3296 & ~n3297 ) | ( n3296 & n3298 ) | ( ~n3297 & n3298 ) ;
  assign n3300 = ~n741 & n3299 ;
  assign n3301 = ( ~n773 & n774 ) | ( ~n773 & n1588 ) | ( n774 & n1588 ) ;
  assign n3302 = ( ~n3295 & n3300 ) | ( ~n3295 & n3301 ) | ( n3300 & n3301 ) ;
  assign n3303 = n3294 & ~n3302 ;
  assign n3304 = ( ~n723 & n1843 ) | ( ~n723 & n2644 ) | ( n1843 & n2644 ) ;
  assign n3305 = ( ~n1849 & n2265 ) | ( ~n1849 & n3304 ) | ( n2265 & n3304 ) ;
  assign n3306 = ( n3295 & ~n3301 ) | ( n3295 & n3305 ) | ( ~n3301 & n3305 ) ;
  assign n3307 = n3294 & n3306 ;
  assign n3308 = ( n3293 & n3303 ) | ( n3293 & n3307 ) | ( n3303 & n3307 ) ;
  assign n3309 = x42 | n1169 ;
  assign n3310 = ~n762 & n3309 ;
  assign n3311 = ( ~n803 & n1595 ) | ( ~n803 & n3310 ) | ( n1595 & n3310 ) ;
  assign n3312 = ( ~n814 & n1859 ) | ( ~n814 & n3311 ) | ( n1859 & n3311 ) ;
  assign n3313 = ( n823 & ~n1863 ) | ( n823 & n3312 ) | ( ~n1863 & n3312 ) ;
  assign n3314 = n898 | n2094 ;
  assign n3315 = ( ~n898 & n902 ) | ( ~n898 & n1872 ) | ( n902 & n1872 ) ;
  assign n3316 = ( n2987 & n3314 ) | ( n2987 & ~n3315 ) | ( n3314 & ~n3315 ) ;
  assign n3317 = ( n859 & ~n3314 ) | ( n859 & n3315 ) | ( ~n3314 & n3315 ) ;
  assign n3318 = ( n3313 & ~n3316 ) | ( n3313 & n3317 ) | ( ~n3316 & n3317 ) ;
  assign n3319 = ~n936 & n2283 ;
  assign n3320 = ( ~n879 & n912 ) | ( ~n879 & n1625 ) | ( n912 & n1625 ) ;
  assign n3321 = ( ~n961 & n3319 ) | ( ~n961 & n3320 ) | ( n3319 & n3320 ) ;
  assign n3322 = ( n961 & n1621 ) | ( n961 & ~n3319 ) | ( n1621 & ~n3319 ) ;
  assign n3323 = ( n3318 & ~n3321 ) | ( n3318 & n3322 ) | ( ~n3321 & n3322 ) ;
  assign n3324 = ( ~n1090 & n1091 ) | ( ~n1090 & n2784 ) | ( n1091 & n2784 ) ;
  assign n3325 = ~n996 & n2291 ;
  assign n3326 = ( n1050 & n1908 ) | ( n1050 & ~n2298 ) | ( n1908 & ~n2298 ) ;
  assign n3327 = ( n1046 & ~n1050 ) | ( n1046 & n2119 ) | ( ~n1050 & n2119 ) ;
  assign n3328 = ( n3325 & n3326 ) | ( n3325 & ~n3327 ) | ( n3326 & ~n3327 ) ;
  assign n3329 = ( n2677 & ~n3324 ) | ( n2677 & n3328 ) | ( ~n3324 & n3328 ) ;
  assign n3330 = ( n2776 & ~n3326 ) | ( n2776 & n3327 ) | ( ~n3326 & n3327 ) ;
  assign n3331 = ( ~n2677 & n3324 ) | ( ~n2677 & n3330 ) | ( n3324 & n3330 ) ;
  assign n3332 = ( n3323 & n3329 ) | ( n3323 & ~n3331 ) | ( n3329 & ~n3331 ) ;
  assign n3333 = x168 & ~n1179 ;
  assign n3334 = n1177 | n1932 ;
  assign n3335 = ( n1109 & ~n1130 ) | ( n1109 & n3115 ) | ( ~n1130 & n3115 ) ;
  assign n3336 = ~n1142 & n2138 ;
  assign n3337 = n1142 | n1680 ;
  assign n3338 = ( n3335 & ~n3336 ) | ( n3335 & n3337 ) | ( ~n3336 & n3337 ) ;
  assign n3339 = ~n1145 & n3338 ;
  assign n3340 = ( ~n1177 & n1178 ) | ( ~n1177 & n1686 ) | ( n1178 & n1686 ) ;
  assign n3341 = ( ~n3334 & n3339 ) | ( ~n3334 & n3340 ) | ( n3339 & n3340 ) ;
  assign n3342 = n3333 & ~n3341 ;
  assign n3343 = ( ~n1127 & n1921 ) | ( ~n1127 & n2679 ) | ( n1921 & n2679 ) ;
  assign n3344 = ( ~n1927 & n2321 ) | ( ~n1927 & n3343 ) | ( n2321 & n3343 ) ;
  assign n3345 = ( n3334 & ~n3340 ) | ( n3334 & n3344 ) | ( ~n3340 & n3344 ) ;
  assign n3346 = n3333 & n3345 ;
  assign n3347 = ( n3332 & n3342 ) | ( n3332 & n3346 ) | ( n3342 & n3346 ) ;
  assign n3348 = x43 | n353 ;
  assign n3349 = ~n1166 & n3348 ;
  assign n3350 = ( ~n1207 & n1693 ) | ( ~n1207 & n3349 ) | ( n1693 & n3349 ) ;
  assign n3351 = ( ~n1218 & n1937 ) | ( ~n1218 & n3350 ) | ( n1937 & n3350 ) ;
  assign n3352 = ( n1227 & ~n1941 ) | ( n1227 & n3351 ) | ( ~n1941 & n3351 ) ;
  assign n3353 = n1302 | n2164 ;
  assign n3354 = ( ~n1302 & n1306 ) | ( ~n1302 & n1950 ) | ( n1306 & n1950 ) ;
  assign n3355 = ( n3023 & n3353 ) | ( n3023 & ~n3354 ) | ( n3353 & ~n3354 ) ;
  assign n3356 = ( n1263 & ~n3353 ) | ( n1263 & n3354 ) | ( ~n3353 & n3354 ) ;
  assign n3357 = ( n3352 & ~n3355 ) | ( n3352 & n3356 ) | ( ~n3355 & n3356 ) ;
  assign n3358 = ~n1340 & n2339 ;
  assign n3359 = ( ~n1283 & n1316 ) | ( ~n1283 & n1723 ) | ( n1316 & n1723 ) ;
  assign n3360 = ( ~n1365 & n3358 ) | ( ~n1365 & n3359 ) | ( n3358 & n3359 ) ;
  assign n3361 = ( n1365 & n1719 ) | ( n1365 & ~n3358 ) | ( n1719 & ~n3358 ) ;
  assign n3362 = ( n3357 & ~n3360 ) | ( n3357 & n3361 ) | ( ~n3360 & n3361 ) ;
  assign n3363 = ( n298 & ~n1477 ) | ( n298 & n2823 ) | ( ~n1477 & n2823 ) ;
  assign n3364 = ~n1400 & n2347 ;
  assign n3365 = ( n1454 & n1986 ) | ( n1454 & ~n2354 ) | ( n1986 & ~n2354 ) ;
  assign n3366 = ( n1450 & ~n1454 ) | ( n1450 & n2189 ) | ( ~n1454 & n2189 ) ;
  assign n3367 = ( n3364 & n3365 ) | ( n3364 & ~n3366 ) | ( n3365 & ~n3366 ) ;
  assign n3368 = ( n2712 & ~n3363 ) | ( n2712 & n3367 ) | ( ~n3363 & n3367 ) ;
  assign n3369 = ( n2815 & ~n3365 ) | ( n2815 & n3366 ) | ( ~n3365 & n3366 ) ;
  assign n3370 = ( ~n2712 & n3363 ) | ( ~n2712 & n3369 ) | ( n3363 & n3369 ) ;
  assign n3371 = ( n3362 & n3368 ) | ( n3362 & ~n3370 ) | ( n3368 & ~n3370 ) ;
  assign n3372 = x169 & ~n356 ;
  assign n3373 = n362 | n383 ;
  assign n3374 = ( ~n322 & n1481 ) | ( ~n322 & n3151 ) | ( n1481 & n3151 ) ;
  assign n3375 = ~n340 & n2209 ;
  assign n3376 = n337 | n340 ;
  assign n3377 = ( n3374 & ~n3375 ) | ( n3374 & n3376 ) | ( ~n3375 & n3376 ) ;
  assign n3378 = ~n330 & n3377 ;
  assign n3379 = ( ~n362 & n373 ) | ( ~n362 & n1774 ) | ( n373 & n1774 ) ;
  assign n3380 = ( ~n3373 & n3378 ) | ( ~n3373 & n3379 ) | ( n3378 & n3379 ) ;
  assign n3381 = n3372 & ~n3380 ;
  assign n3382 = ( ~n1483 & n1998 ) | ( ~n1483 & n2714 ) | ( n1998 & n2714 ) ;
  assign n3383 = ( ~n342 & n2377 ) | ( ~n342 & n3382 ) | ( n2377 & n3382 ) ;
  assign n3384 = ( n3373 & ~n3379 ) | ( n3373 & n3383 ) | ( ~n3379 & n3383 ) ;
  assign n3385 = n3372 & n3384 ;
  assign n3386 = ( n3371 & n3381 ) | ( n3371 & n3385 ) | ( n3381 & n3385 ) ;
  assign n3387 = x44 | n758 ;
  assign n3388 = ~n397 & n3387 ;
  assign n3389 = ( ~n408 & n420 ) | ( ~n408 & n3388 ) | ( n420 & n3388 ) ;
  assign n3390 = ( ~n414 & n2008 ) | ( ~n414 & n3389 ) | ( n2008 & n3389 ) ;
  assign n3391 = ( n1506 & ~n2012 ) | ( n1506 & n3390 ) | ( ~n2012 & n3390 ) ;
  assign n3392 = n490 | n2222 ;
  assign n3393 = ( ~n490 & n501 ) | ( ~n490 & n2021 ) | ( n501 & n2021 ) ;
  assign n3394 = ( n3059 & n3392 ) | ( n3059 & ~n3393 ) | ( n3392 & ~n3393 ) ;
  assign n3395 = ( n1512 & ~n3392 ) | ( n1512 & n3393 ) | ( ~n3392 & n3393 ) ;
  assign n3396 = ( n3391 & ~n3394 ) | ( n3391 & n3395 ) | ( ~n3394 & n3395 ) ;
  assign n3397 = ~n526 & n570 ;
  assign n3398 = ( ~n549 & n1523 ) | ( ~n549 & n1807 ) | ( n1523 & n1807 ) ;
  assign n3399 = ( ~n1534 & n3397 ) | ( ~n1534 & n3398 ) | ( n3397 & n3398 ) ;
  assign n3400 = ( n1534 & n1805 ) | ( n1534 & ~n3397 ) | ( n1805 & ~n3397 ) ;
  assign n3401 = ( n3396 & ~n3399 ) | ( n3396 & n3400 ) | ( ~n3399 & n3400 ) ;
  assign n3402 = ( n703 & ~n1576 ) | ( n703 & n2860 ) | ( ~n1576 & n2860 ) ;
  assign n3403 = ~n588 & n2394 ;
  assign n3404 = ( n649 & n2056 ) | ( n649 & ~n2398 ) | ( n2056 & ~n2398 ) ;
  assign n3405 = ( n638 & ~n649 ) | ( n638 & n2244 ) | ( ~n649 & n2244 ) ;
  assign n3406 = ( n3403 & n3404 ) | ( n3403 & ~n3405 ) | ( n3404 & ~n3405 ) ;
  assign n3407 = ( n2754 & ~n3402 ) | ( n2754 & n3406 ) | ( ~n3402 & n3406 ) ;
  assign n3408 = ( n2852 & ~n3404 ) | ( n2852 & n3405 ) | ( ~n3404 & n3405 ) ;
  assign n3409 = ( ~n2754 & n3402 ) | ( ~n2754 & n3408 ) | ( n3402 & n3408 ) ;
  assign n3410 = ( n3401 & n3407 ) | ( n3401 & ~n3409 ) | ( n3407 & ~n3409 ) ;
  assign n3411 = x170 & ~n761 ;
  assign n3412 = n767 | n788 ;
  assign n3413 = ( ~n727 & n1580 ) | ( ~n727 & n3187 ) | ( n1580 & n3187 ) ;
  assign n3414 = ~n745 & n2265 ;
  assign n3415 = n742 | n745 ;
  assign n3416 = ( n3413 & ~n3414 ) | ( n3413 & n3415 ) | ( ~n3414 & n3415 ) ;
  assign n3417 = ~n735 & n3416 ;
  assign n3418 = ( ~n767 & n778 ) | ( ~n767 & n1852 ) | ( n778 & n1852 ) ;
  assign n3419 = ( ~n3412 & n3417 ) | ( ~n3412 & n3418 ) | ( n3417 & n3418 ) ;
  assign n3420 = n3411 & ~n3419 ;
  assign n3421 = ( ~n1582 & n2068 ) | ( ~n1582 & n2748 ) | ( n2068 & n2748 ) ;
  assign n3422 = ( ~n747 & n2421 ) | ( ~n747 & n3421 ) | ( n2421 & n3421 ) ;
  assign n3423 = ( n3412 & ~n3418 ) | ( n3412 & n3422 ) | ( ~n3418 & n3422 ) ;
  assign n3424 = n3411 & n3423 ;
  assign n3425 = ( n3410 & n3420 ) | ( n3410 & n3424 ) | ( n3420 & n3424 ) ;
  assign n3426 = x45 | n1162 ;
  assign n3427 = ~n802 & n3426 ;
  assign n3428 = ( ~n813 & n825 ) | ( ~n813 & n3427 ) | ( n825 & n3427 ) ;
  assign n3429 = ( ~n819 & n2078 ) | ( ~n819 & n3428 ) | ( n2078 & n3428 ) ;
  assign n3430 = ( n1605 & ~n2082 ) | ( n1605 & n3429 ) | ( ~n2082 & n3429 ) ;
  assign n3431 = n895 | n2278 ;
  assign n3432 = ( ~n895 & n906 ) | ( ~n895 & n2091 ) | ( n906 & n2091 ) ;
  assign n3433 = ( n3095 & n3431 ) | ( n3095 & ~n3432 ) | ( n3431 & ~n3432 ) ;
  assign n3434 = ( n1611 & ~n3431 ) | ( n1611 & n3432 ) | ( ~n3431 & n3432 ) ;
  assign n3435 = ( n3430 & ~n3433 ) | ( n3430 & n3434 ) | ( ~n3433 & n3434 ) ;
  assign n3436 = ~n931 & n975 ;
  assign n3437 = ( ~n954 & n1622 ) | ( ~n954 & n1885 ) | ( n1622 & n1885 ) ;
  assign n3438 = ( ~n1633 & n3436 ) | ( ~n1633 & n3437 ) | ( n3436 & n3437 ) ;
  assign n3439 = ( n1633 & n1883 ) | ( n1633 & ~n3436 ) | ( n1883 & ~n3436 ) ;
  assign n3440 = ( n3435 & ~n3438 ) | ( n3435 & n3439 ) | ( ~n3438 & n3439 ) ;
  assign n3441 = ( n1107 & ~n1674 ) | ( n1107 & n2897 ) | ( ~n1674 & n2897 ) ;
  assign n3442 = ~n993 & n2438 ;
  assign n3443 = ( n1054 & n2126 ) | ( n1054 & ~n2442 ) | ( n2126 & ~n2442 ) ;
  assign n3444 = ( n1043 & ~n1054 ) | ( n1043 & n2300 ) | ( ~n1054 & n2300 ) ;
  assign n3445 = ( n3442 & n3443 ) | ( n3442 & ~n3444 ) | ( n3443 & ~n3444 ) ;
  assign n3446 = ( n2793 & ~n3441 ) | ( n2793 & n3445 ) | ( ~n3441 & n3445 ) ;
  assign n3447 = ( n2889 & ~n3443 ) | ( n2889 & n3444 ) | ( ~n3443 & n3444 ) ;
  assign n3448 = ( ~n2793 & n3441 ) | ( ~n2793 & n3447 ) | ( n3441 & n3447 ) ;
  assign n3449 = ( n3440 & n3446 ) | ( n3440 & ~n3448 ) | ( n3446 & ~n3448 ) ;
  assign n3450 = x171 & ~n1165 ;
  assign n3451 = n1171 | n1192 ;
  assign n3452 = ( ~n1131 & n1678 ) | ( ~n1131 & n3223 ) | ( n1678 & n3223 ) ;
  assign n3453 = ~n1149 & n2321 ;
  assign n3454 = n1146 | n1149 ;
  assign n3455 = ( n3452 & ~n3453 ) | ( n3452 & n3454 ) | ( ~n3453 & n3454 ) ;
  assign n3456 = ~n1139 & n3455 ;
  assign n3457 = ( ~n1171 & n1182 ) | ( ~n1171 & n1930 ) | ( n1182 & n1930 ) ;
  assign n3458 = ( ~n3451 & n3456 ) | ( ~n3451 & n3457 ) | ( n3456 & n3457 ) ;
  assign n3459 = n3450 & ~n3458 ;
  assign n3460 = ( ~n1680 & n2138 ) | ( ~n1680 & n2787 ) | ( n2138 & n2787 ) ;
  assign n3461 = ( ~n1151 & n2465 ) | ( ~n1151 & n3460 ) | ( n2465 & n3460 ) ;
  assign n3462 = ( n3451 & ~n3457 ) | ( n3451 & n3461 ) | ( ~n3457 & n3461 ) ;
  assign n3463 = n3450 & n3462 ;
  assign n3464 = ( n3449 & n3459 ) | ( n3449 & n3463 ) | ( n3459 & n3463 ) ;
  assign n3465 = x46 | n399 ;
  assign n3466 = ~n1206 & n3465 ;
  assign n3467 = ( ~n1217 & n1229 ) | ( ~n1217 & n3466 ) | ( n1229 & n3466 ) ;
  assign n3468 = ( ~n1223 & n2148 ) | ( ~n1223 & n3467 ) | ( n2148 & n3467 ) ;
  assign n3469 = ( n1703 & ~n2152 ) | ( n1703 & n3468 ) | ( ~n2152 & n3468 ) ;
  assign n3470 = n1299 | n2334 ;
  assign n3471 = ( ~n1299 & n1310 ) | ( ~n1299 & n2161 ) | ( n1310 & n2161 ) ;
  assign n3472 = ( n3131 & n3470 ) | ( n3131 & ~n3471 ) | ( n3470 & ~n3471 ) ;
  assign n3473 = ( n1709 & ~n3470 ) | ( n1709 & n3471 ) | ( ~n3470 & n3471 ) ;
  assign n3474 = ( n3469 & ~n3472 ) | ( n3469 & n3473 ) | ( ~n3472 & n3473 ) ;
  assign n3475 = ~n1335 & n1379 ;
  assign n3476 = ( ~n1358 & n1720 ) | ( ~n1358 & n1963 ) | ( n1720 & n1963 ) ;
  assign n3477 = ( ~n1731 & n3475 ) | ( ~n1731 & n3476 ) | ( n3475 & n3476 ) ;
  assign n3478 = ( n1731 & n1961 ) | ( n1731 & ~n3475 ) | ( n1961 & ~n3475 ) ;
  assign n3479 = ( n3474 & ~n3477 ) | ( n3474 & n3478 ) | ( ~n3477 & n3478 ) ;
  assign n3480 = ( ~n294 & n299 ) | ( ~n294 & n2934 ) | ( n299 & n2934 ) ;
  assign n3481 = ~n1397 & n2482 ;
  assign n3482 = ( n1458 & n2196 ) | ( n1458 & ~n2486 ) | ( n2196 & ~n2486 ) ;
  assign n3483 = ( n1447 & ~n1458 ) | ( n1447 & n2356 ) | ( ~n1458 & n2356 ) ;
  assign n3484 = ( n3481 & n3482 ) | ( n3481 & ~n3483 ) | ( n3482 & ~n3483 ) ;
  assign n3485 = ( n2831 & ~n3480 ) | ( n2831 & n3484 ) | ( ~n3480 & n3484 ) ;
  assign n3486 = ( n2926 & ~n3482 ) | ( n2926 & n3483 ) | ( ~n3482 & n3483 ) ;
  assign n3487 = ( ~n2831 & n3480 ) | ( ~n2831 & n3486 ) | ( n3480 & n3486 ) ;
  assign n3488 = ( n3479 & n3485 ) | ( n3479 & ~n3487 ) | ( n3485 & ~n3487 ) ;
  assign n3489 = x172 & ~n396 ;
  assign n3490 = n355 | n1498 ;
  assign n3491 = ( n319 & ~n348 ) | ( n319 & n3259 ) | ( ~n348 & n3259 ) ;
  assign n3492 = ~n327 & n2377 ;
  assign n3493 = n327 | n341 ;
  assign n3494 = ( n3491 & ~n3492 ) | ( n3491 & n3493 ) | ( ~n3492 & n3493 ) ;
  assign n3495 = ~n380 & n3494 ;
  assign n3496 = ( n375 & ~n3490 ) | ( n375 & n3495 ) | ( ~n3490 & n3495 ) ;
  assign n3497 = n3489 & ~n3496 ;
  assign n3498 = ( n323 & ~n337 ) | ( n323 & n2209 ) | ( ~n337 & n2209 ) ;
  assign n3499 = ( ~n1489 & n2509 ) | ( ~n1489 & n3498 ) | ( n2509 & n3498 ) ;
  assign n3500 = ( ~n375 & n3490 ) | ( ~n375 & n3499 ) | ( n3490 & n3499 ) ;
  assign n3501 = n3489 & n3500 ;
  assign n3502 = ( n3488 & n3497 ) | ( n3488 & n3501 ) | ( n3497 & n3501 ) ;
  assign n3503 = x47 | n804 ;
  assign n3504 = ~n407 & n3503 ;
  assign n3505 = ( ~n413 & n421 ) | ( ~n413 & n3504 ) | ( n421 & n3504 ) ;
  assign n3506 = ( n418 & ~n419 ) | ( n418 & n3505 ) | ( ~n419 & n3505 ) ;
  assign n3507 = ( ~n463 & n1789 ) | ( ~n463 & n3506 ) | ( n1789 & n3506 ) ;
  assign n3508 = n481 | n514 ;
  assign n3509 = ( ~n481 & n485 ) | ( ~n481 & n502 ) | ( n485 & n502 ) ;
  assign n3510 = ( n3167 & n3508 ) | ( n3167 & ~n3509 ) | ( n3508 & ~n3509 ) ;
  assign n3511 = ( n1794 & ~n3508 ) | ( n1794 & n3509 ) | ( ~n3508 & n3509 ) ;
  assign n3512 = ( n3507 & ~n3510 ) | ( n3507 & n3511 ) | ( ~n3510 & n3511 ) ;
  assign n3513 = ~n520 & n1539 ;
  assign n3514 = ( n1813 & n2035 ) | ( n1813 & ~n3513 ) | ( n2035 & ~n3513 ) ;
  assign n3515 = ( ~n553 & n567 ) | ( ~n553 & n2029 ) | ( n567 & n2029 ) ;
  assign n3516 = ( ~n1813 & n3513 ) | ( ~n1813 & n3515 ) | ( n3513 & n3515 ) ;
  assign n3517 = ( n3512 & n3514 ) | ( n3512 & ~n3516 ) | ( n3514 & ~n3516 ) ;
  assign n3518 = ( ~n699 & n704 ) | ( ~n699 & n2969 ) | ( n704 & n2969 ) ;
  assign n3519 = ~n581 & n627 ;
  assign n3520 = ( n1562 & n2250 ) | ( n1562 & ~n2251 ) | ( n2250 & ~n2251 ) ;
  assign n3521 = ( n1561 & ~n1562 ) | ( n1561 & n2400 ) | ( ~n1562 & n2400 ) ;
  assign n3522 = ( n3519 & n3520 ) | ( n3519 & ~n3521 ) | ( n3520 & ~n3521 ) ;
  assign n3523 = ( n2868 & ~n3518 ) | ( n2868 & n3522 ) | ( ~n3518 & n3522 ) ;
  assign n3524 = ( n614 & ~n3520 ) | ( n614 & n3521 ) | ( ~n3520 & n3521 ) ;
  assign n3525 = ( ~n2868 & n3518 ) | ( ~n2868 & n3524 ) | ( n3518 & n3524 ) ;
  assign n3526 = ( n3517 & n3523 ) | ( n3517 & ~n3525 ) | ( n3523 & ~n3525 ) ;
  assign n3527 = x173 & ~n801 ;
  assign n3528 = n760 | n1597 ;
  assign n3529 = ( n724 & ~n753 ) | ( n724 & n3298 ) | ( ~n753 & n3298 ) ;
  assign n3530 = ~n732 & n2421 ;
  assign n3531 = n732 | n746 ;
  assign n3532 = ( n3529 & ~n3530 ) | ( n3529 & n3531 ) | ( ~n3530 & n3531 ) ;
  assign n3533 = ~n785 & n3532 ;
  assign n3534 = ( n780 & ~n3528 ) | ( n780 & n3533 ) | ( ~n3528 & n3533 ) ;
  assign n3535 = n3527 & ~n3534 ;
  assign n3536 = ( n728 & ~n742 ) | ( n728 & n2265 ) | ( ~n742 & n2265 ) ;
  assign n3537 = ( ~n1588 & n2546 ) | ( ~n1588 & n3536 ) | ( n2546 & n3536 ) ;
  assign n3538 = ( ~n780 & n3528 ) | ( ~n780 & n3537 ) | ( n3528 & n3537 ) ;
  assign n3539 = n3527 & n3538 ;
  assign n3540 = ( n3526 & n3535 ) | ( n3526 & n3539 ) | ( n3535 & n3539 ) ;
  assign n3541 = x48 | n1208 ;
  assign n3542 = ~n812 & n3541 ;
  assign n3543 = ( ~n818 & n826 ) | ( ~n818 & n3542 ) | ( n826 & n3542 ) ;
  assign n3544 = ( n823 & ~n824 ) | ( n823 & n3543 ) | ( ~n824 & n3543 ) ;
  assign n3545 = ( ~n868 & n1867 ) | ( ~n868 & n3544 ) | ( n1867 & n3544 ) ;
  assign n3546 = n886 | n919 ;
  assign n3547 = ( ~n886 & n890 ) | ( ~n886 & n907 ) | ( n890 & n907 ) ;
  assign n3548 = ( n3203 & n3546 ) | ( n3203 & ~n3547 ) | ( n3546 & ~n3547 ) ;
  assign n3549 = ( n1872 & ~n3546 ) | ( n1872 & n3547 ) | ( ~n3546 & n3547 ) ;
  assign n3550 = ( n3545 & ~n3548 ) | ( n3545 & n3549 ) | ( ~n3548 & n3549 ) ;
  assign n3551 = ~n925 & n1638 ;
  assign n3552 = ( n1891 & n2105 ) | ( n1891 & ~n3551 ) | ( n2105 & ~n3551 ) ;
  assign n3553 = ( ~n958 & n972 ) | ( ~n958 & n2099 ) | ( n972 & n2099 ) ;
  assign n3554 = ( ~n1891 & n3551 ) | ( ~n1891 & n3553 ) | ( n3551 & n3553 ) ;
  assign n3555 = ( n3550 & n3552 ) | ( n3550 & ~n3554 ) | ( n3552 & ~n3554 ) ;
  assign n3556 = ( ~n1103 & n1108 ) | ( ~n1103 & n3005 ) | ( n1108 & n3005 ) ;
  assign n3557 = ~n986 & n1032 ;
  assign n3558 = ( n1661 & n2306 ) | ( n1661 & ~n2307 ) | ( n2306 & ~n2307 ) ;
  assign n3559 = ( n1660 & ~n1661 ) | ( n1660 & n2444 ) | ( ~n1661 & n2444 ) ;
  assign n3560 = ( n3557 & n3558 ) | ( n3557 & ~n3559 ) | ( n3558 & ~n3559 ) ;
  assign n3561 = ( n2905 & ~n3556 ) | ( n2905 & n3560 ) | ( ~n3556 & n3560 ) ;
  assign n3562 = ( n1019 & ~n3558 ) | ( n1019 & n3559 ) | ( ~n3558 & n3559 ) ;
  assign n3563 = ( ~n2905 & n3556 ) | ( ~n2905 & n3562 ) | ( n3556 & n3562 ) ;
  assign n3564 = ( n3555 & n3561 ) | ( n3555 & ~n3563 ) | ( n3561 & ~n3563 ) ;
  assign n3565 = x174 & ~n1205 ;
  assign n3566 = n1164 | n1695 ;
  assign n3567 = ( n1128 & ~n1157 ) | ( n1128 & n3337 ) | ( ~n1157 & n3337 ) ;
  assign n3568 = ~n1136 & n2465 ;
  assign n3569 = n1136 | n1150 ;
  assign n3570 = ( n3567 & ~n3568 ) | ( n3567 & n3569 ) | ( ~n3568 & n3569 ) ;
  assign n3571 = ~n1189 & n3570 ;
  assign n3572 = ( n1184 & ~n3566 ) | ( n1184 & n3571 ) | ( ~n3566 & n3571 ) ;
  assign n3573 = n3565 & ~n3572 ;
  assign n3574 = ( n1132 & ~n1146 ) | ( n1132 & n2321 ) | ( ~n1146 & n2321 ) ;
  assign n3575 = ( ~n1686 & n2583 ) | ( ~n1686 & n3574 ) | ( n2583 & n3574 ) ;
  assign n3576 = ( ~n1184 & n3566 ) | ( ~n1184 & n3575 ) | ( n3566 & n3575 ) ;
  assign n3577 = n3565 & n3576 ;
  assign n3578 = ( n3564 & n3573 ) | ( n3564 & n3577 ) | ( n3573 & n3577 ) ;
  assign n3579 = x49 | n403 ;
  assign n3580 = ~n1216 & n3579 ;
  assign n3581 = ( ~n1222 & n1230 ) | ( ~n1222 & n3580 ) | ( n1230 & n3580 ) ;
  assign n3582 = ( n1227 & ~n1228 ) | ( n1227 & n3581 ) | ( ~n1228 & n3581 ) ;
  assign n3583 = ( ~n1272 & n1945 ) | ( ~n1272 & n3582 ) | ( n1945 & n3582 ) ;
  assign n3584 = n1290 | n1323 ;
  assign n3585 = ( ~n1290 & n1294 ) | ( ~n1290 & n1311 ) | ( n1294 & n1311 ) ;
  assign n3586 = ( n3239 & n3584 ) | ( n3239 & ~n3585 ) | ( n3584 & ~n3585 ) ;
  assign n3587 = ( n1950 & ~n3584 ) | ( n1950 & n3585 ) | ( ~n3584 & n3585 ) ;
  assign n3588 = ( n3583 & ~n3586 ) | ( n3583 & n3587 ) | ( ~n3586 & n3587 ) ;
  assign n3589 = ~n1329 & n1736 ;
  assign n3590 = ( n1969 & n2175 ) | ( n1969 & ~n3589 ) | ( n2175 & ~n3589 ) ;
  assign n3591 = ( ~n1362 & n1376 ) | ( ~n1362 & n2169 ) | ( n1376 & n2169 ) ;
  assign n3592 = ( ~n1969 & n3589 ) | ( ~n1969 & n3591 ) | ( n3589 & n3591 ) ;
  assign n3593 = ( n3588 & n3590 ) | ( n3588 & ~n3592 ) | ( n3590 & ~n3592 ) ;
  assign n3594 = ( n311 & ~n1480 ) | ( n311 & n3042 ) | ( ~n1480 & n3042 ) ;
  assign n3595 = ~n1390 & n1436 ;
  assign n3596 = ( n1756 & n2362 ) | ( n1756 & ~n2363 ) | ( n2362 & ~n2363 ) ;
  assign n3597 = ( n1755 & ~n1756 ) | ( n1755 & n2488 ) | ( ~n1756 & n2488 ) ;
  assign n3598 = ( n3595 & n3596 ) | ( n3595 & ~n3597 ) | ( n3596 & ~n3597 ) ;
  assign n3599 = ( n2942 & ~n3594 ) | ( n2942 & n3598 ) | ( ~n3594 & n3598 ) ;
  assign n3600 = ( n1423 & ~n3596 ) | ( n1423 & n3597 ) | ( ~n3596 & n3597 ) ;
  assign n3601 = ( ~n2942 & n3594 ) | ( ~n2942 & n3600 ) | ( n3594 & n3600 ) ;
  assign n3602 = ( n3593 & n3599 ) | ( n3593 & ~n3601 ) | ( n3599 & ~n3601 ) ;
  assign n3603 = x175 & ~n406 ;
  assign n3604 = n401 | n1782 ;
  assign n3605 = ( ~n349 & n1484 ) | ( ~n349 & n3376 ) | ( n1484 & n3376 ) ;
  assign n3606 = ~n365 & n2509 ;
  assign n3607 = n365 | n1488 ;
  assign n3608 = ( n3605 & ~n3606 ) | ( n3605 & n3607 ) | ( ~n3606 & n3607 ) ;
  assign n3609 = ~n368 & n3608 ;
  assign n3610 = ( n1495 & ~n3604 ) | ( n1495 & n3609 ) | ( ~n3604 & n3609 ) ;
  assign n3611 = n3603 & ~n3610 ;
  assign n3612 = ( ~n341 & n1486 ) | ( ~n341 & n2377 ) | ( n1486 & n2377 ) ;
  assign n3613 = ( ~n1774 & n2618 ) | ( ~n1774 & n3612 ) | ( n2618 & n3612 ) ;
  assign n3614 = ( ~n1495 & n3604 ) | ( ~n1495 & n3613 ) | ( n3604 & n3613 ) ;
  assign n3615 = n3603 & n3614 ;
  assign n3616 = ( n3602 & n3611 ) | ( n3602 & n3615 ) | ( n3611 & n3615 ) ;
  assign n3617 = x50 | n808 ;
  assign n3618 = ~n412 & n3617 ;
  assign n3619 = ( ~n391 & n395 ) | ( ~n391 & n3618 ) | ( n395 & n3618 ) ;
  assign n3620 = ( ~n461 & n1506 ) | ( ~n461 & n3619 ) | ( n1506 & n3619 ) ;
  assign n3621 = ( ~n1515 & n2016 ) | ( ~n1515 & n3620 ) | ( n2016 & n3620 ) ;
  assign n3622 = n506 | n1526 ;
  assign n3623 = ( ~n506 & n511 ) | ( ~n506 & n1521 ) | ( n511 & n1521 ) ;
  assign n3624 = ( n3275 & n3622 ) | ( n3275 & ~n3623 ) | ( n3622 & ~n3623 ) ;
  assign n3625 = ( n2021 & ~n3622 ) | ( n2021 & n3623 ) | ( ~n3622 & n3623 ) ;
  assign n3626 = ( n3621 & ~n3624 ) | ( n3621 & n3625 ) | ( ~n3624 & n3625 ) ;
  assign n3627 = ~n603 & n1818 ;
  assign n3628 = ( ~n537 & n568 ) | ( ~n537 & n2226 ) | ( n568 & n2226 ) ;
  assign n3629 = ( ~n2040 & n3627 ) | ( ~n2040 & n3628 ) | ( n3627 & n3628 ) ;
  assign n3630 = ( n2040 & n2231 ) | ( n2040 & ~n3627 ) | ( n2231 & ~n3627 ) ;
  assign n3631 = ( n3626 & ~n3629 ) | ( n3626 & n3630 ) | ( ~n3629 & n3630 ) ;
  assign n3632 = ( n716 & ~n1579 ) | ( n716 & n3077 ) | ( ~n1579 & n3077 ) ;
  assign n3633 = ~n575 & n1554 ;
  assign n3634 = ( n1834 & n2406 ) | ( n1834 & ~n2407 ) | ( n2406 & ~n2407 ) ;
  assign n3635 = ( n1833 & ~n1834 ) | ( n1833 & n2526 ) | ( ~n1834 & n2526 ) ;
  assign n3636 = ( n3633 & n3634 ) | ( n3633 & ~n3635 ) | ( n3634 & ~n3635 ) ;
  assign n3637 = ( n2978 & ~n3632 ) | ( n2978 & n3636 ) | ( ~n3632 & n3636 ) ;
  assign n3638 = ( n1545 & ~n3634 ) | ( n1545 & n3635 ) | ( ~n3634 & n3635 ) ;
  assign n3639 = ( ~n2978 & n3632 ) | ( ~n2978 & n3638 ) | ( n3632 & n3638 ) ;
  assign n3640 = ( n3631 & n3637 ) | ( n3631 & ~n3639 ) | ( n3637 & ~n3639 ) ;
  assign n3641 = x176 & ~n811 ;
  assign n3642 = n806 | n1860 ;
  assign n3643 = ( ~n754 & n1583 ) | ( ~n754 & n3415 ) | ( n1583 & n3415 ) ;
  assign n3644 = ~n770 & n2546 ;
  assign n3645 = n770 | n1587 ;
  assign n3646 = ( n3643 & ~n3644 ) | ( n3643 & n3645 ) | ( ~n3644 & n3645 ) ;
  assign n3647 = ~n773 & n3646 ;
  assign n3648 = ( n1594 & ~n3642 ) | ( n1594 & n3647 ) | ( ~n3642 & n3647 ) ;
  assign n3649 = n3641 & ~n3648 ;
  assign n3650 = ( ~n746 & n1585 ) | ( ~n746 & n2421 ) | ( n1585 & n2421 ) ;
  assign n3651 = ( ~n1852 & n2653 ) | ( ~n1852 & n3650 ) | ( n2653 & n3650 ) ;
  assign n3652 = ( ~n1594 & n3642 ) | ( ~n1594 & n3651 ) | ( n3642 & n3651 ) ;
  assign n3653 = n3641 & n3652 ;
  assign n3654 = ( n3640 & n3649 ) | ( n3640 & n3653 ) | ( n3649 & n3653 ) ;
  assign n3655 = x51 | n1212 ;
  assign n3656 = ~n817 & n3655 ;
  assign n3657 = ( ~n796 & n800 ) | ( ~n796 & n3656 ) | ( n800 & n3656 ) ;
  assign n3658 = ( ~n866 & n1605 ) | ( ~n866 & n3657 ) | ( n1605 & n3657 ) ;
  assign n3659 = ( ~n1614 & n2086 ) | ( ~n1614 & n3658 ) | ( n2086 & n3658 ) ;
  assign n3660 = n911 | n1625 ;
  assign n3661 = ( ~n911 & n916 ) | ( ~n911 & n1620 ) | ( n916 & n1620 ) ;
  assign n3662 = ( n3314 & n3660 ) | ( n3314 & ~n3661 ) | ( n3660 & ~n3661 ) ;
  assign n3663 = ( n2091 & ~n3660 ) | ( n2091 & n3661 ) | ( ~n3660 & n3661 ) ;
  assign n3664 = ( n3659 & ~n3662 ) | ( n3659 & n3663 ) | ( ~n3662 & n3663 ) ;
  assign n3665 = ~n1008 & n1896 ;
  assign n3666 = ( ~n942 & n973 ) | ( ~n942 & n2282 ) | ( n973 & n2282 ) ;
  assign n3667 = ( ~n2110 & n3665 ) | ( ~n2110 & n3666 ) | ( n3665 & n3666 ) ;
  assign n3668 = ( n2110 & n2287 ) | ( n2110 & ~n3665 ) | ( n2287 & ~n3665 ) ;
  assign n3669 = ( n3664 & ~n3667 ) | ( n3664 & n3668 ) | ( ~n3667 & n3668 ) ;
  assign n3670 = ( n1120 & ~n1677 ) | ( n1120 & n3113 ) | ( ~n1677 & n3113 ) ;
  assign n3671 = ~n980 & n1653 ;
  assign n3672 = ( n1912 & n2450 ) | ( n1912 & ~n2451 ) | ( n2450 & ~n2451 ) ;
  assign n3673 = ( n1911 & ~n1912 ) | ( n1911 & n2563 ) | ( ~n1912 & n2563 ) ;
  assign n3674 = ( n3671 & n3672 ) | ( n3671 & ~n3673 ) | ( n3672 & ~n3673 ) ;
  assign n3675 = ( n3014 & ~n3670 ) | ( n3014 & n3674 ) | ( ~n3670 & n3674 ) ;
  assign n3676 = ( n1644 & ~n3672 ) | ( n1644 & n3673 ) | ( ~n3672 & n3673 ) ;
  assign n3677 = ( ~n3014 & n3670 ) | ( ~n3014 & n3676 ) | ( n3670 & n3676 ) ;
  assign n3678 = ( n3669 & n3675 ) | ( n3669 & ~n3677 ) | ( n3675 & ~n3677 ) ;
  assign n3679 = x177 & ~n1215 ;
  assign n3680 = n1210 | n1938 ;
  assign n3681 = ( ~n1158 & n1681 ) | ( ~n1158 & n3454 ) | ( n1681 & n3454 ) ;
  assign n3682 = ~n1174 & n2583 ;
  assign n3683 = n1174 | n1685 ;
  assign n3684 = ( n3681 & ~n3682 ) | ( n3681 & n3683 ) | ( ~n3682 & n3683 ) ;
  assign n3685 = ~n1177 & n3684 ;
  assign n3686 = ( n1692 & ~n3680 ) | ( n1692 & n3685 ) | ( ~n3680 & n3685 ) ;
  assign n3687 = n3679 & ~n3686 ;
  assign n3688 = ( ~n1150 & n1683 ) | ( ~n1150 & n2465 ) | ( n1683 & n2465 ) ;
  assign n3689 = ( ~n1930 & n2688 ) | ( ~n1930 & n3688 ) | ( n2688 & n3688 ) ;
  assign n3690 = ( ~n1692 & n3680 ) | ( ~n1692 & n3689 ) | ( n3680 & n3689 ) ;
  assign n3691 = n3679 & n3690 ;
  assign n3692 = ( n3678 & n3687 ) | ( n3678 & n3691 ) | ( n3687 & n3691 ) ;
  assign n3693 = x52 | n392 ;
  assign n3694 = ~n1221 & n3693 ;
  assign n3695 = ( ~n1200 & n1204 ) | ( ~n1200 & n3694 ) | ( n1204 & n3694 ) ;
  assign n3696 = ( ~n1270 & n1703 ) | ( ~n1270 & n3695 ) | ( n1703 & n3695 ) ;
  assign n3697 = ( ~n1712 & n2156 ) | ( ~n1712 & n3696 ) | ( n2156 & n3696 ) ;
  assign n3698 = n1315 | n1723 ;
  assign n3699 = ( ~n1315 & n1320 ) | ( ~n1315 & n1718 ) | ( n1320 & n1718 ) ;
  assign n3700 = ( n3353 & n3698 ) | ( n3353 & ~n3699 ) | ( n3698 & ~n3699 ) ;
  assign n3701 = ( n2161 & ~n3698 ) | ( n2161 & n3699 ) | ( ~n3698 & n3699 ) ;
  assign n3702 = ( n3697 & ~n3700 ) | ( n3697 & n3701 ) | ( ~n3700 & n3701 ) ;
  assign n3703 = ~n1412 & n1974 ;
  assign n3704 = ( ~n1346 & n1377 ) | ( ~n1346 & n2338 ) | ( n1377 & n2338 ) ;
  assign n3705 = ( ~n2180 & n3703 ) | ( ~n2180 & n3704 ) | ( n3703 & n3704 ) ;
  assign n3706 = ( n2180 & n2343 ) | ( n2180 & ~n3703 ) | ( n2343 & ~n3703 ) ;
  assign n3707 = ( n3702 & ~n3705 ) | ( n3702 & n3706 ) | ( ~n3705 & n3706 ) ;
  assign n3708 = ( n318 & ~n1765 ) | ( n318 & n3149 ) | ( ~n1765 & n3149 ) ;
  assign n3709 = ~n1384 & n1751 ;
  assign n3710 = ( n269 & n2494 ) | ( n269 & ~n2495 ) | ( n2494 & ~n2495 ) ;
  assign n3711 = ( n265 & ~n269 ) | ( n265 & n2600 ) | ( ~n269 & n2600 ) ;
  assign n3712 = ( n3709 & n3710 ) | ( n3709 & ~n3711 ) | ( n3710 & ~n3711 ) ;
  assign n3713 = ( n3050 & ~n3708 ) | ( n3050 & n3712 ) | ( ~n3708 & n3712 ) ;
  assign n3714 = ( n1742 & ~n3710 ) | ( n1742 & n3711 ) | ( ~n3710 & n3711 ) ;
  assign n3715 = ( ~n3050 & n3708 ) | ( ~n3050 & n3714 ) | ( n3708 & n3714 ) ;
  assign n3716 = ( n3707 & n3713 ) | ( n3707 & ~n3715 ) | ( n3713 & ~n3715 ) ;
  assign n3717 = x178 & ~n411 ;
  assign n3718 = n405 | n2009 ;
  assign n3719 = ( ~n344 & n1771 ) | ( ~n344 & n3493 ) | ( n1771 & n3493 ) ;
  assign n3720 = ~n372 & n2618 ;
  assign n3721 = n369 | n372 ;
  assign n3722 = ( n3719 & ~n3720 ) | ( n3719 & n3721 ) | ( ~n3720 & n3721 ) ;
  assign n3723 = ~n362 & n3722 ;
  assign n3724 = ( n1780 & ~n3718 ) | ( n1780 & n3723 ) | ( ~n3718 & n3723 ) ;
  assign n3725 = n3717 & ~n3724 ;
  assign n3726 = ( n350 & ~n1488 ) | ( n350 & n2509 ) | ( ~n1488 & n2509 ) ;
  assign n3727 = ( ~n374 & n2719 ) | ( ~n374 & n3726 ) | ( n2719 & n3726 ) ;
  assign n3728 = ( ~n1780 & n3718 ) | ( ~n1780 & n3727 ) | ( n3718 & n3727 ) ;
  assign n3729 = n3717 & n3728 ;
  assign n3730 = ( n3716 & n3725 ) | ( n3716 & n3729 ) | ( n3725 & n3729 ) ;
  assign n3731 = x53 | n797 ;
  assign n3732 = ~n390 & n3731 ;
  assign n3733 = ( ~n460 & n1501 ) | ( ~n460 & n3732 ) | ( n1501 & n3732 ) ;
  assign n3734 = ( ~n462 & n1789 ) | ( ~n462 & n3733 ) | ( n1789 & n3733 ) ;
  assign n3735 = ( n438 & ~n1797 ) | ( n438 & n3734 ) | ( ~n1797 & n3734 ) ;
  assign n3736 = n471 | n1807 ;
  assign n3737 = ( ~n471 & n475 ) | ( ~n471 & n1804 ) | ( n475 & n1804 ) ;
  assign n3738 = ( n3392 & n3736 ) | ( n3392 & ~n3737 ) | ( n3736 & ~n3737 ) ;
  assign n3739 = ( n502 & ~n3736 ) | ( n502 & n3737 ) | ( ~n3736 & n3737 ) ;
  assign n3740 = ( n3735 & ~n3738 ) | ( n3735 & n3739 ) | ( ~n3738 & n3739 ) ;
  assign n3741 = ~n607 & n2045 ;
  assign n3742 = ( ~n531 & n540 ) | ( ~n531 & n569 ) | ( n540 & n569 ) ;
  assign n3743 = ( ~n2235 & n3741 ) | ( ~n2235 & n3742 ) | ( n3741 & n3742 ) ;
  assign n3744 = ( n556 & n2235 ) | ( n556 & ~n3741 ) | ( n2235 & ~n3741 ) ;
  assign n3745 = ( n3740 & ~n3743 ) | ( n3740 & n3744 ) | ( ~n3743 & n3744 ) ;
  assign n3746 = ( n723 & ~n1843 ) | ( n723 & n3185 ) | ( ~n1843 & n3185 ) ;
  assign n3747 = ~n655 & n1830 ;
  assign n3748 = ( n674 & n2531 ) | ( n674 & ~n2532 ) | ( n2531 & ~n2532 ) ;
  assign n3749 = ( n670 & ~n674 ) | ( n670 & n2635 ) | ( ~n674 & n2635 ) ;
  assign n3750 = ( n3747 & n3748 ) | ( n3747 & ~n3749 ) | ( n3748 & ~n3749 ) ;
  assign n3751 = ( n3086 & ~n3746 ) | ( n3086 & n3750 ) | ( ~n3746 & n3750 ) ;
  assign n3752 = ( n1823 & ~n3748 ) | ( n1823 & n3749 ) | ( ~n3748 & n3749 ) ;
  assign n3753 = ( ~n3086 & n3746 ) | ( ~n3086 & n3752 ) | ( n3746 & n3752 ) ;
  assign n3754 = ( n3745 & n3751 ) | ( n3745 & ~n3753 ) | ( n3751 & ~n3753 ) ;
  assign n3755 = x179 & ~n816 ;
  assign n3756 = n810 | n2079 ;
  assign n3757 = ( ~n749 & n1849 ) | ( ~n749 & n3531 ) | ( n1849 & n3531 ) ;
  assign n3758 = ~n777 & n2653 ;
  assign n3759 = n774 | n777 ;
  assign n3760 = ( n3757 & ~n3758 ) | ( n3757 & n3759 ) | ( ~n3758 & n3759 ) ;
  assign n3761 = ~n767 & n3760 ;
  assign n3762 = ( n1858 & ~n3756 ) | ( n1858 & n3761 ) | ( ~n3756 & n3761 ) ;
  assign n3763 = n3755 & ~n3762 ;
  assign n3764 = ( n755 & ~n1587 ) | ( n755 & n2546 ) | ( ~n1587 & n2546 ) ;
  assign n3765 = ( ~n779 & n2758 ) | ( ~n779 & n3764 ) | ( n2758 & n3764 ) ;
  assign n3766 = ( ~n1858 & n3756 ) | ( ~n1858 & n3765 ) | ( n3756 & n3765 ) ;
  assign n3767 = n3755 & n3766 ;
  assign n3768 = ( n3754 & n3763 ) | ( n3754 & n3767 ) | ( n3763 & n3767 ) ;
  assign n3769 = x54 | n1201 ;
  assign n3770 = ~n795 & n3769 ;
  assign n3771 = ( ~n865 & n1600 ) | ( ~n865 & n3770 ) | ( n1600 & n3770 ) ;
  assign n3772 = ( ~n867 & n1867 ) | ( ~n867 & n3771 ) | ( n1867 & n3771 ) ;
  assign n3773 = ( n843 & ~n1875 ) | ( n843 & n3772 ) | ( ~n1875 & n3772 ) ;
  assign n3774 = n876 | n1885 ;
  assign n3775 = ( ~n876 & n880 ) | ( ~n876 & n1882 ) | ( n880 & n1882 ) ;
  assign n3776 = ( n3431 & n3774 ) | ( n3431 & ~n3775 ) | ( n3774 & ~n3775 ) ;
  assign n3777 = ( n907 & ~n3774 ) | ( n907 & n3775 ) | ( ~n3774 & n3775 ) ;
  assign n3778 = ( n3773 & ~n3776 ) | ( n3773 & n3777 ) | ( ~n3776 & n3777 ) ;
  assign n3779 = ~n1012 & n2115 ;
  assign n3780 = ( ~n936 & n945 ) | ( ~n936 & n974 ) | ( n945 & n974 ) ;
  assign n3781 = ( ~n2291 & n3779 ) | ( ~n2291 & n3780 ) | ( n3779 & n3780 ) ;
  assign n3782 = ( n961 & n2291 ) | ( n961 & ~n3779 ) | ( n2291 & ~n3779 ) ;
  assign n3783 = ( n3778 & ~n3781 ) | ( n3778 & n3782 ) | ( ~n3781 & n3782 ) ;
  assign n3784 = ( n1127 & ~n1921 ) | ( n1127 & n3221 ) | ( ~n1921 & n3221 ) ;
  assign n3785 = ~n1060 & n1908 ;
  assign n3786 = ( n1078 & n2568 ) | ( n1078 & ~n2569 ) | ( n2568 & ~n2569 ) ;
  assign n3787 = ( n1074 & ~n1078 ) | ( n1074 & n2670 ) | ( ~n1078 & n2670 ) ;
  assign n3788 = ( n3785 & n3786 ) | ( n3785 & ~n3787 ) | ( n3786 & ~n3787 ) ;
  assign n3789 = ( n3122 & ~n3784 ) | ( n3122 & n3788 ) | ( ~n3784 & n3788 ) ;
  assign n3790 = ( n1901 & ~n3786 ) | ( n1901 & n3787 ) | ( ~n3786 & n3787 ) ;
  assign n3791 = ( ~n3122 & n3784 ) | ( ~n3122 & n3790 ) | ( n3784 & n3790 ) ;
  assign n3792 = ( n3783 & n3789 ) | ( n3783 & ~n3791 ) | ( n3789 & ~n3791 ) ;
  assign n3793 = x180 & ~n1220 ;
  assign n3794 = n1214 | n2149 ;
  assign n3795 = ( ~n1153 & n1927 ) | ( ~n1153 & n3569 ) | ( n1927 & n3569 ) ;
  assign n3796 = ~n1181 & n2688 ;
  assign n3797 = n1178 | n1181 ;
  assign n3798 = ( n3795 & ~n3796 ) | ( n3795 & n3797 ) | ( ~n3796 & n3797 ) ;
  assign n3799 = ~n1171 & n3798 ;
  assign n3800 = ( n1936 & ~n3794 ) | ( n1936 & n3799 ) | ( ~n3794 & n3799 ) ;
  assign n3801 = n3793 & ~n3800 ;
  assign n3802 = ( n1159 & ~n1685 ) | ( n1159 & n2583 ) | ( ~n1685 & n2583 ) ;
  assign n3803 = ( ~n1183 & n2797 ) | ( ~n1183 & n3802 ) | ( n2797 & n3802 ) ;
  assign n3804 = ( ~n1936 & n3794 ) | ( ~n1936 & n3803 ) | ( n3794 & n3803 ) ;
  assign n3805 = n3793 & n3804 ;
  assign n3806 = ( n3792 & n3801 ) | ( n3792 & n3805 ) | ( n3801 & n3805 ) ;
  assign n3807 = x55 | n386 ;
  assign n3808 = ~n1199 & n3807 ;
  assign n3809 = ( ~n1269 & n1698 ) | ( ~n1269 & n3808 ) | ( n1698 & n3808 ) ;
  assign n3810 = ( ~n1271 & n1945 ) | ( ~n1271 & n3809 ) | ( n1945 & n3809 ) ;
  assign n3811 = ( n1247 & ~n1953 ) | ( n1247 & n3810 ) | ( ~n1953 & n3810 ) ;
  assign n3812 = n1280 | n1963 ;
  assign n3813 = ( ~n1280 & n1284 ) | ( ~n1280 & n1960 ) | ( n1284 & n1960 ) ;
  assign n3814 = ( n3470 & n3812 ) | ( n3470 & ~n3813 ) | ( n3812 & ~n3813 ) ;
  assign n3815 = ( n1311 & ~n3812 ) | ( n1311 & n3813 ) | ( ~n3812 & n3813 ) ;
  assign n3816 = ( n3811 & ~n3814 ) | ( n3811 & n3815 ) | ( ~n3814 & n3815 ) ;
  assign n3817 = ~n1416 & n2185 ;
  assign n3818 = ( ~n1340 & n1349 ) | ( ~n1340 & n1378 ) | ( n1349 & n1378 ) ;
  assign n3819 = ( ~n2347 & n3817 ) | ( ~n2347 & n3818 ) | ( n3817 & n3818 ) ;
  assign n3820 = ( n1365 & n2347 ) | ( n1365 & ~n3817 ) | ( n2347 & ~n3817 ) ;
  assign n3821 = ( n3816 & ~n3819 ) | ( n3816 & n3820 ) | ( ~n3819 & n3820 ) ;
  assign n3822 = ( n1483 & ~n1998 ) | ( n1483 & n3257 ) | ( ~n1998 & n3257 ) ;
  assign n3823 = ~n1464 & n1986 ;
  assign n3824 = ( n277 & n2604 ) | ( n277 & ~n2605 ) | ( n2604 & ~n2605 ) ;
  assign n3825 = ( n273 & ~n277 ) | ( n273 & n2705 ) | ( ~n277 & n2705 ) ;
  assign n3826 = ( n3823 & n3824 ) | ( n3823 & ~n3825 ) | ( n3824 & ~n3825 ) ;
  assign n3827 = ( n3158 & ~n3822 ) | ( n3158 & n3826 ) | ( ~n3822 & n3826 ) ;
  assign n3828 = ( n1979 & ~n3824 ) | ( n1979 & n3825 ) | ( ~n3824 & n3825 ) ;
  assign n3829 = ( ~n3158 & n3822 ) | ( ~n3158 & n3828 ) | ( n3822 & n3828 ) ;
  assign n3830 = ( n3821 & n3827 ) | ( n3821 & ~n3829 ) | ( n3827 & ~n3829 ) ;
  assign n3831 = x181 & ~n389 ;
  assign n3832 = n394 | n422 ;
  assign n3833 = ( n342 & ~n381 ) | ( n342 & n3607 ) | ( ~n381 & n3607 ) ;
  assign n3834 = ~n358 & n2719 ;
  assign n3835 = n358 | n373 ;
  assign n3836 = ( n3833 & ~n3834 ) | ( n3833 & n3835 ) | ( ~n3834 & n3835 ) ;
  assign n3837 = ~n355 & n3836 ;
  assign n3838 = ( n2007 & ~n3832 ) | ( n2007 & n3837 ) | ( ~n3832 & n3837 ) ;
  assign n3839 = n3831 & ~n3838 ;
  assign n3840 = ( ~n369 & n1491 ) | ( ~n369 & n2618 ) | ( n1491 & n2618 ) ;
  assign n3841 = ( n377 & ~n1494 ) | ( n377 & n3840 ) | ( ~n1494 & n3840 ) ;
  assign n3842 = ( ~n2007 & n3832 ) | ( ~n2007 & n3841 ) | ( n3832 & n3841 ) ;
  assign n3843 = n3831 & n3842 ;
  assign n3844 = ( n3830 & n3839 ) | ( n3830 & n3843 ) | ( n3839 & n3843 ) ;
  assign n3845 = x56 | n791 ;
  assign n3846 = ~n459 & n3845 ;
  assign n3847 = ( ~n445 & n449 ) | ( ~n445 & n3846 ) | ( n449 & n3846 ) ;
  assign n3848 = ( ~n464 & n2016 ) | ( ~n464 & n3847 ) | ( n2016 & n3847 ) ;
  assign n3849 = ( n1510 & ~n2024 ) | ( n1510 & n3848 ) | ( ~n2024 & n3848 ) ;
  assign n3850 = n546 | n2029 ;
  assign n3851 = ( ~n546 & n550 ) | ( ~n546 & n2034 ) | ( n550 & n2034 ) ;
  assign n3852 = ( n3508 & n3850 ) | ( n3508 & ~n3851 ) | ( n3850 & ~n3851 ) ;
  assign n3853 = ( n1521 & ~n3850 ) | ( n1521 & n3851 ) | ( ~n3850 & n3851 ) ;
  assign n3854 = ( n3849 & ~n3852 ) | ( n3849 & n3853 ) | ( ~n3852 & n3853 ) ;
  assign n3855 = ~n594 & n2239 ;
  assign n3856 = ( ~n526 & n560 ) | ( ~n526 & n1538 ) | ( n560 & n1538 ) ;
  assign n3857 = ( ~n2394 & n3855 ) | ( ~n2394 & n3856 ) | ( n3855 & n3856 ) ;
  assign n3858 = ( n1534 & n2394 ) | ( n1534 & ~n3855 ) | ( n2394 & ~n3855 ) ;
  assign n3859 = ( n3854 & ~n3857 ) | ( n3854 & n3858 ) | ( ~n3857 & n3858 ) ;
  assign n3860 = ( n1582 & ~n2068 ) | ( n1582 & n3296 ) | ( ~n2068 & n3296 ) ;
  assign n3861 = ~n641 & n2056 ;
  assign n3862 = ( n678 & ~n682 ) | ( n678 & n2745 ) | ( ~n682 & n2745 ) ;
  assign n3863 = ( n682 & n2639 ) | ( n682 & ~n2640 ) | ( n2639 & ~n2640 ) ;
  assign n3864 = ( n3861 & ~n3862 ) | ( n3861 & n3863 ) | ( ~n3862 & n3863 ) ;
  assign n3865 = ( n3194 & ~n3860 ) | ( n3194 & n3864 ) | ( ~n3860 & n3864 ) ;
  assign n3866 = ( n3288 & n3862 ) | ( n3288 & ~n3863 ) | ( n3862 & ~n3863 ) ;
  assign n3867 = ( ~n3194 & n3860 ) | ( ~n3194 & n3866 ) | ( n3860 & n3866 ) ;
  assign n3868 = ( n3859 & n3865 ) | ( n3859 & ~n3867 ) | ( n3865 & ~n3867 ) ;
  assign n3869 = x182 & ~n794 ;
  assign n3870 = n799 | n827 ;
  assign n3871 = ( n747 & ~n786 ) | ( n747 & n3645 ) | ( ~n786 & n3645 ) ;
  assign n3872 = ~n763 & n2758 ;
  assign n3873 = n763 | n778 ;
  assign n3874 = ( n3871 & ~n3872 ) | ( n3871 & n3873 ) | ( ~n3872 & n3873 ) ;
  assign n3875 = ~n760 & n3874 ;
  assign n3876 = ( n2077 & ~n3870 ) | ( n2077 & n3875 ) | ( ~n3870 & n3875 ) ;
  assign n3877 = n3869 & ~n3876 ;
  assign n3878 = ( ~n774 & n1590 ) | ( ~n774 & n2653 ) | ( n1590 & n2653 ) ;
  assign n3879 = ( n782 & ~n1593 ) | ( n782 & n3878 ) | ( ~n1593 & n3878 ) ;
  assign n3880 = ( ~n2077 & n3870 ) | ( ~n2077 & n3879 ) | ( n3870 & n3879 ) ;
  assign n3881 = n3869 & n3880 ;
  assign n3882 = ( n3868 & n3877 ) | ( n3868 & n3881 ) | ( n3877 & n3881 ) ;
  assign n3883 = x57 | n1195 ;
  assign n3884 = ~n864 & n3883 ;
  assign n3885 = ( ~n850 & n854 ) | ( ~n850 & n3884 ) | ( n854 & n3884 ) ;
  assign n3886 = ( ~n869 & n2086 ) | ( ~n869 & n3885 ) | ( n2086 & n3885 ) ;
  assign n3887 = ( n1609 & ~n2094 ) | ( n1609 & n3886 ) | ( ~n2094 & n3886 ) ;
  assign n3888 = n951 | n2099 ;
  assign n3889 = ( ~n951 & n955 ) | ( ~n951 & n2104 ) | ( n955 & n2104 ) ;
  assign n3890 = ( n3546 & n3888 ) | ( n3546 & ~n3889 ) | ( n3888 & ~n3889 ) ;
  assign n3891 = ( n1620 & ~n3888 ) | ( n1620 & n3889 ) | ( ~n3888 & n3889 ) ;
  assign n3892 = ( n3887 & ~n3890 ) | ( n3887 & n3891 ) | ( ~n3890 & n3891 ) ;
  assign n3893 = ~n999 & n2295 ;
  assign n3894 = ( ~n931 & n965 ) | ( ~n931 & n1637 ) | ( n965 & n1637 ) ;
  assign n3895 = ( ~n2438 & n3893 ) | ( ~n2438 & n3894 ) | ( n3893 & n3894 ) ;
  assign n3896 = ( n1633 & n2438 ) | ( n1633 & ~n3893 ) | ( n2438 & ~n3893 ) ;
  assign n3897 = ( n3892 & ~n3895 ) | ( n3892 & n3896 ) | ( ~n3895 & n3896 ) ;
  assign n3898 = ( n1680 & ~n2138 ) | ( n1680 & n3335 ) | ( ~n2138 & n3335 ) ;
  assign n3899 = ~n1046 & n2126 ;
  assign n3900 = ( n1082 & ~n1086 ) | ( n1082 & n2784 ) | ( ~n1086 & n2784 ) ;
  assign n3901 = ( n1086 & n2674 ) | ( n1086 & ~n2675 ) | ( n2674 & ~n2675 ) ;
  assign n3902 = ( n3899 & ~n3900 ) | ( n3899 & n3901 ) | ( ~n3900 & n3901 ) ;
  assign n3903 = ( n3230 & ~n3898 ) | ( n3230 & n3902 ) | ( ~n3898 & n3902 ) ;
  assign n3904 = ( n3327 & n3900 ) | ( n3327 & ~n3901 ) | ( n3900 & ~n3901 ) ;
  assign n3905 = ( ~n3230 & n3898 ) | ( ~n3230 & n3904 ) | ( n3898 & n3904 ) ;
  assign n3906 = ( n3897 & n3903 ) | ( n3897 & ~n3905 ) | ( n3903 & ~n3905 ) ;
  assign n3907 = x183 & ~n1198 ;
  assign n3908 = n1203 | n1231 ;
  assign n3909 = ( n1151 & ~n1190 ) | ( n1151 & n3683 ) | ( ~n1190 & n3683 ) ;
  assign n3910 = ~n1167 & n2797 ;
  assign n3911 = n1167 | n1182 ;
  assign n3912 = ( n3909 & ~n3910 ) | ( n3909 & n3911 ) | ( ~n3910 & n3911 ) ;
  assign n3913 = ~n1164 & n3912 ;
  assign n3914 = ( n2147 & ~n3908 ) | ( n2147 & n3913 ) | ( ~n3908 & n3913 ) ;
  assign n3915 = n3907 & ~n3914 ;
  assign n3916 = ( ~n1178 & n1688 ) | ( ~n1178 & n2688 ) | ( n1688 & n2688 ) ;
  assign n3917 = ( n1186 & ~n1691 ) | ( n1186 & n3916 ) | ( ~n1691 & n3916 ) ;
  assign n3918 = ( ~n2147 & n3908 ) | ( ~n2147 & n3917 ) | ( n3908 & n3917 ) ;
  assign n3919 = n3907 & n3918 ;
  assign n3920 = ( n3906 & n3915 ) | ( n3906 & n3919 ) | ( n3915 & n3919 ) ;
  assign n3921 = x58 | n446 ;
  assign n3922 = ~n1268 & n3921 ;
  assign n3923 = ( ~n1254 & n1258 ) | ( ~n1254 & n3922 ) | ( n1258 & n3922 ) ;
  assign n3924 = ( ~n1273 & n2156 ) | ( ~n1273 & n3923 ) | ( n2156 & n3923 ) ;
  assign n3925 = ( n1707 & ~n2164 ) | ( n1707 & n3924 ) | ( ~n2164 & n3924 ) ;
  assign n3926 = n1355 | n2169 ;
  assign n3927 = ( ~n1355 & n1359 ) | ( ~n1355 & n2174 ) | ( n1359 & n2174 ) ;
  assign n3928 = ( n3584 & n3926 ) | ( n3584 & ~n3927 ) | ( n3926 & ~n3927 ) ;
  assign n3929 = ( n1718 & ~n3926 ) | ( n1718 & n3927 ) | ( ~n3926 & n3927 ) ;
  assign n3930 = ( n3925 & ~n3928 ) | ( n3925 & n3929 ) | ( ~n3928 & n3929 ) ;
  assign n3931 = ~n1403 & n2351 ;
  assign n3932 = ( ~n1335 & n1369 ) | ( ~n1335 & n1735 ) | ( n1369 & n1735 ) ;
  assign n3933 = ( ~n2482 & n3931 ) | ( ~n2482 & n3932 ) | ( n3931 & n3932 ) ;
  assign n3934 = ( n1731 & n2482 ) | ( n1731 & ~n3931 ) | ( n2482 & ~n3931 ) ;
  assign n3935 = ( n3930 & ~n3933 ) | ( n3930 & n3934 ) | ( ~n3933 & n3934 ) ;
  assign n3936 = ( n337 & ~n2209 ) | ( n337 & n3374 ) | ( ~n2209 & n3374 ) ;
  assign n3937 = ~n1450 & n2196 ;
  assign n3938 = ( n297 & ~n1476 ) | ( n297 & n2823 ) | ( ~n1476 & n2823 ) ;
  assign n3939 = ( n1476 & n2709 ) | ( n1476 & ~n2710 ) | ( n2709 & ~n2710 ) ;
  assign n3940 = ( n3937 & ~n3938 ) | ( n3937 & n3939 ) | ( ~n3938 & n3939 ) ;
  assign n3941 = ( n3266 & ~n3936 ) | ( n3266 & n3940 ) | ( ~n3936 & n3940 ) ;
  assign n3942 = ( n3366 & n3938 ) | ( n3366 & ~n3939 ) | ( n3938 & ~n3939 ) ;
  assign n3943 = ( ~n3266 & n3936 ) | ( ~n3266 & n3942 ) | ( n3936 & n3942 ) ;
  assign n3944 = ( n3935 & n3941 ) | ( n3935 & ~n3943 ) | ( n3941 & ~n3943 ) ;
  assign n3945 = x184 & ~n458 ;
  assign n3946 = n388 | n1507 ;
  assign n3947 = ( ~n382 & n1489 ) | ( ~n382 & n3721 ) | ( n1489 & n3721 ) ;
  assign n3948 = n377 & ~n398 ;
  assign n3949 = n359 | n398 ;
  assign n3950 = ( n3947 & ~n3948 ) | ( n3947 & n3949 ) | ( ~n3948 & n3949 ) ;
  assign n3951 = ~n401 & n3950 ;
  assign n3952 = ( n2218 & ~n3946 ) | ( n2218 & n3951 ) | ( ~n3946 & n3951 ) ;
  assign n3953 = n3945 & ~n3952 ;
  assign n3954 = ( ~n373 & n1776 ) | ( ~n373 & n2719 ) | ( n1776 & n2719 ) ;
  assign n3955 = ( n1497 & ~n1779 ) | ( n1497 & n3954 ) | ( ~n1779 & n3954 ) ;
  assign n3956 = ( ~n2218 & n3946 ) | ( ~n2218 & n3955 ) | ( n3946 & n3955 ) ;
  assign n3957 = n3945 & n3956 ;
  assign n3958 = ( n3944 & n3953 ) | ( n3944 & n3957 ) | ( n3953 & n3957 ) ;
  assign n3959 = x59 | n851 ;
  assign n3960 = ~n444 & n3959 ;
  assign n3961 = ( ~n442 & n453 ) | ( ~n442 & n3960 ) | ( n453 & n3960 ) ;
  assign n3962 = ( n438 & ~n439 ) | ( n438 & n3961 ) | ( ~n439 & n3961 ) ;
  assign n3963 = ( n1793 & ~n2222 ) | ( n1793 & n3962 ) | ( ~n2222 & n3962 ) ;
  assign n3964 = n543 | n2226 ;
  assign n3965 = ( ~n543 & n554 ) | ( ~n543 & n2230 ) | ( n554 & n2230 ) ;
  assign n3966 = ( n3622 & n3964 ) | ( n3622 & ~n3965 ) | ( n3964 & ~n3965 ) ;
  assign n3967 = ( n1804 & ~n3964 ) | ( n1804 & n3965 ) | ( ~n3964 & n3965 ) ;
  assign n3968 = ( n3963 & ~n3966 ) | ( n3963 & n3967 ) | ( ~n3966 & n3967 ) ;
  assign n3969 = ~n584 & n613 ;
  assign n3970 = ( ~n520 & n564 ) | ( ~n520 & n1817 ) | ( n564 & n1817 ) ;
  assign n3971 = ( ~n627 & n3969 ) | ( ~n627 & n3970 ) | ( n3969 & n3970 ) ;
  assign n3972 = ( n627 & n1813 ) | ( n627 & ~n3969 ) | ( n1813 & ~n3969 ) ;
  assign n3973 = ( n3968 & ~n3971 ) | ( n3968 & n3972 ) | ( ~n3971 & n3972 ) ;
  assign n3974 = ( n742 & ~n2265 ) | ( n742 & n3413 ) | ( ~n2265 & n3413 ) ;
  assign n3975 = ~n638 & n2250 ;
  assign n3976 = ( n1575 & ~n2744 ) | ( n1575 & n2753 ) | ( ~n2744 & n2753 ) ;
  assign n3977 = ( n702 & ~n1575 ) | ( n702 & n2860 ) | ( ~n1575 & n2860 ) ;
  assign n3978 = ( n3975 & n3976 ) | ( n3975 & ~n3977 ) | ( n3976 & ~n3977 ) ;
  assign n3979 = ( n3305 & ~n3974 ) | ( n3305 & n3978 ) | ( ~n3974 & n3978 ) ;
  assign n3980 = ( n3405 & ~n3976 ) | ( n3405 & n3977 ) | ( ~n3976 & n3977 ) ;
  assign n3981 = ( ~n3305 & n3974 ) | ( ~n3305 & n3980 ) | ( n3974 & n3980 ) ;
  assign n3982 = ( n3973 & n3979 ) | ( n3973 & ~n3981 ) | ( n3979 & ~n3981 ) ;
  assign n3983 = x185 & ~n863 ;
  assign n3984 = n793 | n1606 ;
  assign n3985 = ( ~n787 & n1588 ) | ( ~n787 & n3759 ) | ( n1588 & n3759 ) ;
  assign n3986 = n782 & ~n803 ;
  assign n3987 = n764 | n803 ;
  assign n3988 = ( n3985 & ~n3986 ) | ( n3985 & n3987 ) | ( ~n3986 & n3987 ) ;
  assign n3989 = ~n806 & n3988 ;
  assign n3990 = ( n2274 & ~n3984 ) | ( n2274 & n3989 ) | ( ~n3984 & n3989 ) ;
  assign n3991 = n3983 & ~n3990 ;
  assign n3992 = ( ~n778 & n1854 ) | ( ~n778 & n2758 ) | ( n1854 & n2758 ) ;
  assign n3993 = ( n1596 & ~n1857 ) | ( n1596 & n3992 ) | ( ~n1857 & n3992 ) ;
  assign n3994 = ( ~n2274 & n3984 ) | ( ~n2274 & n3993 ) | ( n3984 & n3993 ) ;
  assign n3995 = n3983 & n3994 ;
  assign n3996 = ( n3982 & n3991 ) | ( n3982 & n3995 ) | ( n3991 & n3995 ) ;
  assign n3997 = x60 | n1255 ;
  assign n3998 = ~n849 & n3997 ;
  assign n3999 = ( ~n847 & n858 ) | ( ~n847 & n3998 ) | ( n858 & n3998 ) ;
  assign n4000 = ( n843 & ~n844 ) | ( n843 & n3999 ) | ( ~n844 & n3999 ) ;
  assign n4001 = ( n1871 & ~n2278 ) | ( n1871 & n4000 ) | ( ~n2278 & n4000 ) ;
  assign n4002 = n948 | n2282 ;
  assign n4003 = ( ~n948 & n959 ) | ( ~n948 & n2286 ) | ( n959 & n2286 ) ;
  assign n4004 = ( n3660 & n4002 ) | ( n3660 & ~n4003 ) | ( n4002 & ~n4003 ) ;
  assign n4005 = ( n1882 & ~n4002 ) | ( n1882 & n4003 ) | ( ~n4002 & n4003 ) ;
  assign n4006 = ( n4001 & ~n4004 ) | ( n4001 & n4005 ) | ( ~n4004 & n4005 ) ;
  assign n4007 = ~n989 & n1018 ;
  assign n4008 = ( ~n925 & n969 ) | ( ~n925 & n1895 ) | ( n969 & n1895 ) ;
  assign n4009 = ( ~n1032 & n4007 ) | ( ~n1032 & n4008 ) | ( n4007 & n4008 ) ;
  assign n4010 = ( n1032 & n1891 ) | ( n1032 & ~n4007 ) | ( n1891 & ~n4007 ) ;
  assign n4011 = ( n4006 & ~n4009 ) | ( n4006 & n4010 ) | ( ~n4009 & n4010 ) ;
  assign n4012 = ( n1146 & ~n2321 ) | ( n1146 & n3452 ) | ( ~n2321 & n3452 ) ;
  assign n4013 = ~n1043 & n2306 ;
  assign n4014 = ( n1673 & ~n2783 ) | ( n1673 & n2792 ) | ( ~n2783 & n2792 ) ;
  assign n4015 = ( n1106 & ~n1673 ) | ( n1106 & n2897 ) | ( ~n1673 & n2897 ) ;
  assign n4016 = ( n4013 & n4014 ) | ( n4013 & ~n4015 ) | ( n4014 & ~n4015 ) ;
  assign n4017 = ( n3344 & ~n4012 ) | ( n3344 & n4016 ) | ( ~n4012 & n4016 ) ;
  assign n4018 = ( n3444 & ~n4014 ) | ( n3444 & n4015 ) | ( ~n4014 & n4015 ) ;
  assign n4019 = ( ~n3344 & n4012 ) | ( ~n3344 & n4018 ) | ( n4012 & n4018 ) ;
  assign n4020 = ( n4011 & n4017 ) | ( n4011 & ~n4019 ) | ( n4017 & ~n4019 ) ;
  assign n4021 = x186 & ~n1267 ;
  assign n4022 = n1197 | n1704 ;
  assign n4023 = ( ~n1191 & n1686 ) | ( ~n1191 & n3797 ) | ( n1686 & n3797 ) ;
  assign n4024 = n1186 & ~n1207 ;
  assign n4025 = n1168 | n1207 ;
  assign n4026 = ( n4023 & ~n4024 ) | ( n4023 & n4025 ) | ( ~n4024 & n4025 ) ;
  assign n4027 = ~n1210 & n4026 ;
  assign n4028 = ( n2330 & ~n4022 ) | ( n2330 & n4027 ) | ( ~n4022 & n4027 ) ;
  assign n4029 = n4021 & ~n4028 ;
  assign n4030 = ( ~n1182 & n1932 ) | ( ~n1182 & n2797 ) | ( n1932 & n2797 ) ;
  assign n4031 = ( n1694 & ~n1935 ) | ( n1694 & n4030 ) | ( ~n1935 & n4030 ) ;
  assign n4032 = ( ~n2330 & n4022 ) | ( ~n2330 & n4031 ) | ( n4022 & n4031 ) ;
  assign n4033 = n4021 & n4032 ;
  assign n4034 = ( n4020 & n4029 ) | ( n4020 & n4033 ) | ( n4029 & n4033 ) ;
  assign n4035 = x61 | n450 ;
  assign n4036 = ~n1253 & n4035 ;
  assign n4037 = ( ~n1251 & n1262 ) | ( ~n1251 & n4036 ) | ( n1262 & n4036 ) ;
  assign n4038 = ( n1247 & ~n1248 ) | ( n1247 & n4037 ) | ( ~n1248 & n4037 ) ;
  assign n4039 = ( n1949 & ~n2334 ) | ( n1949 & n4038 ) | ( ~n2334 & n4038 ) ;
  assign n4040 = n1352 | n2338 ;
  assign n4041 = ( ~n1352 & n1363 ) | ( ~n1352 & n2342 ) | ( n1363 & n2342 ) ;
  assign n4042 = ( n3698 & n4040 ) | ( n3698 & ~n4041 ) | ( n4040 & ~n4041 ) ;
  assign n4043 = ( n1960 & ~n4040 ) | ( n1960 & n4041 ) | ( ~n4040 & n4041 ) ;
  assign n4044 = ( n4039 & ~n4042 ) | ( n4039 & n4043 ) | ( ~n4042 & n4043 ) ;
  assign n4045 = ~n1393 & n1422 ;
  assign n4046 = ( ~n1329 & n1373 ) | ( ~n1329 & n1973 ) | ( n1373 & n1973 ) ;
  assign n4047 = ( ~n1436 & n4045 ) | ( ~n1436 & n4046 ) | ( n4045 & n4046 ) ;
  assign n4048 = ( n1436 & n1969 ) | ( n1436 & ~n4045 ) | ( n1969 & ~n4045 ) ;
  assign n4049 = ( n4044 & ~n4047 ) | ( n4044 & n4048 ) | ( ~n4047 & n4048 ) ;
  assign n4050 = ( n341 & ~n2377 ) | ( n341 & n3491 ) | ( ~n2377 & n3491 ) ;
  assign n4051 = ~n1447 & n2362 ;
  assign n4052 = ( n293 & ~n2822 ) | ( n293 & n2830 ) | ( ~n2822 & n2830 ) ;
  assign n4053 = ( n289 & ~n293 ) | ( n289 & n2934 ) | ( ~n293 & n2934 ) ;
  assign n4054 = ( n4051 & n4052 ) | ( n4051 & ~n4053 ) | ( n4052 & ~n4053 ) ;
  assign n4055 = ( n3383 & ~n4050 ) | ( n3383 & n4054 ) | ( ~n4050 & n4054 ) ;
  assign n4056 = ( n3483 & ~n4052 ) | ( n3483 & n4053 ) | ( ~n4052 & n4053 ) ;
  assign n4057 = ( ~n3383 & n4050 ) | ( ~n3383 & n4056 ) | ( n4050 & n4056 ) ;
  assign n4058 = ( n4049 & n4055 ) | ( n4049 & ~n4057 ) | ( n4055 & ~n4057 ) ;
  assign n4059 = x187 & ~n443 ;
  assign n4060 = n448 | n1790 ;
  assign n4061 = ( ~n376 & n1774 ) | ( ~n376 & n3835 ) | ( n1774 & n3835 ) ;
  assign n4062 = ~n408 & n1497 ;
  assign n4063 = n402 | n408 ;
  assign n4064 = ( n4061 & ~n4062 ) | ( n4061 & n4063 ) | ( ~n4062 & n4063 ) ;
  assign n4065 = ~n405 & n4064 ;
  assign n4066 = ( n2386 & ~n4060 ) | ( n2386 & n4065 ) | ( ~n4060 & n4065 ) ;
  assign n4067 = n4059 & ~n4066 ;
  assign n4068 = ( n384 & ~n410 ) | ( n384 & n1781 ) | ( ~n410 & n1781 ) ;
  assign n4069 = ( ~n2386 & n4060 ) | ( ~n2386 & n4068 ) | ( n4060 & n4068 ) ;
  assign n4070 = n4059 & n4069 ;
  assign n4071 = ( n4058 & n4067 ) | ( n4058 & n4070 ) | ( n4067 & n4070 ) ;
  assign n4072 = x62 | n855 ;
  assign n4073 = ~n441 & n4072 ;
  assign n4074 = ( ~n433 & n437 ) | ( ~n433 & n4073 ) | ( n437 & n4073 ) ;
  assign n4075 = ( n1510 & ~n1511 ) | ( n1510 & n4074 ) | ( ~n1511 & n4074 ) ;
  assign n4076 = ( ~n514 & n2020 ) | ( ~n514 & n4075 ) | ( n2020 & n4075 ) ;
  assign n4077 = n534 | n569 ;
  assign n4078 = ( ~n534 & n538 ) | ( ~n534 & n555 ) | ( n538 & n555 ) ;
  assign n4079 = ( n3736 & n4077 ) | ( n3736 & ~n4078 ) | ( n4077 & ~n4078 ) ;
  assign n4080 = ( n2034 & ~n4077 ) | ( n2034 & n4078 ) | ( ~n4077 & n4078 ) ;
  assign n4081 = ( n4076 & ~n4079 ) | ( n4076 & n4080 ) | ( ~n4079 & n4080 ) ;
  assign n4082 = ~n578 & n1544 ;
  assign n4083 = ( ~n603 & n604 ) | ( ~n603 & n2044 ) | ( n604 & n2044 ) ;
  assign n4084 = ( ~n1554 & n4082 ) | ( ~n1554 & n4083 ) | ( n4082 & n4083 ) ;
  assign n4085 = ( n1554 & n2040 ) | ( n1554 & ~n4082 ) | ( n2040 & ~n4082 ) ;
  assign n4086 = ( n4081 & ~n4084 ) | ( n4081 & n4085 ) | ( ~n4084 & n4085 ) ;
  assign n4087 = ( n746 & ~n2421 ) | ( n746 & n3529 ) | ( ~n2421 & n3529 ) ;
  assign n4088 = ~n1561 & n2406 ;
  assign n4089 = ( n698 & ~n2859 ) | ( n698 & n2867 ) | ( ~n2859 & n2867 ) ;
  assign n4090 = ( n694 & ~n698 ) | ( n694 & n2969 ) | ( ~n698 & n2969 ) ;
  assign n4091 = ( n4088 & n4089 ) | ( n4088 & ~n4090 ) | ( n4089 & ~n4090 ) ;
  assign n4092 = ( n3422 & ~n4087 ) | ( n3422 & n4091 ) | ( ~n4087 & n4091 ) ;
  assign n4093 = ( n3521 & ~n4089 ) | ( n3521 & n4090 ) | ( ~n4089 & n4090 ) ;
  assign n4094 = ( ~n3422 & n4087 ) | ( ~n3422 & n4093 ) | ( n4087 & n4093 ) ;
  assign n4095 = ( n4086 & n4092 ) | ( n4086 & ~n4094 ) | ( n4092 & ~n4094 ) ;
  assign n4096 = x188 & ~n848 ;
  assign n4097 = n853 | n1868 ;
  assign n4098 = ( ~n781 & n1852 ) | ( ~n781 & n3873 ) | ( n1852 & n3873 ) ;
  assign n4099 = ~n813 & n1596 ;
  assign n4100 = n807 | n813 ;
  assign n4101 = ( n4098 & ~n4099 ) | ( n4098 & n4100 ) | ( ~n4099 & n4100 ) ;
  assign n4102 = ~n810 & n4101 ;
  assign n4103 = ( n2430 & ~n4097 ) | ( n2430 & n4102 ) | ( ~n4097 & n4102 ) ;
  assign n4104 = n4096 & ~n4103 ;
  assign n4105 = ( n789 & ~n815 ) | ( n789 & n1859 ) | ( ~n815 & n1859 ) ;
  assign n4106 = ( ~n2430 & n4097 ) | ( ~n2430 & n4105 ) | ( n4097 & n4105 ) ;
  assign n4107 = n4096 & n4106 ;
  assign n4108 = ( n4095 & n4104 ) | ( n4095 & n4107 ) | ( n4104 & n4107 ) ;
  assign n4109 = x63 | n1259 ;
  assign n4110 = ~n846 & n4109 ;
  assign n4111 = ( ~n838 & n842 ) | ( ~n838 & n4110 ) | ( n842 & n4110 ) ;
  assign n4112 = ( n1609 & ~n1610 ) | ( n1609 & n4111 ) | ( ~n1610 & n4111 ) ;
  assign n4113 = ( ~n919 & n2090 ) | ( ~n919 & n4112 ) | ( n2090 & n4112 ) ;
  assign n4114 = n939 | n974 ;
  assign n4115 = ( ~n939 & n943 ) | ( ~n939 & n960 ) | ( n943 & n960 ) ;
  assign n4116 = ( n3774 & n4114 ) | ( n3774 & ~n4115 ) | ( n4114 & ~n4115 ) ;
  assign n4117 = ( n2104 & ~n4114 ) | ( n2104 & n4115 ) | ( ~n4114 & n4115 ) ;
  assign n4118 = ( n4113 & ~n4116 ) | ( n4113 & n4117 ) | ( ~n4116 & n4117 ) ;
  assign n4119 = ~n983 & n1643 ;
  assign n4120 = ( ~n1008 & n1009 ) | ( ~n1008 & n2114 ) | ( n1009 & n2114 ) ;
  assign n4121 = ( ~n1653 & n4119 ) | ( ~n1653 & n4120 ) | ( n4119 & n4120 ) ;
  assign n4122 = ( n1653 & n2110 ) | ( n1653 & ~n4119 ) | ( n2110 & ~n4119 ) ;
  assign n4123 = ( n4118 & ~n4121 ) | ( n4118 & n4122 ) | ( ~n4121 & n4122 ) ;
  assign n4124 = ( n1150 & ~n2465 ) | ( n1150 & n3567 ) | ( ~n2465 & n3567 ) ;
  assign n4125 = ~n1660 & n2450 ;
  assign n4126 = ( n1102 & ~n2896 ) | ( n1102 & n2904 ) | ( ~n2896 & n2904 ) ;
  assign n4127 = ( n1098 & ~n1102 ) | ( n1098 & n3005 ) | ( ~n1102 & n3005 ) ;
  assign n4128 = ( n4125 & n4126 ) | ( n4125 & ~n4127 ) | ( n4126 & ~n4127 ) ;
  assign n4129 = ( n3461 & ~n4124 ) | ( n3461 & n4128 ) | ( ~n4124 & n4128 ) ;
  assign n4130 = ( n3559 & ~n4126 ) | ( n3559 & n4127 ) | ( ~n4126 & n4127 ) ;
  assign n4131 = ( ~n3461 & n4124 ) | ( ~n3461 & n4130 ) | ( n4124 & n4130 ) ;
  assign n4132 = ( n4123 & n4129 ) | ( n4123 & ~n4131 ) | ( n4129 & ~n4131 ) ;
  assign n4133 = x189 & ~n1252 ;
  assign n4134 = n1257 | n1946 ;
  assign n4135 = ( ~n1185 & n1930 ) | ( ~n1185 & n3911 ) | ( n1930 & n3911 ) ;
  assign n4136 = ~n1217 & n1694 ;
  assign n4137 = n1211 | n1217 ;
  assign n4138 = ( n4135 & ~n4136 ) | ( n4135 & n4137 ) | ( ~n4136 & n4137 ) ;
  assign n4139 = ~n1214 & n4138 ;
  assign n4140 = ( n2474 & ~n4134 ) | ( n2474 & n4139 ) | ( ~n4134 & n4139 ) ;
  assign n4141 = n4133 & ~n4140 ;
  assign n4142 = ( n1193 & ~n1219 ) | ( n1193 & n1937 ) | ( ~n1219 & n1937 ) ;
  assign n4143 = ( ~n2474 & n4134 ) | ( ~n2474 & n4142 ) | ( n4134 & n4142 ) ;
  assign n4144 = n4133 & n4143 ;
  assign n4145 = ( n4132 & n4141 ) | ( n4132 & n4144 ) | ( n4141 & n4144 ) ;
  assign n4146 = x64 | n434 ;
  assign n4147 = ~n1250 & n4146 ;
  assign n4148 = ( ~n1242 & n1246 ) | ( ~n1242 & n4147 ) | ( n1246 & n4147 ) ;
  assign n4149 = ( n1707 & ~n1708 ) | ( n1707 & n4148 ) | ( ~n1708 & n4148 ) ;
  assign n4150 = ( ~n1323 & n2160 ) | ( ~n1323 & n4149 ) | ( n2160 & n4149 ) ;
  assign n4151 = n1343 | n1378 ;
  assign n4152 = ( ~n1343 & n1347 ) | ( ~n1343 & n1364 ) | ( n1347 & n1364 ) ;
  assign n4153 = ( n3812 & n4151 ) | ( n3812 & ~n4152 ) | ( n4151 & ~n4152 ) ;
  assign n4154 = ( n2174 & ~n4151 ) | ( n2174 & n4152 ) | ( ~n4151 & n4152 ) ;
  assign n4155 = ( n4150 & ~n4153 ) | ( n4150 & n4154 ) | ( ~n4153 & n4154 ) ;
  assign n4156 = ~n1387 & n1741 ;
  assign n4157 = ( ~n1412 & n1413 ) | ( ~n1412 & n2184 ) | ( n1413 & n2184 ) ;
  assign n4158 = ( ~n1751 & n4156 ) | ( ~n1751 & n4157 ) | ( n4156 & n4157 ) ;
  assign n4159 = ( n1751 & n2180 ) | ( n1751 & ~n4156 ) | ( n2180 & ~n4156 ) ;
  assign n4160 = ( n4155 & ~n4158 ) | ( n4155 & n4159 ) | ( ~n4158 & n4159 ) ;
  assign n4161 = ( n1488 & ~n2509 ) | ( n1488 & n3605 ) | ( ~n2509 & n3605 ) ;
  assign n4162 = ~n1755 & n2494 ;
  assign n4163 = ( n1479 & ~n2933 ) | ( n1479 & n2941 ) | ( ~n2933 & n2941 ) ;
  assign n4164 = ( n307 & ~n1479 ) | ( n307 & n3042 ) | ( ~n1479 & n3042 ) ;
  assign n4165 = ( n4162 & n4163 ) | ( n4162 & ~n4164 ) | ( n4163 & ~n4164 ) ;
  assign n4166 = ( n3499 & ~n4161 ) | ( n3499 & n4165 ) | ( ~n4161 & n4165 ) ;
  assign n4167 = ( n3597 & ~n4163 ) | ( n3597 & n4164 ) | ( ~n4163 & n4164 ) ;
  assign n4168 = ( ~n3499 & n4161 ) | ( ~n3499 & n4167 ) | ( n4161 & n4167 ) ;
  assign n4169 = ( n4160 & n4166 ) | ( n4160 & ~n4168 ) | ( n4166 & ~n4168 ) ;
  assign n4170 = x190 & ~n440 ;
  assign n4171 = n452 | n2017 ;
  assign n4172 = ( n374 & ~n1496 ) | ( n374 & n3949 ) | ( ~n1496 & n3949 ) ;
  assign n4173 = ~n413 & n1781 ;
  assign n4174 = n409 | n413 ;
  assign n4175 = ( n4172 & ~n4173 ) | ( n4172 & n4174 ) | ( ~n4173 & n4174 ) ;
  assign n4176 = ~n394 & n4175 ;
  assign n4177 = ( n2518 & ~n4171 ) | ( n2518 & n4176 ) | ( ~n4171 & n4176 ) ;
  assign n4178 = n4170 & ~n4177 ;
  assign n4179 = ( n1499 & ~n1502 ) | ( n1499 & n2008 ) | ( ~n1502 & n2008 ) ;
  assign n4180 = ( ~n2518 & n4171 ) | ( ~n2518 & n4179 ) | ( n4171 & n4179 ) ;
  assign n4181 = n4170 & n4180 ;
  assign n4182 = ( n4169 & n4178 ) | ( n4169 & n4181 ) | ( n4178 & n4181 ) ;
  assign n4183 = x65 | n839 ;
  assign n4184 = ~n432 & n4183 ;
  assign n4185 = ( ~n427 & n457 ) | ( ~n427 & n4184 ) | ( n457 & n4184 ) ;
  assign n4186 = ( ~n512 & n1793 ) | ( ~n512 & n4185 ) | ( n1793 & n4185 ) ;
  assign n4187 = ( n486 & ~n1526 ) | ( n486 & n4186 ) | ( ~n1526 & n4186 ) ;
  assign n4188 = n559 | n1538 ;
  assign n4189 = ( ~n559 & n566 ) | ( ~n559 & n1533 ) | ( n566 & n1533 ) ;
  assign n4190 = ( n3850 & n4188 ) | ( n3850 & ~n4189 ) | ( n4188 & ~n4189 ) ;
  assign n4191 = ( n2230 & ~n4188 ) | ( n2230 & n4189 ) | ( ~n4188 & n4189 ) ;
  assign n4192 = ( n4187 & ~n4190 ) | ( n4187 & n4191 ) | ( ~n4190 & n4191 ) ;
  assign n4193 = ~n619 & n1822 ;
  assign n4194 = ( ~n607 & n611 ) | ( ~n607 & n2238 ) | ( n611 & n2238 ) ;
  assign n4195 = ( ~n1830 & n4193 ) | ( ~n1830 & n4194 ) | ( n4193 & n4194 ) ;
  assign n4196 = ( n1830 & n2235 ) | ( n1830 & ~n4193 ) | ( n2235 & ~n4193 ) ;
  assign n4197 = ( n4192 & ~n4195 ) | ( n4192 & n4196 ) | ( ~n4195 & n4196 ) ;
  assign n4198 = ( n1587 & ~n2546 ) | ( n1587 & n3643 ) | ( ~n2546 & n3643 ) ;
  assign n4199 = ~n1833 & n2531 ;
  assign n4200 = ( n1578 & ~n2970 ) | ( n1578 & n2977 ) | ( ~n2970 & n2977 ) ;
  assign n4201 = ( n712 & ~n1578 ) | ( n712 & n3077 ) | ( ~n1578 & n3077 ) ;
  assign n4202 = ( n4199 & n4200 ) | ( n4199 & ~n4201 ) | ( n4200 & ~n4201 ) ;
  assign n4203 = ( n3537 & ~n4198 ) | ( n3537 & n4202 ) | ( ~n4198 & n4202 ) ;
  assign n4204 = ( n3635 & ~n4200 ) | ( n3635 & n4201 ) | ( ~n4200 & n4201 ) ;
  assign n4205 = ( ~n3537 & n4198 ) | ( ~n3537 & n4204 ) | ( n4198 & n4204 ) ;
  assign n4206 = ( n4197 & n4203 ) | ( n4197 & ~n4205 ) | ( n4203 & ~n4205 ) ;
  assign n4207 = x191 & ~n845 ;
  assign n4208 = n857 | n2087 ;
  assign n4209 = ( n779 & ~n1595 ) | ( n779 & n3987 ) | ( ~n1595 & n3987 ) ;
  assign n4210 = ~n818 & n1859 ;
  assign n4211 = n814 | n818 ;
  assign n4212 = ( n4209 & ~n4210 ) | ( n4209 & n4211 ) | ( ~n4210 & n4211 ) ;
  assign n4213 = ~n799 & n4212 ;
  assign n4214 = ( n2555 & ~n4208 ) | ( n2555 & n4213 ) | ( ~n4208 & n4213 ) ;
  assign n4215 = n4207 & ~n4214 ;
  assign n4216 = ( n1598 & ~n1601 ) | ( n1598 & n2078 ) | ( ~n1601 & n2078 ) ;
  assign n4217 = ( ~n2555 & n4208 ) | ( ~n2555 & n4216 ) | ( n4208 & n4216 ) ;
  assign n4218 = n4207 & n4217 ;
  assign n4219 = ( n4206 & n4215 ) | ( n4206 & n4218 ) | ( n4215 & n4218 ) ;
  assign n4220 = x66 | n1243 ;
  assign n4221 = ~n837 & n4220 ;
  assign n4222 = ( ~n832 & n862 ) | ( ~n832 & n4221 ) | ( n862 & n4221 ) ;
  assign n4223 = ( ~n917 & n1871 ) | ( ~n917 & n4222 ) | ( n1871 & n4222 ) ;
  assign n4224 = ( n891 & ~n1625 ) | ( n891 & n4223 ) | ( ~n1625 & n4223 ) ;
  assign n4225 = n964 | n1637 ;
  assign n4226 = ( ~n964 & n971 ) | ( ~n964 & n1632 ) | ( n971 & n1632 ) ;
  assign n4227 = ( n3888 & n4225 ) | ( n3888 & ~n4226 ) | ( n4225 & ~n4226 ) ;
  assign n4228 = ( n2286 & ~n4225 ) | ( n2286 & n4226 ) | ( ~n4225 & n4226 ) ;
  assign n4229 = ( n4224 & ~n4227 ) | ( n4224 & n4228 ) | ( ~n4227 & n4228 ) ;
  assign n4230 = ~n1024 & n1900 ;
  assign n4231 = ( ~n1012 & n1016 ) | ( ~n1012 & n2294 ) | ( n1016 & n2294 ) ;
  assign n4232 = ( ~n1908 & n4230 ) | ( ~n1908 & n4231 ) | ( n4230 & n4231 ) ;
  assign n4233 = ( n1908 & n2291 ) | ( n1908 & ~n4230 ) | ( n2291 & ~n4230 ) ;
  assign n4234 = ( n4229 & ~n4232 ) | ( n4229 & n4233 ) | ( ~n4232 & n4233 ) ;
  assign n4235 = ( n1685 & ~n2583 ) | ( n1685 & n3681 ) | ( ~n2583 & n3681 ) ;
  assign n4236 = ~n1911 & n2568 ;
  assign n4237 = ( n1676 & ~n3006 ) | ( n1676 & n3013 ) | ( ~n3006 & n3013 ) ;
  assign n4238 = ( n1116 & ~n1676 ) | ( n1116 & n3113 ) | ( ~n1676 & n3113 ) ;
  assign n4239 = ( n4236 & n4237 ) | ( n4236 & ~n4238 ) | ( n4237 & ~n4238 ) ;
  assign n4240 = ( n3575 & ~n4235 ) | ( n3575 & n4239 ) | ( ~n4235 & n4239 ) ;
  assign n4241 = ( n3673 & ~n4237 ) | ( n3673 & n4238 ) | ( ~n4237 & n4238 ) ;
  assign n4242 = ( ~n3575 & n4235 ) | ( ~n3575 & n4241 ) | ( n4235 & n4241 ) ;
  assign n4243 = ( n4234 & n4240 ) | ( n4234 & ~n4242 ) | ( n4240 & ~n4242 ) ;
  assign n4244 = x192 & ~n1249 ;
  assign n4245 = n1261 | n2157 ;
  assign n4246 = ( n1183 & ~n1693 ) | ( n1183 & n4025 ) | ( ~n1693 & n4025 ) ;
  assign n4247 = ~n1222 & n1937 ;
  assign n4248 = n1218 | n1222 ;
  assign n4249 = ( n4246 & ~n4247 ) | ( n4246 & n4248 ) | ( ~n4247 & n4248 ) ;
  assign n4250 = ~n1203 & n4249 ;
  assign n4251 = ( n2592 & ~n4245 ) | ( n2592 & n4250 ) | ( ~n4245 & n4250 ) ;
  assign n4252 = n4244 & ~n4251 ;
  assign n4253 = ( n1696 & ~n1699 ) | ( n1696 & n2148 ) | ( ~n1699 & n2148 ) ;
  assign n4254 = ( ~n2592 & n4245 ) | ( ~n2592 & n4253 ) | ( n4245 & n4253 ) ;
  assign n4255 = n4244 & n4254 ;
  assign n4256 = ( n4243 & n4252 ) | ( n4243 & n4255 ) | ( n4252 & n4255 ) ;
  assign n4257 = x67 | n428 ;
  assign n4258 = ~n1241 & n4257 ;
  assign n4259 = ( ~n1236 & n1266 ) | ( ~n1236 & n4258 ) | ( n1266 & n4258 ) ;
  assign n4260 = ( ~n1321 & n1949 ) | ( ~n1321 & n4259 ) | ( n1949 & n4259 ) ;
  assign n4261 = ( n1295 & ~n1723 ) | ( n1295 & n4260 ) | ( ~n1723 & n4260 ) ;
  assign n4262 = n1368 | n1735 ;
  assign n4263 = ( ~n1368 & n1375 ) | ( ~n1368 & n1730 ) | ( n1375 & n1730 ) ;
  assign n4264 = ( n3926 & n4262 ) | ( n3926 & ~n4263 ) | ( n4262 & ~n4263 ) ;
  assign n4265 = ( n2342 & ~n4262 ) | ( n2342 & n4263 ) | ( ~n4262 & n4263 ) ;
  assign n4266 = ( n4261 & ~n4264 ) | ( n4261 & n4265 ) | ( ~n4264 & n4265 ) ;
  assign n4267 = ~n1428 & n1978 ;
  assign n4268 = ( ~n1416 & n1420 ) | ( ~n1416 & n2350 ) | ( n1420 & n2350 ) ;
  assign n4269 = ( ~n1986 & n4267 ) | ( ~n1986 & n4268 ) | ( n4267 & n4268 ) ;
  assign n4270 = ( n1986 & n2347 ) | ( n1986 & ~n4267 ) | ( n2347 & ~n4267 ) ;
  assign n4271 = ( n4266 & ~n4269 ) | ( n4266 & n4270 ) | ( ~n4269 & n4270 ) ;
  assign n4272 = ( n369 & ~n2618 ) | ( n369 & n3719 ) | ( ~n2618 & n3719 ) ;
  assign n4273 = ~n265 & n2604 ;
  assign n4274 = ( n321 & ~n3043 ) | ( n321 & n3049 ) | ( ~n3043 & n3049 ) ;
  assign n4275 = ( n317 & ~n321 ) | ( n317 & n3149 ) | ( ~n321 & n3149 ) ;
  assign n4276 = ( n4273 & n4274 ) | ( n4273 & ~n4275 ) | ( n4274 & ~n4275 ) ;
  assign n4277 = ( n3613 & ~n4272 ) | ( n3613 & n4276 ) | ( ~n4272 & n4276 ) ;
  assign n4278 = ( n3711 & ~n4274 ) | ( n3711 & n4275 ) | ( ~n4274 & n4275 ) ;
  assign n4279 = ( ~n3613 & n4272 ) | ( ~n3613 & n4278 ) | ( n4272 & n4278 ) ;
  assign n4280 = ( n4271 & n4277 ) | ( n4271 & ~n4279 ) | ( n4277 & ~n4279 ) ;
  assign n4281 = x193 & ~n431 ;
  assign n4282 = n436 | n454 ;
  assign n4283 = ( ~n420 & n1494 ) | ( ~n420 & n4063 ) | ( n1494 & n4063 ) ;
  assign n4284 = ~n391 & n2008 ;
  assign n4285 = ( n415 & n4283 ) | ( n415 & ~n4284 ) | ( n4283 & ~n4284 ) ;
  assign n4286 = ~n388 & n4285 ;
  assign n4287 = ( n2627 & ~n4282 ) | ( n2627 & n4286 ) | ( ~n4282 & n4286 ) ;
  assign n4288 = n4281 & ~n4287 ;
  assign n4289 = ( n418 & n1783 ) | ( n418 & ~n1785 ) | ( n1783 & ~n1785 ) ;
  assign n4290 = ( ~n2627 & n4282 ) | ( ~n2627 & n4289 ) | ( n4282 & n4289 ) ;
  assign n4291 = n4281 & n4290 ;
  assign n4292 = ( n4280 & n4288 ) | ( n4280 & n4291 ) | ( n4288 & n4291 ) ;
  assign n4293 = x68 | n833 ;
  assign n4294 = ~n426 & n4293 ;
  assign n4295 = ( ~n493 & n497 ) | ( ~n493 & n4294 ) | ( n497 & n4294 ) ;
  assign n4296 = ( ~n513 & n2020 ) | ( ~n513 & n4295 ) | ( n2020 & n4295 ) ;
  assign n4297 = ( n1520 & ~n1807 ) | ( n1520 & n4296 ) | ( ~n1807 & n4296 ) ;
  assign n4298 = n523 | n1817 ;
  assign n4299 = ( ~n523 & n527 ) | ( ~n523 & n1812 ) | ( n527 & n1812 ) ;
  assign n4300 = ( n3964 & n4298 ) | ( n3964 & ~n4299 ) | ( n4298 & ~n4299 ) ;
  assign n4301 = ( n555 & ~n4298 ) | ( n555 & n4299 ) | ( ~n4298 & n4299 ) ;
  assign n4302 = ( n4297 & ~n4300 ) | ( n4297 & n4301 ) | ( ~n4300 & n4301 ) ;
  assign n4303 = ~n644 & n2049 ;
  assign n4304 = ( n2056 & n2394 ) | ( n2056 & ~n4303 ) | ( n2394 & ~n4303 ) ;
  assign n4305 = ( ~n594 & n595 ) | ( ~n594 & n612 ) | ( n595 & n612 ) ;
  assign n4306 = ( ~n2056 & n4303 ) | ( ~n2056 & n4305 ) | ( n4303 & n4305 ) ;
  assign n4307 = ( n4302 & n4304 ) | ( n4302 & ~n4306 ) | ( n4304 & ~n4306 ) ;
  assign n4308 = ( n774 & ~n2653 ) | ( n774 & n3757 ) | ( ~n2653 & n3757 ) ;
  assign n4309 = ~n670 & n2639 ;
  assign n4310 = ( n726 & ~n3079 ) | ( n726 & n3085 ) | ( ~n3079 & n3085 ) ;
  assign n4311 = ( n722 & ~n726 ) | ( n722 & n3185 ) | ( ~n726 & n3185 ) ;
  assign n4312 = ( n4309 & n4310 ) | ( n4309 & ~n4311 ) | ( n4310 & ~n4311 ) ;
  assign n4313 = ( n3651 & ~n4308 ) | ( n3651 & n4312 ) | ( ~n4308 & n4312 ) ;
  assign n4314 = ( n3749 & ~n4310 ) | ( n3749 & n4311 ) | ( ~n4310 & n4311 ) ;
  assign n4315 = ( ~n3651 & n4308 ) | ( ~n3651 & n4314 ) | ( n4308 & n4314 ) ;
  assign n4316 = ( n4307 & n4313 ) | ( n4307 & ~n4315 ) | ( n4313 & ~n4315 ) ;
  assign n4317 = x194 & ~n836 ;
  assign n4318 = n841 | n859 ;
  assign n4319 = ( ~n825 & n1593 ) | ( ~n825 & n4100 ) | ( n1593 & n4100 ) ;
  assign n4320 = ~n796 & n2078 ;
  assign n4321 = ( n820 & n4319 ) | ( n820 & ~n4320 ) | ( n4319 & ~n4320 ) ;
  assign n4322 = ~n793 & n4321 ;
  assign n4323 = ( n2662 & ~n4318 ) | ( n2662 & n4322 ) | ( ~n4318 & n4322 ) ;
  assign n4324 = n4317 & ~n4323 ;
  assign n4325 = ( n823 & n1861 ) | ( n823 & ~n1863 ) | ( n1861 & ~n1863 ) ;
  assign n4326 = ( ~n2662 & n4318 ) | ( ~n2662 & n4325 ) | ( n4318 & n4325 ) ;
  assign n4327 = n4317 & n4326 ;
  assign n4328 = ( n4316 & n4324 ) | ( n4316 & n4327 ) | ( n4324 & n4327 ) ;
  assign n4329 = x69 | n1237 ;
  assign n4330 = ~n831 & n4329 ;
  assign n4331 = ( ~n898 & n902 ) | ( ~n898 & n4330 ) | ( n902 & n4330 ) ;
  assign n4332 = ( ~n918 & n2090 ) | ( ~n918 & n4331 ) | ( n2090 & n4331 ) ;
  assign n4333 = ( n1619 & ~n1885 ) | ( n1619 & n4332 ) | ( ~n1885 & n4332 ) ;
  assign n4334 = n928 | n1895 ;
  assign n4335 = ( ~n928 & n932 ) | ( ~n928 & n1890 ) | ( n932 & n1890 ) ;
  assign n4336 = ( n4002 & n4334 ) | ( n4002 & ~n4335 ) | ( n4334 & ~n4335 ) ;
  assign n4337 = ( n960 & ~n4334 ) | ( n960 & n4335 ) | ( ~n4334 & n4335 ) ;
  assign n4338 = ( n4333 & ~n4336 ) | ( n4333 & n4337 ) | ( ~n4336 & n4337 ) ;
  assign n4339 = ~n1049 & n2119 ;
  assign n4340 = ( n2126 & n2438 ) | ( n2126 & ~n4339 ) | ( n2438 & ~n4339 ) ;
  assign n4341 = ( ~n999 & n1000 ) | ( ~n999 & n1017 ) | ( n1000 & n1017 ) ;
  assign n4342 = ( ~n2126 & n4339 ) | ( ~n2126 & n4341 ) | ( n4339 & n4341 ) ;
  assign n4343 = ( n4338 & n4340 ) | ( n4338 & ~n4342 ) | ( n4340 & ~n4342 ) ;
  assign n4344 = ( n1178 & ~n2688 ) | ( n1178 & n3795 ) | ( ~n2688 & n3795 ) ;
  assign n4345 = ~n1074 & n2674 ;
  assign n4346 = ( n1130 & ~n3115 ) | ( n1130 & n3121 ) | ( ~n3115 & n3121 ) ;
  assign n4347 = ( n1126 & ~n1130 ) | ( n1126 & n3221 ) | ( ~n1130 & n3221 ) ;
  assign n4348 = ( n4345 & n4346 ) | ( n4345 & ~n4347 ) | ( n4346 & ~n4347 ) ;
  assign n4349 = ( n3689 & ~n4344 ) | ( n3689 & n4348 ) | ( ~n4344 & n4348 ) ;
  assign n4350 = ( n3787 & ~n4346 ) | ( n3787 & n4347 ) | ( ~n4346 & n4347 ) ;
  assign n4351 = ( ~n3689 & n4344 ) | ( ~n3689 & n4350 ) | ( n4344 & n4350 ) ;
  assign n4352 = ( n4343 & n4349 ) | ( n4343 & ~n4351 ) | ( n4349 & ~n4351 ) ;
  assign n4353 = x195 & ~n1240 ;
  assign n4354 = n1245 | n1263 ;
  assign n4355 = ( ~n1229 & n1691 ) | ( ~n1229 & n4137 ) | ( n1691 & n4137 ) ;
  assign n4356 = ~n1200 & n2148 ;
  assign n4357 = ( n1224 & n4355 ) | ( n1224 & ~n4356 ) | ( n4355 & ~n4356 ) ;
  assign n4358 = ~n1197 & n4357 ;
  assign n4359 = ( n2697 & ~n4354 ) | ( n2697 & n4358 ) | ( ~n4354 & n4358 ) ;
  assign n4360 = n4353 & ~n4359 ;
  assign n4361 = ( n1227 & n1939 ) | ( n1227 & ~n1941 ) | ( n1939 & ~n1941 ) ;
  assign n4362 = ( ~n2697 & n4354 ) | ( ~n2697 & n4361 ) | ( n4354 & n4361 ) ;
  assign n4363 = n4353 & n4362 ;
  assign n4364 = ( n4352 & n4360 ) | ( n4352 & n4363 ) | ( n4360 & n4363 ) ;
  assign n4365 = x70 | n494 ;
  assign n4366 = ~n1235 & n4365 ;
  assign n4367 = ( ~n1302 & n1306 ) | ( ~n1302 & n4366 ) | ( n1306 & n4366 ) ;
  assign n4368 = ( ~n1322 & n2160 ) | ( ~n1322 & n4367 ) | ( n2160 & n4367 ) ;
  assign n4369 = ( n1717 & ~n1963 ) | ( n1717 & n4368 ) | ( ~n1963 & n4368 ) ;
  assign n4370 = n1332 | n1973 ;
  assign n4371 = ( ~n1332 & n1336 ) | ( ~n1332 & n1968 ) | ( n1336 & n1968 ) ;
  assign n4372 = ( n4040 & n4370 ) | ( n4040 & ~n4371 ) | ( n4370 & ~n4371 ) ;
  assign n4373 = ( n1364 & ~n4370 ) | ( n1364 & n4371 ) | ( ~n4370 & n4371 ) ;
  assign n4374 = ( n4369 & ~n4372 ) | ( n4369 & n4373 ) | ( ~n4372 & n4373 ) ;
  assign n4375 = ~n1453 & n2189 ;
  assign n4376 = ( n2196 & n2482 ) | ( n2196 & ~n4375 ) | ( n2482 & ~n4375 ) ;
  assign n4377 = ( ~n1403 & n1404 ) | ( ~n1403 & n1421 ) | ( n1404 & n1421 ) ;
  assign n4378 = ( ~n2196 & n4375 ) | ( ~n2196 & n4377 ) | ( n4375 & n4377 ) ;
  assign n4379 = ( n4374 & n4376 ) | ( n4374 & ~n4378 ) | ( n4376 & ~n4378 ) ;
  assign n4380 = ( n373 & ~n2719 ) | ( n373 & n3833 ) | ( ~n2719 & n3833 ) ;
  assign n4381 = ~n273 & n2709 ;
  assign n4382 = ( n322 & ~n3151 ) | ( n322 & n3157 ) | ( ~n3151 & n3157 ) ;
  assign n4383 = ( n304 & ~n322 ) | ( n304 & n3257 ) | ( ~n322 & n3257 ) ;
  assign n4384 = ( n4381 & n4382 ) | ( n4381 & ~n4383 ) | ( n4382 & ~n4383 ) ;
  assign n4385 = ( n3727 & ~n4380 ) | ( n3727 & n4384 ) | ( ~n4380 & n4384 ) ;
  assign n4386 = ( n3825 & ~n4382 ) | ( n3825 & n4383 ) | ( ~n4382 & n4383 ) ;
  assign n4387 = ( ~n3727 & n4380 ) | ( ~n3727 & n4386 ) | ( n4380 & n4386 ) ;
  assign n4388 = ( n4379 & n4385 ) | ( n4379 & ~n4387 ) | ( n4385 & ~n4387 ) ;
  assign n4389 = x196 & ~n425 ;
  assign n4390 = n430 | n1512 ;
  assign n4391 = ( ~n421 & n1779 ) | ( ~n421 & n4174 ) | ( n1779 & n4174 ) ;
  assign n4392 = n418 & ~n460 ;
  assign n4393 = ( n1503 & n4391 ) | ( n1503 & ~n4392 ) | ( n4391 & ~n4392 ) ;
  assign n4394 = ~n448 & n4393 ;
  assign n4395 = ( n2731 & ~n4390 ) | ( n2731 & n4394 ) | ( ~n4390 & n4394 ) ;
  assign n4396 = n4389 & ~n4395 ;
  assign n4397 = ( n1506 & n2010 ) | ( n1506 & ~n2012 ) | ( n2010 & ~n2012 ) ;
  assign n4398 = ( ~n2731 & n4390 ) | ( ~n2731 & n4397 ) | ( n4390 & n4397 ) ;
  assign n4399 = n4389 & n4398 ;
  assign n4400 = ( n4388 & n4396 ) | ( n4388 & n4399 ) | ( n4396 & n4399 ) ;
  assign n4401 = x71 | n899 ;
  assign n4402 = ~n492 & n4401 ;
  assign n4403 = ( ~n490 & n501 ) | ( ~n490 & n4402 ) | ( n501 & n4402 ) ;
  assign n4404 = ( n486 & ~n487 ) | ( n486 & n4403 ) | ( ~n487 & n4403 ) ;
  assign n4405 = ( n1803 & ~n2029 ) | ( n1803 & n4404 ) | ( ~n2029 & n4404 ) ;
  assign n4406 = n600 | n2044 ;
  assign n4407 = ( ~n600 & n1530 ) | ( ~n600 & n2039 ) | ( n1530 & n2039 ) ;
  assign n4408 = ( n4077 & n4406 ) | ( n4077 & ~n4407 ) | ( n4406 & ~n4407 ) ;
  assign n4409 = ( n1533 & ~n4406 ) | ( n1533 & n4407 ) | ( ~n4406 & n4407 ) ;
  assign n4410 = ( n4405 & ~n4408 ) | ( n4405 & n4409 ) | ( ~n4408 & n4409 ) ;
  assign n4411 = ~n648 & n2244 ;
  assign n4412 = ( ~n584 & n623 ) | ( ~n584 & n1543 ) | ( n623 & n1543 ) ;
  assign n4413 = ( ~n2250 & n4411 ) | ( ~n2250 & n4412 ) | ( n4411 & n4412 ) ;
  assign n4414 = ( n627 & n2250 ) | ( n627 & ~n4411 ) | ( n2250 & ~n4411 ) ;
  assign n4415 = ( n4410 & ~n4413 ) | ( n4410 & n4414 ) | ( ~n4413 & n4414 ) ;
  assign n4416 = ( n778 & ~n2758 ) | ( n778 & n3871 ) | ( ~n2758 & n3871 ) ;
  assign n4417 = ~n678 & n2753 ;
  assign n4418 = ( n727 & ~n3187 ) | ( n727 & n3193 ) | ( ~n3187 & n3193 ) ;
  assign n4419 = ( n709 & ~n727 ) | ( n709 & n3296 ) | ( ~n727 & n3296 ) ;
  assign n4420 = ( n4417 & n4418 ) | ( n4417 & ~n4419 ) | ( n4418 & ~n4419 ) ;
  assign n4421 = ( n3765 & ~n4416 ) | ( n3765 & n4420 ) | ( ~n4416 & n4420 ) ;
  assign n4422 = ( n3862 & ~n4418 ) | ( n3862 & n4419 ) | ( ~n4418 & n4419 ) ;
  assign n4423 = ( ~n3765 & n4416 ) | ( ~n3765 & n4422 ) | ( n4416 & n4422 ) ;
  assign n4424 = ( n4415 & n4421 ) | ( n4415 & ~n4423 ) | ( n4421 & ~n4423 ) ;
  assign n4425 = x197 & ~n830 ;
  assign n4426 = n835 | n1611 ;
  assign n4427 = ( ~n826 & n1857 ) | ( ~n826 & n4211 ) | ( n1857 & n4211 ) ;
  assign n4428 = n823 & ~n865 ;
  assign n4429 = ( n1602 & n4427 ) | ( n1602 & ~n4428 ) | ( n4427 & ~n4428 ) ;
  assign n4430 = ~n853 & n4429 ;
  assign n4431 = ( n2770 & ~n4426 ) | ( n2770 & n4430 ) | ( ~n4426 & n4430 ) ;
  assign n4432 = n4425 & ~n4431 ;
  assign n4433 = ( n1605 & n2080 ) | ( n1605 & ~n2082 ) | ( n2080 & ~n2082 ) ;
  assign n4434 = ( ~n2770 & n4426 ) | ( ~n2770 & n4433 ) | ( n4426 & n4433 ) ;
  assign n4435 = n4425 & n4434 ;
  assign n4436 = ( n4424 & n4432 ) | ( n4424 & n4435 ) | ( n4432 & n4435 ) ;
  assign n4437 = x72 | n1303 ;
  assign n4438 = ~n897 & n4437 ;
  assign n4439 = ( ~n895 & n906 ) | ( ~n895 & n4438 ) | ( n906 & n4438 ) ;
  assign n4440 = ( n891 & ~n892 ) | ( n891 & n4439 ) | ( ~n892 & n4439 ) ;
  assign n4441 = ( n1881 & ~n2099 ) | ( n1881 & n4440 ) | ( ~n2099 & n4440 ) ;
  assign n4442 = n1005 | n2114 ;
  assign n4443 = ( ~n1005 & n1629 ) | ( ~n1005 & n2109 ) | ( n1629 & n2109 ) ;
  assign n4444 = ( n4114 & n4442 ) | ( n4114 & ~n4443 ) | ( n4442 & ~n4443 ) ;
  assign n4445 = ( n1632 & ~n4442 ) | ( n1632 & n4443 ) | ( ~n4442 & n4443 ) ;
  assign n4446 = ( n4441 & ~n4444 ) | ( n4441 & n4445 ) | ( ~n4444 & n4445 ) ;
  assign n4447 = ~n1053 & n2300 ;
  assign n4448 = ( ~n989 & n1028 ) | ( ~n989 & n1642 ) | ( n1028 & n1642 ) ;
  assign n4449 = ( ~n2306 & n4447 ) | ( ~n2306 & n4448 ) | ( n4447 & n4448 ) ;
  assign n4450 = ( n1032 & n2306 ) | ( n1032 & ~n4447 ) | ( n2306 & ~n4447 ) ;
  assign n4451 = ( n4446 & ~n4449 ) | ( n4446 & n4450 ) | ( ~n4449 & n4450 ) ;
  assign n4452 = ( n1182 & ~n2797 ) | ( n1182 & n3909 ) | ( ~n2797 & n3909 ) ;
  assign n4453 = ~n1082 & n2792 ;
  assign n4454 = ( n1131 & ~n3223 ) | ( n1131 & n3229 ) | ( ~n3223 & n3229 ) ;
  assign n4455 = ( n1113 & ~n1131 ) | ( n1113 & n3335 ) | ( ~n1131 & n3335 ) ;
  assign n4456 = ( n4453 & n4454 ) | ( n4453 & ~n4455 ) | ( n4454 & ~n4455 ) ;
  assign n4457 = ( n3803 & ~n4452 ) | ( n3803 & n4456 ) | ( ~n4452 & n4456 ) ;
  assign n4458 = ( n3900 & ~n4454 ) | ( n3900 & n4455 ) | ( ~n4454 & n4455 ) ;
  assign n4459 = ( ~n3803 & n4452 ) | ( ~n3803 & n4458 ) | ( n4452 & n4458 ) ;
  assign n4460 = ( n4451 & n4457 ) | ( n4451 & ~n4459 ) | ( n4457 & ~n4459 ) ;
  assign n4461 = x198 & ~n1234 ;
  assign n4462 = n1239 | n1709 ;
  assign n4463 = ( ~n1230 & n1935 ) | ( ~n1230 & n4248 ) | ( n1935 & n4248 ) ;
  assign n4464 = n1227 & ~n1269 ;
  assign n4465 = ( n1700 & n4463 ) | ( n1700 & ~n4464 ) | ( n4463 & ~n4464 ) ;
  assign n4466 = ~n1257 & n4465 ;
  assign n4467 = ( n2809 & ~n4462 ) | ( n2809 & n4466 ) | ( ~n4462 & n4466 ) ;
  assign n4468 = n4461 & ~n4467 ;
  assign n4469 = ( n1703 & n2150 ) | ( n1703 & ~n2152 ) | ( n2150 & ~n2152 ) ;
  assign n4470 = ( ~n2809 & n4462 ) | ( ~n2809 & n4469 ) | ( n4462 & n4469 ) ;
  assign n4471 = n4461 & n4470 ;
  assign n4472 = ( n4460 & n4468 ) | ( n4460 & n4471 ) | ( n4468 & n4471 ) ;
  assign n4473 = x73 | n498 ;
  assign n4474 = ~n1301 & n4473 ;
  assign n4475 = ( ~n1299 & n1310 ) | ( ~n1299 & n4474 ) | ( n1310 & n4474 ) ;
  assign n4476 = ( n1295 & ~n1296 ) | ( n1295 & n4475 ) | ( ~n1296 & n4475 ) ;
  assign n4477 = ( n1959 & ~n2169 ) | ( n1959 & n4476 ) | ( ~n2169 & n4476 ) ;
  assign n4478 = n1409 | n2184 ;
  assign n4479 = ( ~n1409 & n1727 ) | ( ~n1409 & n2179 ) | ( n1727 & n2179 ) ;
  assign n4480 = ( n4151 & n4478 ) | ( n4151 & ~n4479 ) | ( n4478 & ~n4479 ) ;
  assign n4481 = ( n1730 & ~n4478 ) | ( n1730 & n4479 ) | ( ~n4478 & n4479 ) ;
  assign n4482 = ( n4477 & ~n4480 ) | ( n4477 & n4481 ) | ( ~n4480 & n4481 ) ;
  assign n4483 = ~n1457 & n2356 ;
  assign n4484 = ( ~n1393 & n1432 ) | ( ~n1393 & n1740 ) | ( n1432 & n1740 ) ;
  assign n4485 = ( ~n2362 & n4483 ) | ( ~n2362 & n4484 ) | ( n4483 & n4484 ) ;
  assign n4486 = ( n1436 & n2362 ) | ( n1436 & ~n4483 ) | ( n2362 & ~n4483 ) ;
  assign n4487 = ( n4482 & ~n4485 ) | ( n4482 & n4486 ) | ( ~n4485 & n4486 ) ;
  assign n4488 = ( n359 & ~n377 ) | ( n359 & n3947 ) | ( ~n377 & n3947 ) ;
  assign n4489 = ~n297 & n2830 ;
  assign n4490 = ( n348 & ~n3259 ) | ( n348 & n3265 ) | ( ~n3259 & n3265 ) ;
  assign n4491 = ( n333 & ~n348 ) | ( n333 & n3374 ) | ( ~n348 & n3374 ) ;
  assign n4492 = ( n4489 & n4490 ) | ( n4489 & ~n4491 ) | ( n4490 & ~n4491 ) ;
  assign n4493 = ( n3841 & ~n4488 ) | ( n3841 & n4492 ) | ( ~n4488 & n4492 ) ;
  assign n4494 = ( n3938 & ~n4490 ) | ( n3938 & n4491 ) | ( ~n4490 & n4491 ) ;
  assign n4495 = ( ~n3841 & n4488 ) | ( ~n3841 & n4494 ) | ( n4488 & n4494 ) ;
  assign n4496 = ( n4487 & n4493 ) | ( n4487 & ~n4495 ) | ( n4493 & ~n4495 ) ;
  assign n4497 = x199 & ~n491 ;
  assign n4498 = n496 | n1794 ;
  assign n4499 = ~n445 & n1506 ;
  assign n4500 = ( n416 & n1786 ) | ( n416 & ~n4499 ) | ( n1786 & ~n4499 ) ;
  assign n4501 = ~n452 & n4500 ;
  assign n4502 = ( n2846 & ~n4498 ) | ( n2846 & n4501 ) | ( ~n4498 & n4501 ) ;
  assign n4503 = n4497 & ~n4502 ;
  assign n4504 = ( n423 & ~n463 ) | ( n423 & n1789 ) | ( ~n463 & n1789 ) ;
  assign n4505 = ( ~n2846 & n4498 ) | ( ~n2846 & n4504 ) | ( n4498 & n4504 ) ;
  assign n4506 = n4497 & n4505 ;
  assign n4507 = ( n4496 & n4503 ) | ( n4496 & n4506 ) | ( n4503 & n4506 ) ;
  assign n4508 = x74 | n903 ;
  assign n4509 = ~n489 & n4508 ;
  assign n4510 = ( ~n481 & n485 ) | ( ~n481 & n4509 ) | ( n485 & n4509 ) ;
  assign n4511 = ( ~n507 & n1520 ) | ( ~n507 & n4510 ) | ( n1520 & n4510 ) ;
  assign n4512 = ( n2033 & ~n2226 ) | ( n2033 & n4511 ) | ( ~n2226 & n4511 ) ;
  assign n4513 = n610 | n2238 ;
  assign n4514 = ( ~n610 & n624 ) | ( ~n610 & n2234 ) | ( n624 & n2234 ) ;
  assign n4515 = ( n4188 & n4513 ) | ( n4188 & ~n4514 ) | ( n4513 & ~n4514 ) ;
  assign n4516 = ( n1812 & ~n4513 ) | ( n1812 & n4514 ) | ( ~n4513 & n4514 ) ;
  assign n4517 = ( n4512 & ~n4515 ) | ( n4512 & n4516 ) | ( ~n4515 & n4516 ) ;
  assign n4518 = ~n635 & n2400 ;
  assign n4519 = ( ~n578 & n628 ) | ( ~n578 & n1821 ) | ( n628 & n1821 ) ;
  assign n4520 = ( ~n2406 & n4518 ) | ( ~n2406 & n4519 ) | ( n4518 & n4519 ) ;
  assign n4521 = ( n1554 & n2406 ) | ( n1554 & ~n4518 ) | ( n2406 & ~n4518 ) ;
  assign n4522 = ( n4517 & ~n4520 ) | ( n4517 & n4521 ) | ( ~n4520 & n4521 ) ;
  assign n4523 = ( n764 & ~n782 ) | ( n764 & n3985 ) | ( ~n782 & n3985 ) ;
  assign n4524 = ~n702 & n2867 ;
  assign n4525 = ( n753 & ~n3298 ) | ( n753 & n3304 ) | ( ~n3298 & n3304 ) ;
  assign n4526 = ( n738 & ~n753 ) | ( n738 & n3413 ) | ( ~n753 & n3413 ) ;
  assign n4527 = ( n4524 & n4525 ) | ( n4524 & ~n4526 ) | ( n4525 & ~n4526 ) ;
  assign n4528 = ( n3879 & ~n4523 ) | ( n3879 & n4527 ) | ( ~n4523 & n4527 ) ;
  assign n4529 = ( n3977 & ~n4525 ) | ( n3977 & n4526 ) | ( ~n4525 & n4526 ) ;
  assign n4530 = ( ~n3879 & n4523 ) | ( ~n3879 & n4529 ) | ( n4523 & n4529 ) ;
  assign n4531 = ( n4522 & n4528 ) | ( n4522 & ~n4530 ) | ( n4528 & ~n4530 ) ;
  assign n4532 = x200 & ~n896 ;
  assign n4533 = n901 | n1872 ;
  assign n4534 = ~n850 & n1605 ;
  assign n4535 = ( n821 & n1864 ) | ( n821 & ~n4534 ) | ( n1864 & ~n4534 ) ;
  assign n4536 = ~n857 & n4535 ;
  assign n4537 = ( n2883 & ~n4533 ) | ( n2883 & n4536 ) | ( ~n4533 & n4536 ) ;
  assign n4538 = n4532 & ~n4537 ;
  assign n4539 = ( n828 & ~n868 ) | ( n828 & n1867 ) | ( ~n868 & n1867 ) ;
  assign n4540 = ( ~n2883 & n4533 ) | ( ~n2883 & n4539 ) | ( n4533 & n4539 ) ;
  assign n4541 = n4532 & n4540 ;
  assign n4542 = ( n4531 & n4538 ) | ( n4531 & n4541 ) | ( n4538 & n4541 ) ;
  assign n4543 = x75 | n1307 ;
  assign n4544 = ~n894 & n4543 ;
  assign n4545 = ( ~n886 & n890 ) | ( ~n886 & n4544 ) | ( n890 & n4544 ) ;
  assign n4546 = ( ~n912 & n1619 ) | ( ~n912 & n4545 ) | ( n1619 & n4545 ) ;
  assign n4547 = ( n2103 & ~n2282 ) | ( n2103 & n4546 ) | ( ~n2282 & n4546 ) ;
  assign n4548 = n1015 | n2294 ;
  assign n4549 = ( ~n1015 & n1029 ) | ( ~n1015 & n2290 ) | ( n1029 & n2290 ) ;
  assign n4550 = ( n4225 & n4548 ) | ( n4225 & ~n4549 ) | ( n4548 & ~n4549 ) ;
  assign n4551 = ( n1890 & ~n4548 ) | ( n1890 & n4549 ) | ( ~n4548 & n4549 ) ;
  assign n4552 = ( n4547 & ~n4550 ) | ( n4547 & n4551 ) | ( ~n4550 & n4551 ) ;
  assign n4553 = ~n1040 & n2444 ;
  assign n4554 = ( ~n983 & n1033 ) | ( ~n983 & n1899 ) | ( n1033 & n1899 ) ;
  assign n4555 = ( ~n2450 & n4553 ) | ( ~n2450 & n4554 ) | ( n4553 & n4554 ) ;
  assign n4556 = ( n1653 & n2450 ) | ( n1653 & ~n4553 ) | ( n2450 & ~n4553 ) ;
  assign n4557 = ( n4552 & ~n4555 ) | ( n4552 & n4556 ) | ( ~n4555 & n4556 ) ;
  assign n4558 = ( n1168 & ~n1186 ) | ( n1168 & n4023 ) | ( ~n1186 & n4023 ) ;
  assign n4559 = ~n1106 & n2904 ;
  assign n4560 = ( n1157 & ~n3337 ) | ( n1157 & n3343 ) | ( ~n3337 & n3343 ) ;
  assign n4561 = ( n1142 & ~n1157 ) | ( n1142 & n3452 ) | ( ~n1157 & n3452 ) ;
  assign n4562 = ( n4559 & n4560 ) | ( n4559 & ~n4561 ) | ( n4560 & ~n4561 ) ;
  assign n4563 = ( n3917 & ~n4558 ) | ( n3917 & n4562 ) | ( ~n4558 & n4562 ) ;
  assign n4564 = ( n4015 & ~n4560 ) | ( n4015 & n4561 ) | ( ~n4560 & n4561 ) ;
  assign n4565 = ( ~n3917 & n4558 ) | ( ~n3917 & n4564 ) | ( n4558 & n4564 ) ;
  assign n4566 = ( n4557 & n4563 ) | ( n4557 & ~n4565 ) | ( n4563 & ~n4565 ) ;
  assign n4567 = x201 & ~n1300 ;
  assign n4568 = n1305 | n1950 ;
  assign n4569 = ~n1254 & n1703 ;
  assign n4570 = ( n1225 & n1942 ) | ( n1225 & ~n4569 ) | ( n1942 & ~n4569 ) ;
  assign n4571 = ~n1261 & n4570 ;
  assign n4572 = ( n2920 & ~n4568 ) | ( n2920 & n4571 ) | ( ~n4568 & n4571 ) ;
  assign n4573 = n4567 & ~n4572 ;
  assign n4574 = ( n1232 & ~n1272 ) | ( n1232 & n1945 ) | ( ~n1272 & n1945 ) ;
  assign n4575 = ( ~n2920 & n4568 ) | ( ~n2920 & n4574 ) | ( n4568 & n4574 ) ;
  assign n4576 = n4567 & n4575 ;
  assign n4577 = ( n4566 & n4573 ) | ( n4566 & n4576 ) | ( n4573 & n4576 ) ;
  assign n4578 = x76 | n482 ;
  assign n4579 = ~n1298 & n4578 ;
  assign n4580 = ( ~n1290 & n1294 ) | ( ~n1290 & n4579 ) | ( n1294 & n4579 ) ;
  assign n4581 = ( ~n1316 & n1717 ) | ( ~n1316 & n4580 ) | ( n1717 & n4580 ) ;
  assign n4582 = ( n2173 & ~n2338 ) | ( n2173 & n4581 ) | ( ~n2338 & n4581 ) ;
  assign n4583 = n1419 | n2350 ;
  assign n4584 = ( ~n1419 & n1433 ) | ( ~n1419 & n2346 ) | ( n1433 & n2346 ) ;
  assign n4585 = ( n4262 & n4583 ) | ( n4262 & ~n4584 ) | ( n4583 & ~n4584 ) ;
  assign n4586 = ( n1968 & ~n4583 ) | ( n1968 & n4584 ) | ( ~n4583 & n4584 ) ;
  assign n4587 = ( n4582 & ~n4585 ) | ( n4582 & n4586 ) | ( ~n4585 & n4586 ) ;
  assign n4588 = ~n1444 & n2488 ;
  assign n4589 = ( ~n1387 & n1437 ) | ( ~n1387 & n1977 ) | ( n1437 & n1977 ) ;
  assign n4590 = ( ~n2494 & n4588 ) | ( ~n2494 & n4589 ) | ( n4588 & n4589 ) ;
  assign n4591 = ( n1751 & n2494 ) | ( n1751 & ~n4588 ) | ( n2494 & ~n4588 ) ;
  assign n4592 = ( n4587 & ~n4590 ) | ( n4587 & n4591 ) | ( ~n4590 & n4591 ) ;
  assign n4593 = ( n402 & ~n1497 ) | ( n402 & n4061 ) | ( ~n1497 & n4061 ) ;
  assign n4594 = ~n289 & n2941 ;
  assign n4595 = ( n349 & ~n3376 ) | ( n349 & n3382 ) | ( ~n3376 & n3382 ) ;
  assign n4596 = ( n340 & ~n349 ) | ( n340 & n3491 ) | ( ~n349 & n3491 ) ;
  assign n4597 = ( n4594 & n4595 ) | ( n4594 & ~n4596 ) | ( n4595 & ~n4596 ) ;
  assign n4598 = ( n3955 & ~n4593 ) | ( n3955 & n4597 ) | ( ~n4593 & n4597 ) ;
  assign n4599 = ( n4053 & ~n4595 ) | ( n4053 & n4596 ) | ( ~n4595 & n4596 ) ;
  assign n4600 = ( ~n3955 & n4593 ) | ( ~n3955 & n4599 ) | ( n4593 & n4599 ) ;
  assign n4601 = ( n4592 & n4598 ) | ( n4592 & ~n4600 ) | ( n4598 & ~n4600 ) ;
  assign n4602 = x202 & ~n488 ;
  assign n4603 = n500 | n2021 ;
  assign n4604 = ~n442 & n1789 ;
  assign n4605 = ( n1504 & n2013 ) | ( n1504 & ~n4604 ) | ( n2013 & ~n4604 ) ;
  assign n4606 = ~n436 & n4605 ;
  assign n4607 = ( n2957 & ~n4603 ) | ( n2957 & n4606 ) | ( ~n4603 & n4606 ) ;
  assign n4608 = n4602 & ~n4607 ;
  assign n4609 = ( n1508 & ~n1515 ) | ( n1508 & n2016 ) | ( ~n1515 & n2016 ) ;
  assign n4610 = ( ~n2957 & n4603 ) | ( ~n2957 & n4609 ) | ( n4603 & n4609 ) ;
  assign n4611 = n4602 & n4610 ;
  assign n4612 = ( n4601 & n4608 ) | ( n4601 & n4611 ) | ( n4608 & n4611 ) ;
  assign n4613 = x77 | n887 ;
  assign n4614 = ~n480 & n4613 ;
  assign n4615 = ( ~n506 & n511 ) | ( ~n506 & n4614 ) | ( n511 & n4614 ) ;
  assign n4616 = ( ~n1523 & n1803 ) | ( ~n1523 & n4615 ) | ( n1803 & n4615 ) ;
  assign n4617 = ( ~n569 & n2229 ) | ( ~n569 & n4616 ) | ( n2229 & n4616 ) ;
  assign n4618 = n591 | n612 ;
  assign n4619 = ( ~n591 & n625 ) | ( ~n591 & n2393 ) | ( n625 & n2393 ) ;
  assign n4620 = ( n4298 & n4618 ) | ( n4298 & ~n4619 ) | ( n4618 & ~n4619 ) ;
  assign n4621 = ( n2039 & ~n4618 ) | ( n2039 & n4619 ) | ( ~n4618 & n4619 ) ;
  assign n4622 = ( n4617 & ~n4620 ) | ( n4617 & n4621 ) | ( ~n4620 & n4621 ) ;
  assign n4623 = ~n1559 & n2526 ;
  assign n4624 = ( ~n619 & n1549 ) | ( ~n619 & n2048 ) | ( n1549 & n2048 ) ;
  assign n4625 = ( ~n2531 & n4623 ) | ( ~n2531 & n4624 ) | ( n4623 & n4624 ) ;
  assign n4626 = ( n1830 & n2531 ) | ( n1830 & ~n4623 ) | ( n2531 & ~n4623 ) ;
  assign n4627 = ( n4622 & ~n4625 ) | ( n4622 & n4626 ) | ( ~n4625 & n4626 ) ;
  assign n4628 = ( n807 & ~n1596 ) | ( n807 & n4098 ) | ( ~n1596 & n4098 ) ;
  assign n4629 = ~n694 & n2977 ;
  assign n4630 = ( n754 & ~n3415 ) | ( n754 & n3421 ) | ( ~n3415 & n3421 ) ;
  assign n4631 = ( n745 & ~n754 ) | ( n745 & n3529 ) | ( ~n754 & n3529 ) ;
  assign n4632 = ( n4629 & n4630 ) | ( n4629 & ~n4631 ) | ( n4630 & ~n4631 ) ;
  assign n4633 = ( n3993 & ~n4628 ) | ( n3993 & n4632 ) | ( ~n4628 & n4632 ) ;
  assign n4634 = ( n4090 & ~n4630 ) | ( n4090 & n4631 ) | ( ~n4630 & n4631 ) ;
  assign n4635 = ( ~n3993 & n4628 ) | ( ~n3993 & n4634 ) | ( n4628 & n4634 ) ;
  assign n4636 = ( n4627 & n4633 ) | ( n4627 & ~n4635 ) | ( n4633 & ~n4635 ) ;
  assign n4637 = x203 & ~n893 ;
  assign n4638 = n905 | n2091 ;
  assign n4639 = ~n847 & n1867 ;
  assign n4640 = ( n1603 & n2083 ) | ( n1603 & ~n4639 ) | ( n2083 & ~n4639 ) ;
  assign n4641 = ~n841 & n4640 ;
  assign n4642 = ( n2993 & ~n4638 ) | ( n2993 & n4641 ) | ( ~n4638 & n4641 ) ;
  assign n4643 = n4637 & ~n4642 ;
  assign n4644 = ( n1607 & ~n1614 ) | ( n1607 & n2086 ) | ( ~n1614 & n2086 ) ;
  assign n4645 = ( ~n2993 & n4638 ) | ( ~n2993 & n4644 ) | ( n4638 & n4644 ) ;
  assign n4646 = n4637 & n4645 ;
  assign n4647 = ( n4636 & n4643 ) | ( n4636 & n4646 ) | ( n4643 & n4646 ) ;
  assign n4648 = x78 | n1291 ;
  assign n4649 = ~n885 & n4648 ;
  assign n4650 = ( ~n911 & n916 ) | ( ~n911 & n4649 ) | ( n916 & n4649 ) ;
  assign n4651 = ( ~n1622 & n1881 ) | ( ~n1622 & n4650 ) | ( n1881 & n4650 ) ;
  assign n4652 = ( ~n974 & n2285 ) | ( ~n974 & n4651 ) | ( n2285 & n4651 ) ;
  assign n4653 = n996 | n1017 ;
  assign n4654 = ( ~n996 & n1030 ) | ( ~n996 & n2437 ) | ( n1030 & n2437 ) ;
  assign n4655 = ( n4334 & n4653 ) | ( n4334 & ~n4654 ) | ( n4653 & ~n4654 ) ;
  assign n4656 = ( n2109 & ~n4653 ) | ( n2109 & n4654 ) | ( ~n4653 & n4654 ) ;
  assign n4657 = ( n4652 & ~n4655 ) | ( n4652 & n4656 ) | ( ~n4655 & n4656 ) ;
  assign n4658 = ~n1658 & n2563 ;
  assign n4659 = ( ~n1024 & n1648 ) | ( ~n1024 & n2118 ) | ( n1648 & n2118 ) ;
  assign n4660 = ( ~n2568 & n4658 ) | ( ~n2568 & n4659 ) | ( n4658 & n4659 ) ;
  assign n4661 = ( n1908 & n2568 ) | ( n1908 & ~n4658 ) | ( n2568 & ~n4658 ) ;
  assign n4662 = ( n4657 & ~n4660 ) | ( n4657 & n4661 ) | ( ~n4660 & n4661 ) ;
  assign n4663 = ( n1211 & ~n1694 ) | ( n1211 & n4135 ) | ( ~n1694 & n4135 ) ;
  assign n4664 = ~n1098 & n3013 ;
  assign n4665 = ( n1158 & ~n3454 ) | ( n1158 & n3460 ) | ( ~n3454 & n3460 ) ;
  assign n4666 = ( n1149 & ~n1158 ) | ( n1149 & n3567 ) | ( ~n1158 & n3567 ) ;
  assign n4667 = ( n4664 & n4665 ) | ( n4664 & ~n4666 ) | ( n4665 & ~n4666 ) ;
  assign n4668 = ( n4031 & ~n4663 ) | ( n4031 & n4667 ) | ( ~n4663 & n4667 ) ;
  assign n4669 = ( n4127 & ~n4665 ) | ( n4127 & n4666 ) | ( ~n4665 & n4666 ) ;
  assign n4670 = ( ~n4031 & n4663 ) | ( ~n4031 & n4669 ) | ( n4663 & n4669 ) ;
  assign n4671 = ( n4662 & n4668 ) | ( n4662 & ~n4670 ) | ( n4668 & ~n4670 ) ;
  assign n4672 = x204 & ~n1297 ;
  assign n4673 = n1309 | n2161 ;
  assign n4674 = ~n1251 & n1945 ;
  assign n4675 = ( n1701 & n2153 ) | ( n1701 & ~n4674 ) | ( n2153 & ~n4674 ) ;
  assign n4676 = ~n1245 & n4675 ;
  assign n4677 = ( n3029 & ~n4673 ) | ( n3029 & n4676 ) | ( ~n4673 & n4676 ) ;
  assign n4678 = n4672 & ~n4677 ;
  assign n4679 = ( n1705 & ~n1712 ) | ( n1705 & n2156 ) | ( ~n1712 & n2156 ) ;
  assign n4680 = ( ~n3029 & n4673 ) | ( ~n3029 & n4679 ) | ( n4673 & n4679 ) ;
  assign n4681 = n4672 & n4680 ;
  assign n4682 = ( n4671 & n4678 ) | ( n4671 & n4681 ) | ( n4678 & n4681 ) ;
  assign n4683 = x79 | n476 ;
  assign n4684 = ~n1289 & n4683 ;
  assign n4685 = ( ~n1315 & n1320 ) | ( ~n1315 & n4684 ) | ( n1320 & n4684 ) ;
  assign n4686 = ( ~n1720 & n1959 ) | ( ~n1720 & n4685 ) | ( n1959 & n4685 ) ;
  assign n4687 = ( ~n1378 & n2341 ) | ( ~n1378 & n4686 ) | ( n2341 & n4686 ) ;
  assign n4688 = n1400 | n1421 ;
  assign n4689 = ( ~n1400 & n1434 ) | ( ~n1400 & n2481 ) | ( n1434 & n2481 ) ;
  assign n4690 = ( n4370 & n4688 ) | ( n4370 & ~n4689 ) | ( n4688 & ~n4689 ) ;
  assign n4691 = ( n2179 & ~n4688 ) | ( n2179 & n4689 ) | ( ~n4688 & n4689 ) ;
  assign n4692 = ( n4687 & ~n4690 ) | ( n4687 & n4691 ) | ( ~n4690 & n4691 ) ;
  assign n4693 = ~n268 & n2600 ;
  assign n4694 = ( ~n1428 & n1746 ) | ( ~n1428 & n2188 ) | ( n1746 & n2188 ) ;
  assign n4695 = ( ~n2604 & n4693 ) | ( ~n2604 & n4694 ) | ( n4693 & n4694 ) ;
  assign n4696 = ( n1986 & n2604 ) | ( n1986 & ~n4693 ) | ( n2604 & ~n4693 ) ;
  assign n4697 = ( n4692 & ~n4695 ) | ( n4692 & n4696 ) | ( ~n4695 & n4696 ) ;
  assign n4698 = ( n409 & ~n1781 ) | ( n409 & n4172 ) | ( ~n1781 & n4172 ) ;
  assign n4699 = ~n307 & n3049 ;
  assign n4700 = ( n344 & ~n3493 ) | ( n344 & n3498 ) | ( ~n3493 & n3498 ) ;
  assign n4701 = ( n327 & ~n344 ) | ( n327 & n3605 ) | ( ~n344 & n3605 ) ;
  assign n4702 = ( n4699 & n4700 ) | ( n4699 & ~n4701 ) | ( n4700 & ~n4701 ) ;
  assign n4703 = ( n4068 & ~n4698 ) | ( n4068 & n4702 ) | ( ~n4698 & n4702 ) ;
  assign n4704 = ( n4164 & ~n4700 ) | ( n4164 & n4701 ) | ( ~n4700 & n4701 ) ;
  assign n4705 = ( ~n4068 & n4698 ) | ( ~n4068 & n4704 ) | ( n4698 & n4704 ) ;
  assign n4706 = ( n4697 & n4703 ) | ( n4697 & ~n4705 ) | ( n4703 & ~n4705 ) ;
  assign n4707 = x205 & ~n479 ;
  assign n4708 = n484 | n502 ;
  assign n4709 = ~n433 & n2016 ;
  assign n4710 = ( n465 & n1787 ) | ( n465 & ~n4709 ) | ( n1787 & ~n4709 ) ;
  assign n4711 = ~n430 & n4710 ;
  assign n4712 = ( n3066 & ~n4708 ) | ( n3066 & n4711 ) | ( ~n4708 & n4711 ) ;
  assign n4713 = n4707 & ~n4712 ;
  assign n4714 = ( n438 & n1791 ) | ( n438 & ~n1797 ) | ( n1791 & ~n1797 ) ;
  assign n4715 = ( ~n3066 & n4708 ) | ( ~n3066 & n4714 ) | ( n4708 & n4714 ) ;
  assign n4716 = n4707 & n4715 ;
  assign n4717 = ( n4706 & n4713 ) | ( n4706 & n4716 ) | ( n4713 & n4716 ) ;
  assign n4718 = x80 | n881 ;
  assign n4719 = ~n505 & n4718 ;
  assign n4720 = ( ~n471 & n475 ) | ( ~n471 & n4719 ) | ( n475 & n4719 ) ;
  assign n4721 = ( ~n567 & n2033 ) | ( ~n567 & n4720 ) | ( n2033 & n4720 ) ;
  assign n4722 = ( n539 & ~n1538 ) | ( n539 & n4721 ) | ( ~n1538 & n4721 ) ;
  assign n4723 = n588 | n1543 ;
  assign n4724 = ( ~n588 & n597 ) | ( ~n588 & n626 ) | ( n597 & n626 ) ;
  assign n4725 = ( n4406 & n4723 ) | ( n4406 & ~n4724 ) | ( n4723 & ~n4724 ) ;
  assign n4726 = ( n2234 & ~n4723 ) | ( n2234 & n4724 ) | ( ~n4723 & n4724 ) ;
  assign n4727 = ( n4722 & ~n4725 ) | ( n4722 & n4726 ) | ( ~n4725 & n4726 ) ;
  assign n4728 = ~n673 & n2635 ;
  assign n4729 = ( ~n644 & n656 ) | ( ~n644 & n2243 ) | ( n656 & n2243 ) ;
  assign n4730 = ( ~n2639 & n4728 ) | ( ~n2639 & n4729 ) | ( n4728 & n4729 ) ;
  assign n4731 = ( n2056 & n2639 ) | ( n2056 & ~n4728 ) | ( n2639 & ~n4728 ) ;
  assign n4732 = ( n4727 & ~n4730 ) | ( n4727 & n4731 ) | ( ~n4730 & n4731 ) ;
  assign n4733 = ( n814 & ~n1859 ) | ( n814 & n4209 ) | ( ~n1859 & n4209 ) ;
  assign n4734 = ~n712 & n3085 ;
  assign n4735 = ( n749 & ~n3531 ) | ( n749 & n3536 ) | ( ~n3531 & n3536 ) ;
  assign n4736 = ( n732 & ~n749 ) | ( n732 & n3643 ) | ( ~n749 & n3643 ) ;
  assign n4737 = ( n4734 & n4735 ) | ( n4734 & ~n4736 ) | ( n4735 & ~n4736 ) ;
  assign n4738 = ( n4105 & ~n4733 ) | ( n4105 & n4737 ) | ( ~n4733 & n4737 ) ;
  assign n4739 = ( n4201 & ~n4735 ) | ( n4201 & n4736 ) | ( ~n4735 & n4736 ) ;
  assign n4740 = ( ~n4105 & n4733 ) | ( ~n4105 & n4739 ) | ( n4733 & n4739 ) ;
  assign n4741 = ( n4732 & n4738 ) | ( n4732 & ~n4740 ) | ( n4738 & ~n4740 ) ;
  assign n4742 = x206 & ~n884 ;
  assign n4743 = n889 | n907 ;
  assign n4744 = ~n838 & n2086 ;
  assign n4745 = ( n870 & n1865 ) | ( n870 & ~n4744 ) | ( n1865 & ~n4744 ) ;
  assign n4746 = ~n835 & n4745 ;
  assign n4747 = ( n3102 & ~n4743 ) | ( n3102 & n4746 ) | ( ~n4743 & n4746 ) ;
  assign n4748 = n4742 & ~n4747 ;
  assign n4749 = ( n843 & n1869 ) | ( n843 & ~n1875 ) | ( n1869 & ~n1875 ) ;
  assign n4750 = ( ~n3102 & n4743 ) | ( ~n3102 & n4749 ) | ( n4743 & n4749 ) ;
  assign n4751 = n4742 & n4750 ;
  assign n4752 = ( n4741 & n4748 ) | ( n4741 & n4751 ) | ( n4748 & n4751 ) ;
  assign n4753 = x81 | n1285 ;
  assign n4754 = ~n910 & n4753 ;
  assign n4755 = ( ~n876 & n880 ) | ( ~n876 & n4754 ) | ( n880 & n4754 ) ;
  assign n4756 = ( ~n972 & n2103 ) | ( ~n972 & n4755 ) | ( n2103 & n4755 ) ;
  assign n4757 = ( n944 & ~n1637 ) | ( n944 & n4756 ) | ( ~n1637 & n4756 ) ;
  assign n4758 = n993 | n1642 ;
  assign n4759 = ( ~n993 & n1002 ) | ( ~n993 & n1031 ) | ( n1002 & n1031 ) ;
  assign n4760 = ( n4442 & n4758 ) | ( n4442 & ~n4759 ) | ( n4758 & ~n4759 ) ;
  assign n4761 = ( n2290 & ~n4758 ) | ( n2290 & n4759 ) | ( ~n4758 & n4759 ) ;
  assign n4762 = ( n4757 & ~n4760 ) | ( n4757 & n4761 ) | ( ~n4760 & n4761 ) ;
  assign n4763 = ~n1077 & n2670 ;
  assign n4764 = ( ~n1049 & n1061 ) | ( ~n1049 & n2299 ) | ( n1061 & n2299 ) ;
  assign n4765 = ( ~n2674 & n4763 ) | ( ~n2674 & n4764 ) | ( n4763 & n4764 ) ;
  assign n4766 = ( n2126 & n2674 ) | ( n2126 & ~n4763 ) | ( n2674 & ~n4763 ) ;
  assign n4767 = ( n4762 & ~n4765 ) | ( n4762 & n4766 ) | ( ~n4765 & n4766 ) ;
  assign n4768 = ( n1218 & ~n1937 ) | ( n1218 & n4246 ) | ( ~n1937 & n4246 ) ;
  assign n4769 = ~n1116 & n3121 ;
  assign n4770 = ( n1153 & ~n3569 ) | ( n1153 & n3574 ) | ( ~n3569 & n3574 ) ;
  assign n4771 = ( n1136 & ~n1153 ) | ( n1136 & n3681 ) | ( ~n1153 & n3681 ) ;
  assign n4772 = ( n4769 & n4770 ) | ( n4769 & ~n4771 ) | ( n4770 & ~n4771 ) ;
  assign n4773 = ( n4142 & ~n4768 ) | ( n4142 & n4772 ) | ( ~n4768 & n4772 ) ;
  assign n4774 = ( n4238 & ~n4770 ) | ( n4238 & n4771 ) | ( ~n4770 & n4771 ) ;
  assign n4775 = ( ~n4142 & n4768 ) | ( ~n4142 & n4774 ) | ( n4768 & n4774 ) ;
  assign n4776 = ( n4767 & n4773 ) | ( n4767 & ~n4775 ) | ( n4773 & ~n4775 ) ;
  assign n4777 = x207 & ~n1288 ;
  assign n4778 = n1293 | n1311 ;
  assign n4779 = ~n1242 & n2156 ;
  assign n4780 = ( n1274 & n1943 ) | ( n1274 & ~n4779 ) | ( n1943 & ~n4779 ) ;
  assign n4781 = ~n1239 & n4780 ;
  assign n4782 = ( n3138 & ~n4778 ) | ( n3138 & n4781 ) | ( ~n4778 & n4781 ) ;
  assign n4783 = n4777 & ~n4782 ;
  assign n4784 = ( n1247 & n1947 ) | ( n1247 & ~n1953 ) | ( n1947 & ~n1953 ) ;
  assign n4785 = ( ~n3138 & n4778 ) | ( ~n3138 & n4784 ) | ( n4778 & n4784 ) ;
  assign n4786 = n4777 & n4785 ;
  assign n4787 = ( n4776 & n4783 ) | ( n4776 & n4786 ) | ( n4783 & n4786 ) ;
  assign n4788 = x82 | n472 ;
  assign n4789 = ~n1314 & n4788 ;
  assign n4790 = ( ~n1280 & n1284 ) | ( ~n1280 & n4789 ) | ( n1284 & n4789 ) ;
  assign n4791 = ( ~n1376 & n2173 ) | ( ~n1376 & n4790 ) | ( n2173 & n4790 ) ;
  assign n4792 = ( n1348 & ~n1735 ) | ( n1348 & n4791 ) | ( ~n1735 & n4791 ) ;
  assign n4793 = n1397 | n1740 ;
  assign n4794 = ( ~n1397 & n1406 ) | ( ~n1397 & n1435 ) | ( n1406 & n1435 ) ;
  assign n4795 = ( n4478 & n4793 ) | ( n4478 & ~n4794 ) | ( n4793 & ~n4794 ) ;
  assign n4796 = ( n2346 & ~n4793 ) | ( n2346 & n4794 ) | ( ~n4793 & n4794 ) ;
  assign n4797 = ( n4792 & ~n4795 ) | ( n4792 & n4796 ) | ( ~n4795 & n4796 ) ;
  assign n4798 = ~n276 & n2705 ;
  assign n4799 = ( ~n1453 & n1465 ) | ( ~n1453 & n2355 ) | ( n1465 & n2355 ) ;
  assign n4800 = ( ~n2709 & n4798 ) | ( ~n2709 & n4799 ) | ( n4798 & n4799 ) ;
  assign n4801 = ( n2196 & n2709 ) | ( n2196 & ~n4798 ) | ( n2709 & ~n4798 ) ;
  assign n4802 = ( n4797 & ~n4800 ) | ( n4797 & n4801 ) | ( ~n4800 & n4801 ) ;
  assign n4803 = ( n414 & ~n2008 ) | ( n414 & n4283 ) | ( ~n2008 & n4283 ) ;
  assign n4804 = ~n317 & n3157 ;
  assign n4805 = ( n381 & ~n3607 ) | ( n381 & n3612 ) | ( ~n3607 & n3612 ) ;
  assign n4806 = ( n365 & ~n381 ) | ( n365 & n3719 ) | ( ~n381 & n3719 ) ;
  assign n4807 = ( n4804 & n4805 ) | ( n4804 & ~n4806 ) | ( n4805 & ~n4806 ) ;
  assign n4808 = ( n4179 & ~n4803 ) | ( n4179 & n4807 ) | ( ~n4803 & n4807 ) ;
  assign n4809 = ( n4275 & ~n4805 ) | ( n4275 & n4806 ) | ( ~n4805 & n4806 ) ;
  assign n4810 = ( ~n4179 & n4803 ) | ( ~n4179 & n4809 ) | ( n4803 & n4809 ) ;
  assign n4811 = ( n4802 & n4808 ) | ( n4802 & ~n4810 ) | ( n4808 & ~n4810 ) ;
  assign n4812 = x208 & ~n504 ;
  assign n4813 = n478 | n1521 ;
  assign n4814 = ~n427 & n438 ;
  assign n4815 = ( n1516 & n2014 ) | ( n1516 & ~n4814 ) | ( n2014 & ~n4814 ) ;
  assign n4816 = ~n496 & n4815 ;
  assign n4817 = ( n3173 & ~n4813 ) | ( n3173 & n4816 ) | ( ~n4813 & n4816 ) ;
  assign n4818 = n4812 & ~n4817 ;
  assign n4819 = ( n1510 & n2018 ) | ( n1510 & ~n2024 ) | ( n2018 & ~n2024 ) ;
  assign n4820 = ( ~n3173 & n4813 ) | ( ~n3173 & n4819 ) | ( n4813 & n4819 ) ;
  assign n4821 = n4812 & n4820 ;
  assign n4822 = ( n4811 & n4818 ) | ( n4811 & n4821 ) | ( n4818 & n4821 ) ;
  assign n4823 = x83 | n877 ;
  assign n4824 = ~n470 & n4823 ;
  assign n4825 = ( ~n546 & n550 ) | ( ~n546 & n4824 ) | ( n550 & n4824 ) ;
  assign n4826 = ( ~n568 & n2229 ) | ( ~n568 & n4825 ) | ( n2229 & n4825 ) ;
  assign n4827 = ( n1532 & ~n1817 ) | ( n1532 & n4826 ) | ( ~n1817 & n4826 ) ;
  assign n4828 = n581 | n1821 ;
  assign n4829 = ( ~n581 & n585 ) | ( ~n581 & n1553 ) | ( n585 & n1553 ) ;
  assign n4830 = ( n4513 & n4828 ) | ( n4513 & ~n4829 ) | ( n4828 & ~n4829 ) ;
  assign n4831 = ( n2393 & ~n4828 ) | ( n2393 & n4829 ) | ( ~n4828 & n4829 ) ;
  assign n4832 = ( n4827 & ~n4830 ) | ( n4827 & n4831 ) | ( ~n4830 & n4831 ) ;
  assign n4833 = ~n681 & n2745 ;
  assign n4834 = ( ~n648 & n657 ) | ( ~n648 & n2399 ) | ( n657 & n2399 ) ;
  assign n4835 = ( ~n2753 & n4833 ) | ( ~n2753 & n4834 ) | ( n4833 & n4834 ) ;
  assign n4836 = ( n2250 & n2753 ) | ( n2250 & ~n4833 ) | ( n2753 & ~n4833 ) ;
  assign n4837 = ( n4832 & ~n4835 ) | ( n4832 & n4836 ) | ( ~n4835 & n4836 ) ;
  assign n4838 = ( n819 & ~n2078 ) | ( n819 & n4319 ) | ( ~n2078 & n4319 ) ;
  assign n4839 = ~n722 & n3193 ;
  assign n4840 = ( n786 & ~n3645 ) | ( n786 & n3650 ) | ( ~n3645 & n3650 ) ;
  assign n4841 = ( n770 & ~n786 ) | ( n770 & n3757 ) | ( ~n786 & n3757 ) ;
  assign n4842 = ( n4839 & n4840 ) | ( n4839 & ~n4841 ) | ( n4840 & ~n4841 ) ;
  assign n4843 = ( n4216 & ~n4838 ) | ( n4216 & n4842 ) | ( ~n4838 & n4842 ) ;
  assign n4844 = ( n4311 & ~n4840 ) | ( n4311 & n4841 ) | ( ~n4840 & n4841 ) ;
  assign n4845 = ( ~n4216 & n4838 ) | ( ~n4216 & n4844 ) | ( n4838 & n4844 ) ;
  assign n4846 = ( n4837 & n4843 ) | ( n4837 & ~n4845 ) | ( n4843 & ~n4845 ) ;
  assign n4847 = x209 & ~n909 ;
  assign n4848 = n883 | n1620 ;
  assign n4849 = ~n832 & n843 ;
  assign n4850 = ( n1615 & n2084 ) | ( n1615 & ~n4849 ) | ( n2084 & ~n4849 ) ;
  assign n4851 = ~n901 & n4850 ;
  assign n4852 = ( n3209 & ~n4848 ) | ( n3209 & n4851 ) | ( ~n4848 & n4851 ) ;
  assign n4853 = n4847 & ~n4852 ;
  assign n4854 = ( n1609 & n2088 ) | ( n1609 & ~n2094 ) | ( n2088 & ~n2094 ) ;
  assign n4855 = ( ~n3209 & n4848 ) | ( ~n3209 & n4854 ) | ( n4848 & n4854 ) ;
  assign n4856 = n4847 & n4855 ;
  assign n4857 = ( n4846 & n4853 ) | ( n4846 & n4856 ) | ( n4853 & n4856 ) ;
  assign n4858 = x84 | n1281 ;
  assign n4859 = ~n875 & n4858 ;
  assign n4860 = ( ~n951 & n955 ) | ( ~n951 & n4859 ) | ( n955 & n4859 ) ;
  assign n4861 = ( ~n973 & n2285 ) | ( ~n973 & n4860 ) | ( n2285 & n4860 ) ;
  assign n4862 = ( n1631 & ~n1895 ) | ( n1631 & n4861 ) | ( ~n1895 & n4861 ) ;
  assign n4863 = n986 | n1899 ;
  assign n4864 = ( ~n986 & n990 ) | ( ~n986 & n1652 ) | ( n990 & n1652 ) ;
  assign n4865 = ( n4548 & n4863 ) | ( n4548 & ~n4864 ) | ( n4863 & ~n4864 ) ;
  assign n4866 = ( n2437 & ~n4863 ) | ( n2437 & n4864 ) | ( ~n4863 & n4864 ) ;
  assign n4867 = ( n4862 & ~n4865 ) | ( n4862 & n4866 ) | ( ~n4865 & n4866 ) ;
  assign n4868 = ~n1085 & n2784 ;
  assign n4869 = ( ~n1053 & n1062 ) | ( ~n1053 & n2443 ) | ( n1062 & n2443 ) ;
  assign n4870 = ( ~n2792 & n4868 ) | ( ~n2792 & n4869 ) | ( n4868 & n4869 ) ;
  assign n4871 = ( n2306 & n2792 ) | ( n2306 & ~n4868 ) | ( n2792 & ~n4868 ) ;
  assign n4872 = ( n4867 & ~n4870 ) | ( n4867 & n4871 ) | ( ~n4870 & n4871 ) ;
  assign n4873 = ( n1223 & ~n2148 ) | ( n1223 & n4355 ) | ( ~n2148 & n4355 ) ;
  assign n4874 = ~n1126 & n3229 ;
  assign n4875 = ( n1190 & ~n3683 ) | ( n1190 & n3688 ) | ( ~n3683 & n3688 ) ;
  assign n4876 = ( n1174 & ~n1190 ) | ( n1174 & n3795 ) | ( ~n1190 & n3795 ) ;
  assign n4877 = ( n4874 & n4875 ) | ( n4874 & ~n4876 ) | ( n4875 & ~n4876 ) ;
  assign n4878 = ( n4253 & ~n4873 ) | ( n4253 & n4877 ) | ( ~n4873 & n4877 ) ;
  assign n4879 = ( n4347 & ~n4875 ) | ( n4347 & n4876 ) | ( ~n4875 & n4876 ) ;
  assign n4880 = ( ~n4253 & n4873 ) | ( ~n4253 & n4879 ) | ( n4873 & n4879 ) ;
  assign n4881 = ( n4872 & n4878 ) | ( n4872 & ~n4880 ) | ( n4878 & ~n4880 ) ;
  assign n4882 = x210 & ~n1313 ;
  assign n4883 = n1287 | n1718 ;
  assign n4884 = ~n1236 & n1247 ;
  assign n4885 = ( n1713 & n2154 ) | ( n1713 & ~n4884 ) | ( n2154 & ~n4884 ) ;
  assign n4886 = ~n1305 & n4885 ;
  assign n4887 = ( n3245 & ~n4883 ) | ( n3245 & n4886 ) | ( ~n4883 & n4886 ) ;
  assign n4888 = n4882 & ~n4887 ;
  assign n4889 = ( n1707 & n2158 ) | ( n1707 & ~n2164 ) | ( n2158 & ~n2164 ) ;
  assign n4890 = ( ~n3245 & n4883 ) | ( ~n3245 & n4889 ) | ( n4883 & n4889 ) ;
  assign n4891 = n4882 & n4890 ;
  assign n4892 = ( n4881 & n4888 ) | ( n4881 & n4891 ) | ( n4888 & n4891 ) ;
  assign n4893 = x85 | n547 ;
  assign n4894 = ~n1279 & n4893 ;
  assign n4895 = ( ~n1355 & n1359 ) | ( ~n1355 & n4894 ) | ( n1359 & n4894 ) ;
  assign n4896 = ( ~n1377 & n2341 ) | ( ~n1377 & n4895 ) | ( n2341 & n4895 ) ;
  assign n4897 = ( n1729 & ~n1973 ) | ( n1729 & n4896 ) | ( ~n1973 & n4896 ) ;
  assign n4898 = n1390 | n1977 ;
  assign n4899 = ( ~n1390 & n1394 ) | ( ~n1390 & n1750 ) | ( n1394 & n1750 ) ;
  assign n4900 = ( n4583 & n4898 ) | ( n4583 & ~n4899 ) | ( n4898 & ~n4899 ) ;
  assign n4901 = ( n2481 & ~n4898 ) | ( n2481 & n4899 ) | ( ~n4898 & n4899 ) ;
  assign n4902 = ( n4897 & ~n4900 ) | ( n4897 & n4901 ) | ( ~n4900 & n4901 ) ;
  assign n4903 = ~n280 & n2823 ;
  assign n4904 = ( ~n1457 & n1466 ) | ( ~n1457 & n2487 ) | ( n1466 & n2487 ) ;
  assign n4905 = ( ~n2830 & n4903 ) | ( ~n2830 & n4904 ) | ( n4903 & n4904 ) ;
  assign n4906 = ( n2362 & n2830 ) | ( n2362 & ~n4903 ) | ( n2830 & ~n4903 ) ;
  assign n4907 = ( n4902 & ~n4905 ) | ( n4902 & n4906 ) | ( ~n4905 & n4906 ) ;
  assign n4908 = ( ~n418 & n419 ) | ( ~n418 & n4391 ) | ( n419 & n4391 ) ;
  assign n4909 = ~n304 & n3265 ;
  assign n4910 = ( n382 & ~n3721 ) | ( n382 & n3726 ) | ( ~n3721 & n3726 ) ;
  assign n4911 = ( n372 & ~n382 ) | ( n372 & n3833 ) | ( ~n382 & n3833 ) ;
  assign n4912 = ( n4909 & n4910 ) | ( n4909 & ~n4911 ) | ( n4910 & ~n4911 ) ;
  assign n4913 = ( n4289 & ~n4908 ) | ( n4289 & n4912 ) | ( ~n4908 & n4912 ) ;
  assign n4914 = ( n4383 & ~n4910 ) | ( n4383 & n4911 ) | ( ~n4910 & n4911 ) ;
  assign n4915 = ( ~n4289 & n4908 ) | ( ~n4289 & n4914 ) | ( n4908 & n4914 ) ;
  assign n4916 = ( n4907 & n4913 ) | ( n4907 & ~n4915 ) | ( n4913 & ~n4915 ) ;
  assign n4917 = x211 & ~n469 ;
  assign n4918 = n474 | n1804 ;
  assign n4919 = ~n493 & n1510 ;
  assign n4920 = ( n466 & n1798 ) | ( n466 & ~n4919 ) | ( n1798 & ~n4919 ) ;
  assign n4921 = ~n500 & n4920 ;
  assign n4922 = ( n3281 & ~n4918 ) | ( n3281 & n4921 ) | ( ~n4918 & n4921 ) ;
  assign n4923 = n4917 & ~n4922 ;
  assign n4924 = ( n455 & n1793 ) | ( n455 & ~n2222 ) | ( n1793 & ~n2222 ) ;
  assign n4925 = ( ~n3281 & n4918 ) | ( ~n3281 & n4924 ) | ( n4918 & n4924 ) ;
  assign n4926 = n4917 & n4925 ;
  assign n4927 = ( n4916 & n4923 ) | ( n4916 & n4926 ) | ( n4923 & n4926 ) ;
  assign n4928 = x86 | n952 ;
  assign n4929 = ~n545 & n4928 ;
  assign n4930 = ( ~n543 & n554 ) | ( ~n543 & n4929 ) | ( n554 & n4929 ) ;
  assign n4931 = ( n539 & ~n540 ) | ( n539 & n4930 ) | ( ~n540 & n4930 ) ;
  assign n4932 = ( n528 & ~n2044 ) | ( n528 & n4931 ) | ( ~n2044 & n4931 ) ;
  assign n4933 = n575 | n2048 ;
  assign n4934 = ( ~n575 & n621 ) | ( ~n575 & n1829 ) | ( n621 & n1829 ) ;
  assign n4935 = ( n4618 & n4933 ) | ( n4618 & ~n4934 ) | ( n4933 & ~n4934 ) ;
  assign n4936 = ( n626 & ~n4933 ) | ( n626 & n4934 ) | ( ~n4933 & n4934 ) ;
  assign n4937 = ( n4932 & ~n4935 ) | ( n4932 & n4936 ) | ( ~n4935 & n4936 ) ;
  assign n4938 = ~n685 & n2860 ;
  assign n4939 = ( n659 & ~n2867 ) | ( n659 & n4938 ) | ( ~n2867 & n4938 ) ;
  assign n4940 = ( n2406 & n2867 ) | ( n2406 & ~n4938 ) | ( n2867 & ~n4938 ) ;
  assign n4941 = ( n4937 & ~n4939 ) | ( n4937 & n4940 ) | ( ~n4939 & n4940 ) ;
  assign n4942 = ( ~n823 & n824 ) | ( ~n823 & n4427 ) | ( n824 & n4427 ) ;
  assign n4943 = ~n709 & n3304 ;
  assign n4944 = ( n787 & ~n3759 ) | ( n787 & n3764 ) | ( ~n3759 & n3764 ) ;
  assign n4945 = ( n777 & ~n787 ) | ( n777 & n3871 ) | ( ~n787 & n3871 ) ;
  assign n4946 = ( n4943 & n4944 ) | ( n4943 & ~n4945 ) | ( n4944 & ~n4945 ) ;
  assign n4947 = ( n4325 & ~n4942 ) | ( n4325 & n4946 ) | ( ~n4942 & n4946 ) ;
  assign n4948 = ( n4419 & ~n4944 ) | ( n4419 & n4945 ) | ( ~n4944 & n4945 ) ;
  assign n4949 = ( ~n4325 & n4942 ) | ( ~n4325 & n4948 ) | ( n4942 & n4948 ) ;
  assign n4950 = ( n4941 & n4947 ) | ( n4941 & ~n4949 ) | ( n4947 & ~n4949 ) ;
  assign n4951 = x212 & ~n874 ;
  assign n4952 = n879 | n1882 ;
  assign n4953 = ~n898 & n1609 ;
  assign n4954 = ( n871 & n1876 ) | ( n871 & ~n4953 ) | ( n1876 & ~n4953 ) ;
  assign n4955 = ~n905 & n4954 ;
  assign n4956 = ( n3320 & ~n4952 ) | ( n3320 & n4955 ) | ( ~n4952 & n4955 ) ;
  assign n4957 = n4951 & ~n4956 ;
  assign n4958 = ( n860 & n1871 ) | ( n860 & ~n2278 ) | ( n1871 & ~n2278 ) ;
  assign n4959 = ( ~n3320 & n4952 ) | ( ~n3320 & n4958 ) | ( n4952 & n4958 ) ;
  assign n4960 = n4951 & n4959 ;
  assign n4961 = ( n4950 & n4957 ) | ( n4950 & n4960 ) | ( n4957 & n4960 ) ;
  assign n4962 = x87 | n1356 ;
  assign n4963 = ~n950 & n4962 ;
  assign n4964 = ( ~n948 & n959 ) | ( ~n948 & n4963 ) | ( n959 & n4963 ) ;
  assign n4965 = ( n944 & ~n945 ) | ( n944 & n4964 ) | ( ~n945 & n4964 ) ;
  assign n4966 = ( n933 & ~n2114 ) | ( n933 & n4965 ) | ( ~n2114 & n4965 ) ;
  assign n4967 = n980 | n2118 ;
  assign n4968 = ( ~n980 & n1026 ) | ( ~n980 & n1907 ) | ( n1026 & n1907 ) ;
  assign n4969 = ( n4653 & n4967 ) | ( n4653 & ~n4968 ) | ( n4967 & ~n4968 ) ;
  assign n4970 = ( n1031 & ~n4967 ) | ( n1031 & n4968 ) | ( ~n4967 & n4968 ) ;
  assign n4971 = ( n4966 & ~n4969 ) | ( n4966 & n4970 ) | ( ~n4969 & n4970 ) ;
  assign n4972 = ~n1089 & n2897 ;
  assign n4973 = ( n1064 & ~n2904 ) | ( n1064 & n4972 ) | ( ~n2904 & n4972 ) ;
  assign n4974 = ( n2450 & n2904 ) | ( n2450 & ~n4972 ) | ( n2904 & ~n4972 ) ;
  assign n4975 = ( n4971 & ~n4973 ) | ( n4971 & n4974 ) | ( ~n4973 & n4974 ) ;
  assign n4976 = ( ~n1227 & n1228 ) | ( ~n1227 & n4463 ) | ( n1228 & n4463 ) ;
  assign n4977 = ~n1113 & n3343 ;
  assign n4978 = ( n1191 & ~n3797 ) | ( n1191 & n3802 ) | ( ~n3797 & n3802 ) ;
  assign n4979 = ( n1181 & ~n1191 ) | ( n1181 & n3909 ) | ( ~n1191 & n3909 ) ;
  assign n4980 = ( n4977 & n4978 ) | ( n4977 & ~n4979 ) | ( n4978 & ~n4979 ) ;
  assign n4981 = ( n4361 & ~n4976 ) | ( n4361 & n4980 ) | ( ~n4976 & n4980 ) ;
  assign n4982 = ( n4455 & ~n4978 ) | ( n4455 & n4979 ) | ( ~n4978 & n4979 ) ;
  assign n4983 = ( ~n4361 & n4976 ) | ( ~n4361 & n4982 ) | ( n4976 & n4982 ) ;
  assign n4984 = ( n4975 & n4981 ) | ( n4975 & ~n4983 ) | ( n4981 & ~n4983 ) ;
  assign n4985 = x213 & ~n1278 ;
  assign n4986 = n1283 | n1960 ;
  assign n4987 = ~n1302 & n1707 ;
  assign n4988 = ( n1275 & n1954 ) | ( n1275 & ~n4987 ) | ( n1954 & ~n4987 ) ;
  assign n4989 = ~n1309 & n4988 ;
  assign n4990 = ( n3359 & ~n4986 ) | ( n3359 & n4989 ) | ( ~n4986 & n4989 ) ;
  assign n4991 = n4985 & ~n4990 ;
  assign n4992 = ( n1264 & n1949 ) | ( n1264 & ~n2334 ) | ( n1949 & ~n2334 ) ;
  assign n4993 = ( ~n3359 & n4986 ) | ( ~n3359 & n4992 ) | ( n4986 & n4992 ) ;
  assign n4994 = n4985 & n4993 ;
  assign n4995 = ( n4984 & n4991 ) | ( n4984 & n4994 ) | ( n4991 & n4994 ) ;
  assign n4996 = x88 | n551 ;
  assign n4997 = ~n1354 & n4996 ;
  assign n4998 = ( ~n1352 & n1363 ) | ( ~n1352 & n4997 ) | ( n1363 & n4997 ) ;
  assign n4999 = ( n1348 & ~n1349 ) | ( n1348 & n4998 ) | ( ~n1349 & n4998 ) ;
  assign n5000 = ( n1337 & ~n2184 ) | ( n1337 & n4999 ) | ( ~n2184 & n4999 ) ;
  assign n5001 = n1384 | n2188 ;
  assign n5002 = ( ~n1384 & n1430 ) | ( ~n1384 & n1985 ) | ( n1430 & n1985 ) ;
  assign n5003 = ( n4688 & n5001 ) | ( n4688 & ~n5002 ) | ( n5001 & ~n5002 ) ;
  assign n5004 = ( n1435 & ~n5001 ) | ( n1435 & n5002 ) | ( ~n5001 & n5002 ) ;
  assign n5005 = ( n5000 & ~n5003 ) | ( n5000 & n5004 ) | ( ~n5003 & n5004 ) ;
  assign n5006 = ~n292 & n2934 ;
  assign n5007 = ( n1468 & ~n2941 ) | ( n1468 & n5006 ) | ( ~n2941 & n5006 ) ;
  assign n5008 = ( n2494 & n2941 ) | ( n2494 & ~n5006 ) | ( n2941 & ~n5006 ) ;
  assign n5009 = ( n5005 & ~n5007 ) | ( n5005 & n5008 ) | ( ~n5007 & n5008 ) ;
  assign n5010 = ( n416 & n461 ) | ( n416 & ~n1506 ) | ( n461 & ~n1506 ) ;
  assign n5011 = ~n333 & n3382 ;
  assign n5012 = ( n376 & ~n3835 ) | ( n376 & n3840 ) | ( ~n3835 & n3840 ) ;
  assign n5013 = ( n358 & ~n376 ) | ( n358 & n3947 ) | ( ~n376 & n3947 ) ;
  assign n5014 = ( n5011 & n5012 ) | ( n5011 & ~n5013 ) | ( n5012 & ~n5013 ) ;
  assign n5015 = ( n4397 & ~n5010 ) | ( n4397 & n5014 ) | ( ~n5010 & n5014 ) ;
  assign n5016 = ( n4491 & ~n5012 ) | ( n4491 & n5013 ) | ( ~n5012 & n5013 ) ;
  assign n5017 = ( ~n4397 & n5010 ) | ( ~n4397 & n5016 ) | ( n5010 & n5016 ) ;
  assign n5018 = ( n5009 & n5015 ) | ( n5009 & ~n5017 ) | ( n5015 & ~n5017 ) ;
  assign n5019 = x214 & ~n544 ;
  assign n5020 = n549 | n2034 ;
  assign n5021 = ~n490 & n1793 ;
  assign n5022 = ( n1517 & n2025 ) | ( n1517 & ~n5021 ) | ( n2025 & ~n5021 ) ;
  assign n5023 = ~n484 & n5022 ;
  assign n5024 = ( n3398 & ~n5020 ) | ( n3398 & n5023 ) | ( ~n5020 & n5023 ) ;
  assign n5025 = n5019 & ~n5024 ;
  assign n5026 = ( ~n514 & n1513 ) | ( ~n514 & n2020 ) | ( n1513 & n2020 ) ;
  assign n5027 = ( ~n3398 & n5020 ) | ( ~n3398 & n5026 ) | ( n5020 & n5026 ) ;
  assign n5028 = n5019 & n5027 ;
  assign n5029 = ( n5018 & n5025 ) | ( n5018 & n5028 ) | ( n5025 & n5028 ) ;
  assign n5030 = x89 | n956 ;
  assign n5031 = ~n542 & n5030 ;
  assign n5032 = ( ~n534 & n538 ) | ( ~n534 & n5031 ) | ( n538 & n5031 ) ;
  assign n5033 = ( ~n560 & n1532 ) | ( ~n560 & n5032 ) | ( n1532 & n5032 ) ;
  assign n5034 = ( n1531 & ~n2238 ) | ( n1531 & n5033 ) | ( ~n2238 & n5033 ) ;
  assign n5035 = n655 | n2243 ;
  assign n5036 = ( ~n655 & n1551 ) | ( ~n655 & n2055 ) | ( n1551 & n2055 ) ;
  assign n5037 = ( n4723 & n5035 ) | ( n4723 & ~n5036 ) | ( n5035 & ~n5036 ) ;
  assign n5038 = ( n1553 & ~n5035 ) | ( n1553 & n5036 ) | ( ~n5035 & n5036 ) ;
  assign n5039 = ( n5034 & ~n5037 ) | ( n5034 & n5038 ) | ( ~n5037 & n5038 ) ;
  assign n5040 = ~n697 & n2969 ;
  assign n5041 = ( n1567 & ~n2977 ) | ( n1567 & n5040 ) | ( ~n2977 & n5040 ) ;
  assign n5042 = ( n2531 & n2977 ) | ( n2531 & ~n5040 ) | ( n2977 & ~n5040 ) ;
  assign n5043 = ( n5039 & ~n5041 ) | ( n5039 & n5042 ) | ( ~n5041 & n5042 ) ;
  assign n5044 = ( n821 & n866 ) | ( n821 & ~n1605 ) | ( n866 & ~n1605 ) ;
  assign n5045 = ~n738 & n3421 ;
  assign n5046 = ( n781 & ~n3873 ) | ( n781 & n3878 ) | ( ~n3873 & n3878 ) ;
  assign n5047 = ( n763 & ~n781 ) | ( n763 & n3985 ) | ( ~n781 & n3985 ) ;
  assign n5048 = ( n5045 & n5046 ) | ( n5045 & ~n5047 ) | ( n5046 & ~n5047 ) ;
  assign n5049 = ( n4433 & ~n5044 ) | ( n4433 & n5048 ) | ( ~n5044 & n5048 ) ;
  assign n5050 = ( n4526 & ~n5046 ) | ( n4526 & n5047 ) | ( ~n5046 & n5047 ) ;
  assign n5051 = ( ~n4433 & n5044 ) | ( ~n4433 & n5050 ) | ( n5044 & n5050 ) ;
  assign n5052 = ( n5043 & n5049 ) | ( n5043 & ~n5051 ) | ( n5049 & ~n5051 ) ;
  assign n5053 = x215 & ~n949 ;
  assign n5054 = n954 | n2104 ;
  assign n5055 = ~n895 & n1871 ;
  assign n5056 = ( n1616 & n2095 ) | ( n1616 & ~n5055 ) | ( n2095 & ~n5055 ) ;
  assign n5057 = ~n889 & n5056 ;
  assign n5058 = ( n3437 & ~n5054 ) | ( n3437 & n5057 ) | ( ~n5054 & n5057 ) ;
  assign n5059 = n5053 & ~n5058 ;
  assign n5060 = ( ~n919 & n1612 ) | ( ~n919 & n2090 ) | ( n1612 & n2090 ) ;
  assign n5061 = ( ~n3437 & n5054 ) | ( ~n3437 & n5060 ) | ( n5054 & n5060 ) ;
  assign n5062 = n5053 & n5061 ;
  assign n5063 = ( n5052 & n5059 ) | ( n5052 & n5062 ) | ( n5059 & n5062 ) ;
  assign n5064 = x90 | n1360 ;
  assign n5065 = ~n947 & n5064 ;
  assign n5066 = ( ~n939 & n943 ) | ( ~n939 & n5065 ) | ( n943 & n5065 ) ;
  assign n5067 = ( ~n965 & n1631 ) | ( ~n965 & n5066 ) | ( n1631 & n5066 ) ;
  assign n5068 = ( n1630 & ~n2294 ) | ( n1630 & n5067 ) | ( ~n2294 & n5067 ) ;
  assign n5069 = n1060 | n2299 ;
  assign n5070 = ( ~n1060 & n1650 ) | ( ~n1060 & n2125 ) | ( n1650 & n2125 ) ;
  assign n5071 = ( n4758 & n5069 ) | ( n4758 & ~n5070 ) | ( n5069 & ~n5070 ) ;
  assign n5072 = ( n1652 & ~n5069 ) | ( n1652 & n5070 ) | ( ~n5069 & n5070 ) ;
  assign n5073 = ( n5068 & ~n5071 ) | ( n5068 & n5072 ) | ( ~n5071 & n5072 ) ;
  assign n5074 = ~n1101 & n3005 ;
  assign n5075 = ( n1666 & ~n3013 ) | ( n1666 & n5074 ) | ( ~n3013 & n5074 ) ;
  assign n5076 = ( n2568 & n3013 ) | ( n2568 & ~n5074 ) | ( n3013 & ~n5074 ) ;
  assign n5077 = ( n5073 & ~n5075 ) | ( n5073 & n5076 ) | ( ~n5075 & n5076 ) ;
  assign n5078 = ( n1225 & n1270 ) | ( n1225 & ~n1703 ) | ( n1270 & ~n1703 ) ;
  assign n5079 = ~n1142 & n3460 ;
  assign n5080 = ( n1185 & ~n3911 ) | ( n1185 & n3916 ) | ( ~n3911 & n3916 ) ;
  assign n5081 = ( n1167 & ~n1185 ) | ( n1167 & n4023 ) | ( ~n1185 & n4023 ) ;
  assign n5082 = ( n5079 & n5080 ) | ( n5079 & ~n5081 ) | ( n5080 & ~n5081 ) ;
  assign n5083 = ( n4469 & ~n5078 ) | ( n4469 & n5082 ) | ( ~n5078 & n5082 ) ;
  assign n5084 = ( n4561 & ~n5080 ) | ( n4561 & n5081 ) | ( ~n5080 & n5081 ) ;
  assign n5085 = ( ~n4469 & n5078 ) | ( ~n4469 & n5084 ) | ( n5078 & n5084 ) ;
  assign n5086 = ( n5077 & n5083 ) | ( n5077 & ~n5085 ) | ( n5083 & ~n5085 ) ;
  assign n5087 = x216 & ~n1353 ;
  assign n5088 = n1358 | n2174 ;
  assign n5089 = ~n1299 & n1949 ;
  assign n5090 = ( n1714 & n2165 ) | ( n1714 & ~n5089 ) | ( n2165 & ~n5089 ) ;
  assign n5091 = ~n1293 & n5090 ;
  assign n5092 = ( n3476 & ~n5088 ) | ( n3476 & n5091 ) | ( ~n5088 & n5091 ) ;
  assign n5093 = n5087 & ~n5092 ;
  assign n5094 = ( ~n1323 & n1710 ) | ( ~n1323 & n2160 ) | ( n1710 & n2160 ) ;
  assign n5095 = ( ~n3476 & n5088 ) | ( ~n3476 & n5094 ) | ( n5088 & n5094 ) ;
  assign n5096 = n5087 & n5095 ;
  assign n5097 = ( n5086 & n5093 ) | ( n5086 & n5096 ) | ( n5093 & n5096 ) ;
  assign n5098 = x91 | n535 ;
  assign n5099 = ~n1351 & n5098 ;
  assign n5100 = ( ~n1343 & n1347 ) | ( ~n1343 & n5099 ) | ( n1347 & n5099 ) ;
  assign n5101 = ( ~n1369 & n1729 ) | ( ~n1369 & n5100 ) | ( n1729 & n5100 ) ;
  assign n5102 = ( n1728 & ~n2350 ) | ( n1728 & n5101 ) | ( ~n2350 & n5101 ) ;
  assign n5103 = n1464 | n2355 ;
  assign n5104 = ( ~n1464 & n1748 ) | ( ~n1464 & n2195 ) | ( n1748 & n2195 ) ;
  assign n5105 = ( n4793 & n5103 ) | ( n4793 & ~n5104 ) | ( n5103 & ~n5104 ) ;
  assign n5106 = ( n1750 & ~n5103 ) | ( n1750 & n5104 ) | ( ~n5103 & n5104 ) ;
  assign n5107 = ( n5102 & ~n5105 ) | ( n5102 & n5106 ) | ( ~n5105 & n5106 ) ;
  assign n5108 = ~n286 & n3042 ;
  assign n5109 = ( n1761 & ~n3049 ) | ( n1761 & n5108 ) | ( ~n3049 & n5108 ) ;
  assign n5110 = ( n2604 & n3049 ) | ( n2604 & ~n5108 ) | ( n3049 & ~n5108 ) ;
  assign n5111 = ( n5107 & ~n5109 ) | ( n5107 & n5110 ) | ( ~n5109 & n5110 ) ;
  assign n5112 = ( n462 & n1504 ) | ( n462 & ~n1789 ) | ( n1504 & ~n1789 ) ;
  assign n5113 = ~n340 & n3498 ;
  assign n5114 = ( n1496 & ~n3949 ) | ( n1496 & n3954 ) | ( ~n3949 & n3954 ) ;
  assign n5115 = ( n398 & ~n1496 ) | ( n398 & n4061 ) | ( ~n1496 & n4061 ) ;
  assign n5116 = ( n5113 & n5114 ) | ( n5113 & ~n5115 ) | ( n5114 & ~n5115 ) ;
  assign n5117 = ( n4504 & ~n5112 ) | ( n4504 & n5116 ) | ( ~n5112 & n5116 ) ;
  assign n5118 = ( n4596 & ~n5114 ) | ( n4596 & n5115 ) | ( ~n5114 & n5115 ) ;
  assign n5119 = ( ~n4504 & n5112 ) | ( ~n4504 & n5118 ) | ( n5112 & n5118 ) ;
  assign n5120 = ( n5111 & n5117 ) | ( n5111 & ~n5119 ) | ( n5117 & ~n5119 ) ;
  assign n5121 = x217 & ~n541 ;
  assign n5122 = n553 | n2230 ;
  assign n5123 = ~n481 & n2020 ;
  assign n5124 = ( n1799 & n2221 ) | ( n1799 & ~n5123 ) | ( n2221 & ~n5123 ) ;
  assign n5125 = ~n478 & n5124 ;
  assign n5126 = ( n3515 & ~n5122 ) | ( n3515 & n5125 ) | ( ~n5122 & n5125 ) ;
  assign n5127 = n5121 & ~n5126 ;
  assign n5128 = ( n486 & ~n1526 ) | ( n486 & n1795 ) | ( ~n1526 & n1795 ) ;
  assign n5129 = ( ~n3515 & n5122 ) | ( ~n3515 & n5128 ) | ( n5122 & n5128 ) ;
  assign n5130 = n5121 & n5129 ;
  assign n5131 = ( n5120 & n5127 ) | ( n5120 & n5130 ) | ( n5127 & n5130 ) ;
  assign n5132 = x92 | n940 ;
  assign n5133 = ~n533 & n5132 ;
  assign n5134 = ( ~n559 & n566 ) | ( ~n559 & n5133 ) | ( n566 & n5133 ) ;
  assign n5135 = ( n528 & ~n564 ) | ( n528 & n5134 ) | ( ~n564 & n5134 ) ;
  assign n5136 = ( ~n612 & n1811 ) | ( ~n612 & n5135 ) | ( n1811 & n5135 ) ;
  assign n5137 = n641 | n2399 ;
  assign n5138 = ( ~n641 & n645 ) | ( ~n641 & n2249 ) | ( n645 & n2249 ) ;
  assign n5139 = ( n4828 & n5137 ) | ( n4828 & ~n5138 ) | ( n5137 & ~n5138 ) ;
  assign n5140 = ( n1829 & ~n5137 ) | ( n1829 & n5138 ) | ( ~n5137 & n5138 ) ;
  assign n5141 = ( n5136 & ~n5139 ) | ( n5136 & n5140 ) | ( ~n5139 & n5140 ) ;
  assign n5142 = ~n691 & n3077 ;
  assign n5143 = ( n2639 & n3085 ) | ( n2639 & ~n5142 ) | ( n3085 & ~n5142 ) ;
  assign n5144 = ( n1839 & ~n3085 ) | ( n1839 & n5142 ) | ( ~n3085 & n5142 ) ;
  assign n5145 = ( n5141 & n5143 ) | ( n5141 & ~n5144 ) | ( n5143 & ~n5144 ) ;
  assign n5146 = ( n867 & n1603 ) | ( n867 & ~n1867 ) | ( n1603 & ~n1867 ) ;
  assign n5147 = ~n745 & n3536 ;
  assign n5148 = ( n1595 & ~n3987 ) | ( n1595 & n3992 ) | ( ~n3987 & n3992 ) ;
  assign n5149 = ( n803 & ~n1595 ) | ( n803 & n4098 ) | ( ~n1595 & n4098 ) ;
  assign n5150 = ( n5147 & n5148 ) | ( n5147 & ~n5149 ) | ( n5148 & ~n5149 ) ;
  assign n5151 = ( n4539 & ~n5146 ) | ( n4539 & n5150 ) | ( ~n5146 & n5150 ) ;
  assign n5152 = ( n4631 & ~n5148 ) | ( n4631 & n5149 ) | ( ~n5148 & n5149 ) ;
  assign n5153 = ( ~n4539 & n5146 ) | ( ~n4539 & n5152 ) | ( n5146 & n5152 ) ;
  assign n5154 = ( n5145 & n5151 ) | ( n5145 & ~n5153 ) | ( n5151 & ~n5153 ) ;
  assign n5155 = x218 & ~n946 ;
  assign n5156 = n958 | n2286 ;
  assign n5157 = ~n886 & n2090 ;
  assign n5158 = ( n1877 & n2277 ) | ( n1877 & ~n5157 ) | ( n2277 & ~n5157 ) ;
  assign n5159 = ~n883 & n5158 ;
  assign n5160 = ( n3553 & ~n5156 ) | ( n3553 & n5159 ) | ( ~n5156 & n5159 ) ;
  assign n5161 = n5155 & ~n5160 ;
  assign n5162 = ( n891 & ~n1625 ) | ( n891 & n1873 ) | ( ~n1625 & n1873 ) ;
  assign n5163 = ( ~n3553 & n5156 ) | ( ~n3553 & n5162 ) | ( n5156 & n5162 ) ;
  assign n5164 = n5155 & n5163 ;
  assign n5165 = ( n5154 & n5161 ) | ( n5154 & n5164 ) | ( n5161 & n5164 ) ;
  assign n5166 = x93 | n1344 ;
  assign n5167 = ~n938 & n5166 ;
  assign n5168 = ( ~n964 & n971 ) | ( ~n964 & n5167 ) | ( n971 & n5167 ) ;
  assign n5169 = ( n933 & ~n969 ) | ( n933 & n5168 ) | ( ~n969 & n5168 ) ;
  assign n5170 = ( ~n1017 & n1889 ) | ( ~n1017 & n5169 ) | ( n1889 & n5169 ) ;
  assign n5171 = n1046 | n2443 ;
  assign n5172 = ( ~n1046 & n1050 ) | ( ~n1046 & n2305 ) | ( n1050 & n2305 ) ;
  assign n5173 = ( n4863 & n5171 ) | ( n4863 & ~n5172 ) | ( n5171 & ~n5172 ) ;
  assign n5174 = ( n1907 & ~n5171 ) | ( n1907 & n5172 ) | ( ~n5171 & n5172 ) ;
  assign n5175 = ( n5170 & ~n5173 ) | ( n5170 & n5174 ) | ( ~n5173 & n5174 ) ;
  assign n5176 = ~n1095 & n3113 ;
  assign n5177 = ( n2674 & n3121 ) | ( n2674 & ~n5176 ) | ( n3121 & ~n5176 ) ;
  assign n5178 = ( n1917 & ~n3121 ) | ( n1917 & n5176 ) | ( ~n3121 & n5176 ) ;
  assign n5179 = ( n5175 & n5177 ) | ( n5175 & ~n5178 ) | ( n5177 & ~n5178 ) ;
  assign n5180 = ( n1271 & n1701 ) | ( n1271 & ~n1945 ) | ( n1701 & ~n1945 ) ;
  assign n5181 = ~n1149 & n3574 ;
  assign n5182 = ( n1693 & ~n4025 ) | ( n1693 & n4030 ) | ( ~n4025 & n4030 ) ;
  assign n5183 = ( n1207 & ~n1693 ) | ( n1207 & n4135 ) | ( ~n1693 & n4135 ) ;
  assign n5184 = ( n5181 & n5182 ) | ( n5181 & ~n5183 ) | ( n5182 & ~n5183 ) ;
  assign n5185 = ( n4574 & ~n5180 ) | ( n4574 & n5184 ) | ( ~n5180 & n5184 ) ;
  assign n5186 = ( n4666 & ~n5182 ) | ( n4666 & n5183 ) | ( ~n5182 & n5183 ) ;
  assign n5187 = ( ~n4574 & n5180 ) | ( ~n4574 & n5186 ) | ( n5180 & n5186 ) ;
  assign n5188 = ( n5179 & n5185 ) | ( n5179 & ~n5187 ) | ( n5185 & ~n5187 ) ;
  assign n5189 = x219 & ~n1350 ;
  assign n5190 = n1362 | n2342 ;
  assign n5191 = ~n1290 & n2160 ;
  assign n5192 = ( n1955 & n2333 ) | ( n1955 & ~n5191 ) | ( n2333 & ~n5191 ) ;
  assign n5193 = ~n1287 & n5192 ;
  assign n5194 = ( n3591 & ~n5190 ) | ( n3591 & n5193 ) | ( ~n5190 & n5193 ) ;
  assign n5195 = n5189 & ~n5194 ;
  assign n5196 = ( n1295 & ~n1723 ) | ( n1295 & n1951 ) | ( ~n1723 & n1951 ) ;
  assign n5197 = ( ~n3591 & n5190 ) | ( ~n3591 & n5196 ) | ( n5190 & n5196 ) ;
  assign n5198 = n5189 & n5197 ;
  assign n5199 = ( n5188 & n5195 ) | ( n5188 & n5198 ) | ( n5195 & n5198 ) ;
  assign n5200 = x94 | n529 ;
  assign n5201 = ~n1342 & n5200 ;
  assign n5202 = ( ~n1368 & n1375 ) | ( ~n1368 & n5201 ) | ( n1375 & n5201 ) ;
  assign n5203 = ( n1337 & ~n1373 ) | ( n1337 & n5202 ) | ( ~n1373 & n5202 ) ;
  assign n5204 = ( ~n1421 & n1967 ) | ( ~n1421 & n5203 ) | ( n1967 & n5203 ) ;
  assign n5205 = n1450 | n2487 ;
  assign n5206 = ( ~n1450 & n1454 ) | ( ~n1450 & n2361 ) | ( n1454 & n2361 ) ;
  assign n5207 = ( n4898 & n5205 ) | ( n4898 & ~n5206 ) | ( n5205 & ~n5206 ) ;
  assign n5208 = ( n1985 & ~n5205 ) | ( n1985 & n5206 ) | ( ~n5205 & n5206 ) ;
  assign n5209 = ( n5204 & ~n5207 ) | ( n5204 & n5208 ) | ( ~n5207 & n5208 ) ;
  assign n5210 = ~n310 & n3149 ;
  assign n5211 = ( n2709 & n3157 ) | ( n2709 & ~n5210 ) | ( n3157 & ~n5210 ) ;
  assign n5212 = ( n1993 & ~n3157 ) | ( n1993 & n5210 ) | ( ~n3157 & n5210 ) ;
  assign n5213 = ( n5209 & n5211 ) | ( n5209 & ~n5212 ) | ( n5211 & ~n5212 ) ;
  assign n5214 = ( n464 & n1787 ) | ( n464 & ~n2016 ) | ( n1787 & ~n2016 ) ;
  assign n5215 = ~n327 & n3612 ;
  assign n5216 = ( n384 & n420 ) | ( n384 & ~n4063 ) | ( n420 & ~n4063 ) ;
  assign n5217 = ( n408 & ~n420 ) | ( n408 & n4172 ) | ( ~n420 & n4172 ) ;
  assign n5218 = ( n5215 & n5216 ) | ( n5215 & ~n5217 ) | ( n5216 & ~n5217 ) ;
  assign n5219 = ( n4609 & ~n5214 ) | ( n4609 & n5218 ) | ( ~n5214 & n5218 ) ;
  assign n5220 = ( n4701 & ~n5216 ) | ( n4701 & n5217 ) | ( ~n5216 & n5217 ) ;
  assign n5221 = ( ~n4609 & n5214 ) | ( ~n4609 & n5220 ) | ( n5214 & n5220 ) ;
  assign n5222 = ( n5213 & n5219 ) | ( n5213 & ~n5221 ) | ( n5219 & ~n5221 ) ;
  assign n5223 = x220 & ~n532 ;
  assign n5224 = n537 | n555 ;
  assign n5225 = n486 & ~n506 ;
  assign n5226 = ( n510 & n2026 ) | ( n510 & ~n5225 ) | ( n2026 & ~n5225 ) ;
  assign n5227 = ~n474 & n5226 ;
  assign n5228 = ( n3628 & ~n5224 ) | ( n3628 & n5227 ) | ( ~n5224 & n5227 ) ;
  assign n5229 = n5223 & ~n5228 ;
  assign n5230 = ( n1520 & ~n1807 ) | ( n1520 & n2022 ) | ( ~n1807 & n2022 ) ;
  assign n5231 = ( ~n3628 & n5224 ) | ( ~n3628 & n5230 ) | ( n5224 & n5230 ) ;
  assign n5232 = n5223 & n5231 ;
  assign n5233 = ( n5222 & n5229 ) | ( n5222 & n5232 ) | ( n5229 & n5232 ) ;
  assign n5234 = x95 | n934 ;
  assign n5235 = ~n558 & n5234 ;
  assign n5236 = ( ~n523 & n527 ) | ( ~n523 & n5235 ) | ( n527 & n5235 ) ;
  assign n5237 = ( ~n604 & n1531 ) | ( ~n604 & n5236 ) | ( n1531 & n5236 ) ;
  assign n5238 = ( ~n1543 & n2038 ) | ( ~n1543 & n5237 ) | ( n2038 & n5237 ) ;
  assign n5239 = n638 | n658 ;
  assign n5240 = ( ~n638 & n649 ) | ( ~n638 & n2405 ) | ( n649 & n2405 ) ;
  assign n5241 = ( n4933 & n5239 ) | ( n4933 & ~n5240 ) | ( n5239 & ~n5240 ) ;
  assign n5242 = ( n2055 & ~n5239 ) | ( n2055 & n5240 ) | ( ~n5239 & n5240 ) ;
  assign n5243 = ( n5238 & ~n5241 ) | ( n5238 & n5242 ) | ( ~n5241 & n5242 ) ;
  assign n5244 = ~n715 & n3185 ;
  assign n5245 = ( n2063 & ~n3193 ) | ( n2063 & n5244 ) | ( ~n3193 & n5244 ) ;
  assign n5246 = ( n2753 & n3193 ) | ( n2753 & ~n5244 ) | ( n3193 & ~n5244 ) ;
  assign n5247 = ( n5243 & ~n5245 ) | ( n5243 & n5246 ) | ( ~n5245 & n5246 ) ;
  assign n5248 = ( n869 & n1865 ) | ( n869 & ~n2086 ) | ( n1865 & ~n2086 ) ;
  assign n5249 = ~n732 & n3650 ;
  assign n5250 = ( n789 & n825 ) | ( n789 & ~n4100 ) | ( n825 & ~n4100 ) ;
  assign n5251 = ( n813 & ~n825 ) | ( n813 & n4209 ) | ( ~n825 & n4209 ) ;
  assign n5252 = ( n5249 & n5250 ) | ( n5249 & ~n5251 ) | ( n5250 & ~n5251 ) ;
  assign n5253 = ( n4644 & ~n5248 ) | ( n4644 & n5252 ) | ( ~n5248 & n5252 ) ;
  assign n5254 = ( n4736 & ~n5250 ) | ( n4736 & n5251 ) | ( ~n5250 & n5251 ) ;
  assign n5255 = ( ~n4644 & n5248 ) | ( ~n4644 & n5254 ) | ( n5248 & n5254 ) ;
  assign n5256 = ( n5247 & n5253 ) | ( n5247 & ~n5255 ) | ( n5253 & ~n5255 ) ;
  assign n5257 = x221 & ~n937 ;
  assign n5258 = n942 | n960 ;
  assign n5259 = n891 & ~n911 ;
  assign n5260 = ( n915 & n2096 ) | ( n915 & ~n5259 ) | ( n2096 & ~n5259 ) ;
  assign n5261 = ~n879 & n5260 ;
  assign n5262 = ( n3666 & ~n5258 ) | ( n3666 & n5261 ) | ( ~n5258 & n5261 ) ;
  assign n5263 = n5257 & ~n5262 ;
  assign n5264 = ( n1619 & ~n1885 ) | ( n1619 & n2092 ) | ( ~n1885 & n2092 ) ;
  assign n5265 = ( ~n3666 & n5258 ) | ( ~n3666 & n5264 ) | ( n5258 & n5264 ) ;
  assign n5266 = n5257 & n5265 ;
  assign n5267 = ( n5256 & n5263 ) | ( n5256 & n5266 ) | ( n5263 & n5266 ) ;
  assign n5268 = x96 | n1338 ;
  assign n5269 = ~n963 & n5268 ;
  assign n5270 = ( ~n928 & n932 ) | ( ~n928 & n5269 ) | ( n932 & n5269 ) ;
  assign n5271 = ( ~n1009 & n1630 ) | ( ~n1009 & n5270 ) | ( n1630 & n5270 ) ;
  assign n5272 = ( ~n1642 & n2108 ) | ( ~n1642 & n5271 ) | ( n2108 & n5271 ) ;
  assign n5273 = n1043 | n1063 ;
  assign n5274 = ( ~n1043 & n1054 ) | ( ~n1043 & n2449 ) | ( n1054 & n2449 ) ;
  assign n5275 = ( n4967 & n5273 ) | ( n4967 & ~n5274 ) | ( n5273 & ~n5274 ) ;
  assign n5276 = ( n2125 & ~n5273 ) | ( n2125 & n5274 ) | ( ~n5273 & n5274 ) ;
  assign n5277 = ( n5272 & ~n5275 ) | ( n5272 & n5276 ) | ( ~n5275 & n5276 ) ;
  assign n5278 = ~n1119 & n3221 ;
  assign n5279 = ( n2133 & ~n3229 ) | ( n2133 & n5278 ) | ( ~n3229 & n5278 ) ;
  assign n5280 = ( n2792 & n3229 ) | ( n2792 & ~n5278 ) | ( n3229 & ~n5278 ) ;
  assign n5281 = ( n5277 & ~n5279 ) | ( n5277 & n5280 ) | ( ~n5279 & n5280 ) ;
  assign n5282 = ( n1273 & n1943 ) | ( n1273 & ~n2156 ) | ( n1943 & ~n2156 ) ;
  assign n5283 = ~n1136 & n3688 ;
  assign n5284 = ( n1193 & n1229 ) | ( n1193 & ~n4137 ) | ( n1229 & ~n4137 ) ;
  assign n5285 = ( n1217 & ~n1229 ) | ( n1217 & n4246 ) | ( ~n1229 & n4246 ) ;
  assign n5286 = ( n5283 & n5284 ) | ( n5283 & ~n5285 ) | ( n5284 & ~n5285 ) ;
  assign n5287 = ( n4679 & ~n5282 ) | ( n4679 & n5286 ) | ( ~n5282 & n5286 ) ;
  assign n5288 = ( n4771 & ~n5284 ) | ( n4771 & n5285 ) | ( ~n5284 & n5285 ) ;
  assign n5289 = ( ~n4679 & n5282 ) | ( ~n4679 & n5288 ) | ( n5282 & n5288 ) ;
  assign n5290 = ( n5281 & n5287 ) | ( n5281 & ~n5289 ) | ( n5287 & ~n5289 ) ;
  assign n5291 = x222 & ~n1341 ;
  assign n5292 = n1346 | n1364 ;
  assign n5293 = n1295 & ~n1315 ;
  assign n5294 = ( n1319 & n2166 ) | ( n1319 & ~n5293 ) | ( n2166 & ~n5293 ) ;
  assign n5295 = ~n1283 & n5294 ;
  assign n5296 = ( n3704 & ~n5292 ) | ( n3704 & n5295 ) | ( ~n5292 & n5295 ) ;
  assign n5297 = n5291 & ~n5296 ;
  assign n5298 = ( n1717 & ~n1963 ) | ( n1717 & n2162 ) | ( ~n1963 & n2162 ) ;
  assign n5299 = ( ~n3704 & n5292 ) | ( ~n3704 & n5298 ) | ( n5292 & n5298 ) ;
  assign n5300 = n5291 & n5299 ;
  assign n5301 = ( n5290 & n5297 ) | ( n5290 & n5300 ) | ( n5297 & n5300 ) ;
  assign n5302 = x97 | n524 ;
  assign n5303 = ~n1367 & n5302 ;
  assign n5304 = ( ~n1332 & n1336 ) | ( ~n1332 & n5303 ) | ( n1336 & n5303 ) ;
  assign n5305 = ( ~n1413 & n1728 ) | ( ~n1413 & n5304 ) | ( n1728 & n5304 ) ;
  assign n5306 = ( ~n1740 & n2178 ) | ( ~n1740 & n5305 ) | ( n2178 & n5305 ) ;
  assign n5307 = n1447 | n1467 ;
  assign n5308 = ( ~n1447 & n1458 ) | ( ~n1447 & n2493 ) | ( n1458 & n2493 ) ;
  assign n5309 = ( n5001 & n5307 ) | ( n5001 & ~n5308 ) | ( n5307 & ~n5308 ) ;
  assign n5310 = ( n2195 & ~n5307 ) | ( n2195 & n5308 ) | ( ~n5307 & n5308 ) ;
  assign n5311 = ( n5306 & ~n5309 ) | ( n5306 & n5310 ) | ( ~n5309 & n5310 ) ;
  assign n5312 = ~n314 & n3257 ;
  assign n5313 = ( n2202 & ~n3265 ) | ( n2202 & n5312 ) | ( ~n3265 & n5312 ) ;
  assign n5314 = ( n2830 & n3265 ) | ( n2830 & ~n5312 ) | ( n3265 & ~n5312 ) ;
  assign n5315 = ( n5311 & ~n5313 ) | ( n5311 & n5314 ) | ( ~n5313 & n5314 ) ;
  assign n5316 = ( ~n438 & n439 ) | ( ~n438 & n2014 ) | ( n439 & n2014 ) ;
  assign n5317 = ~n365 & n3726 ;
  assign n5318 = ( n421 & n1499 ) | ( n421 & ~n4174 ) | ( n1499 & ~n4174 ) ;
  assign n5319 = ( n413 & ~n421 ) | ( n413 & n4283 ) | ( ~n421 & n4283 ) ;
  assign n5320 = ( n5317 & n5318 ) | ( n5317 & ~n5319 ) | ( n5318 & ~n5319 ) ;
  assign n5321 = ( n4714 & ~n5316 ) | ( n4714 & n5320 ) | ( ~n5316 & n5320 ) ;
  assign n5322 = ( n4806 & ~n5318 ) | ( n4806 & n5319 ) | ( ~n5318 & n5319 ) ;
  assign n5323 = ( ~n4714 & n5316 ) | ( ~n4714 & n5322 ) | ( n5316 & n5322 ) ;
  assign n5324 = ( n5315 & n5321 ) | ( n5315 & ~n5323 ) | ( n5321 & ~n5323 ) ;
  assign n5325 = x223 & ~n557 ;
  assign n5326 = n531 | n1533 ;
  assign n5327 = ~n471 & n1520 ;
  assign n5328 = ( n508 & n2223 ) | ( n508 & ~n5327 ) | ( n2223 & ~n5327 ) ;
  assign n5329 = ~n549 & n5328 ;
  assign n5330 = ( n3742 & ~n5326 ) | ( n3742 & n5329 ) | ( ~n5326 & n5329 ) ;
  assign n5331 = n5325 & ~n5330 ;
  assign n5332 = ( n503 & n1803 ) | ( n503 & ~n2029 ) | ( n1803 & ~n2029 ) ;
  assign n5333 = ( ~n3742 & n5326 ) | ( ~n3742 & n5332 ) | ( n5326 & n5332 ) ;
  assign n5334 = n5325 & n5333 ;
  assign n5335 = ( n5324 & n5331 ) | ( n5324 & n5334 ) | ( n5331 & n5334 ) ;
  assign n5336 = x98 | n929 ;
  assign n5337 = ~n522 & n5336 ;
  assign n5338 = ( ~n600 & n1530 ) | ( ~n600 & n5337 ) | ( n1530 & n5337 ) ;
  assign n5339 = ( ~n611 & n1811 ) | ( ~n611 & n5338 ) | ( n1811 & n5338 ) ;
  assign n5340 = ( n622 & ~n1821 ) | ( n622 & n5339 ) | ( ~n1821 & n5339 ) ;
  assign n5341 = n1561 | n1566 ;
  assign n5342 = ( n650 & ~n1561 ) | ( n650 & n1562 ) | ( ~n1561 & n1562 ) ;
  assign n5343 = ( n5035 & n5341 ) | ( n5035 & ~n5342 ) | ( n5341 & ~n5342 ) ;
  assign n5344 = ( n2249 & ~n5341 ) | ( n2249 & n5342 ) | ( ~n5341 & n5342 ) ;
  assign n5345 = ( n5340 & ~n5343 ) | ( n5340 & n5344 ) | ( ~n5343 & n5344 ) ;
  assign n5346 = ~n719 & n3296 ;
  assign n5347 = ( n2258 & ~n3304 ) | ( n2258 & n5346 ) | ( ~n3304 & n5346 ) ;
  assign n5348 = ( n2867 & n3304 ) | ( n2867 & ~n5346 ) | ( n3304 & ~n5346 ) ;
  assign n5349 = ( n5345 & ~n5347 ) | ( n5345 & n5348 ) | ( ~n5347 & n5348 ) ;
  assign n5350 = ( ~n843 & n844 ) | ( ~n843 & n2084 ) | ( n844 & n2084 ) ;
  assign n5351 = ~n770 & n3764 ;
  assign n5352 = ( n826 & n1598 ) | ( n826 & ~n4211 ) | ( n1598 & ~n4211 ) ;
  assign n5353 = ( n818 & ~n826 ) | ( n818 & n4319 ) | ( ~n826 & n4319 ) ;
  assign n5354 = ( n5351 & n5352 ) | ( n5351 & ~n5353 ) | ( n5352 & ~n5353 ) ;
  assign n5355 = ( n4749 & ~n5350 ) | ( n4749 & n5354 ) | ( ~n5350 & n5354 ) ;
  assign n5356 = ( n4841 & ~n5352 ) | ( n4841 & n5353 ) | ( ~n5352 & n5353 ) ;
  assign n5357 = ( ~n4749 & n5350 ) | ( ~n4749 & n5356 ) | ( n5350 & n5356 ) ;
  assign n5358 = ( n5349 & n5355 ) | ( n5349 & ~n5357 ) | ( n5355 & ~n5357 ) ;
  assign n5359 = x224 & ~n962 ;
  assign n5360 = n936 | n1632 ;
  assign n5361 = ~n876 & n1619 ;
  assign n5362 = ( n913 & n2279 ) | ( n913 & ~n5361 ) | ( n2279 & ~n5361 ) ;
  assign n5363 = ~n954 & n5362 ;
  assign n5364 = ( n3780 & ~n5360 ) | ( n3780 & n5363 ) | ( ~n5360 & n5363 ) ;
  assign n5365 = n5359 & ~n5364 ;
  assign n5366 = ( n908 & n1881 ) | ( n908 & ~n2099 ) | ( n1881 & ~n2099 ) ;
  assign n5367 = ( ~n3780 & n5360 ) | ( ~n3780 & n5366 ) | ( n5360 & n5366 ) ;
  assign n5368 = n5359 & n5367 ;
  assign n5369 = ( n5358 & n5365 ) | ( n5358 & n5368 ) | ( n5365 & n5368 ) ;
  assign n5370 = x99 | n1333 ;
  assign n5371 = ~n927 & n5370 ;
  assign n5372 = ( ~n1005 & n1629 ) | ( ~n1005 & n5371 ) | ( n1629 & n5371 ) ;
  assign n5373 = ( ~n1016 & n1889 ) | ( ~n1016 & n5372 ) | ( n1889 & n5372 ) ;
  assign n5374 = ( n1027 & ~n1899 ) | ( n1027 & n5373 ) | ( ~n1899 & n5373 ) ;
  assign n5375 = n1660 | n1665 ;
  assign n5376 = ( n1055 & ~n1660 ) | ( n1055 & n1661 ) | ( ~n1660 & n1661 ) ;
  assign n5377 = ( n5069 & n5375 ) | ( n5069 & ~n5376 ) | ( n5375 & ~n5376 ) ;
  assign n5378 = ( n2305 & ~n5375 ) | ( n2305 & n5376 ) | ( ~n5375 & n5376 ) ;
  assign n5379 = ( n5374 & ~n5377 ) | ( n5374 & n5378 ) | ( ~n5377 & n5378 ) ;
  assign n5380 = ~n1123 & n3335 ;
  assign n5381 = ( n2314 & ~n3343 ) | ( n2314 & n5380 ) | ( ~n3343 & n5380 ) ;
  assign n5382 = ( n2904 & n3343 ) | ( n2904 & ~n5380 ) | ( n3343 & ~n5380 ) ;
  assign n5383 = ( n5379 & ~n5381 ) | ( n5379 & n5382 ) | ( ~n5381 & n5382 ) ;
  assign n5384 = ( ~n1247 & n1248 ) | ( ~n1247 & n2154 ) | ( n1248 & n2154 ) ;
  assign n5385 = ~n1174 & n3802 ;
  assign n5386 = ( n1230 & n1696 ) | ( n1230 & ~n4248 ) | ( n1696 & ~n4248 ) ;
  assign n5387 = ( n1222 & ~n1230 ) | ( n1222 & n4355 ) | ( ~n1230 & n4355 ) ;
  assign n5388 = ( n5385 & n5386 ) | ( n5385 & ~n5387 ) | ( n5386 & ~n5387 ) ;
  assign n5389 = ( n4784 & ~n5384 ) | ( n4784 & n5388 ) | ( ~n5384 & n5388 ) ;
  assign n5390 = ( n4876 & ~n5386 ) | ( n4876 & n5387 ) | ( ~n5386 & n5387 ) ;
  assign n5391 = ( ~n4784 & n5384 ) | ( ~n4784 & n5390 ) | ( n5384 & n5390 ) ;
  assign n5392 = ( n5383 & n5389 ) | ( n5383 & ~n5391 ) | ( n5389 & ~n5391 ) ;
  assign n5393 = x225 & ~n1366 ;
  assign n5394 = n1340 | n1730 ;
  assign n5395 = ~n1280 & n1717 ;
  assign n5396 = ( n1317 & n2335 ) | ( n1317 & ~n5395 ) | ( n2335 & ~n5395 ) ;
  assign n5397 = ~n1358 & n5396 ;
  assign n5398 = ( n3818 & ~n5394 ) | ( n3818 & n5397 ) | ( ~n5394 & n5397 ) ;
  assign n5399 = n5393 & ~n5398 ;
  assign n5400 = ( n1312 & n1959 ) | ( n1312 & ~n2169 ) | ( n1959 & ~n2169 ) ;
  assign n5401 = ( ~n3818 & n5394 ) | ( ~n3818 & n5400 ) | ( n5394 & n5400 ) ;
  assign n5402 = n5393 & n5401 ;
  assign n5403 = ( n5392 & n5399 ) | ( n5392 & n5402 ) | ( n5399 & n5402 ) ;
  assign n5404 = x100 | n518 ;
  assign n5405 = ~n1331 & n5404 ;
  assign n5406 = ( ~n1409 & n1727 ) | ( ~n1409 & n5405 ) | ( n1727 & n5405 ) ;
  assign n5407 = ( ~n1420 & n1967 ) | ( ~n1420 & n5406 ) | ( n1967 & n5406 ) ;
  assign n5408 = ( n1431 & ~n1977 ) | ( n1431 & n5407 ) | ( ~n1977 & n5407 ) ;
  assign n5409 = n1755 | n1760 ;
  assign n5410 = ( n1459 & ~n1755 ) | ( n1459 & n1756 ) | ( ~n1755 & n1756 ) ;
  assign n5411 = ( n5103 & n5409 ) | ( n5103 & ~n5410 ) | ( n5409 & ~n5410 ) ;
  assign n5412 = ( n2361 & ~n5409 ) | ( n2361 & n5410 ) | ( ~n5409 & n5410 ) ;
  assign n5413 = ( n5408 & ~n5411 ) | ( n5408 & n5412 ) | ( ~n5411 & n5412 ) ;
  assign n5414 = ~n347 & n3374 ;
  assign n5415 = ( n2370 & ~n3382 ) | ( n2370 & n5414 ) | ( ~n3382 & n5414 ) ;
  assign n5416 = ( n2941 & n3382 ) | ( n2941 & ~n5414 ) | ( n3382 & ~n5414 ) ;
  assign n5417 = ( n5413 & ~n5415 ) | ( n5413 & n5416 ) | ( ~n5415 & n5416 ) ;
  assign n5418 = ( n466 & ~n1510 ) | ( n466 & n1511 ) | ( ~n1510 & n1511 ) ;
  assign n5419 = ~n372 & n3840 ;
  assign n5420 = ( n395 & ~n415 ) | ( n395 & n1783 ) | ( ~n415 & n1783 ) ;
  assign n5421 = ( n391 & ~n395 ) | ( n391 & n4391 ) | ( ~n395 & n4391 ) ;
  assign n5422 = ( n5419 & n5420 ) | ( n5419 & ~n5421 ) | ( n5420 & ~n5421 ) ;
  assign n5423 = ( n4819 & ~n5418 ) | ( n4819 & n5422 ) | ( ~n5418 & n5422 ) ;
  assign n5424 = ( n4911 & ~n5420 ) | ( n4911 & n5421 ) | ( ~n5420 & n5421 ) ;
  assign n5425 = ( ~n4819 & n5418 ) | ( ~n4819 & n5424 ) | ( n5418 & n5424 ) ;
  assign n5426 = ( n5417 & n5423 ) | ( n5417 & ~n5425 ) | ( n5423 & ~n5425 ) ;
  assign n5427 = x226 & ~n521 ;
  assign n5428 = n526 | n1812 ;
  assign n5429 = ~n546 & n1803 ;
  assign n5430 = ( n515 & n1524 ) | ( n515 & ~n5429 ) | ( n1524 & ~n5429 ) ;
  assign n5431 = ~n553 & n5430 ;
  assign n5432 = ( n3856 & ~n5428 ) | ( n3856 & n5431 ) | ( ~n5428 & n5431 ) ;
  assign n5433 = n5427 & ~n5432 ;
  assign n5434 = ( n1522 & n2033 ) | ( n1522 & ~n2226 ) | ( n2033 & ~n2226 ) ;
  assign n5435 = ( ~n3856 & n5428 ) | ( ~n3856 & n5434 ) | ( n5428 & n5434 ) ;
  assign n5436 = n5427 & n5435 ;
  assign n5437 = ( n5426 & n5433 ) | ( n5426 & n5436 ) | ( n5433 & n5436 ) ;
  assign n5438 = x101 | n923 ;
  assign n5439 = ~n599 & n5438 ;
  assign n5440 = ( ~n610 & n624 ) | ( ~n610 & n5439 ) | ( n624 & n5439 ) ;
  assign n5441 = ( ~n595 & n2038 ) | ( ~n595 & n5440 ) | ( n2038 & n5440 ) ;
  assign n5442 = ( n1552 & ~n2048 ) | ( n1552 & n5441 ) | ( ~n2048 & n5441 ) ;
  assign n5443 = n1833 | n1838 ;
  assign n5444 = ( n1563 & ~n1833 ) | ( n1563 & n1834 ) | ( ~n1833 & n1834 ) ;
  assign n5445 = ( n5137 & n5443 ) | ( n5137 & ~n5444 ) | ( n5443 & ~n5444 ) ;
  assign n5446 = ( n2405 & ~n5443 ) | ( n2405 & n5444 ) | ( ~n5443 & n5444 ) ;
  assign n5447 = ( n5442 & ~n5445 ) | ( n5442 & n5446 ) | ( ~n5445 & n5446 ) ;
  assign n5448 = ~n752 & n3413 ;
  assign n5449 = ( n2414 & ~n3421 ) | ( n2414 & n5448 ) | ( ~n3421 & n5448 ) ;
  assign n5450 = ( n2977 & n3421 ) | ( n2977 & ~n5448 ) | ( n3421 & ~n5448 ) ;
  assign n5451 = ( n5447 & ~n5449 ) | ( n5447 & n5450 ) | ( ~n5449 & n5450 ) ;
  assign n5452 = ( n871 & ~n1609 ) | ( n871 & n1610 ) | ( ~n1609 & n1610 ) ;
  assign n5453 = ~n777 & n3878 ;
  assign n5454 = ( n800 & ~n820 ) | ( n800 & n1861 ) | ( ~n820 & n1861 ) ;
  assign n5455 = ( n796 & ~n800 ) | ( n796 & n4427 ) | ( ~n800 & n4427 ) ;
  assign n5456 = ( n5453 & n5454 ) | ( n5453 & ~n5455 ) | ( n5454 & ~n5455 ) ;
  assign n5457 = ( n4854 & ~n5452 ) | ( n4854 & n5456 ) | ( ~n5452 & n5456 ) ;
  assign n5458 = ( n4945 & ~n5454 ) | ( n4945 & n5455 ) | ( ~n5454 & n5455 ) ;
  assign n5459 = ( ~n4854 & n5452 ) | ( ~n4854 & n5458 ) | ( n5452 & n5458 ) ;
  assign n5460 = ( n5451 & n5457 ) | ( n5451 & ~n5459 ) | ( n5457 & ~n5459 ) ;
  assign n5461 = x227 & ~n926 ;
  assign n5462 = n931 | n1890 ;
  assign n5463 = ~n951 & n1881 ;
  assign n5464 = ( n920 & n1623 ) | ( n920 & ~n5463 ) | ( n1623 & ~n5463 ) ;
  assign n5465 = ~n958 & n5464 ;
  assign n5466 = ( n3894 & ~n5462 ) | ( n3894 & n5465 ) | ( ~n5462 & n5465 ) ;
  assign n5467 = n5461 & ~n5466 ;
  assign n5468 = ( n1621 & n2103 ) | ( n1621 & ~n2282 ) | ( n2103 & ~n2282 ) ;
  assign n5469 = ( ~n3894 & n5462 ) | ( ~n3894 & n5468 ) | ( n5462 & n5468 ) ;
  assign n5470 = n5461 & n5469 ;
  assign n5471 = ( n5460 & n5467 ) | ( n5460 & n5470 ) | ( n5467 & n5470 ) ;
  assign n5472 = x102 | n1327 ;
  assign n5473 = ~n1004 & n5472 ;
  assign n5474 = ( ~n1015 & n1029 ) | ( ~n1015 & n5473 ) | ( n1029 & n5473 ) ;
  assign n5475 = ( ~n1000 & n2108 ) | ( ~n1000 & n5474 ) | ( n2108 & n5474 ) ;
  assign n5476 = ( n1651 & ~n2118 ) | ( n1651 & n5475 ) | ( ~n2118 & n5475 ) ;
  assign n5477 = n1911 | n1916 ;
  assign n5478 = ( n1662 & ~n1911 ) | ( n1662 & n1912 ) | ( ~n1911 & n1912 ) ;
  assign n5479 = ( n5171 & n5477 ) | ( n5171 & ~n5478 ) | ( n5477 & ~n5478 ) ;
  assign n5480 = ( n2449 & ~n5477 ) | ( n2449 & n5478 ) | ( ~n5477 & n5478 ) ;
  assign n5481 = ( n5476 & ~n5479 ) | ( n5476 & n5480 ) | ( ~n5479 & n5480 ) ;
  assign n5482 = ~n1156 & n3452 ;
  assign n5483 = ( n2458 & ~n3460 ) | ( n2458 & n5482 ) | ( ~n3460 & n5482 ) ;
  assign n5484 = ( n3013 & n3460 ) | ( n3013 & ~n5482 ) | ( n3460 & ~n5482 ) ;
  assign n5485 = ( n5481 & ~n5483 ) | ( n5481 & n5484 ) | ( ~n5483 & n5484 ) ;
  assign n5486 = ( n1275 & ~n1707 ) | ( n1275 & n1708 ) | ( ~n1707 & n1708 ) ;
  assign n5487 = ~n1181 & n3916 ;
  assign n5488 = ( n1204 & ~n1224 ) | ( n1204 & n1939 ) | ( ~n1224 & n1939 ) ;
  assign n5489 = ( n1200 & ~n1204 ) | ( n1200 & n4463 ) | ( ~n1204 & n4463 ) ;
  assign n5490 = ( n5487 & n5488 ) | ( n5487 & ~n5489 ) | ( n5488 & ~n5489 ) ;
  assign n5491 = ( n4889 & ~n5486 ) | ( n4889 & n5490 ) | ( ~n5486 & n5490 ) ;
  assign n5492 = ( n4979 & ~n5488 ) | ( n4979 & n5489 ) | ( ~n5488 & n5489 ) ;
  assign n5493 = ( ~n4889 & n5486 ) | ( ~n4889 & n5492 ) | ( n5486 & n5492 ) ;
  assign n5494 = ( n5485 & n5491 ) | ( n5485 & ~n5493 ) | ( n5491 & ~n5493 ) ;
  assign n5495 = x228 & ~n1330 ;
  assign n5496 = n1335 | n1968 ;
  assign n5497 = ~n1355 & n1959 ;
  assign n5498 = ( n1324 & n1721 ) | ( n1324 & ~n5497 ) | ( n1721 & ~n5497 ) ;
  assign n5499 = ~n1362 & n5498 ;
  assign n5500 = ( n3932 & ~n5496 ) | ( n3932 & n5499 ) | ( ~n5496 & n5499 ) ;
  assign n5501 = n5495 & ~n5500 ;
  assign n5502 = ( n1719 & n2173 ) | ( n1719 & ~n2338 ) | ( n2173 & ~n2338 ) ;
  assign n5503 = ( ~n3932 & n5496 ) | ( ~n3932 & n5502 ) | ( n5496 & n5502 ) ;
  assign n5504 = n5495 & n5503 ;
  assign n5505 = ( n5494 & n5501 ) | ( n5494 & n5504 ) | ( n5501 & n5504 ) ;
  assign n5506 = x103 | n601 ;
  assign n5507 = ~n1408 & n5506 ;
  assign n5508 = ( ~n1419 & n1433 ) | ( ~n1419 & n5507 ) | ( n1433 & n5507 ) ;
  assign n5509 = ( ~n1404 & n2178 ) | ( ~n1404 & n5508 ) | ( n2178 & n5508 ) ;
  assign n5510 = ( n1749 & ~n2188 ) | ( n1749 & n5509 ) | ( ~n2188 & n5509 ) ;
  assign n5511 = n265 | n1992 ;
  assign n5512 = ( ~n265 & n269 ) | ( ~n265 & n1757 ) | ( n269 & n1757 ) ;
  assign n5513 = ( n5205 & n5511 ) | ( n5205 & ~n5512 ) | ( n5511 & ~n5512 ) ;
  assign n5514 = ( n2493 & ~n5511 ) | ( n2493 & n5512 ) | ( ~n5511 & n5512 ) ;
  assign n5515 = ( n5510 & ~n5513 ) | ( n5510 & n5514 ) | ( ~n5513 & n5514 ) ;
  assign n5516 = ~n336 & n3491 ;
  assign n5517 = ( n2502 & ~n3498 ) | ( n2502 & n5516 ) | ( ~n3498 & n5516 ) ;
  assign n5518 = ( n3049 & n3498 ) | ( n3049 & ~n5516 ) | ( n3498 & ~n5516 ) ;
  assign n5519 = ( n5515 & ~n5517 ) | ( n5515 & n5518 ) | ( ~n5517 & n5518 ) ;
  assign n5520 = ( n512 & n1517 ) | ( n512 & ~n1793 ) | ( n1517 & ~n1793 ) ;
  assign n5521 = ~n358 & n3954 ;
  assign n5522 = ( n1501 & ~n1503 ) | ( n1501 & n2010 ) | ( ~n1503 & n2010 ) ;
  assign n5523 = ( n416 & n460 ) | ( n416 & ~n1501 ) | ( n460 & ~n1501 ) ;
  assign n5524 = ( n5521 & n5522 ) | ( n5521 & ~n5523 ) | ( n5522 & ~n5523 ) ;
  assign n5525 = ( n4924 & ~n5520 ) | ( n4924 & n5524 ) | ( ~n5520 & n5524 ) ;
  assign n5526 = ( n5013 & ~n5522 ) | ( n5013 & n5523 ) | ( ~n5522 & n5523 ) ;
  assign n5527 = ( ~n4924 & n5520 ) | ( ~n4924 & n5526 ) | ( n5520 & n5526 ) ;
  assign n5528 = ( n5519 & n5525 ) | ( n5519 & ~n5527 ) | ( n5525 & ~n5527 ) ;
  assign n5529 = x229 & ~n598 ;
  assign n5530 = n520 | n2039 ;
  assign n5531 = ~n543 & n2033 ;
  assign n5532 = ( n1527 & n1802 ) | ( n1527 & ~n5531 ) | ( n1802 & ~n5531 ) ;
  assign n5533 = ~n537 & n5532 ;
  assign n5534 = ( n3970 & ~n5530 ) | ( n3970 & n5533 ) | ( ~n5530 & n5533 ) ;
  assign n5535 = n5529 & ~n5534 ;
  assign n5536 = ( ~n569 & n1805 ) | ( ~n569 & n2229 ) | ( n1805 & n2229 ) ;
  assign n5537 = ( ~n3970 & n5530 ) | ( ~n3970 & n5536 ) | ( n5530 & n5536 ) ;
  assign n5538 = n5529 & n5537 ;
  assign n5539 = ( n5528 & n5535 ) | ( n5528 & n5538 ) | ( n5535 & n5538 ) ;
  assign n5540 = x104 | n1006 ;
  assign n5541 = ~n609 & n5540 ;
  assign n5542 = ( ~n591 & n625 ) | ( ~n591 & n5541 ) | ( n625 & n5541 ) ;
  assign n5543 = ( n622 & ~n623 ) | ( n622 & n5542 ) | ( ~n623 & n5542 ) ;
  assign n5544 = ( n1828 & ~n2243 ) | ( n1828 & n5543 ) | ( ~n2243 & n5543 ) ;
  assign n5545 = n670 | n2062 ;
  assign n5546 = ( ~n670 & n674 ) | ( ~n670 & n1835 ) | ( n674 & n1835 ) ;
  assign n5547 = ( n5239 & n5545 ) | ( n5239 & ~n5546 ) | ( n5545 & ~n5546 ) ;
  assign n5548 = ( n650 & ~n5545 ) | ( n650 & n5546 ) | ( ~n5545 & n5546 ) ;
  assign n5549 = ( n5544 & ~n5547 ) | ( n5544 & n5548 ) | ( ~n5547 & n5548 ) ;
  assign n5550 = ~n741 & n3529 ;
  assign n5551 = ( n2539 & ~n3536 ) | ( n2539 & n5550 ) | ( ~n3536 & n5550 ) ;
  assign n5552 = ( n3085 & n3536 ) | ( n3085 & ~n5550 ) | ( n3536 & ~n5550 ) ;
  assign n5553 = ( n5549 & ~n5551 ) | ( n5549 & n5552 ) | ( ~n5551 & n5552 ) ;
  assign n5554 = ( n917 & n1616 ) | ( n917 & ~n1871 ) | ( n1616 & ~n1871 ) ;
  assign n5555 = ~n763 & n3992 ;
  assign n5556 = ( n1600 & ~n1602 ) | ( n1600 & n2080 ) | ( ~n1602 & n2080 ) ;
  assign n5557 = ( n821 & n865 ) | ( n821 & ~n1600 ) | ( n865 & ~n1600 ) ;
  assign n5558 = ( n5555 & n5556 ) | ( n5555 & ~n5557 ) | ( n5556 & ~n5557 ) ;
  assign n5559 = ( n4958 & ~n5554 ) | ( n4958 & n5558 ) | ( ~n5554 & n5558 ) ;
  assign n5560 = ( n5047 & ~n5556 ) | ( n5047 & n5557 ) | ( ~n5556 & n5557 ) ;
  assign n5561 = ( ~n4958 & n5554 ) | ( ~n4958 & n5560 ) | ( n5554 & n5560 ) ;
  assign n5562 = ( n5553 & n5559 ) | ( n5553 & ~n5561 ) | ( n5559 & ~n5561 ) ;
  assign n5563 = x230 & ~n1003 ;
  assign n5564 = n925 | n2109 ;
  assign n5565 = ~n948 & n2103 ;
  assign n5566 = ( n1626 & n1880 ) | ( n1626 & ~n5565 ) | ( n1880 & ~n5565 ) ;
  assign n5567 = ~n942 & n5566 ;
  assign n5568 = ( n4008 & ~n5564 ) | ( n4008 & n5567 ) | ( ~n5564 & n5567 ) ;
  assign n5569 = n5563 & ~n5568 ;
  assign n5570 = ( ~n974 & n1883 ) | ( ~n974 & n2285 ) | ( n1883 & n2285 ) ;
  assign n5571 = ( ~n4008 & n5564 ) | ( ~n4008 & n5570 ) | ( n5564 & n5570 ) ;
  assign n5572 = n5563 & n5571 ;
  assign n5573 = ( n5562 & n5569 ) | ( n5562 & n5572 ) | ( n5569 & n5572 ) ;
  assign n5574 = x105 | n1410 ;
  assign n5575 = ~n1014 & n5574 ;
  assign n5576 = ( ~n996 & n1030 ) | ( ~n996 & n5575 ) | ( n1030 & n5575 ) ;
  assign n5577 = ( n1027 & ~n1028 ) | ( n1027 & n5576 ) | ( ~n1028 & n5576 ) ;
  assign n5578 = ( n1906 & ~n2299 ) | ( n1906 & n5577 ) | ( ~n2299 & n5577 ) ;
  assign n5579 = n1074 | n2132 ;
  assign n5580 = ( ~n1074 & n1078 ) | ( ~n1074 & n1913 ) | ( n1078 & n1913 ) ;
  assign n5581 = ( n5273 & n5579 ) | ( n5273 & ~n5580 ) | ( n5579 & ~n5580 ) ;
  assign n5582 = ( n1055 & ~n5579 ) | ( n1055 & n5580 ) | ( ~n5579 & n5580 ) ;
  assign n5583 = ( n5578 & ~n5581 ) | ( n5578 & n5582 ) | ( ~n5581 & n5582 ) ;
  assign n5584 = ~n1145 & n3567 ;
  assign n5585 = ( n2576 & ~n3574 ) | ( n2576 & n5584 ) | ( ~n3574 & n5584 ) ;
  assign n5586 = ( n3121 & n3574 ) | ( n3121 & ~n5584 ) | ( n3574 & ~n5584 ) ;
  assign n5587 = ( n5583 & ~n5585 ) | ( n5583 & n5586 ) | ( ~n5585 & n5586 ) ;
  assign n5588 = ( n1321 & n1714 ) | ( n1321 & ~n1949 ) | ( n1714 & ~n1949 ) ;
  assign n5589 = ~n1167 & n4030 ;
  assign n5590 = ( n1698 & ~n1700 ) | ( n1698 & n2150 ) | ( ~n1700 & n2150 ) ;
  assign n5591 = ( n1225 & n1269 ) | ( n1225 & ~n1698 ) | ( n1269 & ~n1698 ) ;
  assign n5592 = ( n5589 & n5590 ) | ( n5589 & ~n5591 ) | ( n5590 & ~n5591 ) ;
  assign n5593 = ( n4992 & ~n5588 ) | ( n4992 & n5592 ) | ( ~n5588 & n5592 ) ;
  assign n5594 = ( n5081 & ~n5590 ) | ( n5081 & n5591 ) | ( ~n5590 & n5591 ) ;
  assign n5595 = ( ~n4992 & n5588 ) | ( ~n4992 & n5594 ) | ( n5588 & n5594 ) ;
  assign n5596 = ( n5587 & n5593 ) | ( n5587 & ~n5595 ) | ( n5593 & ~n5595 ) ;
  assign n5597 = x231 & ~n1407 ;
  assign n5598 = n1329 | n2179 ;
  assign n5599 = ~n1352 & n2173 ;
  assign n5600 = ( n1724 & n1958 ) | ( n1724 & ~n5599 ) | ( n1958 & ~n5599 ) ;
  assign n5601 = ~n1346 & n5600 ;
  assign n5602 = ( n4046 & ~n5598 ) | ( n4046 & n5601 ) | ( ~n5598 & n5601 ) ;
  assign n5603 = n5597 & ~n5602 ;
  assign n5604 = ( ~n1378 & n1961 ) | ( ~n1378 & n2341 ) | ( n1961 & n2341 ) ;
  assign n5605 = ( ~n4046 & n5598 ) | ( ~n4046 & n5604 ) | ( n5598 & n5604 ) ;
  assign n5606 = n5597 & n5605 ;
  assign n5607 = ( n5596 & n5603 ) | ( n5596 & n5606 ) | ( n5603 & n5606 ) ;
  assign n5608 = x106 | n605 ;
  assign n5609 = ~n1418 & n5608 ;
  assign n5610 = ( ~n1400 & n1434 ) | ( ~n1400 & n5609 ) | ( n1434 & n5609 ) ;
  assign n5611 = ( n1431 & ~n1432 ) | ( n1431 & n5610 ) | ( ~n1432 & n5610 ) ;
  assign n5612 = ( n1984 & ~n2355 ) | ( n1984 & n5611 ) | ( ~n2355 & n5611 ) ;
  assign n5613 = n273 | n2201 ;
  assign n5614 = ( ~n273 & n277 ) | ( ~n273 & n1989 ) | ( n277 & n1989 ) ;
  assign n5615 = ( n5307 & n5613 ) | ( n5307 & ~n5614 ) | ( n5613 & ~n5614 ) ;
  assign n5616 = ( n1459 & ~n5613 ) | ( n1459 & n5614 ) | ( ~n5613 & n5614 ) ;
  assign n5617 = ( n5612 & ~n5615 ) | ( n5612 & n5616 ) | ( ~n5615 & n5616 ) ;
  assign n5618 = ~n330 & n3605 ;
  assign n5619 = ( n2611 & ~n3612 ) | ( n2611 & n5618 ) | ( ~n3612 & n5618 ) ;
  assign n5620 = ( n3157 & n3612 ) | ( n3157 & ~n5618 ) | ( n3612 & ~n5618 ) ;
  assign n5621 = ( n5617 & ~n5619 ) | ( n5617 & n5620 ) | ( ~n5619 & n5620 ) ;
  assign n5622 = ( n513 & n1799 ) | ( n513 & ~n2020 ) | ( n1799 & ~n2020 ) ;
  assign n5623 = n384 & ~n398 ;
  assign n5624 = ( n423 & n449 ) | ( n423 & ~n1786 ) | ( n449 & ~n1786 ) ;
  assign n5625 = ( n445 & ~n449 ) | ( n445 & n1504 ) | ( ~n449 & n1504 ) ;
  assign n5626 = ( n5623 & n5624 ) | ( n5623 & ~n5625 ) | ( n5624 & ~n5625 ) ;
  assign n5627 = ( n5026 & ~n5622 ) | ( n5026 & n5626 ) | ( ~n5622 & n5626 ) ;
  assign n5628 = ( n5115 & ~n5624 ) | ( n5115 & n5625 ) | ( ~n5624 & n5625 ) ;
  assign n5629 = ( ~n5026 & n5622 ) | ( ~n5026 & n5628 ) | ( n5622 & n5628 ) ;
  assign n5630 = ( n5621 & n5627 ) | ( n5621 & ~n5629 ) | ( n5627 & ~n5629 ) ;
  assign n5631 = x232 & ~n608 ;
  assign n5632 = n603 | n2234 ;
  assign n5633 = ~n534 & n2229 ;
  assign n5634 = ( n1808 & n2032 ) | ( n1808 & ~n5633 ) | ( n2032 & ~n5633 ) ;
  assign n5635 = ~n531 & n5634 ;
  assign n5636 = ( n4083 & ~n5632 ) | ( n4083 & n5635 ) | ( ~n5632 & n5635 ) ;
  assign n5637 = n5631 & ~n5636 ;
  assign n5638 = ( n539 & ~n1538 ) | ( n539 & n2035 ) | ( ~n1538 & n2035 ) ;
  assign n5639 = ( ~n4083 & n5632 ) | ( ~n4083 & n5638 ) | ( n5632 & n5638 ) ;
  assign n5640 = n5631 & n5639 ;
  assign n5641 = ( n5630 & n5637 ) | ( n5630 & n5640 ) | ( n5637 & n5640 ) ;
  assign n5642 = x107 | n1010 ;
  assign n5643 = ~n590 & n5642 ;
  assign n5644 = ( ~n588 & n597 ) | ( ~n588 & n5643 ) | ( n597 & n5643 ) ;
  assign n5645 = ( ~n628 & n1552 ) | ( ~n628 & n5644 ) | ( n1552 & n5644 ) ;
  assign n5646 = ( n2054 & ~n2399 ) | ( n2054 & n5645 ) | ( ~n2399 & n5645 ) ;
  assign n5647 = n678 | n2257 ;
  assign n5648 = ( ~n678 & n682 ) | ( ~n678 & n2059 ) | ( n682 & n2059 ) ;
  assign n5649 = ( n5341 & n5647 ) | ( n5341 & ~n5648 ) | ( n5647 & ~n5648 ) ;
  assign n5650 = ( n1563 & ~n5647 ) | ( n1563 & n5648 ) | ( ~n5647 & n5648 ) ;
  assign n5651 = ( n5646 & ~n5649 ) | ( n5646 & n5650 ) | ( ~n5649 & n5650 ) ;
  assign n5652 = ~n735 & n3643 ;
  assign n5653 = ( n2646 & ~n3650 ) | ( n2646 & n5652 ) | ( ~n3650 & n5652 ) ;
  assign n5654 = ( n3193 & n3650 ) | ( n3193 & ~n5652 ) | ( n3650 & ~n5652 ) ;
  assign n5655 = ( n5651 & ~n5653 ) | ( n5651 & n5654 ) | ( ~n5653 & n5654 ) ;
  assign n5656 = ( n918 & n1877 ) | ( n918 & ~n2090 ) | ( n1877 & ~n2090 ) ;
  assign n5657 = n789 & ~n803 ;
  assign n5658 = ( n828 & n854 ) | ( n828 & ~n1864 ) | ( n854 & ~n1864 ) ;
  assign n5659 = ( n850 & ~n854 ) | ( n850 & n1603 ) | ( ~n854 & n1603 ) ;
  assign n5660 = ( n5657 & n5658 ) | ( n5657 & ~n5659 ) | ( n5658 & ~n5659 ) ;
  assign n5661 = ( n5060 & ~n5656 ) | ( n5060 & n5660 ) | ( ~n5656 & n5660 ) ;
  assign n5662 = ( n5149 & ~n5658 ) | ( n5149 & n5659 ) | ( ~n5658 & n5659 ) ;
  assign n5663 = ( ~n5060 & n5656 ) | ( ~n5060 & n5662 ) | ( n5656 & n5662 ) ;
  assign n5664 = ( n5655 & n5661 ) | ( n5655 & ~n5663 ) | ( n5661 & ~n5663 ) ;
  assign n5665 = x233 & ~n1013 ;
  assign n5666 = n1008 | n2290 ;
  assign n5667 = ~n939 & n2285 ;
  assign n5668 = ( n1886 & n2102 ) | ( n1886 & ~n5667 ) | ( n2102 & ~n5667 ) ;
  assign n5669 = ~n936 & n5668 ;
  assign n5670 = ( n4120 & ~n5666 ) | ( n4120 & n5669 ) | ( ~n5666 & n5669 ) ;
  assign n5671 = n5665 & ~n5670 ;
  assign n5672 = ( n944 & ~n1637 ) | ( n944 & n2105 ) | ( ~n1637 & n2105 ) ;
  assign n5673 = ( ~n4120 & n5666 ) | ( ~n4120 & n5672 ) | ( n5666 & n5672 ) ;
  assign n5674 = n5665 & n5673 ;
  assign n5675 = ( n5664 & n5671 ) | ( n5664 & n5674 ) | ( n5671 & n5674 ) ;
  assign n5676 = x108 | n1414 ;
  assign n5677 = ~n995 & n5676 ;
  assign n5678 = ( ~n993 & n1002 ) | ( ~n993 & n5677 ) | ( n1002 & n5677 ) ;
  assign n5679 = ( ~n1033 & n1651 ) | ( ~n1033 & n5678 ) | ( n1651 & n5678 ) ;
  assign n5680 = ( n2124 & ~n2443 ) | ( n2124 & n5679 ) | ( ~n2443 & n5679 ) ;
  assign n5681 = n1082 | n2313 ;
  assign n5682 = ( ~n1082 & n1086 ) | ( ~n1082 & n2129 ) | ( n1086 & n2129 ) ;
  assign n5683 = ( n5375 & n5681 ) | ( n5375 & ~n5682 ) | ( n5681 & ~n5682 ) ;
  assign n5684 = ( n1662 & ~n5681 ) | ( n1662 & n5682 ) | ( ~n5681 & n5682 ) ;
  assign n5685 = ( n5680 & ~n5683 ) | ( n5680 & n5684 ) | ( ~n5683 & n5684 ) ;
  assign n5686 = ~n1139 & n3681 ;
  assign n5687 = ( n2681 & ~n3688 ) | ( n2681 & n5686 ) | ( ~n3688 & n5686 ) ;
  assign n5688 = ( n3229 & n3688 ) | ( n3229 & ~n5686 ) | ( n3688 & ~n5686 ) ;
  assign n5689 = ( n5685 & ~n5687 ) | ( n5685 & n5688 ) | ( ~n5687 & n5688 ) ;
  assign n5690 = ( n1322 & n1955 ) | ( n1322 & ~n2160 ) | ( n1955 & ~n2160 ) ;
  assign n5691 = n1193 & ~n1207 ;
  assign n5692 = ( n1232 & n1258 ) | ( n1232 & ~n1942 ) | ( n1258 & ~n1942 ) ;
  assign n5693 = ( n1254 & ~n1258 ) | ( n1254 & n1701 ) | ( ~n1258 & n1701 ) ;
  assign n5694 = ( n5691 & n5692 ) | ( n5691 & ~n5693 ) | ( n5692 & ~n5693 ) ;
  assign n5695 = ( n5094 & ~n5690 ) | ( n5094 & n5694 ) | ( ~n5690 & n5694 ) ;
  assign n5696 = ( n5183 & ~n5692 ) | ( n5183 & n5693 ) | ( ~n5692 & n5693 ) ;
  assign n5697 = ( ~n5094 & n5690 ) | ( ~n5094 & n5696 ) | ( n5690 & n5696 ) ;
  assign n5698 = ( n5689 & n5695 ) | ( n5689 & ~n5697 ) | ( n5695 & ~n5697 ) ;
  assign n5699 = x234 & ~n1417 ;
  assign n5700 = n1412 | n2346 ;
  assign n5701 = ~n1343 & n2341 ;
  assign n5702 = ( n1964 & n2172 ) | ( n1964 & ~n5701 ) | ( n2172 & ~n5701 ) ;
  assign n5703 = ~n1340 & n5702 ;
  assign n5704 = ( n4157 & ~n5700 ) | ( n4157 & n5703 ) | ( ~n5700 & n5703 ) ;
  assign n5705 = n5699 & ~n5704 ;
  assign n5706 = ( n1348 & ~n1735 ) | ( n1348 & n2175 ) | ( ~n1735 & n2175 ) ;
  assign n5707 = ( ~n4157 & n5700 ) | ( ~n4157 & n5706 ) | ( n5700 & n5706 ) ;
  assign n5708 = n5699 & n5707 ;
  assign n5709 = ( n5698 & n5705 ) | ( n5698 & n5708 ) | ( n5705 & n5708 ) ;
  assign n5710 = x109 | n592 ;
  assign n5711 = ~n1399 & n5710 ;
  assign n5712 = ( ~n1397 & n1406 ) | ( ~n1397 & n5711 ) | ( n1406 & n5711 ) ;
  assign n5713 = ( ~n1437 & n1749 ) | ( ~n1437 & n5712 ) | ( n1749 & n5712 ) ;
  assign n5714 = ( n2194 & ~n2487 ) | ( n2194 & n5713 ) | ( ~n2487 & n5713 ) ;
  assign n5715 = n297 | n2369 ;
  assign n5716 = ( ~n297 & n1476 ) | ( ~n297 & n2199 ) | ( n1476 & n2199 ) ;
  assign n5717 = ( n5409 & n5715 ) | ( n5409 & ~n5716 ) | ( n5715 & ~n5716 ) ;
  assign n5718 = ( n1757 & ~n5715 ) | ( n1757 & n5716 ) | ( ~n5715 & n5716 ) ;
  assign n5719 = ( n5714 & ~n5717 ) | ( n5714 & n5718 ) | ( ~n5717 & n5718 ) ;
  assign n5720 = ~n380 & n3719 ;
  assign n5721 = ( n2716 & ~n3726 ) | ( n2716 & n5720 ) | ( ~n3726 & n5720 ) ;
  assign n5722 = ( n3265 & n3726 ) | ( n3265 & ~n5720 ) | ( n3726 & ~n5720 ) ;
  assign n5723 = ( n5719 & ~n5721 ) | ( n5719 & n5722 ) | ( ~n5721 & n5722 ) ;
  assign n5724 = ( ~n486 & n487 ) | ( ~n486 & n2026 ) | ( n487 & n2026 ) ;
  assign n5725 = ~n408 & n1499 ;
  assign n5726 = ( n453 & n1508 ) | ( n453 & ~n2013 ) | ( n1508 & ~n2013 ) ;
  assign n5727 = ( n442 & ~n453 ) | ( n442 & n1787 ) | ( ~n453 & n1787 ) ;
  assign n5728 = ( n5725 & n5726 ) | ( n5725 & ~n5727 ) | ( n5726 & ~n5727 ) ;
  assign n5729 = ( n5128 & ~n5724 ) | ( n5128 & n5728 ) | ( ~n5724 & n5728 ) ;
  assign n5730 = ( n5217 & ~n5726 ) | ( n5217 & n5727 ) | ( ~n5726 & n5727 ) ;
  assign n5731 = ( ~n5128 & n5724 ) | ( ~n5128 & n5730 ) | ( n5724 & n5730 ) ;
  assign n5732 = ( n5723 & n5729 ) | ( n5723 & ~n5731 ) | ( n5729 & ~n5731 ) ;
  assign n5733 = x235 & ~n589 ;
  assign n5734 = n607 | n2393 ;
  assign n5735 = n539 & ~n559 ;
  assign n5736 = ( n565 & n2030 ) | ( n565 & ~n5735 ) | ( n2030 & ~n5735 ) ;
  assign n5737 = ~n526 & n5736 ;
  assign n5738 = ( n4194 & ~n5734 ) | ( n4194 & n5737 ) | ( ~n5734 & n5737 ) ;
  assign n5739 = n5733 & ~n5738 ;
  assign n5740 = ( n1532 & ~n1817 ) | ( n1532 & n2231 ) | ( ~n1817 & n2231 ) ;
  assign n5741 = ( ~n4194 & n5734 ) | ( ~n4194 & n5740 ) | ( n5734 & n5740 ) ;
  assign n5742 = n5733 & n5741 ;
  assign n5743 = ( n5732 & n5739 ) | ( n5732 & n5742 ) | ( n5739 & n5742 ) ;
  assign n5744 = x110 | n997 ;
  assign n5745 = ~n587 & n5744 ;
  assign n5746 = ( ~n581 & n585 ) | ( ~n581 & n5745 ) | ( n585 & n5745 ) ;
  assign n5747 = ( ~n1549 & n1828 ) | ( ~n1549 & n5746 ) | ( n1828 & n5746 ) ;
  assign n5748 = ( ~n658 & n1827 ) | ( ~n658 & n5747 ) | ( n1827 & n5747 ) ;
  assign n5749 = n702 | n2413 ;
  assign n5750 = ( ~n702 & n1575 ) | ( ~n702 & n2255 ) | ( n1575 & n2255 ) ;
  assign n5751 = ( n5443 & n5749 ) | ( n5443 & ~n5750 ) | ( n5749 & ~n5750 ) ;
  assign n5752 = ( n1835 & ~n5749 ) | ( n1835 & n5750 ) | ( ~n5749 & n5750 ) ;
  assign n5753 = ( n5748 & ~n5751 ) | ( n5748 & n5752 ) | ( ~n5751 & n5752 ) ;
  assign n5754 = ~n785 & n3757 ;
  assign n5755 = ( n3304 & n3764 ) | ( n3304 & ~n5754 ) | ( n3764 & ~n5754 ) ;
  assign n5756 = ( n2750 & ~n3764 ) | ( n2750 & n5754 ) | ( ~n3764 & n5754 ) ;
  assign n5757 = ( n5753 & n5755 ) | ( n5753 & ~n5756 ) | ( n5755 & ~n5756 ) ;
  assign n5758 = ( ~n891 & n892 ) | ( ~n891 & n2096 ) | ( n892 & n2096 ) ;
  assign n5759 = ~n813 & n1598 ;
  assign n5760 = ( n858 & n1607 ) | ( n858 & ~n2083 ) | ( n1607 & ~n2083 ) ;
  assign n5761 = ( n847 & ~n858 ) | ( n847 & n1865 ) | ( ~n858 & n1865 ) ;
  assign n5762 = ( n5759 & n5760 ) | ( n5759 & ~n5761 ) | ( n5760 & ~n5761 ) ;
  assign n5763 = ( n5162 & ~n5758 ) | ( n5162 & n5762 ) | ( ~n5758 & n5762 ) ;
  assign n5764 = ( n5251 & ~n5760 ) | ( n5251 & n5761 ) | ( ~n5760 & n5761 ) ;
  assign n5765 = ( ~n5162 & n5758 ) | ( ~n5162 & n5764 ) | ( n5758 & n5764 ) ;
  assign n5766 = ( n5757 & n5763 ) | ( n5757 & ~n5765 ) | ( n5763 & ~n5765 ) ;
  assign n5767 = x236 & ~n994 ;
  assign n5768 = n1012 | n2437 ;
  assign n5769 = n944 & ~n964 ;
  assign n5770 = ( n970 & n2100 ) | ( n970 & ~n5769 ) | ( n2100 & ~n5769 ) ;
  assign n5771 = ~n931 & n5770 ;
  assign n5772 = ( n4231 & ~n5768 ) | ( n4231 & n5771 ) | ( ~n5768 & n5771 ) ;
  assign n5773 = n5767 & ~n5772 ;
  assign n5774 = ( n1631 & ~n1895 ) | ( n1631 & n2287 ) | ( ~n1895 & n2287 ) ;
  assign n5775 = ( ~n4231 & n5768 ) | ( ~n4231 & n5774 ) | ( n5768 & n5774 ) ;
  assign n5776 = n5767 & n5775 ;
  assign n5777 = ( n5766 & n5773 ) | ( n5766 & n5776 ) | ( n5773 & n5776 ) ;
  assign n5778 = x111 | n1401 ;
  assign n5779 = ~n992 & n5778 ;
  assign n5780 = ( ~n986 & n990 ) | ( ~n986 & n5779 ) | ( n990 & n5779 ) ;
  assign n5781 = ( ~n1648 & n1906 ) | ( ~n1648 & n5780 ) | ( n1906 & n5780 ) ;
  assign n5782 = ( ~n1063 & n1905 ) | ( ~n1063 & n5781 ) | ( n1905 & n5781 ) ;
  assign n5783 = n1106 | n2457 ;
  assign n5784 = ( ~n1106 & n1673 ) | ( ~n1106 & n2311 ) | ( n1673 & n2311 ) ;
  assign n5785 = ( n5477 & n5783 ) | ( n5477 & ~n5784 ) | ( n5783 & ~n5784 ) ;
  assign n5786 = ( n1913 & ~n5783 ) | ( n1913 & n5784 ) | ( ~n5783 & n5784 ) ;
  assign n5787 = ( n5782 & ~n5785 ) | ( n5782 & n5786 ) | ( ~n5785 & n5786 ) ;
  assign n5788 = ~n1189 & n3795 ;
  assign n5789 = ( n3343 & n3802 ) | ( n3343 & ~n5788 ) | ( n3802 & ~n5788 ) ;
  assign n5790 = ( n2789 & ~n3802 ) | ( n2789 & n5788 ) | ( ~n3802 & n5788 ) ;
  assign n5791 = ( n5787 & n5789 ) | ( n5787 & ~n5790 ) | ( n5789 & ~n5790 ) ;
  assign n5792 = ( ~n1295 & n1296 ) | ( ~n1295 & n2166 ) | ( n1296 & n2166 ) ;
  assign n5793 = ~n1217 & n1696 ;
  assign n5794 = ( n1262 & n1705 ) | ( n1262 & ~n2153 ) | ( n1705 & ~n2153 ) ;
  assign n5795 = ( n1251 & ~n1262 ) | ( n1251 & n1943 ) | ( ~n1262 & n1943 ) ;
  assign n5796 = ( n5793 & n5794 ) | ( n5793 & ~n5795 ) | ( n5794 & ~n5795 ) ;
  assign n5797 = ( n5196 & ~n5792 ) | ( n5196 & n5796 ) | ( ~n5792 & n5796 ) ;
  assign n5798 = ( n5285 & ~n5794 ) | ( n5285 & n5795 ) | ( ~n5794 & n5795 ) ;
  assign n5799 = ( ~n5196 & n5792 ) | ( ~n5196 & n5798 ) | ( n5792 & n5798 ) ;
  assign n5800 = ( n5791 & n5797 ) | ( n5791 & ~n5799 ) | ( n5797 & ~n5799 ) ;
  assign n5801 = x237 & ~n1398 ;
  assign n5802 = n1416 | n2481 ;
  assign n5803 = n1348 & ~n1368 ;
  assign n5804 = ( n1374 & n2170 ) | ( n1374 & ~n5803 ) | ( n2170 & ~n5803 ) ;
  assign n5805 = ~n1335 & n5804 ;
  assign n5806 = ( n4268 & ~n5802 ) | ( n4268 & n5805 ) | ( ~n5802 & n5805 ) ;
  assign n5807 = n5801 & ~n5806 ;
  assign n5808 = ( n1729 & ~n1973 ) | ( n1729 & n2343 ) | ( ~n1973 & n2343 ) ;
  assign n5809 = ( ~n4268 & n5802 ) | ( ~n4268 & n5808 ) | ( n5802 & n5808 ) ;
  assign n5810 = n5801 & n5809 ;
  assign n5811 = ( n5800 & n5807 ) | ( n5800 & n5810 ) | ( n5807 & n5810 ) ;
  assign n5812 = x112 | n582 ;
  assign n5813 = ~n1396 & n5812 ;
  assign n5814 = ( ~n1390 & n1394 ) | ( ~n1390 & n5813 ) | ( n1394 & n5813 ) ;
  assign n5815 = ( ~n1746 & n1984 ) | ( ~n1746 & n5814 ) | ( n1984 & n5814 ) ;
  assign n5816 = ( ~n1467 & n1983 ) | ( ~n1467 & n5815 ) | ( n1983 & n5815 ) ;
  assign n5817 = n289 | n2501 ;
  assign n5818 = ( ~n289 & n293 ) | ( ~n289 & n2367 ) | ( n293 & n2367 ) ;
  assign n5819 = ( n5511 & n5817 ) | ( n5511 & ~n5818 ) | ( n5817 & ~n5818 ) ;
  assign n5820 = ( n1989 & ~n5817 ) | ( n1989 & n5818 ) | ( ~n5817 & n5818 ) ;
  assign n5821 = ( n5816 & ~n5819 ) | ( n5816 & n5820 ) | ( ~n5819 & n5820 ) ;
  assign n5822 = ~n368 & n3833 ;
  assign n5823 = ( n3382 & n3840 ) | ( n3382 & ~n5822 ) | ( n3840 & ~n5822 ) ;
  assign n5824 = ( n2827 & ~n3840 ) | ( n2827 & n5822 ) | ( ~n3840 & n5822 ) ;
  assign n5825 = ( n5821 & n5823 ) | ( n5821 & ~n5824 ) | ( n5823 & ~n5824 ) ;
  assign n5826 = ( n507 & ~n1520 ) | ( n507 & n2223 ) | ( ~n1520 & n2223 ) ;
  assign n5827 = ~n413 & n1783 ;
  assign n5828 = ( n437 & ~n465 ) | ( n437 & n1791 ) | ( ~n465 & n1791 ) ;
  assign n5829 = ( n433 & ~n437 ) | ( n433 & n2014 ) | ( ~n437 & n2014 ) ;
  assign n5830 = ( n5827 & n5828 ) | ( n5827 & ~n5829 ) | ( n5828 & ~n5829 ) ;
  assign n5831 = ( n5230 & ~n5826 ) | ( n5230 & n5830 ) | ( ~n5826 & n5830 ) ;
  assign n5832 = ( n5319 & ~n5828 ) | ( n5319 & n5829 ) | ( ~n5828 & n5829 ) ;
  assign n5833 = ( ~n5230 & n5826 ) | ( ~n5230 & n5832 ) | ( n5826 & n5832 ) ;
  assign n5834 = ( n5825 & n5831 ) | ( n5825 & ~n5833 ) | ( n5831 & ~n5833 ) ;
  assign n5835 = x238 & ~n586 ;
  assign n5836 = n594 | n626 ;
  assign n5837 = ~n523 & n1532 ;
  assign n5838 = ( n561 & n2227 ) | ( n561 & ~n5837 ) | ( n2227 & ~n5837 ) ;
  assign n5839 = ~n520 & n5838 ;
  assign n5840 = ( n4305 & ~n5836 ) | ( n4305 & n5839 ) | ( ~n5836 & n5839 ) ;
  assign n5841 = n5835 & ~n5840 ;
  assign n5842 = ( n563 & ~n4305 ) | ( n563 & n5836 ) | ( ~n4305 & n5836 ) ;
  assign n5843 = n5835 & n5842 ;
  assign n5844 = ( n5834 & n5841 ) | ( n5834 & n5843 ) | ( n5841 & n5843 ) ;
  assign n5845 = x113 | n987 ;
  assign n5846 = ~n580 & n5845 ;
  assign n5847 = ( ~n575 & n621 ) | ( ~n575 & n5846 ) | ( n621 & n5846 ) ;
  assign n5848 = ( ~n656 & n2054 ) | ( ~n656 & n5847 ) | ( n2054 & n5847 ) ;
  assign n5849 = ( ~n1566 & n2053 ) | ( ~n1566 & n5848 ) | ( n2053 & n5848 ) ;
  assign n5850 = n694 | n2538 ;
  assign n5851 = ( ~n694 & n698 ) | ( ~n694 & n2411 ) | ( n698 & n2411 ) ;
  assign n5852 = ( n5545 & n5850 ) | ( n5545 & ~n5851 ) | ( n5850 & ~n5851 ) ;
  assign n5853 = ( n2059 & ~n5850 ) | ( n2059 & n5851 ) | ( ~n5850 & n5851 ) ;
  assign n5854 = ( n5849 & ~n5852 ) | ( n5849 & n5853 ) | ( ~n5852 & n5853 ) ;
  assign n5855 = ~n773 & n3871 ;
  assign n5856 = ( n3421 & n3878 ) | ( n3421 & ~n5855 ) | ( n3878 & ~n5855 ) ;
  assign n5857 = ( n2864 & ~n3878 ) | ( n2864 & n5855 ) | ( ~n3878 & n5855 ) ;
  assign n5858 = ( n5854 & n5856 ) | ( n5854 & ~n5857 ) | ( n5856 & ~n5857 ) ;
  assign n5859 = ( n912 & ~n1619 ) | ( n912 & n2279 ) | ( ~n1619 & n2279 ) ;
  assign n5860 = ~n818 & n1861 ;
  assign n5861 = ( n842 & ~n870 ) | ( n842 & n1869 ) | ( ~n870 & n1869 ) ;
  assign n5862 = ( n838 & ~n842 ) | ( n838 & n2084 ) | ( ~n842 & n2084 ) ;
  assign n5863 = ( n5860 & n5861 ) | ( n5860 & ~n5862 ) | ( n5861 & ~n5862 ) ;
  assign n5864 = ( n5264 & ~n5859 ) | ( n5264 & n5863 ) | ( ~n5859 & n5863 ) ;
  assign n5865 = ( n5353 & ~n5861 ) | ( n5353 & n5862 ) | ( ~n5861 & n5862 ) ;
  assign n5866 = ( ~n5264 & n5859 ) | ( ~n5264 & n5865 ) | ( n5859 & n5865 ) ;
  assign n5867 = ( n5858 & n5864 ) | ( n5858 & ~n5866 ) | ( n5864 & ~n5866 ) ;
  assign n5868 = x239 & ~n991 ;
  assign n5869 = n999 | n1031 ;
  assign n5870 = ~n928 & n1631 ;
  assign n5871 = ( n966 & n2283 ) | ( n966 & ~n5870 ) | ( n2283 & ~n5870 ) ;
  assign n5872 = ~n925 & n5871 ;
  assign n5873 = ( n4341 & ~n5869 ) | ( n4341 & n5872 ) | ( ~n5869 & n5872 ) ;
  assign n5874 = n5868 & ~n5873 ;
  assign n5875 = ( n968 & ~n4341 ) | ( n968 & n5869 ) | ( ~n4341 & n5869 ) ;
  assign n5876 = n5868 & n5875 ;
  assign n5877 = ( n5867 & n5874 ) | ( n5867 & n5876 ) | ( n5874 & n5876 ) ;
  assign n5878 = x114 | n1391 ;
  assign n5879 = ~n985 & n5878 ;
  assign n5880 = ( ~n980 & n1026 ) | ( ~n980 & n5879 ) | ( n1026 & n5879 ) ;
  assign n5881 = ( ~n1061 & n2124 ) | ( ~n1061 & n5880 ) | ( n2124 & n5880 ) ;
  assign n5882 = ( ~n1665 & n2123 ) | ( ~n1665 & n5881 ) | ( n2123 & n5881 ) ;
  assign n5883 = n1098 | n2575 ;
  assign n5884 = ( ~n1098 & n1102 ) | ( ~n1098 & n2455 ) | ( n1102 & n2455 ) ;
  assign n5885 = ( n5579 & n5883 ) | ( n5579 & ~n5884 ) | ( n5883 & ~n5884 ) ;
  assign n5886 = ( n2129 & ~n5883 ) | ( n2129 & n5884 ) | ( ~n5883 & n5884 ) ;
  assign n5887 = ( n5882 & ~n5885 ) | ( n5882 & n5886 ) | ( ~n5885 & n5886 ) ;
  assign n5888 = ~n1177 & n3909 ;
  assign n5889 = ( n3460 & n3916 ) | ( n3460 & ~n5888 ) | ( n3916 & ~n5888 ) ;
  assign n5890 = ( n2901 & ~n3916 ) | ( n2901 & n5888 ) | ( ~n3916 & n5888 ) ;
  assign n5891 = ( n5887 & n5889 ) | ( n5887 & ~n5890 ) | ( n5889 & ~n5890 ) ;
  assign n5892 = ( n1316 & ~n1717 ) | ( n1316 & n2335 ) | ( ~n1717 & n2335 ) ;
  assign n5893 = ~n1222 & n1939 ;
  assign n5894 = ( n1246 & ~n1274 ) | ( n1246 & n1947 ) | ( ~n1274 & n1947 ) ;
  assign n5895 = ( n1242 & ~n1246 ) | ( n1242 & n2154 ) | ( ~n1246 & n2154 ) ;
  assign n5896 = ( n5893 & n5894 ) | ( n5893 & ~n5895 ) | ( n5894 & ~n5895 ) ;
  assign n5897 = ( n5298 & ~n5892 ) | ( n5298 & n5896 ) | ( ~n5892 & n5896 ) ;
  assign n5898 = ( n5387 & ~n5894 ) | ( n5387 & n5895 ) | ( ~n5894 & n5895 ) ;
  assign n5899 = ( ~n5298 & n5892 ) | ( ~n5298 & n5898 ) | ( n5892 & n5898 ) ;
  assign n5900 = ( n5891 & n5897 ) | ( n5891 & ~n5899 ) | ( n5897 & ~n5899 ) ;
  assign n5901 = x240 & ~n1395 ;
  assign n5902 = n1403 | n1435 ;
  assign n5903 = ~n1332 & n1729 ;
  assign n5904 = ( n1370 & n2339 ) | ( n1370 & ~n5903 ) | ( n2339 & ~n5903 ) ;
  assign n5905 = ~n1329 & n5904 ;
  assign n5906 = ( n4377 & ~n5902 ) | ( n4377 & n5905 ) | ( ~n5902 & n5905 ) ;
  assign n5907 = n5901 & ~n5906 ;
  assign n5908 = ( n1372 & ~n4377 ) | ( n1372 & n5902 ) | ( ~n4377 & n5902 ) ;
  assign n5909 = n5901 & n5908 ;
  assign n5910 = ( n5900 & n5907 ) | ( n5900 & n5909 ) | ( n5907 & n5909 ) ;
  assign n5911 = x115 | n576 ;
  assign n5912 = ~n1389 & n5911 ;
  assign n5913 = ( ~n1384 & n1430 ) | ( ~n1384 & n5912 ) | ( n1430 & n5912 ) ;
  assign n5914 = ( ~n1465 & n2194 ) | ( ~n1465 & n5913 ) | ( n2194 & n5913 ) ;
  assign n5915 = ( ~n1760 & n2193 ) | ( ~n1760 & n5914 ) | ( n2193 & n5914 ) ;
  assign n5916 = n300 | n307 ;
  assign n5917 = ( ~n307 & n1479 ) | ( ~n307 & n2499 ) | ( n1479 & n2499 ) ;
  assign n5918 = ( n5613 & n5916 ) | ( n5613 & ~n5917 ) | ( n5916 & ~n5917 ) ;
  assign n5919 = ( n2199 & ~n5916 ) | ( n2199 & n5917 ) | ( ~n5916 & n5917 ) ;
  assign n5920 = ( n5915 & ~n5918 ) | ( n5915 & n5919 ) | ( ~n5918 & n5919 ) ;
  assign n5921 = ~n362 & n3947 ;
  assign n5922 = ( n3498 & n3954 ) | ( n3498 & ~n5921 ) | ( n3954 & ~n5921 ) ;
  assign n5923 = ( n2938 & ~n3954 ) | ( n2938 & n5921 ) | ( ~n3954 & n5921 ) ;
  assign n5924 = ( n5920 & n5922 ) | ( n5920 & ~n5923 ) | ( n5922 & ~n5923 ) ;
  assign n5925 = ( n515 & n1523 ) | ( n515 & ~n1803 ) | ( n1523 & ~n1803 ) ;
  assign n5926 = ~n391 & n2010 ;
  assign n5927 = ( n457 & ~n1516 ) | ( n457 & n2018 ) | ( ~n1516 & n2018 ) ;
  assign n5928 = ( ~n467 & n5926 ) | ( ~n467 & n5927 ) | ( n5926 & n5927 ) ;
  assign n5929 = ( n5332 & ~n5925 ) | ( n5332 & n5928 ) | ( ~n5925 & n5928 ) ;
  assign n5930 = ( n467 & n5421 ) | ( n467 & ~n5927 ) | ( n5421 & ~n5927 ) ;
  assign n5931 = ( ~n5332 & n5925 ) | ( ~n5332 & n5930 ) | ( n5925 & n5930 ) ;
  assign n5932 = ( n5924 & n5929 ) | ( n5924 & ~n5931 ) | ( n5929 & ~n5931 ) ;
  assign n5933 = x241 & ~n579 ;
  assign n5934 = n584 | n1553 ;
  assign n5935 = n528 & ~n600 ;
  assign n5936 = ( n570 & n1535 ) | ( n570 & ~n5935 ) | ( n1535 & ~n5935 ) ;
  assign n5937 = ~n603 & n5936 ;
  assign n5938 = ( n4412 & ~n5934 ) | ( n4412 & n5937 ) | ( ~n5934 & n5937 ) ;
  assign n5939 = n5933 & ~n5938 ;
  assign n5940 = ( n1537 & ~n4412 ) | ( n1537 & n5934 ) | ( ~n4412 & n5934 ) ;
  assign n5941 = n5933 & n5940 ;
  assign n5942 = ( n5932 & n5939 ) | ( n5932 & n5941 ) | ( n5939 & n5941 ) ;
  assign n5943 = x116 | n981 ;
  assign n5944 = ~n574 & n5943 ;
  assign n5945 = ( ~n655 & n1551 ) | ( ~n655 & n5944 ) | ( n1551 & n5944 ) ;
  assign n5946 = ( ~n657 & n1827 ) | ( ~n657 & n5945 ) | ( n1827 & n5945 ) ;
  assign n5947 = ( ~n1838 & n2248 ) | ( ~n1838 & n5946 ) | ( n2248 & n5946 ) ;
  assign n5948 = n705 | n712 ;
  assign n5949 = ( ~n712 & n1578 ) | ( ~n712 & n2536 ) | ( n1578 & n2536 ) ;
  assign n5950 = ( n5647 & n5948 ) | ( n5647 & ~n5949 ) | ( n5948 & ~n5949 ) ;
  assign n5951 = ( n2255 & ~n5948 ) | ( n2255 & n5949 ) | ( ~n5948 & n5949 ) ;
  assign n5952 = ( n5947 & ~n5950 ) | ( n5947 & n5951 ) | ( ~n5950 & n5951 ) ;
  assign n5953 = ~n767 & n3985 ;
  assign n5954 = ( n3536 & n3992 ) | ( n3536 & ~n5953 ) | ( n3992 & ~n5953 ) ;
  assign n5955 = ( n2974 & ~n3992 ) | ( n2974 & n5953 ) | ( ~n3992 & n5953 ) ;
  assign n5956 = ( n5952 & n5954 ) | ( n5952 & ~n5955 ) | ( n5954 & ~n5955 ) ;
  assign n5957 = ( n920 & n1622 ) | ( n920 & ~n1881 ) | ( n1622 & ~n1881 ) ;
  assign n5958 = ~n796 & n2080 ;
  assign n5959 = ( n862 & ~n1615 ) | ( n862 & n2088 ) | ( ~n1615 & n2088 ) ;
  assign n5960 = ( ~n872 & n5958 ) | ( ~n872 & n5959 ) | ( n5958 & n5959 ) ;
  assign n5961 = ( n5366 & ~n5957 ) | ( n5366 & n5960 ) | ( ~n5957 & n5960 ) ;
  assign n5962 = ( n872 & n5455 ) | ( n872 & ~n5959 ) | ( n5455 & ~n5959 ) ;
  assign n5963 = ( ~n5366 & n5957 ) | ( ~n5366 & n5962 ) | ( n5957 & n5962 ) ;
  assign n5964 = ( n5956 & n5961 ) | ( n5956 & ~n5963 ) | ( n5961 & ~n5963 ) ;
  assign n5965 = x242 & ~n984 ;
  assign n5966 = n989 | n1652 ;
  assign n5967 = n933 & ~n1005 ;
  assign n5968 = ( n975 & n1634 ) | ( n975 & ~n5967 ) | ( n1634 & ~n5967 ) ;
  assign n5969 = ~n1008 & n5968 ;
  assign n5970 = ( n4448 & ~n5966 ) | ( n4448 & n5969 ) | ( ~n5966 & n5969 ) ;
  assign n5971 = n5965 & ~n5970 ;
  assign n5972 = ( n1636 & ~n4448 ) | ( n1636 & n5966 ) | ( ~n4448 & n5966 ) ;
  assign n5973 = n5965 & n5972 ;
  assign n5974 = ( n5964 & n5971 ) | ( n5964 & n5973 ) | ( n5971 & n5973 ) ;
  assign n5975 = x117 | n1385 ;
  assign n5976 = ~n979 & n5975 ;
  assign n5977 = ( ~n1060 & n1650 ) | ( ~n1060 & n5976 ) | ( n1650 & n5976 ) ;
  assign n5978 = ( ~n1062 & n1905 ) | ( ~n1062 & n5977 ) | ( n1905 & n5977 ) ;
  assign n5979 = ( ~n1916 & n2304 ) | ( ~n1916 & n5978 ) | ( n2304 & n5978 ) ;
  assign n5980 = n1109 | n1116 ;
  assign n5981 = ( ~n1116 & n1676 ) | ( ~n1116 & n2573 ) | ( n1676 & n2573 ) ;
  assign n5982 = ( n5681 & n5980 ) | ( n5681 & ~n5981 ) | ( n5980 & ~n5981 ) ;
  assign n5983 = ( n2311 & ~n5980 ) | ( n2311 & n5981 ) | ( ~n5980 & n5981 ) ;
  assign n5984 = ( n5979 & ~n5982 ) | ( n5979 & n5983 ) | ( ~n5982 & n5983 ) ;
  assign n5985 = ~n1171 & n4023 ;
  assign n5986 = ( n3574 & n4030 ) | ( n3574 & ~n5985 ) | ( n4030 & ~n5985 ) ;
  assign n5987 = ( n3010 & ~n4030 ) | ( n3010 & n5985 ) | ( ~n4030 & n5985 ) ;
  assign n5988 = ( n5984 & n5986 ) | ( n5984 & ~n5987 ) | ( n5986 & ~n5987 ) ;
  assign n5989 = ( n1324 & n1720 ) | ( n1324 & ~n1959 ) | ( n1720 & ~n1959 ) ;
  assign n5990 = ~n1200 & n2150 ;
  assign n5991 = ( n1266 & ~n1713 ) | ( n1266 & n2158 ) | ( ~n1713 & n2158 ) ;
  assign n5992 = ( ~n1276 & n5990 ) | ( ~n1276 & n5991 ) | ( n5990 & n5991 ) ;
  assign n5993 = ( n5400 & ~n5989 ) | ( n5400 & n5992 ) | ( ~n5989 & n5992 ) ;
  assign n5994 = ( n1276 & n5489 ) | ( n1276 & ~n5991 ) | ( n5489 & ~n5991 ) ;
  assign n5995 = ( ~n5400 & n5989 ) | ( ~n5400 & n5994 ) | ( n5989 & n5994 ) ;
  assign n5996 = ( n5988 & n5993 ) | ( n5988 & ~n5995 ) | ( n5993 & ~n5995 ) ;
  assign n5997 = x243 & ~n1388 ;
  assign n5998 = n1393 | n1750 ;
  assign n5999 = n1337 & ~n1409 ;
  assign n6000 = ( n1379 & n1732 ) | ( n1379 & ~n5999 ) | ( n1732 & ~n5999 ) ;
  assign n6001 = ~n1412 & n6000 ;
  assign n6002 = ( n4484 & ~n5998 ) | ( n4484 & n6001 ) | ( ~n5998 & n6001 ) ;
  assign n6003 = n5997 & ~n6002 ;
  assign n6004 = ( n1734 & ~n4484 ) | ( n1734 & n5998 ) | ( ~n4484 & n5998 ) ;
  assign n6005 = n5997 & n6004 ;
  assign n6006 = ( n5996 & n6003 ) | ( n5996 & n6005 ) | ( n6003 & n6005 ) ;
  assign n6007 = x118 | n617 ;
  assign n6008 = ~n1383 & n6007 ;
  assign n6009 = ( ~n1464 & n1748 ) | ( ~n1464 & n6008 ) | ( n1748 & n6008 ) ;
  assign n6010 = ( ~n1466 & n1983 ) | ( ~n1466 & n6009 ) | ( n1983 & n6009 ) ;
  assign n6011 = ( ~n1992 & n2360 ) | ( ~n1992 & n6010 ) | ( n2360 & n6010 ) ;
  assign n6012 = n317 | n1481 ;
  assign n6013 = ( ~n317 & n321 ) | ( ~n317 & n2609 ) | ( n321 & n2609 ) ;
  assign n6014 = ( n5715 & n6012 ) | ( n5715 & ~n6013 ) | ( n6012 & ~n6013 ) ;
  assign n6015 = ( n2367 & ~n6012 ) | ( n2367 & n6013 ) | ( ~n6012 & n6013 ) ;
  assign n6016 = ( n6011 & ~n6014 ) | ( n6011 & n6015 ) | ( ~n6014 & n6015 ) ;
  assign n6017 = ~n355 & n4061 ;
  assign n6018 = ( n384 & n3612 ) | ( n384 & ~n6017 ) | ( n3612 & ~n6017 ) ;
  assign n6019 = ( ~n384 & n3046 ) | ( ~n384 & n6017 ) | ( n3046 & n6017 ) ;
  assign n6020 = ( n6016 & n6018 ) | ( n6016 & ~n6019 ) | ( n6018 & ~n6019 ) ;
  assign n6021 = ( n567 & n1527 ) | ( n567 & ~n2033 ) | ( n1527 & ~n2033 ) ;
  assign n6022 = n423 & ~n460 ;
  assign n6023 = ( n455 & n497 ) | ( n455 & ~n1798 ) | ( n497 & ~n1798 ) ;
  assign n6024 = ( ~n1518 & n6022 ) | ( ~n1518 & n6023 ) | ( n6022 & n6023 ) ;
  assign n6025 = ( n5434 & ~n6021 ) | ( n5434 & n6024 ) | ( ~n6021 & n6024 ) ;
  assign n6026 = ( n1518 & n5523 ) | ( n1518 & ~n6023 ) | ( n5523 & ~n6023 ) ;
  assign n6027 = ( ~n5434 & n6021 ) | ( ~n5434 & n6026 ) | ( n6021 & n6026 ) ;
  assign n6028 = ( n6020 & n6025 ) | ( n6020 & ~n6027 ) | ( n6025 & ~n6027 ) ;
  assign n6029 = x244 & ~n573 ;
  assign n6030 = n578 | n1829 ;
  assign n6031 = ~n610 & n1531 ;
  assign n6032 = ( n1539 & n1814 ) | ( n1539 & ~n6031 ) | ( n1814 & ~n6031 ) ;
  assign n6033 = ~n607 & n6032 ;
  assign n6034 = ( n4519 & ~n6030 ) | ( n4519 & n6033 ) | ( ~n6030 & n6033 ) ;
  assign n6035 = n6029 & ~n6034 ;
  assign n6036 = ( n1816 & ~n4519 ) | ( n1816 & n6030 ) | ( ~n4519 & n6030 ) ;
  assign n6037 = n6029 & n6036 ;
  assign n6038 = ( n6028 & n6035 ) | ( n6028 & n6037 ) | ( n6035 & n6037 ) ;
  assign n6039 = x119 | n1022 ;
  assign n6040 = ~n654 & n6039 ;
  assign n6041 = ( ~n641 & n645 ) | ( ~n641 & n6040 ) | ( n645 & n6040 ) ;
  assign n6042 = ( ~n652 & n2053 ) | ( ~n652 & n6041 ) | ( n2053 & n6041 ) ;
  assign n6043 = ( ~n2062 & n2404 ) | ( ~n2062 & n6042 ) | ( n2404 & n6042 ) ;
  assign n6044 = n722 | n1580 ;
  assign n6045 = ( ~n722 & n726 ) | ( ~n722 & n2644 ) | ( n726 & n2644 ) ;
  assign n6046 = ( n5749 & n6044 ) | ( n5749 & ~n6045 ) | ( n6044 & ~n6045 ) ;
  assign n6047 = ( n2411 & ~n6044 ) | ( n2411 & n6045 ) | ( ~n6044 & n6045 ) ;
  assign n6048 = ( n6043 & ~n6046 ) | ( n6043 & n6047 ) | ( ~n6046 & n6047 ) ;
  assign n6049 = ~n760 & n4098 ;
  assign n6050 = ( n789 & n3650 ) | ( n789 & ~n6049 ) | ( n3650 & ~n6049 ) ;
  assign n6051 = ( ~n789 & n3082 ) | ( ~n789 & n6049 ) | ( n3082 & n6049 ) ;
  assign n6052 = ( n6048 & n6050 ) | ( n6048 & ~n6051 ) | ( n6050 & ~n6051 ) ;
  assign n6053 = ( n972 & n1626 ) | ( n972 & ~n2103 ) | ( n1626 & ~n2103 ) ;
  assign n6054 = n828 & ~n865 ;
  assign n6055 = ( n860 & n902 ) | ( n860 & ~n1876 ) | ( n902 & ~n1876 ) ;
  assign n6056 = ( ~n1617 & n6054 ) | ( ~n1617 & n6055 ) | ( n6054 & n6055 ) ;
  assign n6057 = ( n5468 & ~n6053 ) | ( n5468 & n6056 ) | ( ~n6053 & n6056 ) ;
  assign n6058 = ( n1617 & n5557 ) | ( n1617 & ~n6055 ) | ( n5557 & ~n6055 ) ;
  assign n6059 = ( ~n5468 & n6053 ) | ( ~n5468 & n6058 ) | ( n6053 & n6058 ) ;
  assign n6060 = ( n6052 & n6057 ) | ( n6052 & ~n6059 ) | ( n6057 & ~n6059 ) ;
  assign n6061 = x245 & ~n978 ;
  assign n6062 = n983 | n1907 ;
  assign n6063 = ~n1015 & n1630 ;
  assign n6064 = ( n1638 & n1892 ) | ( n1638 & ~n6063 ) | ( n1892 & ~n6063 ) ;
  assign n6065 = ~n1012 & n6064 ;
  assign n6066 = ( n4554 & ~n6062 ) | ( n4554 & n6065 ) | ( ~n6062 & n6065 ) ;
  assign n6067 = n6061 & ~n6066 ;
  assign n6068 = ( n1894 & ~n4554 ) | ( n1894 & n6062 ) | ( ~n4554 & n6062 ) ;
  assign n6069 = n6061 & n6068 ;
  assign n6070 = ( n6060 & n6067 ) | ( n6060 & n6069 ) | ( n6067 & n6069 ) ;
  assign n6071 = x120 | n1426 ;
  assign n6072 = ~n1059 & n6071 ;
  assign n6073 = ( ~n1046 & n1050 ) | ( ~n1046 & n6072 ) | ( n1050 & n6072 ) ;
  assign n6074 = ( ~n1057 & n2123 ) | ( ~n1057 & n6073 ) | ( n2123 & n6073 ) ;
  assign n6075 = ( ~n2132 & n2448 ) | ( ~n2132 & n6074 ) | ( n2448 & n6074 ) ;
  assign n6076 = n1126 | n1678 ;
  assign n6077 = ( ~n1126 & n1130 ) | ( ~n1126 & n2679 ) | ( n1130 & n2679 ) ;
  assign n6078 = ( n5783 & n6076 ) | ( n5783 & ~n6077 ) | ( n6076 & ~n6077 ) ;
  assign n6079 = ( n2455 & ~n6076 ) | ( n2455 & n6077 ) | ( ~n6076 & n6077 ) ;
  assign n6080 = ( n6075 & ~n6078 ) | ( n6075 & n6079 ) | ( ~n6078 & n6079 ) ;
  assign n6081 = ~n1164 & n4135 ;
  assign n6082 = ( n1193 & n3688 ) | ( n1193 & ~n6081 ) | ( n3688 & ~n6081 ) ;
  assign n6083 = ( ~n1193 & n3118 ) | ( ~n1193 & n6081 ) | ( n3118 & n6081 ) ;
  assign n6084 = ( n6080 & n6082 ) | ( n6080 & ~n6083 ) | ( n6082 & ~n6083 ) ;
  assign n6085 = ( n1376 & n1724 ) | ( n1376 & ~n2173 ) | ( n1724 & ~n2173 ) ;
  assign n6086 = n1232 & ~n1269 ;
  assign n6087 = ( n1264 & n1306 ) | ( n1264 & ~n1954 ) | ( n1306 & ~n1954 ) ;
  assign n6088 = ( ~n1715 & n6086 ) | ( ~n1715 & n6087 ) | ( n6086 & n6087 ) ;
  assign n6089 = ( n5502 & ~n6085 ) | ( n5502 & n6088 ) | ( ~n6085 & n6088 ) ;
  assign n6090 = ( n1715 & n5591 ) | ( n1715 & ~n6087 ) | ( n5591 & ~n6087 ) ;
  assign n6091 = ( ~n5502 & n6085 ) | ( ~n5502 & n6090 ) | ( n6085 & n6090 ) ;
  assign n6092 = ( n6084 & n6089 ) | ( n6084 & ~n6091 ) | ( n6089 & ~n6091 ) ;
  assign n6093 = x246 & ~n1382 ;
  assign n6094 = n1387 | n1985 ;
  assign n6095 = ~n1419 & n1728 ;
  assign n6096 = ( n1736 & n1970 ) | ( n1736 & ~n6095 ) | ( n1970 & ~n6095 ) ;
  assign n6097 = ~n1416 & n6096 ;
  assign n6098 = ( n4589 & ~n6094 ) | ( n4589 & n6097 ) | ( ~n6094 & n6097 ) ;
  assign n6099 = n6093 & ~n6098 ;
  assign n6100 = ( n1972 & ~n4589 ) | ( n1972 & n6094 ) | ( ~n4589 & n6094 ) ;
  assign n6101 = n6093 & n6100 ;
  assign n6102 = ( n6092 & n6099 ) | ( n6092 & n6101 ) | ( n6099 & n6101 ) ;
  assign n6103 = x121 | n642 ;
  assign n6104 = ~n1463 & n6103 ;
  assign n6105 = ( ~n1450 & n1454 ) | ( ~n1450 & n6104 ) | ( n1454 & n6104 ) ;
  assign n6106 = ( ~n1461 & n2193 ) | ( ~n1461 & n6105 ) | ( n2193 & n6105 ) ;
  assign n6107 = ( ~n2201 & n2492 ) | ( ~n2201 & n6106 ) | ( n2492 & n6106 ) ;
  assign n6108 = ( ~n304 & n322 ) | ( ~n304 & n2714 ) | ( n322 & n2714 ) ;
  assign n6109 = ( n320 & n5817 ) | ( n320 & ~n6108 ) | ( n5817 & ~n6108 ) ;
  assign n6110 = ( ~n320 & n2499 ) | ( ~n320 & n6108 ) | ( n2499 & n6108 ) ;
  assign n6111 = ( n6107 & ~n6109 ) | ( n6107 & n6110 ) | ( ~n6109 & n6110 ) ;
  assign n6112 = ~n401 & n4172 ;
  assign n6113 = ( n1499 & n3726 ) | ( n1499 & ~n6112 ) | ( n3726 & ~n6112 ) ;
  assign n6114 = ( ~n1499 & n3154 ) | ( ~n1499 & n6112 ) | ( n3154 & n6112 ) ;
  assign n6115 = ( n6111 & n6113 ) | ( n6111 & ~n6114 ) | ( n6113 & ~n6114 ) ;
  assign n6116 = ( n568 & n1808 ) | ( n568 & ~n2229 ) | ( n1808 & ~n2229 ) ;
  assign n6117 = ~n445 & n1508 ;
  assign n6118 = ( n501 & n1513 ) | ( n501 & ~n2025 ) | ( n1513 & ~n2025 ) ;
  assign n6119 = ( ~n1800 & n6117 ) | ( ~n1800 & n6118 ) | ( n6117 & n6118 ) ;
  assign n6120 = ( n5536 & ~n6116 ) | ( n5536 & n6119 ) | ( ~n6116 & n6119 ) ;
  assign n6121 = ( n1800 & n5625 ) | ( n1800 & ~n6118 ) | ( n5625 & ~n6118 ) ;
  assign n6122 = ( ~n5536 & n6116 ) | ( ~n5536 & n6121 ) | ( n6116 & n6121 ) ;
  assign n6123 = ( n6115 & n6120 ) | ( n6115 & ~n6122 ) | ( n6120 & ~n6122 ) ;
  assign n6124 = x247 & ~n653 ;
  assign n6125 = n619 | n2055 ;
  assign n6126 = ~n591 & n1811 ;
  assign n6127 = ( n1818 & n2041 ) | ( n1818 & ~n6126 ) | ( n2041 & ~n6126 ) ;
  assign n6128 = ~n594 & n6127 ;
  assign n6129 = ( n4624 & ~n6125 ) | ( n4624 & n6128 ) | ( ~n6125 & n6128 ) ;
  assign n6130 = n6124 & ~n6129 ;
  assign n6131 = ( n2043 & ~n4624 ) | ( n2043 & n6125 ) | ( ~n4624 & n6125 ) ;
  assign n6132 = n6124 & n6131 ;
  assign n6133 = ( n6123 & n6130 ) | ( n6123 & n6132 ) | ( n6130 & n6132 ) ;
  assign n6134 = x122 | n1047 ;
  assign n6135 = ~n640 & n6134 ;
  assign n6136 = ( ~n638 & n649 ) | ( ~n638 & n6135 ) | ( n649 & n6135 ) ;
  assign n6137 = ( ~n1565 & n2248 ) | ( ~n1565 & n6136 ) | ( n2248 & n6136 ) ;
  assign n6138 = ( ~n2257 & n2530 ) | ( ~n2257 & n6137 ) | ( n2530 & n6137 ) ;
  assign n6139 = ( ~n709 & n727 ) | ( ~n709 & n2748 ) | ( n727 & n2748 ) ;
  assign n6140 = ( n725 & n5850 ) | ( n725 & ~n6139 ) | ( n5850 & ~n6139 ) ;
  assign n6141 = ( ~n725 & n2536 ) | ( ~n725 & n6139 ) | ( n2536 & n6139 ) ;
  assign n6142 = ( n6138 & ~n6140 ) | ( n6138 & n6141 ) | ( ~n6140 & n6141 ) ;
  assign n6143 = ~n806 & n4209 ;
  assign n6144 = ( n1598 & n3764 ) | ( n1598 & ~n6143 ) | ( n3764 & ~n6143 ) ;
  assign n6145 = ( ~n1598 & n3190 ) | ( ~n1598 & n6143 ) | ( n3190 & n6143 ) ;
  assign n6146 = ( n6142 & n6144 ) | ( n6142 & ~n6145 ) | ( n6144 & ~n6145 ) ;
  assign n6147 = ( n973 & n1886 ) | ( n973 & ~n2285 ) | ( n1886 & ~n2285 ) ;
  assign n6148 = ~n850 & n1607 ;
  assign n6149 = ( n906 & n1612 ) | ( n906 & ~n2095 ) | ( n1612 & ~n2095 ) ;
  assign n6150 = ( ~n1878 & n6148 ) | ( ~n1878 & n6149 ) | ( n6148 & n6149 ) ;
  assign n6151 = ( n5570 & ~n6147 ) | ( n5570 & n6150 ) | ( ~n6147 & n6150 ) ;
  assign n6152 = ( n1878 & n5659 ) | ( n1878 & ~n6149 ) | ( n5659 & ~n6149 ) ;
  assign n6153 = ( ~n5570 & n6147 ) | ( ~n5570 & n6152 ) | ( n6147 & n6152 ) ;
  assign n6154 = ( n6146 & n6151 ) | ( n6146 & ~n6153 ) | ( n6151 & ~n6153 ) ;
  assign n6155 = x248 & ~n1058 ;
  assign n6156 = n1024 | n2125 ;
  assign n6157 = ~n996 & n1889 ;
  assign n6158 = ( n1896 & n2111 ) | ( n1896 & ~n6157 ) | ( n2111 & ~n6157 ) ;
  assign n6159 = ~n999 & n6158 ;
  assign n6160 = ( n4659 & ~n6156 ) | ( n4659 & n6159 ) | ( ~n6156 & n6159 ) ;
  assign n6161 = n6155 & ~n6160 ;
  assign n6162 = ( n2113 & ~n4659 ) | ( n2113 & n6156 ) | ( ~n4659 & n6156 ) ;
  assign n6163 = n6155 & n6162 ;
  assign n6164 = ( n6154 & n6161 ) | ( n6154 & n6163 ) | ( n6161 & n6163 ) ;
  assign n6165 = x123 | n1451 ;
  assign n6166 = ~n1045 & n6165 ;
  assign n6167 = ( ~n1043 & n1054 ) | ( ~n1043 & n6166 ) | ( n1054 & n6166 ) ;
  assign n6168 = ( ~n1664 & n2304 ) | ( ~n1664 & n6167 ) | ( n2304 & n6167 ) ;
  assign n6169 = ( ~n2313 & n2567 ) | ( ~n2313 & n6168 ) | ( n2567 & n6168 ) ;
  assign n6170 = ( ~n1113 & n1131 ) | ( ~n1113 & n2787 ) | ( n1131 & n2787 ) ;
  assign n6171 = ( n1129 & n5883 ) | ( n1129 & ~n6170 ) | ( n5883 & ~n6170 ) ;
  assign n6172 = ( ~n1129 & n2573 ) | ( ~n1129 & n6170 ) | ( n2573 & n6170 ) ;
  assign n6173 = ( n6169 & ~n6171 ) | ( n6169 & n6172 ) | ( ~n6171 & n6172 ) ;
  assign n6174 = ~n1210 & n4246 ;
  assign n6175 = ( n1696 & n3802 ) | ( n1696 & ~n6174 ) | ( n3802 & ~n6174 ) ;
  assign n6176 = ( ~n1696 & n3226 ) | ( ~n1696 & n6174 ) | ( n3226 & n6174 ) ;
  assign n6177 = ( n6173 & n6175 ) | ( n6173 & ~n6176 ) | ( n6175 & ~n6176 ) ;
  assign n6178 = ( n1377 & n1964 ) | ( n1377 & ~n2341 ) | ( n1964 & ~n2341 ) ;
  assign n6179 = ~n1254 & n1705 ;
  assign n6180 = ( n1310 & n1710 ) | ( n1310 & ~n2165 ) | ( n1710 & ~n2165 ) ;
  assign n6181 = ( ~n1956 & n6179 ) | ( ~n1956 & n6180 ) | ( n6179 & n6180 ) ;
  assign n6182 = ( n5604 & ~n6178 ) | ( n5604 & n6181 ) | ( ~n6178 & n6181 ) ;
  assign n6183 = ( n1956 & n5693 ) | ( n1956 & ~n6180 ) | ( n5693 & ~n6180 ) ;
  assign n6184 = ( ~n5604 & n6178 ) | ( ~n5604 & n6183 ) | ( n6178 & n6183 ) ;
  assign n6185 = ( n6177 & n6182 ) | ( n6177 & ~n6184 ) | ( n6182 & ~n6184 ) ;
  assign n6186 = x249 & ~n1462 ;
  assign n6187 = n1428 | n2195 ;
  assign n6188 = ~n1400 & n1967 ;
  assign n6189 = ( n1974 & n2181 ) | ( n1974 & ~n6188 ) | ( n2181 & ~n6188 ) ;
  assign n6190 = ~n1403 & n6189 ;
  assign n6191 = ( n4694 & ~n6187 ) | ( n4694 & n6190 ) | ( ~n6187 & n6190 ) ;
  assign n6192 = n6186 & ~n6191 ;
  assign n6193 = ( n2183 & ~n4694 ) | ( n2183 & n6187 ) | ( ~n4694 & n6187 ) ;
  assign n6194 = n6186 & n6193 ;
  assign n6195 = ( n6185 & n6192 ) | ( n6185 & n6194 ) | ( n6192 & n6194 ) ;
  assign n6196 = x124 | n646 ;
  assign n6197 = ~n1449 & n6196 ;
  assign n6198 = ( ~n1447 & n1458 ) | ( ~n1447 & n6197 ) | ( n1458 & n6197 ) ;
  assign n6199 = ( ~n1759 & n2360 ) | ( ~n1759 & n6198 ) | ( n2360 & n6198 ) ;
  assign n6200 = ( n281 & ~n2369 ) | ( n281 & n6199 ) | ( ~n2369 & n6199 ) ;
  assign n6201 = ( n323 & ~n333 ) | ( n323 & n348 ) | ( ~n333 & n348 ) ;
  assign n6202 = ( n1485 & n5916 ) | ( n1485 & ~n6201 ) | ( n5916 & ~n6201 ) ;
  assign n6203 = ( ~n1485 & n2609 ) | ( ~n1485 & n6201 ) | ( n2609 & n6201 ) ;
  assign n6204 = ( n6200 & ~n6202 ) | ( n6200 & n6203 ) | ( ~n6202 & n6203 ) ;
  assign n6205 = ~n405 & n4283 ;
  assign n6206 = ( n1783 & n3840 ) | ( n1783 & ~n6205 ) | ( n3840 & ~n6205 ) ;
  assign n6207 = ( ~n1783 & n3262 ) | ( ~n1783 & n6205 ) | ( n3262 & n6205 ) ;
  assign n6208 = ( n6204 & n6206 ) | ( n6204 & ~n6207 ) | ( n6206 & ~n6207 ) ;
  assign n6209 = ( ~n539 & n540 ) | ( ~n539 & n2030 ) | ( n540 & n2030 ) ;
  assign n6210 = ~n442 & n1791 ;
  assign n6211 = ( n485 & n1795 ) | ( n485 & ~n2221 ) | ( n1795 & ~n2221 ) ;
  assign n6212 = ( ~n2027 & n6210 ) | ( ~n2027 & n6211 ) | ( n6210 & n6211 ) ;
  assign n6213 = ( n5638 & ~n6209 ) | ( n5638 & n6212 ) | ( ~n6209 & n6212 ) ;
  assign n6214 = ( n2027 & n5727 ) | ( n2027 & ~n6211 ) | ( n5727 & ~n6211 ) ;
  assign n6215 = ( ~n5638 & n6209 ) | ( ~n5638 & n6214 ) | ( n6209 & n6214 ) ;
  assign n6216 = ( n6208 & n6213 ) | ( n6208 & ~n6215 ) | ( n6213 & ~n6215 ) ;
  assign n6217 = x250 & ~n639 ;
  assign n6218 = n644 | n2249 ;
  assign n6219 = ~n588 & n2038 ;
  assign n6220 = ( n596 & n2045 ) | ( n596 & ~n6219 ) | ( n2045 & ~n6219 ) ;
  assign n6221 = ~n584 & n6220 ;
  assign n6222 = ( n4729 & ~n6218 ) | ( n4729 & n6221 ) | ( ~n6218 & n6221 ) ;
  assign n6223 = n6217 & ~n6222 ;
  assign n6224 = ( n2237 & ~n4729 ) | ( n2237 & n6218 ) | ( ~n4729 & n6218 ) ;
  assign n6225 = n6217 & n6224 ;
  assign n6226 = ( n6216 & n6223 ) | ( n6216 & n6225 ) | ( n6223 & n6225 ) ;
  assign n6227 = x125 | n1051 ;
  assign n6228 = ~n637 & n6227 ;
  assign n6229 = ( ~n1561 & n1562 ) | ( ~n1561 & n6228 ) | ( n1562 & n6228 ) ;
  assign n6230 = ( ~n1837 & n2404 ) | ( ~n1837 & n6229 ) | ( n2404 & n6229 ) ;
  assign n6231 = ( n686 & ~n2413 ) | ( n686 & n6230 ) | ( ~n2413 & n6230 ) ;
  assign n6232 = ( n728 & ~n738 ) | ( n728 & n753 ) | ( ~n738 & n753 ) ;
  assign n6233 = ( n1584 & n5948 ) | ( n1584 & ~n6232 ) | ( n5948 & ~n6232 ) ;
  assign n6234 = ( ~n1584 & n2644 ) | ( ~n1584 & n6232 ) | ( n2644 & n6232 ) ;
  assign n6235 = ( n6231 & ~n6233 ) | ( n6231 & n6234 ) | ( ~n6233 & n6234 ) ;
  assign n6236 = ~n810 & n4319 ;
  assign n6237 = ( n1861 & n3878 ) | ( n1861 & ~n6236 ) | ( n3878 & ~n6236 ) ;
  assign n6238 = ( ~n1861 & n3301 ) | ( ~n1861 & n6236 ) | ( n3301 & n6236 ) ;
  assign n6239 = ( n6235 & n6237 ) | ( n6235 & ~n6238 ) | ( n6237 & ~n6238 ) ;
  assign n6240 = ( ~n944 & n945 ) | ( ~n944 & n2100 ) | ( n945 & n2100 ) ;
  assign n6241 = ~n847 & n1869 ;
  assign n6242 = ( n890 & n1873 ) | ( n890 & ~n2277 ) | ( n1873 & ~n2277 ) ;
  assign n6243 = ( ~n2097 & n6241 ) | ( ~n2097 & n6242 ) | ( n6241 & n6242 ) ;
  assign n6244 = ( n5672 & ~n6240 ) | ( n5672 & n6243 ) | ( ~n6240 & n6243 ) ;
  assign n6245 = ( n2097 & n5761 ) | ( n2097 & ~n6242 ) | ( n5761 & ~n6242 ) ;
  assign n6246 = ( ~n5672 & n6240 ) | ( ~n5672 & n6245 ) | ( n6240 & n6245 ) ;
  assign n6247 = ( n6239 & n6244 ) | ( n6239 & ~n6246 ) | ( n6244 & ~n6246 ) ;
  assign n6248 = x251 & ~n1044 ;
  assign n6249 = n1049 | n2305 ;
  assign n6250 = ~n993 & n2108 ;
  assign n6251 = ( n1001 & n2115 ) | ( n1001 & ~n6250 ) | ( n2115 & ~n6250 ) ;
  assign n6252 = ~n989 & n6251 ;
  assign n6253 = ( n4764 & ~n6249 ) | ( n4764 & n6252 ) | ( ~n6249 & n6252 ) ;
  assign n6254 = n6248 & ~n6253 ;
  assign n6255 = ( n2293 & ~n4764 ) | ( n2293 & n6249 ) | ( ~n4764 & n6249 ) ;
  assign n6256 = n6248 & n6255 ;
  assign n6257 = ( n6247 & n6254 ) | ( n6247 & n6256 ) | ( n6254 & n6256 ) ;
  assign n6258 = x126 | n1455 ;
  assign n6259 = ~n1042 & n6258 ;
  assign n6260 = ( ~n1660 & n1661 ) | ( ~n1660 & n6259 ) | ( n1661 & n6259 ) ;
  assign n6261 = ( ~n1915 & n2448 ) | ( ~n1915 & n6260 ) | ( n2448 & n6260 ) ;
  assign n6262 = ( n1090 & ~n2457 ) | ( n1090 & n6261 ) | ( ~n2457 & n6261 ) ;
  assign n6263 = ( n1132 & ~n1142 ) | ( n1132 & n1157 ) | ( ~n1142 & n1157 ) ;
  assign n6264 = ( n1682 & n5980 ) | ( n1682 & ~n6263 ) | ( n5980 & ~n6263 ) ;
  assign n6265 = ( ~n1682 & n2679 ) | ( ~n1682 & n6263 ) | ( n2679 & n6263 ) ;
  assign n6266 = ( n6262 & ~n6264 ) | ( n6262 & n6265 ) | ( ~n6264 & n6265 ) ;
  assign n6267 = ~n1214 & n4355 ;
  assign n6268 = ( n1939 & n3916 ) | ( n1939 & ~n6267 ) | ( n3916 & ~n6267 ) ;
  assign n6269 = ( ~n1939 & n3340 ) | ( ~n1939 & n6267 ) | ( n3340 & n6267 ) ;
  assign n6270 = ( n6266 & n6268 ) | ( n6266 & ~n6269 ) | ( n6268 & ~n6269 ) ;
  assign n6271 = ( ~n1348 & n1349 ) | ( ~n1348 & n2170 ) | ( n1349 & n2170 ) ;
  assign n6272 = ~n1251 & n1947 ;
  assign n6273 = ( n1294 & n1951 ) | ( n1294 & ~n2333 ) | ( n1951 & ~n2333 ) ;
  assign n6274 = ( ~n2167 & n6272 ) | ( ~n2167 & n6273 ) | ( n6272 & n6273 ) ;
  assign n6275 = ( n5706 & ~n6271 ) | ( n5706 & n6274 ) | ( ~n6271 & n6274 ) ;
  assign n6276 = ( n2167 & n5795 ) | ( n2167 & ~n6273 ) | ( n5795 & ~n6273 ) ;
  assign n6277 = ( ~n5706 & n6271 ) | ( ~n5706 & n6276 ) | ( n6271 & n6276 ) ;
  assign n6278 = ( n6270 & n6275 ) | ( n6270 & ~n6277 ) | ( n6275 & ~n6277 ) ;
  assign n6279 = x252 & ~n1448 ;
  assign n6280 = n1453 | n2361 ;
  assign n6281 = ~n1397 & n2178 ;
  assign n6282 = ( n1405 & n2185 ) | ( n1405 & ~n6281 ) | ( n2185 & ~n6281 ) ;
  assign n6283 = ~n1393 & n6282 ;
  assign n6284 = ( n4799 & ~n6280 ) | ( n4799 & n6283 ) | ( ~n6280 & n6283 ) ;
  assign n6285 = n6279 & ~n6284 ;
  assign n6286 = ( n2349 & ~n4799 ) | ( n2349 & n6280 ) | ( ~n4799 & n6280 ) ;
  assign n6287 = n6279 & n6286 ;
  assign n6288 = ( n6278 & n6285 ) | ( n6278 & n6287 ) | ( n6285 & n6287 ) ;
  assign n6289 = x127 | n633 ;
  assign n6290 = ~n1446 & n6289 ;
  assign n6291 = ( ~n1755 & n1756 ) | ( ~n1755 & n6290 ) | ( n1756 & n6290 ) ;
  assign n6292 = ( ~n1991 & n2492 ) | ( ~n1991 & n6291 ) | ( n2492 & n6291 ) ;
  assign n6293 = ( n1477 & ~n2501 ) | ( n1477 & n6292 ) | ( ~n2501 & n6292 ) ;
  assign n6294 = ( ~n340 & n349 ) | ( ~n340 & n1486 ) | ( n349 & n1486 ) ;
  assign n6295 = ( n1772 & n6012 ) | ( n1772 & ~n6294 ) | ( n6012 & ~n6294 ) ;
  assign n6296 = ( ~n1772 & n2714 ) | ( ~n1772 & n6294 ) | ( n2714 & n6294 ) ;
  assign n6297 = ( n6293 & ~n6295 ) | ( n6293 & n6296 ) | ( ~n6295 & n6296 ) ;
  assign n6298 = ~n394 & n4391 ;
  assign n6299 = ( n2010 & n3954 ) | ( n2010 & ~n6298 ) | ( n3954 & ~n6298 ) ;
  assign n6300 = ( ~n2010 & n3379 ) | ( ~n2010 & n6298 ) | ( n3379 & n6298 ) ;
  assign n6301 = ( n6297 & n6299 ) | ( n6297 & ~n6300 ) | ( n6299 & ~n6300 ) ;
  assign n6302 = ( n560 & ~n1532 ) | ( n560 & n2227 ) | ( ~n1532 & n2227 ) ;
  assign n6303 = ~n433 & n2018 ;
  assign n6304 = ( ~n510 & n511 ) | ( ~n510 & n2022 ) | ( n511 & n2022 ) ;
  assign n6305 = ( ~n2224 & n6303 ) | ( ~n2224 & n6304 ) | ( n6303 & n6304 ) ;
  assign n6306 = ( n5740 & ~n6302 ) | ( n5740 & n6305 ) | ( ~n6302 & n6305 ) ;
  assign n6307 = ( n2224 & n5829 ) | ( n2224 & ~n6304 ) | ( n5829 & ~n6304 ) ;
  assign n6308 = ( ~n5740 & n6302 ) | ( ~n5740 & n6307 ) | ( n6302 & n6307 ) ;
  assign n6309 = ( n6301 & n6306 ) | ( n6301 & ~n6308 ) | ( n6306 & ~n6308 ) ;
  assign n6310 = x253 & ~n636 ;
  assign n6311 = n648 | n2405 ;
  assign n6312 = ~n581 & n622 ;
  assign n6313 = ( n1542 & n2239 ) | ( n1542 & ~n6312 ) | ( n2239 & ~n6312 ) ;
  assign n6314 = ~n578 & n6313 ;
  assign n6315 = ( n4834 & ~n6311 ) | ( n4834 & n6314 ) | ( ~n6311 & n6314 ) ;
  assign n6316 = n6310 & ~n6315 ;
  assign n6317 = ( n2396 & ~n4834 ) | ( n2396 & n6311 ) | ( ~n4834 & n6311 ) ;
  assign n6318 = n6310 & n6317 ;
  assign n6319 = ( n6309 & n6316 ) | ( n6309 & n6318 ) | ( n6316 & n6318 ) ;
  assign n6320 = x0 | n1038 ;
  assign n6321 = ~n1560 & n6320 ;
  assign n6322 = ( ~n1833 & n1834 ) | ( ~n1833 & n6321 ) | ( n1834 & n6321 ) ;
  assign n6323 = ( ~n2061 & n2530 ) | ( ~n2061 & n6322 ) | ( n2530 & n6322 ) ;
  assign n6324 = ( n1576 & ~n2538 ) | ( n1576 & n6323 ) | ( ~n2538 & n6323 ) ;
  assign n6325 = ( ~n745 & n754 ) | ( ~n745 & n1585 ) | ( n754 & n1585 ) ;
  assign n6326 = ( n1850 & n6044 ) | ( n1850 & ~n6325 ) | ( n6044 & ~n6325 ) ;
  assign n6327 = ( ~n1850 & n2748 ) | ( ~n1850 & n6325 ) | ( n2748 & n6325 ) ;
  assign n6328 = ( n6324 & ~n6326 ) | ( n6324 & n6327 ) | ( ~n6326 & n6327 ) ;
  assign n6329 = ~n799 & n4427 ;
  assign n6330 = ( n2080 & n3992 ) | ( n2080 & ~n6329 ) | ( n3992 & ~n6329 ) ;
  assign n6331 = ( ~n2080 & n3418 ) | ( ~n2080 & n6329 ) | ( n3418 & n6329 ) ;
  assign n6332 = ( n6328 & n6330 ) | ( n6328 & ~n6331 ) | ( n6330 & ~n6331 ) ;
  assign n6333 = ( n965 & ~n1631 ) | ( n965 & n2283 ) | ( ~n1631 & n2283 ) ;
  assign n6334 = ~n838 & n2088 ;
  assign n6335 = ( ~n915 & n916 ) | ( ~n915 & n2092 ) | ( n916 & n2092 ) ;
  assign n6336 = ( ~n2280 & n6334 ) | ( ~n2280 & n6335 ) | ( n6334 & n6335 ) ;
  assign n6337 = ( n5774 & ~n6333 ) | ( n5774 & n6336 ) | ( ~n6333 & n6336 ) ;
  assign n6338 = ( n2280 & n5862 ) | ( n2280 & ~n6335 ) | ( n5862 & ~n6335 ) ;
  assign n6339 = ( ~n5774 & n6333 ) | ( ~n5774 & n6338 ) | ( n6333 & n6338 ) ;
  assign n6340 = ( n6332 & n6337 ) | ( n6332 & ~n6339 ) | ( n6337 & ~n6339 ) ;
  assign n6341 = x254 & ~n1041 ;
  assign n6342 = n1053 | n2449 ;
  assign n6343 = ~n986 & n1027 ;
  assign n6344 = ( n1641 & n2295 ) | ( n1641 & ~n6343 ) | ( n2295 & ~n6343 ) ;
  assign n6345 = ~n983 & n6344 ;
  assign n6346 = ( n4869 & ~n6342 ) | ( n4869 & n6345 ) | ( ~n6342 & n6345 ) ;
  assign n6347 = n6341 & ~n6346 ;
  assign n6348 = ( n2440 & ~n4869 ) | ( n2440 & n6342 ) | ( ~n4869 & n6342 ) ;
  assign n6349 = n6341 & n6348 ;
  assign n6350 = ( n6340 & n6347 ) | ( n6340 & n6349 ) | ( n6347 & n6349 ) ;
  assign n6351 = x1 | n1442 ;
  assign n6352 = ~n1659 & n6351 ;
  assign n6353 = ( ~n1911 & n1912 ) | ( ~n1911 & n6352 ) | ( n1912 & n6352 ) ;
  assign n6354 = ( ~n2131 & n2567 ) | ( ~n2131 & n6353 ) | ( n2567 & n6353 ) ;
  assign n6355 = ( n1674 & ~n2575 ) | ( n1674 & n6354 ) | ( ~n2575 & n6354 ) ;
  assign n6356 = ( ~n1149 & n1158 ) | ( ~n1149 & n1683 ) | ( n1158 & n1683 ) ;
  assign n6357 = ( n1928 & n6076 ) | ( n1928 & ~n6356 ) | ( n6076 & ~n6356 ) ;
  assign n6358 = ( ~n1928 & n2787 ) | ( ~n1928 & n6356 ) | ( n2787 & n6356 ) ;
  assign n6359 = ( n6355 & ~n6357 ) | ( n6355 & n6358 ) | ( ~n6357 & n6358 ) ;
  assign n6360 = ~n1203 & n4463 ;
  assign n6361 = ( n2150 & n4030 ) | ( n2150 & ~n6360 ) | ( n4030 & ~n6360 ) ;
  assign n6362 = ( ~n2150 & n3457 ) | ( ~n2150 & n6360 ) | ( n3457 & n6360 ) ;
  assign n6363 = ( n6359 & n6361 ) | ( n6359 & ~n6362 ) | ( n6361 & ~n6362 ) ;
  assign n6364 = ( n1369 & ~n1729 ) | ( n1369 & n2339 ) | ( ~n1729 & n2339 ) ;
  assign n6365 = ~n1242 & n2158 ;
  assign n6366 = ( ~n1319 & n1320 ) | ( ~n1319 & n2162 ) | ( n1320 & n2162 ) ;
  assign n6367 = ( ~n2336 & n6365 ) | ( ~n2336 & n6366 ) | ( n6365 & n6366 ) ;
  assign n6368 = ( n5808 & ~n6364 ) | ( n5808 & n6367 ) | ( ~n6364 & n6367 ) ;
  assign n6369 = ( n2336 & n5895 ) | ( n2336 & ~n6366 ) | ( n5895 & ~n6366 ) ;
  assign n6370 = ( ~n5808 & n6364 ) | ( ~n5808 & n6369 ) | ( n6364 & n6369 ) ;
  assign n6371 = ( n6363 & n6368 ) | ( n6363 & ~n6370 ) | ( n6368 & ~n6370 ) ;
  assign n6372 = x255 & ~n1445 ;
  assign n6373 = n1457 | n2493 ;
  assign n6374 = ~n1390 & n1431 ;
  assign n6375 = ( n1739 & n2351 ) | ( n1739 & ~n6374 ) | ( n2351 & ~n6374 ) ;
  assign n6376 = ~n1387 & n6375 ;
  assign n6377 = ( n4904 & ~n6373 ) | ( n4904 & n6376 ) | ( ~n6373 & n6376 ) ;
  assign n6378 = n6372 & ~n6377 ;
  assign n6379 = ( n2484 & ~n4904 ) | ( n2484 & n6373 ) | ( ~n4904 & n6373 ) ;
  assign n6380 = n6372 & n6379 ;
  assign n6381 = ( n6371 & n6378 ) | ( n6371 & n6380 ) | ( n6378 & n6380 ) ;
  assign n6382 = n640 | n669 ;
  assign n6383 = n701 | n711 ;
  assign n6384 = n6382 | n6383 ;
  assign n6385 = n522 | n609 ;
  assign n6386 = n574 | n587 ;
  assign n6387 = n6385 | n6386 ;
  assign n6388 = n6384 | n6387 ;
  assign n6389 = n795 | n812 ;
  assign n6390 = n837 | n849 ;
  assign n6391 = n6389 | n6390 ;
  assign n6392 = n708 | n744 ;
  assign n6393 = n762 | n769 ;
  assign n6394 = n6392 | n6393 ;
  assign n6395 = n6391 | n6394 ;
  assign n6396 = n6388 | n6395 ;
  assign n6397 = n326 | n332 ;
  assign n6398 = n371 | n397 ;
  assign n6399 = n6397 | n6398 ;
  assign n6400 = n261 | n272 ;
  assign n6401 = n288 | n316 ;
  assign n6402 = n6400 | n6401 ;
  assign n6403 = n6399 | n6402 ;
  assign n6404 = n489 | n505 ;
  assign n6405 = n533 | n545 ;
  assign n6406 = n6404 | n6405 ;
  assign n6407 = n412 | n459 ;
  assign n6408 = n426 | n441 ;
  assign n6409 = n6407 | n6408 ;
  assign n6410 = n6406 | n6409 ;
  assign n6411 = n6403 | n6410 ;
  assign n6412 = n6396 | n6411 ;
  assign n6413 = n1235 | n1250 ;
  assign n6414 = n1298 | n1314 ;
  assign n6415 = n6413 | n6414 ;
  assign n6416 = n1180 | n1206 ;
  assign n6417 = n1221 | n1268 ;
  assign n6418 = n6416 | n6417 ;
  assign n6419 = n6415 | n6418 ;
  assign n6420 = n1383 | n1396 ;
  assign n6421 = n1449 | n1560 ;
  assign n6422 = n6420 | n6421 ;
  assign n6423 = n1342 | n1354 ;
  assign n6424 = n1331 | n1418 ;
  assign n6425 = n6423 | n6424 ;
  assign n6426 = n6422 | n6425 ;
  assign n6427 = n6419 | n6426 ;
  assign n6428 = n963 | n1004 ;
  assign n6429 = n985 | n995 ;
  assign n6430 = n6428 | n6429 ;
  assign n6431 = n885 | n897 ;
  assign n6432 = n875 | n947 ;
  assign n6433 = n6431 | n6432 ;
  assign n6434 = n6430 | n6433 ;
  assign n6435 = n1097 | n1125 ;
  assign n6436 = n1135 | n1141 ;
  assign n6437 = n6435 | n6436 ;
  assign n6438 = n1042 | n1059 ;
  assign n6439 = n1070 | n1081 ;
  assign n6440 = n6438 | n6439 ;
  assign n6441 = n6437 | n6440 ;
  assign n6442 = n6434 | n6441 ;
  assign n6443 = n6427 | n6442 ;
  assign n6444 = n6412 | n6443 ;
  assign y0 = n661 ;
  assign y1 = n1066 ;
  assign y2 = n1470 ;
  assign y3 = n1569 ;
  assign y4 = n1668 ;
  assign y5 = n1763 ;
  assign y6 = n1841 ;
  assign y7 = n1919 ;
  assign y8 = n1995 ;
  assign y9 = n2065 ;
  assign y10 = n2135 ;
  assign y11 = n2204 ;
  assign y12 = n2260 ;
  assign y13 = n2316 ;
  assign y14 = n2372 ;
  assign y15 = n2416 ;
  assign y16 = n2460 ;
  assign y17 = n2504 ;
  assign y18 = n2541 ;
  assign y19 = n2578 ;
  assign y20 = n2613 ;
  assign y21 = n2648 ;
  assign y22 = n2683 ;
  assign y23 = n2718 ;
  assign y24 = n2757 ;
  assign y25 = n2796 ;
  assign y26 = n2834 ;
  assign y27 = n2871 ;
  assign y28 = n2908 ;
  assign y29 = n2945 ;
  assign y30 = n2981 ;
  assign y31 = n3017 ;
  assign y32 = n3053 ;
  assign y33 = n3089 ;
  assign y34 = n3125 ;
  assign y35 = n3161 ;
  assign y36 = n3197 ;
  assign y37 = n3233 ;
  assign y38 = n3269 ;
  assign y39 = n3308 ;
  assign y40 = n3347 ;
  assign y41 = n3386 ;
  assign y42 = n3425 ;
  assign y43 = n3464 ;
  assign y44 = n3502 ;
  assign y45 = n3540 ;
  assign y46 = n3578 ;
  assign y47 = n3616 ;
  assign y48 = n3654 ;
  assign y49 = n3692 ;
  assign y50 = n3730 ;
  assign y51 = n3768 ;
  assign y52 = n3806 ;
  assign y53 = n3844 ;
  assign y54 = n3882 ;
  assign y55 = n3920 ;
  assign y56 = n3958 ;
  assign y57 = n3996 ;
  assign y58 = n4034 ;
  assign y59 = n4071 ;
  assign y60 = n4108 ;
  assign y61 = n4145 ;
  assign y62 = n4182 ;
  assign y63 = n4219 ;
  assign y64 = n4256 ;
  assign y65 = n4292 ;
  assign y66 = n4328 ;
  assign y67 = n4364 ;
  assign y68 = n4400 ;
  assign y69 = n4436 ;
  assign y70 = n4472 ;
  assign y71 = n4507 ;
  assign y72 = n4542 ;
  assign y73 = n4577 ;
  assign y74 = n4612 ;
  assign y75 = n4647 ;
  assign y76 = n4682 ;
  assign y77 = n4717 ;
  assign y78 = n4752 ;
  assign y79 = n4787 ;
  assign y80 = n4822 ;
  assign y81 = n4857 ;
  assign y82 = n4892 ;
  assign y83 = n4927 ;
  assign y84 = n4961 ;
  assign y85 = n4995 ;
  assign y86 = n5029 ;
  assign y87 = n5063 ;
  assign y88 = n5097 ;
  assign y89 = n5131 ;
  assign y90 = n5165 ;
  assign y91 = n5199 ;
  assign y92 = n5233 ;
  assign y93 = n5267 ;
  assign y94 = n5301 ;
  assign y95 = n5335 ;
  assign y96 = n5369 ;
  assign y97 = n5403 ;
  assign y98 = n5437 ;
  assign y99 = n5471 ;
  assign y100 = n5505 ;
  assign y101 = n5539 ;
  assign y102 = n5573 ;
  assign y103 = n5607 ;
  assign y104 = n5641 ;
  assign y105 = n5675 ;
  assign y106 = n5709 ;
  assign y107 = n5743 ;
  assign y108 = n5777 ;
  assign y109 = n5811 ;
  assign y110 = n5844 ;
  assign y111 = n5877 ;
  assign y112 = n5910 ;
  assign y113 = n5942 ;
  assign y114 = n5974 ;
  assign y115 = n6006 ;
  assign y116 = n6038 ;
  assign y117 = n6070 ;
  assign y118 = n6102 ;
  assign y119 = n6133 ;
  assign y120 = n6164 ;
  assign y121 = n6195 ;
  assign y122 = n6226 ;
  assign y123 = n6257 ;
  assign y124 = n6288 ;
  assign y125 = n6319 ;
  assign y126 = n6350 ;
  assign y127 = n6381 ;
  assign y128 = n6444 ;
endmodule
