module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 , x147 , x148 , x149 , x150 , x151 , x152 , x153 , x154 , x155 , x156 , x157 , x158 , x159 , x160 , x161 , x162 , x163 , x164 , x165 , x166 , x167 , x168 , x169 , x170 , x171 , x172 , x173 , x174 , x175 , x176 , x177 , x178 , x179 , x180 , x181 , x182 , x183 , x184 , x185 , x186 , x187 , x188 , x189 , x190 , x191 , x192 , x193 , x194 , x195 , x196 , x197 , x198 , x199 , x200 , x201 , x202 , x203 , x204 , x205 , x206 , x207 , x208 , x209 , x210 , x211 , x212 , x213 , x214 , x215 , x216 , x217 , x218 , x219 , x220 , x221 , x222 , x223 , x224 , x225 , x226 , x227 , x228 , x229 , x230 , x231 , x232 , x233 , x234 , x235 , x236 , x237 , x238 , x239 , x240 , x241 , x242 , x243 , x244 , x245 , x246 , x247 , x248 , x249 , x250 , x251 , x252 , x253 , x254 , x255 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 , y128 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 , x147 , x148 , x149 , x150 , x151 , x152 , x153 , x154 , x155 , x156 , x157 , x158 , x159 , x160 , x161 , x162 , x163 , x164 , x165 , x166 , x167 , x168 , x169 , x170 , x171 , x172 , x173 , x174 , x175 , x176 , x177 , x178 , x179 , x180 , x181 , x182 , x183 , x184 , x185 , x186 , x187 , x188 , x189 , x190 , x191 , x192 , x193 , x194 , x195 , x196 , x197 , x198 , x199 , x200 , x201 , x202 , x203 , x204 , x205 , x206 , x207 , x208 , x209 , x210 , x211 , x212 , x213 , x214 , x215 , x216 , x217 , x218 , x219 , x220 , x221 , x222 , x223 , x224 , x225 , x226 , x227 , x228 , x229 , x230 , x231 , x232 , x233 , x234 , x235 , x236 , x237 , x238 , x239 , x240 , x241 , x242 , x243 , x244 , x245 , x246 , x247 , x248 , x249 , x250 , x251 , x252 , x253 , x254 , x255 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 , y128 ;
  wire n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , n3931 , n3932 , n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , n3940 , n3941 , n3942 , n3943 , n3944 , n3945 , n3946 , n3947 , n3948 , n3949 , n3950 , n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , n3970 , n3971 , n3972 , n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , n3980 , n3981 , n3982 , n3983 , n3984 , n3985 , n3986 , n3987 , n3988 , n3989 , n3990 , n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , n4000 , n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , n4009 , n4010 , n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , n4019 , n4020 , n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , n4029 , n4030 , n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , n4039 , n4040 , n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4049 , n4050 , n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , n4059 , n4060 , n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , n4070 , n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , n4079 , n4080 , n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , n4089 , n4090 , n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , n4097 , n4098 , n4099 , n4100 , n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , n4109 , n4110 , n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , n4119 , n4120 , n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , n4129 , n4130 , n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , n4139 , n4140 , n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , n4150 , n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , n4159 , n4160 , n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , n4169 , n4170 , n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , n4179 , n4180 , n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , n4189 , n4190 , n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , n4197 , n4198 , n4199 , n4200 , n4201 , n4202 , n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , n4209 , n4210 , n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , n4217 , n4218 , n4219 , n4220 , n4221 , n4222 , n4223 , n4224 , n4225 , n4226 , n4227 , n4228 , n4229 , n4230 , n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , n4237 , n4238 , n4239 , n4240 , n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , n4247 , n4248 , n4249 , n4250 , n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , n4259 , n4260 , n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , n4269 , n4270 , n4271 , n4272 , n4273 , n4274 , n4275 , n4276 , n4277 , n4278 , n4279 , n4280 , n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , n4289 , n4290 , n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , n4299 , n4300 , n4301 , n4302 , n4303 , n4304 , n4305 , n4306 , n4307 , n4308 , n4309 , n4310 , n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , n4319 , n4320 , n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , n4329 , n4330 , n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , n4340 , n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , n4349 , n4350 , n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , n4360 , n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , n4370 , n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , n4380 , n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , n4390 , n4391 , n4392 , n4393 , n4394 , n4395 , n4396 , n4397 , n4398 , n4399 , n4400 , n4401 , n4402 , n4403 , n4404 , n4405 , n4406 , n4407 , n4408 , n4409 , n4410 , n4411 , n4412 , n4413 , n4414 , n4415 , n4416 , n4417 , n4418 , n4419 , n4420 , n4421 , n4422 , n4423 , n4424 , n4425 , n4426 , n4427 , n4428 , n4429 , n4430 , n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , n4437 , n4438 , n4439 , n4440 , n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , n4449 , n4450 , n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , n4459 , n4460 , n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , n4469 , n4470 , n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , n4479 , n4480 , n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , n4487 , n4488 , n4489 , n4490 , n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , n4497 , n4498 , n4499 , n4500 , n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , n4509 , n4510 , n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , n4519 , n4520 , n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , n4529 , n4530 , n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , n4537 , n4538 , n4539 , n4540 , n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , n4547 , n4548 , n4549 , n4550 , n4551 , n4552 , n4553 , n4554 , n4555 , n4556 , n4557 , n4558 , n4559 , n4560 , n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , n4567 , n4568 , n4569 , n4570 , n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , n4579 , n4580 , n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , n4589 , n4590 , n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , n4597 , n4598 , n4599 , n4600 , n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , n4607 , n4608 , n4609 , n4610 , n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , n4617 , n4618 , n4619 , n4620 , n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , n4627 , n4628 , n4629 , n4630 , n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , n4637 , n4638 , n4639 , n4640 , n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , n4647 , n4648 , n4649 , n4650 , n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , n4657 , n4658 , n4659 , n4660 , n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , n4669 , n4670 , n4671 , n4672 , n4673 , n4674 , n4675 , n4676 , n4677 , n4678 , n4679 , n4680 , n4681 , n4682 , n4683 , n4684 , n4685 , n4686 , n4687 , n4688 , n4689 , n4690 , n4691 , n4692 , n4693 , n4694 , n4695 , n4696 , n4697 , n4698 , n4699 , n4700 , n4701 , n4702 , n4703 , n4704 , n4705 , n4706 , n4707 , n4708 , n4709 , n4710 , n4711 , n4712 , n4713 , n4714 , n4715 , n4716 , n4717 , n4718 , n4719 , n4720 , n4721 , n4722 , n4723 , n4724 , n4725 , n4726 , n4727 , n4728 , n4729 , n4730 , n4731 , n4732 , n4733 , n4734 , n4735 , n4736 , n4737 , n4738 , n4739 , n4740 , n4741 , n4742 , n4743 , n4744 , n4745 , n4746 , n4747 , n4748 , n4749 , n4750 , n4751 , n4752 , n4753 , n4754 , n4755 , n4756 , n4757 , n4758 , n4759 , n4760 , n4761 , n4762 , n4763 , n4764 , n4765 , n4766 , n4767 , n4768 , n4769 , n4770 , n4771 , n4772 , n4773 , n4774 , n4775 , n4776 , n4777 , n4778 , n4779 , n4780 , n4781 , n4782 , n4783 , n4784 , n4785 , n4786 , n4787 , n4788 , n4789 , n4790 , n4791 , n4792 , n4793 , n4794 , n4795 , n4796 , n4797 , n4798 , n4799 , n4800 , n4801 , n4802 , n4803 , n4804 , n4805 , n4806 , n4807 , n4808 , n4809 , n4810 , n4811 , n4812 , n4813 , n4814 , n4815 , n4816 , n4817 , n4818 , n4819 , n4820 , n4821 , n4822 , n4823 , n4824 , n4825 , n4826 , n4827 , n4828 , n4829 , n4830 , n4831 , n4832 , n4833 , n4834 , n4835 , n4836 , n4837 , n4838 , n4839 , n4840 , n4841 , n4842 , n4843 , n4844 , n4845 , n4846 , n4847 , n4848 , n4849 , n4850 , n4851 , n4852 , n4853 , n4854 , n4855 , n4856 , n4857 , n4858 , n4859 , n4860 , n4861 , n4862 , n4863 , n4864 , n4865 , n4866 , n4867 , n4868 , n4869 , n4870 , n4871 , n4872 , n4873 , n4874 , n4875 , n4876 , n4877 , n4878 , n4879 , n4880 , n4881 , n4882 , n4883 , n4884 , n4885 , n4886 , n4887 , n4888 , n4889 , n4890 , n4891 , n4892 , n4893 , n4894 , n4895 , n4896 , n4897 , n4898 , n4899 , n4900 , n4901 , n4902 , n4903 , n4904 , n4905 , n4906 , n4907 , n4908 , n4909 , n4910 , n4911 , n4912 , n4913 , n4914 , n4915 , n4916 , n4917 , n4918 , n4919 , n4920 , n4921 , n4922 , n4923 , n4924 , n4925 , n4926 , n4927 , n4928 , n4929 , n4930 , n4931 , n4932 , n4933 , n4934 , n4935 , n4936 , n4937 , n4938 , n4939 , n4940 , n4941 , n4942 , n4943 , n4944 , n4945 , n4946 , n4947 , n4948 , n4949 , n4950 , n4951 , n4952 , n4953 , n4954 , n4955 , n4956 , n4957 , n4958 , n4959 , n4960 , n4961 , n4962 , n4963 , n4964 , n4965 , n4966 , n4967 , n4968 , n4969 , n4970 , n4971 , n4972 , n4973 , n4974 , n4975 , n4976 , n4977 , n4978 , n4979 , n4980 , n4981 , n4982 , n4983 , n4984 , n4985 , n4986 , n4987 , n4988 , n4989 , n4990 , n4991 , n4992 , n4993 , n4994 , n4995 , n4996 , n4997 , n4998 , n4999 , n5000 , n5001 , n5002 , n5003 , n5004 , n5005 , n5006 , n5007 , n5008 , n5009 , n5010 , n5011 , n5012 , n5013 , n5014 , n5015 , n5016 , n5017 , n5018 , n5019 , n5020 , n5021 , n5022 , n5023 , n5024 , n5025 , n5026 , n5027 , n5028 , n5029 , n5030 , n5031 , n5032 , n5033 , n5034 , n5035 , n5036 , n5037 , n5038 , n5039 , n5040 , n5041 , n5042 , n5043 , n5044 , n5045 , n5046 , n5047 , n5048 , n5049 , n5050 , n5051 , n5052 , n5053 , n5054 , n5055 , n5056 , n5057 , n5058 , n5059 , n5060 , n5061 , n5062 , n5063 , n5064 , n5065 , n5066 , n5067 , n5068 , n5069 , n5070 , n5071 , n5072 , n5073 , n5074 , n5075 , n5076 , n5077 , n5078 , n5079 , n5080 , n5081 , n5082 , n5083 , n5084 , n5085 , n5086 , n5087 , n5088 , n5089 , n5090 , n5091 , n5092 , n5093 , n5094 , n5095 , n5096 , n5097 , n5098 , n5099 , n5100 , n5101 , n5102 , n5103 , n5104 , n5105 , n5106 , n5107 , n5108 , n5109 , n5110 , n5111 , n5112 , n5113 , n5114 , n5115 , n5116 , n5117 , n5118 , n5119 , n5120 , n5121 , n5122 , n5123 , n5124 , n5125 , n5126 , n5127 , n5128 , n5129 , n5130 , n5131 , n5132 , n5133 , n5134 , n5135 , n5136 , n5137 , n5138 , n5139 , n5140 , n5141 , n5142 , n5143 , n5144 , n5145 , n5146 , n5147 , n5148 , n5149 , n5150 , n5151 , n5152 , n5153 , n5154 , n5155 , n5156 , n5157 , n5158 , n5159 , n5160 , n5161 , n5162 , n5163 , n5164 , n5165 , n5166 , n5167 , n5168 , n5169 , n5170 , n5171 , n5172 , n5173 , n5174 , n5175 , n5176 , n5177 , n5178 , n5179 , n5180 , n5181 , n5182 , n5183 , n5184 , n5185 , n5186 , n5187 , n5188 , n5189 , n5190 , n5191 , n5192 , n5193 , n5194 , n5195 , n5196 , n5197 , n5198 , n5199 , n5200 , n5201 , n5202 , n5203 , n5204 , n5205 , n5206 , n5207 , n5208 , n5209 , n5210 , n5211 , n5212 , n5213 , n5214 , n5215 , n5216 , n5217 , n5218 , n5219 , n5220 , n5221 , n5222 , n5223 , n5224 , n5225 , n5226 , n5227 , n5228 , n5229 , n5230 , n5231 , n5232 , n5233 , n5234 , n5235 , n5236 , n5237 , n5238 , n5239 , n5240 , n5241 , n5242 , n5243 , n5244 , n5245 , n5246 , n5247 , n5248 , n5249 , n5250 , n5251 , n5252 , n5253 , n5254 , n5255 , n5256 , n5257 , n5258 , n5259 , n5260 , n5261 , n5262 , n5263 , n5264 , n5265 , n5266 , n5267 , n5268 , n5269 , n5270 , n5271 , n5272 , n5273 , n5274 , n5275 , n5276 , n5277 , n5278 , n5279 , n5280 , n5281 , n5282 , n5283 , n5284 , n5285 , n5286 , n5287 , n5288 , n5289 , n5290 , n5291 , n5292 , n5293 , n5294 , n5295 , n5296 , n5297 , n5298 , n5299 , n5300 , n5301 , n5302 , n5303 , n5304 , n5305 , n5306 , n5307 , n5308 , n5309 , n5310 , n5311 , n5312 , n5313 , n5314 , n5315 , n5316 , n5317 , n5318 , n5319 , n5320 , n5321 , n5322 ;
  assign n257 = ~x0 & x255 ;
  assign n258 = x128 & ~n257 ;
  assign n259 = x1 & ~x129 ;
  assign n260 = x2 | n259 ;
  assign n261 = x130 | x131 ;
  assign n262 = n260 & ~n261 ;
  assign n263 = ~x5 & x132 ;
  assign n264 = x133 | x134 ;
  assign n265 = n263 | n264 ;
  assign n266 = x3 & ~x131 ;
  assign n267 = x4 | x5 ;
  assign n268 = n266 | n267 ;
  assign n269 = ~n265 & n268 ;
  assign n270 = ( n262 & ~n265 ) | ( n262 & n269 ) | ( ~n265 & n269 ) ;
  assign n271 = ~x8 & x135 ;
  assign n272 = x136 | x137 ;
  assign n273 = n271 | n272 ;
  assign n274 = x6 & ~x134 ;
  assign n275 = x7 | x8 ;
  assign n276 = n274 | n275 ;
  assign n277 = ~n273 & n276 ;
  assign n278 = x9 & ~x137 ;
  assign n279 = x10 | x11 ;
  assign n280 = n278 | n279 ;
  assign n281 = n277 | n280 ;
  assign n282 = n273 & ~n280 ;
  assign n283 = ( n270 & n281 ) | ( n270 & ~n282 ) | ( n281 & ~n282 ) ;
  assign n284 = ~x14 & x141 ;
  assign n285 = x142 | x143 ;
  assign n286 = n284 | n285 ;
  assign n287 = ~x11 & x138 ;
  assign n288 = x139 | x140 ;
  assign n289 = n287 | n288 ;
  assign n290 = x12 & ~x140 ;
  assign n291 = x13 | x14 ;
  assign n292 = n290 | n291 ;
  assign n293 = n289 & ~n292 ;
  assign n294 = n286 | n293 ;
  assign n295 = x15 & ~x143 ;
  assign n296 = x16 | x17 ;
  assign n297 = n295 | n296 ;
  assign n298 = n294 & ~n297 ;
  assign n299 = ~n286 & n292 ;
  assign n300 = n297 | n299 ;
  assign n301 = ( n283 & ~n298 ) | ( n283 & n300 ) | ( ~n298 & n300 ) ;
  assign n302 = ~x23 & x150 ;
  assign n303 = x151 | x152 ;
  assign n304 = n302 | n303 ;
  assign n305 = ~x20 & x147 ;
  assign n306 = x148 | x149 ;
  assign n307 = n305 | n306 ;
  assign n308 = ~x17 & x144 ;
  assign n309 = x145 | x146 ;
  assign n310 = n308 | n309 ;
  assign n311 = x18 & ~x146 ;
  assign n312 = x19 | x20 ;
  assign n313 = n311 | n312 ;
  assign n314 = n310 & ~n313 ;
  assign n315 = n307 | n314 ;
  assign n316 = x21 & ~x149 ;
  assign n317 = x22 | x23 ;
  assign n318 = n316 | n317 ;
  assign n319 = n315 & ~n318 ;
  assign n320 = n304 | n319 ;
  assign n321 = ~n307 & n313 ;
  assign n322 = n318 | n321 ;
  assign n323 = ~n304 & n322 ;
  assign n324 = ( n301 & ~n320 ) | ( n301 & n323 ) | ( ~n320 & n323 ) ;
  assign n325 = ~x32 & x159 ;
  assign n326 = x160 | x161 ;
  assign n327 = n325 | n326 ;
  assign n328 = ~x29 & x156 ;
  assign n329 = x157 | x158 ;
  assign n330 = n328 | n329 ;
  assign n331 = ~x26 & x153 ;
  assign n332 = x154 | x155 ;
  assign n333 = n331 | n332 ;
  assign n334 = x24 & ~x152 ;
  assign n335 = x25 | x26 ;
  assign n336 = n334 | n335 ;
  assign n337 = ~n333 & n336 ;
  assign n338 = x27 & ~x155 ;
  assign n339 = x28 | x29 ;
  assign n340 = n338 | n339 ;
  assign n341 = n337 | n340 ;
  assign n342 = ~n330 & n341 ;
  assign n343 = x30 & ~x158 ;
  assign n344 = x31 | x32 ;
  assign n345 = n343 | n344 ;
  assign n346 = n342 | n345 ;
  assign n347 = ~n327 & n346 ;
  assign n348 = n333 & ~n340 ;
  assign n349 = n330 & ~n345 ;
  assign n350 = ( ~n345 & n348 ) | ( ~n345 & n349 ) | ( n348 & n349 ) ;
  assign n351 = n327 | n350 ;
  assign n352 = ( n324 & n347 ) | ( n324 & ~n351 ) | ( n347 & ~n351 ) ;
  assign n353 = ~x41 & x168 ;
  assign n354 = x169 | x170 ;
  assign n355 = n353 | n354 ;
  assign n356 = ~x38 & x165 ;
  assign n357 = x166 | x167 ;
  assign n358 = n356 | n357 ;
  assign n359 = ~x35 & x162 ;
  assign n360 = x163 | x164 ;
  assign n361 = n359 | n360 ;
  assign n362 = x33 & ~x161 ;
  assign n363 = x34 | x35 ;
  assign n364 = n362 | n363 ;
  assign n365 = ~n361 & n364 ;
  assign n366 = x36 & ~x164 ;
  assign n367 = x37 | x38 ;
  assign n368 = n366 | n367 ;
  assign n369 = n365 | n368 ;
  assign n370 = ~n358 & n369 ;
  assign n371 = x39 & ~x167 ;
  assign n372 = x40 | x41 ;
  assign n373 = n371 | n372 ;
  assign n374 = n370 | n373 ;
  assign n375 = ~n355 & n374 ;
  assign n376 = x42 & ~x170 ;
  assign n377 = x43 | x44 ;
  assign n378 = n376 | n377 ;
  assign n379 = n375 | n378 ;
  assign n380 = n361 & ~n368 ;
  assign n381 = n358 & ~n373 ;
  assign n382 = ( ~n373 & n380 ) | ( ~n373 & n381 ) | ( n380 & n381 ) ;
  assign n383 = n355 | n382 ;
  assign n384 = ~n378 & n383 ;
  assign n385 = ( n352 & n379 ) | ( n352 & ~n384 ) | ( n379 & ~n384 ) ;
  assign n386 = x54 & ~x182 ;
  assign n387 = x55 | x56 ;
  assign n388 = n386 | n387 ;
  assign n389 = ~x53 & x180 ;
  assign n390 = x181 | x182 ;
  assign n391 = n389 | n390 ;
  assign n392 = x51 & ~x179 ;
  assign n393 = x52 | x53 ;
  assign n394 = n392 | n393 ;
  assign n395 = ~x50 & x177 ;
  assign n396 = x178 | x179 ;
  assign n397 = n395 | n396 ;
  assign n398 = x48 & ~x176 ;
  assign n399 = x49 | x50 ;
  assign n400 = n398 | n399 ;
  assign n401 = ~x47 & x174 ;
  assign n402 = x175 | x176 ;
  assign n403 = n401 | n402 ;
  assign n404 = x45 & ~x173 ;
  assign n405 = x46 | x47 ;
  assign n406 = n404 | n405 ;
  assign n407 = ~n403 & n406 ;
  assign n408 = n400 | n407 ;
  assign n409 = ~n397 & n408 ;
  assign n410 = n394 | n409 ;
  assign n411 = ~n391 & n410 ;
  assign n412 = n388 | n411 ;
  assign n413 = ~x44 & x171 ;
  assign n414 = x172 | x173 ;
  assign n415 = n413 | n414 ;
  assign n416 = ~n406 & n415 ;
  assign n417 = ~n400 & n403 ;
  assign n418 = ( ~n400 & n416 ) | ( ~n400 & n417 ) | ( n416 & n417 ) ;
  assign n419 = n397 | n418 ;
  assign n420 = ~n394 & n419 ;
  assign n421 = ~n388 & n391 ;
  assign n422 = ( ~n388 & n420 ) | ( ~n388 & n421 ) | ( n420 & n421 ) ;
  assign n423 = ( n385 & n412 ) | ( n385 & ~n422 ) | ( n412 & ~n422 ) ;
  assign n424 = ~x68 & x195 ;
  assign n425 = x196 | x197 ;
  assign n426 = n424 | n425 ;
  assign n427 = ~x62 & x189 ;
  assign n428 = x190 | x191 ;
  assign n429 = n427 | n428 ;
  assign n430 = ~x59 & x186 ;
  assign n431 = x187 | x188 ;
  assign n432 = n430 | n431 ;
  assign n433 = ~x56 & x183 ;
  assign n434 = x184 | x185 ;
  assign n435 = n433 | n434 ;
  assign n436 = x57 & ~x185 ;
  assign n437 = x58 | x59 ;
  assign n438 = n436 | n437 ;
  assign n439 = n435 & ~n438 ;
  assign n440 = n432 | n439 ;
  assign n441 = x60 & ~x188 ;
  assign n442 = x61 | x62 ;
  assign n443 = n441 | n442 ;
  assign n444 = n440 & ~n443 ;
  assign n445 = n429 | n444 ;
  assign n446 = x63 & ~x191 ;
  assign n447 = x64 | x65 ;
  assign n448 = n446 | n447 ;
  assign n449 = n445 & ~n448 ;
  assign n450 = x66 & ~x194 ;
  assign n451 = x67 | x68 ;
  assign n452 = n450 | n451 ;
  assign n453 = ~x65 & x192 ;
  assign n454 = x193 | x194 ;
  assign n455 = n453 | n454 ;
  assign n456 = ~n452 & n455 ;
  assign n457 = ( n449 & ~n452 ) | ( n449 & n456 ) | ( ~n452 & n456 ) ;
  assign n458 = n426 | n457 ;
  assign n459 = ~n432 & n438 ;
  assign n460 = n443 | n459 ;
  assign n461 = ~n429 & n460 ;
  assign n462 = n448 | n461 ;
  assign n463 = ~n455 & n462 ;
  assign n464 = n452 | n463 ;
  assign n465 = ~n426 & n464 ;
  assign n466 = ( n423 & ~n458 ) | ( n423 & n465 ) | ( ~n458 & n465 ) ;
  assign n467 = ~x83 & x210 ;
  assign n468 = x211 | x212 ;
  assign n469 = n467 | n468 ;
  assign n470 = x81 & ~x209 ;
  assign n471 = x82 | x83 ;
  assign n472 = n470 | n471 ;
  assign n473 = x78 & ~x206 ;
  assign n474 = x79 | x80 ;
  assign n475 = n473 | n474 ;
  assign n476 = ~x77 & x204 ;
  assign n477 = x205 | x206 ;
  assign n478 = n476 | n477 ;
  assign n479 = x75 & ~x203 ;
  assign n480 = x76 | x77 ;
  assign n481 = n479 | n480 ;
  assign n482 = ~x71 & x198 ;
  assign n483 = x199 | x200 ;
  assign n484 = n482 | n483 ;
  assign n485 = x72 & ~x200 ;
  assign n486 = x73 | x74 ;
  assign n487 = n485 | n486 ;
  assign n488 = n484 & ~n487 ;
  assign n489 = ~x74 & x201 ;
  assign n490 = x202 | x203 ;
  assign n491 = n489 | n490 ;
  assign n492 = ~n481 & n491 ;
  assign n493 = ( ~n481 & n488 ) | ( ~n481 & n492 ) | ( n488 & n492 ) ;
  assign n494 = n478 | n493 ;
  assign n495 = ~n475 & n494 ;
  assign n496 = ~x80 & x207 ;
  assign n497 = x208 | x209 ;
  assign n498 = n496 | n497 ;
  assign n499 = ~n472 & n498 ;
  assign n500 = ( ~n472 & n495 ) | ( ~n472 & n499 ) | ( n495 & n499 ) ;
  assign n501 = n469 | n500 ;
  assign n502 = x69 & ~x197 ;
  assign n503 = x70 | x71 ;
  assign n504 = n502 | n503 ;
  assign n505 = ~n484 & n504 ;
  assign n506 = n487 | n505 ;
  assign n507 = ~n491 & n506 ;
  assign n508 = n481 | n507 ;
  assign n509 = ~n478 & n508 ;
  assign n510 = n475 | n509 ;
  assign n511 = ~n498 & n510 ;
  assign n512 = ~n469 & n472 ;
  assign n513 = ( ~n469 & n511 ) | ( ~n469 & n512 ) | ( n511 & n512 ) ;
  assign n514 = ( n466 & ~n501 ) | ( n466 & n513 ) | ( ~n501 & n513 ) ;
  assign n515 = x99 & ~x227 ;
  assign n516 = x100 | x101 ;
  assign n517 = n515 | n516 ;
  assign n518 = ~x98 & x225 ;
  assign n519 = x226 | x227 ;
  assign n520 = n518 | n519 ;
  assign n521 = ~x95 & x222 ;
  assign n522 = x223 | x224 ;
  assign n523 = n521 | n522 ;
  assign n524 = ~x92 & x219 ;
  assign n525 = x220 | x221 ;
  assign n526 = n524 | n525 ;
  assign n527 = ~x89 & x216 ;
  assign n528 = x217 | x218 ;
  assign n529 = n527 | n528 ;
  assign n530 = ~x86 & x213 ;
  assign n531 = x214 | x215 ;
  assign n532 = n530 | n531 ;
  assign n533 = x84 & ~x212 ;
  assign n534 = x85 | x86 ;
  assign n535 = n533 | n534 ;
  assign n536 = ~n532 & n535 ;
  assign n537 = x87 & ~x215 ;
  assign n538 = x88 | x89 ;
  assign n539 = n537 | n538 ;
  assign n540 = n536 | n539 ;
  assign n541 = ~n529 & n540 ;
  assign n542 = x90 & ~x218 ;
  assign n543 = x91 | x92 ;
  assign n544 = n542 | n543 ;
  assign n545 = n541 | n544 ;
  assign n546 = ~n526 & n545 ;
  assign n547 = x93 & ~x221 ;
  assign n548 = x94 | x95 ;
  assign n549 = n547 | n548 ;
  assign n550 = n546 | n549 ;
  assign n551 = ~n523 & n550 ;
  assign n552 = x96 & ~x224 ;
  assign n553 = x97 | x98 ;
  assign n554 = n552 | n553 ;
  assign n555 = ~n520 & n554 ;
  assign n556 = ( ~n520 & n551 ) | ( ~n520 & n555 ) | ( n551 & n555 ) ;
  assign n557 = n517 | n556 ;
  assign n558 = n532 & ~n539 ;
  assign n559 = n529 & ~n544 ;
  assign n560 = ( ~n544 & n558 ) | ( ~n544 & n559 ) | ( n558 & n559 ) ;
  assign n561 = n526 | n560 ;
  assign n562 = ~n549 & n561 ;
  assign n563 = n523 & ~n554 ;
  assign n564 = ( ~n554 & n562 ) | ( ~n554 & n563 ) | ( n562 & n563 ) ;
  assign n565 = n520 | n564 ;
  assign n566 = ~n517 & n565 ;
  assign n567 = ( n514 & n557 ) | ( n514 & ~n566 ) | ( n557 & ~n566 ) ;
  assign n568 = x117 & ~x245 ;
  assign n569 = x118 | x119 ;
  assign n570 = n568 | n569 ;
  assign n571 = ~x116 & x243 ;
  assign n572 = x244 | x245 ;
  assign n573 = n571 | n572 ;
  assign n574 = ~x113 & x240 ;
  assign n575 = x241 | x242 ;
  assign n576 = n574 | n575 ;
  assign n577 = x111 & ~x239 ;
  assign n578 = x112 | x113 ;
  assign n579 = n577 | n578 ;
  assign n580 = ~x110 & x237 ;
  assign n581 = x238 | x239 ;
  assign n582 = n580 | n581 ;
  assign n583 = x108 & ~x236 ;
  assign n584 = x109 | x110 ;
  assign n585 = n583 | n584 ;
  assign n586 = ~x107 & x234 ;
  assign n587 = x235 | x236 ;
  assign n588 = n586 | n587 ;
  assign n589 = x105 & ~x233 ;
  assign n590 = x106 | x107 ;
  assign n591 = n589 | n590 ;
  assign n592 = ~x104 & x231 ;
  assign n593 = x232 | x233 ;
  assign n594 = n592 | n593 ;
  assign n595 = x102 & ~x230 ;
  assign n596 = x103 | x104 ;
  assign n597 = n595 | n596 ;
  assign n598 = ~n594 & n597 ;
  assign n599 = n591 | n598 ;
  assign n600 = ~n588 & n599 ;
  assign n601 = n585 | n600 ;
  assign n602 = ~n582 & n601 ;
  assign n603 = n579 | n602 ;
  assign n604 = ~n576 & n603 ;
  assign n605 = x114 & ~x242 ;
  assign n606 = x115 | x116 ;
  assign n607 = n605 | n606 ;
  assign n608 = ~n573 & n607 ;
  assign n609 = ( ~n573 & n604 ) | ( ~n573 & n608 ) | ( n604 & n608 ) ;
  assign n610 = n570 | n609 ;
  assign n611 = ~x101 & x228 ;
  assign n612 = x229 | x230 ;
  assign n613 = n611 | n612 ;
  assign n614 = ~n597 & n613 ;
  assign n615 = ~n591 & n594 ;
  assign n616 = ( ~n591 & n614 ) | ( ~n591 & n615 ) | ( n614 & n615 ) ;
  assign n617 = n588 | n616 ;
  assign n618 = ~n585 & n617 ;
  assign n619 = ~n579 & n582 ;
  assign n620 = ( ~n579 & n618 ) | ( ~n579 & n619 ) | ( n618 & n619 ) ;
  assign n621 = n576 | n620 ;
  assign n622 = ~n607 & n621 ;
  assign n623 = ~n570 & n573 ;
  assign n624 = ( ~n570 & n622 ) | ( ~n570 & n623 ) | ( n622 & n623 ) ;
  assign n625 = ( n567 & n610 ) | ( n567 & ~n624 ) | ( n610 & ~n624 ) ;
  assign n626 = ~x125 & x252 ;
  assign n627 = x253 | x254 ;
  assign n628 = n626 | n627 ;
  assign n629 = ~x122 & x249 ;
  assign n630 = x250 | x251 ;
  assign n631 = n629 | n630 ;
  assign n632 = ~x119 & x246 ;
  assign n633 = x247 | x248 ;
  assign n634 = n632 | n633 ;
  assign n635 = x120 & ~x248 ;
  assign n636 = x121 | x122 ;
  assign n637 = n635 | n636 ;
  assign n638 = n634 & ~n637 ;
  assign n639 = n631 | n638 ;
  assign n640 = x123 & ~x251 ;
  assign n641 = x124 | x125 ;
  assign n642 = n640 | n641 ;
  assign n643 = n639 & ~n642 ;
  assign n644 = n628 | n643 ;
  assign n645 = x126 & ~x254 ;
  assign n646 = x127 | n645 ;
  assign n647 = x0 | n646 ;
  assign n648 = n644 & ~n647 ;
  assign n649 = ~n631 & n637 ;
  assign n650 = n642 | n649 ;
  assign n651 = ~n628 & n650 ;
  assign n652 = n647 | n651 ;
  assign n653 = ( n625 & ~n648 ) | ( n625 & n652 ) | ( ~n648 & n652 ) ;
  assign n654 = n258 & n653 ;
  assign n655 = ~x1 & x128 ;
  assign n656 = x129 & ~n655 ;
  assign n657 = x2 & ~x130 ;
  assign n658 = x3 | n657 ;
  assign n659 = x131 | x132 ;
  assign n660 = n658 & ~n659 ;
  assign n661 = ~x6 & x133 ;
  assign n662 = x134 | x135 ;
  assign n663 = n661 | n662 ;
  assign n664 = x4 & ~x132 ;
  assign n665 = x5 | x6 ;
  assign n666 = n664 | n665 ;
  assign n667 = ~n663 & n666 ;
  assign n668 = ( n660 & ~n663 ) | ( n660 & n667 ) | ( ~n663 & n667 ) ;
  assign n669 = ~x9 & x136 ;
  assign n670 = x137 | x138 ;
  assign n671 = n669 | n670 ;
  assign n672 = x7 & ~x135 ;
  assign n673 = x8 | x9 ;
  assign n674 = n672 | n673 ;
  assign n675 = ~n671 & n674 ;
  assign n676 = x10 & ~x138 ;
  assign n677 = x11 | x12 ;
  assign n678 = n676 | n677 ;
  assign n679 = n675 | n678 ;
  assign n680 = n671 & ~n678 ;
  assign n681 = ( n668 & n679 ) | ( n668 & ~n680 ) | ( n679 & ~n680 ) ;
  assign n682 = ~x15 & x142 ;
  assign n683 = x143 | x144 ;
  assign n684 = n682 | n683 ;
  assign n685 = ~x12 & x139 ;
  assign n686 = x140 | x141 ;
  assign n687 = n685 | n686 ;
  assign n688 = x13 & ~x141 ;
  assign n689 = x14 | x15 ;
  assign n690 = n688 | n689 ;
  assign n691 = n687 & ~n690 ;
  assign n692 = n684 | n691 ;
  assign n693 = x16 & ~x144 ;
  assign n694 = x17 | x18 ;
  assign n695 = n693 | n694 ;
  assign n696 = n692 & ~n695 ;
  assign n697 = ~n684 & n690 ;
  assign n698 = n695 | n697 ;
  assign n699 = ( n681 & ~n696 ) | ( n681 & n698 ) | ( ~n696 & n698 ) ;
  assign n700 = ~x24 & x151 ;
  assign n701 = x152 | x153 ;
  assign n702 = n700 | n701 ;
  assign n703 = ~x21 & x148 ;
  assign n704 = x149 | x150 ;
  assign n705 = n703 | n704 ;
  assign n706 = ~x18 & x145 ;
  assign n707 = x146 | x147 ;
  assign n708 = n706 | n707 ;
  assign n709 = x19 & ~x147 ;
  assign n710 = x20 | x21 ;
  assign n711 = n709 | n710 ;
  assign n712 = n708 & ~n711 ;
  assign n713 = n705 | n712 ;
  assign n714 = x22 & ~x150 ;
  assign n715 = x23 | x24 ;
  assign n716 = n714 | n715 ;
  assign n717 = n713 & ~n716 ;
  assign n718 = n702 | n717 ;
  assign n719 = ~n705 & n711 ;
  assign n720 = n716 | n719 ;
  assign n721 = ~n702 & n720 ;
  assign n722 = ( n699 & ~n718 ) | ( n699 & n721 ) | ( ~n718 & n721 ) ;
  assign n723 = ~x33 & x160 ;
  assign n724 = x161 | x162 ;
  assign n725 = n723 | n724 ;
  assign n726 = ~x30 & x157 ;
  assign n727 = x158 | x159 ;
  assign n728 = n726 | n727 ;
  assign n729 = ~x27 & x154 ;
  assign n730 = x155 | x156 ;
  assign n731 = n729 | n730 ;
  assign n732 = x25 & ~x153 ;
  assign n733 = x26 | x27 ;
  assign n734 = n732 | n733 ;
  assign n735 = ~n731 & n734 ;
  assign n736 = x28 & ~x156 ;
  assign n737 = x29 | x30 ;
  assign n738 = n736 | n737 ;
  assign n739 = n735 | n738 ;
  assign n740 = ~n728 & n739 ;
  assign n741 = x31 & ~x159 ;
  assign n742 = x32 | x33 ;
  assign n743 = n741 | n742 ;
  assign n744 = n740 | n743 ;
  assign n745 = ~n725 & n744 ;
  assign n746 = n731 & ~n738 ;
  assign n747 = n728 & ~n743 ;
  assign n748 = ( ~n743 & n746 ) | ( ~n743 & n747 ) | ( n746 & n747 ) ;
  assign n749 = n725 | n748 ;
  assign n750 = ( n722 & n745 ) | ( n722 & ~n749 ) | ( n745 & ~n749 ) ;
  assign n751 = ~x42 & x169 ;
  assign n752 = x170 | x171 ;
  assign n753 = n751 | n752 ;
  assign n754 = ~x39 & x166 ;
  assign n755 = x167 | x168 ;
  assign n756 = n754 | n755 ;
  assign n757 = ~x36 & x163 ;
  assign n758 = x164 | x165 ;
  assign n759 = n757 | n758 ;
  assign n760 = x34 & ~x162 ;
  assign n761 = x35 | x36 ;
  assign n762 = n760 | n761 ;
  assign n763 = ~n759 & n762 ;
  assign n764 = x37 & ~x165 ;
  assign n765 = x38 | x39 ;
  assign n766 = n764 | n765 ;
  assign n767 = n763 | n766 ;
  assign n768 = ~n756 & n767 ;
  assign n769 = x40 & ~x168 ;
  assign n770 = x41 | x42 ;
  assign n771 = n769 | n770 ;
  assign n772 = n768 | n771 ;
  assign n773 = ~n753 & n772 ;
  assign n774 = x43 & ~x171 ;
  assign n775 = x44 | x45 ;
  assign n776 = n774 | n775 ;
  assign n777 = n773 | n776 ;
  assign n778 = n759 & ~n766 ;
  assign n779 = n756 & ~n771 ;
  assign n780 = ( ~n771 & n778 ) | ( ~n771 & n779 ) | ( n778 & n779 ) ;
  assign n781 = n753 | n780 ;
  assign n782 = ~n776 & n781 ;
  assign n783 = ( n750 & n777 ) | ( n750 & ~n782 ) | ( n777 & ~n782 ) ;
  assign n784 = x55 & ~x183 ;
  assign n785 = x56 | x57 ;
  assign n786 = n784 | n785 ;
  assign n787 = ~x54 & x181 ;
  assign n788 = x182 | x183 ;
  assign n789 = n787 | n788 ;
  assign n790 = x52 & ~x180 ;
  assign n791 = x53 | x54 ;
  assign n792 = n790 | n791 ;
  assign n793 = ~x51 & x178 ;
  assign n794 = x179 | x180 ;
  assign n795 = n793 | n794 ;
  assign n796 = x49 & ~x177 ;
  assign n797 = x50 | x51 ;
  assign n798 = n796 | n797 ;
  assign n799 = ~x48 & x175 ;
  assign n800 = x176 | x177 ;
  assign n801 = n799 | n800 ;
  assign n802 = x46 & ~x174 ;
  assign n803 = x47 | x48 ;
  assign n804 = n802 | n803 ;
  assign n805 = ~n801 & n804 ;
  assign n806 = n798 | n805 ;
  assign n807 = ~n795 & n806 ;
  assign n808 = n792 | n807 ;
  assign n809 = ~n789 & n808 ;
  assign n810 = n786 | n809 ;
  assign n811 = ~x45 & x172 ;
  assign n812 = x173 | x174 ;
  assign n813 = n811 | n812 ;
  assign n814 = ~n804 & n813 ;
  assign n815 = ~n798 & n801 ;
  assign n816 = ( ~n798 & n814 ) | ( ~n798 & n815 ) | ( n814 & n815 ) ;
  assign n817 = n795 | n816 ;
  assign n818 = ~n792 & n817 ;
  assign n819 = ~n786 & n789 ;
  assign n820 = ( ~n786 & n818 ) | ( ~n786 & n819 ) | ( n818 & n819 ) ;
  assign n821 = ( n783 & n810 ) | ( n783 & ~n820 ) | ( n810 & ~n820 ) ;
  assign n822 = ~x69 & x196 ;
  assign n823 = x197 | x198 ;
  assign n824 = n822 | n823 ;
  assign n825 = ~x63 & x190 ;
  assign n826 = x191 | x192 ;
  assign n827 = n825 | n826 ;
  assign n828 = ~x60 & x187 ;
  assign n829 = x188 | x189 ;
  assign n830 = n828 | n829 ;
  assign n831 = ~x57 & x184 ;
  assign n832 = x185 | x186 ;
  assign n833 = n831 | n832 ;
  assign n834 = x58 & ~x186 ;
  assign n835 = x59 | x60 ;
  assign n836 = n834 | n835 ;
  assign n837 = n833 & ~n836 ;
  assign n838 = n830 | n837 ;
  assign n839 = x61 & ~x189 ;
  assign n840 = x62 | x63 ;
  assign n841 = n839 | n840 ;
  assign n842 = n838 & ~n841 ;
  assign n843 = n827 | n842 ;
  assign n844 = x64 & ~x192 ;
  assign n845 = x65 | x66 ;
  assign n846 = n844 | n845 ;
  assign n847 = n843 & ~n846 ;
  assign n848 = x67 & ~x195 ;
  assign n849 = x68 | x69 ;
  assign n850 = n848 | n849 ;
  assign n851 = ~x66 & x193 ;
  assign n852 = x194 | x195 ;
  assign n853 = n851 | n852 ;
  assign n854 = ~n850 & n853 ;
  assign n855 = ( n847 & ~n850 ) | ( n847 & n854 ) | ( ~n850 & n854 ) ;
  assign n856 = n824 | n855 ;
  assign n857 = ~n830 & n836 ;
  assign n858 = n841 | n857 ;
  assign n859 = ~n827 & n858 ;
  assign n860 = n846 | n859 ;
  assign n861 = ~n853 & n860 ;
  assign n862 = n850 | n861 ;
  assign n863 = ~n824 & n862 ;
  assign n864 = ( n821 & ~n856 ) | ( n821 & n863 ) | ( ~n856 & n863 ) ;
  assign n865 = ~x84 & x211 ;
  assign n866 = x212 | x213 ;
  assign n867 = n865 | n866 ;
  assign n868 = x82 & ~x210 ;
  assign n869 = x83 | x84 ;
  assign n870 = n868 | n869 ;
  assign n871 = x79 & ~x207 ;
  assign n872 = x80 | x81 ;
  assign n873 = n871 | n872 ;
  assign n874 = ~x78 & x205 ;
  assign n875 = x206 | x207 ;
  assign n876 = n874 | n875 ;
  assign n877 = x76 & ~x204 ;
  assign n878 = x77 | x78 ;
  assign n879 = n877 | n878 ;
  assign n880 = ~x72 & x199 ;
  assign n881 = x200 | x201 ;
  assign n882 = n880 | n881 ;
  assign n883 = x73 & ~x201 ;
  assign n884 = x74 | x75 ;
  assign n885 = n883 | n884 ;
  assign n886 = n882 & ~n885 ;
  assign n887 = ~x75 & x202 ;
  assign n888 = x203 | x204 ;
  assign n889 = n887 | n888 ;
  assign n890 = ~n879 & n889 ;
  assign n891 = ( ~n879 & n886 ) | ( ~n879 & n890 ) | ( n886 & n890 ) ;
  assign n892 = n876 | n891 ;
  assign n893 = ~n873 & n892 ;
  assign n894 = ~x81 & x208 ;
  assign n895 = x209 | x210 ;
  assign n896 = n894 | n895 ;
  assign n897 = ~n870 & n896 ;
  assign n898 = ( ~n870 & n893 ) | ( ~n870 & n897 ) | ( n893 & n897 ) ;
  assign n899 = n867 | n898 ;
  assign n900 = x70 & ~x198 ;
  assign n901 = x71 | x72 ;
  assign n902 = n900 | n901 ;
  assign n903 = ~n882 & n902 ;
  assign n904 = n885 | n903 ;
  assign n905 = ~n889 & n904 ;
  assign n906 = n879 | n905 ;
  assign n907 = ~n876 & n906 ;
  assign n908 = n873 | n907 ;
  assign n909 = ~n896 & n908 ;
  assign n910 = ~n867 & n870 ;
  assign n911 = ( ~n867 & n909 ) | ( ~n867 & n910 ) | ( n909 & n910 ) ;
  assign n912 = ( n864 & ~n899 ) | ( n864 & n911 ) | ( ~n899 & n911 ) ;
  assign n913 = x100 & ~x228 ;
  assign n914 = x101 | x102 ;
  assign n915 = n913 | n914 ;
  assign n916 = ~x99 & x226 ;
  assign n917 = x227 | x228 ;
  assign n918 = n916 | n917 ;
  assign n919 = ~x96 & x223 ;
  assign n920 = x224 | x225 ;
  assign n921 = n919 | n920 ;
  assign n922 = ~x93 & x220 ;
  assign n923 = x221 | x222 ;
  assign n924 = n922 | n923 ;
  assign n925 = ~x90 & x217 ;
  assign n926 = x218 | x219 ;
  assign n927 = n925 | n926 ;
  assign n928 = ~x87 & x214 ;
  assign n929 = x215 | x216 ;
  assign n930 = n928 | n929 ;
  assign n931 = x85 & ~x213 ;
  assign n932 = x86 | x87 ;
  assign n933 = n931 | n932 ;
  assign n934 = ~n930 & n933 ;
  assign n935 = x88 & ~x216 ;
  assign n936 = x89 | x90 ;
  assign n937 = n935 | n936 ;
  assign n938 = n934 | n937 ;
  assign n939 = ~n927 & n938 ;
  assign n940 = x91 & ~x219 ;
  assign n941 = x92 | x93 ;
  assign n942 = n940 | n941 ;
  assign n943 = n939 | n942 ;
  assign n944 = ~n924 & n943 ;
  assign n945 = x94 & ~x222 ;
  assign n946 = x95 | x96 ;
  assign n947 = n945 | n946 ;
  assign n948 = n944 | n947 ;
  assign n949 = ~n921 & n948 ;
  assign n950 = x97 & ~x225 ;
  assign n951 = x98 | x99 ;
  assign n952 = n950 | n951 ;
  assign n953 = ~n918 & n952 ;
  assign n954 = ( ~n918 & n949 ) | ( ~n918 & n953 ) | ( n949 & n953 ) ;
  assign n955 = n915 | n954 ;
  assign n956 = n930 & ~n937 ;
  assign n957 = n927 & ~n942 ;
  assign n958 = ( ~n942 & n956 ) | ( ~n942 & n957 ) | ( n956 & n957 ) ;
  assign n959 = n924 | n958 ;
  assign n960 = ~n947 & n959 ;
  assign n961 = n921 & ~n952 ;
  assign n962 = ( ~n952 & n960 ) | ( ~n952 & n961 ) | ( n960 & n961 ) ;
  assign n963 = n918 | n962 ;
  assign n964 = ~n915 & n963 ;
  assign n965 = ( n912 & n955 ) | ( n912 & ~n964 ) | ( n955 & ~n964 ) ;
  assign n966 = x118 & ~x246 ;
  assign n967 = x119 | x120 ;
  assign n968 = n966 | n967 ;
  assign n969 = ~x117 & x244 ;
  assign n970 = x245 | x246 ;
  assign n971 = n969 | n970 ;
  assign n972 = ~x114 & x241 ;
  assign n973 = x242 | x243 ;
  assign n974 = n972 | n973 ;
  assign n975 = x112 & ~x240 ;
  assign n976 = x113 | x114 ;
  assign n977 = n975 | n976 ;
  assign n978 = ~x111 & x238 ;
  assign n979 = x239 | x240 ;
  assign n980 = n978 | n979 ;
  assign n981 = x109 & ~x237 ;
  assign n982 = x110 | x111 ;
  assign n983 = n981 | n982 ;
  assign n984 = ~x108 & x235 ;
  assign n985 = x236 | x237 ;
  assign n986 = n984 | n985 ;
  assign n987 = x106 & ~x234 ;
  assign n988 = x107 | x108 ;
  assign n989 = n987 | n988 ;
  assign n990 = ~x105 & x232 ;
  assign n991 = x233 | x234 ;
  assign n992 = n990 | n991 ;
  assign n993 = x103 & ~x231 ;
  assign n994 = x104 | x105 ;
  assign n995 = n993 | n994 ;
  assign n996 = ~n992 & n995 ;
  assign n997 = n989 | n996 ;
  assign n998 = ~n986 & n997 ;
  assign n999 = n983 | n998 ;
  assign n1000 = ~n980 & n999 ;
  assign n1001 = n977 | n1000 ;
  assign n1002 = ~n974 & n1001 ;
  assign n1003 = x115 & ~x243 ;
  assign n1004 = x116 | x117 ;
  assign n1005 = n1003 | n1004 ;
  assign n1006 = ~n971 & n1005 ;
  assign n1007 = ( ~n971 & n1002 ) | ( ~n971 & n1006 ) | ( n1002 & n1006 ) ;
  assign n1008 = n968 | n1007 ;
  assign n1009 = ~x102 & x229 ;
  assign n1010 = x230 | x231 ;
  assign n1011 = n1009 | n1010 ;
  assign n1012 = ~n995 & n1011 ;
  assign n1013 = ~n989 & n992 ;
  assign n1014 = ( ~n989 & n1012 ) | ( ~n989 & n1013 ) | ( n1012 & n1013 ) ;
  assign n1015 = n986 | n1014 ;
  assign n1016 = ~n983 & n1015 ;
  assign n1017 = ~n977 & n980 ;
  assign n1018 = ( ~n977 & n1016 ) | ( ~n977 & n1017 ) | ( n1016 & n1017 ) ;
  assign n1019 = n974 | n1018 ;
  assign n1020 = ~n1005 & n1019 ;
  assign n1021 = ~n968 & n971 ;
  assign n1022 = ( ~n968 & n1020 ) | ( ~n968 & n1021 ) | ( n1020 & n1021 ) ;
  assign n1023 = ( n965 & n1008 ) | ( n965 & ~n1022 ) | ( n1008 & ~n1022 ) ;
  assign n1024 = ~x126 & x253 ;
  assign n1025 = x254 | x255 ;
  assign n1026 = n1024 | n1025 ;
  assign n1027 = ~x123 & x250 ;
  assign n1028 = x251 | x252 ;
  assign n1029 = n1027 | n1028 ;
  assign n1030 = ~x120 & x247 ;
  assign n1031 = x248 | x249 ;
  assign n1032 = n1030 | n1031 ;
  assign n1033 = x121 & ~x249 ;
  assign n1034 = x122 | x123 ;
  assign n1035 = n1033 | n1034 ;
  assign n1036 = n1032 & ~n1035 ;
  assign n1037 = n1029 | n1036 ;
  assign n1038 = x124 & ~x252 ;
  assign n1039 = x125 | x126 ;
  assign n1040 = n1038 | n1039 ;
  assign n1041 = n1037 & ~n1040 ;
  assign n1042 = n1026 | n1041 ;
  assign n1043 = x127 & ~x255 ;
  assign n1044 = x0 | x1 ;
  assign n1045 = n1043 | n1044 ;
  assign n1046 = n1042 & ~n1045 ;
  assign n1047 = ~n1029 & n1035 ;
  assign n1048 = n1040 | n1047 ;
  assign n1049 = ~n1026 & n1048 ;
  assign n1050 = n1045 | n1049 ;
  assign n1051 = ( n1023 & ~n1046 ) | ( n1023 & n1050 ) | ( ~n1046 & n1050 ) ;
  assign n1052 = n656 & n1051 ;
  assign n1053 = ~x2 & x129 ;
  assign n1054 = x130 & ~n1053 ;
  assign n1055 = x4 | n266 ;
  assign n1056 = x132 | x133 ;
  assign n1057 = n1055 & ~n1056 ;
  assign n1058 = ~x7 & x134 ;
  assign n1059 = x135 | x136 ;
  assign n1060 = n1058 | n1059 ;
  assign n1061 = x5 & ~x133 ;
  assign n1062 = x6 | x7 ;
  assign n1063 = n1061 | n1062 ;
  assign n1064 = ~n1060 & n1063 ;
  assign n1065 = ( n1057 & ~n1060 ) | ( n1057 & n1064 ) | ( ~n1060 & n1064 ) ;
  assign n1066 = ~x10 & x137 ;
  assign n1067 = x138 | x139 ;
  assign n1068 = n1066 | n1067 ;
  assign n1069 = x8 & ~x136 ;
  assign n1070 = x9 | x10 ;
  assign n1071 = n1069 | n1070 ;
  assign n1072 = ~n1068 & n1071 ;
  assign n1073 = x11 & ~x139 ;
  assign n1074 = x12 | x13 ;
  assign n1075 = n1073 | n1074 ;
  assign n1076 = n1072 | n1075 ;
  assign n1077 = n1068 & ~n1075 ;
  assign n1078 = ( n1065 & n1076 ) | ( n1065 & ~n1077 ) | ( n1076 & ~n1077 ) ;
  assign n1079 = ~x16 & x143 ;
  assign n1080 = x144 | x145 ;
  assign n1081 = n1079 | n1080 ;
  assign n1082 = ~x13 & x140 ;
  assign n1083 = x141 | x142 ;
  assign n1084 = n1082 | n1083 ;
  assign n1085 = x14 & ~x142 ;
  assign n1086 = x15 | x16 ;
  assign n1087 = n1085 | n1086 ;
  assign n1088 = n1084 & ~n1087 ;
  assign n1089 = n1081 | n1088 ;
  assign n1090 = x17 & ~x145 ;
  assign n1091 = x18 | x19 ;
  assign n1092 = n1090 | n1091 ;
  assign n1093 = n1089 & ~n1092 ;
  assign n1094 = ~n1081 & n1087 ;
  assign n1095 = n1092 | n1094 ;
  assign n1096 = ( n1078 & ~n1093 ) | ( n1078 & n1095 ) | ( ~n1093 & n1095 ) ;
  assign n1097 = ~x25 & x152 ;
  assign n1098 = x153 | x154 ;
  assign n1099 = n1097 | n1098 ;
  assign n1100 = ~x22 & x149 ;
  assign n1101 = x150 | x151 ;
  assign n1102 = n1100 | n1101 ;
  assign n1103 = ~x19 & x146 ;
  assign n1104 = x147 | x148 ;
  assign n1105 = n1103 | n1104 ;
  assign n1106 = x20 & ~x148 ;
  assign n1107 = x21 | x22 ;
  assign n1108 = n1106 | n1107 ;
  assign n1109 = n1105 & ~n1108 ;
  assign n1110 = n1102 | n1109 ;
  assign n1111 = x23 & ~x151 ;
  assign n1112 = x24 | x25 ;
  assign n1113 = n1111 | n1112 ;
  assign n1114 = n1110 & ~n1113 ;
  assign n1115 = n1099 | n1114 ;
  assign n1116 = ~n1102 & n1108 ;
  assign n1117 = n1113 | n1116 ;
  assign n1118 = ~n1099 & n1117 ;
  assign n1119 = ( n1096 & ~n1115 ) | ( n1096 & n1118 ) | ( ~n1115 & n1118 ) ;
  assign n1120 = ~x34 & x161 ;
  assign n1121 = x162 | x163 ;
  assign n1122 = n1120 | n1121 ;
  assign n1123 = ~x31 & x158 ;
  assign n1124 = x159 | x160 ;
  assign n1125 = n1123 | n1124 ;
  assign n1126 = ~x28 & x155 ;
  assign n1127 = x156 | x157 ;
  assign n1128 = n1126 | n1127 ;
  assign n1129 = x26 & ~x154 ;
  assign n1130 = x27 | x28 ;
  assign n1131 = n1129 | n1130 ;
  assign n1132 = ~n1128 & n1131 ;
  assign n1133 = x29 & ~x157 ;
  assign n1134 = x30 | x31 ;
  assign n1135 = n1133 | n1134 ;
  assign n1136 = n1132 | n1135 ;
  assign n1137 = ~n1125 & n1136 ;
  assign n1138 = x32 & ~x160 ;
  assign n1139 = x33 | x34 ;
  assign n1140 = n1138 | n1139 ;
  assign n1141 = n1137 | n1140 ;
  assign n1142 = ~n1122 & n1141 ;
  assign n1143 = n1128 & ~n1135 ;
  assign n1144 = n1125 & ~n1140 ;
  assign n1145 = ( ~n1140 & n1143 ) | ( ~n1140 & n1144 ) | ( n1143 & n1144 ) ;
  assign n1146 = n1122 | n1145 ;
  assign n1147 = ( n1119 & n1142 ) | ( n1119 & ~n1146 ) | ( n1142 & ~n1146 ) ;
  assign n1148 = ~x43 & x170 ;
  assign n1149 = x171 | x172 ;
  assign n1150 = n1148 | n1149 ;
  assign n1151 = ~x40 & x167 ;
  assign n1152 = x168 | x169 ;
  assign n1153 = n1151 | n1152 ;
  assign n1154 = ~x37 & x164 ;
  assign n1155 = x165 | x166 ;
  assign n1156 = n1154 | n1155 ;
  assign n1157 = x35 & ~x163 ;
  assign n1158 = x36 | x37 ;
  assign n1159 = n1157 | n1158 ;
  assign n1160 = ~n1156 & n1159 ;
  assign n1161 = x38 & ~x166 ;
  assign n1162 = x39 | x40 ;
  assign n1163 = n1161 | n1162 ;
  assign n1164 = n1160 | n1163 ;
  assign n1165 = ~n1153 & n1164 ;
  assign n1166 = x41 & ~x169 ;
  assign n1167 = x42 | x43 ;
  assign n1168 = n1166 | n1167 ;
  assign n1169 = n1165 | n1168 ;
  assign n1170 = ~n1150 & n1169 ;
  assign n1171 = x44 & ~x172 ;
  assign n1172 = x45 | x46 ;
  assign n1173 = n1171 | n1172 ;
  assign n1174 = n1170 | n1173 ;
  assign n1175 = n1156 & ~n1163 ;
  assign n1176 = n1153 & ~n1168 ;
  assign n1177 = ( ~n1168 & n1175 ) | ( ~n1168 & n1176 ) | ( n1175 & n1176 ) ;
  assign n1178 = n1150 | n1177 ;
  assign n1179 = ~n1173 & n1178 ;
  assign n1180 = ( n1147 & n1174 ) | ( n1147 & ~n1179 ) | ( n1174 & ~n1179 ) ;
  assign n1181 = x56 & ~x184 ;
  assign n1182 = x57 | x58 ;
  assign n1183 = n1181 | n1182 ;
  assign n1184 = ~x55 & x182 ;
  assign n1185 = x183 | x184 ;
  assign n1186 = n1184 | n1185 ;
  assign n1187 = x53 & ~x181 ;
  assign n1188 = x54 | x55 ;
  assign n1189 = n1187 | n1188 ;
  assign n1190 = ~x52 & x179 ;
  assign n1191 = x180 | x181 ;
  assign n1192 = n1190 | n1191 ;
  assign n1193 = x50 & ~x178 ;
  assign n1194 = x51 | x52 ;
  assign n1195 = n1193 | n1194 ;
  assign n1196 = ~x49 & x176 ;
  assign n1197 = x177 | x178 ;
  assign n1198 = n1196 | n1197 ;
  assign n1199 = x47 & ~x175 ;
  assign n1200 = x48 | x49 ;
  assign n1201 = n1199 | n1200 ;
  assign n1202 = ~n1198 & n1201 ;
  assign n1203 = n1195 | n1202 ;
  assign n1204 = ~n1192 & n1203 ;
  assign n1205 = n1189 | n1204 ;
  assign n1206 = ~n1186 & n1205 ;
  assign n1207 = n1183 | n1206 ;
  assign n1208 = ~x46 & x173 ;
  assign n1209 = x174 | x175 ;
  assign n1210 = n1208 | n1209 ;
  assign n1211 = ~n1201 & n1210 ;
  assign n1212 = ~n1195 & n1198 ;
  assign n1213 = ( ~n1195 & n1211 ) | ( ~n1195 & n1212 ) | ( n1211 & n1212 ) ;
  assign n1214 = n1192 | n1213 ;
  assign n1215 = ~n1189 & n1214 ;
  assign n1216 = ~n1183 & n1186 ;
  assign n1217 = ( ~n1183 & n1215 ) | ( ~n1183 & n1216 ) | ( n1215 & n1216 ) ;
  assign n1218 = ( n1180 & n1207 ) | ( n1180 & ~n1217 ) | ( n1207 & ~n1217 ) ;
  assign n1219 = ~x70 & x197 ;
  assign n1220 = x198 | x199 ;
  assign n1221 = n1219 | n1220 ;
  assign n1222 = ~x64 & x191 ;
  assign n1223 = x192 | x193 ;
  assign n1224 = n1222 | n1223 ;
  assign n1225 = ~x61 & x188 ;
  assign n1226 = x189 | x190 ;
  assign n1227 = n1225 | n1226 ;
  assign n1228 = ~x58 & x185 ;
  assign n1229 = x186 | x187 ;
  assign n1230 = n1228 | n1229 ;
  assign n1231 = x59 & ~x187 ;
  assign n1232 = x60 | x61 ;
  assign n1233 = n1231 | n1232 ;
  assign n1234 = n1230 & ~n1233 ;
  assign n1235 = n1227 | n1234 ;
  assign n1236 = x62 & ~x190 ;
  assign n1237 = x63 | x64 ;
  assign n1238 = n1236 | n1237 ;
  assign n1239 = n1235 & ~n1238 ;
  assign n1240 = n1224 | n1239 ;
  assign n1241 = x65 & ~x193 ;
  assign n1242 = x66 | x67 ;
  assign n1243 = n1241 | n1242 ;
  assign n1244 = n1240 & ~n1243 ;
  assign n1245 = x68 & ~x196 ;
  assign n1246 = x69 | x70 ;
  assign n1247 = n1245 | n1246 ;
  assign n1248 = ~x67 & x194 ;
  assign n1249 = x195 | x196 ;
  assign n1250 = n1248 | n1249 ;
  assign n1251 = ~n1247 & n1250 ;
  assign n1252 = ( n1244 & ~n1247 ) | ( n1244 & n1251 ) | ( ~n1247 & n1251 ) ;
  assign n1253 = n1221 | n1252 ;
  assign n1254 = ~n1227 & n1233 ;
  assign n1255 = n1238 | n1254 ;
  assign n1256 = ~n1224 & n1255 ;
  assign n1257 = n1243 | n1256 ;
  assign n1258 = ~n1250 & n1257 ;
  assign n1259 = n1247 | n1258 ;
  assign n1260 = ~n1221 & n1259 ;
  assign n1261 = ( n1218 & ~n1253 ) | ( n1218 & n1260 ) | ( ~n1253 & n1260 ) ;
  assign n1262 = ~x85 & x212 ;
  assign n1263 = x213 | x214 ;
  assign n1264 = n1262 | n1263 ;
  assign n1265 = x83 & ~x211 ;
  assign n1266 = x84 | x85 ;
  assign n1267 = n1265 | n1266 ;
  assign n1268 = x80 & ~x208 ;
  assign n1269 = x81 | x82 ;
  assign n1270 = n1268 | n1269 ;
  assign n1271 = ~x79 & x206 ;
  assign n1272 = x207 | x208 ;
  assign n1273 = n1271 | n1272 ;
  assign n1274 = x77 & ~x205 ;
  assign n1275 = x78 | x79 ;
  assign n1276 = n1274 | n1275 ;
  assign n1277 = ~x73 & x200 ;
  assign n1278 = x201 | x202 ;
  assign n1279 = n1277 | n1278 ;
  assign n1280 = x74 & ~x202 ;
  assign n1281 = x75 | x76 ;
  assign n1282 = n1280 | n1281 ;
  assign n1283 = n1279 & ~n1282 ;
  assign n1284 = ~x76 & x203 ;
  assign n1285 = x204 | x205 ;
  assign n1286 = n1284 | n1285 ;
  assign n1287 = ~n1276 & n1286 ;
  assign n1288 = ( ~n1276 & n1283 ) | ( ~n1276 & n1287 ) | ( n1283 & n1287 ) ;
  assign n1289 = n1273 | n1288 ;
  assign n1290 = ~n1270 & n1289 ;
  assign n1291 = ~x82 & x209 ;
  assign n1292 = x210 | x211 ;
  assign n1293 = n1291 | n1292 ;
  assign n1294 = ~n1267 & n1293 ;
  assign n1295 = ( ~n1267 & n1290 ) | ( ~n1267 & n1294 ) | ( n1290 & n1294 ) ;
  assign n1296 = n1264 | n1295 ;
  assign n1297 = x71 & ~x199 ;
  assign n1298 = x72 | x73 ;
  assign n1299 = n1297 | n1298 ;
  assign n1300 = ~n1279 & n1299 ;
  assign n1301 = n1282 | n1300 ;
  assign n1302 = ~n1286 & n1301 ;
  assign n1303 = n1276 | n1302 ;
  assign n1304 = ~n1273 & n1303 ;
  assign n1305 = n1270 | n1304 ;
  assign n1306 = ~n1293 & n1305 ;
  assign n1307 = ~n1264 & n1267 ;
  assign n1308 = ( ~n1264 & n1306 ) | ( ~n1264 & n1307 ) | ( n1306 & n1307 ) ;
  assign n1309 = ( n1261 & ~n1296 ) | ( n1261 & n1308 ) | ( ~n1296 & n1308 ) ;
  assign n1310 = x101 & ~x229 ;
  assign n1311 = x102 | x103 ;
  assign n1312 = n1310 | n1311 ;
  assign n1313 = ~x100 & x227 ;
  assign n1314 = x228 | x229 ;
  assign n1315 = n1313 | n1314 ;
  assign n1316 = ~x97 & x224 ;
  assign n1317 = x225 | x226 ;
  assign n1318 = n1316 | n1317 ;
  assign n1319 = ~x94 & x221 ;
  assign n1320 = x222 | x223 ;
  assign n1321 = n1319 | n1320 ;
  assign n1322 = ~x91 & x218 ;
  assign n1323 = x219 | x220 ;
  assign n1324 = n1322 | n1323 ;
  assign n1325 = ~x88 & x215 ;
  assign n1326 = x216 | x217 ;
  assign n1327 = n1325 | n1326 ;
  assign n1328 = x86 & ~x214 ;
  assign n1329 = x87 | x88 ;
  assign n1330 = n1328 | n1329 ;
  assign n1331 = ~n1327 & n1330 ;
  assign n1332 = x89 & ~x217 ;
  assign n1333 = x90 | x91 ;
  assign n1334 = n1332 | n1333 ;
  assign n1335 = n1331 | n1334 ;
  assign n1336 = ~n1324 & n1335 ;
  assign n1337 = x92 & ~x220 ;
  assign n1338 = x93 | x94 ;
  assign n1339 = n1337 | n1338 ;
  assign n1340 = n1336 | n1339 ;
  assign n1341 = ~n1321 & n1340 ;
  assign n1342 = x95 & ~x223 ;
  assign n1343 = x96 | x97 ;
  assign n1344 = n1342 | n1343 ;
  assign n1345 = n1341 | n1344 ;
  assign n1346 = ~n1318 & n1345 ;
  assign n1347 = x98 & ~x226 ;
  assign n1348 = x99 | x100 ;
  assign n1349 = n1347 | n1348 ;
  assign n1350 = ~n1315 & n1349 ;
  assign n1351 = ( ~n1315 & n1346 ) | ( ~n1315 & n1350 ) | ( n1346 & n1350 ) ;
  assign n1352 = n1312 | n1351 ;
  assign n1353 = n1327 & ~n1334 ;
  assign n1354 = n1324 & ~n1339 ;
  assign n1355 = ( ~n1339 & n1353 ) | ( ~n1339 & n1354 ) | ( n1353 & n1354 ) ;
  assign n1356 = n1321 | n1355 ;
  assign n1357 = ~n1344 & n1356 ;
  assign n1358 = n1318 & ~n1349 ;
  assign n1359 = ( ~n1349 & n1357 ) | ( ~n1349 & n1358 ) | ( n1357 & n1358 ) ;
  assign n1360 = n1315 | n1359 ;
  assign n1361 = ~n1312 & n1360 ;
  assign n1362 = ( n1309 & n1352 ) | ( n1309 & ~n1361 ) | ( n1352 & ~n1361 ) ;
  assign n1363 = x119 & ~x247 ;
  assign n1364 = x120 | x121 ;
  assign n1365 = n1363 | n1364 ;
  assign n1366 = ~x118 & x245 ;
  assign n1367 = x246 | x247 ;
  assign n1368 = n1366 | n1367 ;
  assign n1369 = ~x115 & x242 ;
  assign n1370 = x243 | x244 ;
  assign n1371 = n1369 | n1370 ;
  assign n1372 = x113 & ~x241 ;
  assign n1373 = x114 | x115 ;
  assign n1374 = n1372 | n1373 ;
  assign n1375 = ~x112 & x239 ;
  assign n1376 = x240 | x241 ;
  assign n1377 = n1375 | n1376 ;
  assign n1378 = x110 & ~x238 ;
  assign n1379 = x111 | x112 ;
  assign n1380 = n1378 | n1379 ;
  assign n1381 = ~x109 & x236 ;
  assign n1382 = x237 | x238 ;
  assign n1383 = n1381 | n1382 ;
  assign n1384 = x107 & ~x235 ;
  assign n1385 = x108 | x109 ;
  assign n1386 = n1384 | n1385 ;
  assign n1387 = ~x106 & x233 ;
  assign n1388 = x234 | x235 ;
  assign n1389 = n1387 | n1388 ;
  assign n1390 = x104 & ~x232 ;
  assign n1391 = x105 | x106 ;
  assign n1392 = n1390 | n1391 ;
  assign n1393 = ~n1389 & n1392 ;
  assign n1394 = n1386 | n1393 ;
  assign n1395 = ~n1383 & n1394 ;
  assign n1396 = n1380 | n1395 ;
  assign n1397 = ~n1377 & n1396 ;
  assign n1398 = n1374 | n1397 ;
  assign n1399 = ~n1371 & n1398 ;
  assign n1400 = x116 & ~x244 ;
  assign n1401 = x117 | x118 ;
  assign n1402 = n1400 | n1401 ;
  assign n1403 = ~n1368 & n1402 ;
  assign n1404 = ( ~n1368 & n1399 ) | ( ~n1368 & n1403 ) | ( n1399 & n1403 ) ;
  assign n1405 = n1365 | n1404 ;
  assign n1406 = ~x103 & x230 ;
  assign n1407 = x231 | x232 ;
  assign n1408 = n1406 | n1407 ;
  assign n1409 = ~n1392 & n1408 ;
  assign n1410 = ~n1386 & n1389 ;
  assign n1411 = ( ~n1386 & n1409 ) | ( ~n1386 & n1410 ) | ( n1409 & n1410 ) ;
  assign n1412 = n1383 | n1411 ;
  assign n1413 = ~n1380 & n1412 ;
  assign n1414 = ~n1374 & n1377 ;
  assign n1415 = ( ~n1374 & n1413 ) | ( ~n1374 & n1414 ) | ( n1413 & n1414 ) ;
  assign n1416 = n1371 | n1415 ;
  assign n1417 = ~n1402 & n1416 ;
  assign n1418 = ~n1365 & n1368 ;
  assign n1419 = ( ~n1365 & n1417 ) | ( ~n1365 & n1418 ) | ( n1417 & n1418 ) ;
  assign n1420 = ( n1362 & n1405 ) | ( n1362 & ~n1419 ) | ( n1405 & ~n1419 ) ;
  assign n1421 = ~x127 & x254 ;
  assign n1422 = x128 | x255 ;
  assign n1423 = n1421 | n1422 ;
  assign n1424 = ~x124 & x251 ;
  assign n1425 = x252 | x253 ;
  assign n1426 = n1424 | n1425 ;
  assign n1427 = ~x121 & x248 ;
  assign n1428 = x249 | x250 ;
  assign n1429 = n1427 | n1428 ;
  assign n1430 = x122 & ~x250 ;
  assign n1431 = x123 | x124 ;
  assign n1432 = n1430 | n1431 ;
  assign n1433 = n1429 & ~n1432 ;
  assign n1434 = n1426 | n1433 ;
  assign n1435 = x125 & ~x253 ;
  assign n1436 = x126 | x127 ;
  assign n1437 = n1435 | n1436 ;
  assign n1438 = n1434 & ~n1437 ;
  assign n1439 = n1423 | n1438 ;
  assign n1440 = x0 & ~x128 ;
  assign n1441 = x1 | x2 ;
  assign n1442 = n1440 | n1441 ;
  assign n1443 = n1439 & ~n1442 ;
  assign n1444 = ~n1426 & n1432 ;
  assign n1445 = n1437 | n1444 ;
  assign n1446 = ~n1423 & n1445 ;
  assign n1447 = n1442 | n1446 ;
  assign n1448 = ( n1420 & ~n1443 ) | ( n1420 & n1447 ) | ( ~n1443 & n1447 ) ;
  assign n1449 = n1054 & n1448 ;
  assign n1450 = ~x3 & x130 ;
  assign n1451 = x131 & ~n1450 ;
  assign n1452 = x5 | n664 ;
  assign n1453 = ~n264 & n1452 ;
  assign n1454 = ( ~n273 & n277 ) | ( ~n273 & n1453 ) | ( n277 & n1453 ) ;
  assign n1455 = n280 & ~n289 ;
  assign n1456 = n292 | n1455 ;
  assign n1457 = ( ~n293 & n1454 ) | ( ~n293 & n1456 ) | ( n1454 & n1456 ) ;
  assign n1458 = n297 & ~n310 ;
  assign n1459 = n313 | n1458 ;
  assign n1460 = n286 & ~n297 ;
  assign n1461 = ( ~n313 & n314 ) | ( ~n313 & n1460 ) | ( n314 & n1460 ) ;
  assign n1462 = ( n1457 & n1459 ) | ( n1457 & ~n1461 ) | ( n1459 & ~n1461 ) ;
  assign n1463 = n307 & ~n318 ;
  assign n1464 = n304 & ~n336 ;
  assign n1465 = ( ~n336 & n1463 ) | ( ~n336 & n1464 ) | ( n1463 & n1464 ) ;
  assign n1466 = n333 | n1465 ;
  assign n1467 = ~n304 & n318 ;
  assign n1468 = n336 | n1467 ;
  assign n1469 = ~n333 & n1468 ;
  assign n1470 = ( n1462 & ~n1466 ) | ( n1462 & n1469 ) | ( ~n1466 & n1469 ) ;
  assign n1471 = ~n330 & n340 ;
  assign n1472 = n345 | n1471 ;
  assign n1473 = ~n327 & n1472 ;
  assign n1474 = n364 | n1473 ;
  assign n1475 = ~n361 & n1474 ;
  assign n1476 = n327 & ~n364 ;
  assign n1477 = ( n349 & ~n364 ) | ( n349 & n1476 ) | ( ~n364 & n1476 ) ;
  assign n1478 = n361 | n1477 ;
  assign n1479 = ( n1470 & n1475 ) | ( n1470 & ~n1478 ) | ( n1475 & ~n1478 ) ;
  assign n1480 = ~n358 & n368 ;
  assign n1481 = n373 | n1480 ;
  assign n1482 = ~n355 & n1481 ;
  assign n1483 = n378 | n1482 ;
  assign n1484 = ~n415 & n1483 ;
  assign n1485 = n406 | n1484 ;
  assign n1486 = n355 & ~n378 ;
  assign n1487 = ( ~n378 & n381 ) | ( ~n378 & n1486 ) | ( n381 & n1486 ) ;
  assign n1488 = n415 | n1487 ;
  assign n1489 = ~n406 & n1488 ;
  assign n1490 = ( n1479 & n1485 ) | ( n1479 & ~n1489 ) | ( n1485 & ~n1489 ) ;
  assign n1491 = ~n397 & n400 ;
  assign n1492 = n394 | n1491 ;
  assign n1493 = ~n391 & n1492 ;
  assign n1494 = n388 | n1493 ;
  assign n1495 = ~n435 & n1494 ;
  assign n1496 = n438 | n1495 ;
  assign n1497 = ~n394 & n397 ;
  assign n1498 = ( ~n394 & n417 ) | ( ~n394 & n1497 ) | ( n417 & n1497 ) ;
  assign n1499 = n391 | n1498 ;
  assign n1500 = ~n388 & n1499 ;
  assign n1501 = ( ~n438 & n439 ) | ( ~n438 & n1500 ) | ( n439 & n1500 ) ;
  assign n1502 = ( n1490 & n1496 ) | ( n1490 & ~n1501 ) | ( n1496 & ~n1501 ) ;
  assign n1503 = n432 & ~n443 ;
  assign n1504 = n429 & ~n448 ;
  assign n1505 = ( ~n448 & n1503 ) | ( ~n448 & n1504 ) | ( n1503 & n1504 ) ;
  assign n1506 = n455 | n1505 ;
  assign n1507 = ~n452 & n1506 ;
  assign n1508 = n426 & ~n504 ;
  assign n1509 = ( ~n504 & n1507 ) | ( ~n504 & n1508 ) | ( n1507 & n1508 ) ;
  assign n1510 = n484 | n1509 ;
  assign n1511 = ~n429 & n443 ;
  assign n1512 = n448 | n1511 ;
  assign n1513 = ~n455 & n1512 ;
  assign n1514 = n452 | n1513 ;
  assign n1515 = ~n426 & n1514 ;
  assign n1516 = n504 | n1515 ;
  assign n1517 = ~n484 & n1516 ;
  assign n1518 = ( n1502 & ~n1510 ) | ( n1502 & n1517 ) | ( ~n1510 & n1517 ) ;
  assign n1519 = ~n475 & n478 ;
  assign n1520 = ( ~n475 & n492 ) | ( ~n475 & n1519 ) | ( n492 & n1519 ) ;
  assign n1521 = n498 | n1520 ;
  assign n1522 = ~n472 & n1521 ;
  assign n1523 = n469 & ~n535 ;
  assign n1524 = ( ~n535 & n1522 ) | ( ~n535 & n1523 ) | ( n1522 & n1523 ) ;
  assign n1525 = n532 | n1524 ;
  assign n1526 = n487 & ~n491 ;
  assign n1527 = n481 | n1526 ;
  assign n1528 = ~n478 & n1527 ;
  assign n1529 = n475 | n1528 ;
  assign n1530 = ~n498 & n1529 ;
  assign n1531 = n472 | n1530 ;
  assign n1532 = ~n469 & n1531 ;
  assign n1533 = ( ~n532 & n536 ) | ( ~n532 & n1532 ) | ( n536 & n1532 ) ;
  assign n1534 = ( n1518 & ~n1525 ) | ( n1518 & n1533 ) | ( ~n1525 & n1533 ) ;
  assign n1535 = ~n529 & n539 ;
  assign n1536 = n544 | n1535 ;
  assign n1537 = ~n526 & n1536 ;
  assign n1538 = n549 | n1537 ;
  assign n1539 = ~n523 & n1538 ;
  assign n1540 = n554 | n1539 ;
  assign n1541 = ~n520 & n1540 ;
  assign n1542 = n517 & ~n613 ;
  assign n1543 = ( ~n613 & n1541 ) | ( ~n613 & n1542 ) | ( n1541 & n1542 ) ;
  assign n1544 = n597 | n1543 ;
  assign n1545 = n526 & ~n549 ;
  assign n1546 = ( ~n549 & n559 ) | ( ~n549 & n1545 ) | ( n559 & n1545 ) ;
  assign n1547 = n523 | n1546 ;
  assign n1548 = ~n554 & n1547 ;
  assign n1549 = ~n517 & n520 ;
  assign n1550 = ( ~n517 & n1548 ) | ( ~n517 & n1549 ) | ( n1548 & n1549 ) ;
  assign n1551 = n613 | n1550 ;
  assign n1552 = ~n597 & n1551 ;
  assign n1553 = ( n1534 & n1544 ) | ( n1534 & ~n1552 ) | ( n1544 & ~n1552 ) ;
  assign n1554 = ~n588 & n591 ;
  assign n1555 = n585 | n1554 ;
  assign n1556 = ~n582 & n1555 ;
  assign n1557 = n579 | n1556 ;
  assign n1558 = ~n576 & n1557 ;
  assign n1559 = n607 | n1558 ;
  assign n1560 = ~n573 & n1559 ;
  assign n1561 = n570 & ~n634 ;
  assign n1562 = ( ~n634 & n1560 ) | ( ~n634 & n1561 ) | ( n1560 & n1561 ) ;
  assign n1563 = n637 | n1562 ;
  assign n1564 = ~n585 & n588 ;
  assign n1565 = ( ~n585 & n615 ) | ( ~n585 & n1564 ) | ( n615 & n1564 ) ;
  assign n1566 = n582 | n1565 ;
  assign n1567 = ~n579 & n1566 ;
  assign n1568 = n576 & ~n607 ;
  assign n1569 = ( ~n607 & n1567 ) | ( ~n607 & n1568 ) | ( n1567 & n1568 ) ;
  assign n1570 = n573 | n1569 ;
  assign n1571 = ~n570 & n1570 ;
  assign n1572 = ( ~n637 & n638 ) | ( ~n637 & n1571 ) | ( n638 & n1571 ) ;
  assign n1573 = ( n1553 & n1563 ) | ( n1553 & ~n1572 ) | ( n1563 & ~n1572 ) ;
  assign n1574 = x128 | x129 ;
  assign n1575 = n257 | n1574 ;
  assign n1576 = n631 & ~n642 ;
  assign n1577 = n628 & ~n647 ;
  assign n1578 = ( ~n647 & n1576 ) | ( ~n647 & n1577 ) | ( n1576 & n1577 ) ;
  assign n1579 = n1575 | n1578 ;
  assign n1580 = x2 | x3 ;
  assign n1581 = n259 | n1580 ;
  assign n1582 = n1579 & ~n1581 ;
  assign n1583 = ~n628 & n642 ;
  assign n1584 = n647 | n1583 ;
  assign n1585 = ~n1575 & n1584 ;
  assign n1586 = n1581 | n1585 ;
  assign n1587 = ( n1573 & ~n1582 ) | ( n1573 & n1586 ) | ( ~n1582 & n1586 ) ;
  assign n1588 = n1451 & n1587 ;
  assign n1589 = ~x4 & x131 ;
  assign n1590 = x132 & ~n1589 ;
  assign n1591 = x6 | n1061 ;
  assign n1592 = ~n662 & n1591 ;
  assign n1593 = ( ~n671 & n675 ) | ( ~n671 & n1592 ) | ( n675 & n1592 ) ;
  assign n1594 = n678 & ~n687 ;
  assign n1595 = n690 | n1594 ;
  assign n1596 = ( ~n691 & n1593 ) | ( ~n691 & n1595 ) | ( n1593 & n1595 ) ;
  assign n1597 = n695 & ~n708 ;
  assign n1598 = n711 | n1597 ;
  assign n1599 = n684 & ~n695 ;
  assign n1600 = ( ~n711 & n712 ) | ( ~n711 & n1599 ) | ( n712 & n1599 ) ;
  assign n1601 = ( n1596 & n1598 ) | ( n1596 & ~n1600 ) | ( n1598 & ~n1600 ) ;
  assign n1602 = n705 & ~n716 ;
  assign n1603 = n702 & ~n734 ;
  assign n1604 = ( ~n734 & n1602 ) | ( ~n734 & n1603 ) | ( n1602 & n1603 ) ;
  assign n1605 = n731 | n1604 ;
  assign n1606 = ~n702 & n716 ;
  assign n1607 = n734 | n1606 ;
  assign n1608 = ~n731 & n1607 ;
  assign n1609 = ( n1601 & ~n1605 ) | ( n1601 & n1608 ) | ( ~n1605 & n1608 ) ;
  assign n1610 = ~n728 & n738 ;
  assign n1611 = n743 | n1610 ;
  assign n1612 = ~n725 & n1611 ;
  assign n1613 = n762 | n1612 ;
  assign n1614 = ~n759 & n1613 ;
  assign n1615 = n725 & ~n762 ;
  assign n1616 = ( n747 & ~n762 ) | ( n747 & n1615 ) | ( ~n762 & n1615 ) ;
  assign n1617 = n759 | n1616 ;
  assign n1618 = ( n1609 & n1614 ) | ( n1609 & ~n1617 ) | ( n1614 & ~n1617 ) ;
  assign n1619 = ~n756 & n766 ;
  assign n1620 = n771 | n1619 ;
  assign n1621 = ~n753 & n1620 ;
  assign n1622 = n776 | n1621 ;
  assign n1623 = ~n813 & n1622 ;
  assign n1624 = n804 | n1623 ;
  assign n1625 = n753 & ~n776 ;
  assign n1626 = ( ~n776 & n779 ) | ( ~n776 & n1625 ) | ( n779 & n1625 ) ;
  assign n1627 = n813 | n1626 ;
  assign n1628 = ~n804 & n1627 ;
  assign n1629 = ( n1618 & n1624 ) | ( n1618 & ~n1628 ) | ( n1624 & ~n1628 ) ;
  assign n1630 = ~n795 & n798 ;
  assign n1631 = n792 | n1630 ;
  assign n1632 = ~n789 & n1631 ;
  assign n1633 = n786 | n1632 ;
  assign n1634 = ~n833 & n1633 ;
  assign n1635 = n836 | n1634 ;
  assign n1636 = ~n792 & n795 ;
  assign n1637 = ( ~n792 & n815 ) | ( ~n792 & n1636 ) | ( n815 & n1636 ) ;
  assign n1638 = n789 | n1637 ;
  assign n1639 = ~n786 & n1638 ;
  assign n1640 = ( ~n836 & n837 ) | ( ~n836 & n1639 ) | ( n837 & n1639 ) ;
  assign n1641 = ( n1629 & n1635 ) | ( n1629 & ~n1640 ) | ( n1635 & ~n1640 ) ;
  assign n1642 = n830 & ~n841 ;
  assign n1643 = n827 & ~n846 ;
  assign n1644 = ( ~n846 & n1642 ) | ( ~n846 & n1643 ) | ( n1642 & n1643 ) ;
  assign n1645 = n853 | n1644 ;
  assign n1646 = ~n850 & n1645 ;
  assign n1647 = n824 & ~n902 ;
  assign n1648 = ( ~n902 & n1646 ) | ( ~n902 & n1647 ) | ( n1646 & n1647 ) ;
  assign n1649 = n882 | n1648 ;
  assign n1650 = ~n827 & n841 ;
  assign n1651 = n846 | n1650 ;
  assign n1652 = ~n853 & n1651 ;
  assign n1653 = n850 | n1652 ;
  assign n1654 = ~n824 & n1653 ;
  assign n1655 = n902 | n1654 ;
  assign n1656 = ~n882 & n1655 ;
  assign n1657 = ( n1641 & ~n1649 ) | ( n1641 & n1656 ) | ( ~n1649 & n1656 ) ;
  assign n1658 = ~n873 & n876 ;
  assign n1659 = ( ~n873 & n890 ) | ( ~n873 & n1658 ) | ( n890 & n1658 ) ;
  assign n1660 = n896 | n1659 ;
  assign n1661 = ~n870 & n1660 ;
  assign n1662 = n867 & ~n933 ;
  assign n1663 = ( ~n933 & n1661 ) | ( ~n933 & n1662 ) | ( n1661 & n1662 ) ;
  assign n1664 = n930 | n1663 ;
  assign n1665 = n885 & ~n889 ;
  assign n1666 = n879 | n1665 ;
  assign n1667 = ~n876 & n1666 ;
  assign n1668 = n873 | n1667 ;
  assign n1669 = ~n896 & n1668 ;
  assign n1670 = n870 | n1669 ;
  assign n1671 = ~n867 & n1670 ;
  assign n1672 = ( ~n930 & n934 ) | ( ~n930 & n1671 ) | ( n934 & n1671 ) ;
  assign n1673 = ( n1657 & ~n1664 ) | ( n1657 & n1672 ) | ( ~n1664 & n1672 ) ;
  assign n1674 = ~n927 & n937 ;
  assign n1675 = n942 | n1674 ;
  assign n1676 = ~n924 & n1675 ;
  assign n1677 = n947 | n1676 ;
  assign n1678 = ~n921 & n1677 ;
  assign n1679 = n952 | n1678 ;
  assign n1680 = ~n918 & n1679 ;
  assign n1681 = n915 & ~n1011 ;
  assign n1682 = ( ~n1011 & n1680 ) | ( ~n1011 & n1681 ) | ( n1680 & n1681 ) ;
  assign n1683 = n995 | n1682 ;
  assign n1684 = n924 & ~n947 ;
  assign n1685 = ( ~n947 & n957 ) | ( ~n947 & n1684 ) | ( n957 & n1684 ) ;
  assign n1686 = n921 | n1685 ;
  assign n1687 = ~n952 & n1686 ;
  assign n1688 = ~n915 & n918 ;
  assign n1689 = ( ~n915 & n1687 ) | ( ~n915 & n1688 ) | ( n1687 & n1688 ) ;
  assign n1690 = n1011 | n1689 ;
  assign n1691 = ~n995 & n1690 ;
  assign n1692 = ( n1673 & n1683 ) | ( n1673 & ~n1691 ) | ( n1683 & ~n1691 ) ;
  assign n1693 = ~n986 & n989 ;
  assign n1694 = n983 | n1693 ;
  assign n1695 = ~n980 & n1694 ;
  assign n1696 = n977 | n1695 ;
  assign n1697 = ~n974 & n1696 ;
  assign n1698 = n1005 | n1697 ;
  assign n1699 = ~n971 & n1698 ;
  assign n1700 = n968 & ~n1032 ;
  assign n1701 = ( ~n1032 & n1699 ) | ( ~n1032 & n1700 ) | ( n1699 & n1700 ) ;
  assign n1702 = n1035 | n1701 ;
  assign n1703 = ~n983 & n986 ;
  assign n1704 = ( ~n983 & n1013 ) | ( ~n983 & n1703 ) | ( n1013 & n1703 ) ;
  assign n1705 = n980 | n1704 ;
  assign n1706 = ~n977 & n1705 ;
  assign n1707 = n974 & ~n1005 ;
  assign n1708 = ( ~n1005 & n1706 ) | ( ~n1005 & n1707 ) | ( n1706 & n1707 ) ;
  assign n1709 = n971 | n1708 ;
  assign n1710 = ~n968 & n1709 ;
  assign n1711 = ( ~n1035 & n1036 ) | ( ~n1035 & n1710 ) | ( n1036 & n1710 ) ;
  assign n1712 = ( n1692 & n1702 ) | ( n1692 & ~n1711 ) | ( n1702 & ~n1711 ) ;
  assign n1713 = x129 | x130 ;
  assign n1714 = n655 | n1713 ;
  assign n1715 = n1029 & ~n1040 ;
  assign n1716 = n1026 & ~n1045 ;
  assign n1717 = ( ~n1045 & n1715 ) | ( ~n1045 & n1716 ) | ( n1715 & n1716 ) ;
  assign n1718 = n1714 | n1717 ;
  assign n1719 = x3 | x4 ;
  assign n1720 = n657 | n1719 ;
  assign n1721 = n1718 & ~n1720 ;
  assign n1722 = ~n1026 & n1040 ;
  assign n1723 = n1045 | n1722 ;
  assign n1724 = ~n1714 & n1723 ;
  assign n1725 = n1720 | n1724 ;
  assign n1726 = ( n1712 & ~n1721 ) | ( n1712 & n1725 ) | ( ~n1721 & n1725 ) ;
  assign n1727 = n1590 & n1726 ;
  assign n1728 = x133 & ~n263 ;
  assign n1729 = x7 | n274 ;
  assign n1730 = ~n1059 & n1729 ;
  assign n1731 = ( ~n1068 & n1072 ) | ( ~n1068 & n1730 ) | ( n1072 & n1730 ) ;
  assign n1732 = n1075 & ~n1084 ;
  assign n1733 = n1087 | n1732 ;
  assign n1734 = ( ~n1088 & n1731 ) | ( ~n1088 & n1733 ) | ( n1731 & n1733 ) ;
  assign n1735 = n1092 & ~n1105 ;
  assign n1736 = n1108 | n1735 ;
  assign n1737 = n1081 & ~n1092 ;
  assign n1738 = ( ~n1108 & n1109 ) | ( ~n1108 & n1737 ) | ( n1109 & n1737 ) ;
  assign n1739 = ( n1734 & n1736 ) | ( n1734 & ~n1738 ) | ( n1736 & ~n1738 ) ;
  assign n1740 = n1102 & ~n1113 ;
  assign n1741 = n1099 & ~n1131 ;
  assign n1742 = ( ~n1131 & n1740 ) | ( ~n1131 & n1741 ) | ( n1740 & n1741 ) ;
  assign n1743 = n1128 | n1742 ;
  assign n1744 = ~n1099 & n1113 ;
  assign n1745 = n1131 | n1744 ;
  assign n1746 = ~n1128 & n1745 ;
  assign n1747 = ( n1739 & ~n1743 ) | ( n1739 & n1746 ) | ( ~n1743 & n1746 ) ;
  assign n1748 = ~n1125 & n1135 ;
  assign n1749 = n1140 | n1748 ;
  assign n1750 = ~n1122 & n1749 ;
  assign n1751 = n1159 | n1750 ;
  assign n1752 = ~n1156 & n1751 ;
  assign n1753 = n1122 & ~n1159 ;
  assign n1754 = ( n1144 & ~n1159 ) | ( n1144 & n1753 ) | ( ~n1159 & n1753 ) ;
  assign n1755 = n1156 | n1754 ;
  assign n1756 = ( n1747 & n1752 ) | ( n1747 & ~n1755 ) | ( n1752 & ~n1755 ) ;
  assign n1757 = ~n1153 & n1163 ;
  assign n1758 = n1168 | n1757 ;
  assign n1759 = ~n1150 & n1758 ;
  assign n1760 = n1173 | n1759 ;
  assign n1761 = ~n1210 & n1760 ;
  assign n1762 = n1201 | n1761 ;
  assign n1763 = n1150 & ~n1173 ;
  assign n1764 = ( ~n1173 & n1176 ) | ( ~n1173 & n1763 ) | ( n1176 & n1763 ) ;
  assign n1765 = n1210 | n1764 ;
  assign n1766 = ~n1201 & n1765 ;
  assign n1767 = ( n1756 & n1762 ) | ( n1756 & ~n1766 ) | ( n1762 & ~n1766 ) ;
  assign n1768 = ~n1192 & n1195 ;
  assign n1769 = n1189 | n1768 ;
  assign n1770 = ~n1186 & n1769 ;
  assign n1771 = n1183 | n1770 ;
  assign n1772 = ~n1230 & n1771 ;
  assign n1773 = n1233 | n1772 ;
  assign n1774 = ~n1189 & n1192 ;
  assign n1775 = ( ~n1189 & n1212 ) | ( ~n1189 & n1774 ) | ( n1212 & n1774 ) ;
  assign n1776 = n1186 | n1775 ;
  assign n1777 = ~n1183 & n1776 ;
  assign n1778 = ( ~n1233 & n1234 ) | ( ~n1233 & n1777 ) | ( n1234 & n1777 ) ;
  assign n1779 = ( n1767 & n1773 ) | ( n1767 & ~n1778 ) | ( n1773 & ~n1778 ) ;
  assign n1780 = n1227 & ~n1238 ;
  assign n1781 = n1224 & ~n1243 ;
  assign n1782 = ( ~n1243 & n1780 ) | ( ~n1243 & n1781 ) | ( n1780 & n1781 ) ;
  assign n1783 = n1250 | n1782 ;
  assign n1784 = ~n1247 & n1783 ;
  assign n1785 = n1221 & ~n1299 ;
  assign n1786 = ( ~n1299 & n1784 ) | ( ~n1299 & n1785 ) | ( n1784 & n1785 ) ;
  assign n1787 = n1279 | n1786 ;
  assign n1788 = ~n1224 & n1238 ;
  assign n1789 = n1243 | n1788 ;
  assign n1790 = ~n1250 & n1789 ;
  assign n1791 = n1247 | n1790 ;
  assign n1792 = ~n1221 & n1791 ;
  assign n1793 = n1299 | n1792 ;
  assign n1794 = ~n1279 & n1793 ;
  assign n1795 = ( n1779 & ~n1787 ) | ( n1779 & n1794 ) | ( ~n1787 & n1794 ) ;
  assign n1796 = ~n1270 & n1273 ;
  assign n1797 = ( ~n1270 & n1287 ) | ( ~n1270 & n1796 ) | ( n1287 & n1796 ) ;
  assign n1798 = n1293 | n1797 ;
  assign n1799 = ~n1267 & n1798 ;
  assign n1800 = n1264 & ~n1330 ;
  assign n1801 = ( ~n1330 & n1799 ) | ( ~n1330 & n1800 ) | ( n1799 & n1800 ) ;
  assign n1802 = n1327 | n1801 ;
  assign n1803 = n1282 & ~n1286 ;
  assign n1804 = n1276 | n1803 ;
  assign n1805 = ~n1273 & n1804 ;
  assign n1806 = n1270 | n1805 ;
  assign n1807 = ~n1293 & n1806 ;
  assign n1808 = n1267 | n1807 ;
  assign n1809 = ~n1264 & n1808 ;
  assign n1810 = ( ~n1327 & n1331 ) | ( ~n1327 & n1809 ) | ( n1331 & n1809 ) ;
  assign n1811 = ( n1795 & ~n1802 ) | ( n1795 & n1810 ) | ( ~n1802 & n1810 ) ;
  assign n1812 = ~n1324 & n1334 ;
  assign n1813 = n1339 | n1812 ;
  assign n1814 = ~n1321 & n1813 ;
  assign n1815 = n1344 | n1814 ;
  assign n1816 = ~n1318 & n1815 ;
  assign n1817 = n1349 | n1816 ;
  assign n1818 = ~n1315 & n1817 ;
  assign n1819 = n1312 & ~n1408 ;
  assign n1820 = ( ~n1408 & n1818 ) | ( ~n1408 & n1819 ) | ( n1818 & n1819 ) ;
  assign n1821 = n1392 | n1820 ;
  assign n1822 = n1321 & ~n1344 ;
  assign n1823 = ( ~n1344 & n1354 ) | ( ~n1344 & n1822 ) | ( n1354 & n1822 ) ;
  assign n1824 = n1318 | n1823 ;
  assign n1825 = ~n1349 & n1824 ;
  assign n1826 = ~n1312 & n1315 ;
  assign n1827 = ( ~n1312 & n1825 ) | ( ~n1312 & n1826 ) | ( n1825 & n1826 ) ;
  assign n1828 = n1408 | n1827 ;
  assign n1829 = ~n1392 & n1828 ;
  assign n1830 = ( n1811 & n1821 ) | ( n1811 & ~n1829 ) | ( n1821 & ~n1829 ) ;
  assign n1831 = ~n1383 & n1386 ;
  assign n1832 = n1380 | n1831 ;
  assign n1833 = ~n1377 & n1832 ;
  assign n1834 = n1374 | n1833 ;
  assign n1835 = ~n1371 & n1834 ;
  assign n1836 = n1402 | n1835 ;
  assign n1837 = ~n1368 & n1836 ;
  assign n1838 = n1365 & ~n1429 ;
  assign n1839 = ( ~n1429 & n1837 ) | ( ~n1429 & n1838 ) | ( n1837 & n1838 ) ;
  assign n1840 = n1432 | n1839 ;
  assign n1841 = ~n1380 & n1383 ;
  assign n1842 = ( ~n1380 & n1410 ) | ( ~n1380 & n1841 ) | ( n1410 & n1841 ) ;
  assign n1843 = n1377 | n1842 ;
  assign n1844 = ~n1374 & n1843 ;
  assign n1845 = n1371 & ~n1402 ;
  assign n1846 = ( ~n1402 & n1844 ) | ( ~n1402 & n1845 ) | ( n1844 & n1845 ) ;
  assign n1847 = n1368 | n1846 ;
  assign n1848 = ~n1365 & n1847 ;
  assign n1849 = ( ~n1432 & n1433 ) | ( ~n1432 & n1848 ) | ( n1433 & n1848 ) ;
  assign n1850 = ( n1830 & n1840 ) | ( n1830 & ~n1849 ) | ( n1840 & ~n1849 ) ;
  assign n1851 = n261 | n1053 ;
  assign n1852 = n1426 & ~n1437 ;
  assign n1853 = n1423 & ~n1442 ;
  assign n1854 = ( ~n1442 & n1852 ) | ( ~n1442 & n1853 ) | ( n1852 & n1853 ) ;
  assign n1855 = n1851 | n1854 ;
  assign n1856 = ~n268 & n1855 ;
  assign n1857 = ~n1423 & n1437 ;
  assign n1858 = n1442 | n1857 ;
  assign n1859 = ~n1851 & n1858 ;
  assign n1860 = n268 | n1859 ;
  assign n1861 = ( n1850 & ~n1856 ) | ( n1850 & n1860 ) | ( ~n1856 & n1860 ) ;
  assign n1862 = n1728 & n1861 ;
  assign n1863 = x134 & ~n661 ;
  assign n1864 = x8 | n672 ;
  assign n1865 = ~n272 & n1864 ;
  assign n1866 = ( ~n289 & n1455 ) | ( ~n289 & n1865 ) | ( n1455 & n1865 ) ;
  assign n1867 = ( n300 & ~n1460 ) | ( n300 & n1866 ) | ( ~n1460 & n1866 ) ;
  assign n1868 = ( ~n319 & n322 ) | ( ~n319 & n1867 ) | ( n322 & n1867 ) ;
  assign n1869 = ( ~n340 & n348 ) | ( ~n340 & n1464 ) | ( n348 & n1464 ) ;
  assign n1870 = n330 | n1869 ;
  assign n1871 = ( n342 & n1868 ) | ( n342 & ~n1870 ) | ( n1868 & ~n1870 ) ;
  assign n1872 = ~n327 & n345 ;
  assign n1873 = n364 | n1872 ;
  assign n1874 = ~n361 & n1873 ;
  assign n1875 = n368 | n1874 ;
  assign n1876 = ~n358 & n1875 ;
  assign n1877 = ( ~n368 & n380 ) | ( ~n368 & n1476 ) | ( n380 & n1476 ) ;
  assign n1878 = n358 | n1877 ;
  assign n1879 = ( n1871 & n1876 ) | ( n1871 & ~n1878 ) | ( n1876 & ~n1878 ) ;
  assign n1880 = ~n355 & n373 ;
  assign n1881 = n378 | n1880 ;
  assign n1882 = ~n415 & n1881 ;
  assign n1883 = n406 | n1882 ;
  assign n1884 = ~n403 & n1883 ;
  assign n1885 = n400 | n1884 ;
  assign n1886 = ( ~n406 & n416 ) | ( ~n406 & n1486 ) | ( n416 & n1486 ) ;
  assign n1887 = n403 | n1886 ;
  assign n1888 = ~n400 & n1887 ;
  assign n1889 = ( n1879 & n1885 ) | ( n1879 & ~n1888 ) | ( n1885 & ~n1888 ) ;
  assign n1890 = ~n391 & n394 ;
  assign n1891 = n388 | n1890 ;
  assign n1892 = ~n435 & n1891 ;
  assign n1893 = n438 | n1892 ;
  assign n1894 = ~n432 & n1893 ;
  assign n1895 = n443 | n1894 ;
  assign n1896 = ( ~n388 & n421 ) | ( ~n388 & n1497 ) | ( n421 & n1497 ) ;
  assign n1897 = n435 | n1896 ;
  assign n1898 = ~n438 & n1897 ;
  assign n1899 = ( ~n443 & n1503 ) | ( ~n443 & n1898 ) | ( n1503 & n1898 ) ;
  assign n1900 = ( n1889 & n1895 ) | ( n1889 & ~n1899 ) | ( n1895 & ~n1899 ) ;
  assign n1901 = ( ~n452 & n456 ) | ( ~n452 & n1504 ) | ( n456 & n1504 ) ;
  assign n1902 = n426 | n1901 ;
  assign n1903 = ~n504 & n1902 ;
  assign n1904 = ( ~n487 & n488 ) | ( ~n487 & n1903 ) | ( n488 & n1903 ) ;
  assign n1905 = n491 | n1904 ;
  assign n1906 = n448 & ~n455 ;
  assign n1907 = n452 | n1906 ;
  assign n1908 = ~n426 & n1907 ;
  assign n1909 = n504 | n1908 ;
  assign n1910 = ~n484 & n1909 ;
  assign n1911 = n487 | n1910 ;
  assign n1912 = ~n491 & n1911 ;
  assign n1913 = ( n1900 & ~n1905 ) | ( n1900 & n1912 ) | ( ~n1905 & n1912 ) ;
  assign n1914 = ( ~n472 & n499 ) | ( ~n472 & n1519 ) | ( n499 & n1519 ) ;
  assign n1915 = n469 | n1914 ;
  assign n1916 = ~n535 & n1915 ;
  assign n1917 = ( ~n539 & n558 ) | ( ~n539 & n1916 ) | ( n558 & n1916 ) ;
  assign n1918 = n529 | n1917 ;
  assign n1919 = ~n478 & n481 ;
  assign n1920 = n475 | n1919 ;
  assign n1921 = ~n498 & n1920 ;
  assign n1922 = n472 | n1921 ;
  assign n1923 = ~n469 & n1922 ;
  assign n1924 = n535 | n1923 ;
  assign n1925 = ~n532 & n1924 ;
  assign n1926 = ( ~n529 & n1535 ) | ( ~n529 & n1925 ) | ( n1535 & n1925 ) ;
  assign n1927 = ( n1913 & ~n1918 ) | ( n1913 & n1926 ) | ( ~n1918 & n1926 ) ;
  assign n1928 = ~n526 & n544 ;
  assign n1929 = n549 | n1928 ;
  assign n1930 = ~n523 & n1929 ;
  assign n1931 = n554 | n1930 ;
  assign n1932 = ~n520 & n1931 ;
  assign n1933 = n517 | n1932 ;
  assign n1934 = ~n613 & n1933 ;
  assign n1935 = ( ~n594 & n598 ) | ( ~n594 & n1934 ) | ( n598 & n1934 ) ;
  assign n1936 = n591 | n1935 ;
  assign n1937 = ( ~n554 & n563 ) | ( ~n554 & n1545 ) | ( n563 & n1545 ) ;
  assign n1938 = n520 | n1937 ;
  assign n1939 = ~n517 & n1938 ;
  assign n1940 = ( ~n597 & n614 ) | ( ~n597 & n1939 ) | ( n614 & n1939 ) ;
  assign n1941 = n594 | n1940 ;
  assign n1942 = ~n591 & n1941 ;
  assign n1943 = ( n1927 & n1936 ) | ( n1927 & ~n1942 ) | ( n1936 & ~n1942 ) ;
  assign n1944 = ~n582 & n585 ;
  assign n1945 = n579 | n1944 ;
  assign n1946 = ~n576 & n1945 ;
  assign n1947 = n607 | n1946 ;
  assign n1948 = ~n573 & n1947 ;
  assign n1949 = n570 | n1948 ;
  assign n1950 = ~n634 & n1949 ;
  assign n1951 = ( ~n631 & n649 ) | ( ~n631 & n1950 ) | ( n649 & n1950 ) ;
  assign n1952 = n642 | n1951 ;
  assign n1953 = ( ~n579 & n619 ) | ( ~n579 & n1564 ) | ( n619 & n1564 ) ;
  assign n1954 = n576 | n1953 ;
  assign n1955 = ~n607 & n1954 ;
  assign n1956 = ( ~n570 & n623 ) | ( ~n570 & n1955 ) | ( n623 & n1955 ) ;
  assign n1957 = n634 | n1956 ;
  assign n1958 = ~n637 & n1957 ;
  assign n1959 = ( ~n642 & n1576 ) | ( ~n642 & n1958 ) | ( n1576 & n1958 ) ;
  assign n1960 = ( n1943 & n1952 ) | ( n1943 & ~n1959 ) | ( n1952 & ~n1959 ) ;
  assign n1961 = n659 | n1450 ;
  assign n1962 = n1575 & ~n1581 ;
  assign n1963 = ( n1577 & ~n1581 ) | ( n1577 & n1962 ) | ( ~n1581 & n1962 ) ;
  assign n1964 = n1961 | n1963 ;
  assign n1965 = ~n666 & n1964 ;
  assign n1966 = n647 & ~n1575 ;
  assign n1967 = n1581 | n1966 ;
  assign n1968 = ~n1961 & n1967 ;
  assign n1969 = n666 | n1968 ;
  assign n1970 = ( n1960 & ~n1965 ) | ( n1960 & n1969 ) | ( ~n1965 & n1969 ) ;
  assign n1971 = n1863 & n1970 ;
  assign n1972 = x135 & ~n1058 ;
  assign n1973 = x9 | n1069 ;
  assign n1974 = ~n670 & n1973 ;
  assign n1975 = ( ~n687 & n1594 ) | ( ~n687 & n1974 ) | ( n1594 & n1974 ) ;
  assign n1976 = ( n698 & ~n1599 ) | ( n698 & n1975 ) | ( ~n1599 & n1975 ) ;
  assign n1977 = ( ~n717 & n720 ) | ( ~n717 & n1976 ) | ( n720 & n1976 ) ;
  assign n1978 = ( ~n738 & n746 ) | ( ~n738 & n1603 ) | ( n746 & n1603 ) ;
  assign n1979 = n728 | n1978 ;
  assign n1980 = ( n740 & n1977 ) | ( n740 & ~n1979 ) | ( n1977 & ~n1979 ) ;
  assign n1981 = ~n725 & n743 ;
  assign n1982 = n762 | n1981 ;
  assign n1983 = ~n759 & n1982 ;
  assign n1984 = n766 | n1983 ;
  assign n1985 = ~n756 & n1984 ;
  assign n1986 = ( ~n766 & n778 ) | ( ~n766 & n1615 ) | ( n778 & n1615 ) ;
  assign n1987 = n756 | n1986 ;
  assign n1988 = ( n1980 & n1985 ) | ( n1980 & ~n1987 ) | ( n1985 & ~n1987 ) ;
  assign n1989 = ~n753 & n771 ;
  assign n1990 = n776 | n1989 ;
  assign n1991 = ~n813 & n1990 ;
  assign n1992 = n804 | n1991 ;
  assign n1993 = ~n801 & n1992 ;
  assign n1994 = n798 | n1993 ;
  assign n1995 = ( ~n804 & n814 ) | ( ~n804 & n1625 ) | ( n814 & n1625 ) ;
  assign n1996 = n801 | n1995 ;
  assign n1997 = ~n798 & n1996 ;
  assign n1998 = ( n1988 & n1994 ) | ( n1988 & ~n1997 ) | ( n1994 & ~n1997 ) ;
  assign n1999 = ~n789 & n792 ;
  assign n2000 = n786 | n1999 ;
  assign n2001 = ~n833 & n2000 ;
  assign n2002 = n836 | n2001 ;
  assign n2003 = ~n830 & n2002 ;
  assign n2004 = n841 | n2003 ;
  assign n2005 = ( ~n786 & n819 ) | ( ~n786 & n1636 ) | ( n819 & n1636 ) ;
  assign n2006 = n833 | n2005 ;
  assign n2007 = ~n836 & n2006 ;
  assign n2008 = ( ~n841 & n1642 ) | ( ~n841 & n2007 ) | ( n1642 & n2007 ) ;
  assign n2009 = ( n1998 & n2004 ) | ( n1998 & ~n2008 ) | ( n2004 & ~n2008 ) ;
  assign n2010 = ( ~n850 & n854 ) | ( ~n850 & n1643 ) | ( n854 & n1643 ) ;
  assign n2011 = n824 | n2010 ;
  assign n2012 = ~n902 & n2011 ;
  assign n2013 = ( ~n885 & n886 ) | ( ~n885 & n2012 ) | ( n886 & n2012 ) ;
  assign n2014 = n889 | n2013 ;
  assign n2015 = n846 & ~n853 ;
  assign n2016 = n850 | n2015 ;
  assign n2017 = ~n824 & n2016 ;
  assign n2018 = n902 | n2017 ;
  assign n2019 = ~n882 & n2018 ;
  assign n2020 = n885 | n2019 ;
  assign n2021 = ~n889 & n2020 ;
  assign n2022 = ( n2009 & ~n2014 ) | ( n2009 & n2021 ) | ( ~n2014 & n2021 ) ;
  assign n2023 = ( ~n870 & n897 ) | ( ~n870 & n1658 ) | ( n897 & n1658 ) ;
  assign n2024 = n867 | n2023 ;
  assign n2025 = ~n933 & n2024 ;
  assign n2026 = ( ~n937 & n956 ) | ( ~n937 & n2025 ) | ( n956 & n2025 ) ;
  assign n2027 = n927 | n2026 ;
  assign n2028 = ~n876 & n879 ;
  assign n2029 = n873 | n2028 ;
  assign n2030 = ~n896 & n2029 ;
  assign n2031 = n870 | n2030 ;
  assign n2032 = ~n867 & n2031 ;
  assign n2033 = n933 | n2032 ;
  assign n2034 = ~n930 & n2033 ;
  assign n2035 = ( ~n927 & n1674 ) | ( ~n927 & n2034 ) | ( n1674 & n2034 ) ;
  assign n2036 = ( n2022 & ~n2027 ) | ( n2022 & n2035 ) | ( ~n2027 & n2035 ) ;
  assign n2037 = ~n924 & n942 ;
  assign n2038 = n947 | n2037 ;
  assign n2039 = ~n921 & n2038 ;
  assign n2040 = n952 | n2039 ;
  assign n2041 = ~n918 & n2040 ;
  assign n2042 = n915 | n2041 ;
  assign n2043 = ~n1011 & n2042 ;
  assign n2044 = ( ~n992 & n996 ) | ( ~n992 & n2043 ) | ( n996 & n2043 ) ;
  assign n2045 = n989 | n2044 ;
  assign n2046 = ( ~n952 & n961 ) | ( ~n952 & n1684 ) | ( n961 & n1684 ) ;
  assign n2047 = n918 | n2046 ;
  assign n2048 = ~n915 & n2047 ;
  assign n2049 = ( ~n995 & n1012 ) | ( ~n995 & n2048 ) | ( n1012 & n2048 ) ;
  assign n2050 = n992 | n2049 ;
  assign n2051 = ~n989 & n2050 ;
  assign n2052 = ( n2036 & n2045 ) | ( n2036 & ~n2051 ) | ( n2045 & ~n2051 ) ;
  assign n2053 = ~n980 & n983 ;
  assign n2054 = n977 | n2053 ;
  assign n2055 = ~n974 & n2054 ;
  assign n2056 = n1005 | n2055 ;
  assign n2057 = ~n971 & n2056 ;
  assign n2058 = n968 | n2057 ;
  assign n2059 = ~n1032 & n2058 ;
  assign n2060 = ( ~n1029 & n1047 ) | ( ~n1029 & n2059 ) | ( n1047 & n2059 ) ;
  assign n2061 = n1040 | n2060 ;
  assign n2062 = ( ~n977 & n1017 ) | ( ~n977 & n1703 ) | ( n1017 & n1703 ) ;
  assign n2063 = n974 | n2062 ;
  assign n2064 = ~n1005 & n2063 ;
  assign n2065 = ( ~n968 & n1021 ) | ( ~n968 & n2064 ) | ( n1021 & n2064 ) ;
  assign n2066 = n1032 | n2065 ;
  assign n2067 = ~n1035 & n2066 ;
  assign n2068 = ( ~n1040 & n1715 ) | ( ~n1040 & n2067 ) | ( n1715 & n2067 ) ;
  assign n2069 = ( n2052 & n2061 ) | ( n2052 & ~n2068 ) | ( n2061 & ~n2068 ) ;
  assign n2070 = n1056 | n1589 ;
  assign n2071 = n1714 & ~n1720 ;
  assign n2072 = ( n1716 & ~n1720 ) | ( n1716 & n2071 ) | ( ~n1720 & n2071 ) ;
  assign n2073 = n2070 | n2072 ;
  assign n2074 = ~n1063 & n2073 ;
  assign n2075 = n1045 & ~n1714 ;
  assign n2076 = n1720 | n2075 ;
  assign n2077 = ~n2070 & n2076 ;
  assign n2078 = n1063 | n2077 ;
  assign n2079 = ( n2069 & ~n2074 ) | ( n2069 & n2078 ) | ( ~n2074 & n2078 ) ;
  assign n2080 = n1972 & n2079 ;
  assign n2081 = x136 & ~n271 ;
  assign n2082 = x10 | n278 ;
  assign n2083 = ~n1067 & n2082 ;
  assign n2084 = ( ~n1084 & n1732 ) | ( ~n1084 & n2083 ) | ( n1732 & n2083 ) ;
  assign n2085 = ( n1095 & ~n1737 ) | ( n1095 & n2084 ) | ( ~n1737 & n2084 ) ;
  assign n2086 = ( ~n1114 & n1117 ) | ( ~n1114 & n2085 ) | ( n1117 & n2085 ) ;
  assign n2087 = ( ~n1135 & n1143 ) | ( ~n1135 & n1741 ) | ( n1143 & n1741 ) ;
  assign n2088 = n1125 | n2087 ;
  assign n2089 = ( n1137 & n2086 ) | ( n1137 & ~n2088 ) | ( n2086 & ~n2088 ) ;
  assign n2090 = ~n1122 & n1140 ;
  assign n2091 = n1159 | n2090 ;
  assign n2092 = ~n1156 & n2091 ;
  assign n2093 = n1163 | n2092 ;
  assign n2094 = ~n1153 & n2093 ;
  assign n2095 = ( ~n1163 & n1175 ) | ( ~n1163 & n1753 ) | ( n1175 & n1753 ) ;
  assign n2096 = n1153 | n2095 ;
  assign n2097 = ( n2089 & n2094 ) | ( n2089 & ~n2096 ) | ( n2094 & ~n2096 ) ;
  assign n2098 = ~n1150 & n1168 ;
  assign n2099 = n1173 | n2098 ;
  assign n2100 = ~n1210 & n2099 ;
  assign n2101 = n1201 | n2100 ;
  assign n2102 = ~n1198 & n2101 ;
  assign n2103 = n1195 | n2102 ;
  assign n2104 = ( ~n1201 & n1211 ) | ( ~n1201 & n1763 ) | ( n1211 & n1763 ) ;
  assign n2105 = n1198 | n2104 ;
  assign n2106 = ~n1195 & n2105 ;
  assign n2107 = ( n2097 & n2103 ) | ( n2097 & ~n2106 ) | ( n2103 & ~n2106 ) ;
  assign n2108 = ~n1186 & n1189 ;
  assign n2109 = n1183 | n2108 ;
  assign n2110 = ~n1230 & n2109 ;
  assign n2111 = n1233 | n2110 ;
  assign n2112 = ~n1227 & n2111 ;
  assign n2113 = n1238 | n2112 ;
  assign n2114 = ( ~n1183 & n1216 ) | ( ~n1183 & n1774 ) | ( n1216 & n1774 ) ;
  assign n2115 = n1230 | n2114 ;
  assign n2116 = ~n1233 & n2115 ;
  assign n2117 = ( ~n1238 & n1780 ) | ( ~n1238 & n2116 ) | ( n1780 & n2116 ) ;
  assign n2118 = ( n2107 & n2113 ) | ( n2107 & ~n2117 ) | ( n2113 & ~n2117 ) ;
  assign n2119 = ( ~n1247 & n1251 ) | ( ~n1247 & n1781 ) | ( n1251 & n1781 ) ;
  assign n2120 = n1221 | n2119 ;
  assign n2121 = ~n1299 & n2120 ;
  assign n2122 = ( ~n1282 & n1283 ) | ( ~n1282 & n2121 ) | ( n1283 & n2121 ) ;
  assign n2123 = n1286 | n2122 ;
  assign n2124 = n1243 & ~n1250 ;
  assign n2125 = n1247 | n2124 ;
  assign n2126 = ~n1221 & n2125 ;
  assign n2127 = n1299 | n2126 ;
  assign n2128 = ~n1279 & n2127 ;
  assign n2129 = n1282 | n2128 ;
  assign n2130 = ~n1286 & n2129 ;
  assign n2131 = ( n2118 & ~n2123 ) | ( n2118 & n2130 ) | ( ~n2123 & n2130 ) ;
  assign n2132 = ( ~n1267 & n1294 ) | ( ~n1267 & n1796 ) | ( n1294 & n1796 ) ;
  assign n2133 = n1264 | n2132 ;
  assign n2134 = ~n1330 & n2133 ;
  assign n2135 = ( ~n1334 & n1353 ) | ( ~n1334 & n2134 ) | ( n1353 & n2134 ) ;
  assign n2136 = n1324 | n2135 ;
  assign n2137 = ~n1273 & n1276 ;
  assign n2138 = n1270 | n2137 ;
  assign n2139 = ~n1293 & n2138 ;
  assign n2140 = n1267 | n2139 ;
  assign n2141 = ~n1264 & n2140 ;
  assign n2142 = n1330 | n2141 ;
  assign n2143 = ~n1327 & n2142 ;
  assign n2144 = ( ~n1324 & n1812 ) | ( ~n1324 & n2143 ) | ( n1812 & n2143 ) ;
  assign n2145 = ( n2131 & ~n2136 ) | ( n2131 & n2144 ) | ( ~n2136 & n2144 ) ;
  assign n2146 = ~n1321 & n1339 ;
  assign n2147 = n1344 | n2146 ;
  assign n2148 = ~n1318 & n2147 ;
  assign n2149 = n1349 | n2148 ;
  assign n2150 = ~n1315 & n2149 ;
  assign n2151 = n1312 | n2150 ;
  assign n2152 = ~n1408 & n2151 ;
  assign n2153 = ( ~n1389 & n1393 ) | ( ~n1389 & n2152 ) | ( n1393 & n2152 ) ;
  assign n2154 = n1386 | n2153 ;
  assign n2155 = ( ~n1349 & n1358 ) | ( ~n1349 & n1822 ) | ( n1358 & n1822 ) ;
  assign n2156 = n1315 | n2155 ;
  assign n2157 = ~n1312 & n2156 ;
  assign n2158 = ( ~n1392 & n1409 ) | ( ~n1392 & n2157 ) | ( n1409 & n2157 ) ;
  assign n2159 = n1389 | n2158 ;
  assign n2160 = ~n1386 & n2159 ;
  assign n2161 = ( n2145 & n2154 ) | ( n2145 & ~n2160 ) | ( n2154 & ~n2160 ) ;
  assign n2162 = ~n1377 & n1380 ;
  assign n2163 = n1374 | n2162 ;
  assign n2164 = ~n1371 & n2163 ;
  assign n2165 = n1402 | n2164 ;
  assign n2166 = ~n1368 & n2165 ;
  assign n2167 = n1365 | n2166 ;
  assign n2168 = ~n1429 & n2167 ;
  assign n2169 = ( ~n1426 & n1444 ) | ( ~n1426 & n2168 ) | ( n1444 & n2168 ) ;
  assign n2170 = n1437 | n2169 ;
  assign n2171 = ( ~n1374 & n1414 ) | ( ~n1374 & n1841 ) | ( n1414 & n1841 ) ;
  assign n2172 = n1371 | n2171 ;
  assign n2173 = ~n1402 & n2172 ;
  assign n2174 = ( ~n1365 & n1418 ) | ( ~n1365 & n2173 ) | ( n1418 & n2173 ) ;
  assign n2175 = n1429 | n2174 ;
  assign n2176 = ~n1432 & n2175 ;
  assign n2177 = ( ~n1437 & n1852 ) | ( ~n1437 & n2176 ) | ( n1852 & n2176 ) ;
  assign n2178 = ( n2161 & n2170 ) | ( n2161 & ~n2177 ) | ( n2170 & ~n2177 ) ;
  assign n2179 = ~n268 & n1851 ;
  assign n2180 = ( ~n268 & n1853 ) | ( ~n268 & n2179 ) | ( n1853 & n2179 ) ;
  assign n2181 = n265 | n2180 ;
  assign n2182 = ~n276 & n2181 ;
  assign n2183 = n1442 & ~n1851 ;
  assign n2184 = n268 | n2183 ;
  assign n2185 = ~n265 & n2184 ;
  assign n2186 = n276 | n2185 ;
  assign n2187 = ( n2178 & ~n2182 ) | ( n2178 & n2186 ) | ( ~n2182 & n2186 ) ;
  assign n2188 = n2081 & n2187 ;
  assign n2189 = x137 & ~n669 ;
  assign n2190 = x11 | n676 ;
  assign n2191 = ~n288 & n2190 ;
  assign n2192 = ( ~n286 & n299 ) | ( ~n286 & n2191 ) | ( n299 & n2191 ) ;
  assign n2193 = ( ~n314 & n1459 ) | ( ~n314 & n2192 ) | ( n1459 & n2192 ) ;
  assign n2194 = ( ~n1465 & n1468 ) | ( ~n1465 & n2193 ) | ( n1468 & n2193 ) ;
  assign n2195 = ( ~n351 & n1473 ) | ( ~n351 & n2194 ) | ( n1473 & n2194 ) ;
  assign n2196 = ( n375 & ~n383 ) | ( n375 & n2195 ) | ( ~n383 & n2195 ) ;
  assign n2197 = n378 & ~n415 ;
  assign n2198 = n406 | n2197 ;
  assign n2199 = ~n403 & n2198 ;
  assign n2200 = n400 | n2199 ;
  assign n2201 = ~n397 & n2200 ;
  assign n2202 = n394 | n2201 ;
  assign n2203 = ( ~n420 & n2196 ) | ( ~n420 & n2202 ) | ( n2196 & n2202 ) ;
  assign n2204 = n388 & ~n435 ;
  assign n2205 = n438 | n2204 ;
  assign n2206 = ~n432 & n2205 ;
  assign n2207 = n443 | n2206 ;
  assign n2208 = ~n429 & n2207 ;
  assign n2209 = n448 | n2208 ;
  assign n2210 = ( n421 & ~n438 ) | ( n421 & n439 ) | ( ~n438 & n439 ) ;
  assign n2211 = n432 | n2210 ;
  assign n2212 = ~n443 & n2211 ;
  assign n2213 = ( ~n448 & n1504 ) | ( ~n448 & n2212 ) | ( n1504 & n2212 ) ;
  assign n2214 = ( n2203 & n2209 ) | ( n2203 & ~n2213 ) | ( n2209 & ~n2213 ) ;
  assign n2215 = ( n456 & ~n504 ) | ( n456 & n1508 ) | ( ~n504 & n1508 ) ;
  assign n2216 = n484 | n2215 ;
  assign n2217 = ~n487 & n2216 ;
  assign n2218 = ( ~n481 & n492 ) | ( ~n481 & n2217 ) | ( n492 & n2217 ) ;
  assign n2219 = n478 | n2218 ;
  assign n2220 = ~n426 & n452 ;
  assign n2221 = n504 | n2220 ;
  assign n2222 = ~n484 & n2221 ;
  assign n2223 = n487 | n2222 ;
  assign n2224 = ~n491 & n2223 ;
  assign n2225 = n481 | n2224 ;
  assign n2226 = ~n478 & n2225 ;
  assign n2227 = ( n2214 & ~n2219 ) | ( n2214 & n2226 ) | ( ~n2219 & n2226 ) ;
  assign n2228 = ( n499 & ~n535 ) | ( n499 & n1523 ) | ( ~n535 & n1523 ) ;
  assign n2229 = n532 | n2228 ;
  assign n2230 = ~n539 & n2229 ;
  assign n2231 = ( ~n544 & n559 ) | ( ~n544 & n2230 ) | ( n559 & n2230 ) ;
  assign n2232 = n526 | n2231 ;
  assign n2233 = n475 & ~n498 ;
  assign n2234 = n472 | n2233 ;
  assign n2235 = ~n469 & n2234 ;
  assign n2236 = n535 | n2235 ;
  assign n2237 = ~n532 & n2236 ;
  assign n2238 = n539 | n2237 ;
  assign n2239 = ~n529 & n2238 ;
  assign n2240 = ( ~n526 & n1928 ) | ( ~n526 & n2239 ) | ( n1928 & n2239 ) ;
  assign n2241 = ( n2227 & ~n2232 ) | ( n2227 & n2240 ) | ( ~n2232 & n2240 ) ;
  assign n2242 = ~n523 & n549 ;
  assign n2243 = n554 | n2242 ;
  assign n2244 = ~n520 & n2243 ;
  assign n2245 = n517 | n2244 ;
  assign n2246 = ~n613 & n2245 ;
  assign n2247 = n597 | n2246 ;
  assign n2248 = ~n594 & n2247 ;
  assign n2249 = ( ~n588 & n1554 ) | ( ~n588 & n2248 ) | ( n1554 & n2248 ) ;
  assign n2250 = n585 | n2249 ;
  assign n2251 = ( ~n517 & n563 ) | ( ~n517 & n1549 ) | ( n563 & n1549 ) ;
  assign n2252 = n613 | n2251 ;
  assign n2253 = ~n597 & n2252 ;
  assign n2254 = ( ~n591 & n615 ) | ( ~n591 & n2253 ) | ( n615 & n2253 ) ;
  assign n2255 = n588 | n2254 ;
  assign n2256 = ~n585 & n2255 ;
  assign n2257 = ( n2241 & n2250 ) | ( n2241 & ~n2256 ) | ( n2250 & ~n2256 ) ;
  assign n2258 = ~n576 & n579 ;
  assign n2259 = n607 | n2258 ;
  assign n2260 = ~n573 & n2259 ;
  assign n2261 = n570 | n2260 ;
  assign n2262 = ~n634 & n2261 ;
  assign n2263 = n637 | n2262 ;
  assign n2264 = ~n631 & n2263 ;
  assign n2265 = ( ~n628 & n1583 ) | ( ~n628 & n2264 ) | ( n1583 & n2264 ) ;
  assign n2266 = n647 | n2265 ;
  assign n2267 = ( ~n607 & n619 ) | ( ~n607 & n1568 ) | ( n619 & n1568 ) ;
  assign n2268 = n573 | n2267 ;
  assign n2269 = ~n570 & n2268 ;
  assign n2270 = ( ~n637 & n638 ) | ( ~n637 & n2269 ) | ( n638 & n2269 ) ;
  assign n2271 = n631 | n2270 ;
  assign n2272 = ~n642 & n2271 ;
  assign n2273 = ( ~n647 & n1577 ) | ( ~n647 & n2272 ) | ( n1577 & n2272 ) ;
  assign n2274 = ( n2257 & n2266 ) | ( n2257 & ~n2273 ) | ( n2266 & ~n2273 ) ;
  assign n2275 = ~n666 & n1961 ;
  assign n2276 = ( ~n666 & n1962 ) | ( ~n666 & n2275 ) | ( n1962 & n2275 ) ;
  assign n2277 = n663 | n2276 ;
  assign n2278 = ~n674 & n2277 ;
  assign n2279 = n1581 & ~n1961 ;
  assign n2280 = n666 | n2279 ;
  assign n2281 = ~n663 & n2280 ;
  assign n2282 = n674 | n2281 ;
  assign n2283 = ( n2274 & ~n2278 ) | ( n2274 & n2282 ) | ( ~n2278 & n2282 ) ;
  assign n2284 = n2189 & n2283 ;
  assign n2285 = x138 & ~n1066 ;
  assign n2286 = x12 | n1073 ;
  assign n2287 = ~n686 & n2286 ;
  assign n2288 = ( ~n684 & n697 ) | ( ~n684 & n2287 ) | ( n697 & n2287 ) ;
  assign n2289 = ( ~n712 & n1598 ) | ( ~n712 & n2288 ) | ( n1598 & n2288 ) ;
  assign n2290 = ( ~n1604 & n1607 ) | ( ~n1604 & n2289 ) | ( n1607 & n2289 ) ;
  assign n2291 = ( ~n749 & n1612 ) | ( ~n749 & n2290 ) | ( n1612 & n2290 ) ;
  assign n2292 = ( n773 & ~n781 ) | ( n773 & n2291 ) | ( ~n781 & n2291 ) ;
  assign n2293 = n776 & ~n813 ;
  assign n2294 = n804 | n2293 ;
  assign n2295 = ~n801 & n2294 ;
  assign n2296 = n798 | n2295 ;
  assign n2297 = ~n795 & n2296 ;
  assign n2298 = n792 | n2297 ;
  assign n2299 = ( ~n818 & n2292 ) | ( ~n818 & n2298 ) | ( n2292 & n2298 ) ;
  assign n2300 = n786 & ~n833 ;
  assign n2301 = n836 | n2300 ;
  assign n2302 = ~n830 & n2301 ;
  assign n2303 = n841 | n2302 ;
  assign n2304 = ~n827 & n2303 ;
  assign n2305 = n846 | n2304 ;
  assign n2306 = ( n819 & ~n836 ) | ( n819 & n837 ) | ( ~n836 & n837 ) ;
  assign n2307 = n830 | n2306 ;
  assign n2308 = ~n841 & n2307 ;
  assign n2309 = ( ~n846 & n1643 ) | ( ~n846 & n2308 ) | ( n1643 & n2308 ) ;
  assign n2310 = ( n2299 & n2305 ) | ( n2299 & ~n2309 ) | ( n2305 & ~n2309 ) ;
  assign n2311 = ( n854 & ~n902 ) | ( n854 & n1647 ) | ( ~n902 & n1647 ) ;
  assign n2312 = n882 | n2311 ;
  assign n2313 = ~n885 & n2312 ;
  assign n2314 = ( ~n879 & n890 ) | ( ~n879 & n2313 ) | ( n890 & n2313 ) ;
  assign n2315 = n876 | n2314 ;
  assign n2316 = ~n824 & n850 ;
  assign n2317 = n902 | n2316 ;
  assign n2318 = ~n882 & n2317 ;
  assign n2319 = n885 | n2318 ;
  assign n2320 = ~n889 & n2319 ;
  assign n2321 = n879 | n2320 ;
  assign n2322 = ~n876 & n2321 ;
  assign n2323 = ( n2310 & ~n2315 ) | ( n2310 & n2322 ) | ( ~n2315 & n2322 ) ;
  assign n2324 = ( n897 & ~n933 ) | ( n897 & n1662 ) | ( ~n933 & n1662 ) ;
  assign n2325 = n930 | n2324 ;
  assign n2326 = ~n937 & n2325 ;
  assign n2327 = ( ~n942 & n957 ) | ( ~n942 & n2326 ) | ( n957 & n2326 ) ;
  assign n2328 = n924 | n2327 ;
  assign n2329 = n873 & ~n896 ;
  assign n2330 = n870 | n2329 ;
  assign n2331 = ~n867 & n2330 ;
  assign n2332 = n933 | n2331 ;
  assign n2333 = ~n930 & n2332 ;
  assign n2334 = n937 | n2333 ;
  assign n2335 = ~n927 & n2334 ;
  assign n2336 = ( ~n924 & n2037 ) | ( ~n924 & n2335 ) | ( n2037 & n2335 ) ;
  assign n2337 = ( n2323 & ~n2328 ) | ( n2323 & n2336 ) | ( ~n2328 & n2336 ) ;
  assign n2338 = ~n921 & n947 ;
  assign n2339 = n952 | n2338 ;
  assign n2340 = ~n918 & n2339 ;
  assign n2341 = n915 | n2340 ;
  assign n2342 = ~n1011 & n2341 ;
  assign n2343 = n995 | n2342 ;
  assign n2344 = ~n992 & n2343 ;
  assign n2345 = ( ~n986 & n1693 ) | ( ~n986 & n2344 ) | ( n1693 & n2344 ) ;
  assign n2346 = n983 | n2345 ;
  assign n2347 = ( ~n915 & n961 ) | ( ~n915 & n1688 ) | ( n961 & n1688 ) ;
  assign n2348 = n1011 | n2347 ;
  assign n2349 = ~n995 & n2348 ;
  assign n2350 = ( ~n989 & n1013 ) | ( ~n989 & n2349 ) | ( n1013 & n2349 ) ;
  assign n2351 = n986 | n2350 ;
  assign n2352 = ~n983 & n2351 ;
  assign n2353 = ( n2337 & n2346 ) | ( n2337 & ~n2352 ) | ( n2346 & ~n2352 ) ;
  assign n2354 = ~n974 & n977 ;
  assign n2355 = n1005 | n2354 ;
  assign n2356 = ~n971 & n2355 ;
  assign n2357 = n968 | n2356 ;
  assign n2358 = ~n1032 & n2357 ;
  assign n2359 = n1035 | n2358 ;
  assign n2360 = ~n1029 & n2359 ;
  assign n2361 = ( ~n1026 & n1722 ) | ( ~n1026 & n2360 ) | ( n1722 & n2360 ) ;
  assign n2362 = n1045 | n2361 ;
  assign n2363 = ( ~n1005 & n1017 ) | ( ~n1005 & n1707 ) | ( n1017 & n1707 ) ;
  assign n2364 = n971 | n2363 ;
  assign n2365 = ~n968 & n2364 ;
  assign n2366 = ( ~n1035 & n1036 ) | ( ~n1035 & n2365 ) | ( n1036 & n2365 ) ;
  assign n2367 = n1029 | n2366 ;
  assign n2368 = ~n1040 & n2367 ;
  assign n2369 = ( ~n1045 & n1716 ) | ( ~n1045 & n2368 ) | ( n1716 & n2368 ) ;
  assign n2370 = ( n2353 & n2362 ) | ( n2353 & ~n2369 ) | ( n2362 & ~n2369 ) ;
  assign n2371 = ~n1063 & n2070 ;
  assign n2372 = ( ~n1063 & n2071 ) | ( ~n1063 & n2371 ) | ( n2071 & n2371 ) ;
  assign n2373 = n1060 | n2372 ;
  assign n2374 = ~n1071 & n2373 ;
  assign n2375 = n1720 & ~n2070 ;
  assign n2376 = n1063 | n2375 ;
  assign n2377 = ~n1060 & n2376 ;
  assign n2378 = n1071 | n2377 ;
  assign n2379 = ( n2370 & ~n2374 ) | ( n2370 & n2378 ) | ( ~n2374 & n2378 ) ;
  assign n2380 = n2285 & n2379 ;
  assign n2381 = x139 & ~n287 ;
  assign n2382 = x13 | n290 ;
  assign n2383 = ~n1083 & n2382 ;
  assign n2384 = ( ~n1081 & n1094 ) | ( ~n1081 & n2383 ) | ( n1094 & n2383 ) ;
  assign n2385 = ( ~n1109 & n1736 ) | ( ~n1109 & n2384 ) | ( n1736 & n2384 ) ;
  assign n2386 = ( ~n1742 & n1745 ) | ( ~n1742 & n2385 ) | ( n1745 & n2385 ) ;
  assign n2387 = ( ~n1146 & n1750 ) | ( ~n1146 & n2386 ) | ( n1750 & n2386 ) ;
  assign n2388 = ( n1170 & ~n1178 ) | ( n1170 & n2387 ) | ( ~n1178 & n2387 ) ;
  assign n2389 = n1173 & ~n1210 ;
  assign n2390 = n1201 | n2389 ;
  assign n2391 = ~n1198 & n2390 ;
  assign n2392 = n1195 | n2391 ;
  assign n2393 = ~n1192 & n2392 ;
  assign n2394 = n1189 | n2393 ;
  assign n2395 = ( ~n1215 & n2388 ) | ( ~n1215 & n2394 ) | ( n2388 & n2394 ) ;
  assign n2396 = n1183 & ~n1230 ;
  assign n2397 = n1233 | n2396 ;
  assign n2398 = ~n1227 & n2397 ;
  assign n2399 = n1238 | n2398 ;
  assign n2400 = ~n1224 & n2399 ;
  assign n2401 = n1243 | n2400 ;
  assign n2402 = ( n1216 & ~n1233 ) | ( n1216 & n1234 ) | ( ~n1233 & n1234 ) ;
  assign n2403 = n1227 | n2402 ;
  assign n2404 = ~n1238 & n2403 ;
  assign n2405 = ( ~n1243 & n1781 ) | ( ~n1243 & n2404 ) | ( n1781 & n2404 ) ;
  assign n2406 = ( n2395 & n2401 ) | ( n2395 & ~n2405 ) | ( n2401 & ~n2405 ) ;
  assign n2407 = ( n1251 & ~n1299 ) | ( n1251 & n1785 ) | ( ~n1299 & n1785 ) ;
  assign n2408 = n1279 | n2407 ;
  assign n2409 = ~n1282 & n2408 ;
  assign n2410 = ( ~n1276 & n1287 ) | ( ~n1276 & n2409 ) | ( n1287 & n2409 ) ;
  assign n2411 = n1273 | n2410 ;
  assign n2412 = ~n1221 & n1247 ;
  assign n2413 = n1299 | n2412 ;
  assign n2414 = ~n1279 & n2413 ;
  assign n2415 = n1282 | n2414 ;
  assign n2416 = ~n1286 & n2415 ;
  assign n2417 = n1276 | n2416 ;
  assign n2418 = ~n1273 & n2417 ;
  assign n2419 = ( n2406 & ~n2411 ) | ( n2406 & n2418 ) | ( ~n2411 & n2418 ) ;
  assign n2420 = ( n1294 & ~n1330 ) | ( n1294 & n1800 ) | ( ~n1330 & n1800 ) ;
  assign n2421 = n1327 | n2420 ;
  assign n2422 = ~n1334 & n2421 ;
  assign n2423 = ( ~n1339 & n1354 ) | ( ~n1339 & n2422 ) | ( n1354 & n2422 ) ;
  assign n2424 = n1321 | n2423 ;
  assign n2425 = n1270 & ~n1293 ;
  assign n2426 = n1267 | n2425 ;
  assign n2427 = ~n1264 & n2426 ;
  assign n2428 = n1330 | n2427 ;
  assign n2429 = ~n1327 & n2428 ;
  assign n2430 = n1334 | n2429 ;
  assign n2431 = ~n1324 & n2430 ;
  assign n2432 = ( ~n1321 & n2146 ) | ( ~n1321 & n2431 ) | ( n2146 & n2431 ) ;
  assign n2433 = ( n2419 & ~n2424 ) | ( n2419 & n2432 ) | ( ~n2424 & n2432 ) ;
  assign n2434 = ~n1318 & n1344 ;
  assign n2435 = n1349 | n2434 ;
  assign n2436 = ~n1315 & n2435 ;
  assign n2437 = n1312 | n2436 ;
  assign n2438 = ~n1408 & n2437 ;
  assign n2439 = n1392 | n2438 ;
  assign n2440 = ~n1389 & n2439 ;
  assign n2441 = ( ~n1383 & n1831 ) | ( ~n1383 & n2440 ) | ( n1831 & n2440 ) ;
  assign n2442 = n1380 | n2441 ;
  assign n2443 = ( ~n1312 & n1358 ) | ( ~n1312 & n1826 ) | ( n1358 & n1826 ) ;
  assign n2444 = n1408 | n2443 ;
  assign n2445 = ~n1392 & n2444 ;
  assign n2446 = ( ~n1386 & n1410 ) | ( ~n1386 & n2445 ) | ( n1410 & n2445 ) ;
  assign n2447 = n1383 | n2446 ;
  assign n2448 = ~n1380 & n2447 ;
  assign n2449 = ( n2433 & n2442 ) | ( n2433 & ~n2448 ) | ( n2442 & ~n2448 ) ;
  assign n2450 = ~n1371 & n1374 ;
  assign n2451 = n1402 | n2450 ;
  assign n2452 = ~n1368 & n2451 ;
  assign n2453 = n1365 | n2452 ;
  assign n2454 = ~n1429 & n2453 ;
  assign n2455 = n1432 | n2454 ;
  assign n2456 = ~n1426 & n2455 ;
  assign n2457 = ( ~n1423 & n1857 ) | ( ~n1423 & n2456 ) | ( n1857 & n2456 ) ;
  assign n2458 = n1442 | n2457 ;
  assign n2459 = ( ~n1402 & n1414 ) | ( ~n1402 & n1845 ) | ( n1414 & n1845 ) ;
  assign n2460 = n1368 | n2459 ;
  assign n2461 = ~n1365 & n2460 ;
  assign n2462 = ( ~n1432 & n1433 ) | ( ~n1432 & n2461 ) | ( n1433 & n2461 ) ;
  assign n2463 = n1426 | n2462 ;
  assign n2464 = ~n1437 & n2463 ;
  assign n2465 = ( ~n1442 & n1853 ) | ( ~n1442 & n2464 ) | ( n1853 & n2464 ) ;
  assign n2466 = ( n2449 & n2458 ) | ( n2449 & ~n2465 ) | ( n2458 & ~n2465 ) ;
  assign n2467 = n265 & ~n276 ;
  assign n2468 = ( ~n276 & n2179 ) | ( ~n276 & n2467 ) | ( n2179 & n2467 ) ;
  assign n2469 = n273 | n2468 ;
  assign n2470 = ~n280 & n2469 ;
  assign n2471 = n269 | n276 ;
  assign n2472 = ~n273 & n2471 ;
  assign n2473 = n280 | n2472 ;
  assign n2474 = ( n2466 & ~n2470 ) | ( n2466 & n2473 ) | ( ~n2470 & n2473 ) ;
  assign n2475 = n2381 & n2474 ;
  assign n2476 = x140 & ~n685 ;
  assign n2477 = x14 | n688 ;
  assign n2478 = ~n285 & n2477 ;
  assign n2479 = ( ~n310 & n1458 ) | ( ~n310 & n2478 ) | ( n1458 & n2478 ) ;
  assign n2480 = ( n322 & ~n1463 ) | ( n322 & n2479 ) | ( ~n1463 & n2479 ) ;
  assign n2481 = ( n341 & ~n1869 ) | ( n341 & n2480 ) | ( ~n1869 & n2480 ) ;
  assign n2482 = ( ~n1478 & n1874 ) | ( ~n1478 & n2481 ) | ( n1874 & n2481 ) ;
  assign n2483 = ( n1484 & ~n1488 ) | ( n1484 & n2482 ) | ( ~n1488 & n2482 ) ;
  assign n2484 = ( n412 & ~n1500 ) | ( n412 & n2483 ) | ( ~n1500 & n2483 ) ;
  assign n2485 = ( ~n457 & n464 ) | ( ~n457 & n2484 ) | ( n464 & n2484 ) ;
  assign n2486 = ( ~n487 & n488 ) | ( ~n487 & n1508 ) | ( n488 & n1508 ) ;
  assign n2487 = n491 | n2486 ;
  assign n2488 = ~n481 & n2487 ;
  assign n2489 = ( ~n475 & n1519 ) | ( ~n475 & n2488 ) | ( n1519 & n2488 ) ;
  assign n2490 = n498 | n2489 ;
  assign n2491 = ( n511 & n2485 ) | ( n511 & ~n2490 ) | ( n2485 & ~n2490 ) ;
  assign n2492 = ( ~n539 & n558 ) | ( ~n539 & n1523 ) | ( n558 & n1523 ) ;
  assign n2493 = n529 | n2492 ;
  assign n2494 = ~n544 & n2493 ;
  assign n2495 = ( ~n549 & n1545 ) | ( ~n549 & n2494 ) | ( n1545 & n2494 ) ;
  assign n2496 = n523 | n2495 ;
  assign n2497 = n512 | n535 ;
  assign n2498 = ~n532 & n2497 ;
  assign n2499 = n539 | n2498 ;
  assign n2500 = ~n529 & n2499 ;
  assign n2501 = n544 | n2500 ;
  assign n2502 = ~n526 & n2501 ;
  assign n2503 = ( ~n523 & n2242 ) | ( ~n523 & n2502 ) | ( n2242 & n2502 ) ;
  assign n2504 = ( n2491 & ~n2496 ) | ( n2491 & n2503 ) | ( ~n2496 & n2503 ) ;
  assign n2505 = n517 | n555 ;
  assign n2506 = ~n613 & n2505 ;
  assign n2507 = n597 | n2506 ;
  assign n2508 = ~n594 & n2507 ;
  assign n2509 = n591 | n2508 ;
  assign n2510 = ~n588 & n2509 ;
  assign n2511 = ( ~n582 & n1944 ) | ( ~n582 & n2510 ) | ( n1944 & n2510 ) ;
  assign n2512 = n579 | n2511 ;
  assign n2513 = ( ~n597 & n614 ) | ( ~n597 & n1549 ) | ( n614 & n1549 ) ;
  assign n2514 = n594 | n2513 ;
  assign n2515 = ~n591 & n2514 ;
  assign n2516 = ( ~n585 & n1564 ) | ( ~n585 & n2515 ) | ( n1564 & n2515 ) ;
  assign n2517 = n582 | n2516 ;
  assign n2518 = ~n579 & n2517 ;
  assign n2519 = ( n2504 & n2512 ) | ( n2504 & ~n2518 ) | ( n2512 & ~n2518 ) ;
  assign n2520 = n570 | n608 ;
  assign n2521 = ~n634 & n2520 ;
  assign n2522 = n637 | n2521 ;
  assign n2523 = ~n631 & n2522 ;
  assign n2524 = n642 | n2523 ;
  assign n2525 = ~n628 & n2524 ;
  assign n2526 = ( ~n1575 & n1966 ) | ( ~n1575 & n2525 ) | ( n1966 & n2525 ) ;
  assign n2527 = n1581 | n2526 ;
  assign n2528 = ( ~n570 & n623 ) | ( ~n570 & n1568 ) | ( n623 & n1568 ) ;
  assign n2529 = n634 | n2528 ;
  assign n2530 = ~n637 & n2529 ;
  assign n2531 = ( ~n642 & n1576 ) | ( ~n642 & n2530 ) | ( n1576 & n2530 ) ;
  assign n2532 = n628 | n2531 ;
  assign n2533 = ~n647 & n2532 ;
  assign n2534 = ( ~n1581 & n1962 ) | ( ~n1581 & n2533 ) | ( n1962 & n2533 ) ;
  assign n2535 = ( n2519 & n2527 ) | ( n2519 & ~n2534 ) | ( n2527 & ~n2534 ) ;
  assign n2536 = n663 & ~n674 ;
  assign n2537 = ( ~n674 & n2275 ) | ( ~n674 & n2536 ) | ( n2275 & n2536 ) ;
  assign n2538 = n671 | n2537 ;
  assign n2539 = ~n678 & n2538 ;
  assign n2540 = n667 | n674 ;
  assign n2541 = ~n671 & n2540 ;
  assign n2542 = n678 | n2541 ;
  assign n2543 = ( n2535 & ~n2539 ) | ( n2535 & n2542 ) | ( ~n2539 & n2542 ) ;
  assign n2544 = n2476 & n2543 ;
  assign n2545 = x141 & ~n1082 ;
  assign n2546 = x15 | n1085 ;
  assign n2547 = ~n683 & n2546 ;
  assign n2548 = ( ~n708 & n1597 ) | ( ~n708 & n2547 ) | ( n1597 & n2547 ) ;
  assign n2549 = ( n720 & ~n1602 ) | ( n720 & n2548 ) | ( ~n1602 & n2548 ) ;
  assign n2550 = ( n739 & ~n1978 ) | ( n739 & n2549 ) | ( ~n1978 & n2549 ) ;
  assign n2551 = ( ~n1617 & n1983 ) | ( ~n1617 & n2550 ) | ( n1983 & n2550 ) ;
  assign n2552 = ( n1623 & ~n1627 ) | ( n1623 & n2551 ) | ( ~n1627 & n2551 ) ;
  assign n2553 = ( n810 & ~n1639 ) | ( n810 & n2552 ) | ( ~n1639 & n2552 ) ;
  assign n2554 = ( ~n855 & n862 ) | ( ~n855 & n2553 ) | ( n862 & n2553 ) ;
  assign n2555 = ( ~n885 & n886 ) | ( ~n885 & n1647 ) | ( n886 & n1647 ) ;
  assign n2556 = n889 | n2555 ;
  assign n2557 = ~n879 & n2556 ;
  assign n2558 = ( ~n873 & n1658 ) | ( ~n873 & n2557 ) | ( n1658 & n2557 ) ;
  assign n2559 = n896 | n2558 ;
  assign n2560 = ( n909 & n2554 ) | ( n909 & ~n2559 ) | ( n2554 & ~n2559 ) ;
  assign n2561 = ( ~n937 & n956 ) | ( ~n937 & n1662 ) | ( n956 & n1662 ) ;
  assign n2562 = n927 | n2561 ;
  assign n2563 = ~n942 & n2562 ;
  assign n2564 = ( ~n947 & n1684 ) | ( ~n947 & n2563 ) | ( n1684 & n2563 ) ;
  assign n2565 = n921 | n2564 ;
  assign n2566 = n910 | n933 ;
  assign n2567 = ~n930 & n2566 ;
  assign n2568 = n937 | n2567 ;
  assign n2569 = ~n927 & n2568 ;
  assign n2570 = n942 | n2569 ;
  assign n2571 = ~n924 & n2570 ;
  assign n2572 = ( ~n921 & n2338 ) | ( ~n921 & n2571 ) | ( n2338 & n2571 ) ;
  assign n2573 = ( n2560 & ~n2565 ) | ( n2560 & n2572 ) | ( ~n2565 & n2572 ) ;
  assign n2574 = n915 | n953 ;
  assign n2575 = ~n1011 & n2574 ;
  assign n2576 = n995 | n2575 ;
  assign n2577 = ~n992 & n2576 ;
  assign n2578 = n989 | n2577 ;
  assign n2579 = ~n986 & n2578 ;
  assign n2580 = ( ~n980 & n2053 ) | ( ~n980 & n2579 ) | ( n2053 & n2579 ) ;
  assign n2581 = n977 | n2580 ;
  assign n2582 = ( ~n995 & n1012 ) | ( ~n995 & n1688 ) | ( n1012 & n1688 ) ;
  assign n2583 = n992 | n2582 ;
  assign n2584 = ~n989 & n2583 ;
  assign n2585 = ( ~n983 & n1703 ) | ( ~n983 & n2584 ) | ( n1703 & n2584 ) ;
  assign n2586 = n980 | n2585 ;
  assign n2587 = ~n977 & n2586 ;
  assign n2588 = ( n2573 & n2581 ) | ( n2573 & ~n2587 ) | ( n2581 & ~n2587 ) ;
  assign n2589 = n968 | n1006 ;
  assign n2590 = ~n1032 & n2589 ;
  assign n2591 = n1035 | n2590 ;
  assign n2592 = ~n1029 & n2591 ;
  assign n2593 = n1040 | n2592 ;
  assign n2594 = ~n1026 & n2593 ;
  assign n2595 = ( ~n1714 & n2075 ) | ( ~n1714 & n2594 ) | ( n2075 & n2594 ) ;
  assign n2596 = n1720 | n2595 ;
  assign n2597 = ( ~n968 & n1021 ) | ( ~n968 & n1707 ) | ( n1021 & n1707 ) ;
  assign n2598 = n1032 | n2597 ;
  assign n2599 = ~n1035 & n2598 ;
  assign n2600 = ( ~n1040 & n1715 ) | ( ~n1040 & n2599 ) | ( n1715 & n2599 ) ;
  assign n2601 = n1026 | n2600 ;
  assign n2602 = ~n1045 & n2601 ;
  assign n2603 = ( ~n1720 & n2071 ) | ( ~n1720 & n2602 ) | ( n2071 & n2602 ) ;
  assign n2604 = ( n2588 & n2596 ) | ( n2588 & ~n2603 ) | ( n2596 & ~n2603 ) ;
  assign n2605 = n1060 & ~n1071 ;
  assign n2606 = ( ~n1071 & n2371 ) | ( ~n1071 & n2605 ) | ( n2371 & n2605 ) ;
  assign n2607 = n1068 | n2606 ;
  assign n2608 = ~n1075 & n2607 ;
  assign n2609 = n1064 | n1071 ;
  assign n2610 = ~n1068 & n2609 ;
  assign n2611 = n1075 | n2610 ;
  assign n2612 = ( n2604 & ~n2608 ) | ( n2604 & n2611 ) | ( ~n2608 & n2611 ) ;
  assign n2613 = n2545 & n2612 ;
  assign n2614 = x142 & ~n284 ;
  assign n2615 = x16 | n295 ;
  assign n2616 = ~n1080 & n2615 ;
  assign n2617 = ( ~n1105 & n1735 ) | ( ~n1105 & n2616 ) | ( n1735 & n2616 ) ;
  assign n2618 = ( n1117 & ~n1740 ) | ( n1117 & n2617 ) | ( ~n1740 & n2617 ) ;
  assign n2619 = ( n1136 & ~n2087 ) | ( n1136 & n2618 ) | ( ~n2087 & n2618 ) ;
  assign n2620 = ( ~n1755 & n2092 ) | ( ~n1755 & n2619 ) | ( n2092 & n2619 ) ;
  assign n2621 = ( n1761 & ~n1765 ) | ( n1761 & n2620 ) | ( ~n1765 & n2620 ) ;
  assign n2622 = ( n1207 & ~n1777 ) | ( n1207 & n2621 ) | ( ~n1777 & n2621 ) ;
  assign n2623 = ( ~n1252 & n1259 ) | ( ~n1252 & n2622 ) | ( n1259 & n2622 ) ;
  assign n2624 = ( ~n1282 & n1283 ) | ( ~n1282 & n1785 ) | ( n1283 & n1785 ) ;
  assign n2625 = n1286 | n2624 ;
  assign n2626 = ~n1276 & n2625 ;
  assign n2627 = ( ~n1270 & n1796 ) | ( ~n1270 & n2626 ) | ( n1796 & n2626 ) ;
  assign n2628 = n1293 | n2627 ;
  assign n2629 = ( n1306 & n2623 ) | ( n1306 & ~n2628 ) | ( n2623 & ~n2628 ) ;
  assign n2630 = ( ~n1334 & n1353 ) | ( ~n1334 & n1800 ) | ( n1353 & n1800 ) ;
  assign n2631 = n1324 | n2630 ;
  assign n2632 = ~n1339 & n2631 ;
  assign n2633 = ( ~n1344 & n1822 ) | ( ~n1344 & n2632 ) | ( n1822 & n2632 ) ;
  assign n2634 = n1318 | n2633 ;
  assign n2635 = n1307 | n1330 ;
  assign n2636 = ~n1327 & n2635 ;
  assign n2637 = n1334 | n2636 ;
  assign n2638 = ~n1324 & n2637 ;
  assign n2639 = n1339 | n2638 ;
  assign n2640 = ~n1321 & n2639 ;
  assign n2641 = ( ~n1318 & n2434 ) | ( ~n1318 & n2640 ) | ( n2434 & n2640 ) ;
  assign n2642 = ( n2629 & ~n2634 ) | ( n2629 & n2641 ) | ( ~n2634 & n2641 ) ;
  assign n2643 = n1312 | n1350 ;
  assign n2644 = ~n1408 & n2643 ;
  assign n2645 = n1392 | n2644 ;
  assign n2646 = ~n1389 & n2645 ;
  assign n2647 = n1386 | n2646 ;
  assign n2648 = ~n1383 & n2647 ;
  assign n2649 = ( ~n1377 & n2162 ) | ( ~n1377 & n2648 ) | ( n2162 & n2648 ) ;
  assign n2650 = n1374 | n2649 ;
  assign n2651 = ( ~n1392 & n1409 ) | ( ~n1392 & n1826 ) | ( n1409 & n1826 ) ;
  assign n2652 = n1389 | n2651 ;
  assign n2653 = ~n1386 & n2652 ;
  assign n2654 = ( ~n1380 & n1841 ) | ( ~n1380 & n2653 ) | ( n1841 & n2653 ) ;
  assign n2655 = n1377 | n2654 ;
  assign n2656 = ~n1374 & n2655 ;
  assign n2657 = ( n2642 & n2650 ) | ( n2642 & ~n2656 ) | ( n2650 & ~n2656 ) ;
  assign n2658 = n1365 | n1403 ;
  assign n2659 = ~n1429 & n2658 ;
  assign n2660 = n1432 | n2659 ;
  assign n2661 = ~n1426 & n2660 ;
  assign n2662 = n1437 | n2661 ;
  assign n2663 = ~n1423 & n2662 ;
  assign n2664 = ( ~n1851 & n2183 ) | ( ~n1851 & n2663 ) | ( n2183 & n2663 ) ;
  assign n2665 = n268 | n2664 ;
  assign n2666 = ( ~n1365 & n1418 ) | ( ~n1365 & n1845 ) | ( n1418 & n1845 ) ;
  assign n2667 = n1429 | n2666 ;
  assign n2668 = ~n1432 & n2667 ;
  assign n2669 = ( ~n1437 & n1852 ) | ( ~n1437 & n2668 ) | ( n1852 & n2668 ) ;
  assign n2670 = n1423 | n2669 ;
  assign n2671 = ~n1442 & n2670 ;
  assign n2672 = ( ~n268 & n2179 ) | ( ~n268 & n2671 ) | ( n2179 & n2671 ) ;
  assign n2673 = ( n2657 & n2665 ) | ( n2657 & ~n2672 ) | ( n2665 & ~n2672 ) ;
  assign n2674 = ( ~n280 & n282 ) | ( ~n280 & n2467 ) | ( n282 & n2467 ) ;
  assign n2675 = n289 | n2674 ;
  assign n2676 = ~n292 & n2675 ;
  assign n2677 = n281 & ~n289 ;
  assign n2678 = n292 | n2677 ;
  assign n2679 = ( n2673 & ~n2676 ) | ( n2673 & n2678 ) | ( ~n2676 & n2678 ) ;
  assign n2680 = n2614 & n2679 ;
  assign n2681 = x143 & ~n682 ;
  assign n2682 = x17 | n693 ;
  assign n2683 = ~n309 & n2682 ;
  assign n2684 = ( ~n307 & n321 ) | ( ~n307 & n2683 ) | ( n321 & n2683 ) ;
  assign n2685 = ( ~n1464 & n1468 ) | ( ~n1464 & n2684 ) | ( n1468 & n2684 ) ;
  assign n2686 = ( ~n350 & n1472 ) | ( ~n350 & n2685 ) | ( n1472 & n2685 ) ;
  assign n2687 = ( n370 & ~n1878 ) | ( n370 & n2686 ) | ( ~n1878 & n2686 ) ;
  assign n2688 = ( n1884 & ~n1887 ) | ( n1884 & n2687 ) | ( ~n1887 & n2687 ) ;
  assign n2689 = ( n1496 & ~n1898 ) | ( n1496 & n2688 ) | ( ~n1898 & n2688 ) ;
  assign n2690 = ( ~n1509 & n1516 ) | ( ~n1509 & n2689 ) | ( n1516 & n2689 ) ;
  assign n2691 = ( ~n501 & n1532 ) | ( ~n501 & n2690 ) | ( n1532 & n2690 ) ;
  assign n2692 = ( n556 & ~n565 ) | ( n556 & n2691 ) | ( ~n565 & n2691 ) ;
  assign n2693 = n597 | n1542 ;
  assign n2694 = ~n594 & n2693 ;
  assign n2695 = n591 | n2694 ;
  assign n2696 = ~n588 & n2695 ;
  assign n2697 = n585 | n2696 ;
  assign n2698 = ~n582 & n2697 ;
  assign n2699 = ( ~n576 & n2258 ) | ( ~n576 & n2698 ) | ( n2258 & n2698 ) ;
  assign n2700 = n607 | n2699 ;
  assign n2701 = ( ~n622 & n2692 ) | ( ~n622 & n2700 ) | ( n2692 & n2700 ) ;
  assign n2702 = n637 | n1561 ;
  assign n2703 = ~n631 & n2702 ;
  assign n2704 = n642 | n2703 ;
  assign n2705 = ~n628 & n2704 ;
  assign n2706 = n647 | n2705 ;
  assign n2707 = ~n1575 & n2706 ;
  assign n2708 = ( ~n1961 & n2279 ) | ( ~n1961 & n2707 ) | ( n2279 & n2707 ) ;
  assign n2709 = n666 | n2708 ;
  assign n2710 = ( n623 & ~n637 ) | ( n623 & n638 ) | ( ~n637 & n638 ) ;
  assign n2711 = n631 | n2710 ;
  assign n2712 = ~n642 & n2711 ;
  assign n2713 = ( ~n647 & n1577 ) | ( ~n647 & n2712 ) | ( n1577 & n2712 ) ;
  assign n2714 = n1575 | n2713 ;
  assign n2715 = ~n1581 & n2714 ;
  assign n2716 = ( ~n666 & n2275 ) | ( ~n666 & n2715 ) | ( n2275 & n2715 ) ;
  assign n2717 = ( n2701 & n2709 ) | ( n2701 & ~n2716 ) | ( n2709 & ~n2716 ) ;
  assign n2718 = ( ~n678 & n680 ) | ( ~n678 & n2536 ) | ( n680 & n2536 ) ;
  assign n2719 = n687 | n2718 ;
  assign n2720 = ~n690 & n2719 ;
  assign n2721 = n679 & ~n687 ;
  assign n2722 = n690 | n2721 ;
  assign n2723 = ( n2717 & ~n2720 ) | ( n2717 & n2722 ) | ( ~n2720 & n2722 ) ;
  assign n2724 = n2681 & n2723 ;
  assign n2725 = x144 & ~n1079 ;
  assign n2726 = x18 | n1090 ;
  assign n2727 = ~n707 & n2726 ;
  assign n2728 = ( ~n705 & n719 ) | ( ~n705 & n2727 ) | ( n719 & n2727 ) ;
  assign n2729 = ( ~n1603 & n1607 ) | ( ~n1603 & n2728 ) | ( n1607 & n2728 ) ;
  assign n2730 = ( ~n748 & n1611 ) | ( ~n748 & n2729 ) | ( n1611 & n2729 ) ;
  assign n2731 = ( n768 & ~n1987 ) | ( n768 & n2730 ) | ( ~n1987 & n2730 ) ;
  assign n2732 = ( n1993 & ~n1996 ) | ( n1993 & n2731 ) | ( ~n1996 & n2731 ) ;
  assign n2733 = ( n1635 & ~n2007 ) | ( n1635 & n2732 ) | ( ~n2007 & n2732 ) ;
  assign n2734 = ( ~n1648 & n1655 ) | ( ~n1648 & n2733 ) | ( n1655 & n2733 ) ;
  assign n2735 = ( ~n899 & n1671 ) | ( ~n899 & n2734 ) | ( n1671 & n2734 ) ;
  assign n2736 = ( n954 & ~n963 ) | ( n954 & n2735 ) | ( ~n963 & n2735 ) ;
  assign n2737 = n995 | n1681 ;
  assign n2738 = ~n992 & n2737 ;
  assign n2739 = n989 | n2738 ;
  assign n2740 = ~n986 & n2739 ;
  assign n2741 = n983 | n2740 ;
  assign n2742 = ~n980 & n2741 ;
  assign n2743 = ( ~n974 & n2354 ) | ( ~n974 & n2742 ) | ( n2354 & n2742 ) ;
  assign n2744 = n1005 | n2743 ;
  assign n2745 = ( ~n1020 & n2736 ) | ( ~n1020 & n2744 ) | ( n2736 & n2744 ) ;
  assign n2746 = n1035 | n1700 ;
  assign n2747 = ~n1029 & n2746 ;
  assign n2748 = n1040 | n2747 ;
  assign n2749 = ~n1026 & n2748 ;
  assign n2750 = n1045 | n2749 ;
  assign n2751 = ~n1714 & n2750 ;
  assign n2752 = ( ~n2070 & n2375 ) | ( ~n2070 & n2751 ) | ( n2375 & n2751 ) ;
  assign n2753 = n1063 | n2752 ;
  assign n2754 = ( n1021 & ~n1035 ) | ( n1021 & n1036 ) | ( ~n1035 & n1036 ) ;
  assign n2755 = n1029 | n2754 ;
  assign n2756 = ~n1040 & n2755 ;
  assign n2757 = ( ~n1045 & n1716 ) | ( ~n1045 & n2756 ) | ( n1716 & n2756 ) ;
  assign n2758 = n1714 | n2757 ;
  assign n2759 = ~n1720 & n2758 ;
  assign n2760 = ( ~n1063 & n2371 ) | ( ~n1063 & n2759 ) | ( n2371 & n2759 ) ;
  assign n2761 = ( n2745 & n2753 ) | ( n2745 & ~n2760 ) | ( n2753 & ~n2760 ) ;
  assign n2762 = ( ~n1075 & n1077 ) | ( ~n1075 & n2605 ) | ( n1077 & n2605 ) ;
  assign n2763 = n1084 | n2762 ;
  assign n2764 = ~n1087 & n2763 ;
  assign n2765 = n1076 & ~n1084 ;
  assign n2766 = n1087 | n2765 ;
  assign n2767 = ( n2761 & ~n2764 ) | ( n2761 & n2766 ) | ( ~n2764 & n2766 ) ;
  assign n2768 = n2725 & n2767 ;
  assign n2769 = x145 & ~n308 ;
  assign n2770 = x19 | n311 ;
  assign n2771 = ~n1104 & n2770 ;
  assign n2772 = ( ~n1102 & n1116 ) | ( ~n1102 & n2771 ) | ( n1116 & n2771 ) ;
  assign n2773 = ( ~n1741 & n1745 ) | ( ~n1741 & n2772 ) | ( n1745 & n2772 ) ;
  assign n2774 = ( ~n1145 & n1749 ) | ( ~n1145 & n2773 ) | ( n1749 & n2773 ) ;
  assign n2775 = ( n1165 & ~n2096 ) | ( n1165 & n2774 ) | ( ~n2096 & n2774 ) ;
  assign n2776 = ( n2102 & ~n2105 ) | ( n2102 & n2775 ) | ( ~n2105 & n2775 ) ;
  assign n2777 = ( n1773 & ~n2116 ) | ( n1773 & n2776 ) | ( ~n2116 & n2776 ) ;
  assign n2778 = ( ~n1786 & n1793 ) | ( ~n1786 & n2777 ) | ( n1793 & n2777 ) ;
  assign n2779 = ( ~n1296 & n1809 ) | ( ~n1296 & n2778 ) | ( n1809 & n2778 ) ;
  assign n2780 = ( n1351 & ~n1360 ) | ( n1351 & n2779 ) | ( ~n1360 & n2779 ) ;
  assign n2781 = n1392 | n1819 ;
  assign n2782 = ~n1389 & n2781 ;
  assign n2783 = n1386 | n2782 ;
  assign n2784 = ~n1383 & n2783 ;
  assign n2785 = n1380 | n2784 ;
  assign n2786 = ~n1377 & n2785 ;
  assign n2787 = ( ~n1371 & n2450 ) | ( ~n1371 & n2786 ) | ( n2450 & n2786 ) ;
  assign n2788 = n1402 | n2787 ;
  assign n2789 = ( ~n1417 & n2780 ) | ( ~n1417 & n2788 ) | ( n2780 & n2788 ) ;
  assign n2790 = n1432 | n1838 ;
  assign n2791 = ~n1426 & n2790 ;
  assign n2792 = n1437 | n2791 ;
  assign n2793 = ~n1423 & n2792 ;
  assign n2794 = n1442 | n2793 ;
  assign n2795 = ~n1851 & n2794 ;
  assign n2796 = ( ~n265 & n269 ) | ( ~n265 & n2795 ) | ( n269 & n2795 ) ;
  assign n2797 = n276 | n2796 ;
  assign n2798 = ( n1418 & ~n1432 ) | ( n1418 & n1433 ) | ( ~n1432 & n1433 ) ;
  assign n2799 = n1426 | n2798 ;
  assign n2800 = ~n1437 & n2799 ;
  assign n2801 = ( ~n1442 & n1853 ) | ( ~n1442 & n2800 ) | ( n1853 & n2800 ) ;
  assign n2802 = n1851 | n2801 ;
  assign n2803 = ~n268 & n2802 ;
  assign n2804 = ( ~n276 & n2467 ) | ( ~n276 & n2803 ) | ( n2467 & n2803 ) ;
  assign n2805 = ( n2789 & n2797 ) | ( n2789 & ~n2804 ) | ( n2797 & ~n2804 ) ;
  assign n2806 = ( n282 & ~n292 ) | ( n282 & n293 ) | ( ~n292 & n293 ) ;
  assign n2807 = n286 | n2806 ;
  assign n2808 = ~n297 & n2807 ;
  assign n2809 = ~n286 & n1456 ;
  assign n2810 = n297 | n2809 ;
  assign n2811 = ( n2805 & ~n2808 ) | ( n2805 & n2810 ) | ( ~n2808 & n2810 ) ;
  assign n2812 = n2769 & n2811 ;
  assign n2813 = x146 & ~n706 ;
  assign n2814 = x20 | n709 ;
  assign n2815 = ~n306 & n2814 ;
  assign n2816 = ( ~n304 & n1467 ) | ( ~n304 & n2815 ) | ( n1467 & n2815 ) ;
  assign n2817 = ( n341 & ~n348 ) | ( n341 & n2816 ) | ( ~n348 & n2816 ) ;
  assign n2818 = ( ~n1477 & n1873 ) | ( ~n1477 & n2817 ) | ( n1873 & n2817 ) ;
  assign n2819 = ( ~n383 & n1482 ) | ( ~n383 & n2818 ) | ( n1482 & n2818 ) ;
  assign n2820 = ( ~n419 & n2201 ) | ( ~n419 & n2819 ) | ( n2201 & n2819 ) ;
  assign n2821 = ( n1895 & ~n2212 ) | ( n1895 & n2820 ) | ( ~n2212 & n2820 ) ;
  assign n2822 = ( ~n1904 & n1911 ) | ( ~n1904 & n2821 ) | ( n1911 & n2821 ) ;
  assign n2823 = ( ~n1525 & n1925 ) | ( ~n1525 & n2822 ) | ( n1925 & n2822 ) ;
  assign n2824 = ( n1543 & ~n1551 ) | ( n1543 & n2823 ) | ( ~n1551 & n2823 ) ;
  assign n2825 = ( n610 & ~n1571 ) | ( n610 & n2824 ) | ( ~n1571 & n2824 ) ;
  assign n2826 = n652 & ~n1575 ;
  assign n2827 = n1581 | n2826 ;
  assign n2828 = ~n1961 & n2827 ;
  assign n2829 = ( ~n663 & n667 ) | ( ~n663 & n2828 ) | ( n667 & n2828 ) ;
  assign n2830 = n674 | n2829 ;
  assign n2831 = ( n648 & ~n1581 ) | ( n648 & n1962 ) | ( ~n1581 & n1962 ) ;
  assign n2832 = n1961 | n2831 ;
  assign n2833 = ~n666 & n2832 ;
  assign n2834 = ( ~n674 & n2536 ) | ( ~n674 & n2833 ) | ( n2536 & n2833 ) ;
  assign n2835 = ( n2825 & n2830 ) | ( n2825 & ~n2834 ) | ( n2830 & ~n2834 ) ;
  assign n2836 = ( n680 & ~n690 ) | ( n680 & n691 ) | ( ~n690 & n691 ) ;
  assign n2837 = n684 | n2836 ;
  assign n2838 = ~n695 & n2837 ;
  assign n2839 = ~n684 & n1595 ;
  assign n2840 = n695 | n2839 ;
  assign n2841 = ( n2835 & ~n2838 ) | ( n2835 & n2840 ) | ( ~n2838 & n2840 ) ;
  assign n2842 = n2813 & n2841 ;
  assign n2843 = x147 & ~n1103 ;
  assign n2844 = x21 | n1106 ;
  assign n2845 = ~n704 & n2844 ;
  assign n2846 = ( ~n702 & n1606 ) | ( ~n702 & n2845 ) | ( n1606 & n2845 ) ;
  assign n2847 = ( n739 & ~n746 ) | ( n739 & n2846 ) | ( ~n746 & n2846 ) ;
  assign n2848 = ( ~n1616 & n1982 ) | ( ~n1616 & n2847 ) | ( n1982 & n2847 ) ;
  assign n2849 = ( ~n781 & n1621 ) | ( ~n781 & n2848 ) | ( n1621 & n2848 ) ;
  assign n2850 = ( ~n817 & n2297 ) | ( ~n817 & n2849 ) | ( n2297 & n2849 ) ;
  assign n2851 = ( n2004 & ~n2308 ) | ( n2004 & n2850 ) | ( ~n2308 & n2850 ) ;
  assign n2852 = ( ~n2013 & n2020 ) | ( ~n2013 & n2851 ) | ( n2020 & n2851 ) ;
  assign n2853 = ( ~n1664 & n2034 ) | ( ~n1664 & n2852 ) | ( n2034 & n2852 ) ;
  assign n2854 = ( n1682 & ~n1690 ) | ( n1682 & n2853 ) | ( ~n1690 & n2853 ) ;
  assign n2855 = ( n1008 & ~n1710 ) | ( n1008 & n2854 ) | ( ~n1710 & n2854 ) ;
  assign n2856 = n1050 & ~n1714 ;
  assign n2857 = n1720 | n2856 ;
  assign n2858 = ~n2070 & n2857 ;
  assign n2859 = ( ~n1060 & n1064 ) | ( ~n1060 & n2858 ) | ( n1064 & n2858 ) ;
  assign n2860 = n1071 | n2859 ;
  assign n2861 = ( n1046 & ~n1720 ) | ( n1046 & n2071 ) | ( ~n1720 & n2071 ) ;
  assign n2862 = n2070 | n2861 ;
  assign n2863 = ~n1063 & n2862 ;
  assign n2864 = ( ~n1071 & n2605 ) | ( ~n1071 & n2863 ) | ( n2605 & n2863 ) ;
  assign n2865 = ( n2855 & n2860 ) | ( n2855 & ~n2864 ) | ( n2860 & ~n2864 ) ;
  assign n2866 = ( n1077 & ~n1087 ) | ( n1077 & n1088 ) | ( ~n1087 & n1088 ) ;
  assign n2867 = n1081 | n2866 ;
  assign n2868 = ~n1092 & n2867 ;
  assign n2869 = ~n1081 & n1733 ;
  assign n2870 = n1092 | n2869 ;
  assign n2871 = ( n2865 & ~n2868 ) | ( n2865 & n2870 ) | ( ~n2868 & n2870 ) ;
  assign n2872 = n2843 & n2871 ;
  assign n2873 = x148 & ~n305 ;
  assign n2874 = x22 | n316 ;
  assign n2875 = ~n1101 & n2874 ;
  assign n2876 = ( ~n1099 & n1744 ) | ( ~n1099 & n2875 ) | ( n1744 & n2875 ) ;
  assign n2877 = ( n1136 & ~n1143 ) | ( n1136 & n2876 ) | ( ~n1143 & n2876 ) ;
  assign n2878 = ( ~n1754 & n2091 ) | ( ~n1754 & n2877 ) | ( n2091 & n2877 ) ;
  assign n2879 = ( ~n1178 & n1759 ) | ( ~n1178 & n2878 ) | ( n1759 & n2878 ) ;
  assign n2880 = ( ~n1214 & n2393 ) | ( ~n1214 & n2879 ) | ( n2393 & n2879 ) ;
  assign n2881 = ( n2113 & ~n2404 ) | ( n2113 & n2880 ) | ( ~n2404 & n2880 ) ;
  assign n2882 = ( ~n2122 & n2129 ) | ( ~n2122 & n2881 ) | ( n2129 & n2881 ) ;
  assign n2883 = ( ~n1802 & n2143 ) | ( ~n1802 & n2882 ) | ( n2143 & n2882 ) ;
  assign n2884 = ( n1820 & ~n1828 ) | ( n1820 & n2883 ) | ( ~n1828 & n2883 ) ;
  assign n2885 = ( n1405 & ~n1848 ) | ( n1405 & n2884 ) | ( ~n1848 & n2884 ) ;
  assign n2886 = n1447 & ~n1851 ;
  assign n2887 = n268 | n2886 ;
  assign n2888 = ~n265 & n2887 ;
  assign n2889 = ( ~n273 & n277 ) | ( ~n273 & n2888 ) | ( n277 & n2888 ) ;
  assign n2890 = n280 | n2889 ;
  assign n2891 = ( ~n268 & n1443 ) | ( ~n268 & n2179 ) | ( n1443 & n2179 ) ;
  assign n2892 = n265 | n2891 ;
  assign n2893 = ~n276 & n2892 ;
  assign n2894 = ( ~n280 & n282 ) | ( ~n280 & n2893 ) | ( n282 & n2893 ) ;
  assign n2895 = ( n2885 & n2890 ) | ( n2885 & ~n2894 ) | ( n2890 & ~n2894 ) ;
  assign n2896 = n298 | n310 ;
  assign n2897 = ~n313 & n2896 ;
  assign n2898 = n300 & ~n310 ;
  assign n2899 = n313 | n2898 ;
  assign n2900 = ( n2895 & ~n2897 ) | ( n2895 & n2899 ) | ( ~n2897 & n2899 ) ;
  assign n2901 = n2873 & n2900 ;
  assign n2902 = x149 & ~n703 ;
  assign n2903 = x23 | n714 ;
  assign n2904 = ~n303 & n2903 ;
  assign n2905 = ( ~n333 & n337 ) | ( ~n333 & n2904 ) | ( n337 & n2904 ) ;
  assign n2906 = ( ~n349 & n1472 ) | ( ~n349 & n2905 ) | ( n1472 & n2905 ) ;
  assign n2907 = ( n369 & ~n1877 ) | ( n369 & n2906 ) | ( ~n1877 & n2906 ) ;
  assign n2908 = ( ~n1488 & n1882 ) | ( ~n1488 & n2907 ) | ( n1882 & n2907 ) ;
  assign n2909 = ( n411 & ~n1499 ) | ( n411 & n2908 ) | ( ~n1499 & n2908 ) ;
  assign n2910 = ( ~n449 & n2209 ) | ( ~n449 & n2909 ) | ( n2209 & n2909 ) ;
  assign n2911 = ( ~n2218 & n2225 ) | ( ~n2218 & n2910 ) | ( n2225 & n2910 ) ;
  assign n2912 = ( ~n1918 & n2239 ) | ( ~n1918 & n2911 ) | ( n2239 & n2911 ) ;
  assign n2913 = ( n1935 & ~n1941 ) | ( n1935 & n2912 ) | ( ~n1941 & n2912 ) ;
  assign n2914 = ( n1563 & ~n1958 ) | ( n1563 & n2913 ) | ( ~n1958 & n2913 ) ;
  assign n2915 = n1586 & ~n1961 ;
  assign n2916 = n666 | n2915 ;
  assign n2917 = ~n663 & n2916 ;
  assign n2918 = ( ~n671 & n675 ) | ( ~n671 & n2917 ) | ( n675 & n2917 ) ;
  assign n2919 = n678 | n2918 ;
  assign n2920 = ( ~n666 & n1582 ) | ( ~n666 & n2275 ) | ( n1582 & n2275 ) ;
  assign n2921 = n663 | n2920 ;
  assign n2922 = ~n674 & n2921 ;
  assign n2923 = ( ~n678 & n680 ) | ( ~n678 & n2922 ) | ( n680 & n2922 ) ;
  assign n2924 = ( n2914 & n2919 ) | ( n2914 & ~n2923 ) | ( n2919 & ~n2923 ) ;
  assign n2925 = n696 | n708 ;
  assign n2926 = ~n711 & n2925 ;
  assign n2927 = n698 & ~n708 ;
  assign n2928 = n711 | n2927 ;
  assign n2929 = ( n2924 & ~n2926 ) | ( n2924 & n2928 ) | ( ~n2926 & n2928 ) ;
  assign n2930 = n2902 & n2929 ;
  assign n2931 = x150 & ~n1100 ;
  assign n2932 = x24 | n1111 ;
  assign n2933 = ~n701 & n2932 ;
  assign n2934 = ( ~n731 & n735 ) | ( ~n731 & n2933 ) | ( n735 & n2933 ) ;
  assign n2935 = ( ~n747 & n1611 ) | ( ~n747 & n2934 ) | ( n1611 & n2934 ) ;
  assign n2936 = ( n767 & ~n1986 ) | ( n767 & n2935 ) | ( ~n1986 & n2935 ) ;
  assign n2937 = ( ~n1627 & n1991 ) | ( ~n1627 & n2936 ) | ( n1991 & n2936 ) ;
  assign n2938 = ( n809 & ~n1638 ) | ( n809 & n2937 ) | ( ~n1638 & n2937 ) ;
  assign n2939 = ( ~n847 & n2305 ) | ( ~n847 & n2938 ) | ( n2305 & n2938 ) ;
  assign n2940 = ( ~n2314 & n2321 ) | ( ~n2314 & n2939 ) | ( n2321 & n2939 ) ;
  assign n2941 = ( ~n2027 & n2335 ) | ( ~n2027 & n2940 ) | ( n2335 & n2940 ) ;
  assign n2942 = ( n2044 & ~n2050 ) | ( n2044 & n2941 ) | ( ~n2050 & n2941 ) ;
  assign n2943 = ( n1702 & ~n2067 ) | ( n1702 & n2942 ) | ( ~n2067 & n2942 ) ;
  assign n2944 = n1725 & ~n2070 ;
  assign n2945 = n1063 | n2944 ;
  assign n2946 = ~n1060 & n2945 ;
  assign n2947 = ( ~n1068 & n1072 ) | ( ~n1068 & n2946 ) | ( n1072 & n2946 ) ;
  assign n2948 = n1075 | n2947 ;
  assign n2949 = ( ~n1063 & n1721 ) | ( ~n1063 & n2371 ) | ( n1721 & n2371 ) ;
  assign n2950 = n1060 | n2949 ;
  assign n2951 = ~n1071 & n2950 ;
  assign n2952 = ( ~n1075 & n1077 ) | ( ~n1075 & n2951 ) | ( n1077 & n2951 ) ;
  assign n2953 = ( n2943 & n2948 ) | ( n2943 & ~n2952 ) | ( n2948 & ~n2952 ) ;
  assign n2954 = n1093 | n1105 ;
  assign n2955 = ~n1108 & n2954 ;
  assign n2956 = n1095 & ~n1105 ;
  assign n2957 = n1108 | n2956 ;
  assign n2958 = ( n2953 & ~n2955 ) | ( n2953 & n2957 ) | ( ~n2955 & n2957 ) ;
  assign n2959 = n2931 & n2958 ;
  assign n2960 = x151 & ~n302 ;
  assign n2961 = x25 | n334 ;
  assign n2962 = ~n1098 & n2961 ;
  assign n2963 = ( ~n1128 & n1132 ) | ( ~n1128 & n2962 ) | ( n1132 & n2962 ) ;
  assign n2964 = ( ~n1144 & n1749 ) | ( ~n1144 & n2963 ) | ( n1749 & n2963 ) ;
  assign n2965 = ( n1164 & ~n2095 ) | ( n1164 & n2964 ) | ( ~n2095 & n2964 ) ;
  assign n2966 = ( ~n1765 & n2100 ) | ( ~n1765 & n2965 ) | ( n2100 & n2965 ) ;
  assign n2967 = ( n1206 & ~n1776 ) | ( n1206 & n2966 ) | ( ~n1776 & n2966 ) ;
  assign n2968 = ( ~n1244 & n2401 ) | ( ~n1244 & n2967 ) | ( n2401 & n2967 ) ;
  assign n2969 = ( ~n2410 & n2417 ) | ( ~n2410 & n2968 ) | ( n2417 & n2968 ) ;
  assign n2970 = ( ~n2136 & n2431 ) | ( ~n2136 & n2969 ) | ( n2431 & n2969 ) ;
  assign n2971 = ( n2153 & ~n2159 ) | ( n2153 & n2970 ) | ( ~n2159 & n2970 ) ;
  assign n2972 = ( n1840 & ~n2176 ) | ( n1840 & n2971 ) | ( ~n2176 & n2971 ) ;
  assign n2973 = ~n265 & n1860 ;
  assign n2974 = n276 | n2973 ;
  assign n2975 = ~n273 & n2974 ;
  assign n2976 = ( ~n289 & n1455 ) | ( ~n289 & n2975 ) | ( n1455 & n2975 ) ;
  assign n2977 = n292 | n2976 ;
  assign n2978 = ( ~n276 & n1856 ) | ( ~n276 & n2467 ) | ( n1856 & n2467 ) ;
  assign n2979 = n273 | n2978 ;
  assign n2980 = ~n280 & n2979 ;
  assign n2981 = ( ~n292 & n293 ) | ( ~n292 & n2980 ) | ( n293 & n2980 ) ;
  assign n2982 = ( n2972 & n2977 ) | ( n2972 & ~n2981 ) | ( n2977 & ~n2981 ) ;
  assign n2983 = n307 | n1461 ;
  assign n2984 = ~n318 & n2983 ;
  assign n2985 = ~n307 & n1459 ;
  assign n2986 = n318 | n2985 ;
  assign n2987 = ( n2982 & ~n2984 ) | ( n2982 & n2986 ) | ( ~n2984 & n2986 ) ;
  assign n2988 = n2960 & n2987 ;
  assign n2989 = x152 & ~n700 ;
  assign n2990 = x26 | n732 ;
  assign n2991 = ~n332 & n2990 ;
  assign n2992 = ( ~n330 & n1471 ) | ( ~n330 & n2991 ) | ( n1471 & n2991 ) ;
  assign n2993 = ( ~n1476 & n1873 ) | ( ~n1476 & n2992 ) | ( n1873 & n2992 ) ;
  assign n2994 = ( ~n382 & n1481 ) | ( ~n382 & n2993 ) | ( n1481 & n2993 ) ;
  assign n2995 = ( ~n1887 & n2199 ) | ( ~n1887 & n2994 ) | ( n2199 & n2994 ) ;
  assign n2996 = ( n1495 & ~n1897 ) | ( n1495 & n2995 ) | ( ~n1897 & n2995 ) ;
  assign n2997 = ( n464 & ~n1507 ) | ( n464 & n2996 ) | ( ~n1507 & n2996 ) ;
  assign n2998 = ( n510 & ~n2489 ) | ( n510 & n2997 ) | ( ~n2489 & n2997 ) ;
  assign n2999 = ( ~n2232 & n2502 ) | ( ~n2232 & n2998 ) | ( n2502 & n2998 ) ;
  assign n3000 = ( n2249 & ~n2255 ) | ( n2249 & n2999 ) | ( ~n2255 & n2999 ) ;
  assign n3001 = ( n1952 & ~n2272 ) | ( n1952 & n3000 ) | ( ~n2272 & n3000 ) ;
  assign n3002 = ~n663 & n1969 ;
  assign n3003 = n674 | n3002 ;
  assign n3004 = ~n671 & n3003 ;
  assign n3005 = ( ~n687 & n1594 ) | ( ~n687 & n3004 ) | ( n1594 & n3004 ) ;
  assign n3006 = n690 | n3005 ;
  assign n3007 = ( ~n674 & n1965 ) | ( ~n674 & n2536 ) | ( n1965 & n2536 ) ;
  assign n3008 = n671 | n3007 ;
  assign n3009 = ~n678 & n3008 ;
  assign n3010 = ( ~n690 & n691 ) | ( ~n690 & n3009 ) | ( n691 & n3009 ) ;
  assign n3011 = ( n3001 & n3006 ) | ( n3001 & ~n3010 ) | ( n3006 & ~n3010 ) ;
  assign n3012 = n705 | n1600 ;
  assign n3013 = ~n716 & n3012 ;
  assign n3014 = ~n705 & n1598 ;
  assign n3015 = n716 | n3014 ;
  assign n3016 = ( n3011 & ~n3013 ) | ( n3011 & n3015 ) | ( ~n3013 & n3015 ) ;
  assign n3017 = n2989 & n3016 ;
  assign n3018 = x153 & ~n1097 ;
  assign n3019 = x27 | n1129 ;
  assign n3020 = ~n730 & n3019 ;
  assign n3021 = ( ~n728 & n1610 ) | ( ~n728 & n3020 ) | ( n1610 & n3020 ) ;
  assign n3022 = ( ~n1615 & n1982 ) | ( ~n1615 & n3021 ) | ( n1982 & n3021 ) ;
  assign n3023 = ( ~n780 & n1620 ) | ( ~n780 & n3022 ) | ( n1620 & n3022 ) ;
  assign n3024 = ( ~n1996 & n2295 ) | ( ~n1996 & n3023 ) | ( n2295 & n3023 ) ;
  assign n3025 = ( n1634 & ~n2006 ) | ( n1634 & n3024 ) | ( ~n2006 & n3024 ) ;
  assign n3026 = ( n862 & ~n1646 ) | ( n862 & n3025 ) | ( ~n1646 & n3025 ) ;
  assign n3027 = ( n908 & ~n2558 ) | ( n908 & n3026 ) | ( ~n2558 & n3026 ) ;
  assign n3028 = ( ~n2328 & n2571 ) | ( ~n2328 & n3027 ) | ( n2571 & n3027 ) ;
  assign n3029 = ( n2345 & ~n2351 ) | ( n2345 & n3028 ) | ( ~n2351 & n3028 ) ;
  assign n3030 = ( n2061 & ~n2368 ) | ( n2061 & n3029 ) | ( ~n2368 & n3029 ) ;
  assign n3031 = ~n1060 & n2078 ;
  assign n3032 = n1071 | n3031 ;
  assign n3033 = ~n1068 & n3032 ;
  assign n3034 = ( ~n1084 & n1732 ) | ( ~n1084 & n3033 ) | ( n1732 & n3033 ) ;
  assign n3035 = n1087 | n3034 ;
  assign n3036 = ( ~n1071 & n2074 ) | ( ~n1071 & n2605 ) | ( n2074 & n2605 ) ;
  assign n3037 = n1068 | n3036 ;
  assign n3038 = ~n1075 & n3037 ;
  assign n3039 = ( ~n1087 & n1088 ) | ( ~n1087 & n3038 ) | ( n1088 & n3038 ) ;
  assign n3040 = ( n3030 & n3035 ) | ( n3030 & ~n3039 ) | ( n3035 & ~n3039 ) ;
  assign n3041 = n1102 | n1738 ;
  assign n3042 = ~n1113 & n3041 ;
  assign n3043 = ~n1102 & n1736 ;
  assign n3044 = n1113 | n3043 ;
  assign n3045 = ( n3040 & ~n3042 ) | ( n3040 & n3044 ) | ( ~n3042 & n3044 ) ;
  assign n3046 = n3018 & n3045 ;
  assign n3047 = x154 & ~n331 ;
  assign n3048 = x28 | n338 ;
  assign n3049 = ~n1127 & n3048 ;
  assign n3050 = ( ~n1125 & n1748 ) | ( ~n1125 & n3049 ) | ( n1748 & n3049 ) ;
  assign n3051 = ( ~n1753 & n2091 ) | ( ~n1753 & n3050 ) | ( n2091 & n3050 ) ;
  assign n3052 = ( ~n1177 & n1758 ) | ( ~n1177 & n3051 ) | ( n1758 & n3051 ) ;
  assign n3053 = ( ~n2105 & n2391 ) | ( ~n2105 & n3052 ) | ( n2391 & n3052 ) ;
  assign n3054 = ( n1772 & ~n2115 ) | ( n1772 & n3053 ) | ( ~n2115 & n3053 ) ;
  assign n3055 = ( n1259 & ~n1784 ) | ( n1259 & n3054 ) | ( ~n1784 & n3054 ) ;
  assign n3056 = ( n1305 & ~n2627 ) | ( n1305 & n3055 ) | ( ~n2627 & n3055 ) ;
  assign n3057 = ( ~n2424 & n2640 ) | ( ~n2424 & n3056 ) | ( n2640 & n3056 ) ;
  assign n3058 = ( n2441 & ~n2447 ) | ( n2441 & n3057 ) | ( ~n2447 & n3057 ) ;
  assign n3059 = ( n2170 & ~n2464 ) | ( n2170 & n3058 ) | ( ~n2464 & n3058 ) ;
  assign n3060 = ~n273 & n2186 ;
  assign n3061 = n280 | n3060 ;
  assign n3062 = ~n289 & n3061 ;
  assign n3063 = ( ~n286 & n299 ) | ( ~n286 & n3062 ) | ( n299 & n3062 ) ;
  assign n3064 = n297 | n3063 ;
  assign n3065 = ( ~n280 & n282 ) | ( ~n280 & n2182 ) | ( n282 & n2182 ) ;
  assign n3066 = n289 | n3065 ;
  assign n3067 = ~n292 & n3066 ;
  assign n3068 = ( ~n297 & n1460 ) | ( ~n297 & n3067 ) | ( n1460 & n3067 ) ;
  assign n3069 = ( n3059 & n3064 ) | ( n3059 & ~n3068 ) | ( n3064 & ~n3068 ) ;
  assign n3070 = n320 & ~n336 ;
  assign n3071 = n323 | n336 ;
  assign n3072 = ( n3069 & ~n3070 ) | ( n3069 & n3071 ) | ( ~n3070 & n3071 ) ;
  assign n3073 = n3047 & n3072 ;
  assign n3074 = x155 & ~n729 ;
  assign n3075 = x29 | n736 ;
  assign n3076 = ~n329 & n3075 ;
  assign n3077 = ( ~n327 & n1872 ) | ( ~n327 & n3076 ) | ( n1872 & n3076 ) ;
  assign n3078 = ( n369 & ~n380 ) | ( n369 & n3077 ) | ( ~n380 & n3077 ) ;
  assign n3079 = ( ~n1487 & n1881 ) | ( ~n1487 & n3078 ) | ( n1881 & n3078 ) ;
  assign n3080 = ( n409 & ~n419 ) | ( n409 & n3079 ) | ( ~n419 & n3079 ) ;
  assign n3081 = ( n1894 & ~n2211 ) | ( n1894 & n3080 ) | ( ~n2211 & n3080 ) ;
  assign n3082 = ( n1516 & ~n1903 ) | ( n1516 & n3081 ) | ( ~n1903 & n3081 ) ;
  assign n3083 = ( ~n500 & n1531 ) | ( ~n500 & n3082 ) | ( n1531 & n3082 ) ;
  assign n3084 = ( n551 & ~n2496 ) | ( n551 & n3083 ) | ( ~n2496 & n3083 ) ;
  assign n3085 = ( n2511 & ~n2517 ) | ( n2511 & n3084 ) | ( ~n2517 & n3084 ) ;
  assign n3086 = ( n2266 & ~n2533 ) | ( n2266 & n3085 ) | ( ~n2533 & n3085 ) ;
  assign n3087 = ~n671 & n2282 ;
  assign n3088 = n678 | n3087 ;
  assign n3089 = ~n687 & n3088 ;
  assign n3090 = ( ~n684 & n697 ) | ( ~n684 & n3089 ) | ( n697 & n3089 ) ;
  assign n3091 = n695 | n3090 ;
  assign n3092 = ( ~n678 & n680 ) | ( ~n678 & n2278 ) | ( n680 & n2278 ) ;
  assign n3093 = n687 | n3092 ;
  assign n3094 = ~n690 & n3093 ;
  assign n3095 = ( ~n695 & n1599 ) | ( ~n695 & n3094 ) | ( n1599 & n3094 ) ;
  assign n3096 = ( n3086 & n3091 ) | ( n3086 & ~n3095 ) | ( n3091 & ~n3095 ) ;
  assign n3097 = n718 & ~n734 ;
  assign n3098 = n721 | n734 ;
  assign n3099 = ( n3096 & ~n3097 ) | ( n3096 & n3098 ) | ( ~n3097 & n3098 ) ;
  assign n3100 = n3074 & n3099 ;
  assign n3101 = x156 & ~n1126 ;
  assign n3102 = x30 | n1133 ;
  assign n3103 = ~n727 & n3102 ;
  assign n3104 = ( ~n725 & n1981 ) | ( ~n725 & n3103 ) | ( n1981 & n3103 ) ;
  assign n3105 = ( n767 & ~n778 ) | ( n767 & n3104 ) | ( ~n778 & n3104 ) ;
  assign n3106 = ( ~n1626 & n1990 ) | ( ~n1626 & n3105 ) | ( n1990 & n3105 ) ;
  assign n3107 = ( n807 & ~n817 ) | ( n807 & n3106 ) | ( ~n817 & n3106 ) ;
  assign n3108 = ( n2003 & ~n2307 ) | ( n2003 & n3107 ) | ( ~n2307 & n3107 ) ;
  assign n3109 = ( n1655 & ~n2012 ) | ( n1655 & n3108 ) | ( ~n2012 & n3108 ) ;
  assign n3110 = ( ~n898 & n1670 ) | ( ~n898 & n3109 ) | ( n1670 & n3109 ) ;
  assign n3111 = ( n949 & ~n2565 ) | ( n949 & n3110 ) | ( ~n2565 & n3110 ) ;
  assign n3112 = ( n2580 & ~n2586 ) | ( n2580 & n3111 ) | ( ~n2586 & n3111 ) ;
  assign n3113 = ( n2362 & ~n2602 ) | ( n2362 & n3112 ) | ( ~n2602 & n3112 ) ;
  assign n3114 = ~n1068 & n2378 ;
  assign n3115 = n1075 | n3114 ;
  assign n3116 = ~n1084 & n3115 ;
  assign n3117 = ( ~n1081 & n1094 ) | ( ~n1081 & n3116 ) | ( n1094 & n3116 ) ;
  assign n3118 = n1092 | n3117 ;
  assign n3119 = ( ~n1075 & n1077 ) | ( ~n1075 & n2374 ) | ( n1077 & n2374 ) ;
  assign n3120 = n1084 | n3119 ;
  assign n3121 = ~n1087 & n3120 ;
  assign n3122 = ( ~n1092 & n1737 ) | ( ~n1092 & n3121 ) | ( n1737 & n3121 ) ;
  assign n3123 = ( n3113 & n3118 ) | ( n3113 & ~n3122 ) | ( n3118 & ~n3122 ) ;
  assign n3124 = n1115 & ~n1131 ;
  assign n3125 = n1118 | n1131 ;
  assign n3126 = ( n3123 & ~n3124 ) | ( n3123 & n3125 ) | ( ~n3124 & n3125 ) ;
  assign n3127 = n3101 & n3126 ;
  assign n3128 = x157 & ~n328 ;
  assign n3129 = x31 | n343 ;
  assign n3130 = ~n1124 & n3129 ;
  assign n3131 = ( ~n1122 & n2090 ) | ( ~n1122 & n3130 ) | ( n2090 & n3130 ) ;
  assign n3132 = ( n1164 & ~n1175 ) | ( n1164 & n3131 ) | ( ~n1175 & n3131 ) ;
  assign n3133 = ( ~n1764 & n2099 ) | ( ~n1764 & n3132 ) | ( n2099 & n3132 ) ;
  assign n3134 = ( n1204 & ~n1214 ) | ( n1204 & n3133 ) | ( ~n1214 & n3133 ) ;
  assign n3135 = ( n2112 & ~n2403 ) | ( n2112 & n3134 ) | ( ~n2403 & n3134 ) ;
  assign n3136 = ( n1793 & ~n2121 ) | ( n1793 & n3135 ) | ( ~n2121 & n3135 ) ;
  assign n3137 = ( ~n1295 & n1808 ) | ( ~n1295 & n3136 ) | ( n1808 & n3136 ) ;
  assign n3138 = ( n1346 & ~n2634 ) | ( n1346 & n3137 ) | ( ~n2634 & n3137 ) ;
  assign n3139 = ( n2649 & ~n2655 ) | ( n2649 & n3138 ) | ( ~n2655 & n3138 ) ;
  assign n3140 = ( n2458 & ~n2671 ) | ( n2458 & n3139 ) | ( ~n2671 & n3139 ) ;
  assign n3141 = ~n289 & n2473 ;
  assign n3142 = n292 | n3141 ;
  assign n3143 = ~n286 & n3142 ;
  assign n3144 = ( ~n310 & n1458 ) | ( ~n310 & n3143 ) | ( n1458 & n3143 ) ;
  assign n3145 = n313 | n3144 ;
  assign n3146 = ( ~n292 & n293 ) | ( ~n292 & n2470 ) | ( n293 & n2470 ) ;
  assign n3147 = n286 | n3146 ;
  assign n3148 = ~n297 & n3147 ;
  assign n3149 = ( ~n313 & n314 ) | ( ~n313 & n3148 ) | ( n314 & n3148 ) ;
  assign n3150 = ( n3140 & n3145 ) | ( n3140 & ~n3149 ) | ( n3145 & ~n3149 ) ;
  assign n3151 = ~n340 & n1466 ;
  assign n3152 = n340 | n1469 ;
  assign n3153 = ( n3150 & ~n3151 ) | ( n3150 & n3152 ) | ( ~n3151 & n3152 ) ;
  assign n3154 = n3128 & n3153 ;
  assign n3155 = x158 & ~n726 ;
  assign n3156 = x32 | n741 ;
  assign n3157 = ~n326 & n3156 ;
  assign n3158 = ( ~n361 & n365 ) | ( ~n361 & n3157 ) | ( n365 & n3157 ) ;
  assign n3159 = ( ~n381 & n1481 ) | ( ~n381 & n3158 ) | ( n1481 & n3158 ) ;
  assign n3160 = ( ~n1886 & n2198 ) | ( ~n1886 & n3159 ) | ( n2198 & n3159 ) ;
  assign n3161 = ( n1493 & ~n1499 ) | ( n1493 & n3160 ) | ( ~n1499 & n3160 ) ;
  assign n3162 = ( ~n445 & n2208 ) | ( ~n445 & n3161 ) | ( n2208 & n3161 ) ;
  assign n3163 = ( n1911 & ~n2217 ) | ( n1911 & n3162 ) | ( ~n2217 & n3162 ) ;
  assign n3164 = ( ~n1524 & n1924 ) | ( ~n1524 & n3163 ) | ( n1924 & n3163 ) ;
  assign n3165 = ( ~n565 & n1541 ) | ( ~n565 & n3164 ) | ( n1541 & n3164 ) ;
  assign n3166 = ( ~n621 & n2699 ) | ( ~n621 & n3165 ) | ( n2699 & n3165 ) ;
  assign n3167 = ( n2527 & ~n2715 ) | ( n2527 & n3166 ) | ( ~n2715 & n3166 ) ;
  assign n3168 = ~n687 & n2542 ;
  assign n3169 = n690 | n3168 ;
  assign n3170 = ~n684 & n3169 ;
  assign n3171 = ( ~n708 & n1597 ) | ( ~n708 & n3170 ) | ( n1597 & n3170 ) ;
  assign n3172 = n711 | n3171 ;
  assign n3173 = ( ~n690 & n691 ) | ( ~n690 & n2539 ) | ( n691 & n2539 ) ;
  assign n3174 = n684 | n3173 ;
  assign n3175 = ~n695 & n3174 ;
  assign n3176 = ( ~n711 & n712 ) | ( ~n711 & n3175 ) | ( n712 & n3175 ) ;
  assign n3177 = ( n3167 & n3172 ) | ( n3167 & ~n3176 ) | ( n3172 & ~n3176 ) ;
  assign n3178 = ~n738 & n1605 ;
  assign n3179 = n738 | n1608 ;
  assign n3180 = ( n3177 & ~n3178 ) | ( n3177 & n3179 ) | ( ~n3178 & n3179 ) ;
  assign n3181 = n3155 & n3180 ;
  assign n3182 = x159 & ~n1123 ;
  assign n3183 = x33 | n1138 ;
  assign n3184 = ~n724 & n3183 ;
  assign n3185 = ( ~n759 & n763 ) | ( ~n759 & n3184 ) | ( n763 & n3184 ) ;
  assign n3186 = ( ~n779 & n1620 ) | ( ~n779 & n3185 ) | ( n1620 & n3185 ) ;
  assign n3187 = ( ~n1995 & n2294 ) | ( ~n1995 & n3186 ) | ( n2294 & n3186 ) ;
  assign n3188 = ( n1632 & ~n1638 ) | ( n1632 & n3187 ) | ( ~n1638 & n3187 ) ;
  assign n3189 = ( ~n843 & n2304 ) | ( ~n843 & n3188 ) | ( n2304 & n3188 ) ;
  assign n3190 = ( n2020 & ~n2313 ) | ( n2020 & n3189 ) | ( ~n2313 & n3189 ) ;
  assign n3191 = ( ~n1663 & n2033 ) | ( ~n1663 & n3190 ) | ( n2033 & n3190 ) ;
  assign n3192 = ( ~n963 & n1680 ) | ( ~n963 & n3191 ) | ( n1680 & n3191 ) ;
  assign n3193 = ( ~n1019 & n2743 ) | ( ~n1019 & n3192 ) | ( n2743 & n3192 ) ;
  assign n3194 = ( n2596 & ~n2759 ) | ( n2596 & n3193 ) | ( ~n2759 & n3193 ) ;
  assign n3195 = ~n1084 & n2611 ;
  assign n3196 = n1087 | n3195 ;
  assign n3197 = ~n1081 & n3196 ;
  assign n3198 = ( ~n1105 & n1735 ) | ( ~n1105 & n3197 ) | ( n1735 & n3197 ) ;
  assign n3199 = n1108 | n3198 ;
  assign n3200 = ( ~n1087 & n1088 ) | ( ~n1087 & n2608 ) | ( n1088 & n2608 ) ;
  assign n3201 = n1081 | n3200 ;
  assign n3202 = ~n1092 & n3201 ;
  assign n3203 = ( ~n1108 & n1109 ) | ( ~n1108 & n3202 ) | ( n1109 & n3202 ) ;
  assign n3204 = ( n3194 & n3199 ) | ( n3194 & ~n3203 ) | ( n3199 & ~n3203 ) ;
  assign n3205 = ~n1135 & n1743 ;
  assign n3206 = n1135 | n1746 ;
  assign n3207 = ( n3204 & ~n3205 ) | ( n3204 & n3206 ) | ( ~n3205 & n3206 ) ;
  assign n3208 = n3182 & n3207 ;
  assign n3209 = x160 & ~n325 ;
  assign n3210 = x34 | n362 ;
  assign n3211 = ~n1121 & n3210 ;
  assign n3212 = ( ~n1156 & n1160 ) | ( ~n1156 & n3211 ) | ( n1160 & n3211 ) ;
  assign n3213 = ( ~n1176 & n1758 ) | ( ~n1176 & n3212 ) | ( n1758 & n3212 ) ;
  assign n3214 = ( ~n2104 & n2390 ) | ( ~n2104 & n3213 ) | ( n2390 & n3213 ) ;
  assign n3215 = ( n1770 & ~n1776 ) | ( n1770 & n3214 ) | ( ~n1776 & n3214 ) ;
  assign n3216 = ( ~n1240 & n2400 ) | ( ~n1240 & n3215 ) | ( n2400 & n3215 ) ;
  assign n3217 = ( n2129 & ~n2409 ) | ( n2129 & n3216 ) | ( ~n2409 & n3216 ) ;
  assign n3218 = ( ~n1801 & n2142 ) | ( ~n1801 & n3217 ) | ( n2142 & n3217 ) ;
  assign n3219 = ( ~n1360 & n1818 ) | ( ~n1360 & n3218 ) | ( n1818 & n3218 ) ;
  assign n3220 = ( ~n1416 & n2787 ) | ( ~n1416 & n3219 ) | ( n2787 & n3219 ) ;
  assign n3221 = ( n2665 & ~n2803 ) | ( n2665 & n3220 ) | ( ~n2803 & n3220 ) ;
  assign n3222 = ~n286 & n2678 ;
  assign n3223 = n297 | n3222 ;
  assign n3224 = ~n310 & n3223 ;
  assign n3225 = ( ~n307 & n321 ) | ( ~n307 & n3224 ) | ( n321 & n3224 ) ;
  assign n3226 = n318 | n3225 ;
  assign n3227 = ( ~n297 & n1460 ) | ( ~n297 & n2676 ) | ( n1460 & n2676 ) ;
  assign n3228 = n310 | n3227 ;
  assign n3229 = ~n313 & n3228 ;
  assign n3230 = ( ~n318 & n1463 ) | ( ~n318 & n3229 ) | ( n1463 & n3229 ) ;
  assign n3231 = ( n3221 & n3226 ) | ( n3221 & ~n3230 ) | ( n3226 & ~n3230 ) ;
  assign n3232 = ~n345 & n1870 ;
  assign n3233 = ( n346 & n3231 ) | ( n346 & ~n3232 ) | ( n3231 & ~n3232 ) ;
  assign n3234 = n3209 & n3233 ;
  assign n3235 = x161 & ~n723 ;
  assign n3236 = x35 | n760 ;
  assign n3237 = ~n360 & n3236 ;
  assign n3238 = ( ~n358 & n1480 ) | ( ~n358 & n3237 ) | ( n1480 & n3237 ) ;
  assign n3239 = ( ~n1486 & n1881 ) | ( ~n1486 & n3238 ) | ( n1881 & n3238 ) ;
  assign n3240 = ( n408 & ~n418 ) | ( n408 & n3239 ) | ( ~n418 & n3239 ) ;
  assign n3241 = ( n1892 & ~n1897 ) | ( n1892 & n3240 ) | ( ~n1897 & n3240 ) ;
  assign n3242 = ( n463 & ~n1506 ) | ( n463 & n3241 ) | ( ~n1506 & n3241 ) ;
  assign n3243 = ( n2225 & ~n2488 ) | ( n2225 & n3242 ) | ( ~n2488 & n3242 ) ;
  assign n3244 = ( ~n1917 & n2238 ) | ( ~n1917 & n3243 ) | ( n2238 & n3243 ) ;
  assign n3245 = ( ~n1551 & n1934 ) | ( ~n1551 & n3244 ) | ( n1934 & n3244 ) ;
  assign n3246 = ( n609 & ~n1570 ) | ( n609 & n3245 ) | ( ~n1570 & n3245 ) ;
  assign n3247 = ( n2709 & ~n2833 ) | ( n2709 & n3246 ) | ( ~n2833 & n3246 ) ;
  assign n3248 = ~n684 & n2722 ;
  assign n3249 = n695 | n3248 ;
  assign n3250 = ~n708 & n3249 ;
  assign n3251 = ( ~n705 & n719 ) | ( ~n705 & n3250 ) | ( n719 & n3250 ) ;
  assign n3252 = n716 | n3251 ;
  assign n3253 = ( ~n695 & n1599 ) | ( ~n695 & n2720 ) | ( n1599 & n2720 ) ;
  assign n3254 = n708 | n3253 ;
  assign n3255 = ~n711 & n3254 ;
  assign n3256 = ( ~n716 & n1602 ) | ( ~n716 & n3255 ) | ( n1602 & n3255 ) ;
  assign n3257 = ( n3247 & n3252 ) | ( n3247 & ~n3256 ) | ( n3252 & ~n3256 ) ;
  assign n3258 = ~n743 & n1979 ;
  assign n3259 = ( n744 & n3257 ) | ( n744 & ~n3258 ) | ( n3257 & ~n3258 ) ;
  assign n3260 = n3235 & n3259 ;
  assign n3261 = x162 & ~n1120 ;
  assign n3262 = x36 | n1157 ;
  assign n3263 = ~n758 & n3262 ;
  assign n3264 = ( ~n756 & n1619 ) | ( ~n756 & n3263 ) | ( n1619 & n3263 ) ;
  assign n3265 = ( ~n1625 & n1990 ) | ( ~n1625 & n3264 ) | ( n1990 & n3264 ) ;
  assign n3266 = ( n806 & ~n816 ) | ( n806 & n3265 ) | ( ~n816 & n3265 ) ;
  assign n3267 = ( n2001 & ~n2006 ) | ( n2001 & n3266 ) | ( ~n2006 & n3266 ) ;
  assign n3268 = ( n861 & ~n1645 ) | ( n861 & n3267 ) | ( ~n1645 & n3267 ) ;
  assign n3269 = ( n2321 & ~n2557 ) | ( n2321 & n3268 ) | ( ~n2557 & n3268 ) ;
  assign n3270 = ( ~n2026 & n2334 ) | ( ~n2026 & n3269 ) | ( n2334 & n3269 ) ;
  assign n3271 = ( ~n1690 & n2043 ) | ( ~n1690 & n3270 ) | ( n2043 & n3270 ) ;
  assign n3272 = ( n1007 & ~n1709 ) | ( n1007 & n3271 ) | ( ~n1709 & n3271 ) ;
  assign n3273 = ( n2753 & ~n2863 ) | ( n2753 & n3272 ) | ( ~n2863 & n3272 ) ;
  assign n3274 = ~n1081 & n2766 ;
  assign n3275 = n1092 | n3274 ;
  assign n3276 = ~n1105 & n3275 ;
  assign n3277 = ( ~n1102 & n1116 ) | ( ~n1102 & n3276 ) | ( n1116 & n3276 ) ;
  assign n3278 = n1113 | n3277 ;
  assign n3279 = ( ~n1092 & n1737 ) | ( ~n1092 & n2764 ) | ( n1737 & n2764 ) ;
  assign n3280 = n1105 | n3279 ;
  assign n3281 = ~n1108 & n3280 ;
  assign n3282 = ( ~n1113 & n1740 ) | ( ~n1113 & n3281 ) | ( n1740 & n3281 ) ;
  assign n3283 = ( n3273 & n3278 ) | ( n3273 & ~n3282 ) | ( n3278 & ~n3282 ) ;
  assign n3284 = ~n1140 & n2088 ;
  assign n3285 = ( n1141 & n3283 ) | ( n1141 & ~n3284 ) | ( n3283 & ~n3284 ) ;
  assign n3286 = n3261 & n3285 ;
  assign n3287 = x163 & ~n359 ;
  assign n3288 = x37 | n366 ;
  assign n3289 = ~n1155 & n3288 ;
  assign n3290 = ( ~n1153 & n1757 ) | ( ~n1153 & n3289 ) | ( n1757 & n3289 ) ;
  assign n3291 = ( ~n1763 & n2099 ) | ( ~n1763 & n3290 ) | ( n2099 & n3290 ) ;
  assign n3292 = ( n1203 & ~n1213 ) | ( n1203 & n3291 ) | ( ~n1213 & n3291 ) ;
  assign n3293 = ( n2110 & ~n2115 ) | ( n2110 & n3292 ) | ( ~n2115 & n3292 ) ;
  assign n3294 = ( n1258 & ~n1783 ) | ( n1258 & n3293 ) | ( ~n1783 & n3293 ) ;
  assign n3295 = ( n2417 & ~n2626 ) | ( n2417 & n3294 ) | ( ~n2626 & n3294 ) ;
  assign n3296 = ( ~n2135 & n2430 ) | ( ~n2135 & n3295 ) | ( n2430 & n3295 ) ;
  assign n3297 = ( ~n1828 & n2152 ) | ( ~n1828 & n3296 ) | ( n2152 & n3296 ) ;
  assign n3298 = ( n1404 & ~n1847 ) | ( n1404 & n3297 ) | ( ~n1847 & n3297 ) ;
  assign n3299 = ( n2797 & ~n2893 ) | ( n2797 & n3298 ) | ( ~n2893 & n3298 ) ;
  assign n3300 = ~n310 & n2810 ;
  assign n3301 = n313 | n3300 ;
  assign n3302 = ~n307 & n3301 ;
  assign n3303 = ( ~n304 & n1467 ) | ( ~n304 & n3302 ) | ( n1467 & n3302 ) ;
  assign n3304 = n336 | n3303 ;
  assign n3305 = ( ~n313 & n314 ) | ( ~n313 & n2808 ) | ( n314 & n2808 ) ;
  assign n3306 = n307 | n3305 ;
  assign n3307 = ~n318 & n3306 ;
  assign n3308 = ( ~n336 & n1464 ) | ( ~n336 & n3307 ) | ( n1464 & n3307 ) ;
  assign n3309 = ( n3299 & n3304 ) | ( n3299 & ~n3308 ) | ( n3304 & ~n3308 ) ;
  assign n3310 = n351 & ~n364 ;
  assign n3311 = ( n1474 & n3309 ) | ( n1474 & ~n3310 ) | ( n3309 & ~n3310 ) ;
  assign n3312 = n3287 & n3311 ;
  assign n3313 = x164 & ~n757 ;
  assign n3314 = x38 | n764 ;
  assign n3315 = ~n357 & n3314 ;
  assign n3316 = ( ~n355 & n1880 ) | ( ~n355 & n3315 ) | ( n1880 & n3315 ) ;
  assign n3317 = ( ~n416 & n2198 ) | ( ~n416 & n3316 ) | ( n2198 & n3316 ) ;
  assign n3318 = ( n1492 & ~n1498 ) | ( n1492 & n3317 ) | ( ~n1498 & n3317 ) ;
  assign n3319 = ( n2206 & ~n2211 ) | ( n2206 & n3318 ) | ( ~n2211 & n3318 ) ;
  assign n3320 = ( n1515 & ~n1902 ) | ( n1515 & n3319 ) | ( ~n1902 & n3319 ) ;
  assign n3321 = ( ~n495 & n510 ) | ( ~n495 & n3320 ) | ( n510 & n3320 ) ;
  assign n3322 = ( ~n2231 & n2501 ) | ( ~n2231 & n3321 ) | ( n2501 & n3321 ) ;
  assign n3323 = ( ~n1941 & n2248 ) | ( ~n1941 & n3322 ) | ( n2248 & n3322 ) ;
  assign n3324 = ( n1562 & ~n1957 ) | ( n1562 & n3323 ) | ( ~n1957 & n3323 ) ;
  assign n3325 = ( n2830 & ~n2922 ) | ( n2830 & n3324 ) | ( ~n2922 & n3324 ) ;
  assign n3326 = ~n708 & n2840 ;
  assign n3327 = n711 | n3326 ;
  assign n3328 = ~n705 & n3327 ;
  assign n3329 = ( ~n702 & n1606 ) | ( ~n702 & n3328 ) | ( n1606 & n3328 ) ;
  assign n3330 = n734 | n3329 ;
  assign n3331 = ( ~n711 & n712 ) | ( ~n711 & n2838 ) | ( n712 & n2838 ) ;
  assign n3332 = n705 | n3331 ;
  assign n3333 = ~n716 & n3332 ;
  assign n3334 = ( ~n734 & n1603 ) | ( ~n734 & n3333 ) | ( n1603 & n3333 ) ;
  assign n3335 = ( n3325 & n3330 ) | ( n3325 & ~n3334 ) | ( n3330 & ~n3334 ) ;
  assign n3336 = n749 & ~n762 ;
  assign n3337 = ( n1613 & n3335 ) | ( n1613 & ~n3336 ) | ( n3335 & ~n3336 ) ;
  assign n3338 = n3313 & n3337 ;
  assign n3339 = x165 & ~n1154 ;
  assign n3340 = x39 | n1161 ;
  assign n3341 = ~n755 & n3340 ;
  assign n3342 = ( ~n753 & n1989 ) | ( ~n753 & n3341 ) | ( n1989 & n3341 ) ;
  assign n3343 = ( ~n814 & n2294 ) | ( ~n814 & n3342 ) | ( n2294 & n3342 ) ;
  assign n3344 = ( n1631 & ~n1637 ) | ( n1631 & n3343 ) | ( ~n1637 & n3343 ) ;
  assign n3345 = ( n2302 & ~n2307 ) | ( n2302 & n3344 ) | ( ~n2307 & n3344 ) ;
  assign n3346 = ( n1654 & ~n2011 ) | ( n1654 & n3345 ) | ( ~n2011 & n3345 ) ;
  assign n3347 = ( ~n893 & n908 ) | ( ~n893 & n3346 ) | ( n908 & n3346 ) ;
  assign n3348 = ( ~n2327 & n2570 ) | ( ~n2327 & n3347 ) | ( n2570 & n3347 ) ;
  assign n3349 = ( ~n2050 & n2344 ) | ( ~n2050 & n3348 ) | ( n2344 & n3348 ) ;
  assign n3350 = ( n1701 & ~n2066 ) | ( n1701 & n3349 ) | ( ~n2066 & n3349 ) ;
  assign n3351 = ( n2860 & ~n2951 ) | ( n2860 & n3350 ) | ( ~n2951 & n3350 ) ;
  assign n3352 = ~n1105 & n2870 ;
  assign n3353 = n1108 | n3352 ;
  assign n3354 = ~n1102 & n3353 ;
  assign n3355 = ( ~n1099 & n1744 ) | ( ~n1099 & n3354 ) | ( n1744 & n3354 ) ;
  assign n3356 = n1131 | n3355 ;
  assign n3357 = ( ~n1108 & n1109 ) | ( ~n1108 & n2868 ) | ( n1109 & n2868 ) ;
  assign n3358 = n1102 | n3357 ;
  assign n3359 = ~n1113 & n3358 ;
  assign n3360 = ( ~n1131 & n1741 ) | ( ~n1131 & n3359 ) | ( n1741 & n3359 ) ;
  assign n3361 = ( n3351 & n3356 ) | ( n3351 & ~n3360 ) | ( n3356 & ~n3360 ) ;
  assign n3362 = n1146 & ~n1159 ;
  assign n3363 = ( n1751 & n3361 ) | ( n1751 & ~n3362 ) | ( n3361 & ~n3362 ) ;
  assign n3364 = n3339 & n3363 ;
  assign n3365 = x166 & ~n356 ;
  assign n3366 = x40 | n371 ;
  assign n3367 = ~n1152 & n3366 ;
  assign n3368 = ( ~n1150 & n2098 ) | ( ~n1150 & n3367 ) | ( n2098 & n3367 ) ;
  assign n3369 = ( ~n1211 & n2390 ) | ( ~n1211 & n3368 ) | ( n2390 & n3368 ) ;
  assign n3370 = ( n1769 & ~n1775 ) | ( n1769 & n3369 ) | ( ~n1775 & n3369 ) ;
  assign n3371 = ( n2398 & ~n2403 ) | ( n2398 & n3370 ) | ( ~n2403 & n3370 ) ;
  assign n3372 = ( n1792 & ~n2120 ) | ( n1792 & n3371 ) | ( ~n2120 & n3371 ) ;
  assign n3373 = ( ~n1290 & n1305 ) | ( ~n1290 & n3372 ) | ( n1305 & n3372 ) ;
  assign n3374 = ( ~n2423 & n2639 ) | ( ~n2423 & n3373 ) | ( n2639 & n3373 ) ;
  assign n3375 = ( ~n2159 & n2440 ) | ( ~n2159 & n3374 ) | ( n2440 & n3374 ) ;
  assign n3376 = ( n1839 & ~n2175 ) | ( n1839 & n3375 ) | ( ~n2175 & n3375 ) ;
  assign n3377 = ( n2890 & ~n2980 ) | ( n2890 & n3376 ) | ( ~n2980 & n3376 ) ;
  assign n3378 = ~n307 & n2899 ;
  assign n3379 = n318 | n3378 ;
  assign n3380 = ~n304 & n3379 ;
  assign n3381 = ( ~n333 & n337 ) | ( ~n333 & n3380 ) | ( n337 & n3380 ) ;
  assign n3382 = n340 | n3381 ;
  assign n3383 = ( ~n318 & n1463 ) | ( ~n318 & n2897 ) | ( n1463 & n2897 ) ;
  assign n3384 = n304 | n3383 ;
  assign n3385 = ~n336 & n3384 ;
  assign n3386 = ( ~n340 & n348 ) | ( ~n340 & n3385 ) | ( n348 & n3385 ) ;
  assign n3387 = ( n3377 & n3382 ) | ( n3377 & ~n3386 ) | ( n3382 & ~n3386 ) ;
  assign n3388 = ~n368 & n1478 ;
  assign n3389 = ( n1875 & n3387 ) | ( n1875 & ~n3388 ) | ( n3387 & ~n3388 ) ;
  assign n3390 = n3365 & n3389 ;
  assign n3391 = x167 & ~n754 ;
  assign n3392 = x41 | n769 ;
  assign n3393 = ~n354 & n3392 ;
  assign n3394 = ( ~n415 & n2197 ) | ( ~n415 & n3393 ) | ( n2197 & n3393 ) ;
  assign n3395 = ( n408 & ~n417 ) | ( n408 & n3394 ) | ( ~n417 & n3394 ) ;
  assign n3396 = ( n1891 & ~n1896 ) | ( n1891 & n3395 ) | ( ~n1896 & n3395 ) ;
  assign n3397 = ( ~n445 & n461 ) | ( ~n445 & n3396 ) | ( n461 & n3396 ) ;
  assign n3398 = ( n1910 & ~n2216 ) | ( n1910 & n3397 ) | ( ~n2216 & n3397 ) ;
  assign n3399 = ( ~n1522 & n1531 ) | ( ~n1522 & n3398 ) | ( n1531 & n3398 ) ;
  assign n3400 = ( n550 & ~n2495 ) | ( n550 & n3399 ) | ( ~n2495 & n3399 ) ;
  assign n3401 = ( ~n2255 & n2510 ) | ( ~n2255 & n3400 ) | ( n2510 & n3400 ) ;
  assign n3402 = ( n1951 & ~n2271 ) | ( n1951 & n3401 ) | ( ~n2271 & n3401 ) ;
  assign n3403 = ( n2919 & ~n3009 ) | ( n2919 & n3402 ) | ( ~n3009 & n3402 ) ;
  assign n3404 = ~n705 & n2928 ;
  assign n3405 = n716 | n3404 ;
  assign n3406 = ~n702 & n3405 ;
  assign n3407 = ( ~n731 & n735 ) | ( ~n731 & n3406 ) | ( n735 & n3406 ) ;
  assign n3408 = n738 | n3407 ;
  assign n3409 = ( ~n716 & n1602 ) | ( ~n716 & n2926 ) | ( n1602 & n2926 ) ;
  assign n3410 = n702 | n3409 ;
  assign n3411 = ~n734 & n3410 ;
  assign n3412 = ( ~n738 & n746 ) | ( ~n738 & n3411 ) | ( n746 & n3411 ) ;
  assign n3413 = ( n3403 & n3408 ) | ( n3403 & ~n3412 ) | ( n3408 & ~n3412 ) ;
  assign n3414 = ~n766 & n1617 ;
  assign n3415 = ( n1984 & n3413 ) | ( n1984 & ~n3414 ) | ( n3413 & ~n3414 ) ;
  assign n3416 = n3391 & n3415 ;
  assign n3417 = x168 & ~n1151 ;
  assign n3418 = x42 | n1166 ;
  assign n3419 = ~n752 & n3418 ;
  assign n3420 = ( ~n813 & n2293 ) | ( ~n813 & n3419 ) | ( n2293 & n3419 ) ;
  assign n3421 = ( n806 & ~n815 ) | ( n806 & n3420 ) | ( ~n815 & n3420 ) ;
  assign n3422 = ( n2000 & ~n2005 ) | ( n2000 & n3421 ) | ( ~n2005 & n3421 ) ;
  assign n3423 = ( ~n843 & n859 ) | ( ~n843 & n3422 ) | ( n859 & n3422 ) ;
  assign n3424 = ( n2019 & ~n2312 ) | ( n2019 & n3423 ) | ( ~n2312 & n3423 ) ;
  assign n3425 = ( ~n1661 & n1670 ) | ( ~n1661 & n3424 ) | ( n1670 & n3424 ) ;
  assign n3426 = ( n948 & ~n2564 ) | ( n948 & n3425 ) | ( ~n2564 & n3425 ) ;
  assign n3427 = ( ~n2351 & n2579 ) | ( ~n2351 & n3426 ) | ( n2579 & n3426 ) ;
  assign n3428 = ( n2060 & ~n2367 ) | ( n2060 & n3427 ) | ( ~n2367 & n3427 ) ;
  assign n3429 = ( n2948 & ~n3038 ) | ( n2948 & n3428 ) | ( ~n3038 & n3428 ) ;
  assign n3430 = ~n1102 & n2957 ;
  assign n3431 = n1113 | n3430 ;
  assign n3432 = ~n1099 & n3431 ;
  assign n3433 = ( ~n1128 & n1132 ) | ( ~n1128 & n3432 ) | ( n1132 & n3432 ) ;
  assign n3434 = n1135 | n3433 ;
  assign n3435 = ( ~n1113 & n1740 ) | ( ~n1113 & n2955 ) | ( n1740 & n2955 ) ;
  assign n3436 = n1099 | n3435 ;
  assign n3437 = ~n1131 & n3436 ;
  assign n3438 = ( ~n1135 & n1143 ) | ( ~n1135 & n3437 ) | ( n1143 & n3437 ) ;
  assign n3439 = ( n3429 & n3434 ) | ( n3429 & ~n3438 ) | ( n3434 & ~n3438 ) ;
  assign n3440 = ~n1163 & n1755 ;
  assign n3441 = ( n2093 & n3439 ) | ( n2093 & ~n3440 ) | ( n3439 & ~n3440 ) ;
  assign n3442 = n3417 & n3441 ;
  assign n3443 = x169 & ~n353 ;
  assign n3444 = x43 | n376 ;
  assign n3445 = ~n1149 & n3444 ;
  assign n3446 = ( ~n1210 & n2389 ) | ( ~n1210 & n3445 ) | ( n2389 & n3445 ) ;
  assign n3447 = ( n1203 & ~n1212 ) | ( n1203 & n3446 ) | ( ~n1212 & n3446 ) ;
  assign n3448 = ( n2109 & ~n2114 ) | ( n2109 & n3447 ) | ( ~n2114 & n3447 ) ;
  assign n3449 = ( ~n1240 & n1256 ) | ( ~n1240 & n3448 ) | ( n1256 & n3448 ) ;
  assign n3450 = ( n2128 & ~n2408 ) | ( n2128 & n3449 ) | ( ~n2408 & n3449 ) ;
  assign n3451 = ( ~n1799 & n1808 ) | ( ~n1799 & n3450 ) | ( n1808 & n3450 ) ;
  assign n3452 = ( n1345 & ~n2633 ) | ( n1345 & n3451 ) | ( ~n2633 & n3451 ) ;
  assign n3453 = ( ~n2447 & n2648 ) | ( ~n2447 & n3452 ) | ( n2648 & n3452 ) ;
  assign n3454 = ( n2169 & ~n2463 ) | ( n2169 & n3453 ) | ( ~n2463 & n3453 ) ;
  assign n3455 = ( n2977 & ~n3067 ) | ( n2977 & n3454 ) | ( ~n3067 & n3454 ) ;
  assign n3456 = ~n304 & n2986 ;
  assign n3457 = n336 | n3456 ;
  assign n3458 = ~n333 & n3457 ;
  assign n3459 = ( ~n330 & n1471 ) | ( ~n330 & n3458 ) | ( n1471 & n3458 ) ;
  assign n3460 = n345 | n3459 ;
  assign n3461 = ( ~n336 & n1464 ) | ( ~n336 & n2984 ) | ( n1464 & n2984 ) ;
  assign n3462 = n333 | n3461 ;
  assign n3463 = ~n340 & n3462 ;
  assign n3464 = ( ~n345 & n349 ) | ( ~n345 & n3463 ) | ( n349 & n3463 ) ;
  assign n3465 = ( n3455 & n3460 ) | ( n3455 & ~n3464 ) | ( n3460 & ~n3464 ) ;
  assign n3466 = ~n373 & n1878 ;
  assign n3467 = ( n374 & n3465 ) | ( n374 & ~n3466 ) | ( n3465 & ~n3466 ) ;
  assign n3468 = n3443 & n3467 ;
  assign n3469 = x170 & ~n751 ;
  assign n3470 = x44 | n774 ;
  assign n3471 = ~n414 & n3470 ;
  assign n3472 = ( ~n403 & n407 ) | ( ~n403 & n3471 ) | ( n407 & n3471 ) ;
  assign n3473 = ( n1492 & ~n1497 ) | ( n1492 & n3472 ) | ( ~n1497 & n3472 ) ;
  assign n3474 = ( n2205 & ~n2210 ) | ( n2205 & n3473 ) | ( ~n2210 & n3473 ) ;
  assign n3475 = ( ~n1506 & n1513 ) | ( ~n1506 & n3474 ) | ( n1513 & n3474 ) ;
  assign n3476 = ( n2224 & ~n2487 ) | ( n2224 & n3475 ) | ( ~n2487 & n3475 ) ;
  assign n3477 = ( ~n1916 & n1924 ) | ( ~n1916 & n3476 ) | ( n1924 & n3476 ) ;
  assign n3478 = ( ~n564 & n1540 ) | ( ~n564 & n3477 ) | ( n1540 & n3477 ) ;
  assign n3479 = ( ~n2517 & n2698 ) | ( ~n2517 & n3478 ) | ( n2698 & n3478 ) ;
  assign n3480 = ( n2265 & ~n2532 ) | ( n2265 & n3479 ) | ( ~n2532 & n3479 ) ;
  assign n3481 = ( n3006 & ~n3094 ) | ( n3006 & n3480 ) | ( ~n3094 & n3480 ) ;
  assign n3482 = ~n702 & n3015 ;
  assign n3483 = n734 | n3482 ;
  assign n3484 = ~n731 & n3483 ;
  assign n3485 = ( ~n728 & n1610 ) | ( ~n728 & n3484 ) | ( n1610 & n3484 ) ;
  assign n3486 = n743 | n3485 ;
  assign n3487 = ( ~n734 & n1603 ) | ( ~n734 & n3013 ) | ( n1603 & n3013 ) ;
  assign n3488 = n731 | n3487 ;
  assign n3489 = ~n738 & n3488 ;
  assign n3490 = ( ~n743 & n747 ) | ( ~n743 & n3489 ) | ( n747 & n3489 ) ;
  assign n3491 = ( n3481 & n3486 ) | ( n3481 & ~n3490 ) | ( n3486 & ~n3490 ) ;
  assign n3492 = ~n771 & n1987 ;
  assign n3493 = ( n772 & n3491 ) | ( n772 & ~n3492 ) | ( n3491 & ~n3492 ) ;
  assign n3494 = n3469 & n3493 ;
  assign n3495 = x171 & ~n1148 ;
  assign n3496 = x45 | n1171 ;
  assign n3497 = ~n812 & n3496 ;
  assign n3498 = ( ~n801 & n805 ) | ( ~n801 & n3497 ) | ( n805 & n3497 ) ;
  assign n3499 = ( n1631 & ~n1636 ) | ( n1631 & n3498 ) | ( ~n1636 & n3498 ) ;
  assign n3500 = ( n2301 & ~n2306 ) | ( n2301 & n3499 ) | ( ~n2306 & n3499 ) ;
  assign n3501 = ( ~n1645 & n1652 ) | ( ~n1645 & n3500 ) | ( n1652 & n3500 ) ;
  assign n3502 = ( n2320 & ~n2556 ) | ( n2320 & n3501 ) | ( ~n2556 & n3501 ) ;
  assign n3503 = ( ~n2025 & n2033 ) | ( ~n2025 & n3502 ) | ( n2033 & n3502 ) ;
  assign n3504 = ( ~n962 & n1679 ) | ( ~n962 & n3503 ) | ( n1679 & n3503 ) ;
  assign n3505 = ( ~n2586 & n2742 ) | ( ~n2586 & n3504 ) | ( n2742 & n3504 ) ;
  assign n3506 = ( n2361 & ~n2601 ) | ( n2361 & n3505 ) | ( ~n2601 & n3505 ) ;
  assign n3507 = ( n3035 & ~n3121 ) | ( n3035 & n3506 ) | ( ~n3121 & n3506 ) ;
  assign n3508 = ~n1099 & n3044 ;
  assign n3509 = n1131 | n3508 ;
  assign n3510 = ~n1128 & n3509 ;
  assign n3511 = ( ~n1125 & n1748 ) | ( ~n1125 & n3510 ) | ( n1748 & n3510 ) ;
  assign n3512 = n1140 | n3511 ;
  assign n3513 = ( ~n1131 & n1741 ) | ( ~n1131 & n3042 ) | ( n1741 & n3042 ) ;
  assign n3514 = n1128 | n3513 ;
  assign n3515 = ~n1135 & n3514 ;
  assign n3516 = ( ~n1140 & n1144 ) | ( ~n1140 & n3515 ) | ( n1144 & n3515 ) ;
  assign n3517 = ( n3507 & n3512 ) | ( n3507 & ~n3516 ) | ( n3512 & ~n3516 ) ;
  assign n3518 = ~n1168 & n2096 ;
  assign n3519 = ( n1169 & n3517 ) | ( n1169 & ~n3518 ) | ( n3517 & ~n3518 ) ;
  assign n3520 = n3495 & n3519 ;
  assign n3521 = x172 & ~n413 ;
  assign n3522 = x46 | n404 ;
  assign n3523 = ~n1209 & n3522 ;
  assign n3524 = ( ~n1198 & n1202 ) | ( ~n1198 & n3523 ) | ( n1202 & n3523 ) ;
  assign n3525 = ( n1769 & ~n1774 ) | ( n1769 & n3524 ) | ( ~n1774 & n3524 ) ;
  assign n3526 = ( n2397 & ~n2402 ) | ( n2397 & n3525 ) | ( ~n2402 & n3525 ) ;
  assign n3527 = ( ~n1783 & n1790 ) | ( ~n1783 & n3526 ) | ( n1790 & n3526 ) ;
  assign n3528 = ( n2416 & ~n2625 ) | ( n2416 & n3527 ) | ( ~n2625 & n3527 ) ;
  assign n3529 = ( ~n2134 & n2142 ) | ( ~n2134 & n3528 ) | ( n2142 & n3528 ) ;
  assign n3530 = ( ~n1359 & n1817 ) | ( ~n1359 & n3529 ) | ( n1817 & n3529 ) ;
  assign n3531 = ( ~n2655 & n2786 ) | ( ~n2655 & n3530 ) | ( n2786 & n3530 ) ;
  assign n3532 = ( n2457 & ~n2670 ) | ( n2457 & n3531 ) | ( ~n2670 & n3531 ) ;
  assign n3533 = ( n3064 & ~n3148 ) | ( n3064 & n3532 ) | ( ~n3148 & n3532 ) ;
  assign n3534 = ~n333 & n3071 ;
  assign n3535 = n340 | n3534 ;
  assign n3536 = ~n330 & n3535 ;
  assign n3537 = ( ~n327 & n1872 ) | ( ~n327 & n3536 ) | ( n1872 & n3536 ) ;
  assign n3538 = n364 | n3537 ;
  assign n3539 = ( ~n340 & n348 ) | ( ~n340 & n3070 ) | ( n348 & n3070 ) ;
  assign n3540 = n330 | n3539 ;
  assign n3541 = ~n345 & n3540 ;
  assign n3542 = ( ~n364 & n1476 ) | ( ~n364 & n3541 ) | ( n1476 & n3541 ) ;
  assign n3543 = ( n3533 & n3538 ) | ( n3533 & ~n3542 ) | ( n3538 & ~n3542 ) ;
  assign n3544 = ( ~n384 & n1483 ) | ( ~n384 & n3543 ) | ( n1483 & n3543 ) ;
  assign n3545 = n3521 & n3544 ;
  assign n3546 = x173 & ~n811 ;
  assign n3547 = x47 | n802 ;
  assign n3548 = ~n402 & n3547 ;
  assign n3549 = ( ~n397 & n1491 ) | ( ~n397 & n3548 ) | ( n1491 & n3548 ) ;
  assign n3550 = ( ~n421 & n1891 ) | ( ~n421 & n3549 ) | ( n1891 & n3549 ) ;
  assign n3551 = ( ~n444 & n460 ) | ( ~n444 & n3550 ) | ( n460 & n3550 ) ;
  assign n3552 = ( ~n1902 & n1908 ) | ( ~n1902 & n3551 ) | ( n1908 & n3551 ) ;
  assign n3553 = ( ~n494 & n509 ) | ( ~n494 & n3552 ) | ( n509 & n3552 ) ;
  assign n3554 = ( ~n2230 & n2238 ) | ( ~n2230 & n3553 ) | ( n2238 & n3553 ) ;
  assign n3555 = ( ~n1550 & n1933 ) | ( ~n1550 & n3554 ) | ( n1933 & n3554 ) ;
  assign n3556 = ( n604 & ~n621 ) | ( n604 & n3555 ) | ( ~n621 & n3555 ) ;
  assign n3557 = ( n2526 & ~n2714 ) | ( n2526 & n3556 ) | ( ~n2714 & n3556 ) ;
  assign n3558 = ( n3091 & ~n3175 ) | ( n3091 & n3557 ) | ( ~n3175 & n3557 ) ;
  assign n3559 = ~n731 & n3098 ;
  assign n3560 = n738 | n3559 ;
  assign n3561 = ~n728 & n3560 ;
  assign n3562 = ( ~n725 & n1981 ) | ( ~n725 & n3561 ) | ( n1981 & n3561 ) ;
  assign n3563 = n762 | n3562 ;
  assign n3564 = ( ~n738 & n746 ) | ( ~n738 & n3097 ) | ( n746 & n3097 ) ;
  assign n3565 = n728 | n3564 ;
  assign n3566 = ~n743 & n3565 ;
  assign n3567 = ( ~n762 & n1615 ) | ( ~n762 & n3566 ) | ( n1615 & n3566 ) ;
  assign n3568 = ( n3558 & n3563 ) | ( n3558 & ~n3567 ) | ( n3563 & ~n3567 ) ;
  assign n3569 = ( ~n782 & n1622 ) | ( ~n782 & n3568 ) | ( n1622 & n3568 ) ;
  assign n3570 = n3546 & n3569 ;
  assign n3571 = x174 & ~n1208 ;
  assign n3572 = x48 | n1199 ;
  assign n3573 = ~n800 & n3572 ;
  assign n3574 = ( ~n795 & n1630 ) | ( ~n795 & n3573 ) | ( n1630 & n3573 ) ;
  assign n3575 = ( ~n819 & n2000 ) | ( ~n819 & n3574 ) | ( n2000 & n3574 ) ;
  assign n3576 = ( ~n842 & n858 ) | ( ~n842 & n3575 ) | ( n858 & n3575 ) ;
  assign n3577 = ( ~n2011 & n2017 ) | ( ~n2011 & n3576 ) | ( n2017 & n3576 ) ;
  assign n3578 = ( ~n892 & n907 ) | ( ~n892 & n3577 ) | ( n907 & n3577 ) ;
  assign n3579 = ( ~n2326 & n2334 ) | ( ~n2326 & n3578 ) | ( n2334 & n3578 ) ;
  assign n3580 = ( ~n1689 & n2042 ) | ( ~n1689 & n3579 ) | ( n2042 & n3579 ) ;
  assign n3581 = ( n1002 & ~n1019 ) | ( n1002 & n3580 ) | ( ~n1019 & n3580 ) ;
  assign n3582 = ( n2595 & ~n2758 ) | ( n2595 & n3581 ) | ( ~n2758 & n3581 ) ;
  assign n3583 = ( n3118 & ~n3202 ) | ( n3118 & n3582 ) | ( ~n3202 & n3582 ) ;
  assign n3584 = ~n1128 & n3125 ;
  assign n3585 = n1135 | n3584 ;
  assign n3586 = ~n1125 & n3585 ;
  assign n3587 = ( ~n1122 & n2090 ) | ( ~n1122 & n3586 ) | ( n2090 & n3586 ) ;
  assign n3588 = n1159 | n3587 ;
  assign n3589 = ( ~n1135 & n1143 ) | ( ~n1135 & n3124 ) | ( n1143 & n3124 ) ;
  assign n3590 = n1125 | n3589 ;
  assign n3591 = ~n1140 & n3590 ;
  assign n3592 = ( ~n1159 & n1753 ) | ( ~n1159 & n3591 ) | ( n1753 & n3591 ) ;
  assign n3593 = ( n3583 & n3588 ) | ( n3583 & ~n3592 ) | ( n3588 & ~n3592 ) ;
  assign n3594 = ( ~n1179 & n1760 ) | ( ~n1179 & n3593 ) | ( n1760 & n3593 ) ;
  assign n3595 = n3571 & n3594 ;
  assign n3596 = x175 & ~n401 ;
  assign n3597 = x49 | n398 ;
  assign n3598 = ~n1197 & n3597 ;
  assign n3599 = ( ~n1192 & n1768 ) | ( ~n1192 & n3598 ) | ( n1768 & n3598 ) ;
  assign n3600 = ( ~n1216 & n2109 ) | ( ~n1216 & n3599 ) | ( n2109 & n3599 ) ;
  assign n3601 = ( ~n1239 & n1255 ) | ( ~n1239 & n3600 ) | ( n1255 & n3600 ) ;
  assign n3602 = ( ~n2120 & n2126 ) | ( ~n2120 & n3601 ) | ( n2126 & n3601 ) ;
  assign n3603 = ( ~n1289 & n1304 ) | ( ~n1289 & n3602 ) | ( n1304 & n3602 ) ;
  assign n3604 = ( ~n2422 & n2430 ) | ( ~n2422 & n3603 ) | ( n2430 & n3603 ) ;
  assign n3605 = ( ~n1827 & n2151 ) | ( ~n1827 & n3604 ) | ( n2151 & n3604 ) ;
  assign n3606 = ( n1399 & ~n1416 ) | ( n1399 & n3605 ) | ( ~n1416 & n3605 ) ;
  assign n3607 = ( n2664 & ~n2802 ) | ( n2664 & n3606 ) | ( ~n2802 & n3606 ) ;
  assign n3608 = ( n3145 & ~n3229 ) | ( n3145 & n3607 ) | ( ~n3229 & n3607 ) ;
  assign n3609 = ~n330 & n3152 ;
  assign n3610 = n345 | n3609 ;
  assign n3611 = ~n327 & n3610 ;
  assign n3612 = ( ~n361 & n365 ) | ( ~n361 & n3611 ) | ( n365 & n3611 ) ;
  assign n3613 = n368 | n3612 ;
  assign n3614 = ( ~n345 & n349 ) | ( ~n345 & n3151 ) | ( n349 & n3151 ) ;
  assign n3615 = n327 | n3614 ;
  assign n3616 = ~n364 & n3615 ;
  assign n3617 = ( ~n368 & n380 ) | ( ~n368 & n3616 ) | ( n380 & n3616 ) ;
  assign n3618 = ( n3608 & n3613 ) | ( n3608 & ~n3617 ) | ( n3613 & ~n3617 ) ;
  assign n3619 = ( ~n1489 & n1883 ) | ( ~n1489 & n3618 ) | ( n1883 & n3618 ) ;
  assign n3620 = n3596 & n3619 ;
  assign n3621 = x176 & ~n799 ;
  assign n3622 = x50 | n796 ;
  assign n3623 = ~n396 & n3622 ;
  assign n3624 = ( ~n391 & n1890 ) | ( ~n391 & n3623 ) | ( n1890 & n3623 ) ;
  assign n3625 = ( ~n439 & n2205 ) | ( ~n439 & n3624 ) | ( n2205 & n3624 ) ;
  assign n3626 = ( ~n1505 & n1512 ) | ( ~n1505 & n3625 ) | ( n1512 & n3625 ) ;
  assign n3627 = ( ~n2216 & n2222 ) | ( ~n2216 & n3626 ) | ( n2222 & n3626 ) ;
  assign n3628 = ( ~n1521 & n1530 ) | ( ~n1521 & n3627 ) | ( n1530 & n3627 ) ;
  assign n3629 = ( ~n2494 & n2501 ) | ( ~n2494 & n3628 ) | ( n2501 & n3628 ) ;
  assign n3630 = ( ~n1940 & n2247 ) | ( ~n1940 & n3629 ) | ( n2247 & n3629 ) ;
  assign n3631 = ( n1560 & ~n1570 ) | ( n1560 & n3630 ) | ( ~n1570 & n3630 ) ;
  assign n3632 = ( n2708 & ~n2832 ) | ( n2708 & n3631 ) | ( ~n2832 & n3631 ) ;
  assign n3633 = ( n3172 & ~n3255 ) | ( n3172 & n3632 ) | ( ~n3255 & n3632 ) ;
  assign n3634 = ~n728 & n3179 ;
  assign n3635 = n743 | n3634 ;
  assign n3636 = ~n725 & n3635 ;
  assign n3637 = ( ~n759 & n763 ) | ( ~n759 & n3636 ) | ( n763 & n3636 ) ;
  assign n3638 = n766 | n3637 ;
  assign n3639 = ( ~n743 & n747 ) | ( ~n743 & n3178 ) | ( n747 & n3178 ) ;
  assign n3640 = n725 | n3639 ;
  assign n3641 = ~n762 & n3640 ;
  assign n3642 = ( ~n766 & n778 ) | ( ~n766 & n3641 ) | ( n778 & n3641 ) ;
  assign n3643 = ( n3633 & n3638 ) | ( n3633 & ~n3642 ) | ( n3638 & ~n3642 ) ;
  assign n3644 = ( ~n1628 & n1992 ) | ( ~n1628 & n3643 ) | ( n1992 & n3643 ) ;
  assign n3645 = n3621 & n3644 ;
  assign n3646 = x177 & ~n1196 ;
  assign n3647 = x51 | n1193 ;
  assign n3648 = ~n794 & n3647 ;
  assign n3649 = ( ~n789 & n1999 ) | ( ~n789 & n3648 ) | ( n1999 & n3648 ) ;
  assign n3650 = ( ~n837 & n2301 ) | ( ~n837 & n3649 ) | ( n2301 & n3649 ) ;
  assign n3651 = ( ~n1644 & n1651 ) | ( ~n1644 & n3650 ) | ( n1651 & n3650 ) ;
  assign n3652 = ( ~n2312 & n2318 ) | ( ~n2312 & n3651 ) | ( n2318 & n3651 ) ;
  assign n3653 = ( ~n1660 & n1669 ) | ( ~n1660 & n3652 ) | ( n1669 & n3652 ) ;
  assign n3654 = ( ~n2563 & n2570 ) | ( ~n2563 & n3653 ) | ( n2570 & n3653 ) ;
  assign n3655 = ( ~n2049 & n2343 ) | ( ~n2049 & n3654 ) | ( n2343 & n3654 ) ;
  assign n3656 = ( n1699 & ~n1709 ) | ( n1699 & n3655 ) | ( ~n1709 & n3655 ) ;
  assign n3657 = ( n2752 & ~n2862 ) | ( n2752 & n3656 ) | ( ~n2862 & n3656 ) ;
  assign n3658 = ( n3199 & ~n3281 ) | ( n3199 & n3657 ) | ( ~n3281 & n3657 ) ;
  assign n3659 = ~n1125 & n3206 ;
  assign n3660 = n1140 | n3659 ;
  assign n3661 = ~n1122 & n3660 ;
  assign n3662 = ( ~n1156 & n1160 ) | ( ~n1156 & n3661 ) | ( n1160 & n3661 ) ;
  assign n3663 = n1163 | n3662 ;
  assign n3664 = ( ~n1140 & n1144 ) | ( ~n1140 & n3205 ) | ( n1144 & n3205 ) ;
  assign n3665 = n1122 | n3664 ;
  assign n3666 = ~n1159 & n3665 ;
  assign n3667 = ( ~n1163 & n1175 ) | ( ~n1163 & n3666 ) | ( n1175 & n3666 ) ;
  assign n3668 = ( n3658 & n3663 ) | ( n3658 & ~n3667 ) | ( n3663 & ~n3667 ) ;
  assign n3669 = ( ~n1766 & n2101 ) | ( ~n1766 & n3668 ) | ( n2101 & n3668 ) ;
  assign n3670 = n3646 & n3669 ;
  assign n3671 = x178 & ~n395 ;
  assign n3672 = x52 | n392 ;
  assign n3673 = ~n1191 & n3672 ;
  assign n3674 = ( ~n1186 & n2108 ) | ( ~n1186 & n3673 ) | ( n2108 & n3673 ) ;
  assign n3675 = ( ~n1234 & n2397 ) | ( ~n1234 & n3674 ) | ( n2397 & n3674 ) ;
  assign n3676 = ( ~n1782 & n1789 ) | ( ~n1782 & n3675 ) | ( n1789 & n3675 ) ;
  assign n3677 = ( ~n2408 & n2414 ) | ( ~n2408 & n3676 ) | ( n2414 & n3676 ) ;
  assign n3678 = ( ~n1798 & n1807 ) | ( ~n1798 & n3677 ) | ( n1807 & n3677 ) ;
  assign n3679 = ( ~n2632 & n2639 ) | ( ~n2632 & n3678 ) | ( n2639 & n3678 ) ;
  assign n3680 = ( ~n2158 & n2439 ) | ( ~n2158 & n3679 ) | ( n2439 & n3679 ) ;
  assign n3681 = ( n1837 & ~n1847 ) | ( n1837 & n3680 ) | ( ~n1847 & n3680 ) ;
  assign n3682 = ( n2796 & ~n2892 ) | ( n2796 & n3681 ) | ( ~n2892 & n3681 ) ;
  assign n3683 = ( n3226 & ~n3307 ) | ( n3226 & n3682 ) | ( ~n3307 & n3682 ) ;
  assign n3684 = n347 | n364 ;
  assign n3685 = ~n361 & n3684 ;
  assign n3686 = ( ~n358 & n1480 ) | ( ~n358 & n3685 ) | ( n1480 & n3685 ) ;
  assign n3687 = n373 | n3686 ;
  assign n3688 = ( ~n364 & n1476 ) | ( ~n364 & n3232 ) | ( n1476 & n3232 ) ;
  assign n3689 = n361 | n3688 ;
  assign n3690 = ~n368 & n3689 ;
  assign n3691 = ( ~n373 & n381 ) | ( ~n373 & n3690 ) | ( n381 & n3690 ) ;
  assign n3692 = ( n3683 & n3687 ) | ( n3683 & ~n3691 ) | ( n3687 & ~n3691 ) ;
  assign n3693 = ( ~n1888 & n2200 ) | ( ~n1888 & n3692 ) | ( n2200 & n3692 ) ;
  assign n3694 = n3671 & n3693 ;
  assign n3695 = x179 & ~n793 ;
  assign n3696 = x53 | n790 ;
  assign n3697 = ~n390 & n3696 ;
  assign n3698 = ( ~n435 & n2204 ) | ( ~n435 & n3697 ) | ( n2204 & n3697 ) ;
  assign n3699 = ( n460 & ~n1503 ) | ( n460 & n3698 ) | ( ~n1503 & n3698 ) ;
  assign n3700 = ( ~n1901 & n1907 ) | ( ~n1901 & n3699 ) | ( n1907 & n3699 ) ;
  assign n3701 = ( n507 & ~n2487 ) | ( n507 & n3700 ) | ( ~n2487 & n3700 ) ;
  assign n3702 = ( ~n1915 & n1923 ) | ( ~n1915 & n3701 ) | ( n1923 & n3701 ) ;
  assign n3703 = ( n550 & ~n562 ) | ( n550 & n3702 ) | ( ~n562 & n3702 ) ;
  assign n3704 = ( ~n2254 & n2509 ) | ( ~n2254 & n3703 ) | ( n2509 & n3703 ) ;
  assign n3705 = ( n1950 & ~n1957 ) | ( n1950 & n3704 ) | ( ~n1957 & n3704 ) ;
  assign n3706 = ( n2829 & ~n2921 ) | ( n2829 & n3705 ) | ( ~n2921 & n3705 ) ;
  assign n3707 = ( n3252 & ~n3333 ) | ( n3252 & n3706 ) | ( ~n3333 & n3706 ) ;
  assign n3708 = n745 | n762 ;
  assign n3709 = ~n759 & n3708 ;
  assign n3710 = ( ~n756 & n1619 ) | ( ~n756 & n3709 ) | ( n1619 & n3709 ) ;
  assign n3711 = n771 | n3710 ;
  assign n3712 = ( ~n762 & n1615 ) | ( ~n762 & n3258 ) | ( n1615 & n3258 ) ;
  assign n3713 = n759 | n3712 ;
  assign n3714 = ~n766 & n3713 ;
  assign n3715 = ( ~n771 & n779 ) | ( ~n771 & n3714 ) | ( n779 & n3714 ) ;
  assign n3716 = ( n3707 & n3711 ) | ( n3707 & ~n3715 ) | ( n3711 & ~n3715 ) ;
  assign n3717 = ( ~n1997 & n2296 ) | ( ~n1997 & n3716 ) | ( n2296 & n3716 ) ;
  assign n3718 = n3695 & n3717 ;
  assign n3719 = x180 & ~n1190 ;
  assign n3720 = x54 | n1187 ;
  assign n3721 = ~n788 & n3720 ;
  assign n3722 = ( ~n833 & n2300 ) | ( ~n833 & n3721 ) | ( n2300 & n3721 ) ;
  assign n3723 = ( n858 & ~n1642 ) | ( n858 & n3722 ) | ( ~n1642 & n3722 ) ;
  assign n3724 = ( ~n2010 & n2016 ) | ( ~n2010 & n3723 ) | ( n2016 & n3723 ) ;
  assign n3725 = ( n905 & ~n2556 ) | ( n905 & n3724 ) | ( ~n2556 & n3724 ) ;
  assign n3726 = ( ~n2024 & n2032 ) | ( ~n2024 & n3725 ) | ( n2032 & n3725 ) ;
  assign n3727 = ( n948 & ~n960 ) | ( n948 & n3726 ) | ( ~n960 & n3726 ) ;
  assign n3728 = ( ~n2350 & n2578 ) | ( ~n2350 & n3727 ) | ( n2578 & n3727 ) ;
  assign n3729 = ( n2059 & ~n2066 ) | ( n2059 & n3728 ) | ( ~n2066 & n3728 ) ;
  assign n3730 = ( n2859 & ~n2950 ) | ( n2859 & n3729 ) | ( ~n2950 & n3729 ) ;
  assign n3731 = ( n3278 & ~n3359 ) | ( n3278 & n3730 ) | ( ~n3359 & n3730 ) ;
  assign n3732 = n1142 | n1159 ;
  assign n3733 = ~n1156 & n3732 ;
  assign n3734 = ( ~n1153 & n1757 ) | ( ~n1153 & n3733 ) | ( n1757 & n3733 ) ;
  assign n3735 = n1168 | n3734 ;
  assign n3736 = ( ~n1159 & n1753 ) | ( ~n1159 & n3284 ) | ( n1753 & n3284 ) ;
  assign n3737 = n1156 | n3736 ;
  assign n3738 = ~n1163 & n3737 ;
  assign n3739 = ( ~n1168 & n1176 ) | ( ~n1168 & n3738 ) | ( n1176 & n3738 ) ;
  assign n3740 = ( n3731 & n3735 ) | ( n3731 & ~n3739 ) | ( n3735 & ~n3739 ) ;
  assign n3741 = ( ~n2106 & n2392 ) | ( ~n2106 & n3740 ) | ( n2392 & n3740 ) ;
  assign n3742 = n3719 & n3741 ;
  assign n3743 = x181 & ~n389 ;
  assign n3744 = x55 | n386 ;
  assign n3745 = ~n1185 & n3744 ;
  assign n3746 = ( ~n1230 & n2396 ) | ( ~n1230 & n3745 ) | ( n2396 & n3745 ) ;
  assign n3747 = ( n1255 & ~n1780 ) | ( n1255 & n3746 ) | ( ~n1780 & n3746 ) ;
  assign n3748 = ( ~n2119 & n2125 ) | ( ~n2119 & n3747 ) | ( n2125 & n3747 ) ;
  assign n3749 = ( n1302 & ~n2625 ) | ( n1302 & n3748 ) | ( ~n2625 & n3748 ) ;
  assign n3750 = ( ~n2133 & n2141 ) | ( ~n2133 & n3749 ) | ( n2141 & n3749 ) ;
  assign n3751 = ( n1345 & ~n1357 ) | ( n1345 & n3750 ) | ( ~n1357 & n3750 ) ;
  assign n3752 = ( ~n2446 & n2647 ) | ( ~n2446 & n3751 ) | ( n2647 & n3751 ) ;
  assign n3753 = ( n2168 & ~n2175 ) | ( n2168 & n3752 ) | ( ~n2175 & n3752 ) ;
  assign n3754 = ( n2889 & ~n2979 ) | ( n2889 & n3753 ) | ( ~n2979 & n3753 ) ;
  assign n3755 = ( n3304 & ~n3385 ) | ( n3304 & n3754 ) | ( ~n3385 & n3754 ) ;
  assign n3756 = n368 | n1475 ;
  assign n3757 = ~n358 & n3756 ;
  assign n3758 = ( ~n355 & n1880 ) | ( ~n355 & n3757 ) | ( n1880 & n3757 ) ;
  assign n3759 = n378 | n3758 ;
  assign n3760 = ( ~n368 & n380 ) | ( ~n368 & n3310 ) | ( n380 & n3310 ) ;
  assign n3761 = n358 | n3760 ;
  assign n3762 = ~n373 & n3761 ;
  assign n3763 = ( ~n378 & n1486 ) | ( ~n378 & n3762 ) | ( n1486 & n3762 ) ;
  assign n3764 = ( n3755 & n3759 ) | ( n3755 & ~n3763 ) | ( n3759 & ~n3763 ) ;
  assign n3765 = ( n410 & ~n420 ) | ( n410 & n3764 ) | ( ~n420 & n3764 ) ;
  assign n3766 = n3743 & n3765 ;
  assign n3767 = x182 & ~n787 ;
  assign n3768 = x56 | n784 ;
  assign n3769 = ~n434 & n3768 ;
  assign n3770 = ( ~n432 & n459 ) | ( ~n432 & n3769 ) | ( n459 & n3769 ) ;
  assign n3771 = ( ~n1504 & n1512 ) | ( ~n1504 & n3770 ) | ( n1512 & n3770 ) ;
  assign n3772 = ( ~n2215 & n2221 ) | ( ~n2215 & n3771 ) | ( n2221 & n3771 ) ;
  assign n3773 = ( ~n494 & n1528 ) | ( ~n494 & n3772 ) | ( n1528 & n3772 ) ;
  assign n3774 = ( ~n2229 & n2237 ) | ( ~n2229 & n3773 ) | ( n2237 & n3773 ) ;
  assign n3775 = ( n1540 & ~n1548 ) | ( n1540 & n3774 ) | ( ~n1548 & n3774 ) ;
  assign n3776 = ( ~n2516 & n2697 ) | ( ~n2516 & n3775 ) | ( n2697 & n3775 ) ;
  assign n3777 = ( n2264 & ~n2271 ) | ( n2264 & n3776 ) | ( ~n2271 & n3776 ) ;
  assign n3778 = ( n2918 & ~n3008 ) | ( n2918 & n3777 ) | ( ~n3008 & n3777 ) ;
  assign n3779 = ( n3330 & ~n3411 ) | ( n3330 & n3778 ) | ( ~n3411 & n3778 ) ;
  assign n3780 = n766 | n1614 ;
  assign n3781 = ~n756 & n3780 ;
  assign n3782 = ( ~n753 & n1989 ) | ( ~n753 & n3781 ) | ( n1989 & n3781 ) ;
  assign n3783 = n776 | n3782 ;
  assign n3784 = ( ~n766 & n778 ) | ( ~n766 & n3336 ) | ( n778 & n3336 ) ;
  assign n3785 = n756 | n3784 ;
  assign n3786 = ~n771 & n3785 ;
  assign n3787 = ( ~n776 & n1625 ) | ( ~n776 & n3786 ) | ( n1625 & n3786 ) ;
  assign n3788 = ( n3779 & n3783 ) | ( n3779 & ~n3787 ) | ( n3783 & ~n3787 ) ;
  assign n3789 = ( n808 & ~n818 ) | ( n808 & n3788 ) | ( ~n818 & n3788 ) ;
  assign n3790 = n3767 & n3789 ;
  assign n3791 = x183 & ~n1184 ;
  assign n3792 = x57 | n1181 ;
  assign n3793 = ~n832 & n3792 ;
  assign n3794 = ( ~n830 & n857 ) | ( ~n830 & n3793 ) | ( n857 & n3793 ) ;
  assign n3795 = ( ~n1643 & n1651 ) | ( ~n1643 & n3794 ) | ( n1651 & n3794 ) ;
  assign n3796 = ( ~n2311 & n2317 ) | ( ~n2311 & n3795 ) | ( n2317 & n3795 ) ;
  assign n3797 = ( ~n892 & n1667 ) | ( ~n892 & n3796 ) | ( n1667 & n3796 ) ;
  assign n3798 = ( ~n2325 & n2333 ) | ( ~n2325 & n3797 ) | ( n2333 & n3797 ) ;
  assign n3799 = ( n1679 & ~n1687 ) | ( n1679 & n3798 ) | ( ~n1687 & n3798 ) ;
  assign n3800 = ( ~n2585 & n2741 ) | ( ~n2585 & n3799 ) | ( n2741 & n3799 ) ;
  assign n3801 = ( n2360 & ~n2367 ) | ( n2360 & n3800 ) | ( ~n2367 & n3800 ) ;
  assign n3802 = ( n2947 & ~n3037 ) | ( n2947 & n3801 ) | ( ~n3037 & n3801 ) ;
  assign n3803 = ( n3356 & ~n3437 ) | ( n3356 & n3802 ) | ( ~n3437 & n3802 ) ;
  assign n3804 = n1163 | n1752 ;
  assign n3805 = ~n1153 & n3804 ;
  assign n3806 = ( ~n1150 & n2098 ) | ( ~n1150 & n3805 ) | ( n2098 & n3805 ) ;
  assign n3807 = n1173 | n3806 ;
  assign n3808 = ( ~n1163 & n1175 ) | ( ~n1163 & n3362 ) | ( n1175 & n3362 ) ;
  assign n3809 = n1153 | n3808 ;
  assign n3810 = ~n1168 & n3809 ;
  assign n3811 = ( ~n1173 & n1763 ) | ( ~n1173 & n3810 ) | ( n1763 & n3810 ) ;
  assign n3812 = ( n3803 & n3807 ) | ( n3803 & ~n3811 ) | ( n3807 & ~n3811 ) ;
  assign n3813 = ( n1205 & ~n1215 ) | ( n1205 & n3812 ) | ( ~n1215 & n3812 ) ;
  assign n3814 = n3791 & n3813 ;
  assign n3815 = x184 & ~n433 ;
  assign n3816 = x58 | n436 ;
  assign n3817 = ~n1229 & n3816 ;
  assign n3818 = ( ~n1227 & n1254 ) | ( ~n1227 & n3817 ) | ( n1254 & n3817 ) ;
  assign n3819 = ( ~n1781 & n1789 ) | ( ~n1781 & n3818 ) | ( n1789 & n3818 ) ;
  assign n3820 = ( ~n2407 & n2413 ) | ( ~n2407 & n3819 ) | ( n2413 & n3819 ) ;
  assign n3821 = ( ~n1289 & n1805 ) | ( ~n1289 & n3820 ) | ( n1805 & n3820 ) ;
  assign n3822 = ( ~n2421 & n2429 ) | ( ~n2421 & n3821 ) | ( n2429 & n3821 ) ;
  assign n3823 = ( n1817 & ~n1825 ) | ( n1817 & n3822 ) | ( ~n1825 & n3822 ) ;
  assign n3824 = ( ~n2654 & n2785 ) | ( ~n2654 & n3823 ) | ( n2785 & n3823 ) ;
  assign n3825 = ( n2456 & ~n2463 ) | ( n2456 & n3824 ) | ( ~n2463 & n3824 ) ;
  assign n3826 = ( n2976 & ~n3066 ) | ( n2976 & n3825 ) | ( ~n3066 & n3825 ) ;
  assign n3827 = ( n3382 & ~n3463 ) | ( n3382 & n3826 ) | ( ~n3463 & n3826 ) ;
  assign n3828 = n373 | n1876 ;
  assign n3829 = ~n355 & n3828 ;
  assign n3830 = ( ~n415 & n2197 ) | ( ~n415 & n3829 ) | ( n2197 & n3829 ) ;
  assign n3831 = n406 | n3830 ;
  assign n3832 = ( ~n373 & n381 ) | ( ~n373 & n3388 ) | ( n381 & n3388 ) ;
  assign n3833 = n355 | n3832 ;
  assign n3834 = ~n378 & n3833 ;
  assign n3835 = ( ~n406 & n416 ) | ( ~n406 & n3834 ) | ( n416 & n3834 ) ;
  assign n3836 = ( n3827 & n3831 ) | ( n3827 & ~n3835 ) | ( n3831 & ~n3835 ) ;
  assign n3837 = ( n1494 & ~n1500 ) | ( n1494 & n3836 ) | ( ~n1500 & n3836 ) ;
  assign n3838 = n3815 & n3837 ;
  assign n3839 = x185 & ~n831 ;
  assign n3840 = x59 | n834 ;
  assign n3841 = ~n431 & n3840 ;
  assign n3842 = ( ~n429 & n1511 ) | ( ~n429 & n3841 ) | ( n1511 & n3841 ) ;
  assign n3843 = ( ~n456 & n1907 ) | ( ~n456 & n3842 ) | ( n1907 & n3842 ) ;
  assign n3844 = ( n506 & ~n2486 ) | ( n506 & n3843 ) | ( ~n2486 & n3843 ) ;
  assign n3845 = ( ~n1521 & n1921 ) | ( ~n1521 & n3844 ) | ( n1921 & n3844 ) ;
  assign n3846 = ( ~n2493 & n2500 ) | ( ~n2493 & n3845 ) | ( n2500 & n3845 ) ;
  assign n3847 = ( n1933 & ~n1939 ) | ( n1933 & n3846 ) | ( ~n1939 & n3846 ) ;
  assign n3848 = ( n603 & ~n620 ) | ( n603 & n3847 ) | ( ~n620 & n3847 ) ;
  assign n3849 = ( n2525 & ~n2532 ) | ( n2525 & n3848 ) | ( ~n2532 & n3848 ) ;
  assign n3850 = ( n3005 & ~n3093 ) | ( n3005 & n3849 ) | ( ~n3093 & n3849 ) ;
  assign n3851 = ( n3408 & ~n3489 ) | ( n3408 & n3850 ) | ( ~n3489 & n3850 ) ;
  assign n3852 = n771 | n1985 ;
  assign n3853 = ~n753 & n3852 ;
  assign n3854 = ( ~n813 & n2293 ) | ( ~n813 & n3853 ) | ( n2293 & n3853 ) ;
  assign n3855 = n804 | n3854 ;
  assign n3856 = ( ~n771 & n779 ) | ( ~n771 & n3414 ) | ( n779 & n3414 ) ;
  assign n3857 = n753 | n3856 ;
  assign n3858 = ~n776 & n3857 ;
  assign n3859 = ( ~n804 & n814 ) | ( ~n804 & n3858 ) | ( n814 & n3858 ) ;
  assign n3860 = ( n3851 & n3855 ) | ( n3851 & ~n3859 ) | ( n3855 & ~n3859 ) ;
  assign n3861 = ( n1633 & ~n1639 ) | ( n1633 & n3860 ) | ( ~n1639 & n3860 ) ;
  assign n3862 = n3839 & n3861 ;
  assign n3863 = x186 & ~n1228 ;
  assign n3864 = x60 | n1231 ;
  assign n3865 = ~n829 & n3864 ;
  assign n3866 = ( ~n827 & n1650 ) | ( ~n827 & n3865 ) | ( n1650 & n3865 ) ;
  assign n3867 = ( ~n854 & n2016 ) | ( ~n854 & n3866 ) | ( n2016 & n3866 ) ;
  assign n3868 = ( n904 & ~n2555 ) | ( n904 & n3867 ) | ( ~n2555 & n3867 ) ;
  assign n3869 = ( ~n1660 & n2030 ) | ( ~n1660 & n3868 ) | ( n2030 & n3868 ) ;
  assign n3870 = ( ~n2562 & n2569 ) | ( ~n2562 & n3869 ) | ( n2569 & n3869 ) ;
  assign n3871 = ( n2042 & ~n2048 ) | ( n2042 & n3870 ) | ( ~n2048 & n3870 ) ;
  assign n3872 = ( n1001 & ~n1018 ) | ( n1001 & n3871 ) | ( ~n1018 & n3871 ) ;
  assign n3873 = ( n2594 & ~n2601 ) | ( n2594 & n3872 ) | ( ~n2601 & n3872 ) ;
  assign n3874 = ( n3034 & ~n3120 ) | ( n3034 & n3873 ) | ( ~n3120 & n3873 ) ;
  assign n3875 = ( n3434 & ~n3515 ) | ( n3434 & n3874 ) | ( ~n3515 & n3874 ) ;
  assign n3876 = n1168 | n2094 ;
  assign n3877 = ~n1150 & n3876 ;
  assign n3878 = ( ~n1210 & n2389 ) | ( ~n1210 & n3877 ) | ( n2389 & n3877 ) ;
  assign n3879 = n1201 | n3878 ;
  assign n3880 = ( ~n1168 & n1176 ) | ( ~n1168 & n3440 ) | ( n1176 & n3440 ) ;
  assign n3881 = n1150 | n3880 ;
  assign n3882 = ~n1173 & n3881 ;
  assign n3883 = ( ~n1201 & n1211 ) | ( ~n1201 & n3882 ) | ( n1211 & n3882 ) ;
  assign n3884 = ( n3875 & n3879 ) | ( n3875 & ~n3883 ) | ( n3879 & ~n3883 ) ;
  assign n3885 = ( n1771 & ~n1777 ) | ( n1771 & n3884 ) | ( ~n1777 & n3884 ) ;
  assign n3886 = n3863 & n3885 ;
  assign n3887 = x187 & ~n430 ;
  assign n3888 = x61 | n441 ;
  assign n3889 = ~n1226 & n3888 ;
  assign n3890 = ( ~n1224 & n1788 ) | ( ~n1224 & n3889 ) | ( n1788 & n3889 ) ;
  assign n3891 = ( ~n1251 & n2125 ) | ( ~n1251 & n3890 ) | ( n2125 & n3890 ) ;
  assign n3892 = ( n1301 & ~n2624 ) | ( n1301 & n3891 ) | ( ~n2624 & n3891 ) ;
  assign n3893 = ( ~n1798 & n2139 ) | ( ~n1798 & n3892 ) | ( n2139 & n3892 ) ;
  assign n3894 = ( ~n2631 & n2638 ) | ( ~n2631 & n3893 ) | ( n2638 & n3893 ) ;
  assign n3895 = ( n2151 & ~n2157 ) | ( n2151 & n3894 ) | ( ~n2157 & n3894 ) ;
  assign n3896 = ( n1398 & ~n1415 ) | ( n1398 & n3895 ) | ( ~n1415 & n3895 ) ;
  assign n3897 = ( n2663 & ~n2670 ) | ( n2663 & n3896 ) | ( ~n2670 & n3896 ) ;
  assign n3898 = ( n3063 & ~n3147 ) | ( n3063 & n3897 ) | ( ~n3147 & n3897 ) ;
  assign n3899 = ( n3460 & ~n3541 ) | ( n3460 & n3898 ) | ( ~n3541 & n3898 ) ;
  assign n3900 = n379 & ~n415 ;
  assign n3901 = ( ~n403 & n407 ) | ( ~n403 & n3900 ) | ( n407 & n3900 ) ;
  assign n3902 = n400 | n3901 ;
  assign n3903 = ( ~n378 & n1486 ) | ( ~n378 & n3466 ) | ( n1486 & n3466 ) ;
  assign n3904 = n415 | n3903 ;
  assign n3905 = ~n406 & n3904 ;
  assign n3906 = ( ~n400 & n417 ) | ( ~n400 & n3905 ) | ( n417 & n3905 ) ;
  assign n3907 = ( n3899 & n3902 ) | ( n3899 & ~n3906 ) | ( n3902 & ~n3906 ) ;
  assign n3908 = ( n1893 & ~n1898 ) | ( n1893 & n3907 ) | ( ~n1898 & n3907 ) ;
  assign n3909 = n3887 & n3908 ;
  assign n3910 = x188 & ~n828 ;
  assign n3911 = x62 | n839 ;
  assign n3912 = ~n428 & n3911 ;
  assign n3913 = ( ~n455 & n1906 ) | ( ~n455 & n3912 ) | ( n1906 & n3912 ) ;
  assign n3914 = ( ~n1508 & n2221 ) | ( ~n1508 & n3913 ) | ( n2221 & n3913 ) ;
  assign n3915 = ( ~n493 & n1527 ) | ( ~n493 & n3914 ) | ( n1527 & n3914 ) ;
  assign n3916 = ( ~n1915 & n2235 ) | ( ~n1915 & n3915 ) | ( n2235 & n3915 ) ;
  assign n3917 = ( n546 & ~n561 ) | ( n546 & n3916 ) | ( ~n561 & n3916 ) ;
  assign n3918 = ( n2247 & ~n2253 ) | ( n2247 & n3917 ) | ( ~n2253 & n3917 ) ;
  assign n3919 = ( n1559 & ~n1569 ) | ( n1559 & n3918 ) | ( ~n1569 & n3918 ) ;
  assign n3920 = ( n2707 & ~n2714 ) | ( n2707 & n3919 ) | ( ~n2714 & n3919 ) ;
  assign n3921 = ( n3090 & ~n3174 ) | ( n3090 & n3920 ) | ( ~n3174 & n3920 ) ;
  assign n3922 = ( n3486 & ~n3566 ) | ( n3486 & n3921 ) | ( ~n3566 & n3921 ) ;
  assign n3923 = n777 & ~n813 ;
  assign n3924 = ( ~n801 & n805 ) | ( ~n801 & n3923 ) | ( n805 & n3923 ) ;
  assign n3925 = n798 | n3924 ;
  assign n3926 = ( ~n776 & n1625 ) | ( ~n776 & n3492 ) | ( n1625 & n3492 ) ;
  assign n3927 = n813 | n3926 ;
  assign n3928 = ~n804 & n3927 ;
  assign n3929 = ( ~n798 & n815 ) | ( ~n798 & n3928 ) | ( n815 & n3928 ) ;
  assign n3930 = ( n3922 & n3925 ) | ( n3922 & ~n3929 ) | ( n3925 & ~n3929 ) ;
  assign n3931 = ( n2002 & ~n2007 ) | ( n2002 & n3930 ) | ( ~n2007 & n3930 ) ;
  assign n3932 = n3910 & n3931 ;
  assign n3933 = x189 & ~n1225 ;
  assign n3934 = x63 | n1236 ;
  assign n3935 = ~n826 & n3934 ;
  assign n3936 = ( ~n853 & n2015 ) | ( ~n853 & n3935 ) | ( n2015 & n3935 ) ;
  assign n3937 = ( ~n1647 & n2317 ) | ( ~n1647 & n3936 ) | ( n2317 & n3936 ) ;
  assign n3938 = ( ~n891 & n1666 ) | ( ~n891 & n3937 ) | ( n1666 & n3937 ) ;
  assign n3939 = ( ~n2024 & n2331 ) | ( ~n2024 & n3938 ) | ( n2331 & n3938 ) ;
  assign n3940 = ( n944 & ~n959 ) | ( n944 & n3939 ) | ( ~n959 & n3939 ) ;
  assign n3941 = ( n2343 & ~n2349 ) | ( n2343 & n3940 ) | ( ~n2349 & n3940 ) ;
  assign n3942 = ( n1698 & ~n1708 ) | ( n1698 & n3941 ) | ( ~n1708 & n3941 ) ;
  assign n3943 = ( n2751 & ~n2758 ) | ( n2751 & n3942 ) | ( ~n2758 & n3942 ) ;
  assign n3944 = ( n3117 & ~n3201 ) | ( n3117 & n3943 ) | ( ~n3201 & n3943 ) ;
  assign n3945 = ( n3512 & ~n3591 ) | ( n3512 & n3944 ) | ( ~n3591 & n3944 ) ;
  assign n3946 = n1174 & ~n1210 ;
  assign n3947 = ( ~n1198 & n1202 ) | ( ~n1198 & n3946 ) | ( n1202 & n3946 ) ;
  assign n3948 = n1195 | n3947 ;
  assign n3949 = ( ~n1173 & n1763 ) | ( ~n1173 & n3518 ) | ( n1763 & n3518 ) ;
  assign n3950 = n1210 | n3949 ;
  assign n3951 = ~n1201 & n3950 ;
  assign n3952 = ( ~n1195 & n1212 ) | ( ~n1195 & n3951 ) | ( n1212 & n3951 ) ;
  assign n3953 = ( n3945 & n3948 ) | ( n3945 & ~n3952 ) | ( n3948 & ~n3952 ) ;
  assign n3954 = ( n2111 & ~n2116 ) | ( n2111 & n3953 ) | ( ~n2116 & n3953 ) ;
  assign n3955 = n3933 & n3954 ;
  assign n3956 = x190 & ~n427 ;
  assign n3957 = x64 | n446 ;
  assign n3958 = ~n1223 & n3957 ;
  assign n3959 = ( ~n1250 & n2124 ) | ( ~n1250 & n3958 ) | ( n2124 & n3958 ) ;
  assign n3960 = ( ~n1785 & n2413 ) | ( ~n1785 & n3959 ) | ( n2413 & n3959 ) ;
  assign n3961 = ( ~n1288 & n1804 ) | ( ~n1288 & n3960 ) | ( n1804 & n3960 ) ;
  assign n3962 = ( ~n2133 & n2427 ) | ( ~n2133 & n3961 ) | ( n2427 & n3961 ) ;
  assign n3963 = ( n1341 & ~n1356 ) | ( n1341 & n3962 ) | ( ~n1356 & n3962 ) ;
  assign n3964 = ( n2439 & ~n2445 ) | ( n2439 & n3963 ) | ( ~n2445 & n3963 ) ;
  assign n3965 = ( n1836 & ~n1846 ) | ( n1836 & n3964 ) | ( ~n1846 & n3964 ) ;
  assign n3966 = ( n2795 & ~n2802 ) | ( n2795 & n3965 ) | ( ~n2802 & n3965 ) ;
  assign n3967 = ( n3144 & ~n3228 ) | ( n3144 & n3966 ) | ( ~n3228 & n3966 ) ;
  assign n3968 = ( n3538 & ~n3616 ) | ( n3538 & n3967 ) | ( ~n3616 & n3967 ) ;
  assign n3969 = ~n403 & n1485 ;
  assign n3970 = ( ~n397 & n1491 ) | ( ~n397 & n3969 ) | ( n1491 & n3969 ) ;
  assign n3971 = n394 | n3970 ;
  assign n3972 = ( n384 & ~n406 ) | ( n384 & n416 ) | ( ~n406 & n416 ) ;
  assign n3973 = n403 | n3972 ;
  assign n3974 = ~n400 & n3973 ;
  assign n3975 = ( ~n394 & n1497 ) | ( ~n394 & n3974 ) | ( n1497 & n3974 ) ;
  assign n3976 = ( n3968 & n3971 ) | ( n3968 & ~n3975 ) | ( n3971 & ~n3975 ) ;
  assign n3977 = ( n2207 & ~n2212 ) | ( n2207 & n3976 ) | ( ~n2212 & n3976 ) ;
  assign n3978 = n3956 & n3977 ;
  assign n3979 = x191 & ~n825 ;
  assign n3980 = x65 | n844 ;
  assign n3981 = ~n454 & n3980 ;
  assign n3982 = ( ~n426 & n2220 ) | ( ~n426 & n3981 ) | ( n2220 & n3981 ) ;
  assign n3983 = ( ~n488 & n506 ) | ( ~n488 & n3982 ) | ( n506 & n3982 ) ;
  assign n3984 = ( ~n1520 & n1920 ) | ( ~n1520 & n3983 ) | ( n1920 & n3983 ) ;
  assign n3985 = ( ~n2229 & n2498 ) | ( ~n2229 & n3984 ) | ( n2498 & n3984 ) ;
  assign n3986 = ( n1539 & ~n1547 ) | ( n1539 & n3985 ) | ( ~n1547 & n3985 ) ;
  assign n3987 = ( n2509 & ~n2515 ) | ( n2509 & n3986 ) | ( ~n2515 & n3986 ) ;
  assign n3988 = ( n1949 & ~n1956 ) | ( n1949 & n3987 ) | ( ~n1956 & n3987 ) ;
  assign n3989 = ( n2828 & ~n2832 ) | ( n2828 & n3988 ) | ( ~n2832 & n3988 ) ;
  assign n3990 = ( n3171 & ~n3254 ) | ( n3171 & n3989 ) | ( ~n3254 & n3989 ) ;
  assign n3991 = ( n3563 & ~n3641 ) | ( n3563 & n3990 ) | ( ~n3641 & n3990 ) ;
  assign n3992 = ~n801 & n1624 ;
  assign n3993 = ( ~n795 & n1630 ) | ( ~n795 & n3992 ) | ( n1630 & n3992 ) ;
  assign n3994 = n792 | n3993 ;
  assign n3995 = ( n782 & ~n804 ) | ( n782 & n814 ) | ( ~n804 & n814 ) ;
  assign n3996 = n801 | n3995 ;
  assign n3997 = ~n798 & n3996 ;
  assign n3998 = ( ~n792 & n1636 ) | ( ~n792 & n3997 ) | ( n1636 & n3997 ) ;
  assign n3999 = ( n3991 & n3994 ) | ( n3991 & ~n3998 ) | ( n3994 & ~n3998 ) ;
  assign n4000 = ( n2303 & ~n2308 ) | ( n2303 & n3999 ) | ( ~n2308 & n3999 ) ;
  assign n4001 = n3979 & n4000 ;
  assign n4002 = x192 & ~n1222 ;
  assign n4003 = x66 | n1241 ;
  assign n4004 = ~n852 & n4003 ;
  assign n4005 = ( ~n824 & n2316 ) | ( ~n824 & n4004 ) | ( n2316 & n4004 ) ;
  assign n4006 = ( ~n886 & n904 ) | ( ~n886 & n4005 ) | ( n904 & n4005 ) ;
  assign n4007 = ( ~n1659 & n2029 ) | ( ~n1659 & n4006 ) | ( n2029 & n4006 ) ;
  assign n4008 = ( ~n2325 & n2567 ) | ( ~n2325 & n4007 ) | ( n2567 & n4007 ) ;
  assign n4009 = ( n1678 & ~n1686 ) | ( n1678 & n4008 ) | ( ~n1686 & n4008 ) ;
  assign n4010 = ( n2578 & ~n2584 ) | ( n2578 & n4009 ) | ( ~n2584 & n4009 ) ;
  assign n4011 = ( n2058 & ~n2065 ) | ( n2058 & n4010 ) | ( ~n2065 & n4010 ) ;
  assign n4012 = ( n2858 & ~n2862 ) | ( n2858 & n4011 ) | ( ~n2862 & n4011 ) ;
  assign n4013 = ( n3198 & ~n3280 ) | ( n3198 & n4012 ) | ( ~n3280 & n4012 ) ;
  assign n4014 = ( n3588 & ~n3666 ) | ( n3588 & n4013 ) | ( ~n3666 & n4013 ) ;
  assign n4015 = ~n1198 & n1762 ;
  assign n4016 = ( ~n1192 & n1768 ) | ( ~n1192 & n4015 ) | ( n1768 & n4015 ) ;
  assign n4017 = n1189 | n4016 ;
  assign n4018 = ( n1179 & ~n1201 ) | ( n1179 & n1211 ) | ( ~n1201 & n1211 ) ;
  assign n4019 = n1198 | n4018 ;
  assign n4020 = ~n1195 & n4019 ;
  assign n4021 = ( ~n1189 & n1774 ) | ( ~n1189 & n4020 ) | ( n1774 & n4020 ) ;
  assign n4022 = ( n4014 & n4017 ) | ( n4014 & ~n4021 ) | ( n4017 & ~n4021 ) ;
  assign n4023 = ( n2399 & ~n2404 ) | ( n2399 & n4022 ) | ( ~n2404 & n4022 ) ;
  assign n4024 = n4002 & n4023 ;
  assign n4025 = x193 & ~n453 ;
  assign n4026 = x67 | n450 ;
  assign n4027 = ~n1249 & n4026 ;
  assign n4028 = ( ~n1221 & n2412 ) | ( ~n1221 & n4027 ) | ( n2412 & n4027 ) ;
  assign n4029 = ( ~n1283 & n1301 ) | ( ~n1283 & n4028 ) | ( n1301 & n4028 ) ;
  assign n4030 = ( ~n1797 & n2138 ) | ( ~n1797 & n4029 ) | ( n2138 & n4029 ) ;
  assign n4031 = ( ~n2421 & n2636 ) | ( ~n2421 & n4030 ) | ( n2636 & n4030 ) ;
  assign n4032 = ( n1816 & ~n1824 ) | ( n1816 & n4031 ) | ( ~n1824 & n4031 ) ;
  assign n4033 = ( n2647 & ~n2653 ) | ( n2647 & n4032 ) | ( ~n2653 & n4032 ) ;
  assign n4034 = ( n2167 & ~n2174 ) | ( n2167 & n4033 ) | ( ~n2174 & n4033 ) ;
  assign n4035 = ( n2888 & ~n2892 ) | ( n2888 & n4034 ) | ( ~n2892 & n4034 ) ;
  assign n4036 = ( n3225 & ~n3306 ) | ( n3225 & n4035 ) | ( ~n3306 & n4035 ) ;
  assign n4037 = ( n3613 & ~n3690 ) | ( n3613 & n4036 ) | ( ~n3690 & n4036 ) ;
  assign n4038 = ~n397 & n1885 ;
  assign n4039 = ( ~n391 & n1890 ) | ( ~n391 & n4038 ) | ( n1890 & n4038 ) ;
  assign n4040 = n388 | n4039 ;
  assign n4041 = ( ~n400 & n417 ) | ( ~n400 & n1489 ) | ( n417 & n1489 ) ;
  assign n4042 = n397 | n4041 ;
  assign n4043 = ~n394 & n4042 ;
  assign n4044 = ( ~n388 & n421 ) | ( ~n388 & n4043 ) | ( n421 & n4043 ) ;
  assign n4045 = ( n4037 & n4040 ) | ( n4037 & ~n4044 ) | ( n4040 & ~n4044 ) ;
  assign n4046 = ( ~n449 & n462 ) | ( ~n449 & n4045 ) | ( n462 & n4045 ) ;
  assign n4047 = n4025 & n4046 ;
  assign n4048 = x194 & ~n851 ;
  assign n4049 = x68 | n848 ;
  assign n4050 = ~n425 & n4049 ;
  assign n4051 = ( ~n484 & n505 ) | ( ~n484 & n4050 ) | ( n505 & n4050 ) ;
  assign n4052 = ( ~n492 & n1527 ) | ( ~n492 & n4051 ) | ( n1527 & n4051 ) ;
  assign n4053 = ( ~n1914 & n2234 ) | ( ~n1914 & n4052 ) | ( n2234 & n4052 ) ;
  assign n4054 = ( n541 & ~n2493 ) | ( n541 & n4053 ) | ( ~n2493 & n4053 ) ;
  assign n4055 = ( n1932 & ~n1938 ) | ( n1932 & n4054 ) | ( ~n1938 & n4054 ) ;
  assign n4056 = ( ~n618 & n2697 ) | ( ~n618 & n4055 ) | ( n2697 & n4055 ) ;
  assign n4057 = ( n2263 & ~n2270 ) | ( n2263 & n4056 ) | ( ~n2270 & n4056 ) ;
  assign n4058 = ( n2917 & ~n2921 ) | ( n2917 & n4057 ) | ( ~n2921 & n4057 ) ;
  assign n4059 = ( n3251 & ~n3332 ) | ( n3251 & n4058 ) | ( ~n3332 & n4058 ) ;
  assign n4060 = ( n3638 & ~n3714 ) | ( n3638 & n4059 ) | ( ~n3714 & n4059 ) ;
  assign n4061 = ~n795 & n1994 ;
  assign n4062 = ( ~n789 & n1999 ) | ( ~n789 & n4061 ) | ( n1999 & n4061 ) ;
  assign n4063 = n786 | n4062 ;
  assign n4064 = ( ~n798 & n815 ) | ( ~n798 & n1628 ) | ( n815 & n1628 ) ;
  assign n4065 = n795 | n4064 ;
  assign n4066 = ~n792 & n4065 ;
  assign n4067 = ( ~n786 & n819 ) | ( ~n786 & n4066 ) | ( n819 & n4066 ) ;
  assign n4068 = ( n4060 & n4063 ) | ( n4060 & ~n4067 ) | ( n4063 & ~n4067 ) ;
  assign n4069 = ( ~n847 & n860 ) | ( ~n847 & n4068 ) | ( n860 & n4068 ) ;
  assign n4070 = n4048 & n4069 ;
  assign n4071 = x195 & ~n1248 ;
  assign n4072 = x69 | n1245 ;
  assign n4073 = ~n823 & n4072 ;
  assign n4074 = ( ~n882 & n903 ) | ( ~n882 & n4073 ) | ( n903 & n4073 ) ;
  assign n4075 = ( ~n890 & n1666 ) | ( ~n890 & n4074 ) | ( n1666 & n4074 ) ;
  assign n4076 = ( ~n2023 & n2330 ) | ( ~n2023 & n4075 ) | ( n2330 & n4075 ) ;
  assign n4077 = ( n939 & ~n2562 ) | ( n939 & n4076 ) | ( ~n2562 & n4076 ) ;
  assign n4078 = ( n2041 & ~n2047 ) | ( n2041 & n4077 ) | ( ~n2047 & n4077 ) ;
  assign n4079 = ( ~n1016 & n2741 ) | ( ~n1016 & n4078 ) | ( n2741 & n4078 ) ;
  assign n4080 = ( n2359 & ~n2366 ) | ( n2359 & n4079 ) | ( ~n2366 & n4079 ) ;
  assign n4081 = ( n2946 & ~n2950 ) | ( n2946 & n4080 ) | ( ~n2950 & n4080 ) ;
  assign n4082 = ( n3277 & ~n3358 ) | ( n3277 & n4081 ) | ( ~n3358 & n4081 ) ;
  assign n4083 = ( n3663 & ~n3738 ) | ( n3663 & n4082 ) | ( ~n3738 & n4082 ) ;
  assign n4084 = ~n1192 & n2103 ;
  assign n4085 = ( ~n1186 & n2108 ) | ( ~n1186 & n4084 ) | ( n2108 & n4084 ) ;
  assign n4086 = n1183 | n4085 ;
  assign n4087 = ( ~n1195 & n1212 ) | ( ~n1195 & n1766 ) | ( n1212 & n1766 ) ;
  assign n4088 = n1192 | n4087 ;
  assign n4089 = ~n1189 & n4088 ;
  assign n4090 = ( ~n1183 & n1216 ) | ( ~n1183 & n4089 ) | ( n1216 & n4089 ) ;
  assign n4091 = ( n4083 & n4086 ) | ( n4083 & ~n4090 ) | ( n4086 & ~n4090 ) ;
  assign n4092 = ( ~n1244 & n1257 ) | ( ~n1244 & n4091 ) | ( n1257 & n4091 ) ;
  assign n4093 = n4071 & n4092 ;
  assign n4094 = x196 & ~n424 ;
  assign n4095 = x70 | n502 ;
  assign n4096 = ~n1220 & n4095 ;
  assign n4097 = ( ~n1279 & n1300 ) | ( ~n1279 & n4096 ) | ( n1300 & n4096 ) ;
  assign n4098 = ( ~n1287 & n1804 ) | ( ~n1287 & n4097 ) | ( n1804 & n4097 ) ;
  assign n4099 = ( ~n2132 & n2426 ) | ( ~n2132 & n4098 ) | ( n2426 & n4098 ) ;
  assign n4100 = ( n1336 & ~n2631 ) | ( n1336 & n4099 ) | ( ~n2631 & n4099 ) ;
  assign n4101 = ( n2150 & ~n2156 ) | ( n2150 & n4100 ) | ( ~n2156 & n4100 ) ;
  assign n4102 = ( ~n1413 & n2785 ) | ( ~n1413 & n4101 ) | ( n2785 & n4101 ) ;
  assign n4103 = ( n2455 & ~n2462 ) | ( n2455 & n4102 ) | ( ~n2462 & n4102 ) ;
  assign n4104 = ( n2975 & ~n2979 ) | ( n2975 & n4103 ) | ( ~n2979 & n4103 ) ;
  assign n4105 = ( n3303 & ~n3384 ) | ( n3303 & n4104 ) | ( ~n3384 & n4104 ) ;
  assign n4106 = ( n3687 & ~n3762 ) | ( n3687 & n4105 ) | ( ~n3762 & n4105 ) ;
  assign n4107 = ~n391 & n2202 ;
  assign n4108 = ( ~n435 & n2204 ) | ( ~n435 & n4107 ) | ( n2204 & n4107 ) ;
  assign n4109 = n438 | n4108 ;
  assign n4110 = ( ~n394 & n1497 ) | ( ~n394 & n1888 ) | ( n1497 & n1888 ) ;
  assign n4111 = n391 | n4110 ;
  assign n4112 = ~n388 & n4111 ;
  assign n4113 = ( ~n438 & n439 ) | ( ~n438 & n4112 ) | ( n439 & n4112 ) ;
  assign n4114 = ( n4106 & n4109 ) | ( n4106 & ~n4113 ) | ( n4109 & ~n4113 ) ;
  assign n4115 = ( ~n1507 & n1514 ) | ( ~n1507 & n4114 ) | ( n1514 & n4114 ) ;
  assign n4116 = n4094 & n4115 ;
  assign n4117 = x197 & ~n822 ;
  assign n4118 = x71 | n900 ;
  assign n4119 = ~n483 & n4118 ;
  assign n4120 = ( ~n491 & n1526 ) | ( ~n491 & n4119 ) | ( n1526 & n4119 ) ;
  assign n4121 = ( ~n1519 & n1920 ) | ( ~n1519 & n4120 ) | ( n1920 & n4120 ) ;
  assign n4122 = ( ~n2228 & n2497 ) | ( ~n2228 & n4121 ) | ( n2497 & n4121 ) ;
  assign n4123 = ( ~n561 & n1537 ) | ( ~n561 & n4122 ) | ( n1537 & n4122 ) ;
  assign n4124 = ( n2246 & ~n2252 ) | ( n2246 & n4123 ) | ( ~n2252 & n4123 ) ;
  assign n4125 = ( n603 & ~n1567 ) | ( n603 & n4124 ) | ( ~n1567 & n4124 ) ;
  assign n4126 = ( n2524 & ~n2531 ) | ( n2524 & n4125 ) | ( ~n2531 & n4125 ) ;
  assign n4127 = ( n3004 & ~n3008 ) | ( n3004 & n4126 ) | ( ~n3008 & n4126 ) ;
  assign n4128 = ( n3329 & ~n3410 ) | ( n3329 & n4127 ) | ( ~n3410 & n4127 ) ;
  assign n4129 = ( n3711 & ~n3786 ) | ( n3711 & n4128 ) | ( ~n3786 & n4128 ) ;
  assign n4130 = ~n789 & n2298 ;
  assign n4131 = ( ~n833 & n2300 ) | ( ~n833 & n4130 ) | ( n2300 & n4130 ) ;
  assign n4132 = n836 | n4131 ;
  assign n4133 = ( ~n792 & n1636 ) | ( ~n792 & n1997 ) | ( n1636 & n1997 ) ;
  assign n4134 = n789 | n4133 ;
  assign n4135 = ~n786 & n4134 ;
  assign n4136 = ( ~n836 & n837 ) | ( ~n836 & n4135 ) | ( n837 & n4135 ) ;
  assign n4137 = ( n4129 & n4132 ) | ( n4129 & ~n4136 ) | ( n4132 & ~n4136 ) ;
  assign n4138 = ( ~n1646 & n1653 ) | ( ~n1646 & n4137 ) | ( n1653 & n4137 ) ;
  assign n4139 = n4117 & n4138 ;
  assign n4140 = x198 & ~n1219 ;
  assign n4141 = x72 | n1297 ;
  assign n4142 = ~n881 & n4141 ;
  assign n4143 = ( ~n889 & n1665 ) | ( ~n889 & n4142 ) | ( n1665 & n4142 ) ;
  assign n4144 = ( ~n1658 & n2029 ) | ( ~n1658 & n4143 ) | ( n2029 & n4143 ) ;
  assign n4145 = ( ~n2324 & n2566 ) | ( ~n2324 & n4144 ) | ( n2566 & n4144 ) ;
  assign n4146 = ( ~n959 & n1676 ) | ( ~n959 & n4145 ) | ( n1676 & n4145 ) ;
  assign n4147 = ( n2342 & ~n2348 ) | ( n2342 & n4146 ) | ( ~n2348 & n4146 ) ;
  assign n4148 = ( n1001 & ~n1706 ) | ( n1001 & n4147 ) | ( ~n1706 & n4147 ) ;
  assign n4149 = ( n2593 & ~n2600 ) | ( n2593 & n4148 ) | ( ~n2600 & n4148 ) ;
  assign n4150 = ( n3033 & ~n3037 ) | ( n3033 & n4149 ) | ( ~n3037 & n4149 ) ;
  assign n4151 = ( n3355 & ~n3436 ) | ( n3355 & n4150 ) | ( ~n3436 & n4150 ) ;
  assign n4152 = ( n3735 & ~n3810 ) | ( n3735 & n4151 ) | ( ~n3810 & n4151 ) ;
  assign n4153 = ~n1186 & n2394 ;
  assign n4154 = ( ~n1230 & n2396 ) | ( ~n1230 & n4153 ) | ( n2396 & n4153 ) ;
  assign n4155 = n1233 | n4154 ;
  assign n4156 = ( ~n1189 & n1774 ) | ( ~n1189 & n2106 ) | ( n1774 & n2106 ) ;
  assign n4157 = n1186 | n4156 ;
  assign n4158 = ~n1183 & n4157 ;
  assign n4159 = ( ~n1233 & n1234 ) | ( ~n1233 & n4158 ) | ( n1234 & n4158 ) ;
  assign n4160 = ( n4152 & n4155 ) | ( n4152 & ~n4159 ) | ( n4155 & ~n4159 ) ;
  assign n4161 = ( ~n1784 & n1791 ) | ( ~n1784 & n4160 ) | ( n1791 & n4160 ) ;
  assign n4162 = n4140 & n4161 ;
  assign n4163 = x199 & ~n482 ;
  assign n4164 = x73 | n485 ;
  assign n4165 = ~n1278 & n4164 ;
  assign n4166 = ( ~n1286 & n1803 ) | ( ~n1286 & n4165 ) | ( n1803 & n4165 ) ;
  assign n4167 = ( ~n1796 & n2138 ) | ( ~n1796 & n4166 ) | ( n2138 & n4166 ) ;
  assign n4168 = ( ~n2420 & n2635 ) | ( ~n2420 & n4167 ) | ( n2635 & n4167 ) ;
  assign n4169 = ( ~n1356 & n1814 ) | ( ~n1356 & n4168 ) | ( n1814 & n4168 ) ;
  assign n4170 = ( n2438 & ~n2444 ) | ( n2438 & n4169 ) | ( ~n2444 & n4169 ) ;
  assign n4171 = ( n1398 & ~n1844 ) | ( n1398 & n4170 ) | ( ~n1844 & n4170 ) ;
  assign n4172 = ( n2662 & ~n2669 ) | ( n2662 & n4171 ) | ( ~n2669 & n4171 ) ;
  assign n4173 = ( n3062 & ~n3066 ) | ( n3062 & n4172 ) | ( ~n3066 & n4172 ) ;
  assign n4174 = ( n3381 & ~n3462 ) | ( n3381 & n4173 ) | ( ~n3462 & n4173 ) ;
  assign n4175 = ( n3759 & ~n3834 ) | ( n3759 & n4174 ) | ( ~n3834 & n4174 ) ;
  assign n4176 = n412 & ~n435 ;
  assign n4177 = ( ~n432 & n459 ) | ( ~n432 & n4176 ) | ( n459 & n4176 ) ;
  assign n4178 = n443 | n4177 ;
  assign n4179 = n422 | n435 ;
  assign n4180 = ~n438 & n4179 ;
  assign n4181 = ( ~n443 & n1503 ) | ( ~n443 & n4180 ) | ( n1503 & n4180 ) ;
  assign n4182 = ( n4175 & n4178 ) | ( n4175 & ~n4181 ) | ( n4178 & ~n4181 ) ;
  assign n4183 = ( ~n1903 & n1909 ) | ( ~n1903 & n4182 ) | ( n1909 & n4182 ) ;
  assign n4184 = n4163 & n4183 ;
  assign n4185 = x200 & ~n880 ;
  assign n4186 = x74 | n883 ;
  assign n4187 = ~n490 & n4186 ;
  assign n4188 = ( ~n478 & n1919 ) | ( ~n478 & n4187 ) | ( n1919 & n4187 ) ;
  assign n4189 = ( ~n499 & n2234 ) | ( ~n499 & n4188 ) | ( n2234 & n4188 ) ;
  assign n4190 = ( n540 & ~n2492 ) | ( n540 & n4189 ) | ( ~n2492 & n4189 ) ;
  assign n4191 = ( ~n1547 & n1930 ) | ( ~n1547 & n4190 ) | ( n1930 & n4190 ) ;
  assign n4192 = ( n2508 & ~n2514 ) | ( n2508 & n4191 ) | ( ~n2514 & n4191 ) ;
  assign n4193 = ( n1559 & ~n1955 ) | ( n1559 & n4192 ) | ( ~n1955 & n4192 ) ;
  assign n4194 = ( n2706 & ~n2713 ) | ( n2706 & n4193 ) | ( ~n2713 & n4193 ) ;
  assign n4195 = ( n3089 & ~n3093 ) | ( n3089 & n4194 ) | ( ~n3093 & n4194 ) ;
  assign n4196 = ( n3407 & ~n3488 ) | ( n3407 & n4195 ) | ( ~n3488 & n4195 ) ;
  assign n4197 = ( n3783 & ~n3858 ) | ( n3783 & n4196 ) | ( ~n3858 & n4196 ) ;
  assign n4198 = n810 & ~n833 ;
  assign n4199 = ( ~n830 & n857 ) | ( ~n830 & n4198 ) | ( n857 & n4198 ) ;
  assign n4200 = n841 | n4199 ;
  assign n4201 = n820 | n833 ;
  assign n4202 = ~n836 & n4201 ;
  assign n4203 = ( ~n841 & n1642 ) | ( ~n841 & n4202 ) | ( n1642 & n4202 ) ;
  assign n4204 = ( n4197 & n4200 ) | ( n4197 & ~n4203 ) | ( n4200 & ~n4203 ) ;
  assign n4205 = ( ~n2012 & n2018 ) | ( ~n2012 & n4204 ) | ( n2018 & n4204 ) ;
  assign n4206 = n4185 & n4205 ;
  assign n4207 = x201 & ~n1277 ;
  assign n4208 = x75 | n1280 ;
  assign n4209 = ~n888 & n4208 ;
  assign n4210 = ( ~n876 & n2028 ) | ( ~n876 & n4209 ) | ( n2028 & n4209 ) ;
  assign n4211 = ( ~n897 & n2330 ) | ( ~n897 & n4210 ) | ( n2330 & n4210 ) ;
  assign n4212 = ( n938 & ~n2561 ) | ( n938 & n4211 ) | ( ~n2561 & n4211 ) ;
  assign n4213 = ( ~n1686 & n2039 ) | ( ~n1686 & n4212 ) | ( n2039 & n4212 ) ;
  assign n4214 = ( n2577 & ~n2583 ) | ( n2577 & n4213 ) | ( ~n2583 & n4213 ) ;
  assign n4215 = ( n1698 & ~n2064 ) | ( n1698 & n4214 ) | ( ~n2064 & n4214 ) ;
  assign n4216 = ( n2750 & ~n2757 ) | ( n2750 & n4215 ) | ( ~n2757 & n4215 ) ;
  assign n4217 = ( n3116 & ~n3120 ) | ( n3116 & n4216 ) | ( ~n3120 & n4216 ) ;
  assign n4218 = ( n3433 & ~n3514 ) | ( n3433 & n4217 ) | ( ~n3514 & n4217 ) ;
  assign n4219 = ( n3807 & ~n3882 ) | ( n3807 & n4218 ) | ( ~n3882 & n4218 ) ;
  assign n4220 = n1207 & ~n1230 ;
  assign n4221 = ( ~n1227 & n1254 ) | ( ~n1227 & n4220 ) | ( n1254 & n4220 ) ;
  assign n4222 = n1238 | n4221 ;
  assign n4223 = n1217 | n1230 ;
  assign n4224 = ~n1233 & n4223 ;
  assign n4225 = ( ~n1238 & n1780 ) | ( ~n1238 & n4224 ) | ( n1780 & n4224 ) ;
  assign n4226 = ( n4219 & n4222 ) | ( n4219 & ~n4225 ) | ( n4222 & ~n4225 ) ;
  assign n4227 = ( ~n2121 & n2127 ) | ( ~n2121 & n4226 ) | ( n2127 & n4226 ) ;
  assign n4228 = n4207 & n4227 ;
  assign n4229 = x202 & ~n489 ;
  assign n4230 = x76 | n479 ;
  assign n4231 = ~n1285 & n4230 ;
  assign n4232 = ( ~n1273 & n2137 ) | ( ~n1273 & n4231 ) | ( n2137 & n4231 ) ;
  assign n4233 = ( ~n1294 & n2426 ) | ( ~n1294 & n4232 ) | ( n2426 & n4232 ) ;
  assign n4234 = ( n1335 & ~n2630 ) | ( n1335 & n4233 ) | ( ~n2630 & n4233 ) ;
  assign n4235 = ( ~n1824 & n2148 ) | ( ~n1824 & n4234 ) | ( n2148 & n4234 ) ;
  assign n4236 = ( n2646 & ~n2652 ) | ( n2646 & n4235 ) | ( ~n2652 & n4235 ) ;
  assign n4237 = ( n1836 & ~n2173 ) | ( n1836 & n4236 ) | ( ~n2173 & n4236 ) ;
  assign n4238 = ( n2794 & ~n2801 ) | ( n2794 & n4237 ) | ( ~n2801 & n4237 ) ;
  assign n4239 = ( n3143 & ~n3147 ) | ( n3143 & n4238 ) | ( ~n3147 & n4238 ) ;
  assign n4240 = ( n3459 & ~n3540 ) | ( n3459 & n4239 ) | ( ~n3540 & n4239 ) ;
  assign n4241 = ( n3831 & ~n3905 ) | ( n3831 & n4240 ) | ( ~n3905 & n4240 ) ;
  assign n4242 = ~n432 & n1496 ;
  assign n4243 = ( ~n429 & n1511 ) | ( ~n429 & n4242 ) | ( n1511 & n4242 ) ;
  assign n4244 = n448 | n4243 ;
  assign n4245 = n432 | n1501 ;
  assign n4246 = ~n443 & n4245 ;
  assign n4247 = ( ~n448 & n1504 ) | ( ~n448 & n4246 ) | ( n1504 & n4246 ) ;
  assign n4248 = ( n4241 & n4244 ) | ( n4241 & ~n4247 ) | ( n4244 & ~n4247 ) ;
  assign n4249 = ( ~n2217 & n2223 ) | ( ~n2217 & n4248 ) | ( n2223 & n4248 ) ;
  assign n4250 = n4229 & n4249 ;
  assign n4251 = x203 & ~n887 ;
  assign n4252 = x77 | n877 ;
  assign n4253 = ~n477 & n4252 ;
  assign n4254 = ( ~n498 & n2233 ) | ( ~n498 & n4253 ) | ( n2233 & n4253 ) ;
  assign n4255 = ( ~n1523 & n2497 ) | ( ~n1523 & n4254 ) | ( n2497 & n4254 ) ;
  assign n4256 = ( ~n560 & n1536 ) | ( ~n560 & n4255 ) | ( n1536 & n4255 ) ;
  assign n4257 = ( ~n1938 & n2244 ) | ( ~n1938 & n4256 ) | ( n2244 & n4256 ) ;
  assign n4258 = ( ~n617 & n2696 ) | ( ~n617 & n4257 ) | ( n2696 & n4257 ) ;
  assign n4259 = ( n1949 & ~n2269 ) | ( n1949 & n4258 ) | ( ~n2269 & n4258 ) ;
  assign n4260 = ( n2827 & ~n2831 ) | ( n2827 & n4259 ) | ( ~n2831 & n4259 ) ;
  assign n4261 = ( n3170 & ~n3174 ) | ( n3170 & n4260 ) | ( ~n3174 & n4260 ) ;
  assign n4262 = ( n3485 & ~n3565 ) | ( n3485 & n4261 ) | ( ~n3565 & n4261 ) ;
  assign n4263 = ( n3855 & ~n3928 ) | ( n3855 & n4262 ) | ( ~n3928 & n4262 ) ;
  assign n4264 = ~n830 & n1635 ;
  assign n4265 = ( ~n827 & n1650 ) | ( ~n827 & n4264 ) | ( n1650 & n4264 ) ;
  assign n4266 = n846 | n4265 ;
  assign n4267 = n830 | n1640 ;
  assign n4268 = ~n841 & n4267 ;
  assign n4269 = ( ~n846 & n1643 ) | ( ~n846 & n4268 ) | ( n1643 & n4268 ) ;
  assign n4270 = ( n4263 & n4266 ) | ( n4263 & ~n4269 ) | ( n4266 & ~n4269 ) ;
  assign n4271 = ( ~n2313 & n2319 ) | ( ~n2313 & n4270 ) | ( n2319 & n4270 ) ;
  assign n4272 = n4251 & n4271 ;
  assign n4273 = x204 & ~n1284 ;
  assign n4274 = x78 | n1274 ;
  assign n4275 = ~n875 & n4274 ;
  assign n4276 = ( ~n896 & n2329 ) | ( ~n896 & n4275 ) | ( n2329 & n4275 ) ;
  assign n4277 = ( ~n1662 & n2566 ) | ( ~n1662 & n4276 ) | ( n2566 & n4276 ) ;
  assign n4278 = ( ~n958 & n1675 ) | ( ~n958 & n4277 ) | ( n1675 & n4277 ) ;
  assign n4279 = ( ~n2047 & n2340 ) | ( ~n2047 & n4278 ) | ( n2340 & n4278 ) ;
  assign n4280 = ( ~n1015 & n2740 ) | ( ~n1015 & n4279 ) | ( n2740 & n4279 ) ;
  assign n4281 = ( n2058 & ~n2365 ) | ( n2058 & n4280 ) | ( ~n2365 & n4280 ) ;
  assign n4282 = ( n2857 & ~n2861 ) | ( n2857 & n4281 ) | ( ~n2861 & n4281 ) ;
  assign n4283 = ( n3197 & ~n3201 ) | ( n3197 & n4282 ) | ( ~n3201 & n4282 ) ;
  assign n4284 = ( n3511 & ~n3590 ) | ( n3511 & n4283 ) | ( ~n3590 & n4283 ) ;
  assign n4285 = ( n3879 & ~n3951 ) | ( n3879 & n4284 ) | ( ~n3951 & n4284 ) ;
  assign n4286 = ~n1227 & n1773 ;
  assign n4287 = ( ~n1224 & n1788 ) | ( ~n1224 & n4286 ) | ( n1788 & n4286 ) ;
  assign n4288 = n1243 | n4287 ;
  assign n4289 = n1227 | n1778 ;
  assign n4290 = ~n1238 & n4289 ;
  assign n4291 = ( ~n1243 & n1781 ) | ( ~n1243 & n4290 ) | ( n1781 & n4290 ) ;
  assign n4292 = ( n4285 & n4288 ) | ( n4285 & ~n4291 ) | ( n4288 & ~n4291 ) ;
  assign n4293 = ( ~n2409 & n2415 ) | ( ~n2409 & n4292 ) | ( n2415 & n4292 ) ;
  assign n4294 = n4273 & n4293 ;
  assign n4295 = x205 & ~n476 ;
  assign n4296 = x79 | n473 ;
  assign n4297 = ~n1272 & n4296 ;
  assign n4298 = ( ~n1293 & n2425 ) | ( ~n1293 & n4297 ) | ( n2425 & n4297 ) ;
  assign n4299 = ( ~n1800 & n2635 ) | ( ~n1800 & n4298 ) | ( n2635 & n4298 ) ;
  assign n4300 = ( ~n1355 & n1813 ) | ( ~n1355 & n4299 ) | ( n1813 & n4299 ) ;
  assign n4301 = ( ~n2156 & n2436 ) | ( ~n2156 & n4300 ) | ( n2436 & n4300 ) ;
  assign n4302 = ( ~n1412 & n2784 ) | ( ~n1412 & n4301 ) | ( n2784 & n4301 ) ;
  assign n4303 = ( n2167 & ~n2461 ) | ( n2167 & n4302 ) | ( ~n2461 & n4302 ) ;
  assign n4304 = ( n2887 & ~n2891 ) | ( n2887 & n4303 ) | ( ~n2891 & n4303 ) ;
  assign n4305 = ( n3224 & ~n3228 ) | ( n3224 & n4304 ) | ( ~n3228 & n4304 ) ;
  assign n4306 = ( n3537 & ~n3615 ) | ( n3537 & n4305 ) | ( ~n3615 & n4305 ) ;
  assign n4307 = ( n3902 & ~n3974 ) | ( n3902 & n4306 ) | ( ~n3974 & n4306 ) ;
  assign n4308 = ~n429 & n1895 ;
  assign n4309 = ( ~n455 & n1906 ) | ( ~n455 & n4308 ) | ( n1906 & n4308 ) ;
  assign n4310 = n452 | n4309 ;
  assign n4311 = n429 | n1899 ;
  assign n4312 = ~n448 & n4311 ;
  assign n4313 = ( ~n452 & n456 ) | ( ~n452 & n4312 ) | ( n456 & n4312 ) ;
  assign n4314 = ( n4307 & n4310 ) | ( n4307 & ~n4313 ) | ( n4310 & ~n4313 ) ;
  assign n4315 = ( n508 & ~n2488 ) | ( n508 & n4314 ) | ( ~n2488 & n4314 ) ;
  assign n4316 = n4295 & n4315 ;
  assign n4317 = x206 & ~n874 ;
  assign n4318 = x80 | n871 ;
  assign n4319 = ~n497 & n4318 ;
  assign n4320 = ( ~n469 & n512 ) | ( ~n469 & n4319 ) | ( n512 & n4319 ) ;
  assign n4321 = ( n540 & ~n558 ) | ( n540 & n4320 ) | ( ~n558 & n4320 ) ;
  assign n4322 = ( ~n1546 & n1929 ) | ( ~n1546 & n4321 ) | ( n1929 & n4321 ) ;
  assign n4323 = ( ~n2252 & n2506 ) | ( ~n2252 & n4322 ) | ( n2506 & n4322 ) ;
  assign n4324 = ( n602 & ~n1566 ) | ( n602 & n4323 ) | ( ~n1566 & n4323 ) ;
  assign n4325 = ( n2263 & ~n2530 ) | ( n2263 & n4324 ) | ( ~n2530 & n4324 ) ;
  assign n4326 = ( n2916 & ~n2920 ) | ( n2916 & n4325 ) | ( ~n2920 & n4325 ) ;
  assign n4327 = ( n3250 & ~n3254 ) | ( n3250 & n4326 ) | ( ~n3254 & n4326 ) ;
  assign n4328 = ( n3562 & ~n3640 ) | ( n3562 & n4327 ) | ( ~n3640 & n4327 ) ;
  assign n4329 = ( n3925 & ~n3997 ) | ( n3925 & n4328 ) | ( ~n3997 & n4328 ) ;
  assign n4330 = ~n827 & n2004 ;
  assign n4331 = ( ~n853 & n2015 ) | ( ~n853 & n4330 ) | ( n2015 & n4330 ) ;
  assign n4332 = n850 | n4331 ;
  assign n4333 = n827 | n2008 ;
  assign n4334 = ~n846 & n4333 ;
  assign n4335 = ( ~n850 & n854 ) | ( ~n850 & n4334 ) | ( n854 & n4334 ) ;
  assign n4336 = ( n4329 & n4332 ) | ( n4329 & ~n4335 ) | ( n4332 & ~n4335 ) ;
  assign n4337 = ( n906 & ~n2557 ) | ( n906 & n4336 ) | ( ~n2557 & n4336 ) ;
  assign n4338 = n4317 & n4337 ;
  assign n4339 = x207 & ~n1271 ;
  assign n4340 = x81 | n1268 ;
  assign n4341 = ~n895 & n4340 ;
  assign n4342 = ( ~n867 & n910 ) | ( ~n867 & n4341 ) | ( n910 & n4341 ) ;
  assign n4343 = ( n938 & ~n956 ) | ( n938 & n4342 ) | ( ~n956 & n4342 ) ;
  assign n4344 = ( ~n1685 & n2038 ) | ( ~n1685 & n4343 ) | ( n2038 & n4343 ) ;
  assign n4345 = ( ~n2348 & n2575 ) | ( ~n2348 & n4344 ) | ( n2575 & n4344 ) ;
  assign n4346 = ( n1000 & ~n1705 ) | ( n1000 & n4345 ) | ( ~n1705 & n4345 ) ;
  assign n4347 = ( n2359 & ~n2599 ) | ( n2359 & n4346 ) | ( ~n2599 & n4346 ) ;
  assign n4348 = ( n2945 & ~n2949 ) | ( n2945 & n4347 ) | ( ~n2949 & n4347 ) ;
  assign n4349 = ( n3276 & ~n3280 ) | ( n3276 & n4348 ) | ( ~n3280 & n4348 ) ;
  assign n4350 = ( n3587 & ~n3665 ) | ( n3587 & n4349 ) | ( ~n3665 & n4349 ) ;
  assign n4351 = ( n3948 & ~n4020 ) | ( n3948 & n4350 ) | ( ~n4020 & n4350 ) ;
  assign n4352 = ~n1224 & n2113 ;
  assign n4353 = ( ~n1250 & n2124 ) | ( ~n1250 & n4352 ) | ( n2124 & n4352 ) ;
  assign n4354 = n1247 | n4353 ;
  assign n4355 = n1224 | n2117 ;
  assign n4356 = ~n1243 & n4355 ;
  assign n4357 = ( ~n1247 & n1251 ) | ( ~n1247 & n4356 ) | ( n1251 & n4356 ) ;
  assign n4358 = ( n4351 & n4354 ) | ( n4351 & ~n4357 ) | ( n4354 & ~n4357 ) ;
  assign n4359 = ( n1303 & ~n2626 ) | ( n1303 & n4358 ) | ( ~n2626 & n4358 ) ;
  assign n4360 = n4339 & n4359 ;
  assign n4361 = x208 & ~n496 ;
  assign n4362 = x82 | n470 ;
  assign n4363 = ~n1292 & n4362 ;
  assign n4364 = ( ~n1264 & n1307 ) | ( ~n1264 & n4363 ) | ( n1307 & n4363 ) ;
  assign n4365 = ( n1335 & ~n1353 ) | ( n1335 & n4364 ) | ( ~n1353 & n4364 ) ;
  assign n4366 = ( ~n1823 & n2147 ) | ( ~n1823 & n4365 ) | ( n2147 & n4365 ) ;
  assign n4367 = ( ~n2444 & n2644 ) | ( ~n2444 & n4366 ) | ( n2644 & n4366 ) ;
  assign n4368 = ( n1397 & ~n1843 ) | ( n1397 & n4367 ) | ( ~n1843 & n4367 ) ;
  assign n4369 = ( n2455 & ~n2668 ) | ( n2455 & n4368 ) | ( ~n2668 & n4368 ) ;
  assign n4370 = ( n2974 & ~n2978 ) | ( n2974 & n4369 ) | ( ~n2978 & n4369 ) ;
  assign n4371 = ( n3302 & ~n3306 ) | ( n3302 & n4370 ) | ( ~n3306 & n4370 ) ;
  assign n4372 = ( n3612 & ~n3689 ) | ( n3612 & n4371 ) | ( ~n3689 & n4371 ) ;
  assign n4373 = ( n3971 & ~n4043 ) | ( n3971 & n4372 ) | ( ~n4043 & n4372 ) ;
  assign n4374 = ~n455 & n2209 ;
  assign n4375 = ( ~n426 & n2220 ) | ( ~n426 & n4374 ) | ( n2220 & n4374 ) ;
  assign n4376 = n504 | n4375 ;
  assign n4377 = n455 | n2213 ;
  assign n4378 = ~n452 & n4377 ;
  assign n4379 = ( ~n504 & n1508 ) | ( ~n504 & n4378 ) | ( n1508 & n4378 ) ;
  assign n4380 = ( n4373 & n4376 ) | ( n4373 & ~n4379 ) | ( n4376 & ~n4379 ) ;
  assign n4381 = ( ~n495 & n1529 ) | ( ~n495 & n4380 ) | ( n1529 & n4380 ) ;
  assign n4382 = n4361 & n4381 ;
  assign n4383 = x209 & ~n894 ;
  assign n4384 = x83 | n868 ;
  assign n4385 = ~n468 & n4384 ;
  assign n4386 = ( ~n532 & n536 ) | ( ~n532 & n4385 ) | ( n536 & n4385 ) ;
  assign n4387 = ( ~n559 & n1536 ) | ( ~n559 & n4386 ) | ( n1536 & n4386 ) ;
  assign n4388 = ( ~n1937 & n2243 ) | ( ~n1937 & n4387 ) | ( n2243 & n4387 ) ;
  assign n4389 = ( ~n2514 & n2694 ) | ( ~n2514 & n4388 ) | ( n2694 & n4388 ) ;
  assign n4390 = ( n1558 & ~n1954 ) | ( n1558 & n4389 ) | ( ~n1954 & n4389 ) ;
  assign n4391 = ( n2524 & ~n2712 ) | ( n2524 & n4390 ) | ( ~n2712 & n4390 ) ;
  assign n4392 = ( n3003 & ~n3007 ) | ( n3003 & n4391 ) | ( ~n3007 & n4391 ) ;
  assign n4393 = ( n3328 & ~n3332 ) | ( n3328 & n4392 ) | ( ~n3332 & n4392 ) ;
  assign n4394 = ( n3637 & ~n3713 ) | ( n3637 & n4393 ) | ( ~n3713 & n4393 ) ;
  assign n4395 = ( n3994 & ~n4066 ) | ( n3994 & n4394 ) | ( ~n4066 & n4394 ) ;
  assign n4396 = ~n853 & n2305 ;
  assign n4397 = ( ~n824 & n2316 ) | ( ~n824 & n4396 ) | ( n2316 & n4396 ) ;
  assign n4398 = n902 | n4397 ;
  assign n4399 = n853 | n2309 ;
  assign n4400 = ~n850 & n4399 ;
  assign n4401 = ( ~n902 & n1647 ) | ( ~n902 & n4400 ) | ( n1647 & n4400 ) ;
  assign n4402 = ( n4395 & n4398 ) | ( n4395 & ~n4401 ) | ( n4398 & ~n4401 ) ;
  assign n4403 = ( ~n893 & n1668 ) | ( ~n893 & n4402 ) | ( n1668 & n4402 ) ;
  assign n4404 = n4383 & n4403 ;
  assign n4405 = x210 & ~n1291 ;
  assign n4406 = x84 | n1265 ;
  assign n4407 = ~n866 & n4406 ;
  assign n4408 = ( ~n930 & n934 ) | ( ~n930 & n4407 ) | ( n934 & n4407 ) ;
  assign n4409 = ( ~n957 & n1675 ) | ( ~n957 & n4408 ) | ( n1675 & n4408 ) ;
  assign n4410 = ( ~n2046 & n2339 ) | ( ~n2046 & n4409 ) | ( n2339 & n4409 ) ;
  assign n4411 = ( ~n2583 & n2738 ) | ( ~n2583 & n4410 ) | ( n2738 & n4410 ) ;
  assign n4412 = ( n1697 & ~n2063 ) | ( n1697 & n4411 ) | ( ~n2063 & n4411 ) ;
  assign n4413 = ( n2593 & ~n2756 ) | ( n2593 & n4412 ) | ( ~n2756 & n4412 ) ;
  assign n4414 = ( n3032 & ~n3036 ) | ( n3032 & n4413 ) | ( ~n3036 & n4413 ) ;
  assign n4415 = ( n3354 & ~n3358 ) | ( n3354 & n4414 ) | ( ~n3358 & n4414 ) ;
  assign n4416 = ( n3662 & ~n3737 ) | ( n3662 & n4415 ) | ( ~n3737 & n4415 ) ;
  assign n4417 = ( n4017 & ~n4089 ) | ( n4017 & n4416 ) | ( ~n4089 & n4416 ) ;
  assign n4418 = ~n1250 & n2401 ;
  assign n4419 = ( ~n1221 & n2412 ) | ( ~n1221 & n4418 ) | ( n2412 & n4418 ) ;
  assign n4420 = n1299 | n4419 ;
  assign n4421 = n1250 | n2405 ;
  assign n4422 = ~n1247 & n4421 ;
  assign n4423 = ( ~n1299 & n1785 ) | ( ~n1299 & n4422 ) | ( n1785 & n4422 ) ;
  assign n4424 = ( n4417 & n4420 ) | ( n4417 & ~n4423 ) | ( n4420 & ~n4423 ) ;
  assign n4425 = ( ~n1290 & n1806 ) | ( ~n1290 & n4424 ) | ( n1806 & n4424 ) ;
  assign n4426 = n4405 & n4425 ;
  assign n4427 = x211 & ~n467 ;
  assign n4428 = x85 | n533 ;
  assign n4429 = ~n1263 & n4428 ;
  assign n4430 = ( ~n1327 & n1331 ) | ( ~n1327 & n4429 ) | ( n1331 & n4429 ) ;
  assign n4431 = ( ~n1354 & n1813 ) | ( ~n1354 & n4430 ) | ( n1813 & n4430 ) ;
  assign n4432 = ( ~n2155 & n2435 ) | ( ~n2155 & n4431 ) | ( n2435 & n4431 ) ;
  assign n4433 = ( ~n2652 & n2782 ) | ( ~n2652 & n4432 ) | ( n2782 & n4432 ) ;
  assign n4434 = ( n1835 & ~n2172 ) | ( n1835 & n4433 ) | ( ~n2172 & n4433 ) ;
  assign n4435 = ( n2662 & ~n2800 ) | ( n2662 & n4434 ) | ( ~n2800 & n4434 ) ;
  assign n4436 = ( n3061 & ~n3065 ) | ( n3061 & n4435 ) | ( ~n3065 & n4435 ) ;
  assign n4437 = ( n3380 & ~n3384 ) | ( n3380 & n4436 ) | ( ~n3384 & n4436 ) ;
  assign n4438 = ( n3686 & ~n3761 ) | ( n3686 & n4437 ) | ( ~n3761 & n4437 ) ;
  assign n4439 = ( n4040 & ~n4112 ) | ( n4040 & n4438 ) | ( ~n4112 & n4438 ) ;
  assign n4440 = ( n465 & ~n484 ) | ( n465 & n505 ) | ( ~n484 & n505 ) ;
  assign n4441 = n487 | n4440 ;
  assign n4442 = n458 & ~n504 ;
  assign n4443 = ( ~n487 & n488 ) | ( ~n487 & n4442 ) | ( n488 & n4442 ) ;
  assign n4444 = ( n4439 & n4441 ) | ( n4439 & ~n4443 ) | ( n4441 & ~n4443 ) ;
  assign n4445 = ( ~n1522 & n1922 ) | ( ~n1522 & n4444 ) | ( n1922 & n4444 ) ;
  assign n4446 = n4427 & n4445 ;
  assign n4447 = x212 & ~n865 ;
  assign n4448 = x86 | n931 ;
  assign n4449 = ~n531 & n4448 ;
  assign n4450 = ( ~n529 & n1535 ) | ( ~n529 & n4449 ) | ( n1535 & n4449 ) ;
  assign n4451 = ( ~n1545 & n1929 ) | ( ~n1545 & n4450 ) | ( n1929 & n4450 ) ;
  assign n4452 = ( ~n2251 & n2505 ) | ( ~n2251 & n4451 ) | ( n2505 & n4451 ) ;
  assign n4453 = ( n600 & ~n617 ) | ( n600 & n4452 ) | ( ~n617 & n4452 ) ;
  assign n4454 = ( n1948 & ~n2268 ) | ( n1948 & n4453 ) | ( ~n2268 & n4453 ) ;
  assign n4455 = ( ~n648 & n2706 ) | ( ~n648 & n4454 ) | ( n2706 & n4454 ) ;
  assign n4456 = ( n3088 & ~n3092 ) | ( n3088 & n4455 ) | ( ~n3092 & n4455 ) ;
  assign n4457 = ( n3406 & ~n3410 ) | ( n3406 & n4456 ) | ( ~n3410 & n4456 ) ;
  assign n4458 = ( n3710 & ~n3785 ) | ( n3710 & n4457 ) | ( ~n3785 & n4457 ) ;
  assign n4459 = ( n4063 & ~n4135 ) | ( n4063 & n4458 ) | ( ~n4135 & n4458 ) ;
  assign n4460 = ( n863 & ~n882 ) | ( n863 & n903 ) | ( ~n882 & n903 ) ;
  assign n4461 = n885 | n4460 ;
  assign n4462 = n856 & ~n902 ;
  assign n4463 = ( ~n885 & n886 ) | ( ~n885 & n4462 ) | ( n886 & n4462 ) ;
  assign n4464 = ( n4459 & n4461 ) | ( n4459 & ~n4463 ) | ( n4461 & ~n4463 ) ;
  assign n4465 = ( ~n1661 & n2031 ) | ( ~n1661 & n4464 ) | ( n2031 & n4464 ) ;
  assign n4466 = n4447 & n4465 ;
  assign n4467 = x213 & ~n1262 ;
  assign n4468 = x87 | n1328 ;
  assign n4469 = ~n929 & n4468 ;
  assign n4470 = ( ~n927 & n1674 ) | ( ~n927 & n4469 ) | ( n1674 & n4469 ) ;
  assign n4471 = ( ~n1684 & n2038 ) | ( ~n1684 & n4470 ) | ( n2038 & n4470 ) ;
  assign n4472 = ( ~n2347 & n2574 ) | ( ~n2347 & n4471 ) | ( n2574 & n4471 ) ;
  assign n4473 = ( n998 & ~n1015 ) | ( n998 & n4472 ) | ( ~n1015 & n4472 ) ;
  assign n4474 = ( n2057 & ~n2364 ) | ( n2057 & n4473 ) | ( ~n2364 & n4473 ) ;
  assign n4475 = ( ~n1046 & n2750 ) | ( ~n1046 & n4474 ) | ( n2750 & n4474 ) ;
  assign n4476 = ( n3115 & ~n3119 ) | ( n3115 & n4475 ) | ( ~n3119 & n4475 ) ;
  assign n4477 = ( n3432 & ~n3436 ) | ( n3432 & n4476 ) | ( ~n3436 & n4476 ) ;
  assign n4478 = ( n3734 & ~n3809 ) | ( n3734 & n4477 ) | ( ~n3809 & n4477 ) ;
  assign n4479 = ( n4086 & ~n4158 ) | ( n4086 & n4478 ) | ( ~n4158 & n4478 ) ;
  assign n4480 = ( n1260 & ~n1279 ) | ( n1260 & n1300 ) | ( ~n1279 & n1300 ) ;
  assign n4481 = n1282 | n4480 ;
  assign n4482 = n1253 & ~n1299 ;
  assign n4483 = ( ~n1282 & n1283 ) | ( ~n1282 & n4482 ) | ( n1283 & n4482 ) ;
  assign n4484 = ( n4479 & n4481 ) | ( n4479 & ~n4483 ) | ( n4481 & ~n4483 ) ;
  assign n4485 = ( ~n1799 & n2140 ) | ( ~n1799 & n4484 ) | ( n2140 & n4484 ) ;
  assign n4486 = n4467 & n4485 ;
  assign n4487 = x214 & ~n530 ;
  assign n4488 = x88 | n537 ;
  assign n4489 = ~n1326 & n4488 ;
  assign n4490 = ( ~n1324 & n1812 ) | ( ~n1324 & n4489 ) | ( n1812 & n4489 ) ;
  assign n4491 = ( ~n1822 & n2147 ) | ( ~n1822 & n4490 ) | ( n2147 & n4490 ) ;
  assign n4492 = ( ~n2443 & n2643 ) | ( ~n2443 & n4491 ) | ( n2643 & n4491 ) ;
  assign n4493 = ( n1395 & ~n1412 ) | ( n1395 & n4492 ) | ( ~n1412 & n4492 ) ;
  assign n4494 = ( n2166 & ~n2460 ) | ( n2166 & n4493 ) | ( ~n2460 & n4493 ) ;
  assign n4495 = ( ~n1443 & n2794 ) | ( ~n1443 & n4494 ) | ( n2794 & n4494 ) ;
  assign n4496 = ( n3142 & ~n3146 ) | ( n3142 & n4495 ) | ( ~n3146 & n4495 ) ;
  assign n4497 = ( n3458 & ~n3462 ) | ( n3458 & n4496 ) | ( ~n3462 & n4496 ) ;
  assign n4498 = ( n3758 & ~n3833 ) | ( n3758 & n4497 ) | ( ~n3833 & n4497 ) ;
  assign n4499 = ( n4109 & ~n4180 ) | ( n4109 & n4498 ) | ( ~n4180 & n4498 ) ;
  assign n4500 = ( ~n491 & n1517 ) | ( ~n491 & n1526 ) | ( n1517 & n1526 ) ;
  assign n4501 = n481 | n4500 ;
  assign n4502 = ~n487 & n1510 ;
  assign n4503 = ( ~n481 & n492 ) | ( ~n481 & n4502 ) | ( n492 & n4502 ) ;
  assign n4504 = ( n4499 & n4501 ) | ( n4499 & ~n4503 ) | ( n4501 & ~n4503 ) ;
  assign n4505 = ( ~n1916 & n2236 ) | ( ~n1916 & n4504 ) | ( n2236 & n4504 ) ;
  assign n4506 = n4487 & n4505 ;
  assign n4507 = x215 & ~n928 ;
  assign n4508 = x89 | n935 ;
  assign n4509 = ~n528 & n4508 ;
  assign n4510 = ( ~n526 & n1928 ) | ( ~n526 & n4509 ) | ( n1928 & n4509 ) ;
  assign n4511 = ( ~n563 & n2243 ) | ( ~n563 & n4510 ) | ( n2243 & n4510 ) ;
  assign n4512 = ( ~n2513 & n2693 ) | ( ~n2513 & n4511 ) | ( n2693 & n4511 ) ;
  assign n4513 = ( n1556 & ~n1566 ) | ( n1556 & n4512 ) | ( ~n1566 & n4512 ) ;
  assign n4514 = ( n2262 & ~n2529 ) | ( n2262 & n4513 ) | ( ~n2529 & n4513 ) ;
  assign n4515 = ( ~n1582 & n2827 ) | ( ~n1582 & n4514 ) | ( n2827 & n4514 ) ;
  assign n4516 = ( n3169 & ~n3173 ) | ( n3169 & n4515 ) | ( ~n3173 & n4515 ) ;
  assign n4517 = ( n3484 & ~n3488 ) | ( n3484 & n4516 ) | ( ~n3488 & n4516 ) ;
  assign n4518 = ( n3782 & ~n3857 ) | ( n3782 & n4517 ) | ( ~n3857 & n4517 ) ;
  assign n4519 = ( n4132 & ~n4202 ) | ( n4132 & n4518 ) | ( ~n4202 & n4518 ) ;
  assign n4520 = ( ~n889 & n1656 ) | ( ~n889 & n1665 ) | ( n1656 & n1665 ) ;
  assign n4521 = n879 | n4520 ;
  assign n4522 = ~n885 & n1649 ;
  assign n4523 = ( ~n879 & n890 ) | ( ~n879 & n4522 ) | ( n890 & n4522 ) ;
  assign n4524 = ( n4519 & n4521 ) | ( n4519 & ~n4523 ) | ( n4521 & ~n4523 ) ;
  assign n4525 = ( ~n2025 & n2332 ) | ( ~n2025 & n4524 ) | ( n2332 & n4524 ) ;
  assign n4526 = n4507 & n4525 ;
  assign n4527 = x216 & ~n1325 ;
  assign n4528 = x90 | n1332 ;
  assign n4529 = ~n926 & n4528 ;
  assign n4530 = ( ~n924 & n2037 ) | ( ~n924 & n4529 ) | ( n2037 & n4529 ) ;
  assign n4531 = ( ~n961 & n2339 ) | ( ~n961 & n4530 ) | ( n2339 & n4530 ) ;
  assign n4532 = ( ~n2582 & n2737 ) | ( ~n2582 & n4531 ) | ( n2737 & n4531 ) ;
  assign n4533 = ( n1695 & ~n1705 ) | ( n1695 & n4532 ) | ( ~n1705 & n4532 ) ;
  assign n4534 = ( n2358 & ~n2598 ) | ( n2358 & n4533 ) | ( ~n2598 & n4533 ) ;
  assign n4535 = ( ~n1721 & n2857 ) | ( ~n1721 & n4534 ) | ( n2857 & n4534 ) ;
  assign n4536 = ( n3196 & ~n3200 ) | ( n3196 & n4535 ) | ( ~n3200 & n4535 ) ;
  assign n4537 = ( n3510 & ~n3514 ) | ( n3510 & n4536 ) | ( ~n3514 & n4536 ) ;
  assign n4538 = ( n3806 & ~n3881 ) | ( n3806 & n4537 ) | ( ~n3881 & n4537 ) ;
  assign n4539 = ( n4155 & ~n4224 ) | ( n4155 & n4538 ) | ( ~n4224 & n4538 ) ;
  assign n4540 = ( ~n1286 & n1794 ) | ( ~n1286 & n1803 ) | ( n1794 & n1803 ) ;
  assign n4541 = n1276 | n4540 ;
  assign n4542 = ~n1282 & n1787 ;
  assign n4543 = ( ~n1276 & n1287 ) | ( ~n1276 & n4542 ) | ( n1287 & n4542 ) ;
  assign n4544 = ( n4539 & n4541 ) | ( n4539 & ~n4543 ) | ( n4541 & ~n4543 ) ;
  assign n4545 = ( ~n2134 & n2428 ) | ( ~n2134 & n4544 ) | ( n2428 & n4544 ) ;
  assign n4546 = n4527 & n4545 ;
  assign n4547 = x217 & ~n527 ;
  assign n4548 = x91 | n542 ;
  assign n4549 = ~n1323 & n4548 ;
  assign n4550 = ( ~n1321 & n2146 ) | ( ~n1321 & n4549 ) | ( n2146 & n4549 ) ;
  assign n4551 = ( ~n1358 & n2435 ) | ( ~n1358 & n4550 ) | ( n2435 & n4550 ) ;
  assign n4552 = ( ~n2651 & n2781 ) | ( ~n2651 & n4551 ) | ( n2781 & n4551 ) ;
  assign n4553 = ( n1833 & ~n1843 ) | ( n1833 & n4552 ) | ( ~n1843 & n4552 ) ;
  assign n4554 = ( n2454 & ~n2667 ) | ( n2454 & n4553 ) | ( ~n2667 & n4553 ) ;
  assign n4555 = ( ~n1856 & n2887 ) | ( ~n1856 & n4554 ) | ( n2887 & n4554 ) ;
  assign n4556 = ( n3223 & ~n3227 ) | ( n3223 & n4555 ) | ( ~n3227 & n4555 ) ;
  assign n4557 = ( n3536 & ~n3540 ) | ( n3536 & n4556 ) | ( ~n3540 & n4556 ) ;
  assign n4558 = ( n3830 & ~n3904 ) | ( n3830 & n4557 ) | ( ~n3904 & n4557 ) ;
  assign n4559 = ( n4178 & ~n4246 ) | ( n4178 & n4558 ) | ( ~n4246 & n4558 ) ;
  assign n4560 = ( ~n478 & n1912 ) | ( ~n478 & n1919 ) | ( n1912 & n1919 ) ;
  assign n4561 = n475 | n4560 ;
  assign n4562 = ~n481 & n1905 ;
  assign n4563 = ( ~n475 & n1519 ) | ( ~n475 & n4562 ) | ( n1519 & n4562 ) ;
  assign n4564 = ( n4559 & n4561 ) | ( n4559 & ~n4563 ) | ( n4561 & ~n4563 ) ;
  assign n4565 = ( ~n2230 & n2499 ) | ( ~n2230 & n4564 ) | ( n2499 & n4564 ) ;
  assign n4566 = n4547 & n4565 ;
  assign n4567 = x218 & ~n925 ;
  assign n4568 = x92 | n940 ;
  assign n4569 = ~n525 & n4568 ;
  assign n4570 = ( ~n523 & n2242 ) | ( ~n523 & n4569 ) | ( n2242 & n4569 ) ;
  assign n4571 = ( ~n1549 & n2505 ) | ( ~n1549 & n4570 ) | ( n2505 & n4570 ) ;
  assign n4572 = ( n599 & ~n616 ) | ( n599 & n4571 ) | ( ~n616 & n4571 ) ;
  assign n4573 = ( n1946 & ~n1954 ) | ( n1946 & n4572 ) | ( ~n1954 & n4572 ) ;
  assign n4574 = ( n2523 & ~n2711 ) | ( n2523 & n4573 ) | ( ~n2711 & n4573 ) ;
  assign n4575 = ( ~n1965 & n2916 ) | ( ~n1965 & n4574 ) | ( n2916 & n4574 ) ;
  assign n4576 = ( n3249 & ~n3253 ) | ( n3249 & n4575 ) | ( ~n3253 & n4575 ) ;
  assign n4577 = ( n3561 & ~n3565 ) | ( n3561 & n4576 ) | ( ~n3565 & n4576 ) ;
  assign n4578 = ( n3854 & ~n3927 ) | ( n3854 & n4577 ) | ( ~n3927 & n4577 ) ;
  assign n4579 = ( n4200 & ~n4268 ) | ( n4200 & n4578 ) | ( ~n4268 & n4578 ) ;
  assign n4580 = ( ~n876 & n2021 ) | ( ~n876 & n2028 ) | ( n2021 & n2028 ) ;
  assign n4581 = n873 | n4580 ;
  assign n4582 = ~n879 & n2014 ;
  assign n4583 = ( ~n873 & n1658 ) | ( ~n873 & n4582 ) | ( n1658 & n4582 ) ;
  assign n4584 = ( n4579 & n4581 ) | ( n4579 & ~n4583 ) | ( n4581 & ~n4583 ) ;
  assign n4585 = ( ~n2326 & n2568 ) | ( ~n2326 & n4584 ) | ( n2568 & n4584 ) ;
  assign n4586 = n4567 & n4585 ;
  assign n4587 = x219 & ~n1322 ;
  assign n4588 = x93 | n1337 ;
  assign n4589 = ~n923 & n4588 ;
  assign n4590 = ( ~n921 & n2338 ) | ( ~n921 & n4589 ) | ( n2338 & n4589 ) ;
  assign n4591 = ( ~n1688 & n2574 ) | ( ~n1688 & n4590 ) | ( n2574 & n4590 ) ;
  assign n4592 = ( n997 & ~n1014 ) | ( n997 & n4591 ) | ( ~n1014 & n4591 ) ;
  assign n4593 = ( n2055 & ~n2063 ) | ( n2055 & n4592 ) | ( ~n2063 & n4592 ) ;
  assign n4594 = ( n2592 & ~n2755 ) | ( n2592 & n4593 ) | ( ~n2755 & n4593 ) ;
  assign n4595 = ( ~n2074 & n2945 ) | ( ~n2074 & n4594 ) | ( n2945 & n4594 ) ;
  assign n4596 = ( n3275 & ~n3279 ) | ( n3275 & n4595 ) | ( ~n3279 & n4595 ) ;
  assign n4597 = ( n3586 & ~n3590 ) | ( n3586 & n4596 ) | ( ~n3590 & n4596 ) ;
  assign n4598 = ( n3878 & ~n3950 ) | ( n3878 & n4597 ) | ( ~n3950 & n4597 ) ;
  assign n4599 = ( n4222 & ~n4290 ) | ( n4222 & n4598 ) | ( ~n4290 & n4598 ) ;
  assign n4600 = ( ~n1273 & n2130 ) | ( ~n1273 & n2137 ) | ( n2130 & n2137 ) ;
  assign n4601 = n1270 | n4600 ;
  assign n4602 = ~n1276 & n2123 ;
  assign n4603 = ( ~n1270 & n1796 ) | ( ~n1270 & n4602 ) | ( n1796 & n4602 ) ;
  assign n4604 = ( n4599 & n4601 ) | ( n4599 & ~n4603 ) | ( n4601 & ~n4603 ) ;
  assign n4605 = ( ~n2422 & n2637 ) | ( ~n2422 & n4604 ) | ( n2637 & n4604 ) ;
  assign n4606 = n4587 & n4605 ;
  assign n4607 = x220 & ~n524 ;
  assign n4608 = x94 | n547 ;
  assign n4609 = ~n1320 & n4608 ;
  assign n4610 = ( ~n1318 & n2434 ) | ( ~n1318 & n4609 ) | ( n2434 & n4609 ) ;
  assign n4611 = ( ~n1826 & n2643 ) | ( ~n1826 & n4610 ) | ( n2643 & n4610 ) ;
  assign n4612 = ( n1394 & ~n1411 ) | ( n1394 & n4611 ) | ( ~n1411 & n4611 ) ;
  assign n4613 = ( n2164 & ~n2172 ) | ( n2164 & n4612 ) | ( ~n2172 & n4612 ) ;
  assign n4614 = ( n2661 & ~n2799 ) | ( n2661 & n4613 ) | ( ~n2799 & n4613 ) ;
  assign n4615 = ( ~n2182 & n2974 ) | ( ~n2182 & n4614 ) | ( n2974 & n4614 ) ;
  assign n4616 = ( n3301 & ~n3305 ) | ( n3301 & n4615 ) | ( ~n3305 & n4615 ) ;
  assign n4617 = ( n3611 & ~n3615 ) | ( n3611 & n4616 ) | ( ~n3615 & n4616 ) ;
  assign n4618 = ( n3901 & ~n3973 ) | ( n3901 & n4617 ) | ( ~n3973 & n4617 ) ;
  assign n4619 = ( n4244 & ~n4312 ) | ( n4244 & n4618 ) | ( ~n4312 & n4618 ) ;
  assign n4620 = ( ~n498 & n2226 ) | ( ~n498 & n2233 ) | ( n2226 & n2233 ) ;
  assign n4621 = n472 | n4620 ;
  assign n4622 = ~n475 & n2219 ;
  assign n4623 = ( ~n472 & n499 ) | ( ~n472 & n4622 ) | ( n499 & n4622 ) ;
  assign n4624 = ( n4619 & n4621 ) | ( n4619 & ~n4623 ) | ( n4621 & ~n4623 ) ;
  assign n4625 = ( n545 & ~n2494 ) | ( n545 & n4624 ) | ( ~n2494 & n4624 ) ;
  assign n4626 = n4607 & n4625 ;
  assign n4627 = x221 & ~n922 ;
  assign n4628 = x95 | n945 ;
  assign n4629 = ~n522 & n4628 ;
  assign n4630 = ( ~n520 & n555 ) | ( ~n520 & n4629 ) | ( n555 & n4629 ) ;
  assign n4631 = ( ~n614 & n2693 ) | ( ~n614 & n4630 ) | ( n2693 & n4630 ) ;
  assign n4632 = ( n1555 & ~n1565 ) | ( n1555 & n4631 ) | ( ~n1565 & n4631 ) ;
  assign n4633 = ( n2260 & ~n2268 ) | ( n2260 & n4632 ) | ( ~n2268 & n4632 ) ;
  assign n4634 = ( ~n644 & n2705 ) | ( ~n644 & n4633 ) | ( n2705 & n4633 ) ;
  assign n4635 = ( ~n2278 & n3003 ) | ( ~n2278 & n4634 ) | ( n3003 & n4634 ) ;
  assign n4636 = ( n3327 & ~n3331 ) | ( n3327 & n4635 ) | ( ~n3331 & n4635 ) ;
  assign n4637 = ( n3636 & ~n3640 ) | ( n3636 & n4636 ) | ( ~n3640 & n4636 ) ;
  assign n4638 = ( n3924 & ~n3996 ) | ( n3924 & n4637 ) | ( ~n3996 & n4637 ) ;
  assign n4639 = ( n4266 & ~n4334 ) | ( n4266 & n4638 ) | ( ~n4334 & n4638 ) ;
  assign n4640 = ( ~n896 & n2322 ) | ( ~n896 & n2329 ) | ( n2322 & n2329 ) ;
  assign n4641 = n870 | n4640 ;
  assign n4642 = ~n873 & n2315 ;
  assign n4643 = ( ~n870 & n897 ) | ( ~n870 & n4642 ) | ( n897 & n4642 ) ;
  assign n4644 = ( n4639 & n4641 ) | ( n4639 & ~n4643 ) | ( n4641 & ~n4643 ) ;
  assign n4645 = ( n943 & ~n2563 ) | ( n943 & n4644 ) | ( ~n2563 & n4644 ) ;
  assign n4646 = n4627 & n4645 ;
  assign n4647 = x222 & ~n1319 ;
  assign n4648 = x96 | n1342 ;
  assign n4649 = ~n920 & n4648 ;
  assign n4650 = ( ~n918 & n953 ) | ( ~n918 & n4649 ) | ( n953 & n4649 ) ;
  assign n4651 = ( ~n1012 & n2737 ) | ( ~n1012 & n4650 ) | ( n2737 & n4650 ) ;
  assign n4652 = ( n1694 & ~n1704 ) | ( n1694 & n4651 ) | ( ~n1704 & n4651 ) ;
  assign n4653 = ( n2356 & ~n2364 ) | ( n2356 & n4652 ) | ( ~n2364 & n4652 ) ;
  assign n4654 = ( ~n1042 & n2749 ) | ( ~n1042 & n4653 ) | ( n2749 & n4653 ) ;
  assign n4655 = ( ~n2374 & n3032 ) | ( ~n2374 & n4654 ) | ( n3032 & n4654 ) ;
  assign n4656 = ( n3353 & ~n3357 ) | ( n3353 & n4655 ) | ( ~n3357 & n4655 ) ;
  assign n4657 = ( n3661 & ~n3665 ) | ( n3661 & n4656 ) | ( ~n3665 & n4656 ) ;
  assign n4658 = ( n3947 & ~n4019 ) | ( n3947 & n4657 ) | ( ~n4019 & n4657 ) ;
  assign n4659 = ( n4288 & ~n4356 ) | ( n4288 & n4658 ) | ( ~n4356 & n4658 ) ;
  assign n4660 = ( ~n1293 & n2418 ) | ( ~n1293 & n2425 ) | ( n2418 & n2425 ) ;
  assign n4661 = n1267 | n4660 ;
  assign n4662 = ~n1270 & n2411 ;
  assign n4663 = ( ~n1267 & n1294 ) | ( ~n1267 & n4662 ) | ( n1294 & n4662 ) ;
  assign n4664 = ( n4659 & n4661 ) | ( n4659 & ~n4663 ) | ( n4661 & ~n4663 ) ;
  assign n4665 = ( n1340 & ~n2632 ) | ( n1340 & n4664 ) | ( ~n2632 & n4664 ) ;
  assign n4666 = n4647 & n4665 ;
  assign n4667 = x223 & ~n521 ;
  assign n4668 = x97 | n552 ;
  assign n4669 = ~n1317 & n4668 ;
  assign n4670 = ( ~n1315 & n1350 ) | ( ~n1315 & n4669 ) | ( n1350 & n4669 ) ;
  assign n4671 = ( ~n1409 & n2781 ) | ( ~n1409 & n4670 ) | ( n2781 & n4670 ) ;
  assign n4672 = ( n1832 & ~n1842 ) | ( n1832 & n4671 ) | ( ~n1842 & n4671 ) ;
  assign n4673 = ( n2452 & ~n2460 ) | ( n2452 & n4672 ) | ( ~n2460 & n4672 ) ;
  assign n4674 = ( ~n1439 & n2793 ) | ( ~n1439 & n4673 ) | ( n2793 & n4673 ) ;
  assign n4675 = ( ~n2470 & n3061 ) | ( ~n2470 & n4674 ) | ( n3061 & n4674 ) ;
  assign n4676 = ( n3379 & ~n3383 ) | ( n3379 & n4675 ) | ( ~n3383 & n4675 ) ;
  assign n4677 = ( n3685 & ~n3689 ) | ( n3685 & n4676 ) | ( ~n3689 & n4676 ) ;
  assign n4678 = ( n3970 & ~n4042 ) | ( n3970 & n4677 ) | ( ~n4042 & n4677 ) ;
  assign n4679 = ( n4310 & ~n4378 ) | ( n4310 & n4678 ) | ( ~n4378 & n4678 ) ;
  assign n4680 = n513 | n535 ;
  assign n4681 = ~n472 & n2490 ;
  assign n4682 = ( ~n535 & n1523 ) | ( ~n535 & n4681 ) | ( n1523 & n4681 ) ;
  assign n4683 = ( n4679 & n4680 ) | ( n4679 & ~n4682 ) | ( n4680 & ~n4682 ) ;
  assign n4684 = ( ~n562 & n1538 ) | ( ~n562 & n4683 ) | ( n1538 & n4683 ) ;
  assign n4685 = n4667 & n4684 ;
  assign n4686 = x224 & ~n919 ;
  assign n4687 = x98 | n950 ;
  assign n4688 = ~n519 & n4687 ;
  assign n4689 = ( ~n613 & n1542 ) | ( ~n613 & n4688 ) | ( n1542 & n4688 ) ;
  assign n4690 = ( n599 & ~n615 ) | ( n599 & n4689 ) | ( ~n615 & n4689 ) ;
  assign n4691 = ( n1945 & ~n1953 ) | ( n1945 & n4690 ) | ( ~n1953 & n4690 ) ;
  assign n4692 = ( n2521 & ~n2529 ) | ( n2521 & n4691 ) | ( ~n2529 & n4691 ) ;
  assign n4693 = ( ~n1579 & n2826 ) | ( ~n1579 & n4692 ) | ( n2826 & n4692 ) ;
  assign n4694 = ( ~n2539 & n3088 ) | ( ~n2539 & n4693 ) | ( n3088 & n4693 ) ;
  assign n4695 = ( n3405 & ~n3409 ) | ( n3405 & n4694 ) | ( ~n3409 & n4694 ) ;
  assign n4696 = ( n3709 & ~n3713 ) | ( n3709 & n4695 ) | ( ~n3713 & n4695 ) ;
  assign n4697 = ( n3993 & ~n4065 ) | ( n3993 & n4696 ) | ( ~n4065 & n4696 ) ;
  assign n4698 = ( n4332 & ~n4400 ) | ( n4332 & n4697 ) | ( ~n4400 & n4697 ) ;
  assign n4699 = n911 | n933 ;
  assign n4700 = ~n870 & n2559 ;
  assign n4701 = ( ~n933 & n1662 ) | ( ~n933 & n4700 ) | ( n1662 & n4700 ) ;
  assign n4702 = ( n4698 & n4699 ) | ( n4698 & ~n4701 ) | ( n4699 & ~n4701 ) ;
  assign n4703 = ( ~n960 & n1677 ) | ( ~n960 & n4702 ) | ( n1677 & n4702 ) ;
  assign n4704 = n4686 & n4703 ;
  assign n4705 = x225 & ~n1316 ;
  assign n4706 = x99 | n1347 ;
  assign n4707 = ~n917 & n4706 ;
  assign n4708 = ( ~n1011 & n1681 ) | ( ~n1011 & n4707 ) | ( n1681 & n4707 ) ;
  assign n4709 = ( n997 & ~n1013 ) | ( n997 & n4708 ) | ( ~n1013 & n4708 ) ;
  assign n4710 = ( n2054 & ~n2062 ) | ( n2054 & n4709 ) | ( ~n2062 & n4709 ) ;
  assign n4711 = ( n2590 & ~n2598 ) | ( n2590 & n4710 ) | ( ~n2598 & n4710 ) ;
  assign n4712 = ( ~n1718 & n2856 ) | ( ~n1718 & n4711 ) | ( n2856 & n4711 ) ;
  assign n4713 = ( ~n2608 & n3115 ) | ( ~n2608 & n4712 ) | ( n3115 & n4712 ) ;
  assign n4714 = ( n3431 & ~n3435 ) | ( n3431 & n4713 ) | ( ~n3435 & n4713 ) ;
  assign n4715 = ( n3733 & ~n3737 ) | ( n3733 & n4714 ) | ( ~n3737 & n4714 ) ;
  assign n4716 = ( n4016 & ~n4088 ) | ( n4016 & n4715 ) | ( ~n4088 & n4715 ) ;
  assign n4717 = ( n4354 & ~n4422 ) | ( n4354 & n4716 ) | ( ~n4422 & n4716 ) ;
  assign n4718 = n1308 | n1330 ;
  assign n4719 = ~n1267 & n2628 ;
  assign n4720 = ( ~n1330 & n1800 ) | ( ~n1330 & n4719 ) | ( n1800 & n4719 ) ;
  assign n4721 = ( n4717 & n4718 ) | ( n4717 & ~n4720 ) | ( n4718 & ~n4720 ) ;
  assign n4722 = ( ~n1357 & n1815 ) | ( ~n1357 & n4721 ) | ( n1815 & n4721 ) ;
  assign n4723 = n4705 & n4722 ;
  assign n4724 = x226 & ~n518 ;
  assign n4725 = x100 | n515 ;
  assign n4726 = ~n1314 & n4725 ;
  assign n4727 = ( ~n1408 & n1819 ) | ( ~n1408 & n4726 ) | ( n1819 & n4726 ) ;
  assign n4728 = ( n1394 & ~n1410 ) | ( n1394 & n4727 ) | ( ~n1410 & n4727 ) ;
  assign n4729 = ( n2163 & ~n2171 ) | ( n2163 & n4728 ) | ( ~n2171 & n4728 ) ;
  assign n4730 = ( n2659 & ~n2667 ) | ( n2659 & n4729 ) | ( ~n2667 & n4729 ) ;
  assign n4731 = ( ~n1855 & n2886 ) | ( ~n1855 & n4730 ) | ( n2886 & n4730 ) ;
  assign n4732 = ( ~n2676 & n3142 ) | ( ~n2676 & n4731 ) | ( n3142 & n4731 ) ;
  assign n4733 = ( n3457 & ~n3461 ) | ( n3457 & n4732 ) | ( ~n3461 & n4732 ) ;
  assign n4734 = ( n3757 & ~n3761 ) | ( n3757 & n4733 ) | ( ~n3761 & n4733 ) ;
  assign n4735 = ( n4039 & ~n4111 ) | ( n4039 & n4734 ) | ( ~n4111 & n4734 ) ;
  assign n4736 = ( n4376 & ~n4442 ) | ( n4376 & n4735 ) | ( ~n4442 & n4735 ) ;
  assign n4737 = n539 | n1533 ;
  assign n4738 = n501 & ~n535 ;
  assign n4739 = ( ~n539 & n558 ) | ( ~n539 & n4738 ) | ( n558 & n4738 ) ;
  assign n4740 = ( n4736 & n4737 ) | ( n4736 & ~n4739 ) | ( n4737 & ~n4739 ) ;
  assign n4741 = ( ~n1548 & n1931 ) | ( ~n1548 & n4740 ) | ( n1931 & n4740 ) ;
  assign n4742 = n4724 & n4741 ;
  assign n4743 = x227 & ~n916 ;
  assign n4744 = x101 | n913 ;
  assign n4745 = ~n612 & n4744 ;
  assign n4746 = ( ~n594 & n598 ) | ( ~n594 & n4745 ) | ( n598 & n4745 ) ;
  assign n4747 = ( n1555 & ~n1564 ) | ( n1555 & n4746 ) | ( ~n1564 & n4746 ) ;
  assign n4748 = ( n2259 & ~n2267 ) | ( n2259 & n4747 ) | ( ~n2267 & n4747 ) ;
  assign n4749 = ( n2703 & ~n2711 ) | ( n2703 & n4748 ) | ( ~n2711 & n4748 ) ;
  assign n4750 = ( ~n1964 & n2915 ) | ( ~n1964 & n4749 ) | ( n2915 & n4749 ) ;
  assign n4751 = ( ~n2720 & n3169 ) | ( ~n2720 & n4750 ) | ( n3169 & n4750 ) ;
  assign n4752 = ( n3483 & ~n3487 ) | ( n3483 & n4751 ) | ( ~n3487 & n4751 ) ;
  assign n4753 = ( n3781 & ~n3785 ) | ( n3781 & n4752 ) | ( ~n3785 & n4752 ) ;
  assign n4754 = ( n4062 & ~n4134 ) | ( n4062 & n4753 ) | ( ~n4134 & n4753 ) ;
  assign n4755 = ( n4398 & ~n4462 ) | ( n4398 & n4754 ) | ( ~n4462 & n4754 ) ;
  assign n4756 = n937 | n1672 ;
  assign n4757 = n899 & ~n933 ;
  assign n4758 = ( ~n937 & n956 ) | ( ~n937 & n4757 ) | ( n956 & n4757 ) ;
  assign n4759 = ( n4755 & n4756 ) | ( n4755 & ~n4758 ) | ( n4756 & ~n4758 ) ;
  assign n4760 = ( ~n1687 & n2040 ) | ( ~n1687 & n4759 ) | ( n2040 & n4759 ) ;
  assign n4761 = n4743 & n4760 ;
  assign n4762 = x228 & ~n1313 ;
  assign n4763 = x102 | n1310 ;
  assign n4764 = ~n1010 & n4763 ;
  assign n4765 = ( ~n992 & n996 ) | ( ~n992 & n4764 ) | ( n996 & n4764 ) ;
  assign n4766 = ( n1694 & ~n1703 ) | ( n1694 & n4765 ) | ( ~n1703 & n4765 ) ;
  assign n4767 = ( n2355 & ~n2363 ) | ( n2355 & n4766 ) | ( ~n2363 & n4766 ) ;
  assign n4768 = ( n2747 & ~n2755 ) | ( n2747 & n4767 ) | ( ~n2755 & n4767 ) ;
  assign n4769 = ( ~n2073 & n2944 ) | ( ~n2073 & n4768 ) | ( n2944 & n4768 ) ;
  assign n4770 = ( ~n2764 & n3196 ) | ( ~n2764 & n4769 ) | ( n3196 & n4769 ) ;
  assign n4771 = ( n3509 & ~n3513 ) | ( n3509 & n4770 ) | ( ~n3513 & n4770 ) ;
  assign n4772 = ( n3805 & ~n3809 ) | ( n3805 & n4771 ) | ( ~n3809 & n4771 ) ;
  assign n4773 = ( n4085 & ~n4157 ) | ( n4085 & n4772 ) | ( ~n4157 & n4772 ) ;
  assign n4774 = ( n4420 & ~n4482 ) | ( n4420 & n4773 ) | ( ~n4482 & n4773 ) ;
  assign n4775 = n1334 | n1810 ;
  assign n4776 = n1296 & ~n1330 ;
  assign n4777 = ( ~n1334 & n1353 ) | ( ~n1334 & n4776 ) | ( n1353 & n4776 ) ;
  assign n4778 = ( n4774 & n4775 ) | ( n4774 & ~n4777 ) | ( n4775 & ~n4777 ) ;
  assign n4779 = ( ~n1825 & n2149 ) | ( ~n1825 & n4778 ) | ( n2149 & n4778 ) ;
  assign n4780 = n4762 & n4779 ;
  assign n4781 = x229 & ~n611 ;
  assign n4782 = x103 | n595 ;
  assign n4783 = ~n1407 & n4782 ;
  assign n4784 = ( ~n1389 & n1393 ) | ( ~n1389 & n4783 ) | ( n1393 & n4783 ) ;
  assign n4785 = ( n1832 & ~n1841 ) | ( n1832 & n4784 ) | ( ~n1841 & n4784 ) ;
  assign n4786 = ( n2451 & ~n2459 ) | ( n2451 & n4785 ) | ( ~n2459 & n4785 ) ;
  assign n4787 = ( n2791 & ~n2799 ) | ( n2791 & n4786 ) | ( ~n2799 & n4786 ) ;
  assign n4788 = ( ~n2181 & n2973 ) | ( ~n2181 & n4787 ) | ( n2973 & n4787 ) ;
  assign n4789 = ( ~n2808 & n3223 ) | ( ~n2808 & n4788 ) | ( n3223 & n4788 ) ;
  assign n4790 = ( n3535 & ~n3539 ) | ( n3535 & n4789 ) | ( ~n3539 & n4789 ) ;
  assign n4791 = ( n3829 & ~n3833 ) | ( n3829 & n4790 ) | ( ~n3833 & n4790 ) ;
  assign n4792 = ( n4108 & ~n4179 ) | ( n4108 & n4791 ) | ( ~n4179 & n4791 ) ;
  assign n4793 = ( n4441 & ~n4502 ) | ( n4441 & n4792 ) | ( ~n4502 & n4792 ) ;
  assign n4794 = n544 | n1926 ;
  assign n4795 = ~n539 & n1525 ;
  assign n4796 = ( ~n544 & n559 ) | ( ~n544 & n4795 ) | ( n559 & n4795 ) ;
  assign n4797 = ( n4793 & n4794 ) | ( n4793 & ~n4796 ) | ( n4794 & ~n4796 ) ;
  assign n4798 = ( ~n1939 & n2245 ) | ( ~n1939 & n4797 ) | ( n2245 & n4797 ) ;
  assign n4799 = n4781 & n4798 ;
  assign n4800 = x230 & ~n1009 ;
  assign n4801 = x104 | n993 ;
  assign n4802 = ~n593 & n4801 ;
  assign n4803 = ( ~n588 & n1554 ) | ( ~n588 & n4802 ) | ( n1554 & n4802 ) ;
  assign n4804 = ( ~n619 & n1945 ) | ( ~n619 & n4803 ) | ( n1945 & n4803 ) ;
  assign n4805 = ( n2520 & ~n2528 ) | ( n2520 & n4804 ) | ( ~n2528 & n4804 ) ;
  assign n4806 = ( ~n644 & n651 ) | ( ~n644 & n4805 ) | ( n651 & n4805 ) ;
  assign n4807 = ( ~n2277 & n3002 ) | ( ~n2277 & n4806 ) | ( n3002 & n4806 ) ;
  assign n4808 = ( ~n2838 & n3249 ) | ( ~n2838 & n4807 ) | ( n3249 & n4807 ) ;
  assign n4809 = ( n3560 & ~n3564 ) | ( n3560 & n4808 ) | ( ~n3564 & n4808 ) ;
  assign n4810 = ( n3853 & ~n3857 ) | ( n3853 & n4809 ) | ( ~n3857 & n4809 ) ;
  assign n4811 = ( n4131 & ~n4201 ) | ( n4131 & n4810 ) | ( ~n4201 & n4810 ) ;
  assign n4812 = ( n4461 & ~n4522 ) | ( n4461 & n4811 ) | ( ~n4522 & n4811 ) ;
  assign n4813 = n942 | n2035 ;
  assign n4814 = ~n937 & n1664 ;
  assign n4815 = ( ~n942 & n957 ) | ( ~n942 & n4814 ) | ( n957 & n4814 ) ;
  assign n4816 = ( n4812 & n4813 ) | ( n4812 & ~n4815 ) | ( n4813 & ~n4815 ) ;
  assign n4817 = ( ~n2048 & n2341 ) | ( ~n2048 & n4816 ) | ( n2341 & n4816 ) ;
  assign n4818 = n4800 & n4817 ;
  assign n4819 = x231 & ~n1406 ;
  assign n4820 = x105 | n1390 ;
  assign n4821 = ~n991 & n4820 ;
  assign n4822 = ( ~n986 & n1693 ) | ( ~n986 & n4821 ) | ( n1693 & n4821 ) ;
  assign n4823 = ( ~n1017 & n2054 ) | ( ~n1017 & n4822 ) | ( n2054 & n4822 ) ;
  assign n4824 = ( n2589 & ~n2597 ) | ( n2589 & n4823 ) | ( ~n2597 & n4823 ) ;
  assign n4825 = ( ~n1042 & n1049 ) | ( ~n1042 & n4824 ) | ( n1049 & n4824 ) ;
  assign n4826 = ( ~n2373 & n3031 ) | ( ~n2373 & n4825 ) | ( n3031 & n4825 ) ;
  assign n4827 = ( ~n2868 & n3275 ) | ( ~n2868 & n4826 ) | ( n3275 & n4826 ) ;
  assign n4828 = ( n3585 & ~n3589 ) | ( n3585 & n4827 ) | ( ~n3589 & n4827 ) ;
  assign n4829 = ( n3877 & ~n3881 ) | ( n3877 & n4828 ) | ( ~n3881 & n4828 ) ;
  assign n4830 = ( n4154 & ~n4223 ) | ( n4154 & n4829 ) | ( ~n4223 & n4829 ) ;
  assign n4831 = ( n4481 & ~n4542 ) | ( n4481 & n4830 ) | ( ~n4542 & n4830 ) ;
  assign n4832 = n1339 | n2144 ;
  assign n4833 = ~n1334 & n1802 ;
  assign n4834 = ( ~n1339 & n1354 ) | ( ~n1339 & n4833 ) | ( n1354 & n4833 ) ;
  assign n4835 = ( n4831 & n4832 ) | ( n4831 & ~n4834 ) | ( n4832 & ~n4834 ) ;
  assign n4836 = ( ~n2157 & n2437 ) | ( ~n2157 & n4835 ) | ( n2437 & n4835 ) ;
  assign n4837 = n4819 & n4836 ;
  assign n4838 = x232 & ~n592 ;
  assign n4839 = x106 | n589 ;
  assign n4840 = ~n1388 & n4839 ;
  assign n4841 = ( ~n1383 & n1831 ) | ( ~n1383 & n4840 ) | ( n1831 & n4840 ) ;
  assign n4842 = ( ~n1414 & n2163 ) | ( ~n1414 & n4841 ) | ( n2163 & n4841 ) ;
  assign n4843 = ( n2658 & ~n2666 ) | ( n2658 & n4842 ) | ( ~n2666 & n4842 ) ;
  assign n4844 = ( ~n1439 & n1446 ) | ( ~n1439 & n4843 ) | ( n1446 & n4843 ) ;
  assign n4845 = ( ~n2469 & n3060 ) | ( ~n2469 & n4844 ) | ( n3060 & n4844 ) ;
  assign n4846 = ( ~n2897 & n3301 ) | ( ~n2897 & n4845 ) | ( n3301 & n4845 ) ;
  assign n4847 = ( n3610 & ~n3614 ) | ( n3610 & n4846 ) | ( ~n3614 & n4846 ) ;
  assign n4848 = ( n3900 & ~n3904 ) | ( n3900 & n4847 ) | ( ~n3904 & n4847 ) ;
  assign n4849 = ( n4177 & ~n4245 ) | ( n4177 & n4848 ) | ( ~n4245 & n4848 ) ;
  assign n4850 = ( n4501 & ~n4562 ) | ( n4501 & n4849 ) | ( ~n4562 & n4849 ) ;
  assign n4851 = n549 | n2240 ;
  assign n4852 = ~n544 & n1918 ;
  assign n4853 = ( ~n549 & n1545 ) | ( ~n549 & n4852 ) | ( n1545 & n4852 ) ;
  assign n4854 = ( n4850 & n4851 ) | ( n4850 & ~n4853 ) | ( n4851 & ~n4853 ) ;
  assign n4855 = ( ~n2253 & n2507 ) | ( ~n2253 & n4854 ) | ( n2507 & n4854 ) ;
  assign n4856 = n4838 & n4855 ;
  assign n4857 = x233 & ~n990 ;
  assign n4858 = x107 | n987 ;
  assign n4859 = ~n587 & n4858 ;
  assign n4860 = ( ~n582 & n1944 ) | ( ~n582 & n4859 ) | ( n1944 & n4859 ) ;
  assign n4861 = ( ~n1568 & n2259 ) | ( ~n1568 & n4860 ) | ( n2259 & n4860 ) ;
  assign n4862 = ( n2702 & ~n2710 ) | ( n2702 & n4861 ) | ( ~n2710 & n4861 ) ;
  assign n4863 = ( ~n1579 & n1585 ) | ( ~n1579 & n4862 ) | ( n1585 & n4862 ) ;
  assign n4864 = ( ~n2538 & n3087 ) | ( ~n2538 & n4863 ) | ( n3087 & n4863 ) ;
  assign n4865 = ( ~n2926 & n3327 ) | ( ~n2926 & n4864 ) | ( n3327 & n4864 ) ;
  assign n4866 = ( n3635 & ~n3639 ) | ( n3635 & n4865 ) | ( ~n3639 & n4865 ) ;
  assign n4867 = ( n3923 & ~n3927 ) | ( n3923 & n4866 ) | ( ~n3927 & n4866 ) ;
  assign n4868 = ( n4199 & ~n4267 ) | ( n4199 & n4867 ) | ( ~n4267 & n4867 ) ;
  assign n4869 = ( n4521 & ~n4582 ) | ( n4521 & n4868 ) | ( ~n4582 & n4868 ) ;
  assign n4870 = n947 | n2336 ;
  assign n4871 = ~n942 & n2027 ;
  assign n4872 = ( ~n947 & n1684 ) | ( ~n947 & n4871 ) | ( n1684 & n4871 ) ;
  assign n4873 = ( n4869 & n4870 ) | ( n4869 & ~n4872 ) | ( n4870 & ~n4872 ) ;
  assign n4874 = ( ~n2349 & n2576 ) | ( ~n2349 & n4873 ) | ( n2576 & n4873 ) ;
  assign n4875 = n4857 & n4874 ;
  assign n4876 = x234 & ~n1387 ;
  assign n4877 = x108 | n1384 ;
  assign n4878 = ~n985 & n4877 ;
  assign n4879 = ( ~n980 & n2053 ) | ( ~n980 & n4878 ) | ( n2053 & n4878 ) ;
  assign n4880 = ( ~n1707 & n2355 ) | ( ~n1707 & n4879 ) | ( n2355 & n4879 ) ;
  assign n4881 = ( n2746 & ~n2754 ) | ( n2746 & n4880 ) | ( ~n2754 & n4880 ) ;
  assign n4882 = ( ~n1718 & n1724 ) | ( ~n1718 & n4881 ) | ( n1724 & n4881 ) ;
  assign n4883 = ( ~n2607 & n3114 ) | ( ~n2607 & n4882 ) | ( n3114 & n4882 ) ;
  assign n4884 = ( ~n2955 & n3353 ) | ( ~n2955 & n4883 ) | ( n3353 & n4883 ) ;
  assign n4885 = ( n3660 & ~n3664 ) | ( n3660 & n4884 ) | ( ~n3664 & n4884 ) ;
  assign n4886 = ( n3946 & ~n3950 ) | ( n3946 & n4885 ) | ( ~n3950 & n4885 ) ;
  assign n4887 = ( n4221 & ~n4289 ) | ( n4221 & n4886 ) | ( ~n4289 & n4886 ) ;
  assign n4888 = ( n4541 & ~n4602 ) | ( n4541 & n4887 ) | ( ~n4602 & n4887 ) ;
  assign n4889 = n1344 | n2432 ;
  assign n4890 = ~n1339 & n2136 ;
  assign n4891 = ( ~n1344 & n1822 ) | ( ~n1344 & n4890 ) | ( n1822 & n4890 ) ;
  assign n4892 = ( n4888 & n4889 ) | ( n4888 & ~n4891 ) | ( n4889 & ~n4891 ) ;
  assign n4893 = ( ~n2445 & n2645 ) | ( ~n2445 & n4892 ) | ( n2645 & n4892 ) ;
  assign n4894 = n4876 & n4893 ;
  assign n4895 = x235 & ~n586 ;
  assign n4896 = x109 | n583 ;
  assign n4897 = ~n1382 & n4896 ;
  assign n4898 = ( ~n1377 & n2162 ) | ( ~n1377 & n4897 ) | ( n2162 & n4897 ) ;
  assign n4899 = ( ~n1845 & n2451 ) | ( ~n1845 & n4898 ) | ( n2451 & n4898 ) ;
  assign n4900 = ( n2790 & ~n2798 ) | ( n2790 & n4899 ) | ( ~n2798 & n4899 ) ;
  assign n4901 = ( ~n1855 & n1859 ) | ( ~n1855 & n4900 ) | ( n1859 & n4900 ) ;
  assign n4902 = ( ~n2675 & n3141 ) | ( ~n2675 & n4901 ) | ( n3141 & n4901 ) ;
  assign n4903 = ( ~n2984 & n3379 ) | ( ~n2984 & n4902 ) | ( n3379 & n4902 ) ;
  assign n4904 = ( n3684 & ~n3688 ) | ( n3684 & n4903 ) | ( ~n3688 & n4903 ) ;
  assign n4905 = ( n3969 & ~n3973 ) | ( n3969 & n4904 ) | ( ~n3973 & n4904 ) ;
  assign n4906 = ( n4243 & ~n4311 ) | ( n4243 & n4905 ) | ( ~n4311 & n4905 ) ;
  assign n4907 = ( n4561 & ~n4622 ) | ( n4561 & n4906 ) | ( ~n4622 & n4906 ) ;
  assign n4908 = n554 | n2503 ;
  assign n4909 = ~n549 & n2232 ;
  assign n4910 = ( ~n554 & n563 ) | ( ~n554 & n4909 ) | ( n563 & n4909 ) ;
  assign n4911 = ( n4907 & n4908 ) | ( n4907 & ~n4910 ) | ( n4908 & ~n4910 ) ;
  assign n4912 = ( ~n2515 & n2695 ) | ( ~n2515 & n4911 ) | ( n2695 & n4911 ) ;
  assign n4913 = n4895 & n4912 ;
  assign n4914 = x236 & ~n984 ;
  assign n4915 = x110 | n981 ;
  assign n4916 = ~n581 & n4915 ;
  assign n4917 = ( ~n576 & n2258 ) | ( ~n576 & n4916 ) | ( n2258 & n4916 ) ;
  assign n4918 = ( ~n623 & n2520 ) | ( ~n623 & n4917 ) | ( n2520 & n4917 ) ;
  assign n4919 = ( ~n643 & n650 ) | ( ~n643 & n4918 ) | ( n650 & n4918 ) ;
  assign n4920 = ( ~n1964 & n1968 ) | ( ~n1964 & n4919 ) | ( n1968 & n4919 ) ;
  assign n4921 = ( ~n2719 & n3168 ) | ( ~n2719 & n4920 ) | ( n3168 & n4920 ) ;
  assign n4922 = ( ~n3013 & n3405 ) | ( ~n3013 & n4921 ) | ( n3405 & n4921 ) ;
  assign n4923 = ( n3708 & ~n3712 ) | ( n3708 & n4922 ) | ( ~n3712 & n4922 ) ;
  assign n4924 = ( n3992 & ~n3996 ) | ( n3992 & n4923 ) | ( ~n3996 & n4923 ) ;
  assign n4925 = ( n4265 & ~n4333 ) | ( n4265 & n4924 ) | ( ~n4333 & n4924 ) ;
  assign n4926 = ( n4581 & ~n4642 ) | ( n4581 & n4925 ) | ( ~n4642 & n4925 ) ;
  assign n4927 = n952 | n2572 ;
  assign n4928 = ~n947 & n2328 ;
  assign n4929 = ( ~n952 & n961 ) | ( ~n952 & n4928 ) | ( n961 & n4928 ) ;
  assign n4930 = ( n4926 & n4927 ) | ( n4926 & ~n4929 ) | ( n4927 & ~n4929 ) ;
  assign n4931 = ( ~n2584 & n2739 ) | ( ~n2584 & n4930 ) | ( n2739 & n4930 ) ;
  assign n4932 = n4914 & n4931 ;
  assign n4933 = x237 & ~n1381 ;
  assign n4934 = x111 | n1378 ;
  assign n4935 = ~n979 & n4934 ;
  assign n4936 = ( ~n974 & n2354 ) | ( ~n974 & n4935 ) | ( n2354 & n4935 ) ;
  assign n4937 = ( ~n1021 & n2589 ) | ( ~n1021 & n4936 ) | ( n2589 & n4936 ) ;
  assign n4938 = ( ~n1041 & n1048 ) | ( ~n1041 & n4937 ) | ( n1048 & n4937 ) ;
  assign n4939 = ( ~n2073 & n2077 ) | ( ~n2073 & n4938 ) | ( n2077 & n4938 ) ;
  assign n4940 = ( ~n2763 & n3195 ) | ( ~n2763 & n4939 ) | ( n3195 & n4939 ) ;
  assign n4941 = ( ~n3042 & n3431 ) | ( ~n3042 & n4940 ) | ( n3431 & n4940 ) ;
  assign n4942 = ( n3732 & ~n3736 ) | ( n3732 & n4941 ) | ( ~n3736 & n4941 ) ;
  assign n4943 = ( n4015 & ~n4019 ) | ( n4015 & n4942 ) | ( ~n4019 & n4942 ) ;
  assign n4944 = ( n4287 & ~n4355 ) | ( n4287 & n4943 ) | ( ~n4355 & n4943 ) ;
  assign n4945 = ( n4601 & ~n4662 ) | ( n4601 & n4944 ) | ( ~n4662 & n4944 ) ;
  assign n4946 = n1349 | n2641 ;
  assign n4947 = ~n1344 & n2424 ;
  assign n4948 = ( ~n1349 & n1358 ) | ( ~n1349 & n4947 ) | ( n1358 & n4947 ) ;
  assign n4949 = ( n4945 & n4946 ) | ( n4945 & ~n4948 ) | ( n4946 & ~n4948 ) ;
  assign n4950 = ( ~n2653 & n2783 ) | ( ~n2653 & n4949 ) | ( n2783 & n4949 ) ;
  assign n4951 = n4933 & n4950 ;
  assign n4952 = x238 & ~n580 ;
  assign n4953 = x112 | n577 ;
  assign n4954 = ~n1376 & n4953 ;
  assign n4955 = ( ~n1371 & n2450 ) | ( ~n1371 & n4954 ) | ( n2450 & n4954 ) ;
  assign n4956 = ( ~n1418 & n2658 ) | ( ~n1418 & n4955 ) | ( n2658 & n4955 ) ;
  assign n4957 = ( ~n1438 & n1445 ) | ( ~n1438 & n4956 ) | ( n1445 & n4956 ) ;
  assign n4958 = ( ~n2181 & n2185 ) | ( ~n2181 & n4957 ) | ( n2185 & n4957 ) ;
  assign n4959 = ( ~n2807 & n3222 ) | ( ~n2807 & n4958 ) | ( n3222 & n4958 ) ;
  assign n4960 = ( ~n3070 & n3457 ) | ( ~n3070 & n4959 ) | ( n3457 & n4959 ) ;
  assign n4961 = ( n3756 & ~n3760 ) | ( n3756 & n4960 ) | ( ~n3760 & n4960 ) ;
  assign n4962 = ( n4038 & ~n4042 ) | ( n4038 & n4961 ) | ( ~n4042 & n4961 ) ;
  assign n4963 = ( n4309 & ~n4377 ) | ( n4309 & n4962 ) | ( ~n4377 & n4962 ) ;
  assign n4964 = ( n4621 & ~n4681 ) | ( n4621 & n4963 ) | ( ~n4681 & n4963 ) ;
  assign n4965 = ~n554 & n2496 ;
  assign n4966 = ( ~n517 & n1549 ) | ( ~n517 & n4965 ) | ( n1549 & n4965 ) ;
  assign n4967 = ( n557 & n4964 ) | ( n557 & ~n4966 ) | ( n4964 & ~n4966 ) ;
  assign n4968 = ( n601 & ~n618 ) | ( n601 & n4967 ) | ( ~n618 & n4967 ) ;
  assign n4969 = n4952 & n4968 ;
  assign n4970 = x239 & ~n978 ;
  assign n4971 = x113 | n975 ;
  assign n4972 = ~n575 & n4971 ;
  assign n4973 = ( ~n573 & n608 ) | ( ~n573 & n4972 ) | ( n608 & n4972 ) ;
  assign n4974 = ( ~n638 & n2702 ) | ( ~n638 & n4973 ) | ( n2702 & n4973 ) ;
  assign n4975 = ( ~n1578 & n1584 ) | ( ~n1578 & n4974 ) | ( n1584 & n4974 ) ;
  assign n4976 = ( ~n2277 & n2281 ) | ( ~n2277 & n4975 ) | ( n2281 & n4975 ) ;
  assign n4977 = ( ~n2837 & n3248 ) | ( ~n2837 & n4976 ) | ( n3248 & n4976 ) ;
  assign n4978 = ( ~n3097 & n3483 ) | ( ~n3097 & n4977 ) | ( n3483 & n4977 ) ;
  assign n4979 = ( n3780 & ~n3784 ) | ( n3780 & n4978 ) | ( ~n3784 & n4978 ) ;
  assign n4980 = ( n4061 & ~n4065 ) | ( n4061 & n4979 ) | ( ~n4065 & n4979 ) ;
  assign n4981 = ( n4331 & ~n4399 ) | ( n4331 & n4980 ) | ( ~n4399 & n4980 ) ;
  assign n4982 = ( n4641 & ~n4700 ) | ( n4641 & n4981 ) | ( ~n4700 & n4981 ) ;
  assign n4983 = ~n952 & n2565 ;
  assign n4984 = ( ~n915 & n1688 ) | ( ~n915 & n4983 ) | ( n1688 & n4983 ) ;
  assign n4985 = ( n955 & n4982 ) | ( n955 & ~n4984 ) | ( n4982 & ~n4984 ) ;
  assign n4986 = ( n999 & ~n1016 ) | ( n999 & n4985 ) | ( ~n1016 & n4985 ) ;
  assign n4987 = n4970 & n4986 ;
  assign n4988 = x240 & ~n1375 ;
  assign n4989 = x114 | n1372 ;
  assign n4990 = ~n973 & n4989 ;
  assign n4991 = ( ~n971 & n1006 ) | ( ~n971 & n4990 ) | ( n1006 & n4990 ) ;
  assign n4992 = ( ~n1036 & n2746 ) | ( ~n1036 & n4991 ) | ( n2746 & n4991 ) ;
  assign n4993 = ( ~n1717 & n1723 ) | ( ~n1717 & n4992 ) | ( n1723 & n4992 ) ;
  assign n4994 = ( ~n2373 & n2377 ) | ( ~n2373 & n4993 ) | ( n2377 & n4993 ) ;
  assign n4995 = ( ~n2867 & n3274 ) | ( ~n2867 & n4994 ) | ( n3274 & n4994 ) ;
  assign n4996 = ( ~n3124 & n3509 ) | ( ~n3124 & n4995 ) | ( n3509 & n4995 ) ;
  assign n4997 = ( n3804 & ~n3808 ) | ( n3804 & n4996 ) | ( ~n3808 & n4996 ) ;
  assign n4998 = ( n4084 & ~n4088 ) | ( n4084 & n4997 ) | ( ~n4088 & n4997 ) ;
  assign n4999 = ( n4353 & ~n4421 ) | ( n4353 & n4998 ) | ( ~n4421 & n4998 ) ;
  assign n5000 = ( n4661 & ~n4719 ) | ( n4661 & n4999 ) | ( ~n4719 & n4999 ) ;
  assign n5001 = ~n1349 & n2634 ;
  assign n5002 = ( ~n1312 & n1826 ) | ( ~n1312 & n5001 ) | ( n1826 & n5001 ) ;
  assign n5003 = ( n1352 & n5000 ) | ( n1352 & ~n5002 ) | ( n5000 & ~n5002 ) ;
  assign n5004 = ( n1396 & ~n1413 ) | ( n1396 & n5003 ) | ( ~n1413 & n5003 ) ;
  assign n5005 = n4988 & n5004 ;
  assign n5006 = x241 & ~n574 ;
  assign n5007 = x115 | n605 ;
  assign n5008 = ~n1370 & n5007 ;
  assign n5009 = ( ~n1368 & n1403 ) | ( ~n1368 & n5008 ) | ( n1403 & n5008 ) ;
  assign n5010 = ( ~n1433 & n2790 ) | ( ~n1433 & n5009 ) | ( n2790 & n5009 ) ;
  assign n5011 = ( ~n1854 & n1858 ) | ( ~n1854 & n5010 ) | ( n1858 & n5010 ) ;
  assign n5012 = ( ~n2469 & n2472 ) | ( ~n2469 & n5011 ) | ( n2472 & n5011 ) ;
  assign n5013 = ( ~n2896 & n3300 ) | ( ~n2896 & n5012 ) | ( n3300 & n5012 ) ;
  assign n5014 = ( ~n3151 & n3535 ) | ( ~n3151 & n5013 ) | ( n3535 & n5013 ) ;
  assign n5015 = ( n3828 & ~n3832 ) | ( n3828 & n5014 ) | ( ~n3832 & n5014 ) ;
  assign n5016 = ( n4107 & ~n4111 ) | ( n4107 & n5015 ) | ( ~n4111 & n5015 ) ;
  assign n5017 = ( ~n458 & n4375 ) | ( ~n458 & n5016 ) | ( n4375 & n5016 ) ;
  assign n5018 = ( n4680 & ~n4738 ) | ( n4680 & n5017 ) | ( ~n4738 & n5017 ) ;
  assign n5019 = ( n566 & ~n597 ) | ( n566 & n614 ) | ( ~n597 & n614 ) ;
  assign n5020 = ( n1544 & n5018 ) | ( n1544 & ~n5019 ) | ( n5018 & ~n5019 ) ;
  assign n5021 = ( n1557 & ~n1567 ) | ( n1557 & n5020 ) | ( ~n1567 & n5020 ) ;
  assign n5022 = n5006 & n5021 ;
  assign n5023 = x242 & ~n972 ;
  assign n5024 = x116 | n1003 ;
  assign n5025 = ~n572 & n5024 ;
  assign n5026 = ( ~n634 & n1561 ) | ( ~n634 & n5025 ) | ( n1561 & n5025 ) ;
  assign n5027 = ( n650 & ~n1576 ) | ( n650 & n5026 ) | ( ~n1576 & n5026 ) ;
  assign n5028 = ( ~n1963 & n1967 ) | ( ~n1963 & n5027 ) | ( n1967 & n5027 ) ;
  assign n5029 = ( ~n2538 & n2541 ) | ( ~n2538 & n5028 ) | ( n2541 & n5028 ) ;
  assign n5030 = ( ~n2925 & n3326 ) | ( ~n2925 & n5029 ) | ( n3326 & n5029 ) ;
  assign n5031 = ( ~n3178 & n3560 ) | ( ~n3178 & n5030 ) | ( n3560 & n5030 ) ;
  assign n5032 = ( n3852 & ~n3856 ) | ( n3852 & n5031 ) | ( ~n3856 & n5031 ) ;
  assign n5033 = ( n4130 & ~n4134 ) | ( n4130 & n5032 ) | ( ~n4134 & n5032 ) ;
  assign n5034 = ( ~n856 & n4397 ) | ( ~n856 & n5033 ) | ( n4397 & n5033 ) ;
  assign n5035 = ( n4699 & ~n4757 ) | ( n4699 & n5034 ) | ( ~n4757 & n5034 ) ;
  assign n5036 = ( n964 & ~n995 ) | ( n964 & n1012 ) | ( ~n995 & n1012 ) ;
  assign n5037 = ( n1683 & n5035 ) | ( n1683 & ~n5036 ) | ( n5035 & ~n5036 ) ;
  assign n5038 = ( n1696 & ~n1706 ) | ( n1696 & n5037 ) | ( ~n1706 & n5037 ) ;
  assign n5039 = n5023 & n5038 ;
  assign n5040 = x243 & ~n1369 ;
  assign n5041 = x117 | n1400 ;
  assign n5042 = ~n970 & n5041 ;
  assign n5043 = ( ~n1032 & n1700 ) | ( ~n1032 & n5042 ) | ( n1700 & n5042 ) ;
  assign n5044 = ( n1048 & ~n1715 ) | ( n1048 & n5043 ) | ( ~n1715 & n5043 ) ;
  assign n5045 = ( ~n2072 & n2076 ) | ( ~n2072 & n5044 ) | ( n2076 & n5044 ) ;
  assign n5046 = ( ~n2607 & n2610 ) | ( ~n2607 & n5045 ) | ( n2610 & n5045 ) ;
  assign n5047 = ( ~n2954 & n3352 ) | ( ~n2954 & n5046 ) | ( n3352 & n5046 ) ;
  assign n5048 = ( ~n3205 & n3585 ) | ( ~n3205 & n5047 ) | ( n3585 & n5047 ) ;
  assign n5049 = ( n3876 & ~n3880 ) | ( n3876 & n5048 ) | ( ~n3880 & n5048 ) ;
  assign n5050 = ( n4153 & ~n4157 ) | ( n4153 & n5049 ) | ( ~n4157 & n5049 ) ;
  assign n5051 = ( ~n1253 & n4419 ) | ( ~n1253 & n5050 ) | ( n4419 & n5050 ) ;
  assign n5052 = ( n4718 & ~n4776 ) | ( n4718 & n5051 ) | ( ~n4776 & n5051 ) ;
  assign n5053 = ( n1361 & ~n1392 ) | ( n1361 & n1409 ) | ( ~n1392 & n1409 ) ;
  assign n5054 = ( n1821 & n5052 ) | ( n1821 & ~n5053 ) | ( n5052 & ~n5053 ) ;
  assign n5055 = ( n1834 & ~n1844 ) | ( n1834 & n5054 ) | ( ~n1844 & n5054 ) ;
  assign n5056 = n5040 & n5055 ;
  assign n5057 = x244 & ~n571 ;
  assign n5058 = x118 | n568 ;
  assign n5059 = ~n1367 & n5058 ;
  assign n5060 = ( ~n1429 & n1838 ) | ( ~n1429 & n5059 ) | ( n1838 & n5059 ) ;
  assign n5061 = ( n1445 & ~n1852 ) | ( n1445 & n5060 ) | ( ~n1852 & n5060 ) ;
  assign n5062 = ( ~n2180 & n2184 ) | ( ~n2180 & n5061 ) | ( n2184 & n5061 ) ;
  assign n5063 = ( ~n2675 & n2677 ) | ( ~n2675 & n5062 ) | ( n2677 & n5062 ) ;
  assign n5064 = ( ~n2983 & n3378 ) | ( ~n2983 & n5063 ) | ( n3378 & n5063 ) ;
  assign n5065 = ( ~n3232 & n3610 ) | ( ~n3232 & n5064 ) | ( n3610 & n5064 ) ;
  assign n5066 = ( n379 & ~n3903 ) | ( n379 & n5065 ) | ( ~n3903 & n5065 ) ;
  assign n5067 = ( n4176 & ~n4179 ) | ( n4176 & n5066 ) | ( ~n4179 & n5066 ) ;
  assign n5068 = ( ~n1510 & n4440 ) | ( ~n1510 & n5067 ) | ( n4440 & n5067 ) ;
  assign n5069 = ( n4737 & ~n4795 ) | ( n4737 & n5068 ) | ( ~n4795 & n5068 ) ;
  assign n5070 = ( ~n591 & n615 ) | ( ~n591 & n1552 ) | ( n615 & n1552 ) ;
  assign n5071 = ( n1936 & n5069 ) | ( n1936 & ~n5070 ) | ( n5069 & ~n5070 ) ;
  assign n5072 = ( n1947 & ~n1955 ) | ( n1947 & n5071 ) | ( ~n1955 & n5071 ) ;
  assign n5073 = n5057 & n5072 ;
  assign n5074 = x245 & ~n969 ;
  assign n5075 = x119 | n966 ;
  assign n5076 = ~n633 & n5075 ;
  assign n5077 = ( ~n631 & n649 ) | ( ~n631 & n5076 ) | ( n649 & n5076 ) ;
  assign n5078 = ( ~n1577 & n1584 ) | ( ~n1577 & n5077 ) | ( n1584 & n5077 ) ;
  assign n5079 = ( ~n2276 & n2280 ) | ( ~n2276 & n5078 ) | ( n2280 & n5078 ) ;
  assign n5080 = ( ~n2719 & n2721 ) | ( ~n2719 & n5079 ) | ( n2721 & n5079 ) ;
  assign n5081 = ( ~n3012 & n3404 ) | ( ~n3012 & n5080 ) | ( n3404 & n5080 ) ;
  assign n5082 = ( ~n3258 & n3635 ) | ( ~n3258 & n5081 ) | ( n3635 & n5081 ) ;
  assign n5083 = ( n777 & ~n3926 ) | ( n777 & n5082 ) | ( ~n3926 & n5082 ) ;
  assign n5084 = ( n4198 & ~n4201 ) | ( n4198 & n5083 ) | ( ~n4201 & n5083 ) ;
  assign n5085 = ( ~n1649 & n4460 ) | ( ~n1649 & n5084 ) | ( n4460 & n5084 ) ;
  assign n5086 = ( n4756 & ~n4814 ) | ( n4756 & n5085 ) | ( ~n4814 & n5085 ) ;
  assign n5087 = ( ~n989 & n1013 ) | ( ~n989 & n1691 ) | ( n1013 & n1691 ) ;
  assign n5088 = ( n2045 & n5086 ) | ( n2045 & ~n5087 ) | ( n5086 & ~n5087 ) ;
  assign n5089 = ( n2056 & ~n2064 ) | ( n2056 & n5088 ) | ( ~n2064 & n5088 ) ;
  assign n5090 = n5074 & n5089 ;
  assign n5091 = x246 & ~n1366 ;
  assign n5092 = x120 | n1363 ;
  assign n5093 = ~n1031 & n5092 ;
  assign n5094 = ( ~n1029 & n1047 ) | ( ~n1029 & n5093 ) | ( n1047 & n5093 ) ;
  assign n5095 = ( ~n1716 & n1723 ) | ( ~n1716 & n5094 ) | ( n1723 & n5094 ) ;
  assign n5096 = ( ~n2372 & n2376 ) | ( ~n2372 & n5095 ) | ( n2376 & n5095 ) ;
  assign n5097 = ( ~n2763 & n2765 ) | ( ~n2763 & n5096 ) | ( n2765 & n5096 ) ;
  assign n5098 = ( ~n3041 & n3430 ) | ( ~n3041 & n5097 ) | ( n3430 & n5097 ) ;
  assign n5099 = ( ~n3284 & n3660 ) | ( ~n3284 & n5098 ) | ( n3660 & n5098 ) ;
  assign n5100 = ( n1174 & ~n3949 ) | ( n1174 & n5099 ) | ( ~n3949 & n5099 ) ;
  assign n5101 = ( n4220 & ~n4223 ) | ( n4220 & n5100 ) | ( ~n4223 & n5100 ) ;
  assign n5102 = ( ~n1787 & n4480 ) | ( ~n1787 & n5101 ) | ( n4480 & n5101 ) ;
  assign n5103 = ( n4775 & ~n4833 ) | ( n4775 & n5102 ) | ( ~n4833 & n5102 ) ;
  assign n5104 = ( ~n1386 & n1410 ) | ( ~n1386 & n1829 ) | ( n1410 & n1829 ) ;
  assign n5105 = ( n2154 & n5103 ) | ( n2154 & ~n5104 ) | ( n5103 & ~n5104 ) ;
  assign n5106 = ( n2165 & ~n2173 ) | ( n2165 & n5105 ) | ( ~n2173 & n5105 ) ;
  assign n5107 = n5091 & n5106 ;
  assign n5108 = x247 & ~n632 ;
  assign n5109 = x121 | n635 ;
  assign n5110 = ~n1428 & n5109 ;
  assign n5111 = ( ~n1426 & n1444 ) | ( ~n1426 & n5110 ) | ( n1444 & n5110 ) ;
  assign n5112 = ( ~n1853 & n1858 ) | ( ~n1853 & n5111 ) | ( n1858 & n5111 ) ;
  assign n5113 = ( ~n2468 & n2471 ) | ( ~n2468 & n5112 ) | ( n2471 & n5112 ) ;
  assign n5114 = ( ~n2807 & n2809 ) | ( ~n2807 & n5113 ) | ( n2809 & n5113 ) ;
  assign n5115 = ( ~n320 & n3456 ) | ( ~n320 & n5114 ) | ( n3456 & n5114 ) ;
  assign n5116 = ( ~n3310 & n3684 ) | ( ~n3310 & n5115 ) | ( n3684 & n5115 ) ;
  assign n5117 = ( n1485 & ~n3972 ) | ( n1485 & n5116 ) | ( ~n3972 & n5116 ) ;
  assign n5118 = ( n4242 & ~n4245 ) | ( n4242 & n5117 ) | ( ~n4245 & n5117 ) ;
  assign n5119 = ( ~n1905 & n4500 ) | ( ~n1905 & n5118 ) | ( n4500 & n5118 ) ;
  assign n5120 = ( n4794 & ~n4852 ) | ( n4794 & n5119 ) | ( ~n4852 & n5119 ) ;
  assign n5121 = ( ~n585 & n1564 ) | ( ~n585 & n1942 ) | ( n1564 & n1942 ) ;
  assign n5122 = ( n2250 & n5120 ) | ( n2250 & ~n5121 ) | ( n5120 & ~n5121 ) ;
  assign n5123 = ( n2261 & ~n2269 ) | ( n2261 & n5122 ) | ( ~n2269 & n5122 ) ;
  assign n5124 = n5108 & n5123 ;
  assign n5125 = x248 & ~n1030 ;
  assign n5126 = x122 | n1033 ;
  assign n5127 = ~n630 & n5126 ;
  assign n5128 = ( ~n628 & n1583 ) | ( ~n628 & n5127 ) | ( n1583 & n5127 ) ;
  assign n5129 = ( ~n1962 & n1967 ) | ( ~n1962 & n5128 ) | ( n1967 & n5128 ) ;
  assign n5130 = ( ~n2537 & n2540 ) | ( ~n2537 & n5129 ) | ( n2540 & n5129 ) ;
  assign n5131 = ( ~n2837 & n2839 ) | ( ~n2837 & n5130 ) | ( n2839 & n5130 ) ;
  assign n5132 = ( ~n718 & n3482 ) | ( ~n718 & n5131 ) | ( n3482 & n5131 ) ;
  assign n5133 = ( ~n3336 & n3708 ) | ( ~n3336 & n5132 ) | ( n3708 & n5132 ) ;
  assign n5134 = ( n1624 & ~n3995 ) | ( n1624 & n5133 ) | ( ~n3995 & n5133 ) ;
  assign n5135 = ( n4264 & ~n4267 ) | ( n4264 & n5134 ) | ( ~n4267 & n5134 ) ;
  assign n5136 = ( ~n2014 & n4520 ) | ( ~n2014 & n5135 ) | ( n4520 & n5135 ) ;
  assign n5137 = ( n4813 & ~n4871 ) | ( n4813 & n5136 ) | ( ~n4871 & n5136 ) ;
  assign n5138 = ( ~n983 & n1703 ) | ( ~n983 & n2051 ) | ( n1703 & n2051 ) ;
  assign n5139 = ( n2346 & n5137 ) | ( n2346 & ~n5138 ) | ( n5137 & ~n5138 ) ;
  assign n5140 = ( n2357 & ~n2365 ) | ( n2357 & n5139 ) | ( ~n2365 & n5139 ) ;
  assign n5141 = n5125 & n5140 ;
  assign n5142 = x249 & ~n1427 ;
  assign n5143 = x123 | n1430 ;
  assign n5144 = ~n1028 & n5143 ;
  assign n5145 = ( ~n1026 & n1722 ) | ( ~n1026 & n5144 ) | ( n1722 & n5144 ) ;
  assign n5146 = ( ~n2071 & n2076 ) | ( ~n2071 & n5145 ) | ( n2076 & n5145 ) ;
  assign n5147 = ( ~n2606 & n2609 ) | ( ~n2606 & n5146 ) | ( n2609 & n5146 ) ;
  assign n5148 = ( ~n2867 & n2869 ) | ( ~n2867 & n5147 ) | ( n2869 & n5147 ) ;
  assign n5149 = ( ~n1115 & n3508 ) | ( ~n1115 & n5148 ) | ( n3508 & n5148 ) ;
  assign n5150 = ( ~n3362 & n3732 ) | ( ~n3362 & n5149 ) | ( n3732 & n5149 ) ;
  assign n5151 = ( n1762 & ~n4018 ) | ( n1762 & n5150 ) | ( ~n4018 & n5150 ) ;
  assign n5152 = ( n4286 & ~n4289 ) | ( n4286 & n5151 ) | ( ~n4289 & n5151 ) ;
  assign n5153 = ( ~n2123 & n4540 ) | ( ~n2123 & n5152 ) | ( n4540 & n5152 ) ;
  assign n5154 = ( n4832 & ~n4890 ) | ( n4832 & n5153 ) | ( ~n4890 & n5153 ) ;
  assign n5155 = ( ~n1380 & n1841 ) | ( ~n1380 & n2160 ) | ( n1841 & n2160 ) ;
  assign n5156 = ( n2442 & n5154 ) | ( n2442 & ~n5155 ) | ( n5154 & ~n5155 ) ;
  assign n5157 = ( n2453 & ~n2461 ) | ( n2453 & n5156 ) | ( ~n2461 & n5156 ) ;
  assign n5158 = n5142 & n5157 ;
  assign n5159 = x250 & ~n629 ;
  assign n5160 = x124 | n640 ;
  assign n5161 = ~n1425 & n5160 ;
  assign n5162 = ( ~n1423 & n1857 ) | ( ~n1423 & n5161 ) | ( n1857 & n5161 ) ;
  assign n5163 = ( ~n2179 & n2184 ) | ( ~n2179 & n5162 ) | ( n2184 & n5162 ) ;
  assign n5164 = ( n281 & ~n2674 ) | ( n281 & n5163 ) | ( ~n2674 & n5163 ) ;
  assign n5165 = ( ~n2896 & n2898 ) | ( ~n2896 & n5164 ) | ( n2898 & n5164 ) ;
  assign n5166 = ( ~n1466 & n3534 ) | ( ~n1466 & n5165 ) | ( n3534 & n5165 ) ;
  assign n5167 = ( ~n3388 & n3756 ) | ( ~n3388 & n5166 ) | ( n3756 & n5166 ) ;
  assign n5168 = ( n1885 & ~n4041 ) | ( n1885 & n5167 ) | ( ~n4041 & n5167 ) ;
  assign n5169 = ( n4308 & ~n4311 ) | ( n4308 & n5168 ) | ( ~n4311 & n5168 ) ;
  assign n5170 = ( ~n2219 & n4560 ) | ( ~n2219 & n5169 ) | ( n4560 & n5169 ) ;
  assign n5171 = ( n4851 & ~n4909 ) | ( n4851 & n5170 ) | ( ~n4909 & n5170 ) ;
  assign n5172 = ( ~n579 & n619 ) | ( ~n579 & n2256 ) | ( n619 & n2256 ) ;
  assign n5173 = ( n2512 & n5171 ) | ( n2512 & ~n5172 ) | ( n5171 & ~n5172 ) ;
  assign n5174 = ( n2522 & ~n2530 ) | ( n2522 & n5173 ) | ( ~n2530 & n5173 ) ;
  assign n5175 = n5159 & n5174 ;
  assign n5176 = x251 & ~n1027 ;
  assign n5177 = x125 | n1038 ;
  assign n5178 = ~n627 & n5177 ;
  assign n5179 = ( ~n1575 & n1966 ) | ( ~n1575 & n5178 ) | ( n1966 & n5178 ) ;
  assign n5180 = ( ~n2275 & n2280 ) | ( ~n2275 & n5179 ) | ( n2280 & n5179 ) ;
  assign n5181 = ( n679 & ~n2718 ) | ( n679 & n5180 ) | ( ~n2718 & n5180 ) ;
  assign n5182 = ( ~n2925 & n2927 ) | ( ~n2925 & n5181 ) | ( n2927 & n5181 ) ;
  assign n5183 = ( ~n1605 & n3559 ) | ( ~n1605 & n5182 ) | ( n3559 & n5182 ) ;
  assign n5184 = ( ~n3414 & n3780 ) | ( ~n3414 & n5183 ) | ( n3780 & n5183 ) ;
  assign n5185 = ( n1994 & ~n4064 ) | ( n1994 & n5184 ) | ( ~n4064 & n5184 ) ;
  assign n5186 = ( n4330 & ~n4333 ) | ( n4330 & n5185 ) | ( ~n4333 & n5185 ) ;
  assign n5187 = ( ~n2315 & n4580 ) | ( ~n2315 & n5186 ) | ( n4580 & n5186 ) ;
  assign n5188 = ( n4870 & ~n4928 ) | ( n4870 & n5187 ) | ( ~n4928 & n5187 ) ;
  assign n5189 = ( ~n977 & n1017 ) | ( ~n977 & n2352 ) | ( n1017 & n2352 ) ;
  assign n5190 = ( n2581 & n5188 ) | ( n2581 & ~n5189 ) | ( n5188 & ~n5189 ) ;
  assign n5191 = ( n2591 & ~n2599 ) | ( n2591 & n5190 ) | ( ~n2599 & n5190 ) ;
  assign n5192 = n5176 & n5191 ;
  assign n5193 = x252 & ~n1424 ;
  assign n5194 = x126 | n1435 ;
  assign n5195 = ~n1025 & n5194 ;
  assign n5196 = ( ~n1714 & n2075 ) | ( ~n1714 & n5195 ) | ( n2075 & n5195 ) ;
  assign n5197 = ( ~n2371 & n2376 ) | ( ~n2371 & n5196 ) | ( n2376 & n5196 ) ;
  assign n5198 = ( n1076 & ~n2762 ) | ( n1076 & n5197 ) | ( ~n2762 & n5197 ) ;
  assign n5199 = ( ~n2954 & n2956 ) | ( ~n2954 & n5198 ) | ( n2956 & n5198 ) ;
  assign n5200 = ( ~n1743 & n3584 ) | ( ~n1743 & n5199 ) | ( n3584 & n5199 ) ;
  assign n5201 = ( ~n3440 & n3804 ) | ( ~n3440 & n5200 ) | ( n3804 & n5200 ) ;
  assign n5202 = ( n2103 & ~n4087 ) | ( n2103 & n5201 ) | ( ~n4087 & n5201 ) ;
  assign n5203 = ( n4352 & ~n4355 ) | ( n4352 & n5202 ) | ( ~n4355 & n5202 ) ;
  assign n5204 = ( ~n2411 & n4600 ) | ( ~n2411 & n5203 ) | ( n4600 & n5203 ) ;
  assign n5205 = ( n4889 & ~n4947 ) | ( n4889 & n5204 ) | ( ~n4947 & n5204 ) ;
  assign n5206 = ( ~n1374 & n1414 ) | ( ~n1374 & n2448 ) | ( n1414 & n2448 ) ;
  assign n5207 = ( n2650 & n5205 ) | ( n2650 & ~n5206 ) | ( n5205 & ~n5206 ) ;
  assign n5208 = ( n2660 & ~n2668 ) | ( n2660 & n5207 ) | ( ~n2668 & n5207 ) ;
  assign n5209 = n5193 & n5208 ;
  assign n5210 = x253 & ~n626 ;
  assign n5211 = n646 & ~n1422 ;
  assign n5212 = ( ~n1851 & n2183 ) | ( ~n1851 & n5211 ) | ( n2183 & n5211 ) ;
  assign n5213 = ( ~n2467 & n2471 ) | ( ~n2467 & n5212 ) | ( n2471 & n5212 ) ;
  assign n5214 = ( n1456 & ~n2806 ) | ( n1456 & n5213 ) | ( ~n2806 & n5213 ) ;
  assign n5215 = ( ~n2983 & n2985 ) | ( ~n2983 & n5214 ) | ( n2985 & n5214 ) ;
  assign n5216 = ( ~n1870 & n3609 ) | ( ~n1870 & n5215 ) | ( n3609 & n5215 ) ;
  assign n5217 = ( ~n3466 & n3828 ) | ( ~n3466 & n5216 ) | ( n3828 & n5216 ) ;
  assign n5218 = ( n2202 & ~n4110 ) | ( n2202 & n5217 ) | ( ~n4110 & n5217 ) ;
  assign n5219 = ( n4374 & ~n4377 ) | ( n4374 & n5218 ) | ( ~n4377 & n5218 ) ;
  assign n5220 = ( ~n2490 & n4620 ) | ( ~n2490 & n5219 ) | ( n4620 & n5219 ) ;
  assign n5221 = ( n4908 & ~n4965 ) | ( n4908 & n5220 ) | ( ~n4965 & n5220 ) ;
  assign n5222 = ( ~n607 & n1568 ) | ( ~n607 & n2518 ) | ( n1568 & n2518 ) ;
  assign n5223 = ( n2700 & n5221 ) | ( n2700 & ~n5222 ) | ( n5221 & ~n5222 ) ;
  assign n5224 = ( n2704 & ~n2712 ) | ( n2704 & n5223 ) | ( ~n2712 & n5223 ) ;
  assign n5225 = n5210 & n5224 ;
  assign n5226 = x254 & ~n1024 ;
  assign n5227 = x0 | n1043 ;
  assign n5228 = ~n1574 & n5227 ;
  assign n5229 = ( ~n1961 & n2279 ) | ( ~n1961 & n5228 ) | ( n2279 & n5228 ) ;
  assign n5230 = ( ~n2536 & n2540 ) | ( ~n2536 & n5229 ) | ( n2540 & n5229 ) ;
  assign n5231 = ( n1595 & ~n2836 ) | ( n1595 & n5230 ) | ( ~n2836 & n5230 ) ;
  assign n5232 = ( ~n3012 & n3014 ) | ( ~n3012 & n5231 ) | ( n3014 & n5231 ) ;
  assign n5233 = ( ~n1979 & n3634 ) | ( ~n1979 & n5232 ) | ( n3634 & n5232 ) ;
  assign n5234 = ( ~n3492 & n3852 ) | ( ~n3492 & n5233 ) | ( n3852 & n5233 ) ;
  assign n5235 = ( n2298 & ~n4133 ) | ( n2298 & n5234 ) | ( ~n4133 & n5234 ) ;
  assign n5236 = ( n4396 & ~n4399 ) | ( n4396 & n5235 ) | ( ~n4399 & n5235 ) ;
  assign n5237 = ( ~n2559 & n4640 ) | ( ~n2559 & n5236 ) | ( n4640 & n5236 ) ;
  assign n5238 = ( n4927 & ~n4983 ) | ( n4927 & n5237 ) | ( ~n4983 & n5237 ) ;
  assign n5239 = ( ~n1005 & n1707 ) | ( ~n1005 & n2587 ) | ( n1707 & n2587 ) ;
  assign n5240 = ( n2744 & n5238 ) | ( n2744 & ~n5239 ) | ( n5238 & ~n5239 ) ;
  assign n5241 = ( n2748 & ~n2756 ) | ( n2748 & n5240 ) | ( ~n2756 & n5240 ) ;
  assign n5242 = n5226 & n5241 ;
  assign n5243 = x255 & ~n1421 ;
  assign n5244 = x1 | n1440 ;
  assign n5245 = ~n1713 & n5244 ;
  assign n5246 = ( ~n2070 & n2375 ) | ( ~n2070 & n5245 ) | ( n2375 & n5245 ) ;
  assign n5247 = ( ~n2605 & n2609 ) | ( ~n2605 & n5246 ) | ( n2609 & n5246 ) ;
  assign n5248 = ( n1733 & ~n2866 ) | ( n1733 & n5247 ) | ( ~n2866 & n5247 ) ;
  assign n5249 = ( ~n3041 & n3043 ) | ( ~n3041 & n5248 ) | ( n3043 & n5248 ) ;
  assign n5250 = ( ~n2088 & n3659 ) | ( ~n2088 & n5249 ) | ( n3659 & n5249 ) ;
  assign n5251 = ( ~n3518 & n3876 ) | ( ~n3518 & n5250 ) | ( n3876 & n5250 ) ;
  assign n5252 = ( n2394 & ~n4156 ) | ( n2394 & n5251 ) | ( ~n4156 & n5251 ) ;
  assign n5253 = ( n4418 & ~n4421 ) | ( n4418 & n5252 ) | ( ~n4421 & n5252 ) ;
  assign n5254 = ( ~n2628 & n4660 ) | ( ~n2628 & n5253 ) | ( n4660 & n5253 ) ;
  assign n5255 = ( n4946 & ~n5001 ) | ( n4946 & n5254 ) | ( ~n5001 & n5254 ) ;
  assign n5256 = ( ~n1402 & n1845 ) | ( ~n1402 & n2656 ) | ( n1845 & n2656 ) ;
  assign n5257 = ( n2788 & n5255 ) | ( n2788 & ~n5256 ) | ( n5255 & ~n5256 ) ;
  assign n5258 = ( n2792 & ~n2800 ) | ( n2792 & n5257 ) | ( ~n2800 & n5257 ) ;
  assign n5259 = n5243 & n5258 ;
  assign n5260 = n630 | n662 ;
  assign n5261 = n686 | n707 ;
  assign n5262 = n5260 | n5261 ;
  assign n5263 = n519 | n593 ;
  assign n5264 = n572 | n581 ;
  assign n5265 = n5263 | n5264 ;
  assign n5266 = n5262 | n5265 ;
  assign n5267 = n788 | n800 ;
  assign n5268 = n829 | n852 ;
  assign n5269 = n5267 | n5268 ;
  assign n5270 = n701 | n727 ;
  assign n5271 = n752 | n758 ;
  assign n5272 = n5270 | n5271 ;
  assign n5273 = n5269 | n5272 ;
  assign n5274 = n5266 | n5273 ;
  assign n5275 = n326 | n332 ;
  assign n5276 = n357 | n414 ;
  assign n5277 = n5275 | n5276 ;
  assign n5278 = n261 | n272 ;
  assign n5279 = n285 | n306 ;
  assign n5280 = n5278 | n5279 ;
  assign n5281 = n5277 | n5280 ;
  assign n5282 = n490 | n497 ;
  assign n5283 = n525 | n531 ;
  assign n5284 = n5282 | n5283 ;
  assign n5285 = n396 | n434 ;
  assign n5286 = n425 | n428 ;
  assign n5287 = n5285 | n5286 ;
  assign n5288 = n5284 | n5287 ;
  assign n5289 = n5281 | n5288 ;
  assign n5290 = n5274 | n5289 ;
  assign n5291 = n1220 | n1223 ;
  assign n5292 = n1285 | n1292 ;
  assign n5293 = n5291 | n5292 ;
  assign n5294 = n1152 | n1209 ;
  assign n5295 = n1191 | n1229 ;
  assign n5296 = n5294 | n5295 ;
  assign n5297 = n5293 | n5296 ;
  assign n5298 = n1367 | n1376 ;
  assign n5299 = n1425 | n1574 ;
  assign n5300 = n5298 | n5299 ;
  assign n5301 = n1320 | n1326 ;
  assign n5302 = n1314 | n1388 ;
  assign n5303 = n5301 | n5302 ;
  assign n5304 = n5300 | n5303 ;
  assign n5305 = n5297 | n5304 ;
  assign n5306 = n920 | n1010 ;
  assign n5307 = n973 | n985 ;
  assign n5308 = n5306 | n5307 ;
  assign n5309 = n875 | n881 ;
  assign n5310 = n866 | n926 ;
  assign n5311 = n5309 | n5310 ;
  assign n5312 = n5308 | n5311 ;
  assign n5313 = n1080 | n1101 ;
  assign n5314 = n1121 | n1127 ;
  assign n5315 = n5313 | n5314 ;
  assign n5316 = n1025 | n1031 ;
  assign n5317 = n1056 | n1067 ;
  assign n5318 = n5316 | n5317 ;
  assign n5319 = n5315 | n5318 ;
  assign n5320 = n5312 | n5319 ;
  assign n5321 = n5305 | n5320 ;
  assign n5322 = n5290 | n5321 ;
  assign y0 = n654 ;
  assign y1 = n1052 ;
  assign y2 = n1449 ;
  assign y3 = n1588 ;
  assign y4 = n1727 ;
  assign y5 = n1862 ;
  assign y6 = n1971 ;
  assign y7 = n2080 ;
  assign y8 = n2188 ;
  assign y9 = n2284 ;
  assign y10 = n2380 ;
  assign y11 = n2475 ;
  assign y12 = n2544 ;
  assign y13 = n2613 ;
  assign y14 = n2680 ;
  assign y15 = n2724 ;
  assign y16 = n2768 ;
  assign y17 = n2812 ;
  assign y18 = n2842 ;
  assign y19 = n2872 ;
  assign y20 = n2901 ;
  assign y21 = n2930 ;
  assign y22 = n2959 ;
  assign y23 = n2988 ;
  assign y24 = n3017 ;
  assign y25 = n3046 ;
  assign y26 = n3073 ;
  assign y27 = n3100 ;
  assign y28 = n3127 ;
  assign y29 = n3154 ;
  assign y30 = n3181 ;
  assign y31 = n3208 ;
  assign y32 = n3234 ;
  assign y33 = n3260 ;
  assign y34 = n3286 ;
  assign y35 = n3312 ;
  assign y36 = n3338 ;
  assign y37 = n3364 ;
  assign y38 = n3390 ;
  assign y39 = n3416 ;
  assign y40 = n3442 ;
  assign y41 = n3468 ;
  assign y42 = n3494 ;
  assign y43 = n3520 ;
  assign y44 = n3545 ;
  assign y45 = n3570 ;
  assign y46 = n3595 ;
  assign y47 = n3620 ;
  assign y48 = n3645 ;
  assign y49 = n3670 ;
  assign y50 = n3694 ;
  assign y51 = n3718 ;
  assign y52 = n3742 ;
  assign y53 = n3766 ;
  assign y54 = n3790 ;
  assign y55 = n3814 ;
  assign y56 = n3838 ;
  assign y57 = n3862 ;
  assign y58 = n3886 ;
  assign y59 = n3909 ;
  assign y60 = n3932 ;
  assign y61 = n3955 ;
  assign y62 = n3978 ;
  assign y63 = n4001 ;
  assign y64 = n4024 ;
  assign y65 = n4047 ;
  assign y66 = n4070 ;
  assign y67 = n4093 ;
  assign y68 = n4116 ;
  assign y69 = n4139 ;
  assign y70 = n4162 ;
  assign y71 = n4184 ;
  assign y72 = n4206 ;
  assign y73 = n4228 ;
  assign y74 = n4250 ;
  assign y75 = n4272 ;
  assign y76 = n4294 ;
  assign y77 = n4316 ;
  assign y78 = n4338 ;
  assign y79 = n4360 ;
  assign y80 = n4382 ;
  assign y81 = n4404 ;
  assign y82 = n4426 ;
  assign y83 = n4446 ;
  assign y84 = n4466 ;
  assign y85 = n4486 ;
  assign y86 = n4506 ;
  assign y87 = n4526 ;
  assign y88 = n4546 ;
  assign y89 = n4566 ;
  assign y90 = n4586 ;
  assign y91 = n4606 ;
  assign y92 = n4626 ;
  assign y93 = n4646 ;
  assign y94 = n4666 ;
  assign y95 = n4685 ;
  assign y96 = n4704 ;
  assign y97 = n4723 ;
  assign y98 = n4742 ;
  assign y99 = n4761 ;
  assign y100 = n4780 ;
  assign y101 = n4799 ;
  assign y102 = n4818 ;
  assign y103 = n4837 ;
  assign y104 = n4856 ;
  assign y105 = n4875 ;
  assign y106 = n4894 ;
  assign y107 = n4913 ;
  assign y108 = n4932 ;
  assign y109 = n4951 ;
  assign y110 = n4969 ;
  assign y111 = n4987 ;
  assign y112 = n5005 ;
  assign y113 = n5022 ;
  assign y114 = n5039 ;
  assign y115 = n5056 ;
  assign y116 = n5073 ;
  assign y117 = n5090 ;
  assign y118 = n5107 ;
  assign y119 = n5124 ;
  assign y120 = n5141 ;
  assign y121 = n5158 ;
  assign y122 = n5175 ;
  assign y123 = n5192 ;
  assign y124 = n5209 ;
  assign y125 = n5225 ;
  assign y126 = n5242 ;
  assign y127 = n5259 ;
  assign y128 = n5322 ;
endmodule
