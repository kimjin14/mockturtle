module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 ;
  wire n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , n3931 , n3932 , n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , n3940 , n3941 , n3942 , n3943 , n3944 , n3945 , n3946 , n3947 , n3948 , n3949 , n3950 , n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , n3970 , n3971 , n3972 , n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , n3980 , n3981 , n3982 , n3983 , n3984 , n3985 , n3986 , n3987 , n3988 , n3989 , n3990 , n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , n4000 , n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , n4009 , n4010 , n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , n4019 , n4020 , n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , n4029 , n4030 , n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , n4039 , n4040 , n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4049 , n4050 , n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , n4059 , n4060 , n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , n4070 , n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , n4079 , n4080 , n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , n4089 , n4090 , n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , n4097 , n4098 , n4099 , n4100 , n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , n4109 , n4110 , n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , n4119 , n4120 , n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , n4129 , n4130 , n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , n4139 , n4140 , n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , n4150 , n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , n4159 , n4160 , n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , n4169 , n4170 , n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , n4179 , n4180 , n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , n4189 , n4190 , n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , n4197 , n4198 , n4199 , n4200 , n4201 , n4202 , n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , n4209 , n4210 , n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , n4217 , n4218 , n4219 , n4220 , n4221 , n4222 , n4223 , n4224 , n4225 , n4226 , n4227 , n4228 , n4229 , n4230 , n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , n4237 , n4238 , n4239 , n4240 , n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , n4247 , n4248 , n4249 , n4250 , n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , n4259 , n4260 , n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , n4269 , n4270 , n4271 , n4272 , n4273 , n4274 , n4275 , n4276 , n4277 , n4278 , n4279 , n4280 , n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , n4289 , n4290 , n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , n4299 , n4300 , n4301 , n4302 , n4303 , n4304 , n4305 , n4306 , n4307 , n4308 , n4309 , n4310 , n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , n4319 , n4320 , n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , n4329 , n4330 , n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , n4340 , n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , n4349 , n4350 , n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , n4360 , n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , n4370 , n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , n4380 , n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , n4390 , n4391 , n4392 , n4393 , n4394 , n4395 , n4396 , n4397 , n4398 , n4399 , n4400 , n4401 , n4402 , n4403 , n4404 , n4405 , n4406 , n4407 , n4408 , n4409 , n4410 , n4411 , n4412 , n4413 , n4414 , n4415 , n4416 , n4417 , n4418 , n4419 , n4420 , n4421 , n4422 , n4423 , n4424 , n4425 , n4426 , n4427 , n4428 , n4429 , n4430 , n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , n4437 , n4438 , n4439 , n4440 , n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , n4449 , n4450 , n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , n4459 , n4460 , n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , n4469 , n4470 , n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , n4479 , n4480 , n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , n4487 , n4488 , n4489 , n4490 , n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , n4497 , n4498 , n4499 , n4500 , n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , n4509 , n4510 , n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , n4519 , n4520 , n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , n4529 , n4530 , n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , n4537 , n4538 , n4539 , n4540 , n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , n4547 , n4548 , n4549 , n4550 , n4551 , n4552 , n4553 , n4554 , n4555 , n4556 , n4557 , n4558 , n4559 , n4560 , n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , n4567 , n4568 , n4569 , n4570 , n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , n4579 , n4580 , n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , n4589 , n4590 , n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , n4597 , n4598 , n4599 , n4600 , n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , n4607 , n4608 , n4609 , n4610 , n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , n4617 , n4618 , n4619 , n4620 , n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , n4627 , n4628 , n4629 , n4630 , n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , n4637 , n4638 , n4639 , n4640 , n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , n4647 , n4648 , n4649 , n4650 , n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , n4657 , n4658 , n4659 , n4660 , n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , n4669 , n4670 , n4671 , n4672 , n4673 , n4674 , n4675 , n4676 , n4677 , n4678 , n4679 , n4680 , n4681 , n4682 , n4683 , n4684 , n4685 , n4686 , n4687 , n4688 , n4689 , n4690 , n4691 , n4692 , n4693 , n4694 , n4695 , n4696 , n4697 , n4698 , n4699 , n4700 , n4701 , n4702 , n4703 , n4704 , n4705 , n4706 , n4707 , n4708 , n4709 , n4710 , n4711 , n4712 , n4713 , n4714 , n4715 , n4716 , n4717 , n4718 , n4719 , n4720 , n4721 , n4722 , n4723 , n4724 , n4725 , n4726 , n4727 , n4728 , n4729 , n4730 , n4731 , n4732 , n4733 , n4734 , n4735 , n4736 , n4737 , n4738 , n4739 , n4740 , n4741 , n4742 , n4743 , n4744 , n4745 , n4746 , n4747 , n4748 , n4749 , n4750 , n4751 , n4752 , n4753 , n4754 , n4755 , n4756 , n4757 , n4758 , n4759 , n4760 , n4761 , n4762 , n4763 , n4764 , n4765 , n4766 , n4767 , n4768 , n4769 , n4770 , n4771 , n4772 , n4773 , n4774 , n4775 , n4776 , n4777 , n4778 , n4779 , n4780 , n4781 , n4782 , n4783 , n4784 , n4785 , n4786 , n4787 , n4788 , n4789 , n4790 , n4791 , n4792 , n4793 , n4794 , n4795 , n4796 , n4797 , n4798 , n4799 , n4800 , n4801 , n4802 , n4803 , n4804 , n4805 , n4806 , n4807 , n4808 , n4809 , n4810 , n4811 , n4812 , n4813 , n4814 , n4815 , n4816 , n4817 , n4818 , n4819 , n4820 , n4821 , n4822 , n4823 , n4824 , n4825 , n4826 , n4827 , n4828 , n4829 , n4830 , n4831 , n4832 , n4833 , n4834 , n4835 , n4836 , n4837 , n4838 , n4839 , n4840 , n4841 , n4842 , n4843 , n4844 , n4845 , n4846 , n4847 , n4848 , n4849 , n4850 , n4851 , n4852 , n4853 , n4854 , n4855 , n4856 , n4857 , n4858 , n4859 , n4860 , n4861 , n4862 , n4863 , n4864 , n4865 , n4866 , n4867 , n4868 , n4869 , n4870 , n4871 , n4872 , n4873 , n4874 , n4875 , n4876 , n4877 , n4878 , n4879 , n4880 , n4881 , n4882 , n4883 , n4884 , n4885 , n4886 , n4887 , n4888 , n4889 , n4890 , n4891 , n4892 , n4893 , n4894 , n4895 , n4896 , n4897 , n4898 , n4899 , n4900 , n4901 , n4902 , n4903 , n4904 , n4905 , n4906 , n4907 , n4908 , n4909 , n4910 , n4911 , n4912 , n4913 , n4914 , n4915 , n4916 , n4917 , n4918 , n4919 , n4920 , n4921 , n4922 , n4923 , n4924 , n4925 , n4926 , n4927 , n4928 , n4929 , n4930 , n4931 , n4932 , n4933 , n4934 , n4935 , n4936 , n4937 , n4938 , n4939 , n4940 , n4941 , n4942 , n4943 , n4944 , n4945 , n4946 , n4947 , n4948 , n4949 , n4950 , n4951 , n4952 , n4953 , n4954 , n4955 , n4956 , n4957 , n4958 , n4959 , n4960 , n4961 , n4962 , n4963 , n4964 , n4965 , n4966 , n4967 , n4968 , n4969 , n4970 , n4971 , n4972 , n4973 , n4974 , n4975 , n4976 , n4977 , n4978 , n4979 , n4980 , n4981 , n4982 , n4983 , n4984 , n4985 , n4986 , n4987 , n4988 , n4989 , n4990 , n4991 , n4992 , n4993 , n4994 , n4995 , n4996 , n4997 , n4998 , n4999 , n5000 , n5001 , n5002 , n5003 , n5004 , n5005 , n5006 , n5007 , n5008 , n5009 , n5010 , n5011 , n5012 , n5013 , n5014 , n5015 , n5016 , n5017 , n5018 , n5019 , n5020 , n5021 , n5022 , n5023 , n5024 , n5025 , n5026 , n5027 , n5028 , n5029 , n5030 , n5031 , n5032 , n5033 , n5034 , n5035 , n5036 , n5037 , n5038 , n5039 , n5040 , n5041 , n5042 , n5043 , n5044 , n5045 , n5046 , n5047 , n5048 , n5049 , n5050 , n5051 , n5052 , n5053 , n5054 , n5055 , n5056 , n5057 , n5058 , n5059 , n5060 , n5061 , n5062 , n5063 , n5064 , n5065 , n5066 , n5067 , n5068 , n5069 , n5070 , n5071 , n5072 , n5073 , n5074 , n5075 , n5076 , n5077 , n5078 , n5079 , n5080 , n5081 , n5082 , n5083 , n5084 , n5085 , n5086 , n5087 , n5088 , n5089 , n5090 , n5091 , n5092 , n5093 , n5094 , n5095 , n5096 , n5097 , n5098 , n5099 , n5100 , n5101 , n5102 , n5103 , n5104 , n5105 , n5106 , n5107 , n5108 , n5109 , n5110 , n5111 , n5112 , n5113 , n5114 , n5115 , n5116 , n5117 , n5118 , n5119 , n5120 , n5121 , n5122 , n5123 , n5124 , n5125 , n5126 , n5127 , n5128 , n5129 , n5130 , n5131 , n5132 , n5133 , n5134 , n5135 , n5136 , n5137 , n5138 , n5139 , n5140 , n5141 , n5142 , n5143 , n5144 , n5145 , n5146 , n5147 , n5148 , n5149 , n5150 , n5151 , n5152 , n5153 , n5154 , n5155 , n5156 , n5157 , n5158 , n5159 , n5160 , n5161 , n5162 , n5163 , n5164 , n5165 , n5166 , n5167 , n5168 , n5169 , n5170 , n5171 , n5172 , n5173 , n5174 , n5175 , n5176 , n5177 , n5178 , n5179 , n5180 , n5181 , n5182 , n5183 , n5184 , n5185 , n5186 , n5187 , n5188 , n5189 , n5190 , n5191 , n5192 , n5193 , n5194 , n5195 , n5196 , n5197 , n5198 , n5199 , n5200 , n5201 , n5202 , n5203 , n5204 , n5205 , n5206 , n5207 , n5208 , n5209 , n5210 , n5211 , n5212 , n5213 , n5214 , n5215 , n5216 , n5217 , n5218 , n5219 , n5220 , n5221 , n5222 , n5223 , n5224 , n5225 , n5226 , n5227 , n5228 , n5229 , n5230 , n5231 , n5232 , n5233 , n5234 , n5235 , n5236 , n5237 , n5238 , n5239 , n5240 , n5241 , n5242 , n5243 , n5244 , n5245 , n5246 , n5247 , n5248 , n5249 , n5250 , n5251 , n5252 , n5253 , n5254 , n5255 , n5256 , n5257 , n5258 , n5259 , n5260 , n5261 , n5262 , n5263 , n5264 , n5265 , n5266 , n5267 , n5268 , n5269 , n5270 , n5271 , n5272 , n5273 , n5274 , n5275 , n5276 , n5277 , n5278 , n5279 , n5280 , n5281 , n5282 , n5283 , n5284 , n5285 , n5286 , n5287 , n5288 , n5289 , n5290 , n5291 , n5292 , n5293 , n5294 , n5295 , n5296 , n5297 , n5298 , n5299 , n5300 , n5301 , n5302 , n5303 , n5304 , n5305 , n5306 , n5307 , n5308 , n5309 , n5310 , n5311 , n5312 , n5313 , n5314 , n5315 , n5316 , n5317 , n5318 , n5319 , n5320 , n5321 , n5322 , n5323 , n5324 , n5325 , n5326 , n5327 , n5328 , n5329 , n5330 , n5331 , n5332 , n5333 , n5334 , n5335 , n5336 , n5337 , n5338 , n5339 , n5340 , n5341 , n5342 , n5343 , n5344 , n5345 , n5346 , n5347 , n5348 , n5349 , n5350 , n5351 , n5352 , n5353 , n5354 , n5355 , n5356 , n5357 , n5358 , n5359 , n5360 , n5361 , n5362 , n5363 , n5364 , n5365 , n5366 , n5367 , n5368 , n5369 , n5370 , n5371 , n5372 , n5373 , n5374 , n5375 , n5376 , n5377 , n5378 , n5379 , n5380 , n5381 , n5382 , n5383 , n5384 , n5385 , n5386 , n5387 , n5388 , n5389 , n5390 , n5391 , n5392 , n5393 , n5394 , n5395 , n5396 , n5397 , n5398 , n5399 , n5400 , n5401 , n5402 , n5403 , n5404 , n5405 , n5406 , n5407 , n5408 , n5409 , n5410 , n5411 , n5412 , n5413 , n5414 , n5415 , n5416 , n5417 , n5418 , n5419 , n5420 , n5421 , n5422 , n5423 , n5424 , n5425 , n5426 , n5427 , n5428 , n5429 , n5430 , n5431 , n5432 , n5433 , n5434 , n5435 , n5436 , n5437 , n5438 , n5439 , n5440 , n5441 , n5442 , n5443 , n5444 , n5445 , n5446 , n5447 , n5448 , n5449 , n5450 , n5451 , n5452 , n5453 , n5454 , n5455 , n5456 , n5457 , n5458 , n5459 , n5460 , n5461 , n5462 , n5463 , n5464 , n5465 , n5466 , n5467 , n5468 , n5469 , n5470 , n5471 , n5472 , n5473 , n5474 , n5475 , n5476 , n5477 , n5478 , n5479 , n5480 , n5481 , n5482 , n5483 , n5484 , n5485 , n5486 , n5487 , n5488 , n5489 , n5490 , n5491 , n5492 , n5493 , n5494 , n5495 , n5496 , n5497 , n5498 , n5499 , n5500 , n5501 , n5502 , n5503 , n5504 , n5505 , n5506 , n5507 , n5508 , n5509 , n5510 , n5511 , n5512 , n5513 , n5514 , n5515 , n5516 , n5517 , n5518 , n5519 , n5520 , n5521 , n5522 , n5523 , n5524 , n5525 , n5526 , n5527 , n5528 , n5529 , n5530 , n5531 , n5532 , n5533 , n5534 , n5535 , n5536 , n5537 , n5538 , n5539 , n5540 , n5541 , n5542 , n5543 , n5544 , n5545 , n5546 , n5547 , n5548 , n5549 , n5550 , n5551 , n5552 , n5553 , n5554 , n5555 , n5556 , n5557 , n5558 , n5559 , n5560 , n5561 , n5562 , n5563 , n5564 , n5565 , n5566 , n5567 , n5568 , n5569 , n5570 , n5571 , n5572 , n5573 , n5574 , n5575 , n5576 , n5577 , n5578 , n5579 , n5580 , n5581 , n5582 , n5583 , n5584 , n5585 , n5586 , n5587 , n5588 , n5589 , n5590 , n5591 , n5592 , n5593 , n5594 , n5595 , n5596 , n5597 , n5598 , n5599 , n5600 , n5601 , n5602 , n5603 , n5604 , n5605 , n5606 , n5607 , n5608 , n5609 , n5610 , n5611 , n5612 , n5613 , n5614 , n5615 , n5616 , n5617 , n5618 , n5619 , n5620 , n5621 , n5622 , n5623 , n5624 , n5625 , n5626 , n5627 , n5628 , n5629 , n5630 , n5631 , n5632 , n5633 , n5634 , n5635 , n5636 , n5637 , n5638 , n5639 , n5640 , n5641 , n5642 , n5643 , n5644 , n5645 , n5646 , n5647 , n5648 , n5649 , n5650 , n5651 , n5652 , n5653 , n5654 , n5655 , n5656 , n5657 , n5658 , n5659 , n5660 , n5661 , n5662 , n5663 , n5664 , n5665 , n5666 , n5667 , n5668 , n5669 , n5670 , n5671 , n5672 , n5673 , n5674 , n5675 , n5676 , n5677 , n5678 , n5679 , n5680 , n5681 , n5682 , n5683 , n5684 , n5685 , n5686 , n5687 , n5688 , n5689 , n5690 , n5691 , n5692 , n5693 , n5694 , n5695 , n5696 , n5697 , n5698 , n5699 , n5700 , n5701 , n5702 , n5703 , n5704 , n5705 , n5706 , n5707 , n5708 , n5709 , n5710 , n5711 , n5712 , n5713 , n5714 , n5715 , n5716 , n5717 , n5718 , n5719 , n5720 , n5721 , n5722 , n5723 , n5724 , n5725 , n5726 , n5727 , n5728 , n5729 , n5730 , n5731 , n5732 , n5733 , n5734 , n5735 , n5736 , n5737 , n5738 , n5739 , n5740 , n5741 , n5742 , n5743 , n5744 , n5745 , n5746 , n5747 , n5748 , n5749 , n5750 , n5751 , n5752 , n5753 , n5754 , n5755 , n5756 , n5757 , n5758 , n5759 , n5760 , n5761 , n5762 , n5763 , n5764 , n5765 , n5766 , n5767 , n5768 , n5769 , n5770 , n5771 , n5772 , n5773 , n5774 , n5775 , n5776 , n5777 , n5778 , n5779 , n5780 , n5781 , n5782 , n5783 , n5784 , n5785 , n5786 , n5787 , n5788 , n5789 , n5790 , n5791 , n5792 , n5793 , n5794 , n5795 , n5796 , n5797 , n5798 , n5799 , n5800 , n5801 , n5802 , n5803 , n5804 , n5805 , n5806 , n5807 , n5808 , n5809 , n5810 , n5811 , n5812 , n5813 , n5814 , n5815 , n5816 , n5817 , n5818 , n5819 , n5820 , n5821 , n5822 , n5823 , n5824 , n5825 , n5826 , n5827 , n5828 , n5829 , n5830 , n5831 , n5832 , n5833 , n5834 , n5835 , n5836 , n5837 , n5838 , n5839 , n5840 , n5841 , n5842 , n5843 , n5844 , n5845 , n5846 , n5847 , n5848 , n5849 , n5850 , n5851 , n5852 , n5853 , n5854 , n5855 , n5856 , n5857 , n5858 , n5859 , n5860 , n5861 , n5862 , n5863 , n5864 , n5865 , n5866 , n5867 , n5868 , n5869 , n5870 , n5871 , n5872 , n5873 , n5874 , n5875 , n5876 , n5877 , n5878 , n5879 , n5880 , n5881 , n5882 , n5883 , n5884 , n5885 , n5886 , n5887 , n5888 , n5889 , n5890 , n5891 , n5892 , n5893 , n5894 , n5895 , n5896 , n5897 , n5898 , n5899 , n5900 , n5901 , n5902 , n5903 , n5904 , n5905 , n5906 , n5907 , n5908 , n5909 , n5910 , n5911 , n5912 , n5913 , n5914 , n5915 , n5916 , n5917 , n5918 , n5919 , n5920 , n5921 , n5922 , n5923 , n5924 , n5925 , n5926 , n5927 , n5928 , n5929 , n5930 , n5931 , n5932 , n5933 , n5934 , n5935 , n5936 , n5937 , n5938 , n5939 , n5940 , n5941 , n5942 , n5943 , n5944 , n5945 , n5946 , n5947 , n5948 , n5949 , n5950 , n5951 , n5952 , n5953 , n5954 , n5955 , n5956 , n5957 , n5958 , n5959 , n5960 , n5961 , n5962 , n5963 , n5964 , n5965 , n5966 , n5967 , n5968 , n5969 , n5970 , n5971 , n5972 , n5973 , n5974 , n5975 , n5976 , n5977 , n5978 , n5979 , n5980 , n5981 , n5982 , n5983 , n5984 , n5985 , n5986 , n5987 , n5988 , n5989 , n5990 , n5991 , n5992 , n5993 , n5994 , n5995 , n5996 , n5997 , n5998 , n5999 , n6000 , n6001 , n6002 , n6003 , n6004 , n6005 , n6006 , n6007 , n6008 , n6009 , n6010 , n6011 , n6012 , n6013 , n6014 , n6015 , n6016 , n6017 , n6018 , n6019 , n6020 , n6021 , n6022 , n6023 , n6024 , n6025 , n6026 , n6027 , n6028 , n6029 , n6030 , n6031 , n6032 , n6033 , n6034 , n6035 , n6036 , n6037 , n6038 , n6039 , n6040 , n6041 , n6042 , n6043 , n6044 , n6045 , n6046 , n6047 , n6048 , n6049 , n6050 , n6051 , n6052 , n6053 , n6054 , n6055 , n6056 , n6057 , n6058 , n6059 , n6060 , n6061 , n6062 , n6063 , n6064 , n6065 , n6066 , n6067 , n6068 , n6069 , n6070 , n6071 , n6072 , n6073 , n6074 , n6075 , n6076 , n6077 , n6078 , n6079 , n6080 , n6081 , n6082 , n6083 , n6084 , n6085 , n6086 , n6087 , n6088 , n6089 , n6090 , n6091 , n6092 , n6093 , n6094 , n6095 , n6096 , n6097 , n6098 , n6099 , n6100 , n6101 , n6102 , n6103 , n6104 , n6105 , n6106 , n6107 , n6108 , n6109 , n6110 , n6111 , n6112 , n6113 , n6114 , n6115 , n6116 , n6117 , n6118 , n6119 , n6120 , n6121 , n6122 , n6123 , n6124 , n6125 , n6126 , n6127 , n6128 , n6129 , n6130 , n6131 , n6132 , n6133 , n6134 , n6135 , n6136 , n6137 , n6138 , n6139 , n6140 , n6141 , n6142 , n6143 , n6144 , n6145 , n6146 , n6147 , n6148 , n6149 , n6150 , n6151 , n6152 , n6153 , n6154 , n6155 , n6156 , n6157 , n6158 , n6159 , n6160 , n6161 , n6162 , n6163 , n6164 , n6165 , n6166 , n6167 , n6168 , n6169 , n6170 , n6171 , n6172 , n6173 , n6174 , n6175 , n6176 , n6177 , n6178 , n6179 , n6180 , n6181 , n6182 , n6183 , n6184 , n6185 , n6186 , n6187 , n6188 , n6189 , n6190 , n6191 , n6192 , n6193 , n6194 , n6195 , n6196 , n6197 , n6198 , n6199 , n6200 , n6201 , n6202 , n6203 , n6204 , n6205 , n6206 , n6207 , n6208 , n6209 , n6210 , n6211 , n6212 , n6213 , n6214 , n6215 , n6216 , n6217 , n6218 , n6219 , n6220 , n6221 , n6222 , n6223 , n6224 , n6225 , n6226 , n6227 , n6228 , n6229 , n6230 , n6231 , n6232 , n6233 , n6234 , n6235 , n6236 , n6237 , n6238 , n6239 , n6240 , n6241 , n6242 , n6243 , n6244 , n6245 , n6246 , n6247 , n6248 , n6249 , n6250 , n6251 , n6252 , n6253 , n6254 , n6255 , n6256 , n6257 , n6258 , n6259 , n6260 , n6261 , n6262 , n6263 , n6264 , n6265 , n6266 , n6267 , n6268 , n6269 , n6270 , n6271 , n6272 , n6273 , n6274 , n6275 , n6276 , n6277 , n6278 , n6279 , n6280 , n6281 , n6282 , n6283 , n6284 , n6285 , n6286 , n6287 , n6288 , n6289 , n6290 , n6291 , n6292 , n6293 , n6294 , n6295 , n6296 , n6297 , n6298 , n6299 , n6300 , n6301 , n6302 , n6303 , n6304 , n6305 , n6306 , n6307 , n6308 , n6309 , n6310 , n6311 , n6312 , n6313 , n6314 , n6315 , n6316 , n6317 , n6318 , n6319 , n6320 , n6321 , n6322 , n6323 , n6324 , n6325 , n6326 , n6327 , n6328 , n6329 , n6330 , n6331 , n6332 , n6333 , n6334 , n6335 , n6336 , n6337 , n6338 , n6339 , n6340 , n6341 , n6342 , n6343 , n6344 , n6345 , n6346 , n6347 , n6348 , n6349 , n6350 , n6351 , n6352 , n6353 , n6354 , n6355 , n6356 , n6357 , n6358 , n6359 , n6360 , n6361 , n6362 , n6363 , n6364 , n6365 , n6366 , n6367 , n6368 , n6369 , n6370 , n6371 , n6372 , n6373 , n6374 , n6375 , n6376 , n6377 , n6378 , n6379 , n6380 , n6381 , n6382 , n6383 , n6384 , n6385 , n6386 , n6387 , n6388 , n6389 , n6390 , n6391 , n6392 , n6393 , n6394 , n6395 , n6396 , n6397 , n6398 , n6399 , n6400 , n6401 , n6402 , n6403 , n6404 , n6405 , n6406 , n6407 , n6408 , n6409 , n6410 , n6411 , n6412 , n6413 , n6414 , n6415 , n6416 , n6417 , n6418 , n6419 , n6420 , n6421 , n6422 , n6423 , n6424 , n6425 , n6426 , n6427 , n6428 , n6429 , n6430 , n6431 , n6432 , n6433 , n6434 , n6435 , n6436 , n6437 , n6438 , n6439 , n6440 , n6441 , n6442 , n6443 , n6444 , n6445 , n6446 , n6447 , n6448 , n6449 , n6450 , n6451 , n6452 , n6453 , n6454 , n6455 , n6456 , n6457 , n6458 , n6459 , n6460 , n6461 , n6462 , n6463 , n6464 , n6465 , n6466 , n6467 , n6468 , n6469 , n6470 , n6471 , n6472 , n6473 , n6474 , n6475 , n6476 , n6477 , n6478 , n6479 , n6480 , n6481 , n6482 , n6483 , n6484 , n6485 , n6486 , n6487 , n6488 , n6489 , n6490 , n6491 , n6492 , n6493 , n6494 , n6495 , n6496 , n6497 , n6498 , n6499 , n6500 , n6501 , n6502 , n6503 , n6504 , n6505 , n6506 , n6507 , n6508 , n6509 , n6510 , n6511 , n6512 , n6513 , n6514 , n6515 , n6516 , n6517 , n6518 , n6519 , n6520 , n6521 , n6522 , n6523 , n6524 , n6525 , n6526 , n6527 , n6528 , n6529 , n6530 , n6531 , n6532 , n6533 , n6534 , n6535 , n6536 , n6537 , n6538 , n6539 , n6540 , n6541 , n6542 , n6543 , n6544 , n6545 , n6546 , n6547 , n6548 , n6549 , n6550 , n6551 , n6552 , n6553 , n6554 , n6555 , n6556 , n6557 , n6558 , n6559 , n6560 , n6561 , n6562 , n6563 , n6564 , n6565 , n6566 , n6567 , n6568 , n6569 , n6570 , n6571 , n6572 , n6573 , n6574 , n6575 , n6576 , n6577 , n6578 , n6579 , n6580 , n6581 , n6582 , n6583 , n6584 , n6585 , n6586 , n6587 , n6588 , n6589 , n6590 , n6591 , n6592 , n6593 , n6594 , n6595 , n6596 , n6597 , n6598 , n6599 , n6600 , n6601 , n6602 , n6603 , n6604 , n6605 , n6606 , n6607 , n6608 , n6609 , n6610 , n6611 , n6612 , n6613 , n6614 , n6615 , n6616 , n6617 , n6618 , n6619 , n6620 , n6621 , n6622 , n6623 , n6624 , n6625 , n6626 , n6627 , n6628 , n6629 , n6630 , n6631 , n6632 , n6633 , n6634 , n6635 , n6636 , n6637 , n6638 , n6639 , n6640 , n6641 , n6642 , n6643 , n6644 , n6645 , n6646 , n6647 , n6648 , n6649 , n6650 , n6651 , n6652 , n6653 , n6654 , n6655 , n6656 , n6657 , n6658 , n6659 , n6660 , n6661 , n6662 , n6663 , n6664 , n6665 , n6666 , n6667 , n6668 , n6669 , n6670 , n6671 , n6672 , n6673 , n6674 , n6675 , n6676 , n6677 , n6678 , n6679 , n6680 , n6681 , n6682 , n6683 , n6684 , n6685 , n6686 , n6687 , n6688 , n6689 , n6690 , n6691 , n6692 , n6693 , n6694 , n6695 , n6696 , n6697 , n6698 , n6699 , n6700 , n6701 , n6702 , n6703 , n6704 , n6705 , n6706 , n6707 , n6708 , n6709 , n6710 , n6711 , n6712 , n6713 , n6714 , n6715 , n6716 , n6717 , n6718 , n6719 , n6720 , n6721 , n6722 , n6723 , n6724 , n6725 , n6726 , n6727 , n6728 , n6729 , n6730 , n6731 , n6732 , n6733 , n6734 , n6735 , n6736 , n6737 , n6738 , n6739 , n6740 , n6741 , n6742 , n6743 , n6744 , n6745 , n6746 , n6747 , n6748 , n6749 , n6750 , n6751 , n6752 , n6753 , n6754 , n6755 , n6756 , n6757 , n6758 , n6759 , n6760 , n6761 , n6762 , n6763 , n6764 , n6765 , n6766 , n6767 , n6768 , n6769 , n6770 , n6771 , n6772 , n6773 , n6774 , n6775 , n6776 , n6777 , n6778 , n6779 , n6780 , n6781 , n6782 , n6783 , n6784 , n6785 , n6786 , n6787 , n6788 , n6789 , n6790 , n6791 , n6792 , n6793 , n6794 , n6795 , n6796 , n6797 , n6798 , n6799 , n6800 , n6801 , n6802 , n6803 , n6804 , n6805 , n6806 , n6807 , n6808 , n6809 , n6810 , n6811 , n6812 , n6813 , n6814 , n6815 , n6816 , n6817 , n6818 , n6819 , n6820 , n6821 , n6822 , n6823 , n6824 , n6825 , n6826 , n6827 , n6828 , n6829 , n6830 , n6831 , n6832 , n6833 , n6834 , n6835 , n6836 , n6837 , n6838 , n6839 , n6840 , n6841 , n6842 , n6843 , n6844 , n6845 , n6846 , n6847 , n6848 , n6849 , n6850 , n6851 , n6852 , n6853 , n6854 , n6855 , n6856 , n6857 , n6858 , n6859 , n6860 , n6861 , n6862 , n6863 , n6864 , n6865 , n6866 , n6867 , n6868 , n6869 , n6870 , n6871 , n6872 , n6873 , n6874 , n6875 , n6876 , n6877 , n6878 , n6879 , n6880 , n6881 , n6882 , n6883 , n6884 , n6885 , n6886 , n6887 , n6888 , n6889 , n6890 , n6891 , n6892 , n6893 , n6894 , n6895 , n6896 , n6897 , n6898 , n6899 , n6900 , n6901 , n6902 , n6903 , n6904 , n6905 , n6906 , n6907 , n6908 , n6909 , n6910 , n6911 , n6912 , n6913 , n6914 , n6915 , n6916 , n6917 , n6918 , n6919 , n6920 , n6921 , n6922 , n6923 , n6924 , n6925 , n6926 , n6927 , n6928 , n6929 , n6930 , n6931 , n6932 , n6933 , n6934 , n6935 , n6936 , n6937 , n6938 , n6939 , n6940 , n6941 , n6942 , n6943 , n6944 , n6945 , n6946 , n6947 , n6948 , n6949 , n6950 , n6951 , n6952 , n6953 , n6954 , n6955 , n6956 , n6957 , n6958 , n6959 , n6960 , n6961 , n6962 , n6963 , n6964 , n6965 , n6966 , n6967 , n6968 , n6969 , n6970 , n6971 , n6972 , n6973 , n6974 , n6975 , n6976 , n6977 , n6978 , n6979 , n6980 , n6981 , n6982 , n6983 , n6984 , n6985 , n6986 , n6987 , n6988 , n6989 , n6990 , n6991 , n6992 , n6993 , n6994 , n6995 , n6996 , n6997 , n6998 , n6999 , n7000 , n7001 , n7002 , n7003 , n7004 , n7005 , n7006 , n7007 , n7008 , n7009 , n7010 , n7011 , n7012 , n7013 , n7014 , n7015 , n7016 , n7017 , n7018 , n7019 , n7020 , n7021 , n7022 , n7023 , n7024 , n7025 , n7026 , n7027 , n7028 , n7029 , n7030 , n7031 , n7032 , n7033 , n7034 , n7035 , n7036 , n7037 , n7038 , n7039 , n7040 , n7041 , n7042 , n7043 , n7044 , n7045 , n7046 , n7047 , n7048 , n7049 , n7050 , n7051 , n7052 , n7053 , n7054 , n7055 , n7056 , n7057 , n7058 , n7059 , n7060 , n7061 , n7062 , n7063 , n7064 , n7065 , n7066 , n7067 , n7068 , n7069 , n7070 , n7071 , n7072 , n7073 , n7074 , n7075 , n7076 , n7077 , n7078 , n7079 , n7080 , n7081 , n7082 , n7083 , n7084 , n7085 , n7086 , n7087 , n7088 , n7089 , n7090 , n7091 , n7092 , n7093 , n7094 , n7095 , n7096 , n7097 , n7098 , n7099 , n7100 , n7101 , n7102 , n7103 , n7104 , n7105 , n7106 , n7107 , n7108 , n7109 , n7110 , n7111 , n7112 , n7113 , n7114 , n7115 , n7116 , n7117 , n7118 , n7119 , n7120 , n7121 , n7122 , n7123 , n7124 , n7125 , n7126 , n7127 , n7128 , n7129 , n7130 , n7131 , n7132 , n7133 , n7134 , n7135 , n7136 , n7137 , n7138 , n7139 , n7140 , n7141 , n7142 , n7143 , n7144 , n7145 , n7146 , n7147 , n7148 , n7149 , n7150 , n7151 , n7152 , n7153 , n7154 , n7155 , n7156 , n7157 , n7158 , n7159 , n7160 , n7161 , n7162 , n7163 , n7164 , n7165 , n7166 , n7167 , n7168 , n7169 , n7170 , n7171 , n7172 , n7173 , n7174 , n7175 , n7176 , n7177 , n7178 , n7179 , n7180 , n7181 , n7182 , n7183 , n7184 , n7185 , n7186 , n7187 , n7188 , n7189 , n7190 , n7191 , n7192 , n7193 , n7194 , n7195 , n7196 , n7197 , n7198 , n7199 , n7200 , n7201 , n7202 , n7203 , n7204 , n7205 , n7206 , n7207 , n7208 , n7209 , n7210 , n7211 , n7212 , n7213 , n7214 , n7215 , n7216 , n7217 , n7218 , n7219 , n7220 , n7221 , n7222 , n7223 , n7224 , n7225 , n7226 , n7227 , n7228 , n7229 , n7230 , n7231 , n7232 , n7233 , n7234 , n7235 , n7236 , n7237 , n7238 , n7239 , n7240 , n7241 , n7242 , n7243 , n7244 , n7245 , n7246 , n7247 , n7248 , n7249 , n7250 , n7251 , n7252 , n7253 , n7254 , n7255 , n7256 , n7257 , n7258 , n7259 , n7260 , n7261 , n7262 , n7263 , n7264 , n7265 , n7266 , n7267 , n7268 , n7269 , n7270 , n7271 , n7272 , n7273 , n7274 , n7275 , n7276 , n7277 , n7278 , n7279 , n7280 , n7281 , n7282 , n7283 , n7284 , n7285 , n7286 , n7287 , n7288 , n7289 , n7290 , n7291 , n7292 , n7293 , n7294 , n7295 , n7296 , n7297 , n7298 , n7299 , n7300 , n7301 , n7302 , n7303 , n7304 , n7305 , n7306 , n7307 , n7308 , n7309 , n7310 , n7311 , n7312 , n7313 , n7314 , n7315 , n7316 , n7317 , n7318 , n7319 , n7320 , n7321 , n7322 , n7323 , n7324 , n7325 , n7326 , n7327 , n7328 , n7329 , n7330 , n7331 , n7332 , n7333 , n7334 , n7335 , n7336 , n7337 , n7338 , n7339 , n7340 , n7341 , n7342 , n7343 , n7344 , n7345 , n7346 , n7347 , n7348 , n7349 , n7350 , n7351 , n7352 , n7353 , n7354 , n7355 , n7356 , n7357 , n7358 , n7359 , n7360 , n7361 , n7362 , n7363 , n7364 , n7365 , n7366 , n7367 , n7368 , n7369 , n7370 , n7371 , n7372 , n7373 , n7374 , n7375 , n7376 , n7377 , n7378 , n7379 , n7380 , n7381 , n7382 , n7383 , n7384 , n7385 , n7386 , n7387 , n7388 , n7389 , n7390 , n7391 , n7392 , n7393 , n7394 , n7395 , n7396 , n7397 , n7398 , n7399 , n7400 , n7401 , n7402 , n7403 , n7404 , n7405 , n7406 , n7407 , n7408 , n7409 , n7410 , n7411 , n7412 , n7413 , n7414 , n7415 , n7416 , n7417 , n7418 , n7419 , n7420 , n7421 , n7422 , n7423 , n7424 , n7425 , n7426 , n7427 , n7428 , n7429 , n7430 , n7431 , n7432 , n7433 , n7434 , n7435 , n7436 , n7437 , n7438 , n7439 , n7440 , n7441 , n7442 , n7443 , n7444 , n7445 , n7446 , n7447 , n7448 , n7449 , n7450 , n7451 , n7452 , n7453 , n7454 , n7455 , n7456 , n7457 , n7458 , n7459 , n7460 , n7461 , n7462 , n7463 , n7464 , n7465 , n7466 , n7467 , n7468 , n7469 , n7470 , n7471 , n7472 , n7473 , n7474 , n7475 , n7476 , n7477 , n7478 , n7479 , n7480 , n7481 , n7482 , n7483 , n7484 , n7485 , n7486 , n7487 , n7488 , n7489 , n7490 , n7491 , n7492 , n7493 , n7494 , n7495 , n7496 , n7497 , n7498 , n7499 , n7500 , n7501 , n7502 , n7503 , n7504 , n7505 , n7506 , n7507 , n7508 , n7509 , n7510 , n7511 , n7512 , n7513 , n7514 , n7515 , n7516 , n7517 , n7518 , n7519 , n7520 , n7521 , n7522 , n7523 , n7524 , n7525 , n7526 , n7527 , n7528 , n7529 , n7530 , n7531 , n7532 , n7533 , n7534 , n7535 , n7536 , n7537 , n7538 , n7539 , n7540 , n7541 , n7542 , n7543 , n7544 , n7545 , n7546 , n7547 , n7548 , n7549 , n7550 , n7551 , n7552 , n7553 , n7554 , n7555 , n7556 , n7557 , n7558 , n7559 , n7560 , n7561 , n7562 , n7563 , n7564 , n7565 , n7566 , n7567 , n7568 , n7569 , n7570 , n7571 , n7572 , n7573 , n7574 , n7575 , n7576 , n7577 , n7578 , n7579 , n7580 , n7581 , n7582 , n7583 , n7584 , n7585 , n7586 , n7587 , n7588 , n7589 , n7590 , n7591 , n7592 , n7593 , n7594 , n7595 , n7596 , n7597 , n7598 , n7599 , n7600 , n7601 , n7602 , n7603 , n7604 , n7605 , n7606 , n7607 , n7608 , n7609 , n7610 , n7611 , n7612 , n7613 , n7614 , n7615 , n7616 , n7617 , n7618 , n7619 , n7620 , n7621 , n7622 , n7623 , n7624 , n7625 , n7626 , n7627 , n7628 , n7629 , n7630 , n7631 , n7632 , n7633 , n7634 , n7635 , n7636 , n7637 , n7638 , n7639 , n7640 , n7641 , n7642 , n7643 , n7644 , n7645 , n7646 , n7647 , n7648 , n7649 , n7650 , n7651 , n7652 , n7653 , n7654 , n7655 , n7656 , n7657 , n7658 , n7659 , n7660 , n7661 , n7662 , n7663 , n7664 , n7665 , n7666 , n7667 , n7668 , n7669 , n7670 , n7671 , n7672 , n7673 , n7674 , n7675 , n7676 , n7677 , n7678 , n7679 , n7680 , n7681 , n7682 , n7683 , n7684 , n7685 , n7686 , n7687 , n7688 , n7689 , n7690 , n7691 , n7692 , n7693 , n7694 , n7695 , n7696 , n7697 , n7698 , n7699 , n7700 , n7701 , n7702 , n7703 , n7704 , n7705 , n7706 , n7707 , n7708 , n7709 , n7710 , n7711 , n7712 , n7713 , n7714 , n7715 , n7716 , n7717 , n7718 , n7719 , n7720 , n7721 , n7722 , n7723 , n7724 , n7725 , n7726 , n7727 , n7728 , n7729 , n7730 , n7731 , n7732 , n7733 , n7734 , n7735 , n7736 , n7737 , n7738 , n7739 , n7740 , n7741 , n7742 , n7743 , n7744 , n7745 , n7746 , n7747 , n7748 , n7749 , n7750 , n7751 , n7752 , n7753 , n7754 , n7755 , n7756 , n7757 , n7758 , n7759 , n7760 , n7761 , n7762 , n7763 , n7764 , n7765 , n7766 , n7767 , n7768 , n7769 , n7770 , n7771 , n7772 , n7773 , n7774 , n7775 , n7776 , n7777 , n7778 , n7779 , n7780 , n7781 , n7782 , n7783 , n7784 , n7785 , n7786 , n7787 , n7788 , n7789 , n7790 , n7791 , n7792 , n7793 , n7794 , n7795 , n7796 , n7797 , n7798 , n7799 , n7800 , n7801 , n7802 , n7803 , n7804 , n7805 , n7806 , n7807 , n7808 , n7809 , n7810 , n7811 , n7812 , n7813 , n7814 , n7815 , n7816 , n7817 , n7818 , n7819 , n7820 , n7821 , n7822 , n7823 , n7824 , n7825 , n7826 , n7827 , n7828 , n7829 , n7830 , n7831 , n7832 , n7833 , n7834 , n7835 , n7836 , n7837 , n7838 , n7839 , n7840 , n7841 , n7842 , n7843 , n7844 , n7845 , n7846 , n7847 , n7848 , n7849 , n7850 , n7851 , n7852 , n7853 , n7854 , n7855 , n7856 , n7857 , n7858 , n7859 , n7860 , n7861 , n7862 , n7863 , n7864 , n7865 , n7866 , n7867 , n7868 , n7869 , n7870 , n7871 , n7872 , n7873 , n7874 , n7875 , n7876 , n7877 , n7878 , n7879 , n7880 , n7881 , n7882 , n7883 , n7884 , n7885 , n7886 , n7887 , n7888 , n7889 , n7890 , n7891 , n7892 , n7893 , n7894 , n7895 , n7896 , n7897 , n7898 , n7899 , n7900 , n7901 , n7902 , n7903 , n7904 , n7905 , n7906 , n7907 , n7908 , n7909 , n7910 , n7911 , n7912 , n7913 , n7914 , n7915 , n7916 , n7917 , n7918 , n7919 , n7920 , n7921 , n7922 , n7923 , n7924 , n7925 , n7926 , n7927 , n7928 , n7929 , n7930 , n7931 , n7932 , n7933 , n7934 , n7935 , n7936 , n7937 , n7938 , n7939 , n7940 , n7941 , n7942 , n7943 , n7944 , n7945 , n7946 , n7947 , n7948 , n7949 , n7950 , n7951 , n7952 , n7953 , n7954 , n7955 , n7956 , n7957 , n7958 , n7959 , n7960 , n7961 , n7962 , n7963 , n7964 , n7965 , n7966 , n7967 , n7968 , n7969 , n7970 , n7971 , n7972 , n7973 , n7974 , n7975 , n7976 , n7977 , n7978 , n7979 , n7980 , n7981 , n7982 , n7983 , n7984 , n7985 , n7986 , n7987 , n7988 , n7989 , n7990 , n7991 , n7992 , n7993 , n7994 , n7995 , n7996 , n7997 , n7998 , n7999 , n8000 , n8001 , n8002 , n8003 , n8004 , n8005 , n8006 , n8007 , n8008 , n8009 , n8010 , n8011 , n8012 , n8013 , n8014 , n8015 , n8016 , n8017 , n8018 , n8019 , n8020 , n8021 , n8022 , n8023 , n8024 , n8025 , n8026 , n8027 , n8028 , n8029 , n8030 , n8031 , n8032 , n8033 , n8034 , n8035 , n8036 , n8037 , n8038 , n8039 , n8040 , n8041 , n8042 , n8043 , n8044 , n8045 , n8046 , n8047 , n8048 , n8049 , n8050 , n8051 , n8052 , n8053 , n8054 , n8055 , n8056 , n8057 , n8058 , n8059 , n8060 , n8061 , n8062 , n8063 , n8064 , n8065 , n8066 , n8067 , n8068 , n8069 , n8070 , n8071 , n8072 , n8073 , n8074 , n8075 , n8076 , n8077 , n8078 , n8079 , n8080 , n8081 , n8082 , n8083 , n8084 , n8085 , n8086 , n8087 , n8088 , n8089 , n8090 , n8091 , n8092 , n8093 , n8094 , n8095 , n8096 , n8097 , n8098 , n8099 , n8100 , n8101 , n8102 , n8103 , n8104 , n8105 , n8106 , n8107 , n8108 , n8109 , n8110 , n8111 , n8112 , n8113 , n8114 , n8115 , n8116 , n8117 , n8118 , n8119 , n8120 , n8121 , n8122 , n8123 , n8124 , n8125 , n8126 , n8127 , n8128 , n8129 , n8130 , n8131 , n8132 , n8133 , n8134 , n8135 , n8136 , n8137 , n8138 , n8139 , n8140 , n8141 , n8142 , n8143 , n8144 , n8145 , n8146 , n8147 , n8148 , n8149 , n8150 , n8151 , n8152 , n8153 , n8154 , n8155 , n8156 , n8157 , n8158 , n8159 , n8160 , n8161 , n8162 , n8163 , n8164 , n8165 , n8166 , n8167 , n8168 , n8169 , n8170 , n8171 , n8172 , n8173 , n8174 , n8175 , n8176 , n8177 , n8178 , n8179 , n8180 , n8181 , n8182 , n8183 , n8184 , n8185 , n8186 , n8187 , n8188 , n8189 , n8190 , n8191 , n8192 , n8193 , n8194 , n8195 , n8196 , n8197 , n8198 , n8199 , n8200 , n8201 , n8202 , n8203 , n8204 , n8205 , n8206 , n8207 , n8208 , n8209 , n8210 , n8211 , n8212 , n8213 , n8214 , n8215 , n8216 , n8217 , n8218 , n8219 , n8220 , n8221 , n8222 , n8223 , n8224 , n8225 , n8226 , n8227 , n8228 , n8229 , n8230 , n8231 , n8232 , n8233 , n8234 , n8235 , n8236 , n8237 , n8238 , n8239 , n8240 , n8241 , n8242 , n8243 , n8244 , n8245 , n8246 , n8247 , n8248 , n8249 , n8250 , n8251 , n8252 , n8253 , n8254 , n8255 , n8256 , n8257 , n8258 , n8259 , n8260 , n8261 , n8262 , n8263 , n8264 , n8265 , n8266 , n8267 , n8268 , n8269 , n8270 , n8271 , n8272 , n8273 , n8274 , n8275 , n8276 , n8277 , n8278 , n8279 , n8280 , n8281 , n8282 , n8283 , n8284 , n8285 , n8286 , n8287 , n8288 , n8289 , n8290 , n8291 , n8292 , n8293 , n8294 , n8295 , n8296 , n8297 , n8298 , n8299 , n8300 , n8301 , n8302 , n8303 , n8304 , n8305 , n8306 , n8307 , n8308 , n8309 , n8310 , n8311 , n8312 , n8313 , n8314 , n8315 , n8316 , n8317 , n8318 , n8319 , n8320 , n8321 , n8322 , n8323 , n8324 , n8325 , n8326 , n8327 , n8328 , n8329 , n8330 , n8331 , n8332 , n8333 , n8334 , n8335 , n8336 , n8337 , n8338 , n8339 , n8340 , n8341 , n8342 , n8343 , n8344 , n8345 , n8346 , n8347 , n8348 , n8349 , n8350 , n8351 , n8352 , n8353 , n8354 , n8355 , n8356 , n8357 , n8358 , n8359 , n8360 , n8361 , n8362 , n8363 , n8364 , n8365 , n8366 , n8367 , n8368 , n8369 , n8370 , n8371 , n8372 , n8373 , n8374 , n8375 , n8376 , n8377 , n8378 , n8379 , n8380 , n8381 , n8382 , n8383 , n8384 , n8385 , n8386 , n8387 , n8388 , n8389 , n8390 , n8391 , n8392 , n8393 , n8394 , n8395 , n8396 , n8397 , n8398 , n8399 , n8400 , n8401 , n8402 , n8403 , n8404 , n8405 , n8406 , n8407 , n8408 , n8409 , n8410 , n8411 , n8412 , n8413 , n8414 , n8415 , n8416 , n8417 , n8418 , n8419 , n8420 , n8421 , n8422 , n8423 , n8424 , n8425 , n8426 , n8427 , n8428 , n8429 , n8430 , n8431 , n8432 , n8433 , n8434 , n8435 , n8436 , n8437 , n8438 , n8439 , n8440 , n8441 , n8442 , n8443 , n8444 , n8445 , n8446 , n8447 , n8448 , n8449 , n8450 , n8451 , n8452 , n8453 , n8454 , n8455 , n8456 , n8457 , n8458 , n8459 , n8460 , n8461 , n8462 , n8463 , n8464 , n8465 , n8466 , n8467 , n8468 , n8469 , n8470 , n8471 , n8472 , n8473 , n8474 , n8475 , n8476 , n8477 , n8478 , n8479 , n8480 , n8481 , n8482 , n8483 , n8484 , n8485 , n8486 , n8487 , n8488 , n8489 , n8490 , n8491 , n8492 , n8493 , n8494 , n8495 , n8496 , n8497 , n8498 , n8499 , n8500 , n8501 , n8502 , n8503 , n8504 , n8505 , n8506 , n8507 , n8508 , n8509 , n8510 , n8511 , n8512 , n8513 , n8514 , n8515 , n8516 , n8517 , n8518 , n8519 , n8520 , n8521 , n8522 , n8523 , n8524 , n8525 , n8526 , n8527 , n8528 , n8529 , n8530 , n8531 , n8532 , n8533 , n8534 , n8535 , n8536 , n8537 , n8538 , n8539 , n8540 , n8541 , n8542 , n8543 , n8544 , n8545 , n8546 , n8547 , n8548 , n8549 , n8550 , n8551 , n8552 , n8553 , n8554 , n8555 , n8556 , n8557 , n8558 , n8559 , n8560 , n8561 , n8562 , n8563 , n8564 , n8565 , n8566 , n8567 , n8568 , n8569 , n8570 , n8571 , n8572 , n8573 , n8574 , n8575 , n8576 , n8577 , n8578 , n8579 , n8580 , n8581 , n8582 , n8583 , n8584 , n8585 , n8586 , n8587 , n8588 , n8589 , n8590 , n8591 , n8592 , n8593 , n8594 , n8595 , n8596 , n8597 , n8598 , n8599 , n8600 , n8601 , n8602 , n8603 , n8604 , n8605 , n8606 , n8607 , n8608 , n8609 , n8610 , n8611 , n8612 , n8613 , n8614 , n8615 , n8616 , n8617 , n8618 , n8619 , n8620 , n8621 , n8622 , n8623 , n8624 , n8625 , n8626 , n8627 , n8628 , n8629 , n8630 , n8631 , n8632 , n8633 , n8634 , n8635 , n8636 , n8637 , n8638 , n8639 , n8640 , n8641 , n8642 , n8643 , n8644 , n8645 , n8646 , n8647 , n8648 , n8649 , n8650 , n8651 , n8652 , n8653 , n8654 , n8655 , n8656 , n8657 , n8658 , n8659 , n8660 , n8661 , n8662 , n8663 , n8664 , n8665 , n8666 , n8667 , n8668 , n8669 , n8670 , n8671 , n8672 , n8673 , n8674 , n8675 , n8676 , n8677 , n8678 , n8679 , n8680 , n8681 , n8682 , n8683 , n8684 , n8685 , n8686 , n8687 , n8688 , n8689 , n8690 , n8691 , n8692 , n8693 , n8694 , n8695 , n8696 , n8697 , n8698 , n8699 , n8700 , n8701 , n8702 , n8703 , n8704 , n8705 , n8706 , n8707 , n8708 , n8709 , n8710 , n8711 , n8712 , n8713 , n8714 , n8715 , n8716 , n8717 , n8718 , n8719 , n8720 , n8721 , n8722 , n8723 , n8724 , n8725 , n8726 , n8727 , n8728 , n8729 , n8730 , n8731 , n8732 , n8733 , n8734 , n8735 , n8736 , n8737 , n8738 , n8739 , n8740 , n8741 , n8742 , n8743 , n8744 , n8745 , n8746 , n8747 , n8748 , n8749 , n8750 , n8751 , n8752 , n8753 , n8754 , n8755 , n8756 , n8757 , n8758 , n8759 , n8760 , n8761 , n8762 , n8763 , n8764 , n8765 , n8766 , n8767 , n8768 , n8769 , n8770 , n8771 , n8772 , n8773 , n8774 , n8775 , n8776 , n8777 , n8778 , n8779 , n8780 , n8781 , n8782 , n8783 , n8784 , n8785 , n8786 , n8787 , n8788 , n8789 , n8790 , n8791 , n8792 , n8793 , n8794 , n8795 , n8796 , n8797 , n8798 , n8799 , n8800 , n8801 , n8802 , n8803 , n8804 , n8805 , n8806 , n8807 , n8808 , n8809 , n8810 , n8811 , n8812 , n8813 , n8814 , n8815 , n8816 , n8817 , n8818 , n8819 , n8820 , n8821 , n8822 , n8823 , n8824 , n8825 , n8826 , n8827 , n8828 , n8829 , n8830 , n8831 , n8832 , n8833 , n8834 , n8835 , n8836 , n8837 , n8838 , n8839 , n8840 , n8841 , n8842 , n8843 , n8844 , n8845 , n8846 , n8847 , n8848 , n8849 , n8850 , n8851 , n8852 , n8853 , n8854 , n8855 , n8856 , n8857 , n8858 , n8859 , n8860 , n8861 , n8862 , n8863 , n8864 , n8865 , n8866 , n8867 , n8868 , n8869 , n8870 , n8871 , n8872 , n8873 , n8874 , n8875 , n8876 , n8877 , n8878 , n8879 , n8880 , n8881 , n8882 , n8883 , n8884 , n8885 , n8886 , n8887 , n8888 , n8889 , n8890 , n8891 , n8892 , n8893 , n8894 , n8895 , n8896 , n8897 , n8898 , n8899 , n8900 , n8901 , n8902 , n8903 , n8904 , n8905 , n8906 , n8907 , n8908 , n8909 , n8910 , n8911 , n8912 , n8913 , n8914 , n8915 , n8916 , n8917 , n8918 , n8919 , n8920 , n8921 , n8922 , n8923 , n8924 , n8925 , n8926 , n8927 , n8928 , n8929 , n8930 , n8931 , n8932 , n8933 , n8934 , n8935 , n8936 , n8937 , n8938 , n8939 , n8940 , n8941 , n8942 , n8943 , n8944 , n8945 , n8946 , n8947 , n8948 , n8949 , n8950 , n8951 , n8952 , n8953 , n8954 , n8955 , n8956 , n8957 , n8958 , n8959 , n8960 , n8961 , n8962 , n8963 , n8964 , n8965 , n8966 , n8967 , n8968 , n8969 , n8970 , n8971 , n8972 , n8973 , n8974 , n8975 , n8976 , n8977 , n8978 , n8979 , n8980 , n8981 , n8982 , n8983 , n8984 , n8985 , n8986 , n8987 , n8988 , n8989 , n8990 , n8991 , n8992 , n8993 , n8994 , n8995 , n8996 , n8997 , n8998 , n8999 , n9000 , n9001 , n9002 , n9003 , n9004 , n9005 , n9006 , n9007 , n9008 , n9009 , n9010 , n9011 , n9012 , n9013 , n9014 , n9015 , n9016 , n9017 , n9018 , n9019 , n9020 , n9021 , n9022 , n9023 , n9024 , n9025 , n9026 , n9027 , n9028 , n9029 , n9030 , n9031 , n9032 , n9033 , n9034 , n9035 , n9036 , n9037 , n9038 , n9039 , n9040 , n9041 , n9042 , n9043 , n9044 , n9045 , n9046 , n9047 , n9048 , n9049 , n9050 , n9051 , n9052 , n9053 , n9054 , n9055 , n9056 , n9057 , n9058 , n9059 , n9060 , n9061 , n9062 , n9063 , n9064 , n9065 , n9066 , n9067 , n9068 , n9069 , n9070 , n9071 , n9072 , n9073 , n9074 , n9075 , n9076 , n9077 , n9078 , n9079 , n9080 , n9081 , n9082 , n9083 , n9084 , n9085 , n9086 , n9087 , n9088 , n9089 , n9090 , n9091 , n9092 , n9093 , n9094 , n9095 , n9096 , n9097 , n9098 , n9099 , n9100 , n9101 , n9102 , n9103 , n9104 , n9105 , n9106 , n9107 , n9108 , n9109 , n9110 , n9111 , n9112 , n9113 , n9114 , n9115 , n9116 , n9117 , n9118 , n9119 , n9120 , n9121 , n9122 , n9123 , n9124 , n9125 , n9126 , n9127 , n9128 , n9129 , n9130 , n9131 , n9132 , n9133 , n9134 , n9135 , n9136 , n9137 , n9138 , n9139 , n9140 , n9141 , n9142 , n9143 , n9144 , n9145 , n9146 , n9147 , n9148 , n9149 , n9150 , n9151 , n9152 , n9153 , n9154 , n9155 , n9156 , n9157 , n9158 , n9159 , n9160 , n9161 , n9162 , n9163 , n9164 , n9165 , n9166 , n9167 , n9168 , n9169 , n9170 , n9171 , n9172 , n9173 , n9174 , n9175 , n9176 , n9177 , n9178 , n9179 , n9180 , n9181 , n9182 , n9183 , n9184 , n9185 , n9186 , n9187 , n9188 , n9189 , n9190 , n9191 , n9192 , n9193 , n9194 , n9195 , n9196 , n9197 , n9198 , n9199 , n9200 , n9201 , n9202 , n9203 , n9204 , n9205 , n9206 , n9207 , n9208 , n9209 , n9210 , n9211 , n9212 , n9213 , n9214 , n9215 , n9216 , n9217 , n9218 , n9219 , n9220 , n9221 , n9222 , n9223 , n9224 , n9225 , n9226 , n9227 , n9228 , n9229 , n9230 , n9231 , n9232 , n9233 , n9234 , n9235 , n9236 , n9237 , n9238 , n9239 , n9240 , n9241 , n9242 , n9243 , n9244 , n9245 , n9246 , n9247 , n9248 , n9249 , n9250 , n9251 , n9252 , n9253 , n9254 , n9255 , n9256 , n9257 , n9258 , n9259 , n9260 , n9261 , n9262 , n9263 , n9264 , n9265 , n9266 , n9267 , n9268 , n9269 , n9270 , n9271 , n9272 , n9273 , n9274 , n9275 , n9276 , n9277 , n9278 , n9279 , n9280 , n9281 , n9282 , n9283 , n9284 , n9285 , n9286 , n9287 , n9288 , n9289 , n9290 , n9291 , n9292 , n9293 , n9294 , n9295 , n9296 , n9297 , n9298 , n9299 , n9300 , n9301 , n9302 , n9303 , n9304 , n9305 , n9306 , n9307 , n9308 , n9309 , n9310 , n9311 , n9312 , n9313 , n9314 , n9315 , n9316 , n9317 , n9318 , n9319 , n9320 , n9321 , n9322 , n9323 , n9324 , n9325 , n9326 , n9327 , n9328 , n9329 , n9330 , n9331 , n9332 , n9333 , n9334 , n9335 , n9336 , n9337 , n9338 , n9339 , n9340 , n9341 , n9342 , n9343 , n9344 , n9345 , n9346 , n9347 , n9348 , n9349 , n9350 , n9351 , n9352 , n9353 , n9354 , n9355 , n9356 , n9357 , n9358 , n9359 , n9360 , n9361 , n9362 , n9363 , n9364 , n9365 , n9366 , n9367 , n9368 , n9369 , n9370 , n9371 , n9372 , n9373 , n9374 , n9375 , n9376 , n9377 , n9378 , n9379 , n9380 , n9381 , n9382 , n9383 , n9384 , n9385 , n9386 , n9387 , n9388 , n9389 , n9390 , n9391 , n9392 , n9393 , n9394 , n9395 , n9396 , n9397 , n9398 , n9399 , n9400 , n9401 , n9402 , n9403 , n9404 , n9405 , n9406 , n9407 , n9408 , n9409 , n9410 , n9411 , n9412 , n9413 , n9414 , n9415 , n9416 , n9417 , n9418 , n9419 , n9420 , n9421 , n9422 , n9423 , n9424 , n9425 , n9426 , n9427 , n9428 , n9429 , n9430 , n9431 , n9432 , n9433 , n9434 , n9435 , n9436 , n9437 , n9438 , n9439 , n9440 , n9441 , n9442 , n9443 , n9444 , n9445 , n9446 , n9447 , n9448 , n9449 , n9450 , n9451 , n9452 , n9453 , n9454 , n9455 , n9456 , n9457 , n9458 , n9459 , n9460 , n9461 , n9462 , n9463 , n9464 , n9465 , n9466 , n9467 , n9468 , n9469 , n9470 , n9471 , n9472 , n9473 , n9474 , n9475 , n9476 , n9477 , n9478 , n9479 , n9480 , n9481 , n9482 , n9483 , n9484 , n9485 , n9486 , n9487 , n9488 , n9489 , n9490 , n9491 , n9492 , n9493 , n9494 , n9495 , n9496 , n9497 , n9498 , n9499 , n9500 , n9501 , n9502 , n9503 , n9504 , n9505 , n9506 , n9507 , n9508 , n9509 , n9510 , n9511 , n9512 , n9513 , n9514 , n9515 , n9516 , n9517 , n9518 , n9519 , n9520 , n9521 , n9522 , n9523 , n9524 , n9525 , n9526 , n9527 , n9528 , n9529 , n9530 , n9531 , n9532 , n9533 , n9534 , n9535 , n9536 , n9537 , n9538 , n9539 , n9540 , n9541 , n9542 , n9543 , n9544 , n9545 , n9546 , n9547 , n9548 , n9549 , n9550 , n9551 , n9552 , n9553 , n9554 , n9555 , n9556 , n9557 , n9558 , n9559 , n9560 , n9561 , n9562 , n9563 , n9564 , n9565 , n9566 , n9567 , n9568 , n9569 , n9570 , n9571 , n9572 , n9573 , n9574 , n9575 , n9576 , n9577 , n9578 , n9579 , n9580 , n9581 , n9582 , n9583 , n9584 , n9585 , n9586 , n9587 , n9588 , n9589 , n9590 , n9591 , n9592 , n9593 , n9594 , n9595 , n9596 , n9597 , n9598 , n9599 , n9600 , n9601 , n9602 , n9603 , n9604 , n9605 , n9606 , n9607 , n9608 , n9609 , n9610 , n9611 , n9612 , n9613 , n9614 , n9615 , n9616 , n9617 , n9618 , n9619 , n9620 , n9621 , n9622 , n9623 , n9624 , n9625 , n9626 , n9627 , n9628 , n9629 , n9630 , n9631 , n9632 , n9633 , n9634 , n9635 , n9636 , n9637 , n9638 , n9639 , n9640 , n9641 , n9642 , n9643 , n9644 , n9645 , n9646 , n9647 , n9648 , n9649 , n9650 , n9651 , n9652 , n9653 , n9654 , n9655 , n9656 , n9657 , n9658 , n9659 , n9660 , n9661 , n9662 , n9663 , n9664 , n9665 , n9666 , n9667 , n9668 , n9669 , n9670 , n9671 , n9672 , n9673 , n9674 , n9675 , n9676 , n9677 , n9678 , n9679 , n9680 , n9681 , n9682 , n9683 , n9684 , n9685 , n9686 , n9687 , n9688 , n9689 , n9690 , n9691 , n9692 , n9693 , n9694 , n9695 , n9696 , n9697 , n9698 , n9699 , n9700 , n9701 , n9702 , n9703 , n9704 , n9705 , n9706 , n9707 , n9708 , n9709 , n9710 , n9711 , n9712 , n9713 , n9714 , n9715 , n9716 , n9717 , n9718 , n9719 , n9720 , n9721 , n9722 , n9723 , n9724 , n9725 , n9726 , n9727 , n9728 , n9729 , n9730 , n9731 , n9732 , n9733 , n9734 , n9735 , n9736 , n9737 , n9738 , n9739 , n9740 , n9741 , n9742 , n9743 , n9744 , n9745 , n9746 , n9747 , n9748 , n9749 , n9750 , n9751 , n9752 , n9753 , n9754 , n9755 , n9756 , n9757 , n9758 , n9759 , n9760 , n9761 , n9762 , n9763 , n9764 , n9765 , n9766 , n9767 , n9768 , n9769 , n9770 , n9771 , n9772 , n9773 , n9774 , n9775 , n9776 , n9777 , n9778 , n9779 , n9780 , n9781 , n9782 , n9783 , n9784 , n9785 , n9786 , n9787 , n9788 , n9789 , n9790 , n9791 , n9792 , n9793 , n9794 , n9795 , n9796 , n9797 , n9798 , n9799 , n9800 , n9801 , n9802 , n9803 , n9804 , n9805 , n9806 , n9807 , n9808 , n9809 , n9810 , n9811 , n9812 , n9813 , n9814 , n9815 , n9816 , n9817 , n9818 , n9819 , n9820 , n9821 , n9822 , n9823 , n9824 , n9825 , n9826 , n9827 , n9828 , n9829 , n9830 , n9831 , n9832 , n9833 , n9834 , n9835 , n9836 , n9837 , n9838 , n9839 , n9840 , n9841 , n9842 , n9843 , n9844 , n9845 , n9846 , n9847 , n9848 , n9849 , n9850 , n9851 , n9852 , n9853 , n9854 , n9855 , n9856 , n9857 , n9858 , n9859 , n9860 , n9861 , n9862 , n9863 , n9864 , n9865 , n9866 , n9867 , n9868 , n9869 , n9870 , n9871 , n9872 , n9873 , n9874 , n9875 , n9876 , n9877 , n9878 , n9879 , n9880 , n9881 , n9882 , n9883 , n9884 , n9885 , n9886 , n9887 , n9888 , n9889 , n9890 , n9891 , n9892 , n9893 , n9894 , n9895 , n9896 , n9897 , n9898 , n9899 , n9900 , n9901 , n9902 , n9903 , n9904 , n9905 , n9906 , n9907 , n9908 , n9909 , n9910 , n9911 , n9912 , n9913 , n9914 , n9915 , n9916 , n9917 , n9918 , n9919 , n9920 , n9921 , n9922 , n9923 , n9924 , n9925 , n9926 , n9927 , n9928 , n9929 , n9930 , n9931 , n9932 , n9933 , n9934 , n9935 , n9936 , n9937 , n9938 , n9939 , n9940 , n9941 , n9942 , n9943 , n9944 , n9945 , n9946 , n9947 , n9948 , n9949 , n9950 , n9951 , n9952 , n9953 , n9954 , n9955 , n9956 , n9957 , n9958 , n9959 , n9960 , n9961 , n9962 , n9963 , n9964 , n9965 , n9966 , n9967 , n9968 , n9969 , n9970 , n9971 , n9972 , n9973 , n9974 , n9975 , n9976 , n9977 , n9978 , n9979 , n9980 , n9981 , n9982 , n9983 , n9984 , n9985 , n9986 , n9987 , n9988 , n9989 , n9990 , n9991 , n9992 , n9993 , n9994 , n9995 , n9996 , n9997 , n9998 , n9999 , n10000 , n10001 , n10002 , n10003 , n10004 , n10005 , n10006 , n10007 , n10008 , n10009 , n10010 , n10011 , n10012 , n10013 , n10014 , n10015 , n10016 , n10017 , n10018 , n10019 , n10020 , n10021 , n10022 , n10023 , n10024 , n10025 , n10026 , n10027 , n10028 , n10029 , n10030 , n10031 , n10032 , n10033 , n10034 , n10035 , n10036 , n10037 , n10038 , n10039 , n10040 , n10041 , n10042 , n10043 , n10044 , n10045 , n10046 , n10047 , n10048 , n10049 , n10050 , n10051 , n10052 , n10053 , n10054 , n10055 , n10056 , n10057 , n10058 , n10059 , n10060 , n10061 , n10062 , n10063 , n10064 , n10065 , n10066 , n10067 , n10068 , n10069 , n10070 , n10071 , n10072 , n10073 , n10074 , n10075 , n10076 , n10077 , n10078 , n10079 , n10080 , n10081 , n10082 , n10083 , n10084 , n10085 , n10086 , n10087 , n10088 , n10089 , n10090 , n10091 , n10092 , n10093 , n10094 , n10095 , n10096 , n10097 , n10098 , n10099 , n10100 , n10101 , n10102 , n10103 , n10104 , n10105 , n10106 , n10107 , n10108 , n10109 , n10110 , n10111 , n10112 , n10113 , n10114 , n10115 , n10116 , n10117 , n10118 , n10119 , n10120 , n10121 , n10122 , n10123 , n10124 , n10125 , n10126 , n10127 , n10128 , n10129 , n10130 , n10131 , n10132 , n10133 , n10134 , n10135 , n10136 , n10137 , n10138 , n10139 , n10140 , n10141 , n10142 , n10143 , n10144 , n10145 , n10146 , n10147 , n10148 , n10149 , n10150 , n10151 , n10152 , n10153 , n10154 , n10155 , n10156 , n10157 , n10158 , n10159 , n10160 , n10161 , n10162 , n10163 , n10164 , n10165 , n10166 , n10167 , n10168 , n10169 , n10170 , n10171 , n10172 , n10173 , n10174 , n10175 , n10176 , n10177 , n10178 , n10179 , n10180 , n10181 , n10182 , n10183 , n10184 , n10185 , n10186 , n10187 , n10188 , n10189 , n10190 , n10191 , n10192 , n10193 , n10194 , n10195 , n10196 , n10197 , n10198 , n10199 , n10200 , n10201 , n10202 , n10203 , n10204 , n10205 , n10206 , n10207 , n10208 , n10209 , n10210 , n10211 , n10212 , n10213 , n10214 , n10215 , n10216 , n10217 , n10218 , n10219 , n10220 , n10221 , n10222 , n10223 , n10224 , n10225 , n10226 , n10227 , n10228 , n10229 , n10230 , n10231 , n10232 , n10233 , n10234 , n10235 , n10236 , n10237 , n10238 , n10239 , n10240 , n10241 , n10242 , n10243 , n10244 , n10245 , n10246 , n10247 , n10248 , n10249 , n10250 , n10251 , n10252 , n10253 , n10254 , n10255 , n10256 , n10257 , n10258 , n10259 , n10260 , n10261 , n10262 , n10263 , n10264 , n10265 , n10266 , n10267 , n10268 , n10269 , n10270 , n10271 , n10272 , n10273 , n10274 , n10275 , n10276 , n10277 , n10278 , n10279 , n10280 , n10281 , n10282 , n10283 , n10284 , n10285 , n10286 , n10287 , n10288 , n10289 , n10290 , n10291 , n10292 , n10293 , n10294 , n10295 , n10296 , n10297 , n10298 , n10299 , n10300 , n10301 , n10302 , n10303 , n10304 , n10305 , n10306 , n10307 , n10308 , n10309 , n10310 , n10311 , n10312 , n10313 , n10314 , n10315 , n10316 , n10317 , n10318 , n10319 , n10320 , n10321 , n10322 , n10323 , n10324 , n10325 , n10326 , n10327 , n10328 , n10329 , n10330 , n10331 , n10332 , n10333 , n10334 , n10335 , n10336 , n10337 , n10338 , n10339 , n10340 , n10341 , n10342 , n10343 , n10344 , n10345 , n10346 , n10347 , n10348 , n10349 , n10350 , n10351 , n10352 , n10353 , n10354 , n10355 , n10356 , n10357 , n10358 , n10359 , n10360 , n10361 , n10362 , n10363 , n10364 , n10365 , n10366 , n10367 , n10368 , n10369 , n10370 , n10371 , n10372 , n10373 , n10374 , n10375 , n10376 , n10377 , n10378 , n10379 , n10380 , n10381 , n10382 , n10383 , n10384 , n10385 , n10386 , n10387 , n10388 , n10389 , n10390 , n10391 , n10392 , n10393 , n10394 , n10395 , n10396 , n10397 , n10398 , n10399 , n10400 , n10401 , n10402 , n10403 , n10404 , n10405 , n10406 , n10407 , n10408 , n10409 , n10410 , n10411 , n10412 , n10413 , n10414 , n10415 , n10416 , n10417 , n10418 , n10419 , n10420 , n10421 , n10422 , n10423 , n10424 , n10425 , n10426 , n10427 , n10428 , n10429 , n10430 , n10431 , n10432 , n10433 , n10434 , n10435 , n10436 , n10437 , n10438 , n10439 , n10440 , n10441 , n10442 , n10443 , n10444 , n10445 , n10446 , n10447 , n10448 , n10449 , n10450 , n10451 , n10452 , n10453 , n10454 , n10455 , n10456 , n10457 , n10458 , n10459 , n10460 , n10461 , n10462 , n10463 , n10464 , n10465 , n10466 , n10467 , n10468 , n10469 , n10470 , n10471 , n10472 , n10473 , n10474 , n10475 , n10476 , n10477 , n10478 , n10479 , n10480 , n10481 , n10482 , n10483 , n10484 , n10485 , n10486 , n10487 , n10488 , n10489 , n10490 , n10491 , n10492 , n10493 , n10494 , n10495 , n10496 , n10497 , n10498 , n10499 , n10500 , n10501 , n10502 , n10503 , n10504 , n10505 , n10506 , n10507 , n10508 , n10509 , n10510 , n10511 , n10512 , n10513 , n10514 , n10515 , n10516 , n10517 , n10518 , n10519 , n10520 , n10521 , n10522 , n10523 , n10524 , n10525 , n10526 , n10527 , n10528 , n10529 , n10530 , n10531 , n10532 , n10533 , n10534 , n10535 , n10536 , n10537 , n10538 , n10539 , n10540 , n10541 , n10542 , n10543 , n10544 , n10545 , n10546 , n10547 , n10548 , n10549 , n10550 , n10551 , n10552 , n10553 , n10554 , n10555 , n10556 , n10557 , n10558 , n10559 , n10560 , n10561 , n10562 , n10563 , n10564 , n10565 , n10566 , n10567 , n10568 , n10569 , n10570 , n10571 , n10572 , n10573 , n10574 , n10575 , n10576 , n10577 , n10578 , n10579 , n10580 , n10581 , n10582 , n10583 , n10584 , n10585 , n10586 , n10587 , n10588 , n10589 , n10590 , n10591 , n10592 , n10593 , n10594 , n10595 , n10596 , n10597 , n10598 , n10599 , n10600 , n10601 , n10602 , n10603 , n10604 , n10605 , n10606 , n10607 , n10608 , n10609 , n10610 , n10611 , n10612 , n10613 , n10614 , n10615 , n10616 , n10617 , n10618 , n10619 , n10620 , n10621 , n10622 , n10623 , n10624 , n10625 , n10626 , n10627 , n10628 , n10629 , n10630 , n10631 , n10632 , n10633 , n10634 , n10635 , n10636 , n10637 , n10638 , n10639 , n10640 , n10641 , n10642 , n10643 , n10644 , n10645 , n10646 , n10647 , n10648 , n10649 , n10650 , n10651 , n10652 , n10653 , n10654 , n10655 , n10656 , n10657 , n10658 , n10659 , n10660 , n10661 , n10662 , n10663 , n10664 , n10665 , n10666 , n10667 , n10668 , n10669 , n10670 , n10671 , n10672 , n10673 , n10674 , n10675 , n10676 , n10677 , n10678 , n10679 , n10680 , n10681 , n10682 , n10683 , n10684 , n10685 , n10686 , n10687 , n10688 , n10689 , n10690 , n10691 , n10692 , n10693 , n10694 , n10695 , n10696 , n10697 , n10698 , n10699 , n10700 , n10701 , n10702 , n10703 , n10704 , n10705 , n10706 , n10707 , n10708 , n10709 , n10710 , n10711 , n10712 , n10713 , n10714 , n10715 , n10716 , n10717 , n10718 , n10719 , n10720 , n10721 , n10722 , n10723 , n10724 , n10725 , n10726 , n10727 , n10728 , n10729 , n10730 , n10731 , n10732 , n10733 , n10734 , n10735 , n10736 , n10737 , n10738 , n10739 , n10740 , n10741 , n10742 , n10743 , n10744 , n10745 , n10746 , n10747 , n10748 , n10749 , n10750 , n10751 , n10752 , n10753 , n10754 , n10755 , n10756 , n10757 , n10758 , n10759 , n10760 , n10761 , n10762 , n10763 , n10764 , n10765 , n10766 , n10767 , n10768 , n10769 , n10770 , n10771 , n10772 , n10773 , n10774 , n10775 , n10776 , n10777 , n10778 , n10779 , n10780 , n10781 , n10782 , n10783 , n10784 , n10785 , n10786 , n10787 , n10788 , n10789 , n10790 , n10791 , n10792 , n10793 , n10794 , n10795 , n10796 , n10797 , n10798 , n10799 , n10800 , n10801 , n10802 , n10803 , n10804 , n10805 , n10806 , n10807 , n10808 , n10809 , n10810 , n10811 , n10812 , n10813 , n10814 , n10815 , n10816 , n10817 , n10818 , n10819 , n10820 , n10821 , n10822 , n10823 , n10824 , n10825 , n10826 , n10827 , n10828 , n10829 , n10830 , n10831 , n10832 , n10833 , n10834 , n10835 , n10836 , n10837 , n10838 , n10839 , n10840 , n10841 , n10842 , n10843 , n10844 , n10845 , n10846 , n10847 , n10848 , n10849 , n10850 , n10851 , n10852 , n10853 , n10854 , n10855 , n10856 , n10857 , n10858 , n10859 , n10860 , n10861 , n10862 , n10863 , n10864 , n10865 , n10866 , n10867 , n10868 , n10869 , n10870 , n10871 , n10872 , n10873 , n10874 , n10875 , n10876 , n10877 , n10878 , n10879 , n10880 , n10881 , n10882 , n10883 , n10884 , n10885 , n10886 , n10887 , n10888 , n10889 , n10890 , n10891 , n10892 , n10893 , n10894 , n10895 , n10896 , n10897 , n10898 , n10899 , n10900 , n10901 , n10902 , n10903 , n10904 , n10905 , n10906 , n10907 , n10908 , n10909 , n10910 , n10911 , n10912 , n10913 , n10914 , n10915 , n10916 , n10917 , n10918 , n10919 , n10920 , n10921 , n10922 , n10923 , n10924 , n10925 , n10926 , n10927 , n10928 , n10929 , n10930 , n10931 , n10932 , n10933 , n10934 , n10935 , n10936 , n10937 , n10938 , n10939 , n10940 , n10941 , n10942 , n10943 , n10944 , n10945 , n10946 , n10947 , n10948 , n10949 , n10950 , n10951 , n10952 , n10953 , n10954 , n10955 , n10956 , n10957 , n10958 , n10959 , n10960 , n10961 , n10962 , n10963 , n10964 , n10965 , n10966 , n10967 , n10968 , n10969 , n10970 , n10971 , n10972 , n10973 , n10974 , n10975 , n10976 , n10977 , n10978 , n10979 , n10980 , n10981 , n10982 , n10983 , n10984 , n10985 , n10986 , n10987 , n10988 , n10989 , n10990 , n10991 , n10992 , n10993 , n10994 , n10995 , n10996 , n10997 , n10998 , n10999 , n11000 , n11001 , n11002 , n11003 , n11004 , n11005 , n11006 , n11007 , n11008 , n11009 , n11010 , n11011 , n11012 , n11013 , n11014 , n11015 , n11016 , n11017 , n11018 , n11019 , n11020 , n11021 , n11022 , n11023 , n11024 , n11025 , n11026 , n11027 , n11028 , n11029 , n11030 , n11031 , n11032 , n11033 , n11034 , n11035 , n11036 , n11037 , n11038 , n11039 , n11040 , n11041 , n11042 , n11043 , n11044 , n11045 , n11046 , n11047 , n11048 , n11049 , n11050 , n11051 , n11052 , n11053 , n11054 , n11055 , n11056 , n11057 , n11058 , n11059 , n11060 , n11061 , n11062 , n11063 , n11064 , n11065 , n11066 , n11067 , n11068 , n11069 , n11070 , n11071 , n11072 , n11073 , n11074 , n11075 , n11076 , n11077 , n11078 , n11079 , n11080 , n11081 , n11082 , n11083 , n11084 , n11085 , n11086 , n11087 , n11088 , n11089 , n11090 , n11091 , n11092 , n11093 , n11094 , n11095 , n11096 , n11097 , n11098 , n11099 , n11100 , n11101 , n11102 , n11103 , n11104 , n11105 , n11106 , n11107 , n11108 , n11109 , n11110 , n11111 , n11112 , n11113 , n11114 , n11115 , n11116 , n11117 , n11118 , n11119 , n11120 , n11121 , n11122 , n11123 , n11124 , n11125 , n11126 , n11127 , n11128 , n11129 , n11130 , n11131 , n11132 , n11133 , n11134 , n11135 , n11136 , n11137 , n11138 , n11139 , n11140 , n11141 , n11142 , n11143 , n11144 , n11145 , n11146 , n11147 , n11148 , n11149 , n11150 , n11151 , n11152 , n11153 , n11154 , n11155 , n11156 , n11157 , n11158 , n11159 , n11160 , n11161 , n11162 , n11163 , n11164 , n11165 , n11166 , n11167 , n11168 , n11169 , n11170 , n11171 , n11172 , n11173 , n11174 , n11175 , n11176 , n11177 , n11178 , n11179 , n11180 , n11181 , n11182 , n11183 , n11184 , n11185 , n11186 , n11187 , n11188 , n11189 , n11190 , n11191 , n11192 , n11193 , n11194 , n11195 , n11196 , n11197 , n11198 , n11199 , n11200 , n11201 , n11202 , n11203 , n11204 , n11205 , n11206 , n11207 , n11208 , n11209 , n11210 , n11211 , n11212 , n11213 , n11214 , n11215 , n11216 , n11217 , n11218 , n11219 , n11220 , n11221 , n11222 , n11223 , n11224 , n11225 , n11226 , n11227 , n11228 , n11229 , n11230 , n11231 , n11232 , n11233 , n11234 , n11235 , n11236 , n11237 , n11238 , n11239 , n11240 , n11241 , n11242 , n11243 , n11244 , n11245 , n11246 , n11247 , n11248 , n11249 , n11250 , n11251 , n11252 , n11253 , n11254 , n11255 , n11256 , n11257 , n11258 , n11259 , n11260 , n11261 , n11262 , n11263 , n11264 , n11265 , n11266 , n11267 , n11268 , n11269 , n11270 , n11271 , n11272 , n11273 , n11274 , n11275 , n11276 , n11277 , n11278 , n11279 , n11280 , n11281 , n11282 , n11283 , n11284 , n11285 , n11286 , n11287 , n11288 , n11289 , n11290 , n11291 , n11292 , n11293 , n11294 , n11295 , n11296 , n11297 , n11298 , n11299 , n11300 , n11301 , n11302 , n11303 , n11304 , n11305 , n11306 , n11307 , n11308 , n11309 , n11310 , n11311 , n11312 , n11313 , n11314 , n11315 , n11316 , n11317 , n11318 , n11319 , n11320 , n11321 , n11322 , n11323 , n11324 , n11325 , n11326 , n11327 , n11328 , n11329 , n11330 , n11331 , n11332 , n11333 , n11334 , n11335 , n11336 , n11337 , n11338 , n11339 , n11340 , n11341 , n11342 , n11343 , n11344 , n11345 , n11346 , n11347 , n11348 , n11349 , n11350 , n11351 , n11352 , n11353 , n11354 , n11355 , n11356 , n11357 , n11358 , n11359 , n11360 , n11361 , n11362 , n11363 , n11364 , n11365 , n11366 , n11367 , n11368 , n11369 , n11370 , n11371 , n11372 , n11373 , n11374 , n11375 , n11376 , n11377 , n11378 , n11379 , n11380 , n11381 , n11382 , n11383 , n11384 , n11385 , n11386 , n11387 , n11388 , n11389 , n11390 , n11391 , n11392 , n11393 , n11394 , n11395 , n11396 , n11397 , n11398 , n11399 , n11400 , n11401 , n11402 , n11403 , n11404 , n11405 , n11406 , n11407 , n11408 , n11409 , n11410 , n11411 , n11412 , n11413 , n11414 , n11415 , n11416 , n11417 , n11418 , n11419 , n11420 , n11421 , n11422 , n11423 , n11424 , n11425 , n11426 , n11427 , n11428 , n11429 , n11430 , n11431 , n11432 , n11433 , n11434 , n11435 , n11436 , n11437 , n11438 , n11439 , n11440 , n11441 , n11442 , n11443 , n11444 , n11445 , n11446 , n11447 , n11448 , n11449 , n11450 , n11451 , n11452 , n11453 , n11454 , n11455 , n11456 , n11457 , n11458 , n11459 , n11460 , n11461 , n11462 , n11463 , n11464 , n11465 , n11466 , n11467 , n11468 , n11469 , n11470 , n11471 , n11472 , n11473 , n11474 , n11475 , n11476 , n11477 , n11478 , n11479 , n11480 , n11481 , n11482 , n11483 , n11484 , n11485 , n11486 , n11487 , n11488 , n11489 , n11490 , n11491 , n11492 , n11493 , n11494 , n11495 , n11496 , n11497 , n11498 , n11499 , n11500 , n11501 , n11502 , n11503 , n11504 , n11505 , n11506 , n11507 , n11508 , n11509 , n11510 , n11511 , n11512 , n11513 , n11514 , n11515 , n11516 , n11517 , n11518 , n11519 , n11520 , n11521 , n11522 , n11523 , n11524 , n11525 , n11526 , n11527 , n11528 , n11529 , n11530 , n11531 , n11532 , n11533 , n11534 , n11535 , n11536 , n11537 , n11538 , n11539 , n11540 , n11541 , n11542 , n11543 , n11544 , n11545 , n11546 , n11547 , n11548 , n11549 , n11550 , n11551 , n11552 , n11553 , n11554 , n11555 , n11556 , n11557 , n11558 , n11559 , n11560 , n11561 , n11562 , n11563 , n11564 , n11565 , n11566 , n11567 , n11568 , n11569 , n11570 , n11571 , n11572 , n11573 , n11574 , n11575 , n11576 , n11577 , n11578 , n11579 , n11580 , n11581 , n11582 , n11583 , n11584 , n11585 , n11586 , n11587 , n11588 , n11589 , n11590 , n11591 , n11592 , n11593 , n11594 , n11595 , n11596 , n11597 , n11598 , n11599 , n11600 , n11601 , n11602 , n11603 , n11604 , n11605 , n11606 , n11607 , n11608 , n11609 , n11610 , n11611 , n11612 , n11613 , n11614 , n11615 , n11616 , n11617 , n11618 , n11619 , n11620 , n11621 , n11622 , n11623 , n11624 , n11625 , n11626 , n11627 , n11628 , n11629 , n11630 , n11631 , n11632 , n11633 , n11634 , n11635 , n11636 , n11637 , n11638 , n11639 , n11640 , n11641 , n11642 , n11643 , n11644 , n11645 , n11646 , n11647 , n11648 , n11649 , n11650 , n11651 , n11652 , n11653 , n11654 , n11655 , n11656 , n11657 , n11658 , n11659 , n11660 , n11661 , n11662 , n11663 , n11664 , n11665 , n11666 , n11667 , n11668 , n11669 , n11670 , n11671 , n11672 , n11673 , n11674 , n11675 , n11676 , n11677 , n11678 , n11679 , n11680 , n11681 , n11682 , n11683 , n11684 , n11685 , n11686 , n11687 , n11688 , n11689 , n11690 , n11691 , n11692 , n11693 , n11694 , n11695 , n11696 , n11697 , n11698 , n11699 , n11700 , n11701 , n11702 , n11703 , n11704 , n11705 , n11706 , n11707 , n11708 , n11709 , n11710 , n11711 , n11712 , n11713 , n11714 , n11715 , n11716 , n11717 , n11718 , n11719 , n11720 , n11721 , n11722 , n11723 , n11724 , n11725 , n11726 , n11727 , n11728 , n11729 , n11730 , n11731 , n11732 , n11733 , n11734 , n11735 , n11736 , n11737 , n11738 , n11739 , n11740 , n11741 , n11742 , n11743 , n11744 , n11745 , n11746 , n11747 , n11748 , n11749 , n11750 , n11751 , n11752 , n11753 , n11754 , n11755 , n11756 , n11757 , n11758 , n11759 , n11760 , n11761 , n11762 , n11763 , n11764 , n11765 , n11766 , n11767 , n11768 , n11769 , n11770 , n11771 , n11772 , n11773 , n11774 , n11775 , n11776 , n11777 , n11778 , n11779 , n11780 , n11781 , n11782 , n11783 , n11784 , n11785 , n11786 , n11787 , n11788 , n11789 , n11790 , n11791 , n11792 , n11793 , n11794 , n11795 , n11796 , n11797 , n11798 , n11799 , n11800 , n11801 , n11802 , n11803 , n11804 , n11805 , n11806 , n11807 , n11808 , n11809 , n11810 , n11811 , n11812 , n11813 , n11814 , n11815 , n11816 , n11817 , n11818 , n11819 , n11820 , n11821 , n11822 , n11823 , n11824 , n11825 , n11826 , n11827 , n11828 , n11829 , n11830 , n11831 , n11832 , n11833 , n11834 , n11835 , n11836 , n11837 , n11838 , n11839 , n11840 , n11841 , n11842 , n11843 , n11844 , n11845 , n11846 , n11847 , n11848 , n11849 , n11850 , n11851 , n11852 , n11853 , n11854 , n11855 , n11856 , n11857 , n11858 , n11859 , n11860 , n11861 , n11862 , n11863 , n11864 , n11865 , n11866 , n11867 , n11868 , n11869 , n11870 , n11871 , n11872 , n11873 , n11874 , n11875 , n11876 , n11877 , n11878 , n11879 , n11880 , n11881 , n11882 , n11883 , n11884 , n11885 , n11886 , n11887 , n11888 , n11889 , n11890 , n11891 , n11892 , n11893 , n11894 , n11895 , n11896 , n11897 , n11898 , n11899 , n11900 , n11901 , n11902 , n11903 , n11904 , n11905 , n11906 , n11907 , n11908 , n11909 , n11910 , n11911 , n11912 , n11913 , n11914 , n11915 , n11916 , n11917 , n11918 , n11919 , n11920 , n11921 , n11922 , n11923 , n11924 , n11925 , n11926 , n11927 , n11928 , n11929 , n11930 , n11931 , n11932 , n11933 , n11934 , n11935 , n11936 , n11937 , n11938 , n11939 , n11940 , n11941 , n11942 , n11943 , n11944 , n11945 , n11946 , n11947 , n11948 , n11949 , n11950 , n11951 , n11952 , n11953 , n11954 , n11955 , n11956 , n11957 , n11958 , n11959 , n11960 , n11961 , n11962 , n11963 , n11964 , n11965 , n11966 , n11967 , n11968 , n11969 , n11970 , n11971 , n11972 , n11973 , n11974 , n11975 , n11976 , n11977 , n11978 , n11979 , n11980 , n11981 , n11982 , n11983 , n11984 , n11985 , n11986 , n11987 , n11988 , n11989 , n11990 , n11991 , n11992 , n11993 , n11994 , n11995 , n11996 , n11997 , n11998 , n11999 , n12000 , n12001 , n12002 , n12003 , n12004 , n12005 , n12006 , n12007 , n12008 , n12009 , n12010 , n12011 , n12012 , n12013 , n12014 , n12015 , n12016 , n12017 , n12018 , n12019 , n12020 , n12021 , n12022 , n12023 , n12024 , n12025 , n12026 , n12027 , n12028 , n12029 , n12030 , n12031 , n12032 , n12033 , n12034 , n12035 , n12036 , n12037 , n12038 , n12039 , n12040 , n12041 , n12042 , n12043 , n12044 , n12045 , n12046 , n12047 , n12048 , n12049 , n12050 , n12051 , n12052 , n12053 , n12054 , n12055 , n12056 , n12057 , n12058 , n12059 , n12060 , n12061 , n12062 , n12063 , n12064 , n12065 , n12066 , n12067 , n12068 , n12069 , n12070 , n12071 , n12072 , n12073 , n12074 , n12075 , n12076 , n12077 , n12078 , n12079 , n12080 , n12081 , n12082 , n12083 , n12084 , n12085 , n12086 , n12087 , n12088 , n12089 , n12090 , n12091 , n12092 , n12093 , n12094 , n12095 , n12096 , n12097 , n12098 , n12099 , n12100 , n12101 , n12102 , n12103 , n12104 , n12105 , n12106 , n12107 , n12108 , n12109 , n12110 , n12111 , n12112 , n12113 , n12114 , n12115 , n12116 , n12117 , n12118 , n12119 , n12120 , n12121 , n12122 , n12123 , n12124 , n12125 , n12126 , n12127 , n12128 , n12129 , n12130 , n12131 , n12132 , n12133 , n12134 , n12135 , n12136 , n12137 , n12138 , n12139 , n12140 , n12141 , n12142 , n12143 , n12144 , n12145 , n12146 , n12147 , n12148 , n12149 , n12150 , n12151 , n12152 , n12153 , n12154 , n12155 , n12156 , n12157 , n12158 , n12159 , n12160 , n12161 , n12162 , n12163 , n12164 , n12165 , n12166 , n12167 , n12168 , n12169 , n12170 , n12171 , n12172 , n12173 , n12174 , n12175 , n12176 , n12177 , n12178 , n12179 , n12180 , n12181 , n12182 , n12183 , n12184 , n12185 , n12186 , n12187 , n12188 , n12189 , n12190 , n12191 , n12192 , n12193 , n12194 , n12195 , n12196 , n12197 , n12198 , n12199 , n12200 , n12201 , n12202 , n12203 , n12204 , n12205 , n12206 , n12207 , n12208 , n12209 , n12210 , n12211 , n12212 , n12213 , n12214 , n12215 , n12216 , n12217 , n12218 , n12219 , n12220 , n12221 , n12222 , n12223 , n12224 , n12225 , n12226 , n12227 , n12228 , n12229 , n12230 , n12231 , n12232 , n12233 , n12234 , n12235 , n12236 , n12237 , n12238 , n12239 , n12240 , n12241 , n12242 , n12243 , n12244 , n12245 , n12246 , n12247 , n12248 , n12249 , n12250 , n12251 , n12252 , n12253 , n12254 , n12255 , n12256 , n12257 , n12258 , n12259 , n12260 , n12261 , n12262 , n12263 , n12264 , n12265 , n12266 , n12267 , n12268 , n12269 , n12270 , n12271 , n12272 , n12273 , n12274 , n12275 , n12276 , n12277 , n12278 , n12279 , n12280 , n12281 , n12282 , n12283 , n12284 , n12285 , n12286 , n12287 , n12288 , n12289 , n12290 , n12291 , n12292 , n12293 , n12294 , n12295 , n12296 , n12297 , n12298 , n12299 , n12300 , n12301 , n12302 , n12303 , n12304 , n12305 , n12306 , n12307 , n12308 , n12309 , n12310 , n12311 , n12312 , n12313 , n12314 , n12315 , n12316 , n12317 , n12318 , n12319 , n12320 , n12321 , n12322 , n12323 , n12324 , n12325 , n12326 , n12327 , n12328 , n12329 , n12330 , n12331 , n12332 , n12333 , n12334 , n12335 , n12336 , n12337 , n12338 , n12339 , n12340 , n12341 , n12342 , n12343 , n12344 , n12345 , n12346 , n12347 , n12348 , n12349 , n12350 , n12351 , n12352 , n12353 , n12354 , n12355 , n12356 , n12357 , n12358 , n12359 , n12360 , n12361 , n12362 , n12363 , n12364 , n12365 , n12366 , n12367 , n12368 , n12369 , n12370 , n12371 , n12372 , n12373 , n12374 , n12375 , n12376 , n12377 , n12378 , n12379 , n12380 , n12381 , n12382 , n12383 , n12384 , n12385 , n12386 , n12387 , n12388 , n12389 , n12390 , n12391 , n12392 , n12393 , n12394 , n12395 , n12396 , n12397 , n12398 , n12399 , n12400 , n12401 , n12402 , n12403 , n12404 , n12405 , n12406 , n12407 , n12408 , n12409 , n12410 , n12411 , n12412 , n12413 , n12414 , n12415 , n12416 , n12417 , n12418 , n12419 , n12420 , n12421 , n12422 , n12423 , n12424 , n12425 , n12426 , n12427 , n12428 , n12429 , n12430 , n12431 , n12432 , n12433 , n12434 , n12435 , n12436 , n12437 , n12438 , n12439 , n12440 , n12441 , n12442 , n12443 , n12444 , n12445 , n12446 , n12447 , n12448 , n12449 , n12450 , n12451 , n12452 , n12453 , n12454 , n12455 , n12456 , n12457 , n12458 , n12459 , n12460 , n12461 , n12462 , n12463 , n12464 , n12465 , n12466 , n12467 , n12468 , n12469 , n12470 , n12471 , n12472 , n12473 , n12474 , n12475 , n12476 , n12477 , n12478 , n12479 , n12480 , n12481 , n12482 , n12483 , n12484 , n12485 , n12486 , n12487 , n12488 , n12489 , n12490 , n12491 , n12492 , n12493 , n12494 , n12495 , n12496 , n12497 , n12498 , n12499 , n12500 , n12501 , n12502 , n12503 , n12504 , n12505 , n12506 , n12507 , n12508 , n12509 , n12510 , n12511 , n12512 , n12513 , n12514 , n12515 , n12516 , n12517 , n12518 , n12519 , n12520 , n12521 , n12522 , n12523 , n12524 , n12525 , n12526 , n12527 , n12528 , n12529 , n12530 , n12531 , n12532 , n12533 , n12534 , n12535 , n12536 , n12537 , n12538 , n12539 , n12540 , n12541 , n12542 , n12543 , n12544 , n12545 , n12546 , n12547 , n12548 , n12549 , n12550 , n12551 , n12552 , n12553 , n12554 , n12555 , n12556 , n12557 , n12558 , n12559 , n12560 , n12561 , n12562 , n12563 , n12564 , n12565 , n12566 , n12567 , n12568 , n12569 , n12570 , n12571 , n12572 , n12573 , n12574 , n12575 , n12576 , n12577 , n12578 , n12579 , n12580 , n12581 , n12582 , n12583 , n12584 , n12585 , n12586 , n12587 , n12588 , n12589 , n12590 , n12591 , n12592 , n12593 , n12594 , n12595 , n12596 , n12597 , n12598 , n12599 , n12600 , n12601 , n12602 , n12603 , n12604 , n12605 , n12606 , n12607 , n12608 , n12609 , n12610 , n12611 , n12612 , n12613 , n12614 , n12615 , n12616 , n12617 , n12618 , n12619 , n12620 , n12621 , n12622 , n12623 , n12624 , n12625 , n12626 , n12627 , n12628 , n12629 , n12630 , n12631 , n12632 , n12633 , n12634 , n12635 , n12636 , n12637 , n12638 , n12639 , n12640 , n12641 , n12642 , n12643 , n12644 , n12645 , n12646 , n12647 , n12648 , n12649 , n12650 , n12651 , n12652 , n12653 , n12654 , n12655 , n12656 , n12657 , n12658 , n12659 , n12660 , n12661 , n12662 , n12663 , n12664 , n12665 , n12666 , n12667 , n12668 , n12669 , n12670 , n12671 , n12672 , n12673 , n12674 , n12675 , n12676 , n12677 , n12678 , n12679 , n12680 , n12681 , n12682 , n12683 , n12684 , n12685 , n12686 , n12687 , n12688 , n12689 , n12690 , n12691 , n12692 , n12693 , n12694 , n12695 , n12696 , n12697 , n12698 , n12699 , n12700 , n12701 , n12702 , n12703 , n12704 , n12705 , n12706 , n12707 , n12708 , n12709 , n12710 , n12711 , n12712 , n12713 , n12714 , n12715 , n12716 , n12717 , n12718 , n12719 , n12720 , n12721 , n12722 , n12723 , n12724 , n12725 , n12726 , n12727 , n12728 , n12729 , n12730 , n12731 , n12732 , n12733 , n12734 , n12735 , n12736 , n12737 , n12738 , n12739 , n12740 , n12741 , n12742 , n12743 , n12744 , n12745 , n12746 , n12747 , n12748 , n12749 , n12750 , n12751 , n12752 , n12753 , n12754 , n12755 , n12756 , n12757 , n12758 , n12759 , n12760 , n12761 , n12762 , n12763 , n12764 , n12765 , n12766 , n12767 , n12768 , n12769 , n12770 , n12771 , n12772 , n12773 , n12774 , n12775 , n12776 , n12777 , n12778 , n12779 , n12780 , n12781 , n12782 , n12783 , n12784 , n12785 , n12786 , n12787 , n12788 , n12789 , n12790 , n12791 , n12792 , n12793 , n12794 , n12795 , n12796 , n12797 , n12798 , n12799 , n12800 , n12801 , n12802 , n12803 , n12804 , n12805 , n12806 , n12807 , n12808 , n12809 , n12810 , n12811 , n12812 , n12813 , n12814 , n12815 , n12816 , n12817 , n12818 , n12819 , n12820 , n12821 , n12822 , n12823 , n12824 , n12825 , n12826 , n12827 , n12828 , n12829 , n12830 , n12831 , n12832 , n12833 , n12834 , n12835 , n12836 , n12837 , n12838 , n12839 , n12840 , n12841 , n12842 , n12843 , n12844 , n12845 , n12846 , n12847 , n12848 , n12849 , n12850 , n12851 , n12852 , n12853 , n12854 , n12855 , n12856 , n12857 , n12858 , n12859 , n12860 , n12861 , n12862 , n12863 , n12864 , n12865 , n12866 , n12867 , n12868 , n12869 , n12870 , n12871 , n12872 , n12873 , n12874 , n12875 , n12876 , n12877 , n12878 , n12879 , n12880 , n12881 , n12882 , n12883 , n12884 , n12885 , n12886 , n12887 , n12888 , n12889 , n12890 , n12891 , n12892 , n12893 , n12894 , n12895 , n12896 , n12897 , n12898 , n12899 , n12900 , n12901 , n12902 , n12903 , n12904 , n12905 , n12906 , n12907 , n12908 , n12909 , n12910 , n12911 , n12912 , n12913 , n12914 , n12915 , n12916 , n12917 , n12918 , n12919 , n12920 , n12921 , n12922 , n12923 , n12924 , n12925 , n12926 , n12927 , n12928 , n12929 , n12930 , n12931 , n12932 , n12933 , n12934 , n12935 , n12936 , n12937 , n12938 , n12939 , n12940 , n12941 , n12942 , n12943 , n12944 , n12945 , n12946 , n12947 , n12948 , n12949 , n12950 , n12951 , n12952 , n12953 , n12954 , n12955 , n12956 , n12957 , n12958 , n12959 , n12960 , n12961 , n12962 , n12963 , n12964 , n12965 , n12966 , n12967 , n12968 , n12969 , n12970 , n12971 , n12972 , n12973 , n12974 , n12975 , n12976 , n12977 , n12978 , n12979 , n12980 , n12981 , n12982 , n12983 , n12984 , n12985 , n12986 , n12987 , n12988 , n12989 , n12990 , n12991 , n12992 , n12993 , n12994 , n12995 , n12996 , n12997 , n12998 , n12999 , n13000 , n13001 , n13002 , n13003 , n13004 , n13005 , n13006 , n13007 , n13008 , n13009 , n13010 , n13011 , n13012 , n13013 , n13014 , n13015 , n13016 , n13017 , n13018 , n13019 , n13020 , n13021 , n13022 , n13023 , n13024 , n13025 , n13026 , n13027 , n13028 , n13029 , n13030 , n13031 , n13032 , n13033 , n13034 , n13035 , n13036 , n13037 , n13038 , n13039 , n13040 , n13041 , n13042 , n13043 , n13044 , n13045 , n13046 , n13047 , n13048 , n13049 , n13050 , n13051 , n13052 , n13053 , n13054 , n13055 , n13056 , n13057 , n13058 , n13059 , n13060 , n13061 , n13062 , n13063 , n13064 , n13065 , n13066 , n13067 , n13068 , n13069 , n13070 , n13071 , n13072 , n13073 , n13074 , n13075 , n13076 , n13077 , n13078 , n13079 , n13080 , n13081 , n13082 , n13083 , n13084 , n13085 , n13086 , n13087 , n13088 , n13089 , n13090 , n13091 , n13092 , n13093 , n13094 , n13095 , n13096 , n13097 , n13098 , n13099 , n13100 , n13101 , n13102 , n13103 , n13104 , n13105 , n13106 , n13107 , n13108 , n13109 , n13110 , n13111 , n13112 , n13113 , n13114 , n13115 , n13116 , n13117 , n13118 , n13119 , n13120 , n13121 , n13122 , n13123 , n13124 , n13125 , n13126 , n13127 , n13128 , n13129 , n13130 , n13131 , n13132 , n13133 , n13134 , n13135 , n13136 , n13137 , n13138 , n13139 , n13140 , n13141 , n13142 , n13143 , n13144 , n13145 , n13146 , n13147 , n13148 , n13149 , n13150 , n13151 , n13152 , n13153 , n13154 , n13155 , n13156 , n13157 , n13158 , n13159 , n13160 , n13161 , n13162 , n13163 , n13164 , n13165 , n13166 , n13167 , n13168 , n13169 , n13170 , n13171 , n13172 , n13173 , n13174 , n13175 , n13176 , n13177 , n13178 , n13179 , n13180 , n13181 , n13182 , n13183 , n13184 , n13185 , n13186 , n13187 , n13188 , n13189 , n13190 , n13191 , n13192 , n13193 , n13194 , n13195 , n13196 , n13197 , n13198 , n13199 , n13200 , n13201 , n13202 , n13203 , n13204 , n13205 , n13206 , n13207 , n13208 , n13209 , n13210 , n13211 , n13212 , n13213 , n13214 , n13215 , n13216 , n13217 , n13218 , n13219 , n13220 , n13221 , n13222 , n13223 , n13224 , n13225 , n13226 , n13227 , n13228 , n13229 , n13230 , n13231 , n13232 , n13233 , n13234 , n13235 , n13236 , n13237 , n13238 , n13239 , n13240 , n13241 , n13242 , n13243 , n13244 , n13245 , n13246 , n13247 , n13248 , n13249 , n13250 , n13251 , n13252 , n13253 , n13254 , n13255 , n13256 , n13257 , n13258 , n13259 , n13260 , n13261 , n13262 , n13263 , n13264 , n13265 , n13266 , n13267 , n13268 , n13269 , n13270 , n13271 , n13272 , n13273 , n13274 , n13275 , n13276 , n13277 , n13278 , n13279 , n13280 , n13281 , n13282 , n13283 , n13284 , n13285 , n13286 , n13287 , n13288 , n13289 , n13290 , n13291 , n13292 , n13293 , n13294 , n13295 , n13296 , n13297 , n13298 , n13299 , n13300 , n13301 , n13302 , n13303 , n13304 , n13305 , n13306 , n13307 , n13308 , n13309 , n13310 , n13311 , n13312 , n13313 , n13314 , n13315 , n13316 , n13317 , n13318 , n13319 , n13320 , n13321 , n13322 , n13323 , n13324 , n13325 , n13326 , n13327 , n13328 , n13329 , n13330 , n13331 , n13332 , n13333 , n13334 , n13335 , n13336 , n13337 , n13338 , n13339 , n13340 , n13341 , n13342 , n13343 , n13344 , n13345 , n13346 , n13347 , n13348 , n13349 , n13350 , n13351 , n13352 , n13353 , n13354 , n13355 , n13356 , n13357 , n13358 , n13359 , n13360 , n13361 , n13362 , n13363 , n13364 , n13365 , n13366 , n13367 , n13368 , n13369 , n13370 , n13371 , n13372 , n13373 , n13374 , n13375 , n13376 , n13377 , n13378 , n13379 , n13380 , n13381 , n13382 , n13383 , n13384 , n13385 , n13386 , n13387 , n13388 , n13389 , n13390 , n13391 , n13392 , n13393 , n13394 , n13395 , n13396 , n13397 , n13398 , n13399 , n13400 , n13401 , n13402 , n13403 , n13404 , n13405 , n13406 , n13407 , n13408 , n13409 , n13410 , n13411 , n13412 , n13413 , n13414 , n13415 , n13416 , n13417 , n13418 , n13419 , n13420 , n13421 , n13422 , n13423 , n13424 , n13425 , n13426 , n13427 , n13428 , n13429 , n13430 , n13431 , n13432 , n13433 , n13434 , n13435 , n13436 , n13437 , n13438 , n13439 , n13440 , n13441 , n13442 , n13443 , n13444 , n13445 , n13446 , n13447 , n13448 , n13449 , n13450 , n13451 , n13452 , n13453 , n13454 , n13455 , n13456 , n13457 , n13458 , n13459 , n13460 , n13461 , n13462 , n13463 , n13464 , n13465 , n13466 , n13467 , n13468 , n13469 , n13470 , n13471 , n13472 , n13473 , n13474 , n13475 , n13476 , n13477 , n13478 , n13479 , n13480 , n13481 , n13482 , n13483 , n13484 , n13485 , n13486 , n13487 , n13488 , n13489 , n13490 , n13491 , n13492 , n13493 , n13494 , n13495 , n13496 , n13497 , n13498 , n13499 , n13500 , n13501 , n13502 , n13503 , n13504 , n13505 , n13506 , n13507 , n13508 , n13509 , n13510 , n13511 , n13512 , n13513 , n13514 , n13515 , n13516 , n13517 , n13518 , n13519 , n13520 , n13521 , n13522 , n13523 , n13524 , n13525 , n13526 , n13527 , n13528 , n13529 , n13530 , n13531 , n13532 , n13533 , n13534 , n13535 , n13536 , n13537 , n13538 , n13539 , n13540 , n13541 , n13542 , n13543 , n13544 , n13545 , n13546 , n13547 , n13548 , n13549 , n13550 , n13551 , n13552 , n13553 , n13554 , n13555 , n13556 , n13557 , n13558 , n13559 , n13560 , n13561 , n13562 , n13563 , n13564 , n13565 , n13566 , n13567 , n13568 , n13569 , n13570 , n13571 , n13572 , n13573 , n13574 , n13575 , n13576 , n13577 , n13578 , n13579 , n13580 , n13581 , n13582 , n13583 , n13584 , n13585 , n13586 , n13587 , n13588 , n13589 , n13590 , n13591 , n13592 , n13593 , n13594 , n13595 , n13596 , n13597 , n13598 , n13599 , n13600 , n13601 , n13602 , n13603 , n13604 , n13605 , n13606 , n13607 , n13608 , n13609 , n13610 , n13611 , n13612 , n13613 , n13614 , n13615 , n13616 , n13617 , n13618 , n13619 , n13620 , n13621 , n13622 , n13623 , n13624 , n13625 , n13626 , n13627 , n13628 , n13629 , n13630 , n13631 , n13632 , n13633 , n13634 , n13635 , n13636 , n13637 , n13638 , n13639 , n13640 , n13641 , n13642 , n13643 , n13644 , n13645 , n13646 , n13647 , n13648 , n13649 , n13650 , n13651 , n13652 , n13653 , n13654 , n13655 , n13656 , n13657 , n13658 , n13659 , n13660 , n13661 , n13662 , n13663 , n13664 , n13665 , n13666 , n13667 , n13668 , n13669 , n13670 , n13671 , n13672 , n13673 , n13674 , n13675 , n13676 , n13677 , n13678 , n13679 , n13680 , n13681 , n13682 , n13683 , n13684 , n13685 , n13686 , n13687 , n13688 , n13689 , n13690 , n13691 , n13692 , n13693 , n13694 , n13695 , n13696 , n13697 , n13698 , n13699 , n13700 , n13701 , n13702 , n13703 , n13704 , n13705 , n13706 , n13707 , n13708 , n13709 , n13710 , n13711 , n13712 , n13713 , n13714 , n13715 , n13716 , n13717 , n13718 , n13719 , n13720 , n13721 , n13722 , n13723 , n13724 , n13725 , n13726 , n13727 , n13728 , n13729 , n13730 , n13731 , n13732 , n13733 , n13734 , n13735 , n13736 , n13737 , n13738 , n13739 , n13740 , n13741 , n13742 , n13743 , n13744 , n13745 , n13746 , n13747 , n13748 , n13749 , n13750 , n13751 , n13752 , n13753 , n13754 , n13755 , n13756 , n13757 , n13758 , n13759 , n13760 , n13761 , n13762 , n13763 , n13764 , n13765 , n13766 , n13767 , n13768 , n13769 , n13770 , n13771 , n13772 , n13773 , n13774 , n13775 , n13776 , n13777 , n13778 , n13779 , n13780 , n13781 , n13782 , n13783 , n13784 , n13785 , n13786 , n13787 , n13788 , n13789 , n13790 , n13791 , n13792 , n13793 , n13794 , n13795 , n13796 , n13797 , n13798 , n13799 , n13800 , n13801 , n13802 , n13803 , n13804 , n13805 , n13806 , n13807 , n13808 , n13809 , n13810 , n13811 , n13812 , n13813 , n13814 , n13815 , n13816 , n13817 , n13818 , n13819 , n13820 , n13821 , n13822 , n13823 , n13824 , n13825 , n13826 , n13827 , n13828 , n13829 , n13830 , n13831 , n13832 , n13833 , n13834 , n13835 , n13836 , n13837 , n13838 , n13839 , n13840 , n13841 , n13842 , n13843 , n13844 , n13845 , n13846 , n13847 , n13848 , n13849 , n13850 , n13851 , n13852 , n13853 , n13854 , n13855 , n13856 , n13857 , n13858 , n13859 , n13860 , n13861 , n13862 , n13863 , n13864 , n13865 , n13866 , n13867 , n13868 , n13869 , n13870 , n13871 , n13872 , n13873 , n13874 , n13875 , n13876 , n13877 , n13878 , n13879 , n13880 , n13881 , n13882 , n13883 , n13884 , n13885 , n13886 , n13887 , n13888 , n13889 , n13890 , n13891 , n13892 , n13893 , n13894 , n13895 , n13896 , n13897 , n13898 , n13899 , n13900 , n13901 , n13902 , n13903 , n13904 , n13905 , n13906 , n13907 , n13908 , n13909 , n13910 , n13911 , n13912 , n13913 , n13914 , n13915 , n13916 , n13917 , n13918 , n13919 , n13920 , n13921 , n13922 , n13923 , n13924 , n13925 , n13926 , n13927 , n13928 , n13929 , n13930 , n13931 , n13932 , n13933 , n13934 , n13935 , n13936 , n13937 , n13938 , n13939 , n13940 , n13941 , n13942 , n13943 , n13944 , n13945 , n13946 , n13947 , n13948 , n13949 , n13950 , n13951 , n13952 , n13953 , n13954 , n13955 , n13956 , n13957 , n13958 , n13959 , n13960 , n13961 , n13962 , n13963 , n13964 , n13965 , n13966 , n13967 , n13968 , n13969 , n13970 , n13971 , n13972 , n13973 , n13974 , n13975 , n13976 , n13977 , n13978 , n13979 , n13980 , n13981 , n13982 , n13983 , n13984 , n13985 , n13986 , n13987 , n13988 , n13989 , n13990 , n13991 , n13992 , n13993 , n13994 , n13995 , n13996 , n13997 , n13998 , n13999 , n14000 , n14001 , n14002 , n14003 , n14004 , n14005 , n14006 , n14007 , n14008 , n14009 , n14010 , n14011 , n14012 , n14013 , n14014 , n14015 , n14016 , n14017 , n14018 , n14019 , n14020 , n14021 , n14022 , n14023 , n14024 , n14025 , n14026 , n14027 , n14028 , n14029 , n14030 , n14031 , n14032 , n14033 , n14034 , n14035 , n14036 , n14037 , n14038 , n14039 , n14040 , n14041 , n14042 , n14043 , n14044 , n14045 , n14046 , n14047 , n14048 , n14049 , n14050 , n14051 , n14052 , n14053 , n14054 , n14055 , n14056 , n14057 , n14058 , n14059 , n14060 , n14061 , n14062 , n14063 , n14064 , n14065 , n14066 , n14067 , n14068 , n14069 , n14070 , n14071 , n14072 , n14073 , n14074 , n14075 , n14076 , n14077 , n14078 , n14079 , n14080 , n14081 , n14082 , n14083 , n14084 , n14085 , n14086 , n14087 , n14088 , n14089 , n14090 , n14091 , n14092 , n14093 , n14094 , n14095 , n14096 , n14097 , n14098 , n14099 , n14100 , n14101 , n14102 , n14103 , n14104 , n14105 , n14106 , n14107 , n14108 , n14109 , n14110 , n14111 , n14112 , n14113 , n14114 , n14115 , n14116 , n14117 , n14118 , n14119 , n14120 , n14121 , n14122 , n14123 , n14124 , n14125 , n14126 , n14127 , n14128 , n14129 , n14130 , n14131 , n14132 , n14133 , n14134 , n14135 , n14136 , n14137 , n14138 , n14139 , n14140 , n14141 , n14142 , n14143 , n14144 , n14145 , n14146 , n14147 , n14148 , n14149 , n14150 , n14151 , n14152 , n14153 , n14154 , n14155 , n14156 , n14157 , n14158 , n14159 , n14160 , n14161 , n14162 , n14163 , n14164 , n14165 , n14166 , n14167 , n14168 , n14169 , n14170 , n14171 , n14172 , n14173 , n14174 , n14175 , n14176 , n14177 , n14178 , n14179 , n14180 , n14181 , n14182 , n14183 , n14184 , n14185 , n14186 , n14187 , n14188 , n14189 , n14190 , n14191 , n14192 , n14193 , n14194 , n14195 , n14196 , n14197 , n14198 , n14199 , n14200 , n14201 , n14202 , n14203 , n14204 , n14205 , n14206 , n14207 , n14208 , n14209 , n14210 , n14211 , n14212 , n14213 , n14214 , n14215 , n14216 , n14217 , n14218 , n14219 , n14220 , n14221 , n14222 , n14223 , n14224 , n14225 , n14226 , n14227 , n14228 , n14229 , n14230 , n14231 , n14232 , n14233 , n14234 , n14235 , n14236 , n14237 , n14238 , n14239 , n14240 , n14241 , n14242 , n14243 , n14244 , n14245 , n14246 , n14247 , n14248 , n14249 , n14250 , n14251 , n14252 , n14253 , n14254 , n14255 , n14256 , n14257 , n14258 , n14259 , n14260 , n14261 , n14262 , n14263 , n14264 , n14265 , n14266 , n14267 , n14268 , n14269 , n14270 , n14271 , n14272 , n14273 , n14274 , n14275 , n14276 , n14277 , n14278 , n14279 , n14280 , n14281 , n14282 , n14283 , n14284 , n14285 , n14286 , n14287 , n14288 , n14289 , n14290 , n14291 , n14292 , n14293 , n14294 , n14295 , n14296 , n14297 , n14298 , n14299 , n14300 , n14301 , n14302 , n14303 , n14304 , n14305 , n14306 , n14307 , n14308 , n14309 , n14310 , n14311 , n14312 , n14313 , n14314 , n14315 , n14316 , n14317 , n14318 , n14319 , n14320 , n14321 , n14322 , n14323 , n14324 , n14325 , n14326 , n14327 , n14328 , n14329 , n14330 , n14331 , n14332 , n14333 , n14334 , n14335 , n14336 , n14337 , n14338 , n14339 , n14340 , n14341 , n14342 , n14343 , n14344 , n14345 , n14346 , n14347 , n14348 , n14349 , n14350 , n14351 , n14352 , n14353 , n14354 , n14355 , n14356 , n14357 , n14358 , n14359 , n14360 , n14361 , n14362 , n14363 , n14364 , n14365 , n14366 , n14367 , n14368 , n14369 , n14370 , n14371 , n14372 , n14373 , n14374 , n14375 , n14376 , n14377 , n14378 , n14379 , n14380 , n14381 , n14382 , n14383 , n14384 , n14385 , n14386 , n14387 , n14388 , n14389 , n14390 , n14391 , n14392 , n14393 , n14394 , n14395 , n14396 , n14397 , n14398 , n14399 , n14400 , n14401 , n14402 , n14403 , n14404 , n14405 , n14406 , n14407 , n14408 , n14409 , n14410 , n14411 , n14412 , n14413 , n14414 , n14415 , n14416 , n14417 , n14418 , n14419 , n14420 , n14421 , n14422 , n14423 , n14424 , n14425 , n14426 , n14427 , n14428 , n14429 , n14430 , n14431 , n14432 , n14433 , n14434 , n14435 , n14436 , n14437 , n14438 , n14439 , n14440 , n14441 , n14442 , n14443 , n14444 , n14445 , n14446 , n14447 , n14448 , n14449 , n14450 , n14451 , n14452 , n14453 , n14454 , n14455 , n14456 , n14457 , n14458 , n14459 , n14460 , n14461 , n14462 , n14463 , n14464 , n14465 , n14466 , n14467 , n14468 , n14469 , n14470 , n14471 , n14472 , n14473 , n14474 , n14475 , n14476 , n14477 , n14478 , n14479 , n14480 , n14481 , n14482 , n14483 , n14484 , n14485 , n14486 , n14487 , n14488 , n14489 , n14490 , n14491 , n14492 , n14493 , n14494 , n14495 , n14496 , n14497 , n14498 , n14499 , n14500 , n14501 , n14502 , n14503 , n14504 , n14505 , n14506 , n14507 , n14508 , n14509 , n14510 , n14511 , n14512 , n14513 , n14514 , n14515 , n14516 , n14517 , n14518 , n14519 , n14520 , n14521 , n14522 , n14523 , n14524 , n14525 , n14526 , n14527 , n14528 , n14529 , n14530 , n14531 , n14532 , n14533 , n14534 , n14535 , n14536 , n14537 , n14538 , n14539 , n14540 , n14541 , n14542 , n14543 , n14544 , n14545 , n14546 , n14547 , n14548 , n14549 , n14550 , n14551 , n14552 , n14553 , n14554 , n14555 , n14556 , n14557 , n14558 , n14559 , n14560 , n14561 , n14562 , n14563 , n14564 , n14565 , n14566 , n14567 , n14568 , n14569 , n14570 , n14571 , n14572 , n14573 , n14574 , n14575 , n14576 , n14577 , n14578 , n14579 , n14580 , n14581 , n14582 , n14583 , n14584 , n14585 , n14586 , n14587 , n14588 , n14589 , n14590 , n14591 , n14592 , n14593 , n14594 , n14595 , n14596 , n14597 , n14598 , n14599 , n14600 , n14601 , n14602 , n14603 , n14604 , n14605 , n14606 , n14607 , n14608 , n14609 , n14610 , n14611 , n14612 , n14613 , n14614 , n14615 , n14616 , n14617 , n14618 , n14619 , n14620 , n14621 , n14622 , n14623 , n14624 , n14625 , n14626 , n14627 , n14628 , n14629 , n14630 , n14631 , n14632 , n14633 , n14634 , n14635 , n14636 , n14637 , n14638 , n14639 , n14640 , n14641 , n14642 , n14643 , n14644 , n14645 , n14646 , n14647 , n14648 , n14649 , n14650 , n14651 , n14652 , n14653 , n14654 , n14655 , n14656 , n14657 , n14658 , n14659 , n14660 , n14661 , n14662 , n14663 , n14664 , n14665 , n14666 , n14667 , n14668 , n14669 , n14670 , n14671 , n14672 , n14673 , n14674 , n14675 , n14676 , n14677 , n14678 , n14679 , n14680 , n14681 , n14682 , n14683 , n14684 , n14685 , n14686 , n14687 , n14688 , n14689 , n14690 , n14691 , n14692 , n14693 , n14694 , n14695 , n14696 , n14697 , n14698 , n14699 , n14700 , n14701 , n14702 , n14703 , n14704 , n14705 , n14706 , n14707 , n14708 , n14709 , n14710 , n14711 , n14712 , n14713 , n14714 , n14715 , n14716 , n14717 , n14718 , n14719 , n14720 , n14721 , n14722 , n14723 , n14724 , n14725 , n14726 , n14727 , n14728 , n14729 , n14730 , n14731 , n14732 , n14733 , n14734 , n14735 , n14736 , n14737 , n14738 , n14739 , n14740 , n14741 , n14742 , n14743 , n14744 , n14745 , n14746 , n14747 , n14748 , n14749 , n14750 , n14751 , n14752 , n14753 , n14754 , n14755 , n14756 , n14757 , n14758 , n14759 , n14760 , n14761 , n14762 , n14763 , n14764 , n14765 , n14766 , n14767 , n14768 , n14769 , n14770 , n14771 , n14772 , n14773 , n14774 , n14775 , n14776 , n14777 , n14778 , n14779 , n14780 , n14781 , n14782 , n14783 , n14784 , n14785 , n14786 , n14787 , n14788 , n14789 , n14790 , n14791 , n14792 , n14793 , n14794 , n14795 , n14796 , n14797 , n14798 , n14799 , n14800 , n14801 , n14802 , n14803 , n14804 , n14805 , n14806 , n14807 , n14808 , n14809 , n14810 , n14811 , n14812 , n14813 , n14814 , n14815 , n14816 , n14817 , n14818 , n14819 , n14820 , n14821 , n14822 , n14823 , n14824 , n14825 , n14826 , n14827 , n14828 , n14829 , n14830 , n14831 , n14832 , n14833 , n14834 , n14835 , n14836 , n14837 , n14838 , n14839 , n14840 , n14841 , n14842 , n14843 , n14844 , n14845 , n14846 , n14847 , n14848 , n14849 , n14850 , n14851 , n14852 , n14853 , n14854 , n14855 , n14856 , n14857 , n14858 , n14859 , n14860 , n14861 , n14862 , n14863 , n14864 , n14865 , n14866 , n14867 , n14868 , n14869 , n14870 , n14871 , n14872 , n14873 , n14874 , n14875 , n14876 , n14877 , n14878 , n14879 , n14880 , n14881 , n14882 , n14883 , n14884 , n14885 , n14886 , n14887 , n14888 , n14889 , n14890 , n14891 , n14892 , n14893 , n14894 , n14895 , n14896 , n14897 , n14898 , n14899 , n14900 , n14901 , n14902 , n14903 , n14904 , n14905 , n14906 , n14907 , n14908 , n14909 , n14910 , n14911 , n14912 , n14913 , n14914 , n14915 , n14916 , n14917 , n14918 , n14919 , n14920 , n14921 , n14922 , n14923 , n14924 , n14925 , n14926 , n14927 , n14928 , n14929 , n14930 , n14931 , n14932 , n14933 , n14934 , n14935 , n14936 , n14937 , n14938 , n14939 , n14940 , n14941 , n14942 , n14943 , n14944 , n14945 , n14946 , n14947 , n14948 , n14949 , n14950 , n14951 , n14952 , n14953 , n14954 , n14955 , n14956 , n14957 , n14958 , n14959 , n14960 , n14961 , n14962 , n14963 , n14964 , n14965 , n14966 , n14967 , n14968 , n14969 , n14970 , n14971 , n14972 , n14973 , n14974 , n14975 , n14976 , n14977 , n14978 , n14979 , n14980 , n14981 , n14982 , n14983 , n14984 , n14985 , n14986 , n14987 , n14988 , n14989 , n14990 , n14991 , n14992 , n14993 , n14994 , n14995 , n14996 , n14997 , n14998 , n14999 , n15000 , n15001 , n15002 , n15003 , n15004 , n15005 , n15006 , n15007 , n15008 , n15009 , n15010 , n15011 , n15012 , n15013 , n15014 , n15015 , n15016 , n15017 , n15018 , n15019 , n15020 , n15021 , n15022 , n15023 , n15024 , n15025 , n15026 , n15027 , n15028 , n15029 , n15030 , n15031 , n15032 , n15033 , n15034 , n15035 , n15036 , n15037 , n15038 , n15039 , n15040 , n15041 , n15042 , n15043 , n15044 , n15045 , n15046 , n15047 , n15048 , n15049 , n15050 , n15051 , n15052 , n15053 , n15054 , n15055 , n15056 , n15057 , n15058 , n15059 , n15060 , n15061 , n15062 , n15063 , n15064 , n15065 , n15066 , n15067 , n15068 , n15069 , n15070 , n15071 , n15072 , n15073 , n15074 , n15075 , n15076 , n15077 , n15078 , n15079 , n15080 , n15081 , n15082 , n15083 , n15084 , n15085 , n15086 , n15087 , n15088 , n15089 , n15090 , n15091 , n15092 , n15093 , n15094 , n15095 , n15096 , n15097 , n15098 , n15099 , n15100 , n15101 , n15102 , n15103 , n15104 , n15105 , n15106 , n15107 , n15108 , n15109 , n15110 , n15111 , n15112 , n15113 , n15114 , n15115 , n15116 , n15117 , n15118 , n15119 , n15120 , n15121 , n15122 , n15123 , n15124 , n15125 , n15126 , n15127 , n15128 , n15129 , n15130 , n15131 , n15132 , n15133 , n15134 , n15135 , n15136 , n15137 , n15138 , n15139 , n15140 , n15141 , n15142 , n15143 , n15144 , n15145 , n15146 , n15147 , n15148 , n15149 , n15150 , n15151 , n15152 , n15153 , n15154 , n15155 , n15156 , n15157 , n15158 , n15159 , n15160 , n15161 , n15162 , n15163 , n15164 , n15165 , n15166 , n15167 , n15168 , n15169 , n15170 , n15171 , n15172 , n15173 , n15174 , n15175 , n15176 , n15177 , n15178 , n15179 , n15180 , n15181 , n15182 , n15183 , n15184 , n15185 , n15186 , n15187 , n15188 , n15189 , n15190 , n15191 , n15192 , n15193 , n15194 , n15195 , n15196 , n15197 , n15198 , n15199 , n15200 , n15201 , n15202 , n15203 , n15204 , n15205 , n15206 , n15207 , n15208 , n15209 , n15210 , n15211 , n15212 , n15213 , n15214 , n15215 , n15216 , n15217 , n15218 , n15219 , n15220 , n15221 , n15222 , n15223 , n15224 , n15225 , n15226 , n15227 , n15228 , n15229 , n15230 , n15231 , n15232 , n15233 , n15234 , n15235 , n15236 , n15237 , n15238 , n15239 , n15240 , n15241 , n15242 , n15243 , n15244 , n15245 , n15246 , n15247 , n15248 , n15249 , n15250 , n15251 , n15252 , n15253 , n15254 , n15255 , n15256 , n15257 , n15258 , n15259 , n15260 , n15261 , n15262 , n15263 , n15264 , n15265 , n15266 , n15267 , n15268 , n15269 , n15270 , n15271 , n15272 , n15273 , n15274 , n15275 , n15276 , n15277 , n15278 , n15279 , n15280 , n15281 , n15282 , n15283 , n15284 , n15285 , n15286 , n15287 , n15288 , n15289 , n15290 , n15291 , n15292 , n15293 , n15294 , n15295 , n15296 , n15297 , n15298 , n15299 , n15300 , n15301 , n15302 , n15303 , n15304 , n15305 , n15306 , n15307 , n15308 , n15309 , n15310 , n15311 , n15312 , n15313 , n15314 , n15315 , n15316 , n15317 , n15318 , n15319 , n15320 , n15321 , n15322 , n15323 , n15324 , n15325 , n15326 , n15327 , n15328 , n15329 , n15330 , n15331 , n15332 , n15333 , n15334 , n15335 , n15336 , n15337 , n15338 , n15339 , n15340 , n15341 , n15342 , n15343 , n15344 , n15345 , n15346 , n15347 , n15348 , n15349 , n15350 , n15351 , n15352 , n15353 , n15354 , n15355 , n15356 , n15357 , n15358 , n15359 , n15360 , n15361 , n15362 , n15363 , n15364 , n15365 , n15366 , n15367 , n15368 , n15369 , n15370 , n15371 , n15372 , n15373 , n15374 , n15375 , n15376 , n15377 , n15378 , n15379 , n15380 , n15381 , n15382 , n15383 , n15384 , n15385 , n15386 , n15387 , n15388 , n15389 , n15390 , n15391 , n15392 , n15393 , n15394 , n15395 , n15396 , n15397 , n15398 , n15399 , n15400 , n15401 , n15402 , n15403 , n15404 , n15405 , n15406 , n15407 , n15408 , n15409 , n15410 , n15411 , n15412 , n15413 , n15414 , n15415 , n15416 , n15417 , n15418 , n15419 , n15420 , n15421 , n15422 , n15423 , n15424 , n15425 , n15426 , n15427 , n15428 , n15429 , n15430 , n15431 , n15432 , n15433 , n15434 , n15435 , n15436 , n15437 , n15438 , n15439 , n15440 , n15441 , n15442 , n15443 , n15444 , n15445 , n15446 , n15447 , n15448 , n15449 , n15450 , n15451 , n15452 , n15453 , n15454 , n15455 , n15456 , n15457 , n15458 , n15459 , n15460 , n15461 , n15462 , n15463 , n15464 , n15465 , n15466 , n15467 , n15468 , n15469 , n15470 , n15471 , n15472 , n15473 , n15474 , n15475 , n15476 , n15477 , n15478 , n15479 , n15480 , n15481 , n15482 , n15483 , n15484 , n15485 , n15486 , n15487 , n15488 , n15489 , n15490 , n15491 , n15492 , n15493 , n15494 , n15495 , n15496 , n15497 , n15498 , n15499 , n15500 , n15501 , n15502 , n15503 , n15504 , n15505 , n15506 , n15507 , n15508 , n15509 , n15510 , n15511 , n15512 , n15513 , n15514 , n15515 , n15516 , n15517 , n15518 , n15519 , n15520 , n15521 , n15522 , n15523 , n15524 , n15525 , n15526 , n15527 , n15528 , n15529 , n15530 , n15531 , n15532 , n15533 , n15534 , n15535 , n15536 , n15537 , n15538 , n15539 , n15540 , n15541 , n15542 , n15543 , n15544 , n15545 , n15546 , n15547 , n15548 , n15549 , n15550 , n15551 , n15552 , n15553 , n15554 , n15555 , n15556 , n15557 , n15558 , n15559 , n15560 , n15561 , n15562 , n15563 , n15564 , n15565 , n15566 , n15567 , n15568 , n15569 , n15570 , n15571 , n15572 , n15573 , n15574 , n15575 , n15576 , n15577 , n15578 , n15579 , n15580 , n15581 , n15582 , n15583 , n15584 , n15585 , n15586 , n15587 , n15588 , n15589 , n15590 , n15591 , n15592 , n15593 , n15594 , n15595 , n15596 , n15597 , n15598 , n15599 , n15600 , n15601 , n15602 , n15603 , n15604 , n15605 , n15606 , n15607 , n15608 , n15609 , n15610 , n15611 , n15612 , n15613 , n15614 , n15615 , n15616 , n15617 , n15618 , n15619 , n15620 , n15621 , n15622 , n15623 , n15624 , n15625 , n15626 , n15627 , n15628 , n15629 , n15630 , n15631 , n15632 , n15633 , n15634 , n15635 , n15636 , n15637 , n15638 , n15639 , n15640 , n15641 , n15642 , n15643 , n15644 , n15645 , n15646 , n15647 , n15648 , n15649 , n15650 , n15651 , n15652 , n15653 , n15654 , n15655 , n15656 , n15657 , n15658 , n15659 , n15660 , n15661 , n15662 , n15663 , n15664 , n15665 , n15666 , n15667 , n15668 , n15669 , n15670 , n15671 , n15672 , n15673 , n15674 , n15675 , n15676 , n15677 , n15678 , n15679 , n15680 , n15681 , n15682 , n15683 , n15684 , n15685 , n15686 , n15687 , n15688 , n15689 , n15690 , n15691 , n15692 , n15693 , n15694 , n15695 , n15696 , n15697 , n15698 , n15699 , n15700 , n15701 , n15702 , n15703 , n15704 , n15705 , n15706 , n15707 , n15708 , n15709 , n15710 , n15711 , n15712 , n15713 , n15714 , n15715 , n15716 , n15717 , n15718 , n15719 , n15720 , n15721 , n15722 , n15723 , n15724 , n15725 , n15726 , n15727 , n15728 , n15729 , n15730 , n15731 , n15732 , n15733 , n15734 , n15735 , n15736 , n15737 , n15738 , n15739 , n15740 , n15741 , n15742 , n15743 , n15744 , n15745 , n15746 , n15747 , n15748 , n15749 , n15750 , n15751 , n15752 , n15753 , n15754 , n15755 , n15756 , n15757 , n15758 , n15759 , n15760 , n15761 , n15762 , n15763 , n15764 , n15765 , n15766 , n15767 , n15768 , n15769 , n15770 , n15771 , n15772 , n15773 , n15774 , n15775 , n15776 , n15777 , n15778 , n15779 , n15780 , n15781 , n15782 , n15783 , n15784 , n15785 , n15786 , n15787 , n15788 , n15789 , n15790 , n15791 , n15792 , n15793 , n15794 , n15795 , n15796 , n15797 , n15798 , n15799 , n15800 , n15801 , n15802 , n15803 , n15804 , n15805 , n15806 , n15807 , n15808 , n15809 , n15810 , n15811 , n15812 , n15813 , n15814 , n15815 , n15816 , n15817 , n15818 , n15819 , n15820 , n15821 , n15822 , n15823 , n15824 , n15825 , n15826 , n15827 , n15828 , n15829 , n15830 , n15831 , n15832 , n15833 , n15834 , n15835 , n15836 , n15837 , n15838 , n15839 , n15840 , n15841 , n15842 , n15843 , n15844 , n15845 , n15846 , n15847 , n15848 , n15849 , n15850 , n15851 , n15852 , n15853 , n15854 , n15855 , n15856 , n15857 , n15858 , n15859 , n15860 , n15861 , n15862 , n15863 , n15864 , n15865 , n15866 , n15867 , n15868 , n15869 , n15870 , n15871 , n15872 , n15873 , n15874 , n15875 , n15876 , n15877 , n15878 , n15879 , n15880 , n15881 , n15882 , n15883 , n15884 , n15885 , n15886 , n15887 , n15888 , n15889 , n15890 , n15891 , n15892 , n15893 , n15894 , n15895 , n15896 , n15897 , n15898 , n15899 , n15900 , n15901 , n15902 , n15903 , n15904 , n15905 , n15906 , n15907 , n15908 , n15909 , n15910 , n15911 , n15912 , n15913 , n15914 , n15915 , n15916 , n15917 , n15918 , n15919 , n15920 , n15921 , n15922 , n15923 , n15924 , n15925 , n15926 , n15927 , n15928 , n15929 , n15930 , n15931 , n15932 , n15933 , n15934 , n15935 , n15936 , n15937 , n15938 , n15939 , n15940 , n15941 , n15942 , n15943 , n15944 , n15945 , n15946 , n15947 , n15948 , n15949 , n15950 , n15951 , n15952 , n15953 , n15954 , n15955 , n15956 , n15957 , n15958 , n15959 , n15960 , n15961 , n15962 , n15963 , n15964 , n15965 , n15966 , n15967 , n15968 , n15969 , n15970 , n15971 , n15972 , n15973 , n15974 , n15975 , n15976 , n15977 , n15978 , n15979 , n15980 , n15981 , n15982 , n15983 , n15984 , n15985 , n15986 , n15987 , n15988 , n15989 , n15990 , n15991 , n15992 , n15993 , n15994 , n15995 , n15996 , n15997 , n15998 , n15999 , n16000 , n16001 , n16002 , n16003 , n16004 , n16005 , n16006 , n16007 , n16008 , n16009 , n16010 , n16011 , n16012 , n16013 , n16014 , n16015 , n16016 , n16017 , n16018 , n16019 , n16020 , n16021 , n16022 , n16023 , n16024 , n16025 , n16026 , n16027 , n16028 , n16029 , n16030 , n16031 , n16032 , n16033 , n16034 , n16035 , n16036 , n16037 , n16038 , n16039 , n16040 , n16041 , n16042 , n16043 , n16044 , n16045 , n16046 , n16047 , n16048 , n16049 , n16050 , n16051 , n16052 , n16053 , n16054 , n16055 , n16056 , n16057 , n16058 , n16059 , n16060 , n16061 , n16062 , n16063 , n16064 , n16065 , n16066 , n16067 , n16068 , n16069 , n16070 , n16071 , n16072 , n16073 , n16074 , n16075 , n16076 , n16077 , n16078 , n16079 , n16080 , n16081 , n16082 , n16083 , n16084 , n16085 , n16086 , n16087 , n16088 , n16089 , n16090 , n16091 , n16092 , n16093 , n16094 , n16095 , n16096 , n16097 , n16098 , n16099 , n16100 , n16101 , n16102 , n16103 , n16104 , n16105 , n16106 , n16107 , n16108 , n16109 , n16110 , n16111 , n16112 , n16113 , n16114 , n16115 , n16116 , n16117 , n16118 , n16119 , n16120 , n16121 , n16122 , n16123 , n16124 , n16125 , n16126 , n16127 , n16128 , n16129 , n16130 , n16131 , n16132 , n16133 , n16134 , n16135 , n16136 , n16137 , n16138 , n16139 , n16140 , n16141 , n16142 , n16143 , n16144 , n16145 , n16146 , n16147 , n16148 , n16149 , n16150 , n16151 , n16152 , n16153 , n16154 , n16155 , n16156 , n16157 , n16158 , n16159 , n16160 , n16161 , n16162 , n16163 , n16164 , n16165 , n16166 , n16167 , n16168 , n16169 , n16170 , n16171 , n16172 , n16173 , n16174 , n16175 , n16176 , n16177 , n16178 , n16179 , n16180 , n16181 , n16182 , n16183 , n16184 , n16185 , n16186 , n16187 , n16188 , n16189 , n16190 , n16191 , n16192 , n16193 , n16194 , n16195 , n16196 , n16197 , n16198 , n16199 , n16200 , n16201 , n16202 , n16203 , n16204 , n16205 , n16206 , n16207 , n16208 , n16209 , n16210 , n16211 , n16212 , n16213 , n16214 , n16215 , n16216 , n16217 , n16218 , n16219 , n16220 , n16221 , n16222 , n16223 , n16224 , n16225 , n16226 , n16227 , n16228 , n16229 , n16230 , n16231 , n16232 , n16233 , n16234 , n16235 , n16236 , n16237 , n16238 , n16239 , n16240 , n16241 , n16242 , n16243 , n16244 , n16245 , n16246 , n16247 , n16248 , n16249 , n16250 , n16251 , n16252 , n16253 , n16254 , n16255 , n16256 , n16257 , n16258 , n16259 , n16260 , n16261 , n16262 , n16263 , n16264 , n16265 , n16266 , n16267 , n16268 , n16269 , n16270 , n16271 , n16272 , n16273 , n16274 , n16275 , n16276 , n16277 , n16278 , n16279 , n16280 , n16281 , n16282 , n16283 , n16284 , n16285 , n16286 , n16287 , n16288 , n16289 , n16290 , n16291 , n16292 , n16293 , n16294 , n16295 , n16296 , n16297 , n16298 , n16299 , n16300 , n16301 , n16302 , n16303 , n16304 , n16305 , n16306 , n16307 , n16308 , n16309 , n16310 , n16311 , n16312 , n16313 , n16314 , n16315 , n16316 , n16317 , n16318 , n16319 , n16320 , n16321 , n16322 , n16323 , n16324 , n16325 , n16326 , n16327 , n16328 , n16329 , n16330 , n16331 , n16332 , n16333 , n16334 , n16335 , n16336 , n16337 , n16338 , n16339 , n16340 , n16341 , n16342 , n16343 , n16344 , n16345 , n16346 , n16347 , n16348 , n16349 , n16350 , n16351 , n16352 , n16353 , n16354 , n16355 , n16356 , n16357 , n16358 , n16359 , n16360 , n16361 , n16362 , n16363 , n16364 , n16365 , n16366 , n16367 , n16368 , n16369 , n16370 , n16371 , n16372 , n16373 , n16374 , n16375 , n16376 , n16377 , n16378 , n16379 , n16380 , n16381 , n16382 , n16383 , n16384 , n16385 , n16386 , n16387 , n16388 , n16389 , n16390 , n16391 , n16392 , n16393 , n16394 , n16395 , n16396 , n16397 , n16398 , n16399 , n16400 , n16401 , n16402 , n16403 , n16404 , n16405 , n16406 , n16407 , n16408 , n16409 , n16410 , n16411 , n16412 , n16413 , n16414 , n16415 , n16416 , n16417 , n16418 , n16419 , n16420 , n16421 , n16422 , n16423 , n16424 , n16425 , n16426 , n16427 , n16428 , n16429 , n16430 , n16431 , n16432 , n16433 , n16434 , n16435 , n16436 , n16437 , n16438 , n16439 , n16440 , n16441 , n16442 , n16443 , n16444 , n16445 , n16446 , n16447 , n16448 , n16449 , n16450 , n16451 , n16452 , n16453 , n16454 , n16455 , n16456 , n16457 , n16458 , n16459 , n16460 , n16461 , n16462 , n16463 , n16464 , n16465 , n16466 , n16467 , n16468 , n16469 , n16470 , n16471 , n16472 , n16473 , n16474 , n16475 , n16476 , n16477 , n16478 , n16479 , n16480 , n16481 , n16482 , n16483 , n16484 , n16485 , n16486 , n16487 , n16488 , n16489 , n16490 , n16491 , n16492 , n16493 , n16494 , n16495 , n16496 , n16497 , n16498 , n16499 , n16500 , n16501 , n16502 , n16503 , n16504 , n16505 , n16506 , n16507 , n16508 , n16509 , n16510 , n16511 , n16512 , n16513 , n16514 , n16515 , n16516 , n16517 , n16518 , n16519 , n16520 , n16521 , n16522 , n16523 , n16524 , n16525 , n16526 , n16527 , n16528 , n16529 , n16530 , n16531 , n16532 , n16533 , n16534 , n16535 , n16536 , n16537 , n16538 , n16539 , n16540 , n16541 , n16542 , n16543 , n16544 , n16545 , n16546 , n16547 , n16548 , n16549 , n16550 , n16551 , n16552 , n16553 , n16554 , n16555 , n16556 , n16557 , n16558 , n16559 , n16560 , n16561 , n16562 , n16563 , n16564 , n16565 , n16566 , n16567 , n16568 , n16569 , n16570 , n16571 , n16572 , n16573 , n16574 , n16575 , n16576 , n16577 , n16578 , n16579 , n16580 , n16581 , n16582 , n16583 , n16584 , n16585 , n16586 , n16587 , n16588 , n16589 , n16590 , n16591 , n16592 , n16593 , n16594 , n16595 , n16596 , n16597 , n16598 , n16599 , n16600 , n16601 , n16602 , n16603 , n16604 , n16605 , n16606 , n16607 , n16608 , n16609 , n16610 , n16611 , n16612 , n16613 , n16614 , n16615 , n16616 , n16617 , n16618 , n16619 , n16620 , n16621 , n16622 , n16623 , n16624 , n16625 , n16626 , n16627 , n16628 , n16629 , n16630 , n16631 , n16632 , n16633 , n16634 , n16635 , n16636 , n16637 , n16638 , n16639 , n16640 , n16641 , n16642 , n16643 , n16644 , n16645 , n16646 , n16647 , n16648 , n16649 , n16650 , n16651 , n16652 , n16653 , n16654 , n16655 , n16656 , n16657 , n16658 , n16659 , n16660 , n16661 , n16662 , n16663 , n16664 , n16665 , n16666 , n16667 , n16668 , n16669 , n16670 , n16671 , n16672 , n16673 , n16674 , n16675 , n16676 , n16677 , n16678 , n16679 , n16680 , n16681 , n16682 , n16683 , n16684 , n16685 , n16686 , n16687 , n16688 , n16689 , n16690 , n16691 , n16692 , n16693 , n16694 , n16695 , n16696 , n16697 , n16698 , n16699 , n16700 , n16701 , n16702 , n16703 , n16704 , n16705 , n16706 , n16707 , n16708 , n16709 , n16710 , n16711 , n16712 , n16713 , n16714 , n16715 , n16716 , n16717 , n16718 , n16719 , n16720 , n16721 , n16722 , n16723 , n16724 , n16725 , n16726 , n16727 , n16728 , n16729 , n16730 , n16731 , n16732 , n16733 , n16734 , n16735 , n16736 , n16737 , n16738 , n16739 , n16740 , n16741 , n16742 , n16743 , n16744 , n16745 , n16746 , n16747 , n16748 , n16749 , n16750 , n16751 , n16752 , n16753 , n16754 , n16755 , n16756 , n16757 , n16758 , n16759 , n16760 , n16761 , n16762 , n16763 , n16764 , n16765 , n16766 , n16767 , n16768 , n16769 , n16770 , n16771 , n16772 , n16773 , n16774 , n16775 , n16776 , n16777 , n16778 , n16779 , n16780 , n16781 , n16782 , n16783 , n16784 , n16785 , n16786 , n16787 , n16788 , n16789 , n16790 , n16791 , n16792 , n16793 , n16794 , n16795 , n16796 , n16797 , n16798 , n16799 , n16800 , n16801 , n16802 , n16803 , n16804 , n16805 , n16806 , n16807 , n16808 , n16809 , n16810 , n16811 , n16812 , n16813 , n16814 , n16815 , n16816 , n16817 , n16818 , n16819 , n16820 , n16821 , n16822 , n16823 , n16824 , n16825 , n16826 , n16827 , n16828 , n16829 , n16830 , n16831 , n16832 , n16833 , n16834 , n16835 , n16836 , n16837 , n16838 , n16839 , n16840 , n16841 , n16842 , n16843 , n16844 , n16845 , n16846 , n16847 , n16848 , n16849 , n16850 , n16851 , n16852 , n16853 , n16854 , n16855 , n16856 , n16857 , n16858 , n16859 , n16860 , n16861 , n16862 , n16863 , n16864 , n16865 , n16866 , n16867 , n16868 , n16869 , n16870 , n16871 , n16872 , n16873 , n16874 , n16875 , n16876 , n16877 , n16878 , n16879 , n16880 , n16881 , n16882 , n16883 , n16884 , n16885 , n16886 , n16887 , n16888 , n16889 , n16890 , n16891 , n16892 , n16893 , n16894 , n16895 , n16896 , n16897 , n16898 , n16899 , n16900 , n16901 , n16902 , n16903 , n16904 , n16905 , n16906 , n16907 , n16908 , n16909 , n16910 , n16911 , n16912 , n16913 , n16914 , n16915 , n16916 , n16917 , n16918 , n16919 , n16920 , n16921 , n16922 , n16923 , n16924 , n16925 , n16926 , n16927 , n16928 , n16929 , n16930 , n16931 , n16932 , n16933 , n16934 , n16935 , n16936 , n16937 , n16938 , n16939 , n16940 , n16941 , n16942 , n16943 , n16944 , n16945 , n16946 , n16947 , n16948 , n16949 , n16950 , n16951 , n16952 , n16953 , n16954 , n16955 , n16956 , n16957 , n16958 , n16959 , n16960 , n16961 , n16962 , n16963 , n16964 , n16965 , n16966 , n16967 , n16968 , n16969 , n16970 , n16971 , n16972 , n16973 , n16974 , n16975 , n16976 , n16977 , n16978 , n16979 , n16980 , n16981 , n16982 , n16983 , n16984 , n16985 , n16986 , n16987 , n16988 , n16989 , n16990 , n16991 , n16992 , n16993 , n16994 , n16995 , n16996 , n16997 , n16998 , n16999 , n17000 , n17001 , n17002 , n17003 , n17004 , n17005 , n17006 , n17007 , n17008 , n17009 , n17010 , n17011 , n17012 , n17013 , n17014 , n17015 , n17016 , n17017 , n17018 , n17019 , n17020 , n17021 , n17022 , n17023 , n17024 , n17025 , n17026 , n17027 , n17028 , n17029 , n17030 , n17031 , n17032 , n17033 , n17034 , n17035 , n17036 , n17037 , n17038 , n17039 , n17040 , n17041 , n17042 , n17043 , n17044 , n17045 , n17046 , n17047 , n17048 , n17049 , n17050 , n17051 , n17052 , n17053 , n17054 , n17055 , n17056 , n17057 , n17058 , n17059 , n17060 , n17061 , n17062 , n17063 , n17064 , n17065 , n17066 , n17067 , n17068 , n17069 , n17070 , n17071 , n17072 , n17073 , n17074 , n17075 , n17076 , n17077 , n17078 , n17079 , n17080 , n17081 , n17082 , n17083 , n17084 , n17085 , n17086 , n17087 , n17088 , n17089 , n17090 , n17091 , n17092 , n17093 , n17094 , n17095 , n17096 , n17097 , n17098 , n17099 , n17100 , n17101 , n17102 , n17103 , n17104 , n17105 , n17106 , n17107 , n17108 , n17109 , n17110 , n17111 , n17112 , n17113 , n17114 , n17115 , n17116 , n17117 , n17118 , n17119 , n17120 , n17121 , n17122 , n17123 , n17124 , n17125 , n17126 , n17127 , n17128 , n17129 , n17130 , n17131 , n17132 , n17133 , n17134 , n17135 , n17136 , n17137 , n17138 , n17139 , n17140 , n17141 , n17142 , n17143 , n17144 , n17145 , n17146 , n17147 , n17148 , n17149 , n17150 , n17151 , n17152 , n17153 , n17154 , n17155 , n17156 , n17157 , n17158 , n17159 , n17160 , n17161 , n17162 , n17163 , n17164 , n17165 , n17166 , n17167 , n17168 , n17169 , n17170 , n17171 , n17172 , n17173 , n17174 , n17175 , n17176 , n17177 , n17178 , n17179 , n17180 , n17181 , n17182 , n17183 , n17184 , n17185 , n17186 , n17187 , n17188 , n17189 , n17190 , n17191 , n17192 , n17193 , n17194 , n17195 , n17196 , n17197 , n17198 , n17199 , n17200 , n17201 , n17202 , n17203 , n17204 , n17205 , n17206 , n17207 , n17208 , n17209 , n17210 , n17211 , n17212 , n17213 , n17214 , n17215 , n17216 , n17217 , n17218 , n17219 , n17220 , n17221 , n17222 , n17223 , n17224 , n17225 , n17226 , n17227 , n17228 , n17229 , n17230 , n17231 , n17232 , n17233 , n17234 , n17235 , n17236 , n17237 , n17238 , n17239 , n17240 , n17241 , n17242 , n17243 , n17244 , n17245 , n17246 , n17247 , n17248 , n17249 , n17250 , n17251 , n17252 , n17253 , n17254 , n17255 , n17256 , n17257 , n17258 , n17259 , n17260 , n17261 , n17262 , n17263 , n17264 , n17265 , n17266 , n17267 , n17268 , n17269 , n17270 , n17271 , n17272 , n17273 , n17274 , n17275 , n17276 , n17277 , n17278 , n17279 , n17280 , n17281 , n17282 , n17283 , n17284 , n17285 , n17286 , n17287 , n17288 , n17289 , n17290 , n17291 , n17292 , n17293 , n17294 , n17295 , n17296 , n17297 , n17298 , n17299 , n17300 , n17301 , n17302 , n17303 , n17304 , n17305 , n17306 , n17307 , n17308 , n17309 , n17310 , n17311 , n17312 , n17313 , n17314 , n17315 , n17316 , n17317 , n17318 , n17319 , n17320 , n17321 , n17322 , n17323 , n17324 , n17325 , n17326 , n17327 , n17328 , n17329 , n17330 , n17331 , n17332 , n17333 , n17334 , n17335 , n17336 , n17337 , n17338 , n17339 , n17340 , n17341 , n17342 , n17343 , n17344 , n17345 , n17346 , n17347 , n17348 , n17349 , n17350 , n17351 , n17352 , n17353 , n17354 , n17355 , n17356 , n17357 , n17358 , n17359 , n17360 , n17361 , n17362 , n17363 , n17364 , n17365 , n17366 , n17367 , n17368 , n17369 , n17370 , n17371 , n17372 , n17373 , n17374 , n17375 , n17376 , n17377 , n17378 , n17379 , n17380 , n17381 , n17382 , n17383 , n17384 , n17385 , n17386 , n17387 , n17388 , n17389 , n17390 , n17391 , n17392 , n17393 , n17394 , n17395 , n17396 , n17397 , n17398 , n17399 , n17400 , n17401 , n17402 , n17403 , n17404 , n17405 , n17406 , n17407 , n17408 , n17409 , n17410 , n17411 , n17412 , n17413 , n17414 , n17415 , n17416 , n17417 , n17418 , n17419 , n17420 , n17421 , n17422 , n17423 , n17424 , n17425 , n17426 , n17427 , n17428 , n17429 , n17430 , n17431 , n17432 , n17433 , n17434 , n17435 , n17436 , n17437 , n17438 , n17439 , n17440 , n17441 , n17442 , n17443 , n17444 , n17445 , n17446 , n17447 , n17448 , n17449 , n17450 , n17451 , n17452 , n17453 , n17454 , n17455 , n17456 , n17457 , n17458 , n17459 , n17460 , n17461 , n17462 , n17463 , n17464 , n17465 , n17466 , n17467 , n17468 , n17469 , n17470 , n17471 , n17472 , n17473 , n17474 , n17475 , n17476 , n17477 , n17478 , n17479 , n17480 , n17481 , n17482 , n17483 , n17484 , n17485 , n17486 , n17487 , n17488 , n17489 , n17490 , n17491 , n17492 , n17493 , n17494 , n17495 , n17496 , n17497 , n17498 , n17499 , n17500 , n17501 , n17502 , n17503 , n17504 , n17505 , n17506 , n17507 , n17508 , n17509 , n17510 , n17511 , n17512 , n17513 , n17514 , n17515 , n17516 , n17517 , n17518 , n17519 , n17520 , n17521 , n17522 , n17523 , n17524 , n17525 , n17526 , n17527 , n17528 , n17529 , n17530 , n17531 , n17532 , n17533 , n17534 , n17535 , n17536 , n17537 , n17538 , n17539 , n17540 , n17541 , n17542 , n17543 , n17544 , n17545 , n17546 , n17547 , n17548 , n17549 , n17550 , n17551 , n17552 , n17553 , n17554 , n17555 , n17556 , n17557 , n17558 , n17559 , n17560 , n17561 , n17562 , n17563 , n17564 , n17565 , n17566 , n17567 , n17568 , n17569 , n17570 , n17571 , n17572 , n17573 , n17574 , n17575 , n17576 , n17577 , n17578 , n17579 , n17580 , n17581 , n17582 , n17583 , n17584 , n17585 , n17586 , n17587 , n17588 , n17589 , n17590 , n17591 , n17592 , n17593 , n17594 , n17595 , n17596 , n17597 , n17598 , n17599 , n17600 , n17601 , n17602 , n17603 , n17604 , n17605 , n17606 , n17607 , n17608 , n17609 , n17610 , n17611 , n17612 , n17613 , n17614 , n17615 , n17616 , n17617 , n17618 , n17619 , n17620 , n17621 , n17622 , n17623 , n17624 , n17625 , n17626 , n17627 , n17628 , n17629 , n17630 , n17631 , n17632 , n17633 , n17634 , n17635 , n17636 , n17637 , n17638 , n17639 , n17640 , n17641 , n17642 , n17643 , n17644 , n17645 , n17646 , n17647 , n17648 , n17649 , n17650 , n17651 , n17652 , n17653 , n17654 , n17655 , n17656 , n17657 , n17658 , n17659 , n17660 , n17661 , n17662 , n17663 , n17664 , n17665 , n17666 , n17667 , n17668 , n17669 , n17670 , n17671 , n17672 , n17673 , n17674 , n17675 , n17676 , n17677 , n17678 , n17679 , n17680 , n17681 , n17682 , n17683 , n17684 , n17685 , n17686 , n17687 , n17688 , n17689 , n17690 , n17691 , n17692 , n17693 , n17694 , n17695 , n17696 , n17697 , n17698 , n17699 , n17700 , n17701 , n17702 , n17703 , n17704 , n17705 , n17706 , n17707 , n17708 , n17709 , n17710 , n17711 , n17712 , n17713 , n17714 , n17715 , n17716 , n17717 , n17718 , n17719 , n17720 , n17721 , n17722 , n17723 , n17724 , n17725 , n17726 , n17727 , n17728 , n17729 , n17730 , n17731 , n17732 , n17733 , n17734 , n17735 , n17736 , n17737 , n17738 , n17739 , n17740 , n17741 , n17742 , n17743 , n17744 , n17745 , n17746 , n17747 , n17748 , n17749 , n17750 , n17751 , n17752 , n17753 , n17754 , n17755 , n17756 , n17757 , n17758 , n17759 , n17760 , n17761 , n17762 , n17763 , n17764 , n17765 , n17766 , n17767 , n17768 , n17769 , n17770 , n17771 , n17772 , n17773 , n17774 , n17775 , n17776 , n17777 , n17778 , n17779 , n17780 , n17781 , n17782 , n17783 , n17784 , n17785 , n17786 , n17787 , n17788 , n17789 , n17790 , n17791 , n17792 , n17793 , n17794 , n17795 , n17796 , n17797 , n17798 , n17799 , n17800 , n17801 , n17802 , n17803 , n17804 , n17805 , n17806 , n17807 , n17808 , n17809 , n17810 , n17811 , n17812 , n17813 , n17814 , n17815 , n17816 , n17817 , n17818 , n17819 , n17820 , n17821 , n17822 , n17823 , n17824 , n17825 , n17826 , n17827 , n17828 , n17829 , n17830 , n17831 , n17832 , n17833 , n17834 , n17835 , n17836 , n17837 , n17838 , n17839 , n17840 , n17841 , n17842 , n17843 , n17844 , n17845 , n17846 , n17847 , n17848 , n17849 , n17850 , n17851 , n17852 , n17853 , n17854 , n17855 , n17856 , n17857 , n17858 , n17859 , n17860 , n17861 , n17862 , n17863 , n17864 , n17865 , n17866 , n17867 , n17868 , n17869 , n17870 , n17871 , n17872 , n17873 , n17874 , n17875 , n17876 , n17877 , n17878 , n17879 , n17880 , n17881 , n17882 , n17883 , n17884 , n17885 , n17886 , n17887 , n17888 , n17889 , n17890 , n17891 , n17892 , n17893 , n17894 , n17895 , n17896 , n17897 , n17898 , n17899 , n17900 , n17901 , n17902 , n17903 , n17904 , n17905 , n17906 , n17907 , n17908 , n17909 , n17910 , n17911 , n17912 , n17913 , n17914 , n17915 , n17916 , n17917 , n17918 , n17919 , n17920 , n17921 , n17922 , n17923 , n17924 , n17925 , n17926 , n17927 , n17928 , n17929 , n17930 , n17931 , n17932 , n17933 , n17934 , n17935 , n17936 , n17937 , n17938 , n17939 , n17940 , n17941 , n17942 , n17943 , n17944 , n17945 , n17946 , n17947 , n17948 , n17949 , n17950 , n17951 , n17952 , n17953 , n17954 , n17955 , n17956 , n17957 , n17958 , n17959 , n17960 , n17961 , n17962 , n17963 , n17964 , n17965 , n17966 , n17967 , n17968 , n17969 , n17970 , n17971 , n17972 , n17973 , n17974 , n17975 , n17976 , n17977 , n17978 , n17979 , n17980 , n17981 , n17982 , n17983 , n17984 , n17985 , n17986 , n17987 , n17988 , n17989 , n17990 , n17991 , n17992 , n17993 , n17994 , n17995 , n17996 , n17997 , n17998 , n17999 , n18000 , n18001 , n18002 , n18003 , n18004 , n18005 , n18006 , n18007 , n18008 , n18009 , n18010 , n18011 , n18012 , n18013 , n18014 , n18015 , n18016 , n18017 , n18018 , n18019 , n18020 , n18021 , n18022 , n18023 , n18024 , n18025 , n18026 , n18027 , n18028 , n18029 , n18030 , n18031 , n18032 , n18033 , n18034 , n18035 , n18036 , n18037 , n18038 , n18039 , n18040 , n18041 , n18042 , n18043 , n18044 , n18045 , n18046 , n18047 , n18048 , n18049 , n18050 , n18051 , n18052 , n18053 , n18054 , n18055 , n18056 , n18057 , n18058 , n18059 , n18060 , n18061 , n18062 , n18063 , n18064 , n18065 , n18066 , n18067 , n18068 , n18069 , n18070 , n18071 , n18072 , n18073 , n18074 , n18075 , n18076 , n18077 , n18078 , n18079 , n18080 , n18081 , n18082 , n18083 , n18084 , n18085 , n18086 , n18087 , n18088 , n18089 , n18090 , n18091 , n18092 , n18093 , n18094 , n18095 , n18096 , n18097 , n18098 , n18099 , n18100 , n18101 , n18102 , n18103 , n18104 , n18105 , n18106 , n18107 , n18108 , n18109 , n18110 , n18111 , n18112 , n18113 , n18114 , n18115 , n18116 , n18117 , n18118 , n18119 , n18120 , n18121 , n18122 , n18123 , n18124 , n18125 , n18126 , n18127 , n18128 , n18129 , n18130 , n18131 , n18132 , n18133 , n18134 , n18135 , n18136 , n18137 , n18138 , n18139 , n18140 , n18141 , n18142 , n18143 , n18144 , n18145 , n18146 , n18147 , n18148 , n18149 , n18150 , n18151 , n18152 , n18153 , n18154 , n18155 , n18156 , n18157 , n18158 , n18159 , n18160 , n18161 , n18162 , n18163 , n18164 , n18165 , n18166 , n18167 , n18168 , n18169 , n18170 , n18171 , n18172 , n18173 , n18174 , n18175 , n18176 , n18177 , n18178 , n18179 , n18180 , n18181 , n18182 , n18183 , n18184 , n18185 , n18186 , n18187 , n18188 , n18189 , n18190 , n18191 , n18192 , n18193 , n18194 , n18195 , n18196 , n18197 , n18198 , n18199 , n18200 , n18201 , n18202 , n18203 , n18204 , n18205 , n18206 , n18207 , n18208 , n18209 , n18210 , n18211 , n18212 , n18213 , n18214 , n18215 , n18216 , n18217 , n18218 , n18219 , n18220 , n18221 , n18222 , n18223 , n18224 , n18225 , n18226 , n18227 , n18228 , n18229 , n18230 , n18231 , n18232 , n18233 , n18234 , n18235 , n18236 , n18237 , n18238 , n18239 , n18240 , n18241 , n18242 , n18243 , n18244 , n18245 , n18246 , n18247 , n18248 , n18249 , n18250 , n18251 , n18252 , n18253 , n18254 , n18255 , n18256 , n18257 , n18258 , n18259 , n18260 , n18261 , n18262 , n18263 , n18264 , n18265 , n18266 , n18267 , n18268 , n18269 , n18270 , n18271 , n18272 , n18273 , n18274 , n18275 , n18276 , n18277 , n18278 , n18279 , n18280 , n18281 , n18282 , n18283 , n18284 , n18285 , n18286 , n18287 , n18288 , n18289 , n18290 , n18291 , n18292 , n18293 , n18294 , n18295 , n18296 , n18297 , n18298 , n18299 , n18300 , n18301 , n18302 , n18303 , n18304 , n18305 , n18306 , n18307 , n18308 , n18309 , n18310 , n18311 , n18312 , n18313 , n18314 , n18315 , n18316 , n18317 , n18318 , n18319 , n18320 , n18321 , n18322 , n18323 , n18324 , n18325 , n18326 , n18327 , n18328 , n18329 , n18330 , n18331 , n18332 , n18333 , n18334 , n18335 , n18336 , n18337 , n18338 , n18339 , n18340 , n18341 , n18342 , n18343 , n18344 , n18345 , n18346 , n18347 , n18348 , n18349 , n18350 , n18351 , n18352 , n18353 , n18354 , n18355 , n18356 , n18357 , n18358 , n18359 , n18360 , n18361 , n18362 , n18363 , n18364 , n18365 , n18366 , n18367 , n18368 , n18369 , n18370 , n18371 , n18372 , n18373 , n18374 , n18375 , n18376 , n18377 , n18378 , n18379 , n18380 , n18381 , n18382 , n18383 , n18384 , n18385 , n18386 , n18387 , n18388 , n18389 , n18390 , n18391 , n18392 , n18393 , n18394 , n18395 , n18396 , n18397 , n18398 , n18399 , n18400 , n18401 , n18402 , n18403 , n18404 , n18405 , n18406 , n18407 , n18408 , n18409 , n18410 , n18411 , n18412 , n18413 , n18414 , n18415 , n18416 , n18417 , n18418 , n18419 , n18420 , n18421 , n18422 , n18423 , n18424 , n18425 , n18426 , n18427 , n18428 , n18429 , n18430 , n18431 , n18432 , n18433 , n18434 , n18435 , n18436 , n18437 , n18438 , n18439 , n18440 , n18441 , n18442 , n18443 , n18444 , n18445 , n18446 , n18447 , n18448 , n18449 , n18450 , n18451 , n18452 , n18453 , n18454 , n18455 , n18456 , n18457 , n18458 , n18459 , n18460 , n18461 , n18462 , n18463 , n18464 , n18465 , n18466 , n18467 , n18468 , n18469 , n18470 , n18471 , n18472 , n18473 , n18474 , n18475 , n18476 , n18477 , n18478 , n18479 , n18480 , n18481 , n18482 , n18483 , n18484 , n18485 , n18486 , n18487 , n18488 , n18489 , n18490 , n18491 , n18492 , n18493 , n18494 , n18495 , n18496 , n18497 , n18498 , n18499 , n18500 , n18501 , n18502 , n18503 , n18504 , n18505 , n18506 , n18507 , n18508 , n18509 , n18510 , n18511 , n18512 , n18513 , n18514 , n18515 , n18516 , n18517 , n18518 , n18519 , n18520 , n18521 , n18522 , n18523 , n18524 , n18525 , n18526 , n18527 , n18528 , n18529 , n18530 , n18531 , n18532 , n18533 , n18534 , n18535 , n18536 , n18537 , n18538 , n18539 , n18540 , n18541 , n18542 , n18543 , n18544 , n18545 , n18546 , n18547 , n18548 , n18549 , n18550 , n18551 , n18552 , n18553 , n18554 , n18555 , n18556 , n18557 , n18558 , n18559 , n18560 , n18561 , n18562 , n18563 , n18564 , n18565 , n18566 , n18567 , n18568 , n18569 , n18570 , n18571 , n18572 , n18573 , n18574 , n18575 , n18576 , n18577 , n18578 , n18579 , n18580 , n18581 , n18582 , n18583 , n18584 , n18585 , n18586 , n18587 , n18588 , n18589 , n18590 , n18591 , n18592 , n18593 , n18594 , n18595 , n18596 , n18597 , n18598 , n18599 , n18600 , n18601 , n18602 , n18603 , n18604 , n18605 , n18606 , n18607 , n18608 , n18609 , n18610 , n18611 , n18612 , n18613 , n18614 , n18615 , n18616 , n18617 , n18618 , n18619 , n18620 , n18621 , n18622 , n18623 , n18624 , n18625 , n18626 , n18627 , n18628 , n18629 , n18630 , n18631 , n18632 , n18633 , n18634 , n18635 , n18636 , n18637 , n18638 , n18639 , n18640 , n18641 , n18642 , n18643 , n18644 , n18645 , n18646 , n18647 , n18648 , n18649 , n18650 , n18651 , n18652 , n18653 , n18654 , n18655 , n18656 , n18657 , n18658 , n18659 , n18660 , n18661 , n18662 , n18663 , n18664 , n18665 , n18666 , n18667 , n18668 , n18669 , n18670 , n18671 , n18672 , n18673 , n18674 , n18675 , n18676 , n18677 , n18678 , n18679 , n18680 , n18681 , n18682 , n18683 , n18684 , n18685 , n18686 , n18687 , n18688 , n18689 , n18690 , n18691 , n18692 , n18693 , n18694 , n18695 , n18696 , n18697 , n18698 , n18699 , n18700 , n18701 , n18702 , n18703 , n18704 , n18705 , n18706 , n18707 , n18708 , n18709 , n18710 , n18711 , n18712 , n18713 , n18714 , n18715 , n18716 , n18717 , n18718 , n18719 , n18720 , n18721 , n18722 , n18723 , n18724 , n18725 , n18726 , n18727 , n18728 , n18729 , n18730 , n18731 , n18732 , n18733 , n18734 , n18735 , n18736 , n18737 , n18738 , n18739 , n18740 , n18741 , n18742 , n18743 , n18744 , n18745 , n18746 , n18747 , n18748 , n18749 , n18750 , n18751 , n18752 , n18753 , n18754 , n18755 , n18756 , n18757 , n18758 , n18759 , n18760 , n18761 , n18762 , n18763 , n18764 , n18765 , n18766 , n18767 , n18768 , n18769 , n18770 , n18771 , n18772 , n18773 , n18774 , n18775 , n18776 , n18777 , n18778 , n18779 , n18780 , n18781 , n18782 , n18783 , n18784 , n18785 , n18786 , n18787 , n18788 , n18789 , n18790 , n18791 , n18792 , n18793 , n18794 , n18795 , n18796 , n18797 , n18798 , n18799 , n18800 , n18801 , n18802 , n18803 , n18804 , n18805 , n18806 , n18807 , n18808 , n18809 , n18810 , n18811 , n18812 , n18813 , n18814 , n18815 , n18816 , n18817 , n18818 , n18819 , n18820 , n18821 , n18822 , n18823 , n18824 , n18825 , n18826 , n18827 , n18828 , n18829 , n18830 , n18831 , n18832 , n18833 , n18834 , n18835 , n18836 , n18837 , n18838 , n18839 , n18840 , n18841 , n18842 , n18843 , n18844 , n18845 , n18846 , n18847 , n18848 , n18849 , n18850 , n18851 , n18852 , n18853 , n18854 , n18855 , n18856 , n18857 , n18858 , n18859 , n18860 , n18861 , n18862 , n18863 , n18864 , n18865 , n18866 , n18867 , n18868 , n18869 , n18870 , n18871 , n18872 , n18873 , n18874 , n18875 , n18876 , n18877 , n18878 , n18879 , n18880 , n18881 , n18882 , n18883 , n18884 , n18885 , n18886 , n18887 , n18888 , n18889 , n18890 , n18891 , n18892 , n18893 , n18894 , n18895 , n18896 , n18897 , n18898 , n18899 , n18900 , n18901 , n18902 , n18903 , n18904 , n18905 , n18906 , n18907 , n18908 , n18909 , n18910 , n18911 , n18912 , n18913 , n18914 , n18915 , n18916 , n18917 , n18918 , n18919 , n18920 , n18921 , n18922 , n18923 , n18924 , n18925 , n18926 , n18927 , n18928 , n18929 , n18930 , n18931 , n18932 , n18933 , n18934 , n18935 , n18936 , n18937 , n18938 , n18939 , n18940 , n18941 , n18942 , n18943 , n18944 , n18945 , n18946 , n18947 , n18948 , n18949 , n18950 , n18951 , n18952 , n18953 , n18954 , n18955 , n18956 , n18957 , n18958 , n18959 , n18960 , n18961 , n18962 , n18963 , n18964 , n18965 , n18966 , n18967 , n18968 , n18969 , n18970 , n18971 , n18972 , n18973 , n18974 , n18975 , n18976 , n18977 , n18978 , n18979 , n18980 , n18981 , n18982 , n18983 , n18984 , n18985 , n18986 , n18987 , n18988 , n18989 , n18990 , n18991 , n18992 , n18993 , n18994 , n18995 , n18996 , n18997 , n18998 , n18999 , n19000 , n19001 , n19002 , n19003 , n19004 , n19005 , n19006 , n19007 , n19008 , n19009 , n19010 , n19011 , n19012 , n19013 , n19014 , n19015 , n19016 , n19017 , n19018 , n19019 , n19020 , n19021 , n19022 , n19023 , n19024 , n19025 , n19026 , n19027 , n19028 , n19029 , n19030 , n19031 , n19032 , n19033 , n19034 , n19035 , n19036 , n19037 , n19038 , n19039 , n19040 , n19041 , n19042 , n19043 , n19044 , n19045 , n19046 , n19047 , n19048 , n19049 , n19050 , n19051 , n19052 , n19053 , n19054 , n19055 , n19056 , n19057 , n19058 , n19059 , n19060 , n19061 , n19062 , n19063 , n19064 , n19065 , n19066 , n19067 , n19068 , n19069 , n19070 , n19071 , n19072 , n19073 , n19074 , n19075 , n19076 , n19077 , n19078 , n19079 , n19080 , n19081 , n19082 , n19083 , n19084 , n19085 , n19086 , n19087 , n19088 , n19089 , n19090 , n19091 , n19092 , n19093 , n19094 , n19095 , n19096 , n19097 , n19098 , n19099 , n19100 , n19101 , n19102 , n19103 , n19104 , n19105 , n19106 , n19107 , n19108 , n19109 , n19110 , n19111 , n19112 , n19113 , n19114 , n19115 , n19116 , n19117 , n19118 , n19119 , n19120 , n19121 , n19122 , n19123 , n19124 , n19125 , n19126 , n19127 , n19128 , n19129 , n19130 , n19131 , n19132 , n19133 , n19134 , n19135 , n19136 , n19137 , n19138 , n19139 , n19140 , n19141 , n19142 , n19143 , n19144 , n19145 , n19146 , n19147 , n19148 , n19149 , n19150 , n19151 , n19152 , n19153 , n19154 , n19155 , n19156 , n19157 , n19158 , n19159 , n19160 , n19161 , n19162 , n19163 , n19164 , n19165 , n19166 , n19167 , n19168 , n19169 , n19170 , n19171 , n19172 , n19173 , n19174 , n19175 , n19176 , n19177 , n19178 , n19179 , n19180 , n19181 , n19182 , n19183 , n19184 , n19185 , n19186 , n19187 , n19188 , n19189 , n19190 , n19191 , n19192 , n19193 , n19194 , n19195 , n19196 , n19197 , n19198 , n19199 , n19200 , n19201 , n19202 , n19203 , n19204 , n19205 , n19206 , n19207 , n19208 , n19209 , n19210 , n19211 , n19212 , n19213 , n19214 , n19215 , n19216 , n19217 , n19218 , n19219 , n19220 , n19221 , n19222 , n19223 , n19224 , n19225 , n19226 , n19227 , n19228 , n19229 , n19230 , n19231 , n19232 , n19233 , n19234 , n19235 , n19236 , n19237 , n19238 , n19239 , n19240 , n19241 , n19242 , n19243 , n19244 , n19245 , n19246 , n19247 , n19248 , n19249 , n19250 , n19251 , n19252 , n19253 , n19254 , n19255 , n19256 , n19257 , n19258 , n19259 , n19260 , n19261 , n19262 , n19263 , n19264 , n19265 , n19266 , n19267 , n19268 , n19269 , n19270 , n19271 , n19272 , n19273 , n19274 , n19275 , n19276 , n19277 , n19278 , n19279 , n19280 , n19281 , n19282 , n19283 , n19284 , n19285 , n19286 , n19287 , n19288 , n19289 , n19290 , n19291 , n19292 , n19293 , n19294 , n19295 , n19296 , n19297 , n19298 , n19299 , n19300 , n19301 , n19302 , n19303 , n19304 , n19305 , n19306 , n19307 , n19308 , n19309 , n19310 , n19311 , n19312 , n19313 , n19314 , n19315 , n19316 , n19317 , n19318 , n19319 , n19320 , n19321 , n19322 , n19323 , n19324 , n19325 , n19326 , n19327 , n19328 , n19329 , n19330 , n19331 , n19332 , n19333 , n19334 , n19335 , n19336 , n19337 , n19338 , n19339 , n19340 , n19341 , n19342 , n19343 , n19344 , n19345 , n19346 , n19347 , n19348 , n19349 , n19350 , n19351 , n19352 , n19353 , n19354 , n19355 , n19356 , n19357 , n19358 , n19359 , n19360 , n19361 , n19362 , n19363 , n19364 , n19365 , n19366 , n19367 , n19368 , n19369 , n19370 , n19371 , n19372 , n19373 , n19374 , n19375 , n19376 , n19377 , n19378 , n19379 , n19380 , n19381 , n19382 , n19383 , n19384 , n19385 , n19386 , n19387 , n19388 , n19389 , n19390 , n19391 , n19392 , n19393 , n19394 , n19395 , n19396 , n19397 , n19398 , n19399 , n19400 , n19401 , n19402 , n19403 , n19404 , n19405 , n19406 , n19407 , n19408 , n19409 , n19410 , n19411 , n19412 , n19413 , n19414 , n19415 , n19416 , n19417 , n19418 , n19419 , n19420 , n19421 , n19422 , n19423 , n19424 , n19425 , n19426 , n19427 , n19428 , n19429 , n19430 , n19431 , n19432 , n19433 , n19434 , n19435 , n19436 , n19437 , n19438 , n19439 , n19440 , n19441 , n19442 , n19443 , n19444 , n19445 , n19446 , n19447 , n19448 , n19449 , n19450 , n19451 , n19452 , n19453 , n19454 , n19455 , n19456 , n19457 , n19458 , n19459 , n19460 , n19461 , n19462 , n19463 , n19464 , n19465 , n19466 , n19467 , n19468 , n19469 , n19470 , n19471 , n19472 , n19473 , n19474 , n19475 , n19476 , n19477 , n19478 , n19479 , n19480 , n19481 , n19482 , n19483 , n19484 , n19485 , n19486 , n19487 , n19488 , n19489 , n19490 , n19491 , n19492 , n19493 , n19494 , n19495 , n19496 , n19497 , n19498 , n19499 , n19500 , n19501 , n19502 , n19503 , n19504 , n19505 , n19506 , n19507 , n19508 , n19509 , n19510 , n19511 , n19512 , n19513 , n19514 , n19515 , n19516 , n19517 , n19518 , n19519 , n19520 , n19521 , n19522 , n19523 , n19524 , n19525 , n19526 , n19527 , n19528 , n19529 , n19530 , n19531 , n19532 , n19533 , n19534 , n19535 , n19536 , n19537 , n19538 , n19539 , n19540 , n19541 , n19542 , n19543 , n19544 , n19545 , n19546 , n19547 , n19548 , n19549 , n19550 , n19551 , n19552 , n19553 , n19554 , n19555 , n19556 , n19557 , n19558 , n19559 , n19560 , n19561 , n19562 , n19563 , n19564 , n19565 , n19566 , n19567 , n19568 , n19569 , n19570 , n19571 , n19572 , n19573 , n19574 , n19575 , n19576 , n19577 , n19578 , n19579 , n19580 , n19581 , n19582 , n19583 , n19584 , n19585 , n19586 , n19587 , n19588 , n19589 , n19590 , n19591 , n19592 , n19593 , n19594 , n19595 , n19596 , n19597 , n19598 , n19599 , n19600 , n19601 , n19602 , n19603 , n19604 , n19605 , n19606 , n19607 , n19608 , n19609 , n19610 , n19611 , n19612 , n19613 , n19614 , n19615 , n19616 , n19617 , n19618 , n19619 , n19620 , n19621 , n19622 , n19623 , n19624 , n19625 , n19626 , n19627 , n19628 , n19629 , n19630 , n19631 , n19632 , n19633 , n19634 , n19635 , n19636 , n19637 , n19638 , n19639 , n19640 , n19641 , n19642 , n19643 , n19644 , n19645 , n19646 , n19647 , n19648 , n19649 , n19650 , n19651 , n19652 , n19653 , n19654 , n19655 , n19656 , n19657 , n19658 , n19659 , n19660 , n19661 , n19662 , n19663 , n19664 , n19665 , n19666 , n19667 , n19668 , n19669 , n19670 , n19671 , n19672 , n19673 , n19674 , n19675 , n19676 , n19677 , n19678 , n19679 , n19680 , n19681 , n19682 , n19683 , n19684 , n19685 , n19686 , n19687 , n19688 , n19689 , n19690 , n19691 , n19692 , n19693 , n19694 , n19695 , n19696 , n19697 , n19698 , n19699 , n19700 , n19701 , n19702 , n19703 , n19704 , n19705 , n19706 , n19707 , n19708 , n19709 , n19710 , n19711 , n19712 , n19713 , n19714 , n19715 , n19716 , n19717 , n19718 , n19719 , n19720 , n19721 , n19722 , n19723 , n19724 , n19725 , n19726 , n19727 , n19728 , n19729 , n19730 , n19731 , n19732 , n19733 , n19734 , n19735 , n19736 , n19737 , n19738 , n19739 , n19740 , n19741 , n19742 , n19743 , n19744 , n19745 , n19746 , n19747 , n19748 , n19749 , n19750 , n19751 , n19752 , n19753 , n19754 , n19755 , n19756 , n19757 , n19758 , n19759 , n19760 , n19761 , n19762 , n19763 , n19764 , n19765 , n19766 , n19767 , n19768 , n19769 , n19770 , n19771 , n19772 , n19773 , n19774 , n19775 , n19776 , n19777 , n19778 , n19779 , n19780 , n19781 , n19782 , n19783 , n19784 , n19785 , n19786 , n19787 , n19788 , n19789 , n19790 , n19791 , n19792 , n19793 , n19794 , n19795 , n19796 , n19797 , n19798 , n19799 , n19800 , n19801 , n19802 , n19803 , n19804 , n19805 , n19806 , n19807 , n19808 , n19809 , n19810 , n19811 , n19812 , n19813 , n19814 , n19815 , n19816 , n19817 , n19818 , n19819 , n19820 , n19821 , n19822 , n19823 , n19824 , n19825 , n19826 , n19827 , n19828 , n19829 , n19830 , n19831 , n19832 , n19833 , n19834 , n19835 , n19836 , n19837 , n19838 , n19839 , n19840 , n19841 , n19842 , n19843 , n19844 , n19845 , n19846 , n19847 , n19848 , n19849 , n19850 , n19851 , n19852 , n19853 , n19854 , n19855 , n19856 , n19857 , n19858 , n19859 , n19860 , n19861 , n19862 , n19863 , n19864 , n19865 , n19866 , n19867 , n19868 , n19869 , n19870 , n19871 , n19872 , n19873 , n19874 , n19875 , n19876 , n19877 , n19878 , n19879 , n19880 , n19881 , n19882 , n19883 , n19884 , n19885 , n19886 , n19887 , n19888 , n19889 , n19890 , n19891 , n19892 , n19893 , n19894 , n19895 , n19896 , n19897 , n19898 , n19899 , n19900 , n19901 , n19902 , n19903 , n19904 , n19905 , n19906 , n19907 , n19908 , n19909 , n19910 , n19911 , n19912 , n19913 , n19914 , n19915 , n19916 , n19917 , n19918 , n19919 , n19920 , n19921 , n19922 , n19923 , n19924 , n19925 , n19926 , n19927 , n19928 , n19929 , n19930 , n19931 , n19932 , n19933 , n19934 , n19935 , n19936 , n19937 , n19938 , n19939 , n19940 , n19941 , n19942 , n19943 , n19944 , n19945 , n19946 , n19947 , n19948 , n19949 , n19950 , n19951 , n19952 , n19953 , n19954 , n19955 , n19956 , n19957 , n19958 , n19959 , n19960 , n19961 , n19962 , n19963 , n19964 , n19965 , n19966 , n19967 , n19968 , n19969 , n19970 , n19971 , n19972 , n19973 , n19974 , n19975 , n19976 , n19977 , n19978 , n19979 , n19980 , n19981 , n19982 , n19983 , n19984 , n19985 , n19986 , n19987 , n19988 , n19989 , n19990 , n19991 , n19992 , n19993 , n19994 , n19995 , n19996 , n19997 , n19998 , n19999 , n20000 , n20001 , n20002 , n20003 , n20004 , n20005 , n20006 , n20007 , n20008 , n20009 , n20010 , n20011 , n20012 , n20013 , n20014 , n20015 , n20016 , n20017 , n20018 , n20019 , n20020 , n20021 , n20022 , n20023 , n20024 , n20025 , n20026 , n20027 , n20028 , n20029 , n20030 , n20031 , n20032 , n20033 , n20034 , n20035 , n20036 , n20037 , n20038 , n20039 , n20040 , n20041 , n20042 , n20043 , n20044 , n20045 , n20046 , n20047 , n20048 , n20049 , n20050 , n20051 , n20052 , n20053 , n20054 , n20055 , n20056 , n20057 , n20058 , n20059 , n20060 , n20061 , n20062 , n20063 , n20064 , n20065 , n20066 , n20067 , n20068 , n20069 , n20070 , n20071 , n20072 , n20073 , n20074 , n20075 , n20076 , n20077 , n20078 , n20079 , n20080 , n20081 , n20082 , n20083 , n20084 , n20085 , n20086 , n20087 , n20088 , n20089 , n20090 , n20091 , n20092 , n20093 , n20094 , n20095 , n20096 , n20097 , n20098 , n20099 , n20100 , n20101 , n20102 , n20103 , n20104 , n20105 , n20106 , n20107 , n20108 , n20109 , n20110 , n20111 , n20112 , n20113 , n20114 , n20115 , n20116 , n20117 , n20118 , n20119 , n20120 , n20121 , n20122 , n20123 , n20124 , n20125 , n20126 , n20127 , n20128 , n20129 , n20130 , n20131 , n20132 , n20133 , n20134 , n20135 , n20136 , n20137 , n20138 , n20139 , n20140 , n20141 , n20142 , n20143 , n20144 , n20145 , n20146 , n20147 , n20148 , n20149 , n20150 , n20151 , n20152 , n20153 , n20154 , n20155 , n20156 , n20157 , n20158 , n20159 , n20160 , n20161 , n20162 , n20163 , n20164 , n20165 , n20166 , n20167 , n20168 , n20169 , n20170 , n20171 , n20172 , n20173 , n20174 , n20175 , n20176 , n20177 , n20178 , n20179 , n20180 , n20181 , n20182 , n20183 , n20184 , n20185 , n20186 , n20187 , n20188 , n20189 , n20190 , n20191 , n20192 , n20193 , n20194 , n20195 , n20196 , n20197 , n20198 , n20199 , n20200 , n20201 , n20202 , n20203 , n20204 , n20205 , n20206 , n20207 , n20208 , n20209 , n20210 , n20211 , n20212 , n20213 , n20214 , n20215 , n20216 , n20217 , n20218 , n20219 , n20220 , n20221 , n20222 , n20223 , n20224 , n20225 , n20226 , n20227 , n20228 , n20229 , n20230 , n20231 , n20232 , n20233 , n20234 , n20235 , n20236 , n20237 , n20238 , n20239 , n20240 , n20241 , n20242 , n20243 , n20244 , n20245 , n20246 , n20247 , n20248 , n20249 , n20250 , n20251 , n20252 , n20253 , n20254 , n20255 , n20256 , n20257 , n20258 , n20259 , n20260 , n20261 , n20262 , n20263 , n20264 , n20265 , n20266 , n20267 , n20268 , n20269 , n20270 , n20271 , n20272 , n20273 , n20274 , n20275 , n20276 , n20277 , n20278 , n20279 , n20280 , n20281 , n20282 , n20283 , n20284 , n20285 , n20286 , n20287 , n20288 , n20289 , n20290 , n20291 , n20292 , n20293 , n20294 , n20295 , n20296 , n20297 , n20298 , n20299 , n20300 , n20301 , n20302 , n20303 , n20304 , n20305 , n20306 , n20307 , n20308 , n20309 , n20310 , n20311 , n20312 , n20313 , n20314 , n20315 , n20316 , n20317 , n20318 , n20319 , n20320 , n20321 , n20322 , n20323 , n20324 , n20325 , n20326 , n20327 , n20328 , n20329 , n20330 , n20331 , n20332 , n20333 , n20334 , n20335 , n20336 , n20337 , n20338 , n20339 , n20340 , n20341 , n20342 , n20343 , n20344 , n20345 , n20346 , n20347 , n20348 , n20349 , n20350 , n20351 , n20352 , n20353 , n20354 , n20355 , n20356 , n20357 , n20358 , n20359 , n20360 , n20361 , n20362 , n20363 , n20364 , n20365 , n20366 , n20367 , n20368 , n20369 , n20370 , n20371 , n20372 , n20373 , n20374 , n20375 , n20376 , n20377 , n20378 , n20379 , n20380 , n20381 , n20382 , n20383 , n20384 , n20385 , n20386 , n20387 , n20388 , n20389 , n20390 , n20391 , n20392 , n20393 , n20394 , n20395 , n20396 , n20397 , n20398 , n20399 , n20400 , n20401 , n20402 , n20403 , n20404 , n20405 , n20406 , n20407 , n20408 , n20409 , n20410 , n20411 , n20412 , n20413 , n20414 , n20415 , n20416 , n20417 , n20418 , n20419 , n20420 , n20421 , n20422 , n20423 , n20424 , n20425 , n20426 , n20427 , n20428 , n20429 , n20430 , n20431 , n20432 , n20433 , n20434 , n20435 , n20436 , n20437 , n20438 , n20439 , n20440 , n20441 , n20442 , n20443 , n20444 , n20445 , n20446 , n20447 , n20448 , n20449 , n20450 , n20451 , n20452 , n20453 , n20454 , n20455 , n20456 , n20457 , n20458 , n20459 , n20460 , n20461 , n20462 , n20463 , n20464 , n20465 , n20466 , n20467 , n20468 , n20469 , n20470 , n20471 , n20472 , n20473 , n20474 , n20475 , n20476 , n20477 , n20478 , n20479 , n20480 , n20481 , n20482 , n20483 , n20484 , n20485 , n20486 , n20487 , n20488 , n20489 , n20490 , n20491 , n20492 , n20493 , n20494 , n20495 , n20496 , n20497 , n20498 , n20499 , n20500 , n20501 , n20502 , n20503 , n20504 , n20505 , n20506 , n20507 , n20508 , n20509 , n20510 , n20511 , n20512 , n20513 , n20514 , n20515 , n20516 , n20517 , n20518 , n20519 , n20520 , n20521 , n20522 , n20523 , n20524 , n20525 , n20526 , n20527 , n20528 , n20529 , n20530 , n20531 , n20532 , n20533 , n20534 , n20535 , n20536 , n20537 , n20538 , n20539 , n20540 , n20541 , n20542 , n20543 , n20544 , n20545 , n20546 , n20547 , n20548 , n20549 , n20550 , n20551 , n20552 , n20553 , n20554 , n20555 , n20556 , n20557 , n20558 , n20559 , n20560 , n20561 , n20562 , n20563 , n20564 , n20565 , n20566 , n20567 , n20568 , n20569 , n20570 , n20571 , n20572 , n20573 , n20574 , n20575 , n20576 , n20577 , n20578 , n20579 , n20580 , n20581 , n20582 , n20583 , n20584 , n20585 , n20586 , n20587 , n20588 , n20589 , n20590 , n20591 , n20592 , n20593 , n20594 , n20595 , n20596 , n20597 , n20598 , n20599 , n20600 , n20601 , n20602 , n20603 , n20604 , n20605 , n20606 , n20607 , n20608 , n20609 , n20610 , n20611 , n20612 , n20613 , n20614 , n20615 , n20616 , n20617 , n20618 , n20619 , n20620 , n20621 , n20622 , n20623 , n20624 , n20625 , n20626 , n20627 , n20628 , n20629 , n20630 , n20631 , n20632 , n20633 , n20634 , n20635 , n20636 , n20637 , n20638 , n20639 , n20640 , n20641 , n20642 , n20643 , n20644 , n20645 , n20646 , n20647 , n20648 , n20649 , n20650 , n20651 , n20652 , n20653 , n20654 , n20655 , n20656 , n20657 , n20658 , n20659 , n20660 , n20661 , n20662 , n20663 , n20664 , n20665 , n20666 , n20667 , n20668 , n20669 , n20670 , n20671 , n20672 , n20673 , n20674 , n20675 , n20676 , n20677 , n20678 , n20679 , n20680 , n20681 , n20682 , n20683 , n20684 , n20685 , n20686 , n20687 , n20688 , n20689 , n20690 , n20691 , n20692 , n20693 , n20694 , n20695 , n20696 , n20697 , n20698 , n20699 , n20700 , n20701 , n20702 , n20703 , n20704 , n20705 , n20706 , n20707 , n20708 , n20709 , n20710 , n20711 , n20712 , n20713 , n20714 , n20715 , n20716 , n20717 , n20718 , n20719 , n20720 , n20721 , n20722 , n20723 , n20724 , n20725 , n20726 , n20727 , n20728 , n20729 , n20730 , n20731 , n20732 , n20733 , n20734 , n20735 , n20736 , n20737 , n20738 , n20739 , n20740 , n20741 , n20742 , n20743 , n20744 , n20745 , n20746 , n20747 , n20748 , n20749 , n20750 , n20751 , n20752 , n20753 , n20754 , n20755 , n20756 , n20757 , n20758 , n20759 , n20760 , n20761 , n20762 , n20763 , n20764 , n20765 , n20766 , n20767 , n20768 , n20769 , n20770 , n20771 , n20772 , n20773 , n20774 , n20775 , n20776 , n20777 , n20778 , n20779 , n20780 , n20781 , n20782 , n20783 , n20784 , n20785 , n20786 , n20787 , n20788 , n20789 , n20790 , n20791 , n20792 , n20793 , n20794 , n20795 , n20796 , n20797 , n20798 , n20799 , n20800 , n20801 , n20802 , n20803 , n20804 , n20805 , n20806 , n20807 , n20808 , n20809 , n20810 , n20811 , n20812 , n20813 , n20814 , n20815 , n20816 , n20817 , n20818 , n20819 , n20820 , n20821 , n20822 , n20823 , n20824 , n20825 , n20826 , n20827 , n20828 , n20829 , n20830 , n20831 , n20832 , n20833 , n20834 , n20835 , n20836 , n20837 , n20838 , n20839 , n20840 , n20841 , n20842 , n20843 , n20844 , n20845 , n20846 , n20847 , n20848 , n20849 , n20850 , n20851 , n20852 , n20853 , n20854 , n20855 , n20856 , n20857 , n20858 , n20859 , n20860 , n20861 , n20862 , n20863 , n20864 , n20865 , n20866 , n20867 , n20868 , n20869 , n20870 , n20871 , n20872 , n20873 , n20874 , n20875 , n20876 , n20877 , n20878 , n20879 , n20880 , n20881 , n20882 , n20883 , n20884 , n20885 , n20886 , n20887 , n20888 , n20889 , n20890 , n20891 , n20892 , n20893 , n20894 , n20895 , n20896 , n20897 , n20898 , n20899 , n20900 , n20901 , n20902 , n20903 , n20904 , n20905 , n20906 , n20907 , n20908 , n20909 , n20910 , n20911 , n20912 , n20913 , n20914 , n20915 , n20916 , n20917 , n20918 , n20919 , n20920 , n20921 , n20922 , n20923 , n20924 , n20925 , n20926 , n20927 , n20928 , n20929 , n20930 , n20931 , n20932 , n20933 , n20934 , n20935 , n20936 , n20937 , n20938 , n20939 , n20940 , n20941 , n20942 , n20943 , n20944 , n20945 , n20946 , n20947 , n20948 , n20949 , n20950 , n20951 , n20952 , n20953 , n20954 , n20955 , n20956 , n20957 , n20958 , n20959 , n20960 , n20961 , n20962 , n20963 , n20964 , n20965 , n20966 , n20967 , n20968 , n20969 , n20970 , n20971 , n20972 , n20973 , n20974 , n20975 , n20976 , n20977 , n20978 , n20979 , n20980 , n20981 , n20982 , n20983 , n20984 , n20985 , n20986 , n20987 , n20988 , n20989 , n20990 , n20991 , n20992 , n20993 , n20994 , n20995 , n20996 , n20997 , n20998 , n20999 , n21000 , n21001 , n21002 , n21003 , n21004 , n21005 , n21006 , n21007 , n21008 , n21009 , n21010 , n21011 , n21012 , n21013 , n21014 , n21015 , n21016 , n21017 , n21018 , n21019 , n21020 , n21021 , n21022 , n21023 , n21024 , n21025 , n21026 , n21027 , n21028 , n21029 , n21030 , n21031 , n21032 , n21033 , n21034 , n21035 , n21036 , n21037 , n21038 , n21039 , n21040 , n21041 , n21042 , n21043 , n21044 , n21045 , n21046 , n21047 , n21048 , n21049 , n21050 , n21051 , n21052 , n21053 , n21054 , n21055 , n21056 , n21057 , n21058 , n21059 , n21060 , n21061 , n21062 , n21063 , n21064 , n21065 , n21066 , n21067 , n21068 , n21069 , n21070 , n21071 , n21072 , n21073 , n21074 , n21075 , n21076 , n21077 , n21078 , n21079 , n21080 , n21081 , n21082 , n21083 , n21084 , n21085 , n21086 , n21087 , n21088 , n21089 , n21090 , n21091 , n21092 , n21093 , n21094 , n21095 , n21096 , n21097 , n21098 , n21099 , n21100 , n21101 , n21102 , n21103 , n21104 , n21105 , n21106 , n21107 , n21108 , n21109 , n21110 , n21111 , n21112 , n21113 , n21114 , n21115 , n21116 , n21117 , n21118 , n21119 , n21120 , n21121 , n21122 , n21123 , n21124 , n21125 , n21126 , n21127 , n21128 , n21129 , n21130 , n21131 , n21132 , n21133 , n21134 , n21135 , n21136 , n21137 , n21138 , n21139 , n21140 , n21141 , n21142 , n21143 , n21144 , n21145 , n21146 , n21147 , n21148 , n21149 , n21150 , n21151 , n21152 , n21153 , n21154 , n21155 , n21156 , n21157 , n21158 , n21159 , n21160 , n21161 , n21162 , n21163 , n21164 , n21165 , n21166 , n21167 , n21168 , n21169 , n21170 , n21171 , n21172 , n21173 , n21174 , n21175 , n21176 , n21177 , n21178 , n21179 , n21180 , n21181 , n21182 , n21183 , n21184 , n21185 , n21186 , n21187 , n21188 , n21189 , n21190 , n21191 , n21192 , n21193 , n21194 , n21195 , n21196 , n21197 , n21198 , n21199 , n21200 , n21201 , n21202 , n21203 , n21204 , n21205 , n21206 , n21207 , n21208 , n21209 , n21210 , n21211 , n21212 , n21213 , n21214 , n21215 , n21216 , n21217 , n21218 , n21219 , n21220 , n21221 , n21222 , n21223 , n21224 , n21225 , n21226 , n21227 , n21228 , n21229 , n21230 , n21231 , n21232 , n21233 , n21234 , n21235 , n21236 , n21237 , n21238 , n21239 , n21240 , n21241 , n21242 , n21243 , n21244 , n21245 , n21246 , n21247 , n21248 , n21249 , n21250 , n21251 , n21252 , n21253 , n21254 , n21255 , n21256 , n21257 , n21258 , n21259 , n21260 , n21261 , n21262 , n21263 , n21264 , n21265 , n21266 , n21267 , n21268 , n21269 , n21270 , n21271 , n21272 , n21273 , n21274 , n21275 , n21276 , n21277 , n21278 , n21279 , n21280 , n21281 , n21282 , n21283 , n21284 , n21285 , n21286 , n21287 , n21288 , n21289 , n21290 , n21291 , n21292 , n21293 , n21294 , n21295 , n21296 , n21297 , n21298 , n21299 , n21300 , n21301 , n21302 , n21303 , n21304 , n21305 , n21306 , n21307 , n21308 , n21309 , n21310 , n21311 , n21312 , n21313 , n21314 , n21315 , n21316 , n21317 , n21318 , n21319 , n21320 , n21321 , n21322 , n21323 , n21324 , n21325 , n21326 , n21327 , n21328 , n21329 , n21330 , n21331 , n21332 , n21333 , n21334 , n21335 , n21336 , n21337 , n21338 , n21339 , n21340 , n21341 , n21342 , n21343 , n21344 , n21345 , n21346 , n21347 , n21348 , n21349 , n21350 , n21351 , n21352 , n21353 , n21354 , n21355 , n21356 , n21357 , n21358 , n21359 , n21360 , n21361 , n21362 , n21363 , n21364 , n21365 , n21366 , n21367 , n21368 , n21369 , n21370 , n21371 , n21372 , n21373 , n21374 , n21375 , n21376 , n21377 , n21378 , n21379 , n21380 , n21381 , n21382 , n21383 , n21384 , n21385 , n21386 , n21387 , n21388 , n21389 , n21390 , n21391 , n21392 , n21393 , n21394 , n21395 , n21396 , n21397 , n21398 , n21399 , n21400 , n21401 , n21402 , n21403 , n21404 , n21405 , n21406 , n21407 , n21408 , n21409 , n21410 , n21411 , n21412 , n21413 , n21414 , n21415 , n21416 , n21417 , n21418 , n21419 , n21420 , n21421 , n21422 , n21423 , n21424 , n21425 , n21426 , n21427 , n21428 , n21429 , n21430 , n21431 , n21432 , n21433 , n21434 , n21435 , n21436 , n21437 , n21438 , n21439 , n21440 , n21441 , n21442 , n21443 , n21444 , n21445 , n21446 , n21447 , n21448 , n21449 , n21450 , n21451 , n21452 , n21453 , n21454 , n21455 , n21456 , n21457 , n21458 , n21459 , n21460 , n21461 , n21462 , n21463 , n21464 , n21465 , n21466 , n21467 , n21468 , n21469 , n21470 , n21471 , n21472 , n21473 , n21474 , n21475 , n21476 , n21477 , n21478 , n21479 , n21480 , n21481 , n21482 , n21483 , n21484 , n21485 , n21486 , n21487 , n21488 , n21489 , n21490 , n21491 , n21492 , n21493 , n21494 , n21495 , n21496 , n21497 , n21498 , n21499 , n21500 , n21501 , n21502 , n21503 , n21504 , n21505 , n21506 , n21507 , n21508 , n21509 , n21510 , n21511 , n21512 , n21513 , n21514 , n21515 , n21516 , n21517 , n21518 , n21519 , n21520 , n21521 , n21522 , n21523 , n21524 , n21525 , n21526 , n21527 , n21528 , n21529 , n21530 , n21531 , n21532 , n21533 , n21534 , n21535 , n21536 , n21537 , n21538 , n21539 , n21540 , n21541 , n21542 , n21543 , n21544 , n21545 , n21546 , n21547 , n21548 , n21549 , n21550 , n21551 , n21552 , n21553 , n21554 , n21555 , n21556 , n21557 , n21558 , n21559 , n21560 , n21561 , n21562 , n21563 , n21564 , n21565 , n21566 , n21567 , n21568 , n21569 , n21570 , n21571 , n21572 , n21573 , n21574 , n21575 , n21576 , n21577 , n21578 , n21579 , n21580 , n21581 , n21582 , n21583 , n21584 , n21585 , n21586 , n21587 , n21588 , n21589 , n21590 , n21591 , n21592 , n21593 , n21594 , n21595 , n21596 , n21597 , n21598 , n21599 , n21600 , n21601 , n21602 , n21603 , n21604 , n21605 , n21606 , n21607 , n21608 , n21609 , n21610 , n21611 , n21612 , n21613 , n21614 , n21615 , n21616 , n21617 , n21618 , n21619 , n21620 , n21621 , n21622 , n21623 , n21624 , n21625 , n21626 , n21627 , n21628 , n21629 , n21630 , n21631 , n21632 , n21633 , n21634 , n21635 , n21636 , n21637 , n21638 , n21639 , n21640 , n21641 , n21642 , n21643 , n21644 , n21645 , n21646 , n21647 , n21648 , n21649 , n21650 , n21651 , n21652 , n21653 , n21654 , n21655 , n21656 , n21657 , n21658 , n21659 , n21660 , n21661 , n21662 , n21663 , n21664 , n21665 , n21666 , n21667 , n21668 , n21669 , n21670 , n21671 , n21672 , n21673 , n21674 , n21675 , n21676 , n21677 , n21678 , n21679 , n21680 , n21681 , n21682 , n21683 , n21684 , n21685 , n21686 , n21687 , n21688 , n21689 , n21690 , n21691 , n21692 , n21693 , n21694 , n21695 , n21696 , n21697 , n21698 , n21699 , n21700 , n21701 , n21702 , n21703 , n21704 , n21705 , n21706 , n21707 , n21708 , n21709 , n21710 , n21711 , n21712 , n21713 , n21714 , n21715 , n21716 , n21717 , n21718 , n21719 , n21720 , n21721 , n21722 , n21723 , n21724 , n21725 , n21726 , n21727 , n21728 , n21729 , n21730 , n21731 , n21732 , n21733 , n21734 , n21735 , n21736 , n21737 , n21738 , n21739 , n21740 , n21741 , n21742 , n21743 , n21744 , n21745 , n21746 , n21747 , n21748 , n21749 , n21750 , n21751 , n21752 , n21753 , n21754 , n21755 , n21756 , n21757 , n21758 , n21759 , n21760 , n21761 , n21762 , n21763 , n21764 , n21765 , n21766 , n21767 , n21768 , n21769 , n21770 , n21771 , n21772 , n21773 , n21774 , n21775 , n21776 , n21777 , n21778 , n21779 , n21780 , n21781 , n21782 , n21783 , n21784 , n21785 , n21786 , n21787 , n21788 , n21789 , n21790 , n21791 , n21792 , n21793 , n21794 , n21795 , n21796 , n21797 , n21798 , n21799 , n21800 , n21801 , n21802 , n21803 , n21804 , n21805 , n21806 , n21807 , n21808 , n21809 , n21810 , n21811 , n21812 , n21813 , n21814 , n21815 , n21816 , n21817 , n21818 , n21819 , n21820 , n21821 , n21822 , n21823 , n21824 , n21825 , n21826 , n21827 , n21828 , n21829 , n21830 , n21831 , n21832 , n21833 , n21834 , n21835 , n21836 , n21837 , n21838 , n21839 , n21840 , n21841 , n21842 , n21843 , n21844 , n21845 , n21846 , n21847 , n21848 , n21849 , n21850 , n21851 , n21852 , n21853 , n21854 , n21855 , n21856 , n21857 , n21858 , n21859 , n21860 , n21861 , n21862 , n21863 , n21864 , n21865 , n21866 , n21867 , n21868 , n21869 , n21870 , n21871 , n21872 , n21873 , n21874 , n21875 , n21876 , n21877 , n21878 , n21879 , n21880 , n21881 , n21882 , n21883 , n21884 , n21885 , n21886 , n21887 , n21888 , n21889 , n21890 , n21891 , n21892 , n21893 , n21894 , n21895 , n21896 , n21897 , n21898 , n21899 , n21900 , n21901 , n21902 , n21903 , n21904 , n21905 , n21906 , n21907 , n21908 , n21909 , n21910 , n21911 , n21912 , n21913 , n21914 , n21915 , n21916 , n21917 , n21918 , n21919 , n21920 , n21921 , n21922 , n21923 , n21924 , n21925 , n21926 , n21927 , n21928 , n21929 , n21930 , n21931 , n21932 , n21933 , n21934 , n21935 , n21936 , n21937 , n21938 , n21939 , n21940 , n21941 , n21942 , n21943 , n21944 , n21945 , n21946 , n21947 , n21948 , n21949 , n21950 , n21951 , n21952 , n21953 , n21954 , n21955 , n21956 , n21957 , n21958 , n21959 , n21960 , n21961 , n21962 , n21963 , n21964 , n21965 , n21966 , n21967 , n21968 , n21969 , n21970 , n21971 , n21972 , n21973 , n21974 , n21975 , n21976 , n21977 , n21978 , n21979 , n21980 , n21981 , n21982 , n21983 , n21984 , n21985 , n21986 , n21987 , n21988 , n21989 , n21990 , n21991 , n21992 , n21993 , n21994 , n21995 , n21996 , n21997 , n21998 , n21999 , n22000 , n22001 , n22002 , n22003 , n22004 , n22005 , n22006 , n22007 , n22008 , n22009 , n22010 , n22011 , n22012 , n22013 , n22014 , n22015 , n22016 , n22017 , n22018 , n22019 , n22020 , n22021 , n22022 , n22023 , n22024 , n22025 , n22026 , n22027 , n22028 , n22029 , n22030 , n22031 , n22032 , n22033 , n22034 , n22035 , n22036 , n22037 , n22038 , n22039 , n22040 , n22041 , n22042 , n22043 , n22044 , n22045 , n22046 , n22047 , n22048 , n22049 , n22050 , n22051 , n22052 , n22053 , n22054 , n22055 , n22056 , n22057 , n22058 , n22059 , n22060 , n22061 , n22062 , n22063 , n22064 , n22065 , n22066 , n22067 , n22068 , n22069 , n22070 , n22071 , n22072 , n22073 , n22074 , n22075 , n22076 , n22077 , n22078 , n22079 , n22080 , n22081 , n22082 , n22083 , n22084 , n22085 , n22086 , n22087 , n22088 , n22089 , n22090 , n22091 , n22092 , n22093 , n22094 , n22095 , n22096 , n22097 , n22098 , n22099 , n22100 , n22101 , n22102 , n22103 , n22104 , n22105 , n22106 , n22107 , n22108 , n22109 , n22110 , n22111 , n22112 , n22113 , n22114 , n22115 , n22116 , n22117 , n22118 , n22119 , n22120 , n22121 , n22122 , n22123 , n22124 , n22125 , n22126 , n22127 , n22128 , n22129 , n22130 , n22131 , n22132 , n22133 , n22134 , n22135 , n22136 , n22137 , n22138 , n22139 , n22140 , n22141 , n22142 , n22143 , n22144 , n22145 , n22146 , n22147 , n22148 , n22149 , n22150 , n22151 , n22152 , n22153 , n22154 , n22155 , n22156 , n22157 , n22158 , n22159 , n22160 , n22161 , n22162 , n22163 , n22164 , n22165 , n22166 , n22167 , n22168 , n22169 , n22170 , n22171 , n22172 , n22173 , n22174 , n22175 , n22176 , n22177 , n22178 , n22179 , n22180 , n22181 , n22182 , n22183 , n22184 , n22185 , n22186 , n22187 , n22188 , n22189 , n22190 , n22191 , n22192 , n22193 , n22194 , n22195 , n22196 , n22197 , n22198 , n22199 , n22200 , n22201 , n22202 , n22203 , n22204 , n22205 , n22206 , n22207 , n22208 , n22209 , n22210 , n22211 , n22212 , n22213 , n22214 , n22215 , n22216 , n22217 , n22218 , n22219 , n22220 , n22221 , n22222 , n22223 , n22224 , n22225 , n22226 , n22227 , n22228 , n22229 , n22230 , n22231 , n22232 , n22233 , n22234 , n22235 , n22236 , n22237 , n22238 , n22239 , n22240 , n22241 , n22242 , n22243 , n22244 , n22245 , n22246 , n22247 , n22248 , n22249 , n22250 , n22251 , n22252 , n22253 , n22254 , n22255 , n22256 , n22257 , n22258 , n22259 , n22260 , n22261 , n22262 , n22263 , n22264 , n22265 , n22266 , n22267 , n22268 , n22269 , n22270 , n22271 , n22272 , n22273 , n22274 , n22275 , n22276 , n22277 , n22278 , n22279 , n22280 , n22281 , n22282 , n22283 , n22284 , n22285 , n22286 , n22287 , n22288 , n22289 , n22290 , n22291 , n22292 , n22293 , n22294 , n22295 , n22296 , n22297 , n22298 , n22299 , n22300 , n22301 , n22302 , n22303 , n22304 , n22305 , n22306 , n22307 , n22308 , n22309 , n22310 , n22311 , n22312 , n22313 , n22314 , n22315 , n22316 , n22317 , n22318 , n22319 , n22320 , n22321 , n22322 , n22323 , n22324 , n22325 , n22326 , n22327 , n22328 , n22329 , n22330 , n22331 , n22332 , n22333 , n22334 , n22335 , n22336 , n22337 , n22338 , n22339 , n22340 , n22341 , n22342 , n22343 , n22344 , n22345 , n22346 , n22347 , n22348 , n22349 , n22350 , n22351 , n22352 , n22353 , n22354 , n22355 , n22356 , n22357 , n22358 , n22359 , n22360 , n22361 , n22362 , n22363 , n22364 , n22365 , n22366 , n22367 , n22368 , n22369 , n22370 , n22371 , n22372 , n22373 , n22374 , n22375 , n22376 , n22377 , n22378 , n22379 , n22380 , n22381 , n22382 , n22383 , n22384 , n22385 , n22386 , n22387 , n22388 , n22389 , n22390 , n22391 , n22392 , n22393 , n22394 , n22395 , n22396 , n22397 , n22398 , n22399 , n22400 , n22401 , n22402 , n22403 , n22404 , n22405 , n22406 , n22407 , n22408 , n22409 , n22410 , n22411 , n22412 , n22413 , n22414 , n22415 , n22416 , n22417 , n22418 , n22419 , n22420 , n22421 , n22422 , n22423 , n22424 , n22425 , n22426 , n22427 , n22428 , n22429 , n22430 , n22431 , n22432 , n22433 , n22434 , n22435 , n22436 , n22437 , n22438 , n22439 , n22440 , n22441 , n22442 , n22443 , n22444 , n22445 , n22446 , n22447 , n22448 , n22449 , n22450 , n22451 , n22452 , n22453 , n22454 , n22455 , n22456 , n22457 , n22458 , n22459 , n22460 , n22461 , n22462 , n22463 , n22464 , n22465 , n22466 , n22467 , n22468 , n22469 , n22470 , n22471 , n22472 , n22473 , n22474 , n22475 , n22476 , n22477 , n22478 , n22479 , n22480 , n22481 , n22482 , n22483 , n22484 , n22485 , n22486 , n22487 , n22488 , n22489 , n22490 , n22491 , n22492 , n22493 , n22494 , n22495 , n22496 , n22497 , n22498 , n22499 , n22500 , n22501 , n22502 , n22503 , n22504 , n22505 , n22506 , n22507 , n22508 , n22509 , n22510 , n22511 , n22512 , n22513 , n22514 , n22515 , n22516 , n22517 , n22518 , n22519 , n22520 , n22521 , n22522 , n22523 , n22524 , n22525 , n22526 , n22527 , n22528 , n22529 , n22530 , n22531 , n22532 , n22533 , n22534 , n22535 , n22536 , n22537 , n22538 , n22539 , n22540 , n22541 , n22542 , n22543 , n22544 , n22545 , n22546 , n22547 , n22548 , n22549 , n22550 , n22551 , n22552 , n22553 , n22554 , n22555 , n22556 , n22557 , n22558 , n22559 , n22560 , n22561 , n22562 , n22563 , n22564 , n22565 , n22566 , n22567 , n22568 , n22569 , n22570 , n22571 , n22572 , n22573 , n22574 , n22575 , n22576 , n22577 , n22578 , n22579 , n22580 , n22581 , n22582 , n22583 , n22584 , n22585 , n22586 , n22587 , n22588 , n22589 , n22590 , n22591 , n22592 , n22593 , n22594 , n22595 , n22596 , n22597 , n22598 , n22599 , n22600 , n22601 , n22602 , n22603 , n22604 , n22605 , n22606 , n22607 , n22608 , n22609 , n22610 , n22611 , n22612 , n22613 , n22614 , n22615 , n22616 , n22617 , n22618 , n22619 , n22620 , n22621 , n22622 , n22623 , n22624 , n22625 , n22626 , n22627 , n22628 , n22629 , n22630 , n22631 , n22632 , n22633 , n22634 , n22635 , n22636 , n22637 , n22638 , n22639 , n22640 , n22641 , n22642 , n22643 , n22644 , n22645 , n22646 , n22647 , n22648 , n22649 , n22650 , n22651 , n22652 , n22653 , n22654 , n22655 , n22656 , n22657 , n22658 , n22659 , n22660 , n22661 , n22662 , n22663 , n22664 , n22665 , n22666 , n22667 , n22668 , n22669 , n22670 , n22671 , n22672 , n22673 , n22674 , n22675 , n22676 , n22677 , n22678 , n22679 , n22680 , n22681 , n22682 , n22683 , n22684 , n22685 , n22686 , n22687 , n22688 , n22689 , n22690 , n22691 , n22692 , n22693 , n22694 , n22695 , n22696 , n22697 , n22698 , n22699 , n22700 , n22701 , n22702 , n22703 , n22704 , n22705 , n22706 , n22707 , n22708 , n22709 , n22710 , n22711 , n22712 , n22713 , n22714 , n22715 , n22716 , n22717 , n22718 , n22719 , n22720 , n22721 , n22722 , n22723 , n22724 , n22725 , n22726 , n22727 , n22728 , n22729 , n22730 , n22731 , n22732 , n22733 , n22734 , n22735 , n22736 , n22737 , n22738 , n22739 , n22740 , n22741 , n22742 , n22743 , n22744 , n22745 , n22746 , n22747 , n22748 , n22749 , n22750 , n22751 , n22752 , n22753 , n22754 , n22755 , n22756 , n22757 , n22758 , n22759 , n22760 , n22761 , n22762 , n22763 , n22764 , n22765 , n22766 , n22767 , n22768 , n22769 , n22770 , n22771 , n22772 , n22773 , n22774 , n22775 , n22776 , n22777 , n22778 , n22779 , n22780 , n22781 , n22782 , n22783 , n22784 , n22785 , n22786 , n22787 , n22788 , n22789 , n22790 , n22791 , n22792 , n22793 , n22794 , n22795 , n22796 , n22797 , n22798 , n22799 , n22800 , n22801 , n22802 , n22803 , n22804 , n22805 , n22806 , n22807 , n22808 , n22809 , n22810 , n22811 , n22812 , n22813 , n22814 , n22815 , n22816 , n22817 , n22818 , n22819 , n22820 , n22821 , n22822 , n22823 , n22824 , n22825 , n22826 , n22827 , n22828 , n22829 , n22830 , n22831 , n22832 , n22833 , n22834 , n22835 , n22836 , n22837 , n22838 , n22839 , n22840 , n22841 , n22842 , n22843 , n22844 , n22845 , n22846 , n22847 , n22848 , n22849 , n22850 , n22851 , n22852 , n22853 , n22854 , n22855 , n22856 , n22857 , n22858 , n22859 , n22860 , n22861 , n22862 , n22863 , n22864 , n22865 , n22866 , n22867 , n22868 , n22869 , n22870 , n22871 , n22872 , n22873 , n22874 , n22875 , n22876 , n22877 , n22878 , n22879 , n22880 , n22881 , n22882 , n22883 , n22884 , n22885 , n22886 , n22887 , n22888 , n22889 , n22890 , n22891 , n22892 , n22893 , n22894 , n22895 , n22896 , n22897 , n22898 , n22899 , n22900 , n22901 , n22902 , n22903 , n22904 , n22905 , n22906 , n22907 , n22908 , n22909 , n22910 , n22911 , n22912 , n22913 , n22914 , n22915 , n22916 , n22917 , n22918 , n22919 , n22920 , n22921 , n22922 , n22923 , n22924 , n22925 , n22926 , n22927 , n22928 , n22929 , n22930 , n22931 , n22932 , n22933 , n22934 , n22935 , n22936 , n22937 , n22938 , n22939 , n22940 , n22941 , n22942 , n22943 , n22944 , n22945 , n22946 , n22947 , n22948 , n22949 , n22950 , n22951 , n22952 , n22953 , n22954 , n22955 , n22956 , n22957 , n22958 , n22959 , n22960 , n22961 , n22962 , n22963 , n22964 , n22965 , n22966 , n22967 , n22968 , n22969 , n22970 , n22971 , n22972 , n22973 , n22974 , n22975 , n22976 , n22977 , n22978 , n22979 , n22980 , n22981 , n22982 , n22983 , n22984 , n22985 , n22986 , n22987 , n22988 , n22989 , n22990 , n22991 , n22992 , n22993 , n22994 , n22995 , n22996 , n22997 , n22998 , n22999 , n23000 , n23001 , n23002 , n23003 , n23004 , n23005 , n23006 , n23007 , n23008 , n23009 , n23010 , n23011 , n23012 , n23013 , n23014 , n23015 , n23016 , n23017 , n23018 , n23019 , n23020 , n23021 , n23022 , n23023 , n23024 , n23025 , n23026 , n23027 , n23028 , n23029 , n23030 , n23031 , n23032 , n23033 , n23034 , n23035 , n23036 , n23037 , n23038 , n23039 , n23040 , n23041 , n23042 , n23043 , n23044 , n23045 , n23046 , n23047 , n23048 , n23049 , n23050 , n23051 , n23052 , n23053 , n23054 , n23055 , n23056 , n23057 , n23058 , n23059 , n23060 , n23061 , n23062 , n23063 , n23064 , n23065 , n23066 , n23067 , n23068 , n23069 , n23070 , n23071 , n23072 , n23073 , n23074 , n23075 , n23076 , n23077 , n23078 , n23079 , n23080 , n23081 , n23082 , n23083 , n23084 , n23085 , n23086 , n23087 , n23088 , n23089 , n23090 , n23091 , n23092 , n23093 , n23094 , n23095 , n23096 , n23097 , n23098 , n23099 , n23100 , n23101 , n23102 , n23103 , n23104 , n23105 , n23106 , n23107 , n23108 , n23109 , n23110 , n23111 , n23112 , n23113 , n23114 , n23115 , n23116 , n23117 , n23118 , n23119 , n23120 , n23121 , n23122 , n23123 , n23124 , n23125 , n23126 , n23127 , n23128 , n23129 , n23130 , n23131 , n23132 , n23133 , n23134 , n23135 , n23136 , n23137 , n23138 , n23139 , n23140 , n23141 , n23142 , n23143 , n23144 , n23145 , n23146 , n23147 , n23148 , n23149 , n23150 , n23151 , n23152 , n23153 , n23154 , n23155 , n23156 , n23157 , n23158 , n23159 , n23160 , n23161 , n23162 , n23163 , n23164 , n23165 , n23166 , n23167 , n23168 , n23169 , n23170 , n23171 , n23172 , n23173 , n23174 , n23175 , n23176 , n23177 , n23178 , n23179 , n23180 , n23181 , n23182 , n23183 , n23184 , n23185 , n23186 , n23187 , n23188 , n23189 , n23190 , n23191 , n23192 , n23193 , n23194 , n23195 , n23196 , n23197 , n23198 , n23199 , n23200 , n23201 , n23202 , n23203 , n23204 , n23205 , n23206 , n23207 , n23208 , n23209 , n23210 , n23211 , n23212 , n23213 , n23214 , n23215 , n23216 , n23217 , n23218 , n23219 , n23220 , n23221 , n23222 , n23223 , n23224 , n23225 , n23226 , n23227 , n23228 , n23229 , n23230 , n23231 , n23232 , n23233 , n23234 , n23235 , n23236 , n23237 , n23238 , n23239 , n23240 , n23241 , n23242 , n23243 , n23244 , n23245 , n23246 , n23247 , n23248 , n23249 , n23250 , n23251 , n23252 , n23253 , n23254 , n23255 , n23256 , n23257 , n23258 , n23259 , n23260 , n23261 , n23262 , n23263 , n23264 , n23265 , n23266 , n23267 , n23268 , n23269 , n23270 , n23271 , n23272 , n23273 , n23274 , n23275 , n23276 , n23277 , n23278 , n23279 , n23280 , n23281 , n23282 , n23283 , n23284 , n23285 , n23286 , n23287 , n23288 , n23289 , n23290 , n23291 , n23292 , n23293 , n23294 , n23295 , n23296 , n23297 , n23298 , n23299 , n23300 , n23301 , n23302 , n23303 , n23304 , n23305 , n23306 , n23307 , n23308 , n23309 , n23310 , n23311 , n23312 , n23313 , n23314 , n23315 , n23316 , n23317 , n23318 , n23319 , n23320 , n23321 , n23322 , n23323 , n23324 , n23325 , n23326 , n23327 , n23328 , n23329 , n23330 , n23331 , n23332 , n23333 , n23334 , n23335 , n23336 , n23337 , n23338 , n23339 , n23340 , n23341 , n23342 , n23343 , n23344 , n23345 , n23346 , n23347 , n23348 , n23349 , n23350 , n23351 , n23352 , n23353 , n23354 , n23355 , n23356 , n23357 , n23358 , n23359 , n23360 , n23361 , n23362 , n23363 , n23364 , n23365 , n23366 , n23367 , n23368 , n23369 , n23370 , n23371 , n23372 , n23373 , n23374 , n23375 , n23376 , n23377 , n23378 , n23379 , n23380 , n23381 , n23382 , n23383 , n23384 , n23385 , n23386 , n23387 , n23388 , n23389 , n23390 , n23391 , n23392 , n23393 , n23394 , n23395 , n23396 , n23397 , n23398 , n23399 , n23400 , n23401 , n23402 , n23403 , n23404 , n23405 , n23406 , n23407 , n23408 , n23409 , n23410 , n23411 , n23412 , n23413 , n23414 , n23415 , n23416 , n23417 , n23418 , n23419 , n23420 , n23421 , n23422 , n23423 , n23424 , n23425 , n23426 , n23427 , n23428 , n23429 , n23430 , n23431 , n23432 , n23433 , n23434 , n23435 , n23436 , n23437 , n23438 , n23439 , n23440 , n23441 , n23442 , n23443 , n23444 , n23445 , n23446 , n23447 , n23448 , n23449 , n23450 , n23451 , n23452 , n23453 , n23454 , n23455 , n23456 , n23457 , n23458 , n23459 , n23460 , n23461 , n23462 , n23463 , n23464 , n23465 , n23466 , n23467 , n23468 , n23469 , n23470 , n23471 , n23472 , n23473 , n23474 , n23475 , n23476 , n23477 , n23478 , n23479 , n23480 , n23481 , n23482 , n23483 , n23484 , n23485 , n23486 , n23487 , n23488 , n23489 , n23490 , n23491 , n23492 , n23493 , n23494 , n23495 , n23496 , n23497 , n23498 , n23499 , n23500 , n23501 , n23502 , n23503 , n23504 , n23505 , n23506 , n23507 , n23508 , n23509 , n23510 , n23511 , n23512 , n23513 , n23514 , n23515 , n23516 , n23517 , n23518 , n23519 , n23520 , n23521 , n23522 , n23523 , n23524 , n23525 , n23526 , n23527 , n23528 , n23529 , n23530 , n23531 , n23532 , n23533 , n23534 , n23535 , n23536 , n23537 , n23538 , n23539 , n23540 , n23541 , n23542 , n23543 , n23544 , n23545 , n23546 , n23547 , n23548 , n23549 , n23550 , n23551 , n23552 , n23553 , n23554 , n23555 , n23556 , n23557 , n23558 , n23559 , n23560 , n23561 , n23562 , n23563 , n23564 , n23565 , n23566 , n23567 , n23568 , n23569 , n23570 , n23571 , n23572 , n23573 , n23574 , n23575 , n23576 , n23577 , n23578 , n23579 , n23580 , n23581 , n23582 , n23583 , n23584 , n23585 , n23586 , n23587 , n23588 , n23589 , n23590 , n23591 , n23592 , n23593 , n23594 , n23595 , n23596 , n23597 , n23598 , n23599 , n23600 , n23601 , n23602 , n23603 , n23604 , n23605 , n23606 , n23607 , n23608 , n23609 , n23610 , n23611 , n23612 , n23613 , n23614 , n23615 , n23616 , n23617 , n23618 , n23619 , n23620 , n23621 , n23622 , n23623 , n23624 , n23625 , n23626 , n23627 , n23628 , n23629 , n23630 , n23631 , n23632 , n23633 , n23634 , n23635 , n23636 , n23637 , n23638 , n23639 , n23640 , n23641 , n23642 , n23643 , n23644 , n23645 , n23646 , n23647 , n23648 , n23649 , n23650 , n23651 , n23652 , n23653 , n23654 , n23655 , n23656 , n23657 , n23658 , n23659 , n23660 , n23661 , n23662 , n23663 , n23664 , n23665 , n23666 , n23667 , n23668 , n23669 , n23670 , n23671 , n23672 , n23673 , n23674 , n23675 , n23676 , n23677 , n23678 , n23679 , n23680 , n23681 , n23682 , n23683 , n23684 , n23685 , n23686 , n23687 , n23688 , n23689 , n23690 , n23691 , n23692 , n23693 , n23694 , n23695 , n23696 , n23697 , n23698 , n23699 , n23700 , n23701 , n23702 , n23703 , n23704 , n23705 , n23706 , n23707 , n23708 , n23709 , n23710 , n23711 , n23712 , n23713 , n23714 , n23715 , n23716 , n23717 , n23718 , n23719 , n23720 , n23721 , n23722 , n23723 , n23724 , n23725 , n23726 , n23727 , n23728 , n23729 , n23730 , n23731 , n23732 , n23733 , n23734 , n23735 , n23736 , n23737 , n23738 , n23739 , n23740 , n23741 , n23742 , n23743 , n23744 , n23745 , n23746 , n23747 , n23748 , n23749 , n23750 , n23751 , n23752 , n23753 , n23754 , n23755 , n23756 , n23757 , n23758 , n23759 , n23760 , n23761 , n23762 , n23763 , n23764 , n23765 , n23766 , n23767 , n23768 , n23769 , n23770 , n23771 , n23772 , n23773 , n23774 , n23775 , n23776 , n23777 , n23778 , n23779 , n23780 , n23781 , n23782 , n23783 , n23784 , n23785 , n23786 , n23787 , n23788 , n23789 , n23790 , n23791 , n23792 , n23793 , n23794 , n23795 , n23796 , n23797 , n23798 , n23799 , n23800 , n23801 , n23802 , n23803 , n23804 , n23805 , n23806 , n23807 , n23808 , n23809 , n23810 , n23811 , n23812 , n23813 , n23814 , n23815 , n23816 , n23817 , n23818 , n23819 , n23820 , n23821 , n23822 , n23823 , n23824 , n23825 , n23826 , n23827 , n23828 , n23829 , n23830 , n23831 , n23832 , n23833 , n23834 , n23835 , n23836 , n23837 , n23838 , n23839 , n23840 , n23841 , n23842 , n23843 , n23844 , n23845 , n23846 , n23847 , n23848 , n23849 , n23850 , n23851 , n23852 , n23853 , n23854 , n23855 , n23856 , n23857 , n23858 , n23859 , n23860 , n23861 , n23862 , n23863 , n23864 , n23865 , n23866 , n23867 , n23868 , n23869 , n23870 , n23871 , n23872 , n23873 , n23874 , n23875 , n23876 , n23877 , n23878 , n23879 , n23880 , n23881 , n23882 , n23883 , n23884 , n23885 , n23886 , n23887 , n23888 , n23889 , n23890 , n23891 , n23892 , n23893 , n23894 , n23895 , n23896 , n23897 , n23898 , n23899 , n23900 , n23901 , n23902 , n23903 , n23904 , n23905 , n23906 , n23907 , n23908 , n23909 , n23910 , n23911 , n23912 , n23913 , n23914 , n23915 , n23916 , n23917 , n23918 , n23919 , n23920 , n23921 , n23922 , n23923 , n23924 , n23925 , n23926 , n23927 , n23928 , n23929 , n23930 , n23931 , n23932 , n23933 , n23934 , n23935 , n23936 , n23937 , n23938 , n23939 , n23940 , n23941 , n23942 , n23943 , n23944 , n23945 , n23946 , n23947 , n23948 , n23949 , n23950 , n23951 , n23952 , n23953 , n23954 , n23955 , n23956 , n23957 , n23958 , n23959 , n23960 , n23961 , n23962 , n23963 , n23964 , n23965 , n23966 , n23967 , n23968 , n23969 , n23970 , n23971 , n23972 , n23973 , n23974 , n23975 , n23976 , n23977 , n23978 , n23979 , n23980 , n23981 , n23982 , n23983 , n23984 , n23985 , n23986 , n23987 , n23988 , n23989 , n23990 , n23991 , n23992 , n23993 , n23994 , n23995 , n23996 , n23997 , n23998 , n23999 , n24000 , n24001 , n24002 , n24003 , n24004 , n24005 , n24006 , n24007 , n24008 , n24009 , n24010 , n24011 , n24012 , n24013 , n24014 , n24015 , n24016 , n24017 , n24018 , n24019 , n24020 , n24021 , n24022 , n24023 , n24024 , n24025 , n24026 , n24027 , n24028 , n24029 , n24030 , n24031 , n24032 , n24033 , n24034 , n24035 , n24036 , n24037 , n24038 , n24039 , n24040 , n24041 , n24042 , n24043 , n24044 , n24045 , n24046 , n24047 , n24048 , n24049 , n24050 , n24051 , n24052 , n24053 , n24054 , n24055 , n24056 , n24057 , n24058 , n24059 , n24060 , n24061 , n24062 , n24063 , n24064 , n24065 , n24066 , n24067 , n24068 , n24069 , n24070 , n24071 , n24072 , n24073 , n24074 , n24075 , n24076 , n24077 , n24078 , n24079 , n24080 , n24081 , n24082 , n24083 , n24084 , n24085 , n24086 , n24087 , n24088 , n24089 , n24090 , n24091 , n24092 , n24093 , n24094 , n24095 , n24096 , n24097 , n24098 , n24099 , n24100 , n24101 , n24102 , n24103 , n24104 , n24105 , n24106 , n24107 , n24108 , n24109 , n24110 , n24111 , n24112 , n24113 , n24114 , n24115 , n24116 , n24117 , n24118 , n24119 , n24120 , n24121 , n24122 , n24123 , n24124 , n24125 , n24126 , n24127 , n24128 , n24129 , n24130 , n24131 , n24132 , n24133 , n24134 , n24135 , n24136 , n24137 , n24138 , n24139 , n24140 , n24141 , n24142 , n24143 , n24144 , n24145 , n24146 , n24147 , n24148 , n24149 , n24150 , n24151 , n24152 , n24153 , n24154 , n24155 , n24156 , n24157 , n24158 , n24159 , n24160 , n24161 , n24162 , n24163 , n24164 , n24165 , n24166 , n24167 , n24168 , n24169 , n24170 , n24171 , n24172 , n24173 , n24174 , n24175 , n24176 , n24177 , n24178 , n24179 , n24180 , n24181 , n24182 , n24183 , n24184 , n24185 , n24186 , n24187 , n24188 , n24189 , n24190 , n24191 , n24192 , n24193 , n24194 , n24195 , n24196 , n24197 , n24198 , n24199 , n24200 , n24201 , n24202 , n24203 , n24204 , n24205 , n24206 , n24207 , n24208 , n24209 , n24210 , n24211 , n24212 , n24213 , n24214 , n24215 , n24216 , n24217 , n24218 , n24219 , n24220 , n24221 , n24222 , n24223 , n24224 , n24225 , n24226 , n24227 , n24228 , n24229 , n24230 , n24231 , n24232 , n24233 , n24234 , n24235 , n24236 , n24237 , n24238 , n24239 , n24240 , n24241 , n24242 , n24243 , n24244 , n24245 , n24246 , n24247 , n24248 , n24249 , n24250 , n24251 , n24252 , n24253 , n24254 , n24255 , n24256 , n24257 , n24258 , n24259 , n24260 , n24261 , n24262 , n24263 , n24264 , n24265 , n24266 , n24267 , n24268 , n24269 , n24270 , n24271 , n24272 , n24273 , n24274 , n24275 , n24276 , n24277 , n24278 , n24279 , n24280 , n24281 , n24282 , n24283 , n24284 , n24285 , n24286 , n24287 , n24288 , n24289 , n24290 , n24291 , n24292 , n24293 , n24294 , n24295 , n24296 , n24297 , n24298 , n24299 , n24300 , n24301 , n24302 , n24303 , n24304 , n24305 , n24306 , n24307 , n24308 , n24309 , n24310 , n24311 , n24312 , n24313 , n24314 , n24315 , n24316 , n24317 , n24318 , n24319 , n24320 , n24321 , n24322 , n24323 , n24324 , n24325 , n24326 , n24327 , n24328 , n24329 , n24330 , n24331 , n24332 , n24333 , n24334 , n24335 , n24336 , n24337 , n24338 , n24339 , n24340 , n24341 , n24342 , n24343 , n24344 , n24345 , n24346 , n24347 , n24348 , n24349 , n24350 , n24351 , n24352 , n24353 , n24354 , n24355 , n24356 , n24357 , n24358 , n24359 , n24360 , n24361 , n24362 , n24363 , n24364 , n24365 , n24366 , n24367 , n24368 , n24369 , n24370 , n24371 , n24372 , n24373 , n24374 , n24375 , n24376 , n24377 , n24378 , n24379 , n24380 , n24381 , n24382 , n24383 , n24384 , n24385 , n24386 , n24387 , n24388 , n24389 , n24390 , n24391 , n24392 , n24393 , n24394 , n24395 , n24396 , n24397 , n24398 , n24399 , n24400 , n24401 , n24402 , n24403 , n24404 , n24405 , n24406 , n24407 , n24408 , n24409 , n24410 , n24411 , n24412 , n24413 , n24414 , n24415 , n24416 , n24417 , n24418 , n24419 , n24420 , n24421 , n24422 , n24423 , n24424 , n24425 , n24426 , n24427 , n24428 , n24429 , n24430 , n24431 , n24432 , n24433 , n24434 , n24435 , n24436 , n24437 , n24438 , n24439 , n24440 , n24441 , n24442 , n24443 , n24444 , n24445 , n24446 , n24447 , n24448 , n24449 , n24450 , n24451 , n24452 , n24453 , n24454 , n24455 , n24456 , n24457 , n24458 , n24459 , n24460 , n24461 , n24462 , n24463 , n24464 , n24465 , n24466 , n24467 , n24468 , n24469 , n24470 , n24471 , n24472 , n24473 , n24474 , n24475 , n24476 , n24477 , n24478 , n24479 , n24480 , n24481 , n24482 , n24483 , n24484 , n24485 , n24486 , n24487 , n24488 , n24489 , n24490 , n24491 , n24492 , n24493 , n24494 , n24495 , n24496 , n24497 , n24498 , n24499 , n24500 , n24501 , n24502 , n24503 , n24504 , n24505 , n24506 , n24507 , n24508 , n24509 , n24510 , n24511 , n24512 , n24513 , n24514 , n24515 , n24516 , n24517 , n24518 , n24519 , n24520 , n24521 , n24522 , n24523 , n24524 , n24525 , n24526 , n24527 , n24528 , n24529 , n24530 , n24531 , n24532 , n24533 , n24534 , n24535 , n24536 , n24537 , n24538 , n24539 , n24540 , n24541 , n24542 , n24543 , n24544 , n24545 , n24546 , n24547 , n24548 , n24549 , n24550 , n24551 , n24552 , n24553 , n24554 , n24555 , n24556 , n24557 , n24558 , n24559 , n24560 , n24561 , n24562 , n24563 , n24564 , n24565 , n24566 , n24567 , n24568 , n24569 , n24570 , n24571 , n24572 , n24573 , n24574 , n24575 , n24576 , n24577 , n24578 , n24579 , n24580 , n24581 , n24582 , n24583 , n24584 , n24585 , n24586 , n24587 , n24588 , n24589 , n24590 , n24591 , n24592 , n24593 , n24594 , n24595 , n24596 , n24597 , n24598 , n24599 , n24600 , n24601 , n24602 , n24603 , n24604 , n24605 , n24606 , n24607 , n24608 , n24609 , n24610 , n24611 , n24612 , n24613 , n24614 , n24615 , n24616 , n24617 , n24618 , n24619 , n24620 , n24621 , n24622 , n24623 , n24624 , n24625 , n24626 , n24627 , n24628 , n24629 , n24630 , n24631 , n24632 , n24633 , n24634 , n24635 , n24636 , n24637 , n24638 , n24639 , n24640 , n24641 , n24642 , n24643 , n24644 , n24645 , n24646 , n24647 , n24648 , n24649 , n24650 , n24651 , n24652 , n24653 , n24654 , n24655 , n24656 , n24657 , n24658 , n24659 , n24660 , n24661 , n24662 , n24663 , n24664 , n24665 , n24666 , n24667 , n24668 , n24669 , n24670 , n24671 , n24672 , n24673 , n24674 , n24675 , n24676 , n24677 , n24678 , n24679 , n24680 , n24681 , n24682 , n24683 , n24684 , n24685 , n24686 , n24687 , n24688 , n24689 , n24690 , n24691 , n24692 , n24693 , n24694 , n24695 , n24696 , n24697 , n24698 , n24699 , n24700 , n24701 , n24702 , n24703 , n24704 , n24705 , n24706 , n24707 , n24708 , n24709 , n24710 , n24711 , n24712 , n24713 , n24714 , n24715 , n24716 , n24717 , n24718 , n24719 , n24720 , n24721 , n24722 , n24723 , n24724 , n24725 , n24726 , n24727 , n24728 , n24729 , n24730 , n24731 , n24732 , n24733 , n24734 , n24735 , n24736 , n24737 , n24738 , n24739 , n24740 , n24741 , n24742 , n24743 , n24744 , n24745 , n24746 , n24747 , n24748 , n24749 , n24750 , n24751 , n24752 , n24753 , n24754 , n24755 , n24756 , n24757 , n24758 , n24759 , n24760 , n24761 , n24762 , n24763 , n24764 , n24765 , n24766 , n24767 , n24768 , n24769 , n24770 , n24771 , n24772 , n24773 , n24774 , n24775 , n24776 , n24777 , n24778 , n24779 , n24780 , n24781 , n24782 , n24783 , n24784 , n24785 , n24786 , n24787 , n24788 , n24789 , n24790 , n24791 , n24792 , n24793 , n24794 , n24795 , n24796 , n24797 , n24798 , n24799 , n24800 , n24801 , n24802 , n24803 , n24804 , n24805 , n24806 , n24807 , n24808 , n24809 , n24810 , n24811 , n24812 , n24813 , n24814 , n24815 , n24816 , n24817 , n24818 , n24819 , n24820 , n24821 , n24822 , n24823 , n24824 , n24825 , n24826 , n24827 , n24828 , n24829 , n24830 , n24831 , n24832 , n24833 , n24834 , n24835 , n24836 , n24837 , n24838 , n24839 , n24840 , n24841 , n24842 , n24843 , n24844 , n24845 , n24846 , n24847 , n24848 , n24849 , n24850 , n24851 , n24852 , n24853 , n24854 , n24855 , n24856 , n24857 , n24858 , n24859 , n24860 , n24861 , n24862 , n24863 , n24864 , n24865 , n24866 , n24867 , n24868 , n24869 , n24870 , n24871 , n24872 , n24873 , n24874 , n24875 , n24876 , n24877 , n24878 , n24879 , n24880 , n24881 , n24882 , n24883 , n24884 , n24885 , n24886 , n24887 , n24888 , n24889 , n24890 , n24891 , n24892 , n24893 , n24894 , n24895 , n24896 , n24897 , n24898 , n24899 , n24900 , n24901 , n24902 , n24903 , n24904 , n24905 , n24906 , n24907 , n24908 , n24909 , n24910 , n24911 , n24912 , n24913 , n24914 , n24915 , n24916 , n24917 , n24918 , n24919 , n24920 , n24921 , n24922 , n24923 , n24924 , n24925 , n24926 , n24927 , n24928 , n24929 , n24930 , n24931 , n24932 , n24933 , n24934 , n24935 , n24936 , n24937 , n24938 , n24939 , n24940 , n24941 , n24942 , n24943 , n24944 , n24945 , n24946 , n24947 , n24948 , n24949 , n24950 , n24951 , n24952 , n24953 , n24954 , n24955 , n24956 , n24957 , n24958 , n24959 , n24960 , n24961 , n24962 , n24963 , n24964 , n24965 , n24966 , n24967 , n24968 , n24969 , n24970 , n24971 , n24972 , n24973 , n24974 , n24975 , n24976 , n24977 , n24978 , n24979 , n24980 , n24981 , n24982 , n24983 , n24984 , n24985 , n24986 , n24987 , n24988 , n24989 , n24990 , n24991 , n24992 , n24993 , n24994 , n24995 , n24996 , n24997 , n24998 , n24999 , n25000 , n25001 , n25002 , n25003 , n25004 , n25005 , n25006 , n25007 , n25008 , n25009 , n25010 , n25011 , n25012 , n25013 , n25014 , n25015 , n25016 , n25017 , n25018 , n25019 , n25020 , n25021 , n25022 , n25023 , n25024 , n25025 , n25026 , n25027 , n25028 , n25029 , n25030 , n25031 , n25032 , n25033 , n25034 , n25035 , n25036 , n25037 , n25038 , n25039 , n25040 , n25041 , n25042 , n25043 , n25044 , n25045 , n25046 , n25047 , n25048 , n25049 , n25050 , n25051 , n25052 , n25053 , n25054 , n25055 , n25056 , n25057 , n25058 , n25059 , n25060 , n25061 , n25062 , n25063 , n25064 , n25065 , n25066 , n25067 , n25068 , n25069 , n25070 , n25071 , n25072 , n25073 , n25074 , n25075 , n25076 , n25077 , n25078 , n25079 , n25080 , n25081 , n25082 , n25083 , n25084 , n25085 , n25086 , n25087 , n25088 , n25089 , n25090 , n25091 , n25092 , n25093 , n25094 , n25095 , n25096 , n25097 , n25098 , n25099 , n25100 , n25101 , n25102 , n25103 , n25104 , n25105 , n25106 , n25107 , n25108 , n25109 , n25110 , n25111 , n25112 , n25113 , n25114 , n25115 , n25116 , n25117 , n25118 , n25119 , n25120 , n25121 , n25122 , n25123 , n25124 , n25125 , n25126 , n25127 , n25128 , n25129 , n25130 , n25131 , n25132 , n25133 , n25134 , n25135 , n25136 , n25137 , n25138 , n25139 , n25140 , n25141 , n25142 , n25143 , n25144 , n25145 , n25146 , n25147 , n25148 , n25149 , n25150 , n25151 , n25152 , n25153 , n25154 , n25155 , n25156 , n25157 , n25158 , n25159 , n25160 , n25161 , n25162 , n25163 , n25164 , n25165 , n25166 , n25167 , n25168 , n25169 , n25170 , n25171 , n25172 , n25173 , n25174 , n25175 , n25176 , n25177 , n25178 , n25179 , n25180 , n25181 , n25182 , n25183 , n25184 , n25185 , n25186 , n25187 , n25188 , n25189 , n25190 , n25191 , n25192 , n25193 , n25194 , n25195 , n25196 , n25197 , n25198 , n25199 , n25200 , n25201 , n25202 , n25203 , n25204 , n25205 , n25206 , n25207 , n25208 , n25209 , n25210 , n25211 , n25212 , n25213 , n25214 , n25215 , n25216 , n25217 , n25218 , n25219 , n25220 , n25221 , n25222 , n25223 , n25224 , n25225 , n25226 , n25227 , n25228 , n25229 , n25230 , n25231 , n25232 , n25233 , n25234 , n25235 , n25236 , n25237 , n25238 , n25239 , n25240 , n25241 , n25242 , n25243 , n25244 , n25245 , n25246 , n25247 , n25248 , n25249 , n25250 , n25251 , n25252 , n25253 , n25254 , n25255 , n25256 , n25257 , n25258 , n25259 , n25260 , n25261 , n25262 , n25263 , n25264 , n25265 , n25266 , n25267 , n25268 , n25269 , n25270 , n25271 , n25272 , n25273 , n25274 , n25275 , n25276 , n25277 , n25278 , n25279 , n25280 , n25281 , n25282 , n25283 , n25284 , n25285 , n25286 , n25287 , n25288 , n25289 , n25290 , n25291 , n25292 , n25293 , n25294 , n25295 , n25296 , n25297 , n25298 , n25299 , n25300 , n25301 , n25302 , n25303 , n25304 , n25305 , n25306 , n25307 , n25308 , n25309 , n25310 , n25311 , n25312 , n25313 , n25314 , n25315 , n25316 , n25317 , n25318 , n25319 , n25320 , n25321 , n25322 , n25323 , n25324 , n25325 , n25326 , n25327 , n25328 , n25329 , n25330 , n25331 , n25332 , n25333 , n25334 , n25335 , n25336 , n25337 , n25338 , n25339 , n25340 , n25341 , n25342 , n25343 , n25344 , n25345 , n25346 , n25347 , n25348 , n25349 , n25350 , n25351 , n25352 , n25353 , n25354 , n25355 , n25356 , n25357 , n25358 , n25359 , n25360 , n25361 , n25362 , n25363 , n25364 , n25365 , n25366 , n25367 , n25368 , n25369 , n25370 , n25371 , n25372 , n25373 , n25374 , n25375 , n25376 , n25377 , n25378 , n25379 , n25380 , n25381 , n25382 , n25383 , n25384 , n25385 , n25386 , n25387 , n25388 , n25389 , n25390 , n25391 , n25392 , n25393 , n25394 , n25395 , n25396 , n25397 , n25398 , n25399 , n25400 , n25401 , n25402 , n25403 , n25404 , n25405 , n25406 , n25407 , n25408 , n25409 , n25410 , n25411 , n25412 , n25413 , n25414 , n25415 , n25416 , n25417 , n25418 , n25419 , n25420 , n25421 , n25422 , n25423 , n25424 , n25425 , n25426 , n25427 , n25428 , n25429 , n25430 , n25431 , n25432 , n25433 , n25434 , n25435 , n25436 , n25437 , n25438 , n25439 , n25440 , n25441 , n25442 , n25443 , n25444 , n25445 , n25446 , n25447 , n25448 , n25449 , n25450 , n25451 , n25452 , n25453 , n25454 , n25455 , n25456 , n25457 , n25458 , n25459 , n25460 , n25461 , n25462 , n25463 , n25464 , n25465 , n25466 , n25467 , n25468 , n25469 , n25470 , n25471 , n25472 , n25473 , n25474 , n25475 , n25476 , n25477 , n25478 , n25479 , n25480 , n25481 , n25482 , n25483 , n25484 , n25485 , n25486 , n25487 , n25488 , n25489 , n25490 , n25491 , n25492 , n25493 , n25494 , n25495 , n25496 , n25497 , n25498 , n25499 , n25500 , n25501 , n25502 , n25503 , n25504 , n25505 , n25506 , n25507 , n25508 , n25509 , n25510 , n25511 , n25512 , n25513 , n25514 , n25515 , n25516 , n25517 , n25518 , n25519 , n25520 , n25521 , n25522 , n25523 , n25524 , n25525 , n25526 , n25527 , n25528 , n25529 , n25530 , n25531 , n25532 , n25533 , n25534 , n25535 , n25536 , n25537 , n25538 , n25539 , n25540 , n25541 , n25542 , n25543 , n25544 , n25545 , n25546 , n25547 , n25548 , n25549 , n25550 , n25551 , n25552 , n25553 , n25554 , n25555 , n25556 , n25557 , n25558 , n25559 , n25560 , n25561 , n25562 , n25563 , n25564 , n25565 , n25566 , n25567 , n25568 , n25569 , n25570 , n25571 , n25572 , n25573 , n25574 , n25575 , n25576 , n25577 , n25578 , n25579 , n25580 , n25581 , n25582 , n25583 , n25584 , n25585 , n25586 , n25587 , n25588 , n25589 , n25590 , n25591 , n25592 , n25593 , n25594 , n25595 , n25596 , n25597 , n25598 , n25599 , n25600 , n25601 , n25602 , n25603 , n25604 , n25605 , n25606 , n25607 , n25608 , n25609 , n25610 , n25611 , n25612 , n25613 , n25614 , n25615 , n25616 , n25617 , n25618 , n25619 , n25620 , n25621 , n25622 , n25623 , n25624 , n25625 , n25626 , n25627 , n25628 , n25629 , n25630 , n25631 , n25632 , n25633 , n25634 , n25635 , n25636 , n25637 , n25638 , n25639 , n25640 , n25641 , n25642 , n25643 , n25644 , n25645 , n25646 , n25647 , n25648 , n25649 , n25650 , n25651 , n25652 , n25653 , n25654 , n25655 , n25656 , n25657 , n25658 , n25659 , n25660 , n25661 , n25662 , n25663 , n25664 , n25665 , n25666 , n25667 , n25668 , n25669 , n25670 , n25671 , n25672 , n25673 , n25674 , n25675 , n25676 , n25677 , n25678 , n25679 , n25680 , n25681 , n25682 , n25683 , n25684 , n25685 , n25686 , n25687 , n25688 , n25689 , n25690 , n25691 , n25692 , n25693 , n25694 , n25695 , n25696 , n25697 , n25698 , n25699 , n25700 , n25701 , n25702 , n25703 , n25704 , n25705 , n25706 , n25707 , n25708 , n25709 , n25710 , n25711 , n25712 , n25713 , n25714 , n25715 , n25716 , n25717 , n25718 , n25719 , n25720 , n25721 , n25722 , n25723 , n25724 , n25725 , n25726 , n25727 , n25728 , n25729 , n25730 , n25731 , n25732 , n25733 , n25734 , n25735 , n25736 , n25737 , n25738 , n25739 , n25740 , n25741 , n25742 , n25743 , n25744 , n25745 , n25746 , n25747 , n25748 , n25749 , n25750 , n25751 , n25752 , n25753 , n25754 , n25755 , n25756 , n25757 , n25758 , n25759 , n25760 , n25761 , n25762 , n25763 , n25764 , n25765 , n25766 , n25767 , n25768 , n25769 , n25770 , n25771 , n25772 , n25773 , n25774 , n25775 , n25776 , n25777 , n25778 , n25779 , n25780 , n25781 , n25782 , n25783 , n25784 , n25785 , n25786 , n25787 , n25788 , n25789 , n25790 , n25791 , n25792 , n25793 , n25794 , n25795 , n25796 , n25797 , n25798 , n25799 , n25800 , n25801 , n25802 , n25803 , n25804 , n25805 , n25806 , n25807 , n25808 , n25809 , n25810 , n25811 , n25812 , n25813 , n25814 , n25815 , n25816 , n25817 , n25818 , n25819 , n25820 , n25821 , n25822 , n25823 , n25824 , n25825 , n25826 , n25827 , n25828 , n25829 , n25830 , n25831 , n25832 , n25833 , n25834 , n25835 , n25836 , n25837 , n25838 , n25839 , n25840 , n25841 , n25842 , n25843 , n25844 , n25845 , n25846 , n25847 , n25848 , n25849 , n25850 , n25851 , n25852 , n25853 , n25854 , n25855 , n25856 , n25857 , n25858 , n25859 , n25860 , n25861 , n25862 , n25863 , n25864 , n25865 , n25866 , n25867 , n25868 , n25869 , n25870 , n25871 , n25872 , n25873 , n25874 , n25875 , n25876 , n25877 , n25878 , n25879 , n25880 , n25881 , n25882 , n25883 , n25884 , n25885 , n25886 , n25887 , n25888 , n25889 , n25890 , n25891 , n25892 , n25893 , n25894 , n25895 , n25896 , n25897 , n25898 , n25899 , n25900 , n25901 , n25902 , n25903 , n25904 , n25905 , n25906 , n25907 , n25908 , n25909 , n25910 , n25911 , n25912 , n25913 , n25914 , n25915 , n25916 , n25917 , n25918 , n25919 , n25920 , n25921 , n25922 , n25923 , n25924 , n25925 , n25926 , n25927 , n25928 , n25929 , n25930 , n25931 , n25932 , n25933 , n25934 , n25935 , n25936 , n25937 , n25938 , n25939 , n25940 , n25941 , n25942 , n25943 , n25944 , n25945 , n25946 , n25947 , n25948 , n25949 , n25950 , n25951 , n25952 , n25953 , n25954 , n25955 , n25956 , n25957 , n25958 , n25959 , n25960 , n25961 , n25962 , n25963 , n25964 , n25965 , n25966 , n25967 , n25968 , n25969 , n25970 , n25971 , n25972 , n25973 , n25974 , n25975 , n25976 , n25977 , n25978 , n25979 , n25980 , n25981 , n25982 , n25983 , n25984 , n25985 , n25986 , n25987 , n25988 , n25989 , n25990 , n25991 , n25992 , n25993 , n25994 , n25995 , n25996 , n25997 , n25998 , n25999 , n26000 , n26001 , n26002 , n26003 , n26004 , n26005 , n26006 , n26007 , n26008 , n26009 , n26010 , n26011 , n26012 , n26013 , n26014 , n26015 , n26016 , n26017 , n26018 , n26019 , n26020 , n26021 , n26022 , n26023 , n26024 , n26025 , n26026 , n26027 , n26028 , n26029 , n26030 , n26031 , n26032 , n26033 , n26034 , n26035 , n26036 , n26037 , n26038 , n26039 , n26040 , n26041 , n26042 , n26043 , n26044 , n26045 , n26046 , n26047 , n26048 , n26049 , n26050 , n26051 , n26052 , n26053 , n26054 , n26055 , n26056 , n26057 , n26058 , n26059 , n26060 , n26061 , n26062 , n26063 , n26064 , n26065 , n26066 , n26067 , n26068 , n26069 , n26070 , n26071 , n26072 , n26073 , n26074 , n26075 , n26076 , n26077 , n26078 , n26079 , n26080 , n26081 , n26082 , n26083 , n26084 , n26085 , n26086 , n26087 , n26088 , n26089 , n26090 , n26091 , n26092 , n26093 , n26094 , n26095 , n26096 , n26097 , n26098 , n26099 , n26100 , n26101 , n26102 , n26103 , n26104 , n26105 , n26106 , n26107 , n26108 , n26109 , n26110 , n26111 , n26112 , n26113 , n26114 , n26115 , n26116 , n26117 , n26118 , n26119 , n26120 , n26121 , n26122 , n26123 , n26124 , n26125 , n26126 , n26127 , n26128 , n26129 , n26130 , n26131 , n26132 , n26133 , n26134 , n26135 , n26136 , n26137 , n26138 , n26139 , n26140 , n26141 , n26142 , n26143 , n26144 , n26145 , n26146 , n26147 , n26148 , n26149 , n26150 , n26151 , n26152 , n26153 , n26154 , n26155 , n26156 , n26157 , n26158 , n26159 , n26160 , n26161 , n26162 , n26163 , n26164 , n26165 , n26166 , n26167 , n26168 , n26169 , n26170 , n26171 , n26172 , n26173 , n26174 , n26175 , n26176 , n26177 , n26178 , n26179 , n26180 , n26181 , n26182 , n26183 , n26184 , n26185 , n26186 , n26187 , n26188 , n26189 , n26190 , n26191 , n26192 , n26193 , n26194 , n26195 , n26196 , n26197 , n26198 , n26199 , n26200 , n26201 , n26202 , n26203 , n26204 , n26205 , n26206 , n26207 , n26208 , n26209 , n26210 , n26211 , n26212 , n26213 , n26214 , n26215 , n26216 , n26217 , n26218 , n26219 , n26220 , n26221 , n26222 , n26223 , n26224 , n26225 , n26226 , n26227 , n26228 , n26229 , n26230 , n26231 , n26232 , n26233 , n26234 , n26235 , n26236 , n26237 , n26238 , n26239 , n26240 , n26241 , n26242 , n26243 , n26244 , n26245 , n26246 , n26247 , n26248 , n26249 , n26250 , n26251 , n26252 , n26253 , n26254 , n26255 , n26256 , n26257 , n26258 , n26259 , n26260 , n26261 , n26262 , n26263 , n26264 , n26265 , n26266 , n26267 , n26268 , n26269 , n26270 , n26271 , n26272 , n26273 , n26274 , n26275 , n26276 , n26277 , n26278 , n26279 , n26280 , n26281 , n26282 , n26283 , n26284 , n26285 , n26286 , n26287 , n26288 , n26289 , n26290 , n26291 , n26292 , n26293 , n26294 , n26295 , n26296 , n26297 , n26298 , n26299 , n26300 , n26301 , n26302 , n26303 , n26304 , n26305 , n26306 , n26307 , n26308 , n26309 , n26310 , n26311 , n26312 , n26313 , n26314 , n26315 , n26316 , n26317 , n26318 , n26319 , n26320 , n26321 , n26322 , n26323 , n26324 , n26325 , n26326 , n26327 , n26328 , n26329 , n26330 , n26331 , n26332 , n26333 , n26334 , n26335 , n26336 , n26337 , n26338 , n26339 , n26340 , n26341 , n26342 , n26343 , n26344 , n26345 , n26346 , n26347 , n26348 , n26349 , n26350 , n26351 , n26352 , n26353 , n26354 , n26355 , n26356 , n26357 , n26358 , n26359 , n26360 , n26361 , n26362 , n26363 , n26364 , n26365 , n26366 , n26367 , n26368 , n26369 , n26370 , n26371 , n26372 , n26373 , n26374 , n26375 , n26376 , n26377 , n26378 , n26379 , n26380 , n26381 , n26382 , n26383 , n26384 , n26385 , n26386 , n26387 , n26388 , n26389 , n26390 , n26391 , n26392 , n26393 , n26394 , n26395 , n26396 , n26397 , n26398 , n26399 , n26400 , n26401 , n26402 , n26403 , n26404 , n26405 , n26406 , n26407 , n26408 , n26409 , n26410 , n26411 , n26412 , n26413 , n26414 , n26415 , n26416 , n26417 , n26418 , n26419 , n26420 , n26421 , n26422 , n26423 , n26424 , n26425 , n26426 , n26427 , n26428 , n26429 , n26430 , n26431 , n26432 , n26433 , n26434 , n26435 , n26436 , n26437 , n26438 , n26439 , n26440 , n26441 , n26442 , n26443 , n26444 , n26445 , n26446 , n26447 , n26448 , n26449 , n26450 , n26451 , n26452 , n26453 , n26454 , n26455 , n26456 , n26457 , n26458 , n26459 , n26460 , n26461 , n26462 , n26463 , n26464 , n26465 , n26466 , n26467 , n26468 , n26469 , n26470 , n26471 , n26472 , n26473 , n26474 , n26475 , n26476 , n26477 , n26478 , n26479 , n26480 , n26481 , n26482 , n26483 , n26484 , n26485 , n26486 , n26487 , n26488 , n26489 , n26490 , n26491 , n26492 , n26493 , n26494 , n26495 , n26496 , n26497 , n26498 , n26499 , n26500 , n26501 , n26502 , n26503 , n26504 , n26505 , n26506 , n26507 , n26508 , n26509 , n26510 , n26511 , n26512 , n26513 , n26514 , n26515 , n26516 , n26517 , n26518 , n26519 , n26520 , n26521 , n26522 , n26523 , n26524 , n26525 , n26526 , n26527 , n26528 , n26529 , n26530 , n26531 , n26532 , n26533 , n26534 , n26535 , n26536 , n26537 , n26538 , n26539 , n26540 , n26541 , n26542 , n26543 , n26544 , n26545 , n26546 , n26547 , n26548 , n26549 , n26550 , n26551 , n26552 , n26553 , n26554 , n26555 , n26556 , n26557 , n26558 , n26559 , n26560 , n26561 , n26562 , n26563 , n26564 , n26565 , n26566 , n26567 , n26568 , n26569 , n26570 , n26571 , n26572 , n26573 , n26574 , n26575 , n26576 , n26577 , n26578 , n26579 , n26580 , n26581 , n26582 , n26583 , n26584 , n26585 , n26586 , n26587 , n26588 , n26589 , n26590 , n26591 , n26592 , n26593 , n26594 , n26595 , n26596 , n26597 , n26598 , n26599 , n26600 , n26601 , n26602 , n26603 , n26604 , n26605 , n26606 , n26607 , n26608 , n26609 , n26610 , n26611 , n26612 , n26613 , n26614 , n26615 , n26616 , n26617 , n26618 , n26619 , n26620 , n26621 , n26622 , n26623 , n26624 , n26625 , n26626 , n26627 , n26628 , n26629 , n26630 , n26631 , n26632 , n26633 , n26634 , n26635 , n26636 , n26637 , n26638 , n26639 , n26640 , n26641 , n26642 , n26643 , n26644 , n26645 , n26646 , n26647 , n26648 , n26649 , n26650 , n26651 , n26652 , n26653 , n26654 , n26655 , n26656 , n26657 , n26658 , n26659 , n26660 , n26661 , n26662 , n26663 , n26664 , n26665 , n26666 , n26667 , n26668 , n26669 , n26670 , n26671 , n26672 , n26673 , n26674 , n26675 , n26676 , n26677 , n26678 , n26679 , n26680 , n26681 , n26682 , n26683 , n26684 , n26685 , n26686 , n26687 , n26688 , n26689 , n26690 , n26691 , n26692 , n26693 , n26694 , n26695 , n26696 , n26697 , n26698 , n26699 , n26700 , n26701 , n26702 , n26703 , n26704 , n26705 , n26706 , n26707 , n26708 , n26709 , n26710 , n26711 , n26712 , n26713 , n26714 , n26715 , n26716 , n26717 , n26718 , n26719 , n26720 , n26721 , n26722 , n26723 , n26724 , n26725 , n26726 , n26727 , n26728 , n26729 , n26730 , n26731 , n26732 , n26733 , n26734 , n26735 , n26736 , n26737 , n26738 , n26739 , n26740 , n26741 , n26742 , n26743 , n26744 , n26745 , n26746 , n26747 , n26748 , n26749 , n26750 , n26751 , n26752 , n26753 , n26754 , n26755 , n26756 , n26757 , n26758 , n26759 , n26760 , n26761 , n26762 , n26763 , n26764 , n26765 , n26766 , n26767 , n26768 , n26769 , n26770 , n26771 , n26772 , n26773 , n26774 , n26775 , n26776 , n26777 , n26778 , n26779 , n26780 , n26781 , n26782 , n26783 , n26784 , n26785 , n26786 , n26787 , n26788 , n26789 , n26790 , n26791 , n26792 , n26793 , n26794 , n26795 , n26796 , n26797 , n26798 , n26799 , n26800 , n26801 , n26802 , n26803 , n26804 , n26805 , n26806 , n26807 , n26808 , n26809 , n26810 , n26811 , n26812 , n26813 , n26814 , n26815 , n26816 , n26817 , n26818 , n26819 , n26820 , n26821 , n26822 , n26823 , n26824 , n26825 , n26826 , n26827 , n26828 , n26829 , n26830 , n26831 , n26832 , n26833 , n26834 , n26835 , n26836 , n26837 , n26838 , n26839 , n26840 , n26841 , n26842 , n26843 , n26844 , n26845 , n26846 , n26847 , n26848 , n26849 , n26850 , n26851 , n26852 , n26853 , n26854 , n26855 , n26856 , n26857 , n26858 , n26859 , n26860 , n26861 , n26862 , n26863 , n26864 , n26865 , n26866 , n26867 , n26868 , n26869 , n26870 , n26871 , n26872 , n26873 , n26874 , n26875 , n26876 , n26877 , n26878 , n26879 , n26880 , n26881 , n26882 , n26883 , n26884 , n26885 , n26886 , n26887 , n26888 , n26889 , n26890 , n26891 , n26892 , n26893 , n26894 , n26895 , n26896 , n26897 , n26898 , n26899 , n26900 , n26901 , n26902 , n26903 , n26904 , n26905 , n26906 , n26907 , n26908 , n26909 , n26910 , n26911 , n26912 , n26913 , n26914 , n26915 , n26916 , n26917 , n26918 , n26919 , n26920 , n26921 , n26922 , n26923 , n26924 , n26925 , n26926 , n26927 , n26928 , n26929 , n26930 , n26931 , n26932 , n26933 , n26934 , n26935 , n26936 , n26937 , n26938 , n26939 , n26940 , n26941 , n26942 , n26943 , n26944 , n26945 , n26946 , n26947 , n26948 , n26949 , n26950 , n26951 , n26952 , n26953 , n26954 , n26955 , n26956 , n26957 , n26958 , n26959 , n26960 , n26961 , n26962 , n26963 , n26964 , n26965 , n26966 , n26967 , n26968 , n26969 , n26970 , n26971 , n26972 , n26973 , n26974 , n26975 , n26976 , n26977 , n26978 , n26979 , n26980 , n26981 , n26982 , n26983 , n26984 , n26985 , n26986 , n26987 , n26988 , n26989 , n26990 , n26991 , n26992 , n26993 , n26994 , n26995 , n26996 , n26997 , n26998 , n26999 , n27000 , n27001 , n27002 , n27003 , n27004 , n27005 , n27006 , n27007 , n27008 , n27009 , n27010 , n27011 , n27012 , n27013 , n27014 , n27015 , n27016 , n27017 , n27018 , n27019 , n27020 , n27021 , n27022 , n27023 , n27024 , n27025 , n27026 , n27027 , n27028 , n27029 , n27030 , n27031 , n27032 , n27033 , n27034 , n27035 , n27036 , n27037 , n27038 , n27039 , n27040 , n27041 , n27042 , n27043 , n27044 , n27045 , n27046 , n27047 , n27048 , n27049 , n27050 , n27051 , n27052 , n27053 , n27054 , n27055 , n27056 , n27057 , n27058 , n27059 , n27060 , n27061 , n27062 , n27063 , n27064 , n27065 , n27066 , n27067 , n27068 , n27069 , n27070 , n27071 , n27072 , n27073 , n27074 , n27075 , n27076 , n27077 , n27078 , n27079 , n27080 , n27081 , n27082 , n27083 , n27084 , n27085 , n27086 , n27087 , n27088 , n27089 , n27090 , n27091 , n27092 , n27093 , n27094 , n27095 , n27096 , n27097 , n27098 , n27099 , n27100 , n27101 , n27102 , n27103 , n27104 , n27105 , n27106 , n27107 , n27108 , n27109 , n27110 , n27111 , n27112 , n27113 , n27114 , n27115 , n27116 , n27117 , n27118 , n27119 , n27120 , n27121 , n27122 , n27123 , n27124 , n27125 , n27126 , n27127 , n27128 , n27129 , n27130 , n27131 , n27132 , n27133 , n27134 , n27135 , n27136 , n27137 , n27138 , n27139 , n27140 , n27141 , n27142 , n27143 , n27144 , n27145 , n27146 , n27147 , n27148 , n27149 , n27150 , n27151 , n27152 , n27153 , n27154 , n27155 , n27156 , n27157 , n27158 , n27159 , n27160 , n27161 , n27162 , n27163 , n27164 , n27165 , n27166 , n27167 , n27168 , n27169 , n27170 , n27171 , n27172 , n27173 , n27174 , n27175 , n27176 , n27177 , n27178 , n27179 , n27180 , n27181 , n27182 , n27183 , n27184 , n27185 , n27186 , n27187 , n27188 , n27189 , n27190 , n27191 , n27192 , n27193 , n27194 , n27195 , n27196 , n27197 , n27198 , n27199 , n27200 , n27201 , n27202 , n27203 , n27204 , n27205 , n27206 , n27207 , n27208 , n27209 , n27210 , n27211 , n27212 , n27213 , n27214 , n27215 , n27216 , n27217 , n27218 , n27219 , n27220 , n27221 , n27222 , n27223 , n27224 , n27225 , n27226 , n27227 , n27228 , n27229 , n27230 , n27231 , n27232 , n27233 , n27234 , n27235 , n27236 , n27237 , n27238 , n27239 , n27240 , n27241 , n27242 , n27243 , n27244 , n27245 , n27246 , n27247 , n27248 , n27249 , n27250 , n27251 , n27252 , n27253 , n27254 , n27255 , n27256 , n27257 , n27258 , n27259 , n27260 , n27261 , n27262 , n27263 , n27264 , n27265 , n27266 , n27267 , n27268 , n27269 , n27270 , n27271 , n27272 , n27273 , n27274 , n27275 , n27276 , n27277 , n27278 , n27279 , n27280 , n27281 , n27282 , n27283 , n27284 , n27285 , n27286 , n27287 , n27288 , n27289 , n27290 , n27291 , n27292 , n27293 , n27294 , n27295 , n27296 , n27297 , n27298 , n27299 , n27300 , n27301 , n27302 , n27303 , n27304 , n27305 , n27306 , n27307 , n27308 , n27309 , n27310 , n27311 , n27312 , n27313 , n27314 , n27315 , n27316 , n27317 , n27318 , n27319 , n27320 , n27321 , n27322 , n27323 , n27324 , n27325 , n27326 , n27327 , n27328 , n27329 , n27330 , n27331 , n27332 , n27333 , n27334 , n27335 , n27336 , n27337 , n27338 , n27339 , n27340 , n27341 , n27342 , n27343 , n27344 , n27345 , n27346 , n27347 , n27348 , n27349 , n27350 , n27351 , n27352 , n27353 , n27354 , n27355 , n27356 , n27357 , n27358 , n27359 , n27360 , n27361 , n27362 , n27363 , n27364 , n27365 , n27366 , n27367 , n27368 , n27369 , n27370 , n27371 , n27372 , n27373 , n27374 , n27375 , n27376 , n27377 , n27378 , n27379 , n27380 , n27381 , n27382 , n27383 , n27384 , n27385 , n27386 , n27387 , n27388 , n27389 , n27390 , n27391 , n27392 , n27393 , n27394 , n27395 , n27396 , n27397 , n27398 , n27399 , n27400 , n27401 , n27402 , n27403 , n27404 , n27405 , n27406 , n27407 , n27408 , n27409 , n27410 , n27411 , n27412 , n27413 , n27414 , n27415 , n27416 , n27417 , n27418 , n27419 , n27420 , n27421 , n27422 , n27423 , n27424 , n27425 , n27426 , n27427 , n27428 , n27429 , n27430 , n27431 , n27432 , n27433 , n27434 , n27435 , n27436 , n27437 , n27438 , n27439 , n27440 , n27441 , n27442 , n27443 , n27444 , n27445 , n27446 , n27447 , n27448 , n27449 , n27450 , n27451 , n27452 , n27453 , n27454 , n27455 , n27456 , n27457 , n27458 , n27459 , n27460 , n27461 , n27462 , n27463 , n27464 , n27465 , n27466 , n27467 , n27468 , n27469 , n27470 , n27471 , n27472 , n27473 , n27474 , n27475 , n27476 , n27477 , n27478 , n27479 , n27480 , n27481 , n27482 , n27483 , n27484 , n27485 , n27486 , n27487 , n27488 , n27489 , n27490 , n27491 , n27492 , n27493 , n27494 , n27495 , n27496 , n27497 , n27498 , n27499 , n27500 , n27501 , n27502 , n27503 , n27504 , n27505 , n27506 , n27507 , n27508 , n27509 , n27510 , n27511 , n27512 , n27513 , n27514 , n27515 , n27516 , n27517 , n27518 , n27519 , n27520 , n27521 , n27522 , n27523 , n27524 , n27525 , n27526 , n27527 , n27528 , n27529 , n27530 , n27531 , n27532 , n27533 , n27534 , n27535 , n27536 , n27537 , n27538 , n27539 , n27540 , n27541 , n27542 , n27543 , n27544 , n27545 , n27546 , n27547 , n27548 , n27549 , n27550 , n27551 , n27552 , n27553 , n27554 , n27555 , n27556 , n27557 , n27558 , n27559 , n27560 , n27561 , n27562 , n27563 , n27564 , n27565 , n27566 , n27567 , n27568 , n27569 , n27570 , n27571 , n27572 , n27573 , n27574 , n27575 , n27576 , n27577 , n27578 , n27579 , n27580 , n27581 , n27582 , n27583 , n27584 , n27585 , n27586 , n27587 , n27588 , n27589 , n27590 , n27591 , n27592 , n27593 , n27594 , n27595 , n27596 , n27597 , n27598 , n27599 , n27600 , n27601 , n27602 , n27603 , n27604 , n27605 , n27606 , n27607 , n27608 , n27609 , n27610 , n27611 , n27612 , n27613 , n27614 , n27615 , n27616 , n27617 , n27618 , n27619 , n27620 , n27621 , n27622 , n27623 , n27624 , n27625 , n27626 , n27627 , n27628 , n27629 , n27630 , n27631 , n27632 , n27633 , n27634 , n27635 , n27636 , n27637 , n27638 , n27639 , n27640 , n27641 , n27642 , n27643 , n27644 , n27645 , n27646 , n27647 , n27648 , n27649 , n27650 , n27651 , n27652 , n27653 , n27654 , n27655 , n27656 , n27657 , n27658 , n27659 , n27660 , n27661 , n27662 , n27663 , n27664 , n27665 , n27666 , n27667 , n27668 , n27669 , n27670 , n27671 , n27672 , n27673 , n27674 , n27675 , n27676 , n27677 , n27678 , n27679 , n27680 , n27681 , n27682 , n27683 , n27684 , n27685 , n27686 , n27687 , n27688 , n27689 , n27690 , n27691 , n27692 , n27693 , n27694 , n27695 , n27696 , n27697 , n27698 , n27699 , n27700 , n27701 , n27702 , n27703 , n27704 , n27705 , n27706 , n27707 , n27708 , n27709 , n27710 , n27711 , n27712 , n27713 , n27714 , n27715 , n27716 , n27717 , n27718 , n27719 , n27720 , n27721 , n27722 , n27723 , n27724 , n27725 , n27726 , n27727 , n27728 , n27729 , n27730 , n27731 , n27732 , n27733 , n27734 , n27735 , n27736 , n27737 , n27738 , n27739 , n27740 , n27741 , n27742 , n27743 , n27744 , n27745 , n27746 , n27747 , n27748 , n27749 , n27750 , n27751 , n27752 , n27753 , n27754 , n27755 , n27756 , n27757 , n27758 , n27759 , n27760 , n27761 , n27762 , n27763 , n27764 , n27765 , n27766 , n27767 , n27768 , n27769 , n27770 , n27771 , n27772 , n27773 , n27774 , n27775 , n27776 , n27777 , n27778 , n27779 , n27780 , n27781 , n27782 , n27783 , n27784 , n27785 , n27786 , n27787 , n27788 , n27789 , n27790 , n27791 , n27792 , n27793 , n27794 , n27795 , n27796 , n27797 , n27798 , n27799 , n27800 , n27801 , n27802 , n27803 , n27804 , n27805 , n27806 , n27807 , n27808 , n27809 , n27810 , n27811 , n27812 , n27813 , n27814 , n27815 , n27816 , n27817 , n27818 , n27819 , n27820 , n27821 , n27822 , n27823 , n27824 , n27825 , n27826 , n27827 , n27828 , n27829 , n27830 , n27831 , n27832 , n27833 , n27834 , n27835 , n27836 , n27837 , n27838 , n27839 , n27840 , n27841 , n27842 , n27843 , n27844 , n27845 , n27846 , n27847 , n27848 , n27849 , n27850 , n27851 , n27852 , n27853 , n27854 , n27855 , n27856 , n27857 , n27858 , n27859 , n27860 , n27861 , n27862 , n27863 , n27864 , n27865 , n27866 , n27867 , n27868 , n27869 , n27870 , n27871 , n27872 , n27873 , n27874 , n27875 , n27876 , n27877 , n27878 , n27879 , n27880 , n27881 , n27882 , n27883 , n27884 , n27885 , n27886 , n27887 , n27888 , n27889 , n27890 , n27891 , n27892 , n27893 , n27894 , n27895 , n27896 , n27897 , n27898 , n27899 , n27900 , n27901 , n27902 , n27903 , n27904 , n27905 , n27906 , n27907 , n27908 , n27909 , n27910 , n27911 , n27912 , n27913 , n27914 , n27915 , n27916 , n27917 , n27918 , n27919 , n27920 , n27921 , n27922 , n27923 , n27924 , n27925 , n27926 , n27927 , n27928 , n27929 , n27930 , n27931 , n27932 , n27933 , n27934 , n27935 , n27936 , n27937 , n27938 , n27939 , n27940 , n27941 , n27942 , n27943 , n27944 , n27945 , n27946 , n27947 , n27948 , n27949 , n27950 , n27951 , n27952 , n27953 , n27954 , n27955 , n27956 , n27957 , n27958 , n27959 , n27960 , n27961 , n27962 , n27963 , n27964 , n27965 , n27966 , n27967 , n27968 , n27969 , n27970 , n27971 , n27972 , n27973 , n27974 , n27975 , n27976 , n27977 , n27978 , n27979 , n27980 , n27981 , n27982 , n27983 , n27984 , n27985 , n27986 , n27987 , n27988 , n27989 , n27990 , n27991 , n27992 , n27993 , n27994 , n27995 , n27996 , n27997 , n27998 , n27999 , n28000 , n28001 , n28002 , n28003 , n28004 , n28005 , n28006 , n28007 , n28008 , n28009 , n28010 , n28011 , n28012 , n28013 , n28014 , n28015 , n28016 , n28017 , n28018 , n28019 , n28020 , n28021 , n28022 , n28023 , n28024 , n28025 , n28026 , n28027 , n28028 , n28029 , n28030 , n28031 , n28032 , n28033 , n28034 , n28035 , n28036 , n28037 , n28038 , n28039 , n28040 , n28041 , n28042 , n28043 , n28044 , n28045 , n28046 , n28047 , n28048 , n28049 , n28050 , n28051 , n28052 , n28053 , n28054 , n28055 , n28056 , n28057 , n28058 , n28059 , n28060 , n28061 , n28062 , n28063 , n28064 , n28065 , n28066 , n28067 , n28068 , n28069 , n28070 , n28071 , n28072 , n28073 , n28074 , n28075 , n28076 , n28077 , n28078 , n28079 , n28080 , n28081 , n28082 , n28083 , n28084 , n28085 , n28086 , n28087 , n28088 , n28089 , n28090 , n28091 , n28092 , n28093 , n28094 , n28095 , n28096 , n28097 , n28098 , n28099 , n28100 , n28101 , n28102 , n28103 , n28104 , n28105 , n28106 , n28107 , n28108 , n28109 , n28110 , n28111 , n28112 , n28113 , n28114 , n28115 , n28116 , n28117 , n28118 , n28119 , n28120 , n28121 , n28122 , n28123 , n28124 , n28125 , n28126 , n28127 , n28128 , n28129 , n28130 , n28131 , n28132 , n28133 , n28134 , n28135 , n28136 , n28137 , n28138 , n28139 , n28140 , n28141 , n28142 , n28143 , n28144 , n28145 , n28146 , n28147 , n28148 , n28149 , n28150 , n28151 , n28152 , n28153 , n28154 , n28155 , n28156 , n28157 , n28158 , n28159 , n28160 , n28161 , n28162 , n28163 , n28164 , n28165 , n28166 , n28167 , n28168 , n28169 , n28170 , n28171 , n28172 , n28173 , n28174 , n28175 , n28176 , n28177 , n28178 , n28179 , n28180 , n28181 , n28182 , n28183 , n28184 , n28185 , n28186 , n28187 , n28188 , n28189 , n28190 , n28191 , n28192 , n28193 , n28194 , n28195 , n28196 , n28197 , n28198 , n28199 , n28200 , n28201 , n28202 , n28203 , n28204 , n28205 , n28206 , n28207 , n28208 , n28209 , n28210 , n28211 , n28212 , n28213 , n28214 , n28215 , n28216 , n28217 , n28218 , n28219 , n28220 , n28221 , n28222 , n28223 , n28224 , n28225 , n28226 , n28227 , n28228 , n28229 , n28230 , n28231 , n28232 , n28233 , n28234 , n28235 , n28236 , n28237 , n28238 , n28239 , n28240 , n28241 , n28242 , n28243 , n28244 , n28245 , n28246 , n28247 , n28248 , n28249 , n28250 , n28251 , n28252 , n28253 , n28254 , n28255 , n28256 , n28257 , n28258 , n28259 , n28260 , n28261 , n28262 , n28263 , n28264 , n28265 , n28266 , n28267 , n28268 , n28269 , n28270 , n28271 , n28272 , n28273 , n28274 , n28275 , n28276 , n28277 , n28278 , n28279 , n28280 , n28281 , n28282 , n28283 , n28284 , n28285 , n28286 , n28287 , n28288 , n28289 , n28290 , n28291 , n28292 , n28293 , n28294 , n28295 , n28296 , n28297 , n28298 , n28299 , n28300 , n28301 , n28302 , n28303 , n28304 , n28305 , n28306 , n28307 , n28308 , n28309 , n28310 , n28311 , n28312 , n28313 , n28314 , n28315 , n28316 , n28317 , n28318 , n28319 , n28320 , n28321 , n28322 , n28323 , n28324 , n28325 , n28326 , n28327 , n28328 , n28329 , n28330 , n28331 , n28332 , n28333 , n28334 , n28335 , n28336 , n28337 , n28338 , n28339 , n28340 , n28341 , n28342 , n28343 , n28344 , n28345 , n28346 , n28347 , n28348 , n28349 , n28350 , n28351 , n28352 , n28353 , n28354 , n28355 , n28356 , n28357 , n28358 , n28359 , n28360 , n28361 , n28362 , n28363 , n28364 , n28365 , n28366 , n28367 , n28368 , n28369 , n28370 , n28371 , n28372 , n28373 , n28374 , n28375 , n28376 , n28377 , n28378 , n28379 , n28380 , n28381 , n28382 , n28383 , n28384 , n28385 , n28386 , n28387 , n28388 , n28389 , n28390 , n28391 , n28392 , n28393 , n28394 , n28395 , n28396 , n28397 , n28398 , n28399 , n28400 , n28401 , n28402 , n28403 , n28404 , n28405 , n28406 , n28407 , n28408 , n28409 , n28410 , n28411 , n28412 , n28413 , n28414 , n28415 , n28416 , n28417 , n28418 , n28419 , n28420 , n28421 , n28422 , n28423 , n28424 , n28425 , n28426 , n28427 , n28428 , n28429 , n28430 , n28431 , n28432 , n28433 , n28434 , n28435 , n28436 , n28437 , n28438 , n28439 , n28440 , n28441 , n28442 , n28443 , n28444 , n28445 , n28446 , n28447 , n28448 , n28449 , n28450 , n28451 , n28452 , n28453 , n28454 , n28455 , n28456 , n28457 , n28458 , n28459 , n28460 , n28461 , n28462 , n28463 , n28464 , n28465 , n28466 , n28467 , n28468 , n28469 , n28470 , n28471 , n28472 , n28473 , n28474 , n28475 , n28476 , n28477 , n28478 , n28479 , n28480 , n28481 , n28482 , n28483 , n28484 , n28485 , n28486 , n28487 , n28488 , n28489 , n28490 , n28491 , n28492 , n28493 , n28494 , n28495 , n28496 , n28497 , n28498 , n28499 , n28500 , n28501 , n28502 , n28503 , n28504 , n28505 , n28506 , n28507 , n28508 , n28509 , n28510 , n28511 , n28512 , n28513 , n28514 , n28515 , n28516 , n28517 , n28518 , n28519 , n28520 , n28521 , n28522 , n28523 , n28524 , n28525 , n28526 , n28527 , n28528 , n28529 , n28530 , n28531 , n28532 , n28533 , n28534 , n28535 , n28536 , n28537 , n28538 , n28539 , n28540 , n28541 , n28542 , n28543 , n28544 , n28545 , n28546 , n28547 , n28548 , n28549 , n28550 , n28551 , n28552 , n28553 , n28554 , n28555 , n28556 , n28557 , n28558 , n28559 , n28560 , n28561 , n28562 , n28563 , n28564 , n28565 , n28566 , n28567 , n28568 , n28569 , n28570 , n28571 , n28572 , n28573 , n28574 , n28575 , n28576 , n28577 , n28578 , n28579 , n28580 , n28581 , n28582 , n28583 , n28584 , n28585 , n28586 , n28587 , n28588 , n28589 , n28590 , n28591 , n28592 , n28593 , n28594 , n28595 , n28596 , n28597 , n28598 , n28599 , n28600 , n28601 , n28602 , n28603 , n28604 , n28605 , n28606 , n28607 , n28608 , n28609 , n28610 , n28611 , n28612 , n28613 , n28614 , n28615 , n28616 , n28617 , n28618 , n28619 , n28620 , n28621 , n28622 , n28623 , n28624 , n28625 , n28626 , n28627 , n28628 , n28629 , n28630 , n28631 , n28632 , n28633 , n28634 , n28635 , n28636 , n28637 , n28638 , n28639 , n28640 , n28641 , n28642 , n28643 , n28644 , n28645 , n28646 , n28647 , n28648 , n28649 , n28650 , n28651 , n28652 , n28653 , n28654 , n28655 , n28656 , n28657 , n28658 , n28659 , n28660 , n28661 , n28662 , n28663 , n28664 , n28665 , n28666 , n28667 , n28668 , n28669 , n28670 , n28671 , n28672 , n28673 , n28674 , n28675 , n28676 , n28677 , n28678 , n28679 , n28680 , n28681 , n28682 , n28683 , n28684 , n28685 , n28686 , n28687 , n28688 , n28689 , n28690 , n28691 , n28692 , n28693 , n28694 , n28695 , n28696 , n28697 , n28698 , n28699 , n28700 , n28701 , n28702 , n28703 , n28704 , n28705 , n28706 , n28707 , n28708 , n28709 , n28710 , n28711 , n28712 , n28713 , n28714 , n28715 , n28716 , n28717 , n28718 , n28719 , n28720 , n28721 , n28722 , n28723 , n28724 , n28725 , n28726 , n28727 , n28728 , n28729 , n28730 , n28731 , n28732 , n28733 , n28734 , n28735 , n28736 , n28737 , n28738 , n28739 , n28740 , n28741 , n28742 , n28743 , n28744 , n28745 , n28746 , n28747 , n28748 , n28749 , n28750 , n28751 , n28752 , n28753 , n28754 , n28755 , n28756 , n28757 , n28758 , n28759 , n28760 , n28761 , n28762 , n28763 , n28764 , n28765 , n28766 , n28767 , n28768 , n28769 , n28770 , n28771 , n28772 , n28773 , n28774 , n28775 , n28776 , n28777 , n28778 , n28779 , n28780 , n28781 , n28782 , n28783 , n28784 , n28785 , n28786 , n28787 , n28788 , n28789 , n28790 , n28791 , n28792 , n28793 , n28794 , n28795 , n28796 , n28797 , n28798 , n28799 , n28800 , n28801 , n28802 , n28803 , n28804 , n28805 , n28806 , n28807 , n28808 , n28809 , n28810 , n28811 , n28812 , n28813 , n28814 , n28815 , n28816 , n28817 , n28818 , n28819 , n28820 , n28821 , n28822 , n28823 , n28824 , n28825 , n28826 , n28827 , n28828 , n28829 , n28830 , n28831 , n28832 , n28833 , n28834 , n28835 , n28836 , n28837 , n28838 , n28839 , n28840 , n28841 , n28842 , n28843 , n28844 , n28845 , n28846 , n28847 , n28848 , n28849 , n28850 , n28851 , n28852 , n28853 , n28854 , n28855 , n28856 , n28857 , n28858 , n28859 , n28860 , n28861 , n28862 , n28863 , n28864 , n28865 , n28866 , n28867 , n28868 , n28869 , n28870 , n28871 , n28872 , n28873 , n28874 , n28875 , n28876 , n28877 , n28878 , n28879 , n28880 , n28881 , n28882 , n28883 , n28884 , n28885 , n28886 , n28887 , n28888 , n28889 , n28890 , n28891 , n28892 , n28893 , n28894 , n28895 , n28896 , n28897 , n28898 , n28899 , n28900 , n28901 , n28902 , n28903 , n28904 , n28905 , n28906 , n28907 , n28908 , n28909 , n28910 , n28911 , n28912 , n28913 , n28914 , n28915 , n28916 , n28917 , n28918 , n28919 , n28920 , n28921 , n28922 , n28923 , n28924 , n28925 , n28926 , n28927 , n28928 , n28929 , n28930 , n28931 , n28932 , n28933 , n28934 , n28935 , n28936 , n28937 , n28938 , n28939 , n28940 , n28941 , n28942 , n28943 , n28944 , n28945 , n28946 , n28947 , n28948 , n28949 , n28950 , n28951 , n28952 , n28953 , n28954 , n28955 , n28956 , n28957 , n28958 , n28959 , n28960 , n28961 , n28962 , n28963 , n28964 , n28965 , n28966 , n28967 , n28968 , n28969 , n28970 , n28971 , n28972 , n28973 , n28974 , n28975 , n28976 , n28977 , n28978 , n28979 , n28980 , n28981 , n28982 , n28983 , n28984 , n28985 , n28986 , n28987 , n28988 , n28989 , n28990 , n28991 , n28992 , n28993 , n28994 , n28995 , n28996 , n28997 , n28998 , n28999 , n29000 , n29001 , n29002 , n29003 , n29004 , n29005 , n29006 , n29007 , n29008 , n29009 , n29010 , n29011 , n29012 , n29013 , n29014 , n29015 , n29016 , n29017 , n29018 , n29019 , n29020 , n29021 , n29022 , n29023 , n29024 , n29025 , n29026 , n29027 , n29028 , n29029 , n29030 , n29031 , n29032 , n29033 , n29034 , n29035 , n29036 , n29037 , n29038 , n29039 , n29040 , n29041 , n29042 , n29043 , n29044 , n29045 , n29046 , n29047 , n29048 , n29049 , n29050 , n29051 , n29052 , n29053 , n29054 , n29055 , n29056 , n29057 , n29058 , n29059 , n29060 , n29061 , n29062 , n29063 , n29064 , n29065 , n29066 , n29067 , n29068 , n29069 , n29070 , n29071 , n29072 , n29073 , n29074 , n29075 , n29076 , n29077 , n29078 , n29079 , n29080 , n29081 , n29082 , n29083 , n29084 , n29085 , n29086 , n29087 , n29088 , n29089 , n29090 , n29091 , n29092 , n29093 , n29094 , n29095 , n29096 , n29097 , n29098 , n29099 , n29100 , n29101 , n29102 , n29103 , n29104 , n29105 , n29106 , n29107 , n29108 , n29109 , n29110 , n29111 , n29112 , n29113 , n29114 , n29115 , n29116 , n29117 , n29118 , n29119 , n29120 , n29121 , n29122 , n29123 , n29124 , n29125 , n29126 , n29127 , n29128 , n29129 , n29130 , n29131 , n29132 , n29133 , n29134 , n29135 , n29136 , n29137 , n29138 , n29139 , n29140 , n29141 , n29142 , n29143 , n29144 , n29145 , n29146 , n29147 , n29148 , n29149 , n29150 , n29151 , n29152 , n29153 , n29154 , n29155 , n29156 , n29157 , n29158 , n29159 , n29160 , n29161 , n29162 , n29163 , n29164 , n29165 , n29166 , n29167 , n29168 , n29169 , n29170 , n29171 , n29172 , n29173 , n29174 , n29175 , n29176 , n29177 , n29178 , n29179 , n29180 , n29181 , n29182 , n29183 , n29184 , n29185 , n29186 , n29187 , n29188 , n29189 , n29190 , n29191 , n29192 , n29193 , n29194 , n29195 , n29196 , n29197 , n29198 , n29199 , n29200 , n29201 , n29202 , n29203 , n29204 , n29205 , n29206 , n29207 , n29208 , n29209 , n29210 , n29211 , n29212 , n29213 , n29214 , n29215 , n29216 , n29217 , n29218 , n29219 , n29220 , n29221 , n29222 , n29223 , n29224 , n29225 , n29226 , n29227 , n29228 , n29229 , n29230 , n29231 , n29232 , n29233 , n29234 , n29235 , n29236 , n29237 , n29238 , n29239 , n29240 , n29241 , n29242 , n29243 , n29244 , n29245 , n29246 , n29247 , n29248 , n29249 , n29250 , n29251 , n29252 , n29253 , n29254 , n29255 , n29256 , n29257 , n29258 , n29259 , n29260 , n29261 , n29262 , n29263 , n29264 , n29265 , n29266 , n29267 , n29268 , n29269 , n29270 , n29271 , n29272 , n29273 , n29274 , n29275 , n29276 , n29277 , n29278 , n29279 , n29280 , n29281 , n29282 , n29283 , n29284 , n29285 , n29286 , n29287 , n29288 , n29289 , n29290 , n29291 , n29292 , n29293 , n29294 , n29295 , n29296 , n29297 , n29298 , n29299 , n29300 , n29301 , n29302 , n29303 , n29304 , n29305 , n29306 , n29307 , n29308 , n29309 , n29310 , n29311 , n29312 , n29313 , n29314 , n29315 , n29316 , n29317 , n29318 , n29319 , n29320 , n29321 , n29322 , n29323 , n29324 , n29325 , n29326 , n29327 , n29328 , n29329 , n29330 , n29331 , n29332 , n29333 , n29334 , n29335 , n29336 , n29337 , n29338 , n29339 , n29340 , n29341 , n29342 , n29343 , n29344 , n29345 , n29346 , n29347 , n29348 , n29349 , n29350 , n29351 , n29352 , n29353 , n29354 , n29355 , n29356 , n29357 , n29358 , n29359 , n29360 , n29361 , n29362 , n29363 , n29364 , n29365 , n29366 , n29367 , n29368 , n29369 , n29370 , n29371 , n29372 , n29373 , n29374 , n29375 , n29376 , n29377 , n29378 , n29379 , n29380 , n29381 , n29382 , n29383 , n29384 , n29385 , n29386 , n29387 , n29388 , n29389 , n29390 , n29391 , n29392 , n29393 , n29394 , n29395 , n29396 , n29397 , n29398 , n29399 , n29400 , n29401 , n29402 , n29403 , n29404 , n29405 , n29406 , n29407 , n29408 , n29409 , n29410 , n29411 , n29412 , n29413 , n29414 , n29415 , n29416 , n29417 , n29418 , n29419 , n29420 , n29421 , n29422 , n29423 , n29424 , n29425 , n29426 , n29427 , n29428 , n29429 , n29430 , n29431 , n29432 , n29433 , n29434 , n29435 , n29436 , n29437 , n29438 , n29439 , n29440 , n29441 , n29442 , n29443 , n29444 , n29445 , n29446 , n29447 , n29448 , n29449 , n29450 , n29451 , n29452 , n29453 , n29454 , n29455 , n29456 , n29457 , n29458 , n29459 , n29460 , n29461 , n29462 , n29463 , n29464 , n29465 , n29466 , n29467 , n29468 , n29469 , n29470 , n29471 , n29472 , n29473 , n29474 , n29475 , n29476 , n29477 , n29478 , n29479 , n29480 , n29481 , n29482 , n29483 , n29484 , n29485 , n29486 , n29487 , n29488 , n29489 , n29490 , n29491 , n29492 , n29493 , n29494 , n29495 , n29496 , n29497 , n29498 , n29499 , n29500 , n29501 , n29502 , n29503 , n29504 , n29505 , n29506 , n29507 , n29508 , n29509 , n29510 , n29511 , n29512 , n29513 , n29514 , n29515 , n29516 , n29517 , n29518 , n29519 , n29520 , n29521 , n29522 , n29523 , n29524 , n29525 , n29526 , n29527 , n29528 , n29529 , n29530 , n29531 , n29532 , n29533 , n29534 , n29535 , n29536 , n29537 , n29538 , n29539 , n29540 , n29541 , n29542 , n29543 , n29544 , n29545 , n29546 , n29547 , n29548 , n29549 , n29550 , n29551 , n29552 , n29553 , n29554 , n29555 , n29556 , n29557 , n29558 , n29559 , n29560 , n29561 , n29562 , n29563 , n29564 , n29565 , n29566 , n29567 , n29568 , n29569 , n29570 , n29571 , n29572 , n29573 , n29574 , n29575 , n29576 , n29577 , n29578 , n29579 , n29580 , n29581 , n29582 , n29583 , n29584 , n29585 , n29586 , n29587 , n29588 , n29589 , n29590 , n29591 , n29592 , n29593 , n29594 , n29595 , n29596 , n29597 , n29598 , n29599 , n29600 , n29601 , n29602 , n29603 , n29604 , n29605 , n29606 , n29607 , n29608 , n29609 , n29610 , n29611 , n29612 , n29613 , n29614 , n29615 , n29616 , n29617 , n29618 , n29619 , n29620 , n29621 , n29622 , n29623 , n29624 , n29625 , n29626 , n29627 , n29628 , n29629 , n29630 , n29631 , n29632 , n29633 , n29634 , n29635 , n29636 , n29637 , n29638 , n29639 , n29640 , n29641 , n29642 , n29643 , n29644 , n29645 , n29646 , n29647 , n29648 , n29649 , n29650 , n29651 , n29652 , n29653 , n29654 , n29655 , n29656 , n29657 , n29658 , n29659 , n29660 , n29661 , n29662 , n29663 , n29664 , n29665 , n29666 , n29667 , n29668 , n29669 , n29670 , n29671 , n29672 , n29673 , n29674 , n29675 , n29676 , n29677 , n29678 , n29679 , n29680 , n29681 , n29682 , n29683 , n29684 , n29685 , n29686 , n29687 , n29688 , n29689 , n29690 , n29691 , n29692 , n29693 , n29694 , n29695 , n29696 , n29697 , n29698 , n29699 , n29700 , n29701 , n29702 , n29703 , n29704 , n29705 , n29706 , n29707 , n29708 , n29709 , n29710 , n29711 , n29712 , n29713 , n29714 , n29715 , n29716 , n29717 , n29718 , n29719 , n29720 , n29721 , n29722 , n29723 , n29724 , n29725 , n29726 , n29727 , n29728 , n29729 , n29730 , n29731 , n29732 , n29733 , n29734 , n29735 , n29736 , n29737 , n29738 , n29739 , n29740 , n29741 , n29742 , n29743 , n29744 , n29745 , n29746 , n29747 , n29748 , n29749 , n29750 , n29751 , n29752 , n29753 , n29754 , n29755 , n29756 , n29757 , n29758 , n29759 , n29760 , n29761 , n29762 , n29763 , n29764 , n29765 , n29766 , n29767 , n29768 , n29769 , n29770 , n29771 , n29772 , n29773 , n29774 , n29775 , n29776 ;
  assign n33 = x11 & ~x12 ;
  assign n34 = ~x11 & x12 ;
  assign n35 = n33 | n34 ;
  assign n36 = x13 & ~x14 ;
  assign n37 = ~x13 & x14 ;
  assign n38 = n36 | n37 ;
  assign n39 = n35 & n38 ;
  assign n40 = x23 & ~x26 ;
  assign n41 = x24 & x25 ;
  assign n42 = n40 & n41 ;
  assign n43 = x27 | x28 ;
  assign n44 = x29 | x30 ;
  assign n45 = n43 | n44 ;
  assign n46 = n42 & ~n45 ;
  assign n47 = x23 & x26 ;
  assign n48 = x24 | x25 ;
  assign n49 = n47 & ~n48 ;
  assign n50 = x27 & x28 ;
  assign n51 = ~n44 & n50 ;
  assign n52 = n49 & n51 ;
  assign n53 = ~x24 & x25 ;
  assign n54 = n47 & n53 ;
  assign n55 = n51 & n54 ;
  assign n56 = n40 & ~n48 ;
  assign n57 = ~n45 & n56 ;
  assign n58 = ~n45 & n49 ;
  assign n59 = n57 | n58 ;
  assign n60 = x24 & ~x25 ;
  assign n61 = n40 & n60 ;
  assign n62 = n51 & n61 ;
  assign n63 = x23 | x26 ;
  assign n64 = n53 & ~n63 ;
  assign n65 = n51 & n64 ;
  assign n66 = n62 | n65 ;
  assign n67 = n59 | n66 ;
  assign n68 = n55 | n67 ;
  assign n69 = n52 | n68 ;
  assign n70 = n46 | n69 ;
  assign n71 = ~x23 & x26 ;
  assign n72 = n60 & n71 ;
  assign n73 = x27 & ~x28 ;
  assign n74 = x29 & ~x30 ;
  assign n75 = n73 & n74 ;
  assign n76 = n72 & n75 ;
  assign n77 = n56 & n75 ;
  assign n78 = n41 & n47 ;
  assign n79 = ~x27 & x28 ;
  assign n80 = n74 & n79 ;
  assign n81 = n78 & n80 ;
  assign n82 = n77 | n81 ;
  assign n83 = n64 & n80 ;
  assign n84 = n41 & n71 ;
  assign n85 = n80 & n84 ;
  assign n86 = n83 | n85 ;
  assign n87 = n82 | n86 ;
  assign n88 = n76 | n87 ;
  assign n89 = n41 & ~n63 ;
  assign n90 = n75 & n89 ;
  assign n91 = n47 & n60 ;
  assign n92 = n75 & n91 ;
  assign n93 = n90 | n92 ;
  assign n94 = n54 & n80 ;
  assign n95 = n40 & n53 ;
  assign n96 = n80 & n95 ;
  assign n97 = n94 | n96 ;
  assign n98 = n93 | n97 ;
  assign n99 = n72 & n80 ;
  assign n100 = n61 & n80 ;
  assign n101 = n99 | n100 ;
  assign n102 = n64 & n75 ;
  assign n103 = n75 & n84 ;
  assign n104 = n102 | n103 ;
  assign n105 = n101 | n104 ;
  assign n106 = n98 | n105 ;
  assign n107 = n88 | n106 ;
  assign n108 = n80 & n89 ;
  assign n109 = ~n48 & n71 ;
  assign n110 = n75 & n109 ;
  assign n111 = n75 & n78 ;
  assign n112 = n56 & n80 ;
  assign n113 = n48 | n63 ;
  assign n114 = n80 & ~n113 ;
  assign n115 = n112 | n114 ;
  assign n116 = n111 | n115 ;
  assign n117 = n110 | n116 ;
  assign n118 = n108 | n117 ;
  assign n119 = n107 | n118 ;
  assign n120 = n75 & ~n113 ;
  assign n121 = ~n43 & n74 ;
  assign n122 = n72 & n121 ;
  assign n123 = n120 | n122 ;
  assign n124 = n119 | n123 ;
  assign n125 = n51 & n84 ;
  assign n126 = n56 & n121 ;
  assign n127 = n125 | n126 ;
  assign n128 = n42 & n121 ;
  assign n129 = n78 & n121 ;
  assign n130 = n128 | n129 ;
  assign n131 = n127 | n130 ;
  assign n132 = n95 & n121 ;
  assign n133 = ~n113 & n121 ;
  assign n134 = n51 & n78 ;
  assign n135 = n133 | n134 ;
  assign n136 = n132 | n135 ;
  assign n137 = n131 | n136 ;
  assign n138 = n53 & n71 ;
  assign n139 = n121 & n138 ;
  assign n140 = n91 & n121 ;
  assign n141 = n139 | n140 ;
  assign n142 = n109 & n121 ;
  assign n143 = n64 & n121 ;
  assign n144 = n142 | n143 ;
  assign n145 = n61 & n121 ;
  assign n146 = n49 & n121 ;
  assign n147 = n145 | n146 ;
  assign n148 = n144 | n147 ;
  assign n149 = n141 | n148 ;
  assign n150 = n137 | n149 ;
  assign n151 = n54 & n121 ;
  assign n152 = n89 & n121 ;
  assign n153 = n151 | n152 ;
  assign n154 = n150 | n153 ;
  assign n155 = n49 & n75 ;
  assign n156 = n50 & n74 ;
  assign n157 = ~n113 & n156 ;
  assign n158 = n155 | n157 ;
  assign n159 = n60 & ~n63 ;
  assign n160 = n75 & n159 ;
  assign n161 = n80 & n159 ;
  assign n162 = n160 | n161 ;
  assign n163 = n158 | n162 ;
  assign n164 = n75 & n95 ;
  assign n165 = n42 & n75 ;
  assign n166 = n164 | n165 ;
  assign n167 = n80 & n109 ;
  assign n168 = n80 & n138 ;
  assign n169 = n167 | n168 ;
  assign n170 = n166 | n169 ;
  assign n171 = n163 | n170 ;
  assign n172 = n42 & n80 ;
  assign n173 = n75 & n138 ;
  assign n174 = n54 & n75 ;
  assign n175 = n61 & n75 ;
  assign n176 = n174 | n175 ;
  assign n177 = n173 | n176 ;
  assign n178 = n172 | n177 ;
  assign n179 = n171 | n178 ;
  assign n180 = n80 & n91 ;
  assign n181 = n49 & n80 ;
  assign n182 = n180 | n181 ;
  assign n183 = n179 | n182 ;
  assign n184 = n154 | n183 ;
  assign n185 = n124 | n184 ;
  assign n186 = n84 & n121 ;
  assign n187 = n121 & n159 ;
  assign n188 = n186 | n187 ;
  assign n189 = n185 | n188 ;
  assign n190 = n51 & n138 ;
  assign n191 = n51 & n72 ;
  assign n192 = n190 | n191 ;
  assign n193 = n51 & n91 ;
  assign n194 = n51 & n89 ;
  assign n195 = n193 | n194 ;
  assign n196 = n192 | n195 ;
  assign n197 = n51 & n95 ;
  assign n198 = n51 & n109 ;
  assign n199 = n42 & n51 ;
  assign n200 = n198 | n199 ;
  assign n201 = n197 | n200 ;
  assign n202 = n196 | n201 ;
  assign n203 = ~n45 & n89 ;
  assign n204 = ~n45 & n95 ;
  assign n205 = n203 | n204 ;
  assign n206 = n89 & n156 ;
  assign n207 = n95 & n156 ;
  assign n208 = n42 & n156 ;
  assign n209 = n207 | n208 ;
  assign n210 = n206 | n209 ;
  assign n211 = n205 | n210 ;
  assign n212 = ~n45 & n61 ;
  assign n213 = ~n45 & n159 ;
  assign n214 = n212 | n213 ;
  assign n215 = ~n45 & n109 ;
  assign n216 = n214 | n215 ;
  assign n217 = n64 & n156 ;
  assign n218 = n109 & n156 ;
  assign n219 = n217 | n218 ;
  assign n220 = n216 | n219 ;
  assign n221 = n211 | n220 ;
  assign n222 = ~n45 & n64 ;
  assign n223 = n56 & n156 ;
  assign n224 = n61 & n156 ;
  assign n225 = n223 | n224 ;
  assign n226 = n45 | n113 ;
  assign n227 = n156 & n159 ;
  assign n228 = n226 & ~n227 ;
  assign n229 = ~n225 & n228 ;
  assign n230 = ~n222 & n229 ;
  assign n231 = ~n221 & n230 ;
  assign n232 = ( n189 & ~n202 ) | ( n189 & n231 ) | ( ~n202 & n231 ) ;
  assign n233 = ~n189 & n232 ;
  assign n234 = ~n70 & n233 ;
  assign n235 = ~x29 & x30 ;
  assign n236 = n50 & n235 ;
  assign n237 = n42 & n236 ;
  assign n238 = x29 & x30 ;
  assign n239 = ~n43 & n238 ;
  assign n240 = n95 & n239 ;
  assign n241 = n64 & n239 ;
  assign n242 = n84 & n236 ;
  assign n243 = n241 | n242 ;
  assign n244 = n138 & n236 ;
  assign n245 = n78 & n236 ;
  assign n246 = n244 | n245 ;
  assign n247 = n243 | n246 ;
  assign n248 = n240 | n247 ;
  assign n249 = ~n113 & n239 ;
  assign n250 = n89 & n239 ;
  assign n251 = n249 | n250 ;
  assign n252 = n159 & n239 ;
  assign n253 = n61 & n239 ;
  assign n254 = n252 | n253 ;
  assign n255 = n251 | n254 ;
  assign n256 = n248 | n255 ;
  assign n257 = n79 & n238 ;
  assign n258 = n42 & n257 ;
  assign n259 = n73 & n238 ;
  assign n260 = n54 & n259 ;
  assign n261 = n258 | n260 ;
  assign n262 = n61 & n257 ;
  assign n263 = ~n113 & n257 ;
  assign n264 = n262 | n263 ;
  assign n265 = n64 & n257 ;
  assign n266 = n49 & n257 ;
  assign n267 = n265 | n266 ;
  assign n268 = n264 | n267 ;
  assign n269 = n78 & n259 ;
  assign n270 = n109 & n257 ;
  assign n271 = n269 | n270 ;
  assign n272 = n268 | n271 ;
  assign n273 = n56 & n257 ;
  assign n274 = n138 & n259 ;
  assign n275 = n273 | n274 ;
  assign n276 = n84 & n259 ;
  assign n277 = n91 & n257 ;
  assign n278 = n276 | n277 ;
  assign n279 = n95 & n257 ;
  assign n280 = n89 & n257 ;
  assign n281 = n279 | n280 ;
  assign n282 = n159 & n257 ;
  assign n283 = n72 & n257 ;
  assign n284 = n282 | n283 ;
  assign n285 = n281 | n284 ;
  assign n286 = n278 | n285 ;
  assign n287 = ( ~n272 & n275 ) | ( ~n272 & n286 ) | ( n275 & n286 ) ;
  assign n288 = n272 | n287 ;
  assign n289 = n261 | n288 ;
  assign n290 = n256 | n289 ;
  assign n291 = n109 & n259 ;
  assign n292 = n42 & n259 ;
  assign n293 = n54 & n239 ;
  assign n294 = n292 | n293 ;
  assign n295 = n109 & n239 ;
  assign n296 = n72 & n259 ;
  assign n297 = n295 | n296 ;
  assign n298 = n294 | n297 ;
  assign n299 = n138 & n239 ;
  assign n300 = n61 & n259 ;
  assign n301 = ~n113 & n259 ;
  assign n302 = n300 | n301 ;
  assign n303 = n299 | n302 ;
  assign n304 = n298 | n303 ;
  assign n305 = n291 | n304 ;
  assign n306 = n89 & n259 ;
  assign n307 = n91 & n259 ;
  assign n308 = n306 | n307 ;
  assign n309 = n159 & n259 ;
  assign n310 = n84 & n239 ;
  assign n311 = n309 | n310 ;
  assign n312 = n308 | n311 ;
  assign n313 = n78 & n239 ;
  assign n314 = n72 & n239 ;
  assign n315 = n91 & n239 ;
  assign n316 = n314 | n315 ;
  assign n317 = n313 | n316 ;
  assign n318 = n312 | n317 ;
  assign n319 = n95 & n259 ;
  assign n320 = n49 & n259 ;
  assign n321 = n64 & n259 ;
  assign n322 = n320 | n321 ;
  assign n323 = n319 | n322 ;
  assign n324 = n318 | n323 ;
  assign n325 = n305 | n324 ;
  assign n326 = n56 & n259 ;
  assign n327 = n49 & n239 ;
  assign n328 = n214 | n327 ;
  assign n329 = n326 | n328 ;
  assign n330 = n57 | n329 ;
  assign n331 = n226 & ~n330 ;
  assign n332 = ~n325 & n331 ;
  assign n333 = ~n290 & n332 ;
  assign n334 = n42 & n239 ;
  assign n335 = n54 & n236 ;
  assign n336 = n334 | n335 ;
  assign n337 = n91 & n236 ;
  assign n338 = n56 & n239 ;
  assign n339 = n337 | n338 ;
  assign n340 = n336 | n339 ;
  assign n341 = n222 | n340 ;
  assign n342 = n333 & ~n341 ;
  assign n343 = n50 & n238 ;
  assign n344 = n42 & n343 ;
  assign n345 = n61 & n343 ;
  assign n346 = n109 & n343 ;
  assign n347 = n345 | n346 ;
  assign n348 = n344 | n347 ;
  assign n349 = n78 & n257 ;
  assign n350 = n54 & n257 ;
  assign n351 = n159 & n343 ;
  assign n352 = n350 | n351 ;
  assign n353 = n349 | n352 ;
  assign n354 = n348 | n353 ;
  assign n355 = n56 & n343 ;
  assign n356 = n64 & n343 ;
  assign n357 = n355 | n356 ;
  assign n358 = n95 & n343 ;
  assign n359 = ~n113 & n343 ;
  assign n360 = ( ~n357 & n358 ) | ( ~n357 & n359 ) | ( n358 & n359 ) ;
  assign n361 = n357 | n360 ;
  assign n362 = n354 | n361 ;
  assign n363 = ~n44 & n79 ;
  assign n364 = n42 & n363 ;
  assign n365 = n46 | n223 ;
  assign n366 = n89 & n343 ;
  assign n367 = n224 | n366 ;
  assign n368 = n365 | n367 ;
  assign n369 = n364 | n368 ;
  assign n370 = n227 | n369 ;
  assign n371 = n362 | n370 ;
  assign n372 = n103 | n217 ;
  assign n373 = n61 & n236 ;
  assign n374 = n100 | n373 ;
  assign n375 = n210 | n374 ;
  assign n376 = n88 | n375 ;
  assign n377 = n54 & n363 ;
  assign n378 = n204 | n377 ;
  assign n379 = n54 & n343 ;
  assign n380 = n84 & n257 ;
  assign n381 = n138 & n257 ;
  assign n382 = n380 | n381 ;
  assign n383 = n49 & n343 ;
  assign n384 = n84 & n343 ;
  assign n385 = n383 | n384 ;
  assign n386 = n382 | n385 ;
  assign n387 = n379 | n386 ;
  assign n388 = n378 | n387 ;
  assign n389 = n376 | n388 ;
  assign n390 = n56 & n363 ;
  assign n391 = n72 & n236 ;
  assign n392 = ~n44 & n73 ;
  assign n393 = n84 & n392 ;
  assign n394 = n391 | n393 ;
  assign n395 = n215 | n394 ;
  assign n396 = n390 | n395 ;
  assign n397 = ( ~n372 & n389 ) | ( ~n372 & n396 ) | ( n389 & n396 ) ;
  assign n398 = n372 | n397 ;
  assign n399 = n58 | n108 ;
  assign n400 = n51 & n56 ;
  assign n401 = n102 | n400 ;
  assign n402 = n399 | n401 ;
  assign n403 = n72 & n363 ;
  assign n404 = n91 & n363 ;
  assign n405 = n403 | n404 ;
  assign n406 = n115 | n405 ;
  assign n407 = n402 | n406 ;
  assign n408 = n61 & n363 ;
  assign n409 = n95 & n236 ;
  assign n410 = n203 | n409 ;
  assign n411 = n408 | n410 ;
  assign n412 = n110 | n411 ;
  assign n413 = n407 | n412 ;
  assign n414 = n99 | n218 ;
  assign n415 = n413 | n414 ;
  assign n416 = n72 & n343 ;
  assign n417 = n138 & n343 ;
  assign n418 = n416 | n417 ;
  assign n419 = n78 & n343 ;
  assign n420 = n91 & n343 ;
  assign n421 = n419 | n420 ;
  assign n422 = n418 | n421 ;
  assign n423 = n98 | n422 ;
  assign n424 = n415 | n423 ;
  assign n425 = n398 | n424 ;
  assign n426 = n371 | n425 ;
  assign n427 = n342 & ~n426 ;
  assign n428 = n89 & n236 ;
  assign n429 = n64 & n236 ;
  assign n430 = n111 | n429 ;
  assign n431 = n49 & n236 ;
  assign n432 = n109 & n236 ;
  assign n433 = n431 | n432 ;
  assign n434 = ~n113 & n363 ;
  assign n435 = n78 & n392 ;
  assign n436 = n434 | n435 ;
  assign n437 = n159 & n363 ;
  assign n438 = n78 & n363 ;
  assign n439 = n437 | n438 ;
  assign n440 = n436 | n439 ;
  assign n441 = n89 & n363 ;
  assign n442 = n64 & n363 ;
  assign n443 = n441 | n442 ;
  assign n444 = n54 & n392 ;
  assign n445 = n84 & n363 ;
  assign n446 = n444 | n445 ;
  assign n447 = n443 | n446 ;
  assign n448 = n440 | n447 ;
  assign n449 = n49 & n363 ;
  assign n450 = n138 & n363 ;
  assign n451 = n51 & ~n113 ;
  assign n452 = n51 & n159 ;
  assign n453 = n451 | n452 ;
  assign n454 = n450 | n453 ;
  assign n455 = n449 | n454 ;
  assign n456 = n448 | n455 ;
  assign n457 = n95 & n363 ;
  assign n458 = n109 & n363 ;
  assign n459 = n457 | n458 ;
  assign n460 = n456 | n459 ;
  assign n461 = n183 | n460 ;
  assign n462 = n433 | n461 ;
  assign n463 = n430 | n462 ;
  assign n464 = n428 | n463 ;
  assign n465 = n427 & ~n464 ;
  assign n466 = ~n237 & n465 ;
  assign n467 = n234 & ~n466 ;
  assign n468 = ~n113 & n236 ;
  assign n469 = n73 & n235 ;
  assign n470 = n56 & n469 ;
  assign n471 = n79 & n235 ;
  assign n472 = n49 & n471 ;
  assign n473 = n470 | n472 ;
  assign n474 = n468 | n473 ;
  assign n475 = n84 & n471 ;
  assign n476 = n89 & n471 ;
  assign n477 = n475 | n476 ;
  assign n478 = n95 & n471 ;
  assign n479 = n91 & n471 ;
  assign n480 = n478 | n479 ;
  assign n481 = n477 | n480 ;
  assign n482 = n56 & n236 ;
  assign n483 = n54 & n471 ;
  assign n484 = n109 & n471 ;
  assign n485 = n483 | n484 ;
  assign n486 = n482 | n485 ;
  assign n487 = n481 | n486 ;
  assign n488 = n138 & n471 ;
  assign n489 = n78 & n471 ;
  assign n490 = n72 & n471 ;
  assign n491 = n489 | n490 ;
  assign n492 = n488 | n491 ;
  assign n493 = n409 | n428 ;
  assign n494 = n433 | n493 ;
  assign n495 = n492 | n494 ;
  assign n496 = n487 | n495 ;
  assign n497 = n474 | n496 ;
  assign n498 = n138 & n469 ;
  assign n499 = n78 & n469 ;
  assign n500 = n109 & n469 ;
  assign n501 = n499 | n500 ;
  assign n502 = n498 | n501 ;
  assign n503 = n61 & n469 ;
  assign n504 = n54 & n469 ;
  assign n505 = n64 & n469 ;
  assign n506 = n504 | n505 ;
  assign n507 = n503 | n506 ;
  assign n508 = n502 | n507 ;
  assign n509 = n56 & n471 ;
  assign n510 = n95 & n469 ;
  assign n511 = n89 & n469 ;
  assign n512 = n510 | n511 ;
  assign n513 = n42 & n469 ;
  assign n514 = ~n113 & n471 ;
  assign n515 = n513 | n514 ;
  assign n516 = n512 | n515 ;
  assign n517 = n509 | n516 ;
  assign n518 = n508 | n517 ;
  assign n519 = n49 & n469 ;
  assign n520 = n84 & n469 ;
  assign n521 = n91 & n469 ;
  assign n522 = n72 & n469 ;
  assign n523 = n521 | n522 ;
  assign n524 = n520 | n523 ;
  assign n525 = n519 | n524 ;
  assign n526 = n518 | n525 ;
  assign n527 = n497 | n526 ;
  assign n528 = n64 & n471 ;
  assign n529 = n42 & n471 ;
  assign n530 = n159 & n471 ;
  assign n531 = n61 & n471 ;
  assign n532 = n530 | n531 ;
  assign n533 = n529 | n532 ;
  assign n534 = n528 | n533 ;
  assign n535 = n391 | n534 ;
  assign n536 = n429 | n535 ;
  assign n537 = n373 | n536 ;
  assign n538 = n527 | n537 ;
  assign n539 = n159 & n469 ;
  assign n540 = n159 & n236 ;
  assign n541 = n237 | n540 ;
  assign n542 = n539 | n541 ;
  assign n543 = n538 | n542 ;
  assign n544 = n342 & ~n543 ;
  assign n545 = n174 | n380 ;
  assign n546 = n93 | n545 ;
  assign n547 = n205 | n381 ;
  assign n548 = n546 | n547 ;
  assign n549 = n76 | n110 ;
  assign n550 = n155 | n549 ;
  assign n551 = n173 | n550 ;
  assign n552 = n548 | n551 ;
  assign n553 = n362 | n366 ;
  assign n554 = n46 | n553 ;
  assign n555 = n77 | n437 ;
  assign n556 = n436 | n555 ;
  assign n557 = n390 | n393 ;
  assign n558 = n120 | n557 ;
  assign n559 = n556 | n558 ;
  assign n560 = n102 | n160 ;
  assign n561 = ( n175 & n186 ) | ( n175 & ~n560 ) | ( n186 & ~n560 ) ;
  assign n562 = n560 | n561 ;
  assign n563 = n559 | n562 ;
  assign n564 = n443 | n563 ;
  assign n565 = n187 | n444 ;
  assign n566 = n154 | n565 ;
  assign n567 = n564 | n566 ;
  assign n568 = n122 | n457 ;
  assign n569 = n138 & n392 ;
  assign n570 = n91 & n392 ;
  assign n571 = n569 | n570 ;
  assign n572 = n568 | n571 ;
  assign n573 = n408 | n572 ;
  assign n574 = n567 | n573 ;
  assign n575 = n554 | n574 ;
  assign n576 = n552 | n575 ;
  assign n577 = n544 & ~n576 ;
  assign n578 = n49 & n392 ;
  assign n579 = n109 & n392 ;
  assign n580 = n89 & n392 ;
  assign n581 = n579 | n580 ;
  assign n582 = n72 & n392 ;
  assign n583 = n42 & n392 ;
  assign n584 = n582 | n583 ;
  assign n585 = n581 | n584 ;
  assign n586 = n578 | n585 ;
  assign n587 = n166 | n586 ;
  assign n588 = n364 | n587 ;
  assign n589 = n577 & ~n588 ;
  assign n590 = ~n45 & n91 ;
  assign n591 = n159 & n392 ;
  assign n592 = n61 & n392 ;
  assign n593 = n591 | n592 ;
  assign n594 = n590 | n593 ;
  assign n595 = ~n45 & n138 ;
  assign n596 = n56 & n392 ;
  assign n597 = ~n113 & n392 ;
  assign n598 = n596 | n597 ;
  assign n599 = n595 | n598 ;
  assign n600 = n594 | n599 ;
  assign n601 = ~n45 & n54 ;
  assign n602 = ~n45 & n72 ;
  assign n603 = n601 | n602 ;
  assign n604 = n205 | n603 ;
  assign n605 = n59 | n604 ;
  assign n606 = n600 | n605 ;
  assign n607 = n64 & n392 ;
  assign n608 = ~n45 & n78 ;
  assign n609 = n607 | n608 ;
  assign n610 = ~n45 & n84 ;
  assign n611 = n222 | n610 ;
  assign n612 = n216 | n611 ;
  assign n613 = n609 | n612 ;
  assign n614 = n606 | n613 ;
  assign n615 = ~n46 & n226 ;
  assign n616 = ~n614 & n615 ;
  assign n617 = ~n43 & n235 ;
  assign n618 = n91 & n617 ;
  assign n619 = n78 & n617 ;
  assign n620 = n618 | n619 ;
  assign n621 = n159 & n617 ;
  assign n622 = n42 & n617 ;
  assign n623 = n621 | n622 ;
  assign n624 = n620 | n623 ;
  assign n625 = n64 & n617 ;
  assign n626 = n61 & n617 ;
  assign n627 = n625 | n626 ;
  assign n628 = n109 & n617 ;
  assign n629 = n84 & n617 ;
  assign n630 = n628 | n629 ;
  assign n631 = n627 | n630 ;
  assign n632 = n624 | n631 ;
  assign n633 = n138 & n617 ;
  assign n634 = n49 & n617 ;
  assign n635 = n633 | n634 ;
  assign n636 = n89 & n617 ;
  assign n637 = n56 & n617 ;
  assign n638 = n636 | n637 ;
  assign n639 = n54 & n617 ;
  assign n640 = n78 & n156 ;
  assign n641 = n639 | n640 ;
  assign n642 = n638 | n641 ;
  assign n643 = n635 | n642 ;
  assign n644 = n632 | n643 ;
  assign n645 = n91 & n156 ;
  assign n646 = n84 & n156 ;
  assign n647 = n138 & n156 ;
  assign n648 = n646 | n647 ;
  assign n649 = n72 & n156 ;
  assign n650 = n54 & n156 ;
  assign n651 = n649 | n650 ;
  assign n652 = n648 | n651 ;
  assign n653 = ~n113 & n617 ;
  assign n654 = n72 & n617 ;
  assign n655 = n95 & n617 ;
  assign n656 = n654 | n655 ;
  assign n657 = n653 | n656 ;
  assign n658 = n652 | n657 ;
  assign n659 = n645 | n658 ;
  assign n660 = n644 | n659 ;
  assign n661 = n49 & n156 ;
  assign n662 = n210 | n661 ;
  assign n663 = n225 | n662 ;
  assign n664 = n219 | n663 ;
  assign n665 = n660 | n664 ;
  assign n666 = n227 | n665 ;
  assign n667 = n616 & ~n666 ;
  assign n668 = ~n189 & n667 ;
  assign n669 = ~n113 & n469 ;
  assign n670 = n95 & n392 ;
  assign n671 = n669 | n670 ;
  assign n672 = n668 & ~n671 ;
  assign n673 = n589 | n672 ;
  assign n674 = n589 & n672 ;
  assign n675 = n673 & ~n674 ;
  assign n676 = n250 | n350 ;
  assign n677 = n451 | n676 ;
  assign n678 = n403 | n470 ;
  assign n679 = n242 | n678 ;
  assign n680 = n677 | n679 ;
  assign n681 = n521 | n569 ;
  assign n682 = n190 | n681 ;
  assign n683 = n125 | n682 ;
  assign n684 = n680 | n683 ;
  assign n685 = n96 | n438 ;
  assign n686 = n684 | n685 ;
  assign n687 = n93 | n277 ;
  assign n688 = n197 | n416 ;
  assign n689 = n687 | n688 ;
  assign n690 = n531 | n540 ;
  assign n691 = n609 | n690 ;
  assign n692 = n504 | n647 ;
  assign n693 = n691 | n692 ;
  assign n694 = n689 | n693 ;
  assign n695 = n568 | n694 ;
  assign n696 = n686 | n695 ;
  assign n697 = n299 | n337 ;
  assign n698 = n625 | n697 ;
  assign n699 = n539 | n698 ;
  assign n700 = n498 | n699 ;
  assign n701 = n314 | n700 ;
  assign n702 = n295 | n701 ;
  assign n703 = n696 | n702 ;
  assign n704 = n198 | n307 ;
  assign n705 = n452 | n704 ;
  assign n706 = n590 | n705 ;
  assign n707 = n703 | n706 ;
  assign n708 = n160 | n193 ;
  assign n709 = n645 | n708 ;
  assign n710 = n274 | n296 ;
  assign n711 = n417 | n476 ;
  assign n712 = n710 | n711 ;
  assign n713 = n709 | n712 ;
  assign n714 = n315 | n489 ;
  assign n715 = n327 | n714 ;
  assign n716 = n292 | n715 ;
  assign n717 = n713 | n716 ;
  assign n718 = n503 | n529 ;
  assign n719 = n258 | n484 ;
  assign n720 = n718 | n719 ;
  assign n721 = n419 | n591 ;
  assign n722 = n582 | n721 ;
  assign n723 = n720 | n722 ;
  assign n724 = n602 | n723 ;
  assign n725 = n244 | n618 ;
  assign n726 = n52 | n520 ;
  assign n727 = n725 | n726 ;
  assign n728 = n522 | n634 ;
  assign n729 = n164 | n291 ;
  assign n730 = n728 | n729 ;
  assign n731 = n145 | n468 ;
  assign n732 = n134 | n650 ;
  assign n733 = n731 | n732 ;
  assign n734 = n132 | n482 ;
  assign n735 = n146 | n734 ;
  assign n736 = n733 | n735 ;
  assign n737 = n730 | n736 ;
  assign n738 = n727 | n737 ;
  assign n739 = n724 | n738 ;
  assign n740 = n398 | n739 ;
  assign n741 = n717 | n740 ;
  assign n742 = n707 | n741 ;
  assign n743 = n601 | n621 ;
  assign n744 = n181 | n458 ;
  assign n745 = n743 | n744 ;
  assign n746 = n187 | n745 ;
  assign n747 = n420 | n478 ;
  assign n748 = n151 | n747 ;
  assign n749 = n180 | n319 ;
  assign n750 = n748 | n749 ;
  assign n751 = n746 | n750 ;
  assign n752 = n213 | n580 ;
  assign n753 = n245 | n306 ;
  assign n754 = n752 | n753 ;
  assign n755 = n408 | n754 ;
  assign n756 = n528 | n579 ;
  assign n757 = n755 | n756 ;
  assign n758 = n751 | n757 ;
  assign n759 = n99 | n654 ;
  assign n760 = n270 | n293 ;
  assign n761 = n759 | n760 ;
  assign n762 = n336 | n761 ;
  assign n763 = n633 | n762 ;
  assign n764 = n280 | n763 ;
  assign n765 = n758 | n764 ;
  assign n766 = n111 | n765 ;
  assign n767 = n475 | n766 ;
  assign n768 = n626 | n767 ;
  assign n769 = n742 | n768 ;
  assign n770 = n283 | n505 ;
  assign n771 = n266 | n770 ;
  assign n772 = n320 | n771 ;
  assign n773 = n62 | n772 ;
  assign n774 = n114 | n773 ;
  assign n775 = n186 | n774 ;
  assign n776 = n152 | n775 ;
  assign n777 = n157 | n776 ;
  assign n778 = n769 | n777 ;
  assign n779 = n146 | n383 ;
  assign n780 = n443 | n779 ;
  assign n781 = n260 | n499 ;
  assign n782 = n338 | n781 ;
  assign n783 = n780 | n782 ;
  assign n784 = n55 | n194 ;
  assign n785 = n445 | n784 ;
  assign n786 = n164 | n785 ;
  assign n787 = n783 | n786 ;
  assign n788 = n77 | n100 ;
  assign n789 = n787 | n788 ;
  assign n790 = n319 | n429 ;
  assign n791 = n301 | n510 ;
  assign n792 = n790 | n791 ;
  assign n793 = n130 | n634 ;
  assign n794 = n792 | n793 ;
  assign n795 = n384 | n654 ;
  assign n796 = n416 | n795 ;
  assign n797 = n76 | n796 ;
  assign n798 = n794 | n797 ;
  assign n799 = n168 | n295 ;
  assign n800 = n365 | n799 ;
  assign n801 = n258 | n404 ;
  assign n802 = n752 | n801 ;
  assign n803 = n800 | n802 ;
  assign n804 = n798 | n803 ;
  assign n805 = n789 | n804 ;
  assign n806 = n227 | n490 ;
  assign n807 = n438 | n592 ;
  assign n808 = n292 | n655 ;
  assign n809 = n807 | n808 ;
  assign n810 = n806 | n809 ;
  assign n811 = n472 | n810 ;
  assign n812 = n629 | n811 ;
  assign n813 = n334 | n812 ;
  assign n814 = n805 | n813 ;
  assign n815 = n263 | n457 ;
  assign n816 = n165 | n815 ;
  assign n817 = n273 | n578 ;
  assign n818 = n219 | n817 ;
  assign n819 = n678 | n818 ;
  assign n820 = n132 | n528 ;
  assign n821 = n269 | n522 ;
  assign n822 = n355 | n821 ;
  assign n823 = n820 | n822 ;
  assign n824 = n819 | n823 ;
  assign n825 = n816 | n824 ;
  assign n826 = n468 | n825 ;
  assign n827 = n204 | n826 ;
  assign n828 = n814 | n827 ;
  assign n829 = n244 | n337 ;
  assign n830 = n393 | n829 ;
  assign n831 = n270 | n345 ;
  assign n832 = n830 | n831 ;
  assign n833 = n310 | n645 ;
  assign n834 = n252 | n489 ;
  assign n835 = n83 | n478 ;
  assign n836 = n834 | n835 ;
  assign n837 = n833 | n836 ;
  assign n838 = n832 | n837 ;
  assign n839 = n266 | n621 ;
  assign n840 = n222 | n435 ;
  assign n841 = n839 | n840 ;
  assign n842 = n250 | n475 ;
  assign n843 = n108 | n327 ;
  assign n844 = n173 | n351 ;
  assign n845 = n843 | n844 ;
  assign n846 = n842 | n845 ;
  assign n847 = n841 | n846 ;
  assign n848 = n838 | n847 ;
  assign n849 = n207 | n514 ;
  assign n850 = n521 | n601 ;
  assign n851 = n849 | n850 ;
  assign n852 = n283 | n670 ;
  assign n853 = n444 | n852 ;
  assign n854 = n851 | n853 ;
  assign n855 = n81 | n111 ;
  assign n856 = n854 | n855 ;
  assign n857 = n349 | n539 ;
  assign n858 = n571 | n857 ;
  assign n859 = n856 | n858 ;
  assign n860 = n848 | n859 ;
  assign n861 = n193 | n590 ;
  assign n862 = n187 | n591 ;
  assign n863 = n861 | n862 ;
  assign n864 = n409 | n863 ;
  assign n865 = n417 | n864 ;
  assign n866 = n125 | n865 ;
  assign n867 = n860 | n866 ;
  assign n868 = n181 | n596 ;
  assign n869 = n359 | n583 ;
  assign n870 = n197 | n646 ;
  assign n871 = n869 | n870 ;
  assign n872 = n868 | n871 ;
  assign n873 = n140 | n313 ;
  assign n874 = n198 | n249 ;
  assign n875 = n103 | n874 ;
  assign n876 = n873 | n875 ;
  assign n877 = n872 | n876 ;
  assign n878 = n175 | n420 ;
  assign n879 = n276 | n391 ;
  assign n880 = n57 | n306 ;
  assign n881 = n879 | n880 ;
  assign n882 = n878 | n881 ;
  assign n883 = n877 | n882 ;
  assign n884 = n595 | n883 ;
  assign n885 = n867 | n884 ;
  assign n886 = n828 | n885 ;
  assign n887 = n379 | n531 ;
  assign n888 = n291 | n636 ;
  assign n889 = n452 | n582 ;
  assign n890 = n513 | n889 ;
  assign n891 = n110 | n112 ;
  assign n892 = n133 | n151 ;
  assign n893 = n511 | n579 ;
  assign n894 = n892 | n893 ;
  assign n895 = ( n215 & ~n891 ) | ( n215 & n894 ) | ( ~n891 & n894 ) ;
  assign n896 = n891 | n895 ;
  assign n897 = n890 | n896 ;
  assign n898 = n888 | n897 ;
  assign n899 = n641 | n898 ;
  assign n900 = n887 | n899 ;
  assign n901 = n280 | n900 ;
  assign n902 = n607 | n901 ;
  assign n903 = n886 | n902 ;
  assign n904 = n85 | n903 ;
  assign n905 = n778 & n904 ;
  assign n906 = n778 | n904 ;
  assign n907 = ~n905 & n906 ;
  assign n908 = n349 | n416 ;
  assign n909 = n224 | n377 ;
  assign n910 = n908 | n909 ;
  assign n911 = n500 | n590 ;
  assign n912 = n488 | n911 ;
  assign n913 = n910 | n912 ;
  assign n914 = n522 | n653 ;
  assign n915 = n241 | n914 ;
  assign n916 = n449 | n915 ;
  assign n917 = n913 | n916 ;
  assign n918 = n94 | n217 ;
  assign n919 = n157 | n918 ;
  assign n920 = n917 | n919 ;
  assign n921 = n381 | n531 ;
  assign n922 = n366 | n921 ;
  assign n923 = n165 | n408 ;
  assign n924 = n314 | n591 ;
  assign n925 = n923 | n924 ;
  assign n926 = n46 | n925 ;
  assign n927 = n199 | n441 ;
  assign n928 = n260 | n355 ;
  assign n929 = n927 | n928 ;
  assign n930 = n926 | n929 ;
  assign n931 = n922 | n930 ;
  assign n932 = n920 | n931 ;
  assign n933 = n175 | n626 ;
  assign n934 = n476 | n933 ;
  assign n935 = n509 | n934 ;
  assign n936 = n634 | n935 ;
  assign n937 = n510 | n936 ;
  assign n938 = n420 | n937 ;
  assign n939 = n932 | n938 ;
  assign n940 = n193 | n400 ;
  assign n941 = n191 | n940 ;
  assign n942 = n172 | n941 ;
  assign n943 = n143 | n942 ;
  assign n944 = n939 | n943 ;
  assign n945 = n134 | n237 ;
  assign n946 = n661 | n945 ;
  assign n947 = n306 | n475 ;
  assign n948 = n125 | n359 ;
  assign n949 = n947 | n948 ;
  assign n950 = n946 | n949 ;
  assign n951 = n624 | n950 ;
  assign n952 = n262 | n528 ;
  assign n953 = n399 | n952 ;
  assign n954 = n391 | n444 ;
  assign n955 = n953 | n954 ;
  assign n956 = n311 | n955 ;
  assign n957 = n951 | n956 ;
  assign n958 = n472 | n639 ;
  assign n959 = n296 | n499 ;
  assign n960 = n358 | n596 ;
  assign n961 = n807 | n960 ;
  assign n962 = n101 | n961 ;
  assign n963 = n959 | n962 ;
  assign n964 = n958 | n963 ;
  assign n965 = n957 | n964 ;
  assign n966 = n164 | n173 ;
  assign n967 = ( n128 & n315 ) | ( n128 & ~n966 ) | ( n315 & ~n966 ) ;
  assign n968 = n966 | n967 ;
  assign n969 = n152 | n968 ;
  assign n970 = n223 | n969 ;
  assign n971 = n965 | n970 ;
  assign n972 = n194 | n428 ;
  assign n973 = n326 | n404 ;
  assign n974 = n142 | n206 ;
  assign n975 = n973 | n974 ;
  assign n976 = n320 | n470 ;
  assign n977 = n356 | n976 ;
  assign n978 = n975 | n977 ;
  assign n979 = n57 | n435 ;
  assign n980 = n226 & ~n979 ;
  assign n981 = ~n112 & n980 ;
  assign n982 = ~n978 & n981 ;
  assign n983 = ~n161 & n982 ;
  assign n984 = n482 | n503 ;
  assign n985 = n251 | n984 ;
  assign n986 = n790 | n985 ;
  assign n987 = n103 | n282 ;
  assign n988 = n336 | n987 ;
  assign n989 = n986 | n988 ;
  assign n990 = n253 | n280 ;
  assign n991 = n611 | n990 ;
  assign n992 = n160 | n393 ;
  assign n993 = n132 | n992 ;
  assign n994 = n991 | n993 ;
  assign n995 = n174 | n498 ;
  assign n996 = n65 | n645 ;
  assign n997 = n995 | n996 ;
  assign n998 = n102 | n655 ;
  assign n999 = n997 | n998 ;
  assign n1000 = n994 | n999 ;
  assign n1001 = n989 | n1000 ;
  assign n1002 = n983 & ~n1001 ;
  assign n1003 = ~n972 & n1002 ;
  assign n1004 = ~n971 & n1003 ;
  assign n1005 = ~n944 & n1004 ;
  assign n1006 = n278 | n648 ;
  assign n1007 = n479 | n1006 ;
  assign n1008 = n258 | n1007 ;
  assign n1009 = n383 | n1008 ;
  assign n1010 = n419 | n1009 ;
  assign n1011 = n437 | n1010 ;
  assign n1012 = n90 | n1011 ;
  assign n1013 = n85 | n1012 ;
  assign n1014 = n1005 & ~n1013 ;
  assign n1015 = n904 & ~n1014 ;
  assign n1016 = n511 | n513 ;
  assign n1017 = n111 | n500 ;
  assign n1018 = n128 | n1017 ;
  assign n1019 = n242 | n637 ;
  assign n1020 = n94 | n1019 ;
  assign n1021 = n1018 | n1020 ;
  assign n1022 = n262 | n582 ;
  assign n1023 = n498 | n654 ;
  assign n1024 = n252 | n314 ;
  assign n1025 = n1023 | n1024 ;
  assign n1026 = n1022 | n1025 ;
  assign n1027 = n1021 | n1026 ;
  assign n1028 = n194 | n351 ;
  assign n1029 = n165 | n1028 ;
  assign n1030 = n640 | n1029 ;
  assign n1031 = n1027 | n1030 ;
  assign n1032 = n199 | n270 ;
  assign n1033 = n946 | n1032 ;
  assign n1034 = n335 | n570 ;
  assign n1035 = n169 | n1034 ;
  assign n1036 = n249 | n366 ;
  assign n1037 = n1035 | n1036 ;
  assign n1038 = n1033 | n1037 ;
  assign n1039 = n580 | n670 ;
  assign n1040 = n458 | n602 ;
  assign n1041 = n1039 | n1040 ;
  assign n1042 = n1038 | n1041 ;
  assign n1043 = n1031 | n1042 ;
  assign n1044 = n419 | n519 ;
  assign n1045 = n266 | n380 ;
  assign n1046 = n1044 | n1045 ;
  assign n1047 = n429 | n1046 ;
  assign n1048 = n653 | n1047 ;
  assign n1049 = ( ~n1016 & n1043 ) | ( ~n1016 & n1048 ) | ( n1043 & n1048 ) ;
  assign n1050 = n1016 | n1049 ;
  assign n1051 = n619 | n669 ;
  assign n1052 = n217 | n384 ;
  assign n1053 = n1051 | n1052 ;
  assign n1054 = n146 | n321 ;
  assign n1055 = n491 | n1054 ;
  assign n1056 = n1053 | n1055 ;
  assign n1057 = n191 | n540 ;
  assign n1058 = n292 | n1057 ;
  assign n1059 = n383 | n1058 ;
  assign n1060 = n1056 | n1059 ;
  assign n1061 = n226 & ~n346 ;
  assign n1062 = ~n133 & n1061 ;
  assign n1063 = ~n1060 & n1062 ;
  assign n1064 = n96 | n595 ;
  assign n1065 = n850 | n1064 ;
  assign n1066 = n164 | n245 ;
  assign n1067 = n710 | n1066 ;
  assign n1068 = n1065 | n1067 ;
  assign n1069 = n81 | n350 ;
  assign n1070 = n250 | n1069 ;
  assign n1071 = n291 | n1070 ;
  assign n1072 = n1068 | n1071 ;
  assign n1073 = n186 | n441 ;
  assign n1074 = n172 | n1073 ;
  assign n1075 = n227 | n1074 ;
  assign n1076 = n1072 | n1075 ;
  assign n1077 = n99 | n505 ;
  assign n1078 = n139 | n530 ;
  assign n1079 = n151 | n240 ;
  assign n1080 = n1078 | n1079 ;
  assign n1081 = n504 | n1080 ;
  assign n1082 = n468 | n514 ;
  assign n1083 = n313 | n1082 ;
  assign n1084 = n472 | n1083 ;
  assign n1085 = n636 | n1084 ;
  assign n1086 = n1081 | n1085 ;
  assign n1087 = n1077 | n1086 ;
  assign n1088 = n1076 | n1087 ;
  assign n1089 = n1063 & ~n1088 ;
  assign n1090 = ~n1050 & n1089 ;
  assign n1091 = ~n158 & n1090 ;
  assign n1092 = n161 | n451 ;
  assign n1093 = n122 | n1092 ;
  assign n1094 = n215 | n279 ;
  assign n1095 = n86 | n1094 ;
  assign n1096 = n1093 | n1095 ;
  assign n1097 = n428 | n655 ;
  assign n1098 = n320 | n1097 ;
  assign n1099 = n269 | n1098 ;
  assign n1100 = n1096 | n1099 ;
  assign n1101 = n222 | n450 ;
  assign n1102 = n132 | n1101 ;
  assign n1103 = n207 | n1102 ;
  assign n1104 = n1100 | n1103 ;
  assign n1105 = n528 | n578 ;
  assign n1106 = n418 | n1105 ;
  assign n1107 = n46 | n173 ;
  assign n1108 = n1106 | n1107 ;
  assign n1109 = n76 | n379 ;
  assign n1110 = n609 | n1109 ;
  assign n1111 = n114 | n1110 ;
  assign n1112 = n830 | n1111 ;
  assign n1113 = n1108 | n1112 ;
  assign n1114 = n1104 | n1113 ;
  assign n1115 = n198 | n263 ;
  assign n1116 = n299 | n478 ;
  assign n1117 = n344 | n1116 ;
  assign n1118 = n295 | n306 ;
  assign n1119 = n634 | n1118 ;
  assign n1120 = n1117 | n1119 ;
  assign n1121 = n307 | n596 ;
  assign n1122 = n58 | n1121 ;
  assign n1123 = n445 | n1122 ;
  assign n1124 = n1120 | n1123 ;
  assign n1125 = n103 | n1124 ;
  assign n1126 = n1115 | n1125 ;
  assign n1127 = n1114 | n1126 ;
  assign n1128 = n120 | n319 ;
  assign n1129 = n479 | n626 ;
  assign n1130 = n300 | n391 ;
  assign n1131 = n1129 | n1130 ;
  assign n1132 = n592 | n1131 ;
  assign n1133 = n127 | n1132 ;
  assign n1134 = n1128 | n1133 ;
  assign n1135 = n277 | n1134 ;
  assign n1136 = n355 | n1135 ;
  assign n1137 = n1127 | n1136 ;
  assign n1138 = n190 | n193 ;
  assign n1139 = n649 | n1138 ;
  assign n1140 = n1137 | n1139 ;
  assign n1141 = n1091 & ~n1140 ;
  assign n1142 = n539 | n621 ;
  assign n1143 = n338 | n1142 ;
  assign n1144 = n420 | n1143 ;
  assign n1145 = n579 | n1144 ;
  assign n1146 = n590 | n1145 ;
  assign n1147 = n377 | n1146 ;
  assign n1148 = n110 | n1147 ;
  assign n1149 = n152 | n1148 ;
  assign n1150 = n647 | n1149 ;
  assign n1151 = n1141 & ~n1150 ;
  assign n1152 = n99 | n186 ;
  assign n1153 = n111 | n125 ;
  assign n1154 = n498 | n510 ;
  assign n1155 = n627 | n1154 ;
  assign n1156 = ( n269 & ~n1153 ) | ( n269 & n1155 ) | ( ~n1153 & n1155 ) ;
  assign n1157 = n1153 | n1156 ;
  assign n1158 = n1152 | n1157 ;
  assign n1159 = n241 | n263 ;
  assign n1160 = n500 | n580 ;
  assign n1161 = n420 | n583 ;
  assign n1162 = n1160 | n1161 ;
  assign n1163 = n1159 | n1162 ;
  assign n1164 = n356 | n428 ;
  assign n1165 = n301 | n337 ;
  assign n1166 = n996 | n1165 ;
  assign n1167 = n1164 | n1166 ;
  assign n1168 = n1163 | n1167 ;
  assign n1169 = n1158 | n1168 ;
  assign n1170 = n381 | n637 ;
  assign n1171 = n1069 | n1170 ;
  assign n1172 = n473 | n1171 ;
  assign n1173 = n482 | n1172 ;
  assign n1174 = n314 | n1173 ;
  assign n1175 = n1169 | n1174 ;
  assign n1176 = n313 | n1175 ;
  assign n1177 = n175 | n610 ;
  assign n1178 = n490 | n636 ;
  assign n1179 = n1177 | n1178 ;
  assign n1180 = n279 | n522 ;
  assign n1181 = n326 | n1180 ;
  assign n1182 = n1179 | n1181 ;
  assign n1183 = n224 | n1182 ;
  assign n1184 = n245 | n622 ;
  assign n1185 = n161 | n582 ;
  assign n1186 = n1184 | n1185 ;
  assign n1187 = n128 | n1186 ;
  assign n1188 = n452 | n591 ;
  assign n1189 = n52 | n94 ;
  assign n1190 = n1188 | n1189 ;
  assign n1191 = n59 | n1190 ;
  assign n1192 = n1187 | n1191 ;
  assign n1193 = n1183 | n1192 ;
  assign n1194 = n133 | n227 ;
  assign n1195 = n1078 | n1194 ;
  assign n1196 = n409 | n1195 ;
  assign n1197 = n334 | n1196 ;
  assign n1198 = n276 | n1197 ;
  assign n1199 = n1193 | n1198 ;
  assign n1200 = n62 | n540 ;
  assign n1201 = n215 | n335 ;
  assign n1202 = n377 | n1201 ;
  assign n1203 = n198 | n511 ;
  assign n1204 = n265 | n628 ;
  assign n1205 = n1203 | n1204 ;
  assign n1206 = n1202 | n1205 ;
  assign n1207 = n1200 | n1206 ;
  assign n1208 = n309 | n602 ;
  assign n1209 = n403 | n1208 ;
  assign n1210 = n640 | n1209 ;
  assign n1211 = n1207 | n1210 ;
  assign n1212 = n1199 | n1211 ;
  assign n1213 = n1176 | n1212 ;
  assign n1214 = n197 | n315 ;
  assign n1215 = n844 | n1214 ;
  assign n1216 = n250 | n479 ;
  assign n1217 = n450 | n1216 ;
  assign n1218 = n1215 | n1217 ;
  assign n1219 = n151 | n1218 ;
  assign n1220 = n181 | n435 ;
  assign n1221 = n344 | n458 ;
  assign n1222 = n432 | n1221 ;
  assign n1223 = n1220 | n1222 ;
  assign n1224 = n857 | n1223 ;
  assign n1225 = n789 | n1224 ;
  assign n1226 = n1219 | n1225 ;
  assign n1227 = n887 | n1226 ;
  assign n1228 = n1213 | n1227 ;
  assign n1229 = n93 | n648 ;
  assign n1230 = n266 | n1229 ;
  assign n1231 = n419 | n1230 ;
  assign n1232 = n364 | n1231 ;
  assign n1233 = n1228 | n1232 ;
  assign n1234 = ~n1151 & n1233 ;
  assign n1235 = n1151 & ~n1233 ;
  assign n1236 = n1234 | n1235 ;
  assign n1237 = n592 | n633 ;
  assign n1238 = n445 | n1237 ;
  assign n1239 = n1131 | n1238 ;
  assign n1240 = n103 | n490 ;
  assign n1241 = n1239 | n1240 ;
  assign n1242 = n216 | n1085 ;
  assign n1243 = n1241 | n1242 ;
  assign n1244 = n241 | n419 ;
  assign n1245 = n579 | n1244 ;
  assign n1246 = n522 | n640 ;
  assign n1247 = n315 | n1246 ;
  assign n1248 = n1245 | n1247 ;
  assign n1249 = n252 | n334 ;
  assign n1250 = n145 | n1249 ;
  assign n1251 = n649 | n1250 ;
  assign n1252 = n1248 | n1251 ;
  assign n1253 = n349 | n482 ;
  assign n1254 = n152 | n578 ;
  assign n1255 = n141 | n1254 ;
  assign n1256 = n1253 | n1255 ;
  assign n1257 = n1252 | n1256 ;
  assign n1258 = n1243 | n1257 ;
  assign n1259 = n263 | n862 ;
  assign n1260 = n186 | n670 ;
  assign n1261 = n218 | n258 ;
  assign n1262 = n1260 | n1261 ;
  assign n1263 = n432 | n1262 ;
  assign n1264 = n1259 | n1263 ;
  assign n1265 = n381 | n1264 ;
  assign n1266 = n293 | n1265 ;
  assign n1267 = n1258 | n1266 ;
  assign n1268 = ( n366 & n435 ) | ( n366 & ~n974 ) | ( n435 & ~n974 ) ;
  assign n1269 = n974 | n1268 ;
  assign n1270 = n1267 | n1269 ;
  assign n1271 = n355 | n409 ;
  assign n1272 = n274 | n476 ;
  assign n1273 = n1271 | n1272 ;
  assign n1274 = n197 | n499 ;
  assign n1275 = n143 | n1274 ;
  assign n1276 = n1273 | n1275 ;
  assign n1277 = n208 | n1276 ;
  assign n1278 = n270 | n618 ;
  assign n1279 = n650 | n1278 ;
  assign n1280 = n108 | n434 ;
  assign n1281 = n611 | n1280 ;
  assign n1282 = n1279 | n1281 ;
  assign n1283 = n590 | n1282 ;
  assign n1284 = n151 | n597 ;
  assign n1285 = n282 | n622 ;
  assign n1286 = n1284 | n1285 ;
  assign n1287 = n111 | n1286 ;
  assign n1288 = n83 | n647 ;
  assign n1289 = n799 | n1288 ;
  assign n1290 = n1287 | n1289 ;
  assign n1291 = n1283 | n1290 ;
  assign n1292 = n364 | n531 ;
  assign n1293 = n408 | n645 ;
  assign n1294 = n1292 | n1293 ;
  assign n1295 = n677 | n1294 ;
  assign n1296 = n428 | n510 ;
  assign n1297 = n157 | n1296 ;
  assign n1298 = n639 | n1297 ;
  assign n1299 = n1295 | n1298 ;
  assign n1300 = n504 | n669 ;
  assign n1301 = n262 | n1300 ;
  assign n1302 = n276 | n1301 ;
  assign n1303 = n345 | n1302 ;
  assign n1304 = n1299 | n1303 ;
  assign n1305 = n126 | n198 ;
  assign n1306 = n1304 | n1305 ;
  assign n1307 = n1291 | n1306 ;
  assign n1308 = n1277 | n1307 ;
  assign n1309 = n1270 | n1308 ;
  assign n1310 = n194 | n629 ;
  assign n1311 = n307 | n602 ;
  assign n1312 = n299 | n511 ;
  assign n1313 = n114 | n384 ;
  assign n1314 = n1312 | n1313 ;
  assign n1315 = n452 | n621 ;
  assign n1316 = n77 | n475 ;
  assign n1317 = n1315 | n1316 ;
  assign n1318 = n1314 | n1317 ;
  assign n1319 = n1311 | n1318 ;
  assign n1320 = n1310 | n1319 ;
  assign n1321 = n528 | n1320 ;
  assign n1322 = n634 | n1321 ;
  assign n1323 = n301 | n1322 ;
  assign n1324 = n344 | n1323 ;
  assign n1325 = n1309 | n1324 ;
  assign n1326 = n122 | n580 ;
  assign n1327 = n1325 | n1326 ;
  assign n1328 = ~n1151 & n1327 ;
  assign n1329 = n76 | n475 ;
  assign n1330 = n1284 | n1329 ;
  assign n1331 = n531 | n1188 ;
  assign n1332 = n1330 | n1331 ;
  assign n1333 = n1108 | n1332 ;
  assign n1334 = n115 | n1333 ;
  assign n1335 = n1063 & ~n1334 ;
  assign n1336 = n218 | n628 ;
  assign n1337 = n327 | n334 ;
  assign n1338 = n1336 | n1337 ;
  assign n1339 = n476 | n1338 ;
  assign n1340 = n479 | n1339 ;
  assign n1341 = n529 | n1340 ;
  assign n1342 = n633 | n1341 ;
  assign n1343 = n1335 & ~n1342 ;
  assign n1344 = n293 | n629 ;
  assign n1345 = n451 | n1344 ;
  assign n1346 = n125 | n1345 ;
  assign n1347 = n215 | n1346 ;
  assign n1348 = n442 | n1347 ;
  assign n1349 = n224 | n1348 ;
  assign n1350 = n1343 & ~n1349 ;
  assign n1351 = n65 | n513 ;
  assign n1352 = n197 | n326 ;
  assign n1353 = n167 | n1352 ;
  assign n1354 = n103 | n661 ;
  assign n1355 = n253 | n438 ;
  assign n1356 = n1354 | n1355 ;
  assign n1357 = n1353 | n1356 ;
  assign n1358 = n249 | n509 ;
  assign n1359 = n128 | n379 ;
  assign n1360 = n1358 | n1359 ;
  assign n1361 = n338 | n522 ;
  assign n1362 = n52 | n450 ;
  assign n1363 = n1361 | n1362 ;
  assign n1364 = n1360 | n1363 ;
  assign n1365 = n1357 | n1364 ;
  assign n1366 = n1351 | n1365 ;
  assign n1367 = n539 | n653 ;
  assign n1368 = n258 | n1367 ;
  assign n1369 = n1283 | n1368 ;
  assign n1370 = n1366 | n1369 ;
  assign n1371 = n142 | n180 ;
  assign n1372 = n206 | n478 ;
  assign n1373 = n1078 | n1372 ;
  assign n1374 = n1371 | n1373 ;
  assign n1375 = n241 | n1374 ;
  assign n1376 = n300 | n1375 ;
  assign n1377 = n393 | n569 ;
  assign n1378 = n126 | n449 ;
  assign n1379 = n1377 | n1378 ;
  assign n1380 = n279 | n602 ;
  assign n1381 = n646 | n1380 ;
  assign n1382 = n277 | n596 ;
  assign n1383 = n165 | n1382 ;
  assign n1384 = n1381 | n1383 ;
  assign n1385 = n1379 | n1384 ;
  assign n1386 = n337 | n511 ;
  assign n1387 = n301 | n356 ;
  assign n1388 = n1386 | n1387 ;
  assign n1389 = n364 | n435 ;
  assign n1390 = n1388 | n1389 ;
  assign n1391 = n1385 | n1390 ;
  assign n1392 = n1376 | n1391 ;
  assign n1393 = n1370 | n1392 ;
  assign n1394 = n100 | n309 ;
  assign n1395 = n208 | n1394 ;
  assign n1396 = n349 | n565 ;
  assign n1397 = n1395 | n1396 ;
  assign n1398 = n351 | n437 ;
  assign n1399 = n143 | n1398 ;
  assign n1400 = n1397 | n1399 ;
  assign n1401 = n1076 | n1400 ;
  assign n1402 = n1393 | n1401 ;
  assign n1403 = n1350 & ~n1402 ;
  assign n1404 = n583 | n625 ;
  assign n1405 = n933 | n1404 ;
  assign n1406 = n237 | n1405 ;
  assign n1407 = n344 | n1406 ;
  assign n1408 = n55 | n1407 ;
  assign n1409 = n90 | n1408 ;
  assign n1410 = n168 | n1409 ;
  assign n1411 = n1403 & ~n1410 ;
  assign n1412 = n365 | n1018 ;
  assign n1413 = n641 | n1093 ;
  assign n1414 = n1412 | n1413 ;
  assign n1415 = n380 | n670 ;
  assign n1416 = n157 | n212 ;
  assign n1417 = n85 | n134 ;
  assign n1418 = ( ~n1415 & n1416 ) | ( ~n1415 & n1417 ) | ( n1416 & n1417 ) ;
  assign n1419 = n1415 | n1418 ;
  assign n1420 = n1414 | n1419 ;
  assign n1421 = n58 | n204 ;
  assign n1422 = n1420 | n1421 ;
  assign n1423 = n126 | n607 ;
  assign n1424 = n711 | n1423 ;
  assign n1425 = n52 | n1424 ;
  assign n1426 = n213 | n444 ;
  assign n1427 = n972 | n1426 ;
  assign n1428 = n186 | n403 ;
  assign n1429 = n1427 | n1428 ;
  assign n1430 = n266 | n337 ;
  assign n1431 = n472 | n482 ;
  assign n1432 = n101 | n1431 ;
  assign n1433 = n1430 | n1432 ;
  assign n1434 = n199 | n520 ;
  assign n1435 = n293 | n628 ;
  assign n1436 = n806 | n1435 ;
  assign n1437 = n1434 | n1436 ;
  assign n1438 = n1433 | n1437 ;
  assign n1439 = n1429 | n1438 ;
  assign n1440 = n1425 | n1439 ;
  assign n1441 = n1422 | n1440 ;
  assign n1442 = n400 | n478 ;
  assign n1443 = n57 | n654 ;
  assign n1444 = n1279 | n1443 ;
  assign n1445 = n284 | n1444 ;
  assign n1446 = n1442 | n1445 ;
  assign n1447 = n431 | n1446 ;
  assign n1448 = n522 | n1447 ;
  assign n1449 = n1441 | n1448 ;
  assign n1450 = n306 | n504 ;
  assign n1451 = n358 | n1450 ;
  assign n1452 = n434 | n1451 ;
  assign n1453 = n187 | n1452 ;
  assign n1454 = n1449 | n1453 ;
  assign n1455 = n252 | n498 ;
  assign n1456 = n320 | n344 ;
  assign n1457 = n1455 | n1456 ;
  assign n1458 = n321 | n648 ;
  assign n1459 = n1457 | n1458 ;
  assign n1460 = n65 | n579 ;
  assign n1461 = n172 | n1460 ;
  assign n1462 = n1459 | n1461 ;
  assign n1463 = n314 | n499 ;
  assign n1464 = n76 | n731 ;
  assign n1465 = n90 | n338 ;
  assign n1466 = n96 | n1465 ;
  assign n1467 = n1464 | n1466 ;
  assign n1468 = n1463 | n1467 ;
  assign n1469 = n237 | n591 ;
  assign n1470 = n164 | n457 ;
  assign n1471 = n1469 | n1470 ;
  assign n1472 = n175 | n206 ;
  assign n1473 = n1471 | n1472 ;
  assign n1474 = n1468 | n1473 ;
  assign n1475 = n291 | n450 ;
  assign n1476 = n155 | n1475 ;
  assign n1477 = n409 | n1352 ;
  assign n1478 = n1476 | n1477 ;
  assign n1479 = n265 | n307 ;
  assign n1480 = n580 | n1479 ;
  assign n1481 = n193 | n1480 ;
  assign n1482 = n1478 | n1481 ;
  assign n1483 = n114 | n217 ;
  assign n1484 = n1482 | n1483 ;
  assign n1485 = n1474 | n1484 ;
  assign n1486 = n292 | n381 ;
  assign n1487 = n435 | n1486 ;
  assign n1488 = n62 | n345 ;
  assign n1489 = n222 | n1488 ;
  assign n1490 = n484 | n1489 ;
  assign n1491 = n1487 | n1490 ;
  assign n1492 = n661 | n1491 ;
  assign n1493 = n1115 | n1492 ;
  assign n1494 = n528 | n1493 ;
  assign n1495 = n1485 | n1494 ;
  assign n1496 = n420 | n458 ;
  assign n1497 = n404 | n1496 ;
  assign n1498 = n779 | n1094 ;
  assign n1499 = n1497 | n1498 ;
  assign n1500 = n429 | n540 ;
  assign n1501 = n276 | n1500 ;
  assign n1502 = n55 | n1501 ;
  assign n1503 = n1499 | n1502 ;
  assign n1504 = n108 | n608 ;
  assign n1505 = n139 | n1504 ;
  assign n1506 = n218 | n1505 ;
  assign n1507 = n645 | n1506 ;
  assign n1508 = n1503 | n1507 ;
  assign n1509 = n510 | n622 ;
  assign n1510 = n503 | n1509 ;
  assign n1511 = n310 | n1510 ;
  assign n1512 = n319 | n1511 ;
  assign n1513 = n240 | n633 ;
  assign n1514 = n302 | n1513 ;
  assign n1515 = n1037 | n1514 ;
  assign n1516 = n1512 | n1515 ;
  assign n1517 = n1508 | n1516 ;
  assign n1518 = n515 | n1517 ;
  assign n1519 = n1495 | n1518 ;
  assign n1520 = n1462 | n1519 ;
  assign n1521 = n1454 | n1520 ;
  assign n1522 = n483 | n629 ;
  assign n1523 = n1284 | n1522 ;
  assign n1524 = n531 | n1523 ;
  assign n1525 = n669 | n1524 ;
  assign n1526 = n350 | n1525 ;
  assign n1527 = n241 | n1526 ;
  assign n1528 = n602 | n1527 ;
  assign n1529 = n377 | n1528 ;
  assign n1530 = n102 | n1529 ;
  assign n1531 = n165 | n1530 ;
  assign n1532 = n1521 | n1531 ;
  assign n1533 = ~n1411 & n1532 ;
  assign n1534 = n1411 & ~n1532 ;
  assign n1535 = n1533 | n1534 ;
  assign n1536 = n158 | n610 ;
  assign n1537 = n555 | n1404 ;
  assign n1538 = n1536 | n1537 ;
  assign n1539 = n1279 | n1315 ;
  assign n1540 = n1538 | n1539 ;
  assign n1541 = n253 | n472 ;
  assign n1542 = n186 | n1541 ;
  assign n1543 = n1540 | n1542 ;
  assign n1544 = n173 | n509 ;
  assign n1545 = n62 | n649 ;
  assign n1546 = n1544 | n1545 ;
  assign n1547 = n134 | n400 ;
  assign n1548 = n92 | n1547 ;
  assign n1549 = n1546 | n1548 ;
  assign n1550 = n878 | n1549 ;
  assign n1551 = n225 | n1550 ;
  assign n1552 = n1543 | n1551 ;
  assign n1553 = n861 | n1079 ;
  assign n1554 = n1115 | n1553 ;
  assign n1555 = n697 | n1554 ;
  assign n1556 = n511 | n1555 ;
  assign n1557 = n500 | n1556 ;
  assign n1558 = n1552 | n1557 ;
  assign n1559 = n358 | n470 ;
  assign n1560 = n1558 | n1559 ;
  assign n1561 = n112 | n580 ;
  assign n1562 = n349 | n431 ;
  assign n1563 = n1561 | n1562 ;
  assign n1564 = n241 | n597 ;
  assign n1565 = n1563 | n1564 ;
  assign n1566 = n55 | n529 ;
  assign n1567 = n94 | n1566 ;
  assign n1568 = n628 | n637 ;
  assign n1569 = n217 | n444 ;
  assign n1570 = n1568 | n1569 ;
  assign n1571 = n227 | n1570 ;
  assign n1572 = n1567 | n1571 ;
  assign n1573 = n1565 | n1572 ;
  assign n1574 = n96 | n633 ;
  assign n1575 = n505 | n540 ;
  assign n1576 = n373 | n442 ;
  assign n1577 = n1575 | n1576 ;
  assign n1578 = n129 | n326 ;
  assign n1579 = n301 | n1578 ;
  assign n1580 = n1577 | n1579 ;
  assign n1581 = n356 | n579 ;
  assign n1582 = n570 | n1581 ;
  assign n1583 = n1580 | n1582 ;
  assign n1584 = n1574 | n1583 ;
  assign n1585 = n1573 | n1584 ;
  assign n1586 = n476 | n514 ;
  assign n1587 = n276 | n1586 ;
  assign n1588 = n359 | n1587 ;
  assign n1589 = n346 | n1588 ;
  assign n1590 = n212 | n1589 ;
  assign n1591 = n377 | n1590 ;
  assign n1592 = n1585 | n1591 ;
  assign n1593 = n265 | n490 ;
  assign n1594 = n110 | n404 ;
  assign n1595 = n1593 | n1594 ;
  assign n1596 = n351 | n384 ;
  assign n1597 = n313 | n435 ;
  assign n1598 = n641 | n1597 ;
  assign n1599 = n1596 | n1598 ;
  assign n1600 = n1595 | n1599 ;
  assign n1601 = n65 | n484 ;
  assign n1602 = n381 | n619 ;
  assign n1603 = n1601 | n1602 ;
  assign n1604 = n126 | n344 ;
  assign n1605 = n1603 | n1604 ;
  assign n1606 = n1600 | n1605 ;
  assign n1607 = n111 | n152 ;
  assign n1608 = ( n74 & n172 ) | ( n74 & n1607 ) | ( n172 & n1607 ) ;
  assign n1609 = n1606 | n1608 ;
  assign n1610 = n842 | n1609 ;
  assign n1611 = n1592 | n1610 ;
  assign n1612 = n1560 | n1611 ;
  assign n1613 = n403 | n669 ;
  assign n1614 = n1311 | n1613 ;
  assign n1615 = n1104 | n1614 ;
  assign n1616 = n284 | n1615 ;
  assign n1617 = n759 | n1616 ;
  assign n1618 = n779 | n1617 ;
  assign n1619 = n1612 | n1618 ;
  assign n1620 = n539 | n721 ;
  assign n1621 = n596 | n1620 ;
  assign n1622 = n58 | n1621 ;
  assign n1623 = n160 | n1622 ;
  assign n1624 = n133 | n1623 ;
  assign n1625 = n1619 | n1624 ;
  assign n1626 = n242 | n504 ;
  assign n1627 = n55 | n345 ;
  assign n1628 = n1626 | n1627 ;
  assign n1629 = n445 | n1628 ;
  assign n1630 = n212 | n299 ;
  assign n1631 = n207 | n1630 ;
  assign n1632 = n338 | n479 ;
  assign n1633 = n83 | n269 ;
  assign n1634 = n1632 | n1633 ;
  assign n1635 = n1631 | n1634 ;
  assign n1636 = n237 | n649 ;
  assign n1637 = n1052 | n1636 ;
  assign n1638 = n1635 | n1637 ;
  assign n1639 = n1629 | n1638 ;
  assign n1640 = n717 | n1639 ;
  assign n1641 = n206 | n1073 ;
  assign n1642 = n1083 | n1641 ;
  assign n1643 = n490 | n591 ;
  assign n1644 = n57 | n1643 ;
  assign n1645 = n1280 | n1644 ;
  assign n1646 = n1642 | n1645 ;
  assign n1647 = n359 | n391 ;
  assign n1648 = n529 | n1647 ;
  assign n1649 = n592 | n1648 ;
  assign n1650 = n578 | n1649 ;
  assign n1651 = n1646 | n1650 ;
  assign n1652 = n102 | n364 ;
  assign n1653 = n650 | n1652 ;
  assign n1654 = n1651 | n1653 ;
  assign n1655 = n1640 | n1654 ;
  assign n1656 = n377 | n608 ;
  assign n1657 = n199 | n215 ;
  assign n1658 = n1463 | n1657 ;
  assign n1659 = n223 | n390 ;
  assign n1660 = n521 | n1659 ;
  assign n1661 = n358 | n1660 ;
  assign n1662 = n226 & ~n1661 ;
  assign n1663 = ~n100 & n1662 ;
  assign n1664 = ~n1658 & n1663 ;
  assign n1665 = ~n1656 & n1664 ;
  assign n1666 = ~n1655 & n1665 ;
  assign n1667 = n625 | n655 ;
  assign n1668 = n307 | n1667 ;
  assign n1669 = n355 | n1668 ;
  assign n1670 = n416 | n1669 ;
  assign n1671 = n595 | n1670 ;
  assign n1672 = n122 | n1671 ;
  assign n1673 = n1666 & ~n1672 ;
  assign n1674 = n90 | n610 ;
  assign n1675 = n161 | n1674 ;
  assign n1676 = n1497 | n1675 ;
  assign n1677 = n431 | n530 ;
  assign n1678 = n634 | n1677 ;
  assign n1679 = n1676 | n1678 ;
  assign n1680 = n194 | n241 ;
  assign n1681 = n142 | n260 ;
  assign n1682 = n151 | n380 ;
  assign n1683 = n1681 | n1682 ;
  assign n1684 = n1680 | n1683 ;
  assign n1685 = n258 | n320 ;
  assign n1686 = n110 | n570 ;
  assign n1687 = n1685 | n1686 ;
  assign n1688 = n126 | n379 ;
  assign n1689 = n1575 | n1688 ;
  assign n1690 = n1687 | n1689 ;
  assign n1691 = n1684 | n1690 ;
  assign n1692 = n488 | n636 ;
  assign n1693 = n438 | n483 ;
  assign n1694 = n1692 | n1693 ;
  assign n1695 = n227 | n1694 ;
  assign n1696 = n128 | n132 ;
  assign n1697 = n531 | n582 ;
  assign n1698 = n1696 | n1697 ;
  assign n1699 = n152 | n400 ;
  assign n1700 = n1698 | n1699 ;
  assign n1701 = n1695 | n1700 ;
  assign n1702 = n1691 | n1701 ;
  assign n1703 = n352 | n1128 ;
  assign n1704 = n409 | n1703 ;
  assign n1705 = n522 | n1704 ;
  assign n1706 = n470 | n1705 ;
  assign n1707 = n1702 | n1706 ;
  assign n1708 = n244 | n270 ;
  assign n1709 = n452 | n601 ;
  assign n1710 = n1708 | n1709 ;
  assign n1711 = n94 | n224 ;
  assign n1712 = n1710 | n1711 ;
  assign n1713 = n478 | n629 ;
  assign n1714 = n66 | n1713 ;
  assign n1715 = n620 | n1203 ;
  assign n1716 = n1714 | n1715 ;
  assign n1717 = n1712 | n1716 ;
  assign n1718 = n250 | n283 ;
  assign n1719 = n58 | n1718 ;
  assign n1720 = n1717 | n1719 ;
  assign n1721 = n1054 | n1720 ;
  assign n1722 = n1707 | n1721 ;
  assign n1723 = n1679 | n1722 ;
  assign n1724 = n1336 | n1723 ;
  assign n1725 = n1673 & ~n1724 ;
  assign n1726 = n626 | n648 ;
  assign n1727 = n301 | n1726 ;
  assign n1728 = n393 | n1727 ;
  assign n1729 = n134 | n1728 ;
  assign n1730 = n125 | n1729 ;
  assign n1731 = n143 | n1730 ;
  assign n1732 = n208 | n1731 ;
  assign n1733 = n1725 & ~n1732 ;
  assign n1734 = n1625 & ~n1733 ;
  assign n1735 = ~n1625 & n1733 ;
  assign n1736 = n1734 | n1735 ;
  assign n1737 = n245 | n505 ;
  assign n1738 = n473 | n1737 ;
  assign n1739 = n295 | n1738 ;
  assign n1740 = n122 | n519 ;
  assign n1741 = n129 | n1740 ;
  assign n1742 = n1631 | n1741 ;
  assign n1743 = n1739 | n1742 ;
  assign n1744 = n1512 | n1743 ;
  assign n1745 = n1400 | n1744 ;
  assign n1746 = n1495 | n1745 ;
  assign n1747 = n540 | n629 ;
  assign n1748 = n270 | n379 ;
  assign n1749 = n1747 | n1748 ;
  assign n1750 = n223 | n1749 ;
  assign n1751 = n337 | n404 ;
  assign n1752 = n296 | n321 ;
  assign n1753 = n458 | n1752 ;
  assign n1754 = n1751 | n1753 ;
  assign n1755 = n1750 | n1754 ;
  assign n1756 = n94 | n301 ;
  assign n1757 = n373 | n490 ;
  assign n1758 = n1756 | n1757 ;
  assign n1759 = n327 | n434 ;
  assign n1760 = n408 | n1759 ;
  assign n1761 = n1758 | n1760 ;
  assign n1762 = n111 | n112 ;
  assign n1763 = n167 | n1762 ;
  assign n1764 = n1761 | n1763 ;
  assign n1765 = n1755 | n1764 ;
  assign n1766 = n890 | n972 ;
  assign n1767 = n995 | n1766 ;
  assign n1768 = n418 | n1767 ;
  assign n1769 = n1765 | n1768 ;
  assign n1770 = n522 | n530 ;
  assign n1771 = n346 | n1770 ;
  assign n1772 = n590 | n1771 ;
  assign n1773 = n602 | n1772 ;
  assign n1774 = n126 | n1773 ;
  assign n1775 = n1769 | n1774 ;
  assign n1776 = n842 | n1775 ;
  assign n1777 = n1746 | n1776 ;
  assign n1778 = n190 | n610 ;
  assign n1779 = n273 | n655 ;
  assign n1780 = n1778 | n1779 ;
  assign n1781 = n482 | n1442 ;
  assign n1782 = n1780 | n1781 ;
  assign n1783 = n46 | n110 ;
  assign n1784 = n1782 | n1783 ;
  assign n1785 = n262 | n619 ;
  assign n1786 = n293 | n595 ;
  assign n1787 = n1785 | n1786 ;
  assign n1788 = n57 | n384 ;
  assign n1789 = n140 | n1788 ;
  assign n1790 = n1787 | n1789 ;
  assign n1791 = n181 | n618 ;
  assign n1792 = n358 | n479 ;
  assign n1793 = n92 | n203 ;
  assign n1794 = n1792 | n1793 ;
  assign n1795 = n1791 | n1794 ;
  assign n1796 = n1790 | n1795 ;
  assign n1797 = n1784 | n1796 ;
  assign n1798 = n520 | n1797 ;
  assign n1799 = n315 | n1798 ;
  assign n1800 = n334 | n1799 ;
  assign n1801 = n355 | n1800 ;
  assign n1802 = n1777 | n1801 ;
  assign n1803 = n173 | n1802 ;
  assign n1804 = n284 | n834 ;
  assign n1805 = n132 | n1804 ;
  assign n1806 = n249 | n706 ;
  assign n1807 = n441 | n1806 ;
  assign n1808 = n1805 | n1807 ;
  assign n1809 = n1177 | n1808 ;
  assign n1810 = n703 | n1809 ;
  assign n1811 = n269 | n519 ;
  assign n1812 = n158 | n1811 ;
  assign n1813 = n748 | n1812 ;
  assign n1814 = n1254 | n1337 ;
  assign n1815 = n472 | n1814 ;
  assign n1816 = n1813 | n1815 ;
  assign n1817 = n300 | n345 ;
  assign n1818 = n81 | n1817 ;
  assign n1819 = n146 | n1818 ;
  assign n1820 = n1816 | n1819 ;
  assign n1821 = n1271 | n1820 ;
  assign n1822 = n1810 | n1821 ;
  assign n1823 = n488 | n621 ;
  assign n1824 = n262 | n628 ;
  assign n1825 = n1823 | n1824 ;
  assign n1826 = n417 | n592 ;
  assign n1827 = n390 | n1826 ;
  assign n1828 = n1825 | n1827 ;
  assign n1829 = n114 | n174 ;
  assign n1830 = n1828 | n1829 ;
  assign n1831 = n267 | n404 ;
  assign n1832 = n172 | n1831 ;
  assign n1833 = n143 | n1832 ;
  assign n1834 = n276 | n522 ;
  assign n1835 = n972 | n1834 ;
  assign n1836 = n226 & ~n1835 ;
  assign n1837 = n133 | n391 ;
  assign n1838 = n1316 | n1544 ;
  assign n1839 = n500 | n1838 ;
  assign n1840 = ( n1836 & n1837 ) | ( n1836 & n1839 ) | ( n1837 & n1839 ) ;
  assign n1841 = n1836 & ~n1840 ;
  assign n1842 = ~n1833 & n1841 ;
  assign n1843 = n293 | n476 ;
  assign n1844 = n344 | n1843 ;
  assign n1845 = n108 | n364 ;
  assign n1846 = n338 | n408 ;
  assign n1847 = n160 | n1846 ;
  assign n1848 = n1845 | n1847 ;
  assign n1849 = n1844 | n1848 ;
  assign n1850 = n727 | n1849 ;
  assign n1851 = n1842 & ~n1850 ;
  assign n1852 = n450 | n649 ;
  assign n1853 = n214 | n1852 ;
  assign n1854 = n240 | n1853 ;
  assign n1855 = n191 | n1854 ;
  assign n1856 = n57 | n1855 ;
  assign n1857 = n601 | n1856 ;
  assign n1858 = n1851 & ~n1857 ;
  assign n1859 = n112 | n437 ;
  assign n1860 = n218 | n1859 ;
  assign n1861 = n646 | n1860 ;
  assign n1862 = n1858 & ~n1861 ;
  assign n1863 = ~n1830 & n1862 ;
  assign n1864 = ~n1822 & n1863 ;
  assign n1865 = n383 | n449 ;
  assign n1866 = n102 | n629 ;
  assign n1867 = n111 | n263 ;
  assign n1868 = n311 | n1867 ;
  assign n1869 = n1866 | n1868 ;
  assign n1870 = n1865 | n1869 ;
  assign n1871 = n759 | n1870 ;
  assign n1872 = n514 | n1871 ;
  assign n1873 = n505 | n1872 ;
  assign n1874 = n346 | n1873 ;
  assign n1875 = n670 | n1874 ;
  assign n1876 = n583 | n1875 ;
  assign n1877 = n1864 & ~n1876 ;
  assign n1878 = n65 | n129 ;
  assign n1879 = n661 | n1878 ;
  assign n1880 = n1877 & ~n1879 ;
  assign n1881 = n1803 & ~n1880 ;
  assign n1882 = ~n1803 & n1880 ;
  assign n1883 = n1881 | n1882 ;
  assign n1884 = n280 | n510 ;
  assign n1885 = n638 | n1884 ;
  assign n1886 = n226 & ~n1885 ;
  assign n1887 = n320 | n503 ;
  assign n1888 = n309 | n1887 ;
  assign n1889 = n597 | n646 ;
  assign n1890 = n1463 | n1889 ;
  assign n1891 = n1888 | n1890 ;
  assign n1892 = n416 | n489 ;
  assign n1893 = n165 | n602 ;
  assign n1894 = n1892 | n1893 ;
  assign n1895 = n1891 | n1894 ;
  assign n1896 = n820 | n1629 ;
  assign n1897 = n1895 | n1896 ;
  assign n1898 = n731 | n807 ;
  assign n1899 = n1647 | n1898 ;
  assign n1900 = n995 | n1899 ;
  assign n1901 = n381 | n1900 ;
  assign n1902 = n1897 | n1901 ;
  assign n1903 = n377 | n607 ;
  assign n1904 = n108 | n1903 ;
  assign n1905 = n187 | n1904 ;
  assign n1906 = n1902 | n1905 ;
  assign n1907 = n192 | n374 ;
  assign n1908 = n162 | n222 ;
  assign n1909 = n1907 | n1908 ;
  assign n1910 = n429 | n634 ;
  assign n1911 = n85 | n295 ;
  assign n1912 = n1910 | n1911 ;
  assign n1913 = ( ~n1906 & n1909 ) | ( ~n1906 & n1912 ) | ( n1909 & n1912 ) ;
  assign n1914 = n1906 | n1913 ;
  assign n1915 = n1886 & ~n1914 ;
  assign n1916 = ~n1560 & n1915 ;
  assign n1917 = n483 | n521 ;
  assign n1918 = n364 | n1917 ;
  assign n1919 = n1741 | n1918 ;
  assign n1920 = n417 | n520 ;
  assign n1921 = n168 | n670 ;
  assign n1922 = n1064 | n1921 ;
  assign n1923 = n1920 | n1922 ;
  assign n1924 = n1919 | n1923 ;
  assign n1925 = n197 | n283 ;
  assign n1926 = n608 | n1925 ;
  assign n1927 = n180 | n1926 ;
  assign n1928 = n152 | n1927 ;
  assign n1929 = n1924 | n1928 ;
  assign n1930 = n208 | n1929 ;
  assign n1931 = n755 | n1337 ;
  assign n1932 = n1930 | n1931 ;
  assign n1933 = n127 | n1932 ;
  assign n1934 = n514 | n1933 ;
  assign n1935 = n1916 & ~n1934 ;
  assign n1936 = n266 | n282 ;
  assign n1937 = n277 | n654 ;
  assign n1938 = n1936 | n1937 ;
  assign n1939 = n292 | n1938 ;
  assign n1940 = n356 | n1939 ;
  assign n1941 = n65 | n1940 ;
  assign n1942 = n164 | n1941 ;
  assign n1943 = n640 | n1942 ;
  assign n1944 = n1935 & ~n1943 ;
  assign n1945 = n1880 | n1944 ;
  assign n1946 = n334 | n373 ;
  assign n1947 = n217 | n1946 ;
  assign n1948 = n502 | n1947 ;
  assign n1949 = n263 | n345 ;
  assign n1950 = n366 | n1949 ;
  assign n1951 = n1779 | n1950 ;
  assign n1952 = n1948 | n1951 ;
  assign n1953 = n443 | n1952 ;
  assign n1954 = n157 | n381 ;
  assign n1955 = n1546 | n1954 ;
  assign n1956 = n190 | n380 ;
  assign n1957 = n1379 | n1956 ;
  assign n1958 = n1955 | n1957 ;
  assign n1959 = n250 | n346 ;
  assign n1960 = n309 | n1959 ;
  assign n1961 = n356 | n1960 ;
  assign n1962 = n650 | n1961 ;
  assign n1963 = n1958 | n1962 ;
  assign n1964 = n1953 | n1963 ;
  assign n1965 = n1254 | n1352 ;
  assign n1966 = n169 | n1965 ;
  assign n1967 = n1522 | n1966 ;
  assign n1968 = n468 | n1967 ;
  assign n1969 = n252 | n1968 ;
  assign n1970 = n1964 | n1969 ;
  assign n1971 = n446 | n635 ;
  assign n1972 = n306 | n1971 ;
  assign n1973 = n350 | n697 ;
  assign n1974 = n1794 | n1973 ;
  assign n1975 = n418 | n1057 ;
  assign n1976 = n1354 | n1975 ;
  assign n1977 = n351 | n451 ;
  assign n1978 = n132 | n1977 ;
  assign n1979 = n611 | n1978 ;
  assign n1980 = n420 | n1979 ;
  assign n1981 = n1976 | n1980 ;
  assign n1982 = n1974 | n1981 ;
  assign n1983 = n1972 | n1982 ;
  assign n1984 = n1970 | n1983 ;
  assign n1985 = n240 | n488 ;
  assign n1986 = n1472 | n1985 ;
  assign n1987 = n1471 | n1986 ;
  assign n1988 = n1790 | n1987 ;
  assign n1989 = n100 | n265 ;
  assign n1990 = n102 | n484 ;
  assign n1991 = n1371 | n1990 ;
  assign n1992 = n243 | n1991 ;
  assign n1993 = n1989 | n1992 ;
  assign n1994 = n1988 | n1993 ;
  assign n1995 = n431 | n531 ;
  assign n1996 = n513 | n1995 ;
  assign n1997 = n327 | n1996 ;
  assign n1998 = n383 | n1997 ;
  assign n1999 = n590 | n1998 ;
  assign n2000 = n1994 | n1999 ;
  assign n2001 = n133 | n2000 ;
  assign n2002 = n266 | n580 ;
  assign n2003 = n81 | n2002 ;
  assign n2004 = n1111 | n1187 ;
  assign n2005 = n2003 | n2004 ;
  assign n2006 = n1647 | n2005 ;
  assign n2007 = n1311 | n2006 ;
  assign n2008 = n2001 | n2007 ;
  assign n2009 = n1984 | n2008 ;
  assign n2010 = n990 | n1442 ;
  assign n2011 = n621 | n2010 ;
  assign n2012 = n194 | n2011 ;
  assign n2013 = n2009 | n2012 ;
  assign n2014 = n307 | n488 ;
  assign n2015 = n1371 | n2014 ;
  assign n2016 = n790 | n2015 ;
  assign n2017 = n1595 | n1778 ;
  assign n2018 = n2016 | n2017 ;
  assign n2019 = n1756 | n2018 ;
  assign n2020 = n245 | n432 ;
  assign n2021 = n499 | n522 ;
  assign n2022 = n2020 | n2021 ;
  assign n2023 = n280 | n503 ;
  assign n2024 = n570 | n2023 ;
  assign n2025 = n2022 | n2024 ;
  assign n2026 = n403 | n2025 ;
  assign n2027 = n807 | n2026 ;
  assign n2028 = n2019 | n2027 ;
  assign n2029 = n260 | n356 ;
  assign n2030 = n1959 | n2029 ;
  assign n2031 = n277 | n2030 ;
  assign n2032 = n839 | n2031 ;
  assign n2033 = n315 | n2032 ;
  assign n2034 = n358 | n2033 ;
  assign n2035 = n2028 | n2034 ;
  assign n2036 = n258 | n569 ;
  assign n2037 = n46 | n313 ;
  assign n2038 = n2036 | n2037 ;
  assign n2039 = n849 | n911 ;
  assign n2040 = n2038 | n2039 ;
  assign n2041 = n489 | n1372 ;
  assign n2042 = n628 | n2041 ;
  assign n2043 = n2040 | n2042 ;
  assign n2044 = n293 | n498 ;
  assign n2045 = n125 | n2044 ;
  assign n2046 = n226 & ~n2045 ;
  assign n2047 = ~n445 & n2046 ;
  assign n2048 = ~n2043 & n2047 ;
  assign n2049 = ~n81 & n2048 ;
  assign n2050 = n374 | n1288 ;
  assign n2051 = n275 | n2050 ;
  assign n2052 = n309 | n483 ;
  assign n2053 = n58 | n595 ;
  assign n2054 = n2052 | n2053 ;
  assign n2055 = n103 | n111 ;
  assign n2056 = n2054 | n2055 ;
  assign n2057 = n2051 | n2056 ;
  assign n2058 = n2049 & ~n2057 ;
  assign n2059 = ~n2035 & n2058 ;
  assign n2060 = n540 | n625 ;
  assign n2061 = n1094 | n2060 ;
  assign n2062 = n618 | n887 ;
  assign n2063 = n2061 | n2062 ;
  assign n2064 = n262 | n579 ;
  assign n2065 = n452 | n2064 ;
  assign n2066 = n203 | n2065 ;
  assign n2067 = n2063 | n2066 ;
  assign n2068 = n217 | n645 ;
  assign n2069 = n2067 | n2068 ;
  assign n2070 = n339 | n520 ;
  assign n2071 = n160 | n269 ;
  assign n2072 = n243 | n2071 ;
  assign n2073 = n2070 | n2072 ;
  assign n2074 = n1024 | n1351 ;
  assign n2075 = n688 | n2074 ;
  assign n2076 = n2073 | n2075 ;
  assign n2077 = n284 | n1417 ;
  assign n2078 = n639 | n655 ;
  assign n2079 = n152 | n2078 ;
  assign n2080 = n2077 | n2079 ;
  assign n2081 = n401 | n1297 ;
  assign n2082 = n2080 | n2081 ;
  assign n2083 = n2076 | n2082 ;
  assign n2084 = n2069 | n2083 ;
  assign n2085 = n653 | n1865 ;
  assign n2086 = n334 | n2085 ;
  assign n2087 = n291 | n2086 ;
  assign n2088 = n55 | n2087 ;
  assign n2089 = n2084 | n2088 ;
  assign n2090 = n1079 | n1425 ;
  assign n2091 = n2089 | n2090 ;
  assign n2092 = n2059 & ~n2091 ;
  assign n2093 = n237 | n635 ;
  assign n2094 = n539 | n2093 ;
  assign n2095 = n299 | n2094 ;
  assign n2096 = n327 | n2095 ;
  assign n2097 = n276 | n2096 ;
  assign n2098 = n419 | n2097 ;
  assign n2099 = n212 | n2098 ;
  assign n2100 = n408 | n2099 ;
  assign n2101 = n2092 & ~n2100 ;
  assign n2102 = n187 | n224 ;
  assign n2103 = n2101 & ~n2102 ;
  assign n2104 = n2013 & ~n2103 ;
  assign n2105 = ~n2013 & n2103 ;
  assign n2106 = n2104 | n2105 ;
  assign n2107 = n801 | n1214 ;
  assign n2108 = n2037 | n2107 ;
  assign n2109 = n301 | n569 ;
  assign n2110 = n208 | n2109 ;
  assign n2111 = ( n482 & ~n1947 ) | ( n482 & n2110 ) | ( ~n1947 & n2110 ) ;
  assign n2112 = n1947 | n2111 ;
  assign n2113 = n2108 | n2112 ;
  assign n2114 = n513 | n633 ;
  assign n2115 = n300 | n2114 ;
  assign n2116 = ( ~n1121 & n2113 ) | ( ~n1121 & n2115 ) | ( n2113 & n2115 ) ;
  assign n2117 = n1121 | n2116 ;
  assign n2118 = n595 | n2117 ;
  assign n2119 = n260 | n393 ;
  assign n2120 = n1714 | n2119 ;
  assign n2121 = n282 | n335 ;
  assign n2122 = n438 | n583 ;
  assign n2123 = n2121 | n2122 ;
  assign n2124 = n2120 | n2123 ;
  assign n2125 = n1041 | n2124 ;
  assign n2126 = n390 | n408 ;
  assign n2127 = n947 | n2126 ;
  assign n2128 = n1844 | n2127 ;
  assign n2129 = n244 | n504 ;
  assign n2130 = n252 | n2129 ;
  assign n2131 = ( ~n1101 & n2128 ) | ( ~n1101 & n2130 ) | ( n2128 & n2130 ) ;
  assign n2132 = n1101 | n2131 ;
  assign n2133 = n2125 | n2132 ;
  assign n2134 = n2118 | n2133 ;
  assign n2135 = n922 | n1920 ;
  assign n2136 = n718 | n2135 ;
  assign n2137 = n278 | n2136 ;
  assign n2138 = n479 | n2137 ;
  assign n2139 = n621 | n2138 ;
  assign n2140 = n2134 | n2139 ;
  assign n2141 = n326 | n500 ;
  assign n2142 = n291 | n2141 ;
  assign n2143 = n269 | n2142 ;
  assign n2144 = n292 | n2143 ;
  assign n2145 = n58 | n2144 ;
  assign n2146 = n207 | n489 ;
  assign n2147 = n55 | n579 ;
  assign n2148 = n383 | n625 ;
  assign n2149 = n2147 | n2148 ;
  assign n2150 = n123 | n2149 ;
  assign n2151 = n2146 | n2150 ;
  assign n2152 = n952 | n2151 ;
  assign n2153 = n119 | n2152 ;
  assign n2154 = n199 | n384 ;
  assign n2155 = n473 | n2154 ;
  assign n2156 = n274 | n310 ;
  assign n2157 = n649 | n2156 ;
  assign n2158 = n2155 | n2157 ;
  assign n2159 = n1429 | n2158 ;
  assign n2160 = n2153 | n2159 ;
  assign n2161 = n2145 | n2160 ;
  assign n2162 = n2140 | n2161 ;
  assign n2163 = n429 | n626 ;
  assign n2164 = n457 | n509 ;
  assign n2165 = n283 | n452 ;
  assign n2166 = n2164 | n2165 ;
  assign n2167 = n959 | n1985 ;
  assign n2168 = n2166 | n2167 ;
  assign n2169 = n400 | n514 ;
  assign n2170 = n243 | n2169 ;
  assign n2171 = n540 | n2170 ;
  assign n2172 = n2168 | n2171 ;
  assign n2173 = n249 | n619 ;
  assign n2174 = n253 | n2173 ;
  assign n2175 = n451 | n2174 ;
  assign n2176 = n2172 | n2175 ;
  assign n2177 = n137 | n147 ;
  assign n2178 = n193 | n204 ;
  assign n2179 = n295 | n607 ;
  assign n2180 = n2178 | n2179 ;
  assign n2181 = n622 | n1246 ;
  assign n2182 = n2180 | n2181 ;
  assign n2183 = n263 | n653 ;
  assign n2184 = n351 | n2183 ;
  assign n2185 = n592 | n2184 ;
  assign n2186 = n2182 | n2185 ;
  assign n2187 = n2177 | n2186 ;
  assign n2188 = n2176 | n2187 ;
  assign n2189 = n2163 | n2188 ;
  assign n2190 = n634 | n2189 ;
  assign n2191 = n639 | n2190 ;
  assign n2192 = n2162 | n2191 ;
  assign n2193 = n637 | n2192 ;
  assign n2194 = n2013 & n2193 ;
  assign n2195 = n2013 | n2193 ;
  assign n2196 = ~n2194 & n2195 ;
  assign n2197 = n237 | n359 ;
  assign n2198 = n590 | n2197 ;
  assign n2199 = n99 | n417 ;
  assign n2200 = n622 | n2199 ;
  assign n2201 = n2198 | n2200 ;
  assign n2202 = n295 | n601 ;
  assign n2203 = n441 | n2202 ;
  assign n2204 = n146 | n2203 ;
  assign n2205 = n2201 | n2204 ;
  assign n2206 = n208 | n2205 ;
  assign n2207 = n187 | n669 ;
  assign n2208 = n320 | n449 ;
  assign n2209 = n114 | n2208 ;
  assign n2210 = n215 | n249 ;
  assign n2211 = n1064 | n2210 ;
  assign n2212 = n2209 | n2211 ;
  assign n2213 = n2207 | n2212 ;
  assign n2214 = n2206 | n2213 ;
  assign n2215 = n1601 | n1681 ;
  assign n2216 = n364 | n431 ;
  assign n2217 = n378 | n2216 ;
  assign n2218 = n2215 | n2217 ;
  assign n2219 = n52 | n393 ;
  assign n2220 = n350 | n2219 ;
  assign n2221 = n191 | n310 ;
  assign n2222 = n520 | n2221 ;
  assign n2223 = n2220 | n2222 ;
  assign n2224 = n2218 | n2223 ;
  assign n2225 = n315 | n349 ;
  assign n2226 = n582 | n2225 ;
  assign n2227 = n437 | n2226 ;
  assign n2228 = n83 | n2227 ;
  assign n2229 = n2224 | n2228 ;
  assign n2230 = n2214 | n2229 ;
  assign n2231 = n435 | n569 ;
  assign n2232 = n174 | n2231 ;
  assign n2233 = n1246 | n2232 ;
  assign n2234 = n55 | n245 ;
  assign n2235 = n217 | n2234 ;
  assign n2236 = n1164 | n2235 ;
  assign n2237 = n2233 | n2236 ;
  assign n2238 = n265 | n476 ;
  assign n2239 = n843 | n2238 ;
  assign n2240 = n175 | n383 ;
  assign n2241 = n647 | n2240 ;
  assign n2242 = n2239 | n2241 ;
  assign n2243 = n1329 | n2242 ;
  assign n2244 = n2237 | n2243 ;
  assign n2245 = n470 | n633 ;
  assign n2246 = n253 | n505 ;
  assign n2247 = n2245 | n2246 ;
  assign n2248 = n326 | n346 ;
  assign n2249 = n607 | n2248 ;
  assign n2250 = n2247 | n2249 ;
  assign n2251 = n58 | n125 ;
  assign n2252 = n2250 | n2251 ;
  assign n2253 = n1254 | n2252 ;
  assign n2254 = n2244 | n2253 ;
  assign n2255 = n335 | n636 ;
  assign n2256 = n299 | n2255 ;
  assign n2257 = n180 | n2256 ;
  assign n2258 = n2254 | n2257 ;
  assign n2259 = n2230 | n2258 ;
  assign n2260 = n528 | n1791 ;
  assign n2261 = n1368 | n2260 ;
  assign n2262 = n1751 | n2261 ;
  assign n2263 = n130 | n1372 ;
  assign n2264 = n592 | n2263 ;
  assign n2265 = n1020 | n2264 ;
  assign n2266 = n2262 | n2265 ;
  assign n2267 = n194 | n300 ;
  assign n2268 = n213 | n351 ;
  assign n2269 = n2267 | n2268 ;
  assign n2270 = n164 | n2269 ;
  assign n2271 = n169 | n308 ;
  assign n2272 = n468 | n498 ;
  assign n2273 = n292 | n2272 ;
  assign n2274 = n2271 | n2273 ;
  assign n2275 = n688 | n849 ;
  assign n2276 = n2274 | n2275 ;
  assign n2277 = n2270 | n2276 ;
  assign n2278 = n2266 | n2277 ;
  assign n2279 = n959 | n2003 ;
  assign n2280 = n432 | n2279 ;
  assign n2281 = n384 | n2280 ;
  assign n2282 = n358 | n2281 ;
  assign n2283 = n2278 | n2282 ;
  assign n2284 = n160 | n442 ;
  assign n2285 = n2283 | n2284 ;
  assign n2286 = n2259 | n2285 ;
  assign n2287 = n1284 | n1659 ;
  assign n2288 = n1417 | n2287 ;
  assign n2289 = n391 | n2288 ;
  assign n2290 = n1747 | n2289 ;
  assign n2291 = n355 | n2290 ;
  assign n2292 = n457 | n2291 ;
  assign n2293 = n143 | n2292 ;
  assign n2294 = n145 | n2293 ;
  assign n2295 = n2286 | n2294 ;
  assign n2296 = n650 | n2295 ;
  assign n2297 = n2193 | n2296 ;
  assign n2298 = n2196 & n2297 ;
  assign n2299 = n2193 & n2296 ;
  assign n2300 = n2196 & n2299 ;
  assign n2301 = n434 | n697 ;
  assign n2302 = n269 | n273 ;
  assign n2303 = n212 | n2302 ;
  assign n2304 = n2301 | n2303 ;
  assign n2305 = n151 | n590 ;
  assign n2306 = n313 | n334 ;
  assign n2307 = n2305 | n2306 ;
  assign n2308 = n2304 | n2307 ;
  assign n2309 = n241 | n520 ;
  assign n2310 = n197 | n437 ;
  assign n2311 = n2309 | n2310 ;
  assign n2312 = n966 | n2311 ;
  assign n2313 = n1368 | n2312 ;
  assign n2314 = n2308 | n2313 ;
  assign n2315 = n133 | n295 ;
  assign n2316 = n1469 | n2315 ;
  assign n2317 = n366 | n420 ;
  assign n2318 = n198 | n2317 ;
  assign n2319 = n2316 | n2318 ;
  assign n2320 = ~n191 & n226 ;
  assign n2321 = ~n364 & n2320 ;
  assign n2322 = ~n2319 & n2321 ;
  assign n2323 = ~n1442 & n2322 ;
  assign n2324 = ~n2314 & n2323 ;
  assign n2325 = n428 | n475 ;
  assign n2326 = n654 | n2325 ;
  assign n2327 = n408 | n2326 ;
  assign n2328 = n227 | n2327 ;
  assign n2329 = n960 | n2328 ;
  assign n2330 = n649 | n2329 ;
  assign n2331 = n2324 & ~n2330 ;
  assign n2332 = n110 | n476 ;
  assign n2333 = n601 | n2332 ;
  assign n2334 = n578 | n2333 ;
  assign n2335 = n175 | n2334 ;
  assign n2336 = n975 | n2335 ;
  assign n2337 = n710 | n2336 ;
  assign n2338 = n2331 & ~n2337 ;
  assign n2339 = n59 | n1906 ;
  assign n2340 = n2338 & ~n2339 ;
  assign n2341 = n83 | n628 ;
  assign n2342 = n1778 | n2341 ;
  assign n2343 = n66 | n2342 ;
  assign n2344 = n167 | n451 ;
  assign n2345 = n635 | n779 ;
  assign n2346 = n282 | n636 ;
  assign n2347 = n2345 | n2346 ;
  assign n2348 = n2344 | n2347 ;
  assign n2349 = n2343 | n2348 ;
  assign n2350 = n244 | n470 ;
  assign n2351 = n530 | n2350 ;
  assign n2352 = n519 | n2351 ;
  assign n2353 = n240 | n2352 ;
  assign n2354 = n2349 | n2353 ;
  assign n2355 = n90 | n213 ;
  assign n2356 = n252 | n292 ;
  assign n2357 = n384 | n2356 ;
  assign n2358 = ( n77 & ~n2355 ) | ( n77 & n2357 ) | ( ~n2355 & n2357 ) ;
  assign n2359 = n2355 | n2358 ;
  assign n2360 = n2354 | n2359 ;
  assign n2361 = n180 | n2360 ;
  assign n2362 = n46 | n155 ;
  assign n2363 = n443 | n2362 ;
  assign n2364 = n1659 | n2363 ;
  assign n2365 = n1253 | n2364 ;
  assign n2366 = n2069 | n2365 ;
  assign n2367 = n2361 | n2366 ;
  assign n2368 = n621 | n2367 ;
  assign n2369 = n2340 & ~n2368 ;
  assign n2370 = n270 | n276 ;
  assign n2371 = ( n457 & ~n2055 ) | ( n457 & n2370 ) | ( ~n2055 & n2370 ) ;
  assign n2372 = n2055 | n2371 ;
  assign n2373 = n99 | n2372 ;
  assign n2374 = n128 | n2373 ;
  assign n2375 = n2369 & ~n2374 ;
  assign n2376 = n2296 & ~n2375 ;
  assign n2377 = ~n2296 & n2375 ;
  assign n2378 = n2376 | n2377 ;
  assign n2379 = n2324 & ~n2328 ;
  assign n2380 = n306 | n315 ;
  assign n2381 = n194 | n416 ;
  assign n2382 = n2380 | n2381 ;
  assign n2383 = n96 | n175 ;
  assign n2384 = n94 | n2383 ;
  assign n2385 = n2382 | n2384 ;
  assign n2386 = n372 | n1989 ;
  assign n2387 = n1220 | n1884 ;
  assign n2388 = n2386 | n2387 ;
  assign n2389 = n409 | n628 ;
  assign n2390 = n669 | n2389 ;
  assign n2391 = n349 | n2390 ;
  assign n2392 = n2388 | n2391 ;
  assign n2393 = n505 | n622 ;
  assign n2394 = n618 | n621 ;
  assign n2395 = n2393 | n2394 ;
  assign n2396 = n650 | n2395 ;
  assign n2397 = n143 | n419 ;
  assign n2398 = n2396 | n2397 ;
  assign n2399 = n2392 | n2398 ;
  assign n2400 = n431 | n438 ;
  assign n2401 = n134 | n335 ;
  assign n2402 = n1160 | n2401 ;
  assign n2403 = n326 | n327 ;
  assign n2404 = n161 | n2403 ;
  assign n2405 = n2402 | n2404 ;
  assign n2406 = n2400 | n2405 ;
  assign n2407 = n2399 | n2406 ;
  assign n2408 = n2385 | n2407 ;
  assign n2409 = n2379 & ~n2408 ;
  assign n2410 = n569 | n582 ;
  assign n2411 = n203 | n338 ;
  assign n2412 = n565 | n2146 ;
  assign n2413 = n2411 | n2412 ;
  assign n2414 = n266 | n379 ;
  assign n2415 = n344 | n442 ;
  assign n2416 = n2414 | n2415 ;
  assign n2417 = n1866 | n2416 ;
  assign n2418 = n2413 | n2417 ;
  assign n2419 = n1170 | n1254 ;
  assign n2420 = n1260 | n2419 ;
  assign n2421 = n488 | n2420 ;
  assign n2422 = n2418 | n2421 ;
  assign n2423 = n262 | n529 ;
  assign n2424 = n249 | n2423 ;
  assign n2425 = n112 | n2424 ;
  assign n2426 = n157 | n2425 ;
  assign n2427 = n2422 | n2426 ;
  assign n2428 = n2410 | n2427 ;
  assign n2429 = n127 | n2428 ;
  assign n2430 = n2409 & ~n2429 ;
  assign n2431 = n546 | n927 ;
  assign n2432 = n1239 | n2431 ;
  assign n2433 = n155 | n320 ;
  assign n2434 = n62 | n165 ;
  assign n2435 = n378 | n2434 ;
  assign n2436 = n2433 | n2435 ;
  assign n2437 = n609 | n2436 ;
  assign n2438 = n2432 | n2437 ;
  assign n2439 = n291 | n958 ;
  assign n2440 = n292 | n2439 ;
  assign n2441 = n57 | n2440 ;
  assign n2442 = n81 | n2441 ;
  assign n2443 = n2438 | n2442 ;
  assign n2444 = n122 | n224 ;
  assign n2445 = n2443 | n2444 ;
  assign n2446 = n504 | n2445 ;
  assign n2447 = n310 | n2446 ;
  assign n2448 = n2430 & ~n2447 ;
  assign n2449 = n252 | n319 ;
  assign n2450 = n597 | n2449 ;
  assign n2451 = n393 | n2450 ;
  assign n2452 = n601 | n2451 ;
  assign n2453 = n168 | n2452 ;
  assign n2454 = n129 | n2453 ;
  assign n2455 = n2448 & ~n2454 ;
  assign n2456 = n2375 | n2455 ;
  assign n2457 = n2375 & n2455 ;
  assign n2458 = n933 | n1315 ;
  assign n2459 = n132 | n2458 ;
  assign n2460 = n191 | n595 ;
  assign n2461 = n437 | n2460 ;
  assign n2462 = n2216 | n2461 ;
  assign n2463 = n2459 | n2462 ;
  assign n2464 = n1852 | n2210 ;
  assign n2465 = n503 | n2464 ;
  assign n2466 = n266 | n2465 ;
  assign n2467 = n2463 | n2466 ;
  assign n2468 = n120 | n327 ;
  assign n2469 = n99 | n2468 ;
  assign n2470 = n218 | n2469 ;
  assign n2471 = n2467 | n2470 ;
  assign n2472 = n381 | n510 ;
  assign n2473 = n597 | n2472 ;
  assign n2474 = n134 | n276 ;
  assign n2475 = n2473 | n2474 ;
  assign n2476 = n213 | n242 ;
  assign n2477 = n81 | n2476 ;
  assign n2478 = n1214 | n2477 ;
  assign n2479 = n2475 | n2478 ;
  assign n2480 = n710 | n2479 ;
  assign n2481 = n377 | n482 ;
  assign n2482 = n911 | n2481 ;
  assign n2483 = n350 | n468 ;
  assign n2484 = n313 | n2483 ;
  assign n2485 = n2482 | n2484 ;
  assign n2486 = n100 | n591 ;
  assign n2487 = n180 | n2486 ;
  assign n2488 = n2485 | n2487 ;
  assign n2489 = n2480 | n2488 ;
  assign n2490 = n2471 | n2489 ;
  assign n2491 = n430 | n1574 ;
  assign n2492 = n209 | n2491 ;
  assign n2493 = n489 | n2492 ;
  assign n2494 = n521 | n2493 ;
  assign n2495 = n282 | n2494 ;
  assign n2496 = n240 | n2495 ;
  assign n2497 = n2490 | n2496 ;
  assign n2498 = n52 | n65 ;
  assign n2499 = n2497 | n2498 ;
  assign n2500 = n472 | n490 ;
  assign n2501 = n1016 | n2500 ;
  assign n2502 = n351 | n608 ;
  assign n2503 = n57 | n2502 ;
  assign n2504 = n2501 | n2503 ;
  assign n2505 = n152 | n165 ;
  assign n2506 = n2504 | n2505 ;
  assign n2507 = n92 | n250 ;
  assign n2508 = n174 | n2507 ;
  assign n2509 = n416 | n2508 ;
  assign n2510 = n146 | n2509 ;
  assign n2511 = n283 | n319 ;
  assign n2512 = n1536 | n2511 ;
  assign n2513 = n2510 | n2512 ;
  assign n2514 = n1680 | n2513 ;
  assign n2515 = n204 | n645 ;
  assign n2516 = n928 | n2515 ;
  assign n2517 = n244 | n1066 ;
  assign n2518 = n2516 | n2517 ;
  assign n2519 = n419 | n619 ;
  assign n2520 = n379 | n2519 ;
  assign n2521 = n198 | n2520 ;
  assign n2522 = n2518 | n2521 ;
  assign n2523 = n46 | n94 ;
  assign n2524 = n133 | n2523 ;
  assign n2525 = n2522 | n2524 ;
  assign n2526 = n2514 | n2525 ;
  assign n2527 = n445 | n530 ;
  assign n2528 = n1023 | n2527 ;
  assign n2529 = n1280 | n2528 ;
  assign n2530 = n2410 | n2529 ;
  assign n2531 = n483 | n2530 ;
  assign n2532 = n356 | n2531 ;
  assign n2533 = n2526 | n2532 ;
  assign n2534 = n458 | n519 ;
  assign n2535 = ( ~n458 & n1222 ) | ( ~n458 & n2534 ) | ( n1222 & n2534 ) ;
  assign n2536 = n408 | n2535 ;
  assign n2537 = n514 | n531 ;
  assign n2538 = n193 | n2537 ;
  assign n2539 = n2207 | n2538 ;
  assign n2540 = n2536 | n2539 ;
  assign n2541 = n383 | n428 ;
  assign n2542 = n110 | n2541 ;
  assign n2543 = n2540 | n2542 ;
  assign n2544 = n869 | n2393 ;
  assign n2545 = n309 | n2544 ;
  assign n2546 = n335 | n499 ;
  assign n2547 = n441 | n451 ;
  assign n2548 = n2546 | n2547 ;
  assign n2549 = n2545 | n2548 ;
  assign n2550 = n76 | n640 ;
  assign n2551 = n224 | n2550 ;
  assign n2552 = n2549 | n2551 ;
  assign n2553 = n2543 | n2552 ;
  assign n2554 = n2533 | n2553 ;
  assign n2555 = n2506 | n2554 ;
  assign n2556 = n2499 | n2555 ;
  assign n2557 = n144 | n568 ;
  assign n2558 = n638 | n2557 ;
  assign n2559 = n127 | n2558 ;
  assign n2560 = n488 | n2559 ;
  assign n2561 = n478 | n2560 ;
  assign n2562 = n237 | n2561 ;
  assign n2563 = n444 | n2562 ;
  assign n2564 = n172 | n2563 ;
  assign n2565 = n167 | n2564 ;
  assign n2566 = n2556 | n2565 ;
  assign n2567 = n85 | n647 ;
  assign n2568 = n650 | n2567 ;
  assign n2569 = n2566 | n2568 ;
  assign n2570 = n833 | n1159 ;
  assign n2571 = n1778 | n1845 ;
  assign n2572 = n2570 | n2571 ;
  assign n2573 = n1077 | n2572 ;
  assign n2574 = n1050 | n2573 ;
  assign n2575 = n1350 & ~n2574 ;
  assign n2576 = n269 | n349 ;
  assign n2577 = n359 | n404 ;
  assign n2578 = n2576 | n2577 ;
  assign n2579 = n204 | n627 ;
  assign n2580 = n2578 | n2579 ;
  assign n2581 = n120 | n408 ;
  assign n2582 = n174 | n2581 ;
  assign n2583 = n132 | n2582 ;
  assign n2584 = n2580 | n2583 ;
  assign n2585 = n428 | n583 ;
  assign n2586 = n457 | n2585 ;
  assign n2587 = n2301 | n2586 ;
  assign n2588 = n315 | n482 ;
  assign n2589 = n446 | n2588 ;
  assign n2590 = n639 | n2589 ;
  assign n2591 = n2587 | n2590 ;
  assign n2592 = n358 | n381 ;
  assign n2593 = n449 | n2592 ;
  assign n2594 = n85 | n2593 ;
  assign n2595 = n650 | n2594 ;
  assign n2596 = n2591 | n2595 ;
  assign n2597 = n2584 | n2596 ;
  assign n2598 = n1990 | n2597 ;
  assign n2599 = n278 | n2598 ;
  assign n2600 = n483 | n2599 ;
  assign n2601 = n2575 & ~n2600 ;
  assign n2602 = n244 | n592 ;
  assign n2603 = ( n260 & n280 ) | ( n260 & ~n2602 ) | ( n280 & ~n2602 ) ;
  assign n2604 = n2602 | n2603 ;
  assign n2605 = n187 | n2604 ;
  assign n2606 = n2601 & ~n2605 ;
  assign n2607 = n2569 & ~n2606 ;
  assign n2608 = ~n2569 & n2606 ;
  assign n2609 = n2607 | n2608 ;
  assign n2610 = n168 | n350 ;
  assign n2611 = n1601 | n2610 ;
  assign n2612 = n55 | n208 ;
  assign n2613 = n2400 | n2612 ;
  assign n2614 = n2611 | n2613 ;
  assign n2615 = n373 | n380 ;
  assign n2616 = n240 | n2615 ;
  assign n2617 = n301 | n2616 ;
  assign n2618 = n2614 | n2617 ;
  assign n2619 = n384 | n450 ;
  assign n2620 = n145 | n2619 ;
  assign n2621 = n661 | n2620 ;
  assign n2622 = n2618 | n2621 ;
  assign n2623 = n173 | n504 ;
  assign n2624 = n222 | n449 ;
  assign n2625 = n2623 | n2624 ;
  assign n2626 = n223 | n2625 ;
  assign n2627 = n393 | n639 ;
  assign n2628 = n186 | n2627 ;
  assign n2629 = n947 | n2628 ;
  assign n2630 = n2261 | n2629 ;
  assign n2631 = n2626 | n2630 ;
  assign n2632 = n2551 | n2631 ;
  assign n2633 = n2622 | n2632 ;
  assign n2634 = n2533 | n2633 ;
  assign n2635 = n81 | n602 ;
  assign n2636 = n272 | n2635 ;
  assign n2637 = n1337 | n2636 ;
  assign n2638 = n2634 | n2637 ;
  assign n2639 = n409 | n513 ;
  assign n2640 = n226 & ~n601 ;
  assign n2641 = ~n2639 & n2640 ;
  assign n2642 = n358 | n646 ;
  assign n2643 = n503 | n2642 ;
  assign n2644 = n275 | n2344 ;
  assign n2645 = n2643 | n2644 ;
  assign n2646 = n2641 & ~n2645 ;
  assign n2647 = n310 | n570 ;
  assign n2648 = n404 | n2647 ;
  assign n2649 = n141 | n442 ;
  assign n2650 = n2648 | n2649 ;
  assign n2651 = n102 | n437 ;
  assign n2652 = n2650 | n2651 ;
  assign n2653 = n2646 & ~n2652 ;
  assign n2654 = n1336 | n2252 ;
  assign n2655 = n2653 & ~n2654 ;
  assign n2656 = n430 | n638 ;
  assign n2657 = n242 | n2656 ;
  assign n2658 = n291 | n2657 ;
  assign n2659 = n160 | n2658 ;
  assign n2660 = n142 | n2659 ;
  assign n2661 = n2655 & ~n2660 ;
  assign n2662 = ~n132 & n2661 ;
  assign n2663 = n134 | n634 ;
  assign n2664 = n114 | n191 ;
  assign n2665 = n2663 | n2664 ;
  assign n2666 = n2662 & ~n2665 ;
  assign n2667 = ~n2638 & n2666 ;
  assign n2668 = n381 | n1284 ;
  assign n2669 = n420 | n2668 ;
  assign n2670 = n90 | n2669 ;
  assign n2671 = n112 | n2670 ;
  assign n2672 = n2667 & ~n2671 ;
  assign n2673 = n1574 | n1751 ;
  assign n2674 = n1078 | n1544 ;
  assign n2675 = n2673 | n2674 ;
  assign n2676 = n429 | n488 ;
  assign n2677 = n295 | n2676 ;
  assign n2678 = n408 | n2677 ;
  assign n2679 = n2675 | n2678 ;
  assign n2680 = n81 | n140 ;
  assign n2681 = n224 | n2680 ;
  assign n2682 = n2679 | n2681 ;
  assign n2683 = n125 | n172 ;
  assign n2684 = n243 | n2683 ;
  assign n2685 = ~n129 & n226 ;
  assign n2686 = ~n2511 & n2685 ;
  assign n2687 = ~n2684 & n2686 ;
  assign n2688 = n143 | n390 ;
  assign n2689 = n145 | n531 ;
  assign n2690 = n2688 | n2689 ;
  assign n2691 = n1657 | n2690 ;
  assign n2692 = n2687 & ~n2691 ;
  assign n2693 = ~n2682 & n2692 ;
  assign n2694 = n580 | n595 ;
  assign n2695 = n834 | n2694 ;
  assign n2696 = n1164 | n2695 ;
  assign n2697 = n687 | n2696 ;
  assign n2698 = n167 | n393 ;
  assign n2699 = n640 | n2698 ;
  assign n2700 = n522 | n1696 ;
  assign n2701 = n2699 | n2700 ;
  assign n2702 = n198 | n300 ;
  assign n2703 = n2701 | n2702 ;
  assign n2704 = n2697 | n2703 ;
  assign n2705 = n373 | n528 ;
  assign n2706 = n322 | n2705 ;
  assign n2707 = n94 | n366 ;
  assign n2708 = n85 | n2707 ;
  assign n2709 = n2706 | n2708 ;
  assign n2710 = n1920 | n2709 ;
  assign n2711 = n1865 | n2710 ;
  assign n2712 = n2704 | n2711 ;
  assign n2713 = n996 | n1522 ;
  assign n2714 = n346 | n2713 ;
  assign n2715 = n193 | n2714 ;
  assign n2716 = n445 | n2715 ;
  assign n2717 = n152 | n2716 ;
  assign n2718 = n2712 | n2717 ;
  assign n2719 = n2693 & ~n2718 ;
  assign n2720 = n208 | n634 ;
  assign n2721 = n1044 | n2720 ;
  assign n2722 = n470 | n539 ;
  assign n2723 = n281 | n2722 ;
  assign n2724 = n2721 | n2723 ;
  assign n2725 = n626 | n1371 ;
  assign n2726 = n262 | n2725 ;
  assign n2727 = n2724 | n2726 ;
  assign n2728 = n313 | n355 ;
  assign n2729 = n597 | n2728 ;
  assign n2730 = n174 | n2729 ;
  assign n2731 = n2727 | n2730 ;
  assign n2732 = n161 | n237 ;
  assign n2733 = n301 | n2732 ;
  assign n2734 = n399 | n2733 ;
  assign n2735 = n2335 | n2734 ;
  assign n2736 = n472 | n625 ;
  assign n2737 = n240 | n2736 ;
  assign n2738 = n1475 | n2737 ;
  assign n2739 = n441 | n569 ;
  assign n2740 = n2588 | n2739 ;
  assign n2741 = n2738 | n2740 ;
  assign n2742 = n2735 | n2741 ;
  assign n2743 = n2731 | n2742 ;
  assign n2744 = n433 | n1416 ;
  assign n2745 = n869 | n2744 ;
  assign n2746 = n1261 | n2745 ;
  assign n2747 = n511 | n2746 ;
  assign n2748 = n669 | n2747 ;
  assign n2749 = n2743 | n2748 ;
  assign n2750 = n338 | n591 ;
  assign n2751 = n194 | n2750 ;
  assign n2752 = n102 | n2751 ;
  assign n2753 = n2749 | n2752 ;
  assign n2754 = n2719 & ~n2753 ;
  assign n2755 = n555 | n1066 ;
  assign n2756 = n1867 | n2755 ;
  assign n2757 = n101 | n2756 ;
  assign n2758 = n336 | n2757 ;
  assign n2759 = n2147 | n2758 ;
  assign n2760 = n654 | n2759 ;
  assign n2761 = n307 | n2760 ;
  assign n2762 = n435 | n2761 ;
  assign n2763 = n2754 & ~n2762 ;
  assign n2764 = ~n400 & n2763 ;
  assign n2765 = ~n2569 & n2764 ;
  assign n2766 = n2672 | n2765 ;
  assign n2767 = n2609 | n2766 ;
  assign n2768 = n2455 & n2606 ;
  assign n2769 = n2455 | n2606 ;
  assign n2770 = ~n2768 & n2769 ;
  assign n2771 = n2607 & n2770 ;
  assign n2772 = n2769 & ~n2771 ;
  assign n2773 = ( n2767 & n2768 ) | ( n2767 & n2772 ) | ( n2768 & n2772 ) ;
  assign n2774 = ( n2456 & n2457 ) | ( n2456 & n2773 ) | ( n2457 & n2773 ) ;
  assign n2775 = n2378 | n2774 ;
  assign n2776 = ~n2376 & n2775 ;
  assign n2777 = ( n2298 & n2300 ) | ( n2298 & ~n2776 ) | ( n2300 & ~n2776 ) ;
  assign n2778 = n2194 | n2777 ;
  assign n2779 = ~n2106 & n2778 ;
  assign n2780 = n1880 & n1944 ;
  assign n2781 = n1945 & ~n2780 ;
  assign n2782 = n1944 | n2103 ;
  assign n2783 = n1944 & n2103 ;
  assign n2784 = n2782 & ~n2783 ;
  assign n2785 = n2104 & n2784 ;
  assign n2786 = n2782 & ~n2785 ;
  assign n2787 = n2781 & ~n2786 ;
  assign n2788 = n2781 & ~n2783 ;
  assign n2789 = ( n2779 & n2787 ) | ( n2779 & n2788 ) | ( n2787 & n2788 ) ;
  assign n2790 = n1945 & ~n2789 ;
  assign n2791 = n1883 | n2790 ;
  assign n2792 = n1659 | n2511 ;
  assign n2793 = n887 | n2154 ;
  assign n2794 = n2792 | n2793 ;
  assign n2795 = n273 | n292 ;
  assign n2796 = n583 | n2795 ;
  assign n2797 = n102 | n2796 ;
  assign n2798 = n2794 | n2797 ;
  assign n2799 = n85 | n187 ;
  assign n2800 = n217 | n2799 ;
  assign n2801 = n2798 | n2800 ;
  assign n2802 = n204 | n483 ;
  assign n2803 = n2210 | n2802 ;
  assign n2804 = n498 | n634 ;
  assign n2805 = n334 | n2804 ;
  assign n2806 = n2803 | n2805 ;
  assign n2807 = n442 | n2806 ;
  assign n2808 = n732 | n2807 ;
  assign n2809 = n2801 | n2808 ;
  assign n2810 = n122 | n139 ;
  assign n2811 = n861 | n2732 ;
  assign n2812 = n1034 | n2811 ;
  assign n2813 = n959 | n2812 ;
  assign n2814 = n2810 | n2813 ;
  assign n2815 = n468 | n2814 ;
  assign n2816 = n2809 | n2815 ;
  assign n2817 = n300 | n432 ;
  assign n2818 = n83 | n2817 ;
  assign n2819 = n513 | n628 ;
  assign n2820 = n263 | n2819 ;
  assign n2821 = n380 | n2820 ;
  assign n2822 = n90 | n2821 ;
  assign n2823 = n420 | n2822 ;
  assign n2824 = n580 | n2823 ;
  assign n2825 = n2818 | n2824 ;
  assign n2826 = n2816 | n2825 ;
  assign n2827 = n478 | n500 ;
  assign n2828 = n277 | n320 ;
  assign n2829 = n2827 | n2828 ;
  assign n2830 = n133 | n208 ;
  assign n2831 = n2829 | n2830 ;
  assign n2832 = n994 | n1051 ;
  assign n2833 = n2831 | n2832 ;
  assign n2834 = n145 | n647 ;
  assign n2835 = n274 | n313 ;
  assign n2836 = n1936 | n2835 ;
  assign n2837 = n207 | n2836 ;
  assign n2838 = n928 | n2739 ;
  assign n2839 = n2473 | n2838 ;
  assign n2840 = n2837 | n2839 ;
  assign n2841 = n1764 | n2840 ;
  assign n2842 = n609 | n1865 ;
  assign n2843 = n479 | n2842 ;
  assign n2844 = n470 | n2843 ;
  assign n2845 = n252 | n2844 ;
  assign n2846 = n2841 | n2845 ;
  assign n2847 = n400 | n670 ;
  assign n2848 = n226 & ~n2847 ;
  assign n2849 = ( n2834 & ~n2846 ) | ( n2834 & n2848 ) | ( ~n2846 & n2848 ) ;
  assign n2850 = ~n2834 & n2849 ;
  assign n2851 = ~n2833 & n2850 ;
  assign n2852 = ~n2826 & n2851 ;
  assign n2853 = n439 | n1254 ;
  assign n2854 = n2070 | n2853 ;
  assign n2855 = n258 | n2623 ;
  assign n2856 = n1708 | n2855 ;
  assign n2857 = n2854 | n2856 ;
  assign n2858 = n306 | n309 ;
  assign n2859 = n435 | n2858 ;
  assign n2860 = n62 | n2859 ;
  assign n2861 = n2857 | n2860 ;
  assign n2862 = n130 | n2861 ;
  assign n2863 = n367 | n2862 ;
  assign n2864 = n101 | n2863 ;
  assign n2865 = n2393 | n2864 ;
  assign n2866 = n2852 & ~n2865 ;
  assign n2867 = n114 | n653 ;
  assign n2868 = n1253 | n2867 ;
  assign n2869 = n625 | n2868 ;
  assign n2870 = n310 | n2869 ;
  assign n2871 = n358 | n2870 ;
  assign n2872 = n126 | n2871 ;
  assign n2873 = n2866 & ~n2872 ;
  assign n2874 = n1733 | n2873 ;
  assign n2875 = n1733 & n2873 ;
  assign n2876 = n2874 & ~n2875 ;
  assign n2877 = n1803 & ~n2873 ;
  assign n2878 = ~n1803 & n2873 ;
  assign n2879 = n2877 | n2878 ;
  assign n2880 = n1881 & ~n2879 ;
  assign n2881 = n2877 | n2880 ;
  assign n2882 = n2876 & n2881 ;
  assign n2883 = n2874 & ~n2882 ;
  assign n2884 = n2876 & ~n2878 ;
  assign n2885 = n2874 & ~n2884 ;
  assign n2886 = ( n2791 & n2883 ) | ( n2791 & n2885 ) | ( n2883 & n2885 ) ;
  assign n2887 = n1736 | n2886 ;
  assign n2888 = ~n1734 & n2887 ;
  assign n2889 = n300 | n579 ;
  assign n2890 = n52 | n186 ;
  assign n2891 = n2889 | n2890 ;
  assign n2892 = n58 | n625 ;
  assign n2893 = n96 | n2892 ;
  assign n2894 = n1980 | n2893 ;
  assign n2895 = n948 | n2894 ;
  assign n2896 = n2891 | n2895 ;
  assign n2897 = n1970 | n2896 ;
  assign n2898 = n253 | n458 ;
  assign n2899 = n296 | n520 ;
  assign n2900 = n90 | n2899 ;
  assign n2901 = n2898 | n2900 ;
  assign n2902 = n1081 | n2901 ;
  assign n2903 = n161 | n637 ;
  assign n2904 = n278 | n2903 ;
  assign n2905 = n436 | n2904 ;
  assign n2906 = n2641 & ~n2905 ;
  assign n2907 = ~n2902 & n2906 ;
  assign n2908 = n432 | n633 ;
  assign n2909 = n2341 | n2908 ;
  assign n2910 = n364 | n670 ;
  assign n2911 = n2909 | n2910 ;
  assign n2912 = n1990 | n2911 ;
  assign n2913 = n933 | n2912 ;
  assign n2914 = n2907 & ~n2913 ;
  assign n2915 = n391 | n1371 ;
  assign n2916 = n618 | n2915 ;
  assign n2917 = n313 | n2916 ;
  assign n2918 = n111 | n2917 ;
  assign n2919 = n2914 & ~n2918 ;
  assign n2920 = ~n2525 & n2919 ;
  assign n2921 = ~n2897 & n2920 ;
  assign n2922 = n55 | n120 ;
  assign n2923 = n282 | n608 ;
  assign n2924 = n77 | n2923 ;
  assign n2925 = n1687 | n2924 ;
  assign n2926 = n405 | n529 ;
  assign n2927 = n295 | n2926 ;
  assign n2928 = n2925 | n2927 ;
  assign n2929 = n293 | n417 ;
  assign n2930 = n2928 | n2929 ;
  assign n2931 = n2922 | n2930 ;
  assign n2932 = n806 | n2931 ;
  assign n2933 = n514 | n2932 ;
  assign n2934 = n429 | n2933 ;
  assign n2935 = n2921 & ~n2934 ;
  assign n2936 = n314 | n321 ;
  assign n2937 = n384 | n2936 ;
  assign n2938 = n390 | n2937 ;
  assign n2939 = n2935 & ~n2938 ;
  assign n2940 = n1532 & ~n2939 ;
  assign n2941 = ~n1532 & n2939 ;
  assign n2942 = n2940 | n2941 ;
  assign n2943 = n313 | n640 ;
  assign n2944 = n648 | n1544 ;
  assign n2945 = n2943 | n2944 ;
  assign n2946 = n265 | n2945 ;
  assign n2947 = n583 | n2946 ;
  assign n2948 = n449 | n2947 ;
  assign n2949 = n114 | n2948 ;
  assign n2950 = n203 | n314 ;
  assign n2951 = n162 | n2950 ;
  assign n2952 = n227 | n419 ;
  assign n2953 = n888 | n2952 ;
  assign n2954 = n1464 | n2953 ;
  assign n2955 = n2264 | n2954 ;
  assign n2956 = n307 | n380 ;
  assign n2957 = n442 | n569 ;
  assign n2958 = n2956 | n2957 ;
  assign n2959 = n152 | n2958 ;
  assign n2960 = n85 | n597 ;
  assign n2961 = n1118 | n2960 ;
  assign n2962 = n2959 | n2961 ;
  assign n2963 = n2955 | n2962 ;
  assign n2964 = ( n1508 & ~n2951 ) | ( n1508 & n2963 ) | ( ~n2951 & n2963 ) ;
  assign n2965 = n2951 | n2964 ;
  assign n2966 = n2949 | n2965 ;
  assign n2967 = n511 | n529 ;
  assign n2968 = n489 | n530 ;
  assign n2969 = n2967 | n2968 ;
  assign n2970 = n349 | n621 ;
  assign n2971 = n250 | n2970 ;
  assign n2972 = n2969 | n2971 ;
  assign n2973 = n191 | n253 ;
  assign n2974 = ( n77 & n366 ) | ( n77 & ~n2973 ) | ( n366 & ~n2973 ) ;
  assign n2975 = n2973 | n2974 ;
  assign n2976 = n2972 | n2975 ;
  assign n2977 = n157 | n2976 ;
  assign n2978 = n93 | n2393 ;
  assign n2979 = n444 | n2169 ;
  assign n2980 = n2978 | n2979 ;
  assign n2981 = n923 | n1837 ;
  assign n2982 = n172 | n222 ;
  assign n2983 = n2981 | n2982 ;
  assign n2984 = n2980 | n2983 ;
  assign n2985 = n81 | n2984 ;
  assign n2986 = n2977 | n2985 ;
  assign n2987 = n1158 | n2986 ;
  assign n2988 = n2966 | n2987 ;
  assign n2989 = n262 | n299 ;
  assign n2990 = n244 | n274 ;
  assign n2991 = n578 | n2990 ;
  assign n2992 = n2989 | n2991 ;
  assign n2993 = n293 | n435 ;
  assign n2994 = n457 | n2993 ;
  assign n2995 = n260 | n373 ;
  assign n2996 = n403 | n2995 ;
  assign n2997 = n327 | n2996 ;
  assign n2998 = n2994 | n2997 ;
  assign n2999 = n140 | n168 ;
  assign n3000 = n2998 | n2999 ;
  assign n3001 = n2992 | n3000 ;
  assign n3002 = n112 | n164 ;
  assign n3003 = n122 | n3002 ;
  assign n3004 = n126 | n174 ;
  assign n3005 = n355 | n654 ;
  assign n3006 = n450 | n3005 ;
  assign n3007 = n390 | n3006 ;
  assign n3008 = ( ~n2911 & n3004 ) | ( ~n2911 & n3007 ) | ( n3004 & n3007 ) ;
  assign n3009 = n2911 | n3008 ;
  assign n3010 = n3003 | n3009 ;
  assign n3011 = n3001 | n3010 ;
  assign n3012 = n225 | n756 ;
  assign n3013 = n348 | n3012 ;
  assign n3014 = n499 | n3013 ;
  assign n3015 = n280 | n3014 ;
  assign n3016 = n451 | n3015 ;
  assign n3017 = n3011 | n3016 ;
  assign n3018 = n175 | n187 ;
  assign n3019 = n661 | n3018 ;
  assign n3020 = n3017 | n3019 ;
  assign n3021 = n1791 | n3020 ;
  assign n3022 = n2988 | n3021 ;
  assign n3023 = n960 | n1644 ;
  assign n3024 = n1990 | n3023 ;
  assign n3025 = n65 | n3024 ;
  assign n3026 = n197 | n3025 ;
  assign n3027 = n213 | n3026 ;
  assign n3028 = n96 | n3027 ;
  assign n3029 = n649 | n3028 ;
  assign n3030 = n3022 | n3029 ;
  assign n3031 = ~n2939 & n3030 ;
  assign n3032 = n1625 | n3030 ;
  assign n3033 = n2939 & ~n3030 ;
  assign n3034 = n3031 | n3033 ;
  assign n3035 = n3032 & ~n3034 ;
  assign n3036 = n3031 | n3035 ;
  assign n3037 = ~n2942 & n3036 ;
  assign n3038 = n2940 | n3037 ;
  assign n3039 = n1625 & n3030 ;
  assign n3040 = ~n3034 & n3039 ;
  assign n3041 = n3031 | n3040 ;
  assign n3042 = ~n2942 & n3041 ;
  assign n3043 = n2940 | n3042 ;
  assign n3044 = ( ~n2888 & n3038 ) | ( ~n2888 & n3043 ) | ( n3038 & n3043 ) ;
  assign n3045 = ~n1535 & n3044 ;
  assign n3046 = n1533 | n3045 ;
  assign n3047 = n1151 & ~n1327 ;
  assign n3048 = n1328 | n3047 ;
  assign n3049 = n528 | n834 ;
  assign n3050 = n250 | n3049 ;
  assign n3051 = n62 | n3050 ;
  assign n3052 = n125 | n3051 ;
  assign n3053 = n103 | n3052 ;
  assign n3054 = n421 | n1128 ;
  assign n3055 = n265 | n1865 ;
  assign n3056 = n1383 | n3055 ;
  assign n3057 = n240 | n444 ;
  assign n3058 = n607 | n3057 ;
  assign n3059 = n451 | n3058 ;
  assign n3060 = n3056 | n3059 ;
  assign n3061 = n314 | n472 ;
  assign n3062 = n366 | n3061 ;
  assign n3063 = n927 | n1845 ;
  assign n3064 = n3062 | n3063 ;
  assign n3065 = n2163 | n3064 ;
  assign n3066 = n3060 | n3065 ;
  assign n3067 = n1329 | n1578 ;
  assign n3068 = n638 | n3067 ;
  assign n3069 = ( ~n3054 & n3066 ) | ( ~n3054 & n3068 ) | ( n3066 & n3068 ) ;
  assign n3070 = n3054 | n3069 ;
  assign n3071 = n3053 | n3070 ;
  assign n3072 = n139 | n3071 ;
  assign n3073 = n479 | n2393 ;
  assign n3074 = n438 | n571 ;
  assign n3075 = n3073 | n3074 ;
  assign n3076 = n862 | n2867 ;
  assign n3077 = n468 | n625 ;
  assign n3078 = n470 | n3077 ;
  assign n3079 = n3076 | n3078 ;
  assign n3080 = ( ~n1775 & n3075 ) | ( ~n1775 & n3079 ) | ( n3075 & n3079 ) ;
  assign n3081 = n1775 | n3080 ;
  assign n3082 = n1852 | n3081 ;
  assign n3083 = n3072 | n3082 ;
  assign n3084 = n2802 | n2967 ;
  assign n3085 = n282 | n293 ;
  assign n3086 = n356 | n3085 ;
  assign n3087 = n3084 | n3086 ;
  assign n3088 = n191 | n3087 ;
  assign n3089 = n338 | n509 ;
  assign n3090 = n219 | n3089 ;
  assign n3091 = n190 | n274 ;
  assign n3092 = n601 | n3091 ;
  assign n3093 = n3090 | n3092 ;
  assign n3094 = n102 | n152 ;
  assign n3095 = n142 | n3094 ;
  assign n3096 = n3093 | n3095 ;
  assign n3097 = n1069 | n3096 ;
  assign n3098 = n3088 | n3097 ;
  assign n3099 = n1260 | n3098 ;
  assign n3100 = n499 | n3099 ;
  assign n3101 = n258 | n3100 ;
  assign n3102 = n3083 | n3101 ;
  assign n3103 = n457 | n578 ;
  assign n3104 = n3102 | n3103 ;
  assign n3105 = n1327 & n3104 ;
  assign n3106 = n1327 | n3104 ;
  assign n3107 = ~n3105 & n3106 ;
  assign n3108 = n46 | n320 ;
  assign n3109 = n129 | n3108 ;
  assign n3110 = n193 | n622 ;
  assign n3111 = n1656 | n3110 ;
  assign n3112 = n3109 | n3111 ;
  assign n3113 = n1051 | n3112 ;
  assign n3114 = n638 | n1057 ;
  assign n3115 = n224 | n390 ;
  assign n3116 = n3114 | n3115 ;
  assign n3117 = n115 | n3116 ;
  assign n3118 = n3113 | n3117 ;
  assign n3119 = n1376 | n3118 ;
  assign n3120 = n1370 | n3119 ;
  assign n3121 = n110 | n2350 ;
  assign n3122 = n157 | n442 ;
  assign n3123 = n162 | n3122 ;
  assign n3124 = n3121 | n3123 ;
  assign n3125 = n479 | n1434 ;
  assign n3126 = n483 | n3125 ;
  assign n3127 = n3124 | n3126 ;
  assign n3128 = n391 | n468 ;
  assign n3129 = n283 | n3128 ;
  assign n3130 = n327 | n3129 ;
  assign n3131 = n345 | n3130 ;
  assign n3132 = n3127 | n3131 ;
  assign n3133 = n140 | n3132 ;
  assign n3134 = n452 | n592 ;
  assign n3135 = n92 | n3134 ;
  assign n3136 = ( n321 & ~n2648 ) | ( n321 & n3135 ) | ( ~n2648 & n3135 ) ;
  assign n3137 = n2648 | n3136 ;
  assign n3138 = n181 | n3137 ;
  assign n3139 = n3133 | n3138 ;
  assign n3140 = n3120 | n3139 ;
  assign n3141 = n59 | n3140 ;
  assign n3142 = n504 | n670 ;
  assign n3143 = n213 | n602 ;
  assign n3144 = n3142 | n3143 ;
  assign n3145 = n155 | n3144 ;
  assign n3146 = n511 | n639 ;
  assign n3147 = n401 | n3146 ;
  assign n3148 = n3145 | n3147 ;
  assign n3149 = n299 | n488 ;
  assign n3150 = n76 | n190 ;
  assign n3151 = n3149 | n3150 ;
  assign n3152 = n174 | n429 ;
  assign n3153 = n476 | n3152 ;
  assign n3154 = n3151 | n3153 ;
  assign n3155 = n314 | n500 ;
  assign n3156 = n260 | n3155 ;
  assign n3157 = n451 | n3156 ;
  assign n3158 = n3154 | n3157 ;
  assign n3159 = n3148 | n3158 ;
  assign n3160 = n1959 | n2112 ;
  assign n3161 = n568 | n3160 ;
  assign n3162 = n3159 | n3161 ;
  assign n3163 = n503 | n862 ;
  assign n3164 = n273 | n3163 ;
  assign n3165 = n203 | n3164 ;
  assign n3166 = n364 | n3165 ;
  assign n3167 = n165 | n3166 ;
  assign n3168 = n3162 | n3167 ;
  assign n3169 = n85 | n100 ;
  assign n3170 = n133 | n3169 ;
  assign n3171 = n3168 | n3170 ;
  assign n3172 = n1254 | n3171 ;
  assign n3173 = n3141 | n3172 ;
  assign n3174 = n472 | n1284 ;
  assign n3175 = n380 | n3174 ;
  assign n3176 = n306 | n3175 ;
  assign n3177 = n640 | n3176 ;
  assign n3178 = n3173 | n3177 ;
  assign n3179 = n3104 & n3178 ;
  assign n3180 = n1411 & ~n3178 ;
  assign n3181 = n3104 | n3178 ;
  assign n3182 = ~n3179 & n3181 ;
  assign n3183 = ~n3180 & n3182 ;
  assign n3184 = n3179 | n3183 ;
  assign n3185 = n3107 & n3184 ;
  assign n3186 = n3105 | n3185 ;
  assign n3187 = ~n3048 & n3186 ;
  assign n3188 = ~n1411 & n3178 ;
  assign n3189 = n3182 & n3188 ;
  assign n3190 = n3179 | n3189 ;
  assign n3191 = n3107 & n3190 ;
  assign n3192 = n3105 | n3191 ;
  assign n3193 = ~n3048 & n3192 ;
  assign n3194 = ( n3046 & n3187 ) | ( n3046 & n3193 ) | ( n3187 & n3193 ) ;
  assign n3195 = n1328 | n3194 ;
  assign n3196 = ~n1236 & n3195 ;
  assign n3197 = ~n904 & n1014 ;
  assign n3198 = n1015 | n3197 ;
  assign n3199 = n711 | n2411 ;
  assign n3200 = n2209 | n3199 ;
  assign n3201 = n1578 | n1921 ;
  assign n3202 = n808 | n3201 ;
  assign n3203 = n3200 | n3202 ;
  assign n3204 = n172 | n619 ;
  assign n3205 = n960 | n1443 ;
  assign n3206 = n2393 | n3205 ;
  assign n3207 = n3204 | n3206 ;
  assign n3208 = n3203 | n3207 ;
  assign n3209 = n253 | n509 ;
  assign n3210 = n400 | n3209 ;
  assign n3211 = n404 | n3210 ;
  assign n3212 = n77 | n3211 ;
  assign n3213 = n133 | n3212 ;
  assign n3214 = n3208 | n3213 ;
  assign n3215 = n661 | n3214 ;
  assign n3216 = n3004 | n3146 ;
  assign n3217 = n570 | n595 ;
  assign n3218 = n223 | n269 ;
  assign n3219 = n3217 | n3218 ;
  assign n3220 = n3216 | n3219 ;
  assign n3221 = n972 | n2221 ;
  assign n3222 = n1329 | n3221 ;
  assign n3223 = n3220 | n3222 ;
  assign n3224 = n351 | n432 ;
  assign n3225 = n1279 | n3224 ;
  assign n3226 = n1128 | n3225 ;
  assign n3227 = n3223 | n3226 ;
  assign n3228 = n313 | n629 ;
  assign n3229 = n646 | n3228 ;
  assign n3230 = n3227 | n3229 ;
  assign n3231 = n212 | n300 ;
  assign n3232 = n165 | n3231 ;
  assign n3233 = ~n85 & n226 ;
  assign n3234 = ~n1221 & n3233 ;
  assign n3235 = ~n3232 & n3234 ;
  assign n3236 = ~n2146 & n3235 ;
  assign n3237 = ~n2347 & n3236 ;
  assign n3238 = n2392 | n2397 ;
  assign n3239 = n3237 & ~n3238 ;
  assign n3240 = ~n3230 & n3239 ;
  assign n3241 = ~n3215 & n3240 ;
  assign n3242 = ~n707 & n3241 ;
  assign n3243 = n46 | n132 ;
  assign n3244 = n1129 | n2126 ;
  assign n3245 = n141 | n530 ;
  assign n3246 = n3244 | n3245 ;
  assign n3247 = n249 | n3246 ;
  assign n3248 = n1079 | n3247 ;
  assign n3249 = n718 | n3248 ;
  assign n3250 = n2029 | n3249 ;
  assign n3251 = n3243 | n3250 ;
  assign n3252 = n359 | n3251 ;
  assign n3253 = n3242 & ~n3252 ;
  assign n3254 = n186 | n218 ;
  assign n3255 = n3253 & ~n3254 ;
  assign n3256 = n1014 | n3255 ;
  assign n3257 = n1014 & n3255 ;
  assign n3258 = n3256 & ~n3257 ;
  assign n3259 = n445 | n450 ;
  assign n3260 = n223 | n3259 ;
  assign n3261 = n194 | n417 ;
  assign n3262 = n92 | n649 ;
  assign n3263 = n889 | n3262 ;
  assign n3264 = n206 | n3263 ;
  assign n3265 = n843 | n2960 ;
  assign n3266 = n490 | n3265 ;
  assign n3267 = n3264 | n3266 ;
  assign n3268 = n522 | n531 ;
  assign n3269 = n505 | n3268 ;
  assign n3270 = n300 | n3269 ;
  assign n3271 = n578 | n3270 ;
  assign n3272 = n3267 | n3271 ;
  assign n3273 = n65 | n3272 ;
  assign n3274 = n377 | n478 ;
  assign n3275 = n166 | n3274 ;
  assign n3276 = n1032 | n1288 ;
  assign n3277 = n3275 | n3276 ;
  assign n3278 = n881 | n3277 ;
  assign n3279 = n326 | n655 ;
  assign n3280 = n611 | n3279 ;
  assign n3281 = n120 | n596 ;
  assign n3282 = n155 | n3281 ;
  assign n3283 = n3280 | n3282 ;
  assign n3284 = n1194 | n3283 ;
  assign n3285 = n3278 | n3284 ;
  assign n3286 = n568 | n3285 ;
  assign n3287 = n3273 | n3286 ;
  assign n3288 = n336 | n1311 ;
  assign n3289 = n834 | n3288 ;
  assign n3290 = n511 | n3289 ;
  assign n3291 = n346 | n3290 ;
  assign n3292 = n217 | n3291 ;
  assign n3293 = n3287 | n3292 ;
  assign n3294 = n203 | n216 ;
  assign n3295 = n146 | n3294 ;
  assign n3296 = n105 | n873 ;
  assign n3297 = n3295 | n3296 ;
  assign n3298 = n82 | n1888 ;
  assign n3299 = n3297 | n3298 ;
  assign n3300 = n96 | n181 ;
  assign n3301 = n1865 | n3300 ;
  assign n3302 = n266 | n2732 ;
  assign n3303 = n3301 | n3302 ;
  assign n3304 = n274 | n400 ;
  assign n3305 = n3303 | n3304 ;
  assign n3306 = n1811 | n3305 ;
  assign n3307 = n3299 | n3306 ;
  assign n3308 = n990 | n2163 ;
  assign n3309 = n1261 | n3308 ;
  assign n3310 = n2029 | n3309 ;
  assign n3311 = n242 | n3310 ;
  assign n3312 = n295 | n3311 ;
  assign n3313 = n3307 | n3312 ;
  assign n3314 = n152 | n379 ;
  assign n3315 = n380 | n579 ;
  assign n3316 = n2739 | n3315 ;
  assign n3317 = n428 | n504 ;
  assign n3318 = n292 | n3317 ;
  assign n3319 = n3316 | n3318 ;
  assign n3320 = n580 | n650 ;
  assign n3321 = n3319 | n3320 ;
  assign n3322 = n58 | n1259 ;
  assign n3323 = n2699 | n3322 ;
  assign n3324 = n514 | n653 ;
  assign n3325 = n172 | n319 ;
  assign n3326 = n3324 | n3325 ;
  assign n3327 = n3323 | n3326 ;
  assign n3328 = n134 | n583 ;
  assign n3329 = n595 | n3328 ;
  assign n3330 = n3327 | n3329 ;
  assign n3331 = n3321 | n3330 ;
  assign n3332 = n3314 | n3331 ;
  assign n3333 = n3313 | n3332 ;
  assign n3334 = n3293 | n3333 ;
  assign n3335 = n791 | n1253 ;
  assign n3336 = n1753 | n3335 ;
  assign n3337 = n483 | n529 ;
  assign n3338 = n250 | n3337 ;
  assign n3339 = n338 | n3338 ;
  assign n3340 = n3336 | n3339 ;
  assign n3341 = n291 | n345 ;
  assign n3342 = n143 | n3341 ;
  assign n3343 = n129 | n3342 ;
  assign n3344 = n3340 | n3343 ;
  assign n3345 = n609 | n3344 ;
  assign n3346 = n625 | n3345 ;
  assign n3347 = ( ~n3261 & n3334 ) | ( ~n3261 & n3346 ) | ( n3334 & n3346 ) ;
  assign n3348 = n3261 | n3347 ;
  assign n3349 = n3260 | n3348 ;
  assign n3350 = ~n3255 & n3349 ;
  assign n3351 = n3255 & ~n3349 ;
  assign n3352 = n3350 | n3351 ;
  assign n3353 = n1233 & n3349 ;
  assign n3354 = n1233 | n3349 ;
  assign n3355 = ~n3353 & n3354 ;
  assign n3356 = n1234 & n3355 ;
  assign n3357 = n3353 | n3356 ;
  assign n3358 = ~n3352 & n3357 ;
  assign n3359 = n3350 | n3358 ;
  assign n3360 = n3258 & n3359 ;
  assign n3361 = n3256 & ~n3360 ;
  assign n3362 = n3198 | n3361 ;
  assign n3363 = ~n3352 & n3354 ;
  assign n3364 = n3350 | n3363 ;
  assign n3365 = n3258 & n3364 ;
  assign n3366 = n3256 & ~n3365 ;
  assign n3367 = n3198 | n3366 ;
  assign n3368 = ( ~n3196 & n3362 ) | ( ~n3196 & n3367 ) | ( n3362 & n3367 ) ;
  assign n3369 = ~n1015 & n3368 ;
  assign n3370 = n907 & ~n3369 ;
  assign n3371 = n143 | n180 ;
  assign n3372 = n2344 | n3371 ;
  assign n3373 = n756 | n2527 ;
  assign n3374 = n3372 | n3373 ;
  assign n3375 = n140 | n172 ;
  assign n3376 = n2810 | n3375 ;
  assign n3377 = n540 | n3376 ;
  assign n3378 = n3374 | n3377 ;
  assign n3379 = n384 | n468 ;
  assign n3380 = n580 | n3379 ;
  assign n3381 = n438 | n3380 ;
  assign n3382 = n403 | n3381 ;
  assign n3383 = n3378 | n3382 ;
  assign n3384 = n94 | n100 ;
  assign n3385 = n108 | n3384 ;
  assign n3386 = n146 | n3385 ;
  assign n3387 = n3383 | n3386 ;
  assign n3388 = n492 | n3301 ;
  assign n3389 = n487 | n3388 ;
  assign n3390 = n529 | n583 ;
  assign n3391 = n450 | n458 ;
  assign n3392 = n3390 | n3391 ;
  assign n3393 = n142 | n3392 ;
  assign n3394 = n86 | n422 ;
  assign n3395 = n3393 | n3394 ;
  assign n3396 = n3389 | n3395 ;
  assign n3397 = n1700 | n3396 ;
  assign n3398 = n3387 | n3397 ;
  assign n3399 = n379 | n472 ;
  assign n3400 = n578 | n3399 ;
  assign n3401 = n377 | n3400 ;
  assign n3402 = n404 | n3401 ;
  assign n3403 = n168 | n3402 ;
  assign n3404 = n99 | n3403 ;
  assign n3405 = n145 | n3404 ;
  assign n3406 = n3398 | n3405 ;
  assign n3407 = ~n115 & n229 ;
  assign n3408 = ~n525 & n3407 ;
  assign n3409 = ~n518 & n3408 ;
  assign n3410 = ~n2722 & n3409 ;
  assign n3411 = n134 | n2635 ;
  assign n3412 = n494 | n3411 ;
  assign n3413 = n590 | n595 ;
  assign n3414 = n601 | n3413 ;
  assign n3415 = n58 | n3414 ;
  assign n3416 = n3412 | n3415 ;
  assign n3417 = n133 | n157 ;
  assign n3418 = n3416 | n3417 ;
  assign n3419 = n3410 & ~n3418 ;
  assign n3420 = ~n187 & n3419 ;
  assign n3421 = ~n3406 & n3420 ;
  assign n3422 = n571 | n2732 ;
  assign n3423 = n430 | n3422 ;
  assign n3424 = n127 | n3423 ;
  assign n3425 = n373 | n3424 ;
  assign n3426 = n444 | n3425 ;
  assign n3427 = n610 | n3426 ;
  assign n3428 = n215 | n3427 ;
  assign n3429 = n57 | n3428 ;
  assign n3430 = n3421 & ~n3429 ;
  assign n3431 = ~n103 & n3430 ;
  assign n3432 = n589 | n3431 ;
  assign n3433 = n589 & n3431 ;
  assign n3434 = n3432 & ~n3433 ;
  assign n3435 = n530 | n650 ;
  assign n3436 = ( n498 & n1161 ) | ( n498 & ~n3435 ) | ( n1161 & ~n3435 ) ;
  assign n3437 = n3435 | n3436 ;
  assign n3438 = n1252 | n3437 ;
  assign n3439 = n245 | n514 ;
  assign n3440 = n2210 | n3439 ;
  assign n3441 = n244 | n653 ;
  assign n3442 = n313 | n3441 ;
  assign n3443 = n3440 | n3442 ;
  assign n3444 = n111 | n3443 ;
  assign n3445 = n791 | n833 ;
  assign n3446 = n3444 | n3445 ;
  assign n3447 = n3438 | n3446 ;
  assign n3448 = n314 | n379 ;
  assign n3449 = n58 | n3448 ;
  assign n3450 = ( n235 & n242 ) | ( n235 & n507 ) | ( n242 & n507 ) ;
  assign n3451 = n3449 | n3450 ;
  assign n3452 = n209 | n3451 ;
  assign n3453 = n127 | n3452 ;
  assign n3454 = n1354 | n3453 ;
  assign n3455 = n3447 | n3454 ;
  assign n3456 = n295 | n519 ;
  assign n3457 = n405 | n1865 ;
  assign n3458 = n513 | n3457 ;
  assign n3459 = ( n250 & ~n3456 ) | ( n250 & n3458 ) | ( ~n3456 & n3458 ) ;
  assign n3460 = n3456 | n3459 ;
  assign n3461 = n578 | n3460 ;
  assign n3462 = n3455 | n3461 ;
  assign n3463 = n219 | n521 ;
  assign n3464 = n648 | n2898 ;
  assign n3465 = n3463 | n3464 ;
  assign n3466 = n240 | n309 ;
  assign n3467 = n3465 | n3466 ;
  assign n3468 = n112 | n602 ;
  assign n3469 = n418 | n3468 ;
  assign n3470 = n187 | n3469 ;
  assign n3471 = n2070 | n3470 ;
  assign n3472 = n3467 | n3471 ;
  assign n3473 = n1314 | n2405 ;
  assign n3474 = n509 | n3473 ;
  assign n3475 = n3472 | n3474 ;
  assign n3476 = n222 | n596 ;
  assign n3477 = n199 | n452 ;
  assign n3478 = n608 | n3477 ;
  assign n3479 = n3476 | n3478 ;
  assign n3480 = n563 | n3479 ;
  assign n3481 = n293 | n499 ;
  assign n3482 = n450 | n3481 ;
  assign n3483 = n143 | n3482 ;
  assign n3484 = n133 | n3483 ;
  assign n3485 = n206 | n3484 ;
  assign n3486 = n3480 | n3485 ;
  assign n3487 = n3475 | n3486 ;
  assign n3488 = n197 | n637 ;
  assign n3489 = n2267 | n3488 ;
  assign n3490 = n83 | n96 ;
  assign n3491 = n100 | n3490 ;
  assign n3492 = n3489 | n3491 ;
  assign n3493 = n108 | n167 ;
  assign n3494 = n3492 | n3493 ;
  assign n3495 = n2722 | n3494 ;
  assign n3496 = n1284 | n3495 ;
  assign n3497 = n3487 | n3496 ;
  assign n3498 = n3462 | n3497 ;
  assign n3499 = n66 | n214 ;
  assign n3500 = n391 | n3499 ;
  assign n3501 = n321 | n3500 ;
  assign n3502 = n172 | n3501 ;
  assign n3503 = n129 | n3502 ;
  assign n3504 = n3498 | n3503 ;
  assign n3505 = ~n3431 & n3504 ;
  assign n3506 = n3431 & ~n3504 ;
  assign n3507 = n3505 | n3506 ;
  assign n3508 = n718 | n1865 ;
  assign n3509 = n3073 | n3508 ;
  assign n3510 = n133 | n207 ;
  assign n3511 = n166 | n3510 ;
  assign n3512 = n436 | n3511 ;
  assign n3513 = n3509 | n3512 ;
  assign n3514 = n1351 | n3513 ;
  assign n3515 = n2411 | n2802 ;
  assign n3516 = n488 | n512 ;
  assign n3517 = n3515 | n3516 ;
  assign n3518 = n274 | n608 ;
  assign n3519 = n110 | n3518 ;
  assign n3520 = n3517 | n3519 ;
  assign n3521 = n248 | n3520 ;
  assign n3522 = n3514 | n3521 ;
  assign n3523 = n888 | n1315 ;
  assign n3524 = n1336 | n3523 ;
  assign n3525 = n127 | n3524 ;
  assign n3526 = n249 | n3525 ;
  assign n3527 = n320 | n3526 ;
  assign n3528 = n3522 | n3527 ;
  assign n3529 = n213 | n282 ;
  assign n3530 = n1354 | n3529 ;
  assign n3531 = n442 | n3530 ;
  assign n3532 = n186 | n191 ;
  assign n3533 = n594 | n3532 ;
  assign n3534 = n3531 | n3533 ;
  assign n3535 = n130 | n1189 ;
  assign n3536 = n377 | n408 ;
  assign n3537 = n180 | n3536 ;
  assign n3538 = n3535 | n3537 ;
  assign n3539 = n132 | n649 ;
  assign n3540 = n3538 | n3539 ;
  assign n3541 = n3534 | n3540 ;
  assign n3542 = n296 | n319 ;
  assign n3543 = n416 | n3542 ;
  assign n3544 = n580 | n3543 ;
  assign n3545 = n3541 | n3544 ;
  assign n3546 = n3528 | n3545 ;
  assign n3547 = n337 | n484 ;
  assign n3548 = n2401 | n3547 ;
  assign n3549 = n252 | n3548 ;
  assign n3550 = n1284 | n1404 ;
  assign n3551 = n500 | n3550 ;
  assign n3552 = n226 & ~n490 ;
  assign n3553 = ~n181 & n3552 ;
  assign n3554 = n1681 | n2898 ;
  assign n3555 = n3553 & ~n3554 ;
  assign n3556 = ~n3551 & n3555 ;
  assign n3557 = ~n3549 & n3556 ;
  assign n3558 = n215 | n307 ;
  assign n3559 = n206 | n476 ;
  assign n3560 = n3558 | n3559 ;
  assign n3561 = n276 | n519 ;
  assign n3562 = n393 | n3561 ;
  assign n3563 = n3560 | n3562 ;
  assign n3564 = n62 | n90 ;
  assign n3565 = n3563 | n3564 ;
  assign n3566 = n808 | n3565 ;
  assign n3567 = n3557 & ~n3566 ;
  assign n3568 = n472 | n626 ;
  assign n3569 = n306 | n3568 ;
  assign n3570 = n155 | n3569 ;
  assign n3571 = n217 | n3570 ;
  assign n3572 = n208 | n3571 ;
  assign n3573 = n3567 & ~n3572 ;
  assign n3574 = ~n2722 & n3573 ;
  assign n3575 = ~n3546 & n3574 ;
  assign n3576 = n279 | n478 ;
  assign n3577 = n112 | n3576 ;
  assign n3578 = n2303 | n3577 ;
  assign n3579 = n531 | n2199 ;
  assign n3580 = n528 | n3579 ;
  assign n3581 = n3578 | n3580 ;
  assign n3582 = n198 | n265 ;
  assign n3583 = n58 | n3582 ;
  assign n3584 = n445 | n3583 ;
  assign n3585 = n3581 | n3584 ;
  assign n3586 = n3217 | n3585 ;
  assign n3587 = n1867 | n3586 ;
  assign n3588 = n3314 | n3587 ;
  assign n3589 = n421 | n3588 ;
  assign n3590 = n3575 & ~n3589 ;
  assign n3591 = n391 | n1022 ;
  assign n3592 = ( n120 & ~n1313 ) | ( n120 & n3591 ) | ( ~n1313 & n3591 ) ;
  assign n3593 = n1313 | n3592 ;
  assign n3594 = n168 | n3593 ;
  assign n3595 = n161 | n3594 ;
  assign n3596 = n3590 & ~n3595 ;
  assign n3597 = n3504 & ~n3596 ;
  assign n3598 = ~n3504 & n3596 ;
  assign n3599 = n3597 | n3598 ;
  assign n3600 = n778 & ~n3596 ;
  assign n3601 = ~n778 & n3596 ;
  assign n3602 = n3600 | n3601 ;
  assign n3603 = n905 & ~n3602 ;
  assign n3604 = n3600 | n3603 ;
  assign n3605 = ~n3599 & n3604 ;
  assign n3606 = n3597 | n3605 ;
  assign n3607 = ~n3507 & n3606 ;
  assign n3608 = n3505 | n3607 ;
  assign n3609 = n3434 & n3608 ;
  assign n3610 = n3432 & ~n3609 ;
  assign n3611 = n3599 | n3601 ;
  assign n3612 = ~n3597 & n3611 ;
  assign n3613 = n3507 | n3612 ;
  assign n3614 = ~n3505 & n3613 ;
  assign n3615 = n3434 & ~n3614 ;
  assign n3616 = n3432 & ~n3615 ;
  assign n3617 = ( ~n3370 & n3610 ) | ( ~n3370 & n3616 ) | ( n3610 & n3616 ) ;
  assign n3618 = n675 & ~n3617 ;
  assign n3619 = n673 & ~n3618 ;
  assign n3620 = ( ~n234 & n466 ) | ( ~n234 & n467 ) | ( n466 & n467 ) ;
  assign n3621 = n459 | n2126 ;
  assign n3622 = n202 | n3621 ;
  assign n3623 = n456 | n3622 ;
  assign n3624 = n571 | n2219 ;
  assign n3625 = n66 | n3624 ;
  assign n3626 = n405 | n3625 ;
  assign n3627 = n400 | n3626 ;
  assign n3628 = n3623 | n3627 ;
  assign n3629 = n364 | n377 ;
  assign n3630 = n586 | n3629 ;
  assign n3631 = n670 | n3630 ;
  assign n3632 = n55 | n3631 ;
  assign n3633 = n3628 | n3632 ;
  assign n3634 = n616 & ~n3633 ;
  assign n3635 = n74 | n235 ;
  assign n3636 = x31 & n3635 ;
  assign n3637 = ~x30 & x31 ;
  assign n3638 = ( x31 & n3635 ) | ( x31 & ~n3637 ) | ( n3635 & ~n3637 ) ;
  assign n3639 = ~n3635 & n3638 ;
  assign n3640 = n3636 | n3639 ;
  assign n3641 = ~n3634 & n3640 ;
  assign n3642 = ~n3620 & n3641 ;
  assign n3643 = ~n467 & n3642 ;
  assign n3644 = n3620 | n3643 ;
  assign n3645 = n672 & n3639 ;
  assign n3646 = ( ~n672 & n3641 ) | ( ~n672 & n3645 ) | ( n3641 & n3645 ) ;
  assign n3647 = ( n3620 & n3644 ) | ( n3620 & n3646 ) | ( n3644 & n3646 ) ;
  assign n3648 = ( ~n3619 & n3644 ) | ( ~n3619 & n3647 ) | ( n3644 & n3647 ) ;
  assign n3649 = n467 | n3648 ;
  assign n3650 = ( ~n3619 & n3641 ) | ( ~n3619 & n3646 ) | ( n3641 & n3646 ) ;
  assign n3651 = ~n3643 & n3650 ;
  assign n3652 = n3649 & ~n3651 ;
  assign n3653 = n203 | n366 ;
  assign n3654 = n408 | n441 ;
  assign n3655 = n3653 | n3654 ;
  assign n3656 = n57 | n484 ;
  assign n3657 = n223 | n3656 ;
  assign n3658 = n291 | n582 ;
  assign n3659 = n301 | n437 ;
  assign n3660 = n3658 | n3659 ;
  assign n3661 = n3657 | n3660 ;
  assign n3662 = n311 | n320 ;
  assign n3663 = n296 | n3662 ;
  assign n3664 = n3661 | n3663 ;
  assign n3665 = n161 | n570 ;
  assign n3666 = n139 | n3665 ;
  assign n3667 = n129 | n3666 ;
  assign n3668 = n3664 | n3667 ;
  assign n3669 = n3655 | n3668 ;
  assign n3670 = n2508 | n3669 ;
  assign n3671 = n2922 | n3670 ;
  assign n3672 = n873 | n2722 ;
  assign n3673 = n210 | n3672 ;
  assign n3674 = n618 | n655 ;
  assign n3675 = n314 | n3674 ;
  assign n3676 = n319 | n3675 ;
  assign n3677 = n3673 | n3676 ;
  assign n3678 = n379 | n579 ;
  assign n3679 = n457 | n3678 ;
  assign n3680 = n111 | n3679 ;
  assign n3681 = n186 | n3680 ;
  assign n3682 = n3677 | n3681 ;
  assign n3683 = n2588 | n3111 ;
  assign n3684 = n157 | n569 ;
  assign n3685 = n190 | n3684 ;
  assign n3686 = n122 | n3685 ;
  assign n3687 = n3683 | n3686 ;
  assign n3688 = n1695 | n3687 ;
  assign n3689 = ( n1350 & n3682 ) | ( n1350 & n3688 ) | ( n3682 & n3688 ) ;
  assign n3690 = n1350 & ~n3689 ;
  assign n3691 = ~n3671 & n3690 ;
  assign n3692 = n1125 | n1417 ;
  assign n3693 = n958 | n3692 ;
  assign n3694 = n421 | n3693 ;
  assign n3695 = n530 | n3694 ;
  assign n3696 = n3691 & ~n3695 ;
  assign n3697 = n468 | n654 ;
  assign n3698 = n300 | n3697 ;
  assign n3699 = n326 | n3698 ;
  assign n3700 = n400 | n3699 ;
  assign n3701 = n81 | n3700 ;
  assign n3702 = n94 | n3701 ;
  assign n3703 = n3696 & ~n3702 ;
  assign n3704 = n221 | n222 ;
  assign n3705 = n1682 | n1954 ;
  assign n3706 = n1423 | n3705 ;
  assign n3707 = n120 | n592 ;
  assign n3708 = n187 | n3707 ;
  assign n3709 = n1260 | n3708 ;
  assign n3710 = n452 | n3709 ;
  assign n3711 = n3706 | n3710 ;
  assign n3712 = n3704 | n3711 ;
  assign n3713 = n526 | n3712 ;
  assign n3714 = n371 | n3713 ;
  assign n3715 = n3406 | n3714 ;
  assign n3716 = n289 | n571 ;
  assign n3717 = n58 | n3716 ;
  assign n3718 = n81 | n3717 ;
  assign n3719 = n129 | n3718 ;
  assign n3720 = n3715 | n3719 ;
  assign n3721 = ( x29 & n3703 ) | ( x29 & ~n3720 ) | ( n3703 & ~n3720 ) ;
  assign n3722 = n466 & ~n3721 ;
  assign n3723 = n672 & ~n3634 ;
  assign n3724 = n672 | n3619 ;
  assign n3725 = n3619 | n3634 ;
  assign n3726 = ( n3723 & ~n3724 ) | ( n3723 & n3725 ) | ( ~n3724 & n3725 ) ;
  assign n3727 = ( x30 & n3637 ) | ( x30 & ~n3638 ) | ( n3637 & ~n3638 ) ;
  assign n3728 = ~n3634 & n3727 ;
  assign n3729 = ( n3639 & ~n3645 ) | ( n3639 & n3728 ) | ( ~n3645 & n3728 ) ;
  assign n3730 = n3636 | n3729 ;
  assign n3731 = ( n3726 & n3729 ) | ( n3726 & n3730 ) | ( n3729 & n3730 ) ;
  assign n3732 = ~n466 & n3721 ;
  assign n3733 = n3722 | n3732 ;
  assign n3734 = n3731 & n3733 ;
  assign n3735 = n3733 & ~n3734 ;
  assign n3736 = ( n3731 & ~n3734 ) | ( n3731 & n3735 ) | ( ~n3734 & n3735 ) ;
  assign n3737 = ( n3722 & n3731 ) | ( n3722 & n3736 ) | ( n3731 & n3736 ) ;
  assign n3738 = ~n3652 & n3737 ;
  assign n3739 = n3652 & ~n3737 ;
  assign n3740 = n3738 | n3739 ;
  assign n3741 = ~n1411 & n3727 ;
  assign n3742 = n3639 | n3741 ;
  assign n3743 = ( n1532 & n3741 ) | ( n1532 & n3742 ) | ( n3741 & n3742 ) ;
  assign n3744 = ~x31 & n3635 ;
  assign n3745 = n3178 & n3744 ;
  assign n3746 = n3743 | n3745 ;
  assign n3747 = n3636 | n3746 ;
  assign n3748 = ( ~n1411 & n3046 ) | ( ~n1411 & n3178 ) | ( n3046 & n3178 ) ;
  assign n3749 = ( n1411 & ~n3178 ) | ( n1411 & n3748 ) | ( ~n3178 & n3748 ) ;
  assign n3750 = ( ~n3046 & n3748 ) | ( ~n3046 & n3749 ) | ( n3748 & n3749 ) ;
  assign n3751 = ( n3746 & n3747 ) | ( n3746 & ~n3750 ) | ( n3747 & ~n3750 ) ;
  assign n3752 = n610 | n626 ;
  assign n3753 = n57 | n3752 ;
  assign n3754 = n799 | n1574 ;
  assign n3755 = n3753 | n3754 ;
  assign n3756 = n337 | n381 ;
  assign n3757 = n249 | n3756 ;
  assign n3758 = n315 | n3757 ;
  assign n3759 = n3755 | n3758 ;
  assign n3760 = n291 | n384 ;
  assign n3761 = n419 | n3760 ;
  assign n3762 = n578 | n3761 ;
  assign n3763 = n203 | n3762 ;
  assign n3764 = n3759 | n3763 ;
  assign n3765 = n601 | n3764 ;
  assign n3766 = n400 | n522 ;
  assign n3767 = n645 | n3766 ;
  assign n3768 = n243 | n2207 ;
  assign n3769 = n3767 | n3768 ;
  assign n3770 = n279 | n519 ;
  assign n3771 = n175 | n3770 ;
  assign n3772 = n3769 | n3771 ;
  assign n3773 = n429 | n607 ;
  assign n3774 = n100 | n3773 ;
  assign n3775 = n270 | n355 ;
  assign n3776 = n253 | n2220 ;
  assign n3777 = n3775 | n3776 ;
  assign n3778 = n3774 | n3777 ;
  assign n3779 = n3772 | n3778 ;
  assign n3780 = n2003 | n2722 ;
  assign n3781 = n3779 | n3780 ;
  assign n3782 = n3765 | n3781 ;
  assign n3783 = n180 | n475 ;
  assign n3784 = n208 | n3783 ;
  assign n3785 = n3074 | n3784 ;
  assign n3786 = n2510 | n3785 ;
  assign n3787 = n46 | n409 ;
  assign n3788 = n1470 | n3787 ;
  assign n3789 = n896 | n3788 ;
  assign n3790 = n3786 | n3789 ;
  assign n3791 = n265 | n344 ;
  assign n3792 = n103 | n3791 ;
  assign n3793 = n433 | n3792 ;
  assign n3794 = n530 | n3793 ;
  assign n3795 = n514 | n3794 ;
  assign n3796 = n3790 | n3795 ;
  assign n3797 = n309 | n314 ;
  assign n3798 = n134 | n3797 ;
  assign n3799 = n404 | n3798 ;
  assign n3800 = n167 | n3799 ;
  assign n3801 = n3796 | n3800 ;
  assign n3802 = n3782 | n3801 ;
  assign n3803 = n207 | n227 ;
  assign n3804 = n911 | n1852 ;
  assign n3805 = n132 | n3804 ;
  assign n3806 = ( n378 & ~n2396 ) | ( n378 & n3805 ) | ( ~n2396 & n3805 ) ;
  assign n3807 = n2396 | n3806 ;
  assign n3808 = n3803 | n3807 ;
  assign n3809 = n299 | n498 ;
  assign n3810 = n3218 | n3809 ;
  assign n3811 = n244 | n321 ;
  assign n3812 = n582 | n3811 ;
  assign n3813 = n3810 | n3812 ;
  assign n3814 = n206 | n3813 ;
  assign n3815 = n334 | n509 ;
  assign n3816 = n65 | n296 ;
  assign n3817 = n3815 | n3816 ;
  assign n3818 = n142 | n403 ;
  assign n3819 = n3817 | n3818 ;
  assign n3820 = n1847 | n2643 ;
  assign n3821 = n3819 | n3820 ;
  assign n3822 = n3814 | n3821 ;
  assign n3823 = n3808 | n3822 ;
  assign n3824 = n1057 | n1867 ;
  assign n3825 = n1522 | n3824 ;
  assign n3826 = n619 | n3825 ;
  assign n3827 = n320 | n3826 ;
  assign n3828 = n307 | n3827 ;
  assign n3829 = n3823 | n3828 ;
  assign n3830 = n356 | n434 ;
  assign n3831 = n90 | n3830 ;
  assign n3832 = n85 | n3831 ;
  assign n3833 = n3829 | n3832 ;
  assign n3834 = n3802 | n3833 ;
  assign n3835 = n1336 | n3314 ;
  assign n3836 = n240 | n3835 ;
  assign n3837 = n62 | n3836 ;
  assign n3838 = n172 | n3837 ;
  assign n3839 = n94 | n3838 ;
  assign n3840 = n186 | n3839 ;
  assign n3841 = n647 | n3840 ;
  assign n3842 = n3834 | n3841 ;
  assign n3843 = n145 | n167 ;
  assign n3844 = n815 | n3843 ;
  assign n3845 = n278 | n1220 ;
  assign n3846 = n227 | n2199 ;
  assign n3847 = n3845 | n3846 ;
  assign n3848 = n3844 | n3847 ;
  assign n3849 = n3247 | n3848 ;
  assign n3850 = n319 | n451 ;
  assign n3851 = n1316 | n1404 ;
  assign n3852 = n219 | n3851 ;
  assign n3853 = n3850 | n3852 ;
  assign n3854 = n2154 | n3853 ;
  assign n3855 = n3849 | n3854 ;
  assign n3856 = n315 | n345 ;
  assign n3857 = n430 | n3856 ;
  assign n3858 = n242 | n3857 ;
  assign n3859 = n596 | n3858 ;
  assign n3860 = n364 | n3859 ;
  assign n3861 = n174 | n3860 ;
  assign n3862 = n3855 | n3861 ;
  assign n3863 = n727 | n3862 ;
  assign n3864 = n129 | n356 ;
  assign n3865 = n66 | n3864 ;
  assign n3866 = n355 | n3865 ;
  assign n3867 = n197 | n253 ;
  assign n3868 = n204 | n223 ;
  assign n3869 = n3867 | n3868 ;
  assign n3870 = n1921 | n3869 ;
  assign n3871 = n3866 | n3870 ;
  assign n3872 = n2960 | n3871 ;
  assign n3873 = n300 | n510 ;
  assign n3874 = n114 | n2534 ;
  assign n3875 = n484 | n1985 ;
  assign n3876 = n3874 | n3875 ;
  assign n3877 = n483 | n504 ;
  assign n3878 = n270 | n3877 ;
  assign n3879 = n96 | n3878 ;
  assign n3880 = n3876 | n3879 ;
  assign n3881 = n3873 | n3880 ;
  assign n3882 = n3872 | n3881 ;
  assign n3883 = n922 | n1280 ;
  assign n3884 = n1989 | n3883 ;
  assign n3885 = n478 | n3884 ;
  assign n3886 = n509 | n3885 ;
  assign n3887 = n3882 | n3886 ;
  assign n3888 = n499 | n653 ;
  assign n3889 = n498 | n3888 ;
  assign n3890 = n346 | n3889 ;
  assign n3891 = n608 | n3890 ;
  assign n3892 = n601 | n3891 ;
  assign n3893 = n3887 | n3892 ;
  assign n3894 = n125 | n514 ;
  assign n3895 = n2355 | n3894 ;
  assign n3896 = n94 | n3895 ;
  assign n3897 = n2481 | n2628 ;
  assign n3898 = n3896 | n3897 ;
  assign n3899 = n352 | n862 ;
  assign n3900 = n373 | n3899 ;
  assign n3901 = n292 | n3900 ;
  assign n3902 = n3898 | n3901 ;
  assign n3903 = n293 | n579 ;
  assign n3904 = n445 | n570 ;
  assign n3905 = ( ~n1805 & n3903 ) | ( ~n1805 & n3904 ) | ( n3903 & n3904 ) ;
  assign n3906 = n1805 | n3905 ;
  assign n3907 = ( ~n3893 & n3902 ) | ( ~n3893 & n3906 ) | ( n3902 & n3906 ) ;
  assign n3908 = n3893 | n3907 ;
  assign n3909 = n3863 | n3908 ;
  assign n3910 = n309 | n540 ;
  assign n3911 = n337 | n472 ;
  assign n3912 = n3910 | n3911 ;
  assign n3913 = n500 | n669 ;
  assign n3914 = n450 | n3913 ;
  assign n3915 = n3912 | n3914 ;
  assign n3916 = n128 | n3915 ;
  assign n3917 = n861 | n3916 ;
  assign n3918 = n1311 | n3917 ;
  assign n3919 = n2433 | n3918 ;
  assign n3920 = n245 | n3919 ;
  assign n3921 = n359 | n3920 ;
  assign n3922 = n3909 | n3921 ;
  assign n3923 = n194 | n215 ;
  assign n3924 = n57 | n3923 ;
  assign n3925 = n76 | n3924 ;
  assign n3926 = n133 | n3925 ;
  assign n3927 = n3922 | n3926 ;
  assign n3928 = ~n3842 & n3927 ;
  assign n3929 = n1535 & ~n3044 ;
  assign n3930 = n3045 | n3929 ;
  assign n3931 = n3842 & ~n3927 ;
  assign n3932 = n1532 & n3727 ;
  assign n3933 = ~n1411 & n3744 ;
  assign n3934 = ~n2939 & n3639 ;
  assign n3935 = n3933 | n3934 ;
  assign n3936 = n3932 | n3935 ;
  assign n3937 = n3636 | n3936 ;
  assign n3938 = ~n3928 & n3937 ;
  assign n3939 = ~n3931 & n3938 ;
  assign n3940 = ~n3928 & n3936 ;
  assign n3941 = ~n3931 & n3940 ;
  assign n3942 = ( ~n3930 & n3939 ) | ( ~n3930 & n3941 ) | ( n3939 & n3941 ) ;
  assign n3943 = n3928 | n3942 ;
  assign n3944 = n1272 | n2179 ;
  assign n3945 = n364 | n450 ;
  assign n3946 = n3204 | n3945 ;
  assign n3947 = n3944 | n3946 ;
  assign n3948 = n374 | n2688 ;
  assign n3949 = n3864 | n3948 ;
  assign n3950 = n3947 | n3949 ;
  assign n3951 = n242 | n540 ;
  assign n3952 = n327 | n3951 ;
  assign n3953 = n3950 | n3952 ;
  assign n3954 = n142 | n579 ;
  assign n3955 = n2434 | n3954 ;
  assign n3956 = n1430 | n2960 ;
  assign n3957 = ( ~n3953 & n3955 ) | ( ~n3953 & n3956 ) | ( n3955 & n3956 ) ;
  assign n3958 = n3953 | n3957 ;
  assign n3959 = n3585 | n3958 ;
  assign n3960 = n490 | n2169 ;
  assign n3961 = n335 | n3960 ;
  assign n3962 = n307 | n3961 ;
  assign n3963 = n670 | n3962 ;
  assign n3964 = n444 | n3963 ;
  assign n3965 = n3959 | n3964 ;
  assign n3966 = n92 | n133 ;
  assign n3967 = n223 | n3966 ;
  assign n3968 = n3965 | n3967 ;
  assign n3969 = n355 | n505 ;
  assign n3970 = n127 | n3969 ;
  assign n3971 = n204 | n590 ;
  assign n3972 = n434 | n3971 ;
  assign n3973 = n3970 | n3972 ;
  assign n3974 = n102 | n1064 ;
  assign n3975 = n3973 | n3974 ;
  assign n3976 = n857 | n2270 ;
  assign n3977 = n3975 | n3976 ;
  assign n3978 = n169 | n731 ;
  assign n3979 = n421 | n3978 ;
  assign n3980 = n648 | n3979 ;
  assign n3981 = n245 | n3980 ;
  assign n3982 = n3977 | n3981 ;
  assign n3983 = n625 | n634 ;
  assign n3984 = n519 | n3983 ;
  assign n3985 = n315 | n3984 ;
  assign n3986 = n241 | n3985 ;
  assign n3987 = n260 | n3986 ;
  assign n3988 = n55 | n3987 ;
  assign n3989 = n3982 | n3988 ;
  assign n3990 = n103 | n442 ;
  assign n3991 = n192 | n1513 ;
  assign n3992 = n3508 | n3991 ;
  assign n3993 = n439 | n3062 ;
  assign n3994 = n3992 | n3993 ;
  assign n3995 = n3990 | n3994 ;
  assign n3996 = n3989 | n3995 ;
  assign n3997 = n3968 | n3996 ;
  assign n3998 = n276 | n655 ;
  assign n3999 = n207 | n3998 ;
  assign n4000 = ( n431 & ~n1641 ) | ( n431 & n3999 ) | ( ~n1641 & n3999 ) ;
  assign n4001 = n1641 | n4000 ;
  assign n4002 = n640 | n4001 ;
  assign n4003 = n1360 | n2232 ;
  assign n4004 = n52 | n484 ;
  assign n4005 = n2867 | n4004 ;
  assign n4006 = n618 | n4005 ;
  assign n4007 = n4003 | n4006 ;
  assign n4008 = n277 | n639 ;
  assign n4009 = n262 | n4008 ;
  assign n4010 = n310 | n4009 ;
  assign n4011 = n226 & ~n4010 ;
  assign n4012 = ~n4007 & n4011 ;
  assign n4013 = ~n4002 & n4012 ;
  assign n4014 = ~n1054 & n4013 ;
  assign n4015 = ~n2635 & n4014 ;
  assign n4016 = ~n1443 & n4015 ;
  assign n4017 = ~n3997 & n4016 ;
  assign n4018 = n475 | n483 ;
  assign n4019 = n510 | n4018 ;
  assign n4020 = n393 | n4019 ;
  assign n4021 = n152 | n4020 ;
  assign n4022 = n4017 & ~n4021 ;
  assign n4023 = ( x14 & ~n3842 ) | ( x14 & n4022 ) | ( ~n3842 & n4022 ) ;
  assign n4024 = ( ~x14 & n3842 ) | ( ~x14 & n4023 ) | ( n3842 & n4023 ) ;
  assign n4025 = ( ~n4022 & n4023 ) | ( ~n4022 & n4024 ) | ( n4023 & n4024 ) ;
  assign n4026 = n3943 & n4025 ;
  assign n4027 = n3943 | n4025 ;
  assign n4028 = ~n4026 & n4027 ;
  assign n4029 = n3751 & n4028 ;
  assign n4030 = n4028 & ~n4029 ;
  assign n4031 = ( n3751 & ~n4029 ) | ( n3751 & n4030 ) | ( ~n4029 & n4030 ) ;
  assign n4032 = ( n3046 & n3186 ) | ( n3046 & n3192 ) | ( n3186 & n3192 ) ;
  assign n4033 = n3048 & ~n4032 ;
  assign n4034 = n3194 | n4033 ;
  assign n4035 = n43 & ~n50 ;
  assign n4036 = x28 & ~x29 ;
  assign n4037 = ~x28 & x29 ;
  assign n4038 = n4036 | n4037 ;
  assign n4039 = x26 & ~x27 ;
  assign n4040 = ~x26 & x27 ;
  assign n4041 = n4039 | n4040 ;
  assign n4042 = n4038 & ~n4041 ;
  assign n4043 = ~n4035 & n4042 ;
  assign n4044 = n3104 & n4043 ;
  assign n4045 = n4035 & ~n4041 ;
  assign n4046 = n1327 & n4045 ;
  assign n4047 = n4044 | n4046 ;
  assign n4048 = ~n4038 & n4041 ;
  assign n4049 = ~n1151 & n4048 ;
  assign n4050 = n4047 | n4049 ;
  assign n4051 = n4038 & n4041 ;
  assign n4052 = n4050 | n4051 ;
  assign n4053 = ( ~n4034 & n4050 ) | ( ~n4034 & n4052 ) | ( n4050 & n4052 ) ;
  assign n4054 = ~x29 & n4053 ;
  assign n4055 = x29 | n4054 ;
  assign n4056 = ( ~n4053 & n4054 ) | ( ~n4053 & n4055 ) | ( n4054 & n4055 ) ;
  assign n4057 = n4031 & n4056 ;
  assign n4058 = n4031 & ~n4057 ;
  assign n4059 = ~n4031 & n4056 ;
  assign n4060 = n4058 | n4059 ;
  assign n4061 = ( ~n3930 & n3936 ) | ( ~n3930 & n3937 ) | ( n3936 & n3937 ) ;
  assign n4062 = ~n3942 & n4061 ;
  assign n4064 = n638 | n2362 ;
  assign n4065 = n488 | n1024 ;
  assign n4066 = n4064 | n4065 ;
  assign n4067 = n114 | n274 ;
  assign n4068 = n126 | n4067 ;
  assign n4069 = n265 | n482 ;
  assign n4070 = n57 | n4069 ;
  assign n4071 = n4068 | n4070 ;
  assign n4072 = n4066 | n4071 ;
  assign n4073 = n3658 | n4072 ;
  assign n4074 = n1583 | n3772 ;
  assign n4075 = n4073 | n4074 ;
  assign n4076 = n971 | n4075 ;
  assign n4077 = n273 | n450 ;
  assign n4078 = n4004 | n4077 ;
  assign n4079 = n2586 | n4078 ;
  assign n4080 = n3375 | n3532 ;
  assign n4081 = n336 | n4080 ;
  assign n4082 = n4079 | n4081 ;
  assign n4083 = n320 | n1522 ;
  assign n4084 = n417 | n4083 ;
  assign n4085 = n364 | n4084 ;
  assign n4086 = n4082 | n4085 ;
  assign n4087 = n142 | n377 ;
  assign n4088 = n4086 | n4087 ;
  assign n4089 = n249 | n489 ;
  assign n4090 = n1657 | n4089 ;
  assign n4091 = n408 | n602 ;
  assign n4092 = n143 | n4091 ;
  assign n4093 = n4090 | n4092 ;
  assign n4094 = n122 | n4093 ;
  assign n4095 = n1464 | n2818 ;
  assign n4096 = n366 | n403 ;
  assign n4097 = n161 | n4096 ;
  assign n4098 = n1023 | n4097 ;
  assign n4099 = n4095 | n4098 ;
  assign n4100 = n4094 | n4099 ;
  assign n4101 = n521 | n578 ;
  assign n4102 = n337 | n4101 ;
  assign n4103 = n626 | n4102 ;
  assign n4104 = n520 | n4103 ;
  assign n4105 = n321 | n4104 ;
  assign n4106 = n4100 | n4105 ;
  assign n4107 = n292 | n344 ;
  assign n4108 = n62 | n4107 ;
  assign n4109 = n650 | n4108 ;
  assign n4110 = n4106 | n4109 ;
  assign n4111 = n4088 | n4110 ;
  assign n4112 = n4076 | n4111 ;
  assign n4113 = n244 | n283 ;
  assign n4114 = n92 | n4113 ;
  assign n4115 = n640 | n4114 ;
  assign n4116 = n4112 | n4115 ;
  assign n4117 = n1183 | n1647 ;
  assign n4118 = n2474 | n3910 ;
  assign n4119 = n519 | n528 ;
  assign n4120 = n57 | n640 ;
  assign n4121 = n4119 | n4120 ;
  assign n4122 = n4118 | n4121 ;
  assign n4123 = n296 | n2419 ;
  assign n4124 = n4122 | n4123 ;
  assign n4125 = n346 | n452 ;
  assign n4126 = n4124 | n4125 ;
  assign n4127 = n468 | n505 ;
  assign n4128 = n321 | n4127 ;
  assign n4129 = n1423 | n3707 ;
  assign n4130 = ( ~n4126 & n4128 ) | ( ~n4126 & n4129 ) | ( n4128 & n4129 ) ;
  assign n4131 = n4126 | n4130 ;
  assign n4132 = n4117 | n4131 ;
  assign n4133 = n635 | n1659 ;
  assign n4134 = n2867 | n4133 ;
  assign n4135 = n472 | n4134 ;
  assign n4136 = n242 | n4135 ;
  assign n4137 = n628 | n4136 ;
  assign n4138 = n4132 | n4137 ;
  assign n4139 = n510 | n513 ;
  assign n4140 = n437 | n4139 ;
  assign n4141 = n458 | n4140 ;
  assign n4142 = n122 | n4141 ;
  assign n4143 = n4138 | n4142 ;
  assign n4144 = n928 | n2893 ;
  assign n4145 = n841 | n3850 ;
  assign n4146 = n4144 | n4145 ;
  assign n4147 = n482 | n618 ;
  assign n4148 = n470 | n4147 ;
  assign n4149 = n338 | n4148 ;
  assign n4150 = n383 | n4149 ;
  assign n4151 = n4146 | n4150 ;
  assign n4152 = n1756 | n3123 ;
  assign n4153 = n212 | n344 ;
  assign n4154 = n132 | n4153 ;
  assign n4155 = n645 | n4154 ;
  assign n4156 = n4152 | n4155 ;
  assign n4157 = n1066 | n4156 ;
  assign n4158 = n4151 | n4157 ;
  assign n4159 = n277 | n601 ;
  assign n4160 = n99 | n4159 ;
  assign n4161 = n857 | n1118 ;
  assign n4162 = n4160 | n4161 ;
  assign n4163 = n431 | n626 ;
  assign n4164 = n669 | n4163 ;
  assign n4165 = n292 | n4164 ;
  assign n4166 = n4162 | n4165 ;
  assign n4167 = n146 | n3971 ;
  assign n4168 = n4166 | n4167 ;
  assign n4169 = n1023 | n4168 ;
  assign n4170 = n4158 | n4169 ;
  assign n4171 = n446 | n3655 ;
  assign n4172 = n4170 | n4171 ;
  assign n4173 = n4143 | n4172 ;
  assign n4174 = n990 | n4088 ;
  assign n4175 = n718 | n4174 ;
  assign n4176 = n834 | n4175 ;
  assign n4177 = n4173 | n4176 ;
  assign n4178 = n258 | n619 ;
  assign n4179 = n315 | n4178 ;
  assign n4180 = n596 | n4179 ;
  assign n4181 = n65 | n4180 ;
  assign n4182 = n434 | n4181 ;
  assign n4183 = n100 | n4182 ;
  assign n4184 = n217 | n4183 ;
  assign n4185 = n649 | n4184 ;
  assign n4186 = n4177 | n4185 ;
  assign n4187 = ( x11 & ~n4116 ) | ( x11 & n4186 ) | ( ~n4116 & n4186 ) ;
  assign n4188 = ( ~x11 & n4116 ) | ( ~x11 & n4187 ) | ( n4116 & n4187 ) ;
  assign n4189 = ~n3842 & n4188 ;
  assign n4190 = ( ~n2888 & n3037 ) | ( ~n2888 & n3042 ) | ( n3037 & n3042 ) ;
  assign n4191 = ( ~n2888 & n3036 ) | ( ~n2888 & n3041 ) | ( n3036 & n3041 ) ;
  assign n4192 = n2942 & ~n4191 ;
  assign n4193 = n4190 | n4192 ;
  assign n4194 = n1532 & n3744 ;
  assign n4195 = n3030 & n3639 ;
  assign n4196 = ~n2939 & n3727 ;
  assign n4197 = n4195 | n4196 ;
  assign n4198 = n4194 | n4197 ;
  assign n4199 = n3636 | n4198 ;
  assign n4200 = ( ~n4193 & n4198 ) | ( ~n4193 & n4199 ) | ( n4198 & n4199 ) ;
  assign n4201 = n3842 & ~n4188 ;
  assign n4202 = n4189 | n4201 ;
  assign n4203 = n4200 & n4202 ;
  assign n4204 = n4202 & ~n4203 ;
  assign n4205 = ( n4200 & ~n4203 ) | ( n4200 & n4204 ) | ( ~n4203 & n4204 ) ;
  assign n4206 = ( n4189 & n4200 ) | ( n4189 & n4205 ) | ( n4200 & n4205 ) ;
  assign n4063 = n3931 | n3943 ;
  assign n4207 = ~n4063 & n4206 ;
  assign n4208 = ( n4062 & n4206 ) | ( n4062 & n4207 ) | ( n4206 & n4207 ) ;
  assign n4209 = n4063 & ~n4206 ;
  assign n4210 = ~n4062 & n4209 ;
  assign n4211 = n4208 | n4210 ;
  assign n4212 = ( ~n2888 & n3035 ) | ( ~n2888 & n3040 ) | ( n3035 & n3040 ) ;
  assign n4213 = ( n1625 & ~n2888 ) | ( n1625 & n3030 ) | ( ~n2888 & n3030 ) ;
  assign n4214 = n3034 & ~n4213 ;
  assign n4215 = n4212 | n4214 ;
  assign n4216 = ~n2939 & n3744 ;
  assign n4217 = n3030 & n3727 ;
  assign n4218 = n1625 & n3639 ;
  assign n4219 = n4217 | n4218 ;
  assign n4220 = n4216 | n4219 ;
  assign n4221 = n3636 | n4220 ;
  assign n4222 = ( ~n4215 & n4220 ) | ( ~n4215 & n4221 ) | ( n4220 & n4221 ) ;
  assign n4223 = ( ~n4186 & n4187 ) | ( ~n4186 & n4188 ) | ( n4187 & n4188 ) ;
  assign n4224 = n4222 & ~n4223 ;
  assign n4225 = n390 | n438 ;
  assign n4226 = n93 | n4225 ;
  assign n4227 = n636 | n653 ;
  assign n4228 = n350 | n4227 ;
  assign n4229 = n4226 | n4228 ;
  assign n4230 = n187 | n194 ;
  assign n4231 = n4229 | n4230 ;
  assign n4232 = n260 | n503 ;
  assign n4233 = n1337 | n4232 ;
  assign n4234 = n167 | n197 ;
  assign n4235 = n4233 | n4234 ;
  assign n4236 = n206 | n661 ;
  assign n4237 = n2950 | n4236 ;
  assign n4238 = n174 | n521 ;
  assign n4239 = n731 | n4238 ;
  assign n4240 = n4237 | n4239 ;
  assign n4241 = n1294 | n4240 ;
  assign n4242 = n4235 | n4241 ;
  assign n4243 = n1608 | n4242 ;
  assign n4244 = n4231 | n4243 ;
  assign n4245 = n1592 | n4244 ;
  assign n4246 = n1543 | n1866 ;
  assign n4247 = n2410 | n4246 ;
  assign n4248 = n4245 | n4247 ;
  assign n4249 = n1140 | n4248 ;
  assign n4250 = n266 | n488 ;
  assign n4251 = n292 | n4250 ;
  assign n4252 = n366 | n4251 ;
  assign n4253 = n52 | n4252 ;
  assign n4254 = n213 | n4253 ;
  assign n4255 = n143 | n4254 ;
  assign n4256 = n4249 | n4255 ;
  assign n4257 = ~n4116 & n4256 ;
  assign n4258 = n4116 & ~n4256 ;
  assign n4259 = n1736 & n2886 ;
  assign n4260 = n2887 & ~n4259 ;
  assign n4261 = n308 | n844 ;
  assign n4262 = n3753 | n4261 ;
  assign n4263 = n1750 | n4262 ;
  assign n4264 = n1368 | n4263 ;
  assign n4265 = n52 | n419 ;
  assign n4266 = n204 | n4265 ;
  assign n4267 = n2123 | n4266 ;
  assign n4268 = n165 | n442 ;
  assign n4269 = n145 | n4268 ;
  assign n4270 = n4267 | n4269 ;
  assign n4271 = n432 | n528 ;
  assign n4272 = n498 | n4271 ;
  assign n4273 = n222 | n350 ;
  assign n4274 = n227 | n4273 ;
  assign n4275 = n475 | n4274 ;
  assign n4276 = n4272 | n4275 ;
  assign n4277 = n194 | n597 ;
  assign n4278 = n226 & ~n4277 ;
  assign n4279 = ~n224 & n4278 ;
  assign n4280 = ~n4276 & n4279 ;
  assign n4281 = ~n4270 & n4280 ;
  assign n4282 = ~n4264 & n4281 ;
  assign n4283 = n529 | n637 ;
  assign n4284 = n252 | n4283 ;
  assign n4285 = n569 | n4284 ;
  assign n4286 = n451 | n4285 ;
  assign n4287 = n111 | n4286 ;
  assign n4288 = n160 | n4287 ;
  assign n4289 = n4282 & ~n4288 ;
  assign n4290 = n83 | n187 ;
  assign n4291 = n1166 | n4128 ;
  assign n4292 = n2831 | n4291 ;
  assign n4293 = n275 | n1692 ;
  assign n4294 = n618 | n639 ;
  assign n4295 = n338 | n4294 ;
  assign n4296 = n4293 | n4295 ;
  assign n4297 = n122 | n309 ;
  assign n4298 = n4296 | n4297 ;
  assign n4299 = n4292 | n4298 ;
  assign n4300 = n415 | n4299 ;
  assign n4301 = n4290 | n4300 ;
  assign n4302 = n4289 & ~n4301 ;
  assign n4303 = n242 | n391 ;
  assign n4304 = n596 | n4303 ;
  assign n4305 = n373 | n2305 ;
  assign n4306 = n4304 | n4305 ;
  assign n4307 = n349 | n4306 ;
  assign n4308 = n358 | n669 ;
  assign n4309 = n1371 | n4308 ;
  assign n4310 = n2149 | n4309 ;
  assign n4311 = n1240 | n4310 ;
  assign n4312 = n4002 | n4311 ;
  assign n4313 = n1078 | n1811 ;
  assign n4314 = n635 | n4313 ;
  assign n4315 = n4101 | n4314 ;
  assign n4316 = n263 | n4315 ;
  assign n4317 = n4312 | n4316 ;
  assign n4318 = n291 | n319 ;
  assign n4319 = n420 | n4318 ;
  assign n4320 = n444 | n4319 ;
  assign n4321 = n90 | n4320 ;
  assign n4322 = n77 | n4321 ;
  assign n4323 = n168 | n4322 ;
  assign n4324 = n4317 | n4323 ;
  assign n4325 = n4307 | n4324 ;
  assign n4326 = n4302 & ~n4325 ;
  assign n4327 = n283 | n621 ;
  assign n4328 = n499 | n4327 ;
  assign n4329 = ( n92 & ~n3582 ) | ( n92 & n4328 ) | ( ~n3582 & n4328 ) ;
  assign n4330 = n3582 | n4329 ;
  assign n4331 = n128 | n4330 ;
  assign n4332 = n217 | n4331 ;
  assign n4333 = n649 | n4332 ;
  assign n4334 = n4326 & ~n4333 ;
  assign n4335 = n102 | n3973 ;
  assign n4336 = n345 | n610 ;
  assign n4337 = n152 | n4336 ;
  assign n4338 = n871 | n4337 ;
  assign n4339 = n2950 | n4338 ;
  assign n4340 = n4335 | n4339 ;
  assign n4341 = n431 | n653 ;
  assign n4342 = n280 | n513 ;
  assign n4343 = n4341 | n4342 ;
  assign n4344 = n309 | n338 ;
  assign n4345 = n420 | n4344 ;
  assign n4346 = n4343 | n4345 ;
  assign n4347 = n81 | n661 ;
  assign n4348 = n4346 | n4347 ;
  assign n4349 = n756 | n4348 ;
  assign n4350 = n4340 | n4349 ;
  assign n4351 = n141 | n1311 ;
  assign n4352 = n1115 | n4351 ;
  assign n4353 = n1261 | n4352 ;
  assign n4354 = n445 | n4353 ;
  assign n4355 = n155 | n4354 ;
  assign n4356 = n4350 | n4355 ;
  assign n4357 = n245 | n337 ;
  assign n4358 = n284 | n4357 ;
  assign n4359 = n364 | n619 ;
  assign n4360 = n110 | n4359 ;
  assign n4361 = n4358 | n4360 ;
  assign n4362 = n103 | n167 ;
  assign n4363 = n146 | n4362 ;
  assign n4364 = n4361 | n4363 ;
  assign n4365 = n128 | n629 ;
  assign n4366 = n216 | n633 ;
  assign n4367 = n4365 | n4366 ;
  assign n4368 = n2538 | n4367 ;
  assign n4369 = n650 | n4368 ;
  assign n4370 = n4364 | n4369 ;
  assign n4371 = n555 | n4370 ;
  assign n4372 = n4356 | n4371 ;
  assign n4373 = n1576 | n2401 ;
  assign n4374 = n59 | n1434 ;
  assign n4375 = n4373 | n4374 ;
  assign n4376 = n260 | n530 ;
  assign n4377 = n320 | n4376 ;
  assign n4378 = n358 | n4377 ;
  assign n4379 = n4375 | n4378 ;
  assign n4380 = n379 | n458 ;
  assign n4381 = n172 | n4380 ;
  assign n4382 = n4379 | n4381 ;
  assign n4383 = n3217 | n4382 ;
  assign n4384 = n641 | n4383 ;
  assign n4385 = n857 | n4384 ;
  assign n4386 = n4372 | n4385 ;
  assign n4387 = n996 | n1284 ;
  assign n4388 = n647 | n2973 ;
  assign n4389 = n4387 | n4388 ;
  assign n4390 = n223 | n4389 ;
  assign n4391 = n1371 | n1959 ;
  assign n4392 = n120 | n4391 ;
  assign n4393 = n206 | n274 ;
  assign n4394 = n93 | n4393 ;
  assign n4395 = n844 | n4394 ;
  assign n4396 = n4392 | n4395 ;
  assign n4397 = n4390 | n4396 ;
  assign n4398 = n2306 | n3476 ;
  assign n4399 = n489 | n807 ;
  assign n4400 = n4398 | n4399 ;
  assign n4401 = n503 | n3983 ;
  assign n4402 = n293 | n4401 ;
  assign n4403 = n4400 | n4402 ;
  assign n4404 = n160 | n608 ;
  assign n4405 = n227 | n4404 ;
  assign n4406 = n4403 | n4405 ;
  assign n4407 = n4397 | n4406 ;
  assign n4408 = n1314 | n1315 ;
  assign n4409 = n2219 | n4408 ;
  assign n4410 = n1613 | n4409 ;
  assign n4411 = n1170 | n4410 ;
  assign n4412 = n4407 | n4411 ;
  assign n4413 = n484 | n654 ;
  assign n4414 = ( n449 & ~n3103 ) | ( n449 & n4413 ) | ( ~n3103 & n4413 ) ;
  assign n4415 = n3103 | n4414 ;
  assign n4416 = n161 | n4415 ;
  assign n4417 = n4412 | n4416 ;
  assign n4418 = n3243 | n4417 ;
  assign n4419 = n4386 | n4418 ;
  assign n4420 = n321 | n510 ;
  assign n4421 = n366 | n4420 ;
  assign n4422 = n670 | n4421 ;
  assign n4423 = n607 | n4422 ;
  assign n4424 = n649 | n4423 ;
  assign n4425 = n4419 | n4424 ;
  assign n4426 = ( x8 & n4334 ) | ( x8 & ~n4425 ) | ( n4334 & ~n4425 ) ;
  assign n4427 = n4116 & n4426 ;
  assign n4428 = ~n2873 & n3639 ;
  assign n4429 = ~n1733 & n3727 ;
  assign n4430 = n4428 | n4429 ;
  assign n4431 = n1625 & n3744 ;
  assign n4432 = n4430 | n4431 ;
  assign n4433 = ( n4116 & n4426 ) | ( n4116 & ~n4432 ) | ( n4426 & ~n4432 ) ;
  assign n4434 = ( ~n3636 & n4427 ) | ( ~n3636 & n4433 ) | ( n4427 & n4433 ) ;
  assign n4435 = n4257 | n4434 ;
  assign n4436 = n4257 | n4433 ;
  assign n4437 = ( ~n4260 & n4435 ) | ( ~n4260 & n4436 ) | ( n4435 & n4436 ) ;
  assign n4438 = n4258 | n4437 ;
  assign n4439 = ~n4257 & n4438 ;
  assign n4440 = ~n4222 & n4223 ;
  assign n4441 = n4224 | n4440 ;
  assign n4442 = n4439 | n4441 ;
  assign n4443 = ~n4224 & n4442 ;
  assign n4444 = n4205 | n4443 ;
  assign n4445 = n4205 & n4443 ;
  assign n4446 = n4444 & ~n4445 ;
  assign n4447 = ( n3046 & n3183 ) | ( n3046 & n3189 ) | ( n3183 & n3189 ) ;
  assign n4448 = n3182 | n3748 ;
  assign n4449 = ~n4447 & n4448 ;
  assign n4450 = ~n1411 & n4043 ;
  assign n4451 = n3178 & n4045 ;
  assign n4452 = n4450 | n4451 ;
  assign n4453 = n3104 & n4048 ;
  assign n4454 = n4452 | n4453 ;
  assign n4455 = n4051 | n4454 ;
  assign n4456 = ( n4449 & n4454 ) | ( n4449 & n4455 ) | ( n4454 & n4455 ) ;
  assign n4457 = x29 & n4456 ;
  assign n4458 = x29 & ~n4457 ;
  assign n4459 = ( n4456 & ~n4457 ) | ( n4456 & n4458 ) | ( ~n4457 & n4458 ) ;
  assign n4460 = n4446 & n4459 ;
  assign n4461 = n4444 & ~n4460 ;
  assign n4462 = n4211 | n4461 ;
  assign n4463 = ~n4208 & n4462 ;
  assign n4464 = n4060 & ~n4463 ;
  assign n4465 = ~n4060 & n4463 ;
  assign n4466 = n4464 | n4465 ;
  assign n4467 = ( n3196 & n3358 ) | ( n3196 & n3363 ) | ( n3358 & n3363 ) ;
  assign n4468 = ( n3196 & n3354 ) | ( n3196 & n3357 ) | ( n3354 & n3357 ) ;
  assign n4469 = n3352 & ~n4468 ;
  assign n4470 = n4467 | n4469 ;
  assign n4471 = ~n41 & n48 ;
  assign n4472 = x23 & ~x24 ;
  assign n4473 = ~x23 & x24 ;
  assign n4474 = n4472 | n4473 ;
  assign n4475 = x25 & ~x26 ;
  assign n4476 = ~x25 & x26 ;
  assign n4477 = n4475 | n4476 ;
  assign n4478 = ~n4474 & n4477 ;
  assign n4479 = ~n4471 & n4478 ;
  assign n4480 = n1233 & n4479 ;
  assign n4481 = n4471 & ~n4474 ;
  assign n4482 = n3349 & n4481 ;
  assign n4483 = n4480 | n4482 ;
  assign n4484 = n4474 & ~n4477 ;
  assign n4485 = ~n3255 & n4484 ;
  assign n4486 = n4483 | n4485 ;
  assign n4487 = n4474 & n4477 ;
  assign n4488 = n4486 | n4487 ;
  assign n4489 = ( ~n4470 & n4486 ) | ( ~n4470 & n4488 ) | ( n4486 & n4488 ) ;
  assign n4490 = ~x26 & n4489 ;
  assign n4491 = x26 | n4490 ;
  assign n4492 = ( ~n4489 & n4490 ) | ( ~n4489 & n4491 ) | ( n4490 & n4491 ) ;
  assign n4493 = ~n4466 & n4492 ;
  assign n4494 = n4466 & ~n4492 ;
  assign n4495 = n4493 | n4494 ;
  assign n4496 = n4211 & n4461 ;
  assign n4497 = n4462 & ~n4496 ;
  assign n4498 = ( n3046 & n3185 ) | ( n3046 & n3191 ) | ( n3185 & n3191 ) ;
  assign n4499 = ( n3046 & n3184 ) | ( n3046 & n3190 ) | ( n3184 & n3190 ) ;
  assign n4500 = n3107 | n4499 ;
  assign n4501 = ~n4498 & n4500 ;
  assign n4502 = n3178 & n4043 ;
  assign n4503 = n3104 & n4045 ;
  assign n4504 = n4502 | n4503 ;
  assign n4505 = n1327 & n4048 ;
  assign n4506 = n4504 | n4505 ;
  assign n4507 = n4051 | n4506 ;
  assign n4508 = ( n4501 & n4506 ) | ( n4501 & n4507 ) | ( n4506 & n4507 ) ;
  assign n4509 = x29 & n4508 ;
  assign n4510 = x29 & ~n4509 ;
  assign n4511 = ( n4508 & ~n4509 ) | ( n4508 & n4510 ) | ( ~n4509 & n4510 ) ;
  assign n4512 = n4497 & n4511 ;
  assign n4513 = n4497 | n4511 ;
  assign n4514 = ~n4512 & n4513 ;
  assign n4515 = ( n3196 & n3355 ) | ( n3196 & n3356 ) | ( n3355 & n3356 ) ;
  assign n4516 = n1234 | n3355 ;
  assign n4517 = n3196 | n4516 ;
  assign n4518 = ~n4515 & n4517 ;
  assign n4519 = ~n1151 & n4479 ;
  assign n4520 = n1233 & n4481 ;
  assign n4521 = n4519 | n4520 ;
  assign n4522 = n3349 & n4484 ;
  assign n4523 = n4521 | n4522 ;
  assign n4524 = n4487 | n4523 ;
  assign n4525 = ( n4518 & n4523 ) | ( n4518 & n4524 ) | ( n4523 & n4524 ) ;
  assign n4526 = x26 & n4525 ;
  assign n4527 = x26 & ~n4526 ;
  assign n4528 = ( n4525 & ~n4526 ) | ( n4525 & n4527 ) | ( ~n4526 & n4527 ) ;
  assign n4529 = n4514 & n4528 ;
  assign n4530 = n4512 | n4529 ;
  assign n4531 = ~n4495 & n4530 ;
  assign n4532 = n4495 & ~n4530 ;
  assign n4533 = n4531 | n4532 ;
  assign n4534 = ~n907 & n3369 ;
  assign n4535 = n3370 | n4534 ;
  assign n4536 = ~x21 & x22 ;
  assign n4537 = x21 & ~x22 ;
  assign n4538 = n4536 | n4537 ;
  assign n4539 = x20 & ~x21 ;
  assign n4540 = ~x20 & x21 ;
  assign n4541 = n4539 | n4540 ;
  assign n4542 = ~x22 & x23 ;
  assign n4543 = x22 & ~x23 ;
  assign n4544 = n4542 | n4543 ;
  assign n4545 = ~n4541 & n4544 ;
  assign n4546 = ~n4538 & n4545 ;
  assign n4547 = ~n1014 & n4546 ;
  assign n4548 = n4538 & ~n4541 ;
  assign n4549 = n904 & n4548 ;
  assign n4550 = n4547 | n4549 ;
  assign n4551 = n4541 & ~n4544 ;
  assign n4552 = n778 & n4551 ;
  assign n4553 = n4550 | n4552 ;
  assign n4554 = n4541 & n4544 ;
  assign n4555 = n4553 | n4554 ;
  assign n4556 = ( ~n4535 & n4553 ) | ( ~n4535 & n4555 ) | ( n4553 & n4555 ) ;
  assign n4557 = ~x23 & n4556 ;
  assign n4558 = x23 | n4557 ;
  assign n4559 = ( ~n4556 & n4557 ) | ( ~n4556 & n4558 ) | ( n4557 & n4558 ) ;
  assign n4560 = ~n4533 & n4559 ;
  assign n4561 = n4533 | n4560 ;
  assign n4562 = n4533 & n4559 ;
  assign n4563 = n4514 & ~n4529 ;
  assign n4564 = ~n4514 & n4528 ;
  assign n4565 = n4446 | n4459 ;
  assign n4566 = ~n4460 & n4565 ;
  assign n4567 = ( ~n4260 & n4433 ) | ( ~n4260 & n4434 ) | ( n4433 & n4434 ) ;
  assign n4568 = n4438 & ~n4567 ;
  assign n4569 = ~n4258 & n4439 ;
  assign n4570 = n4568 | n4569 ;
  assign n4571 = n3030 & n3744 ;
  assign n4572 = n1625 & n3727 ;
  assign n4573 = ~n1733 & n3639 ;
  assign n4574 = n4572 | n4573 ;
  assign n4575 = n3636 | n4574 ;
  assign n4576 = ( n1625 & n2888 ) | ( n1625 & ~n3030 ) | ( n2888 & ~n3030 ) ;
  assign n4577 = ( ~n1625 & n3030 ) | ( ~n1625 & n4576 ) | ( n3030 & n4576 ) ;
  assign n4578 = ( ~n2888 & n4576 ) | ( ~n2888 & n4577 ) | ( n4576 & n4577 ) ;
  assign n4579 = ( n4574 & n4575 ) | ( n4574 & ~n4578 ) | ( n4575 & ~n4578 ) ;
  assign n4580 = n4571 | n4579 ;
  assign n4581 = n4570 & n4580 ;
  assign n4582 = n4570 & ~n4581 ;
  assign n4583 = ~n4570 & n4580 ;
  assign n4584 = n4582 | n4583 ;
  assign n4585 = n1532 & n4045 ;
  assign n4586 = ~n1411 & n4048 ;
  assign n4587 = ~n2939 & n4043 ;
  assign n4588 = n4586 | n4587 ;
  assign n4589 = n4585 | n4588 ;
  assign n4590 = n4051 | n4589 ;
  assign n4591 = ( ~n3930 & n4589 ) | ( ~n3930 & n4590 ) | ( n4589 & n4590 ) ;
  assign n4592 = ~x29 & n4591 ;
  assign n4593 = x29 | n4592 ;
  assign n4594 = ( ~n4591 & n4592 ) | ( ~n4591 & n4593 ) | ( n4592 & n4593 ) ;
  assign n4595 = n4584 & n4594 ;
  assign n4596 = n4439 & n4441 ;
  assign n4597 = n4442 & ~n4596 ;
  assign n4598 = ( n4581 & n4595 ) | ( n4581 & n4597 ) | ( n4595 & n4597 ) ;
  assign n4599 = n4581 | n4597 ;
  assign n4600 = n4595 | n4599 ;
  assign n4601 = ~n4598 & n4600 ;
  assign n4602 = ~n1411 & n4045 ;
  assign n4603 = n4043 | n4602 ;
  assign n4604 = ( n1532 & n4602 ) | ( n1532 & n4603 ) | ( n4602 & n4603 ) ;
  assign n4605 = n3178 & n4048 ;
  assign n4606 = n4604 | n4605 ;
  assign n4607 = n4051 | n4606 ;
  assign n4608 = ( ~n3750 & n4606 ) | ( ~n3750 & n4607 ) | ( n4606 & n4607 ) ;
  assign n4609 = ~x29 & n4608 ;
  assign n4610 = x29 | n4609 ;
  assign n4611 = ( ~n4608 & n4609 ) | ( ~n4608 & n4610 ) | ( n4609 & n4610 ) ;
  assign n4612 = n4601 & n4611 ;
  assign n4613 = n4598 | n4612 ;
  assign n4614 = n1236 & ~n3195 ;
  assign n4615 = n3196 | n4614 ;
  assign n4616 = n1327 & n4479 ;
  assign n4617 = ~n1151 & n4481 ;
  assign n4618 = n4616 | n4617 ;
  assign n4619 = n1233 & n4484 ;
  assign n4620 = n4618 | n4619 ;
  assign n4621 = n4487 | n4620 ;
  assign n4622 = ( ~n4615 & n4620 ) | ( ~n4615 & n4621 ) | ( n4620 & n4621 ) ;
  assign n4623 = ~x26 & n4622 ;
  assign n4624 = x26 | n4623 ;
  assign n4625 = ( ~n4622 & n4623 ) | ( ~n4622 & n4624 ) | ( n4623 & n4624 ) ;
  assign n4626 = ( n4566 & n4613 ) | ( n4566 & n4625 ) | ( n4613 & n4625 ) ;
  assign n4627 = n4564 | n4626 ;
  assign n4628 = n4563 | n4627 ;
  assign n4629 = ( n4563 & n4564 ) | ( n4563 & n4626 ) | ( n4564 & n4626 ) ;
  assign n4630 = ( ~n3196 & n3361 ) | ( ~n3196 & n3366 ) | ( n3361 & n3366 ) ;
  assign n4631 = n3198 & n4630 ;
  assign n4632 = n3368 & ~n4631 ;
  assign n4633 = ~n1014 & n4548 ;
  assign n4634 = ~n3255 & n4546 ;
  assign n4635 = n4633 | n4634 ;
  assign n4636 = n904 & n4551 ;
  assign n4637 = n4635 | n4636 ;
  assign n4638 = n4554 | n4637 ;
  assign n4639 = ( n4632 & n4637 ) | ( n4632 & n4638 ) | ( n4637 & n4638 ) ;
  assign n4640 = x23 & n4639 ;
  assign n4641 = x23 & ~n4640 ;
  assign n4642 = ( n4639 & ~n4640 ) | ( n4639 & n4641 ) | ( ~n4640 & n4641 ) ;
  assign n4643 = ( n4628 & n4629 ) | ( n4628 & n4642 ) | ( n4629 & n4642 ) ;
  assign n4644 = ( ~n4561 & n4562 ) | ( ~n4561 & n4643 ) | ( n4562 & n4643 ) ;
  assign n4645 = n4560 | n4644 ;
  assign n4646 = ( n3370 & ~n3602 ) | ( n3370 & n3603 ) | ( ~n3602 & n3603 ) ;
  assign n4647 = ~n905 & n3602 ;
  assign n4648 = ~n3370 & n4647 ;
  assign n4649 = n4646 | n4648 ;
  assign n4650 = n904 & n4546 ;
  assign n4651 = n778 & n4548 ;
  assign n4652 = n4650 | n4651 ;
  assign n4653 = ~n3596 & n4551 ;
  assign n4654 = n4652 | n4653 ;
  assign n4655 = n4554 | n4654 ;
  assign n4656 = ( ~n4649 & n4654 ) | ( ~n4649 & n4655 ) | ( n4654 & n4655 ) ;
  assign n4657 = ~x23 & n4656 ;
  assign n4658 = x23 | n4657 ;
  assign n4659 = ( ~n4656 & n4657 ) | ( ~n4656 & n4658 ) | ( n4657 & n4658 ) ;
  assign n4660 = n4493 | n4531 ;
  assign n4661 = n4057 | n4464 ;
  assign n4662 = n4026 | n4029 ;
  assign n4663 = ~n1411 & n3639 ;
  assign n4664 = n3178 & n3727 ;
  assign n4665 = n4663 | n4664 ;
  assign n4666 = n3104 & n3744 ;
  assign n4667 = n4665 | n4666 ;
  assign n4668 = n3636 | n4667 ;
  assign n4669 = ( n4449 & n4667 ) | ( n4449 & n4668 ) | ( n4667 & n4668 ) ;
  assign n4670 = n3784 | n4160 ;
  assign n4671 = n3658 | n4670 ;
  assign n4672 = n2056 | n2274 ;
  assign n4673 = n4671 | n4672 ;
  assign n4674 = n2176 | n4673 ;
  assign n4675 = n1045 | n1253 ;
  assign n4676 = n1128 | n4675 ;
  assign n4677 = n1260 | n4676 ;
  assign n4678 = n479 | n4677 ;
  assign n4679 = n245 | n4678 ;
  assign n4680 = n4674 | n4679 ;
  assign n4681 = n504 | n520 ;
  assign n4682 = n110 | n4681 ;
  assign n4683 = n4680 | n4682 ;
  assign n4684 = n146 | n2119 ;
  assign n4685 = n3294 | n4684 ;
  assign n4686 = n2242 | n4685 ;
  assign n4687 = n2400 | n4686 ;
  assign n4688 = n598 | n1052 ;
  assign n4689 = n3955 | n4688 ;
  assign n4690 = n1909 | n4689 ;
  assign n4691 = n697 | n2722 ;
  assign n4692 = n530 | n4691 ;
  assign n4693 = n636 | n4692 ;
  assign n4694 = n4690 | n4693 ;
  assign n4695 = n270 | n503 ;
  assign n4696 = n420 | n4695 ;
  assign n4697 = n578 | n4696 ;
  assign n4698 = n46 | n4697 ;
  assign n4699 = n449 | n4698 ;
  assign n4700 = n4694 | n4699 ;
  assign n4701 = n4687 | n4700 ;
  assign n4702 = n3808 | n4701 ;
  assign n4703 = n4683 | n4702 ;
  assign n4704 = n2508 | n2652 ;
  assign n4705 = n367 | n4704 ;
  assign n4706 = n490 | n4705 ;
  assign n4707 = n276 | n4706 ;
  assign n4708 = n351 | n4707 ;
  assign n4709 = n4703 | n4708 ;
  assign n4710 = n345 | n419 ;
  assign n4711 = n193 | n4710 ;
  assign n4712 = n114 | n4711 ;
  assign n4713 = n128 | n4712 ;
  assign n4714 = n145 | n4713 ;
  assign n4715 = n157 | n4714 ;
  assign n4716 = n4709 | n4715 ;
  assign n4717 = n4023 | n4716 ;
  assign n4718 = n4023 & n4716 ;
  assign n4719 = n4717 & ~n4718 ;
  assign n4720 = n4669 & n4719 ;
  assign n4721 = n4719 & ~n4720 ;
  assign n4722 = ( n4669 & ~n4720 ) | ( n4669 & n4721 ) | ( ~n4720 & n4721 ) ;
  assign n4723 = n4662 & n4722 ;
  assign n4724 = n4662 | n4722 ;
  assign n4725 = ~n4723 & n4724 ;
  assign n4726 = n1327 & n4043 ;
  assign n4727 = ~n1151 & n4045 ;
  assign n4728 = n4726 | n4727 ;
  assign n4729 = n1233 & n4048 ;
  assign n4730 = n4728 | n4729 ;
  assign n4731 = n4051 | n4730 ;
  assign n4732 = ( ~n4615 & n4730 ) | ( ~n4615 & n4731 ) | ( n4730 & n4731 ) ;
  assign n4733 = ~x29 & n4732 ;
  assign n4734 = x29 | n4733 ;
  assign n4735 = ( ~n4732 & n4733 ) | ( ~n4732 & n4734 ) | ( n4733 & n4734 ) ;
  assign n4736 = n4725 & n4735 ;
  assign n4737 = n4725 | n4735 ;
  assign n4738 = ~n4736 & n4737 ;
  assign n4739 = ( n3196 & n3360 ) | ( n3196 & n3365 ) | ( n3360 & n3365 ) ;
  assign n4740 = ( n3196 & n3359 ) | ( n3196 & n3364 ) | ( n3359 & n3364 ) ;
  assign n4741 = n3258 | n4740 ;
  assign n4742 = ~n4739 & n4741 ;
  assign n4743 = ~n1014 & n4484 ;
  assign n4744 = n3349 & n4479 ;
  assign n4745 = ~n3255 & n4481 ;
  assign n4746 = n4744 | n4745 ;
  assign n4747 = n4743 | n4746 ;
  assign n4748 = n4487 | n4747 ;
  assign n4749 = ( n4742 & n4747 ) | ( n4742 & n4748 ) | ( n4747 & n4748 ) ;
  assign n4750 = x26 & n4749 ;
  assign n4751 = x26 & ~n4750 ;
  assign n4752 = ( n4749 & ~n4750 ) | ( n4749 & n4751 ) | ( ~n4750 & n4751 ) ;
  assign n4753 = ( n4661 & n4738 ) | ( n4661 & n4752 ) | ( n4738 & n4752 ) ;
  assign n4754 = ( n4738 & n4752 ) | ( n4738 & ~n4753 ) | ( n4752 & ~n4753 ) ;
  assign n4755 = ( n4661 & ~n4753 ) | ( n4661 & n4754 ) | ( ~n4753 & n4754 ) ;
  assign n4756 = ( n4659 & ~n4660 ) | ( n4659 & n4755 ) | ( ~n4660 & n4755 ) ;
  assign n4757 = ( n4660 & ~n4755 ) | ( n4660 & n4756 ) | ( ~n4755 & n4756 ) ;
  assign n4758 = ( ~n4659 & n4756 ) | ( ~n4659 & n4757 ) | ( n4756 & n4757 ) ;
  assign n4759 = n4645 & n4758 ;
  assign n4760 = n4645 | n4758 ;
  assign n4761 = ~n4759 & n4760 ;
  assign n4762 = ( n3370 & n3609 ) | ( n3370 & n3615 ) | ( n3609 & n3615 ) ;
  assign n4763 = ( n3370 & n3608 ) | ( n3370 & ~n3614 ) | ( n3608 & ~n3614 ) ;
  assign n4764 = n3434 | n4763 ;
  assign n4765 = ~n4762 & n4764 ;
  assign n4766 = ~x18 & x19 ;
  assign n4767 = x18 & ~x19 ;
  assign n4768 = n4766 | n4767 ;
  assign n4769 = x19 & ~x20 ;
  assign n4770 = ~x19 & x20 ;
  assign n4771 = n4769 | n4770 ;
  assign n4772 = x17 & ~x18 ;
  assign n4773 = ~x17 & x18 ;
  assign n4774 = n4772 | n4773 ;
  assign n4775 = n4771 & ~n4774 ;
  assign n4776 = ~n4768 & n4775 ;
  assign n4777 = n3504 & n4776 ;
  assign n4778 = n4768 & ~n4774 ;
  assign n4779 = ~n3431 & n4778 ;
  assign n4780 = n4777 | n4779 ;
  assign n4781 = ~n4771 & n4774 ;
  assign n4782 = ~n589 & n4781 ;
  assign n4783 = n4780 | n4782 ;
  assign n4784 = n4771 & n4774 ;
  assign n4785 = n4783 | n4784 ;
  assign n4786 = ( n4765 & n4783 ) | ( n4765 & n4785 ) | ( n4783 & n4785 ) ;
  assign n4787 = x20 & n4786 ;
  assign n4788 = x20 & ~n4787 ;
  assign n4789 = ( n4786 & ~n4787 ) | ( n4786 & n4788 ) | ( ~n4787 & n4788 ) ;
  assign n4790 = n4761 & n4789 ;
  assign n4791 = n4761 & ~n4790 ;
  assign n4792 = n4562 | n4643 ;
  assign n4793 = n4561 & ~n4792 ;
  assign n4794 = n4644 | n4793 ;
  assign n4795 = ( n3370 & n3607 ) | ( n3370 & ~n3613 ) | ( n3607 & ~n3613 ) ;
  assign n4796 = ( n3370 & n3606 ) | ( n3370 & ~n3612 ) | ( n3606 & ~n3612 ) ;
  assign n4797 = n3507 & ~n4796 ;
  assign n4798 = n4795 | n4797 ;
  assign n4799 = ~n3596 & n4776 ;
  assign n4800 = n3504 & n4778 ;
  assign n4801 = n4799 | n4800 ;
  assign n4802 = ~n3431 & n4781 ;
  assign n4803 = n4801 | n4802 ;
  assign n4804 = n4784 | n4803 ;
  assign n4805 = ( ~n4798 & n4803 ) | ( ~n4798 & n4804 ) | ( n4803 & n4804 ) ;
  assign n4806 = ~x20 & n4805 ;
  assign n4807 = x20 | n4806 ;
  assign n4808 = ( ~n4805 & n4806 ) | ( ~n4805 & n4807 ) | ( n4806 & n4807 ) ;
  assign n4809 = ~n4794 & n4808 ;
  assign n4810 = n4794 & ~n4808 ;
  assign n4811 = n4809 | n4810 ;
  assign n4812 = n4628 & ~n4629 ;
  assign n4813 = ~n4642 & n4812 ;
  assign n4814 = n4642 | n4813 ;
  assign n4815 = ( ~n4812 & n4813 ) | ( ~n4812 & n4814 ) | ( n4813 & n4814 ) ;
  assign n4816 = n4601 & ~n4612 ;
  assign n4817 = ~n4601 & n4611 ;
  assign n4818 = n3104 & n4479 ;
  assign n4819 = n1327 & n4481 ;
  assign n4820 = n4818 | n4819 ;
  assign n4821 = ~n1151 & n4484 ;
  assign n4822 = n4820 | n4821 ;
  assign n4823 = n4487 | n4822 ;
  assign n4824 = ( ~n4034 & n4822 ) | ( ~n4034 & n4823 ) | ( n4822 & n4823 ) ;
  assign n4825 = ~x26 & n4824 ;
  assign n4826 = x26 | n4825 ;
  assign n4827 = ( ~n4824 & n4825 ) | ( ~n4824 & n4826 ) | ( n4825 & n4826 ) ;
  assign n4828 = ( n4816 & n4817 ) | ( n4816 & n4827 ) | ( n4817 & n4827 ) ;
  assign n4829 = n4817 | n4827 ;
  assign n4830 = n4816 | n4829 ;
  assign n4831 = ~n4828 & n4830 ;
  assign n4832 = n4584 | n4594 ;
  assign n4833 = ~n4595 & n4832 ;
  assign n4834 = n3636 | n4432 ;
  assign n4835 = ( n4260 & n4432 ) | ( n4260 & n4834 ) | ( n4432 & n4834 ) ;
  assign n4836 = n4116 | n4426 ;
  assign n4837 = ~n4427 & n4836 ;
  assign n4838 = n4835 & n4837 ;
  assign n4839 = n4837 & ~n4838 ;
  assign n4840 = ( n4835 & ~n4838 ) | ( n4835 & n4839 ) | ( ~n4838 & n4839 ) ;
  assign n4841 = n373 | n1261 ;
  assign n4842 = n409 | n509 ;
  assign n4843 = n625 | n4842 ;
  assign n4844 = n4841 | n4843 ;
  assign n4845 = n948 | n4844 ;
  assign n4846 = n2980 | n2982 ;
  assign n4847 = n4845 | n4846 ;
  assign n4848 = n791 | n2163 ;
  assign n4849 = n529 | n609 ;
  assign n4850 = n4848 | n4849 ;
  assign n4851 = n212 | n277 ;
  assign n4852 = n438 | n4851 ;
  assign n4853 = n404 | n4852 ;
  assign n4854 = n4850 | n4853 ;
  assign n4855 = n76 | n120 ;
  assign n4856 = n168 | n4855 ;
  assign n4857 = n661 | n4856 ;
  assign n4858 = n4854 | n4857 ;
  assign n4859 = n4847 | n4858 ;
  assign n4860 = n959 | n1115 ;
  assign n4861 = n1417 | n4860 ;
  assign n4862 = n266 | n4861 ;
  assign n4863 = n349 | n4862 ;
  assign n4864 = n590 | n4863 ;
  assign n4865 = n4859 | n4864 ;
  assign n4866 = n46 | n4865 ;
  assign n4867 = n489 | n655 ;
  assign n4868 = n358 | n4867 ;
  assign n4869 = n1177 | n4868 ;
  assign n4870 = n4390 | n4869 ;
  assign n4871 = n1031 | n4870 ;
  assign n4872 = n4298 | n4871 ;
  assign n4873 = n101 | n887 ;
  assign n4874 = n670 | n4873 ;
  assign n4875 = n112 | n441 ;
  assign n4876 = n2341 | n4875 ;
  assign n4877 = n730 | n4876 ;
  assign n4878 = n4874 | n4877 ;
  assign n4879 = n143 | n513 ;
  assign n4880 = n1956 | n4879 ;
  assign n4881 = n1852 | n4880 ;
  assign n4882 = n1613 | n4881 ;
  assign n4883 = n4878 | n4882 ;
  assign n4884 = n293 | n478 ;
  assign n4885 = n213 | n4884 ;
  assign n4886 = n437 | n4885 ;
  assign n4887 = n227 | n4886 ;
  assign n4888 = n224 | n4887 ;
  assign n4889 = n4883 | n4888 ;
  assign n4890 = n4872 | n4889 ;
  assign n4891 = n4866 | n4890 ;
  assign n4892 = n2029 | n2527 ;
  assign n4893 = ( n633 & ~n3163 ) | ( n633 & n4892 ) | ( ~n3163 & n4892 ) ;
  assign n4894 = n3163 | n4893 ;
  assign n4895 = n250 | n4894 ;
  assign n4896 = n383 | n4895 ;
  assign n4897 = n393 | n4896 ;
  assign n4898 = n451 | n4897 ;
  assign n4899 = n4891 | n4898 ;
  assign n4900 = n55 | n57 ;
  assign n4901 = n4899 | n4900 ;
  assign n4902 = n4334 & n4901 ;
  assign n4903 = n4334 | n4901 ;
  assign n4904 = n1883 & n2790 ;
  assign n4905 = n2791 & ~n4904 ;
  assign n4906 = n1803 & n3744 ;
  assign n4907 = ~n1944 & n3639 ;
  assign n4908 = n4906 | n4907 ;
  assign n4909 = ~n1880 & n3727 ;
  assign n4910 = n4908 | n4909 ;
  assign n4911 = n3636 | n4910 ;
  assign n4912 = n489 | n582 ;
  assign n4913 = n140 | n4912 ;
  assign n4914 = n622 | n669 ;
  assign n4915 = n277 | n4914 ;
  assign n4916 = n4913 | n4915 ;
  assign n4917 = n428 | n521 ;
  assign n4918 = n293 | n4917 ;
  assign n4919 = n358 | n4918 ;
  assign n4920 = n4916 | n4919 ;
  assign n4921 = n186 | n204 ;
  assign n4922 = n122 | n4921 ;
  assign n4923 = n4920 | n4922 ;
  assign n4924 = n499 | n539 ;
  assign n4925 = n504 | n4924 ;
  assign n4926 = n253 | n519 ;
  assign n4927 = n351 | n4926 ;
  assign n4928 = n155 | n434 ;
  assign n4929 = n207 | n4928 ;
  assign n4930 = n479 | n4929 ;
  assign n4931 = n4927 | n4930 ;
  assign n4932 = n4925 | n4931 ;
  assign n4933 = n1522 | n4932 ;
  assign n4934 = n4923 | n4933 ;
  assign n4935 = n1128 | n3243 ;
  assign n4936 = n2736 | n4935 ;
  assign n4937 = n637 | n4936 ;
  assign n4938 = n258 | n4937 ;
  assign n4939 = n249 | n4938 ;
  assign n4940 = n4934 | n4939 ;
  assign n4941 = n227 | n409 ;
  assign n4942 = n646 | n4941 ;
  assign n4943 = n999 | n4942 ;
  assign n4944 = n309 | n452 ;
  assign n4945 = n441 | n4944 ;
  assign n4946 = n180 | n4945 ;
  assign n4947 = n4943 | n4946 ;
  assign n4948 = n4940 | n4947 ;
  assign n4949 = n3968 | n4948 ;
  assign n4950 = n868 | n2989 ;
  assign n4951 = n134 | n475 ;
  assign n4952 = n197 | n4951 ;
  assign n4953 = n4950 | n4952 ;
  assign n4954 = n128 | n213 ;
  assign n4955 = n4953 | n4954 ;
  assign n4956 = n1222 | n4955 ;
  assign n4957 = n869 | n4956 ;
  assign n4958 = n920 | n4957 ;
  assign n4959 = n2732 | n4958 ;
  assign n4960 = n468 | n4959 ;
  assign n4961 = n4949 | n4960 ;
  assign n4962 = n470 | n621 ;
  assign n4963 = n306 | n4962 ;
  assign n4964 = n435 | n4963 ;
  assign n4965 = n570 | n4964 ;
  assign n4966 = n111 | n4965 ;
  assign n4967 = n218 | n4966 ;
  assign n4968 = n650 | n4967 ;
  assign n4969 = n4961 | n4968 ;
  assign n4970 = ( x2 & x5 ) | ( x2 & ~n4969 ) | ( x5 & ~n4969 ) ;
  assign n4971 = ( n4334 & n4911 ) | ( n4334 & ~n4970 ) | ( n4911 & ~n4970 ) ;
  assign n4972 = ~n4902 & n4971 ;
  assign n4973 = n4334 & ~n4970 ;
  assign n4974 = ~n4334 & n4970 ;
  assign n4975 = n4973 | n4974 ;
  assign n4976 = n4910 & ~n4975 ;
  assign n4977 = n4973 | n4976 ;
  assign n4978 = ~n4902 & n4977 ;
  assign n4979 = ( n4905 & n4972 ) | ( n4905 & n4978 ) | ( n4972 & n4978 ) ;
  assign n4980 = n4903 & n4979 ;
  assign n4981 = n4902 | n4980 ;
  assign n4982 = ( ~n2791 & n2882 ) | ( ~n2791 & n2884 ) | ( n2882 & n2884 ) ;
  assign n4983 = ( n2791 & n2878 ) | ( n2791 & ~n2881 ) | ( n2878 & ~n2881 ) ;
  assign n4984 = ~n2876 & n4983 ;
  assign n4985 = n4982 | n4984 ;
  assign n4986 = n1803 & n3639 ;
  assign n4987 = ~n2873 & n3727 ;
  assign n4988 = n4986 | n4987 ;
  assign n4989 = ~n1733 & n3744 ;
  assign n4990 = n4988 | n4989 ;
  assign n4991 = n3636 | n4990 ;
  assign n4992 = ( ~n4985 & n4990 ) | ( ~n4985 & n4991 ) | ( n4990 & n4991 ) ;
  assign n4993 = ( ~n4334 & n4425 ) | ( ~n4334 & n4426 ) | ( n4425 & n4426 ) ;
  assign n4994 = ( ~x8 & n4426 ) | ( ~x8 & n4993 ) | ( n4426 & n4993 ) ;
  assign n4995 = ( n4981 & n4992 ) | ( n4981 & n4994 ) | ( n4992 & n4994 ) ;
  assign n4996 = n4840 & n4995 ;
  assign n4997 = n4840 | n4995 ;
  assign n4998 = ~n4996 & n4997 ;
  assign n4999 = n1532 & n4048 ;
  assign n5000 = n3030 & n4043 ;
  assign n5001 = ~n2939 & n4045 ;
  assign n5002 = n5000 | n5001 ;
  assign n5003 = n4999 | n5002 ;
  assign n5004 = n4051 | n5003 ;
  assign n5005 = ( ~n4193 & n5003 ) | ( ~n4193 & n5004 ) | ( n5003 & n5004 ) ;
  assign n5006 = ~x29 & n5005 ;
  assign n5007 = x29 | n5006 ;
  assign n5008 = ( ~n5005 & n5006 ) | ( ~n5005 & n5007 ) | ( n5006 & n5007 ) ;
  assign n5009 = n4998 & n5008 ;
  assign n5010 = n4996 | n5009 ;
  assign n5011 = n3178 & n4479 ;
  assign n5012 = n3104 & n4481 ;
  assign n5013 = n5011 | n5012 ;
  assign n5014 = n1327 & n4484 ;
  assign n5015 = n5013 | n5014 ;
  assign n5016 = n4487 | n5015 ;
  assign n5017 = ( n4501 & n5015 ) | ( n4501 & n5016 ) | ( n5015 & n5016 ) ;
  assign n5018 = x26 & n5017 ;
  assign n5019 = x26 & ~n5018 ;
  assign n5020 = ( n5017 & ~n5018 ) | ( n5017 & n5019 ) | ( ~n5018 & n5019 ) ;
  assign n5021 = ( n4833 & n5010 ) | ( n4833 & n5020 ) | ( n5010 & n5020 ) ;
  assign n5022 = n4831 & n5021 ;
  assign n5023 = n4828 | n5022 ;
  assign n5024 = ~n1014 & n4551 ;
  assign n5025 = n3349 & n4546 ;
  assign n5026 = ~n3255 & n4548 ;
  assign n5027 = n5025 | n5026 ;
  assign n5028 = n5024 | n5027 ;
  assign n5029 = n4554 | n5028 ;
  assign n5030 = ( n4742 & n5028 ) | ( n4742 & n5029 ) | ( n5028 & n5029 ) ;
  assign n5031 = x23 & n5030 ;
  assign n5032 = x23 & ~n5031 ;
  assign n5033 = ( n5030 & ~n5031 ) | ( n5030 & n5032 ) | ( ~n5031 & n5032 ) ;
  assign n5034 = ( n4566 & n4625 ) | ( n4566 & ~n4626 ) | ( n4625 & ~n4626 ) ;
  assign n5035 = ( n4613 & ~n4626 ) | ( n4613 & n5034 ) | ( ~n4626 & n5034 ) ;
  assign n5036 = ( n5023 & n5033 ) | ( n5023 & n5035 ) | ( n5033 & n5035 ) ;
  assign n5037 = ( n3370 & n3605 ) | ( n3370 & ~n3611 ) | ( n3605 & ~n3611 ) ;
  assign n5038 = ( n3370 & ~n3601 ) | ( n3370 & n3604 ) | ( ~n3601 & n3604 ) ;
  assign n5039 = n3599 & ~n5038 ;
  assign n5040 = n5037 | n5039 ;
  assign n5041 = n778 & n4776 ;
  assign n5042 = ~n3596 & n4778 ;
  assign n5043 = n5041 | n5042 ;
  assign n5044 = n3504 & n4781 ;
  assign n5045 = n5043 | n5044 ;
  assign n5046 = n4784 | n5045 ;
  assign n5047 = ( ~n5040 & n5045 ) | ( ~n5040 & n5046 ) | ( n5045 & n5046 ) ;
  assign n5048 = ~x20 & n5047 ;
  assign n5049 = x20 | n5048 ;
  assign n5050 = ( ~n5047 & n5048 ) | ( ~n5047 & n5049 ) | ( n5048 & n5049 ) ;
  assign n5051 = ( n4815 & n5036 ) | ( n4815 & n5050 ) | ( n5036 & n5050 ) ;
  assign n5052 = ~n4811 & n5051 ;
  assign n5053 = n4809 | n5052 ;
  assign n5054 = ~n4761 & n4789 ;
  assign n5055 = n5053 | n5054 ;
  assign n5056 = n4791 | n5055 ;
  assign n5057 = ( n4791 & n5053 ) | ( n4791 & n5054 ) | ( n5053 & n5054 ) ;
  assign n5058 = n5056 & ~n5057 ;
  assign n5059 = ~x15 & x16 ;
  assign n5060 = x15 & ~x16 ;
  assign n5061 = n5059 | n5060 ;
  assign n5062 = x14 & ~x15 ;
  assign n5063 = ~x14 & x15 ;
  assign n5064 = n5062 | n5063 ;
  assign n5065 = x16 & ~x17 ;
  assign n5066 = ~x16 & x17 ;
  assign n5067 = n5065 | n5066 ;
  assign n5068 = ~n5064 & n5067 ;
  assign n5069 = ~n5061 & n5068 ;
  assign n5070 = n5061 & ~n5064 ;
  assign n5071 = ~n3634 & n5070 ;
  assign n5072 = n672 & n5069 ;
  assign n5073 = ( n5069 & n5071 ) | ( n5069 & ~n5072 ) | ( n5071 & ~n5072 ) ;
  assign n5074 = n5064 & n5067 ;
  assign n5075 = n5073 | n5074 ;
  assign n5076 = ( n3726 & n5073 ) | ( n3726 & n5075 ) | ( n5073 & n5075 ) ;
  assign n5077 = x17 & n5076 ;
  assign n5078 = x17 & ~n5077 ;
  assign n5079 = ( n5076 & ~n5077 ) | ( n5076 & n5078 ) | ( ~n5077 & n5078 ) ;
  assign n5080 = n5058 & ~n5079 ;
  assign n5081 = n5079 | n5080 ;
  assign n5082 = ( ~n5058 & n5080 ) | ( ~n5058 & n5081 ) | ( n5080 & n5081 ) ;
  assign n5083 = n5064 & ~n5067 ;
  assign n5084 = ~n3634 & n5083 ;
  assign n5085 = ~n672 & n5070 ;
  assign n5086 = n5084 | n5085 ;
  assign n5087 = ~n589 & n5069 ;
  assign n5088 = n5086 | n5087 ;
  assign n5089 = n5074 | n5088 ;
  assign n5090 = ( ~n672 & n3619 ) | ( ~n672 & n3634 ) | ( n3619 & n3634 ) ;
  assign n5091 = ( n672 & ~n3634 ) | ( n672 & n5090 ) | ( ~n3634 & n5090 ) ;
  assign n5092 = ( ~n3619 & n5090 ) | ( ~n3619 & n5091 ) | ( n5090 & n5091 ) ;
  assign n5093 = ( n5088 & n5089 ) | ( n5088 & ~n5092 ) | ( n5089 & ~n5092 ) ;
  assign n5094 = ~x17 & n5093 ;
  assign n5095 = x17 | n5094 ;
  assign n5096 = ( ~n5093 & n5094 ) | ( ~n5093 & n5095 ) | ( n5094 & n5095 ) ;
  assign n5097 = n4831 | n5021 ;
  assign n5098 = ~n5022 & n5097 ;
  assign n5099 = n1233 & n4546 ;
  assign n5100 = n3349 & n4548 ;
  assign n5101 = n5099 | n5100 ;
  assign n5102 = ~n3255 & n4551 ;
  assign n5103 = n5101 | n5102 ;
  assign n5104 = n4554 | n5103 ;
  assign n5105 = ( ~n4470 & n5103 ) | ( ~n4470 & n5104 ) | ( n5103 & n5104 ) ;
  assign n5106 = ~x23 & n5105 ;
  assign n5107 = x23 | n5106 ;
  assign n5108 = ( ~n5105 & n5106 ) | ( ~n5105 & n5107 ) | ( n5106 & n5107 ) ;
  assign n5109 = n5098 & n5108 ;
  assign n5110 = n5108 & ~n5109 ;
  assign n5111 = ( n5098 & ~n5109 ) | ( n5098 & n5110 ) | ( ~n5109 & n5110 ) ;
  assign n5112 = n4998 | n5008 ;
  assign n5113 = ~n5009 & n5112 ;
  assign n5114 = n1625 & n4043 ;
  assign n5115 = n3030 & n4045 ;
  assign n5116 = n5114 | n5115 ;
  assign n5117 = ~n2939 & n4048 ;
  assign n5118 = n5116 | n5117 ;
  assign n5119 = n4051 | n5118 ;
  assign n5120 = ( ~n4215 & n5118 ) | ( ~n4215 & n5119 ) | ( n5118 & n5119 ) ;
  assign n5121 = ~x29 & n5120 ;
  assign n5122 = x29 | n5121 ;
  assign n5123 = ( ~n5120 & n5121 ) | ( ~n5120 & n5122 ) | ( n5121 & n5122 ) ;
  assign n5124 = ( n4981 & n4992 ) | ( n4981 & ~n4994 ) | ( n4992 & ~n4994 ) ;
  assign n5125 = ( ~n4981 & n4994 ) | ( ~n4981 & n5124 ) | ( n4994 & n5124 ) ;
  assign n5126 = ( ~n4992 & n5124 ) | ( ~n4992 & n5125 ) | ( n5124 & n5125 ) ;
  assign n5127 = n5123 & n5126 ;
  assign n5128 = n5126 & ~n5127 ;
  assign n5129 = n5123 & ~n5126 ;
  assign n5130 = n5128 | n5129 ;
  assign n5131 = ( n4905 & n4971 ) | ( n4905 & n4977 ) | ( n4971 & n4977 ) ;
  assign n5132 = ~n4980 & n5131 ;
  assign n5133 = n4903 & ~n4981 ;
  assign n5134 = n5132 | n5133 ;
  assign n5135 = ~n2873 & n3744 ;
  assign n5136 = ( n2791 & n2879 ) | ( n2791 & ~n2880 ) | ( n2879 & ~n2880 ) ;
  assign n5137 = ~n1881 & n2879 ;
  assign n5138 = n2791 & n5137 ;
  assign n5139 = n5136 & ~n5138 ;
  assign n5140 = n1803 & n3727 ;
  assign n5141 = ~n1880 & n3639 ;
  assign n5142 = n5140 | n5141 ;
  assign n5143 = n3636 | n5142 ;
  assign n5144 = ( n5139 & n5142 ) | ( n5139 & n5143 ) | ( n5142 & n5143 ) ;
  assign n5145 = n5135 | n5144 ;
  assign n5146 = n5134 & n5145 ;
  assign n5147 = ( n4905 & n4910 ) | ( n4905 & n4911 ) | ( n4910 & n4911 ) ;
  assign n5148 = n4975 & n5147 ;
  assign n5149 = n4975 & ~n5148 ;
  assign n5150 = ( n5147 & ~n5148 ) | ( n5147 & n5149 ) | ( ~n5148 & n5149 ) ;
  assign n5151 = ( ~x5 & n4969 ) | ( ~x5 & n4970 ) | ( n4969 & n4970 ) ;
  assign n5152 = ( ~x2 & n4970 ) | ( ~x2 & n5151 ) | ( n4970 & n5151 ) ;
  assign n5153 = n3775 | n4239 ;
  assign n5154 = n4121 | n5153 ;
  assign n5155 = n3145 | n5154 ;
  assign n5156 = n398 | n5155 ;
  assign n5157 = n2035 | n5156 ;
  assign n5158 = n1696 | n2610 ;
  assign n5159 = n409 | n833 ;
  assign n5160 = n5158 | n5159 ;
  assign n5161 = n199 | n708 ;
  assign n5162 = n661 | n5161 ;
  assign n5163 = n5160 | n5162 ;
  assign n5164 = n2379 & ~n5163 ;
  assign n5165 = ~n5157 & n5164 ;
  assign n5166 = n637 | n655 ;
  assign n5167 = n2060 | n5166 ;
  assign n5168 = n282 | n450 ;
  assign n5169 = n442 | n5168 ;
  assign n5170 = n5167 | n5169 ;
  assign n5171 = n890 | n5170 ;
  assign n5172 = n3873 | n5171 ;
  assign n5173 = n473 | n5172 ;
  assign n5174 = n194 | n5173 ;
  assign n5175 = n161 | n5174 ;
  assign n5176 = n140 | n5175 ;
  assign n5177 = n5165 & ~n5176 ;
  assign n5178 = x2 | n218 ;
  assign n5179 = n5177 & ~n5178 ;
  assign n5180 = n955 | n3814 ;
  assign n5181 = n443 | n5180 ;
  assign n5182 = n611 | n5181 ;
  assign n5183 = n1311 | n5182 ;
  assign n5184 = n1115 | n5183 ;
  assign n5185 = n1032 | n1561 ;
  assign n5186 = n273 | n335 ;
  assign n5187 = n252 | n5186 ;
  assign n5188 = n5185 | n5187 ;
  assign n5189 = n301 | n346 ;
  assign n5190 = n607 | n5189 ;
  assign n5191 = n393 | n5190 ;
  assign n5192 = n5188 | n5191 ;
  assign n5193 = ( ~n44 & n195 ) | ( ~n44 & n578 ) | ( n195 & n578 ) ;
  assign n5194 = n5192 | n5193 ;
  assign n5195 = n1200 | n3850 ;
  assign n5196 = n473 | n3903 ;
  assign n5197 = n5195 | n5196 ;
  assign n5198 = n687 | n5197 ;
  assign n5199 = ( ~n3215 & n5194 ) | ( ~n3215 & n5198 ) | ( n5194 & n5198 ) ;
  assign n5200 = n3215 | n5199 ;
  assign n5201 = ( ~n2499 & n5184 ) | ( ~n2499 & n5200 ) | ( n5184 & n5200 ) ;
  assign n5202 = n2499 | n5201 ;
  assign n5203 = n314 | n1990 ;
  assign n5204 = n570 | n5203 ;
  assign n5205 = n601 | n5204 ;
  assign n5206 = n173 | n5205 ;
  assign n5207 = n145 | n5206 ;
  assign n5208 = n227 | n5207 ;
  assign n5209 = x2 & n5208 ;
  assign n5210 = ( x2 & n5202 ) | ( x2 & n5209 ) | ( n5202 & n5209 ) ;
  assign n5211 = x2 & n218 ;
  assign n5212 = ( x2 & ~n5177 ) | ( x2 & n5211 ) | ( ~n5177 & n5211 ) ;
  assign n5213 = n5210 | n5212 ;
  assign n5214 = ( n2193 & n2296 ) | ( n2193 & ~n2776 ) | ( n2296 & ~n2776 ) ;
  assign n5215 = n2196 | n5214 ;
  assign n5216 = ~n2777 & n5215 ;
  assign n5217 = n2461 | n4237 ;
  assign n5218 = n168 | n345 ;
  assign n5219 = n1779 | n5218 ;
  assign n5220 = n5217 | n5219 ;
  assign n5221 = n4307 | n5220 ;
  assign n5222 = n842 | n890 ;
  assign n5223 = n611 | n5222 ;
  assign n5224 = n638 | n5223 ;
  assign n5225 = n5221 | n5224 ;
  assign n5226 = n244 | n629 ;
  assign n5227 = n253 | n5226 ;
  assign n5228 = n319 | n5227 ;
  assign n5229 = n155 | n5228 ;
  assign n5230 = n5225 | n5229 ;
  assign n5231 = n442 | n529 ;
  assign n5232 = n3864 | n5231 ;
  assign n5233 = n2119 | n3809 ;
  assign n5234 = n5232 | n5233 ;
  assign n5235 = n2688 | n5234 ;
  assign n5236 = n416 | n488 ;
  assign n5237 = n648 | n5236 ;
  assign n5238 = n62 | n193 ;
  assign n5239 = n83 | n5238 ;
  assign n5240 = n5237 | n5239 ;
  assign n5241 = n5235 | n5240 ;
  assign n5242 = n2731 | n5241 ;
  assign n5243 = n1544 | n1596 ;
  assign n5244 = n310 | n540 ;
  assign n5245 = n241 | n5244 ;
  assign n5246 = n5243 | n5245 ;
  assign n5247 = n320 | n408 ;
  assign n5248 = n112 | n5247 ;
  assign n5249 = n5246 | n5248 ;
  assign n5250 = n5242 | n5249 ;
  assign n5251 = n5230 | n5250 ;
  assign n5252 = n1220 | n5251 ;
  assign n5253 = n1454 | n5252 ;
  assign n5254 = n92 | n3873 ;
  assign n5255 = ( n152 & ~n3843 ) | ( n152 & n5254 ) | ( ~n3843 & n5254 ) ;
  assign n5256 = n3843 | n5255 ;
  assign n5257 = x2 & n5256 ;
  assign n5258 = ( x2 & n5253 ) | ( x2 & n5257 ) | ( n5253 & n5257 ) ;
  assign n5259 = x2 | n5256 ;
  assign n5260 = n5253 | n5259 ;
  assign n5261 = n2296 & n3639 ;
  assign n5262 = n2193 & n3727 ;
  assign n5263 = n5261 | n5262 ;
  assign n5264 = n2013 & n3744 ;
  assign n5265 = n5263 | n5264 ;
  assign n5266 = n3636 | n5265 ;
  assign n5267 = ~n5258 & n5266 ;
  assign n5268 = n5260 & n5267 ;
  assign n5269 = n5258 | n5268 ;
  assign n5270 = ~n5258 & n5265 ;
  assign n5271 = n5260 & n5270 ;
  assign n5272 = n5258 | n5271 ;
  assign n5273 = ( n5216 & n5269 ) | ( n5216 & n5272 ) | ( n5269 & n5272 ) ;
  assign n5274 = x2 | n5208 ;
  assign n5275 = n5202 | n5274 ;
  assign n5276 = ~n5210 & n5275 ;
  assign n5277 = n5273 & n5276 ;
  assign n5278 = ( ~n5179 & n5213 ) | ( ~n5179 & n5277 ) | ( n5213 & n5277 ) ;
  assign n5279 = ( ~n2779 & n2783 ) | ( ~n2779 & n2786 ) | ( n2783 & n2786 ) ;
  assign n5280 = ~n2781 & n5279 ;
  assign n5281 = n2789 | n5280 ;
  assign n5282 = ~n2103 & n3639 ;
  assign n5283 = ~n1944 & n3727 ;
  assign n5284 = n5282 | n5283 ;
  assign n5285 = ~n1880 & n3744 ;
  assign n5286 = n5284 | n5285 ;
  assign n5287 = n3636 | n5286 ;
  assign n5288 = ( ~n5281 & n5286 ) | ( ~n5281 & n5287 ) | ( n5286 & n5287 ) ;
  assign n5289 = ( n5152 & n5278 ) | ( n5152 & n5288 ) | ( n5278 & n5288 ) ;
  assign n5290 = ~n5150 & n5289 ;
  assign n5291 = n5150 & ~n5289 ;
  assign n5292 = n5290 | n5291 ;
  assign n5293 = ~n2873 & n4043 ;
  assign n5294 = ~n1733 & n4045 ;
  assign n5295 = n5293 | n5294 ;
  assign n5296 = n1625 & n4048 ;
  assign n5297 = n5295 | n5296 ;
  assign n5298 = n4051 | n5297 ;
  assign n5299 = ( n4260 & n5297 ) | ( n4260 & n5298 ) | ( n5297 & n5298 ) ;
  assign n5300 = x29 & n5299 ;
  assign n5301 = x29 & ~n5300 ;
  assign n5302 = ( n5299 & ~n5300 ) | ( n5299 & n5301 ) | ( ~n5300 & n5301 ) ;
  assign n5303 = ~n5292 & n5302 ;
  assign n5304 = n5290 | n5303 ;
  assign n5305 = n5134 & ~n5146 ;
  assign n5306 = ~n5134 & n5145 ;
  assign n5307 = n5305 | n5306 ;
  assign n5308 = n5304 & n5307 ;
  assign n5309 = n5146 | n5308 ;
  assign n5310 = n5130 & n5309 ;
  assign n5311 = n5127 | n5310 ;
  assign n5312 = ~n1411 & n4479 ;
  assign n5313 = n3178 & n4481 ;
  assign n5314 = n5312 | n5313 ;
  assign n5315 = n3104 & n4484 ;
  assign n5316 = n5314 | n5315 ;
  assign n5317 = n4487 | n5316 ;
  assign n5318 = ( n4449 & n5316 ) | ( n4449 & n5317 ) | ( n5316 & n5317 ) ;
  assign n5319 = x26 & n5318 ;
  assign n5320 = x26 & ~n5319 ;
  assign n5321 = ( n5318 & ~n5319 ) | ( n5318 & n5320 ) | ( ~n5319 & n5320 ) ;
  assign n5322 = ( n5113 & n5311 ) | ( n5113 & n5321 ) | ( n5311 & n5321 ) ;
  assign n5323 = ~n1151 & n4546 ;
  assign n5324 = n1233 & n4548 ;
  assign n5325 = n5323 | n5324 ;
  assign n5326 = n3349 & n4551 ;
  assign n5327 = n5325 | n5326 ;
  assign n5328 = n4554 | n5327 ;
  assign n5329 = ( n4518 & n5327 ) | ( n4518 & n5328 ) | ( n5327 & n5328 ) ;
  assign n5330 = x23 & n5329 ;
  assign n5331 = x23 & ~n5330 ;
  assign n5332 = ( n5329 & ~n5330 ) | ( n5329 & n5331 ) | ( ~n5330 & n5331 ) ;
  assign n5333 = ( n4833 & n5020 ) | ( n4833 & ~n5021 ) | ( n5020 & ~n5021 ) ;
  assign n5334 = ( n5010 & ~n5021 ) | ( n5010 & n5333 ) | ( ~n5021 & n5333 ) ;
  assign n5335 = ( n5322 & n5332 ) | ( n5322 & n5334 ) | ( n5332 & n5334 ) ;
  assign n5336 = n5111 & n5335 ;
  assign n5337 = n5109 | n5336 ;
  assign n5338 = n904 & n4776 ;
  assign n5339 = n778 & n4778 ;
  assign n5340 = n5338 | n5339 ;
  assign n5341 = ~n3596 & n4781 ;
  assign n5342 = n5340 | n5341 ;
  assign n5343 = n4784 | n5342 ;
  assign n5344 = ( ~n4649 & n5342 ) | ( ~n4649 & n5343 ) | ( n5342 & n5343 ) ;
  assign n5345 = ~x20 & n5344 ;
  assign n5346 = x20 | n5345 ;
  assign n5347 = ( ~n5344 & n5345 ) | ( ~n5344 & n5346 ) | ( n5345 & n5346 ) ;
  assign n5348 = ( ~n5023 & n5033 ) | ( ~n5023 & n5035 ) | ( n5033 & n5035 ) ;
  assign n5349 = ( n5023 & ~n5035 ) | ( n5023 & n5348 ) | ( ~n5035 & n5348 ) ;
  assign n5350 = ( ~n5033 & n5348 ) | ( ~n5033 & n5349 ) | ( n5348 & n5349 ) ;
  assign n5351 = ( n5337 & n5347 ) | ( n5337 & n5350 ) | ( n5347 & n5350 ) ;
  assign n5352 = ~n675 & n3617 ;
  assign n5353 = n3618 | n5352 ;
  assign n5354 = ~n3431 & n5069 ;
  assign n5355 = ~n589 & n5070 ;
  assign n5356 = n5354 | n5355 ;
  assign n5357 = ~n672 & n5083 ;
  assign n5358 = n5356 | n5357 ;
  assign n5359 = n5074 | n5358 ;
  assign n5360 = ( ~n5353 & n5358 ) | ( ~n5353 & n5359 ) | ( n5358 & n5359 ) ;
  assign n5361 = ~x17 & n5360 ;
  assign n5362 = x17 | n5361 ;
  assign n5363 = ( ~n5360 & n5361 ) | ( ~n5360 & n5362 ) | ( n5361 & n5362 ) ;
  assign n5364 = ( n4815 & ~n5036 ) | ( n4815 & n5050 ) | ( ~n5036 & n5050 ) ;
  assign n5365 = ( ~n4815 & n5036 ) | ( ~n4815 & n5364 ) | ( n5036 & n5364 ) ;
  assign n5366 = ( ~n5050 & n5364 ) | ( ~n5050 & n5365 ) | ( n5364 & n5365 ) ;
  assign n5367 = ( n5351 & n5363 ) | ( n5351 & n5366 ) | ( n5363 & n5366 ) ;
  assign n5368 = n5096 & n5367 ;
  assign n5369 = n5096 | n5367 ;
  assign n5370 = ~n5368 & n5369 ;
  assign n5371 = n4811 & ~n5051 ;
  assign n5372 = n5052 | n5371 ;
  assign n5373 = n5370 & ~n5372 ;
  assign n5374 = n5368 | n5373 ;
  assign n5375 = n5082 & n5374 ;
  assign n5376 = n5082 | n5374 ;
  assign n5377 = ~n5375 & n5376 ;
  assign n5378 = ~n5370 & n5372 ;
  assign n5379 = n5373 | n5378 ;
  assign n5380 = ~x12 & x13 ;
  assign n5381 = x12 & ~x13 ;
  assign n5382 = n5380 | n5381 ;
  assign n5383 = ~n35 & n38 ;
  assign n5384 = ~n5382 & n5383 ;
  assign n5385 = n39 | n5384 ;
  assign n5386 = ~n3634 & n5385 ;
  assign n5387 = n672 & n5384 ;
  assign n5388 = ( ~n672 & n5386 ) | ( ~n672 & n5387 ) | ( n5386 & n5387 ) ;
  assign n5389 = ( ~n3619 & n5386 ) | ( ~n3619 & n5388 ) | ( n5386 & n5388 ) ;
  assign n5390 = ~x14 & n5389 ;
  assign n5391 = x14 | n5390 ;
  assign n5392 = ( ~n5389 & n5390 ) | ( ~n5389 & n5391 ) | ( n5390 & n5391 ) ;
  assign n5393 = n5111 | n5335 ;
  assign n5394 = ~n5336 & n5393 ;
  assign n5395 = ~n1014 & n4776 ;
  assign n5396 = n904 & n4778 ;
  assign n5397 = n5395 | n5396 ;
  assign n5398 = n778 & n4781 ;
  assign n5399 = n5397 | n5398 ;
  assign n5400 = n4784 | n5399 ;
  assign n5401 = ( ~n4535 & n5399 ) | ( ~n4535 & n5400 ) | ( n5399 & n5400 ) ;
  assign n5402 = ~x20 & n5401 ;
  assign n5403 = x20 | n5402 ;
  assign n5404 = ( ~n5401 & n5402 ) | ( ~n5401 & n5403 ) | ( n5402 & n5403 ) ;
  assign n5405 = n5394 & n5404 ;
  assign n5406 = n5394 | n5404 ;
  assign n5407 = ~n5405 & n5406 ;
  assign n5408 = n5130 | n5309 ;
  assign n5409 = ~n5310 & n5408 ;
  assign n5410 = ~n1411 & n4481 ;
  assign n5411 = n4479 | n5410 ;
  assign n5412 = ( n1532 & n5410 ) | ( n1532 & n5411 ) | ( n5410 & n5411 ) ;
  assign n5413 = n3178 & n4484 ;
  assign n5414 = n5412 | n5413 ;
  assign n5415 = n4487 | n5414 ;
  assign n5416 = ( ~n3750 & n5414 ) | ( ~n3750 & n5415 ) | ( n5414 & n5415 ) ;
  assign n5417 = ~x26 & n5416 ;
  assign n5418 = x26 | n5417 ;
  assign n5419 = ( ~n5416 & n5417 ) | ( ~n5416 & n5418 ) | ( n5417 & n5418 ) ;
  assign n5420 = n5409 & n5419 ;
  assign n5421 = n5409 | n5419 ;
  assign n5422 = ~n5420 & n5421 ;
  assign n5423 = n5304 & ~n5308 ;
  assign n5424 = n5307 & ~n5308 ;
  assign n5425 = n5423 | n5424 ;
  assign n5426 = ~n1733 & n4043 ;
  assign n5427 = n1625 & n4045 ;
  assign n5428 = n5426 | n5427 ;
  assign n5429 = n3030 & n4048 ;
  assign n5430 = n5428 | n5429 ;
  assign n5431 = n4051 | n5430 ;
  assign n5432 = ( ~n4578 & n5430 ) | ( ~n4578 & n5431 ) | ( n5430 & n5431 ) ;
  assign n5433 = ~x29 & n5432 ;
  assign n5434 = x29 | n5433 ;
  assign n5435 = ( ~n5432 & n5433 ) | ( ~n5432 & n5434 ) | ( n5433 & n5434 ) ;
  assign n5436 = n1532 & n4481 ;
  assign n5437 = ~n1411 & n4484 ;
  assign n5438 = ~n2939 & n4479 ;
  assign n5439 = n5437 | n5438 ;
  assign n5440 = n5436 | n5439 ;
  assign n5441 = n4487 | n5440 ;
  assign n5442 = ( ~n3930 & n5440 ) | ( ~n3930 & n5441 ) | ( n5440 & n5441 ) ;
  assign n5443 = ~x26 & n5442 ;
  assign n5444 = x26 | n5443 ;
  assign n5445 = ( ~n5442 & n5443 ) | ( ~n5442 & n5444 ) | ( n5443 & n5444 ) ;
  assign n5446 = ( n5425 & n5435 ) | ( n5425 & n5445 ) | ( n5435 & n5445 ) ;
  assign n5447 = n5422 & n5446 ;
  assign n5448 = n5420 | n5447 ;
  assign n5449 = n1327 & n4546 ;
  assign n5450 = ~n1151 & n4548 ;
  assign n5451 = n5449 | n5450 ;
  assign n5452 = n1233 & n4551 ;
  assign n5453 = n5451 | n5452 ;
  assign n5454 = n4554 | n5453 ;
  assign n5455 = ( ~n4615 & n5453 ) | ( ~n4615 & n5454 ) | ( n5453 & n5454 ) ;
  assign n5456 = ~x23 & n5455 ;
  assign n5457 = x23 | n5456 ;
  assign n5458 = ( ~n5455 & n5456 ) | ( ~n5455 & n5457 ) | ( n5456 & n5457 ) ;
  assign n5459 = ( n5113 & n5321 ) | ( n5113 & ~n5322 ) | ( n5321 & ~n5322 ) ;
  assign n5460 = ( n5311 & ~n5322 ) | ( n5311 & n5459 ) | ( ~n5322 & n5459 ) ;
  assign n5461 = ( n5448 & n5458 ) | ( n5448 & n5460 ) | ( n5458 & n5460 ) ;
  assign n5462 = ~n1014 & n4778 ;
  assign n5463 = ~n3255 & n4776 ;
  assign n5464 = n5462 | n5463 ;
  assign n5465 = n904 & n4781 ;
  assign n5466 = n5464 | n5465 ;
  assign n5467 = n4784 | n5466 ;
  assign n5468 = ( n4632 & n5466 ) | ( n4632 & n5467 ) | ( n5466 & n5467 ) ;
  assign n5469 = x20 & n5468 ;
  assign n5470 = x20 & ~n5469 ;
  assign n5471 = ( n5468 & ~n5469 ) | ( n5468 & n5470 ) | ( ~n5469 & n5470 ) ;
  assign n5472 = ( ~n5322 & n5332 ) | ( ~n5322 & n5334 ) | ( n5332 & n5334 ) ;
  assign n5473 = ( n5322 & ~n5334 ) | ( n5322 & n5472 ) | ( ~n5334 & n5472 ) ;
  assign n5474 = ( ~n5332 & n5472 ) | ( ~n5332 & n5473 ) | ( n5472 & n5473 ) ;
  assign n5475 = ( n5461 & n5471 ) | ( n5461 & n5474 ) | ( n5471 & n5474 ) ;
  assign n5476 = n5407 & n5475 ;
  assign n5477 = n5405 | n5476 ;
  assign n5478 = n3504 & n5069 ;
  assign n5479 = ~n3431 & n5070 ;
  assign n5480 = n5478 | n5479 ;
  assign n5481 = ~n589 & n5083 ;
  assign n5482 = n5480 | n5481 ;
  assign n5483 = n5074 | n5482 ;
  assign n5484 = ( n4765 & n5482 ) | ( n4765 & n5483 ) | ( n5482 & n5483 ) ;
  assign n5485 = x17 & n5484 ;
  assign n5486 = x17 & ~n5485 ;
  assign n5487 = ( n5484 & ~n5485 ) | ( n5484 & n5486 ) | ( ~n5485 & n5486 ) ;
  assign n5488 = ( ~n5337 & n5347 ) | ( ~n5337 & n5350 ) | ( n5347 & n5350 ) ;
  assign n5489 = ( n5337 & ~n5350 ) | ( n5337 & n5488 ) | ( ~n5350 & n5488 ) ;
  assign n5490 = ( ~n5347 & n5488 ) | ( ~n5347 & n5489 ) | ( n5488 & n5489 ) ;
  assign n5491 = ( n5477 & n5487 ) | ( n5477 & n5490 ) | ( n5487 & n5490 ) ;
  assign n5492 = ( ~n5351 & n5363 ) | ( ~n5351 & n5366 ) | ( n5363 & n5366 ) ;
  assign n5493 = ( n5351 & ~n5366 ) | ( n5351 & n5492 ) | ( ~n5366 & n5492 ) ;
  assign n5494 = ( ~n5363 & n5492 ) | ( ~n5363 & n5493 ) | ( n5492 & n5493 ) ;
  assign n5495 = ( n5392 & n5491 ) | ( n5392 & n5494 ) | ( n5491 & n5494 ) ;
  assign n5496 = ~n5379 & n5495 ;
  assign n5497 = x7 & ~x8 ;
  assign n5498 = ~x7 & x8 ;
  assign n5499 = n5497 | n5498 ;
  assign n5500 = x5 & ~x6 ;
  assign n5501 = ~x5 & x6 ;
  assign n5502 = n5500 | n5501 ;
  assign n5503 = ~n5499 & n5502 ;
  assign n5504 = ~n3634 & n5503 ;
  assign n5505 = ~x6 & x7 ;
  assign n5506 = x6 & ~x7 ;
  assign n5507 = n5505 | n5506 ;
  assign n5508 = ~n5502 & n5507 ;
  assign n5509 = ~n672 & n5508 ;
  assign n5510 = n5504 | n5509 ;
  assign n5511 = n5499 & ~n5502 ;
  assign n5512 = ~n5507 & n5511 ;
  assign n5513 = ~n589 & n5512 ;
  assign n5514 = n5510 | n5513 ;
  assign n5515 = n5499 & n5502 ;
  assign n5516 = n5514 | n5515 ;
  assign n5517 = ( ~n5092 & n5514 ) | ( ~n5092 & n5516 ) | ( n5514 & n5516 ) ;
  assign n5518 = ~x8 & n5517 ;
  assign n5519 = x8 | n5518 ;
  assign n5520 = ( ~n5517 & n5518 ) | ( ~n5517 & n5519 ) | ( n5518 & n5519 ) ;
  assign n5521 = ~n2375 & n3744 ;
  assign n5522 = ~n2455 & n3727 ;
  assign n5523 = ~n2606 & n3639 ;
  assign n5524 = n5522 | n5523 ;
  assign n5525 = n5521 | n5524 ;
  assign n5526 = ( n2375 & ~n2455 ) | ( n2375 & n2773 ) | ( ~n2455 & n2773 ) ;
  assign n5527 = ( ~n2375 & n2455 ) | ( ~n2375 & n5526 ) | ( n2455 & n5526 ) ;
  assign n5528 = ( ~n2773 & n5526 ) | ( ~n2773 & n5527 ) | ( n5526 & n5527 ) ;
  assign n5529 = n3636 | n5525 ;
  assign n5530 = ( n5525 & ~n5528 ) | ( n5525 & n5529 ) | ( ~n5528 & n5529 ) ;
  assign n5531 = n678 | n2989 ;
  assign n5532 = n81 | n514 ;
  assign n5533 = n2002 | n5532 ;
  assign n5534 = n265 | n349 ;
  assign n5535 = n5533 | n5534 ;
  assign n5536 = n5531 | n5535 ;
  assign n5537 = n3467 | n5536 ;
  assign n5538 = n2206 | n5537 ;
  assign n5539 = n4290 | n5538 ;
  assign n5540 = n4289 & ~n5539 ;
  assign n5541 = n2164 | n3204 ;
  assign n5542 = n1297 | n5541 ;
  assign n5543 = n655 | n3243 ;
  assign n5544 = n513 | n5543 ;
  assign n5545 = n5542 | n5544 ;
  assign n5546 = n199 | n570 ;
  assign n5547 = n94 | n5546 ;
  assign n5548 = n5545 | n5547 ;
  assign n5549 = n2602 | n2810 ;
  assign n5550 = n152 | n5549 ;
  assign n5551 = n1548 | n1956 ;
  assign n5552 = n5550 | n5551 ;
  assign n5553 = n291 | n669 ;
  assign n5554 = n1865 | n5553 ;
  assign n5555 = n377 | n5554 ;
  assign n5556 = n4235 | n5555 ;
  assign n5557 = n5552 | n5556 ;
  assign n5558 = n127 | n996 ;
  assign n5559 = n482 | n5558 ;
  assign n5560 = n625 | n5559 ;
  assign n5561 = n633 | n5560 ;
  assign n5562 = n5557 | n5561 ;
  assign n5563 = n346 | n384 ;
  assign n5564 = n212 | n5563 ;
  assign n5565 = n434 | n5564 ;
  assign n5566 = n77 | n5565 ;
  assign n5567 = n110 | n5566 ;
  assign n5568 = n5562 | n5567 ;
  assign n5569 = n5548 | n5568 ;
  assign n5570 = n5540 & ~n5569 ;
  assign n5571 = n300 | n636 ;
  assign n5572 = n366 | n5571 ;
  assign n5573 = ( n120 & ~n1504 ) | ( n120 & n5572 ) | ( ~n1504 & n5572 ) ;
  assign n5574 = n1504 | n5573 ;
  assign n5575 = n5570 & ~n5574 ;
  assign n5576 = n5530 & ~n5575 ;
  assign n5577 = n5530 & ~n5576 ;
  assign n5578 = n5530 | n5575 ;
  assign n5579 = ~n5577 & n5578 ;
  assign n5580 = n2569 & n3744 ;
  assign n5581 = ~n2672 & n2764 ;
  assign n5582 = n2569 | n5581 ;
  assign n5583 = n2569 & n5581 ;
  assign n5584 = n5582 & ~n5583 ;
  assign n5585 = ~n2764 & n3639 ;
  assign n5586 = ~n2672 & n3727 ;
  assign n5587 = n5585 | n5586 ;
  assign n5588 = n3636 | n5587 ;
  assign n5589 = ( n5584 & n5587 ) | ( n5584 & n5588 ) | ( n5587 & n5588 ) ;
  assign n5590 = n5580 | n5589 ;
  assign n5591 = n367 | n1352 ;
  assign n5592 = n428 | n640 ;
  assign n5593 = n5591 | n5592 ;
  assign n5594 = n321 | n346 ;
  assign n5595 = n1404 | n5594 ;
  assign n5596 = n3073 | n5595 ;
  assign n5597 = n1024 | n1636 ;
  assign n5598 = n5596 | n5597 ;
  assign n5599 = n5593 | n5598 ;
  assign n5600 = n345 | n444 ;
  assign n5601 = n3149 | n5600 ;
  assign n5602 = n190 | n434 ;
  assign n5603 = n458 | n5602 ;
  assign n5604 = n5601 | n5603 ;
  assign n5605 = n186 | n5604 ;
  assign n5606 = n3314 | n5605 ;
  assign n5607 = n5599 | n5606 ;
  assign n5608 = n1354 | n1425 ;
  assign n5609 = n530 | n5608 ;
  assign n5610 = n280 | n5609 ;
  assign n5611 = n5607 | n5610 ;
  assign n5612 = n130 | n381 ;
  assign n5613 = n180 | n5612 ;
  assign n5614 = n645 | n5613 ;
  assign n5615 = n878 | n1094 ;
  assign n5616 = n5614 | n5615 ;
  assign n5617 = n283 | n315 ;
  assign n5618 = n309 | n5617 ;
  assign n5619 = ( n160 & ~n3564 ) | ( n160 & n5618 ) | ( ~n3564 & n5618 ) ;
  assign n5620 = n3564 | n5619 ;
  assign n5621 = n5616 | n5620 ;
  assign n5622 = n2049 & ~n5621 ;
  assign n5623 = ~n5611 & n5622 ;
  assign n5624 = n4274 | n4925 ;
  assign n5625 = n96 | n102 ;
  assign n5626 = n114 | n646 ;
  assign n5627 = n5625 | n5626 ;
  assign n5628 = n1032 | n1051 ;
  assign n5629 = n5627 | n5628 ;
  assign n5630 = n5624 | n5629 ;
  assign n5631 = n433 | n1315 ;
  assign n5632 = n755 | n5631 ;
  assign n5633 = n5630 | n5632 ;
  assign n5634 = n243 | n2810 ;
  assign n5635 = n592 | n5634 ;
  assign n5636 = n602 | n5635 ;
  assign n5637 = n450 | n5636 ;
  assign n5638 = n5633 | n5637 ;
  assign n5639 = n142 | n442 ;
  assign n5640 = n5638 | n5639 ;
  assign n5641 = n2411 | n2612 ;
  assign n5642 = n484 | n529 ;
  assign n5643 = n344 | n5642 ;
  assign n5644 = n5641 | n5643 ;
  assign n5645 = n393 | n435 ;
  assign n5646 = n85 | n5645 ;
  assign n5647 = n5644 | n5646 ;
  assign n5648 = n5640 | n5647 ;
  assign n5649 = n5623 & ~n5648 ;
  assign n5650 = n1647 | n2163 ;
  assign n5651 = n960 | n5650 ;
  assign n5652 = n1310 | n5651 ;
  assign n5653 = n958 | n5652 ;
  assign n5654 = n1022 | n5653 ;
  assign n5655 = n475 | n5654 ;
  assign n5656 = n655 | n5655 ;
  assign n5657 = n511 | n5656 ;
  assign n5658 = n5649 & ~n5657 ;
  assign n5659 = n277 | n519 ;
  assign n5660 = n300 | n5659 ;
  assign n5661 = n384 | n5660 ;
  assign n5662 = n570 | n5661 ;
  assign n5663 = n5658 & ~n5662 ;
  assign n5664 = n888 | n2527 ;
  assign n5665 = n1567 | n5664 ;
  assign n5666 = n355 | n3375 ;
  assign n5667 = n226 & ~n5666 ;
  assign n5668 = ~n5665 & n5667 ;
  assign n5669 = n165 | n645 ;
  assign n5670 = n5668 & ~n5669 ;
  assign n5671 = n653 | n2041 ;
  assign n5672 = n2305 | n5671 ;
  assign n5673 = n92 | n390 ;
  assign n5674 = n728 | n5673 ;
  assign n5675 = n1240 | n5674 ;
  assign n5676 = n5672 | n5675 ;
  assign n5677 = n59 | n1791 ;
  assign n5678 = n5676 | n5677 ;
  assign n5679 = n5670 & ~n5678 ;
  assign n5680 = n130 | n1034 ;
  assign n5681 = n1128 | n5680 ;
  assign n5682 = n237 | n5681 ;
  assign n5683 = n283 | n5682 ;
  assign n5684 = n607 | n5683 ;
  assign n5685 = n5679 & ~n5684 ;
  assign n5686 = n83 | n434 ;
  assign n5687 = n99 | n5686 ;
  assign n5688 = n5685 & ~n5687 ;
  assign n5689 = n270 | n452 ;
  assign n5690 = n1260 | n5689 ;
  assign n5691 = n1381 | n5690 ;
  assign n5692 = n1565 | n5691 ;
  assign n5693 = n2543 | n5692 ;
  assign n5694 = n1978 | n5693 ;
  assign n5695 = n1970 | n5694 ;
  assign n5696 = n5688 & ~n5695 ;
  assign n5697 = n476 | n520 ;
  assign n5698 = n2411 | n5697 ;
  assign n5699 = n277 | n419 ;
  assign n5700 = n358 | n5699 ;
  assign n5701 = n5698 | n5700 ;
  assign n5702 = n125 | n198 ;
  assign n5703 = n215 | n5702 ;
  assign n5704 = n807 | n5703 ;
  assign n5705 = n5701 | n5704 ;
  assign n5706 = n435 | n5705 ;
  assign n5707 = n77 | n5706 ;
  assign n5708 = n155 | n5707 ;
  assign n5709 = n160 | n5708 ;
  assign n5710 = n640 | n5709 ;
  assign n5711 = n5696 & ~n5710 ;
  assign n5712 = ~n224 & n5711 ;
  assign n5713 = n5663 | n5712 ;
  assign n5714 = n5590 & ~n5713 ;
  assign n5715 = n2609 & n2766 ;
  assign n5716 = n2767 & ~n5715 ;
  assign n5717 = ~n2606 & n3744 ;
  assign n5718 = ~n2672 & n3639 ;
  assign n5719 = n5717 | n5718 ;
  assign n5720 = n2569 & n3727 ;
  assign n5721 = n5719 | n5720 ;
  assign n5722 = n3636 | n5721 ;
  assign n5723 = ( n5716 & n5721 ) | ( n5716 & n5722 ) | ( n5721 & n5722 ) ;
  assign n5724 = n5590 & ~n5663 ;
  assign n5725 = n5712 & ~n5724 ;
  assign n5726 = n5714 | n5725 ;
  assign n5727 = n5723 & ~n5726 ;
  assign n5728 = n5714 | n5727 ;
  assign n5729 = ( ~n2767 & n2770 ) | ( ~n2767 & n2771 ) | ( n2770 & n2771 ) ;
  assign n5730 = n2607 | n2770 ;
  assign n5731 = n2767 & ~n5730 ;
  assign n5732 = n5729 | n5731 ;
  assign n5733 = ~n2455 & n3744 ;
  assign n5734 = ~n2606 & n3727 ;
  assign n5735 = n2569 & n3639 ;
  assign n5736 = n5734 | n5735 ;
  assign n5737 = n5733 | n5736 ;
  assign n5738 = n3636 | n5737 ;
  assign n5739 = ( ~n5732 & n5737 ) | ( ~n5732 & n5738 ) | ( n5737 & n5738 ) ;
  assign n5740 = n327 | n483 ;
  assign n5741 = n597 | n5740 ;
  assign n5742 = n512 | n749 ;
  assign n5743 = n5741 | n5742 ;
  assign n5744 = n530 | n2951 ;
  assign n5745 = n5743 | n5744 ;
  assign n5746 = n490 | n628 ;
  assign n5747 = n669 | n5746 ;
  assign n5748 = n321 | n5747 ;
  assign n5749 = n582 | n5748 ;
  assign n5750 = n5745 | n5749 ;
  assign n5751 = n100 | n5750 ;
  assign n5752 = n146 | n237 ;
  assign n5753 = n206 | n5752 ;
  assign n5754 = n169 | n449 ;
  assign n5755 = n5753 | n5754 ;
  assign n5756 = n122 | n5755 ;
  assign n5757 = n181 | n505 ;
  assign n5758 = n443 | n5757 ;
  assign n5759 = n1536 | n5758 ;
  assign n5760 = n3809 | n5627 ;
  assign n5761 = n5759 | n5760 ;
  assign n5762 = n5756 | n5761 ;
  assign n5763 = n2145 | n5762 ;
  assign n5764 = n5751 | n5763 ;
  assign n5765 = n1045 | n5764 ;
  assign n5766 = n2140 | n5765 ;
  assign n5767 = n130 | n144 ;
  assign n5768 = n1354 | n5767 ;
  assign n5769 = n421 | n5768 ;
  assign n5770 = n1656 | n5769 ;
  assign n5771 = n636 | n5770 ;
  assign n5772 = n338 | n5771 ;
  assign n5773 = n379 | n5772 ;
  assign n5774 = n591 | n5773 ;
  assign n5775 = n5766 | n5774 ;
  assign n5776 = n1153 | n5775 ;
  assign n5777 = ( n5728 & n5739 ) | ( n5728 & n5776 ) | ( n5739 & n5776 ) ;
  assign n5778 = ~n5579 & n5777 ;
  assign n5779 = n5576 | n5778 ;
  assign n5780 = n2378 & n2774 ;
  assign n5781 = n2775 & ~n5780 ;
  assign n5782 = n2296 & n3744 ;
  assign n5783 = ~n2375 & n3727 ;
  assign n5784 = ~n2455 & n3639 ;
  assign n5785 = n5783 | n5784 ;
  assign n5786 = n5782 | n5785 ;
  assign n5787 = n3636 | n5786 ;
  assign n5788 = ( n5781 & n5786 ) | ( n5781 & n5787 ) | ( n5786 & n5787 ) ;
  assign n5789 = n801 | n1682 ;
  assign n5790 = n3508 | n5789 ;
  assign n5791 = n306 | n654 ;
  assign n5792 = n1371 | n5791 ;
  assign n5793 = n1636 | n5792 ;
  assign n5794 = n5790 | n5793 ;
  assign n5795 = n273 | n293 ;
  assign n5796 = n1311 | n5795 ;
  assign n5797 = n81 | n203 ;
  assign n5798 = n5796 | n5797 ;
  assign n5799 = n1271 | n5798 ;
  assign n5800 = n5794 | n5799 ;
  assign n5801 = n1657 | n5800 ;
  assign n5802 = n3230 | n5801 ;
  assign n5803 = n3864 | n5802 ;
  assign n5804 = n291 | n619 ;
  assign n5805 = n99 | n5804 ;
  assign n5806 = n4097 | n5805 ;
  assign n5807 = n439 | n878 ;
  assign n5808 = n5806 | n5807 ;
  assign n5809 = n5605 | n5808 ;
  assign n5810 = n430 | n3243 ;
  assign n5811 = n245 | n5810 ;
  assign n5812 = n500 | n5811 ;
  assign n5813 = n504 | n5812 ;
  assign n5814 = n5809 | n5813 ;
  assign n5815 = n260 | n384 ;
  assign n5816 = n167 | n5815 ;
  assign n5817 = n218 | n5816 ;
  assign n5818 = n5814 | n5817 ;
  assign n5819 = n4126 | n5818 ;
  assign n5820 = n5803 | n5819 ;
  assign n5821 = n253 | n539 ;
  assign n5822 = n66 | n1194 ;
  assign n5823 = ( n531 & ~n5821 ) | ( n531 & n5822 ) | ( ~n5821 & n5822 ) ;
  assign n5824 = n5821 | n5823 ;
  assign n5825 = ( n90 & ~n2547 ) | ( n90 & n5824 ) | ( ~n2547 & n5824 ) ;
  assign n5826 = n2547 | n5825 ;
  assign n5827 = n5820 | n5826 ;
  assign n5828 = n5788 & n5827 ;
  assign n5829 = n5788 & ~n5828 ;
  assign n5830 = ~n5788 & n5827 ;
  assign n5831 = n5829 | n5830 ;
  assign n5832 = n5779 & n5831 ;
  assign n5833 = n5779 | n5831 ;
  assign n5834 = ~n5832 & n5833 ;
  assign n5835 = n2106 & ~n2778 ;
  assign n5836 = n2779 | n5835 ;
  assign n5837 = n2193 & n4043 ;
  assign n5838 = n2013 & n4045 ;
  assign n5839 = n5837 | n5838 ;
  assign n5840 = ~n2103 & n4048 ;
  assign n5841 = n5839 | n5840 ;
  assign n5842 = n4051 | n5841 ;
  assign n5843 = ( ~n5836 & n5841 ) | ( ~n5836 & n5842 ) | ( n5841 & n5842 ) ;
  assign n5844 = ~x29 & n5843 ;
  assign n5845 = x29 | n5844 ;
  assign n5846 = ( ~n5843 & n5844 ) | ( ~n5843 & n5845 ) | ( n5844 & n5845 ) ;
  assign n5847 = n5834 & n5846 ;
  assign n5848 = n5834 | n5846 ;
  assign n5849 = ~n5847 & n5848 ;
  assign n5850 = n5777 & ~n5778 ;
  assign n5851 = n5579 | n5778 ;
  assign n5852 = ~n5850 & n5851 ;
  assign n5853 = n2296 & n4043 ;
  assign n5854 = n2193 & n4045 ;
  assign n5855 = n5853 | n5854 ;
  assign n5856 = n2013 & n4048 ;
  assign n5857 = n5855 | n5856 ;
  assign n5858 = n4051 | n5857 ;
  assign n5859 = ( n5216 & n5857 ) | ( n5216 & n5858 ) | ( n5857 & n5858 ) ;
  assign n5860 = x29 & n5859 ;
  assign n5861 = x29 & ~n5860 ;
  assign n5862 = ( n5859 & ~n5860 ) | ( n5859 & n5861 ) | ( ~n5860 & n5861 ) ;
  assign n5863 = ~n5852 & n5862 ;
  assign n5864 = n5739 & n5776 ;
  assign n5865 = n5739 & ~n5864 ;
  assign n5866 = ~n5739 & n5776 ;
  assign n5867 = n5865 | n5866 ;
  assign n5868 = n5728 | n5867 ;
  assign n5869 = ~n5867 & n5868 ;
  assign n5870 = ( ~n5728 & n5868 ) | ( ~n5728 & n5869 ) | ( n5868 & n5869 ) ;
  assign n5871 = ~n2375 & n4043 ;
  assign n5872 = n2296 & n4045 ;
  assign n5873 = n5871 | n5872 ;
  assign n5874 = n2193 & n4048 ;
  assign n5875 = n5873 | n5874 ;
  assign n5876 = n4051 | n5875 ;
  assign n5877 = ( n2193 & ~n2296 ) | ( n2193 & n2776 ) | ( ~n2296 & n2776 ) ;
  assign n5878 = ( ~n2193 & n2296 ) | ( ~n2193 & n5877 ) | ( n2296 & n5877 ) ;
  assign n5879 = ( ~n2776 & n5877 ) | ( ~n2776 & n5878 ) | ( n5877 & n5878 ) ;
  assign n5880 = ( n5875 & n5876 ) | ( n5875 & ~n5879 ) | ( n5876 & ~n5879 ) ;
  assign n5881 = ~x29 & n5880 ;
  assign n5882 = x29 | n5881 ;
  assign n5883 = ( ~n5880 & n5881 ) | ( ~n5880 & n5882 ) | ( n5881 & n5882 ) ;
  assign n5884 = n5870 & n5883 ;
  assign n5885 = n5870 & ~n5884 ;
  assign n5886 = ~n5870 & n5883 ;
  assign n5887 = n5885 | n5886 ;
  assign n5888 = ~n2455 & n4043 ;
  assign n5889 = ~n2375 & n4045 ;
  assign n5890 = n5888 | n5889 ;
  assign n5891 = n2296 & n4048 ;
  assign n5892 = n5890 | n5891 ;
  assign n5893 = n4051 | n5892 ;
  assign n5894 = ( n5781 & n5892 ) | ( n5781 & n5893 ) | ( n5892 & n5893 ) ;
  assign n5895 = x29 & n5894 ;
  assign n5896 = x29 & ~n5895 ;
  assign n5897 = ( n5894 & ~n5895 ) | ( n5894 & n5896 ) | ( ~n5895 & n5896 ) ;
  assign n5898 = n5723 & ~n5727 ;
  assign n5899 = n5726 | n5727 ;
  assign n5900 = ~n5898 & n5899 ;
  assign n5901 = n5897 & ~n5900 ;
  assign n5902 = n5897 & ~n5901 ;
  assign n5903 = n5897 | n5900 ;
  assign n5904 = ~n5902 & n5903 ;
  assign n5905 = ~n2606 & n4043 ;
  assign n5906 = ~n2455 & n4045 ;
  assign n5907 = n5905 | n5906 ;
  assign n5908 = ~n2375 & n4048 ;
  assign n5909 = n5907 | n5908 ;
  assign n5910 = n4051 | n5909 ;
  assign n5911 = ( ~n5528 & n5909 ) | ( ~n5528 & n5910 ) | ( n5909 & n5910 ) ;
  assign n5912 = ~x29 & n5911 ;
  assign n5913 = x29 & ~n5911 ;
  assign n5914 = n5912 | n5913 ;
  assign n5915 = n5590 | n5663 ;
  assign n5916 = n5590 & n5663 ;
  assign n5917 = n5915 & ~n5916 ;
  assign n5918 = n5914 & ~n5917 ;
  assign n5919 = ~n5914 & n5917 ;
  assign n5920 = n5918 | n5919 ;
  assign n5921 = ~n2455 & n4048 ;
  assign n5922 = ~n2606 & n4045 ;
  assign n5923 = n5921 | n5922 ;
  assign n5924 = n2569 & n4043 ;
  assign n5925 = n5923 | n5924 ;
  assign n5926 = n4051 | n5925 ;
  assign n5927 = ( ~n5732 & n5925 ) | ( ~n5732 & n5926 ) | ( n5925 & n5926 ) ;
  assign n5928 = ~x29 & n5927 ;
  assign n5929 = x29 & ~n5927 ;
  assign n5930 = n5928 | n5929 ;
  assign n5931 = n2672 & ~n2764 ;
  assign n5932 = n5581 | n5931 ;
  assign n5933 = ~n2764 & n3727 ;
  assign n5934 = ~n2672 & n3744 ;
  assign n5935 = n5933 | n5934 ;
  assign n5936 = n3636 | n5935 ;
  assign n5937 = ( n5932 & n5935 ) | ( n5932 & n5936 ) | ( n5935 & n5936 ) ;
  assign n5938 = n5930 & n5937 ;
  assign n5939 = n5930 | n5937 ;
  assign n5940 = ~n5938 & n5939 ;
  assign n5941 = ~n2764 & n4043 ;
  assign n5942 = ~n2672 & n4045 ;
  assign n5943 = n5941 | n5942 ;
  assign n5944 = n2569 & n4048 ;
  assign n5945 = n5943 | n5944 ;
  assign n5946 = ( n4051 & n5584 ) | ( n4051 & n5945 ) | ( n5584 & n5945 ) ;
  assign n5947 = ( x29 & ~n5945 ) | ( x29 & n5946 ) | ( ~n5945 & n5946 ) ;
  assign n5948 = ~n5946 & n5947 ;
  assign n5949 = n5945 | n5947 ;
  assign n5950 = ( ~x29 & n5948 ) | ( ~x29 & n5949 ) | ( n5948 & n5949 ) ;
  assign n5951 = ~n2764 & n4045 ;
  assign n5952 = ~n2672 & n4048 ;
  assign n5953 = n5951 | n5952 ;
  assign n5954 = n4051 | n5953 ;
  assign n5955 = ( n5932 & n5953 ) | ( n5932 & n5954 ) | ( n5953 & n5954 ) ;
  assign n5956 = ( n400 & ~n2763 ) | ( n400 & n4041 ) | ( ~n2763 & n4041 ) ;
  assign n5957 = x29 & ~n5956 ;
  assign n5958 = ~x29 & n5955 ;
  assign n5959 = ( ~n5955 & n5957 ) | ( ~n5955 & n5958 ) | ( n5957 & n5958 ) ;
  assign n5960 = n5950 & n5959 ;
  assign n5961 = ~n2763 & n3635 ;
  assign n5962 = ~n2606 & n4048 ;
  assign n5963 = ~n2672 & n4043 ;
  assign n5964 = n5962 | n5963 ;
  assign n5965 = n2569 & n4045 ;
  assign n5966 = n5964 | n5965 ;
  assign n5967 = n4051 | n5966 ;
  assign n5968 = ( n5716 & n5966 ) | ( n5716 & n5967 ) | ( n5966 & n5967 ) ;
  assign n5969 = x29 & n5968 ;
  assign n5970 = x29 & ~n5969 ;
  assign n5971 = ( n5968 & ~n5969 ) | ( n5968 & n5970 ) | ( ~n5969 & n5970 ) ;
  assign n5972 = ( n5960 & n5961 ) | ( n5960 & n5971 ) | ( n5961 & n5971 ) ;
  assign n5973 = n5940 & n5972 ;
  assign n5974 = n5938 | n5973 ;
  assign n5975 = ~n5920 & n5974 ;
  assign n5976 = n5918 | n5975 ;
  assign n5977 = ~n5904 & n5976 ;
  assign n5978 = n5901 | n5977 ;
  assign n5979 = n5887 & n5978 ;
  assign n5980 = n5884 | n5979 ;
  assign n5981 = n5852 | n5863 ;
  assign n5982 = ( ~n5862 & n5863 ) | ( ~n5862 & n5981 ) | ( n5863 & n5981 ) ;
  assign n5983 = n5980 & ~n5982 ;
  assign n5984 = n5863 | n5983 ;
  assign n5985 = n5849 & n5984 ;
  assign n5986 = n5828 | n5832 ;
  assign n5987 = n2193 & n3744 ;
  assign n5988 = n2296 & n3727 ;
  assign n5989 = ~n2375 & n3639 ;
  assign n5990 = n5988 | n5989 ;
  assign n5991 = n5987 | n5990 ;
  assign n5992 = n3636 | n5991 ;
  assign n5993 = ( ~n5879 & n5991 ) | ( ~n5879 & n5992 ) | ( n5991 & n5992 ) ;
  assign n5994 = n2474 | n4004 ;
  assign n5995 = n3903 | n5994 ;
  assign n5996 = n3819 | n5995 ;
  assign n5997 = n515 | n5996 ;
  assign n5998 = n2861 | n5997 ;
  assign n5999 = n1316 | n1352 ;
  assign n6000 = n251 | n5999 ;
  assign n6001 = n718 | n6000 ;
  assign n6002 = n472 | n6001 ;
  assign n6003 = n511 | n6002 ;
  assign n6004 = n5998 | n6003 ;
  assign n6005 = n212 | n262 ;
  assign n6006 = n601 | n6005 ;
  assign n6007 = n6004 | n6006 ;
  assign n6008 = n237 | n530 ;
  assign n6009 = n457 | n661 ;
  assign n6010 = n6008 | n6009 ;
  assign n6011 = n868 | n1204 ;
  assign n6012 = n4913 | n6011 ;
  assign n6013 = n6010 | n6012 ;
  assign n6014 = n350 | n416 ;
  assign n6015 = n4327 | n6014 ;
  assign n6016 = n224 | n6015 ;
  assign n6017 = n1657 | n6016 ;
  assign n6018 = n6013 | n6017 ;
  assign n6019 = n3990 | n6018 ;
  assign n6020 = n3953 | n6019 ;
  assign n6021 = n3989 | n6020 ;
  assign n6022 = n6007 | n6021 ;
  assign n6023 = n611 | n1115 ;
  assign n6024 = n348 | n6023 ;
  assign n6025 = n479 | n6024 ;
  assign n6026 = n269 | n6025 ;
  assign n6027 = n203 | n6026 ;
  assign n6028 = n404 | n6027 ;
  assign n6029 = n108 | n6028 ;
  assign n6030 = n6022 | n6029 ;
  assign n6031 = n5993 & n6030 ;
  assign n6032 = n5993 & ~n6031 ;
  assign n6033 = ~n5993 & n6030 ;
  assign n6034 = n6032 | n6033 ;
  assign n6035 = n5986 & n6034 ;
  assign n6036 = n5986 | n6034 ;
  assign n6037 = ~n6035 & n6036 ;
  assign n6038 = ( n2779 & n2784 ) | ( n2779 & n2785 ) | ( n2784 & n2785 ) ;
  assign n6039 = n2104 | n2784 ;
  assign n6040 = n2779 | n6039 ;
  assign n6041 = ~n6038 & n6040 ;
  assign n6042 = n2013 & n4043 ;
  assign n6043 = ~n2103 & n4045 ;
  assign n6044 = n6042 | n6043 ;
  assign n6045 = ~n1944 & n4048 ;
  assign n6046 = n6044 | n6045 ;
  assign n6047 = n4051 | n6046 ;
  assign n6048 = ( n6041 & n6046 ) | ( n6041 & n6047 ) | ( n6046 & n6047 ) ;
  assign n6049 = x29 & n6048 ;
  assign n6050 = x29 & ~n6049 ;
  assign n6051 = ( n6048 & ~n6049 ) | ( n6048 & n6050 ) | ( ~n6049 & n6050 ) ;
  assign n6052 = n6037 & n6051 ;
  assign n6053 = n6037 | n6051 ;
  assign n6054 = ~n6052 & n6053 ;
  assign n6055 = ( n5847 & n5985 ) | ( n5847 & n6054 ) | ( n5985 & n6054 ) ;
  assign n6056 = ( n5216 & n5265 ) | ( n5216 & n5266 ) | ( n5265 & n5266 ) ;
  assign n6057 = ( n5216 & n5268 ) | ( n5216 & n5271 ) | ( n5268 & n5271 ) ;
  assign n6058 = n6056 & ~n6057 ;
  assign n6059 = n5260 & ~n5273 ;
  assign n6060 = n6058 | n6059 ;
  assign n6061 = n6031 | n6060 ;
  assign n6062 = n6035 | n6061 ;
  assign n6063 = ( n6031 & n6035 ) | ( n6031 & n6060 ) | ( n6035 & n6060 ) ;
  assign n6064 = n6062 & ~n6063 ;
  assign n6065 = ~n2103 & n4043 ;
  assign n6066 = ~n1944 & n4045 ;
  assign n6067 = n6065 | n6066 ;
  assign n6068 = ~n1880 & n4048 ;
  assign n6069 = n6067 | n6068 ;
  assign n6070 = n4051 | n6069 ;
  assign n6071 = ( ~n5281 & n6069 ) | ( ~n5281 & n6070 ) | ( n6069 & n6070 ) ;
  assign n6072 = ~x29 & n6071 ;
  assign n6073 = x29 | n6072 ;
  assign n6074 = ( ~n6071 & n6072 ) | ( ~n6071 & n6073 ) | ( n6072 & n6073 ) ;
  assign n6075 = n6064 & n6074 ;
  assign n6076 = n6064 | n6074 ;
  assign n6077 = ~n6075 & n6076 ;
  assign n6078 = n6052 | n6077 ;
  assign n6079 = n6055 | n6078 ;
  assign n6080 = ( n6052 & n6055 ) | ( n6052 & n6077 ) | ( n6055 & n6077 ) ;
  assign n6081 = n6079 & ~n6080 ;
  assign n6082 = n1803 & n4479 ;
  assign n6083 = ~n2873 & n4481 ;
  assign n6084 = n6082 | n6083 ;
  assign n6085 = ~n1733 & n4484 ;
  assign n6086 = n6084 | n6085 ;
  assign n6087 = n4487 | n6086 ;
  assign n6088 = ( ~n4985 & n6086 ) | ( ~n4985 & n6087 ) | ( n6086 & n6087 ) ;
  assign n6089 = ~x26 & n6088 ;
  assign n6090 = x26 | n6089 ;
  assign n6091 = ( ~n6088 & n6089 ) | ( ~n6088 & n6090 ) | ( n6089 & n6090 ) ;
  assign n6092 = n6081 & n6091 ;
  assign n6093 = n6081 | n6091 ;
  assign n6094 = ~n6092 & n6093 ;
  assign n6095 = ( n5847 & n5848 ) | ( n5847 & n5984 ) | ( n5848 & n5984 ) ;
  assign n6096 = n6054 | n6095 ;
  assign n6097 = ~n6055 & n6096 ;
  assign n6098 = ~n2873 & n4484 ;
  assign n6099 = n1803 & n4481 ;
  assign n6100 = n6098 | n6099 ;
  assign n6101 = ~n1880 & n4479 ;
  assign n6102 = n6100 | n6101 ;
  assign n6103 = n4487 | n6102 ;
  assign n6104 = ( n5139 & n6102 ) | ( n5139 & n6103 ) | ( n6102 & n6103 ) ;
  assign n6105 = x26 & n6104 ;
  assign n6106 = x26 & ~n6105 ;
  assign n6107 = ( n6104 & ~n6105 ) | ( n6104 & n6106 ) | ( ~n6105 & n6106 ) ;
  assign n6108 = n6097 & n6107 ;
  assign n6109 = ~n5980 & n5982 ;
  assign n6110 = n5983 | n6109 ;
  assign n6111 = ~n2103 & n4479 ;
  assign n6112 = ~n1944 & n4481 ;
  assign n6113 = n6111 | n6112 ;
  assign n6114 = ~n1880 & n4484 ;
  assign n6115 = n6113 | n6114 ;
  assign n6116 = n4487 | n6115 ;
  assign n6117 = ( ~n5281 & n6115 ) | ( ~n5281 & n6116 ) | ( n6115 & n6116 ) ;
  assign n6118 = ~x26 & n6117 ;
  assign n6119 = x26 | n6118 ;
  assign n6120 = ( ~n6117 & n6118 ) | ( ~n6117 & n6119 ) | ( n6118 & n6119 ) ;
  assign n6121 = ~n6110 & n6120 ;
  assign n6122 = n5904 & ~n5976 ;
  assign n6123 = n5977 | n6122 ;
  assign n6124 = n2193 & n4479 ;
  assign n6125 = n2013 & n4481 ;
  assign n6126 = n6124 | n6125 ;
  assign n6127 = ~n2103 & n4484 ;
  assign n6128 = n6126 | n6127 ;
  assign n6129 = ( n4487 & ~n5836 ) | ( n4487 & n6128 ) | ( ~n5836 & n6128 ) ;
  assign n6130 = n6128 | n6129 ;
  assign n6131 = ~x26 & n6130 ;
  assign n6132 = x26 | n6131 ;
  assign n6133 = ( ~n6130 & n6131 ) | ( ~n6130 & n6132 ) | ( n6131 & n6132 ) ;
  assign n6134 = ~n6123 & n6133 ;
  assign n6135 = n6123 | n6134 ;
  assign n6136 = ( ~n6133 & n6134 ) | ( ~n6133 & n6135 ) | ( n6134 & n6135 ) ;
  assign n6137 = n2296 & n4479 ;
  assign n6138 = n2193 & n4481 ;
  assign n6139 = n6137 | n6138 ;
  assign n6140 = n2013 & n4484 ;
  assign n6141 = n6139 | n6140 ;
  assign n6142 = n4487 | n6141 ;
  assign n6143 = ( n5216 & n6141 ) | ( n5216 & n6142 ) | ( n6141 & n6142 ) ;
  assign n6144 = x26 & n6143 ;
  assign n6145 = x26 & ~n6144 ;
  assign n6146 = ( n6143 & ~n6144 ) | ( n6143 & n6145 ) | ( ~n6144 & n6145 ) ;
  assign n6147 = ~n2375 & n4479 ;
  assign n6148 = n2296 & n4481 ;
  assign n6149 = n6147 | n6148 ;
  assign n6150 = n2193 & n4484 ;
  assign n6151 = n6149 | n6150 ;
  assign n6152 = n4487 | n6151 ;
  assign n6153 = ( ~n5879 & n6151 ) | ( ~n5879 & n6152 ) | ( n6151 & n6152 ) ;
  assign n6154 = ~x26 & n6153 ;
  assign n6155 = x26 | n6154 ;
  assign n6156 = ( ~n6153 & n6154 ) | ( ~n6153 & n6155 ) | ( n6154 & n6155 ) ;
  assign n6157 = n5940 & ~n5973 ;
  assign n6158 = ( n5972 & ~n5973 ) | ( n5972 & n6157 ) | ( ~n5973 & n6157 ) ;
  assign n6159 = n6156 & n6158 ;
  assign n6160 = ~n2455 & n4479 ;
  assign n6161 = ~n2375 & n4481 ;
  assign n6162 = n6160 | n6161 ;
  assign n6163 = n2296 & n4484 ;
  assign n6164 = n6162 | n6163 ;
  assign n6165 = n4487 | n6164 ;
  assign n6166 = ( n5781 & n6164 ) | ( n5781 & n6165 ) | ( n6164 & n6165 ) ;
  assign n6167 = x26 & n6166 ;
  assign n6168 = x26 & ~n6167 ;
  assign n6169 = ( n6166 & ~n6167 ) | ( n6166 & n6168 ) | ( ~n6167 & n6168 ) ;
  assign n6170 = ( n5960 & n5971 ) | ( n5960 & ~n5972 ) | ( n5971 & ~n5972 ) ;
  assign n6171 = ( n5961 & ~n5972 ) | ( n5961 & n6170 ) | ( ~n5972 & n6170 ) ;
  assign n6172 = n6169 & n6171 ;
  assign n6173 = ~n2606 & n4479 ;
  assign n6174 = ~n2455 & n4481 ;
  assign n6175 = n6173 | n6174 ;
  assign n6176 = ~n2375 & n4484 ;
  assign n6177 = n6175 | n6176 ;
  assign n6178 = n4487 | n6177 ;
  assign n6179 = ( ~n5528 & n6177 ) | ( ~n5528 & n6178 ) | ( n6177 & n6178 ) ;
  assign n6180 = ~x26 & n6179 ;
  assign n6181 = x26 & ~n6179 ;
  assign n6182 = n6180 | n6181 ;
  assign n6183 = n5950 | n5959 ;
  assign n6184 = ~n5960 & n6183 ;
  assign n6185 = n6182 & n6184 ;
  assign n6186 = n6182 | n6184 ;
  assign n6187 = ~n6185 & n6186 ;
  assign n6188 = x29 & ~n5955 ;
  assign n6189 = n5957 | n6188 ;
  assign n6190 = n5958 | n6189 ;
  assign n6191 = ~n5959 & n6190 ;
  assign n6192 = ~n2455 & n4484 ;
  assign n6193 = ~n2606 & n4481 ;
  assign n6194 = n6192 | n6193 ;
  assign n6195 = n2569 & n4479 ;
  assign n6196 = n6194 | n6195 ;
  assign n6197 = n4487 | n6196 ;
  assign n6198 = ( ~n5732 & n6196 ) | ( ~n5732 & n6197 ) | ( n6196 & n6197 ) ;
  assign n6199 = ~x26 & n6198 ;
  assign n6200 = x26 | n6199 ;
  assign n6201 = ( ~n6198 & n6199 ) | ( ~n6198 & n6200 ) | ( n6199 & n6200 ) ;
  assign n6202 = n6191 & n6201 ;
  assign n6203 = ~n2764 & n4479 ;
  assign n6204 = ~n2672 & n4481 ;
  assign n6205 = n6203 | n6204 ;
  assign n6206 = n2569 & n4484 ;
  assign n6207 = n6205 | n6206 ;
  assign n6208 = ( n4487 & n5584 ) | ( n4487 & n6207 ) | ( n5584 & n6207 ) ;
  assign n6209 = ( x26 & ~n6207 ) | ( x26 & n6208 ) | ( ~n6207 & n6208 ) ;
  assign n6210 = ~n6208 & n6209 ;
  assign n6211 = n6207 | n6209 ;
  assign n6212 = ( ~x26 & n6210 ) | ( ~x26 & n6211 ) | ( n6210 & n6211 ) ;
  assign n6213 = ~n2764 & n4481 ;
  assign n6214 = ~n2672 & n4484 ;
  assign n6215 = n6213 | n6214 ;
  assign n6216 = n4487 | n6215 ;
  assign n6217 = ( n5932 & n6215 ) | ( n5932 & n6216 ) | ( n6215 & n6216 ) ;
  assign n6218 = ( n400 & ~n2763 ) | ( n400 & n4474 ) | ( ~n2763 & n4474 ) ;
  assign n6219 = x26 & ~n6218 ;
  assign n6220 = ~x26 & n6217 ;
  assign n6221 = ( ~n6217 & n6219 ) | ( ~n6217 & n6220 ) | ( n6219 & n6220 ) ;
  assign n6222 = n6212 & n6221 ;
  assign n6223 = n5956 & n6222 ;
  assign n6224 = ~n2606 & n4484 ;
  assign n6225 = ~n2672 & n4479 ;
  assign n6226 = n6224 | n6225 ;
  assign n6227 = n2569 & n4481 ;
  assign n6228 = n6226 | n6227 ;
  assign n6229 = n4487 | n6228 ;
  assign n6230 = ( n5716 & n6228 ) | ( n5716 & n6229 ) | ( n6228 & n6229 ) ;
  assign n6231 = x26 & n6230 ;
  assign n6232 = x26 & ~n6231 ;
  assign n6233 = ( n6230 & ~n6231 ) | ( n6230 & n6232 ) | ( ~n6231 & n6232 ) ;
  assign n6234 = n6222 & ~n6223 ;
  assign n6235 = ( n5956 & ~n6223 ) | ( n5956 & n6234 ) | ( ~n6223 & n6234 ) ;
  assign n6236 = n6233 & n6235 ;
  assign n6237 = n6223 | n6236 ;
  assign n6238 = n6191 | n6201 ;
  assign n6239 = ~n6202 & n6238 ;
  assign n6240 = n6237 & n6239 ;
  assign n6241 = n6202 | n6240 ;
  assign n6242 = n6187 & n6241 ;
  assign n6243 = n6185 | n6242 ;
  assign n6244 = n6169 & ~n6172 ;
  assign n6245 = ( n6171 & ~n6172 ) | ( n6171 & n6244 ) | ( ~n6172 & n6244 ) ;
  assign n6246 = n6243 & n6245 ;
  assign n6247 = n6172 | n6246 ;
  assign n6248 = n6156 | n6158 ;
  assign n6249 = ~n6159 & n6248 ;
  assign n6250 = n6247 & n6249 ;
  assign n6251 = n6159 | n6250 ;
  assign n6252 = n5920 & ~n5974 ;
  assign n6253 = n5975 | n6252 ;
  assign n6254 = n6146 & ~n6253 ;
  assign n6255 = n6253 | n6254 ;
  assign n6256 = ( ~n6146 & n6254 ) | ( ~n6146 & n6255 ) | ( n6254 & n6255 ) ;
  assign n6257 = n6251 | n6256 ;
  assign n6258 = n6251 & n6256 ;
  assign n6259 = n6257 & ~n6258 ;
  assign n6260 = ( n6146 & n6251 ) | ( n6146 & n6259 ) | ( n6251 & n6259 ) ;
  assign n6261 = ~n6136 & n6260 ;
  assign n6262 = n6134 | n6261 ;
  assign n6263 = n5887 | n5978 ;
  assign n6264 = ~n5979 & n6263 ;
  assign n6265 = n2013 & n4479 ;
  assign n6266 = ~n2103 & n4481 ;
  assign n6267 = n6265 | n6266 ;
  assign n6268 = ~n1944 & n4484 ;
  assign n6269 = n6267 | n6268 ;
  assign n6270 = n4487 | n6269 ;
  assign n6271 = ( n6041 & n6269 ) | ( n6041 & n6270 ) | ( n6269 & n6270 ) ;
  assign n6272 = x26 & n6271 ;
  assign n6273 = x26 & ~n6272 ;
  assign n6274 = ( n6271 & ~n6272 ) | ( n6271 & n6273 ) | ( ~n6272 & n6273 ) ;
  assign n6275 = ( n6262 & n6264 ) | ( n6262 & n6274 ) | ( n6264 & n6274 ) ;
  assign n6276 = n6110 | n6121 ;
  assign n6277 = ( ~n6120 & n6121 ) | ( ~n6120 & n6276 ) | ( n6121 & n6276 ) ;
  assign n6278 = n6275 & ~n6277 ;
  assign n6279 = n6121 | n6278 ;
  assign n6280 = n5849 | n5984 ;
  assign n6281 = ~n5985 & n6280 ;
  assign n6282 = n1803 & n4484 ;
  assign n6283 = ~n1944 & n4479 ;
  assign n6284 = n6282 | n6283 ;
  assign n6285 = ~n1880 & n4481 ;
  assign n6286 = n6284 | n6285 ;
  assign n6287 = n4487 | n6286 ;
  assign n6288 = ( n4905 & n6286 ) | ( n4905 & n6287 ) | ( n6286 & n6287 ) ;
  assign n6289 = x26 & n6288 ;
  assign n6290 = x26 & ~n6289 ;
  assign n6291 = ( n6288 & ~n6289 ) | ( n6288 & n6290 ) | ( ~n6289 & n6290 ) ;
  assign n6292 = ( n6279 & n6281 ) | ( n6279 & n6291 ) | ( n6281 & n6291 ) ;
  assign n6293 = n6097 & ~n6108 ;
  assign n6294 = ~n6097 & n6107 ;
  assign n6295 = n6293 | n6294 ;
  assign n6296 = n6292 & ~n6295 ;
  assign n6297 = ( n6108 & n6292 ) | ( n6108 & ~n6296 ) | ( n6292 & ~n6296 ) ;
  assign n6298 = n6094 & n6297 ;
  assign n6299 = n6094 | n6297 ;
  assign n6300 = ~n6298 & n6299 ;
  assign n6301 = n1625 & n4546 ;
  assign n6302 = n3030 & n4548 ;
  assign n6303 = n6301 | n6302 ;
  assign n6304 = ~n2939 & n4551 ;
  assign n6305 = n6303 | n6304 ;
  assign n6306 = n4554 | n6305 ;
  assign n6307 = ( ~n4215 & n6305 ) | ( ~n4215 & n6306 ) | ( n6305 & n6306 ) ;
  assign n6308 = ~x23 & n6307 ;
  assign n6309 = x23 | n6308 ;
  assign n6310 = ( ~n6307 & n6308 ) | ( ~n6307 & n6309 ) | ( n6308 & n6309 ) ;
  assign n6311 = n6300 & n6310 ;
  assign n6312 = n6300 | n6310 ;
  assign n6313 = ~n6311 & n6312 ;
  assign n6314 = ~n6292 & n6295 ;
  assign n6315 = n6296 | n6314 ;
  assign n6316 = ~n1733 & n4546 ;
  assign n6317 = n1625 & n4548 ;
  assign n6318 = n6316 | n6317 ;
  assign n6319 = n3030 & n4551 ;
  assign n6320 = n6318 | n6319 ;
  assign n6321 = n4554 | n6320 ;
  assign n6322 = ( ~n4578 & n6320 ) | ( ~n4578 & n6321 ) | ( n6320 & n6321 ) ;
  assign n6323 = ~x23 & n6322 ;
  assign n6324 = x23 | n6323 ;
  assign n6325 = ( ~n6322 & n6323 ) | ( ~n6322 & n6324 ) | ( n6323 & n6324 ) ;
  assign n6326 = n6315 & n6325 ;
  assign n6327 = n6315 | n6325 ;
  assign n6328 = ~n6326 & n6327 ;
  assign n6329 = ~n2873 & n4546 ;
  assign n6330 = ~n1733 & n4548 ;
  assign n6331 = n6329 | n6330 ;
  assign n6332 = n1625 & n4551 ;
  assign n6333 = n6331 | n6332 ;
  assign n6334 = n4554 | n6333 ;
  assign n6335 = ( n4260 & n6333 ) | ( n4260 & n6334 ) | ( n6333 & n6334 ) ;
  assign n6336 = x23 & n6335 ;
  assign n6337 = x23 & ~n6336 ;
  assign n6338 = ( n6335 & ~n6336 ) | ( n6335 & n6337 ) | ( ~n6336 & n6337 ) ;
  assign n6339 = ( n6279 & ~n6281 ) | ( n6279 & n6291 ) | ( ~n6281 & n6291 ) ;
  assign n6340 = ( ~n6279 & n6281 ) | ( ~n6279 & n6339 ) | ( n6281 & n6339 ) ;
  assign n6341 = ( ~n6291 & n6339 ) | ( ~n6291 & n6340 ) | ( n6339 & n6340 ) ;
  assign n6342 = n6338 & n6341 ;
  assign n6343 = n6275 & ~n6278 ;
  assign n6344 = n6277 | n6278 ;
  assign n6345 = ~n6343 & n6344 ;
  assign n6346 = n1803 & n4546 ;
  assign n6347 = ~n2873 & n4548 ;
  assign n6348 = n6346 | n6347 ;
  assign n6349 = ~n1733 & n4551 ;
  assign n6350 = n6348 | n6349 ;
  assign n6351 = n4554 | n6350 ;
  assign n6352 = ( ~n4985 & n6350 ) | ( ~n4985 & n6351 ) | ( n6350 & n6351 ) ;
  assign n6353 = ~x23 & n6352 ;
  assign n6354 = x23 | n6353 ;
  assign n6355 = ( ~n6352 & n6353 ) | ( ~n6352 & n6354 ) | ( n6353 & n6354 ) ;
  assign n6356 = ~n6345 & n6355 ;
  assign n6357 = ~n2873 & n4551 ;
  assign n6358 = n1803 & n4548 ;
  assign n6359 = n6357 | n6358 ;
  assign n6360 = ~n1880 & n4546 ;
  assign n6361 = n6359 | n6360 ;
  assign n6362 = n4554 | n6361 ;
  assign n6363 = ( n5139 & n6361 ) | ( n5139 & n6362 ) | ( n6361 & n6362 ) ;
  assign n6364 = x23 & n6363 ;
  assign n6365 = x23 & ~n6364 ;
  assign n6366 = ( n6363 & ~n6364 ) | ( n6363 & n6365 ) | ( ~n6364 & n6365 ) ;
  assign n6367 = ( n6262 & ~n6264 ) | ( n6262 & n6274 ) | ( ~n6264 & n6274 ) ;
  assign n6368 = ( ~n6262 & n6264 ) | ( ~n6262 & n6367 ) | ( n6264 & n6367 ) ;
  assign n6369 = ( ~n6274 & n6367 ) | ( ~n6274 & n6368 ) | ( n6367 & n6368 ) ;
  assign n6370 = n6366 & n6369 ;
  assign n6371 = n6260 & ~n6261 ;
  assign n6372 = n6136 | n6261 ;
  assign n6373 = ~n6371 & n6372 ;
  assign n6374 = n1803 & n4551 ;
  assign n6375 = ~n1944 & n4546 ;
  assign n6376 = n6374 | n6375 ;
  assign n6377 = ~n1880 & n4548 ;
  assign n6378 = n6376 | n6377 ;
  assign n6379 = n4554 | n6378 ;
  assign n6380 = ( n4905 & n6378 ) | ( n4905 & n6379 ) | ( n6378 & n6379 ) ;
  assign n6381 = x23 & n6380 ;
  assign n6382 = x23 & ~n6381 ;
  assign n6383 = ( n6380 & ~n6381 ) | ( n6380 & n6382 ) | ( ~n6381 & n6382 ) ;
  assign n6384 = ~n6373 & n6383 ;
  assign n6385 = ~n2103 & n4546 ;
  assign n6386 = ~n1944 & n4548 ;
  assign n6387 = n6385 | n6386 ;
  assign n6388 = ~n1880 & n4551 ;
  assign n6389 = n6387 | n6388 ;
  assign n6390 = n4554 | n6389 ;
  assign n6391 = ( ~n5281 & n6389 ) | ( ~n5281 & n6390 ) | ( n6389 & n6390 ) ;
  assign n6392 = ~x23 & n6391 ;
  assign n6393 = x23 | n6392 ;
  assign n6394 = ( ~n6391 & n6392 ) | ( ~n6391 & n6393 ) | ( n6392 & n6393 ) ;
  assign n6395 = ~n6259 & n6394 ;
  assign n6396 = n2013 & n4546 ;
  assign n6397 = ~n2103 & n4548 ;
  assign n6398 = n6396 | n6397 ;
  assign n6399 = ~n1944 & n4551 ;
  assign n6400 = n6398 | n6399 ;
  assign n6401 = n4554 | n6400 ;
  assign n6402 = ( n6041 & n6400 ) | ( n6041 & n6401 ) | ( n6400 & n6401 ) ;
  assign n6403 = x23 & n6402 ;
  assign n6404 = x23 & ~n6403 ;
  assign n6405 = ( n6402 & ~n6403 ) | ( n6402 & n6404 ) | ( ~n6403 & n6404 ) ;
  assign n6406 = n6247 & ~n6250 ;
  assign n6407 = ( n6249 & ~n6250 ) | ( n6249 & n6406 ) | ( ~n6250 & n6406 ) ;
  assign n6408 = n6405 & n6407 ;
  assign n6409 = n6407 & ~n6408 ;
  assign n6410 = n6405 & ~n6407 ;
  assign n6411 = n6243 | n6245 ;
  assign n6412 = ~n6246 & n6411 ;
  assign n6413 = n2193 & n4546 ;
  assign n6414 = n2013 & n4548 ;
  assign n6415 = n6413 | n6414 ;
  assign n6416 = ~n2103 & n4551 ;
  assign n6417 = n6415 | n6416 ;
  assign n6418 = n4554 | n6417 ;
  assign n6419 = ( ~n5836 & n6417 ) | ( ~n5836 & n6418 ) | ( n6417 & n6418 ) ;
  assign n6420 = ~x23 & n6419 ;
  assign n6421 = x23 | n6420 ;
  assign n6422 = ( ~n6419 & n6420 ) | ( ~n6419 & n6421 ) | ( n6420 & n6421 ) ;
  assign n6423 = n6412 & n6422 ;
  assign n6424 = n6412 | n6422 ;
  assign n6425 = ~n6423 & n6424 ;
  assign n6426 = n6187 | n6241 ;
  assign n6427 = ~n6242 & n6426 ;
  assign n6428 = n2296 & n4546 ;
  assign n6429 = n2193 & n4548 ;
  assign n6430 = n6428 | n6429 ;
  assign n6431 = n2013 & n4551 ;
  assign n6432 = n6430 | n6431 ;
  assign n6433 = n4554 | n6432 ;
  assign n6434 = ( n5216 & n6432 ) | ( n5216 & n6433 ) | ( n6432 & n6433 ) ;
  assign n6435 = x23 & n6434 ;
  assign n6436 = x23 & ~n6435 ;
  assign n6437 = ( n6434 & ~n6435 ) | ( n6434 & n6436 ) | ( ~n6435 & n6436 ) ;
  assign n6438 = n6237 | n6239 ;
  assign n6439 = ~n6240 & n6438 ;
  assign n6440 = ~n2375 & n4546 ;
  assign n6441 = n2296 & n4548 ;
  assign n6442 = n6440 | n6441 ;
  assign n6443 = n2193 & n4551 ;
  assign n6444 = n6442 | n6443 ;
  assign n6445 = n4554 | n6444 ;
  assign n6446 = ( ~n5879 & n6444 ) | ( ~n5879 & n6445 ) | ( n6444 & n6445 ) ;
  assign n6447 = ~x23 & n6446 ;
  assign n6448 = x23 | n6447 ;
  assign n6449 = ( ~n6446 & n6447 ) | ( ~n6446 & n6448 ) | ( n6447 & n6448 ) ;
  assign n6450 = n6439 & n6449 ;
  assign n6451 = n6233 | n6235 ;
  assign n6452 = ~n6236 & n6451 ;
  assign n6453 = ~n2455 & n4546 ;
  assign n6454 = ~n2375 & n4548 ;
  assign n6455 = n6453 | n6454 ;
  assign n6456 = n2296 & n4551 ;
  assign n6457 = n6455 | n6456 ;
  assign n6458 = n4554 | n6457 ;
  assign n6459 = ( n5781 & n6457 ) | ( n5781 & n6458 ) | ( n6457 & n6458 ) ;
  assign n6460 = x23 & n6459 ;
  assign n6461 = x23 & ~n6460 ;
  assign n6462 = ( n6459 & ~n6460 ) | ( n6459 & n6461 ) | ( ~n6460 & n6461 ) ;
  assign n6463 = n6452 & n6462 ;
  assign n6464 = ~n2606 & n4546 ;
  assign n6465 = ~n2455 & n4548 ;
  assign n6466 = n6464 | n6465 ;
  assign n6467 = ~n2375 & n4551 ;
  assign n6468 = n6466 | n6467 ;
  assign n6469 = n4554 | n6468 ;
  assign n6470 = ( ~n5528 & n6468 ) | ( ~n5528 & n6469 ) | ( n6468 & n6469 ) ;
  assign n6471 = ~x23 & n6470 ;
  assign n6472 = x23 & ~n6470 ;
  assign n6473 = n6471 | n6472 ;
  assign n6474 = n6212 | n6221 ;
  assign n6475 = ~n6222 & n6474 ;
  assign n6476 = n6473 & n6475 ;
  assign n6477 = n6473 | n6475 ;
  assign n6478 = ~n6476 & n6477 ;
  assign n6479 = x26 & ~n6217 ;
  assign n6480 = n6219 | n6479 ;
  assign n6481 = n6220 | n6480 ;
  assign n6482 = ~n6221 & n6481 ;
  assign n6483 = ~n2455 & n4551 ;
  assign n6484 = ~n2606 & n4548 ;
  assign n6485 = n6483 | n6484 ;
  assign n6486 = n2569 & n4546 ;
  assign n6487 = n6485 | n6486 ;
  assign n6488 = n4554 | n6487 ;
  assign n6489 = ( ~n5732 & n6487 ) | ( ~n5732 & n6488 ) | ( n6487 & n6488 ) ;
  assign n6490 = ~x23 & n6489 ;
  assign n6491 = x23 | n6490 ;
  assign n6492 = ( ~n6489 & n6490 ) | ( ~n6489 & n6491 ) | ( n6490 & n6491 ) ;
  assign n6493 = n6482 & n6492 ;
  assign n6494 = ~n2764 & n4546 ;
  assign n6495 = ~n2672 & n4548 ;
  assign n6496 = n6494 | n6495 ;
  assign n6497 = n2569 & n4551 ;
  assign n6498 = n6496 | n6497 ;
  assign n6499 = ( n4554 & n5584 ) | ( n4554 & n6498 ) | ( n5584 & n6498 ) ;
  assign n6500 = ( x23 & ~n6498 ) | ( x23 & n6499 ) | ( ~n6498 & n6499 ) ;
  assign n6501 = ~n6499 & n6500 ;
  assign n6502 = n6498 | n6500 ;
  assign n6503 = ( ~x23 & n6501 ) | ( ~x23 & n6502 ) | ( n6501 & n6502 ) ;
  assign n6504 = ~n2764 & n4548 ;
  assign n6505 = ~n2672 & n4551 ;
  assign n6506 = n6504 | n6505 ;
  assign n6507 = n4554 | n6506 ;
  assign n6508 = ( n5932 & n6506 ) | ( n5932 & n6507 ) | ( n6506 & n6507 ) ;
  assign n6509 = ~n2764 & n4541 ;
  assign n6510 = x23 & ~n6509 ;
  assign n6511 = ~x23 & n6508 ;
  assign n6512 = ( ~n6508 & n6510 ) | ( ~n6508 & n6511 ) | ( n6510 & n6511 ) ;
  assign n6513 = n6503 & n6512 ;
  assign n6514 = n6218 & n6513 ;
  assign n6515 = ~n2606 & n4551 ;
  assign n6516 = ~n2672 & n4546 ;
  assign n6517 = n6515 | n6516 ;
  assign n6518 = n2569 & n4548 ;
  assign n6519 = n6517 | n6518 ;
  assign n6520 = n4554 | n6519 ;
  assign n6521 = ( n5716 & n6519 ) | ( n5716 & n6520 ) | ( n6519 & n6520 ) ;
  assign n6522 = x23 & n6521 ;
  assign n6523 = x23 & ~n6522 ;
  assign n6524 = ( n6521 & ~n6522 ) | ( n6521 & n6523 ) | ( ~n6522 & n6523 ) ;
  assign n6525 = n6513 & ~n6514 ;
  assign n6526 = ( n6218 & ~n6514 ) | ( n6218 & n6525 ) | ( ~n6514 & n6525 ) ;
  assign n6527 = n6524 & n6526 ;
  assign n6528 = n6514 | n6527 ;
  assign n6529 = n6482 | n6492 ;
  assign n6530 = ~n6493 & n6529 ;
  assign n6531 = n6528 & n6530 ;
  assign n6532 = n6493 | n6531 ;
  assign n6533 = n6478 & n6532 ;
  assign n6534 = n6476 | n6533 ;
  assign n6535 = n6452 | n6462 ;
  assign n6536 = ~n6463 & n6535 ;
  assign n6537 = n6534 & n6536 ;
  assign n6538 = n6463 | n6537 ;
  assign n6539 = n6449 & ~n6450 ;
  assign n6540 = ( n6439 & ~n6450 ) | ( n6439 & n6539 ) | ( ~n6450 & n6539 ) ;
  assign n6541 = n6538 & n6540 ;
  assign n6542 = n6450 | n6541 ;
  assign n6543 = ( n6427 & n6437 ) | ( n6427 & n6542 ) | ( n6437 & n6542 ) ;
  assign n6544 = n6425 & n6543 ;
  assign n6545 = n6423 | n6544 ;
  assign n6546 = ( n6409 & n6410 ) | ( n6409 & n6545 ) | ( n6410 & n6545 ) ;
  assign n6547 = n6408 | n6546 ;
  assign n6548 = n6259 & ~n6394 ;
  assign n6549 = n6395 | n6548 ;
  assign n6550 = n6547 & ~n6549 ;
  assign n6551 = n6395 | n6550 ;
  assign n6552 = n6373 | n6384 ;
  assign n6553 = ( ~n6383 & n6384 ) | ( ~n6383 & n6552 ) | ( n6384 & n6552 ) ;
  assign n6554 = n6551 & ~n6553 ;
  assign n6555 = n6384 | n6554 ;
  assign n6556 = n6366 | n6369 ;
  assign n6557 = ~n6370 & n6556 ;
  assign n6558 = n6555 & n6557 ;
  assign n6559 = n6370 | n6558 ;
  assign n6560 = n6345 | n6356 ;
  assign n6561 = ( ~n6355 & n6356 ) | ( ~n6355 & n6560 ) | ( n6356 & n6560 ) ;
  assign n6562 = n6559 & ~n6561 ;
  assign n6563 = n6356 | n6562 ;
  assign n6564 = n6338 | n6341 ;
  assign n6565 = ~n6342 & n6564 ;
  assign n6566 = n6563 & n6565 ;
  assign n6567 = n6342 | n6566 ;
  assign n6568 = n6328 & n6567 ;
  assign n6569 = n6326 | n6568 ;
  assign n6570 = n6313 & n6569 ;
  assign n6571 = n6313 | n6569 ;
  assign n6572 = ~n6570 & n6571 ;
  assign n6573 = ~n1411 & n4778 ;
  assign n6574 = n4776 | n6573 ;
  assign n6575 = ( n1532 & n6573 ) | ( n1532 & n6574 ) | ( n6573 & n6574 ) ;
  assign n6576 = n3178 & n4781 ;
  assign n6577 = n6575 | n6576 ;
  assign n6578 = n4784 | n6577 ;
  assign n6579 = ( ~n3750 & n6577 ) | ( ~n3750 & n6578 ) | ( n6577 & n6578 ) ;
  assign n6580 = ~x20 & n6579 ;
  assign n6581 = x20 | n6580 ;
  assign n6582 = ( ~n6579 & n6580 ) | ( ~n6579 & n6581 ) | ( n6580 & n6581 ) ;
  assign n6583 = n6572 & n6582 ;
  assign n6584 = n6572 | n6582 ;
  assign n6585 = ~n6583 & n6584 ;
  assign n6586 = n6563 | n6565 ;
  assign n6587 = ~n6566 & n6586 ;
  assign n6588 = n1532 & n4781 ;
  assign n6589 = n3030 & n4776 ;
  assign n6590 = ~n2939 & n4778 ;
  assign n6591 = n6589 | n6590 ;
  assign n6592 = n6588 | n6591 ;
  assign n6593 = n4784 | n6592 ;
  assign n6594 = ( ~n4193 & n6592 ) | ( ~n4193 & n6593 ) | ( n6592 & n6593 ) ;
  assign n6595 = ~x20 & n6594 ;
  assign n6596 = x20 | n6595 ;
  assign n6597 = ( ~n6594 & n6595 ) | ( ~n6594 & n6596 ) | ( n6595 & n6596 ) ;
  assign n6598 = n6587 & n6597 ;
  assign n6599 = n6587 & ~n6598 ;
  assign n6600 = ~n6587 & n6597 ;
  assign n6601 = n6599 | n6600 ;
  assign n6602 = n6555 | n6557 ;
  assign n6603 = ~n6558 & n6602 ;
  assign n6604 = ~n1733 & n4776 ;
  assign n6605 = n1625 & n4778 ;
  assign n6606 = n6604 | n6605 ;
  assign n6607 = n3030 & n4781 ;
  assign n6608 = n6606 | n6607 ;
  assign n6609 = ( ~n4578 & n4784 ) | ( ~n4578 & n6608 ) | ( n4784 & n6608 ) ;
  assign n6610 = n6608 | n6609 ;
  assign n6611 = ~x20 & n6610 ;
  assign n6612 = x20 | n6611 ;
  assign n6613 = ( ~n6610 & n6611 ) | ( ~n6610 & n6612 ) | ( n6611 & n6612 ) ;
  assign n6614 = n6603 & n6613 ;
  assign n6615 = ~n6551 & n6553 ;
  assign n6616 = n6554 | n6615 ;
  assign n6617 = ~n2873 & n4776 ;
  assign n6618 = ~n1733 & n4778 ;
  assign n6619 = n6617 | n6618 ;
  assign n6620 = n1625 & n4781 ;
  assign n6621 = n6619 | n6620 ;
  assign n6622 = n4784 | n6621 ;
  assign n6623 = ( n4260 & n6621 ) | ( n4260 & n6622 ) | ( n6621 & n6622 ) ;
  assign n6624 = x20 & n6623 ;
  assign n6625 = x20 & ~n6624 ;
  assign n6626 = ( n6623 & ~n6624 ) | ( n6623 & n6625 ) | ( ~n6624 & n6625 ) ;
  assign n6627 = ~n6616 & n6626 ;
  assign n6628 = ~n6547 & n6549 ;
  assign n6629 = n6550 | n6628 ;
  assign n6630 = n1803 & n4776 ;
  assign n6631 = ~n2873 & n4778 ;
  assign n6632 = n6630 | n6631 ;
  assign n6633 = ~n1733 & n4781 ;
  assign n6634 = n6632 | n6633 ;
  assign n6635 = n4784 | n6634 ;
  assign n6636 = ( ~n4985 & n6634 ) | ( ~n4985 & n6635 ) | ( n6634 & n6635 ) ;
  assign n6637 = ~x20 & n6636 ;
  assign n6638 = x20 | n6637 ;
  assign n6639 = ( ~n6636 & n6637 ) | ( ~n6636 & n6638 ) | ( n6637 & n6638 ) ;
  assign n6640 = ~n6629 & n6639 ;
  assign n6641 = n6410 | n6545 ;
  assign n6642 = n6409 | n6641 ;
  assign n6643 = ~n6546 & n6642 ;
  assign n6644 = ~n2873 & n4781 ;
  assign n6645 = n1803 & n4778 ;
  assign n6646 = n6644 | n6645 ;
  assign n6647 = ~n1880 & n4776 ;
  assign n6648 = n6646 | n6647 ;
  assign n6649 = n4784 | n6648 ;
  assign n6650 = ( n5139 & n6648 ) | ( n5139 & n6649 ) | ( n6648 & n6649 ) ;
  assign n6651 = x20 & n6650 ;
  assign n6652 = x20 & ~n6651 ;
  assign n6653 = ( n6650 & ~n6651 ) | ( n6650 & n6652 ) | ( ~n6651 & n6652 ) ;
  assign n6654 = n6643 & n6653 ;
  assign n6655 = n6425 | n6543 ;
  assign n6656 = ~n6544 & n6655 ;
  assign n6657 = n1803 & n4781 ;
  assign n6658 = ~n1944 & n4776 ;
  assign n6659 = n6657 | n6658 ;
  assign n6660 = ~n1880 & n4778 ;
  assign n6661 = n6659 | n6660 ;
  assign n6662 = n4784 | n6661 ;
  assign n6663 = ( n4905 & n6661 ) | ( n4905 & n6662 ) | ( n6661 & n6662 ) ;
  assign n6664 = x20 & n6663 ;
  assign n6665 = x20 & ~n6664 ;
  assign n6666 = ( n6663 & ~n6664 ) | ( n6663 & n6665 ) | ( ~n6664 & n6665 ) ;
  assign n6667 = n6656 & n6666 ;
  assign n6668 = n6666 & ~n6667 ;
  assign n6669 = ( n6656 & ~n6667 ) | ( n6656 & n6668 ) | ( ~n6667 & n6668 ) ;
  assign n6670 = ~n2103 & n4776 ;
  assign n6671 = ~n1944 & n4778 ;
  assign n6672 = n6670 | n6671 ;
  assign n6673 = ~n1880 & n4781 ;
  assign n6674 = n6672 | n6673 ;
  assign n6675 = n4784 | n6674 ;
  assign n6676 = ( ~n5281 & n6674 ) | ( ~n5281 & n6675 ) | ( n6674 & n6675 ) ;
  assign n6677 = ~x20 & n6676 ;
  assign n6678 = x20 | n6677 ;
  assign n6679 = ( ~n6676 & n6677 ) | ( ~n6676 & n6678 ) | ( n6677 & n6678 ) ;
  assign n6680 = ( n6427 & n6542 ) | ( n6427 & ~n6543 ) | ( n6542 & ~n6543 ) ;
  assign n6681 = ( n6437 & ~n6543 ) | ( n6437 & n6680 ) | ( ~n6543 & n6680 ) ;
  assign n6682 = n6679 & n6681 ;
  assign n6683 = n6679 | n6681 ;
  assign n6684 = ~n6682 & n6683 ;
  assign n6685 = n6538 | n6540 ;
  assign n6686 = ~n6541 & n6685 ;
  assign n6687 = n2013 & n4776 ;
  assign n6688 = ~n2103 & n4778 ;
  assign n6689 = n6687 | n6688 ;
  assign n6690 = ~n1944 & n4781 ;
  assign n6691 = n6689 | n6690 ;
  assign n6692 = n4784 | n6691 ;
  assign n6693 = ( n6041 & n6691 ) | ( n6041 & n6692 ) | ( n6691 & n6692 ) ;
  assign n6694 = x20 & n6693 ;
  assign n6695 = x20 & ~n6694 ;
  assign n6696 = ( n6693 & ~n6694 ) | ( n6693 & n6695 ) | ( ~n6694 & n6695 ) ;
  assign n6697 = n6686 & n6696 ;
  assign n6698 = n6534 | n6536 ;
  assign n6699 = ~n6537 & n6698 ;
  assign n6700 = n2193 & n4776 ;
  assign n6701 = n2013 & n4778 ;
  assign n6702 = n6700 | n6701 ;
  assign n6703 = ~n2103 & n4781 ;
  assign n6704 = n6702 | n6703 ;
  assign n6705 = n4784 | n6704 ;
  assign n6706 = ( ~n5836 & n6704 ) | ( ~n5836 & n6705 ) | ( n6704 & n6705 ) ;
  assign n6707 = ~x20 & n6706 ;
  assign n6708 = x20 | n6707 ;
  assign n6709 = ( ~n6706 & n6707 ) | ( ~n6706 & n6708 ) | ( n6707 & n6708 ) ;
  assign n6710 = n6699 & n6709 ;
  assign n6711 = n6699 & ~n6710 ;
  assign n6712 = ~n6699 & n6709 ;
  assign n6713 = n6711 | n6712 ;
  assign n6714 = n6478 | n6532 ;
  assign n6715 = ~n6533 & n6714 ;
  assign n6716 = n2296 & n4776 ;
  assign n6717 = n2193 & n4778 ;
  assign n6718 = n6716 | n6717 ;
  assign n6719 = n2013 & n4781 ;
  assign n6720 = n6718 | n6719 ;
  assign n6721 = n4784 | n6720 ;
  assign n6722 = ( n5216 & n6720 ) | ( n5216 & n6721 ) | ( n6720 & n6721 ) ;
  assign n6723 = x20 & n6722 ;
  assign n6724 = x20 & ~n6723 ;
  assign n6725 = ( n6722 & ~n6723 ) | ( n6722 & n6724 ) | ( ~n6723 & n6724 ) ;
  assign n6726 = n6528 | n6530 ;
  assign n6727 = ~n6531 & n6726 ;
  assign n6728 = ~n2375 & n4776 ;
  assign n6729 = n2296 & n4778 ;
  assign n6730 = n6728 | n6729 ;
  assign n6731 = n2193 & n4781 ;
  assign n6732 = n6730 | n6731 ;
  assign n6733 = n4784 | n6732 ;
  assign n6734 = ( ~n5879 & n6732 ) | ( ~n5879 & n6733 ) | ( n6732 & n6733 ) ;
  assign n6735 = ~x20 & n6734 ;
  assign n6736 = x20 | n6735 ;
  assign n6737 = ( ~n6734 & n6735 ) | ( ~n6734 & n6736 ) | ( n6735 & n6736 ) ;
  assign n6738 = n6727 & n6737 ;
  assign n6739 = n6524 | n6526 ;
  assign n6740 = ~n6527 & n6739 ;
  assign n6741 = ~n2455 & n4776 ;
  assign n6742 = ~n2375 & n4778 ;
  assign n6743 = n6741 | n6742 ;
  assign n6744 = n2296 & n4781 ;
  assign n6745 = n6743 | n6744 ;
  assign n6746 = n4784 | n6745 ;
  assign n6747 = ( n5781 & n6745 ) | ( n5781 & n6746 ) | ( n6745 & n6746 ) ;
  assign n6748 = x20 & n6747 ;
  assign n6749 = x20 & ~n6748 ;
  assign n6750 = ( n6747 & ~n6748 ) | ( n6747 & n6749 ) | ( ~n6748 & n6749 ) ;
  assign n6751 = n6740 & n6750 ;
  assign n6752 = ~n2606 & n4776 ;
  assign n6753 = ~n2455 & n4778 ;
  assign n6754 = n6752 | n6753 ;
  assign n6755 = ~n2375 & n4781 ;
  assign n6756 = n6754 | n6755 ;
  assign n6757 = n4784 | n6756 ;
  assign n6758 = ( ~n5528 & n6756 ) | ( ~n5528 & n6757 ) | ( n6756 & n6757 ) ;
  assign n6759 = ~x20 & n6758 ;
  assign n6760 = x20 & ~n6758 ;
  assign n6761 = n6759 | n6760 ;
  assign n6762 = n6503 | n6512 ;
  assign n6763 = ~n6513 & n6762 ;
  assign n6764 = n6761 & n6763 ;
  assign n6765 = n6761 | n6763 ;
  assign n6766 = ~n6764 & n6765 ;
  assign n6767 = x23 & ~n6508 ;
  assign n6768 = n6510 | n6767 ;
  assign n6769 = n6511 | n6768 ;
  assign n6770 = ~n6512 & n6769 ;
  assign n6771 = ~n2455 & n4781 ;
  assign n6772 = ~n2606 & n4778 ;
  assign n6773 = n6771 | n6772 ;
  assign n6774 = n2569 & n4776 ;
  assign n6775 = n6773 | n6774 ;
  assign n6776 = n4784 | n6775 ;
  assign n6777 = ( ~n5732 & n6775 ) | ( ~n5732 & n6776 ) | ( n6775 & n6776 ) ;
  assign n6778 = ~x20 & n6777 ;
  assign n6779 = x20 | n6778 ;
  assign n6780 = ( ~n6777 & n6778 ) | ( ~n6777 & n6779 ) | ( n6778 & n6779 ) ;
  assign n6781 = n6770 & n6780 ;
  assign n6782 = ~n2764 & n4776 ;
  assign n6783 = ~n2672 & n4778 ;
  assign n6784 = n6782 | n6783 ;
  assign n6785 = n2569 & n4781 ;
  assign n6786 = n6784 | n6785 ;
  assign n6787 = ( n4784 & n5584 ) | ( n4784 & n6786 ) | ( n5584 & n6786 ) ;
  assign n6788 = ( x20 & ~n6786 ) | ( x20 & n6787 ) | ( ~n6786 & n6787 ) ;
  assign n6789 = ~n6787 & n6788 ;
  assign n6790 = n6786 | n6788 ;
  assign n6791 = ( ~x20 & n6789 ) | ( ~x20 & n6790 ) | ( n6789 & n6790 ) ;
  assign n6792 = ~n2764 & n4778 ;
  assign n6793 = ~n2672 & n4781 ;
  assign n6794 = n6792 | n6793 ;
  assign n6795 = n4784 | n6794 ;
  assign n6796 = ( n5932 & n6794 ) | ( n5932 & n6795 ) | ( n6794 & n6795 ) ;
  assign n6797 = ~n2764 & n4774 ;
  assign n6798 = x20 & ~n6797 ;
  assign n6799 = ~x20 & n6796 ;
  assign n6800 = ( ~n6796 & n6798 ) | ( ~n6796 & n6799 ) | ( n6798 & n6799 ) ;
  assign n6801 = n6791 & n6800 ;
  assign n6802 = n6509 & n6801 ;
  assign n6803 = n6801 & ~n6802 ;
  assign n6804 = n6509 & ~n6801 ;
  assign n6805 = n6803 | n6804 ;
  assign n6806 = ~n2606 & n4781 ;
  assign n6807 = ~n2672 & n4776 ;
  assign n6808 = n6806 | n6807 ;
  assign n6809 = n2569 & n4778 ;
  assign n6810 = n6808 | n6809 ;
  assign n6811 = n4784 | n6810 ;
  assign n6812 = ( n5716 & n6810 ) | ( n5716 & n6811 ) | ( n6810 & n6811 ) ;
  assign n6813 = x20 & n6812 ;
  assign n6814 = x20 & ~n6813 ;
  assign n6815 = ( n6812 & ~n6813 ) | ( n6812 & n6814 ) | ( ~n6813 & n6814 ) ;
  assign n6816 = n6805 & n6815 ;
  assign n6817 = n6802 | n6816 ;
  assign n6818 = n6770 | n6780 ;
  assign n6819 = ~n6781 & n6818 ;
  assign n6820 = n6817 & n6819 ;
  assign n6821 = n6781 | n6820 ;
  assign n6822 = n6766 & n6821 ;
  assign n6823 = n6764 | n6822 ;
  assign n6824 = n6740 | n6750 ;
  assign n6825 = ~n6751 & n6824 ;
  assign n6826 = n6823 & n6825 ;
  assign n6827 = n6751 | n6826 ;
  assign n6828 = n6737 & ~n6738 ;
  assign n6829 = ( n6727 & ~n6738 ) | ( n6727 & n6828 ) | ( ~n6738 & n6828 ) ;
  assign n6830 = n6827 & n6829 ;
  assign n6831 = n6738 | n6830 ;
  assign n6832 = ( n6715 & n6725 ) | ( n6715 & n6831 ) | ( n6725 & n6831 ) ;
  assign n6833 = n6713 & n6832 ;
  assign n6834 = n6710 | n6833 ;
  assign n6835 = n6686 | n6696 ;
  assign n6836 = ~n6697 & n6835 ;
  assign n6837 = n6834 & n6836 ;
  assign n6838 = n6697 | n6837 ;
  assign n6839 = n6684 & n6838 ;
  assign n6840 = n6682 | n6839 ;
  assign n6841 = n6669 & n6840 ;
  assign n6842 = n6667 | n6841 ;
  assign n6843 = n6643 & ~n6654 ;
  assign n6844 = ~n6643 & n6653 ;
  assign n6845 = n6843 | n6844 ;
  assign n6846 = n6842 & n6845 ;
  assign n6847 = n6654 | n6846 ;
  assign n6848 = n6629 | n6640 ;
  assign n6849 = ( ~n6639 & n6640 ) | ( ~n6639 & n6848 ) | ( n6640 & n6848 ) ;
  assign n6850 = n6847 & ~n6849 ;
  assign n6851 = n6640 | n6850 ;
  assign n6852 = n6616 | n6627 ;
  assign n6853 = ( ~n6626 & n6627 ) | ( ~n6626 & n6852 ) | ( n6627 & n6852 ) ;
  assign n6854 = n6851 & ~n6853 ;
  assign n6855 = n6627 | n6854 ;
  assign n6856 = n6603 & ~n6614 ;
  assign n6857 = ~n6603 & n6613 ;
  assign n6858 = n6856 | n6857 ;
  assign n6859 = n6855 & n6858 ;
  assign n6860 = n6614 | n6859 ;
  assign n6861 = n1625 & n4776 ;
  assign n6862 = n3030 & n4778 ;
  assign n6863 = n6861 | n6862 ;
  assign n6864 = ~n2939 & n4781 ;
  assign n6865 = n6863 | n6864 ;
  assign n6866 = n4784 | n6865 ;
  assign n6867 = ( ~n4215 & n6865 ) | ( ~n4215 & n6866 ) | ( n6865 & n6866 ) ;
  assign n6868 = ~x20 & n6867 ;
  assign n6869 = x20 | n6868 ;
  assign n6870 = ( ~n6867 & n6868 ) | ( ~n6867 & n6869 ) | ( n6868 & n6869 ) ;
  assign n6871 = ~n6559 & n6561 ;
  assign n6872 = n6562 | n6871 ;
  assign n6873 = ( n6860 & n6870 ) | ( n6860 & ~n6872 ) | ( n6870 & ~n6872 ) ;
  assign n6874 = n6601 & n6873 ;
  assign n6875 = n6598 | n6874 ;
  assign n6876 = n6328 | n6567 ;
  assign n6877 = ~n6568 & n6876 ;
  assign n6878 = n1532 & n4778 ;
  assign n6879 = ~n1411 & n4781 ;
  assign n6880 = ~n2939 & n4776 ;
  assign n6881 = n6879 | n6880 ;
  assign n6882 = n6878 | n6881 ;
  assign n6883 = n4784 | n6882 ;
  assign n6884 = ( ~n3930 & n6882 ) | ( ~n3930 & n6883 ) | ( n6882 & n6883 ) ;
  assign n6885 = ~x20 & n6884 ;
  assign n6886 = x20 | n6885 ;
  assign n6887 = ( ~n6884 & n6885 ) | ( ~n6884 & n6886 ) | ( n6885 & n6886 ) ;
  assign n6888 = ( n6875 & n6877 ) | ( n6875 & n6887 ) | ( n6877 & n6887 ) ;
  assign n6889 = n6585 & n6888 ;
  assign n6890 = n6585 | n6888 ;
  assign n6891 = ~n6889 & n6890 ;
  assign n6892 = n3104 & n5069 ;
  assign n6893 = n1327 & n5070 ;
  assign n6894 = n6892 | n6893 ;
  assign n6895 = ~n1151 & n5083 ;
  assign n6896 = n6894 | n6895 ;
  assign n6897 = n5074 | n6896 ;
  assign n6898 = ( ~n4034 & n6896 ) | ( ~n4034 & n6897 ) | ( n6896 & n6897 ) ;
  assign n6899 = ~x17 & n6898 ;
  assign n6900 = x17 | n6899 ;
  assign n6901 = ( ~n6898 & n6899 ) | ( ~n6898 & n6900 ) | ( n6899 & n6900 ) ;
  assign n6902 = n6891 & n6901 ;
  assign n6903 = n6891 | n6901 ;
  assign n6904 = ~n6902 & n6903 ;
  assign n6905 = n3178 & n5069 ;
  assign n6906 = n3104 & n5070 ;
  assign n6907 = n6905 | n6906 ;
  assign n6908 = n1327 & n5083 ;
  assign n6909 = n6907 | n6908 ;
  assign n6910 = n5074 | n6909 ;
  assign n6911 = ( n4501 & n6909 ) | ( n4501 & n6910 ) | ( n6909 & n6910 ) ;
  assign n6912 = x17 & n6911 ;
  assign n6913 = x17 & ~n6912 ;
  assign n6914 = ( n6911 & ~n6912 ) | ( n6911 & n6913 ) | ( ~n6912 & n6913 ) ;
  assign n6915 = ( n6875 & ~n6877 ) | ( n6875 & n6887 ) | ( ~n6877 & n6887 ) ;
  assign n6916 = ( ~n6875 & n6877 ) | ( ~n6875 & n6915 ) | ( n6877 & n6915 ) ;
  assign n6917 = ( ~n6887 & n6915 ) | ( ~n6887 & n6916 ) | ( n6915 & n6916 ) ;
  assign n6918 = n6914 & n6917 ;
  assign n6919 = n6873 & ~n6874 ;
  assign n6920 = n6601 & ~n6874 ;
  assign n6921 = n6919 | n6920 ;
  assign n6922 = ~n1411 & n5069 ;
  assign n6923 = n3178 & n5070 ;
  assign n6924 = n6922 | n6923 ;
  assign n6925 = n3104 & n5083 ;
  assign n6926 = n6924 | n6925 ;
  assign n6927 = n5074 | n6926 ;
  assign n6928 = ( n4449 & n6926 ) | ( n4449 & n6927 ) | ( n6926 & n6927 ) ;
  assign n6929 = x17 & n6928 ;
  assign n6930 = x17 & ~n6929 ;
  assign n6931 = ( n6928 & ~n6929 ) | ( n6928 & n6930 ) | ( ~n6929 & n6930 ) ;
  assign n6932 = n6921 & n6931 ;
  assign n6933 = n6921 & ~n6932 ;
  assign n6934 = ~n6921 & n6931 ;
  assign n6935 = n6933 | n6934 ;
  assign n6936 = ( ~n6860 & n6872 ) | ( ~n6860 & n6873 ) | ( n6872 & n6873 ) ;
  assign n6937 = ( ~n6870 & n6873 ) | ( ~n6870 & n6936 ) | ( n6873 & n6936 ) ;
  assign n6938 = ~n1411 & n5070 ;
  assign n6939 = n5069 | n6938 ;
  assign n6940 = ( n1532 & n6938 ) | ( n1532 & n6939 ) | ( n6938 & n6939 ) ;
  assign n6941 = n3178 & n5083 ;
  assign n6942 = n6940 | n6941 ;
  assign n6943 = n5074 | n6942 ;
  assign n6944 = ( ~n3750 & n6942 ) | ( ~n3750 & n6943 ) | ( n6942 & n6943 ) ;
  assign n6945 = ~x17 & n6944 ;
  assign n6946 = x17 | n6945 ;
  assign n6947 = ( ~n6944 & n6945 ) | ( ~n6944 & n6946 ) | ( n6945 & n6946 ) ;
  assign n6948 = ~n6937 & n6947 ;
  assign n6949 = n6937 & ~n6947 ;
  assign n6950 = n6948 | n6949 ;
  assign n6951 = n6855 & ~n6859 ;
  assign n6952 = n6858 & ~n6859 ;
  assign n6953 = n6951 | n6952 ;
  assign n6954 = n1532 & n5070 ;
  assign n6955 = ~n1411 & n5083 ;
  assign n6956 = ~n2939 & n5069 ;
  assign n6957 = n6955 | n6956 ;
  assign n6958 = n6954 | n6957 ;
  assign n6959 = n5074 | n6958 ;
  assign n6960 = ( ~n3930 & n6958 ) | ( ~n3930 & n6959 ) | ( n6958 & n6959 ) ;
  assign n6961 = ~x17 & n6960 ;
  assign n6962 = x17 | n6961 ;
  assign n6963 = ( ~n6960 & n6961 ) | ( ~n6960 & n6962 ) | ( n6961 & n6962 ) ;
  assign n6964 = n6953 & n6963 ;
  assign n6965 = n6953 & ~n6964 ;
  assign n6966 = ~n6953 & n6963 ;
  assign n6967 = n6965 | n6966 ;
  assign n6968 = n6851 & ~n6854 ;
  assign n6969 = n6853 | n6854 ;
  assign n6970 = ~n6968 & n6969 ;
  assign n6971 = n1532 & n5083 ;
  assign n6972 = n3030 & n5069 ;
  assign n6973 = ~n2939 & n5070 ;
  assign n6974 = n6972 | n6973 ;
  assign n6975 = n6971 | n6974 ;
  assign n6976 = n5074 | n6975 ;
  assign n6977 = ( ~n4193 & n6975 ) | ( ~n4193 & n6976 ) | ( n6975 & n6976 ) ;
  assign n6978 = ~x17 & n6977 ;
  assign n6979 = x17 | n6978 ;
  assign n6980 = ( ~n6977 & n6978 ) | ( ~n6977 & n6979 ) | ( n6978 & n6979 ) ;
  assign n6981 = ~n6970 & n6980 ;
  assign n6982 = n6847 & ~n6850 ;
  assign n6983 = n6849 | n6850 ;
  assign n6984 = ~n6982 & n6983 ;
  assign n6985 = n1625 & n5069 ;
  assign n6986 = n3030 & n5070 ;
  assign n6987 = n6985 | n6986 ;
  assign n6988 = ~n2939 & n5083 ;
  assign n6989 = n6987 | n6988 ;
  assign n6990 = n5074 | n6989 ;
  assign n6991 = ( ~n4215 & n6989 ) | ( ~n4215 & n6990 ) | ( n6989 & n6990 ) ;
  assign n6992 = ~x17 & n6991 ;
  assign n6993 = x17 | n6992 ;
  assign n6994 = ( ~n6991 & n6992 ) | ( ~n6991 & n6993 ) | ( n6992 & n6993 ) ;
  assign n6995 = ~n6984 & n6994 ;
  assign n6996 = n6842 & ~n6846 ;
  assign n6997 = n6845 & ~n6846 ;
  assign n6998 = n6996 | n6997 ;
  assign n6999 = ~n1733 & n5069 ;
  assign n7000 = n1625 & n5070 ;
  assign n7001 = n6999 | n7000 ;
  assign n7002 = n3030 & n5083 ;
  assign n7003 = n7001 | n7002 ;
  assign n7004 = n5074 | n7003 ;
  assign n7005 = ( ~n4578 & n7003 ) | ( ~n4578 & n7004 ) | ( n7003 & n7004 ) ;
  assign n7006 = ~x17 & n7005 ;
  assign n7007 = x17 | n7006 ;
  assign n7008 = ( ~n7005 & n7006 ) | ( ~n7005 & n7007 ) | ( n7006 & n7007 ) ;
  assign n7009 = n6998 & n7008 ;
  assign n7010 = n6998 & ~n7009 ;
  assign n7011 = ~n6998 & n7008 ;
  assign n7012 = n7010 | n7011 ;
  assign n7013 = n6669 | n6840 ;
  assign n7014 = ~n6841 & n7013 ;
  assign n7015 = ~n2873 & n5069 ;
  assign n7016 = ~n1733 & n5070 ;
  assign n7017 = n7015 | n7016 ;
  assign n7018 = n1625 & n5083 ;
  assign n7019 = n7017 | n7018 ;
  assign n7020 = n5074 | n7019 ;
  assign n7021 = ( n4260 & n7019 ) | ( n4260 & n7020 ) | ( n7019 & n7020 ) ;
  assign n7022 = x17 & n7021 ;
  assign n7023 = x17 & ~n7022 ;
  assign n7024 = ( n7021 & ~n7022 ) | ( n7021 & n7023 ) | ( ~n7022 & n7023 ) ;
  assign n7025 = n7014 & n7024 ;
  assign n7026 = n6684 | n6838 ;
  assign n7027 = ~n6839 & n7026 ;
  assign n7028 = n1803 & n5069 ;
  assign n7029 = ~n2873 & n5070 ;
  assign n7030 = n7028 | n7029 ;
  assign n7031 = ~n1733 & n5083 ;
  assign n7032 = n7030 | n7031 ;
  assign n7033 = n5074 | n7032 ;
  assign n7034 = ( ~n4985 & n7032 ) | ( ~n4985 & n7033 ) | ( n7032 & n7033 ) ;
  assign n7035 = ~x17 & n7034 ;
  assign n7036 = x17 | n7035 ;
  assign n7037 = ( ~n7034 & n7035 ) | ( ~n7034 & n7036 ) | ( n7035 & n7036 ) ;
  assign n7038 = n7027 & n7037 ;
  assign n7039 = n6834 | n6836 ;
  assign n7040 = ~n6837 & n7039 ;
  assign n7041 = ~n2873 & n5083 ;
  assign n7042 = n1803 & n5070 ;
  assign n7043 = n7041 | n7042 ;
  assign n7044 = ~n1880 & n5069 ;
  assign n7045 = n7043 | n7044 ;
  assign n7046 = n5074 | n7045 ;
  assign n7047 = ( n5139 & n7045 ) | ( n5139 & n7046 ) | ( n7045 & n7046 ) ;
  assign n7048 = x17 & n7047 ;
  assign n7049 = x17 & ~n7048 ;
  assign n7050 = ( n7047 & ~n7048 ) | ( n7047 & n7049 ) | ( ~n7048 & n7049 ) ;
  assign n7051 = n7040 & n7050 ;
  assign n7052 = n7050 & ~n7051 ;
  assign n7053 = ( n7040 & ~n7051 ) | ( n7040 & n7052 ) | ( ~n7051 & n7052 ) ;
  assign n7054 = n1803 & n5083 ;
  assign n7055 = ~n1944 & n5069 ;
  assign n7056 = n7054 | n7055 ;
  assign n7057 = ~n1880 & n5070 ;
  assign n7058 = n7056 | n7057 ;
  assign n7059 = n5074 | n7058 ;
  assign n7060 = ( n4905 & n7058 ) | ( n4905 & n7059 ) | ( n7058 & n7059 ) ;
  assign n7061 = x17 & n7060 ;
  assign n7062 = x17 & ~n7061 ;
  assign n7063 = ( n7060 & ~n7061 ) | ( n7060 & n7062 ) | ( ~n7061 & n7062 ) ;
  assign n7064 = n6713 & ~n6833 ;
  assign n7065 = ( n6832 & ~n6833 ) | ( n6832 & n7064 ) | ( ~n6833 & n7064 ) ;
  assign n7066 = n7063 & n7065 ;
  assign n7067 = n7065 & ~n7066 ;
  assign n7068 = n7063 & ~n7065 ;
  assign n7069 = n7067 | n7068 ;
  assign n7070 = ~n2103 & n5069 ;
  assign n7071 = ~n1944 & n5070 ;
  assign n7072 = n7070 | n7071 ;
  assign n7073 = ~n1880 & n5083 ;
  assign n7074 = n7072 | n7073 ;
  assign n7075 = n5074 | n7074 ;
  assign n7076 = ( ~n5281 & n7074 ) | ( ~n5281 & n7075 ) | ( n7074 & n7075 ) ;
  assign n7077 = ~x17 & n7076 ;
  assign n7078 = x17 | n7077 ;
  assign n7079 = ( ~n7076 & n7077 ) | ( ~n7076 & n7078 ) | ( n7077 & n7078 ) ;
  assign n7080 = ( n6715 & n6831 ) | ( n6715 & ~n6832 ) | ( n6831 & ~n6832 ) ;
  assign n7081 = ( n6725 & ~n6832 ) | ( n6725 & n7080 ) | ( ~n6832 & n7080 ) ;
  assign n7082 = n7079 & n7081 ;
  assign n7083 = n7079 | n7081 ;
  assign n7084 = ~n7082 & n7083 ;
  assign n7085 = n6827 | n6829 ;
  assign n7086 = ~n6830 & n7085 ;
  assign n7087 = n2013 & n5069 ;
  assign n7088 = ~n2103 & n5070 ;
  assign n7089 = n7087 | n7088 ;
  assign n7090 = ~n1944 & n5083 ;
  assign n7091 = n7089 | n7090 ;
  assign n7092 = n5074 | n7091 ;
  assign n7093 = ( n6041 & n7091 ) | ( n6041 & n7092 ) | ( n7091 & n7092 ) ;
  assign n7094 = x17 & n7093 ;
  assign n7095 = x17 & ~n7094 ;
  assign n7096 = ( n7093 & ~n7094 ) | ( n7093 & n7095 ) | ( ~n7094 & n7095 ) ;
  assign n7097 = n7086 & n7096 ;
  assign n7098 = n6823 | n6825 ;
  assign n7099 = ~n6826 & n7098 ;
  assign n7100 = n2193 & n5069 ;
  assign n7101 = n2013 & n5070 ;
  assign n7102 = n7100 | n7101 ;
  assign n7103 = ~n2103 & n5083 ;
  assign n7104 = n7102 | n7103 ;
  assign n7105 = n5074 | n7104 ;
  assign n7106 = ( ~n5836 & n7104 ) | ( ~n5836 & n7105 ) | ( n7104 & n7105 ) ;
  assign n7107 = ~x17 & n7106 ;
  assign n7108 = x17 | n7107 ;
  assign n7109 = ( ~n7106 & n7107 ) | ( ~n7106 & n7108 ) | ( n7107 & n7108 ) ;
  assign n7110 = n7099 & n7109 ;
  assign n7111 = n7099 & ~n7110 ;
  assign n7112 = ~n7099 & n7109 ;
  assign n7113 = n7111 | n7112 ;
  assign n7114 = n6766 | n6821 ;
  assign n7115 = ~n6822 & n7114 ;
  assign n7116 = n2296 & n5069 ;
  assign n7117 = n2193 & n5070 ;
  assign n7118 = n7116 | n7117 ;
  assign n7119 = n2013 & n5083 ;
  assign n7120 = n7118 | n7119 ;
  assign n7121 = n5074 | n7120 ;
  assign n7122 = ( n5216 & n7120 ) | ( n5216 & n7121 ) | ( n7120 & n7121 ) ;
  assign n7123 = x17 & n7122 ;
  assign n7124 = x17 & ~n7123 ;
  assign n7125 = ( n7122 & ~n7123 ) | ( n7122 & n7124 ) | ( ~n7123 & n7124 ) ;
  assign n7126 = n6817 | n6819 ;
  assign n7127 = ~n6820 & n7126 ;
  assign n7128 = ~n2375 & n5069 ;
  assign n7129 = n2296 & n5070 ;
  assign n7130 = n7128 | n7129 ;
  assign n7131 = n2193 & n5083 ;
  assign n7132 = n7130 | n7131 ;
  assign n7133 = n5074 | n7132 ;
  assign n7134 = ( ~n5879 & n7132 ) | ( ~n5879 & n7133 ) | ( n7132 & n7133 ) ;
  assign n7135 = ~x17 & n7134 ;
  assign n7136 = x17 | n7135 ;
  assign n7137 = ( ~n7134 & n7135 ) | ( ~n7134 & n7136 ) | ( n7135 & n7136 ) ;
  assign n7138 = n7127 & n7137 ;
  assign n7139 = n6805 | n6815 ;
  assign n7140 = ~n6816 & n7139 ;
  assign n7141 = ~n2455 & n5069 ;
  assign n7142 = ~n2375 & n5070 ;
  assign n7143 = n7141 | n7142 ;
  assign n7144 = n2296 & n5083 ;
  assign n7145 = n7143 | n7144 ;
  assign n7146 = n5074 | n7145 ;
  assign n7147 = ( n5781 & n7145 ) | ( n5781 & n7146 ) | ( n7145 & n7146 ) ;
  assign n7148 = x17 & n7147 ;
  assign n7149 = x17 & ~n7148 ;
  assign n7150 = ( n7147 & ~n7148 ) | ( n7147 & n7149 ) | ( ~n7148 & n7149 ) ;
  assign n7151 = n7140 & n7150 ;
  assign n7152 = ~n2606 & n5069 ;
  assign n7153 = ~n2455 & n5070 ;
  assign n7154 = n7152 | n7153 ;
  assign n7155 = ~n2375 & n5083 ;
  assign n7156 = n7154 | n7155 ;
  assign n7157 = n5074 | n7156 ;
  assign n7158 = ( ~n5528 & n7156 ) | ( ~n5528 & n7157 ) | ( n7156 & n7157 ) ;
  assign n7159 = ~x17 & n7158 ;
  assign n7160 = x17 & ~n7158 ;
  assign n7161 = n7159 | n7160 ;
  assign n7162 = n6791 | n6800 ;
  assign n7163 = ~n6801 & n7162 ;
  assign n7164 = n7161 & n7163 ;
  assign n7165 = n7161 | n7163 ;
  assign n7166 = ~n7164 & n7165 ;
  assign n7167 = x20 & ~n6796 ;
  assign n7168 = n6798 | n7167 ;
  assign n7169 = n6799 | n7168 ;
  assign n7170 = ~n6800 & n7169 ;
  assign n7171 = ~n2455 & n5083 ;
  assign n7172 = ~n2606 & n5070 ;
  assign n7173 = n7171 | n7172 ;
  assign n7174 = n2569 & n5069 ;
  assign n7175 = n7173 | n7174 ;
  assign n7176 = n5074 | n7175 ;
  assign n7177 = ( ~n5732 & n7175 ) | ( ~n5732 & n7176 ) | ( n7175 & n7176 ) ;
  assign n7178 = ~x17 & n7177 ;
  assign n7179 = x17 | n7178 ;
  assign n7180 = ( ~n7177 & n7178 ) | ( ~n7177 & n7179 ) | ( n7178 & n7179 ) ;
  assign n7181 = n7170 & n7180 ;
  assign n7182 = ~n2764 & n5069 ;
  assign n7183 = ~n2672 & n5070 ;
  assign n7184 = n7182 | n7183 ;
  assign n7185 = n2569 & n5083 ;
  assign n7186 = n7184 | n7185 ;
  assign n7187 = ( n5074 & n5584 ) | ( n5074 & n7186 ) | ( n5584 & n7186 ) ;
  assign n7188 = ( x17 & ~n7186 ) | ( x17 & n7187 ) | ( ~n7186 & n7187 ) ;
  assign n7189 = ~n7187 & n7188 ;
  assign n7190 = n7186 | n7188 ;
  assign n7191 = ( ~x17 & n7189 ) | ( ~x17 & n7190 ) | ( n7189 & n7190 ) ;
  assign n7192 = ~n2764 & n5070 ;
  assign n7193 = ~n2672 & n5083 ;
  assign n7194 = n7192 | n7193 ;
  assign n7195 = n5074 | n7194 ;
  assign n7196 = ( n5932 & n7194 ) | ( n5932 & n7195 ) | ( n7194 & n7195 ) ;
  assign n7197 = ~n2764 & n5064 ;
  assign n7198 = x17 & ~n7197 ;
  assign n7199 = ~x17 & n7196 ;
  assign n7200 = ( ~n7196 & n7198 ) | ( ~n7196 & n7199 ) | ( n7198 & n7199 ) ;
  assign n7201 = n7191 & n7200 ;
  assign n7202 = n6797 & n7201 ;
  assign n7203 = n7201 & ~n7202 ;
  assign n7204 = n6797 & ~n7201 ;
  assign n7205 = n7203 | n7204 ;
  assign n7206 = ~n2606 & n5083 ;
  assign n7207 = ~n2672 & n5069 ;
  assign n7208 = n7206 | n7207 ;
  assign n7209 = n2569 & n5070 ;
  assign n7210 = n7208 | n7209 ;
  assign n7211 = n5074 | n7210 ;
  assign n7212 = ( n5716 & n7210 ) | ( n5716 & n7211 ) | ( n7210 & n7211 ) ;
  assign n7213 = x17 & n7212 ;
  assign n7214 = x17 & ~n7213 ;
  assign n7215 = ( n7212 & ~n7213 ) | ( n7212 & n7214 ) | ( ~n7213 & n7214 ) ;
  assign n7216 = n7205 & n7215 ;
  assign n7217 = n7202 | n7216 ;
  assign n7218 = n7170 | n7180 ;
  assign n7219 = ~n7181 & n7218 ;
  assign n7220 = n7217 & n7219 ;
  assign n7221 = n7181 | n7220 ;
  assign n7222 = n7166 & n7221 ;
  assign n7223 = n7164 | n7222 ;
  assign n7224 = n7140 | n7150 ;
  assign n7225 = ~n7151 & n7224 ;
  assign n7226 = n7223 & n7225 ;
  assign n7227 = n7151 | n7226 ;
  assign n7228 = n7137 & ~n7138 ;
  assign n7229 = ( n7127 & ~n7138 ) | ( n7127 & n7228 ) | ( ~n7138 & n7228 ) ;
  assign n7230 = n7227 & n7229 ;
  assign n7231 = n7138 | n7230 ;
  assign n7232 = ( n7115 & n7125 ) | ( n7115 & n7231 ) | ( n7125 & n7231 ) ;
  assign n7233 = n7113 & n7232 ;
  assign n7234 = n7110 | n7233 ;
  assign n7235 = n7086 | n7096 ;
  assign n7236 = ~n7097 & n7235 ;
  assign n7237 = n7234 & n7236 ;
  assign n7238 = n7097 | n7237 ;
  assign n7239 = n7084 & n7238 ;
  assign n7240 = n7082 | n7239 ;
  assign n7241 = n7069 & n7240 ;
  assign n7242 = n7066 | n7241 ;
  assign n7243 = n7053 & n7242 ;
  assign n7244 = n7051 | n7243 ;
  assign n7245 = n7027 & ~n7038 ;
  assign n7246 = ~n7027 & n7037 ;
  assign n7247 = n7245 | n7246 ;
  assign n7248 = n7244 & n7247 ;
  assign n7249 = n7014 | n7024 ;
  assign n7250 = ~n7025 & n7249 ;
  assign n7251 = ( n7038 & n7248 ) | ( n7038 & n7250 ) | ( n7248 & n7250 ) ;
  assign n7252 = n7025 | n7251 ;
  assign n7253 = n7012 & n7252 ;
  assign n7254 = n7009 | n7253 ;
  assign n7255 = n6984 | n6995 ;
  assign n7256 = ( ~n6994 & n6995 ) | ( ~n6994 & n7255 ) | ( n6995 & n7255 ) ;
  assign n7257 = n7254 & ~n7256 ;
  assign n7258 = n6995 | n7257 ;
  assign n7259 = n6970 | n6981 ;
  assign n7260 = ( ~n6980 & n6981 ) | ( ~n6980 & n7259 ) | ( n6981 & n7259 ) ;
  assign n7261 = n7258 & ~n7260 ;
  assign n7262 = n6981 | n7261 ;
  assign n7263 = n6967 & n7262 ;
  assign n7264 = n6964 | n7263 ;
  assign n7265 = ~n6950 & n7264 ;
  assign n7266 = n6948 | n7265 ;
  assign n7267 = n6935 & n7266 ;
  assign n7268 = n6932 | n7267 ;
  assign n7269 = n6914 | n6917 ;
  assign n7270 = ~n6918 & n7269 ;
  assign n7271 = n7268 & n7270 ;
  assign n7272 = n6918 | n7271 ;
  assign n7273 = n6904 & n7272 ;
  assign n7274 = n6904 | n7272 ;
  assign n7275 = ~n7273 & n7274 ;
  assign n7276 = n1233 & n5384 ;
  assign n7277 = ~n35 & n5382 ;
  assign n7278 = n3349 & n7277 ;
  assign n7279 = n7276 | n7278 ;
  assign n7280 = n35 & ~n38 ;
  assign n7281 = ~n3255 & n7280 ;
  assign n7282 = n7279 | n7281 ;
  assign n7283 = n39 | n7282 ;
  assign n7284 = ( ~n4470 & n7282 ) | ( ~n4470 & n7283 ) | ( n7282 & n7283 ) ;
  assign n7285 = ~x14 & n7284 ;
  assign n7286 = x14 | n7285 ;
  assign n7287 = ( ~n7284 & n7285 ) | ( ~n7284 & n7286 ) | ( n7285 & n7286 ) ;
  assign n7288 = n7275 & n7287 ;
  assign n7289 = n7273 | n7288 ;
  assign n7290 = ~x9 & x10 ;
  assign n7291 = x9 & ~x10 ;
  assign n7292 = n7290 | n7291 ;
  assign n7293 = x10 & ~x11 ;
  assign n7294 = ~x10 & x11 ;
  assign n7295 = n7293 | n7294 ;
  assign n7296 = x8 & ~x9 ;
  assign n7297 = ~x8 & x9 ;
  assign n7298 = n7296 | n7297 ;
  assign n7299 = n7295 & ~n7298 ;
  assign n7300 = ~n7292 & n7299 ;
  assign n7301 = n904 & n7300 ;
  assign n7302 = n7292 & ~n7298 ;
  assign n7303 = n778 & n7302 ;
  assign n7304 = n7301 | n7303 ;
  assign n7305 = ~n7295 & n7298 ;
  assign n7306 = ~n3596 & n7305 ;
  assign n7307 = n7304 | n7306 ;
  assign n7308 = n7295 & n7298 ;
  assign n7309 = n7307 | n7308 ;
  assign n7310 = ( ~n4649 & n7307 ) | ( ~n4649 & n7309 ) | ( n7307 & n7309 ) ;
  assign n7311 = ~x11 & n7310 ;
  assign n7312 = x11 | n7311 ;
  assign n7313 = ( ~n7310 & n7311 ) | ( ~n7310 & n7312 ) | ( n7311 & n7312 ) ;
  assign n7314 = ~n1014 & n7280 ;
  assign n7315 = n3349 & n5384 ;
  assign n7316 = ~n3255 & n7277 ;
  assign n7317 = n7315 | n7316 ;
  assign n7318 = n7314 | n7317 ;
  assign n7319 = n39 | n7318 ;
  assign n7320 = ( n4742 & n7318 ) | ( n4742 & n7319 ) | ( n7318 & n7319 ) ;
  assign n7321 = x14 & n7320 ;
  assign n7322 = x14 & ~n7321 ;
  assign n7323 = ( n7320 & ~n7321 ) | ( n7320 & n7322 ) | ( ~n7321 & n7322 ) ;
  assign n7324 = n6889 | n6902 ;
  assign n7325 = n1327 & n5069 ;
  assign n7326 = ~n1151 & n5070 ;
  assign n7327 = n7325 | n7326 ;
  assign n7328 = n1233 & n5083 ;
  assign n7329 = n7327 | n7328 ;
  assign n7330 = n5074 | n7329 ;
  assign n7331 = ( ~n4615 & n7329 ) | ( ~n4615 & n7330 ) | ( n7329 & n7330 ) ;
  assign n7332 = ~x17 & n7331 ;
  assign n7333 = x17 | n7332 ;
  assign n7334 = ( ~n7331 & n7332 ) | ( ~n7331 & n7333 ) | ( n7332 & n7333 ) ;
  assign n7335 = n6570 | n6583 ;
  assign n7336 = ~n1411 & n4776 ;
  assign n7337 = n3178 & n4778 ;
  assign n7338 = n7336 | n7337 ;
  assign n7339 = n3104 & n4781 ;
  assign n7340 = n7338 | n7339 ;
  assign n7341 = n4784 | n7340 ;
  assign n7342 = ( n4449 & n7340 ) | ( n4449 & n7341 ) | ( n7340 & n7341 ) ;
  assign n7343 = x20 & n7342 ;
  assign n7344 = x20 & ~n7343 ;
  assign n7345 = ( n7342 & ~n7343 ) | ( n7342 & n7344 ) | ( ~n7343 & n7344 ) ;
  assign n7346 = n6298 | n6311 ;
  assign n7347 = n1532 & n4551 ;
  assign n7348 = n3030 & n4546 ;
  assign n7349 = ~n2939 & n4548 ;
  assign n7350 = n7348 | n7349 ;
  assign n7351 = n7347 | n7350 ;
  assign n7352 = n4554 | n7351 ;
  assign n7353 = ( ~n4193 & n7351 ) | ( ~n4193 & n7352 ) | ( n7351 & n7352 ) ;
  assign n7354 = ~x23 & n7353 ;
  assign n7355 = x23 | n7354 ;
  assign n7356 = ( ~n7353 & n7354 ) | ( ~n7353 & n7355 ) | ( n7354 & n7355 ) ;
  assign n7357 = n5273 & ~n5277 ;
  assign n7358 = n5210 | n5277 ;
  assign n7359 = n5275 & ~n7358 ;
  assign n7360 = n7357 | n7359 ;
  assign n7361 = ~n2103 & n3744 ;
  assign n7362 = n2013 & n3727 ;
  assign n7363 = n2193 & n3639 ;
  assign n7364 = n7362 | n7363 ;
  assign n7365 = n3636 | n7364 ;
  assign n7366 = ( ~n5836 & n7364 ) | ( ~n5836 & n7365 ) | ( n7364 & n7365 ) ;
  assign n7367 = n7361 | n7366 ;
  assign n7368 = n7360 & n7367 ;
  assign n7369 = n7360 & ~n7368 ;
  assign n7370 = ~n7360 & n7367 ;
  assign n7371 = n7369 | n7370 ;
  assign n7372 = n6063 | n6075 ;
  assign n7373 = n7371 & ~n7372 ;
  assign n7374 = n1803 & n4048 ;
  assign n7375 = ~n1944 & n4043 ;
  assign n7376 = n7374 | n7375 ;
  assign n7377 = ~n1880 & n4045 ;
  assign n7378 = n7376 | n7377 ;
  assign n7379 = n4051 | n7378 ;
  assign n7380 = ( n4905 & n7378 ) | ( n4905 & n7379 ) | ( n7378 & n7379 ) ;
  assign n7381 = x29 & n7380 ;
  assign n7382 = x29 & ~n7381 ;
  assign n7383 = ( n7380 & ~n7381 ) | ( n7380 & n7382 ) | ( ~n7381 & n7382 ) ;
  assign n7384 = n7373 | n7383 ;
  assign n7385 = ~n7371 & n7372 ;
  assign n7386 = n7384 | n7385 ;
  assign n7387 = ( n7373 & n7383 ) | ( n7373 & n7385 ) | ( n7383 & n7385 ) ;
  assign n7388 = n7386 & ~n7387 ;
  assign n7389 = ~n2873 & n4479 ;
  assign n7390 = ~n1733 & n4481 ;
  assign n7391 = n7389 | n7390 ;
  assign n7392 = n1625 & n4484 ;
  assign n7393 = n7391 | n7392 ;
  assign n7394 = n4487 | n7393 ;
  assign n7395 = ( n4260 & n7393 ) | ( n4260 & n7394 ) | ( n7393 & n7394 ) ;
  assign n7396 = x26 & n7395 ;
  assign n7397 = x26 & ~n7396 ;
  assign n7398 = ( n7395 & ~n7396 ) | ( n7395 & n7397 ) | ( ~n7396 & n7397 ) ;
  assign n7399 = n7388 & ~n7398 ;
  assign n7400 = n7398 | n7399 ;
  assign n7401 = ( ~n7388 & n7399 ) | ( ~n7388 & n7400 ) | ( n7399 & n7400 ) ;
  assign n7402 = n6080 | n6092 ;
  assign n7403 = ( n7356 & n7401 ) | ( n7356 & ~n7402 ) | ( n7401 & ~n7402 ) ;
  assign n7404 = ( ~n7401 & n7402 ) | ( ~n7401 & n7403 ) | ( n7402 & n7403 ) ;
  assign n7405 = ( ~n7356 & n7403 ) | ( ~n7356 & n7404 ) | ( n7403 & n7404 ) ;
  assign n7406 = ( n7345 & ~n7346 ) | ( n7345 & n7405 ) | ( ~n7346 & n7405 ) ;
  assign n7407 = ( n7346 & ~n7405 ) | ( n7346 & n7406 ) | ( ~n7405 & n7406 ) ;
  assign n7408 = ( ~n7345 & n7406 ) | ( ~n7345 & n7407 ) | ( n7406 & n7407 ) ;
  assign n7409 = ( n7334 & ~n7335 ) | ( n7334 & n7408 ) | ( ~n7335 & n7408 ) ;
  assign n7410 = ( n7335 & ~n7408 ) | ( n7335 & n7409 ) | ( ~n7408 & n7409 ) ;
  assign n7411 = ( ~n7334 & n7409 ) | ( ~n7334 & n7410 ) | ( n7409 & n7410 ) ;
  assign n7412 = ( n7323 & ~n7324 ) | ( n7323 & n7411 ) | ( ~n7324 & n7411 ) ;
  assign n7413 = ( n7324 & ~n7411 ) | ( n7324 & n7412 ) | ( ~n7411 & n7412 ) ;
  assign n7414 = ( ~n7323 & n7412 ) | ( ~n7323 & n7413 ) | ( n7412 & n7413 ) ;
  assign n7415 = ( n7289 & n7313 ) | ( n7289 & n7414 ) | ( n7313 & n7414 ) ;
  assign n7416 = n778 & n7300 ;
  assign n7417 = ~n3596 & n7302 ;
  assign n7418 = n7416 | n7417 ;
  assign n7419 = n3504 & n7305 ;
  assign n7420 = n7418 | n7419 ;
  assign n7421 = n7308 | n7420 ;
  assign n7422 = ( ~n5040 & n7420 ) | ( ~n5040 & n7421 ) | ( n7420 & n7421 ) ;
  assign n7423 = ~x11 & n7422 ;
  assign n7424 = x11 | n7423 ;
  assign n7425 = ( ~n7422 & n7423 ) | ( ~n7422 & n7424 ) | ( n7423 & n7424 ) ;
  assign n7426 = ( n7323 & n7324 ) | ( n7323 & n7411 ) | ( n7324 & n7411 ) ;
  assign n7427 = ~n1014 & n7277 ;
  assign n7428 = ~n3255 & n5384 ;
  assign n7429 = n7427 | n7428 ;
  assign n7430 = n904 & n7280 ;
  assign n7431 = n7429 | n7430 ;
  assign n7432 = n39 | n7431 ;
  assign n7433 = ( n4632 & n7431 ) | ( n4632 & n7432 ) | ( n7431 & n7432 ) ;
  assign n7434 = x14 & n7433 ;
  assign n7435 = x14 & ~n7434 ;
  assign n7436 = ( n7433 & ~n7434 ) | ( n7433 & n7435 ) | ( ~n7434 & n7435 ) ;
  assign n7437 = ( n7334 & n7335 ) | ( n7334 & n7408 ) | ( n7335 & n7408 ) ;
  assign n7438 = ~n1151 & n5069 ;
  assign n7439 = n1233 & n5070 ;
  assign n7440 = n7438 | n7439 ;
  assign n7441 = n3349 & n5083 ;
  assign n7442 = n7440 | n7441 ;
  assign n7443 = n5074 | n7442 ;
  assign n7444 = ( n4518 & n7442 ) | ( n4518 & n7443 ) | ( n7442 & n7443 ) ;
  assign n7445 = x17 & n7444 ;
  assign n7446 = x17 & ~n7445 ;
  assign n7447 = ( n7444 & ~n7445 ) | ( n7444 & n7446 ) | ( ~n7445 & n7446 ) ;
  assign n7448 = ( n7356 & n7401 ) | ( n7356 & n7402 ) | ( n7401 & n7402 ) ;
  assign n7449 = ~n1944 & n3744 ;
  assign n7450 = ~n2103 & n3727 ;
  assign n7451 = n2013 & n3639 ;
  assign n7452 = n7450 | n7451 ;
  assign n7453 = n3636 | n7452 ;
  assign n7454 = ( n6041 & n7452 ) | ( n6041 & n7453 ) | ( n7452 & n7453 ) ;
  assign n7455 = n7449 | n7454 ;
  assign n7456 = ( n5179 & n5212 ) | ( n5179 & n7358 ) | ( n5212 & n7358 ) ;
  assign n7457 = ( ~n5179 & n5212 ) | ( ~n5179 & n7358 ) | ( n5212 & n7358 ) ;
  assign n7458 = ( n5179 & ~n7456 ) | ( n5179 & n7457 ) | ( ~n7456 & n7457 ) ;
  assign n7459 = n7455 & ~n7458 ;
  assign n7460 = ~n7455 & n7458 ;
  assign n7461 = n7459 | n7460 ;
  assign n7462 = ( n7368 & n7372 ) | ( n7368 & ~n7385 ) | ( n7372 & ~n7385 ) ;
  assign n7463 = ~n7461 & n7462 ;
  assign n7464 = n7461 & ~n7462 ;
  assign n7465 = n7463 | n7464 ;
  assign n7466 = ~n2873 & n4048 ;
  assign n7467 = n1803 & n4045 ;
  assign n7468 = n7466 | n7467 ;
  assign n7469 = ~n1880 & n4043 ;
  assign n7470 = n7468 | n7469 ;
  assign n7471 = n4051 | n7470 ;
  assign n7472 = ( n5139 & n7470 ) | ( n5139 & n7471 ) | ( n7470 & n7471 ) ;
  assign n7473 = x29 & n7472 ;
  assign n7474 = x29 & ~n7473 ;
  assign n7475 = ( n7472 & ~n7473 ) | ( n7472 & n7474 ) | ( ~n7473 & n7474 ) ;
  assign n7476 = ~n7465 & n7475 ;
  assign n7477 = n7465 & ~n7475 ;
  assign n7478 = n7476 | n7477 ;
  assign n7479 = ~n1733 & n4479 ;
  assign n7480 = n1625 & n4481 ;
  assign n7481 = n7479 | n7480 ;
  assign n7482 = n3030 & n4484 ;
  assign n7483 = n7481 | n7482 ;
  assign n7484 = n4487 | n7483 ;
  assign n7485 = ( ~n4578 & n7483 ) | ( ~n4578 & n7484 ) | ( n7483 & n7484 ) ;
  assign n7486 = ~x26 & n7485 ;
  assign n7487 = x26 | n7486 ;
  assign n7488 = ( ~n7485 & n7486 ) | ( ~n7485 & n7487 ) | ( n7486 & n7487 ) ;
  assign n7489 = ~n7478 & n7488 ;
  assign n7490 = n7478 | n7489 ;
  assign n7491 = n7478 & n7488 ;
  assign n7492 = ( n7386 & n7387 ) | ( n7386 & n7398 ) | ( n7387 & n7398 ) ;
  assign n7493 = n7491 | n7492 ;
  assign n7494 = n7490 & ~n7493 ;
  assign n7495 = ( ~n7490 & n7491 ) | ( ~n7490 & n7492 ) | ( n7491 & n7492 ) ;
  assign n7496 = n7494 | n7495 ;
  assign n7497 = n1532 & n4548 ;
  assign n7498 = ~n1411 & n4551 ;
  assign n7499 = ~n2939 & n4546 ;
  assign n7500 = n7498 | n7499 ;
  assign n7501 = n7497 | n7500 ;
  assign n7502 = n4554 | n7501 ;
  assign n7503 = ( ~n3930 & n7501 ) | ( ~n3930 & n7502 ) | ( n7501 & n7502 ) ;
  assign n7504 = ~x23 & n7503 ;
  assign n7505 = x23 | n7504 ;
  assign n7506 = ( ~n7503 & n7504 ) | ( ~n7503 & n7505 ) | ( n7504 & n7505 ) ;
  assign n7507 = ( n7448 & n7496 ) | ( n7448 & ~n7506 ) | ( n7496 & ~n7506 ) ;
  assign n7508 = ( ~n7496 & n7506 ) | ( ~n7496 & n7507 ) | ( n7506 & n7507 ) ;
  assign n7509 = ( ~n7448 & n7507 ) | ( ~n7448 & n7508 ) | ( n7507 & n7508 ) ;
  assign n7510 = n3178 & n4776 ;
  assign n7511 = n3104 & n4778 ;
  assign n7512 = n7510 | n7511 ;
  assign n7513 = n1327 & n4781 ;
  assign n7514 = n7512 | n7513 ;
  assign n7515 = n4784 | n7514 ;
  assign n7516 = ( n4501 & n7514 ) | ( n4501 & n7515 ) | ( n7514 & n7515 ) ;
  assign n7517 = x20 & n7516 ;
  assign n7518 = x20 & ~n7517 ;
  assign n7519 = ( n7516 & ~n7517 ) | ( n7516 & n7518 ) | ( ~n7517 & n7518 ) ;
  assign n7520 = n7509 | n7519 ;
  assign n7521 = ~n7519 & n7520 ;
  assign n7522 = ( ~n7509 & n7520 ) | ( ~n7509 & n7521 ) | ( n7520 & n7521 ) ;
  assign n7523 = ( n7345 & n7346 ) | ( n7345 & n7405 ) | ( n7346 & n7405 ) ;
  assign n7524 = ( n7447 & n7522 ) | ( n7447 & ~n7523 ) | ( n7522 & ~n7523 ) ;
  assign n7525 = ( ~n7522 & n7523 ) | ( ~n7522 & n7524 ) | ( n7523 & n7524 ) ;
  assign n7526 = ( ~n7447 & n7524 ) | ( ~n7447 & n7525 ) | ( n7524 & n7525 ) ;
  assign n7527 = ( n7436 & ~n7437 ) | ( n7436 & n7526 ) | ( ~n7437 & n7526 ) ;
  assign n7528 = ( n7437 & ~n7526 ) | ( n7437 & n7527 ) | ( ~n7526 & n7527 ) ;
  assign n7529 = ( ~n7436 & n7527 ) | ( ~n7436 & n7528 ) | ( n7527 & n7528 ) ;
  assign n7530 = ( n7425 & ~n7426 ) | ( n7425 & n7529 ) | ( ~n7426 & n7529 ) ;
  assign n7531 = ( n7426 & ~n7529 ) | ( n7426 & n7530 ) | ( ~n7529 & n7530 ) ;
  assign n7532 = ( ~n7425 & n7530 ) | ( ~n7425 & n7531 ) | ( n7530 & n7531 ) ;
  assign n7533 = ~n3431 & n5512 ;
  assign n7534 = ~n589 & n5508 ;
  assign n7535 = n7533 | n7534 ;
  assign n7536 = ~n672 & n5503 ;
  assign n7537 = n7535 | n7536 ;
  assign n7538 = n5515 | n7537 ;
  assign n7539 = ( ~n5353 & n7537 ) | ( ~n5353 & n7538 ) | ( n7537 & n7538 ) ;
  assign n7540 = ~x8 & n7539 ;
  assign n7541 = x8 | n7540 ;
  assign n7542 = ( ~n7539 & n7540 ) | ( ~n7539 & n7541 ) | ( n7540 & n7541 ) ;
  assign n7543 = ( ~n7415 & n7532 ) | ( ~n7415 & n7542 ) | ( n7532 & n7542 ) ;
  assign n7544 = ( n7415 & ~n7532 ) | ( n7415 & n7543 ) | ( ~n7532 & n7543 ) ;
  assign n7545 = n5520 & n7544 ;
  assign n7546 = n7544 & ~n7545 ;
  assign n7547 = ~n3596 & n7300 ;
  assign n7548 = n3504 & n7302 ;
  assign n7549 = n7547 | n7548 ;
  assign n7550 = ~n3431 & n7305 ;
  assign n7551 = n7549 | n7550 ;
  assign n7552 = n7308 | n7551 ;
  assign n7553 = ( ~n4798 & n7551 ) | ( ~n4798 & n7552 ) | ( n7551 & n7552 ) ;
  assign n7554 = ~x11 & n7553 ;
  assign n7555 = x11 | n7554 ;
  assign n7556 = ( ~n7553 & n7554 ) | ( ~n7553 & n7555 ) | ( n7554 & n7555 ) ;
  assign n7557 = n7531 & n7556 ;
  assign n7558 = n7531 | n7556 ;
  assign n7559 = ~n7557 & n7558 ;
  assign n7560 = ( n5152 & ~n5278 ) | ( n5152 & n5288 ) | ( ~n5278 & n5288 ) ;
  assign n7561 = ( ~n5152 & n5278 ) | ( ~n5152 & n7560 ) | ( n5278 & n7560 ) ;
  assign n7562 = ( ~n5288 & n7560 ) | ( ~n5288 & n7561 ) | ( n7560 & n7561 ) ;
  assign n7563 = n7459 | n7562 ;
  assign n7564 = n7463 | n7563 ;
  assign n7565 = ( n7459 & n7463 ) | ( n7459 & n7562 ) | ( n7463 & n7562 ) ;
  assign n7566 = n7564 & ~n7565 ;
  assign n7567 = n1803 & n4043 ;
  assign n7568 = ~n2873 & n4045 ;
  assign n7569 = n7567 | n7568 ;
  assign n7570 = ~n1733 & n4048 ;
  assign n7571 = n7569 | n7570 ;
  assign n7572 = n4051 | n7571 ;
  assign n7573 = ( ~n4985 & n7571 ) | ( ~n4985 & n7572 ) | ( n7571 & n7572 ) ;
  assign n7574 = ~x29 & n7573 ;
  assign n7575 = x29 | n7574 ;
  assign n7576 = ( ~n7573 & n7574 ) | ( ~n7573 & n7575 ) | ( n7574 & n7575 ) ;
  assign n7577 = n7566 & n7576 ;
  assign n7578 = n7566 & ~n7577 ;
  assign n7579 = ~n7566 & n7576 ;
  assign n7580 = n1625 & n4479 ;
  assign n7581 = n3030 & n4481 ;
  assign n7582 = n7580 | n7581 ;
  assign n7583 = ~n2939 & n4484 ;
  assign n7584 = n7582 | n7583 ;
  assign n7585 = n4487 | n7584 ;
  assign n7586 = ( ~n4215 & n7584 ) | ( ~n4215 & n7585 ) | ( n7584 & n7585 ) ;
  assign n7587 = ~x26 & n7586 ;
  assign n7588 = x26 | n7587 ;
  assign n7589 = ( ~n7586 & n7587 ) | ( ~n7586 & n7588 ) | ( n7587 & n7588 ) ;
  assign n7590 = n7579 | n7589 ;
  assign n7591 = n7578 | n7590 ;
  assign n7592 = ( n7578 & n7579 ) | ( n7578 & n7589 ) | ( n7579 & n7589 ) ;
  assign n7593 = n7591 & ~n7592 ;
  assign n7594 = n7476 | n7489 ;
  assign n7595 = n7593 & n7594 ;
  assign n7596 = n7593 | n7594 ;
  assign n7597 = ~n7595 & n7596 ;
  assign n7598 = ~n1411 & n4548 ;
  assign n7599 = n4546 | n7598 ;
  assign n7600 = ( n1532 & n7598 ) | ( n1532 & n7599 ) | ( n7598 & n7599 ) ;
  assign n7601 = n3178 & n4551 ;
  assign n7602 = n7600 | n7601 ;
  assign n7603 = n4554 | n7602 ;
  assign n7604 = ( ~n3750 & n7602 ) | ( ~n3750 & n7603 ) | ( n7602 & n7603 ) ;
  assign n7605 = ~x23 & n7604 ;
  assign n7606 = x23 | n7605 ;
  assign n7607 = ( ~n7604 & n7605 ) | ( ~n7604 & n7606 ) | ( n7605 & n7606 ) ;
  assign n7608 = n7597 & n7607 ;
  assign n7609 = n7597 & ~n7608 ;
  assign n7610 = ~n7597 & n7607 ;
  assign n7611 = ~n7496 & n7506 ;
  assign n7612 = n7495 | n7611 ;
  assign n7613 = n7610 | n7612 ;
  assign n7614 = n7609 | n7613 ;
  assign n7615 = ( n7609 & n7610 ) | ( n7609 & n7612 ) | ( n7610 & n7612 ) ;
  assign n7616 = n7614 & ~n7615 ;
  assign n7617 = n3104 & n4776 ;
  assign n7618 = n1327 & n4778 ;
  assign n7619 = n7617 | n7618 ;
  assign n7620 = ~n1151 & n4781 ;
  assign n7621 = n7619 | n7620 ;
  assign n7622 = n4784 | n7621 ;
  assign n7623 = ( ~n4034 & n7621 ) | ( ~n4034 & n7622 ) | ( n7621 & n7622 ) ;
  assign n7624 = ~x20 & n7623 ;
  assign n7625 = x20 | n7624 ;
  assign n7626 = ( ~n7623 & n7624 ) | ( ~n7623 & n7625 ) | ( n7624 & n7625 ) ;
  assign n7627 = n7616 & n7626 ;
  assign n7628 = n7616 | n7626 ;
  assign n7629 = ~n7627 & n7628 ;
  assign n7630 = ( n7448 & n7519 ) | ( n7448 & n7522 ) | ( n7519 & n7522 ) ;
  assign n7631 = n7629 & n7630 ;
  assign n7632 = n7629 | n7630 ;
  assign n7633 = ~n7631 & n7632 ;
  assign n7634 = n1233 & n5069 ;
  assign n7635 = n3349 & n5070 ;
  assign n7636 = n7634 | n7635 ;
  assign n7637 = ~n3255 & n5083 ;
  assign n7638 = n7636 | n7637 ;
  assign n7639 = n5074 | n7638 ;
  assign n7640 = ( ~n4470 & n7638 ) | ( ~n4470 & n7639 ) | ( n7638 & n7639 ) ;
  assign n7641 = ~x17 & n7640 ;
  assign n7642 = x17 | n7641 ;
  assign n7643 = ( ~n7640 & n7641 ) | ( ~n7640 & n7642 ) | ( n7641 & n7642 ) ;
  assign n7644 = n7633 & n7643 ;
  assign n7645 = n7643 & ~n7644 ;
  assign n7646 = ( n7633 & ~n7644 ) | ( n7633 & n7645 ) | ( ~n7644 & n7645 ) ;
  assign n7647 = n7525 & n7646 ;
  assign n7648 = n7525 | n7646 ;
  assign n7649 = ~n7647 & n7648 ;
  assign n7650 = ~n1014 & n5384 ;
  assign n7651 = n904 & n7277 ;
  assign n7652 = n7650 | n7651 ;
  assign n7653 = n778 & n7280 ;
  assign n7654 = n7652 | n7653 ;
  assign n7655 = n39 | n7654 ;
  assign n7656 = ( ~n4535 & n7654 ) | ( ~n4535 & n7655 ) | ( n7654 & n7655 ) ;
  assign n7657 = ~x14 & n7656 ;
  assign n7658 = x14 | n7657 ;
  assign n7659 = ( ~n7656 & n7657 ) | ( ~n7656 & n7658 ) | ( n7657 & n7658 ) ;
  assign n7660 = n7649 & n7659 ;
  assign n7661 = n7649 | n7659 ;
  assign n7662 = ~n7660 & n7661 ;
  assign n7663 = n7528 & n7662 ;
  assign n7664 = n7528 | n7662 ;
  assign n7665 = ~n7663 & n7664 ;
  assign n7666 = n7559 & n7665 ;
  assign n7667 = n7559 | n7665 ;
  assign n7668 = ~n7666 & n7667 ;
  assign n7669 = n5520 & ~n7544 ;
  assign n7670 = ( n7546 & n7668 ) | ( n7546 & n7669 ) | ( n7668 & n7669 ) ;
  assign n7671 = ~n3634 & n5508 ;
  assign n7672 = n672 & n5512 ;
  assign n7673 = ( n5512 & n7671 ) | ( n5512 & ~n7672 ) | ( n7671 & ~n7672 ) ;
  assign n7674 = n5515 | n7673 ;
  assign n7675 = ( n3726 & n7673 ) | ( n3726 & n7674 ) | ( n7673 & n7674 ) ;
  assign n7676 = x8 & n7675 ;
  assign n7677 = x8 & ~n7676 ;
  assign n7678 = ( n7675 & ~n7676 ) | ( n7675 & n7677 ) | ( ~n7676 & n7677 ) ;
  assign n7679 = n7557 | n7666 ;
  assign n7680 = n7678 & n7679 ;
  assign n7681 = n7678 | n7679 ;
  assign n7682 = ~n7680 & n7681 ;
  assign n7683 = n7644 | n7647 ;
  assign n7684 = n7608 | n7615 ;
  assign n7685 = ~n1411 & n4546 ;
  assign n7686 = n3178 & n4548 ;
  assign n7687 = n7685 | n7686 ;
  assign n7688 = n3104 & n4551 ;
  assign n7689 = n7687 | n7688 ;
  assign n7690 = n4554 | n7689 ;
  assign n7691 = ( n4449 & n7689 ) | ( n4449 & n7690 ) | ( n7689 & n7690 ) ;
  assign n7692 = x23 & n7691 ;
  assign n7693 = x23 & ~n7692 ;
  assign n7694 = ( n7691 & ~n7692 ) | ( n7691 & n7693 ) | ( ~n7692 & n7693 ) ;
  assign n7695 = n7592 | n7595 ;
  assign n7696 = n1532 & n4484 ;
  assign n7697 = n3030 & n4479 ;
  assign n7698 = ~n2939 & n4481 ;
  assign n7699 = n7697 | n7698 ;
  assign n7700 = n7696 | n7699 ;
  assign n7701 = n4487 | n7700 ;
  assign n7702 = ( ~n4193 & n7700 ) | ( ~n4193 & n7701 ) | ( n7700 & n7701 ) ;
  assign n7703 = ~x26 & n7702 ;
  assign n7704 = x26 | n7703 ;
  assign n7705 = ( ~n7702 & n7703 ) | ( ~n7702 & n7704 ) | ( n7703 & n7704 ) ;
  assign n7706 = n5292 & ~n5302 ;
  assign n7707 = n5303 | n7706 ;
  assign n7708 = n7565 | n7577 ;
  assign n7709 = ( n7705 & n7707 ) | ( n7705 & ~n7708 ) | ( n7707 & ~n7708 ) ;
  assign n7710 = ( ~n7707 & n7708 ) | ( ~n7707 & n7709 ) | ( n7708 & n7709 ) ;
  assign n7711 = ( ~n7705 & n7709 ) | ( ~n7705 & n7710 ) | ( n7709 & n7710 ) ;
  assign n7712 = ( n7694 & ~n7695 ) | ( n7694 & n7711 ) | ( ~n7695 & n7711 ) ;
  assign n7713 = ( n7695 & ~n7711 ) | ( n7695 & n7712 ) | ( ~n7711 & n7712 ) ;
  assign n7714 = ( ~n7694 & n7712 ) | ( ~n7694 & n7713 ) | ( n7712 & n7713 ) ;
  assign n7715 = n7684 & ~n7714 ;
  assign n7716 = ~n7684 & n7714 ;
  assign n7717 = n7715 | n7716 ;
  assign n7718 = n1327 & n4776 ;
  assign n7719 = ~n1151 & n4778 ;
  assign n7720 = n7718 | n7719 ;
  assign n7721 = n1233 & n4781 ;
  assign n7722 = n7720 | n7721 ;
  assign n7723 = n4784 | n7722 ;
  assign n7724 = ( ~n4615 & n7722 ) | ( ~n4615 & n7723 ) | ( n7722 & n7723 ) ;
  assign n7725 = ~x20 & n7724 ;
  assign n7726 = x20 | n7725 ;
  assign n7727 = ( ~n7724 & n7725 ) | ( ~n7724 & n7726 ) | ( n7725 & n7726 ) ;
  assign n7728 = ~n7717 & n7727 ;
  assign n7729 = n7717 | n7728 ;
  assign n7730 = n7717 & n7727 ;
  assign n7731 = n7627 | n7631 ;
  assign n7732 = n7730 | n7731 ;
  assign n7733 = n7729 & ~n7732 ;
  assign n7734 = ( ~n7729 & n7730 ) | ( ~n7729 & n7731 ) | ( n7730 & n7731 ) ;
  assign n7735 = n7733 | n7734 ;
  assign n7736 = ~n1014 & n5083 ;
  assign n7737 = n3349 & n5069 ;
  assign n7738 = ~n3255 & n5070 ;
  assign n7739 = n7737 | n7738 ;
  assign n7740 = n7736 | n7739 ;
  assign n7741 = n5074 | n7740 ;
  assign n7742 = ( n4742 & n7740 ) | ( n4742 & n7741 ) | ( n7740 & n7741 ) ;
  assign n7743 = x17 & n7742 ;
  assign n7744 = x17 & ~n7743 ;
  assign n7745 = ( n7742 & ~n7743 ) | ( n7742 & n7744 ) | ( ~n7743 & n7744 ) ;
  assign n7746 = ( n7683 & n7735 ) | ( n7683 & ~n7745 ) | ( n7735 & ~n7745 ) ;
  assign n7747 = ( ~n7735 & n7745 ) | ( ~n7735 & n7746 ) | ( n7745 & n7746 ) ;
  assign n7748 = ( ~n7683 & n7746 ) | ( ~n7683 & n7747 ) | ( n7746 & n7747 ) ;
  assign n7749 = n904 & n5384 ;
  assign n7750 = n778 & n7277 ;
  assign n7751 = n7749 | n7750 ;
  assign n7752 = ~n3596 & n7280 ;
  assign n7753 = n7751 | n7752 ;
  assign n7754 = n39 | n7753 ;
  assign n7755 = ( ~n4649 & n7753 ) | ( ~n4649 & n7754 ) | ( n7753 & n7754 ) ;
  assign n7756 = ~x14 & n7755 ;
  assign n7757 = x14 | n7756 ;
  assign n7758 = ( ~n7755 & n7756 ) | ( ~n7755 & n7757 ) | ( n7756 & n7757 ) ;
  assign n7759 = n7748 | n7758 ;
  assign n7760 = ~n7758 & n7759 ;
  assign n7761 = ( ~n7748 & n7759 ) | ( ~n7748 & n7760 ) | ( n7759 & n7760 ) ;
  assign n7762 = n7660 | n7663 ;
  assign n7763 = n3504 & n7300 ;
  assign n7764 = ~n3431 & n7302 ;
  assign n7765 = n7763 | n7764 ;
  assign n7766 = ~n589 & n7305 ;
  assign n7767 = n7765 | n7766 ;
  assign n7768 = n7308 | n7767 ;
  assign n7769 = ( n4765 & n7767 ) | ( n4765 & n7768 ) | ( n7767 & n7768 ) ;
  assign n7770 = x11 & n7769 ;
  assign n7771 = x11 & ~n7770 ;
  assign n7772 = ( n7769 & ~n7770 ) | ( n7769 & n7771 ) | ( ~n7770 & n7771 ) ;
  assign n7773 = ( n7761 & n7762 ) | ( n7761 & ~n7772 ) | ( n7762 & ~n7772 ) ;
  assign n7774 = ( ~n7762 & n7772 ) | ( ~n7762 & n7773 ) | ( n7772 & n7773 ) ;
  assign n7775 = ( ~n7761 & n7773 ) | ( ~n7761 & n7774 ) | ( n7773 & n7774 ) ;
  assign n7776 = n7682 & ~n7775 ;
  assign n7777 = ~n7682 & n7775 ;
  assign n7778 = n7776 | n7777 ;
  assign n7779 = ( n7545 & n7670 ) | ( n7545 & ~n7778 ) | ( n7670 & ~n7778 ) ;
  assign n7780 = ~n7545 & n7778 ;
  assign n7781 = ~n7670 & n7780 ;
  assign n7782 = n7779 | n7781 ;
  assign n7783 = n6935 | n7266 ;
  assign n7784 = ~n7267 & n7783 ;
  assign n7785 = n1327 & n5384 ;
  assign n7786 = ~n1151 & n7277 ;
  assign n7787 = n7785 | n7786 ;
  assign n7788 = n1233 & n7280 ;
  assign n7789 = n7787 | n7788 ;
  assign n7790 = n39 | n7789 ;
  assign n7791 = ( ~n4615 & n7789 ) | ( ~n4615 & n7790 ) | ( n7789 & n7790 ) ;
  assign n7792 = ~x14 & n7791 ;
  assign n7793 = x14 | n7792 ;
  assign n7794 = ( ~n7791 & n7792 ) | ( ~n7791 & n7793 ) | ( n7792 & n7793 ) ;
  assign n7795 = n7784 & n7794 ;
  assign n7796 = n6950 & ~n7264 ;
  assign n7797 = n7265 | n7796 ;
  assign n7798 = n3104 & n5384 ;
  assign n7799 = n1327 & n7277 ;
  assign n7800 = n7798 | n7799 ;
  assign n7801 = ~n1151 & n7280 ;
  assign n7802 = n7800 | n7801 ;
  assign n7803 = ( n39 & ~n4034 ) | ( n39 & n7802 ) | ( ~n4034 & n7802 ) ;
  assign n7804 = n7802 | n7803 ;
  assign n7805 = ~x14 & n7804 ;
  assign n7806 = x14 | n7805 ;
  assign n7807 = ( ~n7804 & n7805 ) | ( ~n7804 & n7806 ) | ( n7805 & n7806 ) ;
  assign n7808 = ~n7797 & n7807 ;
  assign n7809 = n6967 | n7262 ;
  assign n7810 = ~n7263 & n7809 ;
  assign n7811 = n3178 & n5384 ;
  assign n7812 = n3104 & n7277 ;
  assign n7813 = n7811 | n7812 ;
  assign n7814 = n1327 & n7280 ;
  assign n7815 = n7813 | n7814 ;
  assign n7816 = n39 | n7815 ;
  assign n7817 = ( n4501 & n7815 ) | ( n4501 & n7816 ) | ( n7815 & n7816 ) ;
  assign n7818 = x14 & n7817 ;
  assign n7819 = x14 & ~n7818 ;
  assign n7820 = ( n7817 & ~n7818 ) | ( n7817 & n7819 ) | ( ~n7818 & n7819 ) ;
  assign n7821 = ~n1411 & n5384 ;
  assign n7822 = n3178 & n7277 ;
  assign n7823 = n7821 | n7822 ;
  assign n7824 = n3104 & n7280 ;
  assign n7825 = n7823 | n7824 ;
  assign n7826 = n39 | n7825 ;
  assign n7827 = ( n4449 & n7825 ) | ( n4449 & n7826 ) | ( n7825 & n7826 ) ;
  assign n7828 = x14 & n7827 ;
  assign n7829 = x14 & ~n7828 ;
  assign n7830 = ( n7827 & ~n7828 ) | ( n7827 & n7829 ) | ( ~n7828 & n7829 ) ;
  assign n7831 = ~n1411 & n7277 ;
  assign n7832 = n5384 | n7831 ;
  assign n7833 = ( n1532 & n7831 ) | ( n1532 & n7832 ) | ( n7831 & n7832 ) ;
  assign n7834 = n3178 & n7280 ;
  assign n7835 = n7833 | n7834 ;
  assign n7836 = n39 | n7835 ;
  assign n7837 = ( ~n3750 & n7835 ) | ( ~n3750 & n7836 ) | ( n7835 & n7836 ) ;
  assign n7838 = ~x14 & n7837 ;
  assign n7839 = x14 | n7838 ;
  assign n7840 = ( ~n7837 & n7838 ) | ( ~n7837 & n7839 ) | ( n7838 & n7839 ) ;
  assign n7841 = n7012 | n7252 ;
  assign n7842 = ~n7253 & n7841 ;
  assign n7843 = n1532 & n7277 ;
  assign n7844 = ~n1411 & n7280 ;
  assign n7845 = ~n2939 & n5384 ;
  assign n7846 = n7844 | n7845 ;
  assign n7847 = n7843 | n7846 ;
  assign n7848 = n39 | n7847 ;
  assign n7849 = ( ~n3930 & n7847 ) | ( ~n3930 & n7848 ) | ( n7847 & n7848 ) ;
  assign n7850 = ~x14 & n7849 ;
  assign n7851 = x14 | n7850 ;
  assign n7852 = ( ~n7849 & n7850 ) | ( ~n7849 & n7851 ) | ( n7850 & n7851 ) ;
  assign n7853 = n7038 | n7250 ;
  assign n7854 = n7248 | n7853 ;
  assign n7855 = ~n7251 & n7854 ;
  assign n7856 = n1532 & n7280 ;
  assign n7857 = n3030 & n5384 ;
  assign n7858 = ~n2939 & n7277 ;
  assign n7859 = n7857 | n7858 ;
  assign n7860 = n7856 | n7859 ;
  assign n7861 = n39 | n7860 ;
  assign n7862 = ( ~n4193 & n7860 ) | ( ~n4193 & n7861 ) | ( n7860 & n7861 ) ;
  assign n7863 = ~x14 & n7862 ;
  assign n7864 = x14 | n7863 ;
  assign n7865 = ( ~n7862 & n7863 ) | ( ~n7862 & n7864 ) | ( n7863 & n7864 ) ;
  assign n7866 = n7855 & n7865 ;
  assign n7867 = n7244 & ~n7248 ;
  assign n7868 = n7247 & ~n7248 ;
  assign n7869 = n7867 | n7868 ;
  assign n7870 = n1625 & n5384 ;
  assign n7871 = n3030 & n7277 ;
  assign n7872 = n7870 | n7871 ;
  assign n7873 = ~n2939 & n7280 ;
  assign n7874 = n7872 | n7873 ;
  assign n7875 = n39 | n7874 ;
  assign n7876 = ( ~n4215 & n7874 ) | ( ~n4215 & n7875 ) | ( n7874 & n7875 ) ;
  assign n7877 = ~x14 & n7876 ;
  assign n7878 = x14 | n7877 ;
  assign n7879 = ( ~n7876 & n7877 ) | ( ~n7876 & n7878 ) | ( n7877 & n7878 ) ;
  assign n7880 = n7869 & n7879 ;
  assign n7881 = n7869 & ~n7880 ;
  assign n7882 = ~n7869 & n7879 ;
  assign n7883 = n7881 | n7882 ;
  assign n7884 = n7053 | n7242 ;
  assign n7885 = ~n7243 & n7884 ;
  assign n7886 = ~n1733 & n5384 ;
  assign n7887 = n1625 & n7277 ;
  assign n7888 = n7886 | n7887 ;
  assign n7889 = n3030 & n7280 ;
  assign n7890 = n7888 | n7889 ;
  assign n7891 = n39 | n7890 ;
  assign n7892 = ( ~n4578 & n7890 ) | ( ~n4578 & n7891 ) | ( n7890 & n7891 ) ;
  assign n7893 = ~x14 & n7892 ;
  assign n7894 = x14 | n7893 ;
  assign n7895 = ( ~n7892 & n7893 ) | ( ~n7892 & n7894 ) | ( n7893 & n7894 ) ;
  assign n7896 = n7885 & n7895 ;
  assign n7897 = n7069 | n7240 ;
  assign n7898 = ~n7241 & n7897 ;
  assign n7899 = ~n2873 & n5384 ;
  assign n7900 = ~n1733 & n7277 ;
  assign n7901 = n7899 | n7900 ;
  assign n7902 = n1625 & n7280 ;
  assign n7903 = n7901 | n7902 ;
  assign n7904 = n39 | n7903 ;
  assign n7905 = ( n4260 & n7903 ) | ( n4260 & n7904 ) | ( n7903 & n7904 ) ;
  assign n7906 = x14 & n7905 ;
  assign n7907 = x14 & ~n7906 ;
  assign n7908 = ( n7905 & ~n7906 ) | ( n7905 & n7907 ) | ( ~n7906 & n7907 ) ;
  assign n7909 = n7898 & n7908 ;
  assign n7910 = n7084 | n7238 ;
  assign n7911 = ~n7239 & n7910 ;
  assign n7912 = n1803 & n5384 ;
  assign n7913 = ~n2873 & n7277 ;
  assign n7914 = n7912 | n7913 ;
  assign n7915 = ~n1733 & n7280 ;
  assign n7916 = n7914 | n7915 ;
  assign n7917 = n39 | n7916 ;
  assign n7918 = ( ~n4985 & n7916 ) | ( ~n4985 & n7917 ) | ( n7916 & n7917 ) ;
  assign n7919 = ~x14 & n7918 ;
  assign n7920 = x14 | n7919 ;
  assign n7921 = ( ~n7918 & n7919 ) | ( ~n7918 & n7920 ) | ( n7919 & n7920 ) ;
  assign n7922 = n7911 & n7921 ;
  assign n7923 = n7234 | n7236 ;
  assign n7924 = ~n7237 & n7923 ;
  assign n7925 = ~n2873 & n7280 ;
  assign n7926 = n1803 & n7277 ;
  assign n7927 = n7925 | n7926 ;
  assign n7928 = ~n1880 & n5384 ;
  assign n7929 = n7927 | n7928 ;
  assign n7930 = n39 | n7929 ;
  assign n7931 = ( n5139 & n7929 ) | ( n5139 & n7930 ) | ( n7929 & n7930 ) ;
  assign n7932 = x14 & n7931 ;
  assign n7933 = x14 & ~n7932 ;
  assign n7934 = ( n7931 & ~n7932 ) | ( n7931 & n7933 ) | ( ~n7932 & n7933 ) ;
  assign n7935 = n7924 & n7934 ;
  assign n7936 = n7934 & ~n7935 ;
  assign n7937 = ( n7924 & ~n7935 ) | ( n7924 & n7936 ) | ( ~n7935 & n7936 ) ;
  assign n7938 = n1803 & n7280 ;
  assign n7939 = ~n1944 & n5384 ;
  assign n7940 = n7938 | n7939 ;
  assign n7941 = ~n1880 & n7277 ;
  assign n7942 = n7940 | n7941 ;
  assign n7943 = n39 | n7942 ;
  assign n7944 = ( n4905 & n7942 ) | ( n4905 & n7943 ) | ( n7942 & n7943 ) ;
  assign n7945 = x14 & n7944 ;
  assign n7946 = x14 & ~n7945 ;
  assign n7947 = ( n7944 & ~n7945 ) | ( n7944 & n7946 ) | ( ~n7945 & n7946 ) ;
  assign n7948 = n7113 & ~n7233 ;
  assign n7949 = ( n7232 & ~n7233 ) | ( n7232 & n7948 ) | ( ~n7233 & n7948 ) ;
  assign n7950 = n7947 & n7949 ;
  assign n7951 = n7949 & ~n7950 ;
  assign n7952 = n7947 & ~n7949 ;
  assign n7953 = n7951 | n7952 ;
  assign n7954 = ~n2103 & n5384 ;
  assign n7955 = ~n1944 & n7277 ;
  assign n7956 = n7954 | n7955 ;
  assign n7957 = ~n1880 & n7280 ;
  assign n7958 = n7956 | n7957 ;
  assign n7959 = n39 | n7958 ;
  assign n7960 = ( ~n5281 & n7958 ) | ( ~n5281 & n7959 ) | ( n7958 & n7959 ) ;
  assign n7961 = ~x14 & n7960 ;
  assign n7962 = x14 | n7961 ;
  assign n7963 = ( ~n7960 & n7961 ) | ( ~n7960 & n7962 ) | ( n7961 & n7962 ) ;
  assign n7964 = ( n7115 & n7231 ) | ( n7115 & ~n7232 ) | ( n7231 & ~n7232 ) ;
  assign n7965 = ( n7125 & ~n7232 ) | ( n7125 & n7964 ) | ( ~n7232 & n7964 ) ;
  assign n7966 = n7963 & n7965 ;
  assign n7967 = n7963 | n7965 ;
  assign n7968 = ~n7966 & n7967 ;
  assign n7969 = n7227 | n7229 ;
  assign n7970 = ~n7230 & n7969 ;
  assign n7971 = n2013 & n5384 ;
  assign n7972 = ~n2103 & n7277 ;
  assign n7973 = n7971 | n7972 ;
  assign n7974 = ~n1944 & n7280 ;
  assign n7975 = n7973 | n7974 ;
  assign n7976 = n39 | n7975 ;
  assign n7977 = ( n6041 & n7975 ) | ( n6041 & n7976 ) | ( n7975 & n7976 ) ;
  assign n7978 = x14 & n7977 ;
  assign n7979 = x14 & ~n7978 ;
  assign n7980 = ( n7977 & ~n7978 ) | ( n7977 & n7979 ) | ( ~n7978 & n7979 ) ;
  assign n7981 = n7970 & n7980 ;
  assign n7982 = n7223 | n7225 ;
  assign n7983 = ~n7226 & n7982 ;
  assign n7984 = n2193 & n5384 ;
  assign n7985 = n2013 & n7277 ;
  assign n7986 = n7984 | n7985 ;
  assign n7987 = ~n2103 & n7280 ;
  assign n7988 = n7986 | n7987 ;
  assign n7989 = n39 | n7988 ;
  assign n7990 = ( ~n5836 & n7988 ) | ( ~n5836 & n7989 ) | ( n7988 & n7989 ) ;
  assign n7991 = ~x14 & n7990 ;
  assign n7992 = x14 | n7991 ;
  assign n7993 = ( ~n7990 & n7991 ) | ( ~n7990 & n7992 ) | ( n7991 & n7992 ) ;
  assign n7994 = n7983 & n7993 ;
  assign n7995 = n7983 & ~n7994 ;
  assign n7996 = ~n7983 & n7993 ;
  assign n7997 = n7995 | n7996 ;
  assign n7998 = n7166 | n7221 ;
  assign n7999 = ~n7222 & n7998 ;
  assign n8000 = n2296 & n5384 ;
  assign n8001 = n2193 & n7277 ;
  assign n8002 = n8000 | n8001 ;
  assign n8003 = n2013 & n7280 ;
  assign n8004 = n8002 | n8003 ;
  assign n8005 = n39 | n8004 ;
  assign n8006 = ( n5216 & n8004 ) | ( n5216 & n8005 ) | ( n8004 & n8005 ) ;
  assign n8007 = x14 & n8006 ;
  assign n8008 = x14 & ~n8007 ;
  assign n8009 = ( n8006 & ~n8007 ) | ( n8006 & n8008 ) | ( ~n8007 & n8008 ) ;
  assign n8010 = n7217 | n7219 ;
  assign n8011 = ~n7220 & n8010 ;
  assign n8012 = ~n2375 & n5384 ;
  assign n8013 = n2296 & n7277 ;
  assign n8014 = n8012 | n8013 ;
  assign n8015 = n2193 & n7280 ;
  assign n8016 = n8014 | n8015 ;
  assign n8017 = n39 | n8016 ;
  assign n8018 = ( ~n5879 & n8016 ) | ( ~n5879 & n8017 ) | ( n8016 & n8017 ) ;
  assign n8019 = ~x14 & n8018 ;
  assign n8020 = x14 | n8019 ;
  assign n8021 = ( ~n8018 & n8019 ) | ( ~n8018 & n8020 ) | ( n8019 & n8020 ) ;
  assign n8022 = n8011 & n8021 ;
  assign n8023 = n7205 | n7215 ;
  assign n8024 = ~n7216 & n8023 ;
  assign n8025 = ~n2455 & n5384 ;
  assign n8026 = ~n2375 & n7277 ;
  assign n8027 = n8025 | n8026 ;
  assign n8028 = n2296 & n7280 ;
  assign n8029 = n8027 | n8028 ;
  assign n8030 = n39 | n8029 ;
  assign n8031 = ( n5781 & n8029 ) | ( n5781 & n8030 ) | ( n8029 & n8030 ) ;
  assign n8032 = x14 & n8031 ;
  assign n8033 = x14 & ~n8032 ;
  assign n8034 = ( n8031 & ~n8032 ) | ( n8031 & n8033 ) | ( ~n8032 & n8033 ) ;
  assign n8035 = n8024 & n8034 ;
  assign n8036 = ~n2606 & n5384 ;
  assign n8037 = ~n2455 & n7277 ;
  assign n8038 = n8036 | n8037 ;
  assign n8039 = ~n2375 & n7280 ;
  assign n8040 = n8038 | n8039 ;
  assign n8041 = n39 | n8040 ;
  assign n8042 = ( ~n5528 & n8040 ) | ( ~n5528 & n8041 ) | ( n8040 & n8041 ) ;
  assign n8043 = ~x14 & n8042 ;
  assign n8044 = x14 & ~n8042 ;
  assign n8045 = n8043 | n8044 ;
  assign n8046 = n7191 | n7200 ;
  assign n8047 = ~n7201 & n8046 ;
  assign n8048 = n8045 & n8047 ;
  assign n8049 = n8045 | n8047 ;
  assign n8050 = ~n8048 & n8049 ;
  assign n8051 = x17 & ~n7196 ;
  assign n8052 = n7198 | n8051 ;
  assign n8053 = n7199 | n8052 ;
  assign n8054 = ~n7200 & n8053 ;
  assign n8055 = ~n2455 & n7280 ;
  assign n8056 = ~n2606 & n7277 ;
  assign n8057 = n8055 | n8056 ;
  assign n8058 = n2569 & n5384 ;
  assign n8059 = n8057 | n8058 ;
  assign n8060 = n39 | n8059 ;
  assign n8061 = ( ~n5732 & n8059 ) | ( ~n5732 & n8060 ) | ( n8059 & n8060 ) ;
  assign n8062 = ~x14 & n8061 ;
  assign n8063 = x14 | n8062 ;
  assign n8064 = ( ~n8061 & n8062 ) | ( ~n8061 & n8063 ) | ( n8062 & n8063 ) ;
  assign n8065 = n8054 & n8064 ;
  assign n8066 = ~n2764 & n5384 ;
  assign n8067 = ~n2672 & n7277 ;
  assign n8068 = n8066 | n8067 ;
  assign n8069 = n2569 & n7280 ;
  assign n8070 = n8068 | n8069 ;
  assign n8071 = ( n39 & n5584 ) | ( n39 & n8070 ) | ( n5584 & n8070 ) ;
  assign n8072 = ( x14 & ~n8070 ) | ( x14 & n8071 ) | ( ~n8070 & n8071 ) ;
  assign n8073 = ~n8071 & n8072 ;
  assign n8074 = n8070 | n8072 ;
  assign n8075 = ( ~x14 & n8073 ) | ( ~x14 & n8074 ) | ( n8073 & n8074 ) ;
  assign n8076 = ~n2764 & n7277 ;
  assign n8077 = ~n2672 & n7280 ;
  assign n8078 = n8076 | n8077 ;
  assign n8079 = n39 | n8078 ;
  assign n8080 = ( n5932 & n8078 ) | ( n5932 & n8079 ) | ( n8078 & n8079 ) ;
  assign n8081 = n35 & ~n2764 ;
  assign n8082 = x14 & ~n8081 ;
  assign n8083 = ~x14 & n8080 ;
  assign n8084 = ( ~n8080 & n8082 ) | ( ~n8080 & n8083 ) | ( n8082 & n8083 ) ;
  assign n8085 = n8075 & n8084 ;
  assign n8086 = n7197 & n8085 ;
  assign n8087 = n8085 & ~n8086 ;
  assign n8088 = n7197 & ~n8085 ;
  assign n8089 = n8087 | n8088 ;
  assign n8090 = ~n2606 & n7280 ;
  assign n8091 = ~n2672 & n5384 ;
  assign n8092 = n8090 | n8091 ;
  assign n8093 = n2569 & n7277 ;
  assign n8094 = n8092 | n8093 ;
  assign n8095 = n39 | n8094 ;
  assign n8096 = ( n5716 & n8094 ) | ( n5716 & n8095 ) | ( n8094 & n8095 ) ;
  assign n8097 = x14 & n8096 ;
  assign n8098 = x14 & ~n8097 ;
  assign n8099 = ( n8096 & ~n8097 ) | ( n8096 & n8098 ) | ( ~n8097 & n8098 ) ;
  assign n8100 = n8089 & n8099 ;
  assign n8101 = n8086 | n8100 ;
  assign n8102 = n8054 | n8064 ;
  assign n8103 = ~n8065 & n8102 ;
  assign n8104 = n8101 & n8103 ;
  assign n8105 = n8065 | n8104 ;
  assign n8106 = n8050 & n8105 ;
  assign n8107 = n8048 | n8106 ;
  assign n8108 = n8024 | n8034 ;
  assign n8109 = ~n8035 & n8108 ;
  assign n8110 = n8107 & n8109 ;
  assign n8111 = n8035 | n8110 ;
  assign n8112 = n8021 & ~n8022 ;
  assign n8113 = ( n8011 & ~n8022 ) | ( n8011 & n8112 ) | ( ~n8022 & n8112 ) ;
  assign n8114 = n8111 & n8113 ;
  assign n8115 = n8022 | n8114 ;
  assign n8116 = ( n7999 & n8009 ) | ( n7999 & n8115 ) | ( n8009 & n8115 ) ;
  assign n8117 = n7997 & n8116 ;
  assign n8118 = n7994 | n8117 ;
  assign n8119 = n7970 | n7980 ;
  assign n8120 = ~n7981 & n8119 ;
  assign n8121 = n8118 & n8120 ;
  assign n8122 = n7981 | n8121 ;
  assign n8123 = n7968 & n8122 ;
  assign n8124 = n7966 | n8123 ;
  assign n8125 = n7953 & n8124 ;
  assign n8126 = n7950 | n8125 ;
  assign n8127 = n7937 & n8126 ;
  assign n8128 = n7935 | n8127 ;
  assign n8129 = n7911 & ~n7922 ;
  assign n8130 = ~n7911 & n7921 ;
  assign n8131 = n8129 | n8130 ;
  assign n8132 = n8128 & n8131 ;
  assign n8133 = n7922 | n8132 ;
  assign n8134 = n7898 & ~n7909 ;
  assign n8135 = ~n7898 & n7908 ;
  assign n8136 = n8134 | n8135 ;
  assign n8137 = n8133 & n8136 ;
  assign n8138 = n7885 | n7895 ;
  assign n8139 = ~n7896 & n8138 ;
  assign n8140 = ( n7909 & n8137 ) | ( n7909 & n8139 ) | ( n8137 & n8139 ) ;
  assign n8141 = n7896 | n8140 ;
  assign n8142 = n7883 & n8141 ;
  assign n8143 = n7880 | n8142 ;
  assign n8144 = n7865 & ~n7866 ;
  assign n8145 = ( n7855 & ~n7866 ) | ( n7855 & n8144 ) | ( ~n7866 & n8144 ) ;
  assign n8146 = n8143 & n8145 ;
  assign n8147 = n7866 | n8146 ;
  assign n8148 = ( n7842 & n7852 ) | ( n7842 & n8147 ) | ( n7852 & n8147 ) ;
  assign n8149 = ~n7254 & n7256 ;
  assign n8150 = n7257 | n8149 ;
  assign n8151 = ( n7840 & n8148 ) | ( n7840 & ~n8150 ) | ( n8148 & ~n8150 ) ;
  assign n8152 = ~n7258 & n7260 ;
  assign n8153 = n7261 | n8152 ;
  assign n8154 = ( n7830 & n8151 ) | ( n7830 & ~n8153 ) | ( n8151 & ~n8153 ) ;
  assign n8155 = ( n7810 & n7820 ) | ( n7810 & n8154 ) | ( n7820 & n8154 ) ;
  assign n8156 = n7797 | n7808 ;
  assign n8157 = ( ~n7807 & n7808 ) | ( ~n7807 & n8156 ) | ( n7808 & n8156 ) ;
  assign n8158 = n8155 & ~n8157 ;
  assign n8159 = n7808 | n8158 ;
  assign n8160 = n7784 & ~n7795 ;
  assign n8161 = ~n7784 & n7794 ;
  assign n8162 = n8160 | n8161 ;
  assign n8163 = n8159 & n8162 ;
  assign n8164 = n7795 | n8163 ;
  assign n8165 = n7268 | n7270 ;
  assign n8166 = ~n7271 & n8165 ;
  assign n8167 = ~n1151 & n5384 ;
  assign n8168 = n1233 & n7277 ;
  assign n8169 = n8167 | n8168 ;
  assign n8170 = n3349 & n7280 ;
  assign n8171 = n8169 | n8170 ;
  assign n8172 = n39 | n8171 ;
  assign n8173 = ( n4518 & n8171 ) | ( n4518 & n8172 ) | ( n8171 & n8172 ) ;
  assign n8174 = x14 & n8173 ;
  assign n8175 = x14 & ~n8174 ;
  assign n8176 = ( n8173 & ~n8174 ) | ( n8173 & n8175 ) | ( ~n8174 & n8175 ) ;
  assign n8177 = n8166 & n8176 ;
  assign n8178 = n8166 & ~n8177 ;
  assign n8179 = ~n8166 & n8176 ;
  assign n8180 = n8178 | n8179 ;
  assign n8181 = n8164 & n8180 ;
  assign n8182 = n7275 | n7287 ;
  assign n8183 = ~n7288 & n8182 ;
  assign n8184 = n8177 | n8183 ;
  assign n8185 = n8181 | n8184 ;
  assign n8186 = ( n8177 & n8181 ) | ( n8177 & n8183 ) | ( n8181 & n8183 ) ;
  assign n8187 = n8185 & ~n8186 ;
  assign n8188 = ~n1014 & n7300 ;
  assign n8189 = n904 & n7302 ;
  assign n8190 = n8188 | n8189 ;
  assign n8191 = n778 & n7305 ;
  assign n8192 = n8190 | n8191 ;
  assign n8193 = n7308 | n8192 ;
  assign n8194 = ( ~n4535 & n8192 ) | ( ~n4535 & n8193 ) | ( n8192 & n8193 ) ;
  assign n8195 = ~x11 & n8194 ;
  assign n8196 = x11 | n8195 ;
  assign n8197 = ( ~n8194 & n8195 ) | ( ~n8194 & n8196 ) | ( n8195 & n8196 ) ;
  assign n8198 = n8187 & n8197 ;
  assign n8199 = n8187 | n8197 ;
  assign n8200 = ~n8198 & n8199 ;
  assign n8201 = n8164 & ~n8181 ;
  assign n8202 = n8180 & ~n8181 ;
  assign n8203 = n8201 | n8202 ;
  assign n8204 = ~n1014 & n7302 ;
  assign n8205 = ~n3255 & n7300 ;
  assign n8206 = n8204 | n8205 ;
  assign n8207 = n904 & n7305 ;
  assign n8208 = n8206 | n8207 ;
  assign n8209 = n7308 | n8208 ;
  assign n8210 = ( n4632 & n8208 ) | ( n4632 & n8209 ) | ( n8208 & n8209 ) ;
  assign n8211 = x11 & n8210 ;
  assign n8212 = x11 & ~n8211 ;
  assign n8213 = ( n8210 & ~n8211 ) | ( n8210 & n8212 ) | ( ~n8211 & n8212 ) ;
  assign n8214 = n8203 & n8213 ;
  assign n8215 = n8203 & ~n8214 ;
  assign n8216 = ~n8203 & n8213 ;
  assign n8217 = n8215 | n8216 ;
  assign n8218 = n8159 & ~n8163 ;
  assign n8219 = n8162 & ~n8163 ;
  assign n8220 = n8218 | n8219 ;
  assign n8221 = ~n1014 & n7305 ;
  assign n8222 = n3349 & n7300 ;
  assign n8223 = ~n3255 & n7302 ;
  assign n8224 = n8222 | n8223 ;
  assign n8225 = n8221 | n8224 ;
  assign n8226 = n7308 | n8225 ;
  assign n8227 = ( n4742 & n8225 ) | ( n4742 & n8226 ) | ( n8225 & n8226 ) ;
  assign n8228 = x11 & n8227 ;
  assign n8229 = x11 & ~n8228 ;
  assign n8230 = ( n8227 & ~n8228 ) | ( n8227 & n8229 ) | ( ~n8228 & n8229 ) ;
  assign n8231 = n8220 & n8230 ;
  assign n8232 = n8220 & ~n8231 ;
  assign n8233 = ~n8220 & n8230 ;
  assign n8234 = n8232 | n8233 ;
  assign n8235 = n8155 & ~n8158 ;
  assign n8236 = n8157 | n8158 ;
  assign n8237 = ~n8235 & n8236 ;
  assign n8238 = n1233 & n7300 ;
  assign n8239 = n3349 & n7302 ;
  assign n8240 = n8238 | n8239 ;
  assign n8241 = ~n3255 & n7305 ;
  assign n8242 = n8240 | n8241 ;
  assign n8243 = n7308 | n8242 ;
  assign n8244 = ( ~n4470 & n8242 ) | ( ~n4470 & n8243 ) | ( n8242 & n8243 ) ;
  assign n8245 = ~x11 & n8244 ;
  assign n8246 = x11 | n8245 ;
  assign n8247 = ( ~n8244 & n8245 ) | ( ~n8244 & n8246 ) | ( n8245 & n8246 ) ;
  assign n8248 = ~n8237 & n8247 ;
  assign n8249 = ~n1151 & n7300 ;
  assign n8250 = n1233 & n7302 ;
  assign n8251 = n8249 | n8250 ;
  assign n8252 = n3349 & n7305 ;
  assign n8253 = n8251 | n8252 ;
  assign n8254 = n7308 | n8253 ;
  assign n8255 = ( n4518 & n8253 ) | ( n4518 & n8254 ) | ( n8253 & n8254 ) ;
  assign n8256 = x11 & n8255 ;
  assign n8257 = x11 & ~n8256 ;
  assign n8258 = ( n8255 & ~n8256 ) | ( n8255 & n8257 ) | ( ~n8256 & n8257 ) ;
  assign n8259 = ( n7810 & n8154 ) | ( n7810 & ~n8155 ) | ( n8154 & ~n8155 ) ;
  assign n8260 = ( n7820 & ~n8155 ) | ( n7820 & n8259 ) | ( ~n8155 & n8259 ) ;
  assign n8261 = n8258 & n8260 ;
  assign n8262 = n8258 | n8260 ;
  assign n8263 = ~n8261 & n8262 ;
  assign n8264 = ( ~n7830 & n8153 ) | ( ~n7830 & n8154 ) | ( n8153 & n8154 ) ;
  assign n8265 = ( ~n8151 & n8154 ) | ( ~n8151 & n8264 ) | ( n8154 & n8264 ) ;
  assign n8266 = n1327 & n7300 ;
  assign n8267 = ~n1151 & n7302 ;
  assign n8268 = n8266 | n8267 ;
  assign n8269 = n1233 & n7305 ;
  assign n8270 = n8268 | n8269 ;
  assign n8271 = n7308 | n8270 ;
  assign n8272 = ( ~n4615 & n8270 ) | ( ~n4615 & n8271 ) | ( n8270 & n8271 ) ;
  assign n8273 = ~x11 & n8272 ;
  assign n8274 = x11 | n8273 ;
  assign n8275 = ( ~n8272 & n8273 ) | ( ~n8272 & n8274 ) | ( n8273 & n8274 ) ;
  assign n8276 = ~n8265 & n8275 ;
  assign n8277 = n8265 & ~n8275 ;
  assign n8278 = n8276 | n8277 ;
  assign n8279 = ( ~n7840 & n8150 ) | ( ~n7840 & n8151 ) | ( n8150 & n8151 ) ;
  assign n8280 = ( ~n8148 & n8151 ) | ( ~n8148 & n8279 ) | ( n8151 & n8279 ) ;
  assign n8281 = n3104 & n7300 ;
  assign n8282 = n1327 & n7302 ;
  assign n8283 = n8281 | n8282 ;
  assign n8284 = ~n1151 & n7305 ;
  assign n8285 = n8283 | n8284 ;
  assign n8286 = n7308 | n8285 ;
  assign n8287 = ( ~n4034 & n8285 ) | ( ~n4034 & n8286 ) | ( n8285 & n8286 ) ;
  assign n8288 = ~x11 & n8287 ;
  assign n8289 = x11 | n8288 ;
  assign n8290 = ( ~n8287 & n8288 ) | ( ~n8287 & n8289 ) | ( n8288 & n8289 ) ;
  assign n8291 = ~n8280 & n8290 ;
  assign n8292 = n8280 & ~n8290 ;
  assign n8293 = n8291 | n8292 ;
  assign n8294 = n3178 & n7300 ;
  assign n8295 = n3104 & n7302 ;
  assign n8296 = n8294 | n8295 ;
  assign n8297 = n1327 & n7305 ;
  assign n8298 = n8296 | n8297 ;
  assign n8299 = n7308 | n8298 ;
  assign n8300 = ( n4501 & n8298 ) | ( n4501 & n8299 ) | ( n8298 & n8299 ) ;
  assign n8301 = x11 & n8300 ;
  assign n8302 = x11 & ~n8301 ;
  assign n8303 = ( n8300 & ~n8301 ) | ( n8300 & n8302 ) | ( ~n8301 & n8302 ) ;
  assign n8304 = ( n7842 & n8147 ) | ( n7842 & ~n8148 ) | ( n8147 & ~n8148 ) ;
  assign n8305 = ( n7852 & ~n8148 ) | ( n7852 & n8304 ) | ( ~n8148 & n8304 ) ;
  assign n8306 = n8303 & n8305 ;
  assign n8307 = n8303 | n8305 ;
  assign n8308 = ~n8306 & n8307 ;
  assign n8309 = n8143 | n8145 ;
  assign n8310 = ~n8146 & n8309 ;
  assign n8311 = ~n1411 & n7300 ;
  assign n8312 = n3178 & n7302 ;
  assign n8313 = n8311 | n8312 ;
  assign n8314 = n3104 & n7305 ;
  assign n8315 = n8313 | n8314 ;
  assign n8316 = n7308 | n8315 ;
  assign n8317 = ( n4449 & n8315 ) | ( n4449 & n8316 ) | ( n8315 & n8316 ) ;
  assign n8318 = x11 & n8317 ;
  assign n8319 = x11 & ~n8318 ;
  assign n8320 = ( n8317 & ~n8318 ) | ( n8317 & n8319 ) | ( ~n8318 & n8319 ) ;
  assign n8321 = n8310 & n8320 ;
  assign n8322 = n8310 | n8320 ;
  assign n8323 = ~n8321 & n8322 ;
  assign n8324 = n7883 | n8141 ;
  assign n8325 = ~n8142 & n8324 ;
  assign n8326 = ~n1411 & n7302 ;
  assign n8327 = n7300 | n8326 ;
  assign n8328 = ( n1532 & n8326 ) | ( n1532 & n8327 ) | ( n8326 & n8327 ) ;
  assign n8329 = n3178 & n7305 ;
  assign n8330 = n8328 | n8329 ;
  assign n8331 = n7308 | n8330 ;
  assign n8332 = ( ~n3750 & n8330 ) | ( ~n3750 & n8331 ) | ( n8330 & n8331 ) ;
  assign n8333 = ~x11 & n8332 ;
  assign n8334 = x11 | n8333 ;
  assign n8335 = ( ~n8332 & n8333 ) | ( ~n8332 & n8334 ) | ( n8333 & n8334 ) ;
  assign n8336 = n7909 | n8139 ;
  assign n8337 = n8137 | n8336 ;
  assign n8338 = ~n8140 & n8337 ;
  assign n8339 = n1532 & n7302 ;
  assign n8340 = ~n1411 & n7305 ;
  assign n8341 = ~n2939 & n7300 ;
  assign n8342 = n8340 | n8341 ;
  assign n8343 = n8339 | n8342 ;
  assign n8344 = n7308 | n8343 ;
  assign n8345 = ( ~n3930 & n8343 ) | ( ~n3930 & n8344 ) | ( n8343 & n8344 ) ;
  assign n8346 = ~x11 & n8345 ;
  assign n8347 = x11 | n8346 ;
  assign n8348 = ( ~n8345 & n8346 ) | ( ~n8345 & n8347 ) | ( n8346 & n8347 ) ;
  assign n8349 = n8338 & n8348 ;
  assign n8350 = n8133 & ~n8137 ;
  assign n8351 = n8136 & ~n8137 ;
  assign n8352 = n8350 | n8351 ;
  assign n8353 = n1532 & n7305 ;
  assign n8354 = n3030 & n7300 ;
  assign n8355 = ~n2939 & n7302 ;
  assign n8356 = n8354 | n8355 ;
  assign n8357 = n8353 | n8356 ;
  assign n8358 = n7308 | n8357 ;
  assign n8359 = ( ~n4193 & n8357 ) | ( ~n4193 & n8358 ) | ( n8357 & n8358 ) ;
  assign n8360 = ~x11 & n8359 ;
  assign n8361 = x11 | n8360 ;
  assign n8362 = ( ~n8359 & n8360 ) | ( ~n8359 & n8361 ) | ( n8360 & n8361 ) ;
  assign n8363 = n8352 & n8362 ;
  assign n8364 = n8352 & ~n8363 ;
  assign n8365 = ~n8352 & n8362 ;
  assign n8366 = n8364 | n8365 ;
  assign n8367 = n8128 & ~n8132 ;
  assign n8368 = n8131 & ~n8132 ;
  assign n8369 = n8367 | n8368 ;
  assign n8370 = n1625 & n7300 ;
  assign n8371 = n3030 & n7302 ;
  assign n8372 = n8370 | n8371 ;
  assign n8373 = ~n2939 & n7305 ;
  assign n8374 = n8372 | n8373 ;
  assign n8375 = n7308 | n8374 ;
  assign n8376 = ( ~n4215 & n8374 ) | ( ~n4215 & n8375 ) | ( n8374 & n8375 ) ;
  assign n8377 = ~x11 & n8376 ;
  assign n8378 = x11 | n8377 ;
  assign n8379 = ( ~n8376 & n8377 ) | ( ~n8376 & n8378 ) | ( n8377 & n8378 ) ;
  assign n8380 = n8369 & n8379 ;
  assign n8381 = n8369 & ~n8380 ;
  assign n8382 = ~n8369 & n8379 ;
  assign n8383 = n8381 | n8382 ;
  assign n8384 = n7937 | n8126 ;
  assign n8385 = ~n8127 & n8384 ;
  assign n8386 = ~n1733 & n7300 ;
  assign n8387 = n1625 & n7302 ;
  assign n8388 = n8386 | n8387 ;
  assign n8389 = n3030 & n7305 ;
  assign n8390 = n8388 | n8389 ;
  assign n8391 = n7308 | n8390 ;
  assign n8392 = ( ~n4578 & n8390 ) | ( ~n4578 & n8391 ) | ( n8390 & n8391 ) ;
  assign n8393 = ~x11 & n8392 ;
  assign n8394 = x11 | n8393 ;
  assign n8395 = ( ~n8392 & n8393 ) | ( ~n8392 & n8394 ) | ( n8393 & n8394 ) ;
  assign n8396 = n8385 & n8395 ;
  assign n8397 = n7953 | n8124 ;
  assign n8398 = ~n8125 & n8397 ;
  assign n8399 = ~n2873 & n7300 ;
  assign n8400 = ~n1733 & n7302 ;
  assign n8401 = n8399 | n8400 ;
  assign n8402 = n1625 & n7305 ;
  assign n8403 = n8401 | n8402 ;
  assign n8404 = n7308 | n8403 ;
  assign n8405 = ( n4260 & n8403 ) | ( n4260 & n8404 ) | ( n8403 & n8404 ) ;
  assign n8406 = x11 & n8405 ;
  assign n8407 = x11 & ~n8406 ;
  assign n8408 = ( n8405 & ~n8406 ) | ( n8405 & n8407 ) | ( ~n8406 & n8407 ) ;
  assign n8409 = n8398 & n8408 ;
  assign n8410 = n7968 | n8122 ;
  assign n8411 = ~n8123 & n8410 ;
  assign n8412 = n1803 & n7300 ;
  assign n8413 = ~n2873 & n7302 ;
  assign n8414 = n8412 | n8413 ;
  assign n8415 = ~n1733 & n7305 ;
  assign n8416 = n8414 | n8415 ;
  assign n8417 = n7308 | n8416 ;
  assign n8418 = ( ~n4985 & n8416 ) | ( ~n4985 & n8417 ) | ( n8416 & n8417 ) ;
  assign n8419 = ~x11 & n8418 ;
  assign n8420 = x11 | n8419 ;
  assign n8421 = ( ~n8418 & n8419 ) | ( ~n8418 & n8420 ) | ( n8419 & n8420 ) ;
  assign n8422 = n8411 & n8421 ;
  assign n8423 = n8118 | n8120 ;
  assign n8424 = ~n8121 & n8423 ;
  assign n8425 = ~n2873 & n7305 ;
  assign n8426 = n1803 & n7302 ;
  assign n8427 = n8425 | n8426 ;
  assign n8428 = ~n1880 & n7300 ;
  assign n8429 = n8427 | n8428 ;
  assign n8430 = n7308 | n8429 ;
  assign n8431 = ( n5139 & n8429 ) | ( n5139 & n8430 ) | ( n8429 & n8430 ) ;
  assign n8432 = x11 & n8431 ;
  assign n8433 = x11 & ~n8432 ;
  assign n8434 = ( n8431 & ~n8432 ) | ( n8431 & n8433 ) | ( ~n8432 & n8433 ) ;
  assign n8435 = n8424 & n8434 ;
  assign n8436 = n8434 & ~n8435 ;
  assign n8437 = ( n8424 & ~n8435 ) | ( n8424 & n8436 ) | ( ~n8435 & n8436 ) ;
  assign n8438 = n1803 & n7305 ;
  assign n8439 = ~n1944 & n7300 ;
  assign n8440 = n8438 | n8439 ;
  assign n8441 = ~n1880 & n7302 ;
  assign n8442 = n8440 | n8441 ;
  assign n8443 = n7308 | n8442 ;
  assign n8444 = ( n4905 & n8442 ) | ( n4905 & n8443 ) | ( n8442 & n8443 ) ;
  assign n8445 = x11 & n8444 ;
  assign n8446 = x11 & ~n8445 ;
  assign n8447 = ( n8444 & ~n8445 ) | ( n8444 & n8446 ) | ( ~n8445 & n8446 ) ;
  assign n8448 = n7997 & ~n8117 ;
  assign n8449 = ( n8116 & ~n8117 ) | ( n8116 & n8448 ) | ( ~n8117 & n8448 ) ;
  assign n8450 = n8447 & n8449 ;
  assign n8451 = n8449 & ~n8450 ;
  assign n8452 = n8447 & ~n8449 ;
  assign n8453 = n8451 | n8452 ;
  assign n8454 = ~n2103 & n7300 ;
  assign n8455 = ~n1944 & n7302 ;
  assign n8456 = n8454 | n8455 ;
  assign n8457 = ~n1880 & n7305 ;
  assign n8458 = n8456 | n8457 ;
  assign n8459 = n7308 | n8458 ;
  assign n8460 = ( ~n5281 & n8458 ) | ( ~n5281 & n8459 ) | ( n8458 & n8459 ) ;
  assign n8461 = ~x11 & n8460 ;
  assign n8462 = x11 | n8461 ;
  assign n8463 = ( ~n8460 & n8461 ) | ( ~n8460 & n8462 ) | ( n8461 & n8462 ) ;
  assign n8464 = ( n7999 & n8115 ) | ( n7999 & ~n8116 ) | ( n8115 & ~n8116 ) ;
  assign n8465 = ( n8009 & ~n8116 ) | ( n8009 & n8464 ) | ( ~n8116 & n8464 ) ;
  assign n8466 = n8463 & n8465 ;
  assign n8467 = n8463 | n8465 ;
  assign n8468 = ~n8466 & n8467 ;
  assign n8469 = n8111 | n8113 ;
  assign n8470 = ~n8114 & n8469 ;
  assign n8471 = n2013 & n7300 ;
  assign n8472 = ~n2103 & n7302 ;
  assign n8473 = n8471 | n8472 ;
  assign n8474 = ~n1944 & n7305 ;
  assign n8475 = n8473 | n8474 ;
  assign n8476 = n7308 | n8475 ;
  assign n8477 = ( n6041 & n8475 ) | ( n6041 & n8476 ) | ( n8475 & n8476 ) ;
  assign n8478 = x11 & n8477 ;
  assign n8479 = x11 & ~n8478 ;
  assign n8480 = ( n8477 & ~n8478 ) | ( n8477 & n8479 ) | ( ~n8478 & n8479 ) ;
  assign n8481 = n8470 & n8480 ;
  assign n8482 = n8107 | n8109 ;
  assign n8483 = ~n8110 & n8482 ;
  assign n8484 = n2193 & n7300 ;
  assign n8485 = n2013 & n7302 ;
  assign n8486 = n8484 | n8485 ;
  assign n8487 = ~n2103 & n7305 ;
  assign n8488 = n8486 | n8487 ;
  assign n8489 = n7308 | n8488 ;
  assign n8490 = ( ~n5836 & n8488 ) | ( ~n5836 & n8489 ) | ( n8488 & n8489 ) ;
  assign n8491 = ~x11 & n8490 ;
  assign n8492 = x11 | n8491 ;
  assign n8493 = ( ~n8490 & n8491 ) | ( ~n8490 & n8492 ) | ( n8491 & n8492 ) ;
  assign n8494 = n8483 & n8493 ;
  assign n8495 = n8483 & ~n8494 ;
  assign n8496 = ~n8483 & n8493 ;
  assign n8497 = n8495 | n8496 ;
  assign n8498 = n8050 | n8105 ;
  assign n8499 = ~n8106 & n8498 ;
  assign n8500 = n2296 & n7300 ;
  assign n8501 = n2193 & n7302 ;
  assign n8502 = n8500 | n8501 ;
  assign n8503 = n2013 & n7305 ;
  assign n8504 = n8502 | n8503 ;
  assign n8505 = n7308 | n8504 ;
  assign n8506 = ( n5216 & n8504 ) | ( n5216 & n8505 ) | ( n8504 & n8505 ) ;
  assign n8507 = x11 & n8506 ;
  assign n8508 = x11 & ~n8507 ;
  assign n8509 = ( n8506 & ~n8507 ) | ( n8506 & n8508 ) | ( ~n8507 & n8508 ) ;
  assign n8510 = n8101 | n8103 ;
  assign n8511 = ~n8104 & n8510 ;
  assign n8512 = ~n2375 & n7300 ;
  assign n8513 = n2296 & n7302 ;
  assign n8514 = n8512 | n8513 ;
  assign n8515 = n2193 & n7305 ;
  assign n8516 = n8514 | n8515 ;
  assign n8517 = n7308 | n8516 ;
  assign n8518 = ( ~n5879 & n8516 ) | ( ~n5879 & n8517 ) | ( n8516 & n8517 ) ;
  assign n8519 = ~x11 & n8518 ;
  assign n8520 = x11 | n8519 ;
  assign n8521 = ( ~n8518 & n8519 ) | ( ~n8518 & n8520 ) | ( n8519 & n8520 ) ;
  assign n8522 = n8511 & n8521 ;
  assign n8523 = n8089 | n8099 ;
  assign n8524 = ~n8100 & n8523 ;
  assign n8525 = ~n2455 & n7300 ;
  assign n8526 = ~n2375 & n7302 ;
  assign n8527 = n8525 | n8526 ;
  assign n8528 = n2296 & n7305 ;
  assign n8529 = n8527 | n8528 ;
  assign n8530 = n7308 | n8529 ;
  assign n8531 = ( n5781 & n8529 ) | ( n5781 & n8530 ) | ( n8529 & n8530 ) ;
  assign n8532 = x11 & n8531 ;
  assign n8533 = x11 & ~n8532 ;
  assign n8534 = ( n8531 & ~n8532 ) | ( n8531 & n8533 ) | ( ~n8532 & n8533 ) ;
  assign n8535 = n8524 & n8534 ;
  assign n8536 = ~n2606 & n7300 ;
  assign n8537 = ~n2455 & n7302 ;
  assign n8538 = n8536 | n8537 ;
  assign n8539 = ~n2375 & n7305 ;
  assign n8540 = n8538 | n8539 ;
  assign n8541 = n7308 | n8540 ;
  assign n8542 = ( ~n5528 & n8540 ) | ( ~n5528 & n8541 ) | ( n8540 & n8541 ) ;
  assign n8543 = ~x11 & n8542 ;
  assign n8544 = x11 & ~n8542 ;
  assign n8545 = n8543 | n8544 ;
  assign n8546 = n8075 | n8084 ;
  assign n8547 = ~n8085 & n8546 ;
  assign n8548 = n8545 & n8547 ;
  assign n8549 = n8545 | n8547 ;
  assign n8550 = ~n8548 & n8549 ;
  assign n8551 = x14 & ~n8080 ;
  assign n8552 = n8082 | n8551 ;
  assign n8553 = n8083 | n8552 ;
  assign n8554 = ~n8084 & n8553 ;
  assign n8555 = ~n2455 & n7305 ;
  assign n8556 = ~n2606 & n7302 ;
  assign n8557 = n8555 | n8556 ;
  assign n8558 = n2569 & n7300 ;
  assign n8559 = n8557 | n8558 ;
  assign n8560 = n7308 | n8559 ;
  assign n8561 = ( ~n5732 & n8559 ) | ( ~n5732 & n8560 ) | ( n8559 & n8560 ) ;
  assign n8562 = ~x11 & n8561 ;
  assign n8563 = x11 | n8562 ;
  assign n8564 = ( ~n8561 & n8562 ) | ( ~n8561 & n8563 ) | ( n8562 & n8563 ) ;
  assign n8565 = n8554 & n8564 ;
  assign n8566 = ~n2764 & n7300 ;
  assign n8567 = ~n2672 & n7302 ;
  assign n8568 = n8566 | n8567 ;
  assign n8569 = n2569 & n7305 ;
  assign n8570 = n8568 | n8569 ;
  assign n8571 = ( n5584 & n7308 ) | ( n5584 & n8570 ) | ( n7308 & n8570 ) ;
  assign n8572 = ( x11 & ~n8570 ) | ( x11 & n8571 ) | ( ~n8570 & n8571 ) ;
  assign n8573 = ~n8571 & n8572 ;
  assign n8574 = n8570 | n8572 ;
  assign n8575 = ( ~x11 & n8573 ) | ( ~x11 & n8574 ) | ( n8573 & n8574 ) ;
  assign n8576 = ~n2764 & n7302 ;
  assign n8577 = ~n2672 & n7305 ;
  assign n8578 = n8576 | n8577 ;
  assign n8579 = n7308 | n8578 ;
  assign n8580 = ( n5932 & n8578 ) | ( n5932 & n8579 ) | ( n8578 & n8579 ) ;
  assign n8581 = ~n2764 & n7298 ;
  assign n8582 = x11 & ~n8581 ;
  assign n8583 = ~x11 & n8580 ;
  assign n8584 = ( ~n8580 & n8582 ) | ( ~n8580 & n8583 ) | ( n8582 & n8583 ) ;
  assign n8585 = n8575 & n8584 ;
  assign n8586 = n8081 & n8585 ;
  assign n8587 = n8585 & ~n8586 ;
  assign n8588 = n8081 & ~n8585 ;
  assign n8589 = n8587 | n8588 ;
  assign n8590 = ~n2606 & n7305 ;
  assign n8591 = ~n2672 & n7300 ;
  assign n8592 = n8590 | n8591 ;
  assign n8593 = n2569 & n7302 ;
  assign n8594 = n8592 | n8593 ;
  assign n8595 = n7308 | n8594 ;
  assign n8596 = ( n5716 & n8594 ) | ( n5716 & n8595 ) | ( n8594 & n8595 ) ;
  assign n8597 = x11 & n8596 ;
  assign n8598 = x11 & ~n8597 ;
  assign n8599 = ( n8596 & ~n8597 ) | ( n8596 & n8598 ) | ( ~n8597 & n8598 ) ;
  assign n8600 = n8589 & n8599 ;
  assign n8601 = n8586 | n8600 ;
  assign n8602 = n8554 | n8564 ;
  assign n8603 = ~n8565 & n8602 ;
  assign n8604 = n8601 & n8603 ;
  assign n8605 = n8565 | n8604 ;
  assign n8606 = n8550 & n8605 ;
  assign n8607 = n8548 | n8606 ;
  assign n8608 = n8524 | n8534 ;
  assign n8609 = ~n8535 & n8608 ;
  assign n8610 = n8607 & n8609 ;
  assign n8611 = n8535 | n8610 ;
  assign n8612 = n8521 & ~n8522 ;
  assign n8613 = ( n8511 & ~n8522 ) | ( n8511 & n8612 ) | ( ~n8522 & n8612 ) ;
  assign n8614 = n8611 & n8613 ;
  assign n8615 = n8522 | n8614 ;
  assign n8616 = ( n8499 & n8509 ) | ( n8499 & n8615 ) | ( n8509 & n8615 ) ;
  assign n8617 = n8497 & n8616 ;
  assign n8618 = n8494 | n8617 ;
  assign n8619 = n8470 | n8480 ;
  assign n8620 = ~n8481 & n8619 ;
  assign n8621 = n8618 & n8620 ;
  assign n8622 = n8481 | n8621 ;
  assign n8623 = n8468 & n8622 ;
  assign n8624 = n8466 | n8623 ;
  assign n8625 = n8453 & n8624 ;
  assign n8626 = n8450 | n8625 ;
  assign n8627 = n8437 & n8626 ;
  assign n8628 = n8435 | n8627 ;
  assign n8629 = n8411 & ~n8422 ;
  assign n8630 = ~n8411 & n8421 ;
  assign n8631 = n8629 | n8630 ;
  assign n8632 = n8628 & n8631 ;
  assign n8633 = n8422 | n8632 ;
  assign n8634 = n8398 & ~n8409 ;
  assign n8635 = ~n8398 & n8408 ;
  assign n8636 = n8634 | n8635 ;
  assign n8637 = n8633 & n8636 ;
  assign n8638 = n8385 | n8395 ;
  assign n8639 = ~n8396 & n8638 ;
  assign n8640 = ( n8409 & n8637 ) | ( n8409 & n8639 ) | ( n8637 & n8639 ) ;
  assign n8641 = n8396 | n8640 ;
  assign n8642 = n8383 & n8641 ;
  assign n8643 = n8380 | n8642 ;
  assign n8644 = n8366 & n8643 ;
  assign n8645 = n8363 | n8644 ;
  assign n8646 = n8348 & ~n8349 ;
  assign n8647 = ( n8338 & ~n8349 ) | ( n8338 & n8646 ) | ( ~n8349 & n8646 ) ;
  assign n8648 = n8645 & n8647 ;
  assign n8649 = n8349 | n8648 ;
  assign n8650 = ( n8325 & n8335 ) | ( n8325 & n8649 ) | ( n8335 & n8649 ) ;
  assign n8651 = n8323 & n8650 ;
  assign n8652 = n8321 | n8651 ;
  assign n8653 = n8308 & n8652 ;
  assign n8654 = n8306 | n8653 ;
  assign n8655 = ~n8293 & n8654 ;
  assign n8656 = n8291 | n8655 ;
  assign n8657 = ~n8278 & n8656 ;
  assign n8658 = n8276 | n8657 ;
  assign n8659 = n8263 & n8658 ;
  assign n8660 = n8261 | n8659 ;
  assign n8661 = n8237 | n8248 ;
  assign n8662 = ( ~n8247 & n8248 ) | ( ~n8247 & n8661 ) | ( n8248 & n8661 ) ;
  assign n8663 = n8660 & ~n8662 ;
  assign n8664 = n8248 | n8663 ;
  assign n8665 = n8234 & n8664 ;
  assign n8666 = n8231 | n8665 ;
  assign n8667 = n8217 & n8666 ;
  assign n8668 = n8214 | n8667 ;
  assign n8669 = n8200 & n8668 ;
  assign n8670 = ~x3 & x4 ;
  assign n8671 = x3 & ~x4 ;
  assign n8672 = n8670 | n8671 ;
  assign n8673 = x4 & ~x5 ;
  assign n8674 = ~x4 & x5 ;
  assign n8675 = n8673 | n8674 ;
  assign n8676 = x2 & ~x3 ;
  assign n8677 = ~x2 & x3 ;
  assign n8678 = n8676 | n8677 ;
  assign n8679 = n8675 & ~n8678 ;
  assign n8680 = ~n8672 & n8679 ;
  assign n8681 = n8672 & ~n8678 ;
  assign n8682 = ~n3634 & n8681 ;
  assign n8683 = n672 & n8680 ;
  assign n8684 = ( n8680 & n8682 ) | ( n8680 & ~n8683 ) | ( n8682 & ~n8683 ) ;
  assign n8685 = n8675 & n8678 ;
  assign n8686 = n8684 | n8685 ;
  assign n8687 = ( n3726 & n8684 ) | ( n3726 & n8686 ) | ( n8684 & n8686 ) ;
  assign n8688 = x5 & n8687 ;
  assign n8689 = x5 & ~n8688 ;
  assign n8690 = ( n8687 & ~n8688 ) | ( n8687 & n8689 ) | ( ~n8688 & n8689 ) ;
  assign n8691 = n8669 | n8690 ;
  assign n8692 = n8668 & ~n8669 ;
  assign n8693 = n8200 & ~n8668 ;
  assign n8694 = ~n3596 & n5512 ;
  assign n8695 = n3504 & n5508 ;
  assign n8696 = n8694 | n8695 ;
  assign n8697 = ~n3431 & n5503 ;
  assign n8698 = n8696 | n8697 ;
  assign n8699 = n5515 | n8698 ;
  assign n8700 = ( ~n4798 & n8698 ) | ( ~n4798 & n8699 ) | ( n8698 & n8699 ) ;
  assign n8701 = ~x8 & n8700 ;
  assign n8702 = x8 | n8701 ;
  assign n8703 = ( ~n8700 & n8701 ) | ( ~n8700 & n8702 ) | ( n8701 & n8702 ) ;
  assign n8704 = ( n8692 & n8693 ) | ( n8692 & n8703 ) | ( n8693 & n8703 ) ;
  assign n8705 = n8691 | n8704 ;
  assign n8706 = ( n8669 & n8690 ) | ( n8669 & n8704 ) | ( n8690 & n8704 ) ;
  assign n8707 = n8705 & ~n8706 ;
  assign n8708 = n3504 & n5512 ;
  assign n8709 = ~n3431 & n5508 ;
  assign n8710 = n8708 | n8709 ;
  assign n8711 = ~n589 & n5503 ;
  assign n8712 = n8710 | n8711 ;
  assign n8713 = n5515 | n8712 ;
  assign n8714 = ( n4765 & n8712 ) | ( n4765 & n8713 ) | ( n8712 & n8713 ) ;
  assign n8715 = x8 & n8714 ;
  assign n8716 = x8 & ~n8715 ;
  assign n8717 = ( n8714 & ~n8715 ) | ( n8714 & n8716 ) | ( ~n8715 & n8716 ) ;
  assign n8718 = n8186 | n8198 ;
  assign n8719 = ( ~n7289 & n7313 ) | ( ~n7289 & n7414 ) | ( n7313 & n7414 ) ;
  assign n8720 = ( n7289 & ~n7414 ) | ( n7289 & n8719 ) | ( ~n7414 & n8719 ) ;
  assign n8721 = ( ~n7313 & n8719 ) | ( ~n7313 & n8720 ) | ( n8719 & n8720 ) ;
  assign n8722 = ( n8717 & ~n8718 ) | ( n8717 & n8721 ) | ( ~n8718 & n8721 ) ;
  assign n8723 = ( n8718 & ~n8721 ) | ( n8718 & n8722 ) | ( ~n8721 & n8722 ) ;
  assign n8724 = ( ~n8717 & n8722 ) | ( ~n8717 & n8723 ) | ( n8722 & n8723 ) ;
  assign n8725 = n8707 & n8724 ;
  assign n8726 = n8707 | n8724 ;
  assign n8727 = ~n8725 & n8726 ;
  assign n8728 = n8217 | n8666 ;
  assign n8729 = ~n8667 & n8728 ;
  assign n8730 = n778 & n5512 ;
  assign n8731 = ~n3596 & n5508 ;
  assign n8732 = n8730 | n8731 ;
  assign n8733 = n3504 & n5503 ;
  assign n8734 = n8732 | n8733 ;
  assign n8735 = n5515 | n8734 ;
  assign n8736 = ( ~n5040 & n8734 ) | ( ~n5040 & n8735 ) | ( n8734 & n8735 ) ;
  assign n8737 = ~x8 & n8736 ;
  assign n8738 = x8 | n8737 ;
  assign n8739 = ( ~n8736 & n8737 ) | ( ~n8736 & n8738 ) | ( n8737 & n8738 ) ;
  assign n8740 = n8729 & n8739 ;
  assign n8741 = n8234 | n8664 ;
  assign n8742 = ~n8665 & n8741 ;
  assign n8743 = n904 & n5512 ;
  assign n8744 = n778 & n5508 ;
  assign n8745 = n8743 | n8744 ;
  assign n8746 = ~n3596 & n5503 ;
  assign n8747 = n8745 | n8746 ;
  assign n8748 = ( ~n4649 & n5515 ) | ( ~n4649 & n8747 ) | ( n5515 & n8747 ) ;
  assign n8749 = n8747 | n8748 ;
  assign n8750 = ~x8 & n8749 ;
  assign n8751 = x8 | n8750 ;
  assign n8752 = ( ~n8749 & n8750 ) | ( ~n8749 & n8751 ) | ( n8750 & n8751 ) ;
  assign n8753 = n8742 & n8752 ;
  assign n8754 = ~n8660 & n8662 ;
  assign n8755 = n8663 | n8754 ;
  assign n8756 = ~n1014 & n5512 ;
  assign n8757 = n904 & n5508 ;
  assign n8758 = n8756 | n8757 ;
  assign n8759 = n778 & n5503 ;
  assign n8760 = n8758 | n8759 ;
  assign n8761 = n5515 | n8760 ;
  assign n8762 = ( ~n4535 & n8760 ) | ( ~n4535 & n8761 ) | ( n8760 & n8761 ) ;
  assign n8763 = ~x8 & n8762 ;
  assign n8764 = x8 | n8763 ;
  assign n8765 = ( ~n8762 & n8763 ) | ( ~n8762 & n8764 ) | ( n8763 & n8764 ) ;
  assign n8766 = ~n8755 & n8765 ;
  assign n8767 = n8263 | n8658 ;
  assign n8768 = ~n8659 & n8767 ;
  assign n8769 = ~n1014 & n5508 ;
  assign n8770 = ~n3255 & n5512 ;
  assign n8771 = n8769 | n8770 ;
  assign n8772 = n904 & n5503 ;
  assign n8773 = n8771 | n8772 ;
  assign n8774 = n5515 | n8773 ;
  assign n8775 = ( n4632 & n8773 ) | ( n4632 & n8774 ) | ( n8773 & n8774 ) ;
  assign n8776 = x8 & n8775 ;
  assign n8777 = x8 & ~n8776 ;
  assign n8778 = ( n8775 & ~n8776 ) | ( n8775 & n8777 ) | ( ~n8776 & n8777 ) ;
  assign n8779 = n8768 & n8778 ;
  assign n8780 = n8278 & ~n8656 ;
  assign n8781 = n8657 | n8780 ;
  assign n8782 = ~n1014 & n5503 ;
  assign n8783 = n3349 & n5512 ;
  assign n8784 = ~n3255 & n5508 ;
  assign n8785 = n8783 | n8784 ;
  assign n8786 = n8782 | n8785 ;
  assign n8787 = n5515 | n8786 ;
  assign n8788 = ( n4742 & n8786 ) | ( n4742 & n8787 ) | ( n8786 & n8787 ) ;
  assign n8789 = x8 & n8788 ;
  assign n8790 = x8 & ~n8789 ;
  assign n8791 = ( n8788 & ~n8789 ) | ( n8788 & n8790 ) | ( ~n8789 & n8790 ) ;
  assign n8792 = ~n8781 & n8791 ;
  assign n8793 = n8293 & ~n8654 ;
  assign n8794 = n8655 | n8793 ;
  assign n8795 = n1233 & n5512 ;
  assign n8796 = n3349 & n5508 ;
  assign n8797 = n8795 | n8796 ;
  assign n8798 = ~n3255 & n5503 ;
  assign n8799 = n8797 | n8798 ;
  assign n8800 = n5515 | n8799 ;
  assign n8801 = ( ~n4470 & n8799 ) | ( ~n4470 & n8800 ) | ( n8799 & n8800 ) ;
  assign n8802 = ~x8 & n8801 ;
  assign n8803 = x8 | n8802 ;
  assign n8804 = ( ~n8801 & n8802 ) | ( ~n8801 & n8803 ) | ( n8802 & n8803 ) ;
  assign n8805 = ~n8794 & n8804 ;
  assign n8806 = n8308 | n8652 ;
  assign n8807 = ~n8653 & n8806 ;
  assign n8808 = ~n1151 & n5512 ;
  assign n8809 = n1233 & n5508 ;
  assign n8810 = n8808 | n8809 ;
  assign n8811 = n3349 & n5503 ;
  assign n8812 = n8810 | n8811 ;
  assign n8813 = n5515 | n8812 ;
  assign n8814 = ( n4518 & n8812 ) | ( n4518 & n8813 ) | ( n8812 & n8813 ) ;
  assign n8815 = x8 & n8814 ;
  assign n8816 = x8 & ~n8815 ;
  assign n8817 = ( n8814 & ~n8815 ) | ( n8814 & n8816 ) | ( ~n8815 & n8816 ) ;
  assign n8818 = n8807 & n8817 ;
  assign n8819 = n8323 | n8650 ;
  assign n8820 = ~n8651 & n8819 ;
  assign n8821 = n1327 & n5512 ;
  assign n8822 = ~n1151 & n5508 ;
  assign n8823 = n8821 | n8822 ;
  assign n8824 = n1233 & n5503 ;
  assign n8825 = n8823 | n8824 ;
  assign n8826 = n5515 | n8825 ;
  assign n8827 = ( ~n4615 & n8825 ) | ( ~n4615 & n8826 ) | ( n8825 & n8826 ) ;
  assign n8828 = ~x8 & n8827 ;
  assign n8829 = x8 | n8828 ;
  assign n8830 = ( ~n8827 & n8828 ) | ( ~n8827 & n8829 ) | ( n8828 & n8829 ) ;
  assign n8831 = n8820 & n8830 ;
  assign n8832 = n8830 & ~n8831 ;
  assign n8833 = ( n8820 & ~n8831 ) | ( n8820 & n8832 ) | ( ~n8831 & n8832 ) ;
  assign n8834 = n3104 & n5512 ;
  assign n8835 = n1327 & n5508 ;
  assign n8836 = n8834 | n8835 ;
  assign n8837 = ~n1151 & n5503 ;
  assign n8838 = n8836 | n8837 ;
  assign n8839 = n5515 | n8838 ;
  assign n8840 = ( ~n4034 & n8838 ) | ( ~n4034 & n8839 ) | ( n8838 & n8839 ) ;
  assign n8841 = ~x8 & n8840 ;
  assign n8842 = x8 | n8841 ;
  assign n8843 = ( ~n8840 & n8841 ) | ( ~n8840 & n8842 ) | ( n8841 & n8842 ) ;
  assign n8844 = ( n8325 & n8649 ) | ( n8325 & ~n8650 ) | ( n8649 & ~n8650 ) ;
  assign n8845 = ( n8335 & ~n8650 ) | ( n8335 & n8844 ) | ( ~n8650 & n8844 ) ;
  assign n8846 = n8843 & n8845 ;
  assign n8847 = n8843 | n8845 ;
  assign n8848 = ~n8846 & n8847 ;
  assign n8849 = n8645 | n8647 ;
  assign n8850 = ~n8648 & n8849 ;
  assign n8851 = n3178 & n5512 ;
  assign n8852 = n3104 & n5508 ;
  assign n8853 = n8851 | n8852 ;
  assign n8854 = n1327 & n5503 ;
  assign n8855 = n8853 | n8854 ;
  assign n8856 = n5515 | n8855 ;
  assign n8857 = ( n4501 & n8855 ) | ( n4501 & n8856 ) | ( n8855 & n8856 ) ;
  assign n8858 = x8 & n8857 ;
  assign n8859 = x8 & ~n8858 ;
  assign n8860 = ( n8857 & ~n8858 ) | ( n8857 & n8859 ) | ( ~n8858 & n8859 ) ;
  assign n8861 = n8850 & n8860 ;
  assign n8862 = n8850 | n8860 ;
  assign n8863 = ~n8861 & n8862 ;
  assign n8864 = n8366 | n8643 ;
  assign n8865 = ~n8644 & n8864 ;
  assign n8866 = ~n1411 & n5512 ;
  assign n8867 = n3178 & n5508 ;
  assign n8868 = n8866 | n8867 ;
  assign n8869 = n3104 & n5503 ;
  assign n8870 = n8868 | n8869 ;
  assign n8871 = n5515 | n8870 ;
  assign n8872 = ( n4449 & n8870 ) | ( n4449 & n8871 ) | ( n8870 & n8871 ) ;
  assign n8873 = x8 & n8872 ;
  assign n8874 = x8 & ~n8873 ;
  assign n8875 = ( n8872 & ~n8873 ) | ( n8872 & n8874 ) | ( ~n8873 & n8874 ) ;
  assign n8876 = n8383 | n8641 ;
  assign n8877 = ~n8642 & n8876 ;
  assign n8878 = ~n1411 & n5508 ;
  assign n8879 = n5512 | n8878 ;
  assign n8880 = ( n1532 & n8878 ) | ( n1532 & n8879 ) | ( n8878 & n8879 ) ;
  assign n8881 = n3178 & n5503 ;
  assign n8882 = n8880 | n8881 ;
  assign n8883 = n5515 | n8882 ;
  assign n8884 = ( ~n3750 & n8882 ) | ( ~n3750 & n8883 ) | ( n8882 & n8883 ) ;
  assign n8885 = ~x8 & n8884 ;
  assign n8886 = x8 | n8885 ;
  assign n8887 = ( ~n8884 & n8885 ) | ( ~n8884 & n8886 ) | ( n8885 & n8886 ) ;
  assign n8888 = n8409 | n8639 ;
  assign n8889 = n8637 | n8888 ;
  assign n8890 = ~n8640 & n8889 ;
  assign n8891 = n1532 & n5508 ;
  assign n8892 = ~n1411 & n5503 ;
  assign n8893 = ~n2939 & n5512 ;
  assign n8894 = n8892 | n8893 ;
  assign n8895 = n8891 | n8894 ;
  assign n8896 = n5515 | n8895 ;
  assign n8897 = ( ~n3930 & n8895 ) | ( ~n3930 & n8896 ) | ( n8895 & n8896 ) ;
  assign n8898 = ~x8 & n8897 ;
  assign n8899 = x8 | n8898 ;
  assign n8900 = ( ~n8897 & n8898 ) | ( ~n8897 & n8899 ) | ( n8898 & n8899 ) ;
  assign n8901 = n8890 & n8900 ;
  assign n8902 = n8633 & ~n8637 ;
  assign n8903 = n8636 & ~n8637 ;
  assign n8904 = n8902 | n8903 ;
  assign n8905 = n1532 & n5503 ;
  assign n8906 = n3030 & n5512 ;
  assign n8907 = ~n2939 & n5508 ;
  assign n8908 = n8906 | n8907 ;
  assign n8909 = n8905 | n8908 ;
  assign n8910 = n5515 | n8909 ;
  assign n8911 = ( ~n4193 & n8909 ) | ( ~n4193 & n8910 ) | ( n8909 & n8910 ) ;
  assign n8912 = ~x8 & n8911 ;
  assign n8913 = x8 | n8912 ;
  assign n8914 = ( ~n8911 & n8912 ) | ( ~n8911 & n8913 ) | ( n8912 & n8913 ) ;
  assign n8915 = n8904 & n8914 ;
  assign n8916 = n8904 & ~n8915 ;
  assign n8917 = ~n8904 & n8914 ;
  assign n8918 = n8916 | n8917 ;
  assign n8919 = n8628 & ~n8632 ;
  assign n8920 = n8631 & ~n8632 ;
  assign n8921 = n8919 | n8920 ;
  assign n8922 = n1625 & n5512 ;
  assign n8923 = n3030 & n5508 ;
  assign n8924 = n8922 | n8923 ;
  assign n8925 = ~n2939 & n5503 ;
  assign n8926 = n8924 | n8925 ;
  assign n8927 = n5515 | n8926 ;
  assign n8928 = ( ~n4215 & n8926 ) | ( ~n4215 & n8927 ) | ( n8926 & n8927 ) ;
  assign n8929 = ~x8 & n8928 ;
  assign n8930 = x8 | n8929 ;
  assign n8931 = ( ~n8928 & n8929 ) | ( ~n8928 & n8930 ) | ( n8929 & n8930 ) ;
  assign n8932 = n8921 & n8931 ;
  assign n8933 = n8921 & ~n8932 ;
  assign n8934 = ~n8921 & n8931 ;
  assign n8935 = n8933 | n8934 ;
  assign n8936 = n8437 | n8626 ;
  assign n8937 = ~n8627 & n8936 ;
  assign n8938 = ~n1733 & n5512 ;
  assign n8939 = n1625 & n5508 ;
  assign n8940 = n8938 | n8939 ;
  assign n8941 = n3030 & n5503 ;
  assign n8942 = n8940 | n8941 ;
  assign n8943 = n5515 | n8942 ;
  assign n8944 = ( ~n4578 & n8942 ) | ( ~n4578 & n8943 ) | ( n8942 & n8943 ) ;
  assign n8945 = ~x8 & n8944 ;
  assign n8946 = x8 | n8945 ;
  assign n8947 = ( ~n8944 & n8945 ) | ( ~n8944 & n8946 ) | ( n8945 & n8946 ) ;
  assign n8948 = n8937 & n8947 ;
  assign n8949 = n8453 | n8624 ;
  assign n8950 = ~n8625 & n8949 ;
  assign n8951 = ~n2873 & n5512 ;
  assign n8952 = ~n1733 & n5508 ;
  assign n8953 = n8951 | n8952 ;
  assign n8954 = n1625 & n5503 ;
  assign n8955 = n8953 | n8954 ;
  assign n8956 = n5515 | n8955 ;
  assign n8957 = ( n4260 & n8955 ) | ( n4260 & n8956 ) | ( n8955 & n8956 ) ;
  assign n8958 = x8 & n8957 ;
  assign n8959 = x8 & ~n8958 ;
  assign n8960 = ( n8957 & ~n8958 ) | ( n8957 & n8959 ) | ( ~n8958 & n8959 ) ;
  assign n8961 = n8950 & n8960 ;
  assign n8962 = n8468 | n8622 ;
  assign n8963 = ~n8623 & n8962 ;
  assign n8964 = n1803 & n5512 ;
  assign n8965 = ~n2873 & n5508 ;
  assign n8966 = n8964 | n8965 ;
  assign n8967 = ~n1733 & n5503 ;
  assign n8968 = n8966 | n8967 ;
  assign n8969 = n5515 | n8968 ;
  assign n8970 = ( ~n4985 & n8968 ) | ( ~n4985 & n8969 ) | ( n8968 & n8969 ) ;
  assign n8971 = ~x8 & n8970 ;
  assign n8972 = x8 | n8971 ;
  assign n8973 = ( ~n8970 & n8971 ) | ( ~n8970 & n8972 ) | ( n8971 & n8972 ) ;
  assign n8974 = n8963 & n8973 ;
  assign n8975 = n8618 | n8620 ;
  assign n8976 = ~n8621 & n8975 ;
  assign n8977 = ~n2873 & n5503 ;
  assign n8978 = n1803 & n5508 ;
  assign n8979 = n8977 | n8978 ;
  assign n8980 = ~n1880 & n5512 ;
  assign n8981 = n8979 | n8980 ;
  assign n8982 = n5515 | n8981 ;
  assign n8983 = ( n5139 & n8981 ) | ( n5139 & n8982 ) | ( n8981 & n8982 ) ;
  assign n8984 = x8 & n8983 ;
  assign n8985 = x8 & ~n8984 ;
  assign n8986 = ( n8983 & ~n8984 ) | ( n8983 & n8985 ) | ( ~n8984 & n8985 ) ;
  assign n8987 = n8976 & n8986 ;
  assign n8988 = n8986 & ~n8987 ;
  assign n8989 = ( n8976 & ~n8987 ) | ( n8976 & n8988 ) | ( ~n8987 & n8988 ) ;
  assign n8990 = n1803 & n5503 ;
  assign n8991 = ~n1944 & n5512 ;
  assign n8992 = n8990 | n8991 ;
  assign n8993 = ~n1880 & n5508 ;
  assign n8994 = n8992 | n8993 ;
  assign n8995 = n5515 | n8994 ;
  assign n8996 = ( n4905 & n8994 ) | ( n4905 & n8995 ) | ( n8994 & n8995 ) ;
  assign n8997 = x8 & n8996 ;
  assign n8998 = x8 & ~n8997 ;
  assign n8999 = ( n8996 & ~n8997 ) | ( n8996 & n8998 ) | ( ~n8997 & n8998 ) ;
  assign n9000 = n8497 & ~n8617 ;
  assign n9001 = ( n8616 & ~n8617 ) | ( n8616 & n9000 ) | ( ~n8617 & n9000 ) ;
  assign n9002 = n8999 & n9001 ;
  assign n9003 = n9001 & ~n9002 ;
  assign n9004 = n8999 & ~n9001 ;
  assign n9005 = n9003 | n9004 ;
  assign n9006 = ~n2103 & n5512 ;
  assign n9007 = ~n1944 & n5508 ;
  assign n9008 = n9006 | n9007 ;
  assign n9009 = ~n1880 & n5503 ;
  assign n9010 = n9008 | n9009 ;
  assign n9011 = n5515 | n9010 ;
  assign n9012 = ( ~n5281 & n9010 ) | ( ~n5281 & n9011 ) | ( n9010 & n9011 ) ;
  assign n9013 = ~x8 & n9012 ;
  assign n9014 = x8 | n9013 ;
  assign n9015 = ( ~n9012 & n9013 ) | ( ~n9012 & n9014 ) | ( n9013 & n9014 ) ;
  assign n9016 = ( n8499 & n8615 ) | ( n8499 & ~n8616 ) | ( n8615 & ~n8616 ) ;
  assign n9017 = ( n8509 & ~n8616 ) | ( n8509 & n9016 ) | ( ~n8616 & n9016 ) ;
  assign n9018 = n9015 & n9017 ;
  assign n9019 = n9015 | n9017 ;
  assign n9020 = ~n9018 & n9019 ;
  assign n9021 = n8611 | n8613 ;
  assign n9022 = ~n8614 & n9021 ;
  assign n9023 = n2013 & n5512 ;
  assign n9024 = ~n2103 & n5508 ;
  assign n9025 = n9023 | n9024 ;
  assign n9026 = ~n1944 & n5503 ;
  assign n9027 = n9025 | n9026 ;
  assign n9028 = n5515 | n9027 ;
  assign n9029 = ( n6041 & n9027 ) | ( n6041 & n9028 ) | ( n9027 & n9028 ) ;
  assign n9030 = x8 & n9029 ;
  assign n9031 = x8 & ~n9030 ;
  assign n9032 = ( n9029 & ~n9030 ) | ( n9029 & n9031 ) | ( ~n9030 & n9031 ) ;
  assign n9033 = n9022 & n9032 ;
  assign n9034 = n8607 | n8609 ;
  assign n9035 = ~n8610 & n9034 ;
  assign n9036 = n2193 & n5512 ;
  assign n9037 = n2013 & n5508 ;
  assign n9038 = n9036 | n9037 ;
  assign n9039 = ~n2103 & n5503 ;
  assign n9040 = n9038 | n9039 ;
  assign n9041 = n5515 | n9040 ;
  assign n9042 = ( ~n5836 & n9040 ) | ( ~n5836 & n9041 ) | ( n9040 & n9041 ) ;
  assign n9043 = ~x8 & n9042 ;
  assign n9044 = x8 | n9043 ;
  assign n9045 = ( ~n9042 & n9043 ) | ( ~n9042 & n9044 ) | ( n9043 & n9044 ) ;
  assign n9046 = n9035 & n9045 ;
  assign n9047 = n9035 & ~n9046 ;
  assign n9048 = ~n9035 & n9045 ;
  assign n9049 = n9047 | n9048 ;
  assign n9050 = n8550 | n8605 ;
  assign n9051 = ~n8606 & n9050 ;
  assign n9052 = n2296 & n5512 ;
  assign n9053 = n2193 & n5508 ;
  assign n9054 = n9052 | n9053 ;
  assign n9055 = n2013 & n5503 ;
  assign n9056 = n9054 | n9055 ;
  assign n9057 = n5515 | n9056 ;
  assign n9058 = ( n5216 & n9056 ) | ( n5216 & n9057 ) | ( n9056 & n9057 ) ;
  assign n9059 = x8 & n9058 ;
  assign n9060 = x8 & ~n9059 ;
  assign n9061 = ( n9058 & ~n9059 ) | ( n9058 & n9060 ) | ( ~n9059 & n9060 ) ;
  assign n9062 = n8601 | n8603 ;
  assign n9063 = ~n8604 & n9062 ;
  assign n9064 = ~n2375 & n5512 ;
  assign n9065 = n2296 & n5508 ;
  assign n9066 = n9064 | n9065 ;
  assign n9067 = n2193 & n5503 ;
  assign n9068 = n9066 | n9067 ;
  assign n9069 = n5515 | n9068 ;
  assign n9070 = ( ~n5879 & n9068 ) | ( ~n5879 & n9069 ) | ( n9068 & n9069 ) ;
  assign n9071 = ~x8 & n9070 ;
  assign n9072 = x8 | n9071 ;
  assign n9073 = ( ~n9070 & n9071 ) | ( ~n9070 & n9072 ) | ( n9071 & n9072 ) ;
  assign n9074 = n9063 & n9073 ;
  assign n9075 = n8589 | n8599 ;
  assign n9076 = ~n8600 & n9075 ;
  assign n9077 = ~n2455 & n5512 ;
  assign n9078 = ~n2375 & n5508 ;
  assign n9079 = n9077 | n9078 ;
  assign n9080 = n2296 & n5503 ;
  assign n9081 = n9079 | n9080 ;
  assign n9082 = n5515 | n9081 ;
  assign n9083 = ( n5781 & n9081 ) | ( n5781 & n9082 ) | ( n9081 & n9082 ) ;
  assign n9084 = x8 & n9083 ;
  assign n9085 = x8 & ~n9084 ;
  assign n9086 = ( n9083 & ~n9084 ) | ( n9083 & n9085 ) | ( ~n9084 & n9085 ) ;
  assign n9087 = n9076 & n9086 ;
  assign n9088 = ~n2606 & n5512 ;
  assign n9089 = ~n2455 & n5508 ;
  assign n9090 = n9088 | n9089 ;
  assign n9091 = ~n2375 & n5503 ;
  assign n9092 = n9090 | n9091 ;
  assign n9093 = n5515 | n9092 ;
  assign n9094 = ( ~n5528 & n9092 ) | ( ~n5528 & n9093 ) | ( n9092 & n9093 ) ;
  assign n9095 = ~x8 & n9094 ;
  assign n9096 = x8 & ~n9094 ;
  assign n9097 = n9095 | n9096 ;
  assign n9098 = n8575 | n8584 ;
  assign n9099 = ~n8585 & n9098 ;
  assign n9100 = n9097 & n9099 ;
  assign n9101 = n9097 | n9099 ;
  assign n9102 = ~n9100 & n9101 ;
  assign n9103 = x11 & ~n8580 ;
  assign n9104 = n8582 | n9103 ;
  assign n9105 = n8583 | n9104 ;
  assign n9106 = ~n8584 & n9105 ;
  assign n9107 = ~n2455 & n5503 ;
  assign n9108 = ~n2606 & n5508 ;
  assign n9109 = n9107 | n9108 ;
  assign n9110 = n2569 & n5512 ;
  assign n9111 = n9109 | n9110 ;
  assign n9112 = n5515 | n9111 ;
  assign n9113 = ( ~n5732 & n9111 ) | ( ~n5732 & n9112 ) | ( n9111 & n9112 ) ;
  assign n9114 = ~x8 & n9113 ;
  assign n9115 = x8 | n9114 ;
  assign n9116 = ( ~n9113 & n9114 ) | ( ~n9113 & n9115 ) | ( n9114 & n9115 ) ;
  assign n9117 = n9106 & n9116 ;
  assign n9118 = ~n2764 & n5512 ;
  assign n9119 = ~n2672 & n5508 ;
  assign n9120 = n9118 | n9119 ;
  assign n9121 = n2569 & n5503 ;
  assign n9122 = n9120 | n9121 ;
  assign n9123 = ( n5515 & n5584 ) | ( n5515 & n9122 ) | ( n5584 & n9122 ) ;
  assign n9124 = ( x8 & ~n9122 ) | ( x8 & n9123 ) | ( ~n9122 & n9123 ) ;
  assign n9125 = ~n9123 & n9124 ;
  assign n9126 = n9122 | n9124 ;
  assign n9127 = ( ~x8 & n9125 ) | ( ~x8 & n9126 ) | ( n9125 & n9126 ) ;
  assign n9128 = ~n2764 & n5508 ;
  assign n9129 = ~n2672 & n5503 ;
  assign n9130 = n9128 | n9129 ;
  assign n9131 = n5515 | n9130 ;
  assign n9132 = ( n5932 & n9130 ) | ( n5932 & n9131 ) | ( n9130 & n9131 ) ;
  assign n9133 = ~n2764 & n5502 ;
  assign n9134 = x8 & ~n9133 ;
  assign n9135 = ~x8 & n9132 ;
  assign n9136 = ( ~n9132 & n9134 ) | ( ~n9132 & n9135 ) | ( n9134 & n9135 ) ;
  assign n9137 = n9127 & n9136 ;
  assign n9138 = n8581 & n9137 ;
  assign n9139 = n9137 & ~n9138 ;
  assign n9140 = n8581 & ~n9137 ;
  assign n9141 = n9139 | n9140 ;
  assign n9142 = ~n2606 & n5503 ;
  assign n9143 = ~n2672 & n5512 ;
  assign n9144 = n9142 | n9143 ;
  assign n9145 = n2569 & n5508 ;
  assign n9146 = n9144 | n9145 ;
  assign n9147 = n5515 | n9146 ;
  assign n9148 = ( n5716 & n9146 ) | ( n5716 & n9147 ) | ( n9146 & n9147 ) ;
  assign n9149 = x8 & n9148 ;
  assign n9150 = x8 & ~n9149 ;
  assign n9151 = ( n9148 & ~n9149 ) | ( n9148 & n9150 ) | ( ~n9149 & n9150 ) ;
  assign n9152 = n9141 & n9151 ;
  assign n9153 = n9138 | n9152 ;
  assign n9154 = n9106 | n9116 ;
  assign n9155 = ~n9117 & n9154 ;
  assign n9156 = n9153 & n9155 ;
  assign n9157 = n9117 | n9156 ;
  assign n9158 = n9102 & n9157 ;
  assign n9159 = n9100 | n9158 ;
  assign n9160 = n9076 | n9086 ;
  assign n9161 = ~n9087 & n9160 ;
  assign n9162 = n9159 & n9161 ;
  assign n9163 = n9087 | n9162 ;
  assign n9164 = n9073 & ~n9074 ;
  assign n9165 = ( n9063 & ~n9074 ) | ( n9063 & n9164 ) | ( ~n9074 & n9164 ) ;
  assign n9166 = n9163 & n9165 ;
  assign n9167 = n9074 | n9166 ;
  assign n9168 = ( n9051 & n9061 ) | ( n9051 & n9167 ) | ( n9061 & n9167 ) ;
  assign n9169 = n9049 & n9168 ;
  assign n9170 = n9046 | n9169 ;
  assign n9171 = n9022 | n9032 ;
  assign n9172 = ~n9033 & n9171 ;
  assign n9173 = n9170 & n9172 ;
  assign n9174 = n9033 | n9173 ;
  assign n9175 = n9020 & n9174 ;
  assign n9176 = n9018 | n9175 ;
  assign n9177 = n9005 & n9176 ;
  assign n9178 = n9002 | n9177 ;
  assign n9179 = n8989 & n9178 ;
  assign n9180 = n8987 | n9179 ;
  assign n9181 = n8963 & ~n8974 ;
  assign n9182 = ~n8963 & n8973 ;
  assign n9183 = n9181 | n9182 ;
  assign n9184 = n9180 & n9183 ;
  assign n9185 = n8974 | n9184 ;
  assign n9186 = n8950 & ~n8961 ;
  assign n9187 = ~n8950 & n8960 ;
  assign n9188 = n9186 | n9187 ;
  assign n9189 = n9185 & n9188 ;
  assign n9190 = n8937 | n8947 ;
  assign n9191 = ~n8948 & n9190 ;
  assign n9192 = ( n8961 & n9189 ) | ( n8961 & n9191 ) | ( n9189 & n9191 ) ;
  assign n9193 = n8948 | n9192 ;
  assign n9194 = n8935 & n9193 ;
  assign n9195 = n8932 | n9194 ;
  assign n9196 = n8918 & n9195 ;
  assign n9197 = n8915 | n9196 ;
  assign n9198 = n8900 & ~n8901 ;
  assign n9199 = ( n8890 & ~n8901 ) | ( n8890 & n9198 ) | ( ~n8901 & n9198 ) ;
  assign n9200 = n9197 & n9199 ;
  assign n9201 = n8901 | n9200 ;
  assign n9202 = ( n8877 & n8887 ) | ( n8877 & n9201 ) | ( n8887 & n9201 ) ;
  assign n9203 = ( n8865 & n8875 ) | ( n8865 & n9202 ) | ( n8875 & n9202 ) ;
  assign n9204 = n8863 & n9203 ;
  assign n9205 = n8861 | n9204 ;
  assign n9206 = n8848 & n9205 ;
  assign n9207 = n8846 | n9206 ;
  assign n9208 = n8833 & n9207 ;
  assign n9209 = n8831 | n9208 ;
  assign n9210 = n8807 & ~n8818 ;
  assign n9211 = ~n8807 & n8817 ;
  assign n9212 = n9210 | n9211 ;
  assign n9213 = n9209 & n9212 ;
  assign n9214 = n8818 | n9213 ;
  assign n9215 = n8794 | n8805 ;
  assign n9216 = ( ~n8804 & n8805 ) | ( ~n8804 & n9215 ) | ( n8805 & n9215 ) ;
  assign n9217 = n9214 & ~n9216 ;
  assign n9218 = n8805 | n9217 ;
  assign n9219 = n8781 | n8792 ;
  assign n9220 = ( ~n8791 & n8792 ) | ( ~n8791 & n9219 ) | ( n8792 & n9219 ) ;
  assign n9221 = n9218 & ~n9220 ;
  assign n9222 = n8792 | n9221 ;
  assign n9223 = n8768 & ~n8779 ;
  assign n9224 = ~n8768 & n8778 ;
  assign n9225 = n9223 | n9224 ;
  assign n9226 = n9222 & n9225 ;
  assign n9227 = n8779 | n9226 ;
  assign n9228 = n8755 | n8766 ;
  assign n9229 = ( ~n8765 & n8766 ) | ( ~n8765 & n9228 ) | ( n8766 & n9228 ) ;
  assign n9230 = n9227 & ~n9229 ;
  assign n9231 = n8766 | n9230 ;
  assign n9232 = n8742 & ~n8753 ;
  assign n9233 = ~n8742 & n8752 ;
  assign n9234 = n9232 | n9233 ;
  assign n9235 = n9231 & n9234 ;
  assign n9236 = n8753 | n9235 ;
  assign n9237 = n8729 & ~n8740 ;
  assign n9238 = ~n8729 & n8739 ;
  assign n9239 = n9237 | n9238 ;
  assign n9240 = n9236 & n9239 ;
  assign n9241 = n8740 | n9240 ;
  assign n9242 = n8693 | n8703 ;
  assign n9243 = n8692 | n9242 ;
  assign n9244 = ~n8704 & n9243 ;
  assign n9245 = ~n8675 & n8678 ;
  assign n9246 = ~n3634 & n9245 ;
  assign n9247 = ~n672 & n8681 ;
  assign n9248 = n9246 | n9247 ;
  assign n9249 = ~n589 & n8680 ;
  assign n9250 = n9248 | n9249 ;
  assign n9251 = n8685 | n9250 ;
  assign n9252 = ( ~n5092 & n9250 ) | ( ~n5092 & n9251 ) | ( n9250 & n9251 ) ;
  assign n9253 = ~x5 & n9252 ;
  assign n9254 = x5 | n9253 ;
  assign n9255 = ( ~n9252 & n9253 ) | ( ~n9252 & n9254 ) | ( n9253 & n9254 ) ;
  assign n9256 = ( n9241 & n9244 ) | ( n9241 & n9255 ) | ( n9244 & n9255 ) ;
  assign n9257 = n8727 & n9256 ;
  assign n9258 = n8727 | n9256 ;
  assign n9259 = ~n9257 & n9258 ;
  assign n9260 = n9231 & ~n9235 ;
  assign n9261 = n9234 & ~n9235 ;
  assign n9262 = n9260 | n9261 ;
  assign n9263 = n3504 & n8680 ;
  assign n9264 = ~n3431 & n8681 ;
  assign n9265 = n9263 | n9264 ;
  assign n9266 = ~n589 & n9245 ;
  assign n9267 = n9265 | n9266 ;
  assign n9268 = n8685 | n9267 ;
  assign n9269 = ( n4765 & n9267 ) | ( n4765 & n9268 ) | ( n9267 & n9268 ) ;
  assign n9270 = x5 & n9269 ;
  assign n9271 = x5 & ~n9270 ;
  assign n9272 = ( n9269 & ~n9270 ) | ( n9269 & n9271 ) | ( ~n9270 & n9271 ) ;
  assign n9273 = n9262 & n9272 ;
  assign n9274 = n9262 & ~n9273 ;
  assign n9275 = ~n9262 & n9272 ;
  assign n9276 = n9274 | n9275 ;
  assign n9277 = n9227 & ~n9230 ;
  assign n9278 = n9229 | n9230 ;
  assign n9279 = ~n9277 & n9278 ;
  assign n9280 = ~n3596 & n8680 ;
  assign n9281 = n3504 & n8681 ;
  assign n9282 = n9280 | n9281 ;
  assign n9283 = ~n3431 & n9245 ;
  assign n9284 = n9282 | n9283 ;
  assign n9285 = n8685 | n9284 ;
  assign n9286 = ( ~n4798 & n9284 ) | ( ~n4798 & n9285 ) | ( n9284 & n9285 ) ;
  assign n9287 = ~x5 & n9286 ;
  assign n9288 = x5 | n9287 ;
  assign n9289 = ( ~n9286 & n9287 ) | ( ~n9286 & n9288 ) | ( n9287 & n9288 ) ;
  assign n9290 = ~n9279 & n9289 ;
  assign n9291 = n9222 & ~n9226 ;
  assign n9292 = n9225 & ~n9226 ;
  assign n9293 = n9291 | n9292 ;
  assign n9294 = n778 & n8680 ;
  assign n9295 = ~n3596 & n8681 ;
  assign n9296 = n9294 | n9295 ;
  assign n9297 = n3504 & n9245 ;
  assign n9298 = n9296 | n9297 ;
  assign n9299 = n8685 | n9298 ;
  assign n9300 = ( ~n5040 & n9298 ) | ( ~n5040 & n9299 ) | ( n9298 & n9299 ) ;
  assign n9301 = ~x5 & n9300 ;
  assign n9302 = x5 | n9301 ;
  assign n9303 = ( ~n9300 & n9301 ) | ( ~n9300 & n9302 ) | ( n9301 & n9302 ) ;
  assign n9304 = n9293 & n9303 ;
  assign n9305 = n9293 & ~n9304 ;
  assign n9306 = ~n9293 & n9303 ;
  assign n9307 = n9305 | n9306 ;
  assign n9308 = n9218 & ~n9221 ;
  assign n9309 = n9220 | n9221 ;
  assign n9310 = ~n9308 & n9309 ;
  assign n9311 = n904 & n8680 ;
  assign n9312 = n778 & n8681 ;
  assign n9313 = n9311 | n9312 ;
  assign n9314 = ~n3596 & n9245 ;
  assign n9315 = n9313 | n9314 ;
  assign n9316 = n8685 | n9315 ;
  assign n9317 = ( ~n4649 & n9315 ) | ( ~n4649 & n9316 ) | ( n9315 & n9316 ) ;
  assign n9318 = ~x5 & n9317 ;
  assign n9319 = x5 | n9318 ;
  assign n9320 = ( ~n9317 & n9318 ) | ( ~n9317 & n9319 ) | ( n9318 & n9319 ) ;
  assign n9321 = ~n9310 & n9320 ;
  assign n9322 = n9214 & ~n9217 ;
  assign n9323 = n9216 | n9217 ;
  assign n9324 = ~n9322 & n9323 ;
  assign n9325 = ~n1014 & n8680 ;
  assign n9326 = n904 & n8681 ;
  assign n9327 = n9325 | n9326 ;
  assign n9328 = n778 & n9245 ;
  assign n9329 = n9327 | n9328 ;
  assign n9330 = n8685 | n9329 ;
  assign n9331 = ( ~n4535 & n9329 ) | ( ~n4535 & n9330 ) | ( n9329 & n9330 ) ;
  assign n9332 = ~x5 & n9331 ;
  assign n9333 = x5 | n9332 ;
  assign n9334 = ( ~n9331 & n9332 ) | ( ~n9331 & n9333 ) | ( n9332 & n9333 ) ;
  assign n9335 = ~n9324 & n9334 ;
  assign n9336 = n9209 & ~n9213 ;
  assign n9337 = n9212 & ~n9213 ;
  assign n9338 = n9336 | n9337 ;
  assign n9339 = ~n1014 & n8681 ;
  assign n9340 = ~n3255 & n8680 ;
  assign n9341 = n9339 | n9340 ;
  assign n9342 = n904 & n9245 ;
  assign n9343 = n9341 | n9342 ;
  assign n9344 = n8685 | n9343 ;
  assign n9345 = ( n4632 & n9343 ) | ( n4632 & n9344 ) | ( n9343 & n9344 ) ;
  assign n9346 = x5 & n9345 ;
  assign n9347 = x5 & ~n9346 ;
  assign n9348 = ( n9345 & ~n9346 ) | ( n9345 & n9347 ) | ( ~n9346 & n9347 ) ;
  assign n9349 = n8833 | n9207 ;
  assign n9350 = ~n9208 & n9349 ;
  assign n9351 = ~n1014 & n9245 ;
  assign n9352 = n3349 & n8680 ;
  assign n9353 = ~n3255 & n8681 ;
  assign n9354 = n9352 | n9353 ;
  assign n9355 = n9351 | n9354 ;
  assign n9356 = n8685 | n9355 ;
  assign n9357 = ( n4742 & n9355 ) | ( n4742 & n9356 ) | ( n9355 & n9356 ) ;
  assign n9358 = x5 & n9357 ;
  assign n9359 = x5 & ~n9358 ;
  assign n9360 = ( n9357 & ~n9358 ) | ( n9357 & n9359 ) | ( ~n9358 & n9359 ) ;
  assign n9361 = n9350 & n9360 ;
  assign n9362 = n8848 | n9205 ;
  assign n9363 = ~n9206 & n9362 ;
  assign n9364 = n1233 & n8680 ;
  assign n9365 = n3349 & n8681 ;
  assign n9366 = n9364 | n9365 ;
  assign n9367 = ~n3255 & n9245 ;
  assign n9368 = n9366 | n9367 ;
  assign n9369 = n8685 | n9368 ;
  assign n9370 = ( ~n4470 & n9368 ) | ( ~n4470 & n9369 ) | ( n9368 & n9369 ) ;
  assign n9371 = ~x5 & n9370 ;
  assign n9372 = x5 | n9371 ;
  assign n9373 = ( ~n9370 & n9371 ) | ( ~n9370 & n9372 ) | ( n9371 & n9372 ) ;
  assign n9374 = n9363 & n9373 ;
  assign n9375 = n9350 | n9360 ;
  assign n9376 = ~n9361 & n9375 ;
  assign n9377 = n8863 | n9203 ;
  assign n9378 = ~n9204 & n9377 ;
  assign n9379 = ~n1151 & n8680 ;
  assign n9380 = n1233 & n8681 ;
  assign n9381 = n9379 | n9380 ;
  assign n9382 = n3349 & n9245 ;
  assign n9383 = n9381 | n9382 ;
  assign n9384 = n8685 | n9383 ;
  assign n9385 = ( n4518 & n9383 ) | ( n4518 & n9384 ) | ( n9383 & n9384 ) ;
  assign n9386 = x5 & n9385 ;
  assign n9387 = x5 & ~n9386 ;
  assign n9388 = ( n9385 & ~n9386 ) | ( n9385 & n9387 ) | ( ~n9386 & n9387 ) ;
  assign n9389 = n9378 & n9388 ;
  assign n9390 = n9388 & ~n9389 ;
  assign n9391 = ( n9378 & ~n9389 ) | ( n9378 & n9390 ) | ( ~n9389 & n9390 ) ;
  assign n9392 = n1327 & n8680 ;
  assign n9393 = ~n1151 & n8681 ;
  assign n9394 = n9392 | n9393 ;
  assign n9395 = n1233 & n9245 ;
  assign n9396 = n9394 | n9395 ;
  assign n9397 = n8685 | n9396 ;
  assign n9398 = ( ~n4615 & n9396 ) | ( ~n4615 & n9397 ) | ( n9396 & n9397 ) ;
  assign n9399 = ~x5 & n9398 ;
  assign n9400 = x5 | n9399 ;
  assign n9401 = ( ~n9398 & n9399 ) | ( ~n9398 & n9400 ) | ( n9399 & n9400 ) ;
  assign n9402 = n3104 & n8680 ;
  assign n9403 = n1327 & n8681 ;
  assign n9404 = n9402 | n9403 ;
  assign n9405 = ~n1151 & n9245 ;
  assign n9406 = n9404 | n9405 ;
  assign n9407 = n8685 | n9406 ;
  assign n9408 = ( ~n4034 & n9406 ) | ( ~n4034 & n9407 ) | ( n9406 & n9407 ) ;
  assign n9409 = ~x5 & n9408 ;
  assign n9410 = x5 | n9409 ;
  assign n9411 = ( ~n9408 & n9409 ) | ( ~n9408 & n9410 ) | ( n9409 & n9410 ) ;
  assign n9412 = n9197 | n9199 ;
  assign n9413 = ~n9200 & n9412 ;
  assign n9414 = n3178 & n8680 ;
  assign n9415 = n3104 & n8681 ;
  assign n9416 = n9414 | n9415 ;
  assign n9417 = n1327 & n9245 ;
  assign n9418 = n9416 | n9417 ;
  assign n9419 = n8685 | n9418 ;
  assign n9420 = ( n4501 & n9418 ) | ( n4501 & n9419 ) | ( n9418 & n9419 ) ;
  assign n9421 = x5 & n9420 ;
  assign n9422 = x5 & ~n9421 ;
  assign n9423 = ( n9420 & ~n9421 ) | ( n9420 & n9422 ) | ( ~n9421 & n9422 ) ;
  assign n9424 = n9413 & n9423 ;
  assign n9425 = n9413 | n9423 ;
  assign n9426 = ~n9424 & n9425 ;
  assign n9427 = n8918 | n9195 ;
  assign n9428 = ~n9196 & n9427 ;
  assign n9429 = ~n1411 & n8680 ;
  assign n9430 = n3178 & n8681 ;
  assign n9431 = n9429 | n9430 ;
  assign n9432 = n3104 & n9245 ;
  assign n9433 = n9431 | n9432 ;
  assign n9434 = n8685 | n9433 ;
  assign n9435 = ( n4449 & n9433 ) | ( n4449 & n9434 ) | ( n9433 & n9434 ) ;
  assign n9436 = x5 & n9435 ;
  assign n9437 = x5 & ~n9436 ;
  assign n9438 = ( n9435 & ~n9436 ) | ( n9435 & n9437 ) | ( ~n9436 & n9437 ) ;
  assign n9439 = n8935 | n9193 ;
  assign n9440 = ~n9194 & n9439 ;
  assign n9441 = ~n1411 & n8681 ;
  assign n9442 = n8680 | n9441 ;
  assign n9443 = ( n1532 & n9441 ) | ( n1532 & n9442 ) | ( n9441 & n9442 ) ;
  assign n9444 = n3178 & n9245 ;
  assign n9445 = n9443 | n9444 ;
  assign n9446 = n8685 | n9445 ;
  assign n9447 = ( ~n3750 & n9445 ) | ( ~n3750 & n9446 ) | ( n9445 & n9446 ) ;
  assign n9448 = ~x5 & n9447 ;
  assign n9449 = x5 | n9448 ;
  assign n9450 = ( ~n9447 & n9448 ) | ( ~n9447 & n9449 ) | ( n9448 & n9449 ) ;
  assign n9451 = n8961 | n9191 ;
  assign n9452 = n9189 | n9451 ;
  assign n9453 = ~n9192 & n9452 ;
  assign n9454 = n1532 & n8681 ;
  assign n9455 = ~n1411 & n9245 ;
  assign n9456 = ~n2939 & n8680 ;
  assign n9457 = n9455 | n9456 ;
  assign n9458 = n9454 | n9457 ;
  assign n9459 = n8685 | n9458 ;
  assign n9460 = ( ~n3930 & n9458 ) | ( ~n3930 & n9459 ) | ( n9458 & n9459 ) ;
  assign n9461 = ~x5 & n9460 ;
  assign n9462 = x5 | n9461 ;
  assign n9463 = ( ~n9460 & n9461 ) | ( ~n9460 & n9462 ) | ( n9461 & n9462 ) ;
  assign n9464 = n9185 & ~n9189 ;
  assign n9465 = n9188 & ~n9189 ;
  assign n9466 = n9464 | n9465 ;
  assign n9467 = n1532 & n9245 ;
  assign n9468 = n3030 & n8680 ;
  assign n9469 = ~n2939 & n8681 ;
  assign n9470 = n9468 | n9469 ;
  assign n9471 = n9467 | n9470 ;
  assign n9472 = n8685 | n9471 ;
  assign n9473 = ( ~n4193 & n9471 ) | ( ~n4193 & n9472 ) | ( n9471 & n9472 ) ;
  assign n9474 = ~x5 & n9473 ;
  assign n9475 = x5 | n9474 ;
  assign n9476 = ( ~n9473 & n9474 ) | ( ~n9473 & n9475 ) | ( n9474 & n9475 ) ;
  assign n9477 = n9180 & ~n9184 ;
  assign n9478 = n9183 & ~n9184 ;
  assign n9479 = n9477 | n9478 ;
  assign n9480 = n1625 & n8680 ;
  assign n9481 = n3030 & n8681 ;
  assign n9482 = n9480 | n9481 ;
  assign n9483 = ~n2939 & n9245 ;
  assign n9484 = n9482 | n9483 ;
  assign n9485 = n8685 | n9484 ;
  assign n9486 = ( ~n4215 & n9484 ) | ( ~n4215 & n9485 ) | ( n9484 & n9485 ) ;
  assign n9487 = ~x5 & n9486 ;
  assign n9488 = x5 | n9487 ;
  assign n9489 = ( ~n9486 & n9487 ) | ( ~n9486 & n9488 ) | ( n9487 & n9488 ) ;
  assign n9490 = n8989 | n9178 ;
  assign n9491 = ~n9179 & n9490 ;
  assign n9492 = ~n1733 & n8680 ;
  assign n9493 = n1625 & n8681 ;
  assign n9494 = n9492 | n9493 ;
  assign n9495 = n3030 & n9245 ;
  assign n9496 = n9494 | n9495 ;
  assign n9497 = n8685 | n9496 ;
  assign n9498 = ( ~n4578 & n9496 ) | ( ~n4578 & n9497 ) | ( n9496 & n9497 ) ;
  assign n9499 = ~x5 & n9498 ;
  assign n9500 = x5 | n9499 ;
  assign n9501 = ( ~n9498 & n9499 ) | ( ~n9498 & n9500 ) | ( n9499 & n9500 ) ;
  assign n9502 = n9491 & n9501 ;
  assign n9503 = n9005 | n9176 ;
  assign n9504 = ~n9177 & n9503 ;
  assign n9505 = ~n2873 & n8680 ;
  assign n9506 = ~n1733 & n8681 ;
  assign n9507 = n9505 | n9506 ;
  assign n9508 = n1625 & n9245 ;
  assign n9509 = n9507 | n9508 ;
  assign n9510 = n8685 | n9509 ;
  assign n9511 = ( n4260 & n9509 ) | ( n4260 & n9510 ) | ( n9509 & n9510 ) ;
  assign n9512 = x5 & n9511 ;
  assign n9513 = x5 & ~n9512 ;
  assign n9514 = ( n9511 & ~n9512 ) | ( n9511 & n9513 ) | ( ~n9512 & n9513 ) ;
  assign n9515 = n9504 & n9514 ;
  assign n9516 = n9491 | n9501 ;
  assign n9517 = ~n9502 & n9516 ;
  assign n9518 = n9020 | n9174 ;
  assign n9519 = ~n9175 & n9518 ;
  assign n9520 = n1803 & n8680 ;
  assign n9521 = ~n2873 & n8681 ;
  assign n9522 = n9520 | n9521 ;
  assign n9523 = ~n1733 & n9245 ;
  assign n9524 = n9522 | n9523 ;
  assign n9525 = n8685 | n9524 ;
  assign n9526 = ( ~n4985 & n9524 ) | ( ~n4985 & n9525 ) | ( n9524 & n9525 ) ;
  assign n9527 = ~x5 & n9526 ;
  assign n9528 = x5 | n9527 ;
  assign n9529 = ( ~n9526 & n9527 ) | ( ~n9526 & n9528 ) | ( n9527 & n9528 ) ;
  assign n9530 = n9519 & n9529 ;
  assign n9531 = n9170 | n9172 ;
  assign n9532 = ~n9173 & n9531 ;
  assign n9533 = ~n2873 & n9245 ;
  assign n9534 = n1803 & n8681 ;
  assign n9535 = n9533 | n9534 ;
  assign n9536 = ~n1880 & n8680 ;
  assign n9537 = n9535 | n9536 ;
  assign n9538 = n8685 | n9537 ;
  assign n9539 = ( n5139 & n9537 ) | ( n5139 & n9538 ) | ( n9537 & n9538 ) ;
  assign n9540 = x5 & n9539 ;
  assign n9541 = x5 & ~n9540 ;
  assign n9542 = ( n9539 & ~n9540 ) | ( n9539 & n9541 ) | ( ~n9540 & n9541 ) ;
  assign n9543 = n9532 & n9542 ;
  assign n9544 = n9542 & ~n9543 ;
  assign n9545 = ( n9532 & ~n9543 ) | ( n9532 & n9544 ) | ( ~n9543 & n9544 ) ;
  assign n9546 = n1803 & n9245 ;
  assign n9547 = ~n1944 & n8680 ;
  assign n9548 = n9546 | n9547 ;
  assign n9549 = ~n1880 & n8681 ;
  assign n9550 = n9548 | n9549 ;
  assign n9551 = n8685 | n9550 ;
  assign n9552 = ( n4905 & n9550 ) | ( n4905 & n9551 ) | ( n9550 & n9551 ) ;
  assign n9553 = x5 & n9552 ;
  assign n9554 = x5 & ~n9553 ;
  assign n9555 = ( n9552 & ~n9553 ) | ( n9552 & n9554 ) | ( ~n9553 & n9554 ) ;
  assign n9556 = ~n2103 & n8680 ;
  assign n9557 = ~n1944 & n8681 ;
  assign n9558 = n9556 | n9557 ;
  assign n9559 = ~n1880 & n9245 ;
  assign n9560 = n9558 | n9559 ;
  assign n9561 = n8685 | n9560 ;
  assign n9562 = ( ~n5281 & n9560 ) | ( ~n5281 & n9561 ) | ( n9560 & n9561 ) ;
  assign n9563 = ~x5 & n9562 ;
  assign n9564 = x5 | n9563 ;
  assign n9565 = ( ~n9562 & n9563 ) | ( ~n9562 & n9564 ) | ( n9563 & n9564 ) ;
  assign n9566 = n9163 | n9165 ;
  assign n9567 = ~n9166 & n9566 ;
  assign n9568 = n2013 & n8680 ;
  assign n9569 = ~n2103 & n8681 ;
  assign n9570 = n9568 | n9569 ;
  assign n9571 = ~n1944 & n9245 ;
  assign n9572 = n9570 | n9571 ;
  assign n9573 = n8685 | n9572 ;
  assign n9574 = ( n6041 & n9572 ) | ( n6041 & n9573 ) | ( n9572 & n9573 ) ;
  assign n9575 = x5 & n9574 ;
  assign n9576 = x5 & ~n9575 ;
  assign n9577 = ( n9574 & ~n9575 ) | ( n9574 & n9576 ) | ( ~n9575 & n9576 ) ;
  assign n9578 = n9567 & n9577 ;
  assign n9579 = n9159 | n9161 ;
  assign n9580 = ~n9162 & n9579 ;
  assign n9581 = n2193 & n8680 ;
  assign n9582 = n2013 & n8681 ;
  assign n9583 = n9581 | n9582 ;
  assign n9584 = ~n2103 & n9245 ;
  assign n9585 = n9583 | n9584 ;
  assign n9586 = n8685 | n9585 ;
  assign n9587 = ( ~n5836 & n9585 ) | ( ~n5836 & n9586 ) | ( n9585 & n9586 ) ;
  assign n9588 = ~x5 & n9587 ;
  assign n9589 = x5 | n9588 ;
  assign n9590 = ( ~n9587 & n9588 ) | ( ~n9587 & n9589 ) | ( n9588 & n9589 ) ;
  assign n9591 = n9580 & n9590 ;
  assign n9592 = n9580 & ~n9591 ;
  assign n9593 = ~n9580 & n9590 ;
  assign n9594 = n9592 | n9593 ;
  assign n9595 = n9102 | n9157 ;
  assign n9596 = ~n9158 & n9595 ;
  assign n9597 = n2296 & n8680 ;
  assign n9598 = n2193 & n8681 ;
  assign n9599 = n9597 | n9598 ;
  assign n9600 = n2013 & n9245 ;
  assign n9601 = n9599 | n9600 ;
  assign n9602 = n8685 | n9601 ;
  assign n9603 = ( n5216 & n9601 ) | ( n5216 & n9602 ) | ( n9601 & n9602 ) ;
  assign n9604 = x5 & n9603 ;
  assign n9605 = x5 & ~n9604 ;
  assign n9606 = ( n9603 & ~n9604 ) | ( n9603 & n9605 ) | ( ~n9604 & n9605 ) ;
  assign n9607 = n9596 & n9606 ;
  assign n9608 = n9153 | n9155 ;
  assign n9609 = ~n9156 & n9608 ;
  assign n9610 = ~n2375 & n8680 ;
  assign n9611 = n2296 & n8681 ;
  assign n9612 = n9610 | n9611 ;
  assign n9613 = n2193 & n9245 ;
  assign n9614 = n9612 | n9613 ;
  assign n9615 = n8685 | n9614 ;
  assign n9616 = ( ~n5879 & n9614 ) | ( ~n5879 & n9615 ) | ( n9614 & n9615 ) ;
  assign n9617 = ~x5 & n9616 ;
  assign n9618 = x5 | n9617 ;
  assign n9619 = ( ~n9616 & n9617 ) | ( ~n9616 & n9618 ) | ( n9617 & n9618 ) ;
  assign n9620 = n9609 & n9619 ;
  assign n9621 = n9141 | n9151 ;
  assign n9622 = ~n9152 & n9621 ;
  assign n9623 = ~n2455 & n8680 ;
  assign n9624 = ~n2375 & n8681 ;
  assign n9625 = n9623 | n9624 ;
  assign n9626 = n2296 & n9245 ;
  assign n9627 = n9625 | n9626 ;
  assign n9628 = n8685 | n9627 ;
  assign n9629 = ( n5781 & n9627 ) | ( n5781 & n9628 ) | ( n9627 & n9628 ) ;
  assign n9630 = x5 & n9629 ;
  assign n9631 = x5 & ~n9630 ;
  assign n9632 = ( n9629 & ~n9630 ) | ( n9629 & n9631 ) | ( ~n9630 & n9631 ) ;
  assign n9633 = n9622 & n9632 ;
  assign n9634 = ~n2606 & n8680 ;
  assign n9635 = ~n2455 & n8681 ;
  assign n9636 = n9634 | n9635 ;
  assign n9637 = ~n2375 & n9245 ;
  assign n9638 = n9636 | n9637 ;
  assign n9639 = n8685 | n9638 ;
  assign n9640 = ( ~n5528 & n9638 ) | ( ~n5528 & n9639 ) | ( n9638 & n9639 ) ;
  assign n9641 = ~x5 & n9640 ;
  assign n9642 = x5 & ~n9640 ;
  assign n9643 = n9641 | n9642 ;
  assign n9644 = n9127 | n9136 ;
  assign n9645 = ~n9137 & n9644 ;
  assign n9646 = n9643 & n9645 ;
  assign n9647 = n9643 | n9645 ;
  assign n9648 = ~n9646 & n9647 ;
  assign n9649 = x8 & ~n9132 ;
  assign n9650 = n9134 | n9649 ;
  assign n9651 = n9135 | n9650 ;
  assign n9652 = ~n9136 & n9651 ;
  assign n9653 = ~n2455 & n9245 ;
  assign n9654 = ~n2606 & n8681 ;
  assign n9655 = n9653 | n9654 ;
  assign n9656 = n2569 & n8680 ;
  assign n9657 = n9655 | n9656 ;
  assign n9658 = n8685 | n9657 ;
  assign n9659 = ( ~n5732 & n9657 ) | ( ~n5732 & n9658 ) | ( n9657 & n9658 ) ;
  assign n9660 = ~x5 & n9659 ;
  assign n9661 = x5 | n9660 ;
  assign n9662 = ( ~n9659 & n9660 ) | ( ~n9659 & n9661 ) | ( n9660 & n9661 ) ;
  assign n9663 = n9652 & n9662 ;
  assign n9664 = ~n2764 & n8680 ;
  assign n9665 = ~n2672 & n8681 ;
  assign n9666 = n9664 | n9665 ;
  assign n9667 = n2569 & n9245 ;
  assign n9668 = n9666 | n9667 ;
  assign n9669 = ( n5584 & n8685 ) | ( n5584 & n9668 ) | ( n8685 & n9668 ) ;
  assign n9670 = ( x5 & ~n9668 ) | ( x5 & n9669 ) | ( ~n9668 & n9669 ) ;
  assign n9671 = ~n9669 & n9670 ;
  assign n9672 = n9668 | n9670 ;
  assign n9673 = ( ~x5 & n9671 ) | ( ~x5 & n9672 ) | ( n9671 & n9672 ) ;
  assign n9674 = ~n2764 & n8681 ;
  assign n9675 = ~n2672 & n9245 ;
  assign n9676 = n9674 | n9675 ;
  assign n9677 = n8685 | n9676 ;
  assign n9678 = ( n5932 & n9676 ) | ( n5932 & n9677 ) | ( n9676 & n9677 ) ;
  assign n9679 = ~n2764 & n8678 ;
  assign n9680 = x5 & ~n9679 ;
  assign n9681 = ~x5 & n9678 ;
  assign n9682 = ( ~n9678 & n9680 ) | ( ~n9678 & n9681 ) | ( n9680 & n9681 ) ;
  assign n9683 = n9673 & n9682 ;
  assign n9684 = n9133 & n9683 ;
  assign n9685 = n9683 & ~n9684 ;
  assign n9686 = n9133 & ~n9683 ;
  assign n9687 = ~n2606 & n9245 ;
  assign n9688 = ~n2672 & n8680 ;
  assign n9689 = n9687 | n9688 ;
  assign n9690 = n2569 & n8681 ;
  assign n9691 = n9689 | n9690 ;
  assign n9692 = n8685 | n9691 ;
  assign n9693 = ( n5716 & n9691 ) | ( n5716 & n9692 ) | ( n9691 & n9692 ) ;
  assign n9694 = x5 & n9693 ;
  assign n9695 = x5 & ~n9694 ;
  assign n9696 = ( n9693 & ~n9694 ) | ( n9693 & n9695 ) | ( ~n9694 & n9695 ) ;
  assign n9697 = ( n9685 & n9686 ) | ( n9685 & n9696 ) | ( n9686 & n9696 ) ;
  assign n9698 = n9684 | n9697 ;
  assign n9699 = n9652 | n9662 ;
  assign n9700 = ~n9663 & n9699 ;
  assign n9701 = n9698 & n9700 ;
  assign n9702 = n9663 | n9701 ;
  assign n9703 = n9648 & n9702 ;
  assign n9704 = n9646 | n9703 ;
  assign n9705 = n9622 | n9632 ;
  assign n9706 = ~n9633 & n9705 ;
  assign n9707 = n9704 & n9706 ;
  assign n9708 = n9633 | n9707 ;
  assign n9709 = n9619 & ~n9620 ;
  assign n9710 = ( n9609 & ~n9620 ) | ( n9609 & n9709 ) | ( ~n9620 & n9709 ) ;
  assign n9711 = n9708 & n9710 ;
  assign n9712 = n9596 & ~n9607 ;
  assign n9713 = ~n9596 & n9606 ;
  assign n9714 = n9712 | n9713 ;
  assign n9715 = ( n9620 & n9711 ) | ( n9620 & n9714 ) | ( n9711 & n9714 ) ;
  assign n9716 = n9607 | n9715 ;
  assign n9717 = n9594 & n9716 ;
  assign n9718 = n9591 | n9717 ;
  assign n9719 = n9567 | n9577 ;
  assign n9720 = ~n9578 & n9719 ;
  assign n9721 = n9718 & n9720 ;
  assign n9722 = n9578 | n9721 ;
  assign n9723 = ( n9051 & n9167 ) | ( n9051 & ~n9168 ) | ( n9167 & ~n9168 ) ;
  assign n9724 = ( n9061 & ~n9168 ) | ( n9061 & n9723 ) | ( ~n9168 & n9723 ) ;
  assign n9725 = ( n9565 & n9722 ) | ( n9565 & n9724 ) | ( n9722 & n9724 ) ;
  assign n9726 = n9049 & ~n9169 ;
  assign n9727 = ( n9168 & ~n9169 ) | ( n9168 & n9726 ) | ( ~n9169 & n9726 ) ;
  assign n9728 = ( n9555 & n9725 ) | ( n9555 & n9727 ) | ( n9725 & n9727 ) ;
  assign n9729 = n9545 & n9728 ;
  assign n9730 = n9543 | n9729 ;
  assign n9731 = n9519 & ~n9530 ;
  assign n9732 = ~n9519 & n9529 ;
  assign n9733 = ( n9730 & n9731 ) | ( n9730 & n9732 ) | ( n9731 & n9732 ) ;
  assign n9734 = n9530 | n9733 ;
  assign n9735 = n9504 & ~n9515 ;
  assign n9736 = ~n9504 & n9514 ;
  assign n9737 = ( n9734 & n9735 ) | ( n9734 & n9736 ) | ( n9735 & n9736 ) ;
  assign n9738 = ( n9515 & n9517 ) | ( n9515 & n9737 ) | ( n9517 & n9737 ) ;
  assign n9739 = n9502 | n9738 ;
  assign n9740 = ( n9479 & n9489 ) | ( n9479 & n9739 ) | ( n9489 & n9739 ) ;
  assign n9741 = ( n9466 & n9476 ) | ( n9466 & n9740 ) | ( n9476 & n9740 ) ;
  assign n9742 = ( n9453 & n9463 ) | ( n9453 & n9741 ) | ( n9463 & n9741 ) ;
  assign n9743 = ( n9440 & n9450 ) | ( n9440 & n9742 ) | ( n9450 & n9742 ) ;
  assign n9744 = ( n9428 & n9438 ) | ( n9428 & n9743 ) | ( n9438 & n9743 ) ;
  assign n9745 = n9426 & n9744 ;
  assign n9746 = n9424 | n9745 ;
  assign n9747 = ( n8877 & n9201 ) | ( n8877 & ~n9202 ) | ( n9201 & ~n9202 ) ;
  assign n9748 = ( n8887 & ~n9202 ) | ( n8887 & n9747 ) | ( ~n9202 & n9747 ) ;
  assign n9749 = ( n9411 & n9746 ) | ( n9411 & n9748 ) | ( n9746 & n9748 ) ;
  assign n9750 = ( n8865 & n9202 ) | ( n8865 & ~n9203 ) | ( n9202 & ~n9203 ) ;
  assign n9751 = ( n8875 & ~n9203 ) | ( n8875 & n9750 ) | ( ~n9203 & n9750 ) ;
  assign n9752 = ( n9401 & n9749 ) | ( n9401 & n9751 ) | ( n9749 & n9751 ) ;
  assign n9753 = n9391 & n9752 ;
  assign n9754 = n9389 | n9753 ;
  assign n9755 = n9363 & ~n9374 ;
  assign n9756 = ~n9363 & n9373 ;
  assign n9757 = ( n9754 & n9755 ) | ( n9754 & n9756 ) | ( n9755 & n9756 ) ;
  assign n9758 = ( n9374 & n9376 ) | ( n9374 & n9757 ) | ( n9376 & n9757 ) ;
  assign n9759 = n9361 | n9758 ;
  assign n9760 = ( n9338 & n9348 ) | ( n9338 & n9759 ) | ( n9348 & n9759 ) ;
  assign n9761 = n9324 | n9335 ;
  assign n9762 = ( ~n9334 & n9335 ) | ( ~n9334 & n9761 ) | ( n9335 & n9761 ) ;
  assign n9763 = n9760 & ~n9762 ;
  assign n9764 = n9335 | n9763 ;
  assign n9765 = n9310 | n9321 ;
  assign n9766 = ( ~n9320 & n9321 ) | ( ~n9320 & n9765 ) | ( n9321 & n9765 ) ;
  assign n9767 = n9764 & ~n9766 ;
  assign n9768 = n9321 | n9767 ;
  assign n9769 = n9307 & n9768 ;
  assign n9770 = n9304 | n9769 ;
  assign n9771 = n9279 | n9290 ;
  assign n9772 = ( ~n9289 & n9290 ) | ( ~n9289 & n9771 ) | ( n9290 & n9771 ) ;
  assign n9773 = n9770 & ~n9772 ;
  assign n9774 = n9290 | n9773 ;
  assign n9775 = n9276 & n9774 ;
  assign n9776 = n9276 | n9774 ;
  assign n9777 = ~n9775 & n9776 ;
  assign n9778 = x1 & ~x2 ;
  assign n9779 = ~x1 & x2 ;
  assign n9780 = n9778 | n9779 ;
  assign n9781 = x0 | x1 ;
  assign n9782 = n9780 & ~n9781 ;
  assign n9783 = ~x0 & x1 ;
  assign n9784 = ~n3634 & n9783 ;
  assign n9785 = n672 & n9782 ;
  assign n9786 = ( n9782 & n9784 ) | ( n9782 & ~n9785 ) | ( n9784 & ~n9785 ) ;
  assign n9787 = x0 & n9780 ;
  assign n9788 = n9786 | n9787 ;
  assign n9789 = ( n3726 & n9786 ) | ( n3726 & n9788 ) | ( n9786 & n9788 ) ;
  assign n9790 = x2 & n9789 ;
  assign n9791 = x2 & ~n9790 ;
  assign n9792 = ( n9789 & ~n9790 ) | ( n9789 & n9791 ) | ( ~n9790 & n9791 ) ;
  assign n9793 = n9777 & n9792 ;
  assign n9794 = n9777 | n9792 ;
  assign n9795 = ~n9793 & n9794 ;
  assign n9796 = ~n9770 & n9772 ;
  assign n9797 = n9773 | n9796 ;
  assign n9798 = x0 & ~n9780 ;
  assign n9799 = ~n3634 & n9798 ;
  assign n9800 = ~n672 & n9783 ;
  assign n9801 = n9799 | n9800 ;
  assign n9802 = ~n589 & n9782 ;
  assign n9803 = n9801 | n9802 ;
  assign n9804 = n9787 | n9803 ;
  assign n9805 = ( ~n5092 & n9803 ) | ( ~n5092 & n9804 ) | ( n9803 & n9804 ) ;
  assign n9806 = ~x2 & n9805 ;
  assign n9807 = x2 | n9806 ;
  assign n9808 = ( ~n9805 & n9806 ) | ( ~n9805 & n9807 ) | ( n9806 & n9807 ) ;
  assign n9809 = ~n9797 & n9808 ;
  assign n9810 = n9797 & ~n9808 ;
  assign n9811 = n9809 | n9810 ;
  assign n9812 = n9307 | n9768 ;
  assign n9813 = ~n9769 & n9812 ;
  assign n9814 = ~n3431 & n9782 ;
  assign n9815 = ~n589 & n9783 ;
  assign n9816 = n9814 | n9815 ;
  assign n9817 = ~n672 & n9798 ;
  assign n9818 = n9816 | n9817 ;
  assign n9819 = n9787 | n9818 ;
  assign n9820 = ( ~n5353 & n9818 ) | ( ~n5353 & n9819 ) | ( n9818 & n9819 ) ;
  assign n9821 = ~x2 & n9820 ;
  assign n9822 = x2 | n9821 ;
  assign n9823 = ( ~n9820 & n9821 ) | ( ~n9820 & n9822 ) | ( n9821 & n9822 ) ;
  assign n9824 = n9813 & n9823 ;
  assign n9825 = n9813 | n9823 ;
  assign n9826 = ~n9824 & n9825 ;
  assign n9827 = ~n9764 & n9766 ;
  assign n9828 = n9767 | n9827 ;
  assign n9829 = n3504 & n9782 ;
  assign n9830 = ~n3431 & n9783 ;
  assign n9831 = n9829 | n9830 ;
  assign n9832 = ~n589 & n9798 ;
  assign n9833 = n9831 | n9832 ;
  assign n9834 = n9787 | n9833 ;
  assign n9835 = ( n4765 & n9833 ) | ( n4765 & n9834 ) | ( n9833 & n9834 ) ;
  assign n9836 = x2 & n9835 ;
  assign n9837 = x2 & ~n9836 ;
  assign n9838 = ( n9835 & ~n9836 ) | ( n9835 & n9837 ) | ( ~n9836 & n9837 ) ;
  assign n9839 = n9828 & ~n9838 ;
  assign n9840 = ~n9828 & n9838 ;
  assign n9841 = n9839 | n9840 ;
  assign n9842 = ~n9760 & n9762 ;
  assign n9843 = n9763 | n9842 ;
  assign n9844 = ~n3596 & n9782 ;
  assign n9845 = n3504 & n9783 ;
  assign n9846 = n9844 | n9845 ;
  assign n9847 = ~n3431 & n9798 ;
  assign n9848 = n9846 | n9847 ;
  assign n9849 = n9787 | n9848 ;
  assign n9850 = ( ~n4798 & n9848 ) | ( ~n4798 & n9849 ) | ( n9848 & n9849 ) ;
  assign n9851 = ~x2 & n9850 ;
  assign n9852 = x2 | n9851 ;
  assign n9853 = ( ~n9850 & n9851 ) | ( ~n9850 & n9852 ) | ( n9851 & n9852 ) ;
  assign n9854 = ~n9843 & n9853 ;
  assign n9855 = ~n9841 & n9854 ;
  assign n9856 = n9840 | n9855 ;
  assign n9857 = n9843 | n9854 ;
  assign n9858 = ( ~n9853 & n9854 ) | ( ~n9853 & n9857 ) | ( n9854 & n9857 ) ;
  assign n9859 = n778 & n9782 ;
  assign n9860 = ~n3596 & n9783 ;
  assign n9861 = n9859 | n9860 ;
  assign n9862 = n3504 & n9798 ;
  assign n9863 = n9861 | n9862 ;
  assign n9864 = n9787 | n9863 ;
  assign n9865 = ( ~n5040 & n9863 ) | ( ~n5040 & n9864 ) | ( n9863 & n9864 ) ;
  assign n9866 = ~x2 & n9865 ;
  assign n9867 = x2 | n9866 ;
  assign n9868 = ( ~n9865 & n9866 ) | ( ~n9865 & n9867 ) | ( n9866 & n9867 ) ;
  assign n9869 = n9374 | n9376 ;
  assign n9870 = n9757 | n9869 ;
  assign n9871 = ~n9758 & n9870 ;
  assign n9872 = n9391 | n9752 ;
  assign n9873 = ~n9753 & n9872 ;
  assign n9874 = ~n1014 & n9798 ;
  assign n9875 = n3349 & n9782 ;
  assign n9876 = ~n3255 & n9783 ;
  assign n9877 = n9875 | n9876 ;
  assign n9878 = n9874 | n9877 ;
  assign n9879 = n9787 | n9878 ;
  assign n9880 = ( n4742 & n9878 ) | ( n4742 & n9879 ) | ( n9878 & n9879 ) ;
  assign n9881 = x2 & n9880 ;
  assign n9882 = x2 & ~n9881 ;
  assign n9883 = ( n9880 & ~n9881 ) | ( n9880 & n9882 ) | ( ~n9881 & n9882 ) ;
  assign n9884 = n1233 & n9782 ;
  assign n9885 = n3349 & n9783 ;
  assign n9886 = n9884 | n9885 ;
  assign n9887 = ~n3255 & n9798 ;
  assign n9888 = n9886 | n9887 ;
  assign n9889 = n9787 | n9888 ;
  assign n9890 = ( ~n4470 & n9888 ) | ( ~n4470 & n9889 ) | ( n9888 & n9889 ) ;
  assign n9891 = ~x2 & n9890 ;
  assign n9892 = x2 | n9891 ;
  assign n9893 = ( ~n9890 & n9891 ) | ( ~n9890 & n9892 ) | ( n9891 & n9892 ) ;
  assign n9894 = n9426 | n9744 ;
  assign n9895 = ~n9745 & n9894 ;
  assign n9896 = ( n9428 & n9743 ) | ( n9428 & ~n9744 ) | ( n9743 & ~n9744 ) ;
  assign n9897 = ( n9438 & ~n9744 ) | ( n9438 & n9896 ) | ( ~n9744 & n9896 ) ;
  assign n9898 = ( n9440 & n9742 ) | ( n9440 & ~n9743 ) | ( n9742 & ~n9743 ) ;
  assign n9899 = ( n9450 & ~n9743 ) | ( n9450 & n9898 ) | ( ~n9743 & n9898 ) ;
  assign n9900 = n3178 & n9782 ;
  assign n9901 = n3104 & n9783 ;
  assign n9902 = n9900 | n9901 ;
  assign n9903 = n1327 & n9798 ;
  assign n9904 = n9902 | n9903 ;
  assign n9905 = n9787 | n9904 ;
  assign n9906 = ( n4501 & n9904 ) | ( n4501 & n9905 ) | ( n9904 & n9905 ) ;
  assign n9907 = x2 & n9906 ;
  assign n9908 = x2 & ~n9907 ;
  assign n9909 = ( n9906 & ~n9907 ) | ( n9906 & n9908 ) | ( ~n9907 & n9908 ) ;
  assign n9910 = ~n1411 & n9782 ;
  assign n9911 = n3178 & n9783 ;
  assign n9912 = n9910 | n9911 ;
  assign n9913 = n3104 & n9798 ;
  assign n9914 = n9912 | n9913 ;
  assign n9915 = n9787 | n9914 ;
  assign n9916 = ( n4449 & n9914 ) | ( n4449 & n9915 ) | ( n9914 & n9915 ) ;
  assign n9917 = x2 & n9916 ;
  assign n9918 = x2 & ~n9917 ;
  assign n9919 = ( n9916 & ~n9917 ) | ( n9916 & n9918 ) | ( ~n9917 & n9918 ) ;
  assign n9920 = ~n1411 & n9783 ;
  assign n9921 = n9782 | n9920 ;
  assign n9922 = ( n1532 & n9920 ) | ( n1532 & n9921 ) | ( n9920 & n9921 ) ;
  assign n9923 = n3178 & n9798 ;
  assign n9924 = n9922 | n9923 ;
  assign n9925 = n9787 | n9924 ;
  assign n9926 = ( ~n3750 & n9924 ) | ( ~n3750 & n9925 ) | ( n9924 & n9925 ) ;
  assign n9927 = ~x2 & n9926 ;
  assign n9928 = x2 | n9927 ;
  assign n9929 = ( ~n9926 & n9927 ) | ( ~n9926 & n9928 ) | ( n9927 & n9928 ) ;
  assign n9930 = n9515 | n9517 ;
  assign n9931 = n9737 | n9930 ;
  assign n9932 = ~n9738 & n9931 ;
  assign n9933 = ( ~n9734 & n9735 ) | ( ~n9734 & n9736 ) | ( n9735 & n9736 ) ;
  assign n9934 = n9734 | n9933 ;
  assign n9935 = ~n9737 & n9934 ;
  assign n9936 = n9545 | n9728 ;
  assign n9937 = ~n9729 & n9936 ;
  assign n9938 = ~n2873 & n9782 ;
  assign n9939 = ~n1733 & n9783 ;
  assign n9940 = n9938 | n9939 ;
  assign n9941 = n1625 & n9798 ;
  assign n9942 = n9940 | n9941 ;
  assign n9943 = n9787 | n9942 ;
  assign n9944 = ( n4260 & n9942 ) | ( n4260 & n9943 ) | ( n9942 & n9943 ) ;
  assign n9945 = x2 & n9944 ;
  assign n9946 = x2 & ~n9945 ;
  assign n9947 = ( n9944 & ~n9945 ) | ( n9944 & n9946 ) | ( ~n9945 & n9946 ) ;
  assign n9948 = n1803 & n9782 ;
  assign n9949 = ~n2873 & n9783 ;
  assign n9950 = n9948 | n9949 ;
  assign n9951 = ~n1733 & n9798 ;
  assign n9952 = n9950 | n9951 ;
  assign n9953 = n9787 | n9952 ;
  assign n9954 = ( ~n4985 & n9952 ) | ( ~n4985 & n9953 ) | ( n9952 & n9953 ) ;
  assign n9955 = ~x2 & n9954 ;
  assign n9956 = x2 | n9955 ;
  assign n9957 = ( ~n9954 & n9955 ) | ( ~n9954 & n9956 ) | ( n9955 & n9956 ) ;
  assign n9958 = n9718 | n9720 ;
  assign n9959 = ~n9721 & n9958 ;
  assign n9960 = n9594 | n9716 ;
  assign n9961 = ~n9717 & n9960 ;
  assign n9962 = n9620 | n9714 ;
  assign n9963 = n9711 | n9962 ;
  assign n9964 = ~n9715 & n9963 ;
  assign n9965 = n2193 & n9782 ;
  assign n9966 = n2013 & n9783 ;
  assign n9967 = n9965 | n9966 ;
  assign n9968 = ~n2103 & n9798 ;
  assign n9969 = n9967 | n9968 ;
  assign n9970 = n9787 | n9969 ;
  assign n9971 = ( ~n5836 & n9969 ) | ( ~n5836 & n9970 ) | ( n9969 & n9970 ) ;
  assign n9972 = ~x2 & n9971 ;
  assign n9973 = x2 | n9972 ;
  assign n9974 = ( ~n9971 & n9972 ) | ( ~n9971 & n9973 ) | ( n9972 & n9973 ) ;
  assign n9975 = n2296 & n9782 ;
  assign n9976 = n2193 & n9783 ;
  assign n9977 = n9975 | n9976 ;
  assign n9978 = n2013 & n9798 ;
  assign n9979 = n9977 | n9978 ;
  assign n9980 = n9787 | n9979 ;
  assign n9981 = ( n5216 & n9979 ) | ( n5216 & n9980 ) | ( n9979 & n9980 ) ;
  assign n9982 = x2 & n9981 ;
  assign n9983 = x2 & ~n9982 ;
  assign n9984 = ( n9981 & ~n9982 ) | ( n9981 & n9983 ) | ( ~n9982 & n9983 ) ;
  assign n9985 = n9698 | n9700 ;
  assign n9986 = ~n9701 & n9985 ;
  assign n9987 = ~n2455 & n9782 ;
  assign n9988 = ~n2375 & n9783 ;
  assign n9989 = n9987 | n9988 ;
  assign n9990 = n2296 & n9798 ;
  assign n9991 = n9989 | n9990 ;
  assign n9992 = n9787 | n9991 ;
  assign n9993 = ( n5781 & n9991 ) | ( n5781 & n9992 ) | ( n9991 & n9992 ) ;
  assign n9994 = x2 & n9993 ;
  assign n9995 = x2 & ~n9994 ;
  assign n9996 = ( n9993 & ~n9994 ) | ( n9993 & n9995 ) | ( ~n9994 & n9995 ) ;
  assign n9997 = n9673 | n9682 ;
  assign n9998 = ~n9683 & n9997 ;
  assign n9999 = ~n2455 & n9798 ;
  assign n10000 = ~n2606 & n9783 ;
  assign n10001 = n9999 | n10000 ;
  assign n10002 = n2569 & n9782 ;
  assign n10003 = n10001 | n10002 ;
  assign n10004 = n9787 | n10003 ;
  assign n10005 = ( ~n5732 & n10003 ) | ( ~n5732 & n10004 ) | ( n10003 & n10004 ) ;
  assign n10006 = ~x2 & n10005 ;
  assign n10007 = x2 | n10006 ;
  assign n10008 = ( ~n10005 & n10006 ) | ( ~n10005 & n10007 ) | ( n10006 & n10007 ) ;
  assign n10009 = ~n2606 & n9798 ;
  assign n10010 = ~n2672 & n9782 ;
  assign n10011 = n10009 | n10010 ;
  assign n10012 = n2569 & n9783 ;
  assign n10013 = n10011 | n10012 ;
  assign n10014 = n9787 | n10013 ;
  assign n10015 = ( n5716 & n10013 ) | ( n5716 & n10014 ) | ( n10013 & n10014 ) ;
  assign n10016 = x2 & n10015 ;
  assign n10017 = x2 & ~n10016 ;
  assign n10018 = ( n10015 & ~n10016 ) | ( n10015 & n10017 ) | ( ~n10016 & n10017 ) ;
  assign n10019 = x0 & x2 ;
  assign n10020 = n9780 & n10019 ;
  assign n10021 = n5584 & n10020 ;
  assign n10022 = ~n2764 & n9782 ;
  assign n10023 = ~n2672 & n9783 ;
  assign n10024 = n10022 | n10023 ;
  assign n10025 = n2569 & n9798 ;
  assign n10026 = n10024 | n10025 ;
  assign n10027 = x2 & n10026 ;
  assign n10028 = ~n9780 & n10019 ;
  assign n10029 = n2671 & n10028 ;
  assign n10030 = x2 & ~n10029 ;
  assign n10031 = x2 & ~n10028 ;
  assign n10032 = ( n2667 & n10030 ) | ( n2667 & n10031 ) | ( n10030 & n10031 ) ;
  assign n10033 = x2 & n9783 ;
  assign n10034 = ~n2764 & n10033 ;
  assign n10035 = n10032 & ~n10034 ;
  assign n10036 = ~n10020 & n10035 ;
  assign n10037 = ( ~n5932 & n10035 ) | ( ~n5932 & n10036 ) | ( n10035 & n10036 ) ;
  assign n10038 = ~n10027 & n10037 ;
  assign n10039 = ~n10021 & n10038 ;
  assign n10040 = x0 & ~n2764 ;
  assign n10041 = n10039 & ~n10040 ;
  assign n10042 = ( n9679 & n10018 ) | ( n9679 & n10041 ) | ( n10018 & n10041 ) ;
  assign n10043 = n10008 & n10042 ;
  assign n10044 = n9998 & n10043 ;
  assign n10045 = ( x5 & n9678 ) | ( x5 & ~n9680 ) | ( n9678 & ~n9680 ) ;
  assign n10046 = n10008 | n10042 ;
  assign n10047 = x5 & ~n9680 ;
  assign n10048 = ( n9678 & ~n10046 ) | ( n9678 & n10047 ) | ( ~n10046 & n10047 ) ;
  assign n10049 = n10045 & ~n10048 ;
  assign n10050 = ( n9998 & n10044 ) | ( n9998 & n10049 ) | ( n10044 & n10049 ) ;
  assign n10051 = n9996 & n10050 ;
  assign n10052 = ~n2606 & n9782 ;
  assign n10053 = ~n2455 & n9783 ;
  assign n10054 = n10052 | n10053 ;
  assign n10055 = ~n2375 & n9798 ;
  assign n10056 = n10054 | n10055 ;
  assign n10057 = n9787 | n10056 ;
  assign n10058 = ( ~n5528 & n10056 ) | ( ~n5528 & n10057 ) | ( n10056 & n10057 ) ;
  assign n10059 = ~x2 & n10058 ;
  assign n10060 = n9998 | n10043 ;
  assign n10061 = n10049 | n10060 ;
  assign n10062 = ( ~n10058 & n10059 ) | ( ~n10058 & n10061 ) | ( n10059 & n10061 ) ;
  assign n10063 = ( x2 & n10059 ) | ( x2 & n10062 ) | ( n10059 & n10062 ) ;
  assign n10064 = ( n9996 & n10051 ) | ( n9996 & n10063 ) | ( n10051 & n10063 ) ;
  assign n10065 = n9986 & n10064 ;
  assign n10066 = n9996 | n10050 ;
  assign n10067 = n10063 | n10066 ;
  assign n10068 = n9685 | n9696 ;
  assign n10069 = ( n9686 & n10067 ) | ( n9686 & n10068 ) | ( n10067 & n10068 ) ;
  assign n10070 = ~n9697 & n10069 ;
  assign n10071 = ( n9986 & n10065 ) | ( n9986 & n10070 ) | ( n10065 & n10070 ) ;
  assign n10072 = n9984 & n10071 ;
  assign n10073 = ~n2375 & n9782 ;
  assign n10074 = n2296 & n9783 ;
  assign n10075 = n10073 | n10074 ;
  assign n10076 = n2193 & n9798 ;
  assign n10077 = n10075 | n10076 ;
  assign n10078 = n9787 | n10077 ;
  assign n10079 = ( ~n5879 & n10077 ) | ( ~n5879 & n10078 ) | ( n10077 & n10078 ) ;
  assign n10080 = ~x2 & n10079 ;
  assign n10081 = n9986 | n10064 ;
  assign n10082 = n10070 | n10081 ;
  assign n10083 = ( ~n10079 & n10080 ) | ( ~n10079 & n10082 ) | ( n10080 & n10082 ) ;
  assign n10084 = ( x2 & n10080 ) | ( x2 & n10083 ) | ( n10080 & n10083 ) ;
  assign n10085 = ( n9984 & n10072 ) | ( n9984 & n10084 ) | ( n10072 & n10084 ) ;
  assign n10086 = n9974 | n10085 ;
  assign n10087 = n9984 | n10071 ;
  assign n10088 = n10084 | n10087 ;
  assign n10089 = ( n9648 & n9702 ) | ( n9648 & n10088 ) | ( n9702 & n10088 ) ;
  assign n10090 = ~n9703 & n10089 ;
  assign n10091 = n10086 | n10090 ;
  assign n10092 = ( n9704 & n9706 ) | ( n9704 & n10091 ) | ( n9706 & n10091 ) ;
  assign n10093 = ~n9707 & n10092 ;
  assign n10094 = n2013 & n9782 ;
  assign n10095 = ~n2103 & n9783 ;
  assign n10096 = n10094 | n10095 ;
  assign n10097 = ~n1944 & n9798 ;
  assign n10098 = n10096 | n10097 ;
  assign n10099 = n9787 | n10098 ;
  assign n10100 = ( n6041 & n10098 ) | ( n6041 & n10099 ) | ( n10098 & n10099 ) ;
  assign n10101 = x2 & n10100 ;
  assign n10102 = x2 & ~n10101 ;
  assign n10103 = ( n10100 & ~n10101 ) | ( n10100 & n10102 ) | ( ~n10101 & n10102 ) ;
  assign n10104 = n9974 & n10085 ;
  assign n10105 = ( n9974 & n10090 ) | ( n9974 & n10104 ) | ( n10090 & n10104 ) ;
  assign n10106 = n10103 | n10105 ;
  assign n10107 = n10093 | n10106 ;
  assign n10108 = ( n9708 & n9710 ) | ( n9708 & n10107 ) | ( n9710 & n10107 ) ;
  assign n10109 = ~n9711 & n10108 ;
  assign n10110 = n10103 & n10105 ;
  assign n10111 = ( n10093 & n10103 ) | ( n10093 & n10110 ) | ( n10103 & n10110 ) ;
  assign n10112 = n9964 & n10111 ;
  assign n10113 = ( n9964 & n10109 ) | ( n9964 & n10112 ) | ( n10109 & n10112 ) ;
  assign n10114 = n9961 & n10113 ;
  assign n10115 = ~n2103 & n9782 ;
  assign n10116 = ~n1944 & n9783 ;
  assign n10117 = n10115 | n10116 ;
  assign n10118 = ~n1880 & n9798 ;
  assign n10119 = n10117 | n10118 ;
  assign n10120 = n9787 | n10119 ;
  assign n10121 = ( ~n5281 & n10119 ) | ( ~n5281 & n10120 ) | ( n10119 & n10120 ) ;
  assign n10122 = ~x2 & n10121 ;
  assign n10123 = n9964 | n10111 ;
  assign n10124 = n10109 | n10123 ;
  assign n10125 = ( ~n10121 & n10122 ) | ( ~n10121 & n10124 ) | ( n10122 & n10124 ) ;
  assign n10126 = ( x2 & n10122 ) | ( x2 & n10125 ) | ( n10122 & n10125 ) ;
  assign n10127 = ( n9961 & n10114 ) | ( n9961 & n10126 ) | ( n10114 & n10126 ) ;
  assign n10128 = n9959 & n10127 ;
  assign n10129 = n1803 & n9798 ;
  assign n10130 = ~n1944 & n9782 ;
  assign n10131 = n10129 | n10130 ;
  assign n10132 = ~n1880 & n9783 ;
  assign n10133 = n10131 | n10132 ;
  assign n10134 = n9787 | n10133 ;
  assign n10135 = ( n4905 & n10133 ) | ( n4905 & n10134 ) | ( n10133 & n10134 ) ;
  assign n10136 = ~x2 & n10135 ;
  assign n10137 = n9961 | n10113 ;
  assign n10138 = n10126 | n10137 ;
  assign n10139 = ( ~n10135 & n10136 ) | ( ~n10135 & n10138 ) | ( n10136 & n10138 ) ;
  assign n10140 = ( x2 & n10136 ) | ( x2 & n10139 ) | ( n10136 & n10139 ) ;
  assign n10141 = ( n9959 & n10128 ) | ( n9959 & n10140 ) | ( n10128 & n10140 ) ;
  assign n10142 = n9957 & n10141 ;
  assign n10143 = ~n2873 & n9798 ;
  assign n10144 = n1803 & n9783 ;
  assign n10145 = n10143 | n10144 ;
  assign n10146 = ~n1880 & n9782 ;
  assign n10147 = n10145 | n10146 ;
  assign n10148 = n9787 | n10147 ;
  assign n10149 = ( n5139 & n10147 ) | ( n5139 & n10148 ) | ( n10147 & n10148 ) ;
  assign n10150 = ~x2 & n10149 ;
  assign n10151 = n9959 | n10127 ;
  assign n10152 = n10140 | n10151 ;
  assign n10153 = ( ~n10149 & n10150 ) | ( ~n10149 & n10152 ) | ( n10150 & n10152 ) ;
  assign n10154 = ( x2 & n10150 ) | ( x2 & n10153 ) | ( n10150 & n10153 ) ;
  assign n10155 = ( n9957 & n10142 ) | ( n9957 & n10154 ) | ( n10142 & n10154 ) ;
  assign n10156 = n9947 & n10155 ;
  assign n10157 = n9957 | n10141 ;
  assign n10158 = n10154 | n10157 ;
  assign n10159 = ( n9565 & n9722 ) | ( n9565 & ~n9724 ) | ( n9722 & ~n9724 ) ;
  assign n10160 = ( ~n9565 & n9722 ) | ( ~n9565 & n9724 ) | ( n9722 & n9724 ) ;
  assign n10161 = ( ~n9722 & n10159 ) | ( ~n9722 & n10160 ) | ( n10159 & n10160 ) ;
  assign n10162 = n10158 & n10161 ;
  assign n10163 = ( n9947 & n10156 ) | ( n9947 & n10162 ) | ( n10156 & n10162 ) ;
  assign n10164 = ~n1733 & n9782 ;
  assign n10165 = n1625 & n9783 ;
  assign n10166 = n10164 | n10165 ;
  assign n10167 = n3030 & n9798 ;
  assign n10168 = n10166 | n10167 ;
  assign n10169 = n9787 | n10168 ;
  assign n10170 = ( ~n4578 & n10168 ) | ( ~n4578 & n10169 ) | ( n10168 & n10169 ) ;
  assign n10171 = ~x2 & n10170 ;
  assign n10172 = x2 | n10171 ;
  assign n10173 = ( ~n10170 & n10171 ) | ( ~n10170 & n10172 ) | ( n10171 & n10172 ) ;
  assign n10174 = n10163 | n10173 ;
  assign n10175 = n9947 | n10155 ;
  assign n10176 = n10162 | n10175 ;
  assign n10177 = ( n9555 & n9725 ) | ( n9555 & ~n9727 ) | ( n9725 & ~n9727 ) ;
  assign n10178 = ( ~n9555 & n9725 ) | ( ~n9555 & n9727 ) | ( n9725 & n9727 ) ;
  assign n10179 = ( ~n9725 & n10177 ) | ( ~n9725 & n10178 ) | ( n10177 & n10178 ) ;
  assign n10180 = n10176 & n10179 ;
  assign n10181 = n10174 | n10180 ;
  assign n10182 = n9937 & n10181 ;
  assign n10183 = ( ~n9730 & n9731 ) | ( ~n9730 & n9732 ) | ( n9731 & n9732 ) ;
  assign n10184 = n9730 | n10183 ;
  assign n10185 = ~n9733 & n10184 ;
  assign n10186 = n10163 & n10173 ;
  assign n10187 = ( n10173 & n10180 ) | ( n10173 & n10186 ) | ( n10180 & n10186 ) ;
  assign n10188 = n10185 & n10187 ;
  assign n10189 = ( n10182 & n10185 ) | ( n10182 & n10188 ) | ( n10185 & n10188 ) ;
  assign n10190 = n9935 & n10189 ;
  assign n10191 = n1625 & n9782 ;
  assign n10192 = n3030 & n9783 ;
  assign n10193 = n10191 | n10192 ;
  assign n10194 = ~n2939 & n9798 ;
  assign n10195 = n10193 | n10194 ;
  assign n10196 = n9787 | n10195 ;
  assign n10197 = ( ~n4215 & n10195 ) | ( ~n4215 & n10196 ) | ( n10195 & n10196 ) ;
  assign n10198 = ~x2 & n10197 ;
  assign n10199 = n10185 | n10187 ;
  assign n10200 = n10182 | n10199 ;
  assign n10201 = ( ~n10197 & n10198 ) | ( ~n10197 & n10200 ) | ( n10198 & n10200 ) ;
  assign n10202 = ( x2 & n10198 ) | ( x2 & n10201 ) | ( n10198 & n10201 ) ;
  assign n10203 = ( n9935 & n10190 ) | ( n9935 & n10202 ) | ( n10190 & n10202 ) ;
  assign n10204 = n9932 & n10203 ;
  assign n10205 = n1532 & n9798 ;
  assign n10206 = n3030 & n9782 ;
  assign n10207 = ~n2939 & n9783 ;
  assign n10208 = n10206 | n10207 ;
  assign n10209 = n10205 | n10208 ;
  assign n10210 = n9787 | n10209 ;
  assign n10211 = ( ~n4193 & n10209 ) | ( ~n4193 & n10210 ) | ( n10209 & n10210 ) ;
  assign n10212 = ~x2 & n10211 ;
  assign n10213 = n9935 | n10189 ;
  assign n10214 = n10202 | n10213 ;
  assign n10215 = ( ~n10211 & n10212 ) | ( ~n10211 & n10214 ) | ( n10212 & n10214 ) ;
  assign n10216 = ( x2 & n10212 ) | ( x2 & n10215 ) | ( n10212 & n10215 ) ;
  assign n10217 = ( n9932 & n10204 ) | ( n9932 & n10216 ) | ( n10204 & n10216 ) ;
  assign n10218 = n9929 & n10217 ;
  assign n10219 = n1532 & n9783 ;
  assign n10220 = ~n1411 & n9798 ;
  assign n10221 = ~n2939 & n9782 ;
  assign n10222 = n10220 | n10221 ;
  assign n10223 = n10219 | n10222 ;
  assign n10224 = n9787 | n10223 ;
  assign n10225 = ( ~n3930 & n10223 ) | ( ~n3930 & n10224 ) | ( n10223 & n10224 ) ;
  assign n10226 = ~x2 & n10225 ;
  assign n10227 = n9932 | n10203 ;
  assign n10228 = n10216 | n10227 ;
  assign n10229 = ( ~n10225 & n10226 ) | ( ~n10225 & n10228 ) | ( n10226 & n10228 ) ;
  assign n10230 = ( x2 & n10226 ) | ( x2 & n10229 ) | ( n10226 & n10229 ) ;
  assign n10231 = ( n9929 & n10218 ) | ( n9929 & n10230 ) | ( n10218 & n10230 ) ;
  assign n10232 = n9919 & n10231 ;
  assign n10233 = n9929 | n10217 ;
  assign n10234 = n10230 | n10233 ;
  assign n10235 = ( ~n9479 & n9489 ) | ( ~n9479 & n9739 ) | ( n9489 & n9739 ) ;
  assign n10236 = ( n9479 & ~n9489 ) | ( n9479 & n9739 ) | ( ~n9489 & n9739 ) ;
  assign n10237 = ( ~n9739 & n10235 ) | ( ~n9739 & n10236 ) | ( n10235 & n10236 ) ;
  assign n10238 = n10234 & n10237 ;
  assign n10239 = ( n9919 & n10232 ) | ( n9919 & n10238 ) | ( n10232 & n10238 ) ;
  assign n10240 = n9909 & n10239 ;
  assign n10241 = n9919 | n10231 ;
  assign n10242 = n10238 | n10241 ;
  assign n10243 = ( ~n9466 & n9476 ) | ( ~n9466 & n9740 ) | ( n9476 & n9740 ) ;
  assign n10244 = ( n9466 & ~n9476 ) | ( n9466 & n9740 ) | ( ~n9476 & n9740 ) ;
  assign n10245 = ( ~n9740 & n10243 ) | ( ~n9740 & n10244 ) | ( n10243 & n10244 ) ;
  assign n10246 = n10242 & n10245 ;
  assign n10247 = ( n9909 & n10240 ) | ( n9909 & n10246 ) | ( n10240 & n10246 ) ;
  assign n10248 = n9899 & n10247 ;
  assign n10249 = n9909 | n10239 ;
  assign n10250 = n10246 | n10249 ;
  assign n10251 = ( ~n9453 & n9463 ) | ( ~n9453 & n9741 ) | ( n9463 & n9741 ) ;
  assign n10252 = ( n9453 & ~n9463 ) | ( n9453 & n9741 ) | ( ~n9463 & n9741 ) ;
  assign n10253 = ( ~n9741 & n10251 ) | ( ~n9741 & n10252 ) | ( n10251 & n10252 ) ;
  assign n10254 = n10250 & n10253 ;
  assign n10255 = ( n9899 & n10248 ) | ( n9899 & n10254 ) | ( n10248 & n10254 ) ;
  assign n10256 = n9897 & n10255 ;
  assign n10257 = n3104 & n9782 ;
  assign n10258 = n1327 & n9783 ;
  assign n10259 = n10257 | n10258 ;
  assign n10260 = ~n1151 & n9798 ;
  assign n10261 = n10259 | n10260 ;
  assign n10262 = n9787 | n10261 ;
  assign n10263 = ( ~n4034 & n10261 ) | ( ~n4034 & n10262 ) | ( n10261 & n10262 ) ;
  assign n10264 = ~x2 & n10263 ;
  assign n10265 = n9899 | n10247 ;
  assign n10266 = n10254 | n10265 ;
  assign n10267 = ( ~n10263 & n10264 ) | ( ~n10263 & n10266 ) | ( n10264 & n10266 ) ;
  assign n10268 = ( x2 & n10264 ) | ( x2 & n10267 ) | ( n10264 & n10267 ) ;
  assign n10269 = ( n9897 & n10256 ) | ( n9897 & n10268 ) | ( n10256 & n10268 ) ;
  assign n10270 = n9895 & n10269 ;
  assign n10271 = n1327 & n9782 ;
  assign n10272 = ~n1151 & n9783 ;
  assign n10273 = n10271 | n10272 ;
  assign n10274 = n1233 & n9798 ;
  assign n10275 = n10273 | n10274 ;
  assign n10276 = n9787 | n10275 ;
  assign n10277 = ( ~n4615 & n10275 ) | ( ~n4615 & n10276 ) | ( n10275 & n10276 ) ;
  assign n10278 = ~x2 & n10277 ;
  assign n10279 = n9897 | n10255 ;
  assign n10280 = n10268 | n10279 ;
  assign n10281 = ( ~n10277 & n10278 ) | ( ~n10277 & n10280 ) | ( n10278 & n10280 ) ;
  assign n10282 = ( x2 & n10278 ) | ( x2 & n10281 ) | ( n10278 & n10281 ) ;
  assign n10283 = ( n9895 & n10270 ) | ( n9895 & n10282 ) | ( n10270 & n10282 ) ;
  assign n10284 = n9893 & n10283 ;
  assign n10285 = ~n1151 & n9782 ;
  assign n10286 = n1233 & n9783 ;
  assign n10287 = n10285 | n10286 ;
  assign n10288 = n3349 & n9798 ;
  assign n10289 = n10287 | n10288 ;
  assign n10290 = n9787 | n10289 ;
  assign n10291 = ( n4518 & n10289 ) | ( n4518 & n10290 ) | ( n10289 & n10290 ) ;
  assign n10292 = ~x2 & n10291 ;
  assign n10293 = n9895 | n10269 ;
  assign n10294 = n10282 | n10293 ;
  assign n10295 = ( ~n10291 & n10292 ) | ( ~n10291 & n10294 ) | ( n10292 & n10294 ) ;
  assign n10296 = ( x2 & n10292 ) | ( x2 & n10295 ) | ( n10292 & n10295 ) ;
  assign n10297 = ( n9893 & n10284 ) | ( n9893 & n10296 ) | ( n10284 & n10296 ) ;
  assign n10298 = n9883 & n10297 ;
  assign n10299 = n9893 | n10283 ;
  assign n10300 = n10296 | n10299 ;
  assign n10301 = ( n9411 & n9746 ) | ( n9411 & ~n9748 ) | ( n9746 & ~n9748 ) ;
  assign n10302 = ( ~n9411 & n9746 ) | ( ~n9411 & n9748 ) | ( n9746 & n9748 ) ;
  assign n10303 = ( ~n9746 & n10301 ) | ( ~n9746 & n10302 ) | ( n10301 & n10302 ) ;
  assign n10304 = n10300 & n10303 ;
  assign n10305 = ( n9883 & n10298 ) | ( n9883 & n10304 ) | ( n10298 & n10304 ) ;
  assign n10306 = ~n1014 & n9783 ;
  assign n10307 = ~n3255 & n9782 ;
  assign n10308 = n10306 | n10307 ;
  assign n10309 = n904 & n9798 ;
  assign n10310 = n10308 | n10309 ;
  assign n10311 = n9787 | n10310 ;
  assign n10312 = ( n4632 & n10310 ) | ( n4632 & n10311 ) | ( n10310 & n10311 ) ;
  assign n10313 = x2 & n10312 ;
  assign n10314 = x2 & ~n10313 ;
  assign n10315 = ( n10312 & ~n10313 ) | ( n10312 & n10314 ) | ( ~n10313 & n10314 ) ;
  assign n10316 = n10305 | n10315 ;
  assign n10317 = n9883 | n10297 ;
  assign n10318 = n10304 | n10317 ;
  assign n10319 = ( n9401 & n9749 ) | ( n9401 & ~n9751 ) | ( n9749 & ~n9751 ) ;
  assign n10320 = ( ~n9401 & n9749 ) | ( ~n9401 & n9751 ) | ( n9749 & n9751 ) ;
  assign n10321 = ( ~n9749 & n10319 ) | ( ~n9749 & n10320 ) | ( n10319 & n10320 ) ;
  assign n10322 = n10318 & n10321 ;
  assign n10323 = n10316 | n10322 ;
  assign n10324 = n9873 & n10323 ;
  assign n10325 = ( ~n9754 & n9755 ) | ( ~n9754 & n9756 ) | ( n9755 & n9756 ) ;
  assign n10326 = n9754 | n10325 ;
  assign n10327 = ~n9757 & n10326 ;
  assign n10328 = n10305 & n10315 ;
  assign n10329 = ( n10315 & n10322 ) | ( n10315 & n10328 ) | ( n10322 & n10328 ) ;
  assign n10330 = n10327 & n10329 ;
  assign n10331 = ( n10324 & n10327 ) | ( n10324 & n10330 ) | ( n10327 & n10330 ) ;
  assign n10332 = n9871 & n10331 ;
  assign n10333 = ~n1014 & n9782 ;
  assign n10334 = n904 & n9783 ;
  assign n10335 = n10333 | n10334 ;
  assign n10336 = n778 & n9798 ;
  assign n10337 = n10335 | n10336 ;
  assign n10338 = n9787 | n10337 ;
  assign n10339 = ( ~n4535 & n10337 ) | ( ~n4535 & n10338 ) | ( n10337 & n10338 ) ;
  assign n10340 = ~x2 & n10339 ;
  assign n10341 = n10327 | n10329 ;
  assign n10342 = n10324 | n10341 ;
  assign n10343 = ( ~n10339 & n10340 ) | ( ~n10339 & n10342 ) | ( n10340 & n10342 ) ;
  assign n10344 = ( x2 & n10340 ) | ( x2 & n10343 ) | ( n10340 & n10343 ) ;
  assign n10345 = ( n9871 & n10332 ) | ( n9871 & n10344 ) | ( n10332 & n10344 ) ;
  assign n10346 = n9868 & n10345 ;
  assign n10347 = n904 & n9782 ;
  assign n10348 = n778 & n9783 ;
  assign n10349 = n10347 | n10348 ;
  assign n10350 = ~n3596 & n9798 ;
  assign n10351 = n10349 | n10350 ;
  assign n10352 = n9787 | n10351 ;
  assign n10353 = ( ~n4649 & n10351 ) | ( ~n4649 & n10352 ) | ( n10351 & n10352 ) ;
  assign n10354 = ~x2 & n10353 ;
  assign n10355 = n9871 | n10331 ;
  assign n10356 = n10344 | n10355 ;
  assign n10357 = ( ~n10353 & n10354 ) | ( ~n10353 & n10356 ) | ( n10354 & n10356 ) ;
  assign n10358 = ( x2 & n10354 ) | ( x2 & n10357 ) | ( n10354 & n10357 ) ;
  assign n10359 = ( n9868 & n10346 ) | ( n9868 & n10358 ) | ( n10346 & n10358 ) ;
  assign n10360 = ~n9338 & n9348 ;
  assign n10361 = n9338 & ~n9348 ;
  assign n10362 = n10360 | n10361 ;
  assign n10363 = n9759 | n10362 ;
  assign n10364 = n9868 | n10345 ;
  assign n10365 = n10358 | n10364 ;
  assign n10366 = ( n9759 & n10362 ) | ( n9759 & ~n10365 ) | ( n10362 & ~n10365 ) ;
  assign n10367 = ( n10359 & n10363 ) | ( n10359 & ~n10366 ) | ( n10363 & ~n10366 ) ;
  assign n10368 = ~n9858 & n10367 ;
  assign n10369 = ( ~n9839 & n9856 ) | ( ~n9839 & n10368 ) | ( n9856 & n10368 ) ;
  assign n10370 = n9826 & n10369 ;
  assign n10371 = n9824 | n10370 ;
  assign n10372 = ~n9811 & n10371 ;
  assign n10373 = n9809 | n10372 ;
  assign n10374 = n9795 & n10373 ;
  assign n10375 = n9236 & ~n9240 ;
  assign n10376 = n9239 & ~n9240 ;
  assign n10377 = n10375 | n10376 ;
  assign n10378 = ~n3431 & n8680 ;
  assign n10379 = ~n589 & n8681 ;
  assign n10380 = n10378 | n10379 ;
  assign n10381 = ~n672 & n9245 ;
  assign n10382 = n10380 | n10381 ;
  assign n10383 = n8685 | n10382 ;
  assign n10384 = ( ~n5353 & n10382 ) | ( ~n5353 & n10383 ) | ( n10382 & n10383 ) ;
  assign n10385 = ~x5 & n10384 ;
  assign n10386 = x5 | n10385 ;
  assign n10387 = ( ~n10384 & n10385 ) | ( ~n10384 & n10386 ) | ( n10385 & n10386 ) ;
  assign n10388 = n9782 | n9787 ;
  assign n10389 = ~n3634 & n10388 ;
  assign n10390 = ( ~n672 & n9785 ) | ( ~n672 & n10389 ) | ( n9785 & n10389 ) ;
  assign n10391 = ( ~n3619 & n10389 ) | ( ~n3619 & n10390 ) | ( n10389 & n10390 ) ;
  assign n10392 = ~x2 & n10391 ;
  assign n10393 = x2 | n10392 ;
  assign n10394 = ( ~n10391 & n10392 ) | ( ~n10391 & n10393 ) | ( n10392 & n10393 ) ;
  assign n10395 = n10387 & n10394 ;
  assign n10396 = n10394 & ~n10395 ;
  assign n10397 = ( n10387 & ~n10395 ) | ( n10387 & n10396 ) | ( ~n10395 & n10396 ) ;
  assign n10398 = ~n10377 & n10397 ;
  assign n10399 = n10377 & ~n10397 ;
  assign n10400 = n10398 | n10399 ;
  assign n10401 = n9273 | n9775 ;
  assign n10402 = n10400 & n10401 ;
  assign n10403 = n10400 | n10401 ;
  assign n10404 = ~n10402 & n10403 ;
  assign n10405 = ( n9793 & n10374 ) | ( n9793 & n10404 ) | ( n10374 & n10404 ) ;
  assign n10406 = n9241 & n9244 ;
  assign n10407 = n9256 & ~n10406 ;
  assign n10408 = n9241 & ~n10406 ;
  assign n10409 = n9244 & ~n10406 ;
  assign n10410 = n10408 | n10409 ;
  assign n10411 = n9255 | n10410 ;
  assign n10412 = ( n10377 & n10387 ) | ( n10377 & n10394 ) | ( n10387 & n10394 ) ;
  assign n10413 = ( ~n10407 & n10411 ) | ( ~n10407 & n10412 ) | ( n10411 & n10412 ) ;
  assign n10414 = n10411 & n10412 ;
  assign n10415 = ~n10407 & n10414 ;
  assign n10416 = n10413 & ~n10415 ;
  assign n10417 = n10402 & n10416 ;
  assign n10418 = n10415 | n10417 ;
  assign n10419 = ( n10405 & n10413 ) | ( n10405 & n10418 ) | ( n10413 & n10418 ) ;
  assign n10420 = n9259 & n10419 ;
  assign n10421 = n7668 | n7669 ;
  assign n10422 = n7546 | n10421 ;
  assign n10423 = ~n7670 & n10422 ;
  assign n10424 = n8680 | n8685 ;
  assign n10425 = ~n3634 & n10424 ;
  assign n10426 = ( ~n672 & n8683 ) | ( ~n672 & n10425 ) | ( n8683 & n10425 ) ;
  assign n10427 = ( ~n3619 & n10425 ) | ( ~n3619 & n10426 ) | ( n10425 & n10426 ) ;
  assign n10428 = ~x5 & n10427 ;
  assign n10429 = x5 | n10428 ;
  assign n10430 = ( ~n10427 & n10428 ) | ( ~n10427 & n10429 ) | ( n10428 & n10429 ) ;
  assign n10431 = ( n8717 & n8718 ) | ( n8717 & n8721 ) | ( n8718 & n8721 ) ;
  assign n10432 = n10430 & n10431 ;
  assign n10433 = ( ~n7542 & n7543 ) | ( ~n7542 & n7544 ) | ( n7543 & n7544 ) ;
  assign n10434 = n10430 | n10431 ;
  assign n10435 = ~n10432 & n10434 ;
  assign n10436 = ~n10433 & n10435 ;
  assign n10437 = n10432 | n10436 ;
  assign n10438 = n10423 & n10437 ;
  assign n10439 = n10423 | n10437 ;
  assign n10440 = ~n10438 & n10439 ;
  assign n10441 = n10433 | n10436 ;
  assign n10442 = ( ~n10435 & n10436 ) | ( ~n10435 & n10441 ) | ( n10436 & n10441 ) ;
  assign n10443 = n8706 | n8725 ;
  assign n10444 = ~n10442 & n10443 ;
  assign n10445 = n10442 & ~n10443 ;
  assign n10446 = n10444 | n10445 ;
  assign n10447 = n9257 & ~n10446 ;
  assign n10448 = n10444 | n10447 ;
  assign n10449 = n10440 & n10448 ;
  assign n10450 = n10438 | n10449 ;
  assign n10451 = n10440 & ~n10445 ;
  assign n10452 = n10438 | n10451 ;
  assign n10453 = ( n10420 & n10450 ) | ( n10420 & n10452 ) | ( n10450 & n10452 ) ;
  assign n10454 = ~n7782 & n10453 ;
  assign n10455 = n7779 | n10454 ;
  assign n10456 = n5379 & ~n5495 ;
  assign n10457 = n5496 | n10456 ;
  assign n10458 = n5407 | n5475 ;
  assign n10459 = ~n5476 & n10458 ;
  assign n10460 = ~n3596 & n5069 ;
  assign n10461 = n3504 & n5070 ;
  assign n10462 = n10460 | n10461 ;
  assign n10463 = ~n3431 & n5083 ;
  assign n10464 = n10462 | n10463 ;
  assign n10465 = n5074 | n10464 ;
  assign n10466 = ( ~n4798 & n10464 ) | ( ~n4798 & n10465 ) | ( n10464 & n10465 ) ;
  assign n10467 = ~x17 & n10466 ;
  assign n10468 = x17 | n10467 ;
  assign n10469 = ( ~n10466 & n10467 ) | ( ~n10466 & n10468 ) | ( n10467 & n10468 ) ;
  assign n10470 = n10459 & n10469 ;
  assign n10471 = n10459 & ~n10470 ;
  assign n10472 = ~n10459 & n10469 ;
  assign n10473 = n10471 | n10472 ;
  assign n10474 = n5422 | n5446 ;
  assign n10475 = ~n5447 & n10474 ;
  assign n10476 = n3104 & n4546 ;
  assign n10477 = n1327 & n4548 ;
  assign n10478 = n10476 | n10477 ;
  assign n10479 = ~n1151 & n4551 ;
  assign n10480 = n10478 | n10479 ;
  assign n10481 = n4554 | n10480 ;
  assign n10482 = ( ~n4034 & n10480 ) | ( ~n4034 & n10481 ) | ( n10480 & n10481 ) ;
  assign n10483 = ~x23 & n10482 ;
  assign n10484 = x23 | n10483 ;
  assign n10485 = ( ~n10482 & n10483 ) | ( ~n10482 & n10484 ) | ( n10483 & n10484 ) ;
  assign n10486 = n10475 & n10485 ;
  assign n10487 = n10485 & ~n10486 ;
  assign n10488 = ( n10475 & ~n10486 ) | ( n10475 & n10487 ) | ( ~n10486 & n10487 ) ;
  assign n10489 = n3178 & n4546 ;
  assign n10490 = n3104 & n4548 ;
  assign n10491 = n10489 | n10490 ;
  assign n10492 = n1327 & n4551 ;
  assign n10493 = n10491 | n10492 ;
  assign n10494 = n4554 | n10493 ;
  assign n10495 = ( n4501 & n10493 ) | ( n4501 & n10494 ) | ( n10493 & n10494 ) ;
  assign n10496 = x23 & n10495 ;
  assign n10497 = x23 & ~n10496 ;
  assign n10498 = ( n10495 & ~n10496 ) | ( n10495 & n10497 ) | ( ~n10496 & n10497 ) ;
  assign n10499 = ( n5425 & ~n5435 ) | ( n5425 & n5445 ) | ( ~n5435 & n5445 ) ;
  assign n10500 = ( ~n5425 & n5435 ) | ( ~n5425 & n10499 ) | ( n5435 & n10499 ) ;
  assign n10501 = ( ~n5445 & n10499 ) | ( ~n5445 & n10500 ) | ( n10499 & n10500 ) ;
  assign n10502 = ( n7710 & n10498 ) | ( n7710 & n10501 ) | ( n10498 & n10501 ) ;
  assign n10503 = n10488 & n10502 ;
  assign n10504 = n10486 | n10503 ;
  assign n10505 = ~n1014 & n4781 ;
  assign n10506 = n3349 & n4776 ;
  assign n10507 = ~n3255 & n4778 ;
  assign n10508 = n10506 | n10507 ;
  assign n10509 = n10505 | n10508 ;
  assign n10510 = n4784 | n10509 ;
  assign n10511 = ( n4742 & n10509 ) | ( n4742 & n10510 ) | ( n10509 & n10510 ) ;
  assign n10512 = x20 & n10511 ;
  assign n10513 = x20 & ~n10512 ;
  assign n10514 = ( n10511 & ~n10512 ) | ( n10511 & n10513 ) | ( ~n10512 & n10513 ) ;
  assign n10515 = ( ~n5448 & n5458 ) | ( ~n5448 & n5460 ) | ( n5458 & n5460 ) ;
  assign n10516 = ( n5448 & ~n5460 ) | ( n5448 & n10515 ) | ( ~n5460 & n10515 ) ;
  assign n10517 = ( ~n5458 & n10515 ) | ( ~n5458 & n10516 ) | ( n10515 & n10516 ) ;
  assign n10518 = ( n10504 & n10514 ) | ( n10504 & n10517 ) | ( n10514 & n10517 ) ;
  assign n10519 = n778 & n5069 ;
  assign n10520 = ~n3596 & n5070 ;
  assign n10521 = n10519 | n10520 ;
  assign n10522 = n3504 & n5083 ;
  assign n10523 = n10521 | n10522 ;
  assign n10524 = n5074 | n10523 ;
  assign n10525 = ( ~n5040 & n10523 ) | ( ~n5040 & n10524 ) | ( n10523 & n10524 ) ;
  assign n10526 = ~x17 & n10525 ;
  assign n10527 = x17 | n10526 ;
  assign n10528 = ( ~n10525 & n10526 ) | ( ~n10525 & n10527 ) | ( n10526 & n10527 ) ;
  assign n10529 = ( ~n5461 & n5471 ) | ( ~n5461 & n5474 ) | ( n5471 & n5474 ) ;
  assign n10530 = ( n5461 & ~n5474 ) | ( n5461 & n10529 ) | ( ~n5474 & n10529 ) ;
  assign n10531 = ( ~n5471 & n10529 ) | ( ~n5471 & n10530 ) | ( n10529 & n10530 ) ;
  assign n10532 = ( n10518 & n10528 ) | ( n10518 & n10531 ) | ( n10528 & n10531 ) ;
  assign n10533 = n10473 & n10532 ;
  assign n10534 = ~n3634 & n7277 ;
  assign n10535 = ( n5384 & ~n5387 ) | ( n5384 & n10534 ) | ( ~n5387 & n10534 ) ;
  assign n10536 = n39 | n10535 ;
  assign n10537 = ( n3726 & n10535 ) | ( n3726 & n10536 ) | ( n10535 & n10536 ) ;
  assign n10538 = x14 & n10537 ;
  assign n10539 = x14 & ~n10538 ;
  assign n10540 = ( n10537 & ~n10538 ) | ( n10537 & n10539 ) | ( ~n10538 & n10539 ) ;
  assign n10541 = ( n10470 & n10533 ) | ( n10470 & n10540 ) | ( n10533 & n10540 ) ;
  assign n10542 = n10470 | n10540 ;
  assign n10543 = n10533 | n10542 ;
  assign n10544 = ~n10541 & n10543 ;
  assign n10545 = ( n5477 & n5487 ) | ( n5477 & ~n5490 ) | ( n5487 & ~n5490 ) ;
  assign n10546 = ( ~n5477 & n5490 ) | ( ~n5477 & n10545 ) | ( n5490 & n10545 ) ;
  assign n10547 = ( ~n5487 & n10545 ) | ( ~n5487 & n10546 ) | ( n10545 & n10546 ) ;
  assign n10548 = n10544 & n10547 ;
  assign n10549 = n10541 | n10548 ;
  assign n10550 = ( n5392 & ~n5491 ) | ( n5392 & n5494 ) | ( ~n5491 & n5494 ) ;
  assign n10551 = ( ~n5392 & n5491 ) | ( ~n5392 & n10550 ) | ( n5491 & n10550 ) ;
  assign n10552 = ( ~n5494 & n10550 ) | ( ~n5494 & n10551 ) | ( n10550 & n10551 ) ;
  assign n10553 = n10549 & n10552 ;
  assign n10554 = n10549 | n10552 ;
  assign n10555 = ~n10553 & n10554 ;
  assign n10556 = ~n3634 & n7280 ;
  assign n10557 = ~n672 & n7277 ;
  assign n10558 = n10556 | n10557 ;
  assign n10559 = ~n589 & n5384 ;
  assign n10560 = n10558 | n10559 ;
  assign n10561 = n39 | n10560 ;
  assign n10562 = ( ~n5092 & n10560 ) | ( ~n5092 & n10561 ) | ( n10560 & n10561 ) ;
  assign n10563 = ~x14 & n10562 ;
  assign n10564 = x14 | n10563 ;
  assign n10565 = ( ~n10562 & n10563 ) | ( ~n10562 & n10564 ) | ( n10563 & n10564 ) ;
  assign n10566 = n10488 | n10502 ;
  assign n10567 = ~n10503 & n10566 ;
  assign n10568 = n1233 & n4776 ;
  assign n10569 = n3349 & n4778 ;
  assign n10570 = n10568 | n10569 ;
  assign n10571 = ~n3255 & n4781 ;
  assign n10572 = n10570 | n10571 ;
  assign n10573 = n4784 | n10572 ;
  assign n10574 = ( ~n4470 & n10572 ) | ( ~n4470 & n10573 ) | ( n10572 & n10573 ) ;
  assign n10575 = ~x20 & n10574 ;
  assign n10576 = x20 | n10575 ;
  assign n10577 = ( ~n10574 & n10575 ) | ( ~n10574 & n10576 ) | ( n10575 & n10576 ) ;
  assign n10578 = n10567 & n10577 ;
  assign n10579 = n10567 | n10577 ;
  assign n10580 = ~n10578 & n10579 ;
  assign n10581 = ~n1151 & n4776 ;
  assign n10582 = n1233 & n4778 ;
  assign n10583 = n10581 | n10582 ;
  assign n10584 = n3349 & n4781 ;
  assign n10585 = n10583 | n10584 ;
  assign n10586 = n4784 | n10585 ;
  assign n10587 = ( n4518 & n10585 ) | ( n4518 & n10586 ) | ( n10585 & n10586 ) ;
  assign n10588 = x20 & n10587 ;
  assign n10589 = x20 & ~n10588 ;
  assign n10590 = ( n10587 & ~n10588 ) | ( n10587 & n10589 ) | ( ~n10588 & n10589 ) ;
  assign n10591 = ( ~n7710 & n10498 ) | ( ~n7710 & n10501 ) | ( n10498 & n10501 ) ;
  assign n10592 = ( n7710 & ~n10501 ) | ( n7710 & n10591 ) | ( ~n10501 & n10591 ) ;
  assign n10593 = ( ~n10498 & n10591 ) | ( ~n10498 & n10592 ) | ( n10591 & n10592 ) ;
  assign n10594 = ( n7713 & n10590 ) | ( n7713 & n10593 ) | ( n10590 & n10593 ) ;
  assign n10595 = n10580 & n10594 ;
  assign n10596 = n10578 | n10595 ;
  assign n10597 = n904 & n5069 ;
  assign n10598 = n778 & n5070 ;
  assign n10599 = n10597 | n10598 ;
  assign n10600 = ~n3596 & n5083 ;
  assign n10601 = n10599 | n10600 ;
  assign n10602 = n5074 | n10601 ;
  assign n10603 = ( ~n4649 & n10601 ) | ( ~n4649 & n10602 ) | ( n10601 & n10602 ) ;
  assign n10604 = ~x17 & n10603 ;
  assign n10605 = x17 | n10604 ;
  assign n10606 = ( ~n10603 & n10604 ) | ( ~n10603 & n10605 ) | ( n10604 & n10605 ) ;
  assign n10607 = ( ~n10504 & n10514 ) | ( ~n10504 & n10517 ) | ( n10514 & n10517 ) ;
  assign n10608 = ( n10504 & ~n10517 ) | ( n10504 & n10607 ) | ( ~n10517 & n10607 ) ;
  assign n10609 = ( ~n10514 & n10607 ) | ( ~n10514 & n10608 ) | ( n10607 & n10608 ) ;
  assign n10610 = ( n10596 & n10606 ) | ( n10596 & n10609 ) | ( n10606 & n10609 ) ;
  assign n10611 = ~n3431 & n5384 ;
  assign n10612 = ~n589 & n7277 ;
  assign n10613 = n10611 | n10612 ;
  assign n10614 = ~n672 & n7280 ;
  assign n10615 = n10613 | n10614 ;
  assign n10616 = n39 | n10615 ;
  assign n10617 = ( ~n5353 & n10615 ) | ( ~n5353 & n10616 ) | ( n10615 & n10616 ) ;
  assign n10618 = ~x14 & n10617 ;
  assign n10619 = x14 | n10618 ;
  assign n10620 = ( ~n10617 & n10618 ) | ( ~n10617 & n10619 ) | ( n10618 & n10619 ) ;
  assign n10621 = ( ~n10518 & n10528 ) | ( ~n10518 & n10531 ) | ( n10528 & n10531 ) ;
  assign n10622 = ( n10518 & ~n10531 ) | ( n10518 & n10621 ) | ( ~n10531 & n10621 ) ;
  assign n10623 = ( ~n10528 & n10621 ) | ( ~n10528 & n10622 ) | ( n10621 & n10622 ) ;
  assign n10624 = ( n10610 & n10620 ) | ( n10610 & n10623 ) | ( n10620 & n10623 ) ;
  assign n10625 = n10565 & n10624 ;
  assign n10626 = n10624 & ~n10625 ;
  assign n10627 = n10473 | n10532 ;
  assign n10628 = ~n10533 & n10627 ;
  assign n10629 = n10565 & ~n10624 ;
  assign n10630 = ( n10626 & n10628 ) | ( n10626 & n10629 ) | ( n10628 & n10629 ) ;
  assign n10631 = n10544 | n10547 ;
  assign n10632 = ~n10548 & n10631 ;
  assign n10633 = ( n10625 & n10630 ) | ( n10625 & n10632 ) | ( n10630 & n10632 ) ;
  assign n10634 = n10625 | n10632 ;
  assign n10635 = n10630 | n10634 ;
  assign n10636 = ~n10633 & n10635 ;
  assign n10637 = n10628 | n10629 ;
  assign n10638 = n10626 | n10637 ;
  assign n10639 = ~n10630 & n10638 ;
  assign n10640 = n7300 | n7308 ;
  assign n10641 = ~n3634 & n10640 ;
  assign n10642 = n672 & n7300 ;
  assign n10643 = ( ~n672 & n10641 ) | ( ~n672 & n10642 ) | ( n10641 & n10642 ) ;
  assign n10644 = ( ~n3619 & n10641 ) | ( ~n3619 & n10643 ) | ( n10641 & n10643 ) ;
  assign n10645 = ~x11 & n10644 ;
  assign n10646 = x11 | n10645 ;
  assign n10647 = ( ~n10644 & n10645 ) | ( ~n10644 & n10646 ) | ( n10645 & n10646 ) ;
  assign n10648 = n10580 | n10594 ;
  assign n10649 = ~n10595 & n10648 ;
  assign n10650 = ~n1014 & n5069 ;
  assign n10651 = n904 & n5070 ;
  assign n10652 = n10650 | n10651 ;
  assign n10653 = n778 & n5083 ;
  assign n10654 = n10652 | n10653 ;
  assign n10655 = n5074 | n10654 ;
  assign n10656 = ( ~n4535 & n10654 ) | ( ~n4535 & n10655 ) | ( n10654 & n10655 ) ;
  assign n10657 = ~x17 & n10656 ;
  assign n10658 = x17 | n10657 ;
  assign n10659 = ( ~n10656 & n10657 ) | ( ~n10656 & n10658 ) | ( n10657 & n10658 ) ;
  assign n10660 = n10649 & n10659 ;
  assign n10661 = n10659 & ~n10660 ;
  assign n10662 = ( n10649 & ~n10660 ) | ( n10649 & n10661 ) | ( ~n10660 & n10661 ) ;
  assign n10663 = n7715 | n7728 ;
  assign n10664 = ~n1014 & n5070 ;
  assign n10665 = ~n3255 & n5069 ;
  assign n10666 = n10664 | n10665 ;
  assign n10667 = n904 & n5083 ;
  assign n10668 = n10666 | n10667 ;
  assign n10669 = n5074 | n10668 ;
  assign n10670 = ( n4632 & n10668 ) | ( n4632 & n10669 ) | ( n10668 & n10669 ) ;
  assign n10671 = x17 & n10670 ;
  assign n10672 = x17 & ~n10671 ;
  assign n10673 = ( n10670 & ~n10671 ) | ( n10670 & n10672 ) | ( ~n10671 & n10672 ) ;
  assign n10674 = ( ~n7713 & n10590 ) | ( ~n7713 & n10593 ) | ( n10590 & n10593 ) ;
  assign n10675 = ( n7713 & ~n10593 ) | ( n7713 & n10674 ) | ( ~n10593 & n10674 ) ;
  assign n10676 = ( ~n10590 & n10674 ) | ( ~n10590 & n10675 ) | ( n10674 & n10675 ) ;
  assign n10677 = ( n10663 & n10673 ) | ( n10663 & n10676 ) | ( n10673 & n10676 ) ;
  assign n10678 = n10662 & n10677 ;
  assign n10679 = n10660 | n10678 ;
  assign n10680 = n3504 & n5384 ;
  assign n10681 = ~n3431 & n7277 ;
  assign n10682 = n10680 | n10681 ;
  assign n10683 = ~n589 & n7280 ;
  assign n10684 = n10682 | n10683 ;
  assign n10685 = n39 | n10684 ;
  assign n10686 = ( n4765 & n10684 ) | ( n4765 & n10685 ) | ( n10684 & n10685 ) ;
  assign n10687 = x14 & n10686 ;
  assign n10688 = x14 & ~n10687 ;
  assign n10689 = ( n10686 & ~n10687 ) | ( n10686 & n10688 ) | ( ~n10687 & n10688 ) ;
  assign n10690 = ( n10596 & n10606 ) | ( n10596 & ~n10609 ) | ( n10606 & ~n10609 ) ;
  assign n10691 = ( ~n10596 & n10609 ) | ( ~n10596 & n10690 ) | ( n10609 & n10690 ) ;
  assign n10692 = ( ~n10606 & n10690 ) | ( ~n10606 & n10691 ) | ( n10690 & n10691 ) ;
  assign n10693 = ( n10679 & n10689 ) | ( n10679 & n10692 ) | ( n10689 & n10692 ) ;
  assign n10694 = ( ~n10610 & n10620 ) | ( ~n10610 & n10623 ) | ( n10620 & n10623 ) ;
  assign n10695 = ( n10610 & ~n10623 ) | ( n10610 & n10694 ) | ( ~n10623 & n10694 ) ;
  assign n10696 = ( ~n10620 & n10694 ) | ( ~n10620 & n10695 ) | ( n10694 & n10695 ) ;
  assign n10697 = ( n10647 & n10693 ) | ( n10647 & n10696 ) | ( n10693 & n10696 ) ;
  assign n10698 = n10639 & n10697 ;
  assign n10699 = n10639 | n10697 ;
  assign n10700 = ~n10698 & n10699 ;
  assign n10701 = n10662 | n10677 ;
  assign n10702 = ~n10678 & n10701 ;
  assign n10703 = ~n3596 & n5384 ;
  assign n10704 = n3504 & n7277 ;
  assign n10705 = n10703 | n10704 ;
  assign n10706 = ~n3431 & n7280 ;
  assign n10707 = n10705 | n10706 ;
  assign n10708 = n39 | n10707 ;
  assign n10709 = ( ~n4798 & n10707 ) | ( ~n4798 & n10708 ) | ( n10707 & n10708 ) ;
  assign n10710 = ~x14 & n10709 ;
  assign n10711 = x14 | n10710 ;
  assign n10712 = ( ~n10709 & n10710 ) | ( ~n10709 & n10711 ) | ( n10710 & n10711 ) ;
  assign n10713 = n10702 & n10712 ;
  assign n10714 = ~n7735 & n7745 ;
  assign n10715 = n7734 | n10714 ;
  assign n10716 = ( ~n10663 & n10673 ) | ( ~n10663 & n10676 ) | ( n10673 & n10676 ) ;
  assign n10717 = ( n10663 & ~n10676 ) | ( n10663 & n10716 ) | ( ~n10676 & n10716 ) ;
  assign n10718 = ( ~n10673 & n10716 ) | ( ~n10673 & n10717 ) | ( n10716 & n10717 ) ;
  assign n10719 = n10715 & n10718 ;
  assign n10720 = n10715 | n10718 ;
  assign n10721 = ~n10719 & n10720 ;
  assign n10722 = n778 & n5384 ;
  assign n10723 = ~n3596 & n7277 ;
  assign n10724 = n10722 | n10723 ;
  assign n10725 = n3504 & n7280 ;
  assign n10726 = n10724 | n10725 ;
  assign n10727 = n39 | n10726 ;
  assign n10728 = ( ~n5040 & n10726 ) | ( ~n5040 & n10727 ) | ( n10726 & n10727 ) ;
  assign n10729 = ~x14 & n10728 ;
  assign n10730 = x14 | n10729 ;
  assign n10731 = ( ~n10728 & n10729 ) | ( ~n10728 & n10730 ) | ( n10729 & n10730 ) ;
  assign n10732 = n10721 & n10731 ;
  assign n10733 = n10719 | n10732 ;
  assign n10734 = n10702 & ~n10713 ;
  assign n10735 = ~n10702 & n10712 ;
  assign n10736 = n10734 | n10735 ;
  assign n10737 = n10733 & n10736 ;
  assign n10738 = ~n3634 & n7302 ;
  assign n10739 = ( n7300 & ~n10642 ) | ( n7300 & n10738 ) | ( ~n10642 & n10738 ) ;
  assign n10740 = n7308 | n10739 ;
  assign n10741 = ( n3726 & n10739 ) | ( n3726 & n10740 ) | ( n10739 & n10740 ) ;
  assign n10742 = x11 & n10741 ;
  assign n10743 = x11 & ~n10742 ;
  assign n10744 = ( n10741 & ~n10742 ) | ( n10741 & n10743 ) | ( ~n10742 & n10743 ) ;
  assign n10745 = ( n10713 & n10737 ) | ( n10713 & n10744 ) | ( n10737 & n10744 ) ;
  assign n10746 = n10713 | n10744 ;
  assign n10747 = n10737 | n10746 ;
  assign n10748 = ~n10745 & n10747 ;
  assign n10749 = ( n10679 & n10689 ) | ( n10679 & ~n10692 ) | ( n10689 & ~n10692 ) ;
  assign n10750 = ( ~n10679 & n10692 ) | ( ~n10679 & n10749 ) | ( n10692 & n10749 ) ;
  assign n10751 = ( ~n10689 & n10749 ) | ( ~n10689 & n10750 ) | ( n10749 & n10750 ) ;
  assign n10752 = n10748 & n10751 ;
  assign n10753 = n10745 | n10752 ;
  assign n10754 = ( n10647 & ~n10693 ) | ( n10647 & n10696 ) | ( ~n10693 & n10696 ) ;
  assign n10755 = ( ~n10647 & n10693 ) | ( ~n10647 & n10754 ) | ( n10693 & n10754 ) ;
  assign n10756 = ( ~n10696 & n10754 ) | ( ~n10696 & n10755 ) | ( n10754 & n10755 ) ;
  assign n10757 = n10753 & n10756 ;
  assign n10758 = n10753 | n10756 ;
  assign n10759 = ~n10757 & n10758 ;
  assign n10760 = n10748 | n10751 ;
  assign n10761 = ~n10752 & n10760 ;
  assign n10762 = ~n3634 & n7305 ;
  assign n10763 = ~n672 & n7302 ;
  assign n10764 = n10762 | n10763 ;
  assign n10765 = ~n589 & n7300 ;
  assign n10766 = n10764 | n10765 ;
  assign n10767 = n7308 | n10766 ;
  assign n10768 = ( ~n5092 & n10766 ) | ( ~n5092 & n10767 ) | ( n10766 & n10767 ) ;
  assign n10769 = ~x11 & n10768 ;
  assign n10770 = x11 | n10769 ;
  assign n10771 = ( ~n10768 & n10769 ) | ( ~n10768 & n10770 ) | ( n10769 & n10770 ) ;
  assign n10772 = n10721 & ~n10732 ;
  assign n10773 = ~n10721 & n10731 ;
  assign n10774 = ( n7683 & n7758 ) | ( n7683 & n7761 ) | ( n7758 & n7761 ) ;
  assign n10775 = n10773 | n10774 ;
  assign n10776 = n10772 | n10775 ;
  assign n10777 = ( n10772 & n10773 ) | ( n10772 & n10774 ) | ( n10773 & n10774 ) ;
  assign n10778 = ~n3431 & n7300 ;
  assign n10779 = ~n589 & n7302 ;
  assign n10780 = n10778 | n10779 ;
  assign n10781 = ~n672 & n7305 ;
  assign n10782 = n10780 | n10781 ;
  assign n10783 = n7308 | n10782 ;
  assign n10784 = ( ~n5353 & n10782 ) | ( ~n5353 & n10783 ) | ( n10782 & n10783 ) ;
  assign n10785 = ~x11 & n10784 ;
  assign n10786 = x11 | n10785 ;
  assign n10787 = ( ~n10784 & n10785 ) | ( ~n10784 & n10786 ) | ( n10785 & n10786 ) ;
  assign n10788 = ( n10776 & n10777 ) | ( n10776 & n10787 ) | ( n10777 & n10787 ) ;
  assign n10789 = n10733 & ~n10737 ;
  assign n10790 = n10736 & ~n10737 ;
  assign n10791 = n10789 | n10790 ;
  assign n10792 = ( n10771 & n10788 ) | ( n10771 & n10791 ) | ( n10788 & n10791 ) ;
  assign n10793 = n10761 & n10792 ;
  assign n10794 = n10761 | n10792 ;
  assign n10795 = ~n10793 & n10794 ;
  assign n10796 = n5512 | n5515 ;
  assign n10797 = ~n3634 & n10796 ;
  assign n10798 = ( ~n672 & n7672 ) | ( ~n672 & n10797 ) | ( n7672 & n10797 ) ;
  assign n10799 = ( ~n3619 & n10797 ) | ( ~n3619 & n10798 ) | ( n10797 & n10798 ) ;
  assign n10800 = ~x8 & n10799 ;
  assign n10801 = x8 | n10800 ;
  assign n10802 = ( ~n10799 & n10800 ) | ( ~n10799 & n10801 ) | ( n10800 & n10801 ) ;
  assign n10803 = ( n7762 & n7772 ) | ( n7762 & n7775 ) | ( n7772 & n7775 ) ;
  assign n10804 = n10776 & ~n10777 ;
  assign n10805 = ~n10787 & n10804 ;
  assign n10806 = n10787 | n10805 ;
  assign n10807 = ( ~n10804 & n10805 ) | ( ~n10804 & n10806 ) | ( n10805 & n10806 ) ;
  assign n10808 = ( n10802 & n10803 ) | ( n10802 & n10807 ) | ( n10803 & n10807 ) ;
  assign n10809 = ( n10771 & ~n10788 ) | ( n10771 & n10791 ) | ( ~n10788 & n10791 ) ;
  assign n10810 = ( ~n10771 & n10788 ) | ( ~n10771 & n10809 ) | ( n10788 & n10809 ) ;
  assign n10811 = ( ~n10791 & n10809 ) | ( ~n10791 & n10810 ) | ( n10809 & n10810 ) ;
  assign n10812 = n10808 & n10811 ;
  assign n10813 = n7680 | n7776 ;
  assign n10814 = ( n10802 & ~n10803 ) | ( n10802 & n10807 ) | ( ~n10803 & n10807 ) ;
  assign n10815 = ( ~n10802 & n10803 ) | ( ~n10802 & n10814 ) | ( n10803 & n10814 ) ;
  assign n10816 = ( ~n10807 & n10814 ) | ( ~n10807 & n10815 ) | ( n10814 & n10815 ) ;
  assign n10817 = n10813 | n10816 ;
  assign n10818 = n10808 | n10811 ;
  assign n10819 = ~n10812 & n10818 ;
  assign n10820 = n10817 & n10819 ;
  assign n10821 = n10812 | n10820 ;
  assign n10822 = n10795 & n10821 ;
  assign n10823 = n10793 | n10822 ;
  assign n10824 = n10759 & n10823 ;
  assign n10825 = n10757 | n10824 ;
  assign n10826 = n10700 & n10825 ;
  assign n10827 = n10698 | n10826 ;
  assign n10828 = n10636 & n10827 ;
  assign n10829 = n10633 | n10828 ;
  assign n10830 = n10555 & n10829 ;
  assign n10831 = n10553 | n10830 ;
  assign n10832 = ~n10457 & n10831 ;
  assign n10833 = n10813 & n10816 ;
  assign n10834 = n10819 & n10833 ;
  assign n10835 = n10812 | n10834 ;
  assign n10836 = n10795 & n10835 ;
  assign n10837 = n10793 | n10836 ;
  assign n10838 = n10759 & n10837 ;
  assign n10839 = n10757 | n10838 ;
  assign n10840 = n10700 & n10839 ;
  assign n10841 = n10698 | n10840 ;
  assign n10842 = n10636 & n10841 ;
  assign n10843 = n10633 | n10842 ;
  assign n10844 = n10555 & n10843 ;
  assign n10845 = n10553 | n10844 ;
  assign n10846 = ~n10457 & n10845 ;
  assign n10847 = ( n10455 & n10832 ) | ( n10455 & n10846 ) | ( n10832 & n10846 ) ;
  assign n10848 = n5496 | n10847 ;
  assign n10849 = n5377 & n10848 ;
  assign n10850 = n3463 | n4929 ;
  assign n10851 = n627 | n2739 ;
  assign n10852 = n10850 | n10851 ;
  assign n10853 = n983 & ~n10852 ;
  assign n10854 = n892 | n1170 ;
  assign n10855 = n621 | n1034 ;
  assign n10856 = n10854 | n10855 ;
  assign n10857 = n539 | n669 ;
  assign n10858 = n252 | n10857 ;
  assign n10859 = n300 | n10858 ;
  assign n10860 = n10856 | n10859 ;
  assign n10861 = ( n90 & n359 ) | ( n90 & ~n3115 ) | ( n359 & ~n3115 ) ;
  assign n10862 = n3115 | n10861 ;
  assign n10863 = n10860 | n10862 ;
  assign n10864 = n10853 & ~n10863 ;
  assign n10865 = n1363 | n4337 ;
  assign n10866 = n491 | n960 ;
  assign n10867 = n166 | n10866 ;
  assign n10868 = n10865 | n10867 ;
  assign n10869 = n352 | n2867 ;
  assign n10870 = n244 | n10869 ;
  assign n10871 = n633 | n10870 ;
  assign n10872 = n10868 | n10871 ;
  assign n10873 = n321 | n583 ;
  assign n10874 = n199 | n10873 ;
  assign n10875 = n204 | n10874 ;
  assign n10876 = n181 | n10875 ;
  assign n10877 = n132 | n10876 ;
  assign n10878 = n10872 | n10877 ;
  assign n10879 = n5703 | n10878 ;
  assign n10880 = n10864 & ~n10879 ;
  assign n10881 = ~n4683 & n10880 ;
  assign n10882 = n130 | n641 ;
  assign n10883 = n629 | n10882 ;
  assign n10884 = n355 | n10883 ;
  assign n10885 = n591 | n10884 ;
  assign n10886 = n580 | n10885 ;
  assign n10887 = n134 | n10886 ;
  assign n10888 = n222 | n10887 ;
  assign n10889 = n403 | n10888 ;
  assign n10890 = n10881 & ~n10889 ;
  assign n10891 = n3703 & ~n10890 ;
  assign n10892 = ~n3703 & n10890 ;
  assign n10893 = n3504 & n3639 ;
  assign n10894 = ~n3431 & n3727 ;
  assign n10895 = n10893 | n10894 ;
  assign n10896 = ~n589 & n3744 ;
  assign n10897 = n10895 | n10896 ;
  assign n10898 = n81 | n2966 ;
  assign n10899 = n445 | n618 ;
  assign n10900 = n92 | n10899 ;
  assign n10901 = n1778 | n2199 ;
  assign n10902 = ( ~n5194 & n10900 ) | ( ~n5194 & n10901 ) | ( n10900 & n10901 ) ;
  assign n10903 = n5194 | n10902 ;
  assign n10904 = n4946 | n10903 ;
  assign n10905 = n4940 | n10904 ;
  assign n10906 = n2400 | n10905 ;
  assign n10907 = n10898 | n10906 ;
  assign n10908 = n144 | n555 ;
  assign n10909 = n242 | n531 ;
  assign n10910 = n283 | n513 ;
  assign n10911 = n10909 | n10910 ;
  assign n10912 = n334 | n450 ;
  assign n10913 = ( ~n2383 & n10911 ) | ( ~n2383 & n10912 ) | ( n10911 & n10912 ) ;
  assign n10914 = n2383 | n10913 ;
  assign n10915 = n10908 | n10914 ;
  assign n10916 = n1079 | n10915 ;
  assign n10917 = n3873 | n10916 ;
  assign n10918 = n635 | n10917 ;
  assign n10919 = n718 | n10918 ;
  assign n10920 = n337 | n10919 ;
  assign n10921 = n10907 | n10920 ;
  assign n10922 = n172 | n357 ;
  assign n10923 = n661 | n10922 ;
  assign n10924 = n10921 | n10923 ;
  assign n10925 = n292 | n610 ;
  assign n10926 = n2219 | n10925 ;
  assign n10927 = n449 | n10926 ;
  assign n10928 = n732 | n3869 ;
  assign n10929 = n10927 | n10928 ;
  assign n10930 = n282 | n834 ;
  assign n10931 = n452 | n10930 ;
  assign n10932 = n143 | n10931 ;
  assign n10933 = n10929 | n10932 ;
  assign n10934 = n227 | n10933 ;
  assign n10935 = n307 | n621 ;
  assign n10936 = n140 | n10935 ;
  assign n10937 = n1204 | n5218 ;
  assign n10938 = n10936 | n10937 ;
  assign n10939 = n515 | n10938 ;
  assign n10940 = n5249 | n10939 ;
  assign n10941 = n760 | n1443 ;
  assign n10942 = n959 | n10941 ;
  assign n10943 = n2922 | n10942 ;
  assign n10944 = n475 | n10943 ;
  assign n10945 = n10940 | n10944 ;
  assign n10946 = n484 | n520 ;
  assign n10947 = n358 | n10946 ;
  assign n10948 = n379 | n10947 ;
  assign n10949 = n607 | n10948 ;
  assign n10950 = n570 | n10949 ;
  assign n10951 = n128 | n10950 ;
  assign n10952 = n10945 | n10951 ;
  assign n10953 = n10934 | n10952 ;
  assign n10954 = n139 | n165 ;
  assign n10955 = n648 | n10954 ;
  assign n10956 = n206 | n10955 ;
  assign n10957 = n1837 | n4225 ;
  assign n10958 = n5232 | n10957 ;
  assign n10959 = ( ~n2753 & n10956 ) | ( ~n2753 & n10958 ) | ( n10956 & n10958 ) ;
  assign n10960 = n2753 | n10959 ;
  assign n10961 = n10953 | n10960 ;
  assign n10962 = n731 | n911 ;
  assign n10963 = n2362 | n10962 ;
  assign n10964 = n697 | n10963 ;
  assign n10965 = n3204 | n10964 ;
  assign n10966 = n618 | n10965 ;
  assign n10967 = n349 | n10966 ;
  assign n10968 = n198 | n10967 ;
  assign n10969 = n190 | n10968 ;
  assign n10970 = n10961 | n10969 ;
  assign n10971 = ( x26 & ~n10924 ) | ( x26 & n10970 ) | ( ~n10924 & n10970 ) ;
  assign n10972 = ( ~x26 & n10924 ) | ( ~x26 & n10971 ) | ( n10924 & n10971 ) ;
  assign n10973 = ( n10890 & n10897 ) | ( n10890 & n10972 ) | ( n10897 & n10972 ) ;
  assign n10974 = ~n10891 & n10973 ;
  assign n10975 = ~n10892 & n10974 ;
  assign n10976 = n3636 | n10897 ;
  assign n10977 = ( n10890 & n10972 ) | ( n10890 & n10976 ) | ( n10972 & n10976 ) ;
  assign n10978 = ~n10891 & n10977 ;
  assign n10979 = ~n10892 & n10978 ;
  assign n10980 = ( n4765 & n10975 ) | ( n4765 & n10979 ) | ( n10975 & n10979 ) ;
  assign n10981 = n10891 | n10980 ;
  assign n10982 = ( ~n3703 & n3720 ) | ( ~n3703 & n3721 ) | ( n3720 & n3721 ) ;
  assign n10983 = ( ~x29 & n3721 ) | ( ~x29 & n10982 ) | ( n3721 & n10982 ) ;
  assign n10984 = n10981 & n10983 ;
  assign n10985 = n10981 | n10983 ;
  assign n10986 = ~n10984 & n10985 ;
  assign n10987 = ~n3634 & n3744 ;
  assign n10988 = ~n672 & n3727 ;
  assign n10989 = n10987 | n10988 ;
  assign n10990 = ~n589 & n3639 ;
  assign n10991 = n10989 | n10990 ;
  assign n10992 = n3636 | n10991 ;
  assign n10993 = ( ~n5092 & n10991 ) | ( ~n5092 & n10992 ) | ( n10991 & n10992 ) ;
  assign n10994 = n10986 & n10993 ;
  assign n10995 = n10984 | n10994 ;
  assign n10996 = ~n3736 & n10995 ;
  assign n10997 = n3736 & ~n10995 ;
  assign n10998 = n10996 | n10997 ;
  assign n10999 = n10986 | n10993 ;
  assign n11000 = ~n10994 & n10999 ;
  assign n11001 = ~n3431 & n3639 ;
  assign n11002 = ~n589 & n3727 ;
  assign n11003 = n11001 | n11002 ;
  assign n11004 = ~n672 & n3744 ;
  assign n11005 = n11003 | n11004 ;
  assign n11006 = n3636 | n11005 ;
  assign n11007 = ( ~n5353 & n11005 ) | ( ~n5353 & n11006 ) | ( n11005 & n11006 ) ;
  assign n11008 = n4043 | n4051 ;
  assign n11009 = ~n3634 & n11008 ;
  assign n11010 = n672 & n4043 ;
  assign n11011 = ( ~n672 & n11009 ) | ( ~n672 & n11010 ) | ( n11009 & n11010 ) ;
  assign n11012 = ( ~n3619 & n11009 ) | ( ~n3619 & n11011 ) | ( n11009 & n11011 ) ;
  assign n11013 = ~x29 & n11012 ;
  assign n11014 = x29 | n11013 ;
  assign n11015 = ( ~n11012 & n11013 ) | ( ~n11012 & n11014 ) | ( n11013 & n11014 ) ;
  assign n11016 = n11007 & n11015 ;
  assign n11017 = ( n4765 & n10973 ) | ( n4765 & n10977 ) | ( n10973 & n10977 ) ;
  assign n11018 = ~n10980 & n11017 ;
  assign n11019 = n10892 | n10981 ;
  assign n11020 = ~n11018 & n11019 ;
  assign n11021 = ( ~n11007 & n11015 ) | ( ~n11007 & n11020 ) | ( n11015 & n11020 ) ;
  assign n11022 = ( n11007 & ~n11015 ) | ( n11007 & n11021 ) | ( ~n11015 & n11021 ) ;
  assign n11023 = ~n11020 & n11022 ;
  assign n11024 = ( ~n11020 & n11021 ) | ( ~n11020 & n11023 ) | ( n11021 & n11023 ) ;
  assign n11025 = ( n11000 & n11016 ) | ( n11000 & n11024 ) | ( n11016 & n11024 ) ;
  assign n11026 = n11000 | n11016 ;
  assign n11027 = n11024 | n11026 ;
  assign n11028 = ~n11025 & n11027 ;
  assign n11029 = ( ~n11020 & n11021 ) | ( ~n11020 & n11022 ) | ( n11021 & n11022 ) ;
  assign n11030 = ~n3634 & n4045 ;
  assign n11031 = ( n4043 & ~n11010 ) | ( n4043 & n11030 ) | ( ~n11010 & n11030 ) ;
  assign n11032 = n4051 | n11031 ;
  assign n11033 = ( n3726 & n11031 ) | ( n3726 & n11032 ) | ( n11031 & n11032 ) ;
  assign n11034 = x29 & n11033 ;
  assign n11035 = x29 & ~n11034 ;
  assign n11036 = ( n11033 & ~n11034 ) | ( n11033 & n11035 ) | ( ~n11034 & n11035 ) ;
  assign n11037 = ~n3596 & n3639 ;
  assign n11038 = n3504 & n3727 ;
  assign n11039 = n11037 | n11038 ;
  assign n11040 = ~n3431 & n3744 ;
  assign n11041 = n11039 | n11040 ;
  assign n11042 = n3636 | n11041 ;
  assign n11043 = ( ~n4798 & n11041 ) | ( ~n4798 & n11042 ) | ( n11041 & n11042 ) ;
  assign n11044 = n3326 | n4942 ;
  assign n11045 = n219 | n1791 ;
  assign n11046 = n446 | n11045 ;
  assign n11047 = n11044 | n11046 ;
  assign n11048 = n1442 | n2393 ;
  assign n11049 = n416 | n11048 ;
  assign n11050 = n52 | n11049 ;
  assign n11051 = n11047 | n11050 ;
  assign n11052 = n560 | n11051 ;
  assign n11053 = n258 | n296 ;
  assign n11054 = n55 | n11053 ;
  assign n11055 = n2959 | n11054 ;
  assign n11056 = n245 | n391 ;
  assign n11057 = n273 | n539 ;
  assign n11058 = n11056 | n11057 ;
  assign n11059 = n139 | n155 ;
  assign n11060 = n11058 | n11059 ;
  assign n11061 = n11055 | n11060 ;
  assign n11062 = n3880 | n11061 ;
  assign n11063 = n11052 | n11062 ;
  assign n11064 = ( n93 & n639 ) | ( n93 & ~n5244 ) | ( n639 & ~n5244 ) ;
  assign n11065 = n5244 | n11064 ;
  assign n11066 = n249 | n11065 ;
  assign n11067 = n321 | n11066 ;
  assign n11068 = n358 | n11067 ;
  assign n11069 = n11063 | n11068 ;
  assign n11070 = n161 | n3261 ;
  assign n11071 = n133 | n11070 ;
  assign n11072 = n649 | n11071 ;
  assign n11073 = n280 | n327 ;
  assign n11074 = n174 | n11073 ;
  assign n11075 = n598 | n5218 ;
  assign n11076 = n11074 | n11075 ;
  assign n11077 = n11072 | n11076 ;
  assign n11078 = n11069 | n11077 ;
  assign n11079 = n320 | n629 ;
  assign n11080 = n193 | n11079 ;
  assign n11081 = n313 | n11080 ;
  assign n11082 = n144 | n11081 ;
  assign n11083 = n209 | n11082 ;
  assign n11084 = n509 | n11083 ;
  assign n11085 = n1175 | n11084 ;
  assign n11086 = n306 | n434 ;
  assign n11087 = ( n120 & ~n1594 ) | ( n120 & n11086 ) | ( ~n1594 & n11086 ) ;
  assign n11088 = n1594 | n11087 ;
  assign n11089 = n650 | n11088 ;
  assign n11090 = n11085 | n11089 ;
  assign n11091 = n756 | n11090 ;
  assign n11092 = n11078 | n11091 ;
  assign n11093 = n568 | n1659 ;
  assign n11094 = n862 | n11093 ;
  assign n11095 = n654 | n11094 ;
  assign n11096 = n608 | n11095 ;
  assign n11097 = n610 | n11096 ;
  assign n11098 = n83 | n11097 ;
  assign n11099 = n11092 | n11098 ;
  assign n11100 = ~n10924 & n11099 ;
  assign n11101 = n10924 & ~n11099 ;
  assign n11102 = n778 & n3639 ;
  assign n11103 = ~n3596 & n3727 ;
  assign n11104 = n11102 | n11103 ;
  assign n11105 = n3504 & n3744 ;
  assign n11106 = n11104 | n11105 ;
  assign n11107 = n3636 | n11106 ;
  assign n11108 = ~n11100 & n11107 ;
  assign n11109 = ~n11101 & n11108 ;
  assign n11110 = ~n11100 & n11106 ;
  assign n11111 = ~n11101 & n11110 ;
  assign n11112 = ( ~n5040 & n11109 ) | ( ~n5040 & n11111 ) | ( n11109 & n11111 ) ;
  assign n11113 = n11100 | n11112 ;
  assign n11114 = ( ~n10970 & n10971 ) | ( ~n10970 & n10972 ) | ( n10971 & n10972 ) ;
  assign n11115 = ( ~n11043 & n11113 ) | ( ~n11043 & n11114 ) | ( n11113 & n11114 ) ;
  assign n11116 = ( n11043 & ~n11113 ) | ( n11043 & n11115 ) | ( ~n11113 & n11115 ) ;
  assign n11117 = ( ~n11114 & n11115 ) | ( ~n11114 & n11116 ) | ( n11115 & n11116 ) ;
  assign n11118 = ( n11043 & n11113 ) | ( n11043 & n11117 ) | ( n11113 & n11117 ) ;
  assign n11119 = ( n4765 & n10897 ) | ( n4765 & n10976 ) | ( n10897 & n10976 ) ;
  assign n11120 = ( n10890 & ~n10972 ) | ( n10890 & n11119 ) | ( ~n10972 & n11119 ) ;
  assign n11121 = ( ~n10890 & n10972 ) | ( ~n10890 & n11120 ) | ( n10972 & n11120 ) ;
  assign n11122 = ( ~n11119 & n11120 ) | ( ~n11119 & n11121 ) | ( n11120 & n11121 ) ;
  assign n11123 = ( n11036 & n11118 ) | ( n11036 & n11122 ) | ( n11118 & n11122 ) ;
  assign n11124 = ~n11029 & n11123 ;
  assign n11125 = n11029 & ~n11123 ;
  assign n11126 = n11124 | n11125 ;
  assign n11127 = ( ~n5040 & n11106 ) | ( ~n5040 & n11107 ) | ( n11106 & n11107 ) ;
  assign n11128 = ~n11112 & n11127 ;
  assign n11130 = n4155 | n4231 ;
  assign n11131 = n4151 | n11130 ;
  assign n11132 = n429 | n519 ;
  assign n11133 = n831 | n11132 ;
  assign n11134 = n273 | n279 ;
  assign n11135 = n314 | n11134 ;
  assign n11136 = n11133 | n11135 ;
  assign n11137 = n300 | n595 ;
  assign n11138 = n218 | n11137 ;
  assign n11139 = n11136 | n11138 ;
  assign n11140 = n2506 | n11139 ;
  assign n11141 = n2221 | n11140 ;
  assign n11142 = n11131 | n11141 ;
  assign n11143 = n479 | n5612 ;
  assign n11144 = n578 | n11143 ;
  assign n11145 = n400 | n11144 ;
  assign n11146 = n199 | n11145 ;
  assign n11147 = n602 | n11146 ;
  assign n11148 = n11142 | n11147 ;
  assign n11149 = n134 | n500 ;
  assign n11150 = n77 | n449 ;
  assign n11151 = n11149 | n11150 ;
  assign n11152 = n646 | n11151 ;
  assign n11153 = n2301 | n4876 ;
  assign n11154 = n1118 | n11153 ;
  assign n11155 = n11152 | n11154 ;
  assign n11156 = n1484 | n11155 ;
  assign n11157 = n432 | n488 ;
  assign n11158 = n253 | n276 ;
  assign n11159 = n11157 | n11158 ;
  assign n11160 = n346 | n437 ;
  assign n11161 = n174 | n11160 ;
  assign n11162 = n11159 | n11161 ;
  assign n11163 = n11156 | n11162 ;
  assign n11164 = n103 | n224 ;
  assign n11165 = n11163 | n11164 ;
  assign n11166 = n11148 | n11165 ;
  assign n11167 = n571 | n1866 ;
  assign n11168 = n2922 | n11167 ;
  assign n11169 = n242 | n11168 ;
  assign n11170 = n468 | n11169 ;
  assign n11171 = n539 | n11170 ;
  assign n11172 = n240 | n11171 ;
  assign n11173 = n416 | n11172 ;
  assign n11174 = n610 | n11173 ;
  assign n11175 = n11166 | n11174 ;
  assign n11176 = n449 | n1596 ;
  assign n11177 = n10926 | n11176 ;
  assign n11178 = n101 | n3150 ;
  assign n11179 = n277 | n531 ;
  assign n11180 = ( ~n297 & n11178 ) | ( ~n297 & n11179 ) | ( n11178 & n11179 ) ;
  assign n11181 = n297 | n11180 ;
  assign n11182 = n11177 | n11181 ;
  assign n11183 = n955 | n3000 ;
  assign n11184 = n11182 | n11183 ;
  assign n11185 = n1023 | n1054 ;
  assign n11186 = n1416 | n11185 ;
  assign n11187 = n1920 | n11186 ;
  assign n11188 = n1260 | n11187 ;
  assign n11189 = n509 | n11188 ;
  assign n11190 = n11184 | n11189 ;
  assign n11191 = n2169 | n3659 ;
  assign n11192 = n529 | n655 ;
  assign n11193 = n522 | n11192 ;
  assign n11194 = n11191 | n11193 ;
  assign n11195 = n133 | n164 ;
  assign n11196 = n434 | n11195 ;
  assign n11197 = n11194 | n11196 ;
  assign n11198 = n1117 | n3004 ;
  assign n11199 = n3116 | n11198 ;
  assign n11200 = n476 | n590 ;
  assign n11201 = n167 | n645 ;
  assign n11202 = n11200 | n11201 ;
  assign n11203 = n11199 | n11202 ;
  assign n11204 = n468 | n634 ;
  assign n11205 = n359 | n11204 ;
  assign n11206 = n65 | n11205 ;
  assign n11207 = n155 | n11206 ;
  assign n11208 = n218 | n11207 ;
  assign n11209 = n11203 | n11208 ;
  assign n11210 = n11197 | n11209 ;
  assign n11211 = n11190 | n11210 ;
  assign n11212 = n960 | n2147 ;
  assign n11213 = n3435 | n11212 ;
  assign n11214 = n300 | n380 ;
  assign n11215 = n990 | n11214 ;
  assign n11216 = n197 | n2481 ;
  assign n11217 = n11215 | n11216 ;
  assign n11218 = n11213 | n11217 ;
  assign n11219 = n209 | n470 ;
  assign n11220 = n249 | n11219 ;
  assign n11221 = n438 | n11220 ;
  assign n11222 = n11218 | n11221 ;
  assign n11223 = n5640 | n11222 ;
  assign n11224 = n11211 | n11223 ;
  assign n11225 = n484 | n4101 ;
  assign n11226 = n618 | n11225 ;
  assign n11227 = n263 | n11226 ;
  assign n11228 = n279 | n11227 ;
  assign n11229 = n383 | n11228 ;
  assign n11230 = ( n151 & ~n2799 ) | ( n151 & n11229 ) | ( ~n2799 & n11229 ) ;
  assign n11231 = n2799 | n11230 ;
  assign n11232 = n11224 | n11231 ;
  assign n11233 = n649 | n11232 ;
  assign n11234 = ( x23 & ~n11175 ) | ( x23 & n11233 ) | ( ~n11175 & n11233 ) ;
  assign n11235 = ( ~x23 & n11175 ) | ( ~x23 & n11234 ) | ( n11175 & n11234 ) ;
  assign n11236 = ~n10924 & n11235 ;
  assign n11237 = n904 & n3639 ;
  assign n11238 = n778 & n3727 ;
  assign n11239 = n11237 | n11238 ;
  assign n11240 = ~n3596 & n3744 ;
  assign n11241 = n11239 | n11240 ;
  assign n11242 = n3636 | n11241 ;
  assign n11243 = ( ~n4649 & n11241 ) | ( ~n4649 & n11242 ) | ( n11241 & n11242 ) ;
  assign n11244 = n10924 & ~n11235 ;
  assign n11245 = n11236 | n11244 ;
  assign n11246 = n11243 & n11245 ;
  assign n11247 = n11245 & ~n11246 ;
  assign n11248 = ( n11243 & ~n11246 ) | ( n11243 & n11247 ) | ( ~n11246 & n11247 ) ;
  assign n11249 = ( n11236 & n11243 ) | ( n11236 & n11248 ) | ( n11243 & n11248 ) ;
  assign n11129 = n11101 | n11113 ;
  assign n11250 = ~n11129 & n11249 ;
  assign n11251 = ( n11128 & n11249 ) | ( n11128 & n11250 ) | ( n11249 & n11250 ) ;
  assign n11252 = n11129 & ~n11249 ;
  assign n11253 = ~n11128 & n11252 ;
  assign n11254 = n778 & n3744 ;
  assign n11255 = ~n1014 & n3639 ;
  assign n11256 = n904 & n3727 ;
  assign n11257 = n11255 | n11256 ;
  assign n11258 = n11254 | n11257 ;
  assign n11259 = n3636 | n11258 ;
  assign n11260 = ( ~n4535 & n11258 ) | ( ~n4535 & n11259 ) | ( n11258 & n11259 ) ;
  assign n11261 = ( ~n11233 & n11234 ) | ( ~n11233 & n11235 ) | ( n11234 & n11235 ) ;
  assign n11262 = n11260 & ~n11261 ;
  assign n11263 = ~n11260 & n11261 ;
  assign n11264 = n11262 | n11263 ;
  assign n11265 = n2527 | n4163 ;
  assign n11266 = n640 | n11265 ;
  assign n11267 = ~n1779 & n3233 ;
  assign n11268 = ~n3322 & n11267 ;
  assign n11269 = ~n11266 & n11268 ;
  assign n11270 = ~n2739 & n11269 ;
  assign n11271 = ~n1306 & n11270 ;
  assign n11272 = ~n869 & n11271 ;
  assign n11273 = ~n2285 & n11272 ;
  assign n11274 = n301 | n621 ;
  assign n11275 = n608 | n11274 ;
  assign n11276 = n279 | n647 ;
  assign n11277 = n3910 | n11276 ;
  assign n11278 = n11275 | n11277 ;
  assign n11279 = n3371 | n3476 ;
  assign n11280 = n367 | n11279 ;
  assign n11281 = n11278 | n11280 ;
  assign n11282 = n1443 | n11281 ;
  assign n11283 = n326 | n383 ;
  assign n11284 = n400 | n11283 ;
  assign n11285 = n595 | n11284 ;
  assign n11286 = n253 | n2738 ;
  assign n11287 = n11285 | n11286 ;
  assign n11288 = n1607 | n11287 ;
  assign n11289 = n11282 | n11288 ;
  assign n11290 = n101 | n1354 ;
  assign n11291 = n429 | n11290 ;
  assign n11292 = n245 | n11291 ;
  assign n11293 = n393 | n11292 ;
  assign n11294 = n11289 | n11293 ;
  assign n11295 = n379 | n483 ;
  assign n11296 = n90 | n11295 ;
  assign n11297 = n244 | n500 ;
  assign n11298 = n241 | n11297 ;
  assign n11299 = n509 | n11298 ;
  assign n11300 = n11296 | n11299 ;
  assign n11301 = n96 | n112 ;
  assign n11302 = n11300 | n11301 ;
  assign n11303 = n11294 | n11302 ;
  assign n11304 = n1044 | n11303 ;
  assign n11305 = n11273 & ~n11304 ;
  assign n11306 = n520 | n1178 ;
  assign n11307 = n277 | n11306 ;
  assign n11308 = n191 | n11307 ;
  assign n11309 = n11305 & ~n11308 ;
  assign n11310 = n11175 | n11309 ;
  assign n11311 = n11175 & n11309 ;
  assign n11312 = n240 | n1216 ;
  assign n11313 = n351 | n11312 ;
  assign n11314 = n358 | n11313 ;
  assign n11315 = n583 | n11314 ;
  assign n11316 = n403 | n11315 ;
  assign n11317 = n3315 | n11298 ;
  assign n11318 = n144 | n2635 ;
  assign n11319 = n2154 | n11318 ;
  assign n11320 = n1784 | n11319 ;
  assign n11321 = ( ~n4168 & n11317 ) | ( ~n4168 & n11320 ) | ( n11317 & n11320 ) ;
  assign n11322 = n4168 | n11321 ;
  assign n11323 = n11316 | n11322 ;
  assign n11324 = n128 | n11323 ;
  assign n11325 = n1466 | n3463 ;
  assign n11326 = n1351 | n3776 ;
  assign n11327 = n11325 | n11326 ;
  assign n11328 = n391 | n621 ;
  assign n11329 = n2164 | n11328 ;
  assign n11330 = n451 | n622 ;
  assign n11331 = n437 | n11330 ;
  assign n11332 = n11329 | n11331 ;
  assign n11333 = n1867 | n11332 ;
  assign n11334 = n11327 | n11333 ;
  assign n11335 = n367 | n2665 ;
  assign n11336 = n2922 | n11335 ;
  assign n11337 = n284 | n11336 ;
  assign n11338 = n11334 | n11337 ;
  assign n11339 = n428 | n608 ;
  assign n11340 = n140 | n11339 ;
  assign n11341 = n11338 | n11340 ;
  assign n11342 = n1240 | n2960 ;
  assign n11343 = n474 | n11342 ;
  assign n11344 = n849 | n1200 ;
  assign n11345 = n11343 | n11344 ;
  assign n11346 = n3138 | n11345 ;
  assign n11347 = n3010 | n11346 ;
  assign n11348 = n1811 | n11347 ;
  assign n11349 = n11341 | n11348 ;
  assign n11350 = n11324 | n11349 ;
  assign n11351 = n1522 | n1920 ;
  assign n11352 = n1989 | n11351 ;
  assign n11353 = n484 | n11352 ;
  assign n11354 = n276 | n11353 ;
  assign n11355 = n296 | n11354 ;
  assign n11356 = n580 | n11355 ;
  assign n11357 = n438 | n11356 ;
  assign n11358 = n133 | n11357 ;
  assign n11359 = n11350 | n11358 ;
  assign n11360 = n280 | n391 ;
  assign n11361 = n102 | n11360 ;
  assign n11362 = n141 | n2433 ;
  assign n11363 = n11361 | n11362 ;
  assign n11364 = n199 | n583 ;
  assign n11365 = n161 | n11364 ;
  assign n11366 = n126 | n11365 ;
  assign n11367 = n11363 | n11366 ;
  assign n11368 = n207 | n11367 ;
  assign n11369 = n83 | n646 ;
  assign n11370 = n4101 | n11369 ;
  assign n11371 = n2216 | n11370 ;
  assign n11372 = n418 | n891 ;
  assign n11373 = n4879 | n11372 ;
  assign n11374 = n11371 | n11373 ;
  assign n11375 = n59 | n2527 ;
  assign n11376 = n1959 | n11375 ;
  assign n11377 = n1352 | n11376 ;
  assign n11378 = n11374 | n11377 ;
  assign n11379 = n1272 | n2689 ;
  assign n11380 = n306 | n321 ;
  assign n11381 = n203 | n11380 ;
  assign n11382 = n11379 | n11381 ;
  assign n11383 = n1044 | n11382 ;
  assign n11384 = n1022 | n11383 ;
  assign n11385 = n11378 | n11384 ;
  assign n11386 = n479 | n1989 ;
  assign n11387 = n639 | n11386 ;
  assign n11388 = n279 | n11387 ;
  assign n11389 = n252 | n11388 ;
  assign n11390 = n11385 | n11389 ;
  assign n11391 = n11368 | n11390 ;
  assign n11392 = n831 | n2235 ;
  assign n11393 = n3540 | n11392 ;
  assign n11394 = n269 | n356 ;
  assign n11395 = n366 | n11394 ;
  assign n11396 = n569 | n11395 ;
  assign n11397 = n472 | n475 ;
  assign n11398 = n630 | n11397 ;
  assign n11399 = ( n335 & ~n4113 ) | ( n335 & n11398 ) | ( ~n4113 & n11398 ) ;
  assign n11400 = n4113 | n11399 ;
  assign n11401 = n11396 | n11400 ;
  assign n11402 = n103 | n601 ;
  assign n11403 = n173 | n11402 ;
  assign n11404 = n647 | n11403 ;
  assign n11405 = n11401 | n11404 ;
  assign n11406 = ( ~n4866 & n11393 ) | ( ~n4866 & n11405 ) | ( n11393 & n11405 ) ;
  assign n11407 = n4866 | n11406 ;
  assign n11408 = n11391 | n11407 ;
  assign n11409 = n1079 | n1170 ;
  assign n11410 = n759 | n11409 ;
  assign n11411 = n621 | n11410 ;
  assign n11412 = n146 | n11411 ;
  assign n11413 = n122 | n11412 ;
  assign n11414 = n223 | n11413 ;
  assign n11415 = n11408 | n11414 ;
  assign n11416 = ( x20 & ~n11359 ) | ( x20 & n11415 ) | ( ~n11359 & n11415 ) ;
  assign n11417 = ( ~x20 & n11359 ) | ( ~x20 & n11416 ) | ( n11359 & n11416 ) ;
  assign n11418 = ~n1014 & n3744 ;
  assign n11419 = n3349 & n3639 ;
  assign n11420 = ~n3255 & n3727 ;
  assign n11421 = n11419 | n11420 ;
  assign n11422 = n11418 | n11421 ;
  assign n11423 = n3636 | n11422 ;
  assign n11424 = ( n11309 & n11417 ) | ( n11309 & n11423 ) | ( n11417 & n11423 ) ;
  assign n11425 = n11310 & n11424 ;
  assign n11426 = ~n11311 & n11425 ;
  assign n11427 = ( n11309 & n11417 ) | ( n11309 & n11422 ) | ( n11417 & n11422 ) ;
  assign n11428 = n11310 & n11427 ;
  assign n11429 = ~n11311 & n11428 ;
  assign n11430 = ( n4742 & n11426 ) | ( n4742 & n11429 ) | ( n11426 & n11429 ) ;
  assign n11431 = n11310 & ~n11430 ;
  assign n11432 = n11264 | n11431 ;
  assign n11433 = ~n11262 & n11432 ;
  assign n11434 = n11248 | n11433 ;
  assign n11435 = n11248 & n11433 ;
  assign n11436 = n11434 & ~n11435 ;
  assign n11437 = n3504 & n4043 ;
  assign n11438 = ~n3431 & n4045 ;
  assign n11439 = n11437 | n11438 ;
  assign n11440 = ~n589 & n4048 ;
  assign n11441 = n11439 | n11440 ;
  assign n11442 = n4051 | n11441 ;
  assign n11443 = ( n4765 & n11441 ) | ( n4765 & n11442 ) | ( n11441 & n11442 ) ;
  assign n11444 = x29 & n11443 ;
  assign n11445 = x29 & ~n11444 ;
  assign n11446 = ( n11443 & ~n11444 ) | ( n11443 & n11445 ) | ( ~n11444 & n11445 ) ;
  assign n11447 = n11436 & n11446 ;
  assign n11448 = n11434 & ~n11447 ;
  assign n11449 = ( ~n11251 & n11253 ) | ( ~n11251 & n11448 ) | ( n11253 & n11448 ) ;
  assign n11450 = n11117 | n11449 ;
  assign n11451 = n11117 & n11449 ;
  assign n11452 = n11450 & ~n11451 ;
  assign n11453 = ~n3634 & n4048 ;
  assign n11454 = ~n672 & n4045 ;
  assign n11455 = n11453 | n11454 ;
  assign n11456 = ~n589 & n4043 ;
  assign n11457 = n11455 | n11456 ;
  assign n11458 = n4051 | n11457 ;
  assign n11459 = ( ~n5092 & n11457 ) | ( ~n5092 & n11458 ) | ( n11457 & n11458 ) ;
  assign n11460 = ~x29 & n11459 ;
  assign n11461 = x29 | n11460 ;
  assign n11462 = ( ~n11459 & n11460 ) | ( ~n11459 & n11461 ) | ( n11460 & n11461 ) ;
  assign n11463 = n11452 & ~n11462 ;
  assign n11464 = ( n11450 & ~n11452 ) | ( n11450 & n11463 ) | ( ~n11452 & n11463 ) ;
  assign n11465 = ( ~n11036 & n11118 ) | ( ~n11036 & n11122 ) | ( n11118 & n11122 ) ;
  assign n11466 = ( n11036 & ~n11122 ) | ( n11036 & n11465 ) | ( ~n11122 & n11465 ) ;
  assign n11467 = ( ~n11118 & n11465 ) | ( ~n11118 & n11466 ) | ( n11465 & n11466 ) ;
  assign n11468 = ~n11464 & n11467 ;
  assign n11469 = n11464 & ~n11467 ;
  assign n11470 = n11468 | n11469 ;
  assign n11471 = ~n11452 & n11462 ;
  assign n11472 = n11463 | n11471 ;
  assign n11473 = ~n3431 & n4043 ;
  assign n11474 = ~n589 & n4045 ;
  assign n11475 = n11473 | n11474 ;
  assign n11476 = ~n672 & n4048 ;
  assign n11477 = n11475 | n11476 ;
  assign n11478 = n4051 | n11477 ;
  assign n11479 = ( ~n5353 & n11477 ) | ( ~n5353 & n11478 ) | ( n11477 & n11478 ) ;
  assign n11480 = ~x29 & n11479 ;
  assign n11481 = x29 | n11480 ;
  assign n11482 = ( ~n11479 & n11480 ) | ( ~n11479 & n11481 ) | ( n11480 & n11481 ) ;
  assign n11483 = n4479 | n4487 ;
  assign n11484 = ~n3634 & n11483 ;
  assign n11485 = n672 & n4479 ;
  assign n11486 = ( ~n672 & n11484 ) | ( ~n672 & n11485 ) | ( n11484 & n11485 ) ;
  assign n11487 = ( ~n3619 & n11484 ) | ( ~n3619 & n11486 ) | ( n11484 & n11486 ) ;
  assign n11488 = ~x26 & n11487 ;
  assign n11489 = x26 | n11488 ;
  assign n11490 = ( ~n11487 & n11488 ) | ( ~n11487 & n11489 ) | ( n11488 & n11489 ) ;
  assign n11491 = n11482 & n11490 ;
  assign n11492 = n11251 | n11253 ;
  assign n11493 = n11448 | n11492 ;
  assign n11494 = n11448 & n11492 ;
  assign n11495 = n11493 & ~n11494 ;
  assign n11496 = n11490 & ~n11491 ;
  assign n11497 = ( n11482 & ~n11491 ) | ( n11482 & n11496 ) | ( ~n11491 & n11496 ) ;
  assign n11498 = n11495 & n11497 ;
  assign n11499 = n11491 | n11498 ;
  assign n11500 = n11472 & n11499 ;
  assign n11501 = n11436 | n11446 ;
  assign n11502 = ~n11447 & n11501 ;
  assign n11503 = n11264 & n11431 ;
  assign n11504 = n11432 & ~n11503 ;
  assign n11505 = ( n4742 & n11424 ) | ( n4742 & n11427 ) | ( n11424 & n11427 ) ;
  assign n11506 = ~n11430 & n11505 ;
  assign n11507 = ~n11311 & n11431 ;
  assign n11508 = n11506 | n11507 ;
  assign n11509 = n904 & n3744 ;
  assign n11510 = ~n1014 & n3727 ;
  assign n11511 = ~n3255 & n3639 ;
  assign n11512 = n11510 | n11511 ;
  assign n11513 = n3636 | n11512 ;
  assign n11514 = ( n4632 & n11512 ) | ( n4632 & n11513 ) | ( n11512 & n11513 ) ;
  assign n11515 = n11509 | n11514 ;
  assign n11516 = n11508 & n11515 ;
  assign n11517 = n3511 | n4392 ;
  assign n11518 = n910 | n4367 ;
  assign n11519 = n11517 | n11518 ;
  assign n11520 = n337 | n482 ;
  assign n11521 = n2610 | n11520 ;
  assign n11522 = n279 | n622 ;
  assign n11523 = n241 | n11522 ;
  assign n11524 = n11521 | n11523 ;
  assign n11525 = n601 | n607 ;
  assign n11526 = n11524 | n11525 ;
  assign n11527 = n639 | n2900 ;
  assign n11528 = n404 | n11527 ;
  assign n11529 = n1756 | n11528 ;
  assign n11530 = n11526 | n11529 ;
  assign n11531 = n11519 | n11530 ;
  assign n11532 = n808 | n1057 ;
  assign n11533 = ( n500 & ~n2346 ) | ( n500 & n11532 ) | ( ~n2346 & n11532 ) ;
  assign n11534 = n2346 | n11533 ;
  assign n11535 = n393 | n11534 ;
  assign n11536 = n11531 | n11535 ;
  assign n11537 = n645 | n647 ;
  assign n11538 = n11536 | n11537 ;
  assign n11539 = n3150 | n5741 ;
  assign n11540 = n1836 & ~n11539 ;
  assign n11541 = ~n3305 & n11540 ;
  assign n11542 = ~n2132 & n11541 ;
  assign n11543 = ~n650 & n11542 ;
  assign n11544 = ~n4356 & n11543 ;
  assign n11545 = ~n11538 & n11544 ;
  assign n11546 = n1314 | n3850 ;
  assign n11547 = n1044 | n11546 ;
  assign n11548 = n862 | n11547 ;
  assign n11549 = n270 | n11548 ;
  assign n11550 = n315 | n11549 ;
  assign n11551 = n122 | n11550 ;
  assign n11552 = n11545 & ~n11551 ;
  assign n11553 = n11359 | n11552 ;
  assign n11554 = n11359 & n11552 ;
  assign n11555 = ~n1151 & n3639 ;
  assign n11556 = n1233 & n3727 ;
  assign n11557 = n11555 | n11556 ;
  assign n11558 = n3349 & n3744 ;
  assign n11559 = n11557 | n11558 ;
  assign n11560 = n3636 | n11559 ;
  assign n11561 = n11553 & n11560 ;
  assign n11562 = ~n11554 & n11561 ;
  assign n11563 = n11553 & n11559 ;
  assign n11564 = ~n11554 & n11563 ;
  assign n11565 = ( n4518 & n11562 ) | ( n4518 & n11564 ) | ( n11562 & n11564 ) ;
  assign n11566 = n11553 & ~n11565 ;
  assign n11567 = ( ~n11415 & n11416 ) | ( ~n11415 & n11417 ) | ( n11416 & n11417 ) ;
  assign n11568 = n11566 | n11567 ;
  assign n11569 = n11566 & n11567 ;
  assign n11570 = n11568 & ~n11569 ;
  assign n11571 = n1233 & n3639 ;
  assign n11572 = n3349 & n3727 ;
  assign n11573 = n11571 | n11572 ;
  assign n11574 = ~n3255 & n3744 ;
  assign n11575 = n11573 | n11574 ;
  assign n11576 = n3636 | n11575 ;
  assign n11577 = ( ~n4470 & n11575 ) | ( ~n4470 & n11576 ) | ( n11575 & n11576 ) ;
  assign n11578 = n11570 & ~n11577 ;
  assign n11579 = ( n11566 & n11567 ) | ( n11566 & n11578 ) | ( n11567 & n11578 ) ;
  assign n11580 = ( n4742 & n11422 ) | ( n4742 & n11423 ) | ( n11422 & n11423 ) ;
  assign n11581 = ( n11309 & n11417 ) | ( n11309 & ~n11580 ) | ( n11417 & ~n11580 ) ;
  assign n11582 = ( ~n11417 & n11580 ) | ( ~n11417 & n11581 ) | ( n11580 & n11581 ) ;
  assign n11583 = ( ~n11309 & n11581 ) | ( ~n11309 & n11582 ) | ( n11581 & n11582 ) ;
  assign n11584 = ~n11579 & n11583 ;
  assign n11585 = n11579 & ~n11583 ;
  assign n11586 = n11584 | n11585 ;
  assign n11587 = n904 & n4043 ;
  assign n11588 = n778 & n4045 ;
  assign n11589 = n11587 | n11588 ;
  assign n11590 = ~n3596 & n4048 ;
  assign n11591 = n11589 | n11590 ;
  assign n11592 = n4051 | n11591 ;
  assign n11593 = ( ~n4649 & n11591 ) | ( ~n4649 & n11592 ) | ( n11591 & n11592 ) ;
  assign n11594 = ~x29 & n11593 ;
  assign n11595 = x29 | n11594 ;
  assign n11596 = ( ~n11593 & n11594 ) | ( ~n11593 & n11595 ) | ( n11594 & n11595 ) ;
  assign n11597 = ~n11586 & n11596 ;
  assign n11598 = n11584 | n11597 ;
  assign n11599 = n11508 | n11515 ;
  assign n11600 = ~n11516 & n11599 ;
  assign n11601 = n11598 & n11600 ;
  assign n11602 = n11516 | n11601 ;
  assign n11603 = ~n3596 & n4043 ;
  assign n11604 = n3504 & n4045 ;
  assign n11605 = n11603 | n11604 ;
  assign n11606 = ~n3431 & n4048 ;
  assign n11607 = n11605 | n11606 ;
  assign n11608 = n4051 | n11607 ;
  assign n11609 = ( ~n4798 & n11607 ) | ( ~n4798 & n11608 ) | ( n11607 & n11608 ) ;
  assign n11610 = ~x29 & n11609 ;
  assign n11611 = x29 | n11610 ;
  assign n11612 = ( ~n11609 & n11610 ) | ( ~n11609 & n11611 ) | ( n11610 & n11611 ) ;
  assign n11613 = ( n11504 & n11602 ) | ( n11504 & n11612 ) | ( n11602 & n11612 ) ;
  assign n11614 = n11502 & n11613 ;
  assign n11615 = n11613 & ~n11614 ;
  assign n11616 = n11502 & ~n11613 ;
  assign n11617 = ~n3634 & n4481 ;
  assign n11618 = ( n4479 & ~n11485 ) | ( n4479 & n11617 ) | ( ~n11485 & n11617 ) ;
  assign n11619 = n4487 | n11618 ;
  assign n11620 = ( n3726 & n11618 ) | ( n3726 & n11619 ) | ( n11618 & n11619 ) ;
  assign n11621 = x26 & n11620 ;
  assign n11622 = x26 & ~n11621 ;
  assign n11623 = ( n11620 & ~n11621 ) | ( n11620 & n11622 ) | ( ~n11621 & n11622 ) ;
  assign n11624 = ( n11615 & n11616 ) | ( n11615 & n11623 ) | ( n11616 & n11623 ) ;
  assign n11625 = n11495 | n11497 ;
  assign n11626 = ~n11498 & n11625 ;
  assign n11627 = ( n11614 & n11624 ) | ( n11614 & n11626 ) | ( n11624 & n11626 ) ;
  assign n11628 = n11614 | n11626 ;
  assign n11629 = n11624 | n11628 ;
  assign n11630 = ~n11627 & n11629 ;
  assign n11631 = ~n3634 & n4484 ;
  assign n11632 = ~n672 & n4481 ;
  assign n11633 = n11631 | n11632 ;
  assign n11634 = ~n589 & n4479 ;
  assign n11635 = n11633 | n11634 ;
  assign n11636 = n4487 | n11635 ;
  assign n11637 = ( ~n5092 & n11635 ) | ( ~n5092 & n11636 ) | ( n11635 & n11636 ) ;
  assign n11638 = ~x26 & n11637 ;
  assign n11639 = x26 | n11638 ;
  assign n11640 = ( ~n11637 & n11638 ) | ( ~n11637 & n11639 ) | ( n11638 & n11639 ) ;
  assign n11641 = n11598 & ~n11601 ;
  assign n11642 = ~n11598 & n11600 ;
  assign n11643 = n778 & n4043 ;
  assign n11644 = ~n3596 & n4045 ;
  assign n11645 = n11643 | n11644 ;
  assign n11646 = n3504 & n4048 ;
  assign n11647 = n11645 | n11646 ;
  assign n11648 = n4051 | n11647 ;
  assign n11649 = ( ~n5040 & n11647 ) | ( ~n5040 & n11648 ) | ( n11647 & n11648 ) ;
  assign n11650 = ~x29 & n11649 ;
  assign n11651 = x29 | n11650 ;
  assign n11652 = ( ~n11649 & n11650 ) | ( ~n11649 & n11651 ) | ( n11650 & n11651 ) ;
  assign n11653 = n11642 | n11652 ;
  assign n11654 = n11641 | n11653 ;
  assign n11655 = ( n11641 & n11642 ) | ( n11641 & n11652 ) | ( n11642 & n11652 ) ;
  assign n11656 = ~n3431 & n4479 ;
  assign n11657 = ~n589 & n4481 ;
  assign n11658 = n11656 | n11657 ;
  assign n11659 = ~n672 & n4484 ;
  assign n11660 = n11658 | n11659 ;
  assign n11661 = n4487 | n11660 ;
  assign n11662 = ( ~n5353 & n11660 ) | ( ~n5353 & n11661 ) | ( n11660 & n11661 ) ;
  assign n11663 = ~x26 & n11662 ;
  assign n11664 = x26 | n11663 ;
  assign n11665 = ( ~n11662 & n11663 ) | ( ~n11662 & n11664 ) | ( n11663 & n11664 ) ;
  assign n11666 = ( n11654 & n11655 ) | ( n11654 & n11665 ) | ( n11655 & n11665 ) ;
  assign n11667 = n11640 & n11666 ;
  assign n11668 = n11666 & ~n11667 ;
  assign n11669 = n11640 & ~n11666 ;
  assign n11670 = ( n11504 & n11612 ) | ( n11504 & ~n11613 ) | ( n11612 & ~n11613 ) ;
  assign n11671 = ( n11602 & ~n11613 ) | ( n11602 & n11670 ) | ( ~n11613 & n11670 ) ;
  assign n11672 = ( n11668 & n11669 ) | ( n11668 & n11671 ) | ( n11669 & n11671 ) ;
  assign n11673 = n11667 | n11672 ;
  assign n11674 = n11616 | n11623 ;
  assign n11675 = n11615 | n11674 ;
  assign n11676 = ~n11624 & n11675 ;
  assign n11677 = n11673 & n11676 ;
  assign n11678 = n11673 | n11676 ;
  assign n11679 = ~n11677 & n11678 ;
  assign n11680 = ~n11570 & n11577 ;
  assign n11681 = n11578 | n11680 ;
  assign n11682 = ~n1014 & n4043 ;
  assign n11683 = n904 & n4045 ;
  assign n11684 = n11682 | n11683 ;
  assign n11685 = n778 & n4048 ;
  assign n11686 = n11684 | n11685 ;
  assign n11687 = n4051 | n11686 ;
  assign n11688 = ( ~n4535 & n11686 ) | ( ~n4535 & n11687 ) | ( n11686 & n11687 ) ;
  assign n11689 = ~x29 & n11688 ;
  assign n11690 = x29 | n11689 ;
  assign n11691 = ( ~n11688 & n11689 ) | ( ~n11688 & n11690 ) | ( n11689 & n11690 ) ;
  assign n11692 = n11681 & n11691 ;
  assign n11693 = n11681 | n11691 ;
  assign n11694 = ~n11692 & n11693 ;
  assign n11695 = ( n4518 & n11559 ) | ( n4518 & n11560 ) | ( n11559 & n11560 ) ;
  assign n11696 = ~n11565 & n11695 ;
  assign n11697 = n373 | n633 ;
  assign n11698 = n250 | n300 ;
  assign n11699 = n11697 | n11698 ;
  assign n11700 = n620 | n3218 ;
  assign n11701 = n850 | n2165 ;
  assign n11702 = n11700 | n11701 ;
  assign n11703 = n11699 | n11702 ;
  assign n11704 = n926 | n1271 ;
  assign n11705 = n11703 | n11704 ;
  assign n11706 = n2186 | n11705 ;
  assign n11707 = n3387 | n11706 ;
  assign n11708 = n3573 & ~n11707 ;
  assign n11709 = n1337 | n2427 ;
  assign n11710 = n1261 | n11709 ;
  assign n11711 = n11708 & ~n11710 ;
  assign n11712 = n349 | n3856 ;
  assign n11713 = n326 | n11712 ;
  assign n11714 = n596 | n11713 ;
  assign n11715 = n160 | n11714 ;
  assign n11716 = n11711 & ~n11715 ;
  assign n11717 = n437 | n521 ;
  assign n11718 = n2834 | n11717 ;
  assign n11719 = n3946 | n11718 ;
  assign n11720 = n2207 | n11719 ;
  assign n11721 = n595 | n11720 ;
  assign n11722 = n828 | n11721 ;
  assign n11723 = n5611 | n5620 ;
  assign n11724 = n248 | n11723 ;
  assign n11725 = n11722 | n11724 ;
  assign n11726 = n1057 | n1279 ;
  assign n11727 = n611 | n11726 ;
  assign n11728 = n2867 | n11727 ;
  assign n11729 = n483 | n11728 ;
  assign n11730 = n633 | n11729 ;
  assign n11731 = ( n349 & ~n2899 ) | ( n349 & n11730 ) | ( ~n2899 & n11730 ) ;
  assign n11732 = n2899 | n11731 ;
  assign n11733 = n11725 | n11732 ;
  assign n11734 = n419 | n2956 ;
  assign n11735 = n597 | n11734 ;
  assign n11736 = n92 | n11735 ;
  assign n11737 = ~n11716 & n11736 ;
  assign n11738 = ( ~n11716 & n11733 ) | ( ~n11716 & n11737 ) | ( n11733 & n11737 ) ;
  assign n11739 = n11716 & ~n11736 ;
  assign n11740 = ~n11733 & n11739 ;
  assign n11741 = n11738 | n11740 ;
  assign n11742 = x17 & ~n11738 ;
  assign n11743 = ( ~n11738 & n11741 ) | ( ~n11738 & n11742 ) | ( n11741 & n11742 ) ;
  assign n11744 = n11359 | n11743 ;
  assign n11745 = n1327 & n3639 ;
  assign n11746 = ~n1151 & n3727 ;
  assign n11747 = n11745 | n11746 ;
  assign n11748 = n1233 & n3744 ;
  assign n11749 = n11747 | n11748 ;
  assign n11750 = n3636 | n11749 ;
  assign n11751 = ( ~n4615 & n11749 ) | ( ~n4615 & n11750 ) | ( n11749 & n11750 ) ;
  assign n11752 = n11359 & n11743 ;
  assign n11753 = n11744 & ~n11752 ;
  assign n11754 = n11751 & n11753 ;
  assign n11755 = n11744 & ~n11754 ;
  assign n11756 = ~n11554 & n11566 ;
  assign n11757 = ~n11755 & n11756 ;
  assign n11758 = ( n11696 & ~n11755 ) | ( n11696 & n11757 ) | ( ~n11755 & n11757 ) ;
  assign n11759 = n11755 & ~n11756 ;
  assign n11760 = ~n11696 & n11759 ;
  assign n11761 = n11758 | n11760 ;
  assign n11762 = ~n11740 & n11743 ;
  assign n11763 = ~x17 & n11741 ;
  assign n11764 = n11762 | n11763 ;
  assign n11765 = ~n1151 & n3744 ;
  assign n11766 = n1327 & n3727 ;
  assign n11767 = n3104 & n3639 ;
  assign n11768 = n11766 | n11767 ;
  assign n11769 = n11765 | n11768 ;
  assign n11770 = n3636 | n11769 ;
  assign n11771 = ( ~n4034 & n11769 ) | ( ~n4034 & n11770 ) | ( n11769 & n11770 ) ;
  assign n11772 = n11764 & n11771 ;
  assign n11773 = n11764 | n11771 ;
  assign n11774 = ~n11772 & n11773 ;
  assign n11775 = n4716 & n11716 ;
  assign n11776 = n4716 | n11716 ;
  assign n11777 = ( n4023 & ~n4667 ) | ( n4023 & n4716 ) | ( ~n4667 & n4716 ) ;
  assign n11778 = ( ~n3636 & n4718 ) | ( ~n3636 & n11777 ) | ( n4718 & n11777 ) ;
  assign n11779 = n11775 | n11778 ;
  assign n11780 = n11776 & ~n11779 ;
  assign n11781 = n11775 | n11777 ;
  assign n11782 = n11776 & ~n11781 ;
  assign n11783 = ( n4449 & n11780 ) | ( n4449 & n11782 ) | ( n11780 & n11782 ) ;
  assign n11784 = n11775 | n11783 ;
  assign n11785 = n11774 & n11784 ;
  assign n11786 = n11772 | n11785 ;
  assign n11787 = n11753 & ~n11754 ;
  assign n11788 = ( n11751 & ~n11754 ) | ( n11751 & n11787 ) | ( ~n11754 & n11787 ) ;
  assign n11789 = n11786 & n11788 ;
  assign n11790 = n11786 | n11788 ;
  assign n11791 = ~n11789 & n11790 ;
  assign n11792 = ~n1014 & n4048 ;
  assign n11793 = n3349 & n4043 ;
  assign n11794 = ~n3255 & n4045 ;
  assign n11795 = n11793 | n11794 ;
  assign n11796 = n11792 | n11795 ;
  assign n11797 = n4051 | n11796 ;
  assign n11798 = ( n4742 & n11796 ) | ( n4742 & n11797 ) | ( n11796 & n11797 ) ;
  assign n11799 = x29 & n11798 ;
  assign n11800 = x29 & ~n11799 ;
  assign n11801 = ( n11798 & ~n11799 ) | ( n11798 & n11800 ) | ( ~n11799 & n11800 ) ;
  assign n11802 = n11791 & n11801 ;
  assign n11803 = n11789 | n11802 ;
  assign n11804 = ~n11761 & n11803 ;
  assign n11805 = n11758 | n11804 ;
  assign n11806 = n11694 & n11805 ;
  assign n11807 = n11692 | n11806 ;
  assign n11808 = n11586 & ~n11596 ;
  assign n11809 = n11597 | n11808 ;
  assign n11810 = n11807 & ~n11809 ;
  assign n11811 = n11807 & ~n11810 ;
  assign n11812 = n11807 | n11809 ;
  assign n11813 = n3504 & n4479 ;
  assign n11814 = ~n3431 & n4481 ;
  assign n11815 = n11813 | n11814 ;
  assign n11816 = ~n589 & n4484 ;
  assign n11817 = n11815 | n11816 ;
  assign n11818 = n4487 | n11817 ;
  assign n11819 = ( n4765 & n11817 ) | ( n4765 & n11818 ) | ( n11817 & n11818 ) ;
  assign n11820 = x26 & n11819 ;
  assign n11821 = x26 & ~n11820 ;
  assign n11822 = ( n11819 & ~n11820 ) | ( n11819 & n11821 ) | ( ~n11820 & n11821 ) ;
  assign n11823 = ( n11811 & ~n11812 ) | ( n11811 & n11822 ) | ( ~n11812 & n11822 ) ;
  assign n11824 = n4546 | n4554 ;
  assign n11825 = ~n3634 & n11824 ;
  assign n11826 = n672 & n4546 ;
  assign n11827 = ( ~n672 & n11825 ) | ( ~n672 & n11826 ) | ( n11825 & n11826 ) ;
  assign n11828 = ( ~n3619 & n11825 ) | ( ~n3619 & n11827 ) | ( n11825 & n11827 ) ;
  assign n11829 = ~x23 & n11828 ;
  assign n11830 = x23 | n11829 ;
  assign n11831 = ( ~n11828 & n11829 ) | ( ~n11828 & n11830 ) | ( n11829 & n11830 ) ;
  assign n11832 = ( n11810 & n11823 ) | ( n11810 & n11831 ) | ( n11823 & n11831 ) ;
  assign n11833 = n11810 | n11831 ;
  assign n11834 = n11823 | n11833 ;
  assign n11835 = ~n11832 & n11834 ;
  assign n11836 = n11654 & ~n11655 ;
  assign n11837 = ~n11665 & n11836 ;
  assign n11838 = n11665 | n11837 ;
  assign n11839 = ( ~n11836 & n11837 ) | ( ~n11836 & n11838 ) | ( n11837 & n11838 ) ;
  assign n11840 = n11835 & n11839 ;
  assign n11841 = n11832 | n11840 ;
  assign n11842 = n11669 | n11671 ;
  assign n11843 = n11668 | n11842 ;
  assign n11844 = ~n11672 & n11843 ;
  assign n11845 = n11841 & n11844 ;
  assign n11846 = n11841 | n11844 ;
  assign n11847 = ~n11845 & n11846 ;
  assign n11848 = n11839 & ~n11840 ;
  assign n11849 = ( n11835 & ~n11840 ) | ( n11835 & n11848 ) | ( ~n11840 & n11848 ) ;
  assign n11850 = n11694 | n11805 ;
  assign n11851 = ~n11806 & n11850 ;
  assign n11852 = ~n3596 & n4479 ;
  assign n11853 = n3504 & n4481 ;
  assign n11854 = n11852 | n11853 ;
  assign n11855 = ~n3431 & n4484 ;
  assign n11856 = n11854 | n11855 ;
  assign n11857 = n4487 | n11856 ;
  assign n11858 = ( ~n4798 & n11856 ) | ( ~n4798 & n11857 ) | ( n11856 & n11857 ) ;
  assign n11859 = ~x26 & n11858 ;
  assign n11860 = x26 | n11859 ;
  assign n11861 = ( ~n11858 & n11859 ) | ( ~n11858 & n11860 ) | ( n11859 & n11860 ) ;
  assign n11862 = n11851 & n11861 ;
  assign n11863 = n11851 & ~n11862 ;
  assign n11864 = ~n11851 & n11861 ;
  assign n11865 = n11863 | n11864 ;
  assign n11866 = ~n1014 & n4045 ;
  assign n11867 = ~n3255 & n4043 ;
  assign n11868 = n11866 | n11867 ;
  assign n11869 = n904 & n4048 ;
  assign n11870 = n11868 | n11869 ;
  assign n11871 = n4051 | n11870 ;
  assign n11872 = ( n4632 & n11870 ) | ( n4632 & n11871 ) | ( n11870 & n11871 ) ;
  assign n11873 = x29 & n11872 ;
  assign n11874 = x29 & ~n11873 ;
  assign n11875 = ( n11872 & ~n11873 ) | ( n11872 & n11874 ) | ( ~n11873 & n11874 ) ;
  assign n11876 = n778 & n4479 ;
  assign n11877 = ~n3596 & n4481 ;
  assign n11878 = n11876 | n11877 ;
  assign n11879 = n3504 & n4484 ;
  assign n11880 = n11878 | n11879 ;
  assign n11881 = n4487 | n11880 ;
  assign n11882 = ( ~n5040 & n11880 ) | ( ~n5040 & n11881 ) | ( n11880 & n11881 ) ;
  assign n11883 = ~x26 & n11882 ;
  assign n11884 = x26 | n11883 ;
  assign n11885 = ( ~n11882 & n11883 ) | ( ~n11882 & n11884 ) | ( n11883 & n11884 ) ;
  assign n11886 = n11761 & ~n11803 ;
  assign n11887 = n11804 | n11886 ;
  assign n11888 = ( n11875 & ~n11885 ) | ( n11875 & n11887 ) | ( ~n11885 & n11887 ) ;
  assign n11889 = ( ~n11875 & n11885 ) | ( ~n11875 & n11888 ) | ( n11885 & n11888 ) ;
  assign n11890 = ( ~n11887 & n11888 ) | ( ~n11887 & n11889 ) | ( n11888 & n11889 ) ;
  assign n11891 = ( n11875 & n11885 ) | ( n11875 & n11890 ) | ( n11885 & n11890 ) ;
  assign n11892 = n11865 & n11891 ;
  assign n11893 = n11862 | n11892 ;
  assign n11894 = n11812 & ~n11822 ;
  assign n11895 = ~n11811 & n11894 ;
  assign n11896 = n11823 | n11895 ;
  assign n11897 = n11893 & ~n11896 ;
  assign n11898 = ~n11893 & n11896 ;
  assign n11899 = n11897 | n11898 ;
  assign n11900 = ~n3634 & n4548 ;
  assign n11901 = ( n4546 & ~n11826 ) | ( n4546 & n11900 ) | ( ~n11826 & n11900 ) ;
  assign n11902 = n4554 | n11901 ;
  assign n11903 = ( n3726 & n11901 ) | ( n3726 & n11902 ) | ( n11901 & n11902 ) ;
  assign n11904 = x23 & n11903 ;
  assign n11905 = x23 & ~n11904 ;
  assign n11906 = ( n11903 & ~n11904 ) | ( n11903 & n11905 ) | ( ~n11904 & n11905 ) ;
  assign n11907 = ~n11899 & n11906 ;
  assign n11908 = n11897 | n11907 ;
  assign n11909 = n11849 & n11908 ;
  assign n11910 = n11849 | n11908 ;
  assign n11911 = ~n11909 & n11910 ;
  assign n11912 = n11899 & ~n11906 ;
  assign n11913 = n11907 | n11912 ;
  assign n11914 = ~n3634 & n4551 ;
  assign n11915 = ~n672 & n4548 ;
  assign n11916 = n11914 | n11915 ;
  assign n11917 = ~n589 & n4546 ;
  assign n11918 = n11916 | n11917 ;
  assign n11919 = n4554 | n11918 ;
  assign n11920 = ( ~n5092 & n11918 ) | ( ~n5092 & n11919 ) | ( n11918 & n11919 ) ;
  assign n11921 = ~x23 & n11920 ;
  assign n11922 = x23 | n11921 ;
  assign n11923 = ( ~n11920 & n11921 ) | ( ~n11920 & n11922 ) | ( n11921 & n11922 ) ;
  assign n11924 = n11865 | n11891 ;
  assign n11925 = ~n11892 & n11924 ;
  assign n11926 = ~n3431 & n4546 ;
  assign n11927 = ~n589 & n4548 ;
  assign n11928 = n11926 | n11927 ;
  assign n11929 = ~n672 & n4551 ;
  assign n11930 = n11928 | n11929 ;
  assign n11931 = n4554 | n11930 ;
  assign n11932 = ( ~n5353 & n11930 ) | ( ~n5353 & n11931 ) | ( n11930 & n11931 ) ;
  assign n11933 = ~x23 & n11932 ;
  assign n11934 = x23 | n11933 ;
  assign n11935 = ( ~n11932 & n11933 ) | ( ~n11932 & n11934 ) | ( n11933 & n11934 ) ;
  assign n11936 = n11791 | n11801 ;
  assign n11937 = ~n11802 & n11936 ;
  assign n11938 = n11774 | n11784 ;
  assign n11939 = ~n11785 & n11938 ;
  assign n11940 = ( ~n4449 & n11777 ) | ( ~n4449 & n11778 ) | ( n11777 & n11778 ) ;
  assign n11941 = n11783 | n11940 ;
  assign n11942 = n11776 & ~n11784 ;
  assign n11943 = n11941 & ~n11942 ;
  assign n11944 = n1327 & n3744 ;
  assign n11945 = n3104 & n3727 ;
  assign n11946 = n3178 & n3639 ;
  assign n11947 = n11945 | n11946 ;
  assign n11948 = n3636 | n11947 ;
  assign n11949 = ( n4501 & n11947 ) | ( n4501 & n11948 ) | ( n11947 & n11948 ) ;
  assign n11950 = n11944 | n11949 ;
  assign n11951 = ~n11943 & n11950 ;
  assign n11952 = n11943 & ~n11950 ;
  assign n11953 = n11951 | n11952 ;
  assign n11954 = ~n1151 & n4043 ;
  assign n11955 = n1233 & n4045 ;
  assign n11956 = n11954 | n11955 ;
  assign n11957 = n3349 & n4048 ;
  assign n11958 = n11956 | n11957 ;
  assign n11959 = n4051 | n11958 ;
  assign n11960 = ( n4518 & n11958 ) | ( n4518 & n11959 ) | ( n11958 & n11959 ) ;
  assign n11961 = x29 & n11960 ;
  assign n11962 = x29 & ~n11961 ;
  assign n11963 = ( n11960 & ~n11961 ) | ( n11960 & n11962 ) | ( ~n11961 & n11962 ) ;
  assign n11964 = ~n11953 & n11963 ;
  assign n11965 = n11951 | n11964 ;
  assign n11966 = n11939 & n11965 ;
  assign n11967 = n11939 | n11965 ;
  assign n11968 = ~n11966 & n11967 ;
  assign n11969 = n1233 & n4043 ;
  assign n11970 = n3349 & n4045 ;
  assign n11971 = n11969 | n11970 ;
  assign n11972 = ~n3255 & n4048 ;
  assign n11973 = n11971 | n11972 ;
  assign n11974 = n4051 | n11973 ;
  assign n11975 = ( ~n4470 & n11973 ) | ( ~n4470 & n11974 ) | ( n11973 & n11974 ) ;
  assign n11976 = ~x29 & n11975 ;
  assign n11977 = x29 | n11976 ;
  assign n11978 = ( ~n11975 & n11976 ) | ( ~n11975 & n11977 ) | ( n11976 & n11977 ) ;
  assign n11979 = n11968 & n11978 ;
  assign n11980 = n11966 | n11979 ;
  assign n11981 = n904 & n4479 ;
  assign n11982 = n778 & n4481 ;
  assign n11983 = n11981 | n11982 ;
  assign n11984 = ~n3596 & n4484 ;
  assign n11985 = n11983 | n11984 ;
  assign n11986 = n4487 | n11985 ;
  assign n11987 = ( ~n4649 & n11985 ) | ( ~n4649 & n11986 ) | ( n11985 & n11986 ) ;
  assign n11988 = ~x26 & n11987 ;
  assign n11989 = x26 | n11988 ;
  assign n11990 = ( ~n11987 & n11988 ) | ( ~n11987 & n11989 ) | ( n11988 & n11989 ) ;
  assign n11991 = ( n11937 & n11980 ) | ( n11937 & n11990 ) | ( n11980 & n11990 ) ;
  assign n11992 = ( n11890 & ~n11935 ) | ( n11890 & n11991 ) | ( ~n11935 & n11991 ) ;
  assign n11993 = ( ~n11890 & n11935 ) | ( ~n11890 & n11992 ) | ( n11935 & n11992 ) ;
  assign n11994 = ( n11923 & n11925 ) | ( n11923 & n11993 ) | ( n11925 & n11993 ) ;
  assign n11995 = ~n11913 & n11994 ;
  assign n11996 = n11913 & ~n11994 ;
  assign n11997 = n11995 | n11996 ;
  assign n11998 = n4776 | n4784 ;
  assign n11999 = ~n3634 & n11998 ;
  assign n12000 = n672 & n4776 ;
  assign n12001 = ( ~n672 & n11999 ) | ( ~n672 & n12000 ) | ( n11999 & n12000 ) ;
  assign n12002 = ( ~n3619 & n11999 ) | ( ~n3619 & n12001 ) | ( n11999 & n12001 ) ;
  assign n12003 = ~x20 & n12002 ;
  assign n12004 = x20 | n12003 ;
  assign n12005 = ( ~n12002 & n12003 ) | ( ~n12002 & n12004 ) | ( n12003 & n12004 ) ;
  assign n12006 = n11968 & ~n11979 ;
  assign n12007 = ~n11968 & n11978 ;
  assign n12008 = ~n1014 & n4479 ;
  assign n12009 = n904 & n4481 ;
  assign n12010 = n12008 | n12009 ;
  assign n12011 = n778 & n4484 ;
  assign n12012 = n12010 | n12011 ;
  assign n12013 = n4487 | n12012 ;
  assign n12014 = ( ~n4535 & n12012 ) | ( ~n4535 & n12013 ) | ( n12012 & n12013 ) ;
  assign n12015 = ~x26 & n12014 ;
  assign n12016 = x26 | n12015 ;
  assign n12017 = ( ~n12014 & n12015 ) | ( ~n12014 & n12016 ) | ( n12015 & n12016 ) ;
  assign n12018 = ( n12006 & n12007 ) | ( n12006 & n12017 ) | ( n12007 & n12017 ) ;
  assign n12019 = n12007 | n12017 ;
  assign n12020 = n12006 | n12019 ;
  assign n12021 = ~n12018 & n12020 ;
  assign n12022 = n4723 | n4736 ;
  assign n12023 = ~n1014 & n4481 ;
  assign n12024 = ~n3255 & n4479 ;
  assign n12025 = n12023 | n12024 ;
  assign n12026 = n904 & n4484 ;
  assign n12027 = n12025 | n12026 ;
  assign n12028 = n4487 | n12027 ;
  assign n12029 = ( n4632 & n12027 ) | ( n4632 & n12028 ) | ( n12027 & n12028 ) ;
  assign n12030 = x26 & n12029 ;
  assign n12031 = x26 & ~n12030 ;
  assign n12032 = ( n12029 & ~n12030 ) | ( n12029 & n12031 ) | ( ~n12030 & n12031 ) ;
  assign n12033 = ( n11953 & ~n11963 ) | ( n11953 & n12022 ) | ( ~n11963 & n12022 ) ;
  assign n12034 = ( ~n11953 & n11963 ) | ( ~n11953 & n12033 ) | ( n11963 & n12033 ) ;
  assign n12035 = ( ~n12022 & n12033 ) | ( ~n12022 & n12034 ) | ( n12033 & n12034 ) ;
  assign n12036 = n12032 | n12035 ;
  assign n12037 = ~n12032 & n12036 ;
  assign n12038 = ( ~n12035 & n12036 ) | ( ~n12035 & n12037 ) | ( n12036 & n12037 ) ;
  assign n12039 = ( n12022 & n12032 ) | ( n12022 & n12038 ) | ( n12032 & n12038 ) ;
  assign n12040 = n12021 & n12039 ;
  assign n12041 = n12018 | n12040 ;
  assign n12042 = n3504 & n4546 ;
  assign n12043 = ~n3431 & n4548 ;
  assign n12044 = n12042 | n12043 ;
  assign n12045 = ~n589 & n4551 ;
  assign n12046 = n12044 | n12045 ;
  assign n12047 = n4554 | n12046 ;
  assign n12048 = ( n4765 & n12046 ) | ( n4765 & n12047 ) | ( n12046 & n12047 ) ;
  assign n12049 = x23 & n12048 ;
  assign n12050 = x23 & ~n12049 ;
  assign n12051 = ( n12048 & ~n12049 ) | ( n12048 & n12050 ) | ( ~n12049 & n12050 ) ;
  assign n12052 = ( n11937 & n11990 ) | ( n11937 & ~n11991 ) | ( n11990 & ~n11991 ) ;
  assign n12053 = ( n11980 & ~n11991 ) | ( n11980 & n12052 ) | ( ~n11991 & n12052 ) ;
  assign n12054 = ( n12041 & n12051 ) | ( n12041 & n12053 ) | ( n12051 & n12053 ) ;
  assign n12055 = n12005 & n12054 ;
  assign n12056 = ( ~n11991 & n11992 ) | ( ~n11991 & n11993 ) | ( n11992 & n11993 ) ;
  assign n12057 = n12005 | n12054 ;
  assign n12058 = ~n12055 & n12057 ;
  assign n12059 = ~n12056 & n12058 ;
  assign n12060 = n12055 | n12059 ;
  assign n12061 = ( n11923 & ~n11925 ) | ( n11923 & n11993 ) | ( ~n11925 & n11993 ) ;
  assign n12062 = ( ~n11923 & n11925 ) | ( ~n11923 & n12061 ) | ( n11925 & n12061 ) ;
  assign n12063 = ( ~n11993 & n12061 ) | ( ~n11993 & n12062 ) | ( n12061 & n12062 ) ;
  assign n12064 = n12060 & n12063 ;
  assign n12065 = n12060 | n12063 ;
  assign n12066 = ~n12064 & n12065 ;
  assign n12067 = n12056 | n12059 ;
  assign n12068 = ( ~n12058 & n12059 ) | ( ~n12058 & n12067 ) | ( n12059 & n12067 ) ;
  assign n12069 = n12021 | n12039 ;
  assign n12070 = ~n12040 & n12069 ;
  assign n12071 = ~n3596 & n4546 ;
  assign n12072 = n3504 & n4548 ;
  assign n12073 = n12071 | n12072 ;
  assign n12074 = ~n3431 & n4551 ;
  assign n12075 = n12073 | n12074 ;
  assign n12076 = n4554 | n12075 ;
  assign n12077 = ( ~n4798 & n12075 ) | ( ~n4798 & n12076 ) | ( n12075 & n12076 ) ;
  assign n12078 = ~x23 & n12077 ;
  assign n12079 = x23 | n12078 ;
  assign n12080 = ( ~n12077 & n12078 ) | ( ~n12077 & n12079 ) | ( n12078 & n12079 ) ;
  assign n12081 = n12070 & n12080 ;
  assign n12082 = n12070 & ~n12081 ;
  assign n12083 = ~n12070 & n12080 ;
  assign n12084 = n778 & n4546 ;
  assign n12085 = ~n3596 & n4548 ;
  assign n12086 = n12084 | n12085 ;
  assign n12087 = n3504 & n4551 ;
  assign n12088 = n12086 | n12087 ;
  assign n12089 = n4554 | n12088 ;
  assign n12090 = ( ~n5040 & n12088 ) | ( ~n5040 & n12089 ) | ( n12088 & n12089 ) ;
  assign n12091 = ~x23 & n12090 ;
  assign n12092 = x23 | n12091 ;
  assign n12093 = ( ~n12090 & n12091 ) | ( ~n12090 & n12092 ) | ( n12091 & n12092 ) ;
  assign n12094 = ( ~n4753 & n12038 ) | ( ~n4753 & n12093 ) | ( n12038 & n12093 ) ;
  assign n12095 = ( n4753 & ~n12038 ) | ( n4753 & n12094 ) | ( ~n12038 & n12094 ) ;
  assign n12096 = ( n12082 & n12083 ) | ( n12082 & n12095 ) | ( n12083 & n12095 ) ;
  assign n12097 = n12081 | n12096 ;
  assign n12098 = ~n3634 & n4778 ;
  assign n12099 = ( n4776 & ~n12000 ) | ( n4776 & n12098 ) | ( ~n12000 & n12098 ) ;
  assign n12100 = n4784 | n12099 ;
  assign n12101 = ( n3726 & n12099 ) | ( n3726 & n12100 ) | ( n12099 & n12100 ) ;
  assign n12102 = x20 & n12101 ;
  assign n12103 = x20 & ~n12102 ;
  assign n12104 = ( n12101 & ~n12102 ) | ( n12101 & n12103 ) | ( ~n12102 & n12103 ) ;
  assign n12105 = ( ~n12041 & n12051 ) | ( ~n12041 & n12053 ) | ( n12051 & n12053 ) ;
  assign n12106 = ( n12041 & ~n12053 ) | ( n12041 & n12105 ) | ( ~n12053 & n12105 ) ;
  assign n12107 = ( ~n12051 & n12105 ) | ( ~n12051 & n12106 ) | ( n12105 & n12106 ) ;
  assign n12108 = ( n12097 & n12104 ) | ( n12097 & n12107 ) | ( n12104 & n12107 ) ;
  assign n12109 = ~n12068 & n12108 ;
  assign n12110 = n12068 & ~n12108 ;
  assign n12111 = n12109 | n12110 ;
  assign n12112 = ~n3634 & n4781 ;
  assign n12113 = ~n672 & n4778 ;
  assign n12114 = n12112 | n12113 ;
  assign n12115 = ~n589 & n4776 ;
  assign n12116 = n12114 | n12115 ;
  assign n12117 = n4784 | n12116 ;
  assign n12118 = ( ~n5092 & n12116 ) | ( ~n5092 & n12117 ) | ( n12116 & n12117 ) ;
  assign n12119 = ~x20 & n12118 ;
  assign n12120 = x20 | n12119 ;
  assign n12121 = ( ~n12118 & n12119 ) | ( ~n12118 & n12120 ) | ( n12119 & n12120 ) ;
  assign n12122 = ( ~n12093 & n12094 ) | ( ~n12093 & n12095 ) | ( n12094 & n12095 ) ;
  assign n12123 = ( n4659 & n4660 ) | ( n4659 & n4755 ) | ( n4660 & n4755 ) ;
  assign n12124 = ~n3431 & n4776 ;
  assign n12125 = ~n589 & n4778 ;
  assign n12126 = n12124 | n12125 ;
  assign n12127 = ~n672 & n4781 ;
  assign n12128 = n12126 | n12127 ;
  assign n12129 = n4784 | n12128 ;
  assign n12130 = ( ~n5353 & n12128 ) | ( ~n5353 & n12129 ) | ( n12128 & n12129 ) ;
  assign n12131 = ~x20 & n12130 ;
  assign n12132 = x20 | n12131 ;
  assign n12133 = ( ~n12130 & n12131 ) | ( ~n12130 & n12132 ) | ( n12131 & n12132 ) ;
  assign n12134 = ( n12122 & ~n12123 ) | ( n12122 & n12133 ) | ( ~n12123 & n12133 ) ;
  assign n12135 = ( ~n12122 & n12123 ) | ( ~n12122 & n12134 ) | ( n12123 & n12134 ) ;
  assign n12136 = n12121 & n12135 ;
  assign n12137 = n12121 | n12135 ;
  assign n12138 = ~n12136 & n12137 ;
  assign n12139 = n12083 | n12095 ;
  assign n12140 = n12082 | n12139 ;
  assign n12141 = ~n12096 & n12140 ;
  assign n12142 = n12138 & n12141 ;
  assign n12143 = n12136 | n12142 ;
  assign n12144 = ( n12097 & n12104 ) | ( n12097 & ~n12107 ) | ( n12104 & ~n12107 ) ;
  assign n12145 = ( ~n12097 & n12107 ) | ( ~n12097 & n12144 ) | ( n12107 & n12144 ) ;
  assign n12146 = ( ~n12104 & n12144 ) | ( ~n12104 & n12145 ) | ( n12144 & n12145 ) ;
  assign n12147 = n12143 & n12146 ;
  assign n12148 = n12143 | n12146 ;
  assign n12149 = ~n12147 & n12148 ;
  assign n12150 = n12138 | n12141 ;
  assign n12151 = ~n12142 & n12150 ;
  assign n12152 = n5069 | n5074 ;
  assign n12153 = ~n3634 & n12152 ;
  assign n12154 = ( ~n672 & n5072 ) | ( ~n672 & n12153 ) | ( n5072 & n12153 ) ;
  assign n12155 = ( ~n3619 & n12153 ) | ( ~n3619 & n12154 ) | ( n12153 & n12154 ) ;
  assign n12156 = ~x17 & n12155 ;
  assign n12157 = x17 | n12156 ;
  assign n12158 = ( ~n12155 & n12156 ) | ( ~n12155 & n12157 ) | ( n12156 & n12157 ) ;
  assign n12159 = n4759 | n4790 ;
  assign n12160 = n12158 & n12159 ;
  assign n12161 = ( ~n12133 & n12134 ) | ( ~n12133 & n12135 ) | ( n12134 & n12135 ) ;
  assign n12162 = n12158 | n12159 ;
  assign n12163 = ~n12160 & n12162 ;
  assign n12164 = ~n12161 & n12163 ;
  assign n12165 = n12160 | n12164 ;
  assign n12166 = n12151 & n12165 ;
  assign n12167 = n12151 | n12165 ;
  assign n12168 = ~n12166 & n12167 ;
  assign n12169 = n12161 | n12164 ;
  assign n12170 = ( ~n12163 & n12164 ) | ( ~n12163 & n12169 ) | ( n12164 & n12169 ) ;
  assign n12171 = ( n5056 & n5057 ) | ( n5056 & n5079 ) | ( n5057 & n5079 ) ;
  assign n12172 = ~n12170 & n12171 ;
  assign n12173 = n12170 & ~n12171 ;
  assign n12174 = n12172 | n12173 ;
  assign n12175 = n5375 & ~n12174 ;
  assign n12176 = n12172 | n12175 ;
  assign n12177 = n12168 & n12176 ;
  assign n12178 = n12166 | n12177 ;
  assign n12179 = n12149 & n12178 ;
  assign n12180 = n12147 | n12179 ;
  assign n12181 = ~n12111 & n12180 ;
  assign n12182 = n12109 | n12181 ;
  assign n12183 = n12066 & n12182 ;
  assign n12184 = n12064 | n12183 ;
  assign n12185 = ~n11997 & n12184 ;
  assign n12186 = n11995 | n12185 ;
  assign n12187 = n11911 & n12186 ;
  assign n12188 = n11909 | n12187 ;
  assign n12189 = n11847 & n12188 ;
  assign n12190 = n11845 | n12189 ;
  assign n12191 = n11679 & n12190 ;
  assign n12192 = n11677 | n12191 ;
  assign n12193 = n11630 & n12192 ;
  assign n12194 = n11627 | n12193 ;
  assign n12195 = n11472 | n11499 ;
  assign n12196 = ~n11500 & n12195 ;
  assign n12197 = n12194 & n12196 ;
  assign n12198 = n11500 | n12197 ;
  assign n12199 = ~n11470 & n12198 ;
  assign n12200 = n11468 | n12199 ;
  assign n12201 = ~n11126 & n12200 ;
  assign n12202 = n11124 | n12201 ;
  assign n12203 = n11028 & n12202 ;
  assign n12204 = n11025 | n12203 ;
  assign n12205 = ~n10998 & n12204 ;
  assign n12206 = n10996 | n12205 ;
  assign n12207 = n12168 & ~n12173 ;
  assign n12208 = n12166 | n12207 ;
  assign n12209 = n12149 & n12208 ;
  assign n12210 = n12147 | n12209 ;
  assign n12211 = ~n12111 & n12210 ;
  assign n12212 = n12109 | n12211 ;
  assign n12213 = n12066 & n12212 ;
  assign n12214 = n12064 | n12213 ;
  assign n12215 = ~n11997 & n12214 ;
  assign n12216 = n11995 | n12215 ;
  assign n12217 = n11911 & n12216 ;
  assign n12218 = n11909 | n12217 ;
  assign n12219 = n11847 & n12218 ;
  assign n12220 = n11845 | n12219 ;
  assign n12221 = n11679 & n12220 ;
  assign n12222 = n11677 | n12221 ;
  assign n12223 = n11630 & n12222 ;
  assign n12224 = n11627 | n12223 ;
  assign n12225 = n12196 & n12224 ;
  assign n12226 = n11500 | n12225 ;
  assign n12227 = ~n11470 & n12226 ;
  assign n12228 = n11468 | n12227 ;
  assign n12229 = ~n11126 & n12228 ;
  assign n12230 = n11124 | n12229 ;
  assign n12231 = n11028 & n12230 ;
  assign n12232 = n11025 | n12231 ;
  assign n12233 = ~n10998 & n12232 ;
  assign n12234 = n10996 | n12233 ;
  assign n12235 = ( n10849 & n12206 ) | ( n10849 & n12234 ) | ( n12206 & n12234 ) ;
  assign n12236 = ~n3740 & n12235 ;
  assign n12237 = n3738 | n12236 ;
  assign n12238 = n242 | n266 ;
  assign n12239 = n1329 | n12238 ;
  assign n12240 = n151 | n12239 ;
  assign n12241 = n468 | n636 ;
  assign n12242 = n419 | n12241 ;
  assign n12243 = n62 | n334 ;
  assign n12244 = n441 | n12243 ;
  assign n12245 = n12242 | n12244 ;
  assign n12246 = n1632 | n12245 ;
  assign n12247 = ( ~n11090 & n12240 ) | ( ~n11090 & n12246 ) | ( n12240 & n12246 ) ;
  assign n12248 = n11090 | n12247 ;
  assign n12249 = n3020 | n12248 ;
  assign n12250 = n2400 | n2703 ;
  assign n12251 = n2154 | n12250 ;
  assign n12252 = n284 | n12251 ;
  assign n12253 = n476 | n12252 ;
  assign n12254 = n619 | n12253 ;
  assign n12255 = n12249 | n12254 ;
  assign n12256 = n359 | n503 ;
  assign n12257 = n134 | n12256 ;
  assign n12258 = n108 | n12257 ;
  assign n12259 = n923 | n1240 ;
  assign n12260 = n11718 | n12259 ;
  assign n12261 = n279 | n887 ;
  assign n12262 = n315 | n12261 ;
  assign n12263 = n12260 | n12262 ;
  assign n12264 = n252 | n309 ;
  assign n12265 = n190 | n12264 ;
  assign n12266 = n94 | n12265 ;
  assign n12267 = n129 | n12266 ;
  assign n12268 = n12263 | n12267 ;
  assign n12269 = n1912 | n5753 ;
  assign n12270 = n844 | n12269 ;
  assign n12271 = n5555 | n12270 ;
  assign n12272 = n11072 | n12271 ;
  assign n12273 = n12268 | n12272 ;
  assign n12274 = n2977 | n12273 ;
  assign n12275 = n11069 | n12274 ;
  assign n12276 = n12258 | n12275 ;
  assign n12277 = n12255 | n12276 ;
  assign n12278 = n600 | n603 ;
  assign n12279 = n808 | n890 ;
  assign n12280 = n1352 | n12279 ;
  assign n12281 = n1034 | n12280 ;
  assign n12282 = n278 | n12281 ;
  assign n12283 = n1989 | n12282 ;
  assign n12284 = n520 | n12283 ;
  assign n12285 = n180 | n12284 ;
  assign n12286 = n12278 | n12285 ;
  assign n12287 = n609 | n12286 ;
  assign n12288 = n12277 | n12287 ;
  assign n12289 = n610 | n12288 ;
  assign n12290 = n660 | n661 ;
  assign n12291 = n387 | n422 ;
  assign n12292 = n205 | n554 ;
  assign n12293 = n12291 | n12292 ;
  assign n12294 = n12290 | n12293 ;
  assign n12295 = n544 & ~n12294 ;
  assign n12296 = n215 | n669 ;
  assign n12297 = n58 | n12296 ;
  assign n12298 = n12295 & ~n12297 ;
  assign n12299 = n466 & n12298 ;
  assign n12300 = n12289 & n12299 ;
  assign n12301 = n466 | n12298 ;
  assign n12302 = ~n12299 & n12301 ;
  assign n12303 = n3648 & ~n12302 ;
  assign n12304 = n3648 & ~n12303 ;
  assign n12305 = n3648 | n12302 ;
  assign n12306 = ~n12304 & n12305 ;
  assign n12307 = ~n12303 & n12306 ;
  assign n12308 = n12289 | n12299 ;
  assign n12309 = ~n12307 & n12308 ;
  assign n12310 = ~n12300 & n12309 ;
  assign n12311 = n12289 & n12310 ;
  assign n12312 = ( n12303 & n12307 ) | ( n12303 & n12310 ) | ( n12307 & n12310 ) ;
  assign n12313 = n12289 & n12312 ;
  assign n12314 = ( n12237 & n12311 ) | ( n12237 & n12313 ) | ( n12311 & n12313 ) ;
  assign n12315 = ( n12237 & n12310 ) | ( n12237 & n12312 ) | ( n12310 & n12312 ) ;
  assign n12316 = n12308 & ~n12315 ;
  assign n12317 = ~n12289 & n12316 ;
  assign n12318 = n12314 | n12317 ;
  assign n12319 = n7277 | n7280 ;
  assign n12320 = ~n12314 & n12319 ;
  assign n12321 = n5384 | n12319 ;
  assign n12322 = ( ~n12318 & n12320 ) | ( ~n12318 & n12321 ) | ( n12320 & n12321 ) ;
  assign n12323 = n39 | n12322 ;
  assign n12324 = n3740 & ~n12235 ;
  assign n12325 = n12236 | n12324 ;
  assign n12326 = n12237 & ~n12306 ;
  assign n12327 = ~n12237 & n12306 ;
  assign n12328 = n12326 | n12327 ;
  assign n12329 = n12325 | n12328 ;
  assign n12330 = n12325 & n12328 ;
  assign n12331 = n12329 & ~n12330 ;
  assign n12332 = ( n10849 & n12205 ) | ( n10849 & n12233 ) | ( n12205 & n12233 ) ;
  assign n12333 = ( n10849 & n12204 ) | ( n10849 & n12232 ) | ( n12204 & n12232 ) ;
  assign n12334 = n10998 & ~n12333 ;
  assign n12335 = n12332 | n12334 ;
  assign n12336 = n12325 | n12335 ;
  assign n12337 = ( n10849 & n12197 ) | ( n10849 & n12225 ) | ( n12197 & n12225 ) ;
  assign n12338 = ( n10849 & n12194 ) | ( n10849 & n12224 ) | ( n12194 & n12224 ) ;
  assign n12339 = n12196 | n12338 ;
  assign n12340 = ~n12337 & n12339 ;
  assign n12341 = ( n10849 & n12199 ) | ( n10849 & n12227 ) | ( n12199 & n12227 ) ;
  assign n12342 = ( n10849 & n12198 ) | ( n10849 & n12226 ) | ( n12198 & n12226 ) ;
  assign n12343 = n11470 & ~n12342 ;
  assign n12344 = n12341 | n12343 ;
  assign n12345 = n12340 & ~n12344 ;
  assign n12346 = ~n12340 & n12344 ;
  assign n12347 = n12345 | n12346 ;
  assign n12348 = ( n10849 & n12187 ) | ( n10849 & n12217 ) | ( n12187 & n12217 ) ;
  assign n12349 = ( n10849 & n12186 ) | ( n10849 & n12216 ) | ( n12186 & n12216 ) ;
  assign n12350 = n11911 | n12349 ;
  assign n12351 = ~n12348 & n12350 ;
  assign n12352 = ( n10849 & n12189 ) | ( n10849 & n12219 ) | ( n12189 & n12219 ) ;
  assign n12353 = ( n10849 & n12188 ) | ( n10849 & n12218 ) | ( n12188 & n12218 ) ;
  assign n12354 = n11847 | n12353 ;
  assign n12355 = ~n12352 & n12354 ;
  assign n12356 = n12351 & n12355 ;
  assign n12357 = ( n10849 & n12181 ) | ( n10849 & n12211 ) | ( n12181 & n12211 ) ;
  assign n12358 = ( n10849 & n12180 ) | ( n10849 & n12210 ) | ( n12180 & n12210 ) ;
  assign n12359 = n12111 & ~n12358 ;
  assign n12360 = n12357 | n12359 ;
  assign n12361 = ( n10849 & n12183 ) | ( n10849 & n12213 ) | ( n12183 & n12213 ) ;
  assign n12362 = ( n10849 & n12182 ) | ( n10849 & n12212 ) | ( n12182 & n12212 ) ;
  assign n12363 = n12066 | n12362 ;
  assign n12364 = ~n12361 & n12363 ;
  assign n12365 = ~n12360 & n12364 ;
  assign n12366 = n12360 & ~n12364 ;
  assign n12367 = n12365 | n12366 ;
  assign n12368 = ( n10849 & ~n12174 ) | ( n10849 & n12175 ) | ( ~n12174 & n12175 ) ;
  assign n12369 = ~n5375 & n12174 ;
  assign n12370 = ~n10849 & n12369 ;
  assign n12371 = n12368 | n12370 ;
  assign n12372 = ( n10849 & n12177 ) | ( n10849 & n12207 ) | ( n12177 & n12207 ) ;
  assign n12373 = ( n10849 & ~n12173 ) | ( n10849 & n12176 ) | ( ~n12173 & n12176 ) ;
  assign n12374 = n12168 | n12373 ;
  assign n12375 = ~n12372 & n12374 ;
  assign n12376 = n12371 & ~n12375 ;
  assign n12377 = n5377 | n10848 ;
  assign n12378 = ~n10849 & n12377 ;
  assign n12379 = ~n12371 & n12378 ;
  assign n12380 = ( n10455 & n10828 ) | ( n10455 & n10842 ) | ( n10828 & n10842 ) ;
  assign n12381 = ( n10455 & n10827 ) | ( n10455 & n10841 ) | ( n10827 & n10841 ) ;
  assign n12382 = n10636 | n12381 ;
  assign n12383 = ~n12380 & n12382 ;
  assign n12384 = ( n10455 & n10830 ) | ( n10455 & n10844 ) | ( n10830 & n10844 ) ;
  assign n12385 = ( n10455 & n10829 ) | ( n10455 & n10843 ) | ( n10829 & n10843 ) ;
  assign n12386 = n10555 | n12385 ;
  assign n12387 = ~n12384 & n12386 ;
  assign n12388 = n12383 & n12387 ;
  assign n12389 = ( n10455 & n10826 ) | ( n10455 & n10840 ) | ( n10826 & n10840 ) ;
  assign n12390 = ( n10455 & n10825 ) | ( n10455 & n10839 ) | ( n10825 & n10839 ) ;
  assign n12391 = n10700 | n12390 ;
  assign n12392 = ~n12389 & n12391 ;
  assign n12393 = n12383 | n12392 ;
  assign n12394 = n12383 | n12387 ;
  assign n12395 = n12393 & n12394 ;
  assign n12396 = ~n12388 & n12395 ;
  assign n12397 = n12383 & n12392 ;
  assign n12398 = ( n10455 & n10824 ) | ( n10455 & n10838 ) | ( n10824 & n10838 ) ;
  assign n12399 = ( n10455 & n10823 ) | ( n10455 & n10837 ) | ( n10823 & n10837 ) ;
  assign n12400 = n10759 | n12399 ;
  assign n12401 = ~n12398 & n12400 ;
  assign n12402 = n12392 & n12401 ;
  assign n12403 = n12393 & ~n12397 ;
  assign n12404 = n12402 & n12403 ;
  assign n12405 = ( n12396 & n12397 ) | ( n12396 & n12404 ) | ( n12397 & n12404 ) ;
  assign n12406 = n12392 | n12401 ;
  assign n12407 = ~n12402 & n12406 ;
  assign n12408 = ( n10455 & n10820 ) | ( n10455 & n10834 ) | ( n10820 & n10834 ) ;
  assign n12409 = ( n10455 & n10817 ) | ( n10455 & n10833 ) | ( n10817 & n10833 ) ;
  assign n12410 = n10819 | n12409 ;
  assign n12411 = ~n12408 & n12410 ;
  assign n12412 = ( n10455 & n10822 ) | ( n10455 & n10836 ) | ( n10822 & n10836 ) ;
  assign n12413 = ( n10455 & n10821 ) | ( n10455 & n10835 ) | ( n10821 & n10835 ) ;
  assign n12414 = n10795 | n12413 ;
  assign n12415 = ~n12412 & n12414 ;
  assign n12416 = n12411 | n12415 ;
  assign n12417 = ( n10455 & ~n10813 ) | ( n10455 & n10816 ) | ( ~n10813 & n10816 ) ;
  assign n12418 = ( n10813 & ~n10816 ) | ( n10813 & n12417 ) | ( ~n10816 & n12417 ) ;
  assign n12419 = ( ~n10455 & n12417 ) | ( ~n10455 & n12418 ) | ( n12417 & n12418 ) ;
  assign n12420 = n12411 | n12419 ;
  assign n12421 = n12411 & n12419 ;
  assign n12422 = n7782 & ~n10453 ;
  assign n12423 = n10454 | n12422 ;
  assign n12424 = n12419 & ~n12423 ;
  assign n12425 = n12420 & ~n12421 ;
  assign n12426 = n12424 & n12425 ;
  assign n12427 = n12421 | n12426 ;
  assign n12428 = ~n12419 & n12423 ;
  assign n12429 = n12424 | n12428 ;
  assign n12430 = ( n10420 & n10449 ) | ( n10420 & n10451 ) | ( n10449 & n10451 ) ;
  assign n12431 = ( n10420 & ~n10445 ) | ( n10420 & n10448 ) | ( ~n10445 & n10448 ) ;
  assign n12432 = n10440 | n12431 ;
  assign n12433 = ~n12430 & n12432 ;
  assign n12434 = ~n12423 & n12433 ;
  assign n12435 = ( n10420 & ~n10446 ) | ( n10420 & n10447 ) | ( ~n10446 & n10447 ) ;
  assign n12436 = ~n9257 & n10446 ;
  assign n12437 = ~n10420 & n12436 ;
  assign n12438 = n12435 | n12437 ;
  assign n12439 = n9259 | n10419 ;
  assign n12440 = ~n10420 & n12439 ;
  assign n12441 = ~n12438 & n12440 ;
  assign n12442 = n12438 & ~n12440 ;
  assign n12443 = ( n10405 & n10416 ) | ( n10405 & n10417 ) | ( n10416 & n10417 ) ;
  assign n12444 = n10402 | n10416 ;
  assign n12445 = n10405 | n12444 ;
  assign n12446 = ~n12443 & n12445 ;
  assign n12447 = n12440 & n12446 ;
  assign n12448 = n12440 | n12446 ;
  assign n12449 = ~n12447 & n12448 ;
  assign n12450 = n9793 | n10404 ;
  assign n12451 = n10374 | n12450 ;
  assign n12452 = ~n10405 & n12451 ;
  assign n12453 = n9795 | n10373 ;
  assign n12454 = ~n10374 & n12453 ;
  assign n12455 = n9811 & ~n10371 ;
  assign n12456 = n10372 | n12455 ;
  assign n12457 = n12454 & ~n12456 ;
  assign n12458 = n9826 | n10369 ;
  assign n12459 = ~n10370 & n12458 ;
  assign n12460 = ~n12456 & n12459 ;
  assign n12461 = n12456 & ~n12459 ;
  assign n12462 = n12460 | n12461 ;
  assign n12463 = ( ~n9841 & n9855 ) | ( ~n9841 & n10368 ) | ( n9855 & n10368 ) ;
  assign n12464 = n9841 & ~n9854 ;
  assign n12465 = ~n10368 & n12464 ;
  assign n12466 = n12463 | n12465 ;
  assign n12467 = n9858 & ~n10367 ;
  assign n12468 = n10368 | n12467 ;
  assign n12469 = ~n12466 & n12468 ;
  assign n12470 = ~n12459 & n12469 ;
  assign n12471 = n12466 | n12470 ;
  assign n12472 = n12462 | n12471 ;
  assign n12473 = ~n12460 & n12472 ;
  assign n12474 = ~n12454 & n12456 ;
  assign n12475 = n12457 | n12474 ;
  assign n12476 = n12473 | n12475 ;
  assign n12477 = ~n12457 & n12476 ;
  assign n12478 = ( n12452 & n12454 ) | ( n12452 & ~n12477 ) | ( n12454 & ~n12477 ) ;
  assign n12479 = ( n12446 & n12452 ) | ( n12446 & n12478 ) | ( n12452 & n12478 ) ;
  assign n12480 = n12449 & n12479 ;
  assign n12481 = ( ~n12442 & n12447 ) | ( ~n12442 & n12480 ) | ( n12447 & n12480 ) ;
  assign n12482 = n12441 | n12481 ;
  assign n12483 = ( n12433 & ~n12438 ) | ( n12433 & n12482 ) | ( ~n12438 & n12482 ) ;
  assign n12484 = n12423 & ~n12433 ;
  assign n12485 = n12434 | n12484 ;
  assign n12486 = n12483 & ~n12485 ;
  assign n12487 = ( ~n12429 & n12434 ) | ( ~n12429 & n12486 ) | ( n12434 & n12486 ) ;
  assign n12488 = ( n12420 & n12427 ) | ( n12420 & n12487 ) | ( n12427 & n12487 ) ;
  assign n12489 = n12416 & n12488 ;
  assign n12490 = n12411 & n12415 ;
  assign n12491 = n12401 & n12415 ;
  assign n12492 = n12490 | n12491 ;
  assign n12493 = n12401 | n12415 ;
  assign n12494 = ( n12489 & n12492 ) | ( n12489 & n12493 ) | ( n12492 & n12493 ) ;
  assign n12495 = n12407 & n12494 ;
  assign n12496 = ( n12396 & n12405 ) | ( n12396 & n12495 ) | ( n12405 & n12495 ) ;
  assign n12497 = n12388 | n12496 ;
  assign n12498 = n12371 & ~n12378 ;
  assign n12499 = n12379 | n12498 ;
  assign n12500 = ( n10455 & n10831 ) | ( n10455 & n10845 ) | ( n10831 & n10845 ) ;
  assign n12501 = n10457 & ~n12500 ;
  assign n12502 = n10847 | n12501 ;
  assign n12503 = n12378 & ~n12502 ;
  assign n12504 = ~n12378 & n12502 ;
  assign n12505 = n12503 | n12504 ;
  assign n12506 = ~n12387 & n12502 ;
  assign n12507 = n12505 | n12506 ;
  assign n12508 = ~n12503 & n12507 ;
  assign n12509 = n12499 | n12508 ;
  assign n12510 = n12387 & ~n12502 ;
  assign n12511 = ~n12505 & n12510 ;
  assign n12512 = n12503 | n12511 ;
  assign n12513 = ~n12499 & n12512 ;
  assign n12514 = ( n12497 & ~n12509 ) | ( n12497 & n12513 ) | ( ~n12509 & n12513 ) ;
  assign n12515 = n12379 | n12514 ;
  assign n12516 = ~n12376 & n12515 ;
  assign n12517 = ( n10849 & n12179 ) | ( n10849 & n12209 ) | ( n12179 & n12209 ) ;
  assign n12518 = ( n10849 & n12178 ) | ( n10849 & n12208 ) | ( n12178 & n12208 ) ;
  assign n12519 = n12149 | n12518 ;
  assign n12520 = ~n12517 & n12519 ;
  assign n12521 = ~n12360 & n12520 ;
  assign n12522 = n12360 & ~n12520 ;
  assign n12523 = n12521 | n12522 ;
  assign n12524 = ~n12371 & n12375 ;
  assign n12525 = ( n12375 & n12520 ) | ( n12375 & n12524 ) | ( n12520 & n12524 ) ;
  assign n12526 = ~n12523 & n12525 ;
  assign n12527 = n12521 | n12526 ;
  assign n12528 = n12375 | n12520 ;
  assign n12529 = ~n12523 & n12528 ;
  assign n12530 = n12521 | n12529 ;
  assign n12531 = ( n12516 & n12527 ) | ( n12516 & n12530 ) | ( n12527 & n12530 ) ;
  assign n12532 = ~n12367 & n12531 ;
  assign n12533 = n12365 | n12532 ;
  assign n12534 = ( n10849 & n12185 ) | ( n10849 & n12215 ) | ( n12185 & n12215 ) ;
  assign n12535 = ( n10849 & n12184 ) | ( n10849 & n12214 ) | ( n12184 & n12214 ) ;
  assign n12536 = n11997 & ~n12535 ;
  assign n12537 = n12534 | n12536 ;
  assign n12538 = ~n12364 & n12537 ;
  assign n12539 = ~n12351 & n12537 ;
  assign n12540 = n12538 | n12539 ;
  assign n12541 = n12351 | n12355 ;
  assign n12542 = ~n12540 & n12541 ;
  assign n12543 = ~n12356 & n12542 ;
  assign n12544 = n12351 & ~n12537 ;
  assign n12545 = n12364 & ~n12537 ;
  assign n12546 = ~n12544 & n12545 ;
  assign n12547 = ( n12543 & n12544 ) | ( n12543 & n12546 ) | ( n12544 & n12546 ) ;
  assign n12548 = ( n12533 & n12543 ) | ( n12533 & n12547 ) | ( n12543 & n12547 ) ;
  assign n12549 = n12356 | n12548 ;
  assign n12550 = ( n10849 & n12193 ) | ( n10849 & n12223 ) | ( n12193 & n12223 ) ;
  assign n12551 = ( n10849 & n12192 ) | ( n10849 & n12222 ) | ( n12192 & n12222 ) ;
  assign n12552 = n11630 | n12551 ;
  assign n12553 = ~n12550 & n12552 ;
  assign n12554 = n12340 & n12553 ;
  assign n12555 = ( n10849 & n12191 ) | ( n10849 & n12221 ) | ( n12191 & n12221 ) ;
  assign n12556 = ( n10849 & n12190 ) | ( n10849 & n12220 ) | ( n12190 & n12220 ) ;
  assign n12557 = n11679 | n12556 ;
  assign n12558 = ~n12555 & n12557 ;
  assign n12559 = n12553 & n12558 ;
  assign n12560 = n12355 | n12558 ;
  assign n12561 = n12553 | n12558 ;
  assign n12562 = ~n12559 & n12561 ;
  assign n12563 = n12560 & n12562 ;
  assign n12564 = n12340 | n12553 ;
  assign n12565 = ( n12559 & n12563 ) | ( n12559 & n12564 ) | ( n12563 & n12564 ) ;
  assign n12566 = ~n12554 & n12565 ;
  assign n12567 = n12554 | n12566 ;
  assign n12568 = n12355 & n12558 ;
  assign n12569 = n12562 & n12568 ;
  assign n12570 = ( n12559 & n12566 ) | ( n12559 & n12569 ) | ( n12566 & n12569 ) ;
  assign n12571 = n12554 | n12570 ;
  assign n12572 = ( n12549 & n12567 ) | ( n12549 & n12571 ) | ( n12567 & n12571 ) ;
  assign n12573 = ~n12347 & n12572 ;
  assign n12574 = n12345 | n12573 ;
  assign n12575 = n12325 & n12335 ;
  assign n12576 = n12336 & ~n12575 ;
  assign n12577 = ( n10849 & n12203 ) | ( n10849 & n12231 ) | ( n12203 & n12231 ) ;
  assign n12578 = ( n10849 & n12202 ) | ( n10849 & n12230 ) | ( n12202 & n12230 ) ;
  assign n12579 = n11028 | n12578 ;
  assign n12580 = ~n12577 & n12579 ;
  assign n12581 = ~n12335 & n12580 ;
  assign n12582 = n12335 & ~n12580 ;
  assign n12583 = ( n10849 & n12201 ) | ( n10849 & n12229 ) | ( n12201 & n12229 ) ;
  assign n12584 = ( n10849 & n12200 ) | ( n10849 & n12228 ) | ( n12200 & n12228 ) ;
  assign n12585 = n11126 & ~n12584 ;
  assign n12586 = n12583 | n12585 ;
  assign n12587 = n12580 & ~n12586 ;
  assign n12588 = n12344 & n12586 ;
  assign n12589 = ~n12580 & n12586 ;
  assign n12590 = n12587 | n12589 ;
  assign n12591 = n12588 | n12590 ;
  assign n12592 = ~n12587 & n12591 ;
  assign n12593 = n12582 | n12592 ;
  assign n12594 = n12581 | n12593 ;
  assign n12595 = ~n12581 & n12594 ;
  assign n12596 = n12576 & ~n12595 ;
  assign n12597 = n12344 | n12586 ;
  assign n12598 = n12590 | n12597 ;
  assign n12599 = ( ~n12587 & n12594 ) | ( ~n12587 & n12598 ) | ( n12594 & n12598 ) ;
  assign n12600 = ~n12581 & n12599 ;
  assign n12601 = n12576 & ~n12600 ;
  assign n12602 = ( n12574 & n12596 ) | ( n12574 & n12601 ) | ( n12596 & n12601 ) ;
  assign n12603 = n12336 & ~n12602 ;
  assign n12604 = n12331 & ~n12603 ;
  assign n12605 = ( n12237 & n12303 ) | ( n12237 & ~n12307 ) | ( n12303 & ~n12307 ) ;
  assign n12606 = ~n12315 & n12605 ;
  assign n12607 = ~n12300 & n12316 ;
  assign n12608 = n12606 | n12607 ;
  assign n12609 = ~n12328 & n12608 ;
  assign n12610 = n12329 & ~n12609 ;
  assign n12611 = ~n12318 & n12608 ;
  assign n12612 = n12314 | n12611 ;
  assign n12613 = n12610 | n12612 ;
  assign n12614 = n12317 & ~n12613 ;
  assign n12615 = n12318 & ~n12614 ;
  assign n12616 = ~n12322 & n12615 ;
  assign n12617 = ( n12314 & ~n12604 ) | ( n12314 & n12616 ) | ( ~n12604 & n12616 ) ;
  assign n12618 = n12323 & ~n12617 ;
  assign n12619 = x14 & ~n12618 ;
  assign n12620 = ~x14 & n12618 ;
  assign n12621 = n12619 | n12620 ;
  assign n12622 = n1476 | n3315 ;
  assign n12623 = n2165 | n5595 ;
  assign n12624 = n12622 | n12623 ;
  assign n12625 = n1128 | n1194 ;
  assign n12626 = n513 | n12625 ;
  assign n12627 = n327 | n12626 ;
  assign n12628 = n12624 | n12627 ;
  assign n12629 = n276 | n449 ;
  assign n12630 = n76 | n12629 ;
  assign n12631 = n12628 | n12630 ;
  assign n12632 = n985 | n1889 ;
  assign n12633 = n822 | n12632 ;
  assign n12634 = n2284 | n12633 ;
  assign n12635 = n11332 | n12634 ;
  assign n12636 = n12631 | n12635 ;
  assign n12637 = n2283 | n12636 ;
  assign n12638 = n190 | n240 ;
  assign n12639 = n611 | n12638 ;
  assign n12640 = n378 | n861 ;
  assign n12641 = n12639 | n12640 ;
  assign n12642 = n263 | n315 ;
  assign n12643 = n390 | n12642 ;
  assign n12644 = n112 | n12643 ;
  assign n12645 = n12641 | n12644 ;
  assign n12646 = n661 | n12645 ;
  assign n12647 = n173 | n420 ;
  assign n12648 = n336 | n12647 ;
  assign n12649 = n2386 | n12648 ;
  assign n12650 = n512 | n3152 ;
  assign n12651 = n273 | n12650 ;
  assign n12652 = n12649 | n12651 ;
  assign n12653 = n262 | n435 ;
  assign n12654 = n62 | n12653 ;
  assign n12655 = n52 | n12654 ;
  assign n12656 = n83 | n12655 ;
  assign n12657 = n12652 | n12656 ;
  assign n12658 = n12646 | n12657 ;
  assign n12659 = n2527 | n12658 ;
  assign n12660 = n2333 | n12659 ;
  assign n12661 = n12637 | n12660 ;
  assign n12662 = n127 | n635 ;
  assign n12663 = n933 | n12662 ;
  assign n12664 = n531 | n12663 ;
  assign n12665 = n280 | n12664 ;
  assign n12666 = n139 | n12665 ;
  assign n12667 = n12661 | n12666 ;
  assign n12668 = n1574 | n1634 ;
  assign n12669 = n1886 & ~n12668 ;
  assign n12670 = n539 | n1022 ;
  assign n12671 = n596 | n12670 ;
  assign n12672 = n579 | n12671 ;
  assign n12673 = n12669 & ~n12672 ;
  assign n12674 = ~n77 & n12673 ;
  assign n12675 = n295 | n2267 ;
  assign n12676 = n1738 | n12675 ;
  assign n12677 = n1202 | n4068 ;
  assign n12678 = n12676 | n12677 ;
  assign n12679 = n1636 | n12678 ;
  assign n12680 = n12674 & ~n12679 ;
  assign n12681 = ~n10952 & n12680 ;
  assign n12682 = ~n3171 & n12681 ;
  assign n12683 = n315 | n592 ;
  assign n12684 = n431 | n435 ;
  assign n12685 = n12683 | n12684 ;
  assign n12686 = n309 | n655 ;
  assign n12687 = n92 | n12686 ;
  assign n12688 = n12685 | n12687 ;
  assign n12689 = n1079 | n12688 ;
  assign n12690 = n779 | n12689 ;
  assign n12691 = n490 | n12690 ;
  assign n12692 = n483 | n12691 ;
  assign n12693 = n416 | n12692 ;
  assign n12694 = n583 | n12693 ;
  assign n12695 = n12682 & ~n12694 ;
  assign n12696 = n403 | n441 ;
  assign n12697 = n12695 & ~n12696 ;
  assign n12698 = n12667 & ~n12697 ;
  assign n12699 = ~n12667 & n12697 ;
  assign n12700 = n12698 | n12699 ;
  assign n12701 = n5503 | n5508 ;
  assign n12702 = n5512 | n12701 ;
  assign n12703 = n5515 | n12702 ;
  assign n12704 = ~n12314 & n12703 ;
  assign n12705 = ~x8 & n12704 ;
  assign n12706 = x8 | n12705 ;
  assign n12707 = ( ~n12704 & n12705 ) | ( ~n12704 & n12706 ) | ( n12705 & n12706 ) ;
  assign n12708 = n12700 | n12707 ;
  assign n12709 = n1574 | n2635 ;
  assign n12710 = n1436 | n12709 ;
  assign n12711 = ( ~n63 & n530 ) | ( ~n63 & n2183 ) | ( n530 & n2183 ) ;
  assign n12712 = n274 | n12711 ;
  assign n12713 = n12710 | n12712 ;
  assign n12714 = n379 | n417 ;
  assign n12715 = n608 | n12714 ;
  assign n12716 = n226 & ~n12715 ;
  assign n12717 = ~n12713 & n12716 ;
  assign n12718 = ~n5230 & n12717 ;
  assign n12719 = n1918 | n3657 ;
  assign n12720 = n5593 | n12719 ;
  assign n12721 = n269 | n619 ;
  assign n12722 = n3707 | n12721 ;
  assign n12723 = n125 | n296 ;
  assign n12724 = n165 | n12723 ;
  assign n12725 = n12722 | n12724 ;
  assign n12726 = n820 | n12725 ;
  assign n12727 = ( ~n2753 & n12720 ) | ( ~n2753 & n12726 ) | ( n12720 & n12726 ) ;
  assign n12728 = n2753 | n12727 ;
  assign n12729 = n12718 & ~n12728 ;
  assign n12730 = n405 | n430 ;
  assign n12731 = n278 | n12730 ;
  assign n12732 = n335 | n12731 ;
  assign n12733 = n622 | n12732 ;
  assign n12734 = n3791 | n12733 ;
  assign n12735 = n445 | n12734 ;
  assign n12736 = n77 | n12735 ;
  assign n12737 = n94 | n12736 ;
  assign n12738 = n12729 & ~n12737 ;
  assign n12739 = ~n85 & n12738 ;
  assign n12740 = ( n12698 & ~n12708 ) | ( n12698 & n12739 ) | ( ~n12708 & n12739 ) ;
  assign n12741 = ( ~n12698 & n12699 ) | ( ~n12698 & n12707 ) | ( n12699 & n12707 ) ;
  assign n12742 = ~n12739 & n12741 ;
  assign n12743 = n12740 | n12742 ;
  assign n12744 = n3744 & ~n12502 ;
  assign n12745 = n3727 & n12387 ;
  assign n12746 = n3639 & n12383 ;
  assign n12747 = n12745 | n12746 ;
  assign n12748 = n12744 | n12747 ;
  assign n12749 = ~n12743 & n12748 ;
  assign n12750 = n12740 | n12749 ;
  assign n12751 = n3636 | n12748 ;
  assign n12752 = ~n12743 & n12751 ;
  assign n12753 = n12740 | n12752 ;
  assign n12754 = ( n12387 & n12497 ) | ( n12387 & ~n12502 ) | ( n12497 & ~n12502 ) ;
  assign n12755 = ( ~n12497 & n12502 ) | ( ~n12497 & n12754 ) | ( n12502 & n12754 ) ;
  assign n12756 = ( ~n12387 & n12754 ) | ( ~n12387 & n12755 ) | ( n12754 & n12755 ) ;
  assign n12757 = ( n12750 & n12753 ) | ( n12750 & ~n12756 ) | ( n12753 & ~n12756 ) ;
  assign n12758 = n749 | n1954 ;
  assign n12759 = n2545 | n12758 ;
  assign n12760 = n262 | n591 ;
  assign n12761 = n2163 | n12760 ;
  assign n12762 = n65 | n12761 ;
  assign n12763 = n693 | n12762 ;
  assign n12764 = n12759 | n12763 ;
  assign n12765 = n1842 & ~n12764 ;
  assign n12766 = n55 | n283 ;
  assign n12767 = n126 | n661 ;
  assign n12768 = n12766 | n12767 ;
  assign n12769 = ( n515 & ~n3978 ) | ( n515 & n12768 ) | ( ~n3978 & n12768 ) ;
  assign n12770 = n3978 | n12769 ;
  assign n12771 = n2341 | n12770 ;
  assign n12772 = n12765 & ~n12771 ;
  assign n12773 = n483 | n806 ;
  assign n12774 = n431 | n12773 ;
  assign n12775 = n619 | n12774 ;
  assign n12776 = n132 | n12775 ;
  assign n12777 = n139 | n12776 ;
  assign n12778 = n294 | n1189 ;
  assign n12779 = n1598 | n12778 ;
  assign n12780 = n688 | n12779 ;
  assign n12781 = n12777 | n12780 ;
  assign n12782 = n12772 & ~n12781 ;
  assign n12783 = n565 | n1985 ;
  assign n12784 = n59 | n472 ;
  assign n12785 = n12783 | n12784 ;
  assign n12786 = n242 | n245 ;
  assign n12787 = n321 | n12786 ;
  assign n12788 = n379 | n12787 ;
  assign n12789 = n12785 | n12788 ;
  assign n12790 = n344 | n390 ;
  assign n12791 = n12789 | n12790 ;
  assign n12792 = n4700 | n12791 ;
  assign n12793 = n1069 | n12792 ;
  assign n12794 = n12782 & ~n12793 ;
  assign n12795 = n281 | n568 ;
  assign n12796 = n635 | n12795 ;
  assign n12797 = n432 | n12796 ;
  assign n12798 = n637 | n12797 ;
  assign n12799 = n269 | n12798 ;
  assign n12800 = n346 | n12799 ;
  assign n12801 = n76 | n12800 ;
  assign n12802 = n151 | n12801 ;
  assign n12803 = n12794 & ~n12802 ;
  assign n12804 = ~n12739 & n12803 ;
  assign n12805 = n12739 & ~n12803 ;
  assign n12806 = n12750 & ~n12805 ;
  assign n12807 = n12753 & ~n12805 ;
  assign n12808 = ( ~n12756 & n12806 ) | ( ~n12756 & n12807 ) | ( n12806 & n12807 ) ;
  assign n12809 = ~n12804 & n12808 ;
  assign n12810 = n12757 & ~n12809 ;
  assign n12811 = ( n12757 & n12805 ) | ( n12757 & ~n12810 ) | ( n12805 & ~n12810 ) ;
  assign n12812 = n12804 | n12811 ;
  assign n12813 = ~n12810 & n12812 ;
  assign n12814 = ( n12497 & ~n12507 ) | ( n12497 & n12511 ) | ( ~n12507 & n12511 ) ;
  assign n12815 = n12505 & ~n12754 ;
  assign n12816 = n12814 | n12815 ;
  assign n12817 = n3744 & n12378 ;
  assign n12818 = n3639 & n12387 ;
  assign n12819 = n3727 & ~n12502 ;
  assign n12820 = n12818 | n12819 ;
  assign n12821 = n12817 | n12820 ;
  assign n12822 = n3636 | n12821 ;
  assign n12823 = ( ~n12816 & n12821 ) | ( ~n12816 & n12822 ) | ( n12821 & n12822 ) ;
  assign n12824 = ~n12813 & n12823 ;
  assign n12825 = n12813 & ~n12823 ;
  assign n12826 = n12824 | n12825 ;
  assign n12827 = n4048 & n12520 ;
  assign n12828 = n4043 & ~n12371 ;
  assign n12829 = n4045 & n12375 ;
  assign n12830 = n12828 | n12829 ;
  assign n12831 = n12827 | n12830 ;
  assign n12832 = n12375 & n12520 ;
  assign n12833 = n12528 & ~n12832 ;
  assign n12834 = n12516 | n12524 ;
  assign n12835 = ~n12833 & n12834 ;
  assign n12836 = ~n12525 & n12528 ;
  assign n12837 = ~n12516 & n12836 ;
  assign n12838 = n4051 & ~n12837 ;
  assign n12839 = ~n12835 & n12838 ;
  assign n12840 = ( n4051 & n12831 ) | ( n4051 & ~n12839 ) | ( n12831 & ~n12839 ) ;
  assign n12841 = ~x29 & n12840 ;
  assign n12842 = x29 | n12841 ;
  assign n12843 = ( ~n12840 & n12841 ) | ( ~n12840 & n12842 ) | ( n12841 & n12842 ) ;
  assign n12844 = ~n12826 & n12843 ;
  assign n12845 = n12824 | n12844 ;
  assign n12846 = ( n12497 & ~n12508 ) | ( n12497 & n12512 ) | ( ~n12508 & n12512 ) ;
  assign n12847 = n12499 & ~n12846 ;
  assign n12848 = n12514 | n12847 ;
  assign n12849 = n3744 & ~n12371 ;
  assign n12850 = n3639 & ~n12502 ;
  assign n12851 = n3727 & n12378 ;
  assign n12852 = n12850 | n12851 ;
  assign n12853 = n12849 | n12852 ;
  assign n12854 = n3636 | n12853 ;
  assign n12855 = ( ~n12848 & n12853 ) | ( ~n12848 & n12854 ) | ( n12853 & n12854 ) ;
  assign n12856 = n1245 | n2198 ;
  assign n12857 = n401 | n2588 ;
  assign n12858 = n12856 | n12857 ;
  assign n12859 = n4889 | n12858 ;
  assign n12860 = n3133 | n3230 ;
  assign n12861 = n12859 | n12860 ;
  assign n12862 = ~n841 & n3573 ;
  assign n12863 = ~n12861 & n12862 ;
  assign n12864 = n381 | n2179 ;
  assign n12865 = n1353 | n12864 ;
  assign n12866 = n139 | n457 ;
  assign n12867 = n12865 | n12866 ;
  assign n12868 = n1280 | n12867 ;
  assign n12869 = n3792 | n12868 ;
  assign n12870 = n521 | n12869 ;
  assign n12871 = n301 | n12870 ;
  assign n12872 = n416 | n12871 ;
  assign n12873 = n12863 & ~n12872 ;
  assign n12874 = ~n198 & n12873 ;
  assign n12875 = n12739 | n12874 ;
  assign n12876 = n12739 & n12874 ;
  assign n12877 = n12875 & ~n12876 ;
  assign n12878 = n7302 | n7305 ;
  assign n12879 = n7300 | n12878 ;
  assign n12880 = n7308 | n12879 ;
  assign n12881 = ~n12314 & n12880 ;
  assign n12882 = ~x11 & n12881 ;
  assign n12883 = x11 | n12882 ;
  assign n12884 = ( ~n12881 & n12882 ) | ( ~n12881 & n12883 ) | ( n12882 & n12883 ) ;
  assign n12885 = n12877 & ~n12884 ;
  assign n12886 = ~n12877 & n12884 ;
  assign n12887 = n12885 | n12886 ;
  assign n12888 = n12855 & ~n12887 ;
  assign n12889 = n12855 & ~n12888 ;
  assign n12890 = n12855 | n12887 ;
  assign n12891 = ~n12889 & n12890 ;
  assign n12892 = n12811 & ~n12891 ;
  assign n12893 = ~n12811 & n12891 ;
  assign n12894 = n12892 | n12893 ;
  assign n12895 = n12845 & ~n12894 ;
  assign n12896 = n12845 & ~n12895 ;
  assign n12897 = n12845 | n12894 ;
  assign n12898 = ~n12896 & n12897 ;
  assign n12899 = ( n12516 & n12526 ) | ( n12516 & n12529 ) | ( n12526 & n12529 ) ;
  assign n12900 = ( n12516 & n12525 ) | ( n12516 & n12528 ) | ( n12525 & n12528 ) ;
  assign n12901 = n12523 & ~n12900 ;
  assign n12902 = n12899 | n12901 ;
  assign n12903 = n4048 & ~n12360 ;
  assign n12904 = n4043 & n12375 ;
  assign n12905 = n4045 & n12520 ;
  assign n12906 = n12904 | n12905 ;
  assign n12907 = n12903 | n12906 ;
  assign n12908 = n4051 | n12907 ;
  assign n12909 = ( ~n12902 & n12907 ) | ( ~n12902 & n12908 ) | ( n12907 & n12908 ) ;
  assign n12910 = ~x29 & n12909 ;
  assign n12911 = x29 | n12910 ;
  assign n12912 = ( ~n12909 & n12910 ) | ( ~n12909 & n12911 ) | ( n12910 & n12911 ) ;
  assign n12913 = ~n12898 & n12912 ;
  assign n12914 = n12898 & ~n12912 ;
  assign n12915 = n12913 | n12914 ;
  assign n12916 = n4484 & n12351 ;
  assign n12917 = n4479 & n12364 ;
  assign n12918 = n4481 & ~n12537 ;
  assign n12919 = n12917 | n12918 ;
  assign n12920 = n12916 | n12919 ;
  assign n12921 = n12538 | n12545 ;
  assign n12922 = n12533 & ~n12921 ;
  assign n12923 = n12540 | n12544 ;
  assign n12924 = ( n12533 & n12546 ) | ( n12533 & ~n12923 ) | ( n12546 & ~n12923 ) ;
  assign n12925 = ( n12545 & n12922 ) | ( n12545 & ~n12924 ) | ( n12922 & ~n12924 ) ;
  assign n12926 = n12544 | n12546 ;
  assign n12927 = ( n12533 & ~n12540 ) | ( n12533 & n12926 ) | ( ~n12540 & n12926 ) ;
  assign n12928 = n12539 | n12927 ;
  assign n12929 = n4487 & ~n12928 ;
  assign n12930 = ( n4487 & n12925 ) | ( n4487 & n12929 ) | ( n12925 & n12929 ) ;
  assign n12931 = n12920 | n12930 ;
  assign n12932 = x26 | n12931 ;
  assign n12933 = ~x26 & n12932 ;
  assign n12934 = ( ~n12931 & n12932 ) | ( ~n12931 & n12933 ) | ( n12932 & n12933 ) ;
  assign n12935 = ~n12915 & n12934 ;
  assign n12936 = n12915 | n12935 ;
  assign n12937 = n12915 & n12934 ;
  assign n12938 = ( n12749 & n12752 ) | ( n12749 & ~n12756 ) | ( n12752 & ~n12756 ) ;
  assign n12939 = ( n12748 & n12751 ) | ( n12748 & ~n12756 ) | ( n12751 & ~n12756 ) ;
  assign n12940 = n12743 & ~n12939 ;
  assign n12941 = n12938 | n12940 ;
  assign n12942 = n12700 & n12707 ;
  assign n12943 = n12708 & ~n12942 ;
  assign n12944 = n12397 | n12404 ;
  assign n12945 = ( n12393 & n12495 ) | ( n12393 & n12944 ) | ( n12495 & n12944 ) ;
  assign n12946 = ~n12496 & n12945 ;
  assign n12947 = n12394 & ~n12497 ;
  assign n12948 = n12946 | n12947 ;
  assign n12949 = n3744 & n12387 ;
  assign n12950 = n3639 & n12392 ;
  assign n12951 = n3727 & n12383 ;
  assign n12952 = n12950 | n12951 ;
  assign n12953 = n12949 | n12952 ;
  assign n12954 = n3636 | n12953 ;
  assign n12955 = ( n12948 & n12953 ) | ( n12948 & n12954 ) | ( n12953 & n12954 ) ;
  assign n12956 = n3146 | n4309 ;
  assign n12957 = n145 | n245 ;
  assign n12958 = n1352 | n12957 ;
  assign n12959 = n2037 | n12958 ;
  assign n12960 = n12956 | n12959 ;
  assign n12961 = n1861 | n12960 ;
  assign n12962 = n724 | n12961 ;
  assign n12963 = n433 | n12962 ;
  assign n12964 = n1858 & ~n12963 ;
  assign n12965 = n446 | n686 ;
  assign n12966 = n166 | n12965 ;
  assign n12967 = n12964 & ~n12966 ;
  assign n12968 = n2816 | n2822 ;
  assign n12969 = n490 | n12968 ;
  assign n12970 = n12967 & ~n12969 ;
  assign n12971 = n622 | n655 ;
  assign n12972 = n653 | n12971 ;
  assign n12973 = n76 | n12972 ;
  assign n12974 = n92 | n12973 ;
  assign n12975 = n12970 & ~n12974 ;
  assign n12976 = n12667 | n12975 ;
  assign n12977 = n9780 | n9781 ;
  assign n12978 = ~n12314 & n12977 ;
  assign n12979 = ~x2 & n12978 ;
  assign n12980 = x2 | n12979 ;
  assign n12981 = ( ~n12978 & n12979 ) | ( ~n12978 & n12980 ) | ( n12979 & n12980 ) ;
  assign n12982 = n8681 | n9245 ;
  assign n12983 = n8680 | n12982 ;
  assign n12984 = n8685 | n12983 ;
  assign n12985 = ~n12314 & n12984 ;
  assign n12986 = ~x5 & n12985 ;
  assign n12987 = x5 & ~n12985 ;
  assign n12988 = n12986 | n12987 ;
  assign n12989 = n476 | n869 ;
  assign n12990 = n12768 | n12989 ;
  assign n12991 = n432 | n12990 ;
  assign n12992 = n888 | n1057 ;
  assign n12993 = n4843 | n12992 ;
  assign n12994 = n2119 | n3232 ;
  assign n12995 = n12993 | n12994 ;
  assign n12996 = n12991 | n12995 ;
  assign n12997 = n2488 | n11060 ;
  assign n12998 = n12996 | n12997 ;
  assign n12999 = n367 | n1578 ;
  assign n13000 = n12998 | n12999 ;
  assign n13001 = n1680 | n4225 ;
  assign n13002 = n3152 | n13001 ;
  assign n13003 = n746 | n13002 ;
  assign n13004 = n990 | n2960 ;
  assign n13005 = n521 | n13004 ;
  assign n13006 = n321 | n13005 ;
  assign n13007 = n13003 | n13006 ;
  assign n13008 = n204 | n403 ;
  assign n13009 = n112 | n13008 ;
  assign n13010 = n152 | n13009 ;
  assign n13011 = n157 | n13010 ;
  assign n13012 = n13007 | n13011 ;
  assign n13013 = n278 | n13012 ;
  assign n13014 = n13000 | n13013 ;
  assign n13015 = n1129 | n4841 ;
  assign n13016 = n5240 | n13015 ;
  assign n13017 = n5756 | n13016 ;
  assign n13018 = n12717 & ~n13017 ;
  assign n13019 = ~n11197 & n13018 ;
  assign n13020 = ~n252 & n13019 ;
  assign n13021 = ~n13014 & n13020 ;
  assign n13022 = n2950 | n3217 ;
  assign n13023 = n3850 | n13022 ;
  assign n13024 = n637 | n13023 ;
  assign n13025 = n282 | n13024 ;
  assign n13026 = n240 | n13025 ;
  assign n13027 = n99 | n13026 ;
  assign n13028 = n13021 & ~n13027 ;
  assign n13029 = ( n12981 & n12988 ) | ( n12981 & n13028 ) | ( n12988 & n13028 ) ;
  assign n13030 = n12667 | n13029 ;
  assign n13031 = n12667 & n13029 ;
  assign n13032 = n13030 & ~n13031 ;
  assign n13033 = n12407 | n12494 ;
  assign n13034 = ~n12495 & n13033 ;
  assign n13035 = n3744 & n12392 ;
  assign n13036 = n3727 & n12401 ;
  assign n13037 = n3639 & n12415 ;
  assign n13038 = n13036 | n13037 ;
  assign n13039 = n13035 | n13038 ;
  assign n13040 = n3636 | n13039 ;
  assign n13041 = ( n13034 & n13039 ) | ( n13034 & n13040 ) | ( n13039 & n13040 ) ;
  assign n13042 = n13032 & n13041 ;
  assign n13043 = n13030 & ~n13042 ;
  assign n13044 = n12667 & n12975 ;
  assign n13045 = n12976 & ~n13044 ;
  assign n13046 = ~n13043 & n13045 ;
  assign n13047 = ( n12943 & ~n12976 ) | ( n12943 & n13046 ) | ( ~n12976 & n13046 ) ;
  assign n13048 = ( n12976 & n13043 ) | ( n12976 & n13044 ) | ( n13043 & n13044 ) ;
  assign n13049 = ~n12943 & n13048 ;
  assign n13050 = n13047 | n13049 ;
  assign n13051 = n12955 & n13050 ;
  assign n13052 = n12955 | n13050 ;
  assign n13053 = ~n13051 & n13052 ;
  assign n13054 = ( n12943 & n12955 ) | ( n12943 & n13053 ) | ( n12955 & n13053 ) ;
  assign n13055 = ~n12941 & n13054 ;
  assign n13056 = n12941 & ~n13054 ;
  assign n13057 = n13055 | n13056 ;
  assign n13058 = n4048 & n12375 ;
  assign n13059 = n4043 & n12378 ;
  assign n13060 = n4045 & ~n12371 ;
  assign n13061 = n13059 | n13060 ;
  assign n13062 = n13058 | n13061 ;
  assign n13063 = n12376 | n12524 ;
  assign n13064 = n12515 & n13063 ;
  assign n13065 = n12516 | n13063 ;
  assign n13066 = n4051 & n13065 ;
  assign n13067 = ~n13064 & n13066 ;
  assign n13068 = ( n4051 & n13062 ) | ( n4051 & ~n13067 ) | ( n13062 & ~n13067 ) ;
  assign n13069 = x29 & n13068 ;
  assign n13070 = x29 & ~n13069 ;
  assign n13071 = ( n13068 & ~n13069 ) | ( n13068 & n13070 ) | ( ~n13069 & n13070 ) ;
  assign n13072 = ~n13057 & n13071 ;
  assign n13073 = n13055 | n13072 ;
  assign n13074 = n12826 & ~n12843 ;
  assign n13075 = n12844 | n13074 ;
  assign n13076 = n4484 & ~n12537 ;
  assign n13077 = n4479 & ~n12360 ;
  assign n13078 = n4481 & n12364 ;
  assign n13079 = n13077 | n13078 ;
  assign n13080 = n13076 | n13079 ;
  assign n13081 = n12533 & ~n12922 ;
  assign n13082 = n12533 | n12921 ;
  assign n13083 = ( n4487 & n13081 ) | ( n4487 & ~n13082 ) | ( n13081 & ~n13082 ) ;
  assign n13084 = n13080 | n13083 ;
  assign n13085 = x26 | n13084 ;
  assign n13086 = ~x26 & n13085 ;
  assign n13087 = ( ~n13084 & n13085 ) | ( ~n13084 & n13086 ) | ( n13085 & n13086 ) ;
  assign n13088 = ( ~n13073 & n13075 ) | ( ~n13073 & n13087 ) | ( n13075 & n13087 ) ;
  assign n13089 = ( n13073 & ~n13075 ) | ( n13073 & n13088 ) | ( ~n13075 & n13088 ) ;
  assign n13090 = n12937 | n13089 ;
  assign n13091 = n12936 & ~n13090 ;
  assign n13092 = ( ~n12936 & n12937 ) | ( ~n12936 & n13089 ) | ( n12937 & n13089 ) ;
  assign n13093 = n13091 | n13092 ;
  assign n13094 = ( n12549 & n12563 ) | ( n12549 & n12569 ) | ( n12563 & n12569 ) ;
  assign n13095 = ( n12355 & n12549 ) | ( n12355 & n12558 ) | ( n12549 & n12558 ) ;
  assign n13096 = n12562 | n13095 ;
  assign n13097 = ~n13094 & n13096 ;
  assign n13098 = n4551 & n12553 ;
  assign n13099 = n4546 & n12355 ;
  assign n13100 = n4548 & n12558 ;
  assign n13101 = n13099 | n13100 ;
  assign n13102 = n13098 | n13101 ;
  assign n13103 = n4554 | n13102 ;
  assign n13104 = ( n13097 & n13102 ) | ( n13097 & n13103 ) | ( n13102 & n13103 ) ;
  assign n13105 = x23 & n13104 ;
  assign n13106 = x23 & ~n13105 ;
  assign n13107 = ( n13104 & ~n13105 ) | ( n13104 & n13106 ) | ( ~n13105 & n13106 ) ;
  assign n13108 = ~n13093 & n13107 ;
  assign n13109 = n13093 | n13108 ;
  assign n13110 = n13093 & n13107 ;
  assign n13111 = ( ~n13087 & n13088 ) | ( ~n13087 & n13089 ) | ( n13088 & n13089 ) ;
  assign n13112 = n12367 & ~n12531 ;
  assign n13113 = n12532 | n13112 ;
  assign n13114 = n4484 & n12364 ;
  assign n13115 = n4479 & n12520 ;
  assign n13116 = n4481 & ~n12360 ;
  assign n13117 = n13115 | n13116 ;
  assign n13118 = n13114 | n13117 ;
  assign n13119 = n4487 | n13118 ;
  assign n13120 = ( ~n13113 & n13118 ) | ( ~n13113 & n13119 ) | ( n13118 & n13119 ) ;
  assign n13121 = ~x26 & n13120 ;
  assign n13122 = x26 | n13121 ;
  assign n13123 = ( ~n13120 & n13121 ) | ( ~n13120 & n13122 ) | ( n13121 & n13122 ) ;
  assign n13124 = n4048 & ~n12371 ;
  assign n13125 = n4043 & ~n12502 ;
  assign n13126 = n4045 & n12378 ;
  assign n13127 = n13125 | n13126 ;
  assign n13128 = n13124 | n13127 ;
  assign n13129 = n4051 | n13128 ;
  assign n13130 = ( ~n12848 & n13128 ) | ( ~n12848 & n13129 ) | ( n13128 & n13129 ) ;
  assign n13131 = ~x29 & n13130 ;
  assign n13132 = x29 | n13131 ;
  assign n13133 = ( ~n13130 & n13131 ) | ( ~n13130 & n13132 ) | ( n13131 & n13132 ) ;
  assign n13134 = ~n13053 & n13133 ;
  assign n13135 = n13043 | n13046 ;
  assign n13136 = n13043 & n13045 ;
  assign n13137 = n13135 & ~n13136 ;
  assign n13138 = ( n12403 & n12404 ) | ( n12403 & n12495 ) | ( n12404 & n12495 ) ;
  assign n13139 = n12402 | n12403 ;
  assign n13140 = n12495 | n13139 ;
  assign n13141 = ~n13138 & n13140 ;
  assign n13142 = n3744 & n12383 ;
  assign n13143 = n3639 & n12401 ;
  assign n13144 = n3727 & n12392 ;
  assign n13145 = n13143 | n13144 ;
  assign n13146 = n13142 | n13145 ;
  assign n13147 = n3636 | n13146 ;
  assign n13148 = ( n13141 & n13146 ) | ( n13141 & n13147 ) | ( n13146 & n13147 ) ;
  assign n13149 = ~n13137 & n13148 ;
  assign n13150 = n13137 & ~n13148 ;
  assign n13151 = n13149 | n13150 ;
  assign n13152 = n13032 | n13041 ;
  assign n13153 = ~n13042 & n13152 ;
  assign n13154 = n3744 & n12401 ;
  assign n13155 = n3639 & n12411 ;
  assign n13156 = n3727 & n12415 ;
  assign n13157 = n13155 | n13156 ;
  assign n13158 = n13154 | n13157 ;
  assign n13159 = n12489 | n12490 ;
  assign n13160 = ~n12491 & n12493 ;
  assign n13161 = n13159 & ~n13160 ;
  assign n13162 = ~n12492 & n12493 ;
  assign n13163 = ~n12489 & n13162 ;
  assign n13164 = n3636 & n13163 ;
  assign n13165 = ( n3636 & n13161 ) | ( n3636 & n13164 ) | ( n13161 & n13164 ) ;
  assign n13166 = n13158 | n13165 ;
  assign n13170 = n531 | n2216 ;
  assign n13171 = n1330 | n13170 ;
  assign n13172 = n1737 | n13171 ;
  assign n13173 = n3438 | n13172 ;
  assign n13174 = n11164 | n13173 ;
  assign n13175 = n4923 | n13174 ;
  assign n13176 = n11148 | n13175 ;
  assign n13177 = n933 | n2709 ;
  assign n13178 = n478 | n13177 ;
  assign n13179 = n283 | n13178 ;
  assign n13180 = n274 | n13179 ;
  assign n13181 = n203 | n13180 ;
  assign n13182 = n226 & ~n13181 ;
  assign n13183 = ~n13176 & n13182 ;
  assign n13184 = n160 | n457 ;
  assign n13185 = n173 | n13184 ;
  assign n13186 = n168 | n13185 ;
  assign n13187 = n81 | n13186 ;
  assign n13188 = n13183 & ~n13187 ;
  assign n13189 = n408 | n452 ;
  assign n13190 = n996 | n13189 ;
  assign n13191 = n669 | n13190 ;
  assign n13192 = n12240 | n13191 ;
  assign n13193 = n1657 | n13192 ;
  assign n13194 = n252 | n13193 ;
  assign n13195 = n3321 | n13194 ;
  assign n13196 = n1811 | n13195 ;
  assign n13197 = n13014 | n13196 ;
  assign n13198 = n1337 | n1866 ;
  assign n13199 = n1443 | n13198 ;
  assign n13200 = n1125 | n13199 ;
  assign n13201 = n339 | n13200 ;
  assign n13202 = n93 | n13201 ;
  assign n13203 = n3856 | n13202 ;
  assign n13204 = n13197 | n13203 ;
  assign n13205 = n310 | n528 ;
  assign n13206 = n607 | n13205 ;
  assign n13207 = n222 | n13206 ;
  assign n13208 = n142 | n13207 ;
  assign n13209 = n145 | n13208 ;
  assign n13210 = n217 | n13209 ;
  assign n13211 = n13204 | n13210 ;
  assign n13212 = n12981 | n13211 ;
  assign n13213 = n1463 | n2146 ;
  assign n13214 = n2434 | n13213 ;
  assign n13215 = n3655 | n11202 ;
  assign n13216 = n13214 | n13215 ;
  assign n13217 = n1679 | n13216 ;
  assign n13218 = n1837 | n2178 ;
  assign n13219 = n335 | n619 ;
  assign n13220 = n327 | n13219 ;
  assign n13221 = n13218 | n13220 ;
  assign n13222 = n187 | n364 ;
  assign n13223 = n13221 | n13222 ;
  assign n13224 = n2219 | n13223 ;
  assign n13225 = n13217 | n13224 ;
  assign n13226 = n597 | n5821 ;
  assign n13227 = n437 | n13226 ;
  assign n13228 = n111 | n13227 ;
  assign n13229 = n1636 | n13228 ;
  assign n13230 = n633 | n13229 ;
  assign n13231 = n13225 | n13230 ;
  assign n13232 = n521 | n670 ;
  assign n13233 = n160 | n13232 ;
  assign n13234 = n99 | n13233 ;
  assign n13235 = n13231 | n13234 ;
  assign n13236 = n206 | n484 ;
  assign n13237 = n3558 | n13236 ;
  assign n13238 = n528 | n618 ;
  assign n13239 = n625 | n13238 ;
  assign n13240 = n13237 | n13239 ;
  assign n13241 = n277 | n595 ;
  assign n13242 = n434 | n13241 ;
  assign n13243 = n13240 | n13242 ;
  assign n13244 = ~n1288 & n2685 ;
  assign n13245 = ~n2953 & n13244 ;
  assign n13246 = ~n1712 & n13245 ;
  assign n13247 = ~n13243 & n13246 ;
  assign n13248 = n241 | n299 ;
  assign n13249 = n444 | n13248 ;
  assign n13250 = n450 | n13249 ;
  assign n13251 = n120 | n13250 ;
  assign n13252 = n181 | n13251 ;
  assign n13253 = n381 | n468 ;
  assign n13254 = n873 | n3532 ;
  assign n13255 = n2643 | n13254 ;
  assign n13256 = n1066 | n13255 ;
  assign n13257 = n1830 | n13256 ;
  assign n13258 = n641 | n2154 ;
  assign n13259 = n1656 | n13258 ;
  assign n13260 = ( ~n13253 & n13257 ) | ( ~n13253 & n13259 ) | ( n13257 & n13259 ) ;
  assign n13261 = n13253 | n13260 ;
  assign n13262 = n13252 | n13261 ;
  assign n13263 = n13247 & ~n13262 ;
  assign n13264 = ~n12768 & n13263 ;
  assign n13265 = ~n13235 & n13264 ;
  assign n13266 = n529 | n1522 ;
  assign n13267 = n498 | n13266 ;
  assign n13268 = n263 | n13267 ;
  assign n13269 = n240 | n13268 ;
  assign n13270 = n260 | n13269 ;
  assign n13271 = n596 | n13270 ;
  assign n13272 = n173 | n13271 ;
  assign n13273 = n13265 & ~n13272 ;
  assign n13274 = n3744 & n12419 ;
  assign n13275 = n3639 & n12433 ;
  assign n13276 = n3727 & ~n12423 ;
  assign n13277 = n13275 | n13276 ;
  assign n13278 = n13274 | n13277 ;
  assign n13279 = n3636 | n13278 ;
  assign n13280 = ( n12434 & n12483 ) | ( n12434 & ~n12484 ) | ( n12483 & ~n12484 ) ;
  assign n13281 = n12429 & ~n13280 ;
  assign n13282 = n12487 | n13281 ;
  assign n13283 = ( n13278 & n13279 ) | ( n13278 & ~n13282 ) | ( n13279 & ~n13282 ) ;
  assign n13284 = ( n12981 & ~n13273 ) | ( n12981 & n13283 ) | ( ~n13273 & n13283 ) ;
  assign n13285 = n13212 & n13284 ;
  assign n13286 = n12981 & n13211 ;
  assign n13287 = n13285 | n13286 ;
  assign n13288 = ( n12981 & ~n13188 ) | ( n12981 & n13287 ) | ( ~n13188 & n13287 ) ;
  assign n13167 = ( n12981 & ~n12988 ) | ( n12981 & n13028 ) | ( ~n12988 & n13028 ) ;
  assign n13168 = ( ~n12981 & n12988 ) | ( ~n12981 & n13167 ) | ( n12988 & n13167 ) ;
  assign n13169 = ( ~n13028 & n13167 ) | ( ~n13028 & n13168 ) | ( n13167 & n13168 ) ;
  assign n13289 = ( n13166 & n13169 ) | ( n13166 & ~n13288 ) | ( n13169 & ~n13288 ) ;
  assign n13290 = ( ~n13166 & n13288 ) | ( ~n13166 & n13289 ) | ( n13288 & n13289 ) ;
  assign n13291 = ( ~n13169 & n13289 ) | ( ~n13169 & n13290 ) | ( n13289 & n13290 ) ;
  assign n13292 = ( n13166 & n13288 ) | ( n13166 & n13291 ) | ( n13288 & n13291 ) ;
  assign n13293 = n13153 & n13292 ;
  assign n13294 = n13153 | n13292 ;
  assign n13295 = ~n13293 & n13294 ;
  assign n13296 = n4048 & ~n12502 ;
  assign n13297 = n4043 & n12383 ;
  assign n13298 = n4045 & n12387 ;
  assign n13299 = n13297 | n13298 ;
  assign n13300 = n13296 | n13299 ;
  assign n13301 = n4051 | n13300 ;
  assign n13302 = ( ~n12756 & n13300 ) | ( ~n12756 & n13301 ) | ( n13300 & n13301 ) ;
  assign n13303 = ~x29 & n13302 ;
  assign n13304 = x29 | n13303 ;
  assign n13305 = ( ~n13302 & n13303 ) | ( ~n13302 & n13304 ) | ( n13303 & n13304 ) ;
  assign n13306 = n13295 & n13305 ;
  assign n13307 = n13293 | n13306 ;
  assign n13308 = ~n13151 & n13307 ;
  assign n13309 = n13149 | n13308 ;
  assign n13310 = n13053 & ~n13133 ;
  assign n13311 = n13134 | n13310 ;
  assign n13312 = n13309 & ~n13311 ;
  assign n13313 = n13057 & ~n13071 ;
  assign n13314 = n13072 | n13313 ;
  assign n13315 = ( n13134 & n13312 ) | ( n13134 & ~n13314 ) | ( n13312 & ~n13314 ) ;
  assign n13316 = ~n13134 & n13314 ;
  assign n13317 = ~n13312 & n13316 ;
  assign n13318 = n13315 | n13317 ;
  assign n13319 = n13123 | n13318 ;
  assign n13320 = ~n13123 & n13319 ;
  assign n13321 = ( ~n13318 & n13319 ) | ( ~n13318 & n13320 ) | ( n13319 & n13320 ) ;
  assign n13322 = ( n13123 & n13315 ) | ( n13123 & n13321 ) | ( n13315 & n13321 ) ;
  assign n13323 = n4551 & n12558 ;
  assign n13324 = n4546 & n12351 ;
  assign n13325 = n4548 & n12355 ;
  assign n13326 = n13324 | n13325 ;
  assign n13327 = n13323 | n13326 ;
  assign n13328 = n4554 | n13327 ;
  assign n13329 = ( n12355 & n12558 ) | ( n12355 & ~n13095 ) | ( n12558 & ~n13095 ) ;
  assign n13330 = ( n12549 & ~n13095 ) | ( n12549 & n13329 ) | ( ~n13095 & n13329 ) ;
  assign n13331 = ( n13327 & n13328 ) | ( n13327 & n13330 ) | ( n13328 & n13330 ) ;
  assign n13332 = x23 & n13331 ;
  assign n13333 = x23 & ~n13332 ;
  assign n13334 = ( n13331 & ~n13332 ) | ( n13331 & n13333 ) | ( ~n13332 & n13333 ) ;
  assign n13335 = ( n13111 & ~n13322 ) | ( n13111 & n13334 ) | ( ~n13322 & n13334 ) ;
  assign n13336 = ( ~n13111 & n13322 ) | ( ~n13111 & n13335 ) | ( n13322 & n13335 ) ;
  assign n13337 = ( ~n13109 & n13110 ) | ( ~n13109 & n13336 ) | ( n13110 & n13336 ) ;
  assign n13338 = n13108 | n13337 ;
  assign n13339 = n4551 & n12340 ;
  assign n13340 = n4546 & n12558 ;
  assign n13341 = n4548 & n12553 ;
  assign n13342 = n13340 | n13341 ;
  assign n13343 = n13339 | n13342 ;
  assign n13344 = ( n12549 & n12566 ) | ( n12549 & n12570 ) | ( n12566 & n12570 ) ;
  assign n13345 = n12559 | n13094 ;
  assign n13346 = ~n13344 & n13345 ;
  assign n13347 = n12564 & ~n12572 ;
  assign n13348 = n4554 & n13347 ;
  assign n13349 = ( n4554 & n13346 ) | ( n4554 & n13348 ) | ( n13346 & n13348 ) ;
  assign n13350 = n13343 | n13349 ;
  assign n13351 = x23 | n13350 ;
  assign n13352 = ~x23 & n13351 ;
  assign n13353 = ( ~n13350 & n13351 ) | ( ~n13350 & n13352 ) | ( n13351 & n13352 ) ;
  assign n13354 = n12935 | n13092 ;
  assign n13355 = n12888 | n12892 ;
  assign n13356 = n479 | n4142 ;
  assign n13357 = n293 | n13356 ;
  assign n13358 = n4394 | n13357 ;
  assign n13359 = n4138 | n13358 ;
  assign n13360 = n2622 | n3371 ;
  assign n13361 = n867 | n13360 ;
  assign n13362 = n13359 | n13361 ;
  assign n13363 = n3158 | n3864 ;
  assign n13364 = n237 | n13363 ;
  assign n13365 = n499 | n13364 ;
  assign n13366 = n307 | n13365 ;
  assign n13367 = n1244 | n13366 ;
  assign n13368 = n13362 | n13367 ;
  assign n13369 = n52 | n167 ;
  assign n13370 = n139 | n13369 ;
  assign n13371 = n13368 | n13370 ;
  assign n13372 = ( n12875 & ~n12885 ) | ( n12875 & n13371 ) | ( ~n12885 & n13371 ) ;
  assign n13373 = ( n12875 & n12876 ) | ( n12875 & n12884 ) | ( n12876 & n12884 ) ;
  assign n13374 = n13371 & n13373 ;
  assign n13375 = n13372 & ~n13374 ;
  assign n13376 = n3744 & n12375 ;
  assign n13377 = n3727 & ~n12371 ;
  assign n13378 = n3639 & n12378 ;
  assign n13379 = n13377 | n13378 ;
  assign n13380 = n13376 | n13379 ;
  assign n13381 = n13375 & n13380 ;
  assign n13382 = ( n3636 & n13064 ) | ( n3636 & ~n13065 ) | ( n13064 & ~n13065 ) ;
  assign n13383 = ( n13375 & n13381 ) | ( n13375 & n13382 ) | ( n13381 & n13382 ) ;
  assign n13384 = n13375 | n13380 ;
  assign n13385 = n13382 | n13384 ;
  assign n13386 = ~n13383 & n13385 ;
  assign n13387 = n13355 & n13386 ;
  assign n13388 = n13355 | n13386 ;
  assign n13389 = ~n13387 & n13388 ;
  assign n13390 = n4048 & n12364 ;
  assign n13391 = n4043 & n12520 ;
  assign n13392 = n4045 & ~n12360 ;
  assign n13393 = n13391 | n13392 ;
  assign n13394 = n13390 | n13393 ;
  assign n13395 = n4051 | n13394 ;
  assign n13396 = ( ~n13113 & n13394 ) | ( ~n13113 & n13395 ) | ( n13394 & n13395 ) ;
  assign n13397 = ~x29 & n13396 ;
  assign n13398 = x29 | n13397 ;
  assign n13399 = ( ~n13396 & n13397 ) | ( ~n13396 & n13398 ) | ( n13397 & n13398 ) ;
  assign n13400 = n13389 & n13399 ;
  assign n13401 = n13389 | n13399 ;
  assign n13402 = ~n13400 & n13401 ;
  assign n13403 = n12895 | n13402 ;
  assign n13404 = n12913 | n13403 ;
  assign n13405 = ( n12895 & n12913 ) | ( n12895 & n13402 ) | ( n12913 & n13402 ) ;
  assign n13406 = n13404 & ~n13405 ;
  assign n13407 = ~n12548 & n12927 ;
  assign n13408 = n12541 & ~n12549 ;
  assign n13409 = n13407 | n13408 ;
  assign n13410 = n4484 & n12355 ;
  assign n13411 = n4479 & ~n12537 ;
  assign n13412 = n4481 & n12351 ;
  assign n13413 = n13411 | n13412 ;
  assign n13414 = n13410 | n13413 ;
  assign n13415 = n4487 | n13414 ;
  assign n13416 = ( n13409 & n13414 ) | ( n13409 & n13415 ) | ( n13414 & n13415 ) ;
  assign n13417 = x26 & n13416 ;
  assign n13418 = x26 & ~n13417 ;
  assign n13419 = ( n13416 & ~n13417 ) | ( n13416 & n13418 ) | ( ~n13417 & n13418 ) ;
  assign n13420 = n13406 & ~n13419 ;
  assign n13421 = n13419 | n13420 ;
  assign n13422 = ( ~n13406 & n13420 ) | ( ~n13406 & n13421 ) | ( n13420 & n13421 ) ;
  assign n13423 = ( n13353 & n13354 ) | ( n13353 & ~n13422 ) | ( n13354 & ~n13422 ) ;
  assign n13424 = ( ~n13354 & n13422 ) | ( ~n13354 & n13423 ) | ( n13422 & n13423 ) ;
  assign n13425 = ( ~n13353 & n13423 ) | ( ~n13353 & n13424 ) | ( n13423 & n13424 ) ;
  assign n13426 = n13338 & n13425 ;
  assign n13427 = n13338 | n13425 ;
  assign n13428 = ~n13426 & n13427 ;
  assign n13429 = ( ~n12574 & n12591 ) | ( ~n12574 & n12598 ) | ( n12591 & n12598 ) ;
  assign n13430 = ( ~n12574 & n12588 ) | ( ~n12574 & n12597 ) | ( n12588 & n12597 ) ;
  assign n13431 = n12590 & n13430 ;
  assign n13432 = n13429 & ~n13431 ;
  assign n13433 = n4781 & n12580 ;
  assign n13434 = n4776 & ~n12344 ;
  assign n13435 = n4778 & ~n12586 ;
  assign n13436 = n13434 | n13435 ;
  assign n13437 = n13433 | n13436 ;
  assign n13438 = n4784 | n13437 ;
  assign n13439 = ( n13432 & n13437 ) | ( n13432 & n13438 ) | ( n13437 & n13438 ) ;
  assign n13440 = x20 & n13439 ;
  assign n13441 = x20 & ~n13440 ;
  assign n13442 = ( n13439 & ~n13440 ) | ( n13439 & n13441 ) | ( ~n13440 & n13441 ) ;
  assign n13443 = n13428 & n13442 ;
  assign n13444 = n13428 & ~n13443 ;
  assign n13445 = n13110 | n13336 ;
  assign n13446 = n13109 & ~n13445 ;
  assign n13447 = n13337 | n13446 ;
  assign n13448 = n4781 & ~n12586 ;
  assign n13449 = n4776 & n12340 ;
  assign n13450 = n4778 & ~n12344 ;
  assign n13451 = n13449 | n13450 ;
  assign n13452 = n13448 | n13451 ;
  assign n13453 = ~n12588 & n12597 ;
  assign n13454 = ~n12574 & n13453 ;
  assign n13455 = n12574 & ~n13453 ;
  assign n13456 = ( n4784 & n13454 ) | ( n4784 & n13455 ) | ( n13454 & n13455 ) ;
  assign n13457 = n13452 | n13456 ;
  assign n13458 = x20 | n13457 ;
  assign n13459 = ~x20 & n13458 ;
  assign n13460 = ( ~n13457 & n13458 ) | ( ~n13457 & n13459 ) | ( n13458 & n13459 ) ;
  assign n13461 = ~n13447 & n13460 ;
  assign n13462 = n13447 | n13461 ;
  assign n13463 = n13447 & n13460 ;
  assign n13464 = ( ~n13334 & n13335 ) | ( ~n13334 & n13336 ) | ( n13335 & n13336 ) ;
  assign n13465 = ~n13309 & n13311 ;
  assign n13466 = n13312 | n13465 ;
  assign n13467 = n4484 & ~n12360 ;
  assign n13468 = n4479 & n12375 ;
  assign n13469 = n4481 & n12520 ;
  assign n13470 = n13468 | n13469 ;
  assign n13471 = n13467 | n13470 ;
  assign n13472 = n4487 | n13471 ;
  assign n13473 = ( ~n12902 & n13471 ) | ( ~n12902 & n13472 ) | ( n13471 & n13472 ) ;
  assign n13474 = ~x26 & n13473 ;
  assign n13475 = x26 | n13474 ;
  assign n13476 = ( ~n13473 & n13474 ) | ( ~n13473 & n13475 ) | ( n13474 & n13475 ) ;
  assign n13477 = ~n13466 & n13476 ;
  assign n13478 = n13151 & ~n13307 ;
  assign n13479 = n13308 | n13478 ;
  assign n13480 = n4048 & n12378 ;
  assign n13481 = n4043 & n12387 ;
  assign n13482 = n4045 & ~n12502 ;
  assign n13483 = n13481 | n13482 ;
  assign n13484 = n13480 | n13483 ;
  assign n13485 = n4051 | n13484 ;
  assign n13486 = ( ~n12816 & n13484 ) | ( ~n12816 & n13485 ) | ( n13484 & n13485 ) ;
  assign n13487 = ~x29 & n13486 ;
  assign n13488 = x29 | n13487 ;
  assign n13489 = ( ~n13486 & n13487 ) | ( ~n13486 & n13488 ) | ( n13487 & n13488 ) ;
  assign n13490 = ~n13479 & n13489 ;
  assign n13491 = n4484 & n12520 ;
  assign n13492 = n4479 & ~n12371 ;
  assign n13493 = n4481 & n12375 ;
  assign n13494 = n13492 | n13493 ;
  assign n13495 = n13491 | n13494 ;
  assign n13496 = n4487 & n12837 ;
  assign n13497 = ( n4487 & n12835 ) | ( n4487 & n13496 ) | ( n12835 & n13496 ) ;
  assign n13498 = n13495 | n13497 ;
  assign n13499 = x26 | n13498 ;
  assign n13500 = ~x26 & n13499 ;
  assign n13501 = ( ~n13498 & n13499 ) | ( ~n13498 & n13500 ) | ( n13499 & n13500 ) ;
  assign n13502 = n13479 | n13490 ;
  assign n13503 = ( ~n13489 & n13490 ) | ( ~n13489 & n13502 ) | ( n13490 & n13502 ) ;
  assign n13504 = n13501 & ~n13503 ;
  assign n13505 = n13490 | n13504 ;
  assign n13506 = n13466 | n13477 ;
  assign n13507 = ( ~n13476 & n13477 ) | ( ~n13476 & n13506 ) | ( n13477 & n13506 ) ;
  assign n13508 = n13505 & ~n13507 ;
  assign n13509 = n13477 | n13508 ;
  assign n13510 = n4551 & n12355 ;
  assign n13511 = n4546 & ~n12537 ;
  assign n13512 = n4548 & n12351 ;
  assign n13513 = n13511 | n13512 ;
  assign n13514 = n13510 | n13513 ;
  assign n13515 = n4554 | n13514 ;
  assign n13516 = ( n13409 & n13514 ) | ( n13409 & n13515 ) | ( n13514 & n13515 ) ;
  assign n13517 = x23 & n13516 ;
  assign n13518 = x23 & ~n13517 ;
  assign n13519 = ( n13516 & ~n13517 ) | ( n13516 & n13518 ) | ( ~n13517 & n13518 ) ;
  assign n13520 = ( n13321 & ~n13509 ) | ( n13321 & n13519 ) | ( ~n13509 & n13519 ) ;
  assign n13521 = ( ~n13321 & n13509 ) | ( ~n13321 & n13520 ) | ( n13509 & n13520 ) ;
  assign n13522 = n12347 & ~n12572 ;
  assign n13523 = n12573 | n13522 ;
  assign n13524 = n4781 & ~n12344 ;
  assign n13525 = n4776 & n12553 ;
  assign n13526 = n4778 & n12340 ;
  assign n13527 = n13525 | n13526 ;
  assign n13528 = n13524 | n13527 ;
  assign n13529 = n4784 | n13528 ;
  assign n13530 = ( ~n13523 & n13528 ) | ( ~n13523 & n13529 ) | ( n13528 & n13529 ) ;
  assign n13531 = ~x20 & n13530 ;
  assign n13532 = x20 | n13531 ;
  assign n13533 = ( ~n13530 & n13531 ) | ( ~n13530 & n13532 ) | ( n13531 & n13532 ) ;
  assign n13534 = ( n13464 & ~n13521 ) | ( n13464 & n13533 ) | ( ~n13521 & n13533 ) ;
  assign n13535 = ( ~n13464 & n13521 ) | ( ~n13464 & n13534 ) | ( n13521 & n13534 ) ;
  assign n13536 = ( ~n13462 & n13463 ) | ( ~n13462 & n13535 ) | ( n13463 & n13535 ) ;
  assign n13537 = n13461 | n13536 ;
  assign n13538 = ~n13428 & n13442 ;
  assign n13539 = ( n13444 & n13537 ) | ( n13444 & n13538 ) | ( n13537 & n13538 ) ;
  assign n13540 = n13537 | n13538 ;
  assign n13541 = n13444 | n13540 ;
  assign n13542 = ~n13539 & n13541 ;
  assign n13543 = ~n12331 & n12603 ;
  assign n13544 = n12604 | n13543 ;
  assign n13545 = n5083 & ~n12328 ;
  assign n13546 = n5069 & ~n12335 ;
  assign n13547 = n5070 & ~n12325 ;
  assign n13548 = n13546 | n13547 ;
  assign n13549 = n13545 | n13548 ;
  assign n13550 = n5074 | n13549 ;
  assign n13551 = ( ~n13544 & n13549 ) | ( ~n13544 & n13550 ) | ( n13549 & n13550 ) ;
  assign n13552 = ~x17 & n13551 ;
  assign n13553 = x17 | n13552 ;
  assign n13554 = ( ~n13551 & n13552 ) | ( ~n13551 & n13553 ) | ( n13552 & n13553 ) ;
  assign n13555 = n13542 & n13554 ;
  assign n13556 = n13539 | n13555 ;
  assign n13557 = n12621 & n13556 ;
  assign n13558 = n12621 | n13556 ;
  assign n13559 = ~n13557 & n13558 ;
  assign n13560 = n5069 & ~n12325 ;
  assign n13561 = n5070 & ~n12328 ;
  assign n13562 = n13560 | n13561 ;
  assign n13563 = n5083 & n12608 ;
  assign n13564 = n13562 | n13563 ;
  assign n13565 = n12329 & ~n12604 ;
  assign n13566 = n12328 & ~n12608 ;
  assign n13567 = n12609 | n13566 ;
  assign n13568 = ~n13565 & n13567 ;
  assign n13569 = n12610 & ~n13566 ;
  assign n13570 = ~n12604 & n13569 ;
  assign n13571 = n5074 & n13570 ;
  assign n13572 = ( n5074 & n13568 ) | ( n5074 & n13571 ) | ( n13568 & n13571 ) ;
  assign n13573 = n13564 | n13572 ;
  assign n13574 = x17 | n13573 ;
  assign n13575 = ~x17 & n13574 ;
  assign n13576 = ( ~n13573 & n13574 ) | ( ~n13573 & n13575 ) | ( n13574 & n13575 ) ;
  assign n13577 = n13426 | n13443 ;
  assign n13578 = n4781 & ~n12335 ;
  assign n13579 = n4776 & ~n12586 ;
  assign n13580 = n4778 & n12580 ;
  assign n13581 = n13579 | n13580 ;
  assign n13582 = n13578 | n13581 ;
  assign n13583 = ( ~n12574 & n12594 ) | ( ~n12574 & n12599 ) | ( n12594 & n12599 ) ;
  assign n13584 = ~n12587 & n13429 ;
  assign n13585 = n13583 & ~n13584 ;
  assign n13586 = ( ~n12574 & n12595 ) | ( ~n12574 & n12600 ) | ( n12595 & n12600 ) ;
  assign n13587 = ~n12582 & n13586 ;
  assign n13588 = n4784 & n13587 ;
  assign n13589 = ( n4784 & n13585 ) | ( n4784 & n13588 ) | ( n13585 & n13588 ) ;
  assign n13590 = n13582 | n13589 ;
  assign n13591 = x20 | n13590 ;
  assign n13592 = ~x20 & n13591 ;
  assign n13593 = ( ~n13590 & n13591 ) | ( ~n13590 & n13592 ) | ( n13591 & n13592 ) ;
  assign n13594 = ( n13353 & n13354 ) | ( n13353 & n13422 ) | ( n13354 & n13422 ) ;
  assign n13595 = ( n13404 & n13405 ) | ( n13404 & n13419 ) | ( n13405 & n13419 ) ;
  assign n13596 = n13372 & ~n13383 ;
  assign n13597 = n3636 & n12837 ;
  assign n13598 = ( n3636 & n12835 ) | ( n3636 & n13597 ) | ( n12835 & n13597 ) ;
  assign n13599 = n875 | n3121 ;
  assign n13600 = n4915 | n13599 ;
  assign n13601 = n258 | n590 ;
  assign n13602 = n442 | n602 ;
  assign n13603 = n13601 | n13602 ;
  assign n13604 = n181 | n408 ;
  assign n13605 = n13603 | n13604 ;
  assign n13606 = n820 | n13605 ;
  assign n13607 = n13600 | n13606 ;
  assign n13608 = n1069 | n1316 ;
  assign n13609 = n1054 | n13608 ;
  assign n13610 = n1314 | n13609 ;
  assign n13611 = n635 | n13610 ;
  assign n13612 = n13607 | n13611 ;
  assign n13613 = n296 | n484 ;
  assign n13614 = n96 | n13613 ;
  assign n13615 = n224 | n13614 ;
  assign n13616 = n13612 | n13615 ;
  assign n13617 = n1160 | n2344 ;
  assign n13618 = n11370 | n13617 ;
  assign n13619 = n1845 | n2623 ;
  assign n13620 = n373 | n13619 ;
  assign n13621 = n13618 | n13620 ;
  assign n13622 = n435 | n468 ;
  assign n13623 = n390 | n13622 ;
  assign n13624 = n1888 | n13623 ;
  assign n13625 = n11162 | n13624 ;
  assign n13626 = n13621 | n13625 ;
  assign n13627 = n2270 | n13626 ;
  assign n13628 = n571 | n13627 ;
  assign n13629 = n13616 | n13628 ;
  assign n13630 = n1194 | n1284 ;
  assign n13631 = n2089 | n13630 ;
  assign n13632 = n13629 | n13631 ;
  assign n13633 = n2943 | n3856 ;
  assign n13634 = n479 | n13633 ;
  assign n13635 = n273 | n13634 ;
  assign n13636 = n417 | n13635 ;
  assign n13637 = n607 | n13636 ;
  assign n13638 = n582 | n13637 ;
  assign n13639 = n92 | n13638 ;
  assign n13640 = n175 | n13639 ;
  assign n13641 = n13632 | n13640 ;
  assign n13642 = n122 | n13641 ;
  assign n13643 = n13371 & ~n13642 ;
  assign n13644 = n3744 & n12520 ;
  assign n13645 = n3639 & ~n12371 ;
  assign n13646 = n3727 & n12375 ;
  assign n13647 = n13645 | n13646 ;
  assign n13648 = n13644 | n13647 ;
  assign n13649 = ( ~n13371 & n13642 ) | ( ~n13371 & n13648 ) | ( n13642 & n13648 ) ;
  assign n13650 = n13643 | n13649 ;
  assign n13651 = n13598 | n13650 ;
  assign n13652 = n13596 | n13651 ;
  assign n13653 = ~n13371 & n13642 ;
  assign n13654 = n13643 | n13653 ;
  assign n13655 = n13598 | n13648 ;
  assign n13656 = n13654 & n13655 ;
  assign n13657 = ( n13596 & n13652 ) | ( n13596 & ~n13656 ) | ( n13652 & ~n13656 ) ;
  assign n13658 = n13596 & n13651 ;
  assign n13659 = ~n13656 & n13658 ;
  assign n13660 = n13657 & ~n13659 ;
  assign n13661 = n13387 | n13400 ;
  assign n13662 = n13660 & n13661 ;
  assign n13663 = n13660 | n13661 ;
  assign n13664 = ~n13662 & n13663 ;
  assign n13665 = n4048 & ~n12537 ;
  assign n13666 = n4043 & ~n12360 ;
  assign n13667 = n4045 & n12364 ;
  assign n13668 = n13666 | n13667 ;
  assign n13669 = n13665 | n13668 ;
  assign n13670 = ( n4051 & n13081 ) | ( n4051 & ~n13082 ) | ( n13081 & ~n13082 ) ;
  assign n13671 = n13669 | n13670 ;
  assign n13672 = x29 | n13671 ;
  assign n13673 = ~x29 & n13672 ;
  assign n13674 = ( ~n13671 & n13672 ) | ( ~n13671 & n13673 ) | ( n13672 & n13673 ) ;
  assign n13675 = n13664 & n13674 ;
  assign n13676 = n13664 & ~n13675 ;
  assign n13677 = ~n13664 & n13674 ;
  assign n13678 = n13676 | n13677 ;
  assign n13679 = n4484 & n12558 ;
  assign n13680 = n4479 & n12351 ;
  assign n13681 = n4481 & n12355 ;
  assign n13682 = n13680 | n13681 ;
  assign n13683 = n13679 | n13682 ;
  assign n13684 = n4487 | n13683 ;
  assign n13685 = ( n13330 & n13683 ) | ( n13330 & n13684 ) | ( n13683 & n13684 ) ;
  assign n13686 = x26 & n13685 ;
  assign n13687 = x26 & ~n13686 ;
  assign n13688 = ( n13685 & ~n13686 ) | ( n13685 & n13687 ) | ( ~n13686 & n13687 ) ;
  assign n13689 = n13678 & n13688 ;
  assign n13690 = n13678 | n13688 ;
  assign n13691 = ~n13689 & n13690 ;
  assign n13692 = n4551 & ~n12344 ;
  assign n13693 = n4546 & n12553 ;
  assign n13694 = n4548 & n12340 ;
  assign n13695 = n13693 | n13694 ;
  assign n13696 = n13692 | n13695 ;
  assign n13697 = n4554 | n13696 ;
  assign n13698 = ( ~n13523 & n13696 ) | ( ~n13523 & n13697 ) | ( n13696 & n13697 ) ;
  assign n13699 = ~x23 & n13698 ;
  assign n13700 = x23 | n13699 ;
  assign n13701 = ( ~n13698 & n13699 ) | ( ~n13698 & n13700 ) | ( n13699 & n13700 ) ;
  assign n13702 = ( n13595 & n13691 ) | ( n13595 & n13701 ) | ( n13691 & n13701 ) ;
  assign n13703 = ( n13691 & n13701 ) | ( n13691 & ~n13702 ) | ( n13701 & ~n13702 ) ;
  assign n13704 = ( n13595 & ~n13702 ) | ( n13595 & n13703 ) | ( ~n13702 & n13703 ) ;
  assign n13705 = ( n13593 & ~n13594 ) | ( n13593 & n13704 ) | ( ~n13594 & n13704 ) ;
  assign n13706 = ( n13594 & ~n13704 ) | ( n13594 & n13705 ) | ( ~n13704 & n13705 ) ;
  assign n13707 = ( ~n13593 & n13705 ) | ( ~n13593 & n13706 ) | ( n13705 & n13706 ) ;
  assign n13708 = ( n13576 & ~n13577 ) | ( n13576 & n13707 ) | ( ~n13577 & n13707 ) ;
  assign n13709 = ( n13577 & ~n13707 ) | ( n13577 & n13708 ) | ( ~n13707 & n13708 ) ;
  assign n13710 = ( ~n13576 & n13708 ) | ( ~n13576 & n13709 ) | ( n13708 & n13709 ) ;
  assign n13711 = n13559 & n13710 ;
  assign n13712 = n13710 & ~n13711 ;
  assign n13713 = ( n13559 & ~n13711 ) | ( n13559 & n13712 ) | ( ~n13711 & n13712 ) ;
  assign n13714 = n13542 & ~n13555 ;
  assign n13715 = ~n13542 & n13554 ;
  assign n13716 = n13463 | n13535 ;
  assign n13717 = n13462 & ~n13716 ;
  assign n13718 = n13536 | n13717 ;
  assign n13719 = ~n12576 & n13586 ;
  assign n13720 = n12602 | n13719 ;
  assign n13721 = n5083 & ~n12325 ;
  assign n13722 = n5069 & n12580 ;
  assign n13723 = n5070 & ~n12335 ;
  assign n13724 = n13722 | n13723 ;
  assign n13725 = n13721 | n13724 ;
  assign n13726 = n5074 | n13725 ;
  assign n13727 = ( ~n13720 & n13725 ) | ( ~n13720 & n13726 ) | ( n13725 & n13726 ) ;
  assign n13728 = ~x17 & n13727 ;
  assign n13729 = x17 | n13728 ;
  assign n13730 = ( ~n13727 & n13728 ) | ( ~n13727 & n13729 ) | ( n13728 & n13729 ) ;
  assign n13731 = ~n13718 & n13730 ;
  assign n13732 = ( ~n13533 & n13534 ) | ( ~n13533 & n13535 ) | ( n13534 & n13535 ) ;
  assign n13733 = ( ~n13519 & n13520 ) | ( ~n13519 & n13521 ) | ( n13520 & n13521 ) ;
  assign n13734 = ~n13505 & n13507 ;
  assign n13735 = n13508 | n13734 ;
  assign n13736 = n4551 & n12351 ;
  assign n13737 = n4546 & n12364 ;
  assign n13738 = n4548 & ~n12537 ;
  assign n13739 = n13737 | n13738 ;
  assign n13740 = n13736 | n13739 ;
  assign n13741 = n4554 & ~n12928 ;
  assign n13742 = ( n4554 & n12925 ) | ( n4554 & n13741 ) | ( n12925 & n13741 ) ;
  assign n13743 = n13740 | n13742 ;
  assign n13744 = x23 | n13743 ;
  assign n13745 = ~x23 & n13744 ;
  assign n13746 = ( ~n13743 & n13744 ) | ( ~n13743 & n13745 ) | ( n13744 & n13745 ) ;
  assign n13747 = ~n13735 & n13746 ;
  assign n13748 = n13735 | n13747 ;
  assign n13749 = n13735 & n13746 ;
  assign n13750 = n13295 | n13305 ;
  assign n13751 = ~n13306 & n13750 ;
  assign n13752 = ( n12981 & n13188 ) | ( n12981 & ~n13287 ) | ( n13188 & ~n13287 ) ;
  assign n13753 = ( ~n12981 & n13287 ) | ( ~n12981 & n13752 ) | ( n13287 & n13752 ) ;
  assign n13754 = ( ~n13188 & n13752 ) | ( ~n13188 & n13753 ) | ( n13752 & n13753 ) ;
  assign n13755 = n3744 & n12415 ;
  assign n13756 = n3639 & n12419 ;
  assign n13757 = n3727 & n12411 ;
  assign n13758 = n13756 | n13757 ;
  assign n13759 = n13755 | n13758 ;
  assign n13760 = n12416 & ~n12490 ;
  assign n13761 = ~n12489 & n13760 ;
  assign n13762 = n12488 & ~n13760 ;
  assign n13763 = ( n3636 & n13761 ) | ( n3636 & n13762 ) | ( n13761 & n13762 ) ;
  assign n13764 = n13759 | n13763 ;
  assign n13765 = ~n13754 & n13764 ;
  assign n13766 = n13754 | n13765 ;
  assign n13767 = n13754 & n13764 ;
  assign n13768 = n13766 & ~n13767 ;
  assign n13769 = n13212 & ~n13286 ;
  assign n13770 = ~n13285 & n13769 ;
  assign n13771 = n13284 & ~n13769 ;
  assign n13772 = n13770 | n13771 ;
  assign n13773 = ( n12425 & n12426 ) | ( n12425 & n12487 ) | ( n12426 & n12487 ) ;
  assign n13774 = n12424 | n12425 ;
  assign n13775 = n12487 | n13774 ;
  assign n13776 = ~n13773 & n13775 ;
  assign n13777 = n3744 & n12411 ;
  assign n13778 = n3639 & ~n12423 ;
  assign n13779 = n3727 & n12419 ;
  assign n13780 = n13778 | n13779 ;
  assign n13781 = n13777 | n13780 ;
  assign n13782 = n3636 | n13781 ;
  assign n13783 = ( n13776 & n13781 ) | ( n13776 & n13782 ) | ( n13781 & n13782 ) ;
  assign n13784 = n13772 | n13783 ;
  assign n13785 = ~n12483 & n12485 ;
  assign n13786 = n12486 | n13785 ;
  assign n13787 = n3744 & ~n12423 ;
  assign n13788 = n3727 & n12433 ;
  assign n13789 = n3639 & ~n12438 ;
  assign n13790 = n13788 | n13789 ;
  assign n13791 = n13787 | n13790 ;
  assign n13792 = n3636 | n13791 ;
  assign n13793 = ( ~n13786 & n13791 ) | ( ~n13786 & n13792 ) | ( n13791 & n13792 ) ;
  assign n13794 = n2695 | n11372 ;
  assign n13795 = n2688 | n13794 ;
  assign n13796 = n849 | n2158 ;
  assign n13797 = n13795 | n13796 ;
  assign n13798 = n1210 | n13797 ;
  assign n13799 = n1199 | n13798 ;
  assign n13800 = n12725 | n13799 ;
  assign n13801 = n3893 | n13800 ;
  assign n13802 = n174 | n655 ;
  assign n13803 = n11073 | n13802 ;
  assign n13804 = n345 | n451 ;
  assign n13805 = n449 | n13804 ;
  assign n13806 = n13803 | n13805 ;
  assign n13807 = n661 | n13806 ;
  assign n13808 = n960 | n13807 ;
  assign n13809 = n635 | n13808 ;
  assign n13810 = n718 | n13809 ;
  assign n13811 = n314 | n13810 ;
  assign n13812 = n291 | n13811 ;
  assign n13813 = n13801 | n13812 ;
  assign n13814 = n46 | n569 ;
  assign n13815 = n76 | n13814 ;
  assign n13816 = n13813 | n13815 ;
  assign n13817 = n13793 & n13816 ;
  assign n13818 = n13793 & ~n13817 ;
  assign n13819 = ~n13793 & n13816 ;
  assign n13820 = n13818 | n13819 ;
  assign n13821 = n12449 | n12479 ;
  assign n13822 = ~n12480 & n13821 ;
  assign n13823 = n3744 & n12440 ;
  assign n13824 = n3727 & n12446 ;
  assign n13825 = n3639 & n12452 ;
  assign n13826 = n13824 | n13825 ;
  assign n13827 = n13823 | n13826 ;
  assign n13828 = n3636 | n13827 ;
  assign n13829 = ( n13822 & n13827 ) | ( n13822 & n13828 ) | ( n13827 & n13828 ) ;
  assign n13830 = n878 | n1430 ;
  assign n13831 = n11208 | n13830 ;
  assign n13832 = n11405 | n13831 ;
  assign n13833 = n11190 | n13832 ;
  assign n13834 = n3520 | n5640 ;
  assign n13835 = n13833 | n13834 ;
  assign n13836 = n93 | n1271 ;
  assign n13837 = n265 | n489 ;
  assign n13838 = n441 | n13837 ;
  assign n13839 = n13836 | n13838 ;
  assign n13840 = n120 | n13839 ;
  assign n13841 = n311 | n5703 ;
  assign n13842 = n1644 | n13841 ;
  assign n13843 = n130 | n13842 ;
  assign n13844 = n13840 | n13843 ;
  assign n13845 = n429 | n13844 ;
  assign n13846 = n282 | n13845 ;
  assign n13847 = n276 | n13846 ;
  assign n13848 = n13835 | n13847 ;
  assign n13849 = n46 | n62 ;
  assign n13850 = n172 | n13849 ;
  assign n13851 = n13848 | n13850 ;
  assign n13852 = n13829 & n13851 ;
  assign n13853 = n13829 & ~n13852 ;
  assign n13854 = ~n13829 & n13851 ;
  assign n13855 = n13853 | n13854 ;
  assign n13856 = n3744 & n12446 ;
  assign n13857 = n3727 & n12452 ;
  assign n13858 = n3639 & n12454 ;
  assign n13859 = n13857 | n13858 ;
  assign n13860 = n13856 | n13859 ;
  assign n13861 = ( n12446 & n12452 ) | ( n12446 & ~n12479 ) | ( n12452 & ~n12479 ) ;
  assign n13862 = ( n12478 & ~n12479 ) | ( n12478 & n13861 ) | ( ~n12479 & n13861 ) ;
  assign n13863 = n3636 | n13860 ;
  assign n13864 = ( n13860 & n13862 ) | ( n13860 & n13863 ) | ( n13862 & n13863 ) ;
  assign n13865 = n2178 | n12639 ;
  assign n13866 = n255 | n4304 ;
  assign n13867 = n13865 | n13866 ;
  assign n13868 = n5703 | n13867 ;
  assign n13869 = n144 | n305 ;
  assign n13870 = n13868 | n13869 ;
  assign n13871 = n609 | n1284 ;
  assign n13872 = n862 | n13871 ;
  assign n13873 = n237 | n13872 ;
  assign n13874 = n52 | n13873 ;
  assign n13875 = n140 | n13874 ;
  assign n13876 = n13870 | n13875 ;
  assign n13877 = n146 | n13876 ;
  assign n13878 = n1432 | n2721 ;
  assign n13879 = n218 | n384 ;
  assign n13880 = n10899 | n13879 ;
  assign n13881 = n13878 | n13880 ;
  assign n13882 = n6016 | n13881 ;
  assign n13883 = n13621 | n13623 ;
  assign n13884 = n13882 | n13883 ;
  assign n13885 = n272 | n13884 ;
  assign n13886 = n1866 | n13885 ;
  assign n13887 = n13877 | n13886 ;
  assign n13888 = n344 | n583 ;
  assign n13889 = n437 | n13888 ;
  assign n13890 = n2904 | n13889 ;
  assign n13891 = n1200 | n3856 ;
  assign n13892 = n13890 | n13891 ;
  assign n13893 = n11382 | n13892 ;
  assign n13894 = n5548 | n13893 ;
  assign n13895 = n499 | n2943 ;
  assign n13896 = n310 | n13895 ;
  assign n13897 = n355 | n13896 ;
  assign n13898 = n569 | n13897 ;
  assign n13899 = n103 | n13898 ;
  assign n13900 = n13894 | n13899 ;
  assign n13901 = n168 | n223 ;
  assign n13902 = n13900 | n13901 ;
  assign n13903 = n430 | n1372 ;
  assign n13904 = n93 | n13903 ;
  assign n13905 = n13902 | n13904 ;
  assign n13906 = n13887 | n13905 ;
  assign n13907 = n539 | n636 ;
  assign n13908 = n380 | n13907 ;
  assign n13909 = n458 | n13908 ;
  assign n13910 = n160 | n13909 ;
  assign n13911 = n85 | n13910 ;
  assign n13912 = n13906 | n13911 ;
  assign n13913 = n13864 & n13912 ;
  assign n13914 = n13864 & ~n13913 ;
  assign n13915 = ~n13864 & n13912 ;
  assign n13916 = n13914 | n13915 ;
  assign n13917 = n12452 | n12454 ;
  assign n13918 = ~n12478 & n13917 ;
  assign n13919 = n12452 & n12454 ;
  assign n13920 = n13917 & ~n13919 ;
  assign n13921 = n12477 | n13920 ;
  assign n13922 = ~n13918 & n13921 ;
  assign n13923 = n3744 & n12452 ;
  assign n13924 = n3727 & n12454 ;
  assign n13925 = n3639 & ~n12456 ;
  assign n13926 = n13924 | n13925 ;
  assign n13927 = n13923 | n13926 ;
  assign n13928 = n3636 | n13927 ;
  assign n13929 = ( ~n13922 & n13927 ) | ( ~n13922 & n13928 ) | ( n13927 & n13928 ) ;
  assign n13930 = n498 | n621 ;
  assign n13931 = n364 | n13930 ;
  assign n13932 = n1434 | n2515 ;
  assign n13933 = n13931 | n13932 ;
  assign n13934 = n1041 | n1271 ;
  assign n13935 = n13933 | n13934 ;
  assign n13936 = n225 | n1115 ;
  assign n13937 = n529 | n13936 ;
  assign n13938 = n349 | n13937 ;
  assign n13939 = n13935 | n13938 ;
  assign n13940 = n129 | n582 ;
  assign n13941 = n649 | n13940 ;
  assign n13942 = n13939 | n13941 ;
  assign n13943 = n988 | n11080 ;
  assign n13944 = n512 | n1177 ;
  assign n13945 = ( ~n13942 & n13943 ) | ( ~n13942 & n13944 ) | ( n13943 & n13944 ) ;
  assign n13946 = n13942 | n13945 ;
  assign n13947 = n12777 | n13946 ;
  assign n13948 = n12772 & ~n13947 ;
  assign n13949 = n3655 | n13243 ;
  assign n13950 = n1442 | n13949 ;
  assign n13951 = n834 | n13950 ;
  assign n13952 = n669 | n13951 ;
  assign n13953 = n13948 & ~n13952 ;
  assign n13954 = n326 | n3456 ;
  assign n13955 = n274 | n13954 ;
  assign n13956 = n345 | n13955 ;
  assign n13957 = n592 | n13956 ;
  assign n13958 = n108 | n13957 ;
  assign n13959 = n646 | n13958 ;
  assign n13960 = n13953 & ~n13959 ;
  assign n13961 = n1596 | n2515 ;
  assign n13962 = n1972 | n13961 ;
  assign n13963 = n3470 | n13962 ;
  assign n13964 = n2080 | n13963 ;
  assign n13965 = n5751 | n13964 ;
  assign n13966 = n2331 & ~n13965 ;
  assign n13967 = n474 | n752 ;
  assign n13968 = n10956 | n13967 ;
  assign n13969 = n710 | n3393 ;
  assign n13970 = n13968 | n13969 ;
  assign n13971 = n244 | n2164 ;
  assign n13972 = n3109 | n13971 ;
  assign n13973 = n307 | n310 ;
  assign n13974 = n610 | n13973 ;
  assign n13975 = n96 | n13974 ;
  assign n13976 = n13972 | n13975 ;
  assign n13977 = n13840 | n13976 ;
  assign n13978 = n13970 | n13977 ;
  assign n13979 = n169 | n2393 ;
  assign n13980 = n260 | n13979 ;
  assign n13981 = n419 | n13980 ;
  assign n13982 = n218 | n13981 ;
  assign n13983 = n650 | n13982 ;
  assign n13984 = n13978 | n13983 ;
  assign n13985 = n2026 | n2219 ;
  assign n13986 = n13984 | n13985 ;
  assign n13987 = n13966 & ~n13986 ;
  assign n13988 = n326 | n528 ;
  assign n13989 = n607 | n13988 ;
  assign n13990 = n451 | n13989 ;
  assign n13991 = n108 | n13990 ;
  assign n13992 = n13987 & ~n13991 ;
  assign n13993 = n12466 & ~n12468 ;
  assign n13994 = n12469 | n13993 ;
  assign n13995 = n3727 & ~n12468 ;
  assign n13996 = n3636 | n13995 ;
  assign n13997 = ( n13994 & n13995 ) | ( n13994 & n13996 ) | ( n13995 & n13996 ) ;
  assign n13998 = n3744 & ~n12466 ;
  assign n13999 = n13997 | n13998 ;
  assign n14000 = ~n13992 & n13999 ;
  assign n14001 = ~n13960 & n14000 ;
  assign n14002 = n12459 & ~n12469 ;
  assign n14003 = n12470 | n14002 ;
  assign n14004 = n3636 & n14003 ;
  assign n14005 = n3744 & n12459 ;
  assign n14006 = n3639 & ~n12468 ;
  assign n14007 = n3727 & ~n12466 ;
  assign n14008 = n14006 | n14007 ;
  assign n14009 = n14005 | n14008 ;
  assign n14010 = n14004 | n14009 ;
  assign n14011 = n13960 & ~n14000 ;
  assign n14012 = n14001 | n14011 ;
  assign n14013 = n14010 & ~n14012 ;
  assign n14014 = n14001 | n14013 ;
  assign n14015 = n243 | n311 ;
  assign n14016 = n498 | n14015 ;
  assign n14017 = n393 | n14016 ;
  assign n14018 = n592 | n14017 ;
  assign n14019 = n377 | n14018 ;
  assign n14020 = n1214 | n11361 ;
  assign n14021 = n2536 | n14020 ;
  assign n14022 = n5798 | n14021 ;
  assign n14023 = n4364 | n14022 ;
  assign n14024 = n157 | n3682 ;
  assign n14025 = n10878 | n14024 ;
  assign n14026 = n487 | n14025 ;
  assign n14027 = ( ~n4866 & n14023 ) | ( ~n4866 & n14026 ) | ( n14023 & n14026 ) ;
  assign n14028 = n4866 | n14027 ;
  assign n14029 = n14019 | n14028 ;
  assign n14030 = n12462 & n12471 ;
  assign n14031 = n12472 & ~n14030 ;
  assign n14032 = n3744 & ~n12456 ;
  assign n14033 = n3727 & n12459 ;
  assign n14034 = n3639 & ~n12466 ;
  assign n14035 = n14033 | n14034 ;
  assign n14036 = n14032 | n14035 ;
  assign n14037 = n3636 | n14036 ;
  assign n14038 = ( n14031 & n14036 ) | ( n14031 & n14037 ) | ( n14036 & n14037 ) ;
  assign n14039 = ( n14014 & n14029 ) | ( n14014 & n14038 ) | ( n14029 & n14038 ) ;
  assign n14040 = n12473 & n12475 ;
  assign n14041 = n12476 & ~n14040 ;
  assign n14042 = n3744 & n12454 ;
  assign n14043 = n3727 & ~n12456 ;
  assign n14044 = n3639 & n12459 ;
  assign n14045 = n14043 | n14044 ;
  assign n14046 = n14042 | n14045 ;
  assign n14047 = n3636 | n14046 ;
  assign n14048 = ( n14041 & n14046 ) | ( n14041 & n14047 ) | ( n14046 & n14047 ) ;
  assign n14049 = n436 | n2165 ;
  assign n14050 = n1632 | n14049 ;
  assign n14051 = n3896 | n14050 ;
  assign n14052 = n3283 | n14051 ;
  assign n14053 = n81 | n14052 ;
  assign n14054 = n2229 | n14053 ;
  assign n14055 = n1368 | n14054 ;
  assign n14056 = n2966 | n14055 ;
  assign n14057 = n282 | n409 ;
  assign n14058 = n1036 | n14057 ;
  assign n14059 = n451 | n14058 ;
  assign n14060 = n12790 | n14059 ;
  assign n14061 = n12789 | n14060 ;
  assign n14062 = n373 | n4879 ;
  assign n14063 = n3553 & ~n14062 ;
  assign n14064 = n521 | n580 ;
  assign n14065 = n14063 & ~n14064 ;
  assign n14066 = ~n166 & n14065 ;
  assign n14067 = ~n14061 & n14066 ;
  assign n14068 = n995 | n2333 ;
  assign n14069 = n169 | n14068 ;
  assign n14070 = n528 | n14069 ;
  assign n14071 = n337 | n14070 ;
  assign n14072 = n14067 & ~n14071 ;
  assign n14073 = n241 | n417 ;
  assign n14074 = n400 | n14073 ;
  assign n14075 = n199 | n14074 ;
  assign n14076 = n111 | n14075 ;
  assign n14077 = n207 | n14076 ;
  assign n14078 = n14072 & ~n14077 ;
  assign n14079 = ~n1416 & n14078 ;
  assign n14080 = ~n14056 & n14079 ;
  assign n14081 = n500 | n626 ;
  assign n14082 = n252 | n14081 ;
  assign n14083 = n579 | n14082 ;
  assign n14084 = n193 | n14083 ;
  assign n14085 = n14080 & ~n14084 ;
  assign n14086 = n14048 & ~n14085 ;
  assign n14087 = n14048 & ~n14086 ;
  assign n14088 = n14048 | n14085 ;
  assign n14089 = ( n14039 & ~n14087 ) | ( n14039 & n14088 ) | ( ~n14087 & n14088 ) ;
  assign n14090 = ( n14039 & n14088 ) | ( n14039 & ~n14089 ) | ( n14088 & ~n14089 ) ;
  assign n14091 = ( n14087 & n14089 ) | ( n14087 & ~n14090 ) | ( n14089 & ~n14090 ) ;
  assign n14092 = ( n14039 & n14086 ) | ( n14039 & n14091 ) | ( n14086 & n14091 ) ;
  assign n14093 = n10936 | n11054 ;
  assign n14094 = n77 | n14093 ;
  assign n14095 = n3217 | n14094 ;
  assign n14096 = n12673 & ~n14095 ;
  assign n14097 = ~n1069 & n14096 ;
  assign n14098 = n1337 | n1422 ;
  assign n14099 = n14097 & ~n14098 ;
  assign n14100 = n367 | n1959 ;
  assign n14101 = n2433 | n14100 ;
  assign n14102 = n996 | n14101 ;
  assign n14103 = n634 | n14102 ;
  assign n14104 = n62 | n14103 ;
  assign n14105 = n601 | n14104 ;
  assign n14106 = n450 | n14105 ;
  assign n14107 = n14099 & ~n14106 ;
  assign n14108 = n2332 | n2837 ;
  assign n14109 = n820 | n14108 ;
  assign n14110 = ( ~n11052 & n12268 ) | ( ~n11052 & n14109 ) | ( n12268 & n14109 ) ;
  assign n14111 = n11052 | n14110 ;
  assign n14112 = n1115 | n14111 ;
  assign n14113 = n421 | n14112 ;
  assign n14114 = n14107 & ~n14113 ;
  assign n14115 = n431 | n475 ;
  assign n14116 = n499 | n14115 ;
  assign n14117 = n301 | n14116 ;
  assign n14118 = n607 | n14117 ;
  assign n14119 = n213 | n14118 ;
  assign n14120 = n403 | n14119 ;
  assign n14121 = n14114 & ~n14120 ;
  assign n14122 = n13929 & ~n14121 ;
  assign n14123 = n13929 & ~n14122 ;
  assign n14124 = n13929 | n14121 ;
  assign n14125 = ~n14123 & n14124 ;
  assign n14126 = n14092 & n14125 ;
  assign n14127 = n14092 | n14125 ;
  assign n14128 = ~n14126 & n14127 ;
  assign n14129 = ( n13929 & n14092 ) | ( n13929 & n14128 ) | ( n14092 & n14128 ) ;
  assign n14130 = n13916 & n14129 ;
  assign n14131 = n13913 | n14130 ;
  assign n14132 = n13855 & n14131 ;
  assign n14133 = n13852 | n14132 ;
  assign n14134 = n298 | n2477 ;
  assign n14135 = n1576 | n14134 ;
  assign n14136 = n1719 | n14135 ;
  assign n14137 = n2596 | n14136 ;
  assign n14138 = n1707 | n14137 ;
  assign n14139 = n1316 | n14138 ;
  assign n14140 = n13235 | n14139 ;
  assign n14141 = n1644 | n3792 ;
  assign n14142 = n2867 | n14141 ;
  assign n14143 = n622 | n14142 ;
  assign n14144 = n500 | n14143 ;
  assign n14145 = n403 | n14144 ;
  assign n14146 = n175 | n14145 ;
  assign n14147 = n157 | n14146 ;
  assign n14148 = n14140 | n14147 ;
  assign n14149 = n3744 & ~n12438 ;
  assign n14150 = n3727 & n12440 ;
  assign n14151 = n3639 & n12446 ;
  assign n14152 = n14150 | n14151 ;
  assign n14153 = n14149 | n14152 ;
  assign n14154 = n12442 | n12482 ;
  assign n14155 = ~n12441 & n12481 ;
  assign n14156 = ( n12447 & n12480 ) | ( n12447 & ~n14155 ) | ( n12480 & ~n14155 ) ;
  assign n14157 = ( n3636 & ~n14154 ) | ( n3636 & n14156 ) | ( ~n14154 & n14156 ) ;
  assign n14158 = n14153 | n14157 ;
  assign n14159 = ( n14133 & n14148 ) | ( n14133 & n14158 ) | ( n14148 & n14158 ) ;
  assign n14160 = n3744 & n12433 ;
  assign n14161 = n3727 & ~n12438 ;
  assign n14162 = n3639 & n12440 ;
  assign n14163 = n14161 | n14162 ;
  assign n14164 = n14160 | n14163 ;
  assign n14165 = ( ~n12433 & n12438 ) | ( ~n12433 & n12482 ) | ( n12438 & n12482 ) ;
  assign n14166 = ( n12433 & ~n12482 ) | ( n12433 & n14165 ) | ( ~n12482 & n14165 ) ;
  assign n14167 = ( ~n12438 & n14165 ) | ( ~n12438 & n14166 ) | ( n14165 & n14166 ) ;
  assign n14168 = n3636 | n14164 ;
  assign n14169 = ( n14164 & ~n14167 ) | ( n14164 & n14168 ) | ( ~n14167 & n14168 ) ;
  assign n14170 = n3149 | n11276 ;
  assign n14171 = n2612 | n2689 ;
  assign n14172 = n14170 | n14171 ;
  assign n14173 = n2312 | n14172 ;
  assign n14174 = n5163 | n14173 ;
  assign n14175 = n10863 | n14174 ;
  assign n14176 = n1775 | n14175 ;
  assign n14177 = n3313 | n3329 ;
  assign n14178 = n14176 | n14177 ;
  assign n14179 = n611 | n3224 ;
  assign n14180 = n476 | n14179 ;
  assign n14181 = n283 | n14180 ;
  assign n14182 = n592 | n14181 ;
  assign n14183 = n46 | n14182 ;
  assign n14184 = n186 | n14183 ;
  assign n14185 = n649 | n14184 ;
  assign n14186 = n14178 | n14185 ;
  assign n14187 = n14169 & n14186 ;
  assign n14188 = n14169 & ~n14187 ;
  assign n14189 = ~n14169 & n14186 ;
  assign n14190 = n14188 | n14189 ;
  assign n14191 = n14159 & ~n14190 ;
  assign n14192 = ( n14159 & n14187 ) | ( n14159 & ~n14191 ) | ( n14187 & ~n14191 ) ;
  assign n14193 = n13820 & n14192 ;
  assign n14194 = ~n12981 & n13273 ;
  assign n14195 = n13284 | n14194 ;
  assign n14196 = n12981 & ~n13273 ;
  assign n14197 = ( n13283 & n14194 ) | ( n13283 & n14196 ) | ( n14194 & n14196 ) ;
  assign n14198 = n14195 & ~n14197 ;
  assign n14199 = n13817 & ~n14198 ;
  assign n14200 = ( n14193 & ~n14198 ) | ( n14193 & n14199 ) | ( ~n14198 & n14199 ) ;
  assign n14201 = ~n13817 & n14198 ;
  assign n14202 = ~n14193 & n14201 ;
  assign n14203 = n14200 | n14202 ;
  assign n14204 = n4048 & n12401 ;
  assign n14205 = n4043 & n12411 ;
  assign n14206 = n4045 & n12415 ;
  assign n14207 = n14205 | n14206 ;
  assign n14208 = n14204 | n14207 ;
  assign n14209 = n4051 & ~n13163 ;
  assign n14210 = ~n13161 & n14209 ;
  assign n14211 = ( n4051 & n14208 ) | ( n4051 & ~n14210 ) | ( n14208 & ~n14210 ) ;
  assign n14212 = ~x29 & n14211 ;
  assign n14213 = x29 | n14212 ;
  assign n14214 = ( ~n14211 & n14212 ) | ( ~n14211 & n14213 ) | ( n14212 & n14213 ) ;
  assign n14215 = ~n14203 & n14214 ;
  assign n14216 = n14200 | n14215 ;
  assign n14217 = ( n13772 & ~n13783 ) | ( n13772 & n14216 ) | ( ~n13783 & n14216 ) ;
  assign n14218 = ( ~n13772 & n13783 ) | ( ~n13772 & n14217 ) | ( n13783 & n14217 ) ;
  assign n14219 = ( ~n14216 & n14217 ) | ( ~n14216 & n14218 ) | ( n14217 & n14218 ) ;
  assign n14220 = ( n13784 & n14216 ) | ( n13784 & ~n14219 ) | ( n14216 & ~n14219 ) ;
  assign n14221 = ~n13768 & n14220 ;
  assign n14222 = ( ~n13291 & n13765 ) | ( ~n13291 & n14221 ) | ( n13765 & n14221 ) ;
  assign n14223 = n13291 & ~n13765 ;
  assign n14224 = ~n14221 & n14223 ;
  assign n14225 = n14222 | n14224 ;
  assign n14226 = n4048 & n12387 ;
  assign n14227 = n4043 & n12392 ;
  assign n14228 = n4045 & n12383 ;
  assign n14229 = n14227 | n14228 ;
  assign n14230 = n14226 | n14229 ;
  assign n14231 = n4051 | n14230 ;
  assign n14232 = ( n12948 & n14230 ) | ( n12948 & n14231 ) | ( n14230 & n14231 ) ;
  assign n14233 = x29 & n14232 ;
  assign n14234 = x29 & ~n14233 ;
  assign n14235 = ( n14232 & ~n14233 ) | ( n14232 & n14234 ) | ( ~n14233 & n14234 ) ;
  assign n14236 = ~n14225 & n14235 ;
  assign n14237 = n14222 | n14236 ;
  assign n14238 = n4484 & n12375 ;
  assign n14239 = n4479 & n12378 ;
  assign n14240 = n4481 & ~n12371 ;
  assign n14241 = n14239 | n14240 ;
  assign n14242 = n14238 | n14241 ;
  assign n14243 = ( n4487 & n13064 ) | ( n4487 & ~n13065 ) | ( n13064 & ~n13065 ) ;
  assign n14244 = n14242 | n14243 ;
  assign n14245 = x26 | n14244 ;
  assign n14246 = ~x26 & n14245 ;
  assign n14247 = ( ~n14244 & n14245 ) | ( ~n14244 & n14246 ) | ( n14245 & n14246 ) ;
  assign n14248 = ( n13751 & n14237 ) | ( n13751 & n14247 ) | ( n14237 & n14247 ) ;
  assign n14249 = ~n13501 & n13503 ;
  assign n14250 = n13504 | n14249 ;
  assign n14251 = n4551 & ~n12537 ;
  assign n14252 = n4546 & ~n12360 ;
  assign n14253 = n4548 & n12364 ;
  assign n14254 = n14252 | n14253 ;
  assign n14255 = n14251 | n14254 ;
  assign n14256 = ( n4554 & n13081 ) | ( n4554 & ~n13082 ) | ( n13081 & ~n13082 ) ;
  assign n14257 = n14255 | n14256 ;
  assign n14258 = x23 | n14257 ;
  assign n14259 = ~x23 & n14258 ;
  assign n14260 = ( ~n14257 & n14258 ) | ( ~n14257 & n14259 ) | ( n14258 & n14259 ) ;
  assign n14261 = ( ~n14248 & n14250 ) | ( ~n14248 & n14260 ) | ( n14250 & n14260 ) ;
  assign n14262 = ( n14248 & ~n14250 ) | ( n14248 & n14261 ) | ( ~n14250 & n14261 ) ;
  assign n14263 = ( ~n13748 & n13749 ) | ( ~n13748 & n14262 ) | ( n13749 & n14262 ) ;
  assign n14264 = n13747 | n14263 ;
  assign n14265 = n4781 & n12340 ;
  assign n14266 = n4776 & n12558 ;
  assign n14267 = n4778 & n12553 ;
  assign n14268 = n14266 | n14267 ;
  assign n14269 = n14265 | n14268 ;
  assign n14270 = n4784 & n13347 ;
  assign n14271 = ( n4784 & n13346 ) | ( n4784 & n14270 ) | ( n13346 & n14270 ) ;
  assign n14272 = n14269 | n14271 ;
  assign n14273 = x20 | n14272 ;
  assign n14274 = ~x20 & n14273 ;
  assign n14275 = ( ~n14272 & n14273 ) | ( ~n14272 & n14274 ) | ( n14273 & n14274 ) ;
  assign n14276 = ( n13733 & ~n14264 ) | ( n13733 & n14275 ) | ( ~n14264 & n14275 ) ;
  assign n14277 = ( ~n13733 & n14264 ) | ( ~n13733 & n14276 ) | ( n14264 & n14276 ) ;
  assign n14278 = n5083 & ~n12335 ;
  assign n14279 = n5069 & ~n12586 ;
  assign n14280 = n5070 & n12580 ;
  assign n14281 = n14279 | n14280 ;
  assign n14282 = n14278 | n14281 ;
  assign n14283 = n5074 & n13587 ;
  assign n14284 = ( n5074 & n13585 ) | ( n5074 & n14283 ) | ( n13585 & n14283 ) ;
  assign n14285 = n14282 | n14284 ;
  assign n14286 = x17 | n14285 ;
  assign n14287 = ~x17 & n14286 ;
  assign n14288 = ( ~n14285 & n14286 ) | ( ~n14285 & n14287 ) | ( n14286 & n14287 ) ;
  assign n14289 = ( n13732 & ~n14277 ) | ( n13732 & n14288 ) | ( ~n14277 & n14288 ) ;
  assign n14290 = ( ~n13732 & n14277 ) | ( ~n13732 & n14289 ) | ( n14277 & n14289 ) ;
  assign n14291 = n13718 | n13731 ;
  assign n14292 = ( ~n13730 & n13731 ) | ( ~n13730 & n14291 ) | ( n13731 & n14291 ) ;
  assign n14293 = n14290 & ~n14292 ;
  assign n14294 = n13731 | n14293 ;
  assign n14295 = n13715 | n14294 ;
  assign n14296 = n13714 | n14295 ;
  assign n14297 = ( n12317 & n12604 ) | ( n12317 & n12614 ) | ( n12604 & n12614 ) ;
  assign n14298 = n12612 | n13566 ;
  assign n14299 = ( ~n12604 & n12613 ) | ( ~n12604 & n14298 ) | ( n12613 & n14298 ) ;
  assign n14300 = ~n12611 & n14299 ;
  assign n14301 = ~n12317 & n14300 ;
  assign n14302 = n14297 | n14301 ;
  assign n14303 = n7277 & ~n12318 ;
  assign n14304 = n5384 & n12608 ;
  assign n14305 = n14303 | n14304 ;
  assign n14306 = n7280 & ~n12314 ;
  assign n14307 = n14305 | n14306 ;
  assign n14308 = n39 | n14307 ;
  assign n14309 = ( ~n14302 & n14307 ) | ( ~n14302 & n14308 ) | ( n14307 & n14308 ) ;
  assign n14310 = ~x14 & n14309 ;
  assign n14311 = x14 | n14310 ;
  assign n14312 = ( ~n14309 & n14310 ) | ( ~n14309 & n14311 ) | ( n14310 & n14311 ) ;
  assign n14313 = ( n13714 & n13715 ) | ( n13714 & n14294 ) | ( n13715 & n14294 ) ;
  assign n14314 = ( n14296 & n14312 ) | ( n14296 & n14313 ) | ( n14312 & n14313 ) ;
  assign n14315 = n13713 & n14314 ;
  assign n14316 = n13713 | n14314 ;
  assign n14317 = ~n14315 & n14316 ;
  assign n14318 = ( ~n12604 & n12610 ) | ( ~n12604 & n13566 ) | ( n12610 & n13566 ) ;
  assign n14319 = n12612 & n14318 ;
  assign n14320 = n14299 & ~n14319 ;
  assign n14321 = n7280 & ~n12318 ;
  assign n14322 = n5384 & ~n12328 ;
  assign n14323 = n7277 & n12608 ;
  assign n14324 = n14322 | n14323 ;
  assign n14325 = n14321 | n14324 ;
  assign n14326 = n39 | n14325 ;
  assign n14327 = ( n14320 & n14325 ) | ( n14320 & n14326 ) | ( n14325 & n14326 ) ;
  assign n14328 = x14 & n14327 ;
  assign n14329 = x14 & ~n14328 ;
  assign n14330 = ( n14327 & ~n14328 ) | ( n14327 & n14329 ) | ( ~n14328 & n14329 ) ;
  assign n14331 = ( ~n14288 & n14289 ) | ( ~n14288 & n14290 ) | ( n14289 & n14290 ) ;
  assign n14332 = n5384 & ~n12325 ;
  assign n14333 = n7277 & ~n12328 ;
  assign n14334 = n14332 | n14333 ;
  assign n14335 = n7280 & n12608 ;
  assign n14336 = n14334 | n14335 ;
  assign n14337 = n39 & n13570 ;
  assign n14338 = ( n39 & n13568 ) | ( n39 & n14337 ) | ( n13568 & n14337 ) ;
  assign n14339 = n14336 | n14338 ;
  assign n14340 = x14 | n14339 ;
  assign n14341 = ~x14 & n14340 ;
  assign n14342 = ( ~n14339 & n14340 ) | ( ~n14339 & n14341 ) | ( n14340 & n14341 ) ;
  assign n14343 = ( ~n14275 & n14276 ) | ( ~n14275 & n14277 ) | ( n14276 & n14277 ) ;
  assign n14344 = n13749 | n14262 ;
  assign n14345 = n13748 & ~n14344 ;
  assign n14346 = n14263 | n14345 ;
  assign n14347 = n4781 & n12553 ;
  assign n14348 = n4776 & n12355 ;
  assign n14349 = n4778 & n12558 ;
  assign n14350 = n14348 | n14349 ;
  assign n14351 = n14347 | n14350 ;
  assign n14352 = n4784 | n14351 ;
  assign n14353 = ( n13097 & n14351 ) | ( n13097 & n14352 ) | ( n14351 & n14352 ) ;
  assign n14354 = x20 & n14353 ;
  assign n14355 = x20 & ~n14354 ;
  assign n14356 = ( n14353 & ~n14354 ) | ( n14353 & n14355 ) | ( ~n14354 & n14355 ) ;
  assign n14357 = ~n14346 & n14356 ;
  assign n14358 = ( ~n14260 & n14261 ) | ( ~n14260 & n14262 ) | ( n14261 & n14262 ) ;
  assign n14359 = n4484 & ~n12371 ;
  assign n14360 = n4479 & ~n12502 ;
  assign n14361 = n4481 & n12378 ;
  assign n14362 = n14360 | n14361 ;
  assign n14363 = n14359 | n14362 ;
  assign n14364 = n4487 | n14363 ;
  assign n14365 = ( ~n12848 & n14363 ) | ( ~n12848 & n14364 ) | ( n14363 & n14364 ) ;
  assign n14366 = ~x26 & n14365 ;
  assign n14367 = x26 | n14366 ;
  assign n14368 = ( ~n14365 & n14366 ) | ( ~n14365 & n14367 ) | ( n14366 & n14367 ) ;
  assign n14369 = n14225 | n14236 ;
  assign n14370 = ( ~n14235 & n14236 ) | ( ~n14235 & n14369 ) | ( n14236 & n14369 ) ;
  assign n14371 = n14368 & ~n14370 ;
  assign n14372 = n13768 & ~n14220 ;
  assign n14373 = n14221 | n14372 ;
  assign n14374 = n4048 & n12383 ;
  assign n14375 = n4043 & n12401 ;
  assign n14376 = n4045 & n12392 ;
  assign n14377 = n14375 | n14376 ;
  assign n14378 = n14374 | n14377 ;
  assign n14379 = n4051 | n14378 ;
  assign n14380 = ( n13141 & n14378 ) | ( n13141 & n14379 ) | ( n14378 & n14379 ) ;
  assign n14381 = x29 & n14380 ;
  assign n14382 = x29 & ~n14381 ;
  assign n14383 = ( n14380 & ~n14381 ) | ( n14380 & n14382 ) | ( ~n14381 & n14382 ) ;
  assign n14384 = ~n14373 & n14383 ;
  assign n14385 = n4479 & n12387 ;
  assign n14386 = n4481 & ~n12502 ;
  assign n14387 = n4484 & n12378 ;
  assign n14388 = n14386 | n14387 ;
  assign n14389 = n14385 | n14388 ;
  assign n14390 = n4487 | n14389 ;
  assign n14391 = ( ~n12816 & n14389 ) | ( ~n12816 & n14390 ) | ( n14389 & n14390 ) ;
  assign n14392 = ~x26 & n14391 ;
  assign n14393 = x26 | n14392 ;
  assign n14394 = ( ~n14391 & n14392 ) | ( ~n14391 & n14393 ) | ( n14392 & n14393 ) ;
  assign n14395 = n14373 | n14384 ;
  assign n14396 = ( ~n14383 & n14384 ) | ( ~n14383 & n14395 ) | ( n14384 & n14395 ) ;
  assign n14397 = n14394 & ~n14396 ;
  assign n14398 = n14384 | n14397 ;
  assign n14399 = ~n14368 & n14370 ;
  assign n14400 = n14371 | n14399 ;
  assign n14401 = n14398 & ~n14400 ;
  assign n14402 = n14371 | n14401 ;
  assign n14403 = n4551 & n12364 ;
  assign n14404 = n4546 & n12520 ;
  assign n14405 = n4548 & ~n12360 ;
  assign n14406 = n14404 | n14405 ;
  assign n14407 = n14403 | n14406 ;
  assign n14408 = n4554 | n14407 ;
  assign n14409 = ( ~n13113 & n14407 ) | ( ~n13113 & n14408 ) | ( n14407 & n14408 ) ;
  assign n14410 = ~x23 & n14409 ;
  assign n14411 = x23 | n14410 ;
  assign n14412 = ( ~n14409 & n14410 ) | ( ~n14409 & n14411 ) | ( n14410 & n14411 ) ;
  assign n14413 = ( n13751 & n14247 ) | ( n13751 & ~n14248 ) | ( n14247 & ~n14248 ) ;
  assign n14414 = ( n14237 & ~n14248 ) | ( n14237 & n14413 ) | ( ~n14248 & n14413 ) ;
  assign n14415 = ( n14402 & n14412 ) | ( n14402 & n14414 ) | ( n14412 & n14414 ) ;
  assign n14416 = n4781 & n12558 ;
  assign n14417 = n4776 & n12351 ;
  assign n14418 = n4778 & n12355 ;
  assign n14419 = n14417 | n14418 ;
  assign n14420 = n14416 | n14419 ;
  assign n14421 = n4784 | n14420 ;
  assign n14422 = ( n13330 & n14420 ) | ( n13330 & n14421 ) | ( n14420 & n14421 ) ;
  assign n14423 = x20 & n14422 ;
  assign n14424 = x20 & ~n14423 ;
  assign n14425 = ( n14422 & ~n14423 ) | ( n14422 & n14424 ) | ( ~n14423 & n14424 ) ;
  assign n14426 = ( n14358 & ~n14415 ) | ( n14358 & n14425 ) | ( ~n14415 & n14425 ) ;
  assign n14427 = ( ~n14358 & n14415 ) | ( ~n14358 & n14426 ) | ( n14415 & n14426 ) ;
  assign n14428 = n14346 | n14357 ;
  assign n14429 = ( ~n14356 & n14357 ) | ( ~n14356 & n14428 ) | ( n14357 & n14428 ) ;
  assign n14430 = n14427 & ~n14429 ;
  assign n14431 = n14357 | n14430 ;
  assign n14432 = n5083 & n12580 ;
  assign n14433 = n5069 & ~n12344 ;
  assign n14434 = n5070 & ~n12586 ;
  assign n14435 = n14433 | n14434 ;
  assign n14436 = n14432 | n14435 ;
  assign n14437 = n5074 | n14436 ;
  assign n14438 = ( n13432 & n14436 ) | ( n13432 & n14437 ) | ( n14436 & n14437 ) ;
  assign n14439 = x17 & n14438 ;
  assign n14440 = x17 & ~n14439 ;
  assign n14441 = ( n14438 & ~n14439 ) | ( n14438 & n14440 ) | ( ~n14439 & n14440 ) ;
  assign n14442 = ( n14343 & ~n14431 ) | ( n14343 & n14441 ) | ( ~n14431 & n14441 ) ;
  assign n14443 = ( ~n14343 & n14431 ) | ( ~n14343 & n14442 ) | ( n14431 & n14442 ) ;
  assign n14444 = ( ~n14331 & n14342 ) | ( ~n14331 & n14443 ) | ( n14342 & n14443 ) ;
  assign n14445 = n14330 & n14444 ;
  assign n14446 = n14444 & ~n14445 ;
  assign n14447 = ~n14290 & n14292 ;
  assign n14448 = n14293 | n14447 ;
  assign n14449 = n14330 & ~n14444 ;
  assign n14450 = ( n14446 & ~n14448 ) | ( n14446 & n14449 ) | ( ~n14448 & n14449 ) ;
  assign n14451 = n14445 | n14450 ;
  assign n14452 = n14296 & ~n14313 ;
  assign n14453 = ~n14312 & n14452 ;
  assign n14454 = n14312 | n14453 ;
  assign n14455 = ( ~n14452 & n14453 ) | ( ~n14452 & n14454 ) | ( n14453 & n14454 ) ;
  assign n14456 = n14451 & n14455 ;
  assign n14457 = n14129 & ~n14130 ;
  assign n14458 = n13916 & ~n14130 ;
  assign n14459 = n14457 | n14458 ;
  assign n14460 = n4048 & n12433 ;
  assign n14461 = n4043 & n12440 ;
  assign n14462 = n4045 & ~n12438 ;
  assign n14463 = n14461 | n14462 ;
  assign n14464 = n14460 | n14463 ;
  assign n14465 = n4051 | n14464 ;
  assign n14466 = ( ~n14167 & n14464 ) | ( ~n14167 & n14465 ) | ( n14464 & n14465 ) ;
  assign n14467 = ~x29 & n14466 ;
  assign n14468 = x29 | n14467 ;
  assign n14469 = ( ~n14466 & n14467 ) | ( ~n14466 & n14468 ) | ( n14467 & n14468 ) ;
  assign n14470 = n14459 & n14469 ;
  assign n14471 = n4048 & ~n12438 ;
  assign n14472 = n4043 & n12446 ;
  assign n14473 = n4045 & n12440 ;
  assign n14474 = n14472 | n14473 ;
  assign n14475 = n14471 | n14474 ;
  assign n14476 = ( n4051 & ~n14154 ) | ( n4051 & n14156 ) | ( ~n14154 & n14156 ) ;
  assign n14477 = n14475 | n14476 ;
  assign n14478 = x29 | n14477 ;
  assign n14479 = ~x29 & n14478 ;
  assign n14480 = ( ~n14477 & n14478 ) | ( ~n14477 & n14479 ) | ( n14478 & n14479 ) ;
  assign n14481 = ~n14128 & n14480 ;
  assign n14482 = n14480 & ~n14481 ;
  assign n14483 = n14128 | n14481 ;
  assign n14484 = ~n14482 & n14483 ;
  assign n14485 = n4048 & n12440 ;
  assign n14486 = n4043 & n12452 ;
  assign n14487 = n4045 & n12446 ;
  assign n14488 = n14486 | n14487 ;
  assign n14489 = n14485 | n14488 ;
  assign n14490 = n4051 | n14489 ;
  assign n14491 = ( n13822 & n14489 ) | ( n13822 & n14490 ) | ( n14489 & n14490 ) ;
  assign n14492 = x29 & n14491 ;
  assign n14493 = x29 & ~n14492 ;
  assign n14494 = ( n14491 & ~n14492 ) | ( n14491 & n14493 ) | ( ~n14492 & n14493 ) ;
  assign n14495 = ~n14091 & n14494 ;
  assign n14496 = n4048 & n12446 ;
  assign n14497 = n4043 & n12454 ;
  assign n14498 = n4045 & n12452 ;
  assign n14499 = n14497 | n14498 ;
  assign n14500 = n14496 | n14499 ;
  assign n14501 = n4051 | n14500 ;
  assign n14502 = ( n13862 & n14500 ) | ( n13862 & n14501 ) | ( n14500 & n14501 ) ;
  assign n14503 = ~x29 & n14502 ;
  assign n14504 = x29 & ~n14502 ;
  assign n14505 = n14503 | n14504 ;
  assign n14506 = ( n14014 & ~n14029 ) | ( n14014 & n14038 ) | ( ~n14029 & n14038 ) ;
  assign n14507 = ( ~n14014 & n14029 ) | ( ~n14014 & n14506 ) | ( n14029 & n14506 ) ;
  assign n14508 = ( ~n14038 & n14506 ) | ( ~n14038 & n14507 ) | ( n14506 & n14507 ) ;
  assign n14509 = n14505 & n14508 ;
  assign n14510 = n14505 | n14508 ;
  assign n14511 = ~n14509 & n14510 ;
  assign n14512 = n4048 & n12452 ;
  assign n14513 = n4043 & ~n12456 ;
  assign n14514 = n4045 & n12454 ;
  assign n14515 = n14513 | n14514 ;
  assign n14516 = n14512 | n14515 ;
  assign n14517 = n4051 | n14516 ;
  assign n14518 = ( ~n13922 & n14516 ) | ( ~n13922 & n14517 ) | ( n14516 & n14517 ) ;
  assign n14519 = ~x29 & n14518 ;
  assign n14520 = x29 & ~n14518 ;
  assign n14521 = n14519 | n14520 ;
  assign n14522 = n14010 & ~n14013 ;
  assign n14523 = n14012 | n14013 ;
  assign n14524 = ~n14522 & n14523 ;
  assign n14525 = n14521 & ~n14524 ;
  assign n14526 = ~n14521 & n14524 ;
  assign n14527 = n14525 | n14526 ;
  assign n14528 = n4048 & n12454 ;
  assign n14529 = n4043 & n12459 ;
  assign n14530 = n4045 & ~n12456 ;
  assign n14531 = n14529 | n14530 ;
  assign n14532 = n14528 | n14531 ;
  assign n14533 = n4051 | n14532 ;
  assign n14534 = ( n14041 & n14532 ) | ( n14041 & n14533 ) | ( n14532 & n14533 ) ;
  assign n14535 = ~x29 & n14534 ;
  assign n14536 = x29 & ~n14534 ;
  assign n14537 = n14535 | n14536 ;
  assign n14538 = n13992 | n13999 ;
  assign n14539 = ( ~n13999 & n14000 ) | ( ~n13999 & n14538 ) | ( n14000 & n14538 ) ;
  assign n14540 = n14537 & ~n14539 ;
  assign n14541 = ~n14537 & n14539 ;
  assign n14542 = n14540 | n14541 ;
  assign n14543 = n3635 & ~n12468 ;
  assign n14544 = n4048 & ~n12456 ;
  assign n14545 = n4043 & ~n12466 ;
  assign n14546 = n4045 & n12459 ;
  assign n14547 = n14545 | n14546 ;
  assign n14548 = n14544 | n14547 ;
  assign n14549 = n4051 | n14548 ;
  assign n14550 = ( n14031 & n14548 ) | ( n14031 & n14549 ) | ( n14548 & n14549 ) ;
  assign n14551 = x29 & n14550 ;
  assign n14552 = x29 & ~n14551 ;
  assign n14553 = ( n14550 & ~n14551 ) | ( n14550 & n14552 ) | ( ~n14551 & n14552 ) ;
  assign n14554 = x29 & ~n4041 ;
  assign n14555 = ( x29 & n12468 ) | ( x29 & n14554 ) | ( n12468 & n14554 ) ;
  assign n14556 = n4051 & n13994 ;
  assign n14557 = n4045 & ~n12468 ;
  assign n14558 = n4048 & ~n12466 ;
  assign n14559 = n14557 | n14558 ;
  assign n14560 = n14556 | n14559 ;
  assign n14561 = x29 | n14560 ;
  assign n14562 = ~x29 & n14561 ;
  assign n14563 = ( ~n14560 & n14561 ) | ( ~n14560 & n14562 ) | ( n14561 & n14562 ) ;
  assign n14564 = n14555 & n14563 ;
  assign n14565 = n4048 & n12459 ;
  assign n14566 = n4043 & ~n12468 ;
  assign n14567 = n4045 & ~n12466 ;
  assign n14568 = n14566 | n14567 ;
  assign n14569 = n14565 | n14568 ;
  assign n14570 = n4051 & n14003 ;
  assign n14571 = n14569 | n14570 ;
  assign n14572 = ~x29 & n14571 ;
  assign n14573 = x29 | n14572 ;
  assign n14574 = ( ~n14571 & n14572 ) | ( ~n14571 & n14573 ) | ( n14572 & n14573 ) ;
  assign n14575 = n14564 & n14574 ;
  assign n14576 = ( n14543 & n14553 ) | ( n14543 & n14575 ) | ( n14553 & n14575 ) ;
  assign n14577 = ~n14542 & n14576 ;
  assign n14578 = n14540 | n14577 ;
  assign n14579 = ~n14527 & n14578 ;
  assign n14580 = n14525 | n14579 ;
  assign n14581 = n14511 & n14580 ;
  assign n14582 = n14509 | n14581 ;
  assign n14583 = n14494 & ~n14495 ;
  assign n14584 = n14091 | n14495 ;
  assign n14585 = ~n14583 & n14584 ;
  assign n14586 = n14582 & ~n14585 ;
  assign n14587 = n14495 | n14586 ;
  assign n14588 = ~n14484 & n14587 ;
  assign n14589 = n14459 | n14469 ;
  assign n14590 = ~n14470 & n14589 ;
  assign n14591 = ( n14481 & n14588 ) | ( n14481 & n14590 ) | ( n14588 & n14590 ) ;
  assign n14592 = n13855 | n14131 ;
  assign n14593 = ~n14132 & n14592 ;
  assign n14594 = n4048 & ~n12423 ;
  assign n14595 = n4043 & ~n12438 ;
  assign n14596 = n4045 & n12433 ;
  assign n14597 = n14595 | n14596 ;
  assign n14598 = n14594 | n14597 ;
  assign n14599 = n4051 | n14598 ;
  assign n14600 = ( ~n13786 & n14598 ) | ( ~n13786 & n14599 ) | ( n14598 & n14599 ) ;
  assign n14601 = ~x29 & n14600 ;
  assign n14602 = x29 | n14601 ;
  assign n14603 = ( ~n14600 & n14601 ) | ( ~n14600 & n14602 ) | ( n14601 & n14602 ) ;
  assign n14604 = n14593 & n14603 ;
  assign n14605 = n14593 | n14603 ;
  assign n14606 = ~n14604 & n14605 ;
  assign n14607 = ( n14470 & n14591 ) | ( n14470 & n14606 ) | ( n14591 & n14606 ) ;
  assign n14608 = ~n14148 & n14158 ;
  assign n14609 = n14148 & n14158 ;
  assign n14610 = ( n14148 & n14608 ) | ( n14148 & ~n14609 ) | ( n14608 & ~n14609 ) ;
  assign n14611 = n14133 & ~n14610 ;
  assign n14612 = ~n14133 & n14610 ;
  assign n14613 = n4048 & n12419 ;
  assign n14614 = n4043 & n12433 ;
  assign n14615 = n4045 & ~n12423 ;
  assign n14616 = n14614 | n14615 ;
  assign n14617 = n14613 | n14616 ;
  assign n14618 = n4051 | n14617 ;
  assign n14619 = ( ~n13282 & n14617 ) | ( ~n13282 & n14618 ) | ( n14617 & n14618 ) ;
  assign n14620 = ~x29 & n14619 ;
  assign n14621 = x29 | n14620 ;
  assign n14622 = ( ~n14619 & n14620 ) | ( ~n14619 & n14621 ) | ( n14620 & n14621 ) ;
  assign n14623 = n14612 | n14622 ;
  assign n14624 = n14611 | n14623 ;
  assign n14625 = ( n14611 & n14612 ) | ( n14611 & n14622 ) | ( n14612 & n14622 ) ;
  assign n14626 = n14624 & ~n14625 ;
  assign n14627 = n14604 & n14626 ;
  assign n14628 = ( n14607 & n14626 ) | ( n14607 & n14627 ) | ( n14626 & n14627 ) ;
  assign n14629 = ~n14159 & n14190 ;
  assign n14630 = n4048 & n12411 ;
  assign n14631 = n4043 & ~n12423 ;
  assign n14632 = n4045 & n12419 ;
  assign n14633 = n14631 | n14632 ;
  assign n14634 = n14630 | n14633 ;
  assign n14635 = n4051 | n14634 ;
  assign n14636 = ( n13776 & n14634 ) | ( n13776 & n14635 ) | ( n14634 & n14635 ) ;
  assign n14637 = x29 & n14636 ;
  assign n14638 = x29 & ~n14637 ;
  assign n14639 = ( n14636 & ~n14637 ) | ( n14636 & n14638 ) | ( ~n14637 & n14638 ) ;
  assign n14640 = n14629 | n14639 ;
  assign n14641 = n14191 | n14640 ;
  assign n14642 = ( n14191 & n14629 ) | ( n14191 & n14639 ) | ( n14629 & n14639 ) ;
  assign n14643 = n14641 & ~n14642 ;
  assign n14644 = n14625 | n14643 ;
  assign n14645 = n14628 | n14644 ;
  assign n14646 = ( n14625 & n14628 ) | ( n14625 & n14643 ) | ( n14628 & n14643 ) ;
  assign n14647 = n14645 & ~n14646 ;
  assign n14648 = n4484 & n12392 ;
  assign n14649 = n4479 & n12415 ;
  assign n14650 = n4481 & n12401 ;
  assign n14651 = n14649 | n14650 ;
  assign n14652 = n14648 | n14651 ;
  assign n14653 = n4487 | n14652 ;
  assign n14654 = ( n13034 & n14652 ) | ( n13034 & n14653 ) | ( n14652 & n14653 ) ;
  assign n14655 = x26 & n14654 ;
  assign n14656 = x26 & ~n14655 ;
  assign n14657 = ( n14654 & ~n14655 ) | ( n14654 & n14656 ) | ( ~n14655 & n14656 ) ;
  assign n14658 = ~n14647 & n14657 ;
  assign n14659 = n14647 & ~n14657 ;
  assign n14660 = n14658 | n14659 ;
  assign n14661 = n14604 | n14626 ;
  assign n14662 = n14607 | n14661 ;
  assign n14663 = ~n14628 & n14662 ;
  assign n14664 = n4484 & n12401 ;
  assign n14665 = n4479 & n12411 ;
  assign n14666 = n4481 & n12415 ;
  assign n14667 = n14665 | n14666 ;
  assign n14668 = n14664 | n14667 ;
  assign n14669 = n4487 & ~n13163 ;
  assign n14670 = ~n13161 & n14669 ;
  assign n14671 = ( n4487 & n14668 ) | ( n4487 & ~n14670 ) | ( n14668 & ~n14670 ) ;
  assign n14672 = ~x26 & n14671 ;
  assign n14673 = x26 | n14672 ;
  assign n14674 = ( ~n14671 & n14672 ) | ( ~n14671 & n14673 ) | ( n14672 & n14673 ) ;
  assign n14675 = n14470 | n14606 ;
  assign n14676 = n14591 | n14675 ;
  assign n14677 = ~n14607 & n14676 ;
  assign n14678 = n4484 & n12415 ;
  assign n14679 = n4479 & n12419 ;
  assign n14680 = n4481 & n12411 ;
  assign n14681 = n14679 | n14680 ;
  assign n14682 = n14678 | n14681 ;
  assign n14683 = n4487 & ~n13761 ;
  assign n14684 = ~n13762 & n14683 ;
  assign n14685 = ( n4487 & n14682 ) | ( n4487 & ~n14684 ) | ( n14682 & ~n14684 ) ;
  assign n14686 = ~x26 & n14685 ;
  assign n14687 = x26 | n14686 ;
  assign n14688 = ( ~n14685 & n14686 ) | ( ~n14685 & n14687 ) | ( n14686 & n14687 ) ;
  assign n14689 = n14481 | n14590 ;
  assign n14690 = n14588 | n14689 ;
  assign n14691 = ~n14591 & n14690 ;
  assign n14692 = n4484 & n12411 ;
  assign n14693 = n4479 & ~n12423 ;
  assign n14694 = n4481 & n12419 ;
  assign n14695 = n14693 | n14694 ;
  assign n14696 = n14692 | n14695 ;
  assign n14697 = n4487 | n14696 ;
  assign n14698 = ( n13776 & n14696 ) | ( n13776 & n14697 ) | ( n14696 & n14697 ) ;
  assign n14699 = x26 & n14698 ;
  assign n14700 = x26 & ~n14699 ;
  assign n14701 = ( n14698 & ~n14699 ) | ( n14698 & n14700 ) | ( ~n14699 & n14700 ) ;
  assign n14702 = ~n14582 & n14585 ;
  assign n14703 = n14586 | n14702 ;
  assign n14704 = n4479 & ~n12438 ;
  assign n14705 = n4481 & n12433 ;
  assign n14706 = n4484 & ~n12423 ;
  assign n14707 = n14705 | n14706 ;
  assign n14708 = n14704 | n14707 ;
  assign n14709 = n4487 | n14708 ;
  assign n14710 = ( ~n13786 & n14708 ) | ( ~n13786 & n14709 ) | ( n14708 & n14709 ) ;
  assign n14711 = ~x26 & n14710 ;
  assign n14712 = x26 | n14711 ;
  assign n14713 = ( ~n14710 & n14711 ) | ( ~n14710 & n14712 ) | ( n14711 & n14712 ) ;
  assign n14714 = ~n14703 & n14713 ;
  assign n14715 = n14527 & ~n14578 ;
  assign n14716 = n14579 | n14715 ;
  assign n14717 = n4484 & ~n12438 ;
  assign n14718 = n4481 & n12440 ;
  assign n14719 = n4479 & n12446 ;
  assign n14720 = n14718 | n14719 ;
  assign n14721 = n14717 | n14720 ;
  assign n14722 = n4487 & ~n14156 ;
  assign n14723 = n14154 & n14722 ;
  assign n14724 = ( n4487 & n14721 ) | ( n4487 & ~n14723 ) | ( n14721 & ~n14723 ) ;
  assign n14725 = x26 & n14724 ;
  assign n14726 = x26 & ~n14725 ;
  assign n14727 = ( n14724 & ~n14725 ) | ( n14724 & n14726 ) | ( ~n14725 & n14726 ) ;
  assign n14728 = ~n14716 & n14727 ;
  assign n14729 = n14542 | n14577 ;
  assign n14730 = n14542 & n14576 ;
  assign n14731 = n14729 & ~n14730 ;
  assign n14732 = n4479 & n12452 ;
  assign n14733 = n4481 & n12446 ;
  assign n14734 = n4484 & n12440 ;
  assign n14735 = n14733 | n14734 ;
  assign n14736 = n14732 | n14735 ;
  assign n14737 = n4487 | n14736 ;
  assign n14738 = ( n13822 & n14736 ) | ( n13822 & n14737 ) | ( n14736 & n14737 ) ;
  assign n14739 = x26 & n14738 ;
  assign n14740 = x26 & ~n14739 ;
  assign n14741 = ( n14738 & ~n14739 ) | ( n14738 & n14740 ) | ( ~n14739 & n14740 ) ;
  assign n14742 = ~n14731 & n14741 ;
  assign n14743 = n4481 & n12452 ;
  assign n14744 = n4479 & n12454 ;
  assign n14745 = n4484 | n14744 ;
  assign n14746 = ( n12446 & n14744 ) | ( n12446 & n14745 ) | ( n14744 & n14745 ) ;
  assign n14747 = n14743 | n14746 ;
  assign n14748 = n4487 | n14747 ;
  assign n14749 = ( n13862 & n14747 ) | ( n13862 & n14748 ) | ( n14747 & n14748 ) ;
  assign n14750 = ~x26 & n14749 ;
  assign n14751 = x26 & ~n14749 ;
  assign n14752 = n14750 | n14751 ;
  assign n14753 = ( n14553 & n14575 ) | ( n14553 & ~n14576 ) | ( n14575 & ~n14576 ) ;
  assign n14754 = ( n14543 & ~n14576 ) | ( n14543 & n14753 ) | ( ~n14576 & n14753 ) ;
  assign n14755 = n14752 & n14754 ;
  assign n14756 = n14752 | n14754 ;
  assign n14757 = ~n14755 & n14756 ;
  assign n14758 = n4484 & n12452 ;
  assign n14759 = n4479 & ~n12456 ;
  assign n14760 = n4481 & n12454 ;
  assign n14761 = n14759 | n14760 ;
  assign n14762 = n14758 | n14761 ;
  assign n14763 = n4487 | n14762 ;
  assign n14764 = ( ~n13922 & n14762 ) | ( ~n13922 & n14763 ) | ( n14762 & n14763 ) ;
  assign n14765 = ~x26 & n14764 ;
  assign n14766 = x26 & ~n14764 ;
  assign n14767 = n14765 | n14766 ;
  assign n14768 = n14564 | n14574 ;
  assign n14769 = ~n14575 & n14768 ;
  assign n14770 = n14767 & n14769 ;
  assign n14771 = n14555 | n14563 ;
  assign n14772 = ~n14564 & n14771 ;
  assign n14773 = n4484 & n12454 ;
  assign n14774 = n4479 & n12459 ;
  assign n14775 = n4481 & ~n12456 ;
  assign n14776 = n14774 | n14775 ;
  assign n14777 = n14773 | n14776 ;
  assign n14778 = n4487 | n14777 ;
  assign n14779 = ( n14041 & n14777 ) | ( n14041 & n14778 ) | ( n14777 & n14778 ) ;
  assign n14780 = x26 & n14779 ;
  assign n14781 = x26 & ~n14780 ;
  assign n14782 = ( n14779 & ~n14780 ) | ( n14779 & n14781 ) | ( ~n14780 & n14781 ) ;
  assign n14783 = n14772 & n14782 ;
  assign n14784 = n14772 | n14782 ;
  assign n14785 = ~n14783 & n14784 ;
  assign n14786 = x26 & ~n4474 ;
  assign n14787 = ( x26 & n12468 ) | ( x26 & n14786 ) | ( n12468 & n14786 ) ;
  assign n14788 = n4487 & n13994 ;
  assign n14789 = n4484 & ~n12466 ;
  assign n14790 = n4481 & ~n12468 ;
  assign n14791 = n14789 | n14790 ;
  assign n14792 = n14788 | n14791 ;
  assign n14793 = x26 | n14792 ;
  assign n14794 = ~x26 & n14793 ;
  assign n14795 = ( ~n14792 & n14793 ) | ( ~n14792 & n14794 ) | ( n14793 & n14794 ) ;
  assign n14796 = n14787 & n14795 ;
  assign n14797 = n4041 & ~n12468 ;
  assign n14798 = n4479 & ~n12468 ;
  assign n14799 = n4484 & n12459 ;
  assign n14800 = n4481 & ~n12466 ;
  assign n14801 = n14799 | n14800 ;
  assign n14802 = n14798 | n14801 ;
  assign n14803 = n4487 & n14003 ;
  assign n14804 = n14802 | n14803 ;
  assign n14805 = ~x26 & n14804 ;
  assign n14806 = x26 | n14805 ;
  assign n14807 = ( ~n14804 & n14805 ) | ( ~n14804 & n14806 ) | ( n14805 & n14806 ) ;
  assign n14808 = n14797 & n14807 ;
  assign n14809 = n14796 & n14808 ;
  assign n14810 = n14796 & n14807 ;
  assign n14811 = n14797 | n14810 ;
  assign n14812 = ~n14809 & n14811 ;
  assign n14813 = n4484 & ~n12456 ;
  assign n14814 = n4479 & ~n12466 ;
  assign n14815 = n4481 & n12459 ;
  assign n14816 = n14814 | n14815 ;
  assign n14817 = n14813 | n14816 ;
  assign n14818 = ( n4487 & n14031 ) | ( n4487 & n14817 ) | ( n14031 & n14817 ) ;
  assign n14819 = ( x26 & ~n14817 ) | ( x26 & n14818 ) | ( ~n14817 & n14818 ) ;
  assign n14820 = ~n14818 & n14819 ;
  assign n14821 = n14817 | n14819 ;
  assign n14822 = ( ~x26 & n14820 ) | ( ~x26 & n14821 ) | ( n14820 & n14821 ) ;
  assign n14823 = n14812 & n14822 ;
  assign n14824 = n14809 | n14823 ;
  assign n14825 = n14785 & n14824 ;
  assign n14826 = n14783 | n14825 ;
  assign n14827 = n14767 | n14769 ;
  assign n14828 = ~n14770 & n14827 ;
  assign n14829 = n14826 & n14828 ;
  assign n14830 = n14770 | n14829 ;
  assign n14831 = n14757 & n14830 ;
  assign n14832 = n14755 | n14831 ;
  assign n14833 = n14731 & ~n14741 ;
  assign n14834 = n14742 | n14833 ;
  assign n14835 = n14832 & ~n14834 ;
  assign n14836 = n14742 | n14835 ;
  assign n14837 = n14716 | n14728 ;
  assign n14838 = ( ~n14727 & n14728 ) | ( ~n14727 & n14837 ) | ( n14728 & n14837 ) ;
  assign n14839 = n14836 & ~n14838 ;
  assign n14840 = n14728 | n14839 ;
  assign n14841 = n14511 | n14580 ;
  assign n14842 = ~n14581 & n14841 ;
  assign n14843 = n4479 & n12440 ;
  assign n14844 = n4484 & n12433 ;
  assign n14845 = n4481 & ~n12438 ;
  assign n14846 = n14844 | n14845 ;
  assign n14847 = n14843 | n14846 ;
  assign n14848 = n4487 | n14847 ;
  assign n14849 = ( ~n14167 & n14847 ) | ( ~n14167 & n14848 ) | ( n14847 & n14848 ) ;
  assign n14850 = ~x26 & n14849 ;
  assign n14851 = x26 | n14850 ;
  assign n14852 = ( ~n14849 & n14850 ) | ( ~n14849 & n14851 ) | ( n14850 & n14851 ) ;
  assign n14853 = ( n14840 & n14842 ) | ( n14840 & n14852 ) | ( n14842 & n14852 ) ;
  assign n14854 = n14703 | n14714 ;
  assign n14855 = ( ~n14713 & n14714 ) | ( ~n14713 & n14854 ) | ( n14714 & n14854 ) ;
  assign n14856 = n14853 & ~n14855 ;
  assign n14857 = n14714 | n14856 ;
  assign n14858 = n4484 & n12419 ;
  assign n14859 = n4479 & n12433 ;
  assign n14860 = n4481 & ~n12423 ;
  assign n14861 = n14859 | n14860 ;
  assign n14862 = n14858 | n14861 ;
  assign n14863 = n4487 | n14862 ;
  assign n14864 = ( ~n13282 & n14862 ) | ( ~n13282 & n14863 ) | ( n14862 & n14863 ) ;
  assign n14865 = ~x26 & n14864 ;
  assign n14866 = x26 | n14865 ;
  assign n14867 = ( ~n14864 & n14865 ) | ( ~n14864 & n14866 ) | ( n14865 & n14866 ) ;
  assign n14868 = n14484 & ~n14587 ;
  assign n14869 = n14588 | n14868 ;
  assign n14870 = ( n14857 & n14867 ) | ( n14857 & ~n14869 ) | ( n14867 & ~n14869 ) ;
  assign n14871 = ( n14691 & n14701 ) | ( n14691 & n14870 ) | ( n14701 & n14870 ) ;
  assign n14872 = ( n14677 & n14688 ) | ( n14677 & n14871 ) | ( n14688 & n14871 ) ;
  assign n14873 = ( n14663 & n14674 ) | ( n14663 & n14872 ) | ( n14674 & n14872 ) ;
  assign n14874 = n14660 & ~n14873 ;
  assign n14875 = ~n14660 & n14873 ;
  assign n14876 = n14874 | n14875 ;
  assign n14877 = n4551 & ~n12502 ;
  assign n14878 = n4546 & n12383 ;
  assign n14879 = n4548 & n12387 ;
  assign n14880 = n14878 | n14879 ;
  assign n14881 = n14877 | n14880 ;
  assign n14882 = n4554 | n14881 ;
  assign n14883 = ( ~n12756 & n14881 ) | ( ~n12756 & n14882 ) | ( n14881 & n14882 ) ;
  assign n14884 = ~x23 & n14883 ;
  assign n14885 = x23 | n14884 ;
  assign n14886 = ( ~n14883 & n14884 ) | ( ~n14883 & n14885 ) | ( n14884 & n14885 ) ;
  assign n14887 = n14876 & n14886 ;
  assign n14888 = ~n14663 & n14674 ;
  assign n14889 = n14663 & ~n14674 ;
  assign n14890 = n14888 | n14889 ;
  assign n14891 = ~n14872 & n14890 ;
  assign n14892 = n14872 & ~n14890 ;
  assign n14893 = n14891 | n14892 ;
  assign n14894 = n4551 & n12387 ;
  assign n14895 = n4546 & n12392 ;
  assign n14896 = n4548 & n12383 ;
  assign n14897 = n14895 | n14896 ;
  assign n14898 = n14894 | n14897 ;
  assign n14899 = n4554 | n14898 ;
  assign n14900 = ( n12948 & n14898 ) | ( n12948 & n14899 ) | ( n14898 & n14899 ) ;
  assign n14901 = x23 & n14900 ;
  assign n14902 = x23 & ~n14901 ;
  assign n14903 = ( n14900 & ~n14901 ) | ( n14900 & n14902 ) | ( ~n14901 & n14902 ) ;
  assign n14904 = n14893 & n14903 ;
  assign n14905 = n4551 & n12383 ;
  assign n14906 = n4546 & n12401 ;
  assign n14907 = n4548 & n12392 ;
  assign n14908 = n14906 | n14907 ;
  assign n14909 = n14905 | n14908 ;
  assign n14910 = n4554 | n14909 ;
  assign n14911 = ( n13141 & n14909 ) | ( n13141 & n14910 ) | ( n14909 & n14910 ) ;
  assign n14912 = x23 & n14911 ;
  assign n14913 = x23 & ~n14912 ;
  assign n14914 = ( n14911 & ~n14912 ) | ( n14911 & n14913 ) | ( ~n14912 & n14913 ) ;
  assign n14915 = ~n14677 & n14688 ;
  assign n14916 = n14677 & ~n14688 ;
  assign n14917 = n14915 | n14916 ;
  assign n14918 = n14871 & n14917 ;
  assign n14919 = n14917 & ~n14918 ;
  assign n14920 = ( n14871 & ~n14918 ) | ( n14871 & n14919 ) | ( ~n14918 & n14919 ) ;
  assign n14921 = n14914 & n14920 ;
  assign n14922 = n4551 & n12392 ;
  assign n14923 = n4546 & n12415 ;
  assign n14924 = n4548 & n12401 ;
  assign n14925 = n14923 | n14924 ;
  assign n14926 = n14922 | n14925 ;
  assign n14927 = n4554 | n14926 ;
  assign n14928 = ( n13034 & n14926 ) | ( n13034 & n14927 ) | ( n14926 & n14927 ) ;
  assign n14929 = x23 & n14928 ;
  assign n14930 = x23 & ~n14929 ;
  assign n14931 = ( n14928 & ~n14929 ) | ( n14928 & n14930 ) | ( ~n14929 & n14930 ) ;
  assign n14932 = ( n14691 & n14870 ) | ( n14691 & ~n14871 ) | ( n14870 & ~n14871 ) ;
  assign n14933 = ( n14701 & ~n14871 ) | ( n14701 & n14932 ) | ( ~n14871 & n14932 ) ;
  assign n14934 = n14931 & n14933 ;
  assign n14935 = ( ~n14857 & n14869 ) | ( ~n14857 & n14870 ) | ( n14869 & n14870 ) ;
  assign n14936 = ( ~n14867 & n14870 ) | ( ~n14867 & n14935 ) | ( n14870 & n14935 ) ;
  assign n14937 = n4551 & n12401 ;
  assign n14938 = n4546 & n12411 ;
  assign n14939 = n4548 & n12415 ;
  assign n14940 = n14938 | n14939 ;
  assign n14941 = n14937 | n14940 ;
  assign n14942 = n4554 & n13163 ;
  assign n14943 = ( n4554 & n13161 ) | ( n4554 & n14942 ) | ( n13161 & n14942 ) ;
  assign n14944 = n14941 | n14943 ;
  assign n14945 = x23 | n14944 ;
  assign n14946 = ~x23 & n14945 ;
  assign n14947 = ( ~n14944 & n14945 ) | ( ~n14944 & n14946 ) | ( n14945 & n14946 ) ;
  assign n14948 = ~n14936 & n14947 ;
  assign n14949 = n14853 & ~n14856 ;
  assign n14950 = n14855 | n14856 ;
  assign n14951 = ~n14949 & n14950 ;
  assign n14952 = n4551 & n12415 ;
  assign n14953 = n4546 & n12419 ;
  assign n14954 = n4548 & n12411 ;
  assign n14955 = n14953 | n14954 ;
  assign n14956 = n14952 | n14955 ;
  assign n14957 = ( n4554 & n13761 ) | ( n4554 & n13762 ) | ( n13761 & n13762 ) ;
  assign n14958 = n14956 | n14957 ;
  assign n14959 = x23 | n14958 ;
  assign n14960 = ~x23 & n14959 ;
  assign n14961 = ( ~n14958 & n14959 ) | ( ~n14958 & n14960 ) | ( n14959 & n14960 ) ;
  assign n14962 = ~n14951 & n14961 ;
  assign n14963 = n4551 & n12411 ;
  assign n14964 = n4546 & ~n12423 ;
  assign n14965 = n4548 & n12419 ;
  assign n14966 = n14964 | n14965 ;
  assign n14967 = n14963 | n14966 ;
  assign n14968 = n4554 | n14967 ;
  assign n14969 = ( n13776 & n14967 ) | ( n13776 & n14968 ) | ( n14967 & n14968 ) ;
  assign n14970 = x23 & n14969 ;
  assign n14971 = x23 & ~n14970 ;
  assign n14972 = ( n14969 & ~n14970 ) | ( n14969 & n14971 ) | ( ~n14970 & n14971 ) ;
  assign n14973 = ( n14840 & ~n14842 ) | ( n14840 & n14852 ) | ( ~n14842 & n14852 ) ;
  assign n14974 = ( ~n14840 & n14842 ) | ( ~n14840 & n14973 ) | ( n14842 & n14973 ) ;
  assign n14975 = ( ~n14852 & n14973 ) | ( ~n14852 & n14974 ) | ( n14973 & n14974 ) ;
  assign n14976 = n14972 & n14975 ;
  assign n14977 = n14972 | n14975 ;
  assign n14978 = ~n14976 & n14977 ;
  assign n14979 = n14836 & ~n14839 ;
  assign n14980 = n14838 | n14839 ;
  assign n14981 = ~n14979 & n14980 ;
  assign n14982 = n4551 & n12419 ;
  assign n14983 = n4546 & n12433 ;
  assign n14984 = n4548 & ~n12423 ;
  assign n14985 = n14983 | n14984 ;
  assign n14986 = n14982 | n14985 ;
  assign n14987 = n4554 | n14986 ;
  assign n14988 = ( ~n13282 & n14986 ) | ( ~n13282 & n14987 ) | ( n14986 & n14987 ) ;
  assign n14989 = ~x23 & n14988 ;
  assign n14990 = x23 | n14989 ;
  assign n14991 = ( ~n14988 & n14989 ) | ( ~n14988 & n14990 ) | ( n14989 & n14990 ) ;
  assign n14992 = ~n14981 & n14991 ;
  assign n14993 = n14832 & ~n14835 ;
  assign n14994 = n14834 | n14835 ;
  assign n14995 = ~n14993 & n14994 ;
  assign n14996 = n4551 & ~n12423 ;
  assign n14997 = n4546 & ~n12438 ;
  assign n14998 = n4548 & n12433 ;
  assign n14999 = n14997 | n14998 ;
  assign n15000 = n14996 | n14999 ;
  assign n15001 = n4554 | n15000 ;
  assign n15002 = ( ~n13786 & n15000 ) | ( ~n13786 & n15001 ) | ( n15000 & n15001 ) ;
  assign n15003 = ~x23 & n15002 ;
  assign n15004 = x23 | n15003 ;
  assign n15005 = ( ~n15002 & n15003 ) | ( ~n15002 & n15004 ) | ( n15003 & n15004 ) ;
  assign n15006 = ~n14995 & n15005 ;
  assign n15007 = n14995 | n15006 ;
  assign n15008 = n14995 & n15005 ;
  assign n15009 = n14757 | n14830 ;
  assign n15010 = ~n14831 & n15009 ;
  assign n15011 = n4551 & n12433 ;
  assign n15012 = n4546 & n12440 ;
  assign n15013 = n4548 & ~n12438 ;
  assign n15014 = n15012 | n15013 ;
  assign n15015 = n15011 | n15014 ;
  assign n15016 = n4554 | n15015 ;
  assign n15017 = ( ~n14167 & n15015 ) | ( ~n14167 & n15016 ) | ( n15015 & n15016 ) ;
  assign n15018 = ~x23 & n15017 ;
  assign n15019 = x23 | n15018 ;
  assign n15020 = ( ~n15017 & n15018 ) | ( ~n15017 & n15019 ) | ( n15018 & n15019 ) ;
  assign n15021 = n15010 & n15020 ;
  assign n15022 = n15010 | n15020 ;
  assign n15023 = ~n15021 & n15022 ;
  assign n15024 = n14826 | n14828 ;
  assign n15025 = ~n14829 & n15024 ;
  assign n15026 = n4551 & ~n12438 ;
  assign n15027 = n4546 & n12446 ;
  assign n15028 = n4548 & n12440 ;
  assign n15029 = n15027 | n15028 ;
  assign n15030 = n15026 | n15029 ;
  assign n15031 = n4554 & n14154 ;
  assign n15032 = ~n14156 & n15031 ;
  assign n15033 = ( n4554 & n15030 ) | ( n4554 & ~n15032 ) | ( n15030 & ~n15032 ) ;
  assign n15034 = x23 & n15033 ;
  assign n15035 = x23 & ~n15034 ;
  assign n15036 = ( n15033 & ~n15034 ) | ( n15033 & n15035 ) | ( ~n15034 & n15035 ) ;
  assign n15037 = n14785 | n14824 ;
  assign n15038 = ~n14825 & n15037 ;
  assign n15039 = n4551 & n12440 ;
  assign n15040 = n4546 & n12452 ;
  assign n15041 = n4548 & n12446 ;
  assign n15042 = n15040 | n15041 ;
  assign n15043 = n15039 | n15042 ;
  assign n15044 = n4554 | n15043 ;
  assign n15045 = ( n13822 & n15043 ) | ( n13822 & n15044 ) | ( n15043 & n15044 ) ;
  assign n15046 = x23 & n15045 ;
  assign n15047 = x23 & ~n15046 ;
  assign n15048 = ( n15045 & ~n15046 ) | ( n15045 & n15047 ) | ( ~n15046 & n15047 ) ;
  assign n15049 = n15038 & n15048 ;
  assign n15050 = n4551 & n12446 ;
  assign n15051 = n4546 & n12454 ;
  assign n15052 = n4548 & n12452 ;
  assign n15053 = n15051 | n15052 ;
  assign n15054 = n15050 | n15053 ;
  assign n15055 = n4554 | n15054 ;
  assign n15056 = ( n13862 & n15054 ) | ( n13862 & n15055 ) | ( n15054 & n15055 ) ;
  assign n15057 = x23 & n15056 ;
  assign n15058 = x23 & ~n15057 ;
  assign n15059 = ( n15056 & ~n15057 ) | ( n15056 & n15058 ) | ( ~n15057 & n15058 ) ;
  assign n15060 = n14812 & ~n14823 ;
  assign n15061 = ( n14822 & ~n14823 ) | ( n14822 & n15060 ) | ( ~n14823 & n15060 ) ;
  assign n15062 = n15059 & n15061 ;
  assign n15063 = n15059 | n15061 ;
  assign n15064 = ~n15062 & n15063 ;
  assign n15065 = n4551 & n12452 ;
  assign n15066 = n4546 & ~n12456 ;
  assign n15067 = n4548 & n12454 ;
  assign n15068 = n15066 | n15067 ;
  assign n15069 = n15065 | n15068 ;
  assign n15070 = n4554 | n15069 ;
  assign n15071 = ( ~n13922 & n15069 ) | ( ~n13922 & n15070 ) | ( n15069 & n15070 ) ;
  assign n15072 = ~x23 & n15071 ;
  assign n15073 = x23 & ~n15071 ;
  assign n15074 = n15072 | n15073 ;
  assign n15075 = n14796 | n14807 ;
  assign n15076 = ~n14810 & n15075 ;
  assign n15077 = n15074 & n15076 ;
  assign n15078 = n14787 | n14795 ;
  assign n15079 = ~n14796 & n15078 ;
  assign n15080 = n4551 & n12454 ;
  assign n15081 = n4546 & n12459 ;
  assign n15082 = n4548 & ~n12456 ;
  assign n15083 = n15081 | n15082 ;
  assign n15084 = n15080 | n15083 ;
  assign n15085 = n4554 | n15084 ;
  assign n15086 = ( n14041 & n15084 ) | ( n14041 & n15085 ) | ( n15084 & n15085 ) ;
  assign n15087 = x23 & n15086 ;
  assign n15088 = x23 & ~n15087 ;
  assign n15089 = ( n15086 & ~n15087 ) | ( n15086 & n15088 ) | ( ~n15087 & n15088 ) ;
  assign n15090 = n15079 & n15089 ;
  assign n15091 = n15079 | n15089 ;
  assign n15092 = ~n15090 & n15091 ;
  assign n15093 = x23 & ~n4541 ;
  assign n15094 = ( x23 & n12468 ) | ( x23 & n15093 ) | ( n12468 & n15093 ) ;
  assign n15095 = n4554 & n13994 ;
  assign n15096 = n4548 & ~n12468 ;
  assign n15097 = n4551 & ~n12466 ;
  assign n15098 = n15096 | n15097 ;
  assign n15099 = n15095 | n15098 ;
  assign n15100 = x23 | n15099 ;
  assign n15101 = ~x23 & n15100 ;
  assign n15102 = ( ~n15099 & n15100 ) | ( ~n15099 & n15101 ) | ( n15100 & n15101 ) ;
  assign n15103 = n15094 & n15102 ;
  assign n15104 = n4474 & ~n12468 ;
  assign n15105 = n4551 & n12459 ;
  assign n15106 = n4546 & ~n12468 ;
  assign n15107 = n4548 & ~n12466 ;
  assign n15108 = n15106 | n15107 ;
  assign n15109 = n15105 | n15108 ;
  assign n15110 = n4554 & n14003 ;
  assign n15111 = n15109 | n15110 ;
  assign n15112 = ~x23 & n15111 ;
  assign n15113 = x23 | n15112 ;
  assign n15114 = ( ~n15111 & n15112 ) | ( ~n15111 & n15113 ) | ( n15112 & n15113 ) ;
  assign n15115 = n15104 & n15114 ;
  assign n15116 = n15103 & n15115 ;
  assign n15117 = n15103 & n15114 ;
  assign n15118 = n15104 | n15117 ;
  assign n15119 = ~n15116 & n15118 ;
  assign n15120 = n4551 & ~n12456 ;
  assign n15121 = n4546 & ~n12466 ;
  assign n15122 = n4548 & n12459 ;
  assign n15123 = n15121 | n15122 ;
  assign n15124 = n15120 | n15123 ;
  assign n15125 = ( n4554 & n14031 ) | ( n4554 & n15124 ) | ( n14031 & n15124 ) ;
  assign n15126 = ( x23 & ~n15124 ) | ( x23 & n15125 ) | ( ~n15124 & n15125 ) ;
  assign n15127 = ~n15125 & n15126 ;
  assign n15128 = n15124 | n15126 ;
  assign n15129 = ( ~x23 & n15127 ) | ( ~x23 & n15128 ) | ( n15127 & n15128 ) ;
  assign n15130 = n15119 & n15129 ;
  assign n15131 = n15116 | n15130 ;
  assign n15132 = n15092 & n15131 ;
  assign n15133 = n15090 | n15132 ;
  assign n15134 = n15074 | n15076 ;
  assign n15135 = ~n15077 & n15134 ;
  assign n15136 = n15133 & n15135 ;
  assign n15137 = n15077 | n15136 ;
  assign n15138 = n15064 & n15137 ;
  assign n15139 = n15062 | n15138 ;
  assign n15140 = n15048 & ~n15049 ;
  assign n15141 = ( n15038 & ~n15049 ) | ( n15038 & n15140 ) | ( ~n15049 & n15140 ) ;
  assign n15142 = n15139 & n15141 ;
  assign n15143 = n15049 | n15142 ;
  assign n15144 = ( n15025 & n15036 ) | ( n15025 & n15143 ) | ( n15036 & n15143 ) ;
  assign n15145 = n15023 & n15144 ;
  assign n15146 = n15021 | n15145 ;
  assign n15147 = ( ~n15007 & n15008 ) | ( ~n15007 & n15146 ) | ( n15008 & n15146 ) ;
  assign n15148 = n15006 | n15147 ;
  assign n15149 = n14981 | n14992 ;
  assign n15150 = ( ~n14991 & n14992 ) | ( ~n14991 & n15149 ) | ( n14992 & n15149 ) ;
  assign n15151 = n15148 & ~n15150 ;
  assign n15152 = n14992 | n15151 ;
  assign n15153 = n14978 & n15152 ;
  assign n15154 = n14976 | n15153 ;
  assign n15155 = n14951 | n14962 ;
  assign n15156 = ( ~n14961 & n14962 ) | ( ~n14961 & n15155 ) | ( n14962 & n15155 ) ;
  assign n15157 = n15154 & ~n15156 ;
  assign n15158 = n14962 | n15157 ;
  assign n15159 = n14936 & ~n14947 ;
  assign n15160 = n14948 | n15159 ;
  assign n15161 = n15158 & ~n15160 ;
  assign n15162 = n14948 | n15161 ;
  assign n15163 = n14931 | n14933 ;
  assign n15164 = ~n14934 & n15163 ;
  assign n15165 = n15162 & n15164 ;
  assign n15166 = n14934 | n15165 ;
  assign n15167 = n14914 | n14920 ;
  assign n15168 = ~n14921 & n15167 ;
  assign n15169 = n15166 & n15168 ;
  assign n15170 = n14921 | n15169 ;
  assign n15171 = n14893 | n14903 ;
  assign n15172 = ~n14904 & n15171 ;
  assign n15173 = n15170 & n15172 ;
  assign n15174 = n14904 | n15173 ;
  assign n15175 = n14876 | n14886 ;
  assign n15176 = ~n14887 & n15175 ;
  assign n15177 = n15174 & n15176 ;
  assign n15178 = n14887 | n15177 ;
  assign n15179 = n13820 | n14192 ;
  assign n15180 = ~n14193 & n15179 ;
  assign n15181 = n4048 & n12415 ;
  assign n15182 = n4043 & n12419 ;
  assign n15183 = n4045 & n12411 ;
  assign n15184 = n15182 | n15183 ;
  assign n15185 = n15181 | n15184 ;
  assign n15186 = n4051 & ~n13761 ;
  assign n15187 = ~n13762 & n15186 ;
  assign n15188 = ( n4051 & n15185 ) | ( n4051 & ~n15187 ) | ( n15185 & ~n15187 ) ;
  assign n15189 = ~x29 & n15188 ;
  assign n15190 = x29 | n15189 ;
  assign n15191 = ( ~n15188 & n15189 ) | ( ~n15188 & n15190 ) | ( n15189 & n15190 ) ;
  assign n15192 = n15180 & n15191 ;
  assign n15193 = n15180 | n15191 ;
  assign n15194 = ~n15192 & n15193 ;
  assign n15195 = n14642 | n15194 ;
  assign n15196 = n14646 | n15195 ;
  assign n15197 = ( n14642 & n14646 ) | ( n14642 & n15194 ) | ( n14646 & n15194 ) ;
  assign n15198 = n15196 & ~n15197 ;
  assign n15199 = n4484 & n12383 ;
  assign n15200 = n4479 & n12401 ;
  assign n15201 = n4481 & n12392 ;
  assign n15202 = n15200 | n15201 ;
  assign n15203 = n15199 | n15202 ;
  assign n15204 = n4487 | n15203 ;
  assign n15205 = ( n13141 & n15203 ) | ( n13141 & n15204 ) | ( n15203 & n15204 ) ;
  assign n15206 = x26 & n15205 ;
  assign n15207 = x26 & ~n15206 ;
  assign n15208 = ( n15205 & ~n15206 ) | ( n15205 & n15207 ) | ( ~n15206 & n15207 ) ;
  assign n15209 = n15198 & n15208 ;
  assign n15210 = n15198 | n15208 ;
  assign n15211 = ~n15209 & n15210 ;
  assign n15212 = ( n14647 & n14657 ) | ( n14647 & n14873 ) | ( n14657 & n14873 ) ;
  assign n15213 = n15211 & n15212 ;
  assign n15214 = n15211 | n15212 ;
  assign n15215 = ~n15213 & n15214 ;
  assign n15216 = n4551 & n12378 ;
  assign n15217 = n4546 & n12387 ;
  assign n15218 = n4548 & ~n12502 ;
  assign n15219 = n15217 | n15218 ;
  assign n15220 = n15216 | n15219 ;
  assign n15221 = n4554 | n15220 ;
  assign n15222 = ( ~n12816 & n15220 ) | ( ~n12816 & n15221 ) | ( n15220 & n15221 ) ;
  assign n15223 = ~x23 & n15222 ;
  assign n15224 = x23 | n15223 ;
  assign n15225 = ( ~n15222 & n15223 ) | ( ~n15222 & n15224 ) | ( n15223 & n15224 ) ;
  assign n15226 = n15215 & n15225 ;
  assign n15227 = n15225 & ~n15226 ;
  assign n15228 = ( n15215 & ~n15226 ) | ( n15215 & n15227 ) | ( ~n15226 & n15227 ) ;
  assign n15229 = n15178 & n15228 ;
  assign n15230 = n15178 | n15228 ;
  assign n15231 = ~n15229 & n15230 ;
  assign n15232 = n4781 & n12520 ;
  assign n15233 = n4776 & ~n12371 ;
  assign n15234 = n4778 & n12375 ;
  assign n15235 = n15233 | n15234 ;
  assign n15236 = n15232 | n15235 ;
  assign n15237 = n4784 & ~n12837 ;
  assign n15238 = ~n12835 & n15237 ;
  assign n15239 = ( n4784 & n15236 ) | ( n4784 & ~n15238 ) | ( n15236 & ~n15238 ) ;
  assign n15240 = ~x20 & n15239 ;
  assign n15241 = x20 | n15240 ;
  assign n15242 = ( ~n15239 & n15240 ) | ( ~n15239 & n15241 ) | ( n15240 & n15241 ) ;
  assign n15243 = n15231 & n15242 ;
  assign n15244 = n15231 | n15242 ;
  assign n15245 = ~n15243 & n15244 ;
  assign n15246 = n15174 | n15176 ;
  assign n15247 = ~n15177 & n15246 ;
  assign n15248 = n4781 & n12375 ;
  assign n15249 = n4776 & n12378 ;
  assign n15250 = n4778 & ~n12371 ;
  assign n15251 = n15249 | n15250 ;
  assign n15252 = n15248 | n15251 ;
  assign n15253 = n4784 & n13065 ;
  assign n15254 = ~n13064 & n15253 ;
  assign n15255 = ( n4784 & n15252 ) | ( n4784 & ~n15254 ) | ( n15252 & ~n15254 ) ;
  assign n15256 = x20 & n15255 ;
  assign n15257 = x20 & ~n15256 ;
  assign n15258 = ( n15255 & ~n15256 ) | ( n15255 & n15257 ) | ( ~n15256 & n15257 ) ;
  assign n15259 = n15170 | n15172 ;
  assign n15260 = ~n15173 & n15259 ;
  assign n15261 = n4781 & ~n12371 ;
  assign n15262 = n4776 & ~n12502 ;
  assign n15263 = n4778 & n12378 ;
  assign n15264 = n15262 | n15263 ;
  assign n15265 = n15261 | n15264 ;
  assign n15266 = n4784 | n15265 ;
  assign n15267 = ( ~n12848 & n15265 ) | ( ~n12848 & n15266 ) | ( n15265 & n15266 ) ;
  assign n15268 = ~x20 & n15267 ;
  assign n15269 = x20 | n15268 ;
  assign n15270 = ( ~n15267 & n15268 ) | ( ~n15267 & n15269 ) | ( n15268 & n15269 ) ;
  assign n15271 = n15166 | n15168 ;
  assign n15272 = ~n15169 & n15271 ;
  assign n15273 = n4781 & n12378 ;
  assign n15274 = n4776 & n12387 ;
  assign n15275 = n4778 & ~n12502 ;
  assign n15276 = n15274 | n15275 ;
  assign n15277 = n15273 | n15276 ;
  assign n15278 = n4784 | n15277 ;
  assign n15279 = ( ~n12816 & n15277 ) | ( ~n12816 & n15278 ) | ( n15277 & n15278 ) ;
  assign n15280 = ~x20 & n15279 ;
  assign n15281 = x20 | n15280 ;
  assign n15282 = ( ~n15279 & n15280 ) | ( ~n15279 & n15281 ) | ( n15280 & n15281 ) ;
  assign n15283 = ~n15158 & n15160 ;
  assign n15284 = n15161 | n15283 ;
  assign n15285 = n4781 & n12387 ;
  assign n15286 = n4776 & n12392 ;
  assign n15287 = n4778 & n12383 ;
  assign n15288 = n15286 | n15287 ;
  assign n15289 = n15285 | n15288 ;
  assign n15290 = n4784 | n15289 ;
  assign n15291 = ( n12948 & n15289 ) | ( n12948 & n15290 ) | ( n15289 & n15290 ) ;
  assign n15292 = x20 & n15291 ;
  assign n15293 = x20 & ~n15292 ;
  assign n15294 = ( n15291 & ~n15292 ) | ( n15291 & n15293 ) | ( ~n15292 & n15293 ) ;
  assign n15295 = ~n15284 & n15294 ;
  assign n15296 = ~n15154 & n15156 ;
  assign n15297 = n15157 | n15296 ;
  assign n15298 = n4781 & n12383 ;
  assign n15299 = n4776 & n12401 ;
  assign n15300 = n4778 & n12392 ;
  assign n15301 = n15299 | n15300 ;
  assign n15302 = n15298 | n15301 ;
  assign n15303 = n4784 | n15302 ;
  assign n15304 = ( n13141 & n15302 ) | ( n13141 & n15303 ) | ( n15302 & n15303 ) ;
  assign n15305 = x20 & n15304 ;
  assign n15306 = x20 & ~n15305 ;
  assign n15307 = ( n15304 & ~n15305 ) | ( n15304 & n15306 ) | ( ~n15305 & n15306 ) ;
  assign n15308 = ~n15297 & n15307 ;
  assign n15309 = n14978 | n15152 ;
  assign n15310 = ~n15153 & n15309 ;
  assign n15311 = n4781 & n12392 ;
  assign n15312 = n4776 & n12415 ;
  assign n15313 = n4778 & n12401 ;
  assign n15314 = n15312 | n15313 ;
  assign n15315 = n15311 | n15314 ;
  assign n15316 = n4784 | n15315 ;
  assign n15317 = ( n13034 & n15315 ) | ( n13034 & n15316 ) | ( n15315 & n15316 ) ;
  assign n15318 = x20 & n15317 ;
  assign n15319 = x20 & ~n15318 ;
  assign n15320 = ( n15317 & ~n15318 ) | ( n15317 & n15319 ) | ( ~n15318 & n15319 ) ;
  assign n15321 = n15310 & n15320 ;
  assign n15322 = n15310 & ~n15321 ;
  assign n15323 = ~n15310 & n15320 ;
  assign n15324 = n15322 | n15323 ;
  assign n15325 = n4781 & n12401 ;
  assign n15326 = n4776 & n12411 ;
  assign n15327 = n4778 & n12415 ;
  assign n15328 = n15326 | n15327 ;
  assign n15329 = n15325 | n15328 ;
  assign n15330 = n4784 & ~n13163 ;
  assign n15331 = ~n13161 & n15330 ;
  assign n15332 = ( n4784 & n15329 ) | ( n4784 & ~n15331 ) | ( n15329 & ~n15331 ) ;
  assign n15333 = ~x20 & n15332 ;
  assign n15334 = x20 | n15333 ;
  assign n15335 = ( ~n15332 & n15333 ) | ( ~n15332 & n15334 ) | ( n15333 & n15334 ) ;
  assign n15336 = n15008 | n15146 ;
  assign n15337 = n15007 & ~n15336 ;
  assign n15338 = n15147 | n15337 ;
  assign n15339 = n4781 & n12415 ;
  assign n15340 = n4776 & n12419 ;
  assign n15341 = n4778 & n12411 ;
  assign n15342 = n15340 | n15341 ;
  assign n15343 = n15339 | n15342 ;
  assign n15344 = n4784 & ~n13761 ;
  assign n15345 = ~n13762 & n15344 ;
  assign n15346 = ( n4784 & n15343 ) | ( n4784 & ~n15345 ) | ( n15343 & ~n15345 ) ;
  assign n15347 = ~x20 & n15346 ;
  assign n15348 = x20 | n15347 ;
  assign n15349 = ( ~n15346 & n15347 ) | ( ~n15346 & n15348 ) | ( n15347 & n15348 ) ;
  assign n15350 = ~n15338 & n15349 ;
  assign n15351 = n15023 | n15144 ;
  assign n15352 = ~n15145 & n15351 ;
  assign n15353 = n4781 & n12411 ;
  assign n15354 = n4776 & ~n12423 ;
  assign n15355 = n4778 & n12419 ;
  assign n15356 = n15354 | n15355 ;
  assign n15357 = n15353 | n15356 ;
  assign n15358 = n4784 | n15357 ;
  assign n15359 = ( n13776 & n15357 ) | ( n13776 & n15358 ) | ( n15357 & n15358 ) ;
  assign n15360 = x20 & n15359 ;
  assign n15361 = x20 & ~n15360 ;
  assign n15362 = ( n15359 & ~n15360 ) | ( n15359 & n15361 ) | ( ~n15360 & n15361 ) ;
  assign n15363 = n15352 & n15362 ;
  assign n15364 = n15362 & ~n15363 ;
  assign n15365 = ( n15352 & ~n15363 ) | ( n15352 & n15364 ) | ( ~n15363 & n15364 ) ;
  assign n15366 = n4781 & n12419 ;
  assign n15367 = n4776 & n12433 ;
  assign n15368 = n4778 & ~n12423 ;
  assign n15369 = n15367 | n15368 ;
  assign n15370 = n15366 | n15369 ;
  assign n15371 = n4784 | n15370 ;
  assign n15372 = ( ~n13282 & n15370 ) | ( ~n13282 & n15371 ) | ( n15370 & n15371 ) ;
  assign n15373 = ~x20 & n15372 ;
  assign n15374 = x20 | n15373 ;
  assign n15375 = ( ~n15372 & n15373 ) | ( ~n15372 & n15374 ) | ( n15373 & n15374 ) ;
  assign n15376 = ( n15025 & n15143 ) | ( n15025 & ~n15144 ) | ( n15143 & ~n15144 ) ;
  assign n15377 = ( n15036 & ~n15144 ) | ( n15036 & n15376 ) | ( ~n15144 & n15376 ) ;
  assign n15378 = n15375 & n15377 ;
  assign n15379 = n15375 | n15377 ;
  assign n15380 = ~n15378 & n15379 ;
  assign n15381 = n15139 | n15141 ;
  assign n15382 = ~n15142 & n15381 ;
  assign n15383 = n4781 & ~n12423 ;
  assign n15384 = n4776 & ~n12438 ;
  assign n15385 = n4778 & n12433 ;
  assign n15386 = n15384 | n15385 ;
  assign n15387 = n15383 | n15386 ;
  assign n15388 = n4784 | n15387 ;
  assign n15389 = ( ~n13786 & n15387 ) | ( ~n13786 & n15388 ) | ( n15387 & n15388 ) ;
  assign n15390 = ~x20 & n15389 ;
  assign n15391 = x20 | n15390 ;
  assign n15392 = ( ~n15389 & n15390 ) | ( ~n15389 & n15391 ) | ( n15390 & n15391 ) ;
  assign n15393 = n15382 & n15392 ;
  assign n15394 = n15064 | n15137 ;
  assign n15395 = ~n15138 & n15394 ;
  assign n15396 = n4781 & n12433 ;
  assign n15397 = n4776 & n12440 ;
  assign n15398 = n4778 & ~n12438 ;
  assign n15399 = n15397 | n15398 ;
  assign n15400 = n15396 | n15399 ;
  assign n15401 = n4784 | n15400 ;
  assign n15402 = ( ~n14167 & n15400 ) | ( ~n14167 & n15401 ) | ( n15400 & n15401 ) ;
  assign n15403 = ~x20 & n15402 ;
  assign n15404 = x20 | n15403 ;
  assign n15405 = ( ~n15402 & n15403 ) | ( ~n15402 & n15404 ) | ( n15403 & n15404 ) ;
  assign n15406 = n15395 & n15405 ;
  assign n15407 = n15395 & ~n15406 ;
  assign n15408 = ~n15395 & n15405 ;
  assign n15409 = n15407 | n15408 ;
  assign n15410 = n15133 | n15135 ;
  assign n15411 = ~n15136 & n15410 ;
  assign n15412 = n4781 & ~n12438 ;
  assign n15413 = n4776 & n12446 ;
  assign n15414 = n4778 & n12440 ;
  assign n15415 = n15413 | n15414 ;
  assign n15416 = n15412 | n15415 ;
  assign n15417 = n4784 & n14154 ;
  assign n15418 = ~n14156 & n15417 ;
  assign n15419 = ( n4784 & n15416 ) | ( n4784 & ~n15418 ) | ( n15416 & ~n15418 ) ;
  assign n15420 = x20 & n15419 ;
  assign n15421 = x20 & ~n15420 ;
  assign n15422 = ( n15419 & ~n15420 ) | ( n15419 & n15421 ) | ( ~n15420 & n15421 ) ;
  assign n15423 = n15092 | n15131 ;
  assign n15424 = ~n15132 & n15423 ;
  assign n15425 = n4781 & n12440 ;
  assign n15426 = n4776 & n12452 ;
  assign n15427 = n4778 & n12446 ;
  assign n15428 = n15426 | n15427 ;
  assign n15429 = n15425 | n15428 ;
  assign n15430 = n4784 | n15429 ;
  assign n15431 = ( n13822 & n15429 ) | ( n13822 & n15430 ) | ( n15429 & n15430 ) ;
  assign n15432 = x20 & n15431 ;
  assign n15433 = x20 & ~n15432 ;
  assign n15434 = ( n15431 & ~n15432 ) | ( n15431 & n15433 ) | ( ~n15432 & n15433 ) ;
  assign n15435 = n15424 & n15434 ;
  assign n15436 = n4781 & n12446 ;
  assign n15437 = n4776 & n12454 ;
  assign n15438 = n4778 & n12452 ;
  assign n15439 = n15437 | n15438 ;
  assign n15440 = n15436 | n15439 ;
  assign n15441 = n4784 | n15440 ;
  assign n15442 = ( n13862 & n15440 ) | ( n13862 & n15441 ) | ( n15440 & n15441 ) ;
  assign n15443 = x20 & n15442 ;
  assign n15444 = x20 & ~n15443 ;
  assign n15445 = ( n15442 & ~n15443 ) | ( n15442 & n15444 ) | ( ~n15443 & n15444 ) ;
  assign n15446 = n15119 & ~n15130 ;
  assign n15447 = ( n15129 & ~n15130 ) | ( n15129 & n15446 ) | ( ~n15130 & n15446 ) ;
  assign n15448 = n15445 & n15447 ;
  assign n15449 = n15445 | n15447 ;
  assign n15450 = ~n15448 & n15449 ;
  assign n15451 = n4781 & n12452 ;
  assign n15452 = n4776 & ~n12456 ;
  assign n15453 = n4778 & n12454 ;
  assign n15454 = n15452 | n15453 ;
  assign n15455 = n15451 | n15454 ;
  assign n15456 = n4784 | n15455 ;
  assign n15457 = ( ~n13922 & n15455 ) | ( ~n13922 & n15456 ) | ( n15455 & n15456 ) ;
  assign n15458 = ~x20 & n15457 ;
  assign n15459 = x20 & ~n15457 ;
  assign n15460 = n15458 | n15459 ;
  assign n15461 = n15103 | n15114 ;
  assign n15462 = ~n15117 & n15461 ;
  assign n15463 = n15460 & n15462 ;
  assign n15464 = n15094 | n15102 ;
  assign n15465 = ~n15103 & n15464 ;
  assign n15466 = n4781 & n12454 ;
  assign n15467 = n4776 & n12459 ;
  assign n15468 = n4778 & ~n12456 ;
  assign n15469 = n15467 | n15468 ;
  assign n15470 = n15466 | n15469 ;
  assign n15471 = n4784 | n15470 ;
  assign n15472 = ( n14041 & n15470 ) | ( n14041 & n15471 ) | ( n15470 & n15471 ) ;
  assign n15473 = x20 & n15472 ;
  assign n15474 = x20 & ~n15473 ;
  assign n15475 = ( n15472 & ~n15473 ) | ( n15472 & n15474 ) | ( ~n15473 & n15474 ) ;
  assign n15476 = n15465 & n15475 ;
  assign n15477 = n15465 | n15475 ;
  assign n15478 = ~n15476 & n15477 ;
  assign n15479 = x20 & ~n4774 ;
  assign n15480 = ( x20 & n12468 ) | ( x20 & n15479 ) | ( n12468 & n15479 ) ;
  assign n15481 = n4784 & n13994 ;
  assign n15482 = n4778 & ~n12468 ;
  assign n15483 = n4781 & ~n12466 ;
  assign n15484 = n15482 | n15483 ;
  assign n15485 = n15481 | n15484 ;
  assign n15486 = x20 | n15485 ;
  assign n15487 = ~x20 & n15486 ;
  assign n15488 = ( ~n15485 & n15486 ) | ( ~n15485 & n15487 ) | ( n15486 & n15487 ) ;
  assign n15489 = n15480 & n15488 ;
  assign n15490 = n4541 & ~n12468 ;
  assign n15491 = n4781 & n12459 ;
  assign n15492 = n4776 & ~n12468 ;
  assign n15493 = n4778 & ~n12466 ;
  assign n15494 = n15492 | n15493 ;
  assign n15495 = n15491 | n15494 ;
  assign n15496 = n4784 & n14003 ;
  assign n15497 = n15495 | n15496 ;
  assign n15498 = ~x20 & n15497 ;
  assign n15499 = x20 | n15498 ;
  assign n15500 = ( ~n15497 & n15498 ) | ( ~n15497 & n15499 ) | ( n15498 & n15499 ) ;
  assign n15501 = n15490 & n15500 ;
  assign n15502 = n15489 & n15501 ;
  assign n15503 = n15489 & n15500 ;
  assign n15504 = n15490 | n15503 ;
  assign n15505 = ~n15502 & n15504 ;
  assign n15506 = n4781 & ~n12456 ;
  assign n15507 = n4776 & ~n12466 ;
  assign n15508 = n4778 & n12459 ;
  assign n15509 = n15507 | n15508 ;
  assign n15510 = n15506 | n15509 ;
  assign n15511 = ( n4784 & n14031 ) | ( n4784 & n15510 ) | ( n14031 & n15510 ) ;
  assign n15512 = ( x20 & ~n15510 ) | ( x20 & n15511 ) | ( ~n15510 & n15511 ) ;
  assign n15513 = ~n15511 & n15512 ;
  assign n15514 = n15510 | n15512 ;
  assign n15515 = ( ~x20 & n15513 ) | ( ~x20 & n15514 ) | ( n15513 & n15514 ) ;
  assign n15516 = n15505 & n15515 ;
  assign n15517 = n15502 | n15516 ;
  assign n15518 = n15478 & n15517 ;
  assign n15519 = n15476 | n15518 ;
  assign n15520 = n15460 | n15462 ;
  assign n15521 = ~n15463 & n15520 ;
  assign n15522 = n15519 & n15521 ;
  assign n15523 = n15463 | n15522 ;
  assign n15524 = n15450 & n15523 ;
  assign n15525 = n15448 | n15524 ;
  assign n15526 = n15434 & ~n15435 ;
  assign n15527 = ( n15424 & ~n15435 ) | ( n15424 & n15526 ) | ( ~n15435 & n15526 ) ;
  assign n15528 = n15525 & n15527 ;
  assign n15529 = n15435 | n15528 ;
  assign n15530 = ( n15411 & n15422 ) | ( n15411 & n15529 ) | ( n15422 & n15529 ) ;
  assign n15531 = n15409 & n15530 ;
  assign n15532 = n15406 | n15531 ;
  assign n15533 = n15382 | n15392 ;
  assign n15534 = ~n15393 & n15533 ;
  assign n15535 = n15532 & n15534 ;
  assign n15536 = n15393 | n15535 ;
  assign n15537 = n15380 & n15536 ;
  assign n15538 = n15378 | n15537 ;
  assign n15539 = n15365 & n15538 ;
  assign n15540 = n15363 | n15539 ;
  assign n15541 = n15338 | n15350 ;
  assign n15542 = ( ~n15349 & n15350 ) | ( ~n15349 & n15541 ) | ( n15350 & n15541 ) ;
  assign n15543 = n15540 & ~n15542 ;
  assign n15544 = n15350 | n15543 ;
  assign n15545 = ~n15148 & n15150 ;
  assign n15546 = n15151 | n15545 ;
  assign n15547 = ( n15335 & ~n15544 ) | ( n15335 & n15546 ) | ( ~n15544 & n15546 ) ;
  assign n15548 = ( ~n15335 & n15544 ) | ( ~n15335 & n15547 ) | ( n15544 & n15547 ) ;
  assign n15549 = ( ~n15546 & n15547 ) | ( ~n15546 & n15548 ) | ( n15547 & n15548 ) ;
  assign n15550 = ( n15335 & n15544 ) | ( n15335 & n15549 ) | ( n15544 & n15549 ) ;
  assign n15551 = n15324 & n15550 ;
  assign n15552 = n15321 | n15551 ;
  assign n15553 = n15297 | n15308 ;
  assign n15554 = ( ~n15307 & n15308 ) | ( ~n15307 & n15553 ) | ( n15308 & n15553 ) ;
  assign n15555 = n15552 & ~n15554 ;
  assign n15556 = n15308 | n15555 ;
  assign n15557 = n15284 | n15295 ;
  assign n15558 = ( ~n15294 & n15295 ) | ( ~n15294 & n15557 ) | ( n15295 & n15557 ) ;
  assign n15559 = n15556 & ~n15558 ;
  assign n15560 = n15295 | n15559 ;
  assign n15561 = n15162 | n15164 ;
  assign n15562 = ~n15165 & n15561 ;
  assign n15563 = n4781 & ~n12502 ;
  assign n15564 = n4776 & n12383 ;
  assign n15565 = n4778 & n12387 ;
  assign n15566 = n15564 | n15565 ;
  assign n15567 = n15563 | n15566 ;
  assign n15568 = n4784 | n15567 ;
  assign n15569 = ( ~n12756 & n15567 ) | ( ~n12756 & n15568 ) | ( n15567 & n15568 ) ;
  assign n15570 = ~x20 & n15569 ;
  assign n15571 = x20 | n15570 ;
  assign n15572 = ( ~n15569 & n15570 ) | ( ~n15569 & n15571 ) | ( n15570 & n15571 ) ;
  assign n15573 = ( n15560 & n15562 ) | ( n15560 & n15572 ) | ( n15562 & n15572 ) ;
  assign n15574 = ( n15272 & n15282 ) | ( n15272 & n15573 ) | ( n15282 & n15573 ) ;
  assign n15575 = ( n15260 & n15270 ) | ( n15260 & n15574 ) | ( n15270 & n15574 ) ;
  assign n15576 = ( n15247 & n15258 ) | ( n15247 & n15575 ) | ( n15258 & n15575 ) ;
  assign n15577 = n15245 & n15576 ;
  assign n15578 = n15245 | n15576 ;
  assign n15579 = ~n15577 & n15578 ;
  assign n15580 = n5083 & ~n12537 ;
  assign n15581 = n5069 & ~n12360 ;
  assign n15582 = n5070 & n12364 ;
  assign n15583 = n15581 | n15582 ;
  assign n15584 = n15580 | n15583 ;
  assign n15585 = ( n5074 & n13081 ) | ( n5074 & ~n13082 ) | ( n13081 & ~n13082 ) ;
  assign n15586 = n15584 | n15585 ;
  assign n15587 = x17 | n15586 ;
  assign n15588 = ~x17 & n15587 ;
  assign n15589 = ( ~n15586 & n15587 ) | ( ~n15586 & n15588 ) | ( n15587 & n15588 ) ;
  assign n15590 = n15579 & n15589 ;
  assign n15591 = n5083 & n12364 ;
  assign n15592 = n5069 & n12520 ;
  assign n15593 = n5070 & ~n12360 ;
  assign n15594 = n15592 | n15593 ;
  assign n15595 = n15591 | n15594 ;
  assign n15596 = n5074 | n15595 ;
  assign n15597 = ( ~n13113 & n15595 ) | ( ~n13113 & n15596 ) | ( n15595 & n15596 ) ;
  assign n15598 = ~x17 & n15597 ;
  assign n15599 = x17 | n15598 ;
  assign n15600 = ( ~n15597 & n15598 ) | ( ~n15597 & n15599 ) | ( n15598 & n15599 ) ;
  assign n15601 = ( n15247 & n15575 ) | ( n15247 & ~n15576 ) | ( n15575 & ~n15576 ) ;
  assign n15602 = ( n15258 & ~n15576 ) | ( n15258 & n15601 ) | ( ~n15576 & n15601 ) ;
  assign n15603 = n15600 & n15602 ;
  assign n15604 = n5083 & ~n12360 ;
  assign n15605 = n5069 & n12375 ;
  assign n15606 = n5070 & n12520 ;
  assign n15607 = n15605 | n15606 ;
  assign n15608 = n15604 | n15607 ;
  assign n15609 = n5074 | n15608 ;
  assign n15610 = ( ~n12902 & n15608 ) | ( ~n12902 & n15609 ) | ( n15608 & n15609 ) ;
  assign n15611 = ~x17 & n15610 ;
  assign n15612 = x17 | n15611 ;
  assign n15613 = ( ~n15610 & n15611 ) | ( ~n15610 & n15612 ) | ( n15611 & n15612 ) ;
  assign n15614 = ( n15260 & n15574 ) | ( n15260 & ~n15575 ) | ( n15574 & ~n15575 ) ;
  assign n15615 = ( n15270 & ~n15575 ) | ( n15270 & n15614 ) | ( ~n15575 & n15614 ) ;
  assign n15616 = n15613 & n15615 ;
  assign n15617 = n5083 & n12520 ;
  assign n15618 = n5069 & ~n12371 ;
  assign n15619 = n5070 & n12375 ;
  assign n15620 = n15618 | n15619 ;
  assign n15621 = n15617 | n15620 ;
  assign n15622 = n5074 & n12837 ;
  assign n15623 = ( n5074 & n12835 ) | ( n5074 & n15622 ) | ( n12835 & n15622 ) ;
  assign n15624 = n15621 | n15623 ;
  assign n15625 = x17 | n15624 ;
  assign n15626 = ~x17 & n15625 ;
  assign n15627 = ( ~n15624 & n15625 ) | ( ~n15624 & n15626 ) | ( n15625 & n15626 ) ;
  assign n15628 = ( n15272 & n15573 ) | ( n15272 & ~n15574 ) | ( n15573 & ~n15574 ) ;
  assign n15629 = ( n15282 & ~n15574 ) | ( n15282 & n15628 ) | ( ~n15574 & n15628 ) ;
  assign n15630 = n15627 & n15629 ;
  assign n15631 = n5083 & n12375 ;
  assign n15632 = n5069 & n12378 ;
  assign n15633 = n5070 & ~n12371 ;
  assign n15634 = n15632 | n15633 ;
  assign n15635 = n15631 | n15634 ;
  assign n15636 = ( n5074 & n13064 ) | ( n5074 & ~n13065 ) | ( n13064 & ~n13065 ) ;
  assign n15637 = n15635 | n15636 ;
  assign n15638 = x17 | n15637 ;
  assign n15639 = ~x17 & n15638 ;
  assign n15640 = ( ~n15637 & n15638 ) | ( ~n15637 & n15639 ) | ( n15638 & n15639 ) ;
  assign n15641 = ( n15560 & ~n15562 ) | ( n15560 & n15572 ) | ( ~n15562 & n15572 ) ;
  assign n15642 = ( ~n15560 & n15562 ) | ( ~n15560 & n15641 ) | ( n15562 & n15641 ) ;
  assign n15643 = ( ~n15572 & n15641 ) | ( ~n15572 & n15642 ) | ( n15641 & n15642 ) ;
  assign n15644 = n15640 & n15643 ;
  assign n15645 = n15640 | n15643 ;
  assign n15646 = ~n15644 & n15645 ;
  assign n15647 = n15556 & ~n15559 ;
  assign n15648 = n15558 | n15559 ;
  assign n15649 = ~n15647 & n15648 ;
  assign n15650 = n5083 & ~n12371 ;
  assign n15651 = n5069 & ~n12502 ;
  assign n15652 = n5070 & n12378 ;
  assign n15653 = n15651 | n15652 ;
  assign n15654 = n15650 | n15653 ;
  assign n15655 = n5074 | n15654 ;
  assign n15656 = ( ~n12848 & n15654 ) | ( ~n12848 & n15655 ) | ( n15654 & n15655 ) ;
  assign n15657 = ~x17 & n15656 ;
  assign n15658 = x17 | n15657 ;
  assign n15659 = ( ~n15656 & n15657 ) | ( ~n15656 & n15658 ) | ( n15657 & n15658 ) ;
  assign n15660 = ~n15649 & n15659 ;
  assign n15661 = n15552 & ~n15555 ;
  assign n15662 = n15554 | n15555 ;
  assign n15663 = ~n15661 & n15662 ;
  assign n15664 = n5083 & n12378 ;
  assign n15665 = n5069 & n12387 ;
  assign n15666 = n5070 & ~n12502 ;
  assign n15667 = n15665 | n15666 ;
  assign n15668 = n15664 | n15667 ;
  assign n15669 = n5074 | n15668 ;
  assign n15670 = ( ~n12816 & n15668 ) | ( ~n12816 & n15669 ) | ( n15668 & n15669 ) ;
  assign n15671 = ~x17 & n15670 ;
  assign n15672 = x17 | n15671 ;
  assign n15673 = ( ~n15670 & n15671 ) | ( ~n15670 & n15672 ) | ( n15671 & n15672 ) ;
  assign n15674 = ~n15663 & n15673 ;
  assign n15675 = n15550 & ~n15551 ;
  assign n15676 = n15324 & ~n15551 ;
  assign n15677 = n15675 | n15676 ;
  assign n15678 = n5083 & ~n12502 ;
  assign n15679 = n5069 & n12383 ;
  assign n15680 = n5070 & n12387 ;
  assign n15681 = n15679 | n15680 ;
  assign n15682 = n15678 | n15681 ;
  assign n15683 = n5074 | n15682 ;
  assign n15684 = ( ~n12756 & n15682 ) | ( ~n12756 & n15683 ) | ( n15682 & n15683 ) ;
  assign n15685 = ~x17 & n15684 ;
  assign n15686 = x17 | n15685 ;
  assign n15687 = ( ~n15684 & n15685 ) | ( ~n15684 & n15686 ) | ( n15685 & n15686 ) ;
  assign n15688 = n15677 & n15687 ;
  assign n15689 = n15677 & ~n15688 ;
  assign n15690 = ~n15677 & n15687 ;
  assign n15691 = n15689 | n15690 ;
  assign n15692 = n5083 & n12387 ;
  assign n15693 = n5069 & n12392 ;
  assign n15694 = n5070 & n12383 ;
  assign n15695 = n15693 | n15694 ;
  assign n15696 = n15692 | n15695 ;
  assign n15697 = n5074 | n15696 ;
  assign n15698 = ( n12948 & n15696 ) | ( n12948 & n15697 ) | ( n15696 & n15697 ) ;
  assign n15699 = x17 & n15698 ;
  assign n15700 = x17 & ~n15699 ;
  assign n15701 = ( n15698 & ~n15699 ) | ( n15698 & n15700 ) | ( ~n15699 & n15700 ) ;
  assign n15702 = ~n15549 & n15701 ;
  assign n15703 = n15549 & ~n15701 ;
  assign n15704 = n15702 | n15703 ;
  assign n15705 = n15540 & ~n15543 ;
  assign n15706 = n15542 | n15543 ;
  assign n15707 = ~n15705 & n15706 ;
  assign n15708 = n5083 & n12383 ;
  assign n15709 = n5069 & n12401 ;
  assign n15710 = n5070 & n12392 ;
  assign n15711 = n15709 | n15710 ;
  assign n15712 = n15708 | n15711 ;
  assign n15713 = n5074 | n15712 ;
  assign n15714 = ( n13141 & n15712 ) | ( n13141 & n15713 ) | ( n15712 & n15713 ) ;
  assign n15715 = x17 & n15714 ;
  assign n15716 = x17 & ~n15715 ;
  assign n15717 = ( n15714 & ~n15715 ) | ( n15714 & n15716 ) | ( ~n15715 & n15716 ) ;
  assign n15718 = ~n15707 & n15717 ;
  assign n15719 = n15365 | n15538 ;
  assign n15720 = ~n15539 & n15719 ;
  assign n15721 = n5083 & n12392 ;
  assign n15722 = n5069 & n12415 ;
  assign n15723 = n5070 & n12401 ;
  assign n15724 = n15722 | n15723 ;
  assign n15725 = n15721 | n15724 ;
  assign n15726 = n5074 | n15725 ;
  assign n15727 = ( n13034 & n15725 ) | ( n13034 & n15726 ) | ( n15725 & n15726 ) ;
  assign n15728 = x17 & n15727 ;
  assign n15729 = x17 & ~n15728 ;
  assign n15730 = ( n15727 & ~n15728 ) | ( n15727 & n15729 ) | ( ~n15728 & n15729 ) ;
  assign n15731 = n15720 & n15730 ;
  assign n15732 = n15380 | n15536 ;
  assign n15733 = ~n15537 & n15732 ;
  assign n15734 = n5083 & n12401 ;
  assign n15735 = n5069 & n12411 ;
  assign n15736 = n5070 & n12415 ;
  assign n15737 = n15735 | n15736 ;
  assign n15738 = n15734 | n15737 ;
  assign n15739 = n5074 & ~n13163 ;
  assign n15740 = ~n13161 & n15739 ;
  assign n15741 = ( n5074 & n15738 ) | ( n5074 & ~n15740 ) | ( n15738 & ~n15740 ) ;
  assign n15742 = ~x17 & n15741 ;
  assign n15743 = x17 | n15742 ;
  assign n15744 = ( ~n15741 & n15742 ) | ( ~n15741 & n15743 ) | ( n15742 & n15743 ) ;
  assign n15745 = n15733 & n15744 ;
  assign n15746 = n15532 | n15534 ;
  assign n15747 = ~n15535 & n15746 ;
  assign n15748 = n5083 & n12415 ;
  assign n15749 = n5069 & n12419 ;
  assign n15750 = n5070 & n12411 ;
  assign n15751 = n15749 | n15750 ;
  assign n15752 = n15748 | n15751 ;
  assign n15753 = ( n5074 & n13761 ) | ( n5074 & n13762 ) | ( n13761 & n13762 ) ;
  assign n15754 = n15752 | n15753 ;
  assign n15755 = x17 | n15754 ;
  assign n15756 = ~x17 & n15755 ;
  assign n15757 = ( ~n15754 & n15755 ) | ( ~n15754 & n15756 ) | ( n15755 & n15756 ) ;
  assign n15758 = n15747 & n15757 ;
  assign n15759 = n15757 & ~n15758 ;
  assign n15760 = ( n15747 & ~n15758 ) | ( n15747 & n15759 ) | ( ~n15758 & n15759 ) ;
  assign n15761 = n5083 & n12411 ;
  assign n15762 = n5069 & ~n12423 ;
  assign n15763 = n5070 & n12419 ;
  assign n15764 = n15762 | n15763 ;
  assign n15765 = n15761 | n15764 ;
  assign n15766 = n5074 | n15765 ;
  assign n15767 = ( n13776 & n15765 ) | ( n13776 & n15766 ) | ( n15765 & n15766 ) ;
  assign n15768 = x17 & n15767 ;
  assign n15769 = x17 & ~n15768 ;
  assign n15770 = ( n15767 & ~n15768 ) | ( n15767 & n15769 ) | ( ~n15768 & n15769 ) ;
  assign n15771 = n15409 & ~n15531 ;
  assign n15772 = ( n15530 & ~n15531 ) | ( n15530 & n15771 ) | ( ~n15531 & n15771 ) ;
  assign n15773 = n15770 & n15772 ;
  assign n15774 = n15772 & ~n15773 ;
  assign n15775 = n15770 & ~n15772 ;
  assign n15776 = n15774 | n15775 ;
  assign n15777 = n5083 & n12419 ;
  assign n15778 = n5069 & n12433 ;
  assign n15779 = n5070 & ~n12423 ;
  assign n15780 = n15778 | n15779 ;
  assign n15781 = n15777 | n15780 ;
  assign n15782 = n5074 | n15781 ;
  assign n15783 = ( ~n13282 & n15781 ) | ( ~n13282 & n15782 ) | ( n15781 & n15782 ) ;
  assign n15784 = ~x17 & n15783 ;
  assign n15785 = x17 | n15784 ;
  assign n15786 = ( ~n15783 & n15784 ) | ( ~n15783 & n15785 ) | ( n15784 & n15785 ) ;
  assign n15787 = ( n15411 & n15529 ) | ( n15411 & ~n15530 ) | ( n15529 & ~n15530 ) ;
  assign n15788 = ( n15422 & ~n15530 ) | ( n15422 & n15787 ) | ( ~n15530 & n15787 ) ;
  assign n15789 = n15786 & n15788 ;
  assign n15790 = n15786 | n15788 ;
  assign n15791 = ~n15789 & n15790 ;
  assign n15792 = n15525 | n15527 ;
  assign n15793 = ~n15528 & n15792 ;
  assign n15794 = n5083 & ~n12423 ;
  assign n15795 = n5069 & ~n12438 ;
  assign n15796 = n5070 & n12433 ;
  assign n15797 = n15795 | n15796 ;
  assign n15798 = n15794 | n15797 ;
  assign n15799 = n5074 | n15798 ;
  assign n15800 = ( ~n13786 & n15798 ) | ( ~n13786 & n15799 ) | ( n15798 & n15799 ) ;
  assign n15801 = ~x17 & n15800 ;
  assign n15802 = x17 | n15801 ;
  assign n15803 = ( ~n15800 & n15801 ) | ( ~n15800 & n15802 ) | ( n15801 & n15802 ) ;
  assign n15804 = n15793 & n15803 ;
  assign n15805 = n15450 | n15523 ;
  assign n15806 = ~n15524 & n15805 ;
  assign n15807 = n5083 & n12433 ;
  assign n15808 = n5069 & n12440 ;
  assign n15809 = n5070 & ~n12438 ;
  assign n15810 = n15808 | n15809 ;
  assign n15811 = n15807 | n15810 ;
  assign n15812 = n5074 | n15811 ;
  assign n15813 = ( ~n14167 & n15811 ) | ( ~n14167 & n15812 ) | ( n15811 & n15812 ) ;
  assign n15814 = ~x17 & n15813 ;
  assign n15815 = x17 | n15814 ;
  assign n15816 = ( ~n15813 & n15814 ) | ( ~n15813 & n15815 ) | ( n15814 & n15815 ) ;
  assign n15817 = n15806 & n15816 ;
  assign n15818 = n15806 & ~n15817 ;
  assign n15819 = ~n15806 & n15816 ;
  assign n15820 = n15818 | n15819 ;
  assign n15821 = n15519 | n15521 ;
  assign n15822 = ~n15522 & n15821 ;
  assign n15823 = n5083 & ~n12438 ;
  assign n15824 = n5069 & n12446 ;
  assign n15825 = n5070 & n12440 ;
  assign n15826 = n15824 | n15825 ;
  assign n15827 = n15823 | n15826 ;
  assign n15828 = n5074 & n14154 ;
  assign n15829 = ~n14156 & n15828 ;
  assign n15830 = ( n5074 & n15827 ) | ( n5074 & ~n15829 ) | ( n15827 & ~n15829 ) ;
  assign n15831 = x17 & n15830 ;
  assign n15832 = x17 & ~n15831 ;
  assign n15833 = ( n15830 & ~n15831 ) | ( n15830 & n15832 ) | ( ~n15831 & n15832 ) ;
  assign n15834 = n15478 | n15517 ;
  assign n15835 = ~n15518 & n15834 ;
  assign n15836 = n5083 & n12440 ;
  assign n15837 = n5069 & n12452 ;
  assign n15838 = n5070 & n12446 ;
  assign n15839 = n15837 | n15838 ;
  assign n15840 = n15836 | n15839 ;
  assign n15841 = n5074 | n15840 ;
  assign n15842 = ( n13822 & n15840 ) | ( n13822 & n15841 ) | ( n15840 & n15841 ) ;
  assign n15843 = x17 & n15842 ;
  assign n15844 = x17 & ~n15843 ;
  assign n15845 = ( n15842 & ~n15843 ) | ( n15842 & n15844 ) | ( ~n15843 & n15844 ) ;
  assign n15846 = n15835 & n15845 ;
  assign n15847 = n5083 & n12446 ;
  assign n15848 = n5069 & n12454 ;
  assign n15849 = n5070 & n12452 ;
  assign n15850 = n15848 | n15849 ;
  assign n15851 = n15847 | n15850 ;
  assign n15852 = n5074 | n15851 ;
  assign n15853 = ( n13862 & n15851 ) | ( n13862 & n15852 ) | ( n15851 & n15852 ) ;
  assign n15854 = x17 & n15853 ;
  assign n15855 = x17 & ~n15854 ;
  assign n15856 = ( n15853 & ~n15854 ) | ( n15853 & n15855 ) | ( ~n15854 & n15855 ) ;
  assign n15857 = n15505 & ~n15516 ;
  assign n15858 = ( n15515 & ~n15516 ) | ( n15515 & n15857 ) | ( ~n15516 & n15857 ) ;
  assign n15859 = n15856 & n15858 ;
  assign n15860 = n15856 | n15858 ;
  assign n15861 = ~n15859 & n15860 ;
  assign n15862 = n5083 & n12452 ;
  assign n15863 = n5069 & ~n12456 ;
  assign n15864 = n5070 & n12454 ;
  assign n15865 = n15863 | n15864 ;
  assign n15866 = n15862 | n15865 ;
  assign n15867 = n5074 | n15866 ;
  assign n15868 = ( ~n13922 & n15866 ) | ( ~n13922 & n15867 ) | ( n15866 & n15867 ) ;
  assign n15869 = ~x17 & n15868 ;
  assign n15870 = x17 & ~n15868 ;
  assign n15871 = n15869 | n15870 ;
  assign n15872 = n15489 | n15500 ;
  assign n15873 = ~n15503 & n15872 ;
  assign n15874 = n15871 & n15873 ;
  assign n15875 = n15480 | n15488 ;
  assign n15876 = ~n15489 & n15875 ;
  assign n15877 = n5083 & n12454 ;
  assign n15878 = n5069 & n12459 ;
  assign n15879 = n5070 & ~n12456 ;
  assign n15880 = n15878 | n15879 ;
  assign n15881 = n15877 | n15880 ;
  assign n15882 = n5074 | n15881 ;
  assign n15883 = ( n14041 & n15881 ) | ( n14041 & n15882 ) | ( n15881 & n15882 ) ;
  assign n15884 = x17 & n15883 ;
  assign n15885 = x17 & ~n15884 ;
  assign n15886 = ( n15883 & ~n15884 ) | ( n15883 & n15885 ) | ( ~n15884 & n15885 ) ;
  assign n15887 = n15876 & n15886 ;
  assign n15888 = n15876 | n15886 ;
  assign n15889 = ~n15887 & n15888 ;
  assign n15890 = x17 & ~n5064 ;
  assign n15891 = ( x17 & n12468 ) | ( x17 & n15890 ) | ( n12468 & n15890 ) ;
  assign n15892 = n5074 & n13994 ;
  assign n15893 = n5070 & ~n12468 ;
  assign n15894 = n5083 & ~n12466 ;
  assign n15895 = n15893 | n15894 ;
  assign n15896 = n15892 | n15895 ;
  assign n15897 = x17 | n15896 ;
  assign n15898 = ~x17 & n15897 ;
  assign n15899 = ( ~n15896 & n15897 ) | ( ~n15896 & n15898 ) | ( n15897 & n15898 ) ;
  assign n15900 = n15891 & n15899 ;
  assign n15901 = n4774 & ~n12468 ;
  assign n15902 = n5083 & n12459 ;
  assign n15903 = n5069 & ~n12468 ;
  assign n15904 = n5070 & ~n12466 ;
  assign n15905 = n15903 | n15904 ;
  assign n15906 = n15902 | n15905 ;
  assign n15907 = n5074 & n14003 ;
  assign n15908 = n15906 | n15907 ;
  assign n15909 = ~x17 & n15908 ;
  assign n15910 = x17 | n15909 ;
  assign n15911 = ( ~n15908 & n15909 ) | ( ~n15908 & n15910 ) | ( n15909 & n15910 ) ;
  assign n15912 = n15901 & n15911 ;
  assign n15913 = n15900 & n15912 ;
  assign n15914 = n15900 & n15911 ;
  assign n15915 = n15901 | n15914 ;
  assign n15916 = ~n15913 & n15915 ;
  assign n15917 = n5083 & ~n12456 ;
  assign n15918 = n5069 & ~n12466 ;
  assign n15919 = n5070 & n12459 ;
  assign n15920 = n15918 | n15919 ;
  assign n15921 = n15917 | n15920 ;
  assign n15922 = ( n5074 & n14031 ) | ( n5074 & n15921 ) | ( n14031 & n15921 ) ;
  assign n15923 = ( x17 & ~n15921 ) | ( x17 & n15922 ) | ( ~n15921 & n15922 ) ;
  assign n15924 = ~n15922 & n15923 ;
  assign n15925 = n15921 | n15923 ;
  assign n15926 = ( ~x17 & n15924 ) | ( ~x17 & n15925 ) | ( n15924 & n15925 ) ;
  assign n15927 = n15916 & n15926 ;
  assign n15928 = n15913 | n15927 ;
  assign n15929 = n15889 & n15928 ;
  assign n15930 = n15887 | n15929 ;
  assign n15931 = n15871 | n15873 ;
  assign n15932 = ~n15874 & n15931 ;
  assign n15933 = n15930 & n15932 ;
  assign n15934 = n15874 | n15933 ;
  assign n15935 = n15861 & n15934 ;
  assign n15936 = n15859 | n15935 ;
  assign n15937 = n15845 & ~n15846 ;
  assign n15938 = ( n15835 & ~n15846 ) | ( n15835 & n15937 ) | ( ~n15846 & n15937 ) ;
  assign n15939 = n15936 & n15938 ;
  assign n15940 = n15846 | n15939 ;
  assign n15941 = ( n15822 & n15833 ) | ( n15822 & n15940 ) | ( n15833 & n15940 ) ;
  assign n15942 = n15820 & n15941 ;
  assign n15943 = n15817 | n15942 ;
  assign n15944 = n15793 | n15803 ;
  assign n15945 = ~n15804 & n15944 ;
  assign n15946 = n15943 & n15945 ;
  assign n15947 = n15804 | n15946 ;
  assign n15948 = n15791 & n15947 ;
  assign n15949 = n15789 | n15948 ;
  assign n15950 = n15776 & n15949 ;
  assign n15951 = n15773 | n15950 ;
  assign n15952 = n15760 & n15951 ;
  assign n15953 = n15758 | n15952 ;
  assign n15954 = n15733 & ~n15745 ;
  assign n15955 = ~n15733 & n15744 ;
  assign n15956 = n15954 | n15955 ;
  assign n15957 = n15953 & n15956 ;
  assign n15958 = n15720 | n15730 ;
  assign n15959 = ~n15731 & n15958 ;
  assign n15960 = ( n15745 & n15957 ) | ( n15745 & n15959 ) | ( n15957 & n15959 ) ;
  assign n15961 = n15731 | n15960 ;
  assign n15962 = n15707 | n15718 ;
  assign n15963 = ( ~n15717 & n15718 ) | ( ~n15717 & n15962 ) | ( n15718 & n15962 ) ;
  assign n15964 = n15961 & ~n15963 ;
  assign n15965 = n15718 | n15964 ;
  assign n15966 = ~n15704 & n15965 ;
  assign n15967 = n15702 | n15966 ;
  assign n15968 = n15691 & n15967 ;
  assign n15969 = n15688 | n15968 ;
  assign n15970 = n15663 | n15674 ;
  assign n15971 = ( ~n15673 & n15674 ) | ( ~n15673 & n15970 ) | ( n15674 & n15970 ) ;
  assign n15972 = n15969 & ~n15971 ;
  assign n15973 = n15674 | n15972 ;
  assign n15974 = n15649 | n15660 ;
  assign n15975 = ( ~n15659 & n15660 ) | ( ~n15659 & n15974 ) | ( n15660 & n15974 ) ;
  assign n15976 = n15973 & ~n15975 ;
  assign n15977 = n15660 | n15976 ;
  assign n15978 = n15646 & n15977 ;
  assign n15979 = n15644 | n15978 ;
  assign n15980 = n15627 | n15629 ;
  assign n15981 = ~n15630 & n15980 ;
  assign n15982 = n15979 & n15981 ;
  assign n15983 = n15630 | n15982 ;
  assign n15984 = n15613 | n15615 ;
  assign n15985 = ~n15616 & n15984 ;
  assign n15986 = n15983 & n15985 ;
  assign n15987 = n15616 | n15986 ;
  assign n15988 = n15600 | n15602 ;
  assign n15989 = ~n15603 & n15988 ;
  assign n15990 = n15987 & n15989 ;
  assign n15991 = n15603 | n15990 ;
  assign n15992 = n15589 & ~n15590 ;
  assign n15993 = ( n15579 & ~n15590 ) | ( n15579 & n15992 ) | ( ~n15590 & n15992 ) ;
  assign n15994 = n15991 & n15993 ;
  assign n15995 = n15590 | n15994 ;
  assign n15996 = n5083 & n12351 ;
  assign n15997 = n5069 & n12364 ;
  assign n15998 = n5070 & ~n12537 ;
  assign n15999 = n15997 | n15998 ;
  assign n16000 = n15996 | n15999 ;
  assign n16001 = n5074 & ~n12928 ;
  assign n16002 = ( n5074 & n12925 ) | ( n5074 & n16001 ) | ( n12925 & n16001 ) ;
  assign n16003 = n16000 | n16002 ;
  assign n16004 = x17 | n16003 ;
  assign n16005 = ~x17 & n16004 ;
  assign n16006 = ( ~n16003 & n16004 ) | ( ~n16003 & n16005 ) | ( n16004 & n16005 ) ;
  assign n16007 = n15243 | n15577 ;
  assign n16008 = n4781 & ~n12360 ;
  assign n16009 = n4776 & n12375 ;
  assign n16010 = n4778 & n12520 ;
  assign n16011 = n16009 | n16010 ;
  assign n16012 = n16008 | n16011 ;
  assign n16013 = n4784 | n16012 ;
  assign n16014 = ( ~n12902 & n16012 ) | ( ~n12902 & n16013 ) | ( n16012 & n16013 ) ;
  assign n16015 = ~x20 & n16014 ;
  assign n16016 = x20 | n16015 ;
  assign n16017 = ( ~n16014 & n16015 ) | ( ~n16014 & n16016 ) | ( n16015 & n16016 ) ;
  assign n16018 = n15226 | n15229 ;
  assign n16019 = n4551 & ~n12371 ;
  assign n16020 = n4546 & ~n12502 ;
  assign n16021 = n4548 & n12378 ;
  assign n16022 = n16020 | n16021 ;
  assign n16023 = n16019 | n16022 ;
  assign n16024 = n4554 | n16023 ;
  assign n16025 = ( ~n12848 & n16023 ) | ( ~n12848 & n16024 ) | ( n16023 & n16024 ) ;
  assign n16026 = ~x23 & n16025 ;
  assign n16027 = x23 | n16026 ;
  assign n16028 = ( ~n16025 & n16026 ) | ( ~n16025 & n16027 ) | ( n16026 & n16027 ) ;
  assign n16029 = n15209 | n15213 ;
  assign n16030 = n14203 & ~n14214 ;
  assign n16031 = n14215 | n16030 ;
  assign n16032 = n4484 & n12387 ;
  assign n16033 = n4479 & n12392 ;
  assign n16034 = n4481 & n12383 ;
  assign n16035 = n16033 | n16034 ;
  assign n16036 = n16032 | n16035 ;
  assign n16037 = n4487 | n16036 ;
  assign n16038 = ( n12948 & n16036 ) | ( n12948 & n16037 ) | ( n16036 & n16037 ) ;
  assign n16039 = x26 & n16038 ;
  assign n16040 = x26 & ~n16039 ;
  assign n16041 = ( n16038 & ~n16039 ) | ( n16038 & n16040 ) | ( ~n16039 & n16040 ) ;
  assign n16042 = n15192 | n15197 ;
  assign n16043 = ( n16031 & n16041 ) | ( n16031 & ~n16042 ) | ( n16041 & ~n16042 ) ;
  assign n16044 = ( ~n16041 & n16042 ) | ( ~n16041 & n16043 ) | ( n16042 & n16043 ) ;
  assign n16045 = ( ~n16031 & n16043 ) | ( ~n16031 & n16044 ) | ( n16043 & n16044 ) ;
  assign n16046 = ( n16028 & ~n16029 ) | ( n16028 & n16045 ) | ( ~n16029 & n16045 ) ;
  assign n16047 = ( n16029 & ~n16045 ) | ( n16029 & n16046 ) | ( ~n16045 & n16046 ) ;
  assign n16048 = ( ~n16028 & n16046 ) | ( ~n16028 & n16047 ) | ( n16046 & n16047 ) ;
  assign n16049 = ( n16017 & ~n16018 ) | ( n16017 & n16048 ) | ( ~n16018 & n16048 ) ;
  assign n16050 = ( n16018 & ~n16048 ) | ( n16018 & n16049 ) | ( ~n16048 & n16049 ) ;
  assign n16051 = ( ~n16017 & n16049 ) | ( ~n16017 & n16050 ) | ( n16049 & n16050 ) ;
  assign n16052 = ( n16006 & ~n16007 ) | ( n16006 & n16051 ) | ( ~n16007 & n16051 ) ;
  assign n16053 = ( n16007 & ~n16051 ) | ( n16007 & n16052 ) | ( ~n16051 & n16052 ) ;
  assign n16054 = ( ~n16006 & n16052 ) | ( ~n16006 & n16053 ) | ( n16052 & n16053 ) ;
  assign n16055 = n7280 & n12553 ;
  assign n16056 = n5384 & n12355 ;
  assign n16057 = n7277 & n12558 ;
  assign n16058 = n16056 | n16057 ;
  assign n16059 = n16055 | n16058 ;
  assign n16060 = n39 | n16059 ;
  assign n16061 = ( n13097 & n16059 ) | ( n13097 & n16060 ) | ( n16059 & n16060 ) ;
  assign n16062 = x14 & n16061 ;
  assign n16063 = x14 & ~n16062 ;
  assign n16064 = ( n16061 & ~n16062 ) | ( n16061 & n16063 ) | ( ~n16062 & n16063 ) ;
  assign n16065 = ( ~n15995 & n16054 ) | ( ~n15995 & n16064 ) | ( n16054 & n16064 ) ;
  assign n16066 = ( n15995 & ~n16054 ) | ( n15995 & n16065 ) | ( ~n16054 & n16065 ) ;
  assign n16067 = n7305 & n12580 ;
  assign n16068 = n7300 & ~n12344 ;
  assign n16069 = n7302 & ~n12586 ;
  assign n16070 = n16068 | n16069 ;
  assign n16071 = n16067 | n16070 ;
  assign n16072 = n7308 | n16071 ;
  assign n16073 = ( n13432 & n16071 ) | ( n13432 & n16072 ) | ( n16071 & n16072 ) ;
  assign n16074 = x11 & n16073 ;
  assign n16075 = x11 & ~n16074 ;
  assign n16076 = ( n16073 & ~n16074 ) | ( n16073 & n16075 ) | ( ~n16074 & n16075 ) ;
  assign n16077 = n7280 & n12340 ;
  assign n16078 = n5384 & n12558 ;
  assign n16079 = n7277 & n12553 ;
  assign n16080 = n16078 | n16079 ;
  assign n16081 = n16077 | n16080 ;
  assign n16082 = n39 & n13347 ;
  assign n16083 = ( n39 & n13346 ) | ( n39 & n16082 ) | ( n13346 & n16082 ) ;
  assign n16084 = n16081 | n16083 ;
  assign n16085 = x14 | n16084 ;
  assign n16086 = ~x14 & n16085 ;
  assign n16087 = ( ~n16084 & n16085 ) | ( ~n16084 & n16086 ) | ( n16085 & n16086 ) ;
  assign n16088 = n5083 & n12355 ;
  assign n16089 = n5069 & ~n12537 ;
  assign n16090 = n5070 & n12351 ;
  assign n16091 = n16089 | n16090 ;
  assign n16092 = n16088 | n16091 ;
  assign n16093 = n5074 | n16092 ;
  assign n16094 = ( n13409 & n16092 ) | ( n13409 & n16093 ) | ( n16092 & n16093 ) ;
  assign n16095 = x17 & n16094 ;
  assign n16096 = x17 & ~n16095 ;
  assign n16097 = ( n16094 & ~n16095 ) | ( n16094 & n16096 ) | ( ~n16095 & n16096 ) ;
  assign n16098 = n4781 & n12364 ;
  assign n16099 = n4776 & n12520 ;
  assign n16100 = n4778 & ~n12360 ;
  assign n16101 = n16099 | n16100 ;
  assign n16102 = n16098 | n16101 ;
  assign n16103 = n4784 | n16102 ;
  assign n16104 = ( ~n13113 & n16102 ) | ( ~n13113 & n16103 ) | ( n16102 & n16103 ) ;
  assign n16105 = ~x20 & n16104 ;
  assign n16106 = x20 | n16105 ;
  assign n16107 = ( ~n16104 & n16105 ) | ( ~n16104 & n16106 ) | ( n16105 & n16106 ) ;
  assign n16145 = ( ~n16031 & n16041 ) | ( ~n16031 & n16045 ) | ( n16041 & n16045 ) ;
  assign n16108 = n4048 & n12392 ;
  assign n16109 = n4043 & n12415 ;
  assign n16110 = n4045 & n12401 ;
  assign n16111 = n16109 | n16110 ;
  assign n16112 = n16108 | n16111 ;
  assign n16113 = n4051 | n16112 ;
  assign n16114 = ( n13034 & n16112 ) | ( n13034 & n16113 ) | ( n16112 & n16113 ) ;
  assign n16115 = x29 & n16114 ;
  assign n16116 = x29 & ~n16115 ;
  assign n16117 = ( n16114 & ~n16115 ) | ( n16114 & n16116 ) | ( ~n16115 & n16116 ) ;
  assign n16118 = n14219 & n16117 ;
  assign n16119 = n14219 & ~n16118 ;
  assign n16120 = ~n14219 & n16117 ;
  assign n16121 = n16119 | n16120 ;
  assign n16122 = n4481 & n12387 ;
  assign n16123 = n4484 & ~n12502 ;
  assign n16124 = n4479 & n12383 ;
  assign n16125 = n16123 | n16124 ;
  assign n16126 = n16122 | n16125 ;
  assign n16127 = n4487 | n16126 ;
  assign n16128 = ( ~n12756 & n16126 ) | ( ~n12756 & n16127 ) | ( n16126 & n16127 ) ;
  assign n16129 = ~x26 & n16128 ;
  assign n16130 = x26 | n16129 ;
  assign n16131 = ( ~n16128 & n16129 ) | ( ~n16128 & n16130 ) | ( n16129 & n16130 ) ;
  assign n16132 = n16121 & n16131 ;
  assign n16133 = n16121 | n16131 ;
  assign n16134 = ~n16132 & n16133 ;
  assign n16135 = n4551 & n12375 ;
  assign n16136 = n4546 & n12378 ;
  assign n16137 = n4548 & ~n12371 ;
  assign n16138 = n16136 | n16137 ;
  assign n16139 = n16135 | n16138 ;
  assign n16140 = ( n4554 & n13064 ) | ( n4554 & ~n13065 ) | ( n13064 & ~n13065 ) ;
  assign n16141 = n16139 | n16140 ;
  assign n16142 = x23 | n16141 ;
  assign n16143 = ~x23 & n16142 ;
  assign n16144 = ( ~n16141 & n16142 ) | ( ~n16141 & n16143 ) | ( n16142 & n16143 ) ;
  assign n16146 = ( n16134 & n16144 ) | ( n16134 & n16145 ) | ( n16144 & n16145 ) ;
  assign n16147 = ( n16134 & n16144 ) | ( n16134 & ~n16146 ) | ( n16144 & ~n16146 ) ;
  assign n16148 = ( n16145 & ~n16146 ) | ( n16145 & n16147 ) | ( ~n16146 & n16147 ) ;
  assign n16149 = ( ~n16047 & n16107 ) | ( ~n16047 & n16148 ) | ( n16107 & n16148 ) ;
  assign n16150 = ( n16047 & ~n16148 ) | ( n16047 & n16149 ) | ( ~n16148 & n16149 ) ;
  assign n16151 = ( ~n16107 & n16149 ) | ( ~n16107 & n16150 ) | ( n16149 & n16150 ) ;
  assign n16152 = ( ~n16050 & n16097 ) | ( ~n16050 & n16151 ) | ( n16097 & n16151 ) ;
  assign n16153 = ( n16050 & ~n16151 ) | ( n16050 & n16152 ) | ( ~n16151 & n16152 ) ;
  assign n16154 = ( ~n16097 & n16152 ) | ( ~n16097 & n16153 ) | ( n16152 & n16153 ) ;
  assign n16155 = ( ~n16053 & n16087 ) | ( ~n16053 & n16154 ) | ( n16087 & n16154 ) ;
  assign n16156 = ( n16053 & ~n16154 ) | ( n16053 & n16155 ) | ( ~n16154 & n16155 ) ;
  assign n16157 = ( ~n16087 & n16155 ) | ( ~n16087 & n16156 ) | ( n16155 & n16156 ) ;
  assign n16158 = ( n16066 & n16076 ) | ( n16066 & n16157 ) | ( n16076 & n16157 ) ;
  assign n16159 = n7305 & ~n12335 ;
  assign n16160 = n7300 & ~n12586 ;
  assign n16161 = n7302 & n12580 ;
  assign n16162 = n16160 | n16161 ;
  assign n16163 = n16159 | n16162 ;
  assign n16164 = n7308 & n13587 ;
  assign n16165 = ( n7308 & n13585 ) | ( n7308 & n16164 ) | ( n13585 & n16164 ) ;
  assign n16166 = n16163 | n16165 ;
  assign n16167 = x11 | n16166 ;
  assign n16168 = ~x11 & n16167 ;
  assign n16169 = ( ~n16166 & n16167 ) | ( ~n16166 & n16168 ) | ( n16167 & n16168 ) ;
  assign n16170 = ( n16053 & n16087 ) | ( n16053 & n16154 ) | ( n16087 & n16154 ) ;
  assign n16171 = n7280 & ~n12344 ;
  assign n16172 = n5384 & n12553 ;
  assign n16173 = n7277 & n12340 ;
  assign n16174 = n16172 | n16173 ;
  assign n16175 = n16171 | n16174 ;
  assign n16176 = n39 | n16175 ;
  assign n16177 = ( ~n13523 & n16175 ) | ( ~n13523 & n16176 ) | ( n16175 & n16176 ) ;
  assign n16178 = ~x14 & n16177 ;
  assign n16179 = x14 | n16178 ;
  assign n16180 = ( ~n16177 & n16178 ) | ( ~n16177 & n16179 ) | ( n16178 & n16179 ) ;
  assign n16181 = ( n16050 & n16097 ) | ( n16050 & n16151 ) | ( n16097 & n16151 ) ;
  assign n16182 = n5083 & n12558 ;
  assign n16183 = n5069 & n12351 ;
  assign n16184 = n5070 & n12355 ;
  assign n16185 = n16183 | n16184 ;
  assign n16186 = n16182 | n16185 ;
  assign n16187 = n5074 | n16186 ;
  assign n16188 = ( n13330 & n16186 ) | ( n13330 & n16187 ) | ( n16186 & n16187 ) ;
  assign n16189 = x17 & n16188 ;
  assign n16190 = x17 & ~n16189 ;
  assign n16191 = ( n16188 & ~n16189 ) | ( n16188 & n16190 ) | ( ~n16189 & n16190 ) ;
  assign n16192 = n16118 | n16132 ;
  assign n16193 = ~n14394 & n14396 ;
  assign n16194 = n14397 | n16193 ;
  assign n16195 = n16192 & ~n16194 ;
  assign n16196 = ~n16192 & n16194 ;
  assign n16197 = n16195 | n16196 ;
  assign n16198 = n4551 & n12520 ;
  assign n16199 = n4546 & ~n12371 ;
  assign n16200 = n4548 & n12375 ;
  assign n16201 = n16199 | n16200 ;
  assign n16202 = n16198 | n16201 ;
  assign n16203 = n4554 & n12837 ;
  assign n16204 = ( n4554 & n12835 ) | ( n4554 & n16203 ) | ( n12835 & n16203 ) ;
  assign n16205 = n16202 | n16204 ;
  assign n16206 = x23 | n16205 ;
  assign n16207 = ~x23 & n16206 ;
  assign n16208 = ( ~n16205 & n16206 ) | ( ~n16205 & n16207 ) | ( n16206 & n16207 ) ;
  assign n16209 = ( n16146 & n16197 ) | ( n16146 & ~n16208 ) | ( n16197 & ~n16208 ) ;
  assign n16210 = ( ~n16197 & n16208 ) | ( ~n16197 & n16209 ) | ( n16208 & n16209 ) ;
  assign n16211 = ( ~n16146 & n16209 ) | ( ~n16146 & n16210 ) | ( n16209 & n16210 ) ;
  assign n16212 = n4781 & ~n12537 ;
  assign n16213 = n4776 & ~n12360 ;
  assign n16214 = n4778 & n12364 ;
  assign n16215 = n16213 | n16214 ;
  assign n16216 = n16212 | n16215 ;
  assign n16217 = ( n4784 & n13081 ) | ( n4784 & ~n13082 ) | ( n13081 & ~n13082 ) ;
  assign n16218 = n16216 | n16217 ;
  assign n16219 = x20 | n16218 ;
  assign n16220 = ~x20 & n16219 ;
  assign n16221 = ( ~n16218 & n16219 ) | ( ~n16218 & n16220 ) | ( n16219 & n16220 ) ;
  assign n16222 = n16211 | n16221 ;
  assign n16223 = ~n16221 & n16222 ;
  assign n16224 = ( ~n16211 & n16222 ) | ( ~n16211 & n16223 ) | ( n16222 & n16223 ) ;
  assign n16225 = ( n16047 & n16107 ) | ( n16047 & n16148 ) | ( n16107 & n16148 ) ;
  assign n16226 = ( n16191 & n16224 ) | ( n16191 & ~n16225 ) | ( n16224 & ~n16225 ) ;
  assign n16227 = ( ~n16224 & n16225 ) | ( ~n16224 & n16226 ) | ( n16225 & n16226 ) ;
  assign n16228 = ( ~n16191 & n16226 ) | ( ~n16191 & n16227 ) | ( n16226 & n16227 ) ;
  assign n16229 = ( n16180 & ~n16181 ) | ( n16180 & n16228 ) | ( ~n16181 & n16228 ) ;
  assign n16230 = ( n16181 & ~n16228 ) | ( n16181 & n16229 ) | ( ~n16228 & n16229 ) ;
  assign n16231 = ( ~n16180 & n16229 ) | ( ~n16180 & n16230 ) | ( n16229 & n16230 ) ;
  assign n16232 = ( n16169 & ~n16170 ) | ( n16169 & n16231 ) | ( ~n16170 & n16231 ) ;
  assign n16233 = ( n16170 & ~n16231 ) | ( n16170 & n16232 ) | ( ~n16231 & n16232 ) ;
  assign n16234 = ( ~n16169 & n16232 ) | ( ~n16169 & n16233 ) | ( n16232 & n16233 ) ;
  assign n16235 = n5512 & ~n12325 ;
  assign n16236 = n5508 & ~n12328 ;
  assign n16237 = n16235 | n16236 ;
  assign n16238 = n5503 & n12608 ;
  assign n16239 = n16237 | n16238 ;
  assign n16240 = n5515 & n13570 ;
  assign n16241 = ( n5515 & n13568 ) | ( n5515 & n16240 ) | ( n13568 & n16240 ) ;
  assign n16242 = n16239 | n16241 ;
  assign n16243 = x8 | n16242 ;
  assign n16244 = ~x8 & n16243 ;
  assign n16245 = ( ~n16242 & n16243 ) | ( ~n16242 & n16244 ) | ( n16243 & n16244 ) ;
  assign n16246 = ( ~n16158 & n16234 ) | ( ~n16158 & n16245 ) | ( n16234 & n16245 ) ;
  assign n16247 = ( n16158 & ~n16234 ) | ( n16158 & n16246 ) | ( ~n16234 & n16246 ) ;
  assign n16248 = n5503 & ~n12318 ;
  assign n16249 = n5512 & ~n12328 ;
  assign n16250 = n5508 & n12608 ;
  assign n16251 = n16249 | n16250 ;
  assign n16252 = n16248 | n16251 ;
  assign n16253 = n5515 | n16252 ;
  assign n16254 = ( n14320 & n16252 ) | ( n14320 & n16253 ) | ( n16252 & n16253 ) ;
  assign n16255 = x8 & n16254 ;
  assign n16256 = x8 & ~n16255 ;
  assign n16257 = ( n16254 & ~n16255 ) | ( n16254 & n16256 ) | ( ~n16255 & n16256 ) ;
  assign n16258 = n16247 & n16257 ;
  assign n16259 = n16247 & ~n16258 ;
  assign n16260 = n7305 & ~n12325 ;
  assign n16261 = n7300 & n12580 ;
  assign n16262 = n7302 & ~n12335 ;
  assign n16263 = n16261 | n16262 ;
  assign n16264 = n16260 | n16263 ;
  assign n16265 = n7308 | n16264 ;
  assign n16266 = ( ~n13720 & n16264 ) | ( ~n13720 & n16265 ) | ( n16264 & n16265 ) ;
  assign n16267 = ~x11 & n16266 ;
  assign n16268 = x11 | n16267 ;
  assign n16269 = ( ~n16266 & n16267 ) | ( ~n16266 & n16268 ) | ( n16267 & n16268 ) ;
  assign n16270 = n7280 & ~n12586 ;
  assign n16271 = n5384 & n12340 ;
  assign n16272 = n7277 & ~n12344 ;
  assign n16273 = n16271 | n16272 ;
  assign n16274 = n16270 | n16273 ;
  assign n16275 = ( n39 & n13454 ) | ( n39 & n13455 ) | ( n13454 & n13455 ) ;
  assign n16276 = n16274 | n16275 ;
  assign n16277 = x14 | n16276 ;
  assign n16278 = ~x14 & n16277 ;
  assign n16279 = ( ~n16276 & n16277 ) | ( ~n16276 & n16278 ) | ( n16277 & n16278 ) ;
  assign n16280 = ~n14398 & n14400 ;
  assign n16281 = n14401 | n16280 ;
  assign n16282 = n4551 & ~n12360 ;
  assign n16283 = n4546 & n12375 ;
  assign n16284 = n4548 & n12520 ;
  assign n16285 = n16283 | n16284 ;
  assign n16286 = n16282 | n16285 ;
  assign n16287 = n4554 | n16286 ;
  assign n16288 = ( ~n12902 & n16286 ) | ( ~n12902 & n16287 ) | ( n16286 & n16287 ) ;
  assign n16289 = ~x23 & n16288 ;
  assign n16290 = x23 | n16289 ;
  assign n16291 = ( ~n16288 & n16289 ) | ( ~n16288 & n16290 ) | ( n16289 & n16290 ) ;
  assign n16292 = ~n16281 & n16291 ;
  assign n16293 = n16281 | n16292 ;
  assign n16294 = n16281 & n16291 ;
  assign n16295 = ~n16197 & n16208 ;
  assign n16296 = n16195 | n16295 ;
  assign n16297 = n16294 | n16296 ;
  assign n16298 = n16293 & ~n16297 ;
  assign n16299 = ( ~n16293 & n16294 ) | ( ~n16293 & n16296 ) | ( n16294 & n16296 ) ;
  assign n16300 = n16298 | n16299 ;
  assign n16301 = n4781 & n12351 ;
  assign n16302 = n4776 & n12364 ;
  assign n16303 = n4778 & ~n12537 ;
  assign n16304 = n16302 | n16303 ;
  assign n16305 = n16301 | n16304 ;
  assign n16306 = n4784 & ~n12928 ;
  assign n16307 = ( n4784 & n12925 ) | ( n4784 & n16306 ) | ( n12925 & n16306 ) ;
  assign n16308 = n16305 | n16307 ;
  assign n16309 = x20 | n16308 ;
  assign n16310 = ~x20 & n16309 ;
  assign n16311 = ( ~n16308 & n16309 ) | ( ~n16308 & n16310 ) | ( n16309 & n16310 ) ;
  assign n16312 = ~n16300 & n16311 ;
  assign n16313 = n16300 | n16312 ;
  assign n16314 = n16300 & n16311 ;
  assign n16315 = ( n16146 & n16221 ) | ( n16146 & n16224 ) | ( n16221 & n16224 ) ;
  assign n16316 = n16314 | n16315 ;
  assign n16317 = n16313 & ~n16316 ;
  assign n16318 = ( ~n16313 & n16314 ) | ( ~n16313 & n16315 ) | ( n16314 & n16315 ) ;
  assign n16319 = n16317 | n16318 ;
  assign n16320 = n5083 & n12553 ;
  assign n16321 = n5069 & n12355 ;
  assign n16322 = n5070 & n12558 ;
  assign n16323 = n16321 | n16322 ;
  assign n16324 = n16320 | n16323 ;
  assign n16325 = n5074 | n16324 ;
  assign n16326 = ( n13097 & n16324 ) | ( n13097 & n16325 ) | ( n16324 & n16325 ) ;
  assign n16327 = x17 & n16326 ;
  assign n16328 = x17 & ~n16327 ;
  assign n16329 = ( n16326 & ~n16327 ) | ( n16326 & n16328 ) | ( ~n16327 & n16328 ) ;
  assign n16330 = ~n16319 & n16329 ;
  assign n16331 = n16319 | n16330 ;
  assign n16332 = n16319 & n16329 ;
  assign n16333 = n16227 | n16332 ;
  assign n16334 = n16331 & ~n16333 ;
  assign n16335 = ( n16227 & ~n16331 ) | ( n16227 & n16332 ) | ( ~n16331 & n16332 ) ;
  assign n16336 = n16334 | n16335 ;
  assign n16337 = n16279 & ~n16336 ;
  assign n16338 = n16336 | n16337 ;
  assign n16339 = ( ~n16279 & n16337 ) | ( ~n16279 & n16338 ) | ( n16337 & n16338 ) ;
  assign n16340 = n16230 & ~n16339 ;
  assign n16341 = ~n16230 & n16339 ;
  assign n16342 = n16340 | n16341 ;
  assign n16343 = n16269 & ~n16342 ;
  assign n16344 = n16342 | n16343 ;
  assign n16345 = ( ~n16269 & n16343 ) | ( ~n16269 & n16344 ) | ( n16343 & n16344 ) ;
  assign n16346 = n16233 & ~n16345 ;
  assign n16347 = ~n16233 & n16345 ;
  assign n16348 = n16346 | n16347 ;
  assign n16349 = ~n16247 & n16257 ;
  assign n16350 = ( n16259 & ~n16348 ) | ( n16259 & n16349 ) | ( ~n16348 & n16349 ) ;
  assign n16351 = n16348 & ~n16349 ;
  assign n16352 = ~n16259 & n16351 ;
  assign n16353 = n16350 | n16352 ;
  assign n16354 = ~n12314 & n12982 ;
  assign n16355 = ( ~n12318 & n12983 ) | ( ~n12318 & n16354 ) | ( n12983 & n16354 ) ;
  assign n16356 = n8685 | n16355 ;
  assign n16357 = n12615 & ~n16355 ;
  assign n16358 = ( n12314 & ~n12604 ) | ( n12314 & n16357 ) | ( ~n12604 & n16357 ) ;
  assign n16359 = n16356 & ~n16358 ;
  assign n16360 = x5 & ~n16359 ;
  assign n16361 = ~x5 & n16359 ;
  assign n16362 = n16360 | n16361 ;
  assign n16363 = ( ~n16064 & n16065 ) | ( ~n16064 & n16066 ) | ( n16065 & n16066 ) ;
  assign n16364 = n15991 | n15993 ;
  assign n16365 = ~n15994 & n16364 ;
  assign n16366 = n7280 & n12558 ;
  assign n16367 = n5384 & n12351 ;
  assign n16368 = n7277 & n12355 ;
  assign n16369 = n16367 | n16368 ;
  assign n16370 = n16366 | n16369 ;
  assign n16371 = n39 | n16370 ;
  assign n16372 = ( n13330 & n16370 ) | ( n13330 & n16371 ) | ( n16370 & n16371 ) ;
  assign n16373 = x14 & n16372 ;
  assign n16374 = x14 & ~n16373 ;
  assign n16375 = ( n16372 & ~n16373 ) | ( n16372 & n16374 ) | ( ~n16373 & n16374 ) ;
  assign n16376 = n16365 & n16375 ;
  assign n16377 = n16365 | n16375 ;
  assign n16378 = ~n16376 & n16377 ;
  assign n16379 = n15987 | n15989 ;
  assign n16380 = ~n15990 & n16379 ;
  assign n16381 = n7280 & n12355 ;
  assign n16382 = n5384 & ~n12537 ;
  assign n16383 = n7277 & n12351 ;
  assign n16384 = n16382 | n16383 ;
  assign n16385 = n16381 | n16384 ;
  assign n16386 = n39 | n16385 ;
  assign n16387 = ( n13409 & n16385 ) | ( n13409 & n16386 ) | ( n16385 & n16386 ) ;
  assign n16388 = x14 & n16387 ;
  assign n16389 = x14 & ~n16388 ;
  assign n16390 = ( n16387 & ~n16388 ) | ( n16387 & n16389 ) | ( ~n16388 & n16389 ) ;
  assign n16391 = n15979 | n15981 ;
  assign n16392 = ~n15982 & n16391 ;
  assign n16393 = n7280 & ~n12537 ;
  assign n16394 = n5384 & ~n12360 ;
  assign n16395 = n7277 & n12364 ;
  assign n16396 = n16394 | n16395 ;
  assign n16397 = n16393 | n16396 ;
  assign n16398 = n39 & ~n13081 ;
  assign n16399 = n13082 & n16398 ;
  assign n16400 = ( n39 & n16397 ) | ( n39 & ~n16399 ) | ( n16397 & ~n16399 ) ;
  assign n16401 = x14 & n16400 ;
  assign n16402 = x14 & ~n16401 ;
  assign n16403 = ( n16400 & ~n16401 ) | ( n16400 & n16402 ) | ( ~n16401 & n16402 ) ;
  assign n16404 = n16392 & n16403 ;
  assign n16405 = n15646 | n15977 ;
  assign n16406 = ~n15978 & n16405 ;
  assign n16407 = n7280 & n12364 ;
  assign n16408 = n5384 & n12520 ;
  assign n16409 = n7277 & ~n12360 ;
  assign n16410 = n16408 | n16409 ;
  assign n16411 = n16407 | n16410 ;
  assign n16412 = n39 | n16411 ;
  assign n16413 = ( ~n13113 & n16411 ) | ( ~n13113 & n16412 ) | ( n16411 & n16412 ) ;
  assign n16414 = ~x14 & n16413 ;
  assign n16415 = x14 | n16414 ;
  assign n16416 = ( ~n16413 & n16414 ) | ( ~n16413 & n16415 ) | ( n16414 & n16415 ) ;
  assign n16417 = n16406 & n16416 ;
  assign n16418 = n16406 & ~n16417 ;
  assign n16419 = ~n16406 & n16416 ;
  assign n16420 = n16418 | n16419 ;
  assign n16421 = n7280 & ~n12360 ;
  assign n16422 = n5384 & n12375 ;
  assign n16423 = n7277 & n12520 ;
  assign n16424 = n16422 | n16423 ;
  assign n16425 = n16421 | n16424 ;
  assign n16426 = n39 | n16425 ;
  assign n16427 = ( ~n12902 & n16425 ) | ( ~n12902 & n16426 ) | ( n16425 & n16426 ) ;
  assign n16428 = ~x14 & n16427 ;
  assign n16429 = x14 | n16428 ;
  assign n16430 = ( ~n16427 & n16428 ) | ( ~n16427 & n16429 ) | ( n16428 & n16429 ) ;
  assign n16431 = ~n15973 & n15975 ;
  assign n16432 = n15976 | n16431 ;
  assign n16433 = n7280 & n12520 ;
  assign n16434 = n5384 & ~n12371 ;
  assign n16435 = n7277 & n12375 ;
  assign n16436 = n16434 | n16435 ;
  assign n16437 = n16433 | n16436 ;
  assign n16438 = n39 & ~n12837 ;
  assign n16439 = ~n12835 & n16438 ;
  assign n16440 = ( n39 & n16437 ) | ( n39 & ~n16439 ) | ( n16437 & ~n16439 ) ;
  assign n16441 = ~x14 & n16440 ;
  assign n16442 = x14 | n16441 ;
  assign n16443 = ( ~n16440 & n16441 ) | ( ~n16440 & n16442 ) | ( n16441 & n16442 ) ;
  assign n16444 = n15691 | n15967 ;
  assign n16445 = ~n15968 & n16444 ;
  assign n16446 = n7280 & n12375 ;
  assign n16447 = n5384 & n12378 ;
  assign n16448 = n7277 & ~n12371 ;
  assign n16449 = n16447 | n16448 ;
  assign n16450 = n16446 | n16449 ;
  assign n16451 = n39 & n13065 ;
  assign n16452 = ~n13064 & n16451 ;
  assign n16453 = ( n39 & n16450 ) | ( n39 & ~n16452 ) | ( n16450 & ~n16452 ) ;
  assign n16454 = x14 & n16453 ;
  assign n16455 = x14 & ~n16454 ;
  assign n16456 = ( n16453 & ~n16454 ) | ( n16453 & n16455 ) | ( ~n16454 & n16455 ) ;
  assign n16457 = n7280 & ~n12371 ;
  assign n16458 = n5384 & ~n12502 ;
  assign n16459 = n7277 & n12378 ;
  assign n16460 = n16458 | n16459 ;
  assign n16461 = n16457 | n16460 ;
  assign n16462 = n39 | n16461 ;
  assign n16463 = ( ~n12848 & n16461 ) | ( ~n12848 & n16462 ) | ( n16461 & n16462 ) ;
  assign n16464 = ~x14 & n16463 ;
  assign n16465 = x14 | n16464 ;
  assign n16466 = ( ~n16463 & n16464 ) | ( ~n16463 & n16465 ) | ( n16464 & n16465 ) ;
  assign n16467 = n7280 & n12378 ;
  assign n16468 = n5384 & n12387 ;
  assign n16469 = n7277 & ~n12502 ;
  assign n16470 = n16468 | n16469 ;
  assign n16471 = n16467 | n16470 ;
  assign n16472 = n39 | n16471 ;
  assign n16473 = ( ~n12816 & n16471 ) | ( ~n12816 & n16472 ) | ( n16471 & n16472 ) ;
  assign n16474 = ~x14 & n16473 ;
  assign n16475 = x14 | n16474 ;
  assign n16476 = ( ~n16473 & n16474 ) | ( ~n16473 & n16475 ) | ( n16474 & n16475 ) ;
  assign n16477 = n15745 | n15959 ;
  assign n16478 = n15957 | n16477 ;
  assign n16479 = ~n15960 & n16478 ;
  assign n16480 = n7280 & ~n12502 ;
  assign n16481 = n5384 & n12383 ;
  assign n16482 = n7277 & n12387 ;
  assign n16483 = n16481 | n16482 ;
  assign n16484 = n16480 | n16483 ;
  assign n16485 = n39 | n16484 ;
  assign n16486 = ( ~n12756 & n16484 ) | ( ~n12756 & n16485 ) | ( n16484 & n16485 ) ;
  assign n16487 = ~x14 & n16486 ;
  assign n16488 = x14 | n16487 ;
  assign n16489 = ( ~n16486 & n16487 ) | ( ~n16486 & n16488 ) | ( n16487 & n16488 ) ;
  assign n16490 = n16479 & n16489 ;
  assign n16491 = n15953 & ~n15957 ;
  assign n16492 = n15956 & ~n15957 ;
  assign n16493 = n16491 | n16492 ;
  assign n16494 = n7280 & n12387 ;
  assign n16495 = n5384 & n12392 ;
  assign n16496 = n7277 & n12383 ;
  assign n16497 = n16495 | n16496 ;
  assign n16498 = n16494 | n16497 ;
  assign n16499 = n39 | n16498 ;
  assign n16500 = ( n12948 & n16498 ) | ( n12948 & n16499 ) | ( n16498 & n16499 ) ;
  assign n16501 = x14 & n16500 ;
  assign n16502 = x14 & ~n16501 ;
  assign n16503 = ( n16500 & ~n16501 ) | ( n16500 & n16502 ) | ( ~n16501 & n16502 ) ;
  assign n16504 = n16493 & n16503 ;
  assign n16505 = n16493 & ~n16504 ;
  assign n16506 = ~n16493 & n16503 ;
  assign n16507 = n16505 | n16506 ;
  assign n16508 = n15760 | n15951 ;
  assign n16509 = ~n15952 & n16508 ;
  assign n16510 = n7280 & n12383 ;
  assign n16511 = n5384 & n12401 ;
  assign n16512 = n7277 & n12392 ;
  assign n16513 = n16511 | n16512 ;
  assign n16514 = n16510 | n16513 ;
  assign n16515 = n39 | n16514 ;
  assign n16516 = ( n13141 & n16514 ) | ( n13141 & n16515 ) | ( n16514 & n16515 ) ;
  assign n16517 = x14 & n16516 ;
  assign n16518 = x14 & ~n16517 ;
  assign n16519 = ( n16516 & ~n16517 ) | ( n16516 & n16518 ) | ( ~n16517 & n16518 ) ;
  assign n16520 = n16509 & n16519 ;
  assign n16521 = n15776 | n15949 ;
  assign n16522 = ~n15950 & n16521 ;
  assign n16523 = n7280 & n12392 ;
  assign n16524 = n5384 & n12415 ;
  assign n16525 = n7277 & n12401 ;
  assign n16526 = n16524 | n16525 ;
  assign n16527 = n16523 | n16526 ;
  assign n16528 = n39 | n16527 ;
  assign n16529 = ( n13034 & n16527 ) | ( n13034 & n16528 ) | ( n16527 & n16528 ) ;
  assign n16530 = x14 & n16529 ;
  assign n16531 = x14 & ~n16530 ;
  assign n16532 = ( n16529 & ~n16530 ) | ( n16529 & n16531 ) | ( ~n16530 & n16531 ) ;
  assign n16533 = n16522 & n16532 ;
  assign n16534 = n15791 | n15947 ;
  assign n16535 = ~n15948 & n16534 ;
  assign n16536 = n7280 & n12401 ;
  assign n16537 = n5384 & n12411 ;
  assign n16538 = n7277 & n12415 ;
  assign n16539 = n16537 | n16538 ;
  assign n16540 = n16536 | n16539 ;
  assign n16541 = n39 & ~n13163 ;
  assign n16542 = ~n13161 & n16541 ;
  assign n16543 = ( n39 & n16540 ) | ( n39 & ~n16542 ) | ( n16540 & ~n16542 ) ;
  assign n16544 = ~x14 & n16543 ;
  assign n16545 = x14 | n16544 ;
  assign n16546 = ( ~n16543 & n16544 ) | ( ~n16543 & n16545 ) | ( n16544 & n16545 ) ;
  assign n16547 = n16535 & n16546 ;
  assign n16548 = n15943 | n15945 ;
  assign n16549 = ~n15946 & n16548 ;
  assign n16550 = n7280 & n12415 ;
  assign n16551 = n5384 & n12419 ;
  assign n16552 = n7277 & n12411 ;
  assign n16553 = n16551 | n16552 ;
  assign n16554 = n16550 | n16553 ;
  assign n16555 = ( n39 & n13761 ) | ( n39 & n13762 ) | ( n13761 & n13762 ) ;
  assign n16556 = n16554 | n16555 ;
  assign n16557 = x14 | n16556 ;
  assign n16558 = ~x14 & n16557 ;
  assign n16559 = ( ~n16556 & n16557 ) | ( ~n16556 & n16558 ) | ( n16557 & n16558 ) ;
  assign n16560 = n16549 & n16559 ;
  assign n16561 = n16559 & ~n16560 ;
  assign n16562 = ( n16549 & ~n16560 ) | ( n16549 & n16561 ) | ( ~n16560 & n16561 ) ;
  assign n16563 = n7280 & n12411 ;
  assign n16564 = n5384 & ~n12423 ;
  assign n16565 = n7277 & n12419 ;
  assign n16566 = n16564 | n16565 ;
  assign n16567 = n16563 | n16566 ;
  assign n16568 = n39 | n16567 ;
  assign n16569 = ( n13776 & n16567 ) | ( n13776 & n16568 ) | ( n16567 & n16568 ) ;
  assign n16570 = x14 & n16569 ;
  assign n16571 = x14 & ~n16570 ;
  assign n16572 = ( n16569 & ~n16570 ) | ( n16569 & n16571 ) | ( ~n16570 & n16571 ) ;
  assign n16573 = n15820 & ~n15942 ;
  assign n16574 = ( n15941 & ~n15942 ) | ( n15941 & n16573 ) | ( ~n15942 & n16573 ) ;
  assign n16575 = n16572 & n16574 ;
  assign n16576 = n16574 & ~n16575 ;
  assign n16577 = n16572 & ~n16574 ;
  assign n16578 = n16576 | n16577 ;
  assign n16579 = n7280 & n12419 ;
  assign n16580 = n5384 & n12433 ;
  assign n16581 = n7277 & ~n12423 ;
  assign n16582 = n16580 | n16581 ;
  assign n16583 = n16579 | n16582 ;
  assign n16584 = n39 | n16583 ;
  assign n16585 = ( ~n13282 & n16583 ) | ( ~n13282 & n16584 ) | ( n16583 & n16584 ) ;
  assign n16586 = ~x14 & n16585 ;
  assign n16587 = x14 | n16586 ;
  assign n16588 = ( ~n16585 & n16586 ) | ( ~n16585 & n16587 ) | ( n16586 & n16587 ) ;
  assign n16589 = ( n15822 & n15940 ) | ( n15822 & ~n15941 ) | ( n15940 & ~n15941 ) ;
  assign n16590 = ( n15833 & ~n15941 ) | ( n15833 & n16589 ) | ( ~n15941 & n16589 ) ;
  assign n16591 = n16588 & n16590 ;
  assign n16592 = n16588 | n16590 ;
  assign n16593 = ~n16591 & n16592 ;
  assign n16594 = n15936 | n15938 ;
  assign n16595 = ~n15939 & n16594 ;
  assign n16596 = n7280 & ~n12423 ;
  assign n16597 = n5384 & ~n12438 ;
  assign n16598 = n7277 & n12433 ;
  assign n16599 = n16597 | n16598 ;
  assign n16600 = n16596 | n16599 ;
  assign n16601 = n39 | n16600 ;
  assign n16602 = ( ~n13786 & n16600 ) | ( ~n13786 & n16601 ) | ( n16600 & n16601 ) ;
  assign n16603 = ~x14 & n16602 ;
  assign n16604 = x14 | n16603 ;
  assign n16605 = ( ~n16602 & n16603 ) | ( ~n16602 & n16604 ) | ( n16603 & n16604 ) ;
  assign n16606 = n16595 & n16605 ;
  assign n16607 = n15861 | n15934 ;
  assign n16608 = ~n15935 & n16607 ;
  assign n16609 = n7280 & n12433 ;
  assign n16610 = n5384 & n12440 ;
  assign n16611 = n7277 & ~n12438 ;
  assign n16612 = n16610 | n16611 ;
  assign n16613 = n16609 | n16612 ;
  assign n16614 = n39 | n16613 ;
  assign n16615 = ( ~n14167 & n16613 ) | ( ~n14167 & n16614 ) | ( n16613 & n16614 ) ;
  assign n16616 = ~x14 & n16615 ;
  assign n16617 = x14 | n16616 ;
  assign n16618 = ( ~n16615 & n16616 ) | ( ~n16615 & n16617 ) | ( n16616 & n16617 ) ;
  assign n16619 = n16608 & n16618 ;
  assign n16620 = n16608 & ~n16619 ;
  assign n16621 = ~n16608 & n16618 ;
  assign n16622 = n16620 | n16621 ;
  assign n16623 = n15930 | n15932 ;
  assign n16624 = ~n15933 & n16623 ;
  assign n16625 = n7280 & ~n12438 ;
  assign n16626 = n5384 & n12446 ;
  assign n16627 = n7277 & n12440 ;
  assign n16628 = n16626 | n16627 ;
  assign n16629 = n16625 | n16628 ;
  assign n16630 = n39 & n14154 ;
  assign n16631 = ~n14156 & n16630 ;
  assign n16632 = ( n39 & n16629 ) | ( n39 & ~n16631 ) | ( n16629 & ~n16631 ) ;
  assign n16633 = x14 & n16632 ;
  assign n16634 = x14 & ~n16633 ;
  assign n16635 = ( n16632 & ~n16633 ) | ( n16632 & n16634 ) | ( ~n16633 & n16634 ) ;
  assign n16636 = n15889 | n15928 ;
  assign n16637 = ~n15929 & n16636 ;
  assign n16638 = n7280 & n12440 ;
  assign n16639 = n5384 & n12452 ;
  assign n16640 = n7277 & n12446 ;
  assign n16641 = n16639 | n16640 ;
  assign n16642 = n16638 | n16641 ;
  assign n16643 = n39 | n16642 ;
  assign n16644 = ( n13822 & n16642 ) | ( n13822 & n16643 ) | ( n16642 & n16643 ) ;
  assign n16645 = x14 & n16644 ;
  assign n16646 = x14 & ~n16645 ;
  assign n16647 = ( n16644 & ~n16645 ) | ( n16644 & n16646 ) | ( ~n16645 & n16646 ) ;
  assign n16648 = n16637 & n16647 ;
  assign n16649 = n7280 & n12446 ;
  assign n16650 = n5384 & n12454 ;
  assign n16651 = n7277 & n12452 ;
  assign n16652 = n16650 | n16651 ;
  assign n16653 = n16649 | n16652 ;
  assign n16654 = n39 | n16653 ;
  assign n16655 = ( n13862 & n16653 ) | ( n13862 & n16654 ) | ( n16653 & n16654 ) ;
  assign n16656 = x14 & n16655 ;
  assign n16657 = x14 & ~n16656 ;
  assign n16658 = ( n16655 & ~n16656 ) | ( n16655 & n16657 ) | ( ~n16656 & n16657 ) ;
  assign n16659 = n15916 & ~n15927 ;
  assign n16660 = ( n15926 & ~n15927 ) | ( n15926 & n16659 ) | ( ~n15927 & n16659 ) ;
  assign n16661 = n16658 & n16660 ;
  assign n16662 = n16658 | n16660 ;
  assign n16663 = ~n16661 & n16662 ;
  assign n16664 = n7280 & n12452 ;
  assign n16665 = n5384 & ~n12456 ;
  assign n16666 = n7277 & n12454 ;
  assign n16667 = n16665 | n16666 ;
  assign n16668 = n16664 | n16667 ;
  assign n16669 = n39 | n16668 ;
  assign n16670 = ( ~n13922 & n16668 ) | ( ~n13922 & n16669 ) | ( n16668 & n16669 ) ;
  assign n16671 = ~x14 & n16670 ;
  assign n16672 = x14 & ~n16670 ;
  assign n16673 = n16671 | n16672 ;
  assign n16674 = n15900 | n15911 ;
  assign n16675 = ~n15914 & n16674 ;
  assign n16676 = n16673 & n16675 ;
  assign n16677 = n15891 | n15899 ;
  assign n16678 = ~n15900 & n16677 ;
  assign n16679 = n7280 & n12454 ;
  assign n16680 = n5384 & n12459 ;
  assign n16681 = n7277 & ~n12456 ;
  assign n16682 = n16680 | n16681 ;
  assign n16683 = n16679 | n16682 ;
  assign n16684 = n39 | n16683 ;
  assign n16685 = ( n14041 & n16683 ) | ( n14041 & n16684 ) | ( n16683 & n16684 ) ;
  assign n16686 = x14 & n16685 ;
  assign n16687 = x14 & ~n16686 ;
  assign n16688 = ( n16685 & ~n16686 ) | ( n16685 & n16687 ) | ( ~n16686 & n16687 ) ;
  assign n16689 = n16678 & n16688 ;
  assign n16690 = n16678 | n16688 ;
  assign n16691 = ~n16689 & n16690 ;
  assign n16692 = x14 & ~n35 ;
  assign n16693 = ( x14 & n12468 ) | ( x14 & n16692 ) | ( n12468 & n16692 ) ;
  assign n16694 = n39 & n13994 ;
  assign n16695 = n7277 & ~n12468 ;
  assign n16696 = n7280 & ~n12466 ;
  assign n16697 = n16695 | n16696 ;
  assign n16698 = n16694 | n16697 ;
  assign n16699 = x14 | n16698 ;
  assign n16700 = ~x14 & n16699 ;
  assign n16701 = ( ~n16698 & n16699 ) | ( ~n16698 & n16700 ) | ( n16699 & n16700 ) ;
  assign n16702 = n16693 & n16701 ;
  assign n16703 = n5064 & ~n12468 ;
  assign n16704 = n7280 & n12459 ;
  assign n16705 = n5384 & ~n12468 ;
  assign n16706 = n7277 & ~n12466 ;
  assign n16707 = n16705 | n16706 ;
  assign n16708 = n16704 | n16707 ;
  assign n16709 = n39 & n14003 ;
  assign n16710 = n16708 | n16709 ;
  assign n16711 = ~x14 & n16710 ;
  assign n16712 = x14 | n16711 ;
  assign n16713 = ( ~n16710 & n16711 ) | ( ~n16710 & n16712 ) | ( n16711 & n16712 ) ;
  assign n16714 = n16703 & n16713 ;
  assign n16715 = n16702 & n16714 ;
  assign n16716 = n16702 & n16713 ;
  assign n16717 = n16703 | n16716 ;
  assign n16718 = ~n16715 & n16717 ;
  assign n16719 = n7280 & ~n12456 ;
  assign n16720 = n5384 & ~n12466 ;
  assign n16721 = n7277 & n12459 ;
  assign n16722 = n16720 | n16721 ;
  assign n16723 = n16719 | n16722 ;
  assign n16724 = ( n39 & n14031 ) | ( n39 & n16723 ) | ( n14031 & n16723 ) ;
  assign n16725 = ( x14 & ~n16723 ) | ( x14 & n16724 ) | ( ~n16723 & n16724 ) ;
  assign n16726 = ~n16724 & n16725 ;
  assign n16727 = n16723 | n16725 ;
  assign n16728 = ( ~x14 & n16726 ) | ( ~x14 & n16727 ) | ( n16726 & n16727 ) ;
  assign n16729 = n16718 & n16728 ;
  assign n16730 = n16715 | n16729 ;
  assign n16731 = n16691 & n16730 ;
  assign n16732 = n16689 | n16731 ;
  assign n16733 = n16673 | n16675 ;
  assign n16734 = ~n16676 & n16733 ;
  assign n16735 = n16732 & n16734 ;
  assign n16736 = n16676 | n16735 ;
  assign n16737 = n16663 & n16736 ;
  assign n16738 = n16661 | n16737 ;
  assign n16739 = n16647 & ~n16648 ;
  assign n16740 = ( n16637 & ~n16648 ) | ( n16637 & n16739 ) | ( ~n16648 & n16739 ) ;
  assign n16741 = n16738 & n16740 ;
  assign n16742 = n16648 | n16741 ;
  assign n16743 = ( n16624 & n16635 ) | ( n16624 & n16742 ) | ( n16635 & n16742 ) ;
  assign n16744 = n16622 & n16743 ;
  assign n16745 = n16619 | n16744 ;
  assign n16746 = n16595 | n16605 ;
  assign n16747 = ~n16606 & n16746 ;
  assign n16748 = n16745 & n16747 ;
  assign n16749 = n16606 | n16748 ;
  assign n16750 = n16593 & n16749 ;
  assign n16751 = n16591 | n16750 ;
  assign n16752 = n16578 & n16751 ;
  assign n16753 = n16575 | n16752 ;
  assign n16754 = n16562 & n16753 ;
  assign n16755 = n16560 | n16754 ;
  assign n16756 = n16535 & ~n16547 ;
  assign n16757 = ~n16535 & n16546 ;
  assign n16758 = n16756 | n16757 ;
  assign n16759 = n16755 & n16758 ;
  assign n16760 = n16547 | n16759 ;
  assign n16761 = n16522 & ~n16533 ;
  assign n16762 = ~n16522 & n16532 ;
  assign n16763 = n16761 | n16762 ;
  assign n16764 = n16760 & n16763 ;
  assign n16765 = n16509 | n16519 ;
  assign n16766 = ~n16520 & n16765 ;
  assign n16767 = ( n16533 & n16764 ) | ( n16533 & n16766 ) | ( n16764 & n16766 ) ;
  assign n16768 = n16520 | n16767 ;
  assign n16769 = n16507 & n16768 ;
  assign n16770 = n16504 | n16769 ;
  assign n16771 = n16489 & ~n16490 ;
  assign n16772 = ( n16479 & ~n16490 ) | ( n16479 & n16771 ) | ( ~n16490 & n16771 ) ;
  assign n16773 = n16770 & n16772 ;
  assign n16774 = n16490 | n16773 ;
  assign n16775 = ~n15961 & n15963 ;
  assign n16776 = n15964 | n16775 ;
  assign n16777 = ( n16476 & ~n16774 ) | ( n16476 & n16776 ) | ( ~n16774 & n16776 ) ;
  assign n16778 = ( ~n16476 & n16774 ) | ( ~n16476 & n16777 ) | ( n16774 & n16777 ) ;
  assign n16779 = ( ~n16776 & n16777 ) | ( ~n16776 & n16778 ) | ( n16777 & n16778 ) ;
  assign n16780 = ( n16476 & n16774 ) | ( n16476 & n16779 ) | ( n16774 & n16779 ) ;
  assign n16781 = n15704 & ~n15965 ;
  assign n16782 = n15966 | n16781 ;
  assign n16783 = ( n16466 & n16780 ) | ( n16466 & ~n16782 ) | ( n16780 & ~n16782 ) ;
  assign n16784 = ( n16445 & n16456 ) | ( n16445 & n16783 ) | ( n16456 & n16783 ) ;
  assign n16785 = ~n15969 & n15971 ;
  assign n16786 = n15972 | n16785 ;
  assign n16787 = n16443 & ~n16786 ;
  assign n16788 = n16786 | n16787 ;
  assign n16789 = ( ~n16443 & n16787 ) | ( ~n16443 & n16788 ) | ( n16787 & n16788 ) ;
  assign n16790 = n16784 & n16789 ;
  assign n16791 = n16784 | n16789 ;
  assign n16792 = ~n16790 & n16791 ;
  assign n16793 = ( n16443 & n16784 ) | ( n16443 & n16792 ) | ( n16784 & n16792 ) ;
  assign n16794 = ( ~n16430 & n16432 ) | ( ~n16430 & n16793 ) | ( n16432 & n16793 ) ;
  assign n16795 = ( n16430 & ~n16432 ) | ( n16430 & n16794 ) | ( ~n16432 & n16794 ) ;
  assign n16796 = n16420 & n16795 ;
  assign n16797 = n16417 | n16796 ;
  assign n16798 = n16392 & ~n16404 ;
  assign n16799 = ~n16392 & n16403 ;
  assign n16800 = n16798 | n16799 ;
  assign n16801 = n16797 & n16800 ;
  assign n16802 = n16404 | n16801 ;
  assign n16803 = n15983 | n15985 ;
  assign n16804 = ~n15986 & n16803 ;
  assign n16805 = n7280 & n12351 ;
  assign n16806 = n5384 & n12364 ;
  assign n16807 = n7277 & ~n12537 ;
  assign n16808 = n16806 | n16807 ;
  assign n16809 = n16805 | n16808 ;
  assign n16810 = n39 & n12928 ;
  assign n16811 = ~n12925 & n16810 ;
  assign n16812 = ( n39 & n16809 ) | ( n39 & ~n16811 ) | ( n16809 & ~n16811 ) ;
  assign n16813 = x14 & n16812 ;
  assign n16814 = x14 & ~n16813 ;
  assign n16815 = ( n16812 & ~n16813 ) | ( n16812 & n16814 ) | ( ~n16813 & n16814 ) ;
  assign n16816 = ( n16802 & n16804 ) | ( n16802 & n16815 ) | ( n16804 & n16815 ) ;
  assign n16817 = ( n16380 & n16390 ) | ( n16380 & n16816 ) | ( n16390 & n16816 ) ;
  assign n16818 = n16378 & n16817 ;
  assign n16819 = n16376 | n16818 ;
  assign n16820 = n7305 & ~n12586 ;
  assign n16821 = n7300 & n12340 ;
  assign n16822 = n7302 & ~n12344 ;
  assign n16823 = n16821 | n16822 ;
  assign n16824 = n16820 | n16823 ;
  assign n16825 = ( n7308 & n13454 ) | ( n7308 & n13455 ) | ( n13454 & n13455 ) ;
  assign n16826 = n16824 | n16825 ;
  assign n16827 = x11 | n16826 ;
  assign n16828 = ~x11 & n16827 ;
  assign n16829 = ( ~n16826 & n16827 ) | ( ~n16826 & n16828 ) | ( n16827 & n16828 ) ;
  assign n16830 = ( n16363 & ~n16819 ) | ( n16363 & n16829 ) | ( ~n16819 & n16829 ) ;
  assign n16831 = ( ~n16363 & n16819 ) | ( ~n16363 & n16830 ) | ( n16819 & n16830 ) ;
  assign n16832 = n5503 & ~n12328 ;
  assign n16833 = n5512 & ~n12335 ;
  assign n16834 = n5508 & ~n12325 ;
  assign n16835 = n16833 | n16834 ;
  assign n16836 = n16832 | n16835 ;
  assign n16837 = n5515 | n16836 ;
  assign n16838 = ( ~n13544 & n16836 ) | ( ~n13544 & n16837 ) | ( n16836 & n16837 ) ;
  assign n16839 = ~x8 & n16838 ;
  assign n16840 = x8 | n16839 ;
  assign n16841 = ( ~n16838 & n16839 ) | ( ~n16838 & n16840 ) | ( n16839 & n16840 ) ;
  assign n16842 = ( ~n16066 & n16076 ) | ( ~n16066 & n16157 ) | ( n16076 & n16157 ) ;
  assign n16843 = ( n16066 & ~n16157 ) | ( n16066 & n16842 ) | ( ~n16157 & n16842 ) ;
  assign n16844 = ( ~n16076 & n16842 ) | ( ~n16076 & n16843 ) | ( n16842 & n16843 ) ;
  assign n16845 = ( n16831 & n16841 ) | ( n16831 & n16844 ) | ( n16841 & n16844 ) ;
  assign n16846 = n16362 & n16845 ;
  assign n16847 = ( ~n16245 & n16246 ) | ( ~n16245 & n16247 ) | ( n16246 & n16247 ) ;
  assign n16848 = n16362 | n16845 ;
  assign n16849 = ~n16846 & n16848 ;
  assign n16850 = ~n16847 & n16849 ;
  assign n16851 = n16846 | n16850 ;
  assign n16852 = ~n16353 & n16851 ;
  assign n16853 = n16353 & ~n16851 ;
  assign n16854 = n16852 | n16853 ;
  assign n16855 = n7305 & n12553 ;
  assign n16856 = n7300 & n12355 ;
  assign n16857 = n7302 & n12558 ;
  assign n16858 = n16856 | n16857 ;
  assign n16859 = n16855 | n16858 ;
  assign n16860 = n7308 | n16859 ;
  assign n16861 = ( n13097 & n16859 ) | ( n13097 & n16860 ) | ( n16859 & n16860 ) ;
  assign n16862 = x11 & n16861 ;
  assign n16863 = x11 & ~n16862 ;
  assign n16864 = ( n16861 & ~n16862 ) | ( n16861 & n16863 ) | ( ~n16862 & n16863 ) ;
  assign n16865 = ( n16802 & ~n16804 ) | ( n16802 & n16815 ) | ( ~n16804 & n16815 ) ;
  assign n16866 = ( ~n16802 & n16804 ) | ( ~n16802 & n16865 ) | ( n16804 & n16865 ) ;
  assign n16867 = ( ~n16815 & n16865 ) | ( ~n16815 & n16866 ) | ( n16865 & n16866 ) ;
  assign n16868 = n16864 & n16867 ;
  assign n16869 = n16864 | n16867 ;
  assign n16870 = ~n16868 & n16869 ;
  assign n16871 = n16797 & ~n16801 ;
  assign n16872 = n16800 & ~n16801 ;
  assign n16873 = n16871 | n16872 ;
  assign n16874 = n7305 & n12558 ;
  assign n16875 = n7300 & n12351 ;
  assign n16876 = n7302 & n12355 ;
  assign n16877 = n16875 | n16876 ;
  assign n16878 = n16874 | n16877 ;
  assign n16879 = n7308 | n16878 ;
  assign n16880 = ( n13330 & n16878 ) | ( n13330 & n16879 ) | ( n16878 & n16879 ) ;
  assign n16881 = x11 & n16880 ;
  assign n16882 = x11 & ~n16881 ;
  assign n16883 = ( n16880 & ~n16881 ) | ( n16880 & n16882 ) | ( ~n16881 & n16882 ) ;
  assign n16884 = n16873 & n16883 ;
  assign n16885 = n16873 & ~n16884 ;
  assign n16886 = ~n16873 & n16883 ;
  assign n16887 = n16885 | n16886 ;
  assign n16888 = n16795 & ~n16796 ;
  assign n16889 = n16420 & ~n16796 ;
  assign n16890 = n16888 | n16889 ;
  assign n16891 = n7305 & n12355 ;
  assign n16892 = n7300 & ~n12537 ;
  assign n16893 = n7302 & n12351 ;
  assign n16894 = n16892 | n16893 ;
  assign n16895 = n16891 | n16894 ;
  assign n16896 = n7308 | n16895 ;
  assign n16897 = ( n13409 & n16895 ) | ( n13409 & n16896 ) | ( n16895 & n16896 ) ;
  assign n16898 = x11 & n16897 ;
  assign n16899 = x11 & ~n16898 ;
  assign n16900 = ( n16897 & ~n16898 ) | ( n16897 & n16899 ) | ( ~n16898 & n16899 ) ;
  assign n16901 = n16890 & n16900 ;
  assign n16902 = n16890 & ~n16901 ;
  assign n16903 = ~n16890 & n16900 ;
  assign n16904 = n16902 | n16903 ;
  assign n16905 = ( ~n16793 & n16794 ) | ( ~n16793 & n16795 ) | ( n16794 & n16795 ) ;
  assign n16906 = n7305 & n12351 ;
  assign n16907 = n7300 & n12364 ;
  assign n16908 = n7302 & ~n12537 ;
  assign n16909 = n16907 | n16908 ;
  assign n16910 = n16906 | n16909 ;
  assign n16911 = n7308 & ~n12928 ;
  assign n16912 = ( n7308 & n12925 ) | ( n7308 & n16911 ) | ( n12925 & n16911 ) ;
  assign n16913 = n16910 | n16912 ;
  assign n16914 = x11 | n16913 ;
  assign n16915 = ~x11 & n16914 ;
  assign n16916 = ( ~n16913 & n16914 ) | ( ~n16913 & n16915 ) | ( n16914 & n16915 ) ;
  assign n16917 = ~n16905 & n16916 ;
  assign n16918 = n16905 & ~n16916 ;
  assign n16919 = n16917 | n16918 ;
  assign n16920 = n7305 & ~n12537 ;
  assign n16921 = n7300 & ~n12360 ;
  assign n16922 = n7302 & n12364 ;
  assign n16923 = n16921 | n16922 ;
  assign n16924 = n16920 | n16923 ;
  assign n16925 = ( n7308 & n13081 ) | ( n7308 & ~n13082 ) | ( n13081 & ~n13082 ) ;
  assign n16926 = n16924 | n16925 ;
  assign n16927 = x11 | n16926 ;
  assign n16928 = ~x11 & n16927 ;
  assign n16929 = ( ~n16926 & n16927 ) | ( ~n16926 & n16928 ) | ( n16927 & n16928 ) ;
  assign n16930 = ~n16792 & n16929 ;
  assign n16931 = n16792 & ~n16929 ;
  assign n16932 = n16930 | n16931 ;
  assign n16933 = n7305 & n12364 ;
  assign n16934 = n7300 & n12520 ;
  assign n16935 = n7302 & ~n12360 ;
  assign n16936 = n16934 | n16935 ;
  assign n16937 = n16933 | n16936 ;
  assign n16938 = n7308 | n16937 ;
  assign n16939 = ( ~n13113 & n16937 ) | ( ~n13113 & n16938 ) | ( n16937 & n16938 ) ;
  assign n16940 = ~x11 & n16939 ;
  assign n16941 = x11 | n16940 ;
  assign n16942 = ( ~n16939 & n16940 ) | ( ~n16939 & n16941 ) | ( n16940 & n16941 ) ;
  assign n16943 = ( n16445 & n16783 ) | ( n16445 & ~n16784 ) | ( n16783 & ~n16784 ) ;
  assign n16944 = ( n16456 & ~n16784 ) | ( n16456 & n16943 ) | ( ~n16784 & n16943 ) ;
  assign n16945 = n16942 & n16944 ;
  assign n16946 = n16942 | n16944 ;
  assign n16947 = ~n16945 & n16946 ;
  assign n16948 = ( ~n16466 & n16782 ) | ( ~n16466 & n16783 ) | ( n16782 & n16783 ) ;
  assign n16949 = ( ~n16780 & n16783 ) | ( ~n16780 & n16948 ) | ( n16783 & n16948 ) ;
  assign n16950 = n7305 & ~n12360 ;
  assign n16951 = n7300 & n12375 ;
  assign n16952 = n7302 & n12520 ;
  assign n16953 = n16951 | n16952 ;
  assign n16954 = n16950 | n16953 ;
  assign n16955 = n7308 | n16954 ;
  assign n16956 = ( ~n12902 & n16954 ) | ( ~n12902 & n16955 ) | ( n16954 & n16955 ) ;
  assign n16957 = ~x11 & n16956 ;
  assign n16958 = x11 | n16957 ;
  assign n16959 = ( ~n16956 & n16957 ) | ( ~n16956 & n16958 ) | ( n16957 & n16958 ) ;
  assign n16960 = ~n16949 & n16959 ;
  assign n16961 = n16949 & ~n16959 ;
  assign n16962 = n16960 | n16961 ;
  assign n16963 = n7305 & n12520 ;
  assign n16964 = n7300 & ~n12371 ;
  assign n16965 = n7302 & n12375 ;
  assign n16966 = n16964 | n16965 ;
  assign n16967 = n16963 | n16966 ;
  assign n16968 = n7308 & n12837 ;
  assign n16969 = ( n7308 & n12835 ) | ( n7308 & n16968 ) | ( n12835 & n16968 ) ;
  assign n16970 = n16967 | n16969 ;
  assign n16971 = x11 | n16970 ;
  assign n16972 = ~x11 & n16971 ;
  assign n16973 = ( ~n16970 & n16971 ) | ( ~n16970 & n16972 ) | ( n16971 & n16972 ) ;
  assign n16974 = ~n16779 & n16973 ;
  assign n16975 = n16779 & ~n16973 ;
  assign n16976 = n16974 | n16975 ;
  assign n16977 = n16770 | n16772 ;
  assign n16978 = ~n16773 & n16977 ;
  assign n16979 = n7305 & n12375 ;
  assign n16980 = n7300 & n12378 ;
  assign n16981 = n7302 & ~n12371 ;
  assign n16982 = n16980 | n16981 ;
  assign n16983 = n16979 | n16982 ;
  assign n16984 = n7308 & n13065 ;
  assign n16985 = ~n13064 & n16984 ;
  assign n16986 = ( n7308 & n16983 ) | ( n7308 & ~n16985 ) | ( n16983 & ~n16985 ) ;
  assign n16987 = x11 & n16986 ;
  assign n16988 = x11 & ~n16987 ;
  assign n16989 = ( n16986 & ~n16987 ) | ( n16986 & n16988 ) | ( ~n16987 & n16988 ) ;
  assign n16990 = n16978 & n16989 ;
  assign n16991 = n16978 | n16989 ;
  assign n16992 = ~n16990 & n16991 ;
  assign n16993 = n16507 | n16768 ;
  assign n16994 = ~n16769 & n16993 ;
  assign n16995 = n7305 & ~n12371 ;
  assign n16996 = n7300 & ~n12502 ;
  assign n16997 = n7302 & n12378 ;
  assign n16998 = n16996 | n16997 ;
  assign n16999 = n16995 | n16998 ;
  assign n17000 = n7308 | n16999 ;
  assign n17001 = ( ~n12848 & n16999 ) | ( ~n12848 & n17000 ) | ( n16999 & n17000 ) ;
  assign n17002 = ~x11 & n17001 ;
  assign n17003 = x11 | n17002 ;
  assign n17004 = ( ~n17001 & n17002 ) | ( ~n17001 & n17003 ) | ( n17002 & n17003 ) ;
  assign n17005 = n16533 | n16766 ;
  assign n17006 = n16764 | n17005 ;
  assign n17007 = ~n16767 & n17006 ;
  assign n17008 = n7305 & n12378 ;
  assign n17009 = n7300 & n12387 ;
  assign n17010 = n7302 & ~n12502 ;
  assign n17011 = n17009 | n17010 ;
  assign n17012 = n17008 | n17011 ;
  assign n17013 = n7308 | n17012 ;
  assign n17014 = ( ~n12816 & n17012 ) | ( ~n12816 & n17013 ) | ( n17012 & n17013 ) ;
  assign n17015 = ~x11 & n17014 ;
  assign n17016 = x11 | n17015 ;
  assign n17017 = ( ~n17014 & n17015 ) | ( ~n17014 & n17016 ) | ( n17015 & n17016 ) ;
  assign n17018 = n17007 & n17017 ;
  assign n17019 = n16760 & ~n16764 ;
  assign n17020 = n16763 & ~n16764 ;
  assign n17021 = n17019 | n17020 ;
  assign n17022 = n7305 & ~n12502 ;
  assign n17023 = n7300 & n12383 ;
  assign n17024 = n7302 & n12387 ;
  assign n17025 = n17023 | n17024 ;
  assign n17026 = n17022 | n17025 ;
  assign n17027 = n7308 | n17026 ;
  assign n17028 = ( ~n12756 & n17026 ) | ( ~n12756 & n17027 ) | ( n17026 & n17027 ) ;
  assign n17029 = ~x11 & n17028 ;
  assign n17030 = x11 | n17029 ;
  assign n17031 = ( ~n17028 & n17029 ) | ( ~n17028 & n17030 ) | ( n17029 & n17030 ) ;
  assign n17032 = n17021 & n17031 ;
  assign n17033 = n17021 & ~n17032 ;
  assign n17034 = ~n17021 & n17031 ;
  assign n17035 = n17033 | n17034 ;
  assign n17036 = n16755 & ~n16759 ;
  assign n17037 = n16758 & ~n16759 ;
  assign n17038 = n17036 | n17037 ;
  assign n17039 = n7305 & n12387 ;
  assign n17040 = n7300 & n12392 ;
  assign n17041 = n7302 & n12383 ;
  assign n17042 = n17040 | n17041 ;
  assign n17043 = n17039 | n17042 ;
  assign n17044 = n7308 | n17043 ;
  assign n17045 = ( n12948 & n17043 ) | ( n12948 & n17044 ) | ( n17043 & n17044 ) ;
  assign n17046 = x11 & n17045 ;
  assign n17047 = x11 & ~n17046 ;
  assign n17048 = ( n17045 & ~n17046 ) | ( n17045 & n17047 ) | ( ~n17046 & n17047 ) ;
  assign n17049 = n17038 & n17048 ;
  assign n17050 = n17038 & ~n17049 ;
  assign n17051 = ~n17038 & n17048 ;
  assign n17052 = n17050 | n17051 ;
  assign n17053 = n16562 | n16753 ;
  assign n17054 = ~n16754 & n17053 ;
  assign n17055 = n7305 & n12383 ;
  assign n17056 = n7300 & n12401 ;
  assign n17057 = n7302 & n12392 ;
  assign n17058 = n17056 | n17057 ;
  assign n17059 = n17055 | n17058 ;
  assign n17060 = n7308 | n17059 ;
  assign n17061 = ( n13141 & n17059 ) | ( n13141 & n17060 ) | ( n17059 & n17060 ) ;
  assign n17062 = x11 & n17061 ;
  assign n17063 = x11 & ~n17062 ;
  assign n17064 = ( n17061 & ~n17062 ) | ( n17061 & n17063 ) | ( ~n17062 & n17063 ) ;
  assign n17065 = n17054 & n17064 ;
  assign n17066 = n16578 | n16751 ;
  assign n17067 = ~n16752 & n17066 ;
  assign n17068 = n7305 & n12392 ;
  assign n17069 = n7300 & n12415 ;
  assign n17070 = n7302 & n12401 ;
  assign n17071 = n17069 | n17070 ;
  assign n17072 = n17068 | n17071 ;
  assign n17073 = n7308 | n17072 ;
  assign n17074 = ( n13034 & n17072 ) | ( n13034 & n17073 ) | ( n17072 & n17073 ) ;
  assign n17075 = x11 & n17074 ;
  assign n17076 = x11 & ~n17075 ;
  assign n17077 = ( n17074 & ~n17075 ) | ( n17074 & n17076 ) | ( ~n17075 & n17076 ) ;
  assign n17078 = n17067 & n17077 ;
  assign n17079 = n16593 | n16749 ;
  assign n17080 = ~n16750 & n17079 ;
  assign n17081 = n7305 & n12401 ;
  assign n17082 = n7300 & n12411 ;
  assign n17083 = n7302 & n12415 ;
  assign n17084 = n17082 | n17083 ;
  assign n17085 = n17081 | n17084 ;
  assign n17086 = n7308 & ~n13163 ;
  assign n17087 = ~n13161 & n17086 ;
  assign n17088 = ( n7308 & n17085 ) | ( n7308 & ~n17087 ) | ( n17085 & ~n17087 ) ;
  assign n17089 = ~x11 & n17088 ;
  assign n17090 = x11 | n17089 ;
  assign n17091 = ( ~n17088 & n17089 ) | ( ~n17088 & n17090 ) | ( n17089 & n17090 ) ;
  assign n17092 = n17080 & n17091 ;
  assign n17093 = n16745 | n16747 ;
  assign n17094 = ~n16748 & n17093 ;
  assign n17095 = n7305 & n12415 ;
  assign n17096 = n7300 & n12419 ;
  assign n17097 = n7302 & n12411 ;
  assign n17098 = n17096 | n17097 ;
  assign n17099 = n17095 | n17098 ;
  assign n17100 = ( n7308 & n13761 ) | ( n7308 & n13762 ) | ( n13761 & n13762 ) ;
  assign n17101 = n17099 | n17100 ;
  assign n17102 = x11 | n17101 ;
  assign n17103 = ~x11 & n17102 ;
  assign n17104 = ( ~n17101 & n17102 ) | ( ~n17101 & n17103 ) | ( n17102 & n17103 ) ;
  assign n17105 = n17094 & n17104 ;
  assign n17106 = n17104 & ~n17105 ;
  assign n17107 = ( n17094 & ~n17105 ) | ( n17094 & n17106 ) | ( ~n17105 & n17106 ) ;
  assign n17108 = n7305 & n12411 ;
  assign n17109 = n7300 & ~n12423 ;
  assign n17110 = n7302 & n12419 ;
  assign n17111 = n17109 | n17110 ;
  assign n17112 = n17108 | n17111 ;
  assign n17113 = n7308 | n17112 ;
  assign n17114 = ( n13776 & n17112 ) | ( n13776 & n17113 ) | ( n17112 & n17113 ) ;
  assign n17115 = x11 & n17114 ;
  assign n17116 = x11 & ~n17115 ;
  assign n17117 = ( n17114 & ~n17115 ) | ( n17114 & n17116 ) | ( ~n17115 & n17116 ) ;
  assign n17118 = n16622 & ~n16744 ;
  assign n17119 = ( n16743 & ~n16744 ) | ( n16743 & n17118 ) | ( ~n16744 & n17118 ) ;
  assign n17120 = n17117 & n17119 ;
  assign n17121 = n17119 & ~n17120 ;
  assign n17122 = n17117 & ~n17119 ;
  assign n17123 = n17121 | n17122 ;
  assign n17124 = n7305 & n12419 ;
  assign n17125 = n7300 & n12433 ;
  assign n17126 = n7302 & ~n12423 ;
  assign n17127 = n17125 | n17126 ;
  assign n17128 = n17124 | n17127 ;
  assign n17129 = n7308 | n17128 ;
  assign n17130 = ( ~n13282 & n17128 ) | ( ~n13282 & n17129 ) | ( n17128 & n17129 ) ;
  assign n17131 = ~x11 & n17130 ;
  assign n17132 = x11 | n17131 ;
  assign n17133 = ( ~n17130 & n17131 ) | ( ~n17130 & n17132 ) | ( n17131 & n17132 ) ;
  assign n17134 = ( n16624 & n16742 ) | ( n16624 & ~n16743 ) | ( n16742 & ~n16743 ) ;
  assign n17135 = ( n16635 & ~n16743 ) | ( n16635 & n17134 ) | ( ~n16743 & n17134 ) ;
  assign n17136 = n17133 & n17135 ;
  assign n17137 = n17133 | n17135 ;
  assign n17138 = ~n17136 & n17137 ;
  assign n17139 = n16738 | n16740 ;
  assign n17140 = ~n16741 & n17139 ;
  assign n17141 = n7305 & ~n12423 ;
  assign n17142 = n7300 & ~n12438 ;
  assign n17143 = n7302 & n12433 ;
  assign n17144 = n17142 | n17143 ;
  assign n17145 = n17141 | n17144 ;
  assign n17146 = n7308 | n17145 ;
  assign n17147 = ( ~n13786 & n17145 ) | ( ~n13786 & n17146 ) | ( n17145 & n17146 ) ;
  assign n17148 = ~x11 & n17147 ;
  assign n17149 = x11 | n17148 ;
  assign n17150 = ( ~n17147 & n17148 ) | ( ~n17147 & n17149 ) | ( n17148 & n17149 ) ;
  assign n17151 = n17140 & n17150 ;
  assign n17152 = n16663 | n16736 ;
  assign n17153 = ~n16737 & n17152 ;
  assign n17154 = n7305 & n12433 ;
  assign n17155 = n7300 & n12440 ;
  assign n17156 = n7302 & ~n12438 ;
  assign n17157 = n17155 | n17156 ;
  assign n17158 = n17154 | n17157 ;
  assign n17159 = n7308 | n17158 ;
  assign n17160 = ( ~n14167 & n17158 ) | ( ~n14167 & n17159 ) | ( n17158 & n17159 ) ;
  assign n17161 = ~x11 & n17160 ;
  assign n17162 = x11 | n17161 ;
  assign n17163 = ( ~n17160 & n17161 ) | ( ~n17160 & n17162 ) | ( n17161 & n17162 ) ;
  assign n17164 = n17153 & n17163 ;
  assign n17165 = n17153 & ~n17164 ;
  assign n17166 = ~n17153 & n17163 ;
  assign n17167 = n17165 | n17166 ;
  assign n17168 = n16732 | n16734 ;
  assign n17169 = ~n16735 & n17168 ;
  assign n17170 = n7305 & ~n12438 ;
  assign n17171 = n7300 & n12446 ;
  assign n17172 = n7302 & n12440 ;
  assign n17173 = n17171 | n17172 ;
  assign n17174 = n17170 | n17173 ;
  assign n17175 = n7308 & n14154 ;
  assign n17176 = ~n14156 & n17175 ;
  assign n17177 = ( n7308 & n17174 ) | ( n7308 & ~n17176 ) | ( n17174 & ~n17176 ) ;
  assign n17178 = x11 & n17177 ;
  assign n17179 = x11 & ~n17178 ;
  assign n17180 = ( n17177 & ~n17178 ) | ( n17177 & n17179 ) | ( ~n17178 & n17179 ) ;
  assign n17181 = n16691 | n16730 ;
  assign n17182 = ~n16731 & n17181 ;
  assign n17183 = n7305 & n12440 ;
  assign n17184 = n7300 & n12452 ;
  assign n17185 = n7302 & n12446 ;
  assign n17186 = n17184 | n17185 ;
  assign n17187 = n17183 | n17186 ;
  assign n17188 = n7308 | n17187 ;
  assign n17189 = ( n13822 & n17187 ) | ( n13822 & n17188 ) | ( n17187 & n17188 ) ;
  assign n17190 = x11 & n17189 ;
  assign n17191 = x11 & ~n17190 ;
  assign n17192 = ( n17189 & ~n17190 ) | ( n17189 & n17191 ) | ( ~n17190 & n17191 ) ;
  assign n17193 = n17182 & n17192 ;
  assign n17194 = n7305 & n12446 ;
  assign n17195 = n7300 & n12454 ;
  assign n17196 = n7302 & n12452 ;
  assign n17197 = n17195 | n17196 ;
  assign n17198 = n17194 | n17197 ;
  assign n17199 = n7308 | n17198 ;
  assign n17200 = ( n13862 & n17198 ) | ( n13862 & n17199 ) | ( n17198 & n17199 ) ;
  assign n17201 = x11 & n17200 ;
  assign n17202 = x11 & ~n17201 ;
  assign n17203 = ( n17200 & ~n17201 ) | ( n17200 & n17202 ) | ( ~n17201 & n17202 ) ;
  assign n17204 = n16718 & ~n16729 ;
  assign n17205 = ( n16728 & ~n16729 ) | ( n16728 & n17204 ) | ( ~n16729 & n17204 ) ;
  assign n17206 = n17203 & n17205 ;
  assign n17207 = n17203 | n17205 ;
  assign n17208 = ~n17206 & n17207 ;
  assign n17209 = n7305 & n12452 ;
  assign n17210 = n7300 & ~n12456 ;
  assign n17211 = n7302 & n12454 ;
  assign n17212 = n17210 | n17211 ;
  assign n17213 = n17209 | n17212 ;
  assign n17214 = n7308 | n17213 ;
  assign n17215 = ( ~n13922 & n17213 ) | ( ~n13922 & n17214 ) | ( n17213 & n17214 ) ;
  assign n17216 = ~x11 & n17215 ;
  assign n17217 = x11 & ~n17215 ;
  assign n17218 = n17216 | n17217 ;
  assign n17219 = n16702 | n16713 ;
  assign n17220 = ~n16716 & n17219 ;
  assign n17221 = n17218 & n17220 ;
  assign n17222 = n16693 | n16701 ;
  assign n17223 = ~n16702 & n17222 ;
  assign n17224 = n7305 & n12454 ;
  assign n17225 = n7300 & n12459 ;
  assign n17226 = n7302 & ~n12456 ;
  assign n17227 = n17225 | n17226 ;
  assign n17228 = n17224 | n17227 ;
  assign n17229 = n7308 | n17228 ;
  assign n17230 = ( n14041 & n17228 ) | ( n14041 & n17229 ) | ( n17228 & n17229 ) ;
  assign n17231 = x11 & n17230 ;
  assign n17232 = x11 & ~n17231 ;
  assign n17233 = ( n17230 & ~n17231 ) | ( n17230 & n17232 ) | ( ~n17231 & n17232 ) ;
  assign n17234 = n17223 & n17233 ;
  assign n17235 = n17223 | n17233 ;
  assign n17236 = ~n17234 & n17235 ;
  assign n17237 = x11 & ~n7298 ;
  assign n17238 = ( x11 & n12468 ) | ( x11 & n17237 ) | ( n12468 & n17237 ) ;
  assign n17239 = n7308 & n13994 ;
  assign n17240 = n7302 & ~n12468 ;
  assign n17241 = n7305 & ~n12466 ;
  assign n17242 = n17240 | n17241 ;
  assign n17243 = n17239 | n17242 ;
  assign n17244 = x11 | n17243 ;
  assign n17245 = ~x11 & n17244 ;
  assign n17246 = ( ~n17243 & n17244 ) | ( ~n17243 & n17245 ) | ( n17244 & n17245 ) ;
  assign n17247 = n17238 & n17246 ;
  assign n17248 = n35 & ~n12468 ;
  assign n17249 = n7305 & n12459 ;
  assign n17250 = n7300 & ~n12468 ;
  assign n17251 = n7302 & ~n12466 ;
  assign n17252 = n17250 | n17251 ;
  assign n17253 = n17249 | n17252 ;
  assign n17254 = n7308 & n14003 ;
  assign n17255 = n17253 | n17254 ;
  assign n17256 = ~x11 & n17255 ;
  assign n17257 = x11 | n17256 ;
  assign n17258 = ( ~n17255 & n17256 ) | ( ~n17255 & n17257 ) | ( n17256 & n17257 ) ;
  assign n17259 = n17248 & n17258 ;
  assign n17260 = n17247 & n17259 ;
  assign n17261 = n17247 & n17258 ;
  assign n17262 = n17248 | n17261 ;
  assign n17263 = ~n17260 & n17262 ;
  assign n17264 = n7305 & ~n12456 ;
  assign n17265 = n7300 & ~n12466 ;
  assign n17266 = n7302 & n12459 ;
  assign n17267 = n17265 | n17266 ;
  assign n17268 = n17264 | n17267 ;
  assign n17269 = ( n7308 & n14031 ) | ( n7308 & n17268 ) | ( n14031 & n17268 ) ;
  assign n17270 = ( x11 & ~n17268 ) | ( x11 & n17269 ) | ( ~n17268 & n17269 ) ;
  assign n17271 = ~n17269 & n17270 ;
  assign n17272 = n17268 | n17270 ;
  assign n17273 = ( ~x11 & n17271 ) | ( ~x11 & n17272 ) | ( n17271 & n17272 ) ;
  assign n17274 = n17263 & n17273 ;
  assign n17275 = n17260 | n17274 ;
  assign n17276 = n17236 & n17275 ;
  assign n17277 = n17234 | n17276 ;
  assign n17278 = n17218 | n17220 ;
  assign n17279 = ~n17221 & n17278 ;
  assign n17280 = n17277 & n17279 ;
  assign n17281 = n17221 | n17280 ;
  assign n17282 = n17208 & n17281 ;
  assign n17283 = n17206 | n17282 ;
  assign n17284 = n17192 & ~n17193 ;
  assign n17285 = ( n17182 & ~n17193 ) | ( n17182 & n17284 ) | ( ~n17193 & n17284 ) ;
  assign n17286 = n17283 & n17285 ;
  assign n17287 = n17193 | n17286 ;
  assign n17288 = ( n17169 & n17180 ) | ( n17169 & n17287 ) | ( n17180 & n17287 ) ;
  assign n17289 = n17167 & n17288 ;
  assign n17290 = n17164 | n17289 ;
  assign n17291 = n17140 | n17150 ;
  assign n17292 = ~n17151 & n17291 ;
  assign n17293 = n17290 & n17292 ;
  assign n17294 = n17151 | n17293 ;
  assign n17295 = n17138 & n17294 ;
  assign n17296 = n17136 | n17295 ;
  assign n17297 = n17123 & n17296 ;
  assign n17298 = n17120 | n17297 ;
  assign n17299 = n17107 & n17298 ;
  assign n17300 = n17105 | n17299 ;
  assign n17301 = n17080 & ~n17092 ;
  assign n17302 = ~n17080 & n17091 ;
  assign n17303 = n17301 | n17302 ;
  assign n17304 = n17300 & n17303 ;
  assign n17305 = n17092 | n17304 ;
  assign n17306 = n17067 & ~n17078 ;
  assign n17307 = ~n17067 & n17077 ;
  assign n17308 = n17306 | n17307 ;
  assign n17309 = n17305 & n17308 ;
  assign n17310 = n17054 | n17064 ;
  assign n17311 = ~n17065 & n17310 ;
  assign n17312 = ( n17078 & n17309 ) | ( n17078 & n17311 ) | ( n17309 & n17311 ) ;
  assign n17313 = n17065 | n17312 ;
  assign n17314 = n17052 & n17313 ;
  assign n17315 = n17049 | n17314 ;
  assign n17316 = n17035 & n17315 ;
  assign n17317 = n17032 | n17316 ;
  assign n17318 = n17017 & ~n17018 ;
  assign n17319 = ( n17007 & ~n17018 ) | ( n17007 & n17318 ) | ( ~n17018 & n17318 ) ;
  assign n17320 = n17317 & n17319 ;
  assign n17321 = n17018 | n17320 ;
  assign n17322 = ( n16994 & n17004 ) | ( n16994 & n17321 ) | ( n17004 & n17321 ) ;
  assign n17323 = n16992 & n17322 ;
  assign n17324 = n16990 | n17323 ;
  assign n17325 = ~n16976 & n17324 ;
  assign n17326 = n16974 | n17325 ;
  assign n17327 = ~n16962 & n17326 ;
  assign n17328 = n16960 | n17327 ;
  assign n17329 = n16947 & n17328 ;
  assign n17330 = n16945 | n17329 ;
  assign n17331 = ~n16932 & n17330 ;
  assign n17332 = n16930 | n17331 ;
  assign n17333 = ~n16919 & n17332 ;
  assign n17334 = n16917 | n17333 ;
  assign n17335 = n16904 & n17334 ;
  assign n17336 = n16901 | n17335 ;
  assign n17337 = n16887 & n17336 ;
  assign n17338 = n16884 | n17337 ;
  assign n17339 = n16870 & n17338 ;
  assign n17340 = n16868 | n17339 ;
  assign n17341 = n7305 & n12340 ;
  assign n17342 = n7300 & n12558 ;
  assign n17343 = n7302 & n12553 ;
  assign n17344 = n17342 | n17343 ;
  assign n17345 = n17341 | n17344 ;
  assign n17346 = n7308 & n13347 ;
  assign n17347 = ( n7308 & n13346 ) | ( n7308 & n17346 ) | ( n13346 & n17346 ) ;
  assign n17348 = n17345 | n17347 ;
  assign n17349 = x11 | n17348 ;
  assign n17350 = ~x11 & n17349 ;
  assign n17351 = ( ~n17348 & n17349 ) | ( ~n17348 & n17350 ) | ( n17349 & n17350 ) ;
  assign n17352 = ( n16380 & n16816 ) | ( n16380 & ~n16817 ) | ( n16816 & ~n16817 ) ;
  assign n17353 = ( n16390 & ~n16817 ) | ( n16390 & n17352 ) | ( ~n16817 & n17352 ) ;
  assign n17354 = n17351 & n17353 ;
  assign n17355 = n17351 | n17353 ;
  assign n17356 = ~n17354 & n17355 ;
  assign n17357 = n17340 & n17356 ;
  assign n17358 = n17340 | n17356 ;
  assign n17359 = ~n17357 & n17358 ;
  assign n17360 = n5503 & n12580 ;
  assign n17361 = n5512 & ~n12344 ;
  assign n17362 = n5508 & ~n12586 ;
  assign n17363 = n17361 | n17362 ;
  assign n17364 = n17360 | n17363 ;
  assign n17365 = n5515 | n17364 ;
  assign n17366 = ( n13432 & n17364 ) | ( n13432 & n17365 ) | ( n17364 & n17365 ) ;
  assign n17367 = x8 & n17366 ;
  assign n17368 = x8 & ~n17367 ;
  assign n17369 = ( n17366 & ~n17367 ) | ( n17366 & n17368 ) | ( ~n17367 & n17368 ) ;
  assign n17370 = n17359 & n17369 ;
  assign n17371 = n17359 & ~n17370 ;
  assign n17372 = ~n17359 & n17369 ;
  assign n17373 = n17371 | n17372 ;
  assign n17374 = n16887 | n17336 ;
  assign n17375 = ~n17337 & n17374 ;
  assign n17376 = n5503 & ~n12344 ;
  assign n17377 = n5512 & n12553 ;
  assign n17378 = n5508 & n12340 ;
  assign n17379 = n17377 | n17378 ;
  assign n17380 = n17376 | n17379 ;
  assign n17381 = n5515 | n17380 ;
  assign n17382 = ( ~n13523 & n17380 ) | ( ~n13523 & n17381 ) | ( n17380 & n17381 ) ;
  assign n17383 = ~x8 & n17382 ;
  assign n17384 = x8 | n17383 ;
  assign n17385 = ( ~n17382 & n17383 ) | ( ~n17382 & n17384 ) | ( n17383 & n17384 ) ;
  assign n17386 = n17375 & n17385 ;
  assign n17387 = n16904 | n17334 ;
  assign n17388 = ~n17335 & n17387 ;
  assign n17389 = n5503 & n12340 ;
  assign n17390 = n5512 & n12558 ;
  assign n17391 = n5508 & n12553 ;
  assign n17392 = n17390 | n17391 ;
  assign n17393 = n17389 | n17392 ;
  assign n17394 = n5515 & ~n13346 ;
  assign n17395 = ~n13347 & n17394 ;
  assign n17396 = ( n5515 & n17393 ) | ( n5515 & ~n17395 ) | ( n17393 & ~n17395 ) ;
  assign n17397 = ~x8 & n17396 ;
  assign n17398 = x8 | n17397 ;
  assign n17399 = ( ~n17396 & n17397 ) | ( ~n17396 & n17398 ) | ( n17397 & n17398 ) ;
  assign n17400 = n17388 & n17399 ;
  assign n17401 = n16919 & ~n17332 ;
  assign n17402 = n17333 | n17401 ;
  assign n17403 = n5503 & n12553 ;
  assign n17404 = n5512 & n12355 ;
  assign n17405 = n5508 & n12558 ;
  assign n17406 = n17404 | n17405 ;
  assign n17407 = n17403 | n17406 ;
  assign n17408 = n5515 | n17407 ;
  assign n17409 = ( n13097 & n17407 ) | ( n13097 & n17408 ) | ( n17407 & n17408 ) ;
  assign n17410 = x8 & n17409 ;
  assign n17411 = x8 & ~n17410 ;
  assign n17412 = ( n17409 & ~n17410 ) | ( n17409 & n17411 ) | ( ~n17410 & n17411 ) ;
  assign n17413 = ~n17402 & n17412 ;
  assign n17414 = n16932 & ~n17330 ;
  assign n17415 = n17331 | n17414 ;
  assign n17416 = n5503 & n12558 ;
  assign n17417 = n5512 & n12351 ;
  assign n17418 = n5508 & n12355 ;
  assign n17419 = n17417 | n17418 ;
  assign n17420 = n17416 | n17419 ;
  assign n17421 = n5515 | n17420 ;
  assign n17422 = ( n13330 & n17420 ) | ( n13330 & n17421 ) | ( n17420 & n17421 ) ;
  assign n17423 = x8 & n17422 ;
  assign n17424 = x8 & ~n17423 ;
  assign n17425 = ( n17422 & ~n17423 ) | ( n17422 & n17424 ) | ( ~n17423 & n17424 ) ;
  assign n17426 = ~n17415 & n17425 ;
  assign n17427 = n16947 | n17328 ;
  assign n17428 = ~n17329 & n17427 ;
  assign n17429 = n5503 & n12355 ;
  assign n17430 = n5512 & ~n12537 ;
  assign n17431 = n5508 & n12351 ;
  assign n17432 = n17430 | n17431 ;
  assign n17433 = n17429 | n17432 ;
  assign n17434 = n5515 | n17433 ;
  assign n17435 = ( n13409 & n17433 ) | ( n13409 & n17434 ) | ( n17433 & n17434 ) ;
  assign n17436 = x8 & n17435 ;
  assign n17437 = x8 & ~n17436 ;
  assign n17438 = ( n17435 & ~n17436 ) | ( n17435 & n17437 ) | ( ~n17436 & n17437 ) ;
  assign n17439 = n17428 & n17438 ;
  assign n17440 = n16962 & ~n17326 ;
  assign n17441 = n17327 | n17440 ;
  assign n17442 = n5503 & n12351 ;
  assign n17443 = n5512 & n12364 ;
  assign n17444 = n5508 & ~n12537 ;
  assign n17445 = n17443 | n17444 ;
  assign n17446 = n17442 | n17445 ;
  assign n17447 = n5515 & ~n12925 ;
  assign n17448 = n12928 & n17447 ;
  assign n17449 = ( n5515 & n17446 ) | ( n5515 & ~n17448 ) | ( n17446 & ~n17448 ) ;
  assign n17450 = x8 & n17449 ;
  assign n17451 = x8 & ~n17450 ;
  assign n17452 = ( n17449 & ~n17450 ) | ( n17449 & n17451 ) | ( ~n17450 & n17451 ) ;
  assign n17453 = ~n17441 & n17452 ;
  assign n17454 = n16976 & ~n17324 ;
  assign n17455 = n17325 | n17454 ;
  assign n17456 = n5503 & ~n12537 ;
  assign n17457 = n5512 & ~n12360 ;
  assign n17458 = n5508 & n12364 ;
  assign n17459 = n17457 | n17458 ;
  assign n17460 = n17456 | n17459 ;
  assign n17461 = n5515 & ~n13081 ;
  assign n17462 = n13082 & n17461 ;
  assign n17463 = ( n5515 & n17460 ) | ( n5515 & ~n17462 ) | ( n17460 & ~n17462 ) ;
  assign n17464 = x8 & n17463 ;
  assign n17465 = x8 & ~n17464 ;
  assign n17466 = ( n17463 & ~n17464 ) | ( n17463 & n17465 ) | ( ~n17464 & n17465 ) ;
  assign n17467 = ~n17455 & n17466 ;
  assign n17468 = n16992 | n17322 ;
  assign n17469 = ~n17323 & n17468 ;
  assign n17470 = n5503 & n12364 ;
  assign n17471 = n5512 & n12520 ;
  assign n17472 = n5508 & ~n12360 ;
  assign n17473 = n17471 | n17472 ;
  assign n17474 = n17470 | n17473 ;
  assign n17475 = n5515 | n17474 ;
  assign n17476 = ( ~n13113 & n17474 ) | ( ~n13113 & n17475 ) | ( n17474 & n17475 ) ;
  assign n17477 = ~x8 & n17476 ;
  assign n17478 = x8 | n17477 ;
  assign n17479 = ( ~n17476 & n17477 ) | ( ~n17476 & n17478 ) | ( n17477 & n17478 ) ;
  assign n17480 = n17469 & n17479 ;
  assign n17481 = n17479 & ~n17480 ;
  assign n17482 = ( n17469 & ~n17480 ) | ( n17469 & n17481 ) | ( ~n17480 & n17481 ) ;
  assign n17483 = n5503 & ~n12360 ;
  assign n17484 = n5512 & n12375 ;
  assign n17485 = n5508 & n12520 ;
  assign n17486 = n17484 | n17485 ;
  assign n17487 = n17483 | n17486 ;
  assign n17488 = n5515 | n17487 ;
  assign n17489 = ( ~n12902 & n17487 ) | ( ~n12902 & n17488 ) | ( n17487 & n17488 ) ;
  assign n17490 = ~x8 & n17489 ;
  assign n17491 = x8 | n17490 ;
  assign n17492 = ( ~n17489 & n17490 ) | ( ~n17489 & n17491 ) | ( n17490 & n17491 ) ;
  assign n17493 = ( n16994 & n17321 ) | ( n16994 & ~n17322 ) | ( n17321 & ~n17322 ) ;
  assign n17494 = ( n17004 & ~n17322 ) | ( n17004 & n17493 ) | ( ~n17322 & n17493 ) ;
  assign n17495 = n17492 & n17494 ;
  assign n17496 = n17492 | n17494 ;
  assign n17497 = ~n17495 & n17496 ;
  assign n17498 = n17317 | n17319 ;
  assign n17499 = ~n17320 & n17498 ;
  assign n17500 = n5503 & n12520 ;
  assign n17501 = n5512 & ~n12371 ;
  assign n17502 = n5508 & n12375 ;
  assign n17503 = n17501 | n17502 ;
  assign n17504 = n17500 | n17503 ;
  assign n17505 = n5515 & ~n12837 ;
  assign n17506 = ~n12835 & n17505 ;
  assign n17507 = ( n5515 & n17504 ) | ( n5515 & ~n17506 ) | ( n17504 & ~n17506 ) ;
  assign n17508 = ~x8 & n17507 ;
  assign n17509 = x8 | n17508 ;
  assign n17510 = ( ~n17507 & n17508 ) | ( ~n17507 & n17509 ) | ( n17508 & n17509 ) ;
  assign n17511 = n17499 & n17510 ;
  assign n17512 = n17499 | n17510 ;
  assign n17513 = ~n17511 & n17512 ;
  assign n17514 = n17035 | n17315 ;
  assign n17515 = ~n17316 & n17514 ;
  assign n17516 = n5503 & n12375 ;
  assign n17517 = n5512 & n12378 ;
  assign n17518 = n5508 & ~n12371 ;
  assign n17519 = n17517 | n17518 ;
  assign n17520 = n17516 | n17519 ;
  assign n17521 = n5515 & n13065 ;
  assign n17522 = ~n13064 & n17521 ;
  assign n17523 = ( n5515 & n17520 ) | ( n5515 & ~n17522 ) | ( n17520 & ~n17522 ) ;
  assign n17524 = x8 & n17523 ;
  assign n17525 = x8 & ~n17524 ;
  assign n17526 = ( n17523 & ~n17524 ) | ( n17523 & n17525 ) | ( ~n17524 & n17525 ) ;
  assign n17527 = n17052 | n17313 ;
  assign n17528 = ~n17314 & n17527 ;
  assign n17529 = n5503 & ~n12371 ;
  assign n17530 = n5512 & ~n12502 ;
  assign n17531 = n5508 & n12378 ;
  assign n17532 = n17530 | n17531 ;
  assign n17533 = n17529 | n17532 ;
  assign n17534 = n5515 | n17533 ;
  assign n17535 = ( ~n12848 & n17533 ) | ( ~n12848 & n17534 ) | ( n17533 & n17534 ) ;
  assign n17536 = ~x8 & n17535 ;
  assign n17537 = x8 | n17536 ;
  assign n17538 = ( ~n17535 & n17536 ) | ( ~n17535 & n17537 ) | ( n17536 & n17537 ) ;
  assign n17539 = n17078 | n17311 ;
  assign n17540 = n17309 | n17539 ;
  assign n17541 = ~n17312 & n17540 ;
  assign n17542 = n5503 & n12378 ;
  assign n17543 = n5512 & n12387 ;
  assign n17544 = n5508 & ~n12502 ;
  assign n17545 = n17543 | n17544 ;
  assign n17546 = n17542 | n17545 ;
  assign n17547 = n5515 | n17546 ;
  assign n17548 = ( ~n12816 & n17546 ) | ( ~n12816 & n17547 ) | ( n17546 & n17547 ) ;
  assign n17549 = ~x8 & n17548 ;
  assign n17550 = x8 | n17549 ;
  assign n17551 = ( ~n17548 & n17549 ) | ( ~n17548 & n17550 ) | ( n17549 & n17550 ) ;
  assign n17552 = n17541 & n17551 ;
  assign n17553 = n17305 & ~n17309 ;
  assign n17554 = n17308 & ~n17309 ;
  assign n17555 = n17553 | n17554 ;
  assign n17556 = n5503 & ~n12502 ;
  assign n17557 = n5512 & n12383 ;
  assign n17558 = n5508 & n12387 ;
  assign n17559 = n17557 | n17558 ;
  assign n17560 = n17556 | n17559 ;
  assign n17561 = n5515 | n17560 ;
  assign n17562 = ( ~n12756 & n17560 ) | ( ~n12756 & n17561 ) | ( n17560 & n17561 ) ;
  assign n17563 = ~x8 & n17562 ;
  assign n17564 = x8 | n17563 ;
  assign n17565 = ( ~n17562 & n17563 ) | ( ~n17562 & n17564 ) | ( n17563 & n17564 ) ;
  assign n17566 = n17555 & n17565 ;
  assign n17567 = n17555 & ~n17566 ;
  assign n17568 = ~n17555 & n17565 ;
  assign n17569 = n17567 | n17568 ;
  assign n17570 = n17300 & ~n17304 ;
  assign n17571 = n17303 & ~n17304 ;
  assign n17572 = n17570 | n17571 ;
  assign n17573 = n5503 & n12387 ;
  assign n17574 = n5512 & n12392 ;
  assign n17575 = n5508 & n12383 ;
  assign n17576 = n17574 | n17575 ;
  assign n17577 = n17573 | n17576 ;
  assign n17578 = n5515 | n17577 ;
  assign n17579 = ( n12948 & n17577 ) | ( n12948 & n17578 ) | ( n17577 & n17578 ) ;
  assign n17580 = x8 & n17579 ;
  assign n17581 = x8 & ~n17580 ;
  assign n17582 = ( n17579 & ~n17580 ) | ( n17579 & n17581 ) | ( ~n17580 & n17581 ) ;
  assign n17583 = n17572 & n17582 ;
  assign n17584 = n17572 & ~n17583 ;
  assign n17585 = ~n17572 & n17582 ;
  assign n17586 = n17584 | n17585 ;
  assign n17587 = n17107 | n17298 ;
  assign n17588 = ~n17299 & n17587 ;
  assign n17589 = n5503 & n12383 ;
  assign n17590 = n5512 & n12401 ;
  assign n17591 = n5508 & n12392 ;
  assign n17592 = n17590 | n17591 ;
  assign n17593 = n17589 | n17592 ;
  assign n17594 = n5515 | n17593 ;
  assign n17595 = ( n13141 & n17593 ) | ( n13141 & n17594 ) | ( n17593 & n17594 ) ;
  assign n17596 = x8 & n17595 ;
  assign n17597 = x8 & ~n17596 ;
  assign n17598 = ( n17595 & ~n17596 ) | ( n17595 & n17597 ) | ( ~n17596 & n17597 ) ;
  assign n17599 = n17588 & n17598 ;
  assign n17600 = n17123 | n17296 ;
  assign n17601 = ~n17297 & n17600 ;
  assign n17602 = n5503 & n12392 ;
  assign n17603 = n5512 & n12415 ;
  assign n17604 = n5508 & n12401 ;
  assign n17605 = n17603 | n17604 ;
  assign n17606 = n17602 | n17605 ;
  assign n17607 = n5515 | n17606 ;
  assign n17608 = ( n13034 & n17606 ) | ( n13034 & n17607 ) | ( n17606 & n17607 ) ;
  assign n17609 = x8 & n17608 ;
  assign n17610 = x8 & ~n17609 ;
  assign n17611 = ( n17608 & ~n17609 ) | ( n17608 & n17610 ) | ( ~n17609 & n17610 ) ;
  assign n17612 = n17601 & n17611 ;
  assign n17613 = n17138 | n17294 ;
  assign n17614 = ~n17295 & n17613 ;
  assign n17615 = n5503 & n12401 ;
  assign n17616 = n5512 & n12411 ;
  assign n17617 = n5508 & n12415 ;
  assign n17618 = n17616 | n17617 ;
  assign n17619 = n17615 | n17618 ;
  assign n17620 = n5515 & ~n13163 ;
  assign n17621 = ~n13161 & n17620 ;
  assign n17622 = ( n5515 & n17619 ) | ( n5515 & ~n17621 ) | ( n17619 & ~n17621 ) ;
  assign n17623 = ~x8 & n17622 ;
  assign n17624 = x8 | n17623 ;
  assign n17625 = ( ~n17622 & n17623 ) | ( ~n17622 & n17624 ) | ( n17623 & n17624 ) ;
  assign n17626 = n17614 & n17625 ;
  assign n17627 = n17290 | n17292 ;
  assign n17628 = ~n17293 & n17627 ;
  assign n17629 = n5503 & n12415 ;
  assign n17630 = n5512 & n12419 ;
  assign n17631 = n5508 & n12411 ;
  assign n17632 = n17630 | n17631 ;
  assign n17633 = n17629 | n17632 ;
  assign n17634 = ( n5515 & n13761 ) | ( n5515 & n13762 ) | ( n13761 & n13762 ) ;
  assign n17635 = n17633 | n17634 ;
  assign n17636 = x8 | n17635 ;
  assign n17637 = ~x8 & n17636 ;
  assign n17638 = ( ~n17635 & n17636 ) | ( ~n17635 & n17637 ) | ( n17636 & n17637 ) ;
  assign n17639 = n17628 & n17638 ;
  assign n17640 = n17638 & ~n17639 ;
  assign n17641 = ( n17628 & ~n17639 ) | ( n17628 & n17640 ) | ( ~n17639 & n17640 ) ;
  assign n17642 = n5503 & n12411 ;
  assign n17643 = n5512 & ~n12423 ;
  assign n17644 = n5508 & n12419 ;
  assign n17645 = n17643 | n17644 ;
  assign n17646 = n17642 | n17645 ;
  assign n17647 = n5515 | n17646 ;
  assign n17648 = ( n13776 & n17646 ) | ( n13776 & n17647 ) | ( n17646 & n17647 ) ;
  assign n17649 = x8 & n17648 ;
  assign n17650 = x8 & ~n17649 ;
  assign n17651 = ( n17648 & ~n17649 ) | ( n17648 & n17650 ) | ( ~n17649 & n17650 ) ;
  assign n17652 = n17167 & ~n17289 ;
  assign n17653 = ( n17288 & ~n17289 ) | ( n17288 & n17652 ) | ( ~n17289 & n17652 ) ;
  assign n17654 = n17651 & n17653 ;
  assign n17655 = n17653 & ~n17654 ;
  assign n17656 = n17651 & ~n17653 ;
  assign n17657 = n17655 | n17656 ;
  assign n17658 = n5503 & n12419 ;
  assign n17659 = n5512 & n12433 ;
  assign n17660 = n5508 & ~n12423 ;
  assign n17661 = n17659 | n17660 ;
  assign n17662 = n17658 | n17661 ;
  assign n17663 = n5515 | n17662 ;
  assign n17664 = ( ~n13282 & n17662 ) | ( ~n13282 & n17663 ) | ( n17662 & n17663 ) ;
  assign n17665 = ~x8 & n17664 ;
  assign n17666 = x8 | n17665 ;
  assign n17667 = ( ~n17664 & n17665 ) | ( ~n17664 & n17666 ) | ( n17665 & n17666 ) ;
  assign n17668 = ( n17169 & n17287 ) | ( n17169 & ~n17288 ) | ( n17287 & ~n17288 ) ;
  assign n17669 = ( n17180 & ~n17288 ) | ( n17180 & n17668 ) | ( ~n17288 & n17668 ) ;
  assign n17670 = n17667 & n17669 ;
  assign n17671 = n17667 | n17669 ;
  assign n17672 = ~n17670 & n17671 ;
  assign n17673 = n17283 | n17285 ;
  assign n17674 = ~n17286 & n17673 ;
  assign n17675 = n5503 & ~n12423 ;
  assign n17676 = n5512 & ~n12438 ;
  assign n17677 = n5508 & n12433 ;
  assign n17678 = n17676 | n17677 ;
  assign n17679 = n17675 | n17678 ;
  assign n17680 = n5515 | n17679 ;
  assign n17681 = ( ~n13786 & n17679 ) | ( ~n13786 & n17680 ) | ( n17679 & n17680 ) ;
  assign n17682 = ~x8 & n17681 ;
  assign n17683 = x8 | n17682 ;
  assign n17684 = ( ~n17681 & n17682 ) | ( ~n17681 & n17683 ) | ( n17682 & n17683 ) ;
  assign n17685 = n17674 & n17684 ;
  assign n17686 = n17208 | n17281 ;
  assign n17687 = ~n17282 & n17686 ;
  assign n17688 = n5503 & n12433 ;
  assign n17689 = n5512 & n12440 ;
  assign n17690 = n5508 & ~n12438 ;
  assign n17691 = n17689 | n17690 ;
  assign n17692 = n17688 | n17691 ;
  assign n17693 = n5515 | n17692 ;
  assign n17694 = ( ~n14167 & n17692 ) | ( ~n14167 & n17693 ) | ( n17692 & n17693 ) ;
  assign n17695 = ~x8 & n17694 ;
  assign n17696 = x8 | n17695 ;
  assign n17697 = ( ~n17694 & n17695 ) | ( ~n17694 & n17696 ) | ( n17695 & n17696 ) ;
  assign n17698 = n17687 & n17697 ;
  assign n17699 = n17687 & ~n17698 ;
  assign n17700 = ~n17687 & n17697 ;
  assign n17701 = n17699 | n17700 ;
  assign n17702 = n17277 | n17279 ;
  assign n17703 = ~n17280 & n17702 ;
  assign n17704 = n5503 & ~n12438 ;
  assign n17705 = n5512 & n12446 ;
  assign n17706 = n5508 & n12440 ;
  assign n17707 = n17705 | n17706 ;
  assign n17708 = n17704 | n17707 ;
  assign n17709 = n5515 & n14154 ;
  assign n17710 = ~n14156 & n17709 ;
  assign n17711 = ( n5515 & n17708 ) | ( n5515 & ~n17710 ) | ( n17708 & ~n17710 ) ;
  assign n17712 = x8 & n17711 ;
  assign n17713 = x8 & ~n17712 ;
  assign n17714 = ( n17711 & ~n17712 ) | ( n17711 & n17713 ) | ( ~n17712 & n17713 ) ;
  assign n17715 = n17236 | n17275 ;
  assign n17716 = ~n17276 & n17715 ;
  assign n17717 = n5503 & n12440 ;
  assign n17718 = n5512 & n12452 ;
  assign n17719 = n5508 & n12446 ;
  assign n17720 = n17718 | n17719 ;
  assign n17721 = n17717 | n17720 ;
  assign n17722 = n5515 | n17721 ;
  assign n17723 = ( n13822 & n17721 ) | ( n13822 & n17722 ) | ( n17721 & n17722 ) ;
  assign n17724 = x8 & n17723 ;
  assign n17725 = x8 & ~n17724 ;
  assign n17726 = ( n17723 & ~n17724 ) | ( n17723 & n17725 ) | ( ~n17724 & n17725 ) ;
  assign n17727 = n17716 & n17726 ;
  assign n17728 = n5503 & n12446 ;
  assign n17729 = n5512 & n12454 ;
  assign n17730 = n5508 & n12452 ;
  assign n17731 = n17729 | n17730 ;
  assign n17732 = n17728 | n17731 ;
  assign n17733 = n5515 | n17732 ;
  assign n17734 = ( n13862 & n17732 ) | ( n13862 & n17733 ) | ( n17732 & n17733 ) ;
  assign n17735 = x8 & n17734 ;
  assign n17736 = x8 & ~n17735 ;
  assign n17737 = ( n17734 & ~n17735 ) | ( n17734 & n17736 ) | ( ~n17735 & n17736 ) ;
  assign n17738 = n17263 & ~n17274 ;
  assign n17739 = ( n17273 & ~n17274 ) | ( n17273 & n17738 ) | ( ~n17274 & n17738 ) ;
  assign n17740 = n17737 & n17739 ;
  assign n17741 = n17737 | n17739 ;
  assign n17742 = ~n17740 & n17741 ;
  assign n17743 = n5503 & n12452 ;
  assign n17744 = n5512 & ~n12456 ;
  assign n17745 = n5508 & n12454 ;
  assign n17746 = n17744 | n17745 ;
  assign n17747 = n17743 | n17746 ;
  assign n17748 = n5515 | n17747 ;
  assign n17749 = ( ~n13922 & n17747 ) | ( ~n13922 & n17748 ) | ( n17747 & n17748 ) ;
  assign n17750 = ~x8 & n17749 ;
  assign n17751 = x8 & ~n17749 ;
  assign n17752 = n17750 | n17751 ;
  assign n17753 = n17247 | n17258 ;
  assign n17754 = ~n17261 & n17753 ;
  assign n17755 = n17752 & n17754 ;
  assign n17756 = n17238 | n17246 ;
  assign n17757 = ~n17247 & n17756 ;
  assign n17758 = n5503 & n12454 ;
  assign n17759 = n5512 & n12459 ;
  assign n17760 = n5508 & ~n12456 ;
  assign n17761 = n17759 | n17760 ;
  assign n17762 = n17758 | n17761 ;
  assign n17763 = n5515 | n17762 ;
  assign n17764 = ( n14041 & n17762 ) | ( n14041 & n17763 ) | ( n17762 & n17763 ) ;
  assign n17765 = x8 & n17764 ;
  assign n17766 = x8 & ~n17765 ;
  assign n17767 = ( n17764 & ~n17765 ) | ( n17764 & n17766 ) | ( ~n17765 & n17766 ) ;
  assign n17768 = n17757 & n17767 ;
  assign n17769 = n17757 | n17767 ;
  assign n17770 = ~n17768 & n17769 ;
  assign n17771 = x8 & ~n5502 ;
  assign n17772 = ( x8 & n12468 ) | ( x8 & n17771 ) | ( n12468 & n17771 ) ;
  assign n17773 = n5515 & n13994 ;
  assign n17774 = n5508 & ~n12468 ;
  assign n17775 = n5503 & ~n12466 ;
  assign n17776 = n17774 | n17775 ;
  assign n17777 = n17773 | n17776 ;
  assign n17778 = x8 | n17777 ;
  assign n17779 = ~x8 & n17778 ;
  assign n17780 = ( ~n17777 & n17778 ) | ( ~n17777 & n17779 ) | ( n17778 & n17779 ) ;
  assign n17781 = n17772 & n17780 ;
  assign n17782 = n7298 & ~n12468 ;
  assign n17783 = n5503 & n12459 ;
  assign n17784 = n5512 & ~n12468 ;
  assign n17785 = n5508 & ~n12466 ;
  assign n17786 = n17784 | n17785 ;
  assign n17787 = n17783 | n17786 ;
  assign n17788 = n5515 & n14003 ;
  assign n17789 = n17787 | n17788 ;
  assign n17790 = ~x8 & n17789 ;
  assign n17791 = x8 | n17790 ;
  assign n17792 = ( ~n17789 & n17790 ) | ( ~n17789 & n17791 ) | ( n17790 & n17791 ) ;
  assign n17793 = n17782 & n17792 ;
  assign n17794 = n17781 & n17793 ;
  assign n17795 = n17781 & n17792 ;
  assign n17796 = n17782 | n17795 ;
  assign n17797 = ~n17794 & n17796 ;
  assign n17798 = n5503 & ~n12456 ;
  assign n17799 = n5512 & ~n12466 ;
  assign n17800 = n5508 & n12459 ;
  assign n17801 = n17799 | n17800 ;
  assign n17802 = n17798 | n17801 ;
  assign n17803 = ( n5515 & n14031 ) | ( n5515 & n17802 ) | ( n14031 & n17802 ) ;
  assign n17804 = ( x8 & ~n17802 ) | ( x8 & n17803 ) | ( ~n17802 & n17803 ) ;
  assign n17805 = ~n17803 & n17804 ;
  assign n17806 = n17802 | n17804 ;
  assign n17807 = ( ~x8 & n17805 ) | ( ~x8 & n17806 ) | ( n17805 & n17806 ) ;
  assign n17808 = n17797 & n17807 ;
  assign n17809 = n17794 | n17808 ;
  assign n17810 = n17770 & n17809 ;
  assign n17811 = n17768 | n17810 ;
  assign n17812 = n17752 | n17754 ;
  assign n17813 = ~n17755 & n17812 ;
  assign n17814 = n17811 & n17813 ;
  assign n17815 = n17755 | n17814 ;
  assign n17816 = n17742 & n17815 ;
  assign n17817 = n17740 | n17816 ;
  assign n17818 = n17726 & ~n17727 ;
  assign n17819 = ( n17716 & ~n17727 ) | ( n17716 & n17818 ) | ( ~n17727 & n17818 ) ;
  assign n17820 = n17817 & n17819 ;
  assign n17821 = n17727 | n17820 ;
  assign n17822 = ( n17703 & n17714 ) | ( n17703 & n17821 ) | ( n17714 & n17821 ) ;
  assign n17823 = n17701 & n17822 ;
  assign n17824 = n17698 | n17823 ;
  assign n17825 = n17674 | n17684 ;
  assign n17826 = ~n17685 & n17825 ;
  assign n17827 = n17824 & n17826 ;
  assign n17828 = n17685 | n17827 ;
  assign n17829 = n17672 & n17828 ;
  assign n17830 = n17670 | n17829 ;
  assign n17831 = n17657 & n17830 ;
  assign n17832 = n17654 | n17831 ;
  assign n17833 = n17641 & n17832 ;
  assign n17834 = n17639 | n17833 ;
  assign n17835 = n17614 & ~n17626 ;
  assign n17836 = ~n17614 & n17625 ;
  assign n17837 = n17835 | n17836 ;
  assign n17838 = n17834 & n17837 ;
  assign n17839 = n17626 | n17838 ;
  assign n17840 = n17601 & ~n17612 ;
  assign n17841 = ~n17601 & n17611 ;
  assign n17842 = n17840 | n17841 ;
  assign n17843 = n17839 & n17842 ;
  assign n17844 = n17588 | n17598 ;
  assign n17845 = ~n17599 & n17844 ;
  assign n17846 = ( n17612 & n17843 ) | ( n17612 & n17845 ) | ( n17843 & n17845 ) ;
  assign n17847 = n17599 | n17846 ;
  assign n17848 = n17586 & n17847 ;
  assign n17849 = n17583 | n17848 ;
  assign n17850 = n17569 & n17849 ;
  assign n17851 = n17566 | n17850 ;
  assign n17852 = n17551 & ~n17552 ;
  assign n17853 = ( n17541 & ~n17552 ) | ( n17541 & n17852 ) | ( ~n17552 & n17852 ) ;
  assign n17854 = n17851 & n17853 ;
  assign n17855 = n17552 | n17854 ;
  assign n17856 = ( n17528 & n17538 ) | ( n17528 & n17855 ) | ( n17538 & n17855 ) ;
  assign n17857 = ( n17515 & n17526 ) | ( n17515 & n17856 ) | ( n17526 & n17856 ) ;
  assign n17858 = n17513 & n17857 ;
  assign n17859 = n17511 | n17858 ;
  assign n17860 = n17497 & n17859 ;
  assign n17861 = n17495 | n17860 ;
  assign n17862 = n17482 & n17861 ;
  assign n17863 = n17480 | n17862 ;
  assign n17864 = n17455 | n17467 ;
  assign n17865 = ( ~n17466 & n17467 ) | ( ~n17466 & n17864 ) | ( n17467 & n17864 ) ;
  assign n17866 = n17863 & ~n17865 ;
  assign n17867 = n17467 | n17866 ;
  assign n17868 = n17441 | n17453 ;
  assign n17869 = ( ~n17452 & n17453 ) | ( ~n17452 & n17868 ) | ( n17453 & n17868 ) ;
  assign n17870 = n17867 & ~n17869 ;
  assign n17871 = n17453 | n17870 ;
  assign n17872 = n17428 & ~n17439 ;
  assign n17873 = ~n17428 & n17438 ;
  assign n17874 = n17872 | n17873 ;
  assign n17875 = n17871 & n17874 ;
  assign n17876 = n17439 | n17875 ;
  assign n17877 = n17415 | n17426 ;
  assign n17878 = ( ~n17425 & n17426 ) | ( ~n17425 & n17877 ) | ( n17426 & n17877 ) ;
  assign n17879 = n17876 & ~n17878 ;
  assign n17880 = n17426 | n17879 ;
  assign n17881 = n17402 | n17413 ;
  assign n17882 = ( ~n17412 & n17413 ) | ( ~n17412 & n17881 ) | ( n17413 & n17881 ) ;
  assign n17883 = n17880 & ~n17882 ;
  assign n17884 = n17413 | n17883 ;
  assign n17885 = n17388 & ~n17400 ;
  assign n17886 = ~n17388 & n17399 ;
  assign n17887 = n17885 | n17886 ;
  assign n17888 = n17884 & n17887 ;
  assign n17889 = n17400 | n17888 ;
  assign n17890 = n17375 & ~n17386 ;
  assign n17891 = ~n17375 & n17385 ;
  assign n17892 = n17890 | n17891 ;
  assign n17893 = n17889 & n17892 ;
  assign n17894 = n17386 | n17893 ;
  assign n17895 = n16870 | n17338 ;
  assign n17896 = ~n17339 & n17895 ;
  assign n17897 = n5503 & ~n12586 ;
  assign n17898 = n5512 & n12340 ;
  assign n17899 = n5508 & ~n12344 ;
  assign n17900 = n17898 | n17899 ;
  assign n17901 = n17897 | n17900 ;
  assign n17902 = n5515 & ~n13454 ;
  assign n17903 = ~n13455 & n17902 ;
  assign n17904 = ( n5515 & n17901 ) | ( n5515 & ~n17903 ) | ( n17901 & ~n17903 ) ;
  assign n17905 = ~x8 & n17904 ;
  assign n17906 = x8 | n17905 ;
  assign n17907 = ( ~n17904 & n17905 ) | ( ~n17904 & n17906 ) | ( n17905 & n17906 ) ;
  assign n17908 = ( n17894 & n17896 ) | ( n17894 & n17907 ) | ( n17896 & n17907 ) ;
  assign n17909 = n17373 & n17908 ;
  assign n17910 = n17354 | n17357 ;
  assign n17911 = n16378 | n16817 ;
  assign n17912 = ~n16818 & n17911 ;
  assign n17913 = n7305 & ~n12344 ;
  assign n17914 = n7300 & n12553 ;
  assign n17915 = n7302 & n12340 ;
  assign n17916 = n17914 | n17915 ;
  assign n17917 = n17913 | n17916 ;
  assign n17918 = n7308 | n17917 ;
  assign n17919 = ( ~n13523 & n17917 ) | ( ~n13523 & n17918 ) | ( n17917 & n17918 ) ;
  assign n17920 = ~x11 & n17919 ;
  assign n17921 = x11 | n17920 ;
  assign n17922 = ( ~n17919 & n17920 ) | ( ~n17919 & n17921 ) | ( n17920 & n17921 ) ;
  assign n17923 = n17912 & n17922 ;
  assign n17924 = n17922 & ~n17923 ;
  assign n17925 = ( n17912 & ~n17923 ) | ( n17912 & n17924 ) | ( ~n17923 & n17924 ) ;
  assign n17926 = n17910 & n17925 ;
  assign n17927 = n17910 | n17925 ;
  assign n17928 = ~n17926 & n17927 ;
  assign n17929 = n5503 & ~n12335 ;
  assign n17930 = n5512 & ~n12586 ;
  assign n17931 = n5508 & n12580 ;
  assign n17932 = n17930 | n17931 ;
  assign n17933 = n17929 | n17932 ;
  assign n17934 = n5515 & ~n13585 ;
  assign n17935 = ~n13587 & n17934 ;
  assign n17936 = ( n5515 & n17933 ) | ( n5515 & ~n17935 ) | ( n17933 & ~n17935 ) ;
  assign n17937 = ~x8 & n17936 ;
  assign n17938 = x8 | n17937 ;
  assign n17939 = ( ~n17936 & n17937 ) | ( ~n17936 & n17938 ) | ( n17937 & n17938 ) ;
  assign n17940 = n17928 & n17939 ;
  assign n17941 = n17928 | n17939 ;
  assign n17942 = ~n17940 & n17941 ;
  assign n17943 = n17370 | n17942 ;
  assign n17944 = n17909 | n17943 ;
  assign n17945 = ( n17370 & n17909 ) | ( n17370 & n17942 ) | ( n17909 & n17942 ) ;
  assign n17946 = n17944 & ~n17945 ;
  assign n17947 = n8680 & ~n12325 ;
  assign n17948 = n8681 & ~n12328 ;
  assign n17949 = n17947 | n17948 ;
  assign n17950 = n9245 & n12608 ;
  assign n17951 = n17949 | n17950 ;
  assign n17952 = n8685 & n13570 ;
  assign n17953 = ( n8685 & n13568 ) | ( n8685 & n17952 ) | ( n13568 & n17952 ) ;
  assign n17954 = n17951 | n17953 ;
  assign n17955 = x5 | n17954 ;
  assign n17956 = ~x5 & n17955 ;
  assign n17957 = ( ~n17954 & n17955 ) | ( ~n17954 & n17956 ) | ( n17955 & n17956 ) ;
  assign n17958 = n17946 & n17957 ;
  assign n17959 = n17946 & ~n17958 ;
  assign n17960 = ~n17946 & n17957 ;
  assign n17961 = n17959 | n17960 ;
  assign n17962 = n9783 | n9798 ;
  assign n17963 = ~n12314 & n17962 ;
  assign n17964 = n9782 | n17963 ;
  assign n17965 = ( ~n12318 & n17963 ) | ( ~n12318 & n17964 ) | ( n17963 & n17964 ) ;
  assign n17966 = ( n12314 & ~n12604 ) | ( n12314 & n12615 ) | ( ~n12604 & n12615 ) ;
  assign n17967 = n9787 & ~n17966 ;
  assign n17968 = n17965 | n17967 ;
  assign n17969 = x2 & ~n17968 ;
  assign n17970 = ~x2 & n17968 ;
  assign n17971 = n17969 | n17970 ;
  assign n17972 = n17961 & n17971 ;
  assign n17973 = n17958 | n17972 ;
  assign n17974 = n9245 & ~n12318 ;
  assign n17975 = n8680 & ~n12328 ;
  assign n17976 = n8681 & n12608 ;
  assign n17977 = n17975 | n17976 ;
  assign n17978 = n17974 | n17977 ;
  assign n17979 = n8685 | n17978 ;
  assign n17980 = ( n14320 & n17978 ) | ( n14320 & n17979 ) | ( n17978 & n17979 ) ;
  assign n17981 = x5 & n17980 ;
  assign n17982 = x5 & ~n17981 ;
  assign n17983 = ( n17980 & ~n17981 ) | ( n17980 & n17982 ) | ( ~n17981 & n17982 ) ;
  assign n17984 = n17940 | n17945 ;
  assign n17985 = n5503 & ~n12325 ;
  assign n17986 = n5512 & n12580 ;
  assign n17987 = n5508 & ~n12335 ;
  assign n17988 = n17986 | n17987 ;
  assign n17989 = n17985 | n17988 ;
  assign n17990 = n5515 | n17989 ;
  assign n17991 = ( ~n13720 & n17989 ) | ( ~n13720 & n17990 ) | ( n17989 & n17990 ) ;
  assign n17992 = ~x8 & n17991 ;
  assign n17993 = x8 | n17992 ;
  assign n17994 = ( ~n17991 & n17992 ) | ( ~n17991 & n17993 ) | ( n17992 & n17993 ) ;
  assign n17995 = ( ~n16829 & n16830 ) | ( ~n16829 & n16831 ) | ( n16830 & n16831 ) ;
  assign n17996 = n17923 | n17926 ;
  assign n17997 = ( n17994 & n17995 ) | ( n17994 & ~n17996 ) | ( n17995 & ~n17996 ) ;
  assign n17998 = ( ~n17995 & n17996 ) | ( ~n17995 & n17997 ) | ( n17996 & n17997 ) ;
  assign n17999 = ( ~n17994 & n17997 ) | ( ~n17994 & n17998 ) | ( n17997 & n17998 ) ;
  assign n18000 = ( n17983 & ~n17984 ) | ( n17983 & n17999 ) | ( ~n17984 & n17999 ) ;
  assign n18001 = ( n17984 & ~n17999 ) | ( n17984 & n18000 ) | ( ~n17999 & n18000 ) ;
  assign n18002 = ( ~n17983 & n18000 ) | ( ~n17983 & n18001 ) | ( n18000 & n18001 ) ;
  assign n18003 = n17973 & ~n18002 ;
  assign n18004 = n9245 & ~n12328 ;
  assign n18005 = n8680 & ~n12335 ;
  assign n18006 = n8681 & ~n12325 ;
  assign n18007 = n18005 | n18006 ;
  assign n18008 = n18004 | n18007 ;
  assign n18009 = n8685 | n18008 ;
  assign n18010 = ( ~n13544 & n18008 ) | ( ~n13544 & n18009 ) | ( n18008 & n18009 ) ;
  assign n18011 = ~x5 & n18010 ;
  assign n18012 = x5 | n18011 ;
  assign n18013 = ( ~n18010 & n18011 ) | ( ~n18010 & n18012 ) | ( n18011 & n18012 ) ;
  assign n18014 = n17373 & ~n17909 ;
  assign n18015 = ( n17908 & ~n17909 ) | ( n17908 & n18014 ) | ( ~n17909 & n18014 ) ;
  assign n18016 = n18013 & n18015 ;
  assign n18017 = n18015 & ~n18016 ;
  assign n18018 = n18013 & ~n18015 ;
  assign n18019 = n18017 | n18018 ;
  assign n18020 = n9245 & ~n12325 ;
  assign n18021 = n8680 & n12580 ;
  assign n18022 = n8681 & ~n12335 ;
  assign n18023 = n18021 | n18022 ;
  assign n18024 = n18020 | n18023 ;
  assign n18025 = n8685 | n18024 ;
  assign n18026 = ( ~n13720 & n18024 ) | ( ~n13720 & n18025 ) | ( n18024 & n18025 ) ;
  assign n18027 = ~x5 & n18026 ;
  assign n18028 = x5 | n18027 ;
  assign n18029 = ( ~n18026 & n18027 ) | ( ~n18026 & n18028 ) | ( n18027 & n18028 ) ;
  assign n18030 = ( n17894 & ~n17896 ) | ( n17894 & n17907 ) | ( ~n17896 & n17907 ) ;
  assign n18031 = ( ~n17894 & n17896 ) | ( ~n17894 & n18030 ) | ( n17896 & n18030 ) ;
  assign n18032 = ( ~n17907 & n18030 ) | ( ~n17907 & n18031 ) | ( n18030 & n18031 ) ;
  assign n18033 = n18029 & n18032 ;
  assign n18034 = n18029 | n18032 ;
  assign n18035 = ~n18033 & n18034 ;
  assign n18036 = n17889 & ~n17893 ;
  assign n18037 = n17892 & ~n17893 ;
  assign n18038 = n18036 | n18037 ;
  assign n18039 = n9245 & ~n12335 ;
  assign n18040 = n8680 & ~n12586 ;
  assign n18041 = n8681 & n12580 ;
  assign n18042 = n18040 | n18041 ;
  assign n18043 = n18039 | n18042 ;
  assign n18044 = n8685 & n13587 ;
  assign n18045 = ( n8685 & n13585 ) | ( n8685 & n18044 ) | ( n13585 & n18044 ) ;
  assign n18046 = n18043 | n18045 ;
  assign n18047 = x5 | n18046 ;
  assign n18048 = ~x5 & n18047 ;
  assign n18049 = ( ~n18046 & n18047 ) | ( ~n18046 & n18048 ) | ( n18047 & n18048 ) ;
  assign n18050 = n18038 & n18049 ;
  assign n18051 = n18038 & ~n18050 ;
  assign n18052 = ~n18038 & n18049 ;
  assign n18053 = n18051 | n18052 ;
  assign n18054 = n17884 & ~n17888 ;
  assign n18055 = n17887 & ~n17888 ;
  assign n18056 = n18054 | n18055 ;
  assign n18057 = n9245 & n12580 ;
  assign n18058 = n8680 & ~n12344 ;
  assign n18059 = n8681 & ~n12586 ;
  assign n18060 = n18058 | n18059 ;
  assign n18061 = n18057 | n18060 ;
  assign n18062 = n8685 | n18061 ;
  assign n18063 = ( n13432 & n18061 ) | ( n13432 & n18062 ) | ( n18061 & n18062 ) ;
  assign n18064 = x5 & n18063 ;
  assign n18065 = x5 & ~n18064 ;
  assign n18066 = ( n18063 & ~n18064 ) | ( n18063 & n18065 ) | ( ~n18064 & n18065 ) ;
  assign n18067 = n18056 & n18066 ;
  assign n18068 = n18056 & ~n18067 ;
  assign n18069 = ~n18056 & n18066 ;
  assign n18070 = n18068 | n18069 ;
  assign n18071 = n17880 & ~n17883 ;
  assign n18072 = n17882 | n17883 ;
  assign n18073 = ~n18071 & n18072 ;
  assign n18074 = n9245 & ~n12586 ;
  assign n18075 = n8680 & n12340 ;
  assign n18076 = n8681 & ~n12344 ;
  assign n18077 = n18075 | n18076 ;
  assign n18078 = n18074 | n18077 ;
  assign n18079 = ( n8685 & n13454 ) | ( n8685 & n13455 ) | ( n13454 & n13455 ) ;
  assign n18080 = n18078 | n18079 ;
  assign n18081 = x5 | n18080 ;
  assign n18082 = ~x5 & n18081 ;
  assign n18083 = ( ~n18080 & n18081 ) | ( ~n18080 & n18082 ) | ( n18081 & n18082 ) ;
  assign n18084 = ~n18073 & n18083 ;
  assign n18085 = n17876 & ~n17879 ;
  assign n18086 = n17878 | n17879 ;
  assign n18087 = ~n18085 & n18086 ;
  assign n18088 = n9245 & ~n12344 ;
  assign n18089 = n8680 & n12553 ;
  assign n18090 = n8681 & n12340 ;
  assign n18091 = n18089 | n18090 ;
  assign n18092 = n18088 | n18091 ;
  assign n18093 = n8685 | n18092 ;
  assign n18094 = ( ~n13523 & n18092 ) | ( ~n13523 & n18093 ) | ( n18092 & n18093 ) ;
  assign n18095 = ~x5 & n18094 ;
  assign n18096 = x5 | n18095 ;
  assign n18097 = ( ~n18094 & n18095 ) | ( ~n18094 & n18096 ) | ( n18095 & n18096 ) ;
  assign n18098 = ~n18087 & n18097 ;
  assign n18099 = n17871 & ~n17875 ;
  assign n18100 = n17874 & ~n17875 ;
  assign n18101 = n18099 | n18100 ;
  assign n18102 = n9245 & n12340 ;
  assign n18103 = n8680 & n12558 ;
  assign n18104 = n8681 & n12553 ;
  assign n18105 = n18103 | n18104 ;
  assign n18106 = n18102 | n18105 ;
  assign n18107 = n8685 & n13347 ;
  assign n18108 = ( n8685 & n13346 ) | ( n8685 & n18107 ) | ( n13346 & n18107 ) ;
  assign n18109 = n18106 | n18108 ;
  assign n18110 = x5 | n18109 ;
  assign n18111 = ~x5 & n18110 ;
  assign n18112 = ( ~n18109 & n18110 ) | ( ~n18109 & n18111 ) | ( n18110 & n18111 ) ;
  assign n18113 = n18101 & n18112 ;
  assign n18114 = n18101 & ~n18113 ;
  assign n18115 = ~n18101 & n18112 ;
  assign n18116 = n18114 | n18115 ;
  assign n18117 = n17867 & ~n17870 ;
  assign n18118 = n17869 | n17870 ;
  assign n18119 = ~n18117 & n18118 ;
  assign n18120 = n9245 & n12553 ;
  assign n18121 = n8680 & n12355 ;
  assign n18122 = n8681 & n12558 ;
  assign n18123 = n18121 | n18122 ;
  assign n18124 = n18120 | n18123 ;
  assign n18125 = n8685 | n18124 ;
  assign n18126 = ( n13097 & n18124 ) | ( n13097 & n18125 ) | ( n18124 & n18125 ) ;
  assign n18127 = x5 & n18126 ;
  assign n18128 = x5 & ~n18127 ;
  assign n18129 = ( n18126 & ~n18127 ) | ( n18126 & n18128 ) | ( ~n18127 & n18128 ) ;
  assign n18130 = ~n18119 & n18129 ;
  assign n18131 = n17863 & ~n17866 ;
  assign n18132 = n17865 | n17866 ;
  assign n18133 = ~n18131 & n18132 ;
  assign n18134 = n9245 & n12558 ;
  assign n18135 = n8680 & n12351 ;
  assign n18136 = n8681 & n12355 ;
  assign n18137 = n18135 | n18136 ;
  assign n18138 = n18134 | n18137 ;
  assign n18139 = n8685 | n18138 ;
  assign n18140 = ( n13330 & n18138 ) | ( n13330 & n18139 ) | ( n18138 & n18139 ) ;
  assign n18141 = x5 & n18140 ;
  assign n18142 = x5 & ~n18141 ;
  assign n18143 = ( n18140 & ~n18141 ) | ( n18140 & n18142 ) | ( ~n18141 & n18142 ) ;
  assign n18144 = ~n18133 & n18143 ;
  assign n18145 = n17482 | n17861 ;
  assign n18146 = ~n17862 & n18145 ;
  assign n18147 = n9245 & n12355 ;
  assign n18148 = n8680 & ~n12537 ;
  assign n18149 = n8681 & n12351 ;
  assign n18150 = n18148 | n18149 ;
  assign n18151 = n18147 | n18150 ;
  assign n18152 = n8685 | n18151 ;
  assign n18153 = ( n13409 & n18151 ) | ( n13409 & n18152 ) | ( n18151 & n18152 ) ;
  assign n18154 = x5 & n18153 ;
  assign n18155 = x5 & ~n18154 ;
  assign n18156 = ( n18153 & ~n18154 ) | ( n18153 & n18155 ) | ( ~n18154 & n18155 ) ;
  assign n18157 = n18146 & n18156 ;
  assign n18158 = n17497 | n17859 ;
  assign n18159 = ~n17860 & n18158 ;
  assign n18160 = n9245 & n12351 ;
  assign n18161 = n8680 & n12364 ;
  assign n18162 = n8681 & ~n12537 ;
  assign n18163 = n18161 | n18162 ;
  assign n18164 = n18160 | n18163 ;
  assign n18165 = n8685 & n12928 ;
  assign n18166 = ~n12925 & n18165 ;
  assign n18167 = ( n8685 & n18164 ) | ( n8685 & ~n18166 ) | ( n18164 & ~n18166 ) ;
  assign n18168 = x5 & n18167 ;
  assign n18169 = x5 & ~n18168 ;
  assign n18170 = ( n18167 & ~n18168 ) | ( n18167 & n18169 ) | ( ~n18168 & n18169 ) ;
  assign n18171 = n18159 & n18170 ;
  assign n18172 = n18146 | n18156 ;
  assign n18173 = ~n18157 & n18172 ;
  assign n18174 = n17513 | n17857 ;
  assign n18175 = ~n17858 & n18174 ;
  assign n18176 = n9245 & ~n12537 ;
  assign n18177 = n8680 & ~n12360 ;
  assign n18178 = n8681 & n12364 ;
  assign n18179 = n18177 | n18178 ;
  assign n18180 = n18176 | n18179 ;
  assign n18181 = ( n8685 & n13081 ) | ( n8685 & ~n13082 ) | ( n13081 & ~n13082 ) ;
  assign n18182 = n18180 | n18181 ;
  assign n18183 = x5 | n18182 ;
  assign n18184 = ~x5 & n18183 ;
  assign n18185 = ( ~n18182 & n18183 ) | ( ~n18182 & n18184 ) | ( n18183 & n18184 ) ;
  assign n18186 = n18175 & n18185 ;
  assign n18187 = n18185 & ~n18186 ;
  assign n18188 = ( n18175 & ~n18186 ) | ( n18175 & n18187 ) | ( ~n18186 & n18187 ) ;
  assign n18189 = n9245 & n12364 ;
  assign n18190 = n8680 & n12520 ;
  assign n18191 = n8681 & ~n12360 ;
  assign n18192 = n18190 | n18191 ;
  assign n18193 = n18189 | n18192 ;
  assign n18194 = n8685 | n18193 ;
  assign n18195 = ( ~n13113 & n18193 ) | ( ~n13113 & n18194 ) | ( n18193 & n18194 ) ;
  assign n18196 = ~x5 & n18195 ;
  assign n18197 = x5 | n18196 ;
  assign n18198 = ( ~n18195 & n18196 ) | ( ~n18195 & n18197 ) | ( n18196 & n18197 ) ;
  assign n18199 = n9245 & ~n12360 ;
  assign n18200 = n8680 & n12375 ;
  assign n18201 = n8681 & n12520 ;
  assign n18202 = n18200 | n18201 ;
  assign n18203 = n18199 | n18202 ;
  assign n18204 = n8685 | n18203 ;
  assign n18205 = ( ~n12902 & n18203 ) | ( ~n12902 & n18204 ) | ( n18203 & n18204 ) ;
  assign n18206 = ~x5 & n18205 ;
  assign n18207 = x5 | n18206 ;
  assign n18208 = ( ~n18205 & n18206 ) | ( ~n18205 & n18207 ) | ( n18206 & n18207 ) ;
  assign n18209 = n17851 | n17853 ;
  assign n18210 = ~n17854 & n18209 ;
  assign n18211 = n9245 & n12520 ;
  assign n18212 = n8680 & ~n12371 ;
  assign n18213 = n8681 & n12375 ;
  assign n18214 = n18212 | n18213 ;
  assign n18215 = n18211 | n18214 ;
  assign n18216 = n8685 & ~n12837 ;
  assign n18217 = ~n12835 & n18216 ;
  assign n18218 = ( n8685 & n18215 ) | ( n8685 & ~n18217 ) | ( n18215 & ~n18217 ) ;
  assign n18219 = ~x5 & n18218 ;
  assign n18220 = x5 | n18219 ;
  assign n18221 = ( ~n18218 & n18219 ) | ( ~n18218 & n18220 ) | ( n18219 & n18220 ) ;
  assign n18222 = n18210 & n18221 ;
  assign n18223 = n18210 | n18221 ;
  assign n18224 = ~n18222 & n18223 ;
  assign n18225 = n17569 | n17849 ;
  assign n18226 = ~n17850 & n18225 ;
  assign n18227 = n9245 & n12375 ;
  assign n18228 = n8680 & n12378 ;
  assign n18229 = n8681 & ~n12371 ;
  assign n18230 = n18228 | n18229 ;
  assign n18231 = n18227 | n18230 ;
  assign n18232 = n8685 & n13065 ;
  assign n18233 = ~n13064 & n18232 ;
  assign n18234 = ( n8685 & n18231 ) | ( n8685 & ~n18233 ) | ( n18231 & ~n18233 ) ;
  assign n18235 = x5 & n18234 ;
  assign n18236 = x5 & ~n18235 ;
  assign n18237 = ( n18234 & ~n18235 ) | ( n18234 & n18236 ) | ( ~n18235 & n18236 ) ;
  assign n18238 = n17586 | n17847 ;
  assign n18239 = ~n17848 & n18238 ;
  assign n18240 = n9245 & ~n12371 ;
  assign n18241 = n8680 & ~n12502 ;
  assign n18242 = n8681 & n12378 ;
  assign n18243 = n18241 | n18242 ;
  assign n18244 = n18240 | n18243 ;
  assign n18245 = n8685 | n18244 ;
  assign n18246 = ( ~n12848 & n18244 ) | ( ~n12848 & n18245 ) | ( n18244 & n18245 ) ;
  assign n18247 = ~x5 & n18246 ;
  assign n18248 = x5 | n18247 ;
  assign n18249 = ( ~n18246 & n18247 ) | ( ~n18246 & n18248 ) | ( n18247 & n18248 ) ;
  assign n18250 = n17612 | n17845 ;
  assign n18251 = n17843 | n18250 ;
  assign n18252 = ~n17846 & n18251 ;
  assign n18253 = n9245 & n12378 ;
  assign n18254 = n8680 & n12387 ;
  assign n18255 = n8681 & ~n12502 ;
  assign n18256 = n18254 | n18255 ;
  assign n18257 = n18253 | n18256 ;
  assign n18258 = n8685 | n18257 ;
  assign n18259 = ( ~n12816 & n18257 ) | ( ~n12816 & n18258 ) | ( n18257 & n18258 ) ;
  assign n18260 = ~x5 & n18259 ;
  assign n18261 = x5 | n18260 ;
  assign n18262 = ( ~n18259 & n18260 ) | ( ~n18259 & n18261 ) | ( n18260 & n18261 ) ;
  assign n18263 = n17839 & ~n17843 ;
  assign n18264 = n17842 & ~n17843 ;
  assign n18265 = n18263 | n18264 ;
  assign n18266 = n9245 & ~n12502 ;
  assign n18267 = n8680 & n12383 ;
  assign n18268 = n8681 & n12387 ;
  assign n18269 = n18267 | n18268 ;
  assign n18270 = n18266 | n18269 ;
  assign n18271 = n8685 | n18270 ;
  assign n18272 = ( ~n12756 & n18270 ) | ( ~n12756 & n18271 ) | ( n18270 & n18271 ) ;
  assign n18273 = ~x5 & n18272 ;
  assign n18274 = x5 | n18273 ;
  assign n18275 = ( ~n18272 & n18273 ) | ( ~n18272 & n18274 ) | ( n18273 & n18274 ) ;
  assign n18276 = n17834 & ~n17838 ;
  assign n18277 = n17837 & ~n17838 ;
  assign n18278 = n18276 | n18277 ;
  assign n18279 = n9245 & n12387 ;
  assign n18280 = n8680 & n12392 ;
  assign n18281 = n8681 & n12383 ;
  assign n18282 = n18280 | n18281 ;
  assign n18283 = n18279 | n18282 ;
  assign n18284 = n8685 | n18283 ;
  assign n18285 = ( n12948 & n18283 ) | ( n12948 & n18284 ) | ( n18283 & n18284 ) ;
  assign n18286 = x5 & n18285 ;
  assign n18287 = x5 & ~n18286 ;
  assign n18288 = ( n18285 & ~n18286 ) | ( n18285 & n18287 ) | ( ~n18286 & n18287 ) ;
  assign n18289 = n17641 | n17832 ;
  assign n18290 = ~n17833 & n18289 ;
  assign n18291 = n9245 & n12383 ;
  assign n18292 = n8680 & n12401 ;
  assign n18293 = n8681 & n12392 ;
  assign n18294 = n18292 | n18293 ;
  assign n18295 = n18291 | n18294 ;
  assign n18296 = n8685 | n18295 ;
  assign n18297 = ( n13141 & n18295 ) | ( n13141 & n18296 ) | ( n18295 & n18296 ) ;
  assign n18298 = x5 & n18297 ;
  assign n18299 = x5 & ~n18298 ;
  assign n18300 = ( n18297 & ~n18298 ) | ( n18297 & n18299 ) | ( ~n18298 & n18299 ) ;
  assign n18301 = n18290 & n18300 ;
  assign n18302 = n17657 | n17830 ;
  assign n18303 = ~n17831 & n18302 ;
  assign n18304 = n9245 & n12392 ;
  assign n18305 = n8680 & n12415 ;
  assign n18306 = n8681 & n12401 ;
  assign n18307 = n18305 | n18306 ;
  assign n18308 = n18304 | n18307 ;
  assign n18309 = n8685 | n18308 ;
  assign n18310 = ( n13034 & n18308 ) | ( n13034 & n18309 ) | ( n18308 & n18309 ) ;
  assign n18311 = x5 & n18310 ;
  assign n18312 = x5 & ~n18311 ;
  assign n18313 = ( n18310 & ~n18311 ) | ( n18310 & n18312 ) | ( ~n18311 & n18312 ) ;
  assign n18314 = n18303 & n18313 ;
  assign n18315 = n18290 | n18300 ;
  assign n18316 = ~n18301 & n18315 ;
  assign n18317 = n17672 | n17828 ;
  assign n18318 = ~n17829 & n18317 ;
  assign n18319 = n9245 & n12401 ;
  assign n18320 = n8680 & n12411 ;
  assign n18321 = n8681 & n12415 ;
  assign n18322 = n18320 | n18321 ;
  assign n18323 = n18319 | n18322 ;
  assign n18324 = n8685 & ~n13163 ;
  assign n18325 = ~n13161 & n18324 ;
  assign n18326 = ( n8685 & n18323 ) | ( n8685 & ~n18325 ) | ( n18323 & ~n18325 ) ;
  assign n18327 = ~x5 & n18326 ;
  assign n18328 = x5 | n18327 ;
  assign n18329 = ( ~n18326 & n18327 ) | ( ~n18326 & n18328 ) | ( n18327 & n18328 ) ;
  assign n18330 = n18318 & n18329 ;
  assign n18331 = n17824 | n17826 ;
  assign n18332 = ~n17827 & n18331 ;
  assign n18333 = n9245 & n12415 ;
  assign n18334 = n8680 & n12419 ;
  assign n18335 = n8681 & n12411 ;
  assign n18336 = n18334 | n18335 ;
  assign n18337 = n18333 | n18336 ;
  assign n18338 = ( n8685 & n13761 ) | ( n8685 & n13762 ) | ( n13761 & n13762 ) ;
  assign n18339 = n18337 | n18338 ;
  assign n18340 = x5 | n18339 ;
  assign n18341 = ~x5 & n18340 ;
  assign n18342 = ( ~n18339 & n18340 ) | ( ~n18339 & n18341 ) | ( n18340 & n18341 ) ;
  assign n18343 = n18332 & n18342 ;
  assign n18344 = n18342 & ~n18343 ;
  assign n18345 = ( n18332 & ~n18343 ) | ( n18332 & n18344 ) | ( ~n18343 & n18344 ) ;
  assign n18346 = n9245 & n12411 ;
  assign n18347 = n8680 & ~n12423 ;
  assign n18348 = n8681 & n12419 ;
  assign n18349 = n18347 | n18348 ;
  assign n18350 = n18346 | n18349 ;
  assign n18351 = n8685 | n18350 ;
  assign n18352 = ( n13776 & n18350 ) | ( n13776 & n18351 ) | ( n18350 & n18351 ) ;
  assign n18353 = x5 & n18352 ;
  assign n18354 = x5 & ~n18353 ;
  assign n18355 = ( n18352 & ~n18353 ) | ( n18352 & n18354 ) | ( ~n18353 & n18354 ) ;
  assign n18356 = n9245 & n12419 ;
  assign n18357 = n8680 & n12433 ;
  assign n18358 = n8681 & ~n12423 ;
  assign n18359 = n18357 | n18358 ;
  assign n18360 = n18356 | n18359 ;
  assign n18361 = n8685 | n18360 ;
  assign n18362 = ( ~n13282 & n18360 ) | ( ~n13282 & n18361 ) | ( n18360 & n18361 ) ;
  assign n18363 = ~x5 & n18362 ;
  assign n18364 = x5 | n18363 ;
  assign n18365 = ( ~n18362 & n18363 ) | ( ~n18362 & n18364 ) | ( n18363 & n18364 ) ;
  assign n18366 = n17817 | n17819 ;
  assign n18367 = ~n17820 & n18366 ;
  assign n18368 = n9245 & ~n12423 ;
  assign n18369 = n8680 & ~n12438 ;
  assign n18370 = n8681 & n12433 ;
  assign n18371 = n18369 | n18370 ;
  assign n18372 = n18368 | n18371 ;
  assign n18373 = n8685 | n18372 ;
  assign n18374 = ( ~n13786 & n18372 ) | ( ~n13786 & n18373 ) | ( n18372 & n18373 ) ;
  assign n18375 = ~x5 & n18374 ;
  assign n18376 = x5 | n18375 ;
  assign n18377 = ( ~n18374 & n18375 ) | ( ~n18374 & n18376 ) | ( n18375 & n18376 ) ;
  assign n18378 = n18367 & n18377 ;
  assign n18379 = n17742 | n17815 ;
  assign n18380 = ~n17816 & n18379 ;
  assign n18381 = n9245 & n12433 ;
  assign n18382 = n8680 & n12440 ;
  assign n18383 = n8681 & ~n12438 ;
  assign n18384 = n18382 | n18383 ;
  assign n18385 = n18381 | n18384 ;
  assign n18386 = n8685 | n18385 ;
  assign n18387 = ( ~n14167 & n18385 ) | ( ~n14167 & n18386 ) | ( n18385 & n18386 ) ;
  assign n18388 = ~x5 & n18387 ;
  assign n18389 = x5 | n18388 ;
  assign n18390 = ( ~n18387 & n18388 ) | ( ~n18387 & n18389 ) | ( n18388 & n18389 ) ;
  assign n18391 = n18380 & n18390 ;
  assign n18392 = n18380 & ~n18391 ;
  assign n18393 = ~n18380 & n18390 ;
  assign n18394 = n18392 | n18393 ;
  assign n18395 = n17811 | n17813 ;
  assign n18396 = ~n17814 & n18395 ;
  assign n18397 = n9245 & ~n12438 ;
  assign n18398 = n8680 & n12446 ;
  assign n18399 = n8681 & n12440 ;
  assign n18400 = n18398 | n18399 ;
  assign n18401 = n18397 | n18400 ;
  assign n18402 = n8685 & n14154 ;
  assign n18403 = ~n14156 & n18402 ;
  assign n18404 = ( n8685 & n18401 ) | ( n8685 & ~n18403 ) | ( n18401 & ~n18403 ) ;
  assign n18405 = x5 & n18404 ;
  assign n18406 = x5 & ~n18405 ;
  assign n18407 = ( n18404 & ~n18405 ) | ( n18404 & n18406 ) | ( ~n18405 & n18406 ) ;
  assign n18408 = n17770 | n17809 ;
  assign n18409 = ~n17810 & n18408 ;
  assign n18410 = n9245 & n12440 ;
  assign n18411 = n8680 & n12452 ;
  assign n18412 = n8681 & n12446 ;
  assign n18413 = n18411 | n18412 ;
  assign n18414 = n18410 | n18413 ;
  assign n18415 = n8685 | n18414 ;
  assign n18416 = ( n13822 & n18414 ) | ( n13822 & n18415 ) | ( n18414 & n18415 ) ;
  assign n18417 = x5 & n18416 ;
  assign n18418 = x5 & ~n18417 ;
  assign n18419 = ( n18416 & ~n18417 ) | ( n18416 & n18418 ) | ( ~n18417 & n18418 ) ;
  assign n18420 = n9245 & n12446 ;
  assign n18421 = n8680 & n12454 ;
  assign n18422 = n8681 & n12452 ;
  assign n18423 = n18421 | n18422 ;
  assign n18424 = n18420 | n18423 ;
  assign n18425 = n8685 | n18424 ;
  assign n18426 = ( n13862 & n18424 ) | ( n13862 & n18425 ) | ( n18424 & n18425 ) ;
  assign n18427 = x5 & n18426 ;
  assign n18428 = x5 & ~n18427 ;
  assign n18429 = ( n18426 & ~n18427 ) | ( n18426 & n18428 ) | ( ~n18427 & n18428 ) ;
  assign n18430 = n17797 & ~n17808 ;
  assign n18431 = ( n17807 & ~n17808 ) | ( n17807 & n18430 ) | ( ~n17808 & n18430 ) ;
  assign n18432 = n18429 & n18431 ;
  assign n18433 = n18429 | n18431 ;
  assign n18434 = ~n18432 & n18433 ;
  assign n18435 = n17772 | n17780 ;
  assign n18436 = ~n17781 & n18435 ;
  assign n18437 = n9245 & n12454 ;
  assign n18438 = n8680 & n12459 ;
  assign n18439 = n8681 & ~n12456 ;
  assign n18440 = n18438 | n18439 ;
  assign n18441 = n18437 | n18440 ;
  assign n18442 = n8685 | n18441 ;
  assign n18443 = ( n14041 & n18441 ) | ( n14041 & n18442 ) | ( n18441 & n18442 ) ;
  assign n18444 = x5 & n18443 ;
  assign n18445 = x5 & ~n18444 ;
  assign n18446 = ( n18443 & ~n18444 ) | ( n18443 & n18445 ) | ( ~n18444 & n18445 ) ;
  assign n18447 = n18436 & n18446 ;
  assign n18448 = n18436 | n18446 ;
  assign n18449 = ~n18447 & n18448 ;
  assign n18450 = n5502 & ~n12468 ;
  assign n18451 = x5 & ~n8678 ;
  assign n18452 = ( x5 & n12468 ) | ( x5 & n18451 ) | ( n12468 & n18451 ) ;
  assign n18453 = n8685 & n13994 ;
  assign n18454 = n8681 & ~n12468 ;
  assign n18455 = n9245 & ~n12466 ;
  assign n18456 = n18454 | n18455 ;
  assign n18457 = n18453 | n18456 ;
  assign n18458 = x5 | n18457 ;
  assign n18459 = ~x5 & n18458 ;
  assign n18460 = ( ~n18457 & n18458 ) | ( ~n18457 & n18459 ) | ( n18458 & n18459 ) ;
  assign n18461 = n18452 & n18460 ;
  assign n18462 = n9245 & n12459 ;
  assign n18463 = n8680 & ~n12468 ;
  assign n18464 = n8681 & ~n12466 ;
  assign n18465 = n18463 | n18464 ;
  assign n18466 = n18462 | n18465 ;
  assign n18467 = n8685 & n14003 ;
  assign n18468 = n18466 | n18467 ;
  assign n18469 = ~x5 & n18468 ;
  assign n18470 = x5 | n18469 ;
  assign n18471 = ( ~n18468 & n18469 ) | ( ~n18468 & n18470 ) | ( n18469 & n18470 ) ;
  assign n18472 = n18461 & n18471 ;
  assign n18473 = n9245 & ~n12456 ;
  assign n18474 = n8680 & ~n12466 ;
  assign n18475 = n8681 & n12459 ;
  assign n18476 = n18474 | n18475 ;
  assign n18477 = n18473 | n18476 ;
  assign n18478 = ( n8685 & n14031 ) | ( n8685 & n18477 ) | ( n14031 & n18477 ) ;
  assign n18479 = ( x5 & ~n18477 ) | ( x5 & n18478 ) | ( ~n18477 & n18478 ) ;
  assign n18480 = ~n18478 & n18479 ;
  assign n18481 = n18477 | n18479 ;
  assign n18482 = ( ~x5 & n18480 ) | ( ~x5 & n18481 ) | ( n18480 & n18481 ) ;
  assign n18483 = ( n18450 & n18472 ) | ( n18450 & n18482 ) | ( n18472 & n18482 ) ;
  assign n18484 = n18449 & n18483 ;
  assign n18485 = n18447 | n18484 ;
  assign n18486 = n9245 & n12452 ;
  assign n18487 = n8680 & ~n12456 ;
  assign n18488 = n8681 & n12454 ;
  assign n18489 = n18487 | n18488 ;
  assign n18490 = n18486 | n18489 ;
  assign n18491 = n8685 | n18490 ;
  assign n18492 = ( ~n13922 & n18490 ) | ( ~n13922 & n18491 ) | ( n18490 & n18491 ) ;
  assign n18493 = ~x5 & n18492 ;
  assign n18494 = x5 & ~n18492 ;
  assign n18495 = n18493 | n18494 ;
  assign n18496 = n17781 | n17792 ;
  assign n18497 = ~n17795 & n18496 ;
  assign n18498 = ( n18485 & n18495 ) | ( n18485 & n18497 ) | ( n18495 & n18497 ) ;
  assign n18499 = n18434 & n18498 ;
  assign n18500 = n18432 | n18499 ;
  assign n18501 = ( n18409 & n18419 ) | ( n18409 & n18500 ) | ( n18419 & n18500 ) ;
  assign n18502 = ( n18396 & n18407 ) | ( n18396 & n18501 ) | ( n18407 & n18501 ) ;
  assign n18503 = n18394 & n18502 ;
  assign n18504 = n18391 | n18503 ;
  assign n18505 = n18367 | n18377 ;
  assign n18506 = ~n18378 & n18505 ;
  assign n18507 = n18504 & n18506 ;
  assign n18508 = n18378 | n18507 ;
  assign n18509 = ( n17703 & n17821 ) | ( n17703 & ~n17822 ) | ( n17821 & ~n17822 ) ;
  assign n18510 = ( n17714 & ~n17822 ) | ( n17714 & n18509 ) | ( ~n17822 & n18509 ) ;
  assign n18511 = ( n18365 & n18508 ) | ( n18365 & n18510 ) | ( n18508 & n18510 ) ;
  assign n18512 = n17701 & ~n17823 ;
  assign n18513 = ( n17822 & ~n17823 ) | ( n17822 & n18512 ) | ( ~n17823 & n18512 ) ;
  assign n18514 = ( n18355 & n18511 ) | ( n18355 & n18513 ) | ( n18511 & n18513 ) ;
  assign n18515 = n18345 & n18514 ;
  assign n18516 = n18343 | n18515 ;
  assign n18517 = n18318 & ~n18330 ;
  assign n18518 = ~n18318 & n18329 ;
  assign n18519 = ( n18516 & n18517 ) | ( n18516 & n18518 ) | ( n18517 & n18518 ) ;
  assign n18520 = n18330 | n18519 ;
  assign n18521 = n18303 & ~n18314 ;
  assign n18522 = ~n18303 & n18313 ;
  assign n18523 = ( n18520 & n18521 ) | ( n18520 & n18522 ) | ( n18521 & n18522 ) ;
  assign n18524 = ( n18314 & n18316 ) | ( n18314 & n18523 ) | ( n18316 & n18523 ) ;
  assign n18525 = n18301 | n18524 ;
  assign n18526 = ( n18278 & n18288 ) | ( n18278 & n18525 ) | ( n18288 & n18525 ) ;
  assign n18527 = ( n18265 & n18275 ) | ( n18265 & n18526 ) | ( n18275 & n18526 ) ;
  assign n18528 = ( n18252 & n18262 ) | ( n18252 & n18527 ) | ( n18262 & n18527 ) ;
  assign n18529 = ( n18239 & n18249 ) | ( n18239 & n18528 ) | ( n18249 & n18528 ) ;
  assign n18530 = ( n18226 & n18237 ) | ( n18226 & n18529 ) | ( n18237 & n18529 ) ;
  assign n18531 = n18224 & n18530 ;
  assign n18532 = n18222 | n18531 ;
  assign n18533 = ( n17528 & n17855 ) | ( n17528 & ~n17856 ) | ( n17855 & ~n17856 ) ;
  assign n18534 = ( n17538 & ~n17856 ) | ( n17538 & n18533 ) | ( ~n17856 & n18533 ) ;
  assign n18535 = ( n18208 & n18532 ) | ( n18208 & n18534 ) | ( n18532 & n18534 ) ;
  assign n18536 = ( n17515 & n17856 ) | ( n17515 & ~n17857 ) | ( n17856 & ~n17857 ) ;
  assign n18537 = ( n17526 & ~n17857 ) | ( n17526 & n18536 ) | ( ~n17857 & n18536 ) ;
  assign n18538 = ( n18198 & n18535 ) | ( n18198 & n18537 ) | ( n18535 & n18537 ) ;
  assign n18539 = n18188 & n18538 ;
  assign n18540 = n18186 | n18539 ;
  assign n18541 = n18159 & ~n18171 ;
  assign n18542 = ~n18159 & n18170 ;
  assign n18543 = ( n18540 & n18541 ) | ( n18540 & n18542 ) | ( n18541 & n18542 ) ;
  assign n18544 = ( n18171 & n18173 ) | ( n18171 & n18543 ) | ( n18173 & n18543 ) ;
  assign n18545 = n18157 | n18544 ;
  assign n18546 = n18133 | n18144 ;
  assign n18547 = ( ~n18143 & n18144 ) | ( ~n18143 & n18546 ) | ( n18144 & n18546 ) ;
  assign n18548 = n18545 & ~n18547 ;
  assign n18549 = n18144 | n18548 ;
  assign n18550 = n18119 | n18130 ;
  assign n18551 = ( ~n18129 & n18130 ) | ( ~n18129 & n18550 ) | ( n18130 & n18550 ) ;
  assign n18552 = n18549 & ~n18551 ;
  assign n18553 = n18130 | n18552 ;
  assign n18554 = n18116 & n18553 ;
  assign n18555 = n18113 | n18554 ;
  assign n18556 = n18087 | n18098 ;
  assign n18557 = ( ~n18097 & n18098 ) | ( ~n18097 & n18556 ) | ( n18098 & n18556 ) ;
  assign n18558 = n18555 & ~n18557 ;
  assign n18559 = n18098 | n18558 ;
  assign n18560 = n18073 | n18084 ;
  assign n18561 = ( ~n18083 & n18084 ) | ( ~n18083 & n18560 ) | ( n18084 & n18560 ) ;
  assign n18562 = n18559 & ~n18561 ;
  assign n18563 = n18084 | n18562 ;
  assign n18564 = n18070 & n18563 ;
  assign n18565 = n18067 | n18564 ;
  assign n18566 = n18053 & n18565 ;
  assign n18567 = n18050 | n18566 ;
  assign n18568 = n18035 & n18567 ;
  assign n18569 = n18033 | n18568 ;
  assign n18570 = n18019 & n18569 ;
  assign n18571 = n18016 | n18570 ;
  assign n18572 = n17961 | n17971 ;
  assign n18573 = ~n17972 & n18572 ;
  assign n18574 = n18571 & n18573 ;
  assign n18575 = n18019 | n18569 ;
  assign n18576 = ~n18570 & n18575 ;
  assign n18577 = n9783 & ~n12318 ;
  assign n18578 = n9782 & n12608 ;
  assign n18579 = n18577 | n18578 ;
  assign n18580 = n9798 & ~n12314 ;
  assign n18581 = n18579 | n18580 ;
  assign n18582 = n9787 | n18581 ;
  assign n18583 = ( ~n14302 & n18581 ) | ( ~n14302 & n18582 ) | ( n18581 & n18582 ) ;
  assign n18584 = ~x2 & n18583 ;
  assign n18585 = x2 | n18584 ;
  assign n18586 = ( ~n18583 & n18584 ) | ( ~n18583 & n18585 ) | ( n18584 & n18585 ) ;
  assign n18587 = n18576 & n18586 ;
  assign n18588 = n18576 | n18586 ;
  assign n18589 = ~n18587 & n18588 ;
  assign n18590 = n18035 | n18567 ;
  assign n18591 = ~n18568 & n18590 ;
  assign n18592 = n9798 & ~n12318 ;
  assign n18593 = n9782 & ~n12328 ;
  assign n18594 = n9783 & n12608 ;
  assign n18595 = n18593 | n18594 ;
  assign n18596 = n18592 | n18595 ;
  assign n18597 = n9787 | n18596 ;
  assign n18598 = ( n14320 & n18596 ) | ( n14320 & n18597 ) | ( n18596 & n18597 ) ;
  assign n18599 = x2 & n18598 ;
  assign n18600 = x2 & ~n18599 ;
  assign n18601 = ( n18598 & ~n18599 ) | ( n18598 & n18600 ) | ( ~n18599 & n18600 ) ;
  assign n18602 = n18591 & n18601 ;
  assign n18603 = n18053 | n18565 ;
  assign n18604 = ~n18566 & n18603 ;
  assign n18605 = n9782 & ~n12325 ;
  assign n18606 = n9783 & ~n12328 ;
  assign n18607 = n18605 | n18606 ;
  assign n18608 = n9798 & n12608 ;
  assign n18609 = n18607 | n18608 ;
  assign n18610 = n9787 & ~n13570 ;
  assign n18611 = ~n13568 & n18610 ;
  assign n18612 = ( n9787 & n18609 ) | ( n9787 & ~n18611 ) | ( n18609 & ~n18611 ) ;
  assign n18613 = ~x2 & n18612 ;
  assign n18614 = x2 | n18613 ;
  assign n18615 = ( ~n18612 & n18613 ) | ( ~n18612 & n18614 ) | ( n18613 & n18614 ) ;
  assign n18616 = n18604 & n18615 ;
  assign n18617 = n18070 | n18563 ;
  assign n18618 = ~n18564 & n18617 ;
  assign n18619 = n9798 & ~n12328 ;
  assign n18620 = n9782 & ~n12335 ;
  assign n18621 = n9783 & ~n12325 ;
  assign n18622 = n18620 | n18621 ;
  assign n18623 = n18619 | n18622 ;
  assign n18624 = n9787 | n18623 ;
  assign n18625 = ( ~n13544 & n18623 ) | ( ~n13544 & n18624 ) | ( n18623 & n18624 ) ;
  assign n18626 = ~x2 & n18625 ;
  assign n18627 = x2 | n18626 ;
  assign n18628 = ( ~n18625 & n18626 ) | ( ~n18625 & n18627 ) | ( n18626 & n18627 ) ;
  assign n18629 = n18618 & n18628 ;
  assign n18630 = ~n18559 & n18561 ;
  assign n18631 = n18562 | n18630 ;
  assign n18632 = n9798 & ~n12325 ;
  assign n18633 = n9782 & n12580 ;
  assign n18634 = n9783 & ~n12335 ;
  assign n18635 = n18633 | n18634 ;
  assign n18636 = n18632 | n18635 ;
  assign n18637 = n9787 | n18636 ;
  assign n18638 = ( ~n13720 & n18636 ) | ( ~n13720 & n18637 ) | ( n18636 & n18637 ) ;
  assign n18639 = ~x2 & n18638 ;
  assign n18640 = x2 | n18639 ;
  assign n18641 = ( ~n18638 & n18639 ) | ( ~n18638 & n18640 ) | ( n18639 & n18640 ) ;
  assign n18642 = ~n18631 & n18641 ;
  assign n18643 = n18631 & ~n18641 ;
  assign n18644 = n18642 | n18643 ;
  assign n18645 = ~n18555 & n18557 ;
  assign n18646 = n18558 | n18645 ;
  assign n18647 = n9798 & ~n12335 ;
  assign n18648 = n9782 & ~n12586 ;
  assign n18649 = n9783 & n12580 ;
  assign n18650 = n18648 | n18649 ;
  assign n18651 = n18647 | n18650 ;
  assign n18652 = n9787 & ~n13585 ;
  assign n18653 = ~n13587 & n18652 ;
  assign n18654 = ( n9787 & n18651 ) | ( n9787 & ~n18653 ) | ( n18651 & ~n18653 ) ;
  assign n18655 = ~x2 & n18654 ;
  assign n18656 = x2 | n18655 ;
  assign n18657 = ( ~n18654 & n18655 ) | ( ~n18654 & n18656 ) | ( n18655 & n18656 ) ;
  assign n18658 = ~n18646 & n18657 ;
  assign n18659 = n18646 & ~n18657 ;
  assign n18660 = n18658 | n18659 ;
  assign n18661 = n18116 | n18553 ;
  assign n18662 = ~n18554 & n18661 ;
  assign n18663 = n9798 & n12580 ;
  assign n18664 = n9782 & ~n12344 ;
  assign n18665 = n9783 & ~n12586 ;
  assign n18666 = n18664 | n18665 ;
  assign n18667 = n18663 | n18666 ;
  assign n18668 = n9787 | n18667 ;
  assign n18669 = ( n13432 & n18667 ) | ( n13432 & n18668 ) | ( n18667 & n18668 ) ;
  assign n18670 = x2 & n18669 ;
  assign n18671 = x2 & ~n18670 ;
  assign n18672 = ( n18669 & ~n18670 ) | ( n18669 & n18671 ) | ( ~n18670 & n18671 ) ;
  assign n18673 = n18662 & n18672 ;
  assign n18674 = n18662 | n18672 ;
  assign n18675 = ~n18673 & n18674 ;
  assign n18676 = ~n18549 & n18551 ;
  assign n18677 = n18552 | n18676 ;
  assign n18678 = n9798 & ~n12586 ;
  assign n18679 = n9782 & n12340 ;
  assign n18680 = n9783 & ~n12344 ;
  assign n18681 = n18679 | n18680 ;
  assign n18682 = n18678 | n18681 ;
  assign n18683 = n9787 & ~n13454 ;
  assign n18684 = ~n13455 & n18683 ;
  assign n18685 = ( n9787 & n18682 ) | ( n9787 & ~n18684 ) | ( n18682 & ~n18684 ) ;
  assign n18686 = ~x2 & n18685 ;
  assign n18687 = x2 | n18686 ;
  assign n18688 = ( ~n18685 & n18686 ) | ( ~n18685 & n18687 ) | ( n18686 & n18687 ) ;
  assign n18689 = n18677 & ~n18688 ;
  assign n18690 = ~n18677 & n18688 ;
  assign n18691 = n18689 | n18690 ;
  assign n18692 = ~n18545 & n18547 ;
  assign n18693 = n18548 | n18692 ;
  assign n18694 = n9798 & ~n12344 ;
  assign n18695 = n9782 & n12553 ;
  assign n18696 = n9783 & n12340 ;
  assign n18697 = n18695 | n18696 ;
  assign n18698 = n18694 | n18697 ;
  assign n18699 = n9787 | n18698 ;
  assign n18700 = ( ~n13523 & n18698 ) | ( ~n13523 & n18699 ) | ( n18698 & n18699 ) ;
  assign n18701 = ~x2 & n18700 ;
  assign n18702 = x2 | n18701 ;
  assign n18703 = ( ~n18700 & n18701 ) | ( ~n18700 & n18702 ) | ( n18701 & n18702 ) ;
  assign n18704 = ~n18693 & n18703 ;
  assign n18705 = ~n18691 & n18704 ;
  assign n18706 = n18690 | n18705 ;
  assign n18707 = n18693 | n18704 ;
  assign n18708 = ( ~n18703 & n18704 ) | ( ~n18703 & n18707 ) | ( n18704 & n18707 ) ;
  assign n18709 = n18171 | n18173 ;
  assign n18710 = n18543 | n18709 ;
  assign n18711 = ~n18544 & n18710 ;
  assign n18712 = n18188 | n18538 ;
  assign n18713 = ~n18539 & n18712 ;
  assign n18714 = n9798 & n12355 ;
  assign n18715 = n9782 & ~n12537 ;
  assign n18716 = n9783 & n12351 ;
  assign n18717 = n18715 | n18716 ;
  assign n18718 = n18714 | n18717 ;
  assign n18719 = n9787 | n18718 ;
  assign n18720 = ( n13409 & n18718 ) | ( n13409 & n18719 ) | ( n18718 & n18719 ) ;
  assign n18721 = x2 & n18720 ;
  assign n18722 = x2 & ~n18721 ;
  assign n18723 = ( n18720 & ~n18721 ) | ( n18720 & n18722 ) | ( ~n18721 & n18722 ) ;
  assign n18724 = n9798 & n12351 ;
  assign n18725 = n9782 & n12364 ;
  assign n18726 = n9783 & ~n12537 ;
  assign n18727 = n18725 | n18726 ;
  assign n18728 = n18724 | n18727 ;
  assign n18729 = n9787 & n12928 ;
  assign n18730 = ~n12925 & n18729 ;
  assign n18731 = ( n9787 & n18728 ) | ( n9787 & ~n18730 ) | ( n18728 & ~n18730 ) ;
  assign n18732 = x2 & n18731 ;
  assign n18733 = x2 & ~n18732 ;
  assign n18734 = ( n18731 & ~n18732 ) | ( n18731 & n18733 ) | ( ~n18732 & n18733 ) ;
  assign n18735 = n18224 | n18530 ;
  assign n18736 = ~n18531 & n18735 ;
  assign n18737 = ( n18226 & n18529 ) | ( n18226 & ~n18530 ) | ( n18529 & ~n18530 ) ;
  assign n18738 = ( n18237 & ~n18530 ) | ( n18237 & n18737 ) | ( ~n18530 & n18737 ) ;
  assign n18739 = ( n18239 & n18528 ) | ( n18239 & ~n18529 ) | ( n18528 & ~n18529 ) ;
  assign n18740 = ( n18249 & ~n18529 ) | ( n18249 & n18739 ) | ( ~n18529 & n18739 ) ;
  assign n18741 = n9798 & n12520 ;
  assign n18742 = n9782 & ~n12371 ;
  assign n18743 = n9783 & n12375 ;
  assign n18744 = n18742 | n18743 ;
  assign n18745 = n18741 | n18744 ;
  assign n18746 = n9787 & ~n12837 ;
  assign n18747 = ~n12835 & n18746 ;
  assign n18748 = ( n9787 & n18745 ) | ( n9787 & ~n18747 ) | ( n18745 & ~n18747 ) ;
  assign n18749 = ~x2 & n18748 ;
  assign n18750 = x2 | n18749 ;
  assign n18751 = ( ~n18748 & n18749 ) | ( ~n18748 & n18750 ) | ( n18749 & n18750 ) ;
  assign n18752 = n9798 & n12375 ;
  assign n18753 = n9782 & n12378 ;
  assign n18754 = n9783 & ~n12371 ;
  assign n18755 = n18753 | n18754 ;
  assign n18756 = n18752 | n18755 ;
  assign n18757 = n9787 & n13065 ;
  assign n18758 = ~n13064 & n18757 ;
  assign n18759 = ( n9787 & n18756 ) | ( n9787 & ~n18758 ) | ( n18756 & ~n18758 ) ;
  assign n18760 = x2 & n18759 ;
  assign n18761 = x2 & ~n18760 ;
  assign n18762 = ( n18759 & ~n18760 ) | ( n18759 & n18761 ) | ( ~n18760 & n18761 ) ;
  assign n18763 = n9798 & ~n12371 ;
  assign n18764 = n9782 & ~n12502 ;
  assign n18765 = n9783 & n12378 ;
  assign n18766 = n18764 | n18765 ;
  assign n18767 = n18763 | n18766 ;
  assign n18768 = n9787 | n18767 ;
  assign n18769 = ( ~n12848 & n18767 ) | ( ~n12848 & n18768 ) | ( n18767 & n18768 ) ;
  assign n18770 = ~x2 & n18769 ;
  assign n18771 = x2 | n18770 ;
  assign n18772 = ( ~n18769 & n18770 ) | ( ~n18769 & n18771 ) | ( n18770 & n18771 ) ;
  assign n18773 = n18314 | n18316 ;
  assign n18774 = n18523 | n18773 ;
  assign n18775 = ~n18524 & n18774 ;
  assign n18776 = ( ~n18520 & n18521 ) | ( ~n18520 & n18522 ) | ( n18521 & n18522 ) ;
  assign n18777 = n18520 | n18776 ;
  assign n18778 = ~n18523 & n18777 ;
  assign n18779 = n18345 | n18514 ;
  assign n18780 = ~n18515 & n18779 ;
  assign n18781 = n9798 & n12392 ;
  assign n18782 = n9782 & n12415 ;
  assign n18783 = n9783 & n12401 ;
  assign n18784 = n18782 | n18783 ;
  assign n18785 = n18781 | n18784 ;
  assign n18786 = n9787 | n18785 ;
  assign n18787 = ( n13034 & n18785 ) | ( n13034 & n18786 ) | ( n18785 & n18786 ) ;
  assign n18788 = x2 & n18787 ;
  assign n18789 = x2 & ~n18788 ;
  assign n18790 = ( n18787 & ~n18788 ) | ( n18787 & n18789 ) | ( ~n18788 & n18789 ) ;
  assign n18791 = n9798 & n12401 ;
  assign n18792 = n9782 & n12411 ;
  assign n18793 = n9783 & n12415 ;
  assign n18794 = n18792 | n18793 ;
  assign n18795 = n18791 | n18794 ;
  assign n18796 = n9787 & ~n13163 ;
  assign n18797 = ~n13161 & n18796 ;
  assign n18798 = ( n9787 & n18795 ) | ( n9787 & ~n18797 ) | ( n18795 & ~n18797 ) ;
  assign n18799 = ~x2 & n18798 ;
  assign n18800 = x2 | n18799 ;
  assign n18801 = ( ~n18798 & n18799 ) | ( ~n18798 & n18800 ) | ( n18799 & n18800 ) ;
  assign n18802 = n18504 | n18506 ;
  assign n18803 = ~n18507 & n18802 ;
  assign n18804 = n18394 | n18502 ;
  assign n18805 = ~n18503 & n18804 ;
  assign n18806 = ( n18396 & n18501 ) | ( n18396 & ~n18502 ) | ( n18501 & ~n18502 ) ;
  assign n18807 = ( n18407 & ~n18502 ) | ( n18407 & n18806 ) | ( ~n18502 & n18806 ) ;
  assign n18808 = n18434 | n18498 ;
  assign n18809 = ~n18499 & n18808 ;
  assign n18810 = n9798 & ~n12438 ;
  assign n18811 = n9782 & n12446 ;
  assign n18812 = n9783 & n12440 ;
  assign n18813 = n18811 | n18812 ;
  assign n18814 = n18810 | n18813 ;
  assign n18815 = n9787 & n14154 ;
  assign n18816 = ~n14156 & n18815 ;
  assign n18817 = ( n9787 & n18814 ) | ( n9787 & ~n18816 ) | ( n18814 & ~n18816 ) ;
  assign n18818 = x2 & n18817 ;
  assign n18819 = x2 & ~n18818 ;
  assign n18820 = ( n18817 & ~n18818 ) | ( n18817 & n18819 ) | ( ~n18818 & n18819 ) ;
  assign n18821 = n18449 | n18483 ;
  assign n18822 = ~n18484 & n18821 ;
  assign n18823 = n18450 | n18472 ;
  assign n18824 = n18450 & n18472 ;
  assign n18825 = n18823 & ~n18824 ;
  assign n18826 = ~n18482 & n18825 ;
  assign n18827 = n9798 & n12446 ;
  assign n18828 = n9782 & n12454 ;
  assign n18829 = n9783 & n12452 ;
  assign n18830 = n18828 | n18829 ;
  assign n18831 = n18827 | n18830 ;
  assign n18832 = n9787 | n18831 ;
  assign n18833 = ( n13862 & n18831 ) | ( n13862 & n18832 ) | ( n18831 & n18832 ) ;
  assign n18834 = x2 & n18833 ;
  assign n18835 = x2 & ~n18834 ;
  assign n18836 = ( n18833 & ~n18834 ) | ( n18833 & n18835 ) | ( ~n18834 & n18835 ) ;
  assign n18837 = n8678 & ~n12468 ;
  assign n18838 = n10020 & n13994 ;
  assign n18839 = n10033 & ~n12468 ;
  assign n18840 = ( x2 & n10031 ) | ( x2 & n12466 ) | ( n10031 & n12466 ) ;
  assign n18841 = ~n18839 & n18840 ;
  assign n18842 = ~n18838 & n18841 ;
  assign n18843 = n9782 & ~n12468 ;
  assign n18844 = n9783 & ~n12466 ;
  assign n18845 = n18843 | n18844 ;
  assign n18846 = n9798 & n12459 ;
  assign n18847 = x2 & n18846 ;
  assign n18848 = ( x2 & n18845 ) | ( x2 & n18847 ) | ( n18845 & n18847 ) ;
  assign n18849 = n18842 & ~n18848 ;
  assign n18850 = x0 & ~n12468 ;
  assign n18851 = n10020 & n14003 ;
  assign n18852 = n18850 | n18851 ;
  assign n18853 = n18849 & ~n18852 ;
  assign n18854 = n9798 & ~n12456 ;
  assign n18855 = n9782 & ~n12466 ;
  assign n18856 = n9783 & n12459 ;
  assign n18857 = n18855 | n18856 ;
  assign n18858 = n18854 | n18857 ;
  assign n18859 = n9787 | n18858 ;
  assign n18860 = ( n14031 & n18858 ) | ( n14031 & n18859 ) | ( n18858 & n18859 ) ;
  assign n18861 = x2 & n18860 ;
  assign n18862 = x2 & ~n18861 ;
  assign n18863 = ( n18860 & ~n18861 ) | ( n18860 & n18862 ) | ( ~n18861 & n18862 ) ;
  assign n18864 = ( n18837 & n18853 ) | ( n18837 & n18863 ) | ( n18853 & n18863 ) ;
  assign n18865 = n9798 & n12454 ;
  assign n18866 = n9782 & n12459 ;
  assign n18867 = n9783 & ~n12456 ;
  assign n18868 = n18866 | n18867 ;
  assign n18869 = n18865 | n18868 ;
  assign n18870 = n9787 | n18869 ;
  assign n18871 = ( n14041 & n18869 ) | ( n14041 & n18870 ) | ( n18869 & n18870 ) ;
  assign n18872 = x2 & n18871 ;
  assign n18873 = x2 & ~n18872 ;
  assign n18874 = ( n18871 & ~n18872 ) | ( n18871 & n18873 ) | ( ~n18872 & n18873 ) ;
  assign n18875 = n18864 | n18874 ;
  assign n18876 = n18452 | n18460 ;
  assign n18877 = ~n18461 & n18876 ;
  assign n18878 = n18875 & n18877 ;
  assign n18879 = n18461 | n18471 ;
  assign n18880 = ~n18472 & n18879 ;
  assign n18881 = n18864 & n18874 ;
  assign n18882 = n18880 & n18881 ;
  assign n18883 = ( n18878 & n18880 ) | ( n18878 & n18882 ) | ( n18880 & n18882 ) ;
  assign n18884 = n18836 | n18883 ;
  assign n18885 = n9798 & n12452 ;
  assign n18886 = n9782 & ~n12456 ;
  assign n18887 = n9783 & n12454 ;
  assign n18888 = n18886 | n18887 ;
  assign n18889 = n18885 | n18888 ;
  assign n18890 = n9787 | n18889 ;
  assign n18891 = ( ~n13922 & n18889 ) | ( ~n13922 & n18890 ) | ( n18889 & n18890 ) ;
  assign n18892 = ~x2 & n18891 ;
  assign n18893 = n18880 | n18881 ;
  assign n18894 = n18878 | n18893 ;
  assign n18895 = ( ~n18891 & n18892 ) | ( ~n18891 & n18894 ) | ( n18892 & n18894 ) ;
  assign n18896 = ( x2 & n18892 ) | ( x2 & n18895 ) | ( n18892 & n18895 ) ;
  assign n18897 = n18884 | n18896 ;
  assign n18898 = ( n18482 & n18826 ) | ( n18482 & n18897 ) | ( n18826 & n18897 ) ;
  assign n18899 = ( ~n18825 & n18826 ) | ( ~n18825 & n18898 ) | ( n18826 & n18898 ) ;
  assign n18900 = n18836 & n18883 ;
  assign n18901 = ( n18836 & n18896 ) | ( n18836 & n18900 ) | ( n18896 & n18900 ) ;
  assign n18902 = n18822 & n18901 ;
  assign n18903 = ( n18822 & n18899 ) | ( n18822 & n18902 ) | ( n18899 & n18902 ) ;
  assign n18904 = n18820 & n18903 ;
  assign n18905 = n9798 & n12440 ;
  assign n18906 = n9782 & n12452 ;
  assign n18907 = n9783 & n12446 ;
  assign n18908 = n18906 | n18907 ;
  assign n18909 = n18905 | n18908 ;
  assign n18910 = n9787 | n18909 ;
  assign n18911 = ( n13822 & n18909 ) | ( n13822 & n18910 ) | ( n18909 & n18910 ) ;
  assign n18912 = ~x2 & n18911 ;
  assign n18913 = n18822 | n18901 ;
  assign n18914 = n18899 | n18913 ;
  assign n18915 = ( ~n18911 & n18912 ) | ( ~n18911 & n18914 ) | ( n18912 & n18914 ) ;
  assign n18916 = ( x2 & n18912 ) | ( x2 & n18915 ) | ( n18912 & n18915 ) ;
  assign n18917 = ( n18820 & n18904 ) | ( n18820 & n18916 ) | ( n18904 & n18916 ) ;
  assign n18918 = n9798 & n12433 ;
  assign n18919 = n9782 & n12440 ;
  assign n18920 = n9783 & ~n12438 ;
  assign n18921 = n18919 | n18920 ;
  assign n18922 = n18918 | n18921 ;
  assign n18923 = n9787 | n18922 ;
  assign n18924 = ( ~n14167 & n18922 ) | ( ~n14167 & n18923 ) | ( n18922 & n18923 ) ;
  assign n18925 = ~x2 & n18924 ;
  assign n18926 = x2 | n18925 ;
  assign n18927 = ( ~n18924 & n18925 ) | ( ~n18924 & n18926 ) | ( n18925 & n18926 ) ;
  assign n18928 = n18917 | n18927 ;
  assign n18929 = n18820 | n18903 ;
  assign n18930 = n18916 | n18929 ;
  assign n18931 = ( n18485 & ~n18495 ) | ( n18485 & n18497 ) | ( ~n18495 & n18497 ) ;
  assign n18932 = ( ~n18485 & n18495 ) | ( ~n18485 & n18497 ) | ( n18495 & n18497 ) ;
  assign n18933 = ( ~n18497 & n18931 ) | ( ~n18497 & n18932 ) | ( n18931 & n18932 ) ;
  assign n18934 = n18930 & n18933 ;
  assign n18935 = n18928 | n18934 ;
  assign n18936 = n18809 & n18935 ;
  assign n18937 = n9798 & ~n12423 ;
  assign n18938 = n9782 & ~n12438 ;
  assign n18939 = n9783 & n12433 ;
  assign n18940 = n18938 | n18939 ;
  assign n18941 = n18937 | n18940 ;
  assign n18942 = n9787 | n18941 ;
  assign n18943 = ( ~n13786 & n18941 ) | ( ~n13786 & n18942 ) | ( n18941 & n18942 ) ;
  assign n18944 = ~x2 & n18943 ;
  assign n18945 = x2 | n18944 ;
  assign n18946 = ( ~n18943 & n18944 ) | ( ~n18943 & n18945 ) | ( n18944 & n18945 ) ;
  assign n18947 = n18917 & n18927 ;
  assign n18948 = ( n18927 & n18934 ) | ( n18927 & n18947 ) | ( n18934 & n18947 ) ;
  assign n18949 = n18946 & n18948 ;
  assign n18950 = ( n18936 & n18946 ) | ( n18936 & n18949 ) | ( n18946 & n18949 ) ;
  assign n18951 = n18807 & n18950 ;
  assign n18952 = n18946 | n18948 ;
  assign n18953 = n18936 | n18952 ;
  assign n18954 = ( ~n18409 & n18419 ) | ( ~n18409 & n18500 ) | ( n18419 & n18500 ) ;
  assign n18955 = ( n18409 & ~n18419 ) | ( n18409 & n18500 ) | ( ~n18419 & n18500 ) ;
  assign n18956 = ( ~n18500 & n18954 ) | ( ~n18500 & n18955 ) | ( n18954 & n18955 ) ;
  assign n18957 = n18953 & n18956 ;
  assign n18958 = ( n18807 & n18951 ) | ( n18807 & n18957 ) | ( n18951 & n18957 ) ;
  assign n18959 = n18805 & n18958 ;
  assign n18960 = n9798 & n12419 ;
  assign n18961 = n9782 & n12433 ;
  assign n18962 = n9783 & ~n12423 ;
  assign n18963 = n18961 | n18962 ;
  assign n18964 = n18960 | n18963 ;
  assign n18965 = n9787 | n18964 ;
  assign n18966 = ( ~n13282 & n18964 ) | ( ~n13282 & n18965 ) | ( n18964 & n18965 ) ;
  assign n18967 = ~x2 & n18966 ;
  assign n18968 = n18807 | n18950 ;
  assign n18969 = n18957 | n18968 ;
  assign n18970 = ( ~n18966 & n18967 ) | ( ~n18966 & n18969 ) | ( n18967 & n18969 ) ;
  assign n18971 = ( x2 & n18967 ) | ( x2 & n18970 ) | ( n18967 & n18970 ) ;
  assign n18972 = ( n18805 & n18959 ) | ( n18805 & n18971 ) | ( n18959 & n18971 ) ;
  assign n18973 = n18803 & n18972 ;
  assign n18974 = n9798 & n12411 ;
  assign n18975 = n9782 & ~n12423 ;
  assign n18976 = n9783 & n12419 ;
  assign n18977 = n18975 | n18976 ;
  assign n18978 = n18974 | n18977 ;
  assign n18979 = n9787 | n18978 ;
  assign n18980 = ( n13776 & n18978 ) | ( n13776 & n18979 ) | ( n18978 & n18979 ) ;
  assign n18981 = ~x2 & n18980 ;
  assign n18982 = n18805 | n18958 ;
  assign n18983 = n18971 | n18982 ;
  assign n18984 = ( ~n18980 & n18981 ) | ( ~n18980 & n18983 ) | ( n18981 & n18983 ) ;
  assign n18985 = ( x2 & n18981 ) | ( x2 & n18984 ) | ( n18981 & n18984 ) ;
  assign n18986 = ( n18803 & n18973 ) | ( n18803 & n18985 ) | ( n18973 & n18985 ) ;
  assign n18987 = n18801 & n18986 ;
  assign n18988 = n9798 & n12415 ;
  assign n18989 = n9782 & n12419 ;
  assign n18990 = n9783 & n12411 ;
  assign n18991 = n18989 | n18990 ;
  assign n18992 = n18988 | n18991 ;
  assign n18993 = ( n9787 & n13761 ) | ( n9787 & n13762 ) | ( n13761 & n13762 ) ;
  assign n18994 = n18992 | n18993 ;
  assign n18995 = x2 & n18994 ;
  assign n18996 = n18803 | n18972 ;
  assign n18997 = n18985 | n18996 ;
  assign n18998 = ( x2 & n18994 ) | ( x2 & n18997 ) | ( n18994 & n18997 ) ;
  assign n18999 = ~n18995 & n18998 ;
  assign n19000 = ( n18801 & n18987 ) | ( n18801 & n18999 ) | ( n18987 & n18999 ) ;
  assign n19001 = n18790 & n19000 ;
  assign n19002 = n18801 | n18986 ;
  assign n19003 = n18999 | n19002 ;
  assign n19004 = ( n18365 & n18508 ) | ( n18365 & ~n18510 ) | ( n18508 & ~n18510 ) ;
  assign n19005 = ( ~n18365 & n18508 ) | ( ~n18365 & n18510 ) | ( n18508 & n18510 ) ;
  assign n19006 = ( ~n18508 & n19004 ) | ( ~n18508 & n19005 ) | ( n19004 & n19005 ) ;
  assign n19007 = n19003 & n19006 ;
  assign n19008 = ( n18790 & n19001 ) | ( n18790 & n19007 ) | ( n19001 & n19007 ) ;
  assign n19009 = n9798 & n12383 ;
  assign n19010 = n9782 & n12401 ;
  assign n19011 = n9783 & n12392 ;
  assign n19012 = n19010 | n19011 ;
  assign n19013 = n19009 | n19012 ;
  assign n19014 = n9787 | n19013 ;
  assign n19015 = ( n13141 & n19013 ) | ( n13141 & n19014 ) | ( n19013 & n19014 ) ;
  assign n19016 = x2 & n19015 ;
  assign n19017 = x2 & ~n19016 ;
  assign n19018 = ( n19015 & ~n19016 ) | ( n19015 & n19017 ) | ( ~n19016 & n19017 ) ;
  assign n19019 = n19008 | n19018 ;
  assign n19020 = n18790 | n19000 ;
  assign n19021 = n19007 | n19020 ;
  assign n19022 = ( n18355 & n18511 ) | ( n18355 & ~n18513 ) | ( n18511 & ~n18513 ) ;
  assign n19023 = ( ~n18355 & n18511 ) | ( ~n18355 & n18513 ) | ( n18511 & n18513 ) ;
  assign n19024 = ( ~n18511 & n19022 ) | ( ~n18511 & n19023 ) | ( n19022 & n19023 ) ;
  assign n19025 = n19021 & n19024 ;
  assign n19026 = n19019 | n19025 ;
  assign n19027 = n18780 & n19026 ;
  assign n19028 = ( ~n18516 & n18517 ) | ( ~n18516 & n18518 ) | ( n18517 & n18518 ) ;
  assign n19029 = n18516 | n19028 ;
  assign n19030 = ~n18519 & n19029 ;
  assign n19031 = n19008 & n19018 ;
  assign n19032 = ( n19018 & n19025 ) | ( n19018 & n19031 ) | ( n19025 & n19031 ) ;
  assign n19033 = n19030 & n19032 ;
  assign n19034 = ( n19027 & n19030 ) | ( n19027 & n19033 ) | ( n19030 & n19033 ) ;
  assign n19035 = n18778 & n19034 ;
  assign n19036 = n9798 & n12387 ;
  assign n19037 = n9782 & n12392 ;
  assign n19038 = n9783 & n12383 ;
  assign n19039 = n19037 | n19038 ;
  assign n19040 = n19036 | n19039 ;
  assign n19041 = n9787 | n19040 ;
  assign n19042 = ( n12948 & n19040 ) | ( n12948 & n19041 ) | ( n19040 & n19041 ) ;
  assign n19043 = ~x2 & n19042 ;
  assign n19044 = n19030 | n19032 ;
  assign n19045 = n19027 | n19044 ;
  assign n19046 = ( ~n19042 & n19043 ) | ( ~n19042 & n19045 ) | ( n19043 & n19045 ) ;
  assign n19047 = ( x2 & n19043 ) | ( x2 & n19046 ) | ( n19043 & n19046 ) ;
  assign n19048 = ( n18778 & n19035 ) | ( n18778 & n19047 ) | ( n19035 & n19047 ) ;
  assign n19049 = n18775 & n19048 ;
  assign n19050 = n9798 & ~n12502 ;
  assign n19051 = n9782 & n12383 ;
  assign n19052 = n9783 & n12387 ;
  assign n19053 = n19051 | n19052 ;
  assign n19054 = n19050 | n19053 ;
  assign n19055 = n9787 | n19054 ;
  assign n19056 = ( ~n12756 & n19054 ) | ( ~n12756 & n19055 ) | ( n19054 & n19055 ) ;
  assign n19057 = ~x2 & n19056 ;
  assign n19058 = n18778 | n19034 ;
  assign n19059 = n19047 | n19058 ;
  assign n19060 = ( ~n19056 & n19057 ) | ( ~n19056 & n19059 ) | ( n19057 & n19059 ) ;
  assign n19061 = ( x2 & n19057 ) | ( x2 & n19060 ) | ( n19057 & n19060 ) ;
  assign n19062 = ( n18775 & n19049 ) | ( n18775 & n19061 ) | ( n19049 & n19061 ) ;
  assign n19063 = n18772 & n19062 ;
  assign n19064 = n9798 & n12378 ;
  assign n19065 = n9782 & n12387 ;
  assign n19066 = n9783 & ~n12502 ;
  assign n19067 = n19065 | n19066 ;
  assign n19068 = n19064 | n19067 ;
  assign n19069 = n9787 | n19068 ;
  assign n19070 = ( ~n12816 & n19068 ) | ( ~n12816 & n19069 ) | ( n19068 & n19069 ) ;
  assign n19071 = ~x2 & n19070 ;
  assign n19072 = n18775 | n19048 ;
  assign n19073 = n19061 | n19072 ;
  assign n19074 = ( ~n19070 & n19071 ) | ( ~n19070 & n19073 ) | ( n19071 & n19073 ) ;
  assign n19075 = ( x2 & n19071 ) | ( x2 & n19074 ) | ( n19071 & n19074 ) ;
  assign n19076 = ( n18772 & n19063 ) | ( n18772 & n19075 ) | ( n19063 & n19075 ) ;
  assign n19077 = n18762 & n19076 ;
  assign n19078 = n18772 | n19062 ;
  assign n19079 = n19075 | n19078 ;
  assign n19080 = ( ~n18278 & n18288 ) | ( ~n18278 & n18525 ) | ( n18288 & n18525 ) ;
  assign n19081 = ( n18278 & ~n18288 ) | ( n18278 & n18525 ) | ( ~n18288 & n18525 ) ;
  assign n19082 = ( ~n18525 & n19080 ) | ( ~n18525 & n19081 ) | ( n19080 & n19081 ) ;
  assign n19083 = n19079 & n19082 ;
  assign n19084 = ( n18762 & n19077 ) | ( n18762 & n19083 ) | ( n19077 & n19083 ) ;
  assign n19085 = n18751 & n19084 ;
  assign n19086 = n18762 | n19076 ;
  assign n19087 = n19083 | n19086 ;
  assign n19088 = ( ~n18265 & n18275 ) | ( ~n18265 & n18526 ) | ( n18275 & n18526 ) ;
  assign n19089 = ( n18265 & ~n18275 ) | ( n18265 & n18526 ) | ( ~n18275 & n18526 ) ;
  assign n19090 = ( ~n18526 & n19088 ) | ( ~n18526 & n19089 ) | ( n19088 & n19089 ) ;
  assign n19091 = n19087 & n19090 ;
  assign n19092 = ( n18751 & n19085 ) | ( n18751 & n19091 ) | ( n19085 & n19091 ) ;
  assign n19093 = n18740 & n19092 ;
  assign n19094 = n18751 | n19084 ;
  assign n19095 = n19091 | n19094 ;
  assign n19096 = ( ~n18252 & n18262 ) | ( ~n18252 & n18527 ) | ( n18262 & n18527 ) ;
  assign n19097 = ( n18252 & ~n18262 ) | ( n18252 & n18527 ) | ( ~n18262 & n18527 ) ;
  assign n19098 = ( ~n18527 & n19096 ) | ( ~n18527 & n19097 ) | ( n19096 & n19097 ) ;
  assign n19099 = n19095 & n19098 ;
  assign n19100 = ( n18740 & n19093 ) | ( n18740 & n19099 ) | ( n19093 & n19099 ) ;
  assign n19101 = n18738 & n19100 ;
  assign n19102 = n9798 & ~n12360 ;
  assign n19103 = n9782 & n12375 ;
  assign n19104 = n9783 & n12520 ;
  assign n19105 = n19103 | n19104 ;
  assign n19106 = n19102 | n19105 ;
  assign n19107 = n9787 | n19106 ;
  assign n19108 = ( ~n12902 & n19106 ) | ( ~n12902 & n19107 ) | ( n19106 & n19107 ) ;
  assign n19109 = ~x2 & n19108 ;
  assign n19110 = n18740 | n19092 ;
  assign n19111 = n19099 | n19110 ;
  assign n19112 = ( ~n19108 & n19109 ) | ( ~n19108 & n19111 ) | ( n19109 & n19111 ) ;
  assign n19113 = ( x2 & n19109 ) | ( x2 & n19112 ) | ( n19109 & n19112 ) ;
  assign n19114 = ( n18738 & n19101 ) | ( n18738 & n19113 ) | ( n19101 & n19113 ) ;
  assign n19115 = n18736 & n19114 ;
  assign n19116 = n9798 & n12364 ;
  assign n19117 = n9782 & n12520 ;
  assign n19118 = n9783 & ~n12360 ;
  assign n19119 = n19117 | n19118 ;
  assign n19120 = n19116 | n19119 ;
  assign n19121 = n9787 | n19120 ;
  assign n19122 = ( ~n13113 & n19120 ) | ( ~n13113 & n19121 ) | ( n19120 & n19121 ) ;
  assign n19123 = ~x2 & n19122 ;
  assign n19124 = n18738 | n19100 ;
  assign n19125 = n19113 | n19124 ;
  assign n19126 = ( ~n19122 & n19123 ) | ( ~n19122 & n19125 ) | ( n19123 & n19125 ) ;
  assign n19127 = ( x2 & n19123 ) | ( x2 & n19126 ) | ( n19123 & n19126 ) ;
  assign n19128 = ( n18736 & n19115 ) | ( n18736 & n19127 ) | ( n19115 & n19127 ) ;
  assign n19129 = n18734 & n19128 ;
  assign n19130 = n9798 & ~n12537 ;
  assign n19131 = n9782 & ~n12360 ;
  assign n19132 = n9783 & n12364 ;
  assign n19133 = n19131 | n19132 ;
  assign n19134 = n19130 | n19133 ;
  assign n19135 = ( n9787 & n13081 ) | ( n9787 & ~n13082 ) | ( n13081 & ~n13082 ) ;
  assign n19136 = n19134 | n19135 ;
  assign n19137 = x2 & n19136 ;
  assign n19138 = n18736 | n19114 ;
  assign n19139 = n19127 | n19138 ;
  assign n19140 = ( x2 & n19136 ) | ( x2 & n19139 ) | ( n19136 & n19139 ) ;
  assign n19141 = ~n19137 & n19140 ;
  assign n19142 = ( n18734 & n19129 ) | ( n18734 & n19141 ) | ( n19129 & n19141 ) ;
  assign n19143 = n18723 & n19142 ;
  assign n19144 = n18734 | n19128 ;
  assign n19145 = n19141 | n19144 ;
  assign n19146 = ( n18208 & n18532 ) | ( n18208 & ~n18534 ) | ( n18532 & ~n18534 ) ;
  assign n19147 = ( ~n18208 & n18532 ) | ( ~n18208 & n18534 ) | ( n18532 & n18534 ) ;
  assign n19148 = ( ~n18532 & n19146 ) | ( ~n18532 & n19147 ) | ( n19146 & n19147 ) ;
  assign n19149 = n19145 & n19148 ;
  assign n19150 = ( n18723 & n19143 ) | ( n18723 & n19149 ) | ( n19143 & n19149 ) ;
  assign n19151 = n9798 & n12558 ;
  assign n19152 = n9782 & n12351 ;
  assign n19153 = n9783 & n12355 ;
  assign n19154 = n19152 | n19153 ;
  assign n19155 = n19151 | n19154 ;
  assign n19156 = n9787 | n19155 ;
  assign n19157 = ( n13330 & n19155 ) | ( n13330 & n19156 ) | ( n19155 & n19156 ) ;
  assign n19158 = x2 & n19157 ;
  assign n19159 = x2 & ~n19158 ;
  assign n19160 = ( n19157 & ~n19158 ) | ( n19157 & n19159 ) | ( ~n19158 & n19159 ) ;
  assign n19161 = n19150 | n19160 ;
  assign n19162 = n18723 | n19142 ;
  assign n19163 = n19149 | n19162 ;
  assign n19164 = ( n18198 & n18535 ) | ( n18198 & ~n18537 ) | ( n18535 & ~n18537 ) ;
  assign n19165 = ( ~n18198 & n18535 ) | ( ~n18198 & n18537 ) | ( n18535 & n18537 ) ;
  assign n19166 = ( ~n18535 & n19164 ) | ( ~n18535 & n19165 ) | ( n19164 & n19165 ) ;
  assign n19167 = n19163 & n19166 ;
  assign n19168 = n19161 | n19167 ;
  assign n19169 = n18713 & n19168 ;
  assign n19170 = ( ~n18540 & n18541 ) | ( ~n18540 & n18542 ) | ( n18541 & n18542 ) ;
  assign n19171 = n18540 | n19170 ;
  assign n19172 = ~n18543 & n19171 ;
  assign n19173 = n19150 & n19160 ;
  assign n19174 = ( n19160 & n19167 ) | ( n19160 & n19173 ) | ( n19167 & n19173 ) ;
  assign n19175 = n19172 & n19174 ;
  assign n19176 = ( n19169 & n19172 ) | ( n19169 & n19175 ) | ( n19172 & n19175 ) ;
  assign n19177 = n18711 & n19176 ;
  assign n19178 = n9798 & n12553 ;
  assign n19179 = n9782 & n12355 ;
  assign n19180 = n9783 & n12558 ;
  assign n19181 = n19179 | n19180 ;
  assign n19182 = n19178 | n19181 ;
  assign n19183 = n9787 | n19182 ;
  assign n19184 = ( n13097 & n19182 ) | ( n13097 & n19183 ) | ( n19182 & n19183 ) ;
  assign n19185 = ~x2 & n19184 ;
  assign n19186 = n19172 | n19174 ;
  assign n19187 = n19169 | n19186 ;
  assign n19188 = ( ~n19184 & n19185 ) | ( ~n19184 & n19187 ) | ( n19185 & n19187 ) ;
  assign n19189 = ( x2 & n19185 ) | ( x2 & n19188 ) | ( n19185 & n19188 ) ;
  assign n19190 = ( n18711 & n19177 ) | ( n18711 & n19189 ) | ( n19177 & n19189 ) ;
  assign n19191 = n9787 & n13347 ;
  assign n19192 = ( n9787 & n13346 ) | ( n9787 & n19191 ) | ( n13346 & n19191 ) ;
  assign n19193 = n9798 & n12340 ;
  assign n19194 = n9782 & n12558 ;
  assign n19195 = n9783 & n12553 ;
  assign n19196 = n19194 | n19195 ;
  assign n19197 = n19193 | n19196 ;
  assign n19198 = n19192 | n19197 ;
  assign n19199 = n18711 | n19176 ;
  assign n19200 = n19189 | n19199 ;
  assign n19201 = ( x2 & n19198 ) | ( x2 & ~n19200 ) | ( n19198 & ~n19200 ) ;
  assign n19202 = x2 | n19198 ;
  assign n19203 = ( n19190 & ~n19201 ) | ( n19190 & n19202 ) | ( ~n19201 & n19202 ) ;
  assign n19204 = ~n18708 & n19203 ;
  assign n19205 = ( ~n18689 & n18706 ) | ( ~n18689 & n19204 ) | ( n18706 & n19204 ) ;
  assign n19206 = n18675 & n19205 ;
  assign n19207 = n18673 | n19206 ;
  assign n19208 = ~n18660 & n19207 ;
  assign n19209 = n18658 | n19208 ;
  assign n19210 = ~n18644 & n19209 ;
  assign n19211 = n18642 | n19210 ;
  assign n19212 = n18618 | n18628 ;
  assign n19213 = ~n18629 & n19212 ;
  assign n19214 = n19211 & n19213 ;
  assign n19215 = n18629 | n19214 ;
  assign n19216 = n18604 | n18615 ;
  assign n19217 = ~n18616 & n19216 ;
  assign n19218 = n19215 & n19217 ;
  assign n19219 = n18616 | n19218 ;
  assign n19220 = n18591 | n18601 ;
  assign n19221 = ~n18602 & n19220 ;
  assign n19222 = n19219 & n19221 ;
  assign n19223 = n18602 | n19222 ;
  assign n19224 = n18589 & n19223 ;
  assign n19225 = n18571 | n18573 ;
  assign n19226 = ~n18574 & n19225 ;
  assign n19227 = ( n18587 & n19224 ) | ( n18587 & n19226 ) | ( n19224 & n19226 ) ;
  assign n19228 = ~n17973 & n18002 ;
  assign n19229 = n18003 | n19228 ;
  assign n19230 = ( n18574 & n19227 ) | ( n18574 & ~n19229 ) | ( n19227 & ~n19229 ) ;
  assign n19231 = n18003 | n19230 ;
  assign n19232 = n16847 | n16850 ;
  assign n19233 = ( ~n16849 & n16850 ) | ( ~n16849 & n19232 ) | ( n16850 & n19232 ) ;
  assign n19234 = n8681 & ~n12318 ;
  assign n19235 = n8680 & n12608 ;
  assign n19236 = n19234 | n19235 ;
  assign n19237 = n9245 & ~n12314 ;
  assign n19238 = n19236 | n19237 ;
  assign n19239 = n8685 | n19238 ;
  assign n19240 = ( ~n14302 & n19238 ) | ( ~n14302 & n19239 ) | ( n19238 & n19239 ) ;
  assign n19241 = ~x5 & n19240 ;
  assign n19242 = x5 | n19241 ;
  assign n19243 = ( ~n19240 & n19241 ) | ( ~n19240 & n19242 ) | ( n19241 & n19242 ) ;
  assign n19244 = ( ~n16831 & n16841 ) | ( ~n16831 & n16844 ) | ( n16841 & n16844 ) ;
  assign n19245 = ( n16831 & ~n16844 ) | ( n16831 & n19244 ) | ( ~n16844 & n19244 ) ;
  assign n19246 = ( ~n16841 & n19244 ) | ( ~n16841 & n19245 ) | ( n19244 & n19245 ) ;
  assign n19247 = ( n17998 & n19243 ) | ( n17998 & n19246 ) | ( n19243 & n19246 ) ;
  assign n19248 = ~n19233 & n19247 ;
  assign n19249 = ( ~n17998 & n19243 ) | ( ~n17998 & n19246 ) | ( n19243 & n19246 ) ;
  assign n19250 = ( n17998 & ~n19246 ) | ( n17998 & n19249 ) | ( ~n19246 & n19249 ) ;
  assign n19251 = ( ~n19243 & n19249 ) | ( ~n19243 & n19250 ) | ( n19249 & n19250 ) ;
  assign n19252 = n18001 | n19251 ;
  assign n19253 = n19233 & ~n19247 ;
  assign n19254 = n19248 | n19253 ;
  assign n19255 = n19252 & ~n19254 ;
  assign n19256 = n19248 | n19255 ;
  assign n19257 = n18001 & n19251 ;
  assign n19258 = ~n19254 & n19257 ;
  assign n19259 = n19248 | n19258 ;
  assign n19260 = ( n19231 & n19256 ) | ( n19231 & n19259 ) | ( n19256 & n19259 ) ;
  assign n19261 = ~n16854 & n19260 ;
  assign n19262 = n16852 | n19261 ;
  assign n19263 = n14451 & ~n14456 ;
  assign n19264 = ~n14451 & n14455 ;
  assign n19265 = n19263 | n19264 ;
  assign n19266 = n14448 & ~n14449 ;
  assign n19267 = ~n14446 & n19266 ;
  assign n19268 = n14450 | n19267 ;
  assign n19269 = ~n12314 & n12878 ;
  assign n19270 = ( ~n12318 & n12879 ) | ( ~n12318 & n19269 ) | ( n12879 & n19269 ) ;
  assign n19271 = n7308 | n19270 ;
  assign n19272 = n12615 & ~n19270 ;
  assign n19273 = ( n12314 & ~n12604 ) | ( n12314 & n19272 ) | ( ~n12604 & n19272 ) ;
  assign n19274 = n19271 & ~n19273 ;
  assign n19275 = x11 & ~n19274 ;
  assign n19276 = ~x11 & n19274 ;
  assign n19277 = n19275 | n19276 ;
  assign n19278 = ( ~n14441 & n14442 ) | ( ~n14441 & n14443 ) | ( n14442 & n14443 ) ;
  assign n19279 = ~n14427 & n14429 ;
  assign n19280 = n14430 | n19279 ;
  assign n19281 = n5083 & ~n12586 ;
  assign n19282 = n5069 & n12340 ;
  assign n19283 = n5070 & ~n12344 ;
  assign n19284 = n19282 | n19283 ;
  assign n19285 = n19281 | n19284 ;
  assign n19286 = ( n5074 & n13454 ) | ( n5074 & n13455 ) | ( n13454 & n13455 ) ;
  assign n19287 = n19285 | n19286 ;
  assign n19288 = x17 | n19287 ;
  assign n19289 = ~x17 & n19288 ;
  assign n19290 = ( ~n19287 & n19288 ) | ( ~n19287 & n19289 ) | ( n19288 & n19289 ) ;
  assign n19291 = ~n19280 & n19290 ;
  assign n19292 = ( ~n14425 & n14426 ) | ( ~n14425 & n14427 ) | ( n14426 & n14427 ) ;
  assign n19293 = n16292 | n16299 ;
  assign n19294 = n4781 & n12355 ;
  assign n19295 = n4776 & ~n12537 ;
  assign n19296 = n4778 & n12351 ;
  assign n19297 = n19295 | n19296 ;
  assign n19298 = n19294 | n19297 ;
  assign n19299 = n4784 | n19298 ;
  assign n19300 = ( n13409 & n19298 ) | ( n13409 & n19299 ) | ( n19298 & n19299 ) ;
  assign n19301 = x20 & n19300 ;
  assign n19302 = x20 & ~n19301 ;
  assign n19303 = ( n19300 & ~n19301 ) | ( n19300 & n19302 ) | ( ~n19301 & n19302 ) ;
  assign n19304 = ( ~n14402 & n14412 ) | ( ~n14402 & n14414 ) | ( n14412 & n14414 ) ;
  assign n19305 = ( n14402 & ~n14414 ) | ( n14402 & n19304 ) | ( ~n14414 & n19304 ) ;
  assign n19306 = ( ~n14412 & n19304 ) | ( ~n14412 & n19305 ) | ( n19304 & n19305 ) ;
  assign n19307 = ( n19293 & n19303 ) | ( n19293 & n19306 ) | ( n19303 & n19306 ) ;
  assign n19308 = n5083 & ~n12344 ;
  assign n19309 = n5069 & n12553 ;
  assign n19310 = n5070 & n12340 ;
  assign n19311 = n19309 | n19310 ;
  assign n19312 = n19308 | n19311 ;
  assign n19313 = n5074 | n19312 ;
  assign n19314 = ( ~n13523 & n19312 ) | ( ~n13523 & n19313 ) | ( n19312 & n19313 ) ;
  assign n19315 = ~x17 & n19314 ;
  assign n19316 = x17 | n19315 ;
  assign n19317 = ( ~n19314 & n19315 ) | ( ~n19314 & n19316 ) | ( n19315 & n19316 ) ;
  assign n19318 = ( n19292 & ~n19307 ) | ( n19292 & n19317 ) | ( ~n19307 & n19317 ) ;
  assign n19319 = ( ~n19292 & n19307 ) | ( ~n19292 & n19318 ) | ( n19307 & n19318 ) ;
  assign n19320 = n19280 | n19291 ;
  assign n19321 = ( ~n19290 & n19291 ) | ( ~n19290 & n19320 ) | ( n19291 & n19320 ) ;
  assign n19322 = n19319 & ~n19321 ;
  assign n19323 = n19291 | n19322 ;
  assign n19324 = n7280 & ~n12328 ;
  assign n19325 = n5384 & ~n12335 ;
  assign n19326 = n7277 & ~n12325 ;
  assign n19327 = n19325 | n19326 ;
  assign n19328 = n19324 | n19327 ;
  assign n19329 = n39 | n19328 ;
  assign n19330 = ( ~n13544 & n19328 ) | ( ~n13544 & n19329 ) | ( n19328 & n19329 ) ;
  assign n19331 = ~x14 & n19330 ;
  assign n19332 = x14 | n19331 ;
  assign n19333 = ( ~n19330 & n19331 ) | ( ~n19330 & n19332 ) | ( n19331 & n19332 ) ;
  assign n19334 = ( n19278 & ~n19323 ) | ( n19278 & n19333 ) | ( ~n19323 & n19333 ) ;
  assign n19335 = ( ~n19278 & n19323 ) | ( ~n19278 & n19334 ) | ( n19323 & n19334 ) ;
  assign n19336 = n19277 & n19335 ;
  assign n19337 = ( n14331 & ~n14342 ) | ( n14331 & n14444 ) | ( ~n14342 & n14444 ) ;
  assign n19338 = ( ~n14443 & n14444 ) | ( ~n14443 & n19337 ) | ( n14444 & n19337 ) ;
  assign n19339 = n19277 | n19335 ;
  assign n19340 = ~n19336 & n19339 ;
  assign n19341 = ~n19338 & n19340 ;
  assign n19342 = n19336 | n19341 ;
  assign n19343 = ~n19268 & n19342 ;
  assign n19344 = n19268 & ~n19342 ;
  assign n19345 = n19343 | n19344 ;
  assign n19346 = n19338 | n19341 ;
  assign n19347 = ( ~n19340 & n19341 ) | ( ~n19340 & n19346 ) | ( n19341 & n19346 ) ;
  assign n19348 = ( ~n19333 & n19334 ) | ( ~n19333 & n19335 ) | ( n19334 & n19335 ) ;
  assign n19349 = ~n19319 & n19321 ;
  assign n19350 = n19322 | n19349 ;
  assign n19351 = n7280 & ~n12325 ;
  assign n19352 = n5384 & n12580 ;
  assign n19353 = n7277 & ~n12335 ;
  assign n19354 = n19352 | n19353 ;
  assign n19355 = n19351 | n19354 ;
  assign n19356 = n39 | n19355 ;
  assign n19357 = ( ~n13720 & n19355 ) | ( ~n13720 & n19356 ) | ( n19355 & n19356 ) ;
  assign n19358 = ~x14 & n19357 ;
  assign n19359 = x14 | n19358 ;
  assign n19360 = ( ~n19357 & n19358 ) | ( ~n19357 & n19359 ) | ( n19358 & n19359 ) ;
  assign n19361 = ~n19350 & n19360 ;
  assign n19362 = ( ~n19317 & n19318 ) | ( ~n19317 & n19319 ) | ( n19318 & n19319 ) ;
  assign n19363 = n16312 | n16318 ;
  assign n19364 = ( n19293 & n19303 ) | ( n19293 & ~n19306 ) | ( n19303 & ~n19306 ) ;
  assign n19365 = ( ~n19293 & n19306 ) | ( ~n19293 & n19364 ) | ( n19306 & n19364 ) ;
  assign n19366 = ( ~n19303 & n19364 ) | ( ~n19303 & n19365 ) | ( n19364 & n19365 ) ;
  assign n19367 = n19363 & n19366 ;
  assign n19368 = n19363 | n19366 ;
  assign n19369 = ~n19367 & n19368 ;
  assign n19370 = n5083 & n12340 ;
  assign n19371 = n5069 & n12558 ;
  assign n19372 = n5070 & n12553 ;
  assign n19373 = n19371 | n19372 ;
  assign n19374 = n19370 | n19373 ;
  assign n19375 = n5074 & n13347 ;
  assign n19376 = ( n5074 & n13346 ) | ( n5074 & n19375 ) | ( n13346 & n19375 ) ;
  assign n19377 = n19374 | n19376 ;
  assign n19378 = x17 | n19377 ;
  assign n19379 = ~x17 & n19378 ;
  assign n19380 = ( ~n19377 & n19378 ) | ( ~n19377 & n19379 ) | ( n19378 & n19379 ) ;
  assign n19381 = n19369 & n19380 ;
  assign n19382 = n19367 | n19381 ;
  assign n19383 = n7280 & ~n12335 ;
  assign n19384 = n5384 & ~n12586 ;
  assign n19385 = n7277 & n12580 ;
  assign n19386 = n19384 | n19385 ;
  assign n19387 = n19383 | n19386 ;
  assign n19388 = n39 & n13587 ;
  assign n19389 = ( n39 & n13585 ) | ( n39 & n19388 ) | ( n13585 & n19388 ) ;
  assign n19390 = n19387 | n19389 ;
  assign n19391 = x14 | n19390 ;
  assign n19392 = ~x14 & n19391 ;
  assign n19393 = ( ~n19390 & n19391 ) | ( ~n19390 & n19392 ) | ( n19391 & n19392 ) ;
  assign n19394 = ( n19362 & ~n19382 ) | ( n19362 & n19393 ) | ( ~n19382 & n19393 ) ;
  assign n19395 = ( ~n19362 & n19382 ) | ( ~n19362 & n19394 ) | ( n19382 & n19394 ) ;
  assign n19396 = n19350 | n19361 ;
  assign n19397 = ( ~n19360 & n19361 ) | ( ~n19360 & n19396 ) | ( n19361 & n19396 ) ;
  assign n19398 = n19395 & ~n19397 ;
  assign n19399 = n19361 | n19398 ;
  assign n19400 = n7302 & ~n12318 ;
  assign n19401 = n7300 & n12608 ;
  assign n19402 = n19400 | n19401 ;
  assign n19403 = n7305 & ~n12314 ;
  assign n19404 = n19402 | n19403 ;
  assign n19405 = n7308 | n19404 ;
  assign n19406 = ( ~n14302 & n19404 ) | ( ~n14302 & n19405 ) | ( n19404 & n19405 ) ;
  assign n19407 = ~x11 & n19406 ;
  assign n19408 = x11 | n19407 ;
  assign n19409 = ( ~n19406 & n19407 ) | ( ~n19406 & n19408 ) | ( n19407 & n19408 ) ;
  assign n19410 = ( n19348 & ~n19399 ) | ( n19348 & n19409 ) | ( ~n19399 & n19409 ) ;
  assign n19411 = ( ~n19348 & n19399 ) | ( ~n19348 & n19410 ) | ( n19399 & n19410 ) ;
  assign n19412 = ~n19347 & n19411 ;
  assign n19413 = n19347 & ~n19411 ;
  assign n19414 = n19412 | n19413 ;
  assign n19415 = ( ~n19409 & n19410 ) | ( ~n19409 & n19411 ) | ( n19410 & n19411 ) ;
  assign n19416 = n7305 & ~n12318 ;
  assign n19417 = n7300 & ~n12328 ;
  assign n19418 = n7302 & n12608 ;
  assign n19419 = n19417 | n19418 ;
  assign n19420 = n19416 | n19419 ;
  assign n19421 = n7308 | n19420 ;
  assign n19422 = ( n14320 & n19420 ) | ( n14320 & n19421 ) | ( n19420 & n19421 ) ;
  assign n19423 = x11 & n19422 ;
  assign n19424 = x11 & ~n19423 ;
  assign n19425 = ( n19422 & ~n19423 ) | ( n19422 & n19424 ) | ( ~n19423 & n19424 ) ;
  assign n19426 = ( ~n19393 & n19394 ) | ( ~n19393 & n19395 ) | ( n19394 & n19395 ) ;
  assign n19427 = n19369 & ~n19381 ;
  assign n19428 = n16330 | n16335 ;
  assign n19429 = ~n19369 & n19380 ;
  assign n19432 = ( n19427 & n19428 ) | ( n19427 & n19429 ) | ( n19428 & n19429 ) ;
  assign n19430 = n19428 | n19429 ;
  assign n19431 = n19427 | n19430 ;
  assign n19433 = n19431 & ~n19432 ;
  assign n19434 = n7280 & n12580 ;
  assign n19435 = n5384 & ~n12344 ;
  assign n19436 = n7277 & ~n12586 ;
  assign n19437 = n19435 | n19436 ;
  assign n19438 = n19434 | n19437 ;
  assign n19439 = n39 | n19438 ;
  assign n19440 = ( n13432 & n19438 ) | ( n13432 & n19439 ) | ( n19438 & n19439 ) ;
  assign n19441 = x14 & n19440 ;
  assign n19442 = x14 & ~n19441 ;
  assign n19443 = ( n19440 & ~n19441 ) | ( n19440 & n19442 ) | ( ~n19441 & n19442 ) ;
  assign n19444 = n19433 & n19443 ;
  assign n19445 = n19432 | n19444 ;
  assign n19446 = n7300 & ~n12325 ;
  assign n19447 = n7302 & ~n12328 ;
  assign n19448 = n19446 | n19447 ;
  assign n19449 = n7305 & n12608 ;
  assign n19450 = n19448 | n19449 ;
  assign n19451 = n7308 & n13570 ;
  assign n19452 = ( n7308 & n13568 ) | ( n7308 & n19451 ) | ( n13568 & n19451 ) ;
  assign n19453 = n19450 | n19452 ;
  assign n19454 = x11 | n19453 ;
  assign n19455 = ~x11 & n19454 ;
  assign n19456 = ( ~n19453 & n19454 ) | ( ~n19453 & n19455 ) | ( n19454 & n19455 ) ;
  assign n19457 = ( ~n19426 & n19445 ) | ( ~n19426 & n19456 ) | ( n19445 & n19456 ) ;
  assign n19458 = n19425 & n19457 ;
  assign n19459 = n19457 & ~n19458 ;
  assign n19460 = ~n19395 & n19397 ;
  assign n19461 = n19398 | n19460 ;
  assign n19462 = n19425 & ~n19457 ;
  assign n19463 = ( n19459 & ~n19461 ) | ( n19459 & n19462 ) | ( ~n19461 & n19462 ) ;
  assign n19464 = n19458 | n19463 ;
  assign n19465 = ~n19415 & n19464 ;
  assign n19466 = n19464 & ~n19465 ;
  assign n19467 = n19415 | n19464 ;
  assign n19468 = ~n19466 & n19467 ;
  assign n19469 = ~n12314 & n12701 ;
  assign n19470 = ( ~n12318 & n12702 ) | ( ~n12318 & n19469 ) | ( n12702 & n19469 ) ;
  assign n19471 = n5515 | n19470 ;
  assign n19472 = n12615 & ~n19470 ;
  assign n19473 = ( n12314 & ~n12604 ) | ( n12314 & n19472 ) | ( ~n12604 & n19472 ) ;
  assign n19474 = n19471 & ~n19473 ;
  assign n19475 = x8 & ~n19474 ;
  assign n19476 = ~x8 & n19474 ;
  assign n19477 = n19475 | n19476 ;
  assign n19478 = n19433 & ~n19444 ;
  assign n19479 = n16337 | n16340 ;
  assign n19480 = ~n19433 & n19443 ;
  assign n19481 = n19479 | n19480 ;
  assign n19482 = n19478 | n19481 ;
  assign n19483 = n7305 & ~n12328 ;
  assign n19484 = n7300 & ~n12335 ;
  assign n19485 = n7302 & ~n12325 ;
  assign n19486 = n19484 | n19485 ;
  assign n19487 = n19483 | n19486 ;
  assign n19488 = n7308 | n19487 ;
  assign n19489 = ( ~n13544 & n19487 ) | ( ~n13544 & n19488 ) | ( n19487 & n19488 ) ;
  assign n19490 = ~x11 & n19489 ;
  assign n19491 = x11 | n19490 ;
  assign n19492 = ( ~n19489 & n19490 ) | ( ~n19489 & n19491 ) | ( n19490 & n19491 ) ;
  assign n19493 = ( n19478 & n19479 ) | ( n19478 & n19480 ) | ( n19479 & n19480 ) ;
  assign n19494 = ( n19482 & n19492 ) | ( n19482 & n19493 ) | ( n19492 & n19493 ) ;
  assign n19495 = n19477 & n19494 ;
  assign n19496 = ( n19426 & ~n19445 ) | ( n19426 & n19457 ) | ( ~n19445 & n19457 ) ;
  assign n19497 = ( ~n19456 & n19457 ) | ( ~n19456 & n19496 ) | ( n19457 & n19496 ) ;
  assign n19498 = n19477 | n19494 ;
  assign n19499 = ~n19495 & n19498 ;
  assign n19500 = ~n19497 & n19499 ;
  assign n19501 = n19495 | n19500 ;
  assign n19502 = n19461 & ~n19462 ;
  assign n19503 = ~n19459 & n19502 ;
  assign n19504 = n19463 | n19503 ;
  assign n19505 = n19501 & ~n19504 ;
  assign n19506 = ~n19501 & n19504 ;
  assign n19507 = n19505 | n19506 ;
  assign n19508 = n19497 | n19500 ;
  assign n19509 = n19499 & ~n19500 ;
  assign n19510 = n19508 & ~n19509 ;
  assign n19511 = n16343 | n16346 ;
  assign n19512 = n19482 & ~n19493 ;
  assign n19513 = ~n19492 & n19512 ;
  assign n19514 = n19492 | n19513 ;
  assign n19515 = ( ~n19512 & n19513 ) | ( ~n19512 & n19514 ) | ( n19513 & n19514 ) ;
  assign n19516 = n5508 & ~n12318 ;
  assign n19517 = n5512 & n12608 ;
  assign n19518 = n19516 | n19517 ;
  assign n19519 = n5503 & ~n12314 ;
  assign n19520 = n19518 | n19519 ;
  assign n19521 = n5515 | n19520 ;
  assign n19522 = ( ~n14302 & n19520 ) | ( ~n14302 & n19521 ) | ( n19520 & n19521 ) ;
  assign n19523 = ~x8 & n19522 ;
  assign n19524 = x8 | n19523 ;
  assign n19525 = ( ~n19522 & n19523 ) | ( ~n19522 & n19524 ) | ( n19523 & n19524 ) ;
  assign n19526 = ( n19511 & n19515 ) | ( n19511 & n19525 ) | ( n19515 & n19525 ) ;
  assign n19527 = ~n19510 & n19526 ;
  assign n19528 = n19510 & ~n19526 ;
  assign n19529 = n19527 | n19528 ;
  assign n19530 = ( n19511 & ~n19515 ) | ( n19511 & n19525 ) | ( ~n19515 & n19525 ) ;
  assign n19531 = ( ~n19511 & n19515 ) | ( ~n19511 & n19530 ) | ( n19515 & n19530 ) ;
  assign n19532 = ( ~n19525 & n19530 ) | ( ~n19525 & n19531 ) | ( n19530 & n19531 ) ;
  assign n19533 = ( n16258 & n16350 ) | ( n16258 & n19532 ) | ( n16350 & n19532 ) ;
  assign n19534 = ( n16258 & n16350 ) | ( n16258 & ~n19532 ) | ( n16350 & ~n19532 ) ;
  assign n19535 = ( n19532 & ~n19533 ) | ( n19532 & n19534 ) | ( ~n19533 & n19534 ) ;
  assign n19536 = n19533 | n19535 ;
  assign n19537 = ~n19529 & n19536 ;
  assign n19538 = n19527 | n19537 ;
  assign n19539 = ~n19507 & n19538 ;
  assign n19540 = n19505 | n19539 ;
  assign n19541 = ~n19468 & n19540 ;
  assign n19542 = n19465 | n19541 ;
  assign n19543 = ~n19414 & n19542 ;
  assign n19544 = n19412 | n19543 ;
  assign n19545 = ~n19345 & n19544 ;
  assign n19546 = n19343 | n19545 ;
  assign n19547 = n19265 & n19546 ;
  assign n19548 = ~n19529 & n19533 ;
  assign n19549 = n19527 | n19548 ;
  assign n19550 = ~n19507 & n19549 ;
  assign n19551 = n19505 | n19550 ;
  assign n19552 = ~n19468 & n19551 ;
  assign n19553 = n19465 | n19552 ;
  assign n19554 = ~n19414 & n19553 ;
  assign n19555 = n19412 | n19554 ;
  assign n19556 = ~n19345 & n19555 ;
  assign n19557 = n19343 | n19556 ;
  assign n19558 = n19265 & n19557 ;
  assign n19559 = ( n19262 & n19547 ) | ( n19262 & n19558 ) | ( n19547 & n19558 ) ;
  assign n19560 = n14456 | n19559 ;
  assign n19561 = n14317 & n19560 ;
  assign n19562 = n4551 & ~n12318 ;
  assign n19563 = n4546 & ~n12328 ;
  assign n19564 = n4548 & n12608 ;
  assign n19565 = n19563 | n19564 ;
  assign n19566 = n19562 | n19565 ;
  assign n19567 = n4554 | n19566 ;
  assign n19568 = ( n14320 & n19566 ) | ( n14320 & n19567 ) | ( n19566 & n19567 ) ;
  assign n19569 = x23 & n19568 ;
  assign n19570 = x23 & ~n19569 ;
  assign n19571 = ( n19568 & ~n19569 ) | ( n19568 & n19570 ) | ( ~n19569 & n19570 ) ;
  assign n19572 = n4546 & ~n12325 ;
  assign n19573 = n4548 & ~n12328 ;
  assign n19574 = n19572 | n19573 ;
  assign n19575 = n4551 & n12608 ;
  assign n19576 = n19574 | n19575 ;
  assign n19577 = n4554 & n13570 ;
  assign n19578 = ( n4554 & n13568 ) | ( n4554 & n19577 ) | ( n13568 & n19577 ) ;
  assign n19579 = n19576 | n19578 ;
  assign n19580 = x23 | n19579 ;
  assign n19581 = ~x23 & n19580 ;
  assign n19582 = ( ~n19579 & n19580 ) | ( ~n19579 & n19581 ) | ( n19580 & n19581 ) ;
  assign n19583 = n1311 | n2922 ;
  assign n19584 = n213 | n539 ;
  assign n19585 = n458 | n19584 ;
  assign n19586 = n19583 | n19585 ;
  assign n19587 = n646 | n19586 ;
  assign n19588 = n1513 | n12992 ;
  assign n19589 = n3788 | n19588 ;
  assign n19590 = n3264 | n11266 ;
  assign n19591 = n19589 | n19590 ;
  assign n19592 = n19587 | n19591 ;
  assign n19593 = n2850 & ~n19592 ;
  assign n19594 = ~n6007 & n19593 ;
  assign n19595 = n1054 | n2801 ;
  assign n19596 = n618 | n19595 ;
  assign n19597 = n241 | n19596 ;
  assign n19598 = n351 | n19597 ;
  assign n19599 = n19594 & ~n19598 ;
  assign n19600 = n203 | n417 ;
  assign n19601 = ( n2999 & n19599 ) | ( n2999 & ~n19600 ) | ( n19599 & ~n19600 ) ;
  assign n19602 = ~n2999 & n19601 ;
  assign n19603 = n13371 & ~n19602 ;
  assign n19604 = ~n13371 & n19602 ;
  assign n19605 = n19603 | n19604 ;
  assign n19606 = n39 | n12321 ;
  assign n19607 = ~n12314 & n19606 ;
  assign n19608 = ~x14 & n19607 ;
  assign n19609 = x14 | n19608 ;
  assign n19610 = ( ~n19607 & n19608 ) | ( ~n19607 & n19609 ) | ( n19608 & n19609 ) ;
  assign n19611 = n19605 | n19610 ;
  assign n19612 = n2922 | n5170 ;
  assign n19613 = n245 | n19612 ;
  assign n19614 = n618 | n19613 ;
  assign n19615 = n4879 | n13189 ;
  assign n19616 = n472 | n484 ;
  assign n19617 = n244 | n499 ;
  assign n19618 = n19616 | n19617 ;
  assign n19619 = n99 | n596 ;
  assign n19620 = n19618 | n19619 ;
  assign n19621 = ( ~n3765 & n19615 ) | ( ~n3765 & n19620 ) | ( n19615 & n19620 ) ;
  assign n19622 = n3765 | n19621 ;
  assign n19623 = n19614 | n19622 ;
  assign n19624 = n327 | n380 ;
  assign n19625 = n269 | n19624 ;
  assign n19626 = n359 | n19625 ;
  assign n19627 = n77 | n19626 ;
  assign n19628 = n145 | n19627 ;
  assign n19629 = n2642 | n19628 ;
  assign n19630 = n521 | n19629 ;
  assign n19631 = n19623 | n19630 ;
  assign n19632 = n1489 | n1844 ;
  assign n19633 = n4931 | n19632 ;
  assign n19634 = n2718 | n19633 ;
  assign n19635 = n19631 | n19634 ;
  assign n19636 = n281 | n1416 ;
  assign n19637 = n911 | n1329 ;
  assign n19638 = n19636 | n19637 ;
  assign n19639 = n490 | n510 ;
  assign n19640 = n505 | n19639 ;
  assign n19641 = n310 | n19640 ;
  assign n19642 = n19638 | n19641 ;
  assign n19643 = n175 | n306 ;
  assign n19644 = n186 | n19643 ;
  assign n19645 = n19642 | n19644 ;
  assign n19646 = n1613 | n19645 ;
  assign n19647 = n2410 | n19646 ;
  assign n19648 = n568 | n19647 ;
  assign n19649 = n1656 | n19648 ;
  assign n19650 = n19635 | n19649 ;
  assign n19651 = n432 | n628 ;
  assign n19652 = n636 | n19651 ;
  assign n19653 = n420 | n19652 ;
  assign n19654 = n58 | n19653 ;
  assign n19655 = n110 | n19654 ;
  assign n19656 = n114 | n19655 ;
  assign n19657 = n19650 | n19656 ;
  assign n19658 = ( ~n19603 & n19611 ) | ( ~n19603 & n19657 ) | ( n19611 & n19657 ) ;
  assign n19659 = ( ~n19603 & n19604 ) | ( ~n19603 & n19610 ) | ( n19604 & n19610 ) ;
  assign n19660 = n19657 & n19659 ;
  assign n19661 = n19658 & ~n19660 ;
  assign n19662 = n3744 & n12364 ;
  assign n19663 = n3727 & ~n12360 ;
  assign n19664 = n3639 & n12520 ;
  assign n19665 = n19663 | n19664 ;
  assign n19666 = n19662 | n19665 ;
  assign n19667 = n3636 | n19666 ;
  assign n19668 = n19661 & n19667 ;
  assign n19669 = n19658 & ~n19668 ;
  assign n19670 = n19661 & n19666 ;
  assign n19671 = n19658 & ~n19670 ;
  assign n19672 = ( n13113 & n19669 ) | ( n13113 & n19671 ) | ( n19669 & n19671 ) ;
  assign n19673 = n468 | n488 ;
  assign n19674 = n2685 & ~n19673 ;
  assign n19675 = n252 | n653 ;
  assign n19676 = n591 | n19675 ;
  assign n19677 = n19674 & ~n19676 ;
  assign n19678 = ~n197 & n19677 ;
  assign n19679 = n801 | n1950 ;
  assign n19680 = n2416 | n19679 ;
  assign n19681 = ( n2258 & n19678 ) | ( n2258 & ~n19680 ) | ( n19678 & ~n19680 ) ;
  assign n19682 = ~n2258 & n19681 ;
  assign n19683 = ~n158 & n19682 ;
  assign n19684 = ~n11324 & n19683 ;
  assign n19685 = n3873 | n4406 ;
  assign n19686 = n2810 | n19685 ;
  assign n19687 = n430 | n19686 ;
  assign n19688 = n958 | n19687 ;
  assign n19689 = n19684 & ~n19688 ;
  assign n19690 = n504 | n14057 ;
  assign n19691 = n279 | n19690 ;
  assign n19692 = n580 | n19691 ;
  assign n19693 = n92 | n19692 ;
  assign n19694 = n164 | n19693 ;
  assign n19695 = n186 | n19694 ;
  assign n19696 = n19689 & ~n19695 ;
  assign n19697 = n19657 & n19696 ;
  assign n19698 = n19657 | n19696 ;
  assign n19699 = ~n19669 & n19698 ;
  assign n19700 = ~n19697 & n19699 ;
  assign n19701 = ~n19671 & n19698 ;
  assign n19702 = ~n19697 & n19701 ;
  assign n19703 = ( ~n13113 & n19700 ) | ( ~n13113 & n19702 ) | ( n19700 & n19702 ) ;
  assign n19704 = n19672 | n19703 ;
  assign n19705 = n19697 | n19703 ;
  assign n19706 = n19698 & ~n19705 ;
  assign n19707 = n19704 & ~n19706 ;
  assign n19708 = n3744 & ~n12537 ;
  assign n19709 = n3639 & ~n12360 ;
  assign n19710 = n3727 & n12364 ;
  assign n19711 = n19709 | n19710 ;
  assign n19712 = n19708 | n19711 ;
  assign n19713 = ( n3636 & n13081 ) | ( n3636 & ~n13082 ) | ( n13081 & ~n13082 ) ;
  assign n19714 = n19712 | n19713 ;
  assign n19715 = ~n19707 & n19714 ;
  assign n19716 = n19707 | n19715 ;
  assign n19717 = n19714 & ~n19715 ;
  assign n19718 = n19716 & ~n19717 ;
  assign n19719 = n4048 & n12558 ;
  assign n19720 = n4043 & n12351 ;
  assign n19721 = n4045 & n12355 ;
  assign n19722 = n19720 | n19721 ;
  assign n19723 = n19719 | n19722 ;
  assign n19724 = n4051 | n19723 ;
  assign n19725 = ( n13330 & n19723 ) | ( n13330 & n19724 ) | ( n19723 & n19724 ) ;
  assign n19726 = x29 & n19725 ;
  assign n19727 = x29 & ~n19726 ;
  assign n19728 = ( n19725 & ~n19726 ) | ( n19725 & n19727 ) | ( ~n19726 & n19727 ) ;
  assign n19729 = ~n19718 & n19728 ;
  assign n19730 = n19715 | n19729 ;
  assign n19731 = n2733 | n12648 ;
  assign n19732 = n5758 | n19731 ;
  assign n19733 = n3686 | n19732 ;
  assign n19734 = n3682 | n19733 ;
  assign n19735 = n1561 | n3767 ;
  assign n19736 = n3224 | n11150 ;
  assign n19737 = n299 | n19736 ;
  assign n19738 = n19735 | n19737 ;
  assign n19739 = n160 | n321 ;
  assign n19740 = n142 | n19739 ;
  assign n19741 = n217 | n19740 ;
  assign n19742 = n647 | n19741 ;
  assign n19743 = n19738 | n19742 ;
  assign n19744 = n262 | n279 ;
  assign n19745 = n152 | n198 ;
  assign n19746 = n19744 | n19745 ;
  assign n19747 = n19743 | n19746 ;
  assign n19748 = n19734 | n19747 ;
  assign n19749 = n2471 | n19748 ;
  assign n19750 = n3893 | n19749 ;
  assign n19751 = n1613 | n2362 ;
  assign n19752 = n93 | n19751 ;
  assign n19753 = n2341 | n19752 ;
  assign n19754 = n479 | n19753 ;
  assign n19755 = n349 | n19754 ;
  assign n19756 = n445 | n19755 ;
  assign n19757 = n661 | n19756 ;
  assign n19758 = n19750 | n19757 ;
  assign n19759 = ~n19696 & n19758 ;
  assign n19760 = n19696 & ~n19758 ;
  assign n19761 = n19759 | n19760 ;
  assign n19762 = n5070 | n5083 ;
  assign n19763 = n5069 | n19762 ;
  assign n19764 = n5074 | n19763 ;
  assign n19765 = ~n12314 & n19764 ;
  assign n19766 = ~x17 & n19765 ;
  assign n19767 = x17 | n19766 ;
  assign n19768 = ( ~n19765 & n19766 ) | ( ~n19765 & n19767 ) | ( n19766 & n19767 ) ;
  assign n19769 = n19761 | n19768 ;
  assign n19770 = n19761 & n19768 ;
  assign n19771 = n19769 & ~n19770 ;
  assign n19772 = n3636 & ~n12928 ;
  assign n19773 = ( n3636 & n12925 ) | ( n3636 & n19772 ) | ( n12925 & n19772 ) ;
  assign n19774 = n3744 & n12351 ;
  assign n19775 = n3639 & n12364 ;
  assign n19776 = n3727 & ~n12537 ;
  assign n19777 = n19775 | n19776 ;
  assign n19778 = n19774 | n19777 ;
  assign n19779 = n19771 & n19778 ;
  assign n19780 = ( n19771 & n19773 ) | ( n19771 & n19779 ) | ( n19773 & n19779 ) ;
  assign n19781 = n19773 | n19778 ;
  assign n19782 = ~n19771 & n19781 ;
  assign n19783 = ( n19771 & ~n19780 ) | ( n19771 & n19782 ) | ( ~n19780 & n19782 ) ;
  assign n19784 = n19705 & n19783 ;
  assign n19785 = n19705 | n19783 ;
  assign n19786 = ~n19784 & n19785 ;
  assign n19787 = n19730 & n19786 ;
  assign n19788 = n19730 & ~n19787 ;
  assign n19789 = ( n19786 & ~n19787 ) | ( n19786 & n19788 ) | ( ~n19787 & n19788 ) ;
  assign n19790 = n4048 & n12553 ;
  assign n19791 = n4043 & n12355 ;
  assign n19792 = n4045 & n12558 ;
  assign n19793 = n19791 | n19792 ;
  assign n19794 = n19790 | n19793 ;
  assign n19795 = n4051 | n19794 ;
  assign n19796 = ( n13097 & n19794 ) | ( n13097 & n19795 ) | ( n19794 & n19795 ) ;
  assign n19797 = x29 & n19796 ;
  assign n19798 = x29 & ~n19797 ;
  assign n19799 = ( n19796 & ~n19797 ) | ( n19796 & n19798 ) | ( ~n19797 & n19798 ) ;
  assign n19800 = n19789 & ~n19799 ;
  assign n19801 = ( n19787 & n19789 ) | ( n19787 & ~n19800 ) | ( n19789 & ~n19800 ) ;
  assign n19802 = n245 | n509 ;
  assign n19803 = n283 | n540 ;
  assign n19804 = n19802 | n19803 ;
  assign n19805 = n222 | n291 ;
  assign n19806 = n602 | n19805 ;
  assign n19807 = n19804 | n19806 ;
  assign n19808 = n390 | n19807 ;
  assign n19809 = n19743 | n19808 ;
  assign n19810 = n1372 | n19809 ;
  assign n19811 = n3792 | n19810 ;
  assign n19812 = n409 | n19811 ;
  assign n19813 = n373 | n634 ;
  assign n19814 = n470 | n19813 ;
  assign n19815 = ~n1522 & n3233 ;
  assign n19816 = ~n19814 & n19815 ;
  assign n19817 = ~n167 & n19816 ;
  assign n19818 = n947 | n1159 ;
  assign n19819 = n1423 | n2434 ;
  assign n19820 = n19818 | n19819 ;
  assign n19821 = n19817 & ~n19820 ;
  assign n19822 = ~n147 & n19821 ;
  assign n19823 = n1920 | n2623 ;
  assign n19824 = n6010 | n19823 ;
  assign n19825 = n428 | n529 ;
  assign n19826 = n349 | n19825 ;
  assign n19827 = n295 | n19826 ;
  assign n19828 = n19824 | n19827 ;
  assign n19829 = n186 | n345 ;
  assign n19830 = n19828 | n19829 ;
  assign n19831 = n488 | n1161 ;
  assign n19832 = n4064 | n19831 ;
  assign n19833 = n310 | n366 ;
  assign n19834 = n2036 | n19833 ;
  assign n19835 = n55 | n58 ;
  assign n19836 = n129 | n19835 ;
  assign n19837 = n19834 | n19836 ;
  assign n19838 = n2333 | n19837 ;
  assign n19839 = n479 | n19838 ;
  assign n19840 = ( ~n19830 & n19832 ) | ( ~n19830 & n19839 ) | ( n19832 & n19839 ) ;
  assign n19841 = n19830 | n19840 ;
  assign n19842 = ( n2499 & n19822 ) | ( n2499 & ~n19841 ) | ( n19822 & ~n19841 ) ;
  assign n19843 = ~n2499 & n19842 ;
  assign n19844 = ~n19812 & n19843 ;
  assign n19845 = n326 | n511 ;
  assign n19846 = n359 | n19845 ;
  assign n19847 = n19844 & ~n19846 ;
  assign n19848 = ( n19759 & ~n19769 ) | ( n19759 & n19847 ) | ( ~n19769 & n19847 ) ;
  assign n19849 = ( ~n19759 & n19760 ) | ( ~n19759 & n19768 ) | ( n19760 & n19768 ) ;
  assign n19850 = ~n19847 & n19849 ;
  assign n19851 = n19848 | n19850 ;
  assign n19852 = n3744 & n12355 ;
  assign n19853 = n3727 & n12351 ;
  assign n19854 = n3639 & ~n12537 ;
  assign n19855 = n19853 | n19854 ;
  assign n19856 = n19852 | n19855 ;
  assign n19857 = n3636 | n19856 ;
  assign n19858 = ( n13409 & n19856 ) | ( n13409 & n19857 ) | ( n19856 & n19857 ) ;
  assign n19859 = n19851 & ~n19858 ;
  assign n19860 = ~n19851 & n19858 ;
  assign n19861 = n19859 | n19860 ;
  assign n19862 = ~n19780 & n19861 ;
  assign n19863 = ~n19784 & n19862 ;
  assign n19864 = ( n19780 & n19784 ) | ( n19780 & ~n19861 ) | ( n19784 & ~n19861 ) ;
  assign n19865 = n19863 | n19864 ;
  assign n19866 = n4048 & n12340 ;
  assign n19867 = n4043 & n12558 ;
  assign n19868 = n4045 & n12553 ;
  assign n19869 = n19867 | n19868 ;
  assign n19870 = n19866 | n19869 ;
  assign n19871 = n4051 & ~n13346 ;
  assign n19872 = ~n13347 & n19871 ;
  assign n19873 = ( n4051 & n19870 ) | ( n4051 & ~n19872 ) | ( n19870 & ~n19872 ) ;
  assign n19874 = ~x29 & n19873 ;
  assign n19875 = x29 | n19874 ;
  assign n19876 = ( ~n19873 & n19874 ) | ( ~n19873 & n19875 ) | ( n19874 & n19875 ) ;
  assign n19877 = ~n19865 & n19876 ;
  assign n19878 = n19865 & ~n19876 ;
  assign n19879 = n19877 | n19878 ;
  assign n19880 = n4484 & n12580 ;
  assign n19881 = n4479 & ~n12344 ;
  assign n19882 = n4481 & ~n12586 ;
  assign n19883 = n19881 | n19882 ;
  assign n19884 = n19880 | n19883 ;
  assign n19885 = n4487 | n19884 ;
  assign n19886 = ( n13432 & n19884 ) | ( n13432 & n19885 ) | ( n19884 & n19885 ) ;
  assign n19887 = x26 & n19886 ;
  assign n19888 = x26 & ~n19887 ;
  assign n19889 = ( n19886 & ~n19887 ) | ( n19886 & n19888 ) | ( ~n19887 & n19888 ) ;
  assign n19890 = ( ~n19801 & n19879 ) | ( ~n19801 & n19889 ) | ( n19879 & n19889 ) ;
  assign n19891 = ( n19801 & ~n19879 ) | ( n19801 & n19890 ) | ( ~n19879 & n19890 ) ;
  assign n19892 = n4484 & ~n12335 ;
  assign n19893 = n4479 & ~n12586 ;
  assign n19894 = n4481 & n12580 ;
  assign n19895 = n19893 | n19894 ;
  assign n19896 = n19892 | n19895 ;
  assign n19897 = n4487 & n13587 ;
  assign n19898 = ( n4487 & n13585 ) | ( n4487 & n19897 ) | ( n13585 & n19897 ) ;
  assign n19899 = n19896 | n19898 ;
  assign n19900 = x26 | n19899 ;
  assign n19901 = ~x26 & n19900 ;
  assign n19902 = ( ~n19899 & n19900 ) | ( ~n19899 & n19901 ) | ( n19900 & n19901 ) ;
  assign n19903 = n4048 & ~n12344 ;
  assign n19904 = n4043 & n12553 ;
  assign n19905 = n4045 & n12340 ;
  assign n19906 = n19904 | n19905 ;
  assign n19907 = n19903 | n19906 ;
  assign n19908 = n4051 | n19907 ;
  assign n19909 = ( ~n13523 & n19907 ) | ( ~n13523 & n19908 ) | ( n19907 & n19908 ) ;
  assign n19910 = ~x29 & n19909 ;
  assign n19911 = x29 | n19910 ;
  assign n19912 = ( ~n19909 & n19910 ) | ( ~n19909 & n19911 ) | ( n19910 & n19911 ) ;
  assign n19913 = n3744 & n12558 ;
  assign n19914 = n3639 & n12351 ;
  assign n19915 = n3727 & n12355 ;
  assign n19916 = n19914 | n19915 ;
  assign n19917 = n19913 | n19916 ;
  assign n19918 = n3636 | n19917 ;
  assign n19919 = ( n13330 & n19917 ) | ( n13330 & n19918 ) | ( n19917 & n19918 ) ;
  assign n19920 = n522 | n622 ;
  assign n19921 = n276 | n504 ;
  assign n19922 = n19920 | n19921 ;
  assign n19923 = n650 | n19922 ;
  assign n19924 = n294 | n3774 ;
  assign n19925 = n19923 | n19924 ;
  assign n19926 = n1390 | n19925 ;
  assign n19927 = n4290 | n19926 ;
  assign n19928 = n1820 | n19927 ;
  assign n19929 = n4289 & ~n19928 ;
  assign n19930 = n2950 | n13262 ;
  assign n19931 = n19929 & ~n19930 ;
  assign n19932 = n959 | n2527 ;
  assign n19933 = n1417 | n19932 ;
  assign n19934 = n428 | n19933 ;
  assign n19935 = n634 | n19934 ;
  assign n19936 = n380 | n19935 ;
  assign n19937 = n570 | n19936 ;
  assign n19938 = n5702 | n19937 ;
  assign n19939 = n458 | n19938 ;
  assign n19940 = n19931 & ~n19939 ;
  assign n19941 = n76 | n167 ;
  assign n19942 = n19940 & ~n19941 ;
  assign n19943 = ~n19847 & n19942 ;
  assign n19944 = n19847 & ~n19942 ;
  assign n19945 = n19918 & ~n19944 ;
  assign n19946 = ~n19943 & n19945 ;
  assign n19947 = n19917 & ~n19944 ;
  assign n19948 = ~n19943 & n19947 ;
  assign n19949 = ( n13330 & n19946 ) | ( n13330 & n19948 ) | ( n19946 & n19948 ) ;
  assign n19950 = n19919 & ~n19949 ;
  assign n19951 = n19848 | n19860 ;
  assign n19952 = n19944 | n19949 ;
  assign n19953 = n19943 | n19952 ;
  assign n19954 = n19951 & ~n19953 ;
  assign n19955 = ( n19950 & n19951 ) | ( n19950 & n19954 ) | ( n19951 & n19954 ) ;
  assign n19956 = ~n19951 & n19953 ;
  assign n19957 = ~n19950 & n19956 ;
  assign n19958 = n19955 | n19957 ;
  assign n19959 = n19864 | n19877 ;
  assign n19960 = ~n19958 & n19959 ;
  assign n19961 = n19958 & ~n19959 ;
  assign n19962 = n19960 | n19961 ;
  assign n19963 = n19912 & ~n19962 ;
  assign n19964 = n19962 | n19963 ;
  assign n19965 = ( ~n19912 & n19963 ) | ( ~n19912 & n19964 ) | ( n19963 & n19964 ) ;
  assign n19966 = n19902 & ~n19965 ;
  assign n19967 = ~n19902 & n19965 ;
  assign n19968 = n19966 | n19967 ;
  assign n19969 = ( n19582 & n19891 ) | ( n19582 & ~n19968 ) | ( n19891 & ~n19968 ) ;
  assign n19970 = n19571 & n19969 ;
  assign n19971 = n19963 | n19966 ;
  assign n19972 = n4484 & ~n12325 ;
  assign n19973 = n4479 & n12580 ;
  assign n19974 = n4481 & ~n12335 ;
  assign n19975 = n19973 | n19974 ;
  assign n19976 = n19972 | n19975 ;
  assign n19977 = n4487 | n19976 ;
  assign n19978 = ( ~n13720 & n19976 ) | ( ~n13720 & n19977 ) | ( n19976 & n19977 ) ;
  assign n19979 = ~x26 & n19978 ;
  assign n19980 = x26 | n19979 ;
  assign n19981 = ( ~n19978 & n19979 ) | ( ~n19978 & n19980 ) | ( n19979 & n19980 ) ;
  assign n19982 = n4048 & ~n12586 ;
  assign n19983 = n4043 & n12340 ;
  assign n19984 = n4045 & ~n12344 ;
  assign n19985 = n19983 | n19984 ;
  assign n19986 = n19982 | n19985 ;
  assign n19987 = ( n4051 & n13454 ) | ( n4051 & n13455 ) | ( n13454 & n13455 ) ;
  assign n19988 = n19986 | n19987 ;
  assign n19989 = x29 | n19988 ;
  assign n19990 = ~x29 & n19989 ;
  assign n19991 = ( ~n19988 & n19989 ) | ( ~n19988 & n19990 ) | ( n19989 & n19990 ) ;
  assign n19992 = n3744 & n12553 ;
  assign n19993 = n3639 & n12355 ;
  assign n19994 = n3727 & n12558 ;
  assign n19995 = n19993 | n19994 ;
  assign n19996 = n19992 | n19995 ;
  assign n19997 = n3636 | n19996 ;
  assign n19998 = ( n13097 & n19996 ) | ( n13097 & n19997 ) | ( n19996 & n19997 ) ;
  assign n19999 = ~n1655 & n1663 ;
  assign n20000 = n1884 | n4077 ;
  assign n20001 = n2459 | n20000 ;
  assign n20002 = n1737 | n3531 ;
  assign n20003 = n20001 | n20002 ;
  assign n20004 = n1462 | n2221 ;
  assign n20005 = n20003 | n20004 ;
  assign n20006 = n1417 | n1578 ;
  assign n20007 = n432 | n20006 ;
  assign n20008 = n618 | n20007 ;
  assign n20009 = n654 | n20008 ;
  assign n20010 = n110 | n20009 ;
  assign n20011 = n20005 | n20010 ;
  assign n20012 = n1045 | n3060 ;
  assign n20013 = ( n1203 & ~n2682 ) | ( n1203 & n4841 ) | ( ~n2682 & n4841 ) ;
  assign n20014 = n2682 | n20013 ;
  assign n20015 = n20012 | n20014 ;
  assign n20016 = n640 | n20015 ;
  assign n20017 = n20011 | n20016 ;
  assign n20018 = n19999 & ~n20017 ;
  assign n20019 = n1170 | n1194 ;
  assign n20020 = n1310 | n20019 ;
  assign n20021 = n653 | n20020 ;
  assign n20022 = n639 | n20021 ;
  assign n20023 = n174 | n20022 ;
  assign n20024 = n142 | n20023 ;
  assign n20025 = n187 | n20024 ;
  assign n20026 = n157 | n20025 ;
  assign n20027 = n20018 & ~n20026 ;
  assign n20028 = ~n208 & n20027 ;
  assign n20029 = n19847 & n20028 ;
  assign n20030 = n19847 | n20028 ;
  assign n20031 = ~n20029 & n20030 ;
  assign n20032 = n4778 | n4781 ;
  assign n20033 = n4776 | n20032 ;
  assign n20034 = n4784 | n20033 ;
  assign n20035 = ~n12314 & n20034 ;
  assign n20036 = ~x20 & n20035 ;
  assign n20037 = x20 | n20036 ;
  assign n20038 = ( ~n20035 & n20036 ) | ( ~n20035 & n20037 ) | ( n20036 & n20037 ) ;
  assign n20039 = n20031 & ~n20038 ;
  assign n20040 = ~n20031 & n20038 ;
  assign n20041 = n20039 | n20040 ;
  assign n20042 = ( n19952 & n19998 ) | ( n19952 & ~n20041 ) | ( n19998 & ~n20041 ) ;
  assign n20043 = ( ~n19952 & n20041 ) | ( ~n19952 & n20042 ) | ( n20041 & n20042 ) ;
  assign n20044 = ( ~n19998 & n20042 ) | ( ~n19998 & n20043 ) | ( n20042 & n20043 ) ;
  assign n20045 = ( n19955 & n19960 ) | ( n19955 & ~n20044 ) | ( n19960 & ~n20044 ) ;
  assign n20046 = ( n19955 & ~n19957 ) | ( n19955 & n19959 ) | ( ~n19957 & n19959 ) ;
  assign n20047 = n20044 & ~n20046 ;
  assign n20048 = n20045 | n20047 ;
  assign n20049 = n19991 & ~n20048 ;
  assign n20050 = n20048 | n20049 ;
  assign n20051 = ( ~n19991 & n20049 ) | ( ~n19991 & n20050 ) | ( n20049 & n20050 ) ;
  assign n20052 = n19981 & ~n20051 ;
  assign n20053 = ~n19981 & n20051 ;
  assign n20054 = n20052 | n20053 ;
  assign n20055 = n19971 & ~n20054 ;
  assign n20056 = ~n19971 & n20054 ;
  assign n20057 = n20055 | n20056 ;
  assign n20058 = n19969 & ~n19970 ;
  assign n20059 = n19571 & ~n19969 ;
  assign n20060 = ( ~n20057 & n20058 ) | ( ~n20057 & n20059 ) | ( n20058 & n20059 ) ;
  assign n20061 = n19970 | n20060 ;
  assign n20062 = n4548 & ~n12318 ;
  assign n20063 = n4546 & n12608 ;
  assign n20064 = n20062 | n20063 ;
  assign n20065 = n4551 & ~n12314 ;
  assign n20066 = n20064 | n20065 ;
  assign n20067 = n4554 | n20066 ;
  assign n20068 = ( ~n14302 & n20066 ) | ( ~n14302 & n20067 ) | ( n20066 & n20067 ) ;
  assign n20069 = ~x23 & n20068 ;
  assign n20070 = x23 | n20069 ;
  assign n20071 = ( ~n20068 & n20069 ) | ( ~n20068 & n20070 ) | ( n20069 & n20070 ) ;
  assign n20072 = n20052 | n20055 ;
  assign n20073 = n20045 | n20049 ;
  assign n20074 = n12255 | n12258 ;
  assign n20075 = ( n20030 & ~n20039 ) | ( n20030 & n20074 ) | ( ~n20039 & n20074 ) ;
  assign n20076 = ( n20029 & n20030 ) | ( n20029 & n20038 ) | ( n20030 & n20038 ) ;
  assign n20077 = n20074 & n20076 ;
  assign n20078 = n20075 & ~n20077 ;
  assign n20079 = n3636 & n13347 ;
  assign n20080 = ( n3636 & n13346 ) | ( n3636 & n20079 ) | ( n13346 & n20079 ) ;
  assign n20081 = n3744 & n12340 ;
  assign n20082 = n3727 & n12553 ;
  assign n20083 = n3639 & n12558 ;
  assign n20084 = n20082 | n20083 ;
  assign n20085 = n20081 | n20084 ;
  assign n20086 = n20078 & n20085 ;
  assign n20087 = ( n20078 & n20080 ) | ( n20078 & n20086 ) | ( n20080 & n20086 ) ;
  assign n20088 = n20078 | n20085 ;
  assign n20089 = n20080 | n20088 ;
  assign n20090 = ~n20087 & n20089 ;
  assign n20091 = n20042 & n20090 ;
  assign n20092 = n20042 | n20090 ;
  assign n20093 = ~n20091 & n20092 ;
  assign n20094 = n4048 & n12580 ;
  assign n20095 = n4043 & ~n12344 ;
  assign n20096 = n4045 & ~n12586 ;
  assign n20097 = n20095 | n20096 ;
  assign n20098 = n20094 | n20097 ;
  assign n20099 = n4051 | n20098 ;
  assign n20100 = ( n13432 & n20098 ) | ( n13432 & n20099 ) | ( n20098 & n20099 ) ;
  assign n20101 = x29 & n20100 ;
  assign n20102 = x29 & ~n20101 ;
  assign n20103 = ( n20100 & ~n20101 ) | ( n20100 & n20102 ) | ( ~n20101 & n20102 ) ;
  assign n20104 = n20093 & n20103 ;
  assign n20105 = n20093 | n20103 ;
  assign n20106 = ~n20104 & n20105 ;
  assign n20107 = n4484 & ~n12328 ;
  assign n20108 = n4479 & ~n12335 ;
  assign n20109 = n4481 & ~n12325 ;
  assign n20110 = n20108 | n20109 ;
  assign n20111 = n20107 | n20110 ;
  assign n20112 = n4487 | n20111 ;
  assign n20113 = ( ~n13544 & n20111 ) | ( ~n13544 & n20112 ) | ( n20111 & n20112 ) ;
  assign n20114 = ~x26 & n20113 ;
  assign n20115 = x26 | n20114 ;
  assign n20116 = ( ~n20113 & n20114 ) | ( ~n20113 & n20115 ) | ( n20114 & n20115 ) ;
  assign n20117 = ( n20073 & n20106 ) | ( n20073 & n20116 ) | ( n20106 & n20116 ) ;
  assign n20118 = ( n20106 & n20116 ) | ( n20106 & ~n20117 ) | ( n20116 & ~n20117 ) ;
  assign n20119 = ( n20073 & ~n20117 ) | ( n20073 & n20118 ) | ( ~n20117 & n20118 ) ;
  assign n20120 = ( n20071 & ~n20072 ) | ( n20071 & n20119 ) | ( ~n20072 & n20119 ) ;
  assign n20121 = ( n20072 & ~n20119 ) | ( n20072 & n20120 ) | ( ~n20119 & n20120 ) ;
  assign n20122 = ( ~n20071 & n20120 ) | ( ~n20071 & n20121 ) | ( n20120 & n20121 ) ;
  assign n20123 = n20061 & n20122 ;
  assign n20124 = n20061 & ~n20123 ;
  assign n20125 = ~n20061 & n20122 ;
  assign n20126 = n20124 | n20125 ;
  assign n20127 = n20057 & ~n20059 ;
  assign n20128 = ~n20058 & n20127 ;
  assign n20129 = n20060 | n20128 ;
  assign n20130 = ~n12314 & n20032 ;
  assign n20131 = ( ~n12318 & n20033 ) | ( ~n12318 & n20130 ) | ( n20033 & n20130 ) ;
  assign n20132 = n4784 | n20131 ;
  assign n20133 = n12615 & ~n20131 ;
  assign n20134 = ( n12314 & ~n12604 ) | ( n12314 & n20133 ) | ( ~n12604 & n20133 ) ;
  assign n20135 = n20132 & ~n20134 ;
  assign n20136 = x20 & ~n20135 ;
  assign n20137 = ~x20 & n20135 ;
  assign n20138 = n20136 | n20137 ;
  assign n20139 = ( ~n19889 & n19890 ) | ( ~n19889 & n19891 ) | ( n19890 & n19891 ) ;
  assign n20140 = ~n19789 & n19799 ;
  assign n20141 = n19800 | n20140 ;
  assign n20142 = n4484 & ~n12586 ;
  assign n20143 = n4479 & n12340 ;
  assign n20144 = n4481 & ~n12344 ;
  assign n20145 = n20143 | n20144 ;
  assign n20146 = n20142 | n20145 ;
  assign n20147 = ( n4487 & n13454 ) | ( n4487 & n13455 ) | ( n13454 & n13455 ) ;
  assign n20148 = n20146 | n20147 ;
  assign n20149 = x26 | n20148 ;
  assign n20150 = ~x26 & n20149 ;
  assign n20151 = ( ~n20148 & n20149 ) | ( ~n20148 & n20150 ) | ( n20149 & n20150 ) ;
  assign n20152 = n20141 & n20151 ;
  assign n20153 = n20141 | n20151 ;
  assign n20154 = ~n20152 & n20153 ;
  assign n20155 = ( ~n13113 & n19668 ) | ( ~n13113 & n19670 ) | ( n19668 & n19670 ) ;
  assign n20156 = ( ~n13113 & n19666 ) | ( ~n13113 & n19667 ) | ( n19666 & n19667 ) ;
  assign n20157 = n19661 | n20156 ;
  assign n20158 = ~n20155 & n20157 ;
  assign n20159 = n19605 & n19610 ;
  assign n20160 = n19611 & ~n20159 ;
  assign n20161 = ( n13598 & ~n13643 ) | ( n13598 & n13649 ) | ( ~n13643 & n13649 ) ;
  assign n20162 = n3744 & ~n12360 ;
  assign n20163 = n3639 & n12375 ;
  assign n20164 = n3727 & n12520 ;
  assign n20165 = n20163 | n20164 ;
  assign n20166 = n20162 | n20165 ;
  assign n20167 = n3636 | n20166 ;
  assign n20168 = ( ~n12902 & n20166 ) | ( ~n12902 & n20167 ) | ( n20166 & n20167 ) ;
  assign n20169 = ( n20160 & n20161 ) | ( n20160 & n20168 ) | ( n20161 & n20168 ) ;
  assign n20170 = n20158 & n20169 ;
  assign n20171 = n20158 | n20169 ;
  assign n20172 = ~n20170 & n20171 ;
  assign n20173 = n4048 & n12355 ;
  assign n20174 = n4043 & ~n12537 ;
  assign n20175 = n4045 & n12351 ;
  assign n20176 = n20174 | n20175 ;
  assign n20177 = n20173 | n20176 ;
  assign n20178 = n4051 | n20177 ;
  assign n20179 = ( n13409 & n20177 ) | ( n13409 & n20178 ) | ( n20177 & n20178 ) ;
  assign n20180 = x29 & n20179 ;
  assign n20181 = x29 & ~n20180 ;
  assign n20182 = ( n20179 & ~n20180 ) | ( n20179 & n20181 ) | ( ~n20180 & n20181 ) ;
  assign n20183 = n20172 & n20182 ;
  assign n20184 = n20170 | n20183 ;
  assign n20185 = n4484 & ~n12344 ;
  assign n20186 = n4479 & n12553 ;
  assign n20187 = n4481 & n12340 ;
  assign n20188 = n20186 | n20187 ;
  assign n20189 = n20185 | n20188 ;
  assign n20190 = n4487 | n20189 ;
  assign n20191 = ( ~n13523 & n20189 ) | ( ~n13523 & n20190 ) | ( n20189 & n20190 ) ;
  assign n20192 = ~x26 & n20191 ;
  assign n20193 = x26 | n20192 ;
  assign n20194 = ( ~n20191 & n20192 ) | ( ~n20191 & n20193 ) | ( n20192 & n20193 ) ;
  assign n20195 = n19718 & ~n19728 ;
  assign n20196 = n19729 | n20195 ;
  assign n20197 = ( n20184 & ~n20194 ) | ( n20184 & n20196 ) | ( ~n20194 & n20196 ) ;
  assign n20198 = ( ~n20184 & n20194 ) | ( ~n20184 & n20197 ) | ( n20194 & n20197 ) ;
  assign n20199 = ( ~n20196 & n20197 ) | ( ~n20196 & n20198 ) | ( n20197 & n20198 ) ;
  assign n20200 = ( n20184 & n20194 ) | ( n20184 & n20199 ) | ( n20194 & n20199 ) ;
  assign n20201 = n20154 & n20200 ;
  assign n20202 = n20152 | n20201 ;
  assign n20203 = n4551 & ~n12328 ;
  assign n20204 = n4546 & ~n12335 ;
  assign n20205 = n4548 & ~n12325 ;
  assign n20206 = n20204 | n20205 ;
  assign n20207 = n20203 | n20206 ;
  assign n20208 = n4554 | n20207 ;
  assign n20209 = ( ~n13544 & n20207 ) | ( ~n13544 & n20208 ) | ( n20207 & n20208 ) ;
  assign n20210 = ~x23 & n20209 ;
  assign n20211 = x23 | n20210 ;
  assign n20212 = ( ~n20209 & n20210 ) | ( ~n20209 & n20211 ) | ( n20210 & n20211 ) ;
  assign n20213 = ( n20139 & ~n20202 ) | ( n20139 & n20212 ) | ( ~n20202 & n20212 ) ;
  assign n20214 = ( ~n20139 & n20202 ) | ( ~n20139 & n20213 ) | ( n20202 & n20213 ) ;
  assign n20215 = n20138 & n20214 ;
  assign n20216 = ( ~n19582 & n19968 ) | ( ~n19582 & n19969 ) | ( n19968 & n19969 ) ;
  assign n20217 = ( ~n19891 & n19969 ) | ( ~n19891 & n20216 ) | ( n19969 & n20216 ) ;
  assign n20218 = n20138 | n20214 ;
  assign n20219 = ~n20215 & n20218 ;
  assign n20220 = ~n20217 & n20219 ;
  assign n20221 = n20215 | n20220 ;
  assign n20222 = ~n20129 & n20221 ;
  assign n20223 = n20129 & ~n20221 ;
  assign n20224 = n20222 | n20223 ;
  assign n20225 = n20217 | n20220 ;
  assign n20226 = ( ~n20219 & n20220 ) | ( ~n20219 & n20225 ) | ( n20220 & n20225 ) ;
  assign n20227 = ( ~n20212 & n20213 ) | ( ~n20212 & n20214 ) | ( n20213 & n20214 ) ;
  assign n20228 = n20154 | n20200 ;
  assign n20229 = ~n20201 & n20228 ;
  assign n20230 = n4551 & ~n12325 ;
  assign n20231 = n4546 & n12580 ;
  assign n20232 = n4548 & ~n12335 ;
  assign n20233 = n20231 | n20232 ;
  assign n20234 = n20230 | n20233 ;
  assign n20235 = n4554 | n20234 ;
  assign n20236 = ( ~n13720 & n20234 ) | ( ~n13720 & n20235 ) | ( n20234 & n20235 ) ;
  assign n20237 = ~x23 & n20236 ;
  assign n20238 = x23 | n20237 ;
  assign n20239 = ( ~n20236 & n20237 ) | ( ~n20236 & n20238 ) | ( n20237 & n20238 ) ;
  assign n20240 = n20229 & n20239 ;
  assign n20241 = n20229 & ~n20240 ;
  assign n20242 = ~n20229 & n20239 ;
  assign n20243 = n4551 & ~n12335 ;
  assign n20244 = n4546 & ~n12586 ;
  assign n20245 = n4548 & n12580 ;
  assign n20246 = n20244 | n20245 ;
  assign n20247 = n20243 | n20246 ;
  assign n20248 = n4554 & n13587 ;
  assign n20249 = ( n4554 & n13585 ) | ( n4554 & n20248 ) | ( n13585 & n20248 ) ;
  assign n20250 = n20247 | n20249 ;
  assign n20251 = x23 | n20250 ;
  assign n20252 = ~x23 & n20251 ;
  assign n20253 = ( ~n20250 & n20251 ) | ( ~n20250 & n20252 ) | ( n20251 & n20252 ) ;
  assign n20254 = ( n20160 & n20168 ) | ( n20160 & ~n20169 ) | ( n20168 & ~n20169 ) ;
  assign n20255 = ( n20161 & ~n20169 ) | ( n20161 & n20254 ) | ( ~n20169 & n20254 ) ;
  assign n20256 = n4048 & n12351 ;
  assign n20257 = n4043 & n12364 ;
  assign n20258 = n4045 & ~n12537 ;
  assign n20259 = n20257 | n20258 ;
  assign n20260 = n20256 | n20259 ;
  assign n20261 = n4051 & ~n12928 ;
  assign n20262 = ( n4051 & n12925 ) | ( n4051 & n20261 ) | ( n12925 & n20261 ) ;
  assign n20263 = n20260 | n20262 ;
  assign n20264 = x29 | n20263 ;
  assign n20265 = ~x29 & n20264 ;
  assign n20266 = ( ~n20263 & n20264 ) | ( ~n20263 & n20265 ) | ( n20264 & n20265 ) ;
  assign n20267 = n20255 & n20266 ;
  assign n20268 = n20255 & ~n20267 ;
  assign n20269 = ~n20255 & n20266 ;
  assign n20270 = n13657 & ~n13662 ;
  assign n20271 = ( n20268 & n20269 ) | ( n20268 & ~n20270 ) | ( n20269 & ~n20270 ) ;
  assign n20272 = n20172 | n20182 ;
  assign n20273 = ~n20183 & n20272 ;
  assign n20274 = n20267 | n20273 ;
  assign n20275 = n20271 | n20274 ;
  assign n20276 = ( n20267 & n20271 ) | ( n20267 & n20273 ) | ( n20271 & n20273 ) ;
  assign n20277 = n4484 & n12340 ;
  assign n20278 = n4479 & n12558 ;
  assign n20279 = n4481 & n12553 ;
  assign n20280 = n20278 | n20279 ;
  assign n20281 = n20277 | n20280 ;
  assign n20282 = n4487 & n13347 ;
  assign n20283 = ( n4487 & n13346 ) | ( n4487 & n20282 ) | ( n13346 & n20282 ) ;
  assign n20284 = n20281 | n20283 ;
  assign n20285 = x26 | n20284 ;
  assign n20286 = ~x26 & n20285 ;
  assign n20287 = ( ~n20284 & n20285 ) | ( ~n20284 & n20286 ) | ( n20285 & n20286 ) ;
  assign n20288 = ( n20275 & n20276 ) | ( n20275 & n20287 ) | ( n20276 & n20287 ) ;
  assign n20289 = ( n20199 & ~n20253 ) | ( n20199 & n20288 ) | ( ~n20253 & n20288 ) ;
  assign n20290 = ( ~n20199 & n20253 ) | ( ~n20199 & n20289 ) | ( n20253 & n20289 ) ;
  assign n20291 = ( n20241 & n20242 ) | ( n20241 & n20290 ) | ( n20242 & n20290 ) ;
  assign n20292 = n20240 | n20291 ;
  assign n20293 = n4778 & ~n12318 ;
  assign n20294 = n4776 & n12608 ;
  assign n20295 = n20293 | n20294 ;
  assign n20296 = n4781 & ~n12314 ;
  assign n20297 = n20295 | n20296 ;
  assign n20298 = n4784 | n20297 ;
  assign n20299 = ( ~n14302 & n20297 ) | ( ~n14302 & n20298 ) | ( n20297 & n20298 ) ;
  assign n20300 = ~x20 & n20299 ;
  assign n20301 = x20 | n20300 ;
  assign n20302 = ( ~n20299 & n20300 ) | ( ~n20299 & n20301 ) | ( n20300 & n20301 ) ;
  assign n20303 = ( ~n20227 & n20292 ) | ( ~n20227 & n20302 ) | ( n20292 & n20302 ) ;
  assign n20304 = ~n20226 & n20303 ;
  assign n20305 = n20226 & ~n20303 ;
  assign n20306 = n20304 | n20305 ;
  assign n20307 = ( n20227 & ~n20292 ) | ( n20227 & n20303 ) | ( ~n20292 & n20303 ) ;
  assign n20308 = ( ~n20302 & n20303 ) | ( ~n20302 & n20307 ) | ( n20303 & n20307 ) ;
  assign n20309 = n4781 & ~n12318 ;
  assign n20310 = n4776 & ~n12328 ;
  assign n20311 = n4778 & n12608 ;
  assign n20312 = n20310 | n20311 ;
  assign n20313 = n20309 | n20312 ;
  assign n20314 = n4784 | n20313 ;
  assign n20315 = ( n14320 & n20313 ) | ( n14320 & n20314 ) | ( n20313 & n20314 ) ;
  assign n20316 = x20 & n20315 ;
  assign n20317 = x20 & ~n20316 ;
  assign n20318 = ( n20315 & ~n20316 ) | ( n20315 & n20317 ) | ( ~n20316 & n20317 ) ;
  assign n20319 = ( ~n20288 & n20289 ) | ( ~n20288 & n20290 ) | ( n20289 & n20290 ) ;
  assign n20320 = n4776 & ~n12325 ;
  assign n20321 = n4778 & ~n12328 ;
  assign n20322 = n20320 | n20321 ;
  assign n20323 = n4781 & n12608 ;
  assign n20324 = n20322 | n20323 ;
  assign n20325 = n4784 & n13570 ;
  assign n20326 = ( n4784 & n13568 ) | ( n4784 & n20325 ) | ( n13568 & n20325 ) ;
  assign n20327 = n20324 | n20326 ;
  assign n20328 = x20 | n20327 ;
  assign n20329 = ~x20 & n20328 ;
  assign n20330 = ( ~n20327 & n20328 ) | ( ~n20327 & n20329 ) | ( n20328 & n20329 ) ;
  assign n20331 = n20275 & ~n20276 ;
  assign n20332 = ~n20287 & n20331 ;
  assign n20333 = n20287 | n20332 ;
  assign n20334 = ( ~n20331 & n20332 ) | ( ~n20331 & n20333 ) | ( n20332 & n20333 ) ;
  assign n20335 = ~n20269 & n20270 ;
  assign n20336 = ~n20268 & n20335 ;
  assign n20337 = n20271 | n20336 ;
  assign n20338 = n4484 & n12553 ;
  assign n20339 = n4479 & n12355 ;
  assign n20340 = n4481 & n12558 ;
  assign n20341 = n20339 | n20340 ;
  assign n20342 = n20338 | n20341 ;
  assign n20343 = n4487 | n20342 ;
  assign n20344 = ( n13097 & n20342 ) | ( n13097 & n20343 ) | ( n20342 & n20343 ) ;
  assign n20345 = x26 & n20344 ;
  assign n20346 = x26 & ~n20345 ;
  assign n20347 = ( n20344 & ~n20345 ) | ( n20344 & n20346 ) | ( ~n20345 & n20346 ) ;
  assign n20348 = ~n20337 & n20347 ;
  assign n20349 = n13675 | n13689 ;
  assign n20350 = n20337 | n20348 ;
  assign n20351 = ( ~n20347 & n20348 ) | ( ~n20347 & n20350 ) | ( n20348 & n20350 ) ;
  assign n20352 = n20349 & ~n20351 ;
  assign n20353 = n20348 | n20352 ;
  assign n20354 = n4551 & n12580 ;
  assign n20355 = n4546 & ~n12344 ;
  assign n20356 = n4548 & ~n12586 ;
  assign n20357 = n20355 | n20356 ;
  assign n20358 = n20354 | n20357 ;
  assign n20359 = n4554 | n20358 ;
  assign n20360 = ( n13432 & n20358 ) | ( n13432 & n20359 ) | ( n20358 & n20359 ) ;
  assign n20361 = x23 & n20360 ;
  assign n20362 = x23 & ~n20361 ;
  assign n20363 = ( n20360 & ~n20361 ) | ( n20360 & n20362 ) | ( ~n20361 & n20362 ) ;
  assign n20364 = ( n20334 & n20353 ) | ( n20334 & n20363 ) | ( n20353 & n20363 ) ;
  assign n20365 = ( n20319 & ~n20330 ) | ( n20319 & n20364 ) | ( ~n20330 & n20364 ) ;
  assign n20366 = ( ~n20319 & n20330 ) | ( ~n20319 & n20365 ) | ( n20330 & n20365 ) ;
  assign n20367 = n20318 & n20366 ;
  assign n20368 = n20242 | n20290 ;
  assign n20369 = n20241 | n20368 ;
  assign n20370 = ~n20291 & n20369 ;
  assign n20371 = n20366 & ~n20367 ;
  assign n20372 = n20318 & ~n20366 ;
  assign n20373 = ( n20370 & n20371 ) | ( n20370 & n20372 ) | ( n20371 & n20372 ) ;
  assign n20374 = n20367 | n20373 ;
  assign n20375 = ~n20308 & n20374 ;
  assign n20376 = n20308 | n20375 ;
  assign n20377 = n20308 & n20374 ;
  assign n20378 = n20376 & ~n20377 ;
  assign n20379 = n20370 | n20372 ;
  assign n20380 = n20371 | n20379 ;
  assign n20381 = ~n20373 & n20380 ;
  assign n20382 = ~n12314 & n19762 ;
  assign n20383 = ( ~n12318 & n19763 ) | ( ~n12318 & n20382 ) | ( n19763 & n20382 ) ;
  assign n20384 = n5074 | n20383 ;
  assign n20385 = n12615 & ~n20383 ;
  assign n20386 = ( n12314 & ~n12604 ) | ( n12314 & n20385 ) | ( ~n12604 & n20385 ) ;
  assign n20387 = n20384 & ~n20386 ;
  assign n20388 = x17 & ~n20387 ;
  assign n20389 = ~x17 & n20387 ;
  assign n20390 = n20388 | n20389 ;
  assign n20391 = ~n20349 & n20351 ;
  assign n20392 = n20352 | n20391 ;
  assign n20393 = n4551 & ~n12586 ;
  assign n20394 = n4546 & n12340 ;
  assign n20395 = n4548 & ~n12344 ;
  assign n20396 = n20394 | n20395 ;
  assign n20397 = n20393 | n20396 ;
  assign n20398 = ( n4554 & n13454 ) | ( n4554 & n13455 ) | ( n13454 & n13455 ) ;
  assign n20399 = n20397 | n20398 ;
  assign n20400 = x23 | n20399 ;
  assign n20401 = ~x23 & n20400 ;
  assign n20402 = ( ~n20399 & n20400 ) | ( ~n20399 & n20401 ) | ( n20400 & n20401 ) ;
  assign n20403 = ~n20392 & n20402 ;
  assign n20404 = n20392 | n20403 ;
  assign n20405 = n20392 & n20402 ;
  assign n20406 = ( n13702 & ~n20404 ) | ( n13702 & n20405 ) | ( ~n20404 & n20405 ) ;
  assign n20407 = n20403 | n20406 ;
  assign n20408 = n4781 & ~n12328 ;
  assign n20409 = n4776 & ~n12335 ;
  assign n20410 = n4778 & ~n12325 ;
  assign n20411 = n20409 | n20410 ;
  assign n20412 = n20408 | n20411 ;
  assign n20413 = n4784 | n20412 ;
  assign n20414 = ( ~n13544 & n20412 ) | ( ~n13544 & n20413 ) | ( n20412 & n20413 ) ;
  assign n20415 = ~x20 & n20414 ;
  assign n20416 = x20 | n20415 ;
  assign n20417 = ( ~n20414 & n20415 ) | ( ~n20414 & n20416 ) | ( n20415 & n20416 ) ;
  assign n20418 = ( n20334 & ~n20353 ) | ( n20334 & n20363 ) | ( ~n20353 & n20363 ) ;
  assign n20419 = ( ~n20334 & n20353 ) | ( ~n20334 & n20418 ) | ( n20353 & n20418 ) ;
  assign n20420 = ( ~n20363 & n20418 ) | ( ~n20363 & n20419 ) | ( n20418 & n20419 ) ;
  assign n20421 = ( n20407 & n20417 ) | ( n20407 & n20420 ) | ( n20417 & n20420 ) ;
  assign n20422 = n20390 & n20421 ;
  assign n20423 = ( ~n20364 & n20365 ) | ( ~n20364 & n20366 ) | ( n20365 & n20366 ) ;
  assign n20424 = n20390 | n20421 ;
  assign n20425 = ~n20422 & n20424 ;
  assign n20426 = ~n20423 & n20425 ;
  assign n20427 = n20422 | n20426 ;
  assign n20428 = n20381 & n20427 ;
  assign n20429 = n20381 | n20427 ;
  assign n20430 = ~n20428 & n20429 ;
  assign n20431 = n20423 | n20426 ;
  assign n20432 = ( ~n20425 & n20426 ) | ( ~n20425 & n20431 ) | ( n20426 & n20431 ) ;
  assign n20433 = n13702 | n20405 ;
  assign n20434 = n20404 & ~n20433 ;
  assign n20435 = n20406 | n20434 ;
  assign n20436 = n4781 & ~n12325 ;
  assign n20437 = n4776 & n12580 ;
  assign n20438 = n4778 & ~n12335 ;
  assign n20439 = n20437 | n20438 ;
  assign n20440 = n20436 | n20439 ;
  assign n20441 = n4784 | n20440 ;
  assign n20442 = ( ~n13720 & n20440 ) | ( ~n13720 & n20441 ) | ( n20440 & n20441 ) ;
  assign n20443 = ~x20 & n20442 ;
  assign n20444 = x20 | n20443 ;
  assign n20445 = ( ~n20442 & n20443 ) | ( ~n20442 & n20444 ) | ( n20443 & n20444 ) ;
  assign n20446 = ~n20435 & n20445 ;
  assign n20447 = ( n13593 & n13594 ) | ( n13593 & n13704 ) | ( n13594 & n13704 ) ;
  assign n20448 = n20435 | n20446 ;
  assign n20449 = ( ~n20445 & n20446 ) | ( ~n20445 & n20448 ) | ( n20446 & n20448 ) ;
  assign n20450 = n20447 & ~n20449 ;
  assign n20451 = n20446 | n20450 ;
  assign n20452 = n5070 & ~n12318 ;
  assign n20453 = n5069 & n12608 ;
  assign n20454 = n20452 | n20453 ;
  assign n20455 = n5083 & ~n12314 ;
  assign n20456 = n20454 | n20455 ;
  assign n20457 = n5074 | n20456 ;
  assign n20458 = ( ~n14302 & n20456 ) | ( ~n14302 & n20457 ) | ( n20456 & n20457 ) ;
  assign n20459 = ~x17 & n20458 ;
  assign n20460 = x17 | n20459 ;
  assign n20461 = ( ~n20458 & n20459 ) | ( ~n20458 & n20460 ) | ( n20459 & n20460 ) ;
  assign n20462 = ( n20407 & n20417 ) | ( n20407 & ~n20420 ) | ( n20417 & ~n20420 ) ;
  assign n20463 = ( ~n20407 & n20420 ) | ( ~n20407 & n20462 ) | ( n20420 & n20462 ) ;
  assign n20464 = ( ~n20417 & n20462 ) | ( ~n20417 & n20463 ) | ( n20462 & n20463 ) ;
  assign n20465 = ( n20451 & n20461 ) | ( n20451 & n20464 ) | ( n20461 & n20464 ) ;
  assign n20466 = ~n20432 & n20465 ;
  assign n20467 = n20432 & ~n20465 ;
  assign n20468 = n20466 | n20467 ;
  assign n20469 = n5083 & ~n12318 ;
  assign n20470 = n5069 & ~n12328 ;
  assign n20471 = n5070 & n12608 ;
  assign n20472 = n20470 | n20471 ;
  assign n20473 = n20469 | n20472 ;
  assign n20474 = n5074 | n20473 ;
  assign n20475 = ( n14320 & n20473 ) | ( n14320 & n20474 ) | ( n20473 & n20474 ) ;
  assign n20476 = x17 & n20475 ;
  assign n20477 = x17 & ~n20476 ;
  assign n20478 = ( n20475 & ~n20476 ) | ( n20475 & n20477 ) | ( ~n20476 & n20477 ) ;
  assign n20479 = ( n13576 & n13577 ) | ( n13576 & n13707 ) | ( n13577 & n13707 ) ;
  assign n20480 = n20478 & n20479 ;
  assign n20481 = n20479 & ~n20480 ;
  assign n20482 = ~n20447 & n20449 ;
  assign n20483 = n20450 | n20482 ;
  assign n20484 = n20478 & ~n20479 ;
  assign n20485 = ( n20481 & ~n20483 ) | ( n20481 & n20484 ) | ( ~n20483 & n20484 ) ;
  assign n20486 = n20480 | n20485 ;
  assign n20487 = ( ~n20451 & n20461 ) | ( ~n20451 & n20464 ) | ( n20461 & n20464 ) ;
  assign n20488 = ( n20451 & ~n20464 ) | ( n20451 & n20487 ) | ( ~n20464 & n20487 ) ;
  assign n20489 = ( ~n20461 & n20487 ) | ( ~n20461 & n20488 ) | ( n20487 & n20488 ) ;
  assign n20490 = n20486 & n20489 ;
  assign n20491 = n20486 & ~n20490 ;
  assign n20492 = ~n20486 & n20489 ;
  assign n20493 = n20491 | n20492 ;
  assign n20494 = n13557 | n13711 ;
  assign n20495 = n20483 & ~n20484 ;
  assign n20496 = ~n20481 & n20495 ;
  assign n20497 = n20485 | n20496 ;
  assign n20498 = n20494 & ~n20497 ;
  assign n20499 = ~n20494 & n20497 ;
  assign n20500 = n20498 | n20499 ;
  assign n20501 = n14315 & ~n20500 ;
  assign n20502 = n20498 | n20501 ;
  assign n20503 = n20493 & n20502 ;
  assign n20504 = n20490 | n20503 ;
  assign n20505 = ~n20468 & n20504 ;
  assign n20506 = n20466 | n20505 ;
  assign n20507 = n20430 & n20506 ;
  assign n20508 = n20428 | n20507 ;
  assign n20509 = ~n20378 & n20508 ;
  assign n20510 = n20375 | n20509 ;
  assign n20511 = ~n20306 & n20510 ;
  assign n20512 = n20304 | n20511 ;
  assign n20513 = ~n20224 & n20512 ;
  assign n20514 = n20222 | n20513 ;
  assign n20515 = n20126 & n20514 ;
  assign n20516 = n20493 & ~n20499 ;
  assign n20517 = n20490 | n20516 ;
  assign n20518 = ~n20468 & n20517 ;
  assign n20519 = n20466 | n20518 ;
  assign n20520 = n20430 & n20519 ;
  assign n20521 = n20428 | n20520 ;
  assign n20522 = ~n20378 & n20521 ;
  assign n20523 = n20375 | n20522 ;
  assign n20524 = ~n20306 & n20523 ;
  assign n20525 = n20304 | n20524 ;
  assign n20526 = ~n20224 & n20525 ;
  assign n20527 = n20222 | n20526 ;
  assign n20528 = n20126 & n20527 ;
  assign n20529 = ( n19561 & n20515 ) | ( n19561 & n20528 ) | ( n20515 & n20528 ) ;
  assign n20530 = ( n19561 & n20514 ) | ( n19561 & n20527 ) | ( n20514 & n20527 ) ;
  assign n20531 = n20126 | n20530 ;
  assign n20532 = ~n20529 & n20531 ;
  assign n20533 = ( n19561 & n20513 ) | ( n19561 & n20526 ) | ( n20513 & n20526 ) ;
  assign n20534 = ( n19561 & n20512 ) | ( n19561 & n20525 ) | ( n20512 & n20525 ) ;
  assign n20535 = n20224 & ~n20534 ;
  assign n20536 = n20533 | n20535 ;
  assign n20537 = n20532 & ~n20536 ;
  assign n20538 = ~n20532 & n20536 ;
  assign n20539 = ( n19561 & n20509 ) | ( n19561 & n20522 ) | ( n20509 & n20522 ) ;
  assign n20540 = ( n19561 & n20508 ) | ( n19561 & n20521 ) | ( n20508 & n20521 ) ;
  assign n20541 = n20378 & ~n20540 ;
  assign n20542 = n20539 | n20541 ;
  assign n20543 = ( n19561 & n20507 ) | ( n19561 & n20520 ) | ( n20507 & n20520 ) ;
  assign n20544 = ( n19561 & n20506 ) | ( n19561 & n20519 ) | ( n20506 & n20519 ) ;
  assign n20545 = n20430 | n20544 ;
  assign n20546 = ~n20543 & n20545 ;
  assign n20547 = ~n20542 & n20546 ;
  assign n20548 = n20542 & ~n20546 ;
  assign n20549 = ( n19561 & ~n20500 ) | ( n19561 & n20501 ) | ( ~n20500 & n20501 ) ;
  assign n20550 = ~n14315 & n20500 ;
  assign n20551 = ~n19561 & n20550 ;
  assign n20552 = n20549 | n20551 ;
  assign n20553 = ( n19561 & n20503 ) | ( n19561 & n20516 ) | ( n20503 & n20516 ) ;
  assign n20554 = ( n19561 & ~n20499 ) | ( n19561 & n20502 ) | ( ~n20499 & n20502 ) ;
  assign n20555 = n20493 | n20554 ;
  assign n20556 = ~n20553 & n20555 ;
  assign n20557 = ~n20552 & n20556 ;
  assign n20558 = ( n19262 & n19546 ) | ( n19262 & n19557 ) | ( n19546 & n19557 ) ;
  assign n20559 = n19265 | n20558 ;
  assign n20560 = ~n19559 & n20559 ;
  assign n20561 = n14317 | n19560 ;
  assign n20562 = ~n19561 & n20561 ;
  assign n20563 = n20560 & n20562 ;
  assign n20564 = n20560 | n20562 ;
  assign n20565 = ~n20563 & n20564 ;
  assign n20566 = ( n19262 & n19541 ) | ( n19262 & n19552 ) | ( n19541 & n19552 ) ;
  assign n20567 = ( n19262 & n19540 ) | ( n19262 & n19551 ) | ( n19540 & n19551 ) ;
  assign n20568 = n19468 & ~n20567 ;
  assign n20569 = n20566 | n20568 ;
  assign n20570 = ( n19262 & n19543 ) | ( n19262 & n19554 ) | ( n19543 & n19554 ) ;
  assign n20571 = ( n19262 & n19542 ) | ( n19262 & n19553 ) | ( n19542 & n19553 ) ;
  assign n20572 = n19414 & ~n20571 ;
  assign n20573 = n20570 | n20572 ;
  assign n20574 = n20569 | n20573 ;
  assign n20575 = n20569 & n20573 ;
  assign n20576 = n20574 & ~n20575 ;
  assign n20577 = ( n19262 & n19537 ) | ( n19262 & n19548 ) | ( n19537 & n19548 ) ;
  assign n20578 = ( n19262 & n19533 ) | ( n19262 & n19536 ) | ( n19533 & n19536 ) ;
  assign n20579 = n19529 & ~n20578 ;
  assign n20580 = n20577 | n20579 ;
  assign n20581 = ( n19262 & n19539 ) | ( n19262 & n19550 ) | ( n19539 & n19550 ) ;
  assign n20582 = ( n19262 & n19538 ) | ( n19262 & n19549 ) | ( n19538 & n19549 ) ;
  assign n20583 = n19507 & ~n20582 ;
  assign n20584 = n20581 | n20583 ;
  assign n20585 = n20580 | n20584 ;
  assign n20586 = n19262 & n19535 ;
  assign n20587 = n19262 | n19535 ;
  assign n20588 = ~n20586 & n20587 ;
  assign n20589 = ~n20580 & n20588 ;
  assign n20590 = n16854 & ~n19260 ;
  assign n20591 = n19261 | n20590 ;
  assign n20592 = ( n19231 & n19255 ) | ( n19231 & n19258 ) | ( n19255 & n19258 ) ;
  assign n20593 = ( n19231 & n19252 ) | ( n19231 & n19257 ) | ( n19252 & n19257 ) ;
  assign n20594 = n19254 & ~n20593 ;
  assign n20595 = n20592 | n20594 ;
  assign n20596 = n20591 | n20595 ;
  assign n20597 = n20591 & n20595 ;
  assign n20598 = ( ~n18001 & n19231 ) | ( ~n18001 & n19251 ) | ( n19231 & n19251 ) ;
  assign n20599 = ( n18001 & ~n19251 ) | ( n18001 & n20598 ) | ( ~n19251 & n20598 ) ;
  assign n20600 = ( ~n19231 & n20598 ) | ( ~n19231 & n20599 ) | ( n20598 & n20599 ) ;
  assign n20601 = ~n20595 & n20600 ;
  assign n20602 = n20595 & ~n20600 ;
  assign n20603 = ~n18574 & n19229 ;
  assign n20604 = ~n19227 & n20603 ;
  assign n20605 = n19230 | n20604 ;
  assign n20606 = n20600 & ~n20605 ;
  assign n20607 = ~n20600 & n20605 ;
  assign n20608 = n20606 | n20607 ;
  assign n20609 = n18587 | n19226 ;
  assign n20610 = n19224 | n20609 ;
  assign n20611 = ~n19227 & n20610 ;
  assign n20612 = ~n20605 & n20611 ;
  assign n20613 = n18589 | n19223 ;
  assign n20614 = ~n19224 & n20613 ;
  assign n20615 = n19219 | n19221 ;
  assign n20616 = ~n19222 & n20615 ;
  assign n20617 = n20614 & n20616 ;
  assign n20618 = n19215 | n19217 ;
  assign n20619 = ~n19218 & n20618 ;
  assign n20620 = n20616 & n20619 ;
  assign n20621 = n19211 | n19213 ;
  assign n20622 = ~n19214 & n20621 ;
  assign n20623 = n20619 & n20622 ;
  assign n20624 = n18644 & ~n19209 ;
  assign n20625 = n19210 | n20624 ;
  assign n20626 = n20622 & ~n20625 ;
  assign n20627 = ~n20622 & n20625 ;
  assign n20628 = n20626 | n20627 ;
  assign n20629 = n18660 & ~n19207 ;
  assign n20630 = n19208 | n20629 ;
  assign n20631 = n20625 | n20630 ;
  assign n20632 = n18675 | n19205 ;
  assign n20633 = ~n19206 & n20632 ;
  assign n20634 = ~n20630 & n20633 ;
  assign n20635 = n20630 & ~n20633 ;
  assign n20636 = n20634 | n20635 ;
  assign n20637 = ( ~n18691 & n18705 ) | ( ~n18691 & n19204 ) | ( n18705 & n19204 ) ;
  assign n20638 = n18691 & ~n18704 ;
  assign n20639 = ~n19204 & n20638 ;
  assign n20640 = n20637 | n20639 ;
  assign n20641 = n18708 & ~n19203 ;
  assign n20642 = n19204 | n20641 ;
  assign n20643 = ~n20640 & n20642 ;
  assign n20644 = ~n20633 & n20643 ;
  assign n20645 = n20640 | n20644 ;
  assign n20646 = n20636 | n20645 ;
  assign n20647 = ~n20634 & n20646 ;
  assign n20648 = n20625 & n20630 ;
  assign n20649 = n20631 & ~n20648 ;
  assign n20650 = ~n20647 & n20649 ;
  assign n20651 = n20631 & ~n20650 ;
  assign n20652 = n20628 | n20651 ;
  assign n20653 = ~n20626 & n20652 ;
  assign n20654 = n20619 | n20622 ;
  assign n20655 = ~n20623 & n20654 ;
  assign n20656 = ~n20653 & n20655 ;
  assign n20657 = n20623 | n20656 ;
  assign n20658 = n20616 | n20619 ;
  assign n20659 = ~n20620 & n20658 ;
  assign n20660 = n20657 & n20659 ;
  assign n20661 = n20620 | n20660 ;
  assign n20662 = n20614 | n20616 ;
  assign n20663 = ~n20617 & n20662 ;
  assign n20664 = n20661 & n20663 ;
  assign n20665 = n20617 | n20664 ;
  assign n20666 = ( n20611 & n20614 ) | ( n20611 & n20665 ) | ( n20614 & n20665 ) ;
  assign n20667 = n20605 & ~n20611 ;
  assign n20668 = n20612 | n20667 ;
  assign n20669 = n20666 & ~n20668 ;
  assign n20670 = n20612 | n20669 ;
  assign n20671 = ~n20608 & n20670 ;
  assign n20672 = n20606 | n20671 ;
  assign n20673 = ( n20601 & ~n20602 ) | ( n20601 & n20672 ) | ( ~n20602 & n20672 ) ;
  assign n20674 = ~n20597 & n20673 ;
  assign n20675 = n20596 & ~n20674 ;
  assign n20676 = ( ~n20588 & n20591 ) | ( ~n20588 & n20675 ) | ( n20591 & n20675 ) ;
  assign n20677 = n20580 & ~n20588 ;
  assign n20678 = ( n20580 & n20584 ) | ( n20580 & n20677 ) | ( n20584 & n20677 ) ;
  assign n20679 = ( ~n20589 & n20676 ) | ( ~n20589 & n20678 ) | ( n20676 & n20678 ) ;
  assign n20680 = n20585 & ~n20679 ;
  assign n20681 = n20569 & n20584 ;
  assign n20682 = ( n20569 & n20584 ) | ( n20569 & n20585 ) | ( n20584 & n20585 ) ;
  assign n20683 = ( ~n20680 & n20681 ) | ( ~n20680 & n20682 ) | ( n20681 & n20682 ) ;
  assign n20684 = n20576 & ~n20683 ;
  assign n20685 = n20574 & ~n20684 ;
  assign n20686 = ( n19262 & n19545 ) | ( n19262 & n19556 ) | ( n19545 & n19556 ) ;
  assign n20687 = ( n19262 & n19544 ) | ( n19262 & n19555 ) | ( n19544 & n19555 ) ;
  assign n20688 = n19345 & ~n20687 ;
  assign n20689 = n20686 | n20688 ;
  assign n20690 = n20573 & n20689 ;
  assign n20691 = ~n20560 & n20689 ;
  assign n20692 = n20690 | n20691 ;
  assign n20693 = n20560 & ~n20689 ;
  assign n20694 = n20573 | n20689 ;
  assign n20695 = ~n20693 & n20694 ;
  assign n20696 = ( n20685 & n20692 ) | ( n20685 & n20695 ) | ( n20692 & n20695 ) ;
  assign n20697 = n20565 & ~n20696 ;
  assign n20698 = ~n20552 & n20562 ;
  assign n20699 = n20563 | n20698 ;
  assign n20700 = n20552 & ~n20556 ;
  assign n20701 = n20699 & ~n20700 ;
  assign n20702 = n20552 & ~n20562 ;
  assign n20703 = n20700 | n20702 ;
  assign n20704 = ( n20697 & n20701 ) | ( n20697 & ~n20703 ) | ( n20701 & ~n20703 ) ;
  assign n20705 = ~n20557 & n20704 ;
  assign n20706 = n20557 | n20705 ;
  assign n20707 = ( n19561 & n20505 ) | ( n19561 & n20518 ) | ( n20505 & n20518 ) ;
  assign n20708 = ( n19561 & n20504 ) | ( n19561 & n20517 ) | ( n20504 & n20517 ) ;
  assign n20709 = n20468 & ~n20708 ;
  assign n20710 = n20707 | n20709 ;
  assign n20711 = ~n20546 & n20710 ;
  assign n20712 = ~n20556 & n20710 ;
  assign n20713 = n20711 | n20712 ;
  assign n20714 = n20546 & ~n20710 ;
  assign n20715 = n20556 & ~n20710 ;
  assign n20716 = ~n20714 & n20715 ;
  assign n20717 = n20714 | n20716 ;
  assign n20718 = ( n20706 & ~n20713 ) | ( n20706 & n20717 ) | ( ~n20713 & n20717 ) ;
  assign n20719 = ~n20548 & n20718 ;
  assign n20720 = ~n20547 & n20719 ;
  assign n20721 = ( n19561 & n20511 ) | ( n19561 & n20524 ) | ( n20511 & n20524 ) ;
  assign n20722 = ( n19561 & n20510 ) | ( n19561 & n20523 ) | ( n20510 & n20523 ) ;
  assign n20723 = n20306 & ~n20722 ;
  assign n20724 = n20721 | n20723 ;
  assign n20725 = n20542 & n20724 ;
  assign n20726 = n20536 & n20724 ;
  assign n20727 = n20725 | n20726 ;
  assign n20728 = n20542 | n20724 ;
  assign n20729 = ~n20725 & n20728 ;
  assign n20730 = n20547 & n20729 ;
  assign n20731 = n20728 & ~n20730 ;
  assign n20732 = ( n20536 & n20724 ) | ( n20536 & n20731 ) | ( n20724 & n20731 ) ;
  assign n20733 = ( ~n20720 & n20727 ) | ( ~n20720 & n20732 ) | ( n20727 & n20732 ) ;
  assign n20734 = n20538 | n20733 ;
  assign n20735 = n20537 | n20734 ;
  assign n20736 = ( n20071 & n20072 ) | ( n20071 & n20119 ) | ( n20072 & n20119 ) ;
  assign n20737 = n4548 | n4551 ;
  assign n20738 = n4546 | n20737 ;
  assign n20739 = ~n12314 & n20737 ;
  assign n20740 = ( ~n12318 & n20738 ) | ( ~n12318 & n20739 ) | ( n20738 & n20739 ) ;
  assign n20741 = n4554 | n20740 ;
  assign n20742 = n12615 & ~n20740 ;
  assign n20743 = ( n12314 & ~n12604 ) | ( n12314 & n20742 ) | ( ~n12604 & n20742 ) ;
  assign n20744 = n20741 & ~n20743 ;
  assign n20745 = x23 & ~n20744 ;
  assign n20746 = ~x23 & n20744 ;
  assign n20747 = n20745 | n20746 ;
  assign n20748 = n20091 | n20104 ;
  assign n20749 = n3478 | n3874 ;
  assign n20750 = n1845 | n2207 ;
  assign n20751 = n760 | n20750 ;
  assign n20752 = n20749 | n20751 ;
  assign n20753 = n482 | n1443 ;
  assign n20754 = n273 | n20753 ;
  assign n20755 = n381 | n20754 ;
  assign n20756 = n20752 | n20755 ;
  assign n20757 = n139 | n11195 ;
  assign n20758 = n20756 | n20757 ;
  assign n20759 = n197 | n11215 ;
  assign n20760 = n670 | n749 ;
  assign n20761 = n4873 | n20760 ;
  assign n20762 = n20759 | n20761 ;
  assign n20763 = n3549 | n20762 ;
  assign n20764 = n147 | n20763 ;
  assign n20765 = n19841 | n20764 ;
  assign n20766 = n20758 | n20765 ;
  assign n20767 = n3833 | n20766 ;
  assign n20768 = n807 | n1254 ;
  assign n20769 = ( ~n2483 & n3375 ) | ( ~n2483 & n20768 ) | ( n3375 & n20768 ) ;
  assign n20770 = n2483 | n20769 ;
  assign n20771 = n596 | n20770 ;
  assign n20772 = n393 | n20771 ;
  assign n20773 = n212 | n20772 ;
  assign n20774 = n20767 | n20773 ;
  assign n20775 = ~n20074 & n20774 ;
  assign n20776 = n20074 & ~n20774 ;
  assign n20777 = n20077 | n20775 ;
  assign n20778 = n20776 | n20777 ;
  assign n20779 = ( ~n20085 & n20088 ) | ( ~n20085 & n20778 ) | ( n20088 & n20778 ) ;
  assign n20780 = ( ~n20080 & n20777 ) | ( ~n20080 & n20779 ) | ( n20777 & n20779 ) ;
  assign n20781 = ~n20776 & n20780 ;
  assign n20782 = ~n20775 & n20781 ;
  assign n20783 = n20075 & ~n20086 ;
  assign n20784 = ( n20077 & ~n20080 ) | ( n20077 & n20783 ) | ( ~n20080 & n20783 ) ;
  assign n20785 = n20778 & ~n20784 ;
  assign n20786 = n20782 | n20785 ;
  assign n20787 = n3744 & ~n12344 ;
  assign n20788 = n3639 & n12553 ;
  assign n20789 = n3727 & n12340 ;
  assign n20790 = n20788 | n20789 ;
  assign n20791 = n20787 | n20790 ;
  assign n20792 = n3636 | n20791 ;
  assign n20793 = ( ~n13523 & n20791 ) | ( ~n13523 & n20792 ) | ( n20791 & n20792 ) ;
  assign n20794 = n20786 & n20793 ;
  assign n20795 = n20786 | n20793 ;
  assign n20796 = ~n20794 & n20795 ;
  assign n20797 = n4048 & ~n12335 ;
  assign n20798 = n4043 & ~n12586 ;
  assign n20799 = n4045 & n12580 ;
  assign n20800 = n20798 | n20799 ;
  assign n20801 = n20797 | n20800 ;
  assign n20802 = n4051 & ~n13585 ;
  assign n20803 = ~n13587 & n20802 ;
  assign n20804 = ( n4051 & n20801 ) | ( n4051 & ~n20803 ) | ( n20801 & ~n20803 ) ;
  assign n20805 = ~x29 & n20804 ;
  assign n20806 = x29 | n20805 ;
  assign n20807 = ( ~n20804 & n20805 ) | ( ~n20804 & n20806 ) | ( n20805 & n20806 ) ;
  assign n20808 = n20796 & n20807 ;
  assign n20809 = n20796 | n20807 ;
  assign n20810 = ~n20808 & n20809 ;
  assign n20811 = n4479 & ~n12325 ;
  assign n20812 = n4481 & ~n12328 ;
  assign n20813 = n20811 | n20812 ;
  assign n20814 = n4484 & n12608 ;
  assign n20815 = n20813 | n20814 ;
  assign n20816 = n4487 & n13570 ;
  assign n20817 = ( n4487 & n13568 ) | ( n4487 & n20816 ) | ( n13568 & n20816 ) ;
  assign n20818 = n20815 | n20817 ;
  assign n20819 = x26 | n20818 ;
  assign n20820 = ~x26 & n20819 ;
  assign n20821 = ( ~n20818 & n20819 ) | ( ~n20818 & n20820 ) | ( n20819 & n20820 ) ;
  assign n20822 = ( n20748 & n20810 ) | ( n20748 & n20821 ) | ( n20810 & n20821 ) ;
  assign n20823 = ( n20810 & n20821 ) | ( n20810 & ~n20822 ) | ( n20821 & ~n20822 ) ;
  assign n20824 = ( n20748 & ~n20822 ) | ( n20748 & n20823 ) | ( ~n20822 & n20823 ) ;
  assign n20825 = ( n20117 & n20747 ) | ( n20117 & ~n20824 ) | ( n20747 & ~n20824 ) ;
  assign n20826 = ( ~n20747 & n20824 ) | ( ~n20747 & n20825 ) | ( n20824 & n20825 ) ;
  assign n20827 = ( ~n20117 & n20825 ) | ( ~n20117 & n20826 ) | ( n20825 & n20826 ) ;
  assign n20828 = n20736 & n20827 ;
  assign n20829 = n20736 | n20827 ;
  assign n20830 = ~n20828 & n20829 ;
  assign n20831 = n20123 | n20515 ;
  assign n20832 = n20830 & n20831 ;
  assign n20833 = n20123 | n20528 ;
  assign n20834 = n20830 & n20833 ;
  assign n20835 = ( n19561 & n20832 ) | ( n19561 & n20834 ) | ( n20832 & n20834 ) ;
  assign n20836 = ( n19561 & n20831 ) | ( n19561 & n20833 ) | ( n20831 & n20833 ) ;
  assign n20837 = n20830 | n20836 ;
  assign n20838 = ~n20835 & n20837 ;
  assign n20839 = n20532 | n20838 ;
  assign n20840 = n4048 & ~n12325 ;
  assign n20841 = n4043 & n12580 ;
  assign n20842 = n4045 & ~n12335 ;
  assign n20843 = n20841 | n20842 ;
  assign n20844 = n20840 | n20843 ;
  assign n20845 = n4051 | n20844 ;
  assign n20846 = ( ~n13720 & n20844 ) | ( ~n13720 & n20845 ) | ( n20844 & n20845 ) ;
  assign n20847 = ~x29 & n20846 ;
  assign n20848 = x29 | n20847 ;
  assign n20849 = ( ~n20846 & n20847 ) | ( ~n20846 & n20848 ) | ( n20847 & n20848 ) ;
  assign n20850 = n19623 | n19628 ;
  assign n20851 = n711 | n11276 ;
  assign n20852 = n5792 | n20851 ;
  assign n20853 = n3904 | n20852 ;
  assign n20854 = n3902 | n20853 ;
  assign n20855 = n13942 | n20854 ;
  assign n20856 = n12657 | n20855 ;
  assign n20857 = n20850 | n20856 ;
  assign n20858 = n166 | n1054 ;
  assign n20859 = n3451 | n20858 ;
  assign n20860 = n806 | n20859 ;
  assign n20861 = n468 | n20860 ;
  assign n20862 = n300 | n20861 ;
  assign n20863 = n319 | n20862 ;
  assign n20864 = n449 | n20863 ;
  assign n20865 = n20857 | n20864 ;
  assign n20866 = n122 | n661 ;
  assign n20867 = n20865 | n20866 ;
  assign n20868 = n20774 | n20867 ;
  assign n20869 = n20774 & n20867 ;
  assign n20870 = n20868 & ~n20869 ;
  assign n20871 = n4554 | n20738 ;
  assign n20872 = ~n12314 & n20871 ;
  assign n20873 = ~x23 & n20872 ;
  assign n20874 = x23 | n20873 ;
  assign n20875 = ( ~n20872 & n20873 ) | ( ~n20872 & n20874 ) | ( n20873 & n20874 ) ;
  assign n20876 = n20870 & ~n20875 ;
  assign n20877 = ~n20870 & n20875 ;
  assign n20878 = n20876 | n20877 ;
  assign n20879 = n20781 | n20878 ;
  assign n20880 = n20781 & n20878 ;
  assign n20881 = n20879 & ~n20880 ;
  assign n20882 = n3744 & ~n12586 ;
  assign n20883 = n3639 & n12340 ;
  assign n20884 = n3727 & ~n12344 ;
  assign n20885 = n20883 | n20884 ;
  assign n20886 = n20882 | n20885 ;
  assign n20887 = ( n3636 & n13454 ) | ( n3636 & n13455 ) | ( n13454 & n13455 ) ;
  assign n20888 = n20886 | n20887 ;
  assign n20889 = n20881 & n20888 ;
  assign n20890 = n20881 & ~n20889 ;
  assign n20891 = n20888 & ~n20889 ;
  assign n20892 = n20890 | n20891 ;
  assign n20893 = n20794 | n20808 ;
  assign n20894 = ( n20849 & n20892 ) | ( n20849 & ~n20893 ) | ( n20892 & ~n20893 ) ;
  assign n20895 = ( ~n20892 & n20893 ) | ( ~n20892 & n20894 ) | ( n20893 & n20894 ) ;
  assign n20896 = ( ~n20849 & n20894 ) | ( ~n20849 & n20895 ) | ( n20894 & n20895 ) ;
  assign n20897 = n4484 & ~n12318 ;
  assign n20898 = n4479 & ~n12328 ;
  assign n20899 = n4481 & n12608 ;
  assign n20900 = n20898 | n20899 ;
  assign n20901 = n20897 | n20900 ;
  assign n20902 = n4487 | n20901 ;
  assign n20903 = ( n14320 & n20901 ) | ( n14320 & n20902 ) | ( n20901 & n20902 ) ;
  assign n20904 = x26 & n20903 ;
  assign n20905 = x26 & ~n20904 ;
  assign n20906 = ( n20903 & ~n20904 ) | ( n20903 & n20905 ) | ( ~n20904 & n20905 ) ;
  assign n20907 = ( ~n20822 & n20896 ) | ( ~n20822 & n20906 ) | ( n20896 & n20906 ) ;
  assign n20908 = ( n20822 & ~n20906 ) | ( n20822 & n20907 ) | ( ~n20906 & n20907 ) ;
  assign n20909 = ( ~n20896 & n20907 ) | ( ~n20896 & n20908 ) | ( n20907 & n20908 ) ;
  assign n20910 = ( n20117 & n20747 ) | ( n20117 & n20824 ) | ( n20747 & n20824 ) ;
  assign n20911 = n20909 & n20910 ;
  assign n20912 = n20909 | n20910 ;
  assign n20913 = ~n20911 & n20912 ;
  assign n20914 = n20828 | n20832 ;
  assign n20915 = n20913 & n20914 ;
  assign n20916 = n20828 | n20834 ;
  assign n20917 = n20913 & n20916 ;
  assign n20918 = ( n19561 & n20915 ) | ( n19561 & n20917 ) | ( n20915 & n20917 ) ;
  assign n20919 = ( n19561 & n20914 ) | ( n19561 & n20916 ) | ( n20914 & n20916 ) ;
  assign n20920 = n20913 | n20919 ;
  assign n20921 = ~n20918 & n20920 ;
  assign n20922 = n20838 | n20921 ;
  assign n20923 = n20839 & n20922 ;
  assign n20924 = n20532 & n20838 ;
  assign n20925 = n20839 & ~n20924 ;
  assign n20926 = n20537 & n20925 ;
  assign n20927 = n20924 | n20926 ;
  assign n20928 = ( n20838 & n20921 ) | ( n20838 & n20927 ) | ( n20921 & n20927 ) ;
  assign n20929 = ( ~n20735 & n20923 ) | ( ~n20735 & n20928 ) | ( n20923 & n20928 ) ;
  assign n20930 = n4481 & ~n12318 ;
  assign n20931 = n4479 & n12608 ;
  assign n20932 = n20930 | n20931 ;
  assign n20933 = n4484 & ~n12314 ;
  assign n20934 = n20932 | n20933 ;
  assign n20935 = n4487 | n20934 ;
  assign n20936 = ( ~n14302 & n20934 ) | ( ~n14302 & n20935 ) | ( n20934 & n20935 ) ;
  assign n20937 = ~x26 & n20936 ;
  assign n20938 = x26 | n20937 ;
  assign n20939 = ( ~n20936 & n20937 ) | ( ~n20936 & n20938 ) | ( n20937 & n20938 ) ;
  assign n20940 = ( n20849 & n20892 ) | ( n20849 & n20893 ) | ( n20892 & n20893 ) ;
  assign n20941 = n371 | n850 ;
  assign n20942 = n3544 | n20941 ;
  assign n20943 = n3528 | n20942 ;
  assign n20944 = ~n3494 & n3573 ;
  assign n20945 = ~n20943 & n20944 ;
  assign n20946 = n1054 | n2810 ;
  assign n20947 = n5674 | n20946 ;
  assign n20948 = n381 | n3375 ;
  assign n20949 = n610 | n20948 ;
  assign n20950 = n20947 | n20949 ;
  assign n20951 = n76 | n437 ;
  assign n20952 = n20950 | n20951 ;
  assign n20953 = n842 | n20952 ;
  assign n20954 = n2147 | n20953 ;
  assign n20955 = n405 | n20954 ;
  assign n20956 = n489 | n20955 ;
  assign n20957 = n20945 & ~n20956 ;
  assign n20958 = ~n1415 & n20957 ;
  assign n20959 = ( n20869 & n20876 ) | ( n20869 & n20958 ) | ( n20876 & n20958 ) ;
  assign n20960 = ( n20868 & n20869 ) | ( n20868 & ~n20875 ) | ( n20869 & ~n20875 ) ;
  assign n20961 = n20958 | n20960 ;
  assign n20962 = ~n20959 & n20961 ;
  assign n20963 = n3744 & n12580 ;
  assign n20964 = n3727 & ~n12586 ;
  assign n20965 = n3639 & ~n12344 ;
  assign n20966 = n20964 | n20965 ;
  assign n20967 = n20963 | n20966 ;
  assign n20968 = n3636 | n20967 ;
  assign n20969 = ( n13432 & n20967 ) | ( n13432 & n20968 ) | ( n20967 & n20968 ) ;
  assign n20970 = n20962 | n20969 ;
  assign n20971 = n20962 & n20969 ;
  assign n20972 = n20970 & ~n20971 ;
  assign n20973 = n20879 & ~n20972 ;
  assign n20974 = ~n20889 & n20973 ;
  assign n20975 = ( ~n20879 & n20889 ) | ( ~n20879 & n20972 ) | ( n20889 & n20972 ) ;
  assign n20976 = n20974 | n20975 ;
  assign n20977 = n4048 & ~n12328 ;
  assign n20978 = n4043 & ~n12335 ;
  assign n20979 = n4045 & ~n12325 ;
  assign n20980 = n20978 | n20979 ;
  assign n20981 = n20977 | n20980 ;
  assign n20982 = n4051 | n20981 ;
  assign n20983 = ( ~n13544 & n20981 ) | ( ~n13544 & n20982 ) | ( n20981 & n20982 ) ;
  assign n20984 = ~x29 & n20983 ;
  assign n20985 = x29 | n20984 ;
  assign n20986 = ( ~n20983 & n20984 ) | ( ~n20983 & n20985 ) | ( n20984 & n20985 ) ;
  assign n20987 = ~n20976 & n20986 ;
  assign n20988 = n20976 & ~n20986 ;
  assign n20989 = n20987 | n20988 ;
  assign n20990 = ( n20939 & n20940 ) | ( n20939 & ~n20989 ) | ( n20940 & ~n20989 ) ;
  assign n20991 = ( ~n20940 & n20989 ) | ( ~n20940 & n20990 ) | ( n20989 & n20990 ) ;
  assign n20992 = ( ~n20939 & n20990 ) | ( ~n20939 & n20991 ) | ( n20990 & n20991 ) ;
  assign n20993 = ( n20822 & n20896 ) | ( n20822 & n20906 ) | ( n20896 & n20906 ) ;
  assign n20994 = ~n20992 & n20993 ;
  assign n20995 = n20992 | n20994 ;
  assign n20996 = n20993 & ~n20994 ;
  assign n20997 = n20995 & ~n20996 ;
  assign n20998 = n20911 | n20915 ;
  assign n20999 = ~n20997 & n20998 ;
  assign n21000 = n20911 | n20917 ;
  assign n21001 = ~n20997 & n21000 ;
  assign n21002 = ( n19561 & n20999 ) | ( n19561 & n21001 ) | ( n20999 & n21001 ) ;
  assign n21003 = ( n19561 & n20998 ) | ( n19561 & n21000 ) | ( n20998 & n21000 ) ;
  assign n21004 = n20997 & ~n21003 ;
  assign n21005 = n21002 | n21004 ;
  assign n21006 = n20921 & ~n21005 ;
  assign n21007 = ~n20921 & n21005 ;
  assign n21008 = n20928 & ~n21007 ;
  assign n21009 = n20923 & ~n21007 ;
  assign n21010 = ( ~n20735 & n21008 ) | ( ~n20735 & n21009 ) | ( n21008 & n21009 ) ;
  assign n21011 = ~n21006 & n21010 ;
  assign n21012 = n20929 & ~n21011 ;
  assign n21013 = n21006 | n21011 ;
  assign n21014 = n21007 | n21013 ;
  assign n21015 = ~n21012 & n21014 ;
  assign n21016 = n9245 & ~n21005 ;
  assign n21017 = n8680 & n20838 ;
  assign n21018 = n8681 & n20921 ;
  assign n21019 = n21017 | n21018 ;
  assign n21020 = n21016 | n21019 ;
  assign n21021 = n8685 | n21020 ;
  assign n21022 = ( ~n21015 & n21020 ) | ( ~n21015 & n21021 ) | ( n21020 & n21021 ) ;
  assign n21023 = ~x5 & n21022 ;
  assign n21024 = x5 | n21023 ;
  assign n21025 = ( ~n21022 & n21023 ) | ( ~n21022 & n21024 ) | ( n21023 & n21024 ) ;
  assign n23208 = n5503 & ~n20536 ;
  assign n23209 = n5512 & ~n20542 ;
  assign n23210 = n5508 & ~n20724 ;
  assign n23211 = n23209 | n23210 ;
  assign n23212 = n23208 | n23211 ;
  assign n23213 = ~n20726 & n20733 ;
  assign n23214 = n20536 | n20724 ;
  assign n23215 = ~n20727 & n23214 ;
  assign n23216 = ( ~n20720 & n20725 ) | ( ~n20720 & n20731 ) | ( n20725 & n20731 ) ;
  assign n23217 = n23215 | n23216 ;
  assign n23218 = n5515 & n23217 ;
  assign n23219 = ~n23213 & n23218 ;
  assign n23220 = ( n5515 & n23212 ) | ( n5515 & ~n23219 ) | ( n23212 & ~n23219 ) ;
  assign n23221 = x8 & n23220 ;
  assign n23222 = x8 & ~n23221 ;
  assign n23223 = ( n23220 & ~n23221 ) | ( n23220 & n23222 ) | ( ~n23221 & n23222 ) ;
  assign n22635 = n7305 & ~n20710 ;
  assign n22636 = n7300 & ~n20552 ;
  assign n22637 = n7302 & n20556 ;
  assign n22638 = n22636 | n22637 ;
  assign n22639 = n22635 | n22638 ;
  assign n21033 = n20712 | n20715 ;
  assign n21034 = n20706 & ~n21033 ;
  assign n22640 = ~n20706 & n21033 ;
  assign n22641 = n21034 | n22640 ;
  assign n22642 = n7308 | n22639 ;
  assign n22643 = ( n22639 & ~n22641 ) | ( n22639 & n22642 ) | ( ~n22641 & n22642 ) ;
  assign n22644 = ~x11 & n22643 ;
  assign n22645 = x11 | n22644 ;
  assign n22646 = ( ~n22643 & n22644 ) | ( ~n22643 & n22645 ) | ( n22644 & n22645 ) ;
  assign n21043 = ~n20565 & n20696 ;
  assign n21044 = n20697 | n21043 ;
  assign n21045 = n7280 & n20562 ;
  assign n21046 = n5384 & ~n20689 ;
  assign n21047 = n7277 & n20560 ;
  assign n21048 = n21046 | n21047 ;
  assign n21049 = n21045 | n21048 ;
  assign n21050 = n39 | n21049 ;
  assign n21051 = ( ~n21044 & n21049 ) | ( ~n21044 & n21050 ) | ( n21049 & n21050 ) ;
  assign n21052 = ~x14 & n21051 ;
  assign n21053 = x14 | n21052 ;
  assign n21054 = ( ~n21051 & n21052 ) | ( ~n21051 & n21053 ) | ( n21052 & n21053 ) ;
  assign n21055 = n20653 & ~n20655 ;
  assign n21056 = n20656 | n21055 ;
  assign n21057 = n4479 & ~n20625 ;
  assign n21058 = n4481 | n21057 ;
  assign n21059 = ( n20622 & n21057 ) | ( n20622 & n21058 ) | ( n21057 & n21058 ) ;
  assign n21060 = n4484 | n21059 ;
  assign n21061 = ( n20619 & n21059 ) | ( n20619 & n21060 ) | ( n21059 & n21060 ) ;
  assign n21062 = n4487 | n21061 ;
  assign n21063 = ( ~n21056 & n21061 ) | ( ~n21056 & n21062 ) | ( n21061 & n21062 ) ;
  assign n21064 = ~x26 & n21063 ;
  assign n21065 = x26 & ~n21063 ;
  assign n21066 = n21064 | n21065 ;
  assign n21067 = ( x29 & n14554 ) | ( x29 & n20642 ) | ( n14554 & n20642 ) ;
  assign n21068 = n20640 & ~n20642 ;
  assign n21069 = n20643 | n21068 ;
  assign n21070 = n4051 & n21069 ;
  assign n21071 = n4045 & ~n20642 ;
  assign n21072 = n4048 & ~n20640 ;
  assign n21073 = n21071 | n21072 ;
  assign n21074 = n21070 | n21073 ;
  assign n21075 = x29 | n21074 ;
  assign n21076 = ~x29 & n21075 ;
  assign n21077 = ( ~n21074 & n21075 ) | ( ~n21074 & n21076 ) | ( n21075 & n21076 ) ;
  assign n21078 = n21067 & n21077 ;
  assign n21079 = n4048 & n20633 ;
  assign n21080 = n4043 & ~n20642 ;
  assign n21081 = n4045 & ~n20640 ;
  assign n21082 = n21080 | n21081 ;
  assign n21083 = n21079 | n21082 ;
  assign n21084 = n20633 & ~n20643 ;
  assign n21085 = n20644 | n21084 ;
  assign n21086 = n4051 & n21085 ;
  assign n21087 = n21083 | n21086 ;
  assign n21088 = ~x29 & n21087 ;
  assign n21089 = x29 | n21088 ;
  assign n21090 = ( ~n21087 & n21088 ) | ( ~n21087 & n21089 ) | ( n21088 & n21089 ) ;
  assign n21091 = n21078 & n21090 ;
  assign n21092 = n3635 & ~n20642 ;
  assign n21093 = n4048 & ~n20630 ;
  assign n21094 = n4043 & ~n20640 ;
  assign n21095 = n4045 & n20633 ;
  assign n21096 = n21094 | n21095 ;
  assign n21097 = n21093 | n21096 ;
  assign n21098 = n20636 & n20645 ;
  assign n21099 = n20646 & ~n21098 ;
  assign n21100 = n4051 | n21097 ;
  assign n21101 = ( n21097 & n21099 ) | ( n21097 & n21100 ) | ( n21099 & n21100 ) ;
  assign n21102 = x29 & n21101 ;
  assign n21103 = x29 & ~n21102 ;
  assign n21104 = ( n21101 & ~n21102 ) | ( n21101 & n21103 ) | ( ~n21102 & n21103 ) ;
  assign n21105 = ( n21091 & n21092 ) | ( n21091 & n21104 ) | ( n21092 & n21104 ) ;
  assign n21106 = ( n21092 & n21104 ) | ( n21092 & ~n21105 ) | ( n21104 & ~n21105 ) ;
  assign n21107 = ( n21091 & ~n21105 ) | ( n21091 & n21106 ) | ( ~n21105 & n21106 ) ;
  assign n21108 = n21066 & n21107 ;
  assign n21109 = n21066 | n21107 ;
  assign n21110 = ~n21108 & n21109 ;
  assign n21111 = n21078 | n21090 ;
  assign n21112 = ~n21091 & n21111 ;
  assign n21113 = n20628 & n20651 ;
  assign n21114 = n20652 & ~n21113 ;
  assign n21115 = n4484 & n20622 ;
  assign n21116 = n4479 & ~n20630 ;
  assign n21117 = n4481 & ~n20625 ;
  assign n21118 = n21116 | n21117 ;
  assign n21119 = n21115 | n21118 ;
  assign n21120 = n4487 | n21119 ;
  assign n21121 = ( n21114 & n21119 ) | ( n21114 & n21120 ) | ( n21119 & n21120 ) ;
  assign n21122 = x26 & n21121 ;
  assign n21123 = x26 | n21121 ;
  assign n21124 = ~n21122 & n21123 ;
  assign n21125 = n21112 & n21124 ;
  assign n21126 = n21067 | n21077 ;
  assign n21127 = ~n21078 & n21126 ;
  assign n21128 = n20647 & ~n20649 ;
  assign n21129 = n20650 | n21128 ;
  assign n21130 = n4484 & ~n20625 ;
  assign n21131 = n4479 & n20633 ;
  assign n21132 = n4481 & ~n20630 ;
  assign n21133 = n21131 | n21132 ;
  assign n21134 = n21130 | n21133 ;
  assign n21135 = n4487 | n21134 ;
  assign n21136 = ( ~n21129 & n21134 ) | ( ~n21129 & n21135 ) | ( n21134 & n21135 ) ;
  assign n21137 = ~x26 & n21136 ;
  assign n21138 = x26 | n21137 ;
  assign n21139 = ( ~n21136 & n21137 ) | ( ~n21136 & n21138 ) | ( n21137 & n21138 ) ;
  assign n21140 = n21127 & n21139 ;
  assign n21141 = n21127 | n21139 ;
  assign n21142 = ~n21140 & n21141 ;
  assign n21143 = ( x26 & n14786 ) | ( x26 & n20642 ) | ( n14786 & n20642 ) ;
  assign n21144 = n4487 & n21069 ;
  assign n21145 = n4481 & ~n20642 ;
  assign n21146 = n4484 & ~n20640 ;
  assign n21147 = n21145 | n21146 ;
  assign n21148 = n21144 | n21147 ;
  assign n21149 = x26 | n21148 ;
  assign n21150 = ~x26 & n21149 ;
  assign n21151 = ( ~n21148 & n21149 ) | ( ~n21148 & n21150 ) | ( n21149 & n21150 ) ;
  assign n21152 = n21143 & n21151 ;
  assign n21153 = n4041 & ~n20642 ;
  assign n21154 = n4484 & n20633 ;
  assign n21155 = n4479 & ~n20642 ;
  assign n21156 = n4481 & ~n20640 ;
  assign n21157 = n21155 | n21156 ;
  assign n21158 = n21154 | n21157 ;
  assign n21159 = n4487 & n21085 ;
  assign n21160 = n21158 | n21159 ;
  assign n21161 = ~x26 & n21160 ;
  assign n21162 = x26 | n21161 ;
  assign n21163 = ( ~n21160 & n21161 ) | ( ~n21160 & n21162 ) | ( n21161 & n21162 ) ;
  assign n21164 = n21153 & n21163 ;
  assign n21165 = n21152 & n21164 ;
  assign n21166 = n21152 & n21163 ;
  assign n21167 = n21153 | n21166 ;
  assign n21168 = ~n21165 & n21167 ;
  assign n21169 = n4484 & ~n20630 ;
  assign n21170 = n4479 & ~n20640 ;
  assign n21171 = n4481 & n20633 ;
  assign n21172 = n21170 | n21171 ;
  assign n21173 = n21169 | n21172 ;
  assign n21174 = n4487 | n21173 ;
  assign n21175 = ( n21099 & n21173 ) | ( n21099 & n21174 ) | ( n21173 & n21174 ) ;
  assign n21176 = x26 & n21175 ;
  assign n21177 = x26 | n21175 ;
  assign n21178 = ~n21176 & n21177 ;
  assign n21179 = n21168 & n21178 ;
  assign n21180 = n21165 | n21179 ;
  assign n21181 = n21142 & n21180 ;
  assign n21182 = n21140 | n21181 ;
  assign n21183 = n21124 & ~n21125 ;
  assign n21184 = ( n21112 & ~n21125 ) | ( n21112 & n21183 ) | ( ~n21125 & n21183 ) ;
  assign n21185 = n21182 & n21184 ;
  assign n21186 = n21125 | n21185 ;
  assign n21187 = n21110 & n21186 ;
  assign n21188 = n21108 | n21187 ;
  assign n21189 = n20657 | n20659 ;
  assign n21190 = ~n20660 & n21189 ;
  assign n21191 = n4479 & n20622 ;
  assign n21192 = n4481 | n21191 ;
  assign n21193 = ( n20619 & n21191 ) | ( n20619 & n21192 ) | ( n21191 & n21192 ) ;
  assign n21194 = n4484 | n21193 ;
  assign n21195 = ( n20616 & n21193 ) | ( n20616 & n21194 ) | ( n21193 & n21194 ) ;
  assign n21196 = n4487 | n21195 ;
  assign n21197 = ( n21190 & n21195 ) | ( n21190 & n21196 ) | ( n21195 & n21196 ) ;
  assign n21198 = x26 & n21197 ;
  assign n21199 = x26 & ~n21198 ;
  assign n21200 = ( n21197 & ~n21198 ) | ( n21197 & n21199 ) | ( ~n21198 & n21199 ) ;
  assign n21201 = n4048 & ~n20625 ;
  assign n21202 = n4043 & n20633 ;
  assign n21203 = n4045 & ~n20630 ;
  assign n21204 = n21202 | n21203 ;
  assign n21205 = n21201 | n21204 ;
  assign n21206 = n4051 | n21205 ;
  assign n21207 = ( ~n21129 & n21205 ) | ( ~n21129 & n21206 ) | ( n21205 & n21206 ) ;
  assign n21208 = ~x29 & n21207 ;
  assign n21209 = x29 & ~n21207 ;
  assign n21210 = n21208 | n21209 ;
  assign n21211 = n3727 & ~n20642 ;
  assign n21212 = n3636 | n21211 ;
  assign n21213 = ( n21069 & n21211 ) | ( n21069 & n21212 ) | ( n21211 & n21212 ) ;
  assign n21214 = n3744 & ~n20640 ;
  assign n21215 = n21213 | n21214 ;
  assign n21216 = n843 | n849 ;
  assign n21217 = n1260 | n2029 ;
  assign n21218 = n21216 | n21217 ;
  assign n21219 = n391 | n405 ;
  assign n21220 = n314 | n21219 ;
  assign n21221 = n21218 | n21220 ;
  assign n21222 = n346 | n351 ;
  assign n21223 = n444 | n21222 ;
  assign n21224 = n601 | n21223 ;
  assign n21225 = n110 | n21224 ;
  assign n21226 = n21221 | n21225 ;
  assign n21227 = ~n630 & n2685 ;
  assign n21228 = ~n652 & n21227 ;
  assign n21229 = ~n11699 & n21228 ;
  assign n21230 = n1044 | n13605 ;
  assign n21231 = n21229 & ~n21230 ;
  assign n21232 = n2147 | n4101 ;
  assign n21233 = n996 | n21232 ;
  assign n21234 = n834 | n21233 ;
  assign n21235 = n214 | n21234 ;
  assign n21236 = n21231 & ~n21235 ;
  assign n21237 = n1094 | n2072 ;
  assign n21238 = n3079 | n21237 ;
  assign n21239 = n14059 | n21238 ;
  assign n21240 = n364 | n379 ;
  assign n21241 = n438 | n21240 ;
  assign n21242 = n155 | n21241 ;
  assign n21243 = n21239 | n21242 ;
  assign n21244 = n21236 & ~n21243 ;
  assign n21245 = ~n21226 & n21244 ;
  assign n21246 = ~n13902 & n21245 ;
  assign n21247 = n806 | n1656 ;
  assign n21248 = n933 | n21247 ;
  assign n21249 = n1022 | n21248 ;
  assign n21250 = n1371 | n21249 ;
  assign n21251 = ( n1989 & ~n3877 ) | ( n1989 & n21250 ) | ( ~n3877 & n21250 ) ;
  assign n21252 = n3877 | n21251 ;
  assign n21253 = n435 | n21252 ;
  assign n21254 = n21246 & ~n21253 ;
  assign n21255 = n165 | n452 ;
  assign n21256 = n21254 & ~n21255 ;
  assign n21257 = n21215 | n21256 ;
  assign n21258 = ~n21256 & n21257 ;
  assign n21259 = ( ~n21215 & n21257 ) | ( ~n21215 & n21258 ) | ( n21257 & n21258 ) ;
  assign n21260 = n21210 & ~n21259 ;
  assign n21261 = ~n21210 & n21259 ;
  assign n21262 = n21260 | n21261 ;
  assign n21263 = ( ~n21105 & n21200 ) | ( ~n21105 & n21262 ) | ( n21200 & n21262 ) ;
  assign n21264 = ( n21105 & ~n21262 ) | ( n21105 & n21263 ) | ( ~n21262 & n21263 ) ;
  assign n21265 = ( ~n21200 & n21263 ) | ( ~n21200 & n21264 ) | ( n21263 & n21264 ) ;
  assign n21266 = n21188 & n21265 ;
  assign n21267 = n21188 | n21265 ;
  assign n21268 = ~n21266 & n21267 ;
  assign n21269 = n4551 & ~n20605 ;
  assign n21270 = n4546 & n20614 ;
  assign n21271 = n4548 & n20611 ;
  assign n21272 = n21270 | n21271 ;
  assign n21273 = n21269 | n21272 ;
  assign n21274 = ~n20666 & n20668 ;
  assign n21275 = n20669 | n21274 ;
  assign n21276 = n4554 | n21273 ;
  assign n21277 = ( n21273 & ~n21275 ) | ( n21273 & n21276 ) | ( ~n21275 & n21276 ) ;
  assign n21278 = ~x23 & n21277 ;
  assign n21279 = x23 | n21278 ;
  assign n21280 = ( ~n21277 & n21278 ) | ( ~n21277 & n21279 ) | ( n21278 & n21279 ) ;
  assign n21281 = ~n21268 & n21280 ;
  assign n21282 = n21268 & ~n21280 ;
  assign n21283 = n21281 | n21282 ;
  assign n21284 = n21110 | n21186 ;
  assign n21285 = ~n21187 & n21284 ;
  assign n21286 = n4551 & n20611 ;
  assign n21287 = n4546 & n20616 ;
  assign n21288 = n4548 & n20614 ;
  assign n21289 = n21287 | n21288 ;
  assign n21290 = n21286 | n21289 ;
  assign n21291 = n4554 | n21290 ;
  assign n21292 = ( n20614 & n20665 ) | ( n20614 & ~n20666 ) | ( n20665 & ~n20666 ) ;
  assign n21293 = ( n20611 & ~n20666 ) | ( n20611 & n21292 ) | ( ~n20666 & n21292 ) ;
  assign n21294 = ( n21290 & n21291 ) | ( n21290 & n21293 ) | ( n21291 & n21293 ) ;
  assign n21295 = x23 & n21294 ;
  assign n21296 = x23 & ~n21295 ;
  assign n21297 = ( n21294 & ~n21295 ) | ( n21294 & n21296 ) | ( ~n21295 & n21296 ) ;
  assign n21298 = n21285 & n21297 ;
  assign n21299 = n21182 | n21184 ;
  assign n21300 = ~n21185 & n21299 ;
  assign n21301 = n20661 | n20663 ;
  assign n21302 = ~n20664 & n21301 ;
  assign n21303 = n4551 & n20614 ;
  assign n21304 = n4546 & n20619 ;
  assign n21305 = n4548 | n21304 ;
  assign n21306 = ( n20616 & n21304 ) | ( n20616 & n21305 ) | ( n21304 & n21305 ) ;
  assign n21307 = n21303 | n21306 ;
  assign n21308 = n4554 | n21307 ;
  assign n21309 = ( n21302 & n21307 ) | ( n21302 & n21308 ) | ( n21307 & n21308 ) ;
  assign n21310 = x23 & n21309 ;
  assign n21311 = x23 & ~n21310 ;
  assign n21312 = ( n21309 & ~n21310 ) | ( n21309 & n21311 ) | ( ~n21310 & n21311 ) ;
  assign n21313 = n21300 & n21312 ;
  assign n21314 = n4546 & n20622 ;
  assign n21315 = n4548 | n21314 ;
  assign n21316 = ( n20619 & n21314 ) | ( n20619 & n21315 ) | ( n21314 & n21315 ) ;
  assign n21317 = n4551 | n21316 ;
  assign n21318 = ( n20616 & n21316 ) | ( n20616 & n21317 ) | ( n21316 & n21317 ) ;
  assign n21319 = n4554 | n21318 ;
  assign n21320 = ( n21190 & n21318 ) | ( n21190 & n21319 ) | ( n21318 & n21319 ) ;
  assign n21321 = ~x23 & n21320 ;
  assign n21322 = x23 & ~n21320 ;
  assign n21323 = n21321 | n21322 ;
  assign n21324 = n21142 | n21180 ;
  assign n21325 = ~n21181 & n21324 ;
  assign n21326 = n21323 & n21325 ;
  assign n21327 = n4546 & ~n20625 ;
  assign n21328 = n4548 | n21327 ;
  assign n21329 = ( n20622 & n21327 ) | ( n20622 & n21328 ) | ( n21327 & n21328 ) ;
  assign n21330 = n4551 | n21329 ;
  assign n21331 = ( n20619 & n21329 ) | ( n20619 & n21330 ) | ( n21329 & n21330 ) ;
  assign n21332 = n4554 | n21331 ;
  assign n21333 = ( ~n21056 & n21331 ) | ( ~n21056 & n21332 ) | ( n21331 & n21332 ) ;
  assign n21334 = ~x23 & n21333 ;
  assign n21335 = x23 | n21334 ;
  assign n21336 = ( ~n21333 & n21334 ) | ( ~n21333 & n21335 ) | ( n21334 & n21335 ) ;
  assign n21337 = n21168 & ~n21179 ;
  assign n21338 = ( n21178 & ~n21179 ) | ( n21178 & n21337 ) | ( ~n21179 & n21337 ) ;
  assign n21339 = n21336 & n21338 ;
  assign n21340 = n21336 | n21338 ;
  assign n21341 = ~n21339 & n21340 ;
  assign n21342 = n21152 | n21163 ;
  assign n21343 = ~n21166 & n21342 ;
  assign n21344 = n4551 & n20622 ;
  assign n21345 = n4546 & ~n20630 ;
  assign n21346 = n4548 & ~n20625 ;
  assign n21347 = n21345 | n21346 ;
  assign n21348 = n21344 | n21347 ;
  assign n21349 = n4554 | n21348 ;
  assign n21350 = ( n21114 & n21348 ) | ( n21114 & n21349 ) | ( n21348 & n21349 ) ;
  assign n21351 = x23 & n21350 ;
  assign n21352 = x23 | n21350 ;
  assign n21353 = ~n21351 & n21352 ;
  assign n21354 = n21343 & n21353 ;
  assign n21355 = n21143 | n21151 ;
  assign n21356 = ~n21152 & n21355 ;
  assign n21357 = n4551 & ~n20625 ;
  assign n21358 = n4546 & n20633 ;
  assign n21359 = n4548 & ~n20630 ;
  assign n21360 = n21358 | n21359 ;
  assign n21361 = n21357 | n21360 ;
  assign n21362 = n4554 | n21361 ;
  assign n21363 = ( ~n21129 & n21361 ) | ( ~n21129 & n21362 ) | ( n21361 & n21362 ) ;
  assign n21364 = ~x23 & n21363 ;
  assign n21365 = x23 | n21364 ;
  assign n21366 = ( ~n21363 & n21364 ) | ( ~n21363 & n21365 ) | ( n21364 & n21365 ) ;
  assign n21367 = n21356 & n21366 ;
  assign n21368 = n21356 | n21366 ;
  assign n21369 = ~n21367 & n21368 ;
  assign n21370 = ( x23 & n15093 ) | ( x23 & n20642 ) | ( n15093 & n20642 ) ;
  assign n21371 = n4554 & n21069 ;
  assign n21372 = n4548 & ~n20642 ;
  assign n21373 = n4551 & ~n20640 ;
  assign n21374 = n21372 | n21373 ;
  assign n21375 = n21371 | n21374 ;
  assign n21376 = x23 | n21375 ;
  assign n21377 = ~x23 & n21376 ;
  assign n21378 = ( ~n21375 & n21376 ) | ( ~n21375 & n21377 ) | ( n21376 & n21377 ) ;
  assign n21379 = n21370 & n21378 ;
  assign n21380 = n4474 & ~n20642 ;
  assign n21381 = n4551 & n20633 ;
  assign n21382 = n4546 & ~n20642 ;
  assign n21383 = n4548 & ~n20640 ;
  assign n21384 = n21382 | n21383 ;
  assign n21385 = n21381 | n21384 ;
  assign n21386 = n4554 & n21085 ;
  assign n21387 = n21385 | n21386 ;
  assign n21388 = ~x23 & n21387 ;
  assign n21389 = x23 | n21388 ;
  assign n21390 = ( ~n21387 & n21388 ) | ( ~n21387 & n21389 ) | ( n21388 & n21389 ) ;
  assign n21391 = n21380 & n21390 ;
  assign n21392 = n21379 & n21391 ;
  assign n21393 = n21379 & n21390 ;
  assign n21394 = n21380 | n21393 ;
  assign n21395 = ~n21392 & n21394 ;
  assign n21396 = n4551 & ~n20630 ;
  assign n21397 = n4546 & ~n20640 ;
  assign n21398 = n4548 & n20633 ;
  assign n21399 = n21397 | n21398 ;
  assign n21400 = n21396 | n21399 ;
  assign n21401 = n4554 | n21400 ;
  assign n21402 = ( n21099 & n21400 ) | ( n21099 & n21401 ) | ( n21400 & n21401 ) ;
  assign n21403 = x23 & n21402 ;
  assign n21404 = x23 | n21402 ;
  assign n21405 = ~n21403 & n21404 ;
  assign n21406 = n21395 & n21405 ;
  assign n21407 = n21392 | n21406 ;
  assign n21408 = n21369 & n21407 ;
  assign n21409 = n21367 | n21408 ;
  assign n21410 = n21353 & ~n21354 ;
  assign n21411 = ( n21343 & ~n21354 ) | ( n21343 & n21410 ) | ( ~n21354 & n21410 ) ;
  assign n21412 = n21409 & n21411 ;
  assign n21413 = n21354 | n21412 ;
  assign n21414 = n21341 & n21413 ;
  assign n21415 = n21339 | n21414 ;
  assign n21416 = n21323 | n21325 ;
  assign n21417 = ~n21326 & n21416 ;
  assign n21418 = n21415 & n21417 ;
  assign n21419 = n21326 | n21418 ;
  assign n21420 = n21300 & ~n21313 ;
  assign n21421 = n21312 & ~n21313 ;
  assign n21422 = n21420 | n21421 ;
  assign n21423 = n21419 & n21422 ;
  assign n21424 = n21313 | n21423 ;
  assign n21425 = n21285 | n21297 ;
  assign n21426 = ~n21298 & n21425 ;
  assign n21427 = n21424 & n21426 ;
  assign n21428 = n21298 | n21427 ;
  assign n21429 = ~n21283 & n21428 ;
  assign n21430 = n21281 | n21429 ;
  assign n21431 = n20608 & ~n20670 ;
  assign n21432 = n20671 | n21431 ;
  assign n21433 = n4551 & n20600 ;
  assign n21434 = n4546 & n20611 ;
  assign n21435 = n4548 & ~n20605 ;
  assign n21436 = n21434 | n21435 ;
  assign n21437 = n21433 | n21436 ;
  assign n21438 = n4554 | n21437 ;
  assign n21439 = ( ~n21432 & n21437 ) | ( ~n21432 & n21438 ) | ( n21437 & n21438 ) ;
  assign n21440 = ~x23 & n21439 ;
  assign n21441 = x23 | n21440 ;
  assign n21442 = ( ~n21439 & n21440 ) | ( ~n21439 & n21441 ) | ( n21440 & n21441 ) ;
  assign n21443 = ( n21188 & n21200 ) | ( n21188 & n21268 ) | ( n21200 & n21268 ) ;
  assign n21444 = n4484 & n20614 ;
  assign n21445 = n4479 & n20619 ;
  assign n21446 = n4481 | n21445 ;
  assign n21447 = ( n20616 & n21445 ) | ( n20616 & n21446 ) | ( n21445 & n21446 ) ;
  assign n21448 = n21444 | n21447 ;
  assign n21449 = n4487 | n21448 ;
  assign n21450 = ( n21302 & n21448 ) | ( n21302 & n21449 ) | ( n21448 & n21449 ) ;
  assign n21451 = x26 & n21450 ;
  assign n21452 = x26 & ~n21451 ;
  assign n21453 = ( n21450 & ~n21451 ) | ( n21450 & n21452 ) | ( ~n21451 & n21452 ) ;
  assign n21454 = n4048 & n20622 ;
  assign n21455 = n4043 & ~n20630 ;
  assign n21456 = n4045 & ~n20625 ;
  assign n21457 = n21455 | n21456 ;
  assign n21458 = n21454 | n21457 ;
  assign n21459 = n4051 | n21458 ;
  assign n21460 = ( n21114 & n21458 ) | ( n21114 & n21459 ) | ( n21458 & n21459 ) ;
  assign n21461 = x29 & n21460 ;
  assign n21462 = x29 | n21460 ;
  assign n21463 = ~n21461 & n21462 ;
  assign n21464 = n3636 & n21085 ;
  assign n21465 = n3744 & n20633 ;
  assign n21466 = n3639 & ~n20642 ;
  assign n21467 = n3727 & ~n20640 ;
  assign n21468 = n21466 | n21467 ;
  assign n21469 = n21465 | n21468 ;
  assign n21470 = n21464 | n21469 ;
  assign n21471 = ~n3088 & n4280 ;
  assign n21472 = ~n1578 & n21471 ;
  assign n21473 = ~n1372 & n21472 ;
  assign n21474 = n181 | n270 ;
  assign n21475 = n186 | n21474 ;
  assign n21476 = n3371 | n13189 ;
  assign n21477 = n21475 | n21476 ;
  assign n21478 = n11213 | n21477 ;
  assign n21479 = n86 | n11528 ;
  assign n21480 = ( ~n5568 & n21478 ) | ( ~n5568 & n21479 ) | ( n21478 & n21479 ) ;
  assign n21481 = n5568 | n21480 ;
  assign n21482 = n21473 & ~n21481 ;
  assign n21483 = ~n1115 & n21482 ;
  assign n21484 = n335 | n13902 ;
  assign n21485 = n21483 & ~n21484 ;
  assign n21486 = n351 | n505 ;
  assign n21487 = n444 | n21486 ;
  assign n21488 = n52 | n21487 ;
  assign n21489 = n58 | n21488 ;
  assign n21490 = n21485 & ~n21489 ;
  assign n21491 = n21258 & ~n21490 ;
  assign n21492 = ~n21258 & n21490 ;
  assign n21493 = n21491 | n21492 ;
  assign n21494 = n21470 & ~n21493 ;
  assign n21495 = n21470 & ~n21494 ;
  assign n21496 = n21493 | n21494 ;
  assign n21497 = ~n21495 & n21496 ;
  assign n21498 = n21463 & ~n21497 ;
  assign n21499 = n21497 | n21498 ;
  assign n21500 = ( ~n21463 & n21498 ) | ( ~n21463 & n21499 ) | ( n21498 & n21499 ) ;
  assign n21501 = ( n21105 & n21210 ) | ( n21105 & ~n21259 ) | ( n21210 & ~n21259 ) ;
  assign n21502 = n21500 & ~n21501 ;
  assign n21503 = ~n21500 & n21501 ;
  assign n21504 = n21502 | n21503 ;
  assign n21505 = n21453 & ~n21504 ;
  assign n21506 = n21504 | n21505 ;
  assign n21507 = ( ~n21453 & n21505 ) | ( ~n21453 & n21506 ) | ( n21505 & n21506 ) ;
  assign n21508 = n21443 & ~n21507 ;
  assign n21509 = n21443 & ~n21508 ;
  assign n21510 = n21507 | n21508 ;
  assign n21511 = ~n21509 & n21510 ;
  assign n21512 = n21442 & ~n21511 ;
  assign n21513 = n21511 | n21512 ;
  assign n21514 = ( ~n21442 & n21512 ) | ( ~n21442 & n21513 ) | ( n21512 & n21513 ) ;
  assign n21515 = n21430 & ~n21514 ;
  assign n21516 = ~n21430 & n21514 ;
  assign n21517 = n21515 | n21516 ;
  assign n21518 = n4781 & n20588 ;
  assign n21519 = n4776 & ~n20595 ;
  assign n21520 = n4778 & ~n20591 ;
  assign n21521 = n21519 | n21520 ;
  assign n21522 = n21518 | n21521 ;
  assign n21523 = n4784 | n21522 ;
  assign n21524 = ( n20588 & ~n20591 ) | ( n20588 & n20675 ) | ( ~n20591 & n20675 ) ;
  assign n21525 = ( n20591 & ~n20675 ) | ( n20591 & n21524 ) | ( ~n20675 & n21524 ) ;
  assign n21526 = ( ~n20588 & n21524 ) | ( ~n20588 & n21525 ) | ( n21524 & n21525 ) ;
  assign n21527 = ( n21522 & n21523 ) | ( n21522 & n21526 ) | ( n21523 & n21526 ) ;
  assign n21528 = x20 & n21527 ;
  assign n21529 = x20 & ~n21528 ;
  assign n21530 = ( n21527 & ~n21528 ) | ( n21527 & n21529 ) | ( ~n21528 & n21529 ) ;
  assign n21531 = ~n21517 & n21530 ;
  assign n21532 = n21283 & ~n21428 ;
  assign n21533 = n21429 | n21532 ;
  assign n21534 = n4781 & ~n20591 ;
  assign n21535 = n4776 & n20600 ;
  assign n21536 = n4778 & ~n20595 ;
  assign n21537 = n21535 | n21536 ;
  assign n21538 = n21534 | n21537 ;
  assign n21539 = ~n20597 & n20675 ;
  assign n21540 = n20601 | n20602 ;
  assign n21541 = n20672 & ~n21540 ;
  assign n21542 = n20596 & n20674 ;
  assign n21543 = ( n20601 & n21541 ) | ( n20601 & ~n21542 ) | ( n21541 & ~n21542 ) ;
  assign n21544 = n4784 & ~n21543 ;
  assign n21545 = ~n21539 & n21544 ;
  assign n21546 = ( n4784 & n21538 ) | ( n4784 & ~n21545 ) | ( n21538 & ~n21545 ) ;
  assign n21547 = ~x20 & n21546 ;
  assign n21548 = x20 | n21547 ;
  assign n21549 = ( ~n21546 & n21547 ) | ( ~n21546 & n21548 ) | ( n21547 & n21548 ) ;
  assign n21550 = ~n21533 & n21549 ;
  assign n21551 = n21424 | n21426 ;
  assign n21552 = ~n21427 & n21551 ;
  assign n21553 = ~n20672 & n21540 ;
  assign n21554 = n21541 | n21553 ;
  assign n21555 = n4781 & ~n20595 ;
  assign n21556 = n4776 & ~n20605 ;
  assign n21557 = n4778 & n20600 ;
  assign n21558 = n21556 | n21557 ;
  assign n21559 = n21555 | n21558 ;
  assign n21560 = n4784 | n21559 ;
  assign n21561 = ( ~n21554 & n21559 ) | ( ~n21554 & n21560 ) | ( n21559 & n21560 ) ;
  assign n21562 = ~x20 & n21561 ;
  assign n21563 = x20 | n21562 ;
  assign n21564 = ( ~n21561 & n21562 ) | ( ~n21561 & n21563 ) | ( n21562 & n21563 ) ;
  assign n21565 = n21552 & n21564 ;
  assign n21566 = n21564 & ~n21565 ;
  assign n21567 = ( n21552 & ~n21565 ) | ( n21552 & n21566 ) | ( ~n21565 & n21566 ) ;
  assign n21568 = n21419 & ~n21423 ;
  assign n21569 = n21422 & ~n21423 ;
  assign n21570 = n21568 | n21569 ;
  assign n21571 = n4781 & n20600 ;
  assign n21572 = n4776 & n20611 ;
  assign n21573 = n4778 & ~n20605 ;
  assign n21574 = n21572 | n21573 ;
  assign n21575 = n21571 | n21574 ;
  assign n21576 = n4784 | n21575 ;
  assign n21577 = ( ~n21432 & n21575 ) | ( ~n21432 & n21576 ) | ( n21575 & n21576 ) ;
  assign n21578 = ~x20 & n21577 ;
  assign n21579 = x20 | n21578 ;
  assign n21580 = ( ~n21577 & n21578 ) | ( ~n21577 & n21579 ) | ( n21578 & n21579 ) ;
  assign n21581 = n21570 & n21580 ;
  assign n21582 = n21570 & ~n21581 ;
  assign n21583 = ~n21570 & n21580 ;
  assign n21584 = n21582 | n21583 ;
  assign n21585 = n21415 | n21417 ;
  assign n21586 = ~n21418 & n21585 ;
  assign n21587 = n4781 & ~n20605 ;
  assign n21588 = n4776 & n20614 ;
  assign n21589 = n4778 & n20611 ;
  assign n21590 = n21588 | n21589 ;
  assign n21591 = n21587 | n21590 ;
  assign n21592 = n4784 | n21591 ;
  assign n21593 = ( ~n21275 & n21591 ) | ( ~n21275 & n21592 ) | ( n21591 & n21592 ) ;
  assign n21594 = ~x20 & n21593 ;
  assign n21595 = x20 | n21594 ;
  assign n21596 = ( ~n21593 & n21594 ) | ( ~n21593 & n21595 ) | ( n21594 & n21595 ) ;
  assign n21597 = n21586 & n21596 ;
  assign n21598 = n21341 | n21413 ;
  assign n21599 = ~n21414 & n21598 ;
  assign n21600 = n4781 & n20611 ;
  assign n21601 = n4776 & n20616 ;
  assign n21602 = n4778 & n20614 ;
  assign n21603 = n21601 | n21602 ;
  assign n21604 = n21600 | n21603 ;
  assign n21605 = n4784 | n21604 ;
  assign n21606 = ( n21293 & n21604 ) | ( n21293 & n21605 ) | ( n21604 & n21605 ) ;
  assign n21607 = x20 & n21606 ;
  assign n21608 = x20 & ~n21607 ;
  assign n21609 = ( n21606 & ~n21607 ) | ( n21606 & n21608 ) | ( ~n21607 & n21608 ) ;
  assign n21610 = n21599 & n21609 ;
  assign n21611 = n21409 | n21411 ;
  assign n21612 = ~n21412 & n21611 ;
  assign n21613 = n4781 & n20614 ;
  assign n21614 = n4776 & n20619 ;
  assign n21615 = n4778 | n21614 ;
  assign n21616 = ( n20616 & n21614 ) | ( n20616 & n21615 ) | ( n21614 & n21615 ) ;
  assign n21617 = n21613 | n21616 ;
  assign n21618 = n4784 | n21617 ;
  assign n21619 = ( n21302 & n21617 ) | ( n21302 & n21618 ) | ( n21617 & n21618 ) ;
  assign n21620 = x20 & n21619 ;
  assign n21621 = x20 & ~n21620 ;
  assign n21622 = ( n21619 & ~n21620 ) | ( n21619 & n21621 ) | ( ~n21620 & n21621 ) ;
  assign n21623 = n21612 & n21622 ;
  assign n21624 = n4776 & n20622 ;
  assign n21625 = n4778 | n21624 ;
  assign n21626 = ( n20619 & n21624 ) | ( n20619 & n21625 ) | ( n21624 & n21625 ) ;
  assign n21627 = n4781 | n21626 ;
  assign n21628 = ( n20616 & n21626 ) | ( n20616 & n21627 ) | ( n21626 & n21627 ) ;
  assign n21629 = n4784 | n21628 ;
  assign n21630 = ( n21190 & n21628 ) | ( n21190 & n21629 ) | ( n21628 & n21629 ) ;
  assign n21631 = ~x20 & n21630 ;
  assign n21632 = x20 & ~n21630 ;
  assign n21633 = n21631 | n21632 ;
  assign n21634 = n21369 | n21407 ;
  assign n21635 = ~n21408 & n21634 ;
  assign n21636 = n21633 & n21635 ;
  assign n21637 = n4776 & ~n20625 ;
  assign n21638 = n4778 | n21637 ;
  assign n21639 = ( n20622 & n21637 ) | ( n20622 & n21638 ) | ( n21637 & n21638 ) ;
  assign n21640 = n4781 | n21639 ;
  assign n21641 = ( n20619 & n21639 ) | ( n20619 & n21640 ) | ( n21639 & n21640 ) ;
  assign n21642 = n4784 | n21641 ;
  assign n21643 = ( ~n21056 & n21641 ) | ( ~n21056 & n21642 ) | ( n21641 & n21642 ) ;
  assign n21644 = ~x20 & n21643 ;
  assign n21645 = x20 | n21644 ;
  assign n21646 = ( ~n21643 & n21644 ) | ( ~n21643 & n21645 ) | ( n21644 & n21645 ) ;
  assign n21647 = n21395 & ~n21406 ;
  assign n21648 = ( n21405 & ~n21406 ) | ( n21405 & n21647 ) | ( ~n21406 & n21647 ) ;
  assign n21649 = n21646 & n21648 ;
  assign n21650 = n21646 | n21648 ;
  assign n21651 = ~n21649 & n21650 ;
  assign n21652 = n21379 | n21390 ;
  assign n21653 = ~n21393 & n21652 ;
  assign n21654 = n4781 & n20622 ;
  assign n21655 = n4776 & ~n20630 ;
  assign n21656 = n4778 & ~n20625 ;
  assign n21657 = n21655 | n21656 ;
  assign n21658 = n21654 | n21657 ;
  assign n21659 = n4784 | n21658 ;
  assign n21660 = ( n21114 & n21658 ) | ( n21114 & n21659 ) | ( n21658 & n21659 ) ;
  assign n21661 = x20 & n21660 ;
  assign n21662 = x20 | n21660 ;
  assign n21663 = ~n21661 & n21662 ;
  assign n21664 = n21653 & n21663 ;
  assign n21665 = n21370 | n21378 ;
  assign n21666 = ~n21379 & n21665 ;
  assign n21667 = n4781 & ~n20625 ;
  assign n21668 = n4776 & n20633 ;
  assign n21669 = n4778 & ~n20630 ;
  assign n21670 = n21668 | n21669 ;
  assign n21671 = n21667 | n21670 ;
  assign n21672 = n4784 | n21671 ;
  assign n21673 = ( ~n21129 & n21671 ) | ( ~n21129 & n21672 ) | ( n21671 & n21672 ) ;
  assign n21674 = ~x20 & n21673 ;
  assign n21675 = x20 | n21674 ;
  assign n21676 = ( ~n21673 & n21674 ) | ( ~n21673 & n21675 ) | ( n21674 & n21675 ) ;
  assign n21677 = n21666 & n21676 ;
  assign n21678 = n21666 | n21676 ;
  assign n21679 = ~n21677 & n21678 ;
  assign n21680 = ( x20 & n15479 ) | ( x20 & n20642 ) | ( n15479 & n20642 ) ;
  assign n21681 = n4784 & n21069 ;
  assign n21682 = n4778 & ~n20642 ;
  assign n21683 = n4781 & ~n20640 ;
  assign n21684 = n21682 | n21683 ;
  assign n21685 = n21681 | n21684 ;
  assign n21686 = x20 | n21685 ;
  assign n21687 = ~x20 & n21686 ;
  assign n21688 = ( ~n21685 & n21686 ) | ( ~n21685 & n21687 ) | ( n21686 & n21687 ) ;
  assign n21689 = n21680 & n21688 ;
  assign n21690 = n4541 & ~n20642 ;
  assign n21691 = n4781 & n20633 ;
  assign n21692 = n4776 & ~n20642 ;
  assign n21693 = n4778 & ~n20640 ;
  assign n21694 = n21692 | n21693 ;
  assign n21695 = n21691 | n21694 ;
  assign n21696 = n4784 & n21085 ;
  assign n21697 = n21695 | n21696 ;
  assign n21698 = ~x20 & n21697 ;
  assign n21699 = x20 | n21698 ;
  assign n21700 = ( ~n21697 & n21698 ) | ( ~n21697 & n21699 ) | ( n21698 & n21699 ) ;
  assign n21701 = n21690 & n21700 ;
  assign n21702 = n21689 & n21701 ;
  assign n21703 = n21689 & n21700 ;
  assign n21704 = n21690 | n21703 ;
  assign n21705 = ~n21702 & n21704 ;
  assign n21706 = n4781 & ~n20630 ;
  assign n21707 = n4776 & ~n20640 ;
  assign n21708 = n4778 & n20633 ;
  assign n21709 = n21707 | n21708 ;
  assign n21710 = n21706 | n21709 ;
  assign n21711 = n4784 | n21710 ;
  assign n21712 = ( n21099 & n21710 ) | ( n21099 & n21711 ) | ( n21710 & n21711 ) ;
  assign n21713 = x20 & n21712 ;
  assign n21714 = x20 | n21712 ;
  assign n21715 = ~n21713 & n21714 ;
  assign n21716 = n21705 & n21715 ;
  assign n21717 = n21702 | n21716 ;
  assign n21718 = n21679 & n21717 ;
  assign n21719 = n21677 | n21718 ;
  assign n21720 = n21663 & ~n21664 ;
  assign n21721 = ( n21653 & ~n21664 ) | ( n21653 & n21720 ) | ( ~n21664 & n21720 ) ;
  assign n21722 = n21719 & n21721 ;
  assign n21723 = n21664 | n21722 ;
  assign n21724 = n21651 & n21723 ;
  assign n21725 = n21649 | n21724 ;
  assign n21726 = n21633 | n21635 ;
  assign n21727 = ~n21636 & n21726 ;
  assign n21728 = n21725 & n21727 ;
  assign n21729 = n21636 | n21728 ;
  assign n21730 = n21612 & ~n21623 ;
  assign n21731 = n21622 & ~n21623 ;
  assign n21732 = n21730 | n21731 ;
  assign n21733 = n21729 & n21732 ;
  assign n21734 = n21623 | n21733 ;
  assign n21735 = n21609 & ~n21610 ;
  assign n21736 = ( n21599 & ~n21610 ) | ( n21599 & n21735 ) | ( ~n21610 & n21735 ) ;
  assign n21737 = n21734 & n21736 ;
  assign n21738 = n21586 | n21596 ;
  assign n21739 = ~n21597 & n21738 ;
  assign n21740 = ( n21610 & n21737 ) | ( n21610 & n21739 ) | ( n21737 & n21739 ) ;
  assign n21741 = n21597 | n21740 ;
  assign n21742 = n21584 & n21741 ;
  assign n21743 = n21581 | n21742 ;
  assign n21744 = n21567 & n21743 ;
  assign n21745 = n21565 | n21744 ;
  assign n21746 = n21533 | n21550 ;
  assign n21747 = ( ~n21549 & n21550 ) | ( ~n21549 & n21746 ) | ( n21550 & n21746 ) ;
  assign n21748 = n21745 & ~n21747 ;
  assign n21749 = n21550 | n21748 ;
  assign n21750 = n21517 | n21531 ;
  assign n21751 = ( ~n21530 & n21531 ) | ( ~n21530 & n21750 ) | ( n21531 & n21750 ) ;
  assign n21752 = n21749 & ~n21751 ;
  assign n21753 = n21531 | n21752 ;
  assign n21754 = n21505 | n21508 ;
  assign n21755 = n4043 & ~n20625 ;
  assign n21756 = n4045 | n21755 ;
  assign n21757 = ( n20622 & n21755 ) | ( n20622 & n21756 ) | ( n21755 & n21756 ) ;
  assign n21758 = n4048 | n21757 ;
  assign n21759 = ( n20619 & n21757 ) | ( n20619 & n21758 ) | ( n21757 & n21758 ) ;
  assign n21760 = n4051 | n21759 ;
  assign n21761 = ( ~n21056 & n21759 ) | ( ~n21056 & n21760 ) | ( n21759 & n21760 ) ;
  assign n21762 = ~x29 & n21761 ;
  assign n21763 = x29 & ~n21761 ;
  assign n21764 = n21762 | n21763 ;
  assign n21765 = n3744 & ~n20630 ;
  assign n21766 = n3727 & n20633 ;
  assign n21767 = n3639 & ~n20640 ;
  assign n21768 = n21766 | n21767 ;
  assign n21769 = n21765 | n21768 ;
  assign n21770 = n3636 | n21769 ;
  assign n21771 = ( n21099 & n21769 ) | ( n21099 & n21770 ) | ( n21769 & n21770 ) ;
  assign n21772 = n21491 | n21494 ;
  assign n21773 = n266 | n519 ;
  assign n21774 = n718 | n21773 ;
  assign n21775 = n1807 | n4077 ;
  assign n21776 = n21774 | n21775 ;
  assign n21777 = n703 | n21776 ;
  assign n21778 = n1571 | n3658 ;
  assign n21779 = n4382 | n21778 ;
  assign n21780 = n21777 | n21779 ;
  assign n21781 = n1270 | n4348 ;
  assign n21782 = n21780 | n21781 ;
  assign n21783 = n808 | n2219 ;
  assign n21784 = n166 | n21783 ;
  assign n21785 = n130 | n21784 ;
  assign n21786 = n2732 | n21785 ;
  assign n21787 = n240 | n21786 ;
  assign n21788 = n356 | n21787 ;
  assign n21789 = n601 | n21788 ;
  assign n21790 = n120 | n21789 ;
  assign n21791 = n21782 | n21790 ;
  assign n21792 = ( n21771 & n21772 ) | ( n21771 & ~n21791 ) | ( n21772 & ~n21791 ) ;
  assign n21793 = ( ~n21772 & n21791 ) | ( ~n21772 & n21792 ) | ( n21791 & n21792 ) ;
  assign n21794 = ( ~n21771 & n21792 ) | ( ~n21771 & n21793 ) | ( n21792 & n21793 ) ;
  assign n21795 = n21764 & n21794 ;
  assign n21796 = n21764 | n21794 ;
  assign n21797 = ~n21795 & n21796 ;
  assign n21798 = n21498 | n21503 ;
  assign n21799 = n21797 | n21798 ;
  assign n21800 = n21797 & n21798 ;
  assign n21801 = n21799 & ~n21800 ;
  assign n21802 = n4484 & n20611 ;
  assign n21803 = n4479 & n20616 ;
  assign n21804 = n4481 & n20614 ;
  assign n21805 = n21803 | n21804 ;
  assign n21806 = n21802 | n21805 ;
  assign n21807 = n4487 | n21806 ;
  assign n21808 = ( n21293 & n21806 ) | ( n21293 & n21807 ) | ( n21806 & n21807 ) ;
  assign n21809 = x26 & n21808 ;
  assign n21810 = x26 & ~n21809 ;
  assign n21811 = ( n21808 & ~n21809 ) | ( n21808 & n21810 ) | ( ~n21809 & n21810 ) ;
  assign n21812 = n21801 & n21811 ;
  assign n21813 = n21811 & ~n21812 ;
  assign n21814 = ( n21801 & ~n21812 ) | ( n21801 & n21813 ) | ( ~n21812 & n21813 ) ;
  assign n21815 = n21754 & n21814 ;
  assign n21816 = n21754 & ~n21815 ;
  assign n21817 = n21814 & ~n21815 ;
  assign n21818 = n21816 | n21817 ;
  assign n21819 = n4551 & ~n20595 ;
  assign n21820 = n4546 & ~n20605 ;
  assign n21821 = n4548 & n20600 ;
  assign n21822 = n21820 | n21821 ;
  assign n21823 = n21819 | n21822 ;
  assign n21824 = n4554 | n21823 ;
  assign n21825 = ( ~n21554 & n21823 ) | ( ~n21554 & n21824 ) | ( n21823 & n21824 ) ;
  assign n21826 = ~x23 & n21825 ;
  assign n21827 = x23 | n21826 ;
  assign n21828 = ( ~n21825 & n21826 ) | ( ~n21825 & n21827 ) | ( n21826 & n21827 ) ;
  assign n21829 = n21818 & n21828 ;
  assign n21830 = n21818 & ~n21829 ;
  assign n21831 = ~n21818 & n21828 ;
  assign n21832 = n21830 | n21831 ;
  assign n21833 = n21512 | n21515 ;
  assign n21834 = n21832 | n21833 ;
  assign n21835 = n21832 & n21833 ;
  assign n21836 = n21834 & ~n21835 ;
  assign n21837 = n20589 | n20677 ;
  assign n21838 = n20676 | n21837 ;
  assign n21839 = n20676 & n21837 ;
  assign n21840 = n21838 & ~n21839 ;
  assign n21841 = n4781 & ~n20580 ;
  assign n21842 = n4776 & ~n20591 ;
  assign n21843 = n4778 & n20588 ;
  assign n21844 = n21842 | n21843 ;
  assign n21845 = n21841 | n21844 ;
  assign n21846 = n4784 | n21845 ;
  assign n21847 = ( n21840 & n21845 ) | ( n21840 & n21846 ) | ( n21845 & n21846 ) ;
  assign n21848 = x20 & n21847 ;
  assign n21849 = x20 & ~n21848 ;
  assign n21850 = ( n21847 & ~n21848 ) | ( n21847 & n21849 ) | ( ~n21848 & n21849 ) ;
  assign n21851 = n21836 & n21850 ;
  assign n21852 = n21836 & ~n21851 ;
  assign n21853 = ~n21836 & n21850 ;
  assign n21854 = n21852 | n21853 ;
  assign n21855 = n21753 & n21854 ;
  assign n21856 = n21753 & ~n21855 ;
  assign n21857 = n21854 & ~n21855 ;
  assign n21858 = n21856 | n21857 ;
  assign n21859 = ~n20576 & n20683 ;
  assign n21860 = n20684 | n21859 ;
  assign n21861 = n5083 & ~n20573 ;
  assign n21862 = n5069 & ~n20584 ;
  assign n21863 = n5070 & ~n20569 ;
  assign n21864 = n21862 | n21863 ;
  assign n21865 = n21861 | n21864 ;
  assign n21866 = n5074 | n21865 ;
  assign n21867 = ( ~n21860 & n21865 ) | ( ~n21860 & n21866 ) | ( n21865 & n21866 ) ;
  assign n21868 = ~x17 & n21867 ;
  assign n21869 = x17 | n21868 ;
  assign n21870 = ( ~n21867 & n21868 ) | ( ~n21867 & n21869 ) | ( n21868 & n21869 ) ;
  assign n21871 = n21858 & n21870 ;
  assign n21872 = n21858 & ~n21871 ;
  assign n21873 = ~n21858 & n21870 ;
  assign n21874 = n21872 | n21873 ;
  assign n21875 = n21749 & ~n21752 ;
  assign n21876 = n21751 | n21752 ;
  assign n21877 = ~n21875 & n21876 ;
  assign n21878 = n5083 & ~n20569 ;
  assign n21879 = n5069 & ~n20580 ;
  assign n21880 = n5070 & ~n20584 ;
  assign n21881 = n21879 | n21880 ;
  assign n21882 = n21878 | n21881 ;
  assign n21883 = ~n20681 & n20682 ;
  assign n21884 = ~n20680 & n21883 ;
  assign n21885 = n5074 & n21884 ;
  assign n21886 = n20569 | n20584 ;
  assign n21887 = ~n20681 & n21886 ;
  assign n21888 = n20585 & ~n20680 ;
  assign n21889 = n21887 | n21888 ;
  assign n21890 = ( n5074 & n21885 ) | ( n5074 & ~n21889 ) | ( n21885 & ~n21889 ) ;
  assign n21891 = n21882 | n21890 ;
  assign n21892 = x17 | n21891 ;
  assign n21893 = ~x17 & n21892 ;
  assign n21894 = ( ~n21891 & n21892 ) | ( ~n21891 & n21893 ) | ( n21892 & n21893 ) ;
  assign n21895 = ~n21877 & n21894 ;
  assign n21896 = n21745 & ~n21748 ;
  assign n21897 = n21747 | n21748 ;
  assign n21898 = ~n21896 & n21897 ;
  assign n21899 = ( ~n20589 & n20680 ) | ( ~n20589 & n21838 ) | ( n20680 & n21838 ) ;
  assign n21900 = ( n20580 & n20584 ) | ( n20580 & n20680 ) | ( n20584 & n20680 ) ;
  assign n21901 = ( ~n20585 & n21899 ) | ( ~n20585 & n21900 ) | ( n21899 & n21900 ) ;
  assign n21902 = n5083 & ~n20584 ;
  assign n21903 = n5069 & n20588 ;
  assign n21904 = n5070 & ~n20580 ;
  assign n21905 = n21903 | n21904 ;
  assign n21906 = n21902 | n21905 ;
  assign n21907 = n5074 | n21906 ;
  assign n21908 = ( ~n21901 & n21906 ) | ( ~n21901 & n21907 ) | ( n21906 & n21907 ) ;
  assign n21909 = ~x17 & n21908 ;
  assign n21910 = x17 | n21909 ;
  assign n21911 = ( ~n21908 & n21909 ) | ( ~n21908 & n21910 ) | ( n21909 & n21910 ) ;
  assign n21912 = ~n21898 & n21911 ;
  assign n21913 = n21898 | n21912 ;
  assign n21914 = n21898 & n21911 ;
  assign n21915 = n21567 | n21743 ;
  assign n21916 = ~n21744 & n21915 ;
  assign n21917 = n5083 & ~n20580 ;
  assign n21918 = n5069 & ~n20591 ;
  assign n21919 = n5070 & n20588 ;
  assign n21920 = n21918 | n21919 ;
  assign n21921 = n21917 | n21920 ;
  assign n21922 = n5074 | n21921 ;
  assign n21923 = ( n21840 & n21921 ) | ( n21840 & n21922 ) | ( n21921 & n21922 ) ;
  assign n21924 = x17 & n21923 ;
  assign n21925 = x17 & ~n21924 ;
  assign n21926 = ( n21923 & ~n21924 ) | ( n21923 & n21925 ) | ( ~n21924 & n21925 ) ;
  assign n21927 = n21916 & n21926 ;
  assign n21928 = n21916 | n21926 ;
  assign n21929 = ~n21927 & n21928 ;
  assign n21930 = n21584 | n21741 ;
  assign n21931 = ~n21742 & n21930 ;
  assign n21932 = n5083 & n20588 ;
  assign n21933 = n5069 & ~n20595 ;
  assign n21934 = n5070 & ~n20591 ;
  assign n21935 = n21933 | n21934 ;
  assign n21936 = n21932 | n21935 ;
  assign n21937 = n5074 | n21936 ;
  assign n21938 = ( n21526 & n21936 ) | ( n21526 & n21937 ) | ( n21936 & n21937 ) ;
  assign n21939 = x17 & n21938 ;
  assign n21940 = x17 & ~n21939 ;
  assign n21941 = ( n21938 & ~n21939 ) | ( n21938 & n21940 ) | ( ~n21939 & n21940 ) ;
  assign n21942 = n21610 | n21739 ;
  assign n21943 = n21737 | n21942 ;
  assign n21944 = ~n21740 & n21943 ;
  assign n21945 = n5083 & ~n20591 ;
  assign n21946 = n5069 & n20600 ;
  assign n21947 = n5070 & ~n20595 ;
  assign n21948 = n21946 | n21947 ;
  assign n21949 = n21945 | n21948 ;
  assign n21950 = n5074 & n21539 ;
  assign n21951 = ( n5074 & n21543 ) | ( n5074 & n21950 ) | ( n21543 & n21950 ) ;
  assign n21952 = n21949 | n21951 ;
  assign n21953 = x17 | n21952 ;
  assign n21954 = ~x17 & n21953 ;
  assign n21955 = ( ~n21952 & n21953 ) | ( ~n21952 & n21954 ) | ( n21953 & n21954 ) ;
  assign n21956 = n21944 & n21955 ;
  assign n21957 = n21734 & ~n21737 ;
  assign n21958 = n21736 & ~n21737 ;
  assign n21959 = n21957 | n21958 ;
  assign n21960 = n5083 & ~n20595 ;
  assign n21961 = n5069 & ~n20605 ;
  assign n21962 = n5070 & n20600 ;
  assign n21963 = n21961 | n21962 ;
  assign n21964 = n21960 | n21963 ;
  assign n21965 = n5074 | n21964 ;
  assign n21966 = ( ~n21554 & n21964 ) | ( ~n21554 & n21965 ) | ( n21964 & n21965 ) ;
  assign n21967 = ~x17 & n21966 ;
  assign n21968 = x17 | n21967 ;
  assign n21969 = ( ~n21966 & n21967 ) | ( ~n21966 & n21968 ) | ( n21967 & n21968 ) ;
  assign n21970 = n21959 & n21969 ;
  assign n21971 = n21959 & ~n21970 ;
  assign n21972 = ~n21959 & n21969 ;
  assign n21973 = n21971 | n21972 ;
  assign n21974 = n21729 & ~n21733 ;
  assign n21975 = n21732 & ~n21733 ;
  assign n21976 = n21974 | n21975 ;
  assign n21977 = n5083 & n20600 ;
  assign n21978 = n5069 & n20611 ;
  assign n21979 = n5070 & ~n20605 ;
  assign n21980 = n21978 | n21979 ;
  assign n21981 = n21977 | n21980 ;
  assign n21982 = n5074 | n21981 ;
  assign n21983 = ( ~n21432 & n21981 ) | ( ~n21432 & n21982 ) | ( n21981 & n21982 ) ;
  assign n21984 = ~x17 & n21983 ;
  assign n21985 = x17 | n21984 ;
  assign n21986 = ( ~n21983 & n21984 ) | ( ~n21983 & n21985 ) | ( n21984 & n21985 ) ;
  assign n21987 = n21976 & n21986 ;
  assign n21988 = n21976 & ~n21987 ;
  assign n21989 = ~n21976 & n21986 ;
  assign n21990 = n21988 | n21989 ;
  assign n21991 = n21725 | n21727 ;
  assign n21992 = ~n21728 & n21991 ;
  assign n21993 = n5083 & ~n20605 ;
  assign n21994 = n5069 & n20614 ;
  assign n21995 = n5070 & n20611 ;
  assign n21996 = n21994 | n21995 ;
  assign n21997 = n21993 | n21996 ;
  assign n21998 = n5074 | n21997 ;
  assign n21999 = ( ~n21275 & n21997 ) | ( ~n21275 & n21998 ) | ( n21997 & n21998 ) ;
  assign n22000 = ~x17 & n21999 ;
  assign n22001 = x17 | n22000 ;
  assign n22002 = ( ~n21999 & n22000 ) | ( ~n21999 & n22001 ) | ( n22000 & n22001 ) ;
  assign n22003 = n21992 & n22002 ;
  assign n22004 = n21651 | n21723 ;
  assign n22005 = ~n21724 & n22004 ;
  assign n22006 = n5083 & n20611 ;
  assign n22007 = n5069 & n20616 ;
  assign n22008 = n5070 & n20614 ;
  assign n22009 = n22007 | n22008 ;
  assign n22010 = n22006 | n22009 ;
  assign n22011 = n5074 | n22010 ;
  assign n22012 = ( n21293 & n22010 ) | ( n21293 & n22011 ) | ( n22010 & n22011 ) ;
  assign n22013 = x17 & n22012 ;
  assign n22014 = x17 & ~n22013 ;
  assign n22015 = ( n22012 & ~n22013 ) | ( n22012 & n22014 ) | ( ~n22013 & n22014 ) ;
  assign n22016 = n22005 & n22015 ;
  assign n22017 = n21719 | n21721 ;
  assign n22018 = ~n21722 & n22017 ;
  assign n22019 = n5083 & n20614 ;
  assign n22020 = n5069 & n20619 ;
  assign n22021 = n5070 | n22020 ;
  assign n22022 = ( n20616 & n22020 ) | ( n20616 & n22021 ) | ( n22020 & n22021 ) ;
  assign n22023 = n22019 | n22022 ;
  assign n22024 = n5074 | n22023 ;
  assign n22025 = ( n21302 & n22023 ) | ( n21302 & n22024 ) | ( n22023 & n22024 ) ;
  assign n22026 = x17 & n22025 ;
  assign n22027 = x17 & ~n22026 ;
  assign n22028 = ( n22025 & ~n22026 ) | ( n22025 & n22027 ) | ( ~n22026 & n22027 ) ;
  assign n22029 = n22018 & n22028 ;
  assign n22030 = n5069 & n20622 ;
  assign n22031 = n5070 | n22030 ;
  assign n22032 = ( n20619 & n22030 ) | ( n20619 & n22031 ) | ( n22030 & n22031 ) ;
  assign n22033 = n5083 | n22032 ;
  assign n22034 = ( n20616 & n22032 ) | ( n20616 & n22033 ) | ( n22032 & n22033 ) ;
  assign n22035 = n5074 | n22034 ;
  assign n22036 = ( n21190 & n22034 ) | ( n21190 & n22035 ) | ( n22034 & n22035 ) ;
  assign n22037 = ~x17 & n22036 ;
  assign n22038 = x17 & ~n22036 ;
  assign n22039 = n22037 | n22038 ;
  assign n22040 = n21679 | n21717 ;
  assign n22041 = ~n21718 & n22040 ;
  assign n22042 = n22039 & n22041 ;
  assign n22043 = n5069 & ~n20625 ;
  assign n22044 = n5070 | n22043 ;
  assign n22045 = ( n20622 & n22043 ) | ( n20622 & n22044 ) | ( n22043 & n22044 ) ;
  assign n22046 = n5083 | n22045 ;
  assign n22047 = ( n20619 & n22045 ) | ( n20619 & n22046 ) | ( n22045 & n22046 ) ;
  assign n22048 = n5074 | n22047 ;
  assign n22049 = ( ~n21056 & n22047 ) | ( ~n21056 & n22048 ) | ( n22047 & n22048 ) ;
  assign n22050 = ~x17 & n22049 ;
  assign n22051 = x17 | n22050 ;
  assign n22052 = ( ~n22049 & n22050 ) | ( ~n22049 & n22051 ) | ( n22050 & n22051 ) ;
  assign n22053 = n21705 & ~n21716 ;
  assign n22054 = ( n21715 & ~n21716 ) | ( n21715 & n22053 ) | ( ~n21716 & n22053 ) ;
  assign n22055 = n22052 & n22054 ;
  assign n22056 = n22052 | n22054 ;
  assign n22057 = ~n22055 & n22056 ;
  assign n22058 = n21689 | n21700 ;
  assign n22059 = ~n21703 & n22058 ;
  assign n22060 = n5083 & n20622 ;
  assign n22061 = n5069 & ~n20630 ;
  assign n22062 = n5070 & ~n20625 ;
  assign n22063 = n22061 | n22062 ;
  assign n22064 = n22060 | n22063 ;
  assign n22065 = n5074 | n22064 ;
  assign n22066 = ( n21114 & n22064 ) | ( n21114 & n22065 ) | ( n22064 & n22065 ) ;
  assign n22067 = x17 & n22066 ;
  assign n22068 = x17 | n22066 ;
  assign n22069 = ~n22067 & n22068 ;
  assign n22070 = n22059 & n22069 ;
  assign n22071 = n21680 | n21688 ;
  assign n22072 = ~n21689 & n22071 ;
  assign n22073 = n5083 & ~n20625 ;
  assign n22074 = n5069 & n20633 ;
  assign n22075 = n5070 & ~n20630 ;
  assign n22076 = n22074 | n22075 ;
  assign n22077 = n22073 | n22076 ;
  assign n22078 = n5074 | n22077 ;
  assign n22079 = ( ~n21129 & n22077 ) | ( ~n21129 & n22078 ) | ( n22077 & n22078 ) ;
  assign n22080 = ~x17 & n22079 ;
  assign n22081 = x17 | n22080 ;
  assign n22082 = ( ~n22079 & n22080 ) | ( ~n22079 & n22081 ) | ( n22080 & n22081 ) ;
  assign n22083 = n22072 & n22082 ;
  assign n22084 = n22072 | n22082 ;
  assign n22085 = ~n22083 & n22084 ;
  assign n22086 = ( x17 & n15890 ) | ( x17 & n20642 ) | ( n15890 & n20642 ) ;
  assign n22087 = n5074 & n21069 ;
  assign n22088 = n5070 & ~n20642 ;
  assign n22089 = n5083 & ~n20640 ;
  assign n22090 = n22088 | n22089 ;
  assign n22091 = n22087 | n22090 ;
  assign n22092 = x17 | n22091 ;
  assign n22093 = ~x17 & n22092 ;
  assign n22094 = ( ~n22091 & n22092 ) | ( ~n22091 & n22093 ) | ( n22092 & n22093 ) ;
  assign n22095 = n22086 & n22094 ;
  assign n22096 = n4774 & ~n20642 ;
  assign n22097 = n5083 & n20633 ;
  assign n22098 = n5069 & ~n20642 ;
  assign n22099 = n5070 & ~n20640 ;
  assign n22100 = n22098 | n22099 ;
  assign n22101 = n22097 | n22100 ;
  assign n22102 = n5074 & n21085 ;
  assign n22103 = n22101 | n22102 ;
  assign n22104 = ~x17 & n22103 ;
  assign n22105 = x17 | n22104 ;
  assign n22106 = ( ~n22103 & n22104 ) | ( ~n22103 & n22105 ) | ( n22104 & n22105 ) ;
  assign n22107 = n22096 & n22106 ;
  assign n22108 = n22095 & n22107 ;
  assign n22109 = n22095 & n22106 ;
  assign n22110 = n22096 | n22109 ;
  assign n22111 = ~n22108 & n22110 ;
  assign n22112 = n5083 & ~n20630 ;
  assign n22113 = n5069 & ~n20640 ;
  assign n22114 = n5070 & n20633 ;
  assign n22115 = n22113 | n22114 ;
  assign n22116 = n22112 | n22115 ;
  assign n22117 = n5074 | n22116 ;
  assign n22118 = ( n21099 & n22116 ) | ( n21099 & n22117 ) | ( n22116 & n22117 ) ;
  assign n22119 = x17 & n22118 ;
  assign n22120 = x17 | n22118 ;
  assign n22121 = ~n22119 & n22120 ;
  assign n22122 = n22111 & n22121 ;
  assign n22123 = n22108 | n22122 ;
  assign n22124 = n22085 & n22123 ;
  assign n22125 = n22083 | n22124 ;
  assign n22126 = n22069 & ~n22070 ;
  assign n22127 = ( n22059 & ~n22070 ) | ( n22059 & n22126 ) | ( ~n22070 & n22126 ) ;
  assign n22128 = n22125 & n22127 ;
  assign n22129 = n22070 | n22128 ;
  assign n22130 = n22057 & n22129 ;
  assign n22131 = n22055 | n22130 ;
  assign n22132 = n22039 | n22041 ;
  assign n22133 = ~n22042 & n22132 ;
  assign n22134 = n22131 & n22133 ;
  assign n22135 = n22042 | n22134 ;
  assign n22136 = n22018 & ~n22029 ;
  assign n22137 = n22028 & ~n22029 ;
  assign n22138 = n22136 | n22137 ;
  assign n22139 = n22135 & n22138 ;
  assign n22140 = n22029 | n22139 ;
  assign n22141 = n22015 & ~n22016 ;
  assign n22142 = ( n22005 & ~n22016 ) | ( n22005 & n22141 ) | ( ~n22016 & n22141 ) ;
  assign n22143 = n22140 & n22142 ;
  assign n22144 = n21992 | n22002 ;
  assign n22145 = ~n22003 & n22144 ;
  assign n22146 = ( n22016 & n22143 ) | ( n22016 & n22145 ) | ( n22143 & n22145 ) ;
  assign n22147 = n22003 | n22146 ;
  assign n22148 = n21990 & n22147 ;
  assign n22149 = n21987 | n22148 ;
  assign n22150 = n21973 & n22149 ;
  assign n22151 = n21970 | n22150 ;
  assign n22152 = n21955 & ~n21956 ;
  assign n22153 = ( n21944 & ~n21956 ) | ( n21944 & n22152 ) | ( ~n21956 & n22152 ) ;
  assign n22154 = n22151 & n22153 ;
  assign n22155 = n21956 | n22154 ;
  assign n22156 = ( n21931 & n21941 ) | ( n21931 & n22155 ) | ( n21941 & n22155 ) ;
  assign n22157 = n21929 & n22156 ;
  assign n22158 = n21927 | n22157 ;
  assign n22159 = ( ~n21913 & n21914 ) | ( ~n21913 & n22158 ) | ( n21914 & n22158 ) ;
  assign n22160 = n21912 | n22159 ;
  assign n22161 = n21877 | n21895 ;
  assign n22162 = ( ~n21894 & n21895 ) | ( ~n21894 & n22161 ) | ( n21895 & n22161 ) ;
  assign n22163 = n22160 & ~n22162 ;
  assign n22164 = n21895 | n22163 ;
  assign n22165 = n21874 & n22164 ;
  assign n22166 = n21874 | n22164 ;
  assign n22167 = ~n22165 & n22166 ;
  assign n22168 = n7280 & n20560 ;
  assign n22169 = n5384 & ~n20573 ;
  assign n22170 = n7277 & ~n20689 ;
  assign n22171 = n22169 | n22170 ;
  assign n22172 = n22168 | n22171 ;
  assign n22173 = ~n20691 & n20696 ;
  assign n22174 = ( n20560 & n20685 ) | ( n20560 & n20689 ) | ( n20685 & n20689 ) ;
  assign n22175 = ( n20560 & ~n20573 ) | ( n20560 & n20689 ) | ( ~n20573 & n20689 ) ;
  assign n22176 = ( n20693 & ~n22174 ) | ( n20693 & n22175 ) | ( ~n22174 & n22175 ) ;
  assign n22177 = n39 & ~n22176 ;
  assign n22178 = ~n22173 & n22177 ;
  assign n22179 = ( n39 & n22172 ) | ( n39 & ~n22178 ) | ( n22172 & ~n22178 ) ;
  assign n22180 = ~x14 & n22179 ;
  assign n22181 = x14 | n22180 ;
  assign n22182 = ( ~n22179 & n22180 ) | ( ~n22179 & n22181 ) | ( n22180 & n22181 ) ;
  assign n22183 = n21914 | n22158 ;
  assign n22184 = n21913 & ~n22183 ;
  assign n22185 = n22159 | n22184 ;
  assign n22186 = n7280 & ~n20689 ;
  assign n22187 = n5384 & ~n20569 ;
  assign n22188 = n7277 & ~n20573 ;
  assign n22189 = n22187 | n22188 ;
  assign n22190 = n22186 | n22189 ;
  assign n22191 = ~n20690 & n20694 ;
  assign n22192 = n20685 | n22191 ;
  assign n22193 = n20685 & n22191 ;
  assign n22194 = n39 & ~n22193 ;
  assign n22195 = n22192 & n22194 ;
  assign n22196 = ( n39 & n22190 ) | ( n39 & ~n22195 ) | ( n22190 & ~n22195 ) ;
  assign n22197 = x14 & n22196 ;
  assign n22198 = x14 & ~n22197 ;
  assign n22199 = ( n22196 & ~n22197 ) | ( n22196 & n22198 ) | ( ~n22197 & n22198 ) ;
  assign n22200 = ~n22185 & n22199 ;
  assign n22201 = n21929 | n22156 ;
  assign n22202 = ~n22157 & n22201 ;
  assign n22203 = n7280 & ~n20573 ;
  assign n22204 = n5384 & ~n20584 ;
  assign n22205 = n7277 & ~n20569 ;
  assign n22206 = n22204 | n22205 ;
  assign n22207 = n22203 | n22206 ;
  assign n22208 = n39 | n22207 ;
  assign n22209 = ( ~n21860 & n22207 ) | ( ~n21860 & n22208 ) | ( n22207 & n22208 ) ;
  assign n22210 = ~x14 & n22209 ;
  assign n22211 = x14 | n22210 ;
  assign n22212 = ( ~n22209 & n22210 ) | ( ~n22209 & n22211 ) | ( n22210 & n22211 ) ;
  assign n22213 = n22202 & n22212 ;
  assign n22214 = n22212 & ~n22213 ;
  assign n22215 = ( n22202 & ~n22213 ) | ( n22202 & n22214 ) | ( ~n22213 & n22214 ) ;
  assign n22216 = n7280 & ~n20569 ;
  assign n22217 = n5384 & ~n20580 ;
  assign n22218 = n7277 & ~n20584 ;
  assign n22219 = n22217 | n22218 ;
  assign n22220 = n22216 | n22219 ;
  assign n22221 = n39 & n21884 ;
  assign n22222 = ( n39 & ~n21889 ) | ( n39 & n22221 ) | ( ~n21889 & n22221 ) ;
  assign n22223 = n22220 | n22222 ;
  assign n22224 = x14 | n22223 ;
  assign n22225 = ~x14 & n22224 ;
  assign n22226 = ( ~n22223 & n22224 ) | ( ~n22223 & n22225 ) | ( n22224 & n22225 ) ;
  assign n22227 = ( n21931 & n22155 ) | ( n21931 & ~n22156 ) | ( n22155 & ~n22156 ) ;
  assign n22228 = ( n21941 & ~n22156 ) | ( n21941 & n22227 ) | ( ~n22156 & n22227 ) ;
  assign n22229 = n22226 & n22228 ;
  assign n22230 = n22226 | n22228 ;
  assign n22231 = ~n22229 & n22230 ;
  assign n22232 = n22151 | n22153 ;
  assign n22233 = ~n22154 & n22232 ;
  assign n22234 = n7280 & ~n20584 ;
  assign n22235 = n5384 & n20588 ;
  assign n22236 = n7277 & ~n20580 ;
  assign n22237 = n22235 | n22236 ;
  assign n22238 = n22234 | n22237 ;
  assign n22239 = n39 | n22238 ;
  assign n22240 = ( ~n21901 & n22238 ) | ( ~n21901 & n22239 ) | ( n22238 & n22239 ) ;
  assign n22241 = ~x14 & n22240 ;
  assign n22242 = x14 | n22241 ;
  assign n22243 = ( ~n22240 & n22241 ) | ( ~n22240 & n22242 ) | ( n22241 & n22242 ) ;
  assign n22244 = n22233 & n22243 ;
  assign n22245 = n22233 | n22243 ;
  assign n22246 = ~n22244 & n22245 ;
  assign n22247 = n21973 | n22149 ;
  assign n22248 = ~n22150 & n22247 ;
  assign n22249 = n7280 & ~n20580 ;
  assign n22250 = n5384 & ~n20591 ;
  assign n22251 = n7277 & n20588 ;
  assign n22252 = n22250 | n22251 ;
  assign n22253 = n22249 | n22252 ;
  assign n22254 = n39 | n22253 ;
  assign n22255 = ( n21840 & n22253 ) | ( n21840 & n22254 ) | ( n22253 & n22254 ) ;
  assign n22256 = x14 & n22255 ;
  assign n22257 = x14 & ~n22256 ;
  assign n22258 = ( n22255 & ~n22256 ) | ( n22255 & n22257 ) | ( ~n22256 & n22257 ) ;
  assign n22259 = n21990 | n22147 ;
  assign n22260 = ~n22148 & n22259 ;
  assign n22261 = n7280 & n20588 ;
  assign n22262 = n5384 & ~n20595 ;
  assign n22263 = n7277 & ~n20591 ;
  assign n22264 = n22262 | n22263 ;
  assign n22265 = n22261 | n22264 ;
  assign n22266 = n39 | n22265 ;
  assign n22267 = ( n21526 & n22265 ) | ( n21526 & n22266 ) | ( n22265 & n22266 ) ;
  assign n22268 = x14 & n22267 ;
  assign n22269 = x14 & ~n22268 ;
  assign n22270 = ( n22267 & ~n22268 ) | ( n22267 & n22269 ) | ( ~n22268 & n22269 ) ;
  assign n22271 = n22016 | n22145 ;
  assign n22272 = n22143 | n22271 ;
  assign n22273 = ~n22146 & n22272 ;
  assign n22274 = n7280 & ~n20591 ;
  assign n22275 = n5384 & n20600 ;
  assign n22276 = n7277 & ~n20595 ;
  assign n22277 = n22275 | n22276 ;
  assign n22278 = n22274 | n22277 ;
  assign n22279 = n39 & n21539 ;
  assign n22280 = ( n39 & n21543 ) | ( n39 & n22279 ) | ( n21543 & n22279 ) ;
  assign n22281 = n22278 | n22280 ;
  assign n22282 = x14 | n22281 ;
  assign n22283 = ~x14 & n22282 ;
  assign n22284 = ( ~n22281 & n22282 ) | ( ~n22281 & n22283 ) | ( n22282 & n22283 ) ;
  assign n22285 = n22273 & n22284 ;
  assign n22286 = n22140 & ~n22143 ;
  assign n22287 = n22142 & ~n22143 ;
  assign n22288 = n22286 | n22287 ;
  assign n22289 = n7280 & ~n20595 ;
  assign n22290 = n5384 & ~n20605 ;
  assign n22291 = n7277 & n20600 ;
  assign n22292 = n22290 | n22291 ;
  assign n22293 = n22289 | n22292 ;
  assign n22294 = n39 | n22293 ;
  assign n22295 = ( ~n21554 & n22293 ) | ( ~n21554 & n22294 ) | ( n22293 & n22294 ) ;
  assign n22296 = ~x14 & n22295 ;
  assign n22297 = x14 | n22296 ;
  assign n22298 = ( ~n22295 & n22296 ) | ( ~n22295 & n22297 ) | ( n22296 & n22297 ) ;
  assign n22299 = n22288 & n22298 ;
  assign n22300 = n22288 & ~n22299 ;
  assign n22301 = ~n22288 & n22298 ;
  assign n22302 = n22300 | n22301 ;
  assign n22303 = n22135 & ~n22139 ;
  assign n22304 = n22138 & ~n22139 ;
  assign n22305 = n22303 | n22304 ;
  assign n22306 = n7280 & n20600 ;
  assign n22307 = n5384 & n20611 ;
  assign n22308 = n7277 & ~n20605 ;
  assign n22309 = n22307 | n22308 ;
  assign n22310 = n22306 | n22309 ;
  assign n22311 = n39 | n22310 ;
  assign n22312 = ( ~n21432 & n22310 ) | ( ~n21432 & n22311 ) | ( n22310 & n22311 ) ;
  assign n22313 = ~x14 & n22312 ;
  assign n22314 = x14 | n22313 ;
  assign n22315 = ( ~n22312 & n22313 ) | ( ~n22312 & n22314 ) | ( n22313 & n22314 ) ;
  assign n22316 = n22305 & n22315 ;
  assign n22317 = n22305 & ~n22316 ;
  assign n22318 = ~n22305 & n22315 ;
  assign n22319 = n22317 | n22318 ;
  assign n22320 = n22131 | n22133 ;
  assign n22321 = ~n22134 & n22320 ;
  assign n22322 = n7280 & ~n20605 ;
  assign n22323 = n5384 & n20614 ;
  assign n22324 = n7277 & n20611 ;
  assign n22325 = n22323 | n22324 ;
  assign n22326 = n22322 | n22325 ;
  assign n22327 = n39 | n22326 ;
  assign n22328 = ( ~n21275 & n22326 ) | ( ~n21275 & n22327 ) | ( n22326 & n22327 ) ;
  assign n22329 = ~x14 & n22328 ;
  assign n22330 = x14 | n22329 ;
  assign n22331 = ( ~n22328 & n22329 ) | ( ~n22328 & n22330 ) | ( n22329 & n22330 ) ;
  assign n22332 = n22321 & n22331 ;
  assign n22333 = n22057 | n22129 ;
  assign n22334 = ~n22130 & n22333 ;
  assign n22335 = n7280 & n20611 ;
  assign n22336 = n5384 & n20616 ;
  assign n22337 = n7277 & n20614 ;
  assign n22338 = n22336 | n22337 ;
  assign n22339 = n22335 | n22338 ;
  assign n22340 = n39 | n22339 ;
  assign n22341 = ( n21293 & n22339 ) | ( n21293 & n22340 ) | ( n22339 & n22340 ) ;
  assign n22342 = x14 & n22341 ;
  assign n22343 = x14 & ~n22342 ;
  assign n22344 = ( n22341 & ~n22342 ) | ( n22341 & n22343 ) | ( ~n22342 & n22343 ) ;
  assign n22345 = n22334 & n22344 ;
  assign n22346 = n22125 | n22127 ;
  assign n22347 = ~n22128 & n22346 ;
  assign n22348 = n7280 & n20614 ;
  assign n22349 = n5384 & n20619 ;
  assign n22350 = n7277 | n22349 ;
  assign n22351 = ( n20616 & n22349 ) | ( n20616 & n22350 ) | ( n22349 & n22350 ) ;
  assign n22352 = n22348 | n22351 ;
  assign n22353 = n39 | n22352 ;
  assign n22354 = ( n21302 & n22352 ) | ( n21302 & n22353 ) | ( n22352 & n22353 ) ;
  assign n22355 = x14 & n22354 ;
  assign n22356 = x14 & ~n22355 ;
  assign n22357 = ( n22354 & ~n22355 ) | ( n22354 & n22356 ) | ( ~n22355 & n22356 ) ;
  assign n22358 = n22347 & n22357 ;
  assign n22359 = n5384 & n20622 ;
  assign n22360 = n7277 | n22359 ;
  assign n22361 = ( n20619 & n22359 ) | ( n20619 & n22360 ) | ( n22359 & n22360 ) ;
  assign n22362 = n7280 | n22361 ;
  assign n22363 = ( n20616 & n22361 ) | ( n20616 & n22362 ) | ( n22361 & n22362 ) ;
  assign n22364 = n39 | n22363 ;
  assign n22365 = ( n21190 & n22363 ) | ( n21190 & n22364 ) | ( n22363 & n22364 ) ;
  assign n22366 = ~x14 & n22365 ;
  assign n22367 = x14 & ~n22365 ;
  assign n22368 = n22366 | n22367 ;
  assign n22369 = n22085 | n22123 ;
  assign n22370 = ~n22124 & n22369 ;
  assign n22371 = n22368 & n22370 ;
  assign n22372 = n5384 & ~n20625 ;
  assign n22373 = n7277 | n22372 ;
  assign n22374 = ( n20622 & n22372 ) | ( n20622 & n22373 ) | ( n22372 & n22373 ) ;
  assign n22375 = n7280 | n22374 ;
  assign n22376 = ( n20619 & n22374 ) | ( n20619 & n22375 ) | ( n22374 & n22375 ) ;
  assign n22377 = n39 | n22376 ;
  assign n22378 = ( ~n21056 & n22376 ) | ( ~n21056 & n22377 ) | ( n22376 & n22377 ) ;
  assign n22379 = ~x14 & n22378 ;
  assign n22380 = x14 | n22379 ;
  assign n22381 = ( ~n22378 & n22379 ) | ( ~n22378 & n22380 ) | ( n22379 & n22380 ) ;
  assign n22382 = n22111 & ~n22122 ;
  assign n22383 = ( n22121 & ~n22122 ) | ( n22121 & n22382 ) | ( ~n22122 & n22382 ) ;
  assign n22384 = n22381 & n22383 ;
  assign n22385 = n22381 | n22383 ;
  assign n22386 = ~n22384 & n22385 ;
  assign n22387 = n22095 | n22106 ;
  assign n22388 = ~n22109 & n22387 ;
  assign n22389 = n7280 & n20622 ;
  assign n22390 = n5384 & ~n20630 ;
  assign n22391 = n7277 & ~n20625 ;
  assign n22392 = n22390 | n22391 ;
  assign n22393 = n22389 | n22392 ;
  assign n22394 = n39 | n22393 ;
  assign n22395 = ( n21114 & n22393 ) | ( n21114 & n22394 ) | ( n22393 & n22394 ) ;
  assign n22396 = x14 & n22395 ;
  assign n22397 = x14 | n22395 ;
  assign n22398 = ~n22396 & n22397 ;
  assign n22399 = n22388 & n22398 ;
  assign n22400 = n22086 | n22094 ;
  assign n22401 = ~n22095 & n22400 ;
  assign n22402 = n7280 & ~n20625 ;
  assign n22403 = n5384 & n20633 ;
  assign n22404 = n7277 & ~n20630 ;
  assign n22405 = n22403 | n22404 ;
  assign n22406 = n22402 | n22405 ;
  assign n22407 = n39 | n22406 ;
  assign n22408 = ( ~n21129 & n22406 ) | ( ~n21129 & n22407 ) | ( n22406 & n22407 ) ;
  assign n22409 = ~x14 & n22408 ;
  assign n22410 = x14 | n22409 ;
  assign n22411 = ( ~n22408 & n22409 ) | ( ~n22408 & n22410 ) | ( n22409 & n22410 ) ;
  assign n22412 = n22401 & n22411 ;
  assign n22413 = n22401 | n22411 ;
  assign n22414 = ~n22412 & n22413 ;
  assign n22415 = ( x14 & n16692 ) | ( x14 & n20642 ) | ( n16692 & n20642 ) ;
  assign n22416 = n39 & n21069 ;
  assign n22417 = n7277 & ~n20642 ;
  assign n22418 = n7280 & ~n20640 ;
  assign n22419 = n22417 | n22418 ;
  assign n22420 = n22416 | n22419 ;
  assign n22421 = x14 | n22420 ;
  assign n22422 = ~x14 & n22421 ;
  assign n22423 = ( ~n22420 & n22421 ) | ( ~n22420 & n22422 ) | ( n22421 & n22422 ) ;
  assign n22424 = n22415 & n22423 ;
  assign n22425 = n5064 & ~n20642 ;
  assign n22426 = n7280 & n20633 ;
  assign n22427 = n5384 & ~n20642 ;
  assign n22428 = n7277 & ~n20640 ;
  assign n22429 = n22427 | n22428 ;
  assign n22430 = n22426 | n22429 ;
  assign n22431 = n39 & n21085 ;
  assign n22432 = n22430 | n22431 ;
  assign n22433 = ~x14 & n22432 ;
  assign n22434 = x14 | n22433 ;
  assign n22435 = ( ~n22432 & n22433 ) | ( ~n22432 & n22434 ) | ( n22433 & n22434 ) ;
  assign n22436 = n22425 & n22435 ;
  assign n22437 = n22424 & n22436 ;
  assign n22438 = n22424 & n22435 ;
  assign n22439 = n22425 | n22438 ;
  assign n22440 = ~n22437 & n22439 ;
  assign n22441 = n7280 & ~n20630 ;
  assign n22442 = n5384 & ~n20640 ;
  assign n22443 = n7277 & n20633 ;
  assign n22444 = n22442 | n22443 ;
  assign n22445 = n22441 | n22444 ;
  assign n22446 = n39 | n22445 ;
  assign n22447 = ( n21099 & n22445 ) | ( n21099 & n22446 ) | ( n22445 & n22446 ) ;
  assign n22448 = x14 & n22447 ;
  assign n22449 = x14 | n22447 ;
  assign n22450 = ~n22448 & n22449 ;
  assign n22451 = n22440 & n22450 ;
  assign n22452 = n22437 | n22451 ;
  assign n22453 = n22414 & n22452 ;
  assign n22454 = n22412 | n22453 ;
  assign n22455 = n22398 & ~n22399 ;
  assign n22456 = ( n22388 & ~n22399 ) | ( n22388 & n22455 ) | ( ~n22399 & n22455 ) ;
  assign n22457 = n22454 & n22456 ;
  assign n22458 = n22399 | n22457 ;
  assign n22459 = n22386 & n22458 ;
  assign n22460 = n22384 | n22459 ;
  assign n22461 = n22368 | n22370 ;
  assign n22462 = ~n22371 & n22461 ;
  assign n22463 = n22460 & n22462 ;
  assign n22464 = n22371 | n22463 ;
  assign n22465 = n22347 & ~n22358 ;
  assign n22466 = n22357 & ~n22358 ;
  assign n22467 = n22465 | n22466 ;
  assign n22468 = n22464 & n22467 ;
  assign n22469 = n22358 | n22468 ;
  assign n22470 = n22344 & ~n22345 ;
  assign n22471 = ( n22334 & ~n22345 ) | ( n22334 & n22470 ) | ( ~n22345 & n22470 ) ;
  assign n22472 = n22469 & n22471 ;
  assign n22473 = n22321 | n22331 ;
  assign n22474 = ~n22332 & n22473 ;
  assign n22475 = ( n22345 & n22472 ) | ( n22345 & n22474 ) | ( n22472 & n22474 ) ;
  assign n22476 = n22332 | n22475 ;
  assign n22477 = n22319 & n22476 ;
  assign n22478 = n22316 | n22477 ;
  assign n22479 = n22302 & n22478 ;
  assign n22480 = n22299 | n22479 ;
  assign n22481 = n22284 & ~n22285 ;
  assign n22482 = ( n22273 & ~n22285 ) | ( n22273 & n22481 ) | ( ~n22285 & n22481 ) ;
  assign n22483 = n22480 & n22482 ;
  assign n22484 = n22285 | n22483 ;
  assign n22485 = ( n22260 & n22270 ) | ( n22260 & n22484 ) | ( n22270 & n22484 ) ;
  assign n22486 = ( n22248 & n22258 ) | ( n22248 & n22485 ) | ( n22258 & n22485 ) ;
  assign n22487 = n22246 & n22486 ;
  assign n22488 = n22244 | n22487 ;
  assign n22489 = n22231 & n22488 ;
  assign n22490 = n22229 | n22489 ;
  assign n22491 = n22215 & n22490 ;
  assign n22492 = n22213 | n22491 ;
  assign n22493 = n22185 | n22200 ;
  assign n22494 = ( ~n22199 & n22200 ) | ( ~n22199 & n22493 ) | ( n22200 & n22493 ) ;
  assign n22495 = n22492 & ~n22494 ;
  assign n22496 = n22200 | n22495 ;
  assign n22497 = ~n22160 & n22162 ;
  assign n22498 = n22163 | n22497 ;
  assign n22499 = ( n22182 & ~n22496 ) | ( n22182 & n22498 ) | ( ~n22496 & n22498 ) ;
  assign n22500 = ( ~n22182 & n22496 ) | ( ~n22182 & n22499 ) | ( n22496 & n22499 ) ;
  assign n22501 = ( ~n22498 & n22499 ) | ( ~n22498 & n22500 ) | ( n22499 & n22500 ) ;
  assign n22502 = ( n22182 & n22496 ) | ( n22182 & n22501 ) | ( n22496 & n22501 ) ;
  assign n22503 = ( n21054 & n22167 ) | ( n21054 & n22502 ) | ( n22167 & n22502 ) ;
  assign n22647 = ( n22167 & n22502 ) | ( n22167 & ~n22503 ) | ( n22502 & ~n22503 ) ;
  assign n22648 = ( n21054 & ~n22503 ) | ( n21054 & n22647 ) | ( ~n22503 & n22647 ) ;
  assign n22649 = n22646 & n22648 ;
  assign n22650 = n22646 | n22648 ;
  assign n22651 = ~n22649 & n22650 ;
  assign n22652 = ( n20697 & n20699 ) | ( n20697 & ~n20702 ) | ( n20699 & ~n20702 ) ;
  assign n22653 = ~n20705 & n22652 ;
  assign n22654 = n20700 | n20706 ;
  assign n22655 = ~n22653 & n22654 ;
  assign n22656 = n7305 & n20556 ;
  assign n22657 = n7300 & n20562 ;
  assign n22658 = n7302 & ~n20552 ;
  assign n22659 = n22657 | n22658 ;
  assign n22660 = n22656 | n22659 ;
  assign n22661 = n7308 | n22660 ;
  assign n22662 = ( ~n22655 & n22660 ) | ( ~n22655 & n22661 ) | ( n22660 & n22661 ) ;
  assign n22663 = ~x11 & n22662 ;
  assign n22664 = x11 | n22663 ;
  assign n22665 = ( ~n22662 & n22663 ) | ( ~n22662 & n22664 ) | ( n22663 & n22664 ) ;
  assign n22666 = ~n22501 & n22665 ;
  assign n22667 = n22501 & ~n22665 ;
  assign n22668 = n22666 | n22667 ;
  assign n22669 = n22492 & ~n22495 ;
  assign n22670 = n22494 | n22495 ;
  assign n22671 = ~n22669 & n22670 ;
  assign n22672 = n7305 & ~n20552 ;
  assign n22673 = n7300 & n20560 ;
  assign n22674 = n7302 & n20562 ;
  assign n22675 = n22673 | n22674 ;
  assign n22676 = n22672 | n22675 ;
  assign n22511 = n20698 | n20702 ;
  assign n22512 = ( n20563 & n20697 ) | ( n20563 & n22511 ) | ( n20697 & n22511 ) ;
  assign n22509 = n20699 | n20702 ;
  assign n22510 = n20697 | n22509 ;
  assign n22677 = n7308 & ~n22510 ;
  assign n22678 = ( n7308 & n22512 ) | ( n7308 & n22677 ) | ( n22512 & n22677 ) ;
  assign n22679 = n22676 | n22678 ;
  assign n22680 = x11 | n22679 ;
  assign n22681 = ~x11 & n22680 ;
  assign n22682 = ( ~n22679 & n22680 ) | ( ~n22679 & n22681 ) | ( n22680 & n22681 ) ;
  assign n22683 = ~n22671 & n22682 ;
  assign n22684 = n22215 | n22490 ;
  assign n22685 = ~n22491 & n22684 ;
  assign n22686 = n7305 & n20562 ;
  assign n22687 = n7300 & ~n20689 ;
  assign n22688 = n7302 & n20560 ;
  assign n22689 = n22687 | n22688 ;
  assign n22690 = n22686 | n22689 ;
  assign n22691 = n7308 | n22690 ;
  assign n22692 = ( ~n21044 & n22690 ) | ( ~n21044 & n22691 ) | ( n22690 & n22691 ) ;
  assign n22693 = ~x11 & n22692 ;
  assign n22694 = x11 | n22693 ;
  assign n22695 = ( ~n22692 & n22693 ) | ( ~n22692 & n22694 ) | ( n22693 & n22694 ) ;
  assign n22696 = n22685 & n22695 ;
  assign n22697 = n22231 | n22488 ;
  assign n22698 = ~n22489 & n22697 ;
  assign n22699 = n7305 & n20560 ;
  assign n22700 = n7300 & ~n20573 ;
  assign n22701 = n7302 & ~n20689 ;
  assign n22702 = n22700 | n22701 ;
  assign n22703 = n22699 | n22702 ;
  assign n22704 = n7308 & ~n22176 ;
  assign n22705 = ~n22173 & n22704 ;
  assign n22706 = ( n7308 & n22703 ) | ( n7308 & ~n22705 ) | ( n22703 & ~n22705 ) ;
  assign n22707 = ~x11 & n22706 ;
  assign n22708 = x11 | n22707 ;
  assign n22709 = ( ~n22706 & n22707 ) | ( ~n22706 & n22708 ) | ( n22707 & n22708 ) ;
  assign n22710 = n22698 & n22709 ;
  assign n22711 = n22246 | n22486 ;
  assign n22712 = ~n22487 & n22711 ;
  assign n22713 = n7305 & ~n20689 ;
  assign n22714 = n7300 & ~n20569 ;
  assign n22715 = n7302 & ~n20573 ;
  assign n22716 = n22714 | n22715 ;
  assign n22717 = n22713 | n22716 ;
  assign n22718 = ( n7308 & ~n22192 ) | ( n7308 & n22193 ) | ( ~n22192 & n22193 ) ;
  assign n22719 = n22717 | n22718 ;
  assign n22720 = x11 | n22719 ;
  assign n22721 = ~x11 & n22720 ;
  assign n22722 = ( ~n22719 & n22720 ) | ( ~n22719 & n22721 ) | ( n22720 & n22721 ) ;
  assign n22723 = n22712 & n22722 ;
  assign n22724 = n22722 & ~n22723 ;
  assign n22725 = ( n22712 & ~n22723 ) | ( n22712 & n22724 ) | ( ~n22723 & n22724 ) ;
  assign n22726 = n7305 & ~n20573 ;
  assign n22727 = n7300 & ~n20584 ;
  assign n22728 = n7302 & ~n20569 ;
  assign n22729 = n22727 | n22728 ;
  assign n22730 = n22726 | n22729 ;
  assign n22731 = n7308 | n22730 ;
  assign n22732 = ( ~n21860 & n22730 ) | ( ~n21860 & n22731 ) | ( n22730 & n22731 ) ;
  assign n22733 = ~x11 & n22732 ;
  assign n22734 = x11 | n22733 ;
  assign n22735 = ( ~n22732 & n22733 ) | ( ~n22732 & n22734 ) | ( n22733 & n22734 ) ;
  assign n22736 = ( n22248 & n22485 ) | ( n22248 & ~n22486 ) | ( n22485 & ~n22486 ) ;
  assign n22737 = ( n22258 & ~n22486 ) | ( n22258 & n22736 ) | ( ~n22486 & n22736 ) ;
  assign n22738 = n22735 & n22737 ;
  assign n22739 = n22735 | n22737 ;
  assign n22740 = ~n22738 & n22739 ;
  assign n22741 = n7305 & ~n20569 ;
  assign n22742 = n7300 & ~n20580 ;
  assign n22743 = n7302 & ~n20584 ;
  assign n22744 = n22742 | n22743 ;
  assign n22745 = n22741 | n22744 ;
  assign n22746 = n7308 & n21884 ;
  assign n22747 = ( n7308 & ~n21889 ) | ( n7308 & n22746 ) | ( ~n21889 & n22746 ) ;
  assign n22748 = n22745 | n22747 ;
  assign n22749 = x11 | n22748 ;
  assign n22750 = ~x11 & n22749 ;
  assign n22751 = ( ~n22748 & n22749 ) | ( ~n22748 & n22750 ) | ( n22749 & n22750 ) ;
  assign n22752 = ( n22260 & n22484 ) | ( n22260 & ~n22485 ) | ( n22484 & ~n22485 ) ;
  assign n22753 = ( n22270 & ~n22485 ) | ( n22270 & n22752 ) | ( ~n22485 & n22752 ) ;
  assign n22754 = n22751 & n22753 ;
  assign n22755 = n22751 | n22753 ;
  assign n22756 = ~n22754 & n22755 ;
  assign n22757 = n22480 | n22482 ;
  assign n22758 = ~n22483 & n22757 ;
  assign n22759 = n7305 & ~n20584 ;
  assign n22760 = n7300 & n20588 ;
  assign n22761 = n7302 & ~n20580 ;
  assign n22762 = n22760 | n22761 ;
  assign n22763 = n22759 | n22762 ;
  assign n22764 = n7308 | n22763 ;
  assign n22765 = ( ~n21901 & n22763 ) | ( ~n21901 & n22764 ) | ( n22763 & n22764 ) ;
  assign n22766 = ~x11 & n22765 ;
  assign n22767 = x11 | n22766 ;
  assign n22768 = ( ~n22765 & n22766 ) | ( ~n22765 & n22767 ) | ( n22766 & n22767 ) ;
  assign n22769 = n22758 & n22768 ;
  assign n22770 = n22758 | n22768 ;
  assign n22771 = ~n22769 & n22770 ;
  assign n22772 = n22302 | n22478 ;
  assign n22773 = ~n22479 & n22772 ;
  assign n22774 = n7305 & ~n20580 ;
  assign n22775 = n7300 & ~n20591 ;
  assign n22776 = n7302 & n20588 ;
  assign n22777 = n22775 | n22776 ;
  assign n22778 = n22774 | n22777 ;
  assign n22779 = n7308 | n22778 ;
  assign n22780 = ( n21840 & n22778 ) | ( n21840 & n22779 ) | ( n22778 & n22779 ) ;
  assign n22781 = x11 & n22780 ;
  assign n22782 = x11 & ~n22781 ;
  assign n22783 = ( n22780 & ~n22781 ) | ( n22780 & n22782 ) | ( ~n22781 & n22782 ) ;
  assign n22784 = n22319 | n22476 ;
  assign n22785 = ~n22477 & n22784 ;
  assign n22786 = n7305 & n20588 ;
  assign n22787 = n7300 & ~n20595 ;
  assign n22788 = n7302 & ~n20591 ;
  assign n22789 = n22787 | n22788 ;
  assign n22790 = n22786 | n22789 ;
  assign n22791 = n7308 | n22790 ;
  assign n22792 = ( n21526 & n22790 ) | ( n21526 & n22791 ) | ( n22790 & n22791 ) ;
  assign n22793 = x11 & n22792 ;
  assign n22794 = x11 & ~n22793 ;
  assign n22795 = ( n22792 & ~n22793 ) | ( n22792 & n22794 ) | ( ~n22793 & n22794 ) ;
  assign n22796 = n22345 | n22474 ;
  assign n22797 = n22472 | n22796 ;
  assign n22798 = ~n22475 & n22797 ;
  assign n22799 = n7305 & ~n20591 ;
  assign n22800 = n7300 & n20600 ;
  assign n22801 = n7302 & ~n20595 ;
  assign n22802 = n22800 | n22801 ;
  assign n22803 = n22799 | n22802 ;
  assign n22804 = n7308 & n21539 ;
  assign n22805 = ( n7308 & n21543 ) | ( n7308 & n22804 ) | ( n21543 & n22804 ) ;
  assign n22806 = n22803 | n22805 ;
  assign n22807 = x11 | n22806 ;
  assign n22808 = ~x11 & n22807 ;
  assign n22809 = ( ~n22806 & n22807 ) | ( ~n22806 & n22808 ) | ( n22807 & n22808 ) ;
  assign n22810 = n22798 & n22809 ;
  assign n22811 = n22469 & ~n22472 ;
  assign n22812 = n22471 & ~n22472 ;
  assign n22813 = n22811 | n22812 ;
  assign n22814 = n7305 & ~n20595 ;
  assign n22815 = n7300 & ~n20605 ;
  assign n22816 = n7302 & n20600 ;
  assign n22817 = n22815 | n22816 ;
  assign n22818 = n22814 | n22817 ;
  assign n22819 = n7308 | n22818 ;
  assign n22820 = ( ~n21554 & n22818 ) | ( ~n21554 & n22819 ) | ( n22818 & n22819 ) ;
  assign n22821 = ~x11 & n22820 ;
  assign n22822 = x11 | n22821 ;
  assign n22823 = ( ~n22820 & n22821 ) | ( ~n22820 & n22822 ) | ( n22821 & n22822 ) ;
  assign n22824 = n22813 & n22823 ;
  assign n22825 = n22813 & ~n22824 ;
  assign n22826 = ~n22813 & n22823 ;
  assign n22827 = n22825 | n22826 ;
  assign n22828 = n22464 & ~n22468 ;
  assign n22829 = n22467 & ~n22468 ;
  assign n22830 = n22828 | n22829 ;
  assign n22831 = n7305 & n20600 ;
  assign n22832 = n7300 & n20611 ;
  assign n22833 = n7302 & ~n20605 ;
  assign n22834 = n22832 | n22833 ;
  assign n22835 = n22831 | n22834 ;
  assign n22836 = n7308 | n22835 ;
  assign n22837 = ( ~n21432 & n22835 ) | ( ~n21432 & n22836 ) | ( n22835 & n22836 ) ;
  assign n22838 = ~x11 & n22837 ;
  assign n22839 = x11 | n22838 ;
  assign n22840 = ( ~n22837 & n22838 ) | ( ~n22837 & n22839 ) | ( n22838 & n22839 ) ;
  assign n22841 = n22830 & n22840 ;
  assign n22842 = n22830 & ~n22841 ;
  assign n22843 = ~n22830 & n22840 ;
  assign n22844 = n22842 | n22843 ;
  assign n22845 = n22460 | n22462 ;
  assign n22846 = ~n22463 & n22845 ;
  assign n22847 = n7305 & ~n20605 ;
  assign n22848 = n7300 & n20614 ;
  assign n22849 = n7302 & n20611 ;
  assign n22850 = n22848 | n22849 ;
  assign n22851 = n22847 | n22850 ;
  assign n22852 = n7308 | n22851 ;
  assign n22853 = ( ~n21275 & n22851 ) | ( ~n21275 & n22852 ) | ( n22851 & n22852 ) ;
  assign n22854 = ~x11 & n22853 ;
  assign n22855 = x11 | n22854 ;
  assign n22856 = ( ~n22853 & n22854 ) | ( ~n22853 & n22855 ) | ( n22854 & n22855 ) ;
  assign n22857 = n22846 & n22856 ;
  assign n22858 = n22386 | n22458 ;
  assign n22859 = ~n22459 & n22858 ;
  assign n22860 = n7305 & n20611 ;
  assign n22861 = n7300 & n20616 ;
  assign n22862 = n7302 & n20614 ;
  assign n22863 = n22861 | n22862 ;
  assign n22864 = n22860 | n22863 ;
  assign n22865 = n7308 | n22864 ;
  assign n22866 = ( n21293 & n22864 ) | ( n21293 & n22865 ) | ( n22864 & n22865 ) ;
  assign n22867 = x11 & n22866 ;
  assign n22868 = x11 & ~n22867 ;
  assign n22869 = ( n22866 & ~n22867 ) | ( n22866 & n22868 ) | ( ~n22867 & n22868 ) ;
  assign n22870 = n22859 & n22869 ;
  assign n22871 = n22454 | n22456 ;
  assign n22872 = ~n22457 & n22871 ;
  assign n22873 = n7305 & n20614 ;
  assign n22874 = n7300 & n20619 ;
  assign n22875 = n7302 | n22874 ;
  assign n22876 = ( n20616 & n22874 ) | ( n20616 & n22875 ) | ( n22874 & n22875 ) ;
  assign n22877 = n22873 | n22876 ;
  assign n22878 = n7308 | n22877 ;
  assign n22879 = ( n21302 & n22877 ) | ( n21302 & n22878 ) | ( n22877 & n22878 ) ;
  assign n22880 = x11 & n22879 ;
  assign n22881 = x11 & ~n22880 ;
  assign n22882 = ( n22879 & ~n22880 ) | ( n22879 & n22881 ) | ( ~n22880 & n22881 ) ;
  assign n22883 = n22872 & n22882 ;
  assign n22884 = n7300 & n20622 ;
  assign n22885 = n7302 | n22884 ;
  assign n22886 = ( n20619 & n22884 ) | ( n20619 & n22885 ) | ( n22884 & n22885 ) ;
  assign n22887 = n7305 | n22886 ;
  assign n22888 = ( n20616 & n22886 ) | ( n20616 & n22887 ) | ( n22886 & n22887 ) ;
  assign n22889 = n7308 | n22888 ;
  assign n22890 = ( n21190 & n22888 ) | ( n21190 & n22889 ) | ( n22888 & n22889 ) ;
  assign n22891 = ~x11 & n22890 ;
  assign n22892 = x11 & ~n22890 ;
  assign n22893 = n22891 | n22892 ;
  assign n22894 = n22414 | n22452 ;
  assign n22895 = ~n22453 & n22894 ;
  assign n22896 = n22893 & n22895 ;
  assign n22897 = n7300 & ~n20625 ;
  assign n22898 = n7302 | n22897 ;
  assign n22899 = ( n20622 & n22897 ) | ( n20622 & n22898 ) | ( n22897 & n22898 ) ;
  assign n22900 = n7305 | n22899 ;
  assign n22901 = ( n20619 & n22899 ) | ( n20619 & n22900 ) | ( n22899 & n22900 ) ;
  assign n22902 = n7308 | n22901 ;
  assign n22903 = ( ~n21056 & n22901 ) | ( ~n21056 & n22902 ) | ( n22901 & n22902 ) ;
  assign n22904 = ~x11 & n22903 ;
  assign n22905 = x11 | n22904 ;
  assign n22906 = ( ~n22903 & n22904 ) | ( ~n22903 & n22905 ) | ( n22904 & n22905 ) ;
  assign n22907 = n22440 & ~n22451 ;
  assign n22908 = ( n22450 & ~n22451 ) | ( n22450 & n22907 ) | ( ~n22451 & n22907 ) ;
  assign n22909 = n22906 & n22908 ;
  assign n22910 = n22906 | n22908 ;
  assign n22911 = ~n22909 & n22910 ;
  assign n22912 = n22424 | n22435 ;
  assign n22913 = ~n22438 & n22912 ;
  assign n22914 = n7305 & n20622 ;
  assign n22915 = n7300 & ~n20630 ;
  assign n22916 = n7302 & ~n20625 ;
  assign n22917 = n22915 | n22916 ;
  assign n22918 = n22914 | n22917 ;
  assign n22919 = n7308 | n22918 ;
  assign n22920 = ( n21114 & n22918 ) | ( n21114 & n22919 ) | ( n22918 & n22919 ) ;
  assign n22921 = x11 & n22920 ;
  assign n22922 = x11 | n22920 ;
  assign n22923 = ~n22921 & n22922 ;
  assign n22924 = n22913 & n22923 ;
  assign n22925 = n22415 | n22423 ;
  assign n22926 = ~n22424 & n22925 ;
  assign n22927 = n7305 & ~n20625 ;
  assign n22928 = n7300 & n20633 ;
  assign n22929 = n7302 & ~n20630 ;
  assign n22930 = n22928 | n22929 ;
  assign n22931 = n22927 | n22930 ;
  assign n22932 = n7308 | n22931 ;
  assign n22933 = ( ~n21129 & n22931 ) | ( ~n21129 & n22932 ) | ( n22931 & n22932 ) ;
  assign n22934 = ~x11 & n22933 ;
  assign n22935 = x11 | n22934 ;
  assign n22936 = ( ~n22933 & n22934 ) | ( ~n22933 & n22935 ) | ( n22934 & n22935 ) ;
  assign n22937 = n22926 & n22936 ;
  assign n22938 = n22926 | n22936 ;
  assign n22939 = ~n22937 & n22938 ;
  assign n22940 = ( x11 & n17237 ) | ( x11 & n20642 ) | ( n17237 & n20642 ) ;
  assign n22941 = n7308 & n21069 ;
  assign n22942 = n7302 & ~n20642 ;
  assign n22943 = n7305 & ~n20640 ;
  assign n22944 = n22942 | n22943 ;
  assign n22945 = n22941 | n22944 ;
  assign n22946 = x11 | n22945 ;
  assign n22947 = ~x11 & n22946 ;
  assign n22948 = ( ~n22945 & n22946 ) | ( ~n22945 & n22947 ) | ( n22946 & n22947 ) ;
  assign n22949 = n22940 & n22948 ;
  assign n22950 = n35 & ~n20642 ;
  assign n22951 = n7305 & n20633 ;
  assign n22952 = n7300 & ~n20642 ;
  assign n22953 = n7302 & ~n20640 ;
  assign n22954 = n22952 | n22953 ;
  assign n22955 = n22951 | n22954 ;
  assign n22956 = n7308 & n21085 ;
  assign n22957 = n22955 | n22956 ;
  assign n22958 = ~x11 & n22957 ;
  assign n22959 = x11 | n22958 ;
  assign n22960 = ( ~n22957 & n22958 ) | ( ~n22957 & n22959 ) | ( n22958 & n22959 ) ;
  assign n22961 = n22950 & n22960 ;
  assign n22962 = n22949 & n22961 ;
  assign n22963 = n22949 & n22960 ;
  assign n22964 = n22950 | n22963 ;
  assign n22965 = ~n22962 & n22964 ;
  assign n22966 = n7305 & ~n20630 ;
  assign n22967 = n7300 & ~n20640 ;
  assign n22968 = n7302 & n20633 ;
  assign n22969 = n22967 | n22968 ;
  assign n22970 = n22966 | n22969 ;
  assign n22971 = n7308 | n22970 ;
  assign n22972 = ( n21099 & n22970 ) | ( n21099 & n22971 ) | ( n22970 & n22971 ) ;
  assign n22973 = x11 & n22972 ;
  assign n22974 = x11 | n22972 ;
  assign n22975 = ~n22973 & n22974 ;
  assign n22976 = n22965 & n22975 ;
  assign n22977 = n22962 | n22976 ;
  assign n22978 = n22939 & n22977 ;
  assign n22979 = n22937 | n22978 ;
  assign n22980 = n22923 & ~n22924 ;
  assign n22981 = ( n22913 & ~n22924 ) | ( n22913 & n22980 ) | ( ~n22924 & n22980 ) ;
  assign n22982 = n22979 & n22981 ;
  assign n22983 = n22924 | n22982 ;
  assign n22984 = n22911 & n22983 ;
  assign n22985 = n22909 | n22984 ;
  assign n22986 = n22893 | n22895 ;
  assign n22987 = ~n22896 & n22986 ;
  assign n22988 = n22985 & n22987 ;
  assign n22989 = n22896 | n22988 ;
  assign n22990 = n22872 & ~n22883 ;
  assign n22991 = n22882 & ~n22883 ;
  assign n22992 = n22990 | n22991 ;
  assign n22993 = n22989 & n22992 ;
  assign n22994 = n22883 | n22993 ;
  assign n22995 = n22869 & ~n22870 ;
  assign n22996 = ( n22859 & ~n22870 ) | ( n22859 & n22995 ) | ( ~n22870 & n22995 ) ;
  assign n22997 = n22994 & n22996 ;
  assign n22998 = n22846 | n22856 ;
  assign n22999 = ~n22857 & n22998 ;
  assign n23000 = ( n22870 & n22997 ) | ( n22870 & n22999 ) | ( n22997 & n22999 ) ;
  assign n23001 = n22857 | n23000 ;
  assign n23002 = n22844 & n23001 ;
  assign n23003 = n22841 | n23002 ;
  assign n23004 = n22827 & n23003 ;
  assign n23005 = n22824 | n23004 ;
  assign n23006 = n22809 & ~n22810 ;
  assign n23007 = ( n22798 & ~n22810 ) | ( n22798 & n23006 ) | ( ~n22810 & n23006 ) ;
  assign n23008 = n23005 & n23007 ;
  assign n23009 = n22810 | n23008 ;
  assign n23010 = ( n22785 & n22795 ) | ( n22785 & n23009 ) | ( n22795 & n23009 ) ;
  assign n23011 = ( n22773 & n22783 ) | ( n22773 & n23010 ) | ( n22783 & n23010 ) ;
  assign n23012 = n22771 & n23011 ;
  assign n23013 = n22769 | n23012 ;
  assign n23014 = n22756 & n23013 ;
  assign n23015 = n22754 | n23014 ;
  assign n23016 = n22740 & n23015 ;
  assign n23017 = n22738 | n23016 ;
  assign n23018 = n22725 & n23017 ;
  assign n23019 = n22723 | n23018 ;
  assign n23020 = n22698 & ~n22710 ;
  assign n23021 = ~n22698 & n22709 ;
  assign n23022 = n23020 | n23021 ;
  assign n23023 = n23019 & n23022 ;
  assign n23024 = n22685 | n22695 ;
  assign n23025 = ~n22696 & n23024 ;
  assign n23026 = ( n22710 & n23023 ) | ( n22710 & n23025 ) | ( n23023 & n23025 ) ;
  assign n23027 = n22696 | n23026 ;
  assign n23028 = n22671 | n22683 ;
  assign n23029 = ( ~n22682 & n22683 ) | ( ~n22682 & n23028 ) | ( n22683 & n23028 ) ;
  assign n23030 = n23027 & ~n23029 ;
  assign n23031 = n22683 | n23030 ;
  assign n23032 = ~n22668 & n23031 ;
  assign n23033 = n22666 | n23032 ;
  assign n23034 = n22651 & n23033 ;
  assign n23224 = n22651 | n23033 ;
  assign n23225 = ~n23034 & n23224 ;
  assign n23226 = ( n20720 & n20729 ) | ( n20720 & n20730 ) | ( n20729 & n20730 ) ;
  assign n23227 = n20547 | n20729 ;
  assign n23228 = n20720 | n23227 ;
  assign n23229 = ~n23226 & n23228 ;
  assign n23230 = n5503 & ~n20724 ;
  assign n23231 = n5512 & n20546 ;
  assign n23232 = n5508 & ~n20542 ;
  assign n23233 = n23231 | n23232 ;
  assign n23234 = n23230 | n23233 ;
  assign n23235 = n5515 | n23234 ;
  assign n23236 = ( n23229 & n23234 ) | ( n23229 & n23235 ) | ( n23234 & n23235 ) ;
  assign n23237 = x8 & n23236 ;
  assign n23238 = x8 & ~n23237 ;
  assign n23239 = ( n23236 & ~n23237 ) | ( n23236 & n23238 ) | ( ~n23237 & n23238 ) ;
  assign n23040 = n20547 | n20548 ;
  assign n23041 = ~n20718 & n23040 ;
  assign n23042 = n20720 | n23041 ;
  assign n23240 = n5503 & ~n20542 ;
  assign n23241 = n5512 & ~n20710 ;
  assign n23242 = n5508 & n20546 ;
  assign n23243 = n23241 | n23242 ;
  assign n23244 = n23240 | n23243 ;
  assign n23245 = n5515 | n23244 ;
  assign n23246 = ( ~n23042 & n23244 ) | ( ~n23042 & n23245 ) | ( n23244 & n23245 ) ;
  assign n23247 = ~x8 & n23246 ;
  assign n23248 = x8 | n23247 ;
  assign n23249 = ( ~n23246 & n23247 ) | ( ~n23246 & n23248 ) | ( n23247 & n23248 ) ;
  assign n23250 = n5503 & n20546 ;
  assign n23251 = n5512 & n20556 ;
  assign n23252 = n5508 & ~n20710 ;
  assign n23253 = n23251 | n23252 ;
  assign n23254 = n23250 | n23253 ;
  assign n21035 = n20713 | n20714 ;
  assign n21036 = ( n20706 & n20716 ) | ( n20706 & ~n21035 ) | ( n20716 & ~n21035 ) ;
  assign n21037 = ( n20715 & n21034 ) | ( n20715 & ~n21036 ) | ( n21034 & ~n21036 ) ;
  assign n21031 = n20711 | n20718 ;
  assign n23255 = n5515 & n21031 ;
  assign n23256 = ~n21037 & n23255 ;
  assign n23257 = ( n5515 & n23254 ) | ( n5515 & ~n23256 ) | ( n23254 & ~n23256 ) ;
  assign n23258 = x8 & n23257 ;
  assign n23259 = x8 & ~n23258 ;
  assign n23260 = ( n23257 & ~n23258 ) | ( n23257 & n23259 ) | ( ~n23258 & n23259 ) ;
  assign n23261 = n22710 | n23025 ;
  assign n23262 = n23023 | n23261 ;
  assign n23263 = ~n23026 & n23262 ;
  assign n23264 = n5503 & ~n20710 ;
  assign n23265 = n5512 & ~n20552 ;
  assign n23266 = n5508 & n20556 ;
  assign n23267 = n23265 | n23266 ;
  assign n23268 = n23264 | n23267 ;
  assign n23269 = n5515 | n23268 ;
  assign n23270 = ( ~n22641 & n23268 ) | ( ~n22641 & n23269 ) | ( n23268 & n23269 ) ;
  assign n23271 = ~x8 & n23270 ;
  assign n23272 = x8 | n23271 ;
  assign n23273 = ( ~n23270 & n23271 ) | ( ~n23270 & n23272 ) | ( n23271 & n23272 ) ;
  assign n23274 = n23263 & n23273 ;
  assign n23275 = n23019 & ~n23023 ;
  assign n23276 = n23022 & ~n23023 ;
  assign n23277 = n23275 | n23276 ;
  assign n23278 = n5503 & n20556 ;
  assign n23279 = n5512 & n20562 ;
  assign n23280 = n5508 & ~n20552 ;
  assign n23281 = n23279 | n23280 ;
  assign n23282 = n23278 | n23281 ;
  assign n23283 = n5515 | n23282 ;
  assign n23284 = ( ~n22655 & n23282 ) | ( ~n22655 & n23283 ) | ( n23282 & n23283 ) ;
  assign n23285 = ~x8 & n23284 ;
  assign n23286 = x8 | n23285 ;
  assign n23287 = ( ~n23284 & n23285 ) | ( ~n23284 & n23286 ) | ( n23285 & n23286 ) ;
  assign n23288 = n23277 & n23287 ;
  assign n23289 = n23277 & ~n23288 ;
  assign n23290 = ~n23277 & n23287 ;
  assign n23291 = n23289 | n23290 ;
  assign n23292 = n22725 | n23017 ;
  assign n23293 = ~n23018 & n23292 ;
  assign n23294 = n5503 & ~n20552 ;
  assign n23295 = n5512 & n20560 ;
  assign n23296 = n5508 & n20562 ;
  assign n23297 = n23295 | n23296 ;
  assign n23298 = n23294 | n23297 ;
  assign n23299 = n5515 & n22510 ;
  assign n23300 = ~n22512 & n23299 ;
  assign n23301 = ( n5515 & n23298 ) | ( n5515 & ~n23300 ) | ( n23298 & ~n23300 ) ;
  assign n23302 = x8 & n23301 ;
  assign n23303 = x8 & ~n23302 ;
  assign n23304 = ( n23301 & ~n23302 ) | ( n23301 & n23303 ) | ( ~n23302 & n23303 ) ;
  assign n23305 = n23293 & n23304 ;
  assign n23306 = n22740 | n23015 ;
  assign n23307 = ~n23016 & n23306 ;
  assign n23308 = n5503 & n20562 ;
  assign n23309 = n5512 & ~n20689 ;
  assign n23310 = n5508 & n20560 ;
  assign n23311 = n23309 | n23310 ;
  assign n23312 = n23308 | n23311 ;
  assign n23313 = n5515 | n23312 ;
  assign n23314 = ( ~n21044 & n23312 ) | ( ~n21044 & n23313 ) | ( n23312 & n23313 ) ;
  assign n23315 = ~x8 & n23314 ;
  assign n23316 = x8 | n23315 ;
  assign n23317 = ( ~n23314 & n23315 ) | ( ~n23314 & n23316 ) | ( n23315 & n23316 ) ;
  assign n23318 = n23307 & n23317 ;
  assign n23319 = n22756 | n23013 ;
  assign n23320 = ~n23014 & n23319 ;
  assign n23321 = n5503 & n20560 ;
  assign n23322 = n5512 & ~n20573 ;
  assign n23323 = n5508 & ~n20689 ;
  assign n23324 = n23322 | n23323 ;
  assign n23325 = n23321 | n23324 ;
  assign n23326 = n5515 & ~n22176 ;
  assign n23327 = ~n22173 & n23326 ;
  assign n23328 = ( n5515 & n23325 ) | ( n5515 & ~n23327 ) | ( n23325 & ~n23327 ) ;
  assign n23329 = ~x8 & n23328 ;
  assign n23330 = x8 | n23329 ;
  assign n23331 = ( ~n23328 & n23329 ) | ( ~n23328 & n23330 ) | ( n23329 & n23330 ) ;
  assign n23332 = n23320 & n23331 ;
  assign n23333 = n22771 | n23011 ;
  assign n23334 = ~n23012 & n23333 ;
  assign n23335 = n5503 & ~n20689 ;
  assign n23336 = n5512 & ~n20569 ;
  assign n23337 = n5508 & ~n20573 ;
  assign n23338 = n23336 | n23337 ;
  assign n23339 = n23335 | n23338 ;
  assign n23340 = ( n5515 & ~n22192 ) | ( n5515 & n22193 ) | ( ~n22192 & n22193 ) ;
  assign n23341 = n23339 | n23340 ;
  assign n23342 = x8 | n23341 ;
  assign n23343 = ~x8 & n23342 ;
  assign n23344 = ( ~n23341 & n23342 ) | ( ~n23341 & n23343 ) | ( n23342 & n23343 ) ;
  assign n23345 = n23334 & n23344 ;
  assign n23346 = n23344 & ~n23345 ;
  assign n23347 = ( n23334 & ~n23345 ) | ( n23334 & n23346 ) | ( ~n23345 & n23346 ) ;
  assign n23348 = n5503 & ~n20573 ;
  assign n23349 = n5512 & ~n20584 ;
  assign n23350 = n5508 & ~n20569 ;
  assign n23351 = n23349 | n23350 ;
  assign n23352 = n23348 | n23351 ;
  assign n23353 = n5515 | n23352 ;
  assign n23354 = ( ~n21860 & n23352 ) | ( ~n21860 & n23353 ) | ( n23352 & n23353 ) ;
  assign n23355 = ~x8 & n23354 ;
  assign n23356 = x8 | n23355 ;
  assign n23357 = ( ~n23354 & n23355 ) | ( ~n23354 & n23356 ) | ( n23355 & n23356 ) ;
  assign n23358 = ( n22773 & n23010 ) | ( n22773 & ~n23011 ) | ( n23010 & ~n23011 ) ;
  assign n23359 = ( n22783 & ~n23011 ) | ( n22783 & n23358 ) | ( ~n23011 & n23358 ) ;
  assign n23360 = n23357 & n23359 ;
  assign n23361 = n23357 | n23359 ;
  assign n23362 = ~n23360 & n23361 ;
  assign n23363 = n5503 & ~n20569 ;
  assign n23364 = n5512 & ~n20580 ;
  assign n23365 = n5508 & ~n20584 ;
  assign n23366 = n23364 | n23365 ;
  assign n23367 = n23363 | n23366 ;
  assign n23368 = n5515 & n21884 ;
  assign n23369 = ( n5515 & ~n21889 ) | ( n5515 & n23368 ) | ( ~n21889 & n23368 ) ;
  assign n23370 = n23367 | n23369 ;
  assign n23371 = x8 | n23370 ;
  assign n23372 = ~x8 & n23371 ;
  assign n23373 = ( ~n23370 & n23371 ) | ( ~n23370 & n23372 ) | ( n23371 & n23372 ) ;
  assign n23374 = ( n22785 & n23009 ) | ( n22785 & ~n23010 ) | ( n23009 & ~n23010 ) ;
  assign n23375 = ( n22795 & ~n23010 ) | ( n22795 & n23374 ) | ( ~n23010 & n23374 ) ;
  assign n23376 = n23373 & n23375 ;
  assign n23377 = n23373 | n23375 ;
  assign n23378 = ~n23376 & n23377 ;
  assign n23379 = n23005 | n23007 ;
  assign n23380 = ~n23008 & n23379 ;
  assign n23381 = n5503 & ~n20584 ;
  assign n23382 = n5512 & n20588 ;
  assign n23383 = n5508 & ~n20580 ;
  assign n23384 = n23382 | n23383 ;
  assign n23385 = n23381 | n23384 ;
  assign n23386 = n5515 | n23385 ;
  assign n23387 = ( ~n21901 & n23385 ) | ( ~n21901 & n23386 ) | ( n23385 & n23386 ) ;
  assign n23388 = ~x8 & n23387 ;
  assign n23389 = x8 | n23388 ;
  assign n23390 = ( ~n23387 & n23388 ) | ( ~n23387 & n23389 ) | ( n23388 & n23389 ) ;
  assign n23391 = n23380 & n23390 ;
  assign n23392 = n23380 | n23390 ;
  assign n23393 = ~n23391 & n23392 ;
  assign n23394 = n22827 | n23003 ;
  assign n23395 = ~n23004 & n23394 ;
  assign n23396 = n5503 & ~n20580 ;
  assign n23397 = n5512 & ~n20591 ;
  assign n23398 = n5508 & n20588 ;
  assign n23399 = n23397 | n23398 ;
  assign n23400 = n23396 | n23399 ;
  assign n23401 = n5515 | n23400 ;
  assign n23402 = ( n21840 & n23400 ) | ( n21840 & n23401 ) | ( n23400 & n23401 ) ;
  assign n23403 = x8 & n23402 ;
  assign n23404 = x8 & ~n23403 ;
  assign n23405 = ( n23402 & ~n23403 ) | ( n23402 & n23404 ) | ( ~n23403 & n23404 ) ;
  assign n23406 = n22844 | n23001 ;
  assign n23407 = ~n23002 & n23406 ;
  assign n23408 = n5503 & n20588 ;
  assign n23409 = n5512 & ~n20595 ;
  assign n23410 = n5508 & ~n20591 ;
  assign n23411 = n23409 | n23410 ;
  assign n23412 = n23408 | n23411 ;
  assign n23413 = n5515 | n23412 ;
  assign n23414 = ( n21526 & n23412 ) | ( n21526 & n23413 ) | ( n23412 & n23413 ) ;
  assign n23415 = x8 & n23414 ;
  assign n23416 = x8 & ~n23415 ;
  assign n23417 = ( n23414 & ~n23415 ) | ( n23414 & n23416 ) | ( ~n23415 & n23416 ) ;
  assign n23418 = n22870 | n22999 ;
  assign n23419 = n22997 | n23418 ;
  assign n23420 = ~n23000 & n23419 ;
  assign n23421 = n5503 & ~n20591 ;
  assign n23422 = n5512 & n20600 ;
  assign n23423 = n5508 & ~n20595 ;
  assign n23424 = n23422 | n23423 ;
  assign n23425 = n23421 | n23424 ;
  assign n23426 = n5515 & n21539 ;
  assign n23427 = ( n5515 & n21543 ) | ( n5515 & n23426 ) | ( n21543 & n23426 ) ;
  assign n23428 = n23425 | n23427 ;
  assign n23429 = x8 | n23428 ;
  assign n23430 = ~x8 & n23429 ;
  assign n23431 = ( ~n23428 & n23429 ) | ( ~n23428 & n23430 ) | ( n23429 & n23430 ) ;
  assign n23432 = n23420 & n23431 ;
  assign n23433 = n22994 & ~n22997 ;
  assign n23434 = n22996 & ~n22997 ;
  assign n23435 = n23433 | n23434 ;
  assign n23436 = n5503 & ~n20595 ;
  assign n23437 = n5512 & ~n20605 ;
  assign n23438 = n5508 & n20600 ;
  assign n23439 = n23437 | n23438 ;
  assign n23440 = n23436 | n23439 ;
  assign n23441 = n5515 | n23440 ;
  assign n23442 = ( ~n21554 & n23440 ) | ( ~n21554 & n23441 ) | ( n23440 & n23441 ) ;
  assign n23443 = ~x8 & n23442 ;
  assign n23444 = x8 | n23443 ;
  assign n23445 = ( ~n23442 & n23443 ) | ( ~n23442 & n23444 ) | ( n23443 & n23444 ) ;
  assign n23446 = n23435 & n23445 ;
  assign n23447 = n23435 & ~n23446 ;
  assign n23448 = ~n23435 & n23445 ;
  assign n23449 = n23447 | n23448 ;
  assign n23450 = n22989 & ~n22993 ;
  assign n23451 = n22992 & ~n22993 ;
  assign n23452 = n23450 | n23451 ;
  assign n23453 = n5503 & n20600 ;
  assign n23454 = n5512 & n20611 ;
  assign n23455 = n5508 & ~n20605 ;
  assign n23456 = n23454 | n23455 ;
  assign n23457 = n23453 | n23456 ;
  assign n23458 = n5515 | n23457 ;
  assign n23459 = ( ~n21432 & n23457 ) | ( ~n21432 & n23458 ) | ( n23457 & n23458 ) ;
  assign n23460 = ~x8 & n23459 ;
  assign n23461 = x8 | n23460 ;
  assign n23462 = ( ~n23459 & n23460 ) | ( ~n23459 & n23461 ) | ( n23460 & n23461 ) ;
  assign n23463 = n23452 & n23462 ;
  assign n23464 = n23452 & ~n23463 ;
  assign n23465 = ~n23452 & n23462 ;
  assign n23466 = n23464 | n23465 ;
  assign n23467 = n22985 | n22987 ;
  assign n23468 = ~n22988 & n23467 ;
  assign n23469 = n5503 & ~n20605 ;
  assign n23470 = n5512 & n20614 ;
  assign n23471 = n5508 & n20611 ;
  assign n23472 = n23470 | n23471 ;
  assign n23473 = n23469 | n23472 ;
  assign n23474 = n5515 | n23473 ;
  assign n23475 = ( ~n21275 & n23473 ) | ( ~n21275 & n23474 ) | ( n23473 & n23474 ) ;
  assign n23476 = ~x8 & n23475 ;
  assign n23477 = x8 | n23476 ;
  assign n23478 = ( ~n23475 & n23476 ) | ( ~n23475 & n23477 ) | ( n23476 & n23477 ) ;
  assign n23479 = n23468 & n23478 ;
  assign n23480 = n22911 | n22983 ;
  assign n23481 = ~n22984 & n23480 ;
  assign n23482 = n5503 & n20611 ;
  assign n23483 = n5512 & n20616 ;
  assign n23484 = n5508 & n20614 ;
  assign n23485 = n23483 | n23484 ;
  assign n23486 = n23482 | n23485 ;
  assign n23487 = n5515 | n23486 ;
  assign n23488 = ( n21293 & n23486 ) | ( n21293 & n23487 ) | ( n23486 & n23487 ) ;
  assign n23489 = x8 & n23488 ;
  assign n23490 = x8 & ~n23489 ;
  assign n23491 = ( n23488 & ~n23489 ) | ( n23488 & n23490 ) | ( ~n23489 & n23490 ) ;
  assign n23492 = n23481 & n23491 ;
  assign n23493 = n22979 | n22981 ;
  assign n23494 = ~n22982 & n23493 ;
  assign n23495 = n5503 & n20614 ;
  assign n23496 = n5512 & n20619 ;
  assign n23497 = n5508 | n23496 ;
  assign n23498 = ( n20616 & n23496 ) | ( n20616 & n23497 ) | ( n23496 & n23497 ) ;
  assign n23499 = n23495 | n23498 ;
  assign n23500 = n5515 | n23499 ;
  assign n23501 = ( n21302 & n23499 ) | ( n21302 & n23500 ) | ( n23499 & n23500 ) ;
  assign n23502 = x8 & n23501 ;
  assign n23503 = x8 & ~n23502 ;
  assign n23504 = ( n23501 & ~n23502 ) | ( n23501 & n23503 ) | ( ~n23502 & n23503 ) ;
  assign n23505 = n23494 & n23504 ;
  assign n23506 = n5512 & n20622 ;
  assign n23507 = n5508 | n23506 ;
  assign n23508 = ( n20619 & n23506 ) | ( n20619 & n23507 ) | ( n23506 & n23507 ) ;
  assign n23509 = n5503 | n23508 ;
  assign n23510 = ( n20616 & n23508 ) | ( n20616 & n23509 ) | ( n23508 & n23509 ) ;
  assign n23511 = n5515 | n23510 ;
  assign n23512 = ( n21190 & n23510 ) | ( n21190 & n23511 ) | ( n23510 & n23511 ) ;
  assign n23513 = ~x8 & n23512 ;
  assign n23514 = x8 & ~n23512 ;
  assign n23515 = n23513 | n23514 ;
  assign n23516 = n22939 | n22977 ;
  assign n23517 = ~n22978 & n23516 ;
  assign n23518 = n23515 & n23517 ;
  assign n23519 = n5512 & ~n20625 ;
  assign n23520 = n5508 | n23519 ;
  assign n23521 = ( n20622 & n23519 ) | ( n20622 & n23520 ) | ( n23519 & n23520 ) ;
  assign n23522 = n5503 | n23521 ;
  assign n23523 = ( n20619 & n23521 ) | ( n20619 & n23522 ) | ( n23521 & n23522 ) ;
  assign n23524 = n5515 | n23523 ;
  assign n23525 = ( ~n21056 & n23523 ) | ( ~n21056 & n23524 ) | ( n23523 & n23524 ) ;
  assign n23526 = ~x8 & n23525 ;
  assign n23527 = x8 | n23526 ;
  assign n23528 = ( ~n23525 & n23526 ) | ( ~n23525 & n23527 ) | ( n23526 & n23527 ) ;
  assign n23529 = n22965 & ~n22976 ;
  assign n23530 = ( n22975 & ~n22976 ) | ( n22975 & n23529 ) | ( ~n22976 & n23529 ) ;
  assign n23531 = n23528 & n23530 ;
  assign n23532 = n23528 | n23530 ;
  assign n23533 = ~n23531 & n23532 ;
  assign n23534 = n22949 | n22960 ;
  assign n23535 = ~n22963 & n23534 ;
  assign n23536 = n5503 & n20622 ;
  assign n23537 = n5512 & ~n20630 ;
  assign n23538 = n5508 & ~n20625 ;
  assign n23539 = n23537 | n23538 ;
  assign n23540 = n23536 | n23539 ;
  assign n23541 = n5515 | n23540 ;
  assign n23542 = ( n21114 & n23540 ) | ( n21114 & n23541 ) | ( n23540 & n23541 ) ;
  assign n23543 = x8 & n23542 ;
  assign n23544 = x8 | n23542 ;
  assign n23545 = ~n23543 & n23544 ;
  assign n23546 = n23535 & n23545 ;
  assign n23547 = n22940 | n22948 ;
  assign n23548 = ~n22949 & n23547 ;
  assign n23549 = n5503 & ~n20625 ;
  assign n23550 = n5512 & n20633 ;
  assign n23551 = n5508 & ~n20630 ;
  assign n23552 = n23550 | n23551 ;
  assign n23553 = n23549 | n23552 ;
  assign n23554 = n5515 | n23553 ;
  assign n23555 = ( ~n21129 & n23553 ) | ( ~n21129 & n23554 ) | ( n23553 & n23554 ) ;
  assign n23556 = ~x8 & n23555 ;
  assign n23557 = x8 | n23556 ;
  assign n23558 = ( ~n23555 & n23556 ) | ( ~n23555 & n23557 ) | ( n23556 & n23557 ) ;
  assign n23559 = n23548 & n23558 ;
  assign n23560 = n23548 | n23558 ;
  assign n23561 = ~n23559 & n23560 ;
  assign n23562 = ( x8 & n17771 ) | ( x8 & n20642 ) | ( n17771 & n20642 ) ;
  assign n23563 = n5515 & n21069 ;
  assign n23564 = n5508 & ~n20642 ;
  assign n23565 = n5503 & ~n20640 ;
  assign n23566 = n23564 | n23565 ;
  assign n23567 = n23563 | n23566 ;
  assign n23568 = x8 | n23567 ;
  assign n23569 = ~x8 & n23568 ;
  assign n23570 = ( ~n23567 & n23568 ) | ( ~n23567 & n23569 ) | ( n23568 & n23569 ) ;
  assign n23571 = n23562 & n23570 ;
  assign n23572 = n7298 & ~n20642 ;
  assign n23573 = n5503 & n20633 ;
  assign n23574 = n5512 & ~n20642 ;
  assign n23575 = n5508 & ~n20640 ;
  assign n23576 = n23574 | n23575 ;
  assign n23577 = n23573 | n23576 ;
  assign n23578 = n5515 & n21085 ;
  assign n23579 = n23577 | n23578 ;
  assign n23580 = ~x8 & n23579 ;
  assign n23581 = x8 | n23580 ;
  assign n23582 = ( ~n23579 & n23580 ) | ( ~n23579 & n23581 ) | ( n23580 & n23581 ) ;
  assign n23583 = n23572 & n23582 ;
  assign n23584 = n23571 & n23583 ;
  assign n23585 = n23571 & n23582 ;
  assign n23586 = n23572 | n23585 ;
  assign n23587 = ~n23584 & n23586 ;
  assign n23588 = n5503 & ~n20630 ;
  assign n23589 = n5512 & ~n20640 ;
  assign n23590 = n5508 & n20633 ;
  assign n23591 = n23589 | n23590 ;
  assign n23592 = n23588 | n23591 ;
  assign n23593 = n5515 | n23592 ;
  assign n23594 = ( n21099 & n23592 ) | ( n21099 & n23593 ) | ( n23592 & n23593 ) ;
  assign n23595 = x8 & n23594 ;
  assign n23596 = x8 | n23594 ;
  assign n23597 = ~n23595 & n23596 ;
  assign n23598 = n23587 & n23597 ;
  assign n23599 = n23584 | n23598 ;
  assign n23600 = n23561 & n23599 ;
  assign n23601 = n23559 | n23600 ;
  assign n23602 = n23545 & ~n23546 ;
  assign n23603 = ( n23535 & ~n23546 ) | ( n23535 & n23602 ) | ( ~n23546 & n23602 ) ;
  assign n23604 = n23601 & n23603 ;
  assign n23605 = n23546 | n23604 ;
  assign n23606 = n23533 & n23605 ;
  assign n23607 = n23531 | n23606 ;
  assign n23608 = n23515 | n23517 ;
  assign n23609 = ~n23518 & n23608 ;
  assign n23610 = n23607 & n23609 ;
  assign n23611 = n23518 | n23610 ;
  assign n23612 = n23494 & ~n23505 ;
  assign n23613 = n23504 & ~n23505 ;
  assign n23614 = n23612 | n23613 ;
  assign n23615 = n23611 & n23614 ;
  assign n23616 = n23505 | n23615 ;
  assign n23617 = n23491 & ~n23492 ;
  assign n23618 = ( n23481 & ~n23492 ) | ( n23481 & n23617 ) | ( ~n23492 & n23617 ) ;
  assign n23619 = n23616 & n23618 ;
  assign n23620 = n23468 | n23478 ;
  assign n23621 = ~n23479 & n23620 ;
  assign n23622 = ( n23492 & n23619 ) | ( n23492 & n23621 ) | ( n23619 & n23621 ) ;
  assign n23623 = n23479 | n23622 ;
  assign n23624 = n23466 & n23623 ;
  assign n23625 = n23463 | n23624 ;
  assign n23626 = n23449 & n23625 ;
  assign n23627 = n23446 | n23626 ;
  assign n23628 = n23431 & ~n23432 ;
  assign n23629 = ( n23420 & ~n23432 ) | ( n23420 & n23628 ) | ( ~n23432 & n23628 ) ;
  assign n23630 = n23627 & n23629 ;
  assign n23631 = n23432 | n23630 ;
  assign n23632 = ( n23407 & n23417 ) | ( n23407 & n23631 ) | ( n23417 & n23631 ) ;
  assign n23633 = ( n23395 & n23405 ) | ( n23395 & n23632 ) | ( n23405 & n23632 ) ;
  assign n23634 = n23393 & n23633 ;
  assign n23635 = n23391 | n23634 ;
  assign n23636 = n23378 & n23635 ;
  assign n23637 = n23376 | n23636 ;
  assign n23638 = n23362 & n23637 ;
  assign n23639 = n23360 | n23638 ;
  assign n23640 = n23347 & n23639 ;
  assign n23641 = n23345 | n23640 ;
  assign n23642 = n23320 & ~n23332 ;
  assign n23643 = ~n23320 & n23331 ;
  assign n23644 = n23642 | n23643 ;
  assign n23645 = n23641 & n23644 ;
  assign n23646 = n23332 | n23645 ;
  assign n23647 = n23307 & ~n23318 ;
  assign n23648 = ~n23307 & n23317 ;
  assign n23649 = n23647 | n23648 ;
  assign n23650 = n23646 & n23649 ;
  assign n23651 = n23293 | n23304 ;
  assign n23652 = ~n23305 & n23651 ;
  assign n23653 = ( n23318 & n23650 ) | ( n23318 & n23652 ) | ( n23650 & n23652 ) ;
  assign n23654 = n23305 | n23653 ;
  assign n23655 = n23291 & n23654 ;
  assign n23656 = n23288 | n23655 ;
  assign n23657 = n23273 & ~n23274 ;
  assign n23658 = ( n23263 & ~n23274 ) | ( n23263 & n23657 ) | ( ~n23274 & n23657 ) ;
  assign n23659 = n23656 & n23658 ;
  assign n23660 = n23274 | n23659 ;
  assign n23661 = ~n23027 & n23029 ;
  assign n23662 = n23030 | n23661 ;
  assign n23663 = ( n23260 & ~n23660 ) | ( n23260 & n23662 ) | ( ~n23660 & n23662 ) ;
  assign n23664 = ( ~n23260 & n23660 ) | ( ~n23260 & n23663 ) | ( n23660 & n23663 ) ;
  assign n23665 = ( ~n23662 & n23663 ) | ( ~n23662 & n23664 ) | ( n23663 & n23664 ) ;
  assign n23666 = ( n23260 & n23660 ) | ( n23260 & n23665 ) | ( n23660 & n23665 ) ;
  assign n23667 = n22668 & ~n23031 ;
  assign n23668 = n23032 | n23667 ;
  assign n23669 = ( n23249 & n23666 ) | ( n23249 & ~n23668 ) | ( n23666 & ~n23668 ) ;
  assign n23670 = ( n23225 & n23239 ) | ( n23225 & n23669 ) | ( n23239 & n23669 ) ;
  assign n23035 = n22649 | n23034 ;
  assign n21026 = n7305 & n20546 ;
  assign n21027 = n7300 & n20556 ;
  assign n21028 = n7302 & ~n20710 ;
  assign n21029 = n21027 | n21028 ;
  assign n21030 = n21026 | n21029 ;
  assign n21032 = n7308 & ~n21031 ;
  assign n21038 = ( n7308 & n21032 ) | ( n7308 & n21037 ) | ( n21032 & n21037 ) ;
  assign n21039 = n21030 | n21038 ;
  assign n21040 = x11 | n21039 ;
  assign n21041 = ~x11 & n21040 ;
  assign n21042 = ( ~n21039 & n21040 ) | ( ~n21039 & n21041 ) | ( n21040 & n21041 ) ;
  assign n22504 = n7280 & ~n20552 ;
  assign n22505 = n5384 & n20560 ;
  assign n22506 = n7277 & n20562 ;
  assign n22507 = n22505 | n22506 ;
  assign n22508 = n22504 | n22507 ;
  assign n22513 = n39 & ~n22512 ;
  assign n22514 = n22510 & n22513 ;
  assign n22515 = ( n39 & n22508 ) | ( n39 & ~n22514 ) | ( n22508 & ~n22514 ) ;
  assign n22516 = x14 & n22515 ;
  assign n22517 = x14 & ~n22516 ;
  assign n22518 = ( n22515 & ~n22516 ) | ( n22515 & n22517 ) | ( ~n22516 & n22517 ) ;
  assign n22519 = n5083 & ~n20689 ;
  assign n22520 = n5069 & ~n20569 ;
  assign n22521 = n5070 & ~n20573 ;
  assign n22522 = n22520 | n22521 ;
  assign n22523 = n22519 | n22522 ;
  assign n22524 = ( n5074 & ~n22192 ) | ( n5074 & n22193 ) | ( ~n22192 & n22193 ) ;
  assign n22525 = n22523 | n22524 ;
  assign n22526 = x17 | n22525 ;
  assign n22527 = ~x17 & n22526 ;
  assign n22528 = ( ~n22525 & n22526 ) | ( ~n22525 & n22527 ) | ( n22526 & n22527 ) ;
  assign n22529 = n4781 & ~n20584 ;
  assign n22530 = n4776 & n20588 ;
  assign n22531 = n4778 & ~n20580 ;
  assign n22532 = n22530 | n22531 ;
  assign n22533 = n22529 | n22532 ;
  assign n22534 = n4784 | n22533 ;
  assign n22535 = ( ~n21901 & n22533 ) | ( ~n21901 & n22534 ) | ( n22533 & n22534 ) ;
  assign n22536 = ~x20 & n22535 ;
  assign n22537 = x20 | n22536 ;
  assign n22538 = ( ~n22535 & n22536 ) | ( ~n22535 & n22537 ) | ( n22536 & n22537 ) ;
  assign n22539 = n21851 | n21855 ;
  assign n22540 = n4551 & ~n20591 ;
  assign n22541 = n4546 & n20600 ;
  assign n22542 = n4548 & ~n20595 ;
  assign n22543 = n22541 | n22542 ;
  assign n22544 = n22540 | n22543 ;
  assign n22545 = n4554 & n21539 ;
  assign n22546 = ( n4554 & n21543 ) | ( n4554 & n22545 ) | ( n21543 & n22545 ) ;
  assign n22547 = n22544 | n22546 ;
  assign n22548 = x23 | n22547 ;
  assign n22549 = ~x23 & n22548 ;
  assign n22550 = ( ~n22547 & n22548 ) | ( ~n22547 & n22549 ) | ( n22548 & n22549 ) ;
  assign n22551 = n4484 & ~n20605 ;
  assign n22552 = n4479 & n20614 ;
  assign n22553 = n4481 & n20611 ;
  assign n22554 = n22552 | n22553 ;
  assign n22555 = n22551 | n22554 ;
  assign n22556 = n4487 | n22555 ;
  assign n22557 = ( ~n21275 & n22555 ) | ( ~n21275 & n22556 ) | ( n22555 & n22556 ) ;
  assign n22558 = ~x26 & n22557 ;
  assign n22559 = x26 | n22558 ;
  assign n22560 = ( ~n22557 & n22558 ) | ( ~n22557 & n22559 ) | ( n22558 & n22559 ) ;
  assign n22561 = n21812 | n21815 ;
  assign n22562 = n21795 | n21800 ;
  assign n22563 = n4043 & n20622 ;
  assign n22564 = n4045 | n22563 ;
  assign n22565 = ( n20619 & n22563 ) | ( n20619 & n22564 ) | ( n22563 & n22564 ) ;
  assign n22566 = n4048 | n22565 ;
  assign n22567 = ( n20616 & n22565 ) | ( n20616 & n22566 ) | ( n22565 & n22566 ) ;
  assign n22568 = n4051 | n22567 ;
  assign n22569 = ( n21190 & n22567 ) | ( n21190 & n22568 ) | ( n22567 & n22568 ) ;
  assign n22570 = ~x29 & n22569 ;
  assign n22571 = x29 & ~n22569 ;
  assign n22572 = n22570 | n22571 ;
  assign n22573 = n3744 & ~n20625 ;
  assign n22574 = n3727 & ~n20630 ;
  assign n22575 = n3639 & n20633 ;
  assign n22576 = n22574 | n22575 ;
  assign n22577 = n22573 | n22576 ;
  assign n22578 = n3636 | n22577 ;
  assign n22579 = ( ~n21129 & n22577 ) | ( ~n21129 & n22578 ) | ( n22577 & n22578 ) ;
  assign n22580 = n19808 | n19830 ;
  assign n22581 = n1561 | n3809 ;
  assign n22582 = n4868 | n22581 ;
  assign n22583 = n687 | n1204 ;
  assign n22584 = ( ~n20758 & n22582 ) | ( ~n20758 & n22583 ) | ( n22582 & n22583 ) ;
  assign n22585 = n20758 | n22584 ;
  assign n22586 = n22580 | n22585 ;
  assign n22587 = n1865 | n22586 ;
  assign n22588 = n619 | n22587 ;
  assign n22589 = n14107 & ~n22588 ;
  assign n22590 = n591 | n626 ;
  assign n22591 = n435 | n22590 ;
  assign n22592 = n120 | n22591 ;
  assign n22593 = n22589 & ~n22592 ;
  assign n22594 = n22579 & ~n22593 ;
  assign n22595 = n22579 & ~n22594 ;
  assign n22596 = n22579 | n22593 ;
  assign n22597 = ( n21771 & n21772 ) | ( n21771 & n21791 ) | ( n21772 & n21791 ) ;
  assign n22598 = ( ~n22595 & n22596 ) | ( ~n22595 & n22597 ) | ( n22596 & n22597 ) ;
  assign n22599 = ( n22596 & n22597 ) | ( n22596 & ~n22598 ) | ( n22597 & ~n22598 ) ;
  assign n22600 = ( n22595 & n22598 ) | ( n22595 & ~n22599 ) | ( n22598 & ~n22599 ) ;
  assign n22601 = n22572 & ~n22600 ;
  assign n22602 = ~n22572 & n22600 ;
  assign n22603 = n22601 | n22602 ;
  assign n22604 = ~n22562 & n22603 ;
  assign n22605 = n22562 & ~n22603 ;
  assign n22606 = n22604 | n22605 ;
  assign n22607 = ( n22560 & n22561 ) | ( n22560 & ~n22606 ) | ( n22561 & ~n22606 ) ;
  assign n22608 = ( ~n22561 & n22606 ) | ( ~n22561 & n22607 ) | ( n22606 & n22607 ) ;
  assign n22609 = ( ~n22560 & n22607 ) | ( ~n22560 & n22608 ) | ( n22607 & n22608 ) ;
  assign n22610 = n22550 & ~n22609 ;
  assign n22611 = ~n22550 & n22609 ;
  assign n22612 = n22610 | n22611 ;
  assign n22613 = n21829 | n21835 ;
  assign n22614 = n22612 & ~n22613 ;
  assign n22615 = ~n22612 & n22613 ;
  assign n22616 = n22614 | n22615 ;
  assign n22617 = ( n22538 & n22539 ) | ( n22538 & ~n22616 ) | ( n22539 & ~n22616 ) ;
  assign n22618 = ( ~n22539 & n22616 ) | ( ~n22539 & n22617 ) | ( n22616 & n22617 ) ;
  assign n22619 = ( ~n22538 & n22617 ) | ( ~n22538 & n22618 ) | ( n22617 & n22618 ) ;
  assign n22620 = n22528 & ~n22619 ;
  assign n22621 = ~n22528 & n22619 ;
  assign n22622 = n22620 | n22621 ;
  assign n22623 = n21871 | n22165 ;
  assign n22624 = n22622 & ~n22623 ;
  assign n22625 = ~n22622 & n22623 ;
  assign n22626 = n22624 | n22625 ;
  assign n22627 = n22518 & ~n22626 ;
  assign n22628 = n22626 | n22627 ;
  assign n22629 = ( ~n22518 & n22627 ) | ( ~n22518 & n22628 ) | ( n22627 & n22628 ) ;
  assign n22630 = n22503 & ~n22629 ;
  assign n22631 = n22503 & ~n22630 ;
  assign n22632 = n22629 | n22630 ;
  assign n22633 = ~n22631 & n22632 ;
  assign n22634 = n21042 & ~n22633 ;
  assign n23036 = n22633 | n22634 ;
  assign n23037 = ( ~n21042 & n22634 ) | ( ~n21042 & n23036 ) | ( n22634 & n23036 ) ;
  assign n23038 = n23035 & ~n23037 ;
  assign n23671 = ~n23035 & n23037 ;
  assign n23672 = n23038 | n23671 ;
  assign n23673 = n23223 & ~n23672 ;
  assign n23674 = n23672 | n23673 ;
  assign n23675 = ( ~n23223 & n23673 ) | ( ~n23223 & n23674 ) | ( n23673 & n23674 ) ;
  assign n23676 = n23670 & n23675 ;
  assign n23677 = n23670 | n23675 ;
  assign n23678 = ~n23676 & n23677 ;
  assign n23679 = ( n23223 & n23670 ) | ( n23223 & n23678 ) | ( n23670 & n23678 ) ;
  assign n23039 = n22634 | n23038 ;
  assign n23043 = n7305 & ~n20542 ;
  assign n23044 = n7300 & ~n20710 ;
  assign n23045 = n7302 & n20546 ;
  assign n23046 = n23044 | n23045 ;
  assign n23047 = n23043 | n23046 ;
  assign n23048 = n7308 | n23047 ;
  assign n23049 = ( ~n23042 & n23047 ) | ( ~n23042 & n23048 ) | ( n23047 & n23048 ) ;
  assign n23050 = ~x11 & n23049 ;
  assign n23051 = x11 | n23050 ;
  assign n23052 = ( ~n23049 & n23050 ) | ( ~n23049 & n23051 ) | ( n23050 & n23051 ) ;
  assign n23053 = n22627 | n22630 ;
  assign n23054 = n7280 & n20556 ;
  assign n23055 = n5384 & n20562 ;
  assign n23056 = n7277 & ~n20552 ;
  assign n23057 = n23055 | n23056 ;
  assign n23058 = n23054 | n23057 ;
  assign n23059 = n39 | n23058 ;
  assign n23060 = ( ~n22655 & n23058 ) | ( ~n22655 & n23059 ) | ( n23058 & n23059 ) ;
  assign n23061 = ~x14 & n23060 ;
  assign n23062 = x14 | n23061 ;
  assign n23063 = ( ~n23060 & n23061 ) | ( ~n23060 & n23062 ) | ( n23061 & n23062 ) ;
  assign n23064 = n22620 | n22625 ;
  assign n23065 = n5083 & n20560 ;
  assign n23066 = n5069 & ~n20573 ;
  assign n23067 = n5070 & ~n20689 ;
  assign n23068 = n23066 | n23067 ;
  assign n23069 = n23065 | n23068 ;
  assign n23070 = ( n5074 & n22173 ) | ( n5074 & n22176 ) | ( n22173 & n22176 ) ;
  assign n23071 = n23069 | n23070 ;
  assign n23072 = x17 | n23071 ;
  assign n23073 = ~x17 & n23072 ;
  assign n23074 = ( ~n23071 & n23072 ) | ( ~n23071 & n23073 ) | ( n23072 & n23073 ) ;
  assign n23075 = n4781 & ~n20569 ;
  assign n23076 = n4776 & ~n20580 ;
  assign n23077 = n4778 & ~n20584 ;
  assign n23078 = n23076 | n23077 ;
  assign n23079 = n23075 | n23078 ;
  assign n23080 = n4784 & ~n21884 ;
  assign n23081 = n21889 & n23080 ;
  assign n23082 = ( n4784 & n23079 ) | ( n4784 & ~n23081 ) | ( n23079 & ~n23081 ) ;
  assign n23083 = x20 & n23082 ;
  assign n23084 = x20 & ~n23083 ;
  assign n23085 = ( n23082 & ~n23083 ) | ( n23082 & n23084 ) | ( ~n23083 & n23084 ) ;
  assign n23086 = n22610 | n22615 ;
  assign n23087 = n4551 & n20588 ;
  assign n23088 = n4546 & ~n20595 ;
  assign n23089 = n4548 & ~n20591 ;
  assign n23090 = n23088 | n23089 ;
  assign n23091 = n23087 | n23090 ;
  assign n23092 = n4554 | n23091 ;
  assign n23093 = ( n21526 & n23091 ) | ( n21526 & n23092 ) | ( n23091 & n23092 ) ;
  assign n23094 = x23 & n23093 ;
  assign n23095 = x23 & ~n23094 ;
  assign n23096 = ( n23093 & ~n23094 ) | ( n23093 & n23095 ) | ( ~n23094 & n23095 ) ;
  assign n23097 = n4484 & n20600 ;
  assign n23098 = n4479 & n20611 ;
  assign n23099 = n4481 & ~n20605 ;
  assign n23100 = n23098 | n23099 ;
  assign n23101 = n23097 | n23100 ;
  assign n23102 = n4487 | n23101 ;
  assign n23103 = ( ~n21432 & n23101 ) | ( ~n21432 & n23102 ) | ( n23101 & n23102 ) ;
  assign n23104 = ~x26 & n23103 ;
  assign n23105 = x26 | n23104 ;
  assign n23106 = ( ~n23103 & n23104 ) | ( ~n23103 & n23105 ) | ( n23104 & n23105 ) ;
  assign n23107 = n22601 | n22605 ;
  assign n23108 = n4048 & n20614 ;
  assign n23109 = n4043 & n20619 ;
  assign n23110 = n4045 | n23109 ;
  assign n23111 = ( n20616 & n23109 ) | ( n20616 & n23110 ) | ( n23109 & n23110 ) ;
  assign n23112 = n23108 | n23111 ;
  assign n23113 = n4051 | n23112 ;
  assign n23114 = ( n21302 & n23112 ) | ( n21302 & n23113 ) | ( n23112 & n23113 ) ;
  assign n23115 = ~x29 & n23114 ;
  assign n23116 = x29 & ~n23114 ;
  assign n23117 = n23115 | n23116 ;
  assign n23118 = ( n22594 & n22597 ) | ( n22594 & n22600 ) | ( n22597 & n22600 ) ;
  assign n23119 = n3744 & n20622 ;
  assign n23120 = n3727 & ~n20625 ;
  assign n23121 = n3639 & ~n20630 ;
  assign n23122 = n23120 | n23121 ;
  assign n23123 = n23119 | n23122 ;
  assign n23124 = n3636 | n23123 ;
  assign n23125 = ( n21114 & n23123 ) | ( n21114 & n23124 ) | ( n23123 & n23124 ) ;
  assign n23126 = n227 | n3845 ;
  assign n23127 = n3659 | n23126 ;
  assign n23128 = n1787 | n23127 ;
  assign n23129 = n710 | n23128 ;
  assign n23130 = n19678 & ~n23129 ;
  assign n23131 = ~n3801 & n23130 ;
  assign n23132 = ~n19631 & n23131 ;
  assign n23133 = n972 | n11368 ;
  assign n23134 = n1280 | n23133 ;
  assign n23135 = n1522 | n23134 ;
  assign n23136 = n718 | n23135 ;
  assign n23137 = n23132 & ~n23136 ;
  assign n23138 = n283 | n602 ;
  assign n23139 = n441 | n23138 ;
  assign n23140 = n206 | n23139 ;
  assign n23141 = n23137 & ~n23140 ;
  assign n23142 = n23125 & ~n23141 ;
  assign n23143 = n23125 & ~n23142 ;
  assign n23144 = n23125 | n23141 ;
  assign n23145 = ~n23143 & n23144 ;
  assign n23146 = n23118 & ~n23145 ;
  assign n23147 = n23118 & ~n23146 ;
  assign n23148 = n23145 | n23146 ;
  assign n23149 = ~n23147 & n23148 ;
  assign n23150 = n23117 & ~n23149 ;
  assign n23151 = ~n23117 & n23149 ;
  assign n23152 = n23150 | n23151 ;
  assign n23153 = ~n23107 & n23152 ;
  assign n23154 = n23107 & ~n23152 ;
  assign n23155 = n23153 | n23154 ;
  assign n23156 = n23106 & ~n23155 ;
  assign n23157 = n23155 | n23156 ;
  assign n23158 = ( ~n23106 & n23156 ) | ( ~n23106 & n23157 ) | ( n23156 & n23157 ) ;
  assign n23159 = n22607 & ~n23158 ;
  assign n23160 = n22607 & ~n23159 ;
  assign n23161 = n23158 | n23159 ;
  assign n23162 = ~n23160 & n23161 ;
  assign n23163 = n23096 & ~n23162 ;
  assign n23164 = n23162 | n23163 ;
  assign n23165 = ( ~n23096 & n23163 ) | ( ~n23096 & n23164 ) | ( n23163 & n23164 ) ;
  assign n23166 = ~n23086 & n23165 ;
  assign n23167 = n23086 & ~n23165 ;
  assign n23168 = n23166 | n23167 ;
  assign n23169 = n23085 & ~n23168 ;
  assign n23170 = n23168 | n23169 ;
  assign n23171 = ( ~n23085 & n23169 ) | ( ~n23085 & n23170 ) | ( n23169 & n23170 ) ;
  assign n23172 = n22617 & ~n23171 ;
  assign n23173 = n22617 & ~n23172 ;
  assign n23174 = n23171 | n23172 ;
  assign n23175 = ~n23173 & n23174 ;
  assign n23176 = n23074 & ~n23175 ;
  assign n23177 = n23175 | n23176 ;
  assign n23178 = ( ~n23074 & n23176 ) | ( ~n23074 & n23177 ) | ( n23176 & n23177 ) ;
  assign n23179 = ~n23064 & n23178 ;
  assign n23180 = n23064 & ~n23178 ;
  assign n23181 = n23179 | n23180 ;
  assign n23182 = n23063 & ~n23181 ;
  assign n23183 = n23181 | n23182 ;
  assign n23184 = ( ~n23063 & n23182 ) | ( ~n23063 & n23183 ) | ( n23182 & n23183 ) ;
  assign n23185 = n23053 & ~n23184 ;
  assign n23186 = n23053 & ~n23185 ;
  assign n23187 = n23184 | n23185 ;
  assign n23188 = ~n23186 & n23187 ;
  assign n23189 = n23052 & ~n23188 ;
  assign n23190 = n23188 | n23189 ;
  assign n23191 = ( ~n23052 & n23189 ) | ( ~n23052 & n23190 ) | ( n23189 & n23190 ) ;
  assign n23192 = ~n23039 & n23191 ;
  assign n23193 = n23039 & ~n23191 ;
  assign n23194 = n23192 | n23193 ;
  assign n23195 = n5503 & n20532 ;
  assign n23196 = n5512 & ~n20724 ;
  assign n23197 = n5508 & ~n20536 ;
  assign n23198 = n23196 | n23197 ;
  assign n23199 = n23195 | n23198 ;
  assign n23200 = n5515 | n23199 ;
  assign n23201 = n20537 | n20538 ;
  assign n23202 = n20733 & n23201 ;
  assign n23203 = n20735 & ~n23202 ;
  assign n23204 = ( n23199 & n23200 ) | ( n23199 & n23203 ) | ( n23200 & n23203 ) ;
  assign n23205 = x8 & n23204 ;
  assign n23206 = x8 & ~n23205 ;
  assign n23207 = ( n23204 & ~n23205 ) | ( n23204 & n23206 ) | ( ~n23205 & n23206 ) ;
  assign n23680 = ( n23194 & ~n23207 ) | ( n23194 & n23679 ) | ( ~n23207 & n23679 ) ;
  assign n23681 = ( ~n23194 & n23207 ) | ( ~n23194 & n23680 ) | ( n23207 & n23680 ) ;
  assign n23682 = ( ~n23679 & n23680 ) | ( ~n23679 & n23681 ) | ( n23680 & n23681 ) ;
  assign n23683 = n21025 & ~n23682 ;
  assign n23684 = ~n21025 & n23682 ;
  assign n23685 = n23683 | n23684 ;
  assign n23686 = n9245 & n20921 ;
  assign n23687 = n8680 & n20532 ;
  assign n23688 = n8681 & n20838 ;
  assign n23689 = n23687 | n23688 ;
  assign n23690 = n23686 | n23689 ;
  assign n23691 = n20922 & ~n20929 ;
  assign n23692 = n20838 & n20921 ;
  assign n23693 = n20923 & ~n23692 ;
  assign n23694 = ( ~n20735 & n20839 ) | ( ~n20735 & n20927 ) | ( n20839 & n20927 ) ;
  assign n23695 = ~n23693 & n23694 ;
  assign n23696 = ( n8685 & n23691 ) | ( n8685 & n23695 ) | ( n23691 & n23695 ) ;
  assign n23697 = n23690 | n23696 ;
  assign n23698 = x5 | n23697 ;
  assign n23699 = ~x5 & n23698 ;
  assign n23700 = ( ~n23697 & n23698 ) | ( ~n23697 & n23699 ) | ( n23698 & n23699 ) ;
  assign n23701 = ~n23678 & n23700 ;
  assign n23702 = n23678 & ~n23700 ;
  assign n23703 = n23701 | n23702 ;
  assign n23704 = n9245 & n20838 ;
  assign n23705 = n8680 & ~n20536 ;
  assign n23706 = n8681 & n20532 ;
  assign n23707 = n23705 | n23706 ;
  assign n23708 = n23704 | n23707 ;
  assign n23709 = ( ~n20735 & n20925 ) | ( ~n20735 & n20926 ) | ( n20925 & n20926 ) ;
  assign n23710 = n20537 | n20925 ;
  assign n23711 = n20735 & ~n23710 ;
  assign n23712 = n23709 | n23711 ;
  assign n23713 = n8685 | n23708 ;
  assign n23714 = ( n23708 & ~n23712 ) | ( n23708 & n23713 ) | ( ~n23712 & n23713 ) ;
  assign n23715 = ~x5 & n23714 ;
  assign n23716 = x5 | n23715 ;
  assign n23717 = ( ~n23714 & n23715 ) | ( ~n23714 & n23716 ) | ( n23715 & n23716 ) ;
  assign n23718 = ( n23225 & n23669 ) | ( n23225 & ~n23670 ) | ( n23669 & ~n23670 ) ;
  assign n23719 = ( n23239 & ~n23670 ) | ( n23239 & n23718 ) | ( ~n23670 & n23718 ) ;
  assign n23720 = ( ~n23249 & n23668 ) | ( ~n23249 & n23669 ) | ( n23668 & n23669 ) ;
  assign n23721 = ( ~n23666 & n23669 ) | ( ~n23666 & n23720 ) | ( n23669 & n23720 ) ;
  assign n23722 = n9245 & n20532 ;
  assign n23723 = n8680 & ~n20724 ;
  assign n23724 = n8681 & ~n20536 ;
  assign n23725 = n23723 | n23724 ;
  assign n23726 = n23722 | n23725 ;
  assign n23727 = n8685 | n23726 ;
  assign n23728 = ( n23203 & n23726 ) | ( n23203 & n23727 ) | ( n23726 & n23727 ) ;
  assign n23729 = x5 & n23728 ;
  assign n23730 = x5 & ~n23729 ;
  assign n23731 = ( n23728 & ~n23729 ) | ( n23728 & n23730 ) | ( ~n23729 & n23730 ) ;
  assign n23732 = n9245 & ~n20536 ;
  assign n23733 = n8680 & ~n20542 ;
  assign n23734 = n8681 & ~n20724 ;
  assign n23735 = n23733 | n23734 ;
  assign n23736 = n23732 | n23735 ;
  assign n23737 = ( n8685 & n23213 ) | ( n8685 & ~n23217 ) | ( n23213 & ~n23217 ) ;
  assign n23738 = n23736 | n23737 ;
  assign n23739 = x5 | n23738 ;
  assign n23740 = ~x5 & n23739 ;
  assign n23741 = ( ~n23738 & n23739 ) | ( ~n23738 & n23740 ) | ( n23739 & n23740 ) ;
  assign n23742 = n23656 | n23658 ;
  assign n23743 = ~n23659 & n23742 ;
  assign n23744 = n9245 & ~n20724 ;
  assign n23745 = n8680 & n20546 ;
  assign n23746 = n8681 & ~n20542 ;
  assign n23747 = n23745 | n23746 ;
  assign n23748 = n23744 | n23747 ;
  assign n23749 = n8685 | n23748 ;
  assign n23750 = ( n23229 & n23748 ) | ( n23229 & n23749 ) | ( n23748 & n23749 ) ;
  assign n23751 = x5 & n23750 ;
  assign n23752 = x5 & ~n23751 ;
  assign n23753 = ( n23750 & ~n23751 ) | ( n23750 & n23752 ) | ( ~n23751 & n23752 ) ;
  assign n23754 = n23743 & n23753 ;
  assign n23755 = n23743 | n23753 ;
  assign n23756 = ~n23754 & n23755 ;
  assign n23757 = n23291 | n23654 ;
  assign n23758 = ~n23655 & n23757 ;
  assign n23759 = n9245 & ~n20542 ;
  assign n23760 = n8680 & ~n20710 ;
  assign n23761 = n8681 & n20546 ;
  assign n23762 = n23760 | n23761 ;
  assign n23763 = n23759 | n23762 ;
  assign n23764 = n8685 | n23763 ;
  assign n23765 = ( ~n23042 & n23763 ) | ( ~n23042 & n23764 ) | ( n23763 & n23764 ) ;
  assign n23766 = ~x5 & n23765 ;
  assign n23767 = x5 | n23766 ;
  assign n23768 = ( ~n23765 & n23766 ) | ( ~n23765 & n23767 ) | ( n23766 & n23767 ) ;
  assign n23769 = n23318 | n23652 ;
  assign n23770 = n23650 | n23769 ;
  assign n23771 = ~n23653 & n23770 ;
  assign n23772 = n9245 & n20546 ;
  assign n23773 = n8680 & n20556 ;
  assign n23774 = n8681 & ~n20710 ;
  assign n23775 = n23773 | n23774 ;
  assign n23776 = n23772 | n23775 ;
  assign n23777 = n8685 & ~n21031 ;
  assign n23778 = ( n8685 & n21037 ) | ( n8685 & n23777 ) | ( n21037 & n23777 ) ;
  assign n23779 = n23776 | n23778 ;
  assign n23780 = x5 | n23779 ;
  assign n23781 = ~x5 & n23780 ;
  assign n23782 = ( ~n23779 & n23780 ) | ( ~n23779 & n23781 ) | ( n23780 & n23781 ) ;
  assign n23783 = n23646 & ~n23650 ;
  assign n23784 = n23649 & ~n23650 ;
  assign n23785 = n23783 | n23784 ;
  assign n23786 = n9245 & ~n20710 ;
  assign n23787 = n8680 & ~n20552 ;
  assign n23788 = n8681 & n20556 ;
  assign n23789 = n23787 | n23788 ;
  assign n23790 = n23786 | n23789 ;
  assign n23791 = n8685 | n23790 ;
  assign n23792 = ( ~n22641 & n23790 ) | ( ~n22641 & n23791 ) | ( n23790 & n23791 ) ;
  assign n23793 = ~x5 & n23792 ;
  assign n23794 = x5 | n23793 ;
  assign n23795 = ( ~n23792 & n23793 ) | ( ~n23792 & n23794 ) | ( n23793 & n23794 ) ;
  assign n23796 = n23641 & ~n23645 ;
  assign n23797 = n23644 & ~n23645 ;
  assign n23798 = n23796 | n23797 ;
  assign n23799 = n9245 & n20556 ;
  assign n23800 = n8680 & n20562 ;
  assign n23801 = n8681 & ~n20552 ;
  assign n23802 = n23800 | n23801 ;
  assign n23803 = n23799 | n23802 ;
  assign n23804 = n8685 | n23803 ;
  assign n23805 = ( ~n22655 & n23803 ) | ( ~n22655 & n23804 ) | ( n23803 & n23804 ) ;
  assign n23806 = ~x5 & n23805 ;
  assign n23807 = x5 | n23806 ;
  assign n23808 = ( ~n23805 & n23806 ) | ( ~n23805 & n23807 ) | ( n23806 & n23807 ) ;
  assign n23809 = n23347 | n23639 ;
  assign n23810 = ~n23640 & n23809 ;
  assign n23811 = n9245 & ~n20552 ;
  assign n23812 = n8680 & n20560 ;
  assign n23813 = n8681 & n20562 ;
  assign n23814 = n23812 | n23813 ;
  assign n23815 = n23811 | n23814 ;
  assign n23816 = n8685 & n22510 ;
  assign n23817 = ~n22512 & n23816 ;
  assign n23818 = ( n8685 & n23815 ) | ( n8685 & ~n23817 ) | ( n23815 & ~n23817 ) ;
  assign n23819 = x5 & n23818 ;
  assign n23820 = x5 & ~n23819 ;
  assign n23821 = ( n23818 & ~n23819 ) | ( n23818 & n23820 ) | ( ~n23819 & n23820 ) ;
  assign n23822 = n23810 & n23821 ;
  assign n23823 = n23362 | n23637 ;
  assign n23824 = ~n23638 & n23823 ;
  assign n23825 = n9245 & n20562 ;
  assign n23826 = n8680 & ~n20689 ;
  assign n23827 = n8681 & n20560 ;
  assign n23828 = n23826 | n23827 ;
  assign n23829 = n23825 | n23828 ;
  assign n23830 = n8685 | n23829 ;
  assign n23831 = ( ~n21044 & n23829 ) | ( ~n21044 & n23830 ) | ( n23829 & n23830 ) ;
  assign n23832 = ~x5 & n23831 ;
  assign n23833 = x5 | n23832 ;
  assign n23834 = ( ~n23831 & n23832 ) | ( ~n23831 & n23833 ) | ( n23832 & n23833 ) ;
  assign n23835 = n23824 & n23834 ;
  assign n23836 = n23810 | n23821 ;
  assign n23837 = ~n23822 & n23836 ;
  assign n23838 = n23378 | n23635 ;
  assign n23839 = ~n23636 & n23838 ;
  assign n23840 = n9245 & n20560 ;
  assign n23841 = n8680 & ~n20573 ;
  assign n23842 = n8681 & ~n20689 ;
  assign n23843 = n23841 | n23842 ;
  assign n23844 = n23840 | n23843 ;
  assign n23845 = n8685 & ~n22176 ;
  assign n23846 = ~n22173 & n23845 ;
  assign n23847 = ( n8685 & n23844 ) | ( n8685 & ~n23846 ) | ( n23844 & ~n23846 ) ;
  assign n23848 = ~x5 & n23847 ;
  assign n23849 = x5 | n23848 ;
  assign n23850 = ( ~n23847 & n23848 ) | ( ~n23847 & n23849 ) | ( n23848 & n23849 ) ;
  assign n23851 = n23839 & n23850 ;
  assign n23852 = n23393 | n23633 ;
  assign n23853 = ~n23634 & n23852 ;
  assign n23854 = n9245 & ~n20689 ;
  assign n23855 = n8680 & ~n20569 ;
  assign n23856 = n8681 & ~n20573 ;
  assign n23857 = n23855 | n23856 ;
  assign n23858 = n23854 | n23857 ;
  assign n23859 = ( n8685 & ~n22192 ) | ( n8685 & n22193 ) | ( ~n22192 & n22193 ) ;
  assign n23860 = n23858 | n23859 ;
  assign n23861 = x5 | n23860 ;
  assign n23862 = ~x5 & n23861 ;
  assign n23863 = ( ~n23860 & n23861 ) | ( ~n23860 & n23862 ) | ( n23861 & n23862 ) ;
  assign n23864 = n23853 & n23863 ;
  assign n23865 = n23863 & ~n23864 ;
  assign n23866 = ( n23853 & ~n23864 ) | ( n23853 & n23865 ) | ( ~n23864 & n23865 ) ;
  assign n23867 = n9245 & ~n20573 ;
  assign n23868 = n8680 & ~n20584 ;
  assign n23869 = n8681 & ~n20569 ;
  assign n23870 = n23868 | n23869 ;
  assign n23871 = n23867 | n23870 ;
  assign n23872 = n8685 | n23871 ;
  assign n23873 = ( ~n21860 & n23871 ) | ( ~n21860 & n23872 ) | ( n23871 & n23872 ) ;
  assign n23874 = ~x5 & n23873 ;
  assign n23875 = x5 | n23874 ;
  assign n23876 = ( ~n23873 & n23874 ) | ( ~n23873 & n23875 ) | ( n23874 & n23875 ) ;
  assign n23877 = n9245 & ~n20569 ;
  assign n23878 = n8680 & ~n20580 ;
  assign n23879 = n8681 & ~n20584 ;
  assign n23880 = n23878 | n23879 ;
  assign n23881 = n23877 | n23880 ;
  assign n23882 = n8685 & n21884 ;
  assign n23883 = ( n8685 & ~n21889 ) | ( n8685 & n23882 ) | ( ~n21889 & n23882 ) ;
  assign n23884 = n23881 | n23883 ;
  assign n23885 = x5 | n23884 ;
  assign n23886 = ~x5 & n23885 ;
  assign n23887 = ( ~n23884 & n23885 ) | ( ~n23884 & n23886 ) | ( n23885 & n23886 ) ;
  assign n23888 = n23627 | n23629 ;
  assign n23889 = ~n23630 & n23888 ;
  assign n23890 = n9245 & ~n20584 ;
  assign n23891 = n8680 & n20588 ;
  assign n23892 = n8681 & ~n20580 ;
  assign n23893 = n23891 | n23892 ;
  assign n23894 = n23890 | n23893 ;
  assign n23895 = n8685 | n23894 ;
  assign n23896 = ( ~n21901 & n23894 ) | ( ~n21901 & n23895 ) | ( n23894 & n23895 ) ;
  assign n23897 = ~x5 & n23896 ;
  assign n23898 = x5 | n23897 ;
  assign n23899 = ( ~n23896 & n23897 ) | ( ~n23896 & n23898 ) | ( n23897 & n23898 ) ;
  assign n23900 = n23889 & n23899 ;
  assign n23901 = n23889 | n23899 ;
  assign n23902 = ~n23900 & n23901 ;
  assign n23903 = n23449 | n23625 ;
  assign n23904 = ~n23626 & n23903 ;
  assign n23905 = n9245 & ~n20580 ;
  assign n23906 = n8680 & ~n20591 ;
  assign n23907 = n8681 & n20588 ;
  assign n23908 = n23906 | n23907 ;
  assign n23909 = n23905 | n23908 ;
  assign n23910 = n8685 | n23909 ;
  assign n23911 = ( n21840 & n23909 ) | ( n21840 & n23910 ) | ( n23909 & n23910 ) ;
  assign n23912 = x5 & n23911 ;
  assign n23913 = x5 & ~n23912 ;
  assign n23914 = ( n23911 & ~n23912 ) | ( n23911 & n23913 ) | ( ~n23912 & n23913 ) ;
  assign n23915 = n23466 | n23623 ;
  assign n23916 = ~n23624 & n23915 ;
  assign n23917 = n9245 & n20588 ;
  assign n23918 = n8680 & ~n20595 ;
  assign n23919 = n8681 & ~n20591 ;
  assign n23920 = n23918 | n23919 ;
  assign n23921 = n23917 | n23920 ;
  assign n23922 = n8685 | n23921 ;
  assign n23923 = ( n21526 & n23921 ) | ( n21526 & n23922 ) | ( n23921 & n23922 ) ;
  assign n23924 = x5 & n23923 ;
  assign n23925 = x5 & ~n23924 ;
  assign n23926 = ( n23923 & ~n23924 ) | ( n23923 & n23925 ) | ( ~n23924 & n23925 ) ;
  assign n23927 = n23492 | n23621 ;
  assign n23928 = n23619 | n23927 ;
  assign n23929 = ~n23622 & n23928 ;
  assign n23930 = n9245 & ~n20591 ;
  assign n23931 = n8680 & n20600 ;
  assign n23932 = n8681 & ~n20595 ;
  assign n23933 = n23931 | n23932 ;
  assign n23934 = n23930 | n23933 ;
  assign n23935 = n8685 & n21539 ;
  assign n23936 = ( n8685 & n21543 ) | ( n8685 & n23935 ) | ( n21543 & n23935 ) ;
  assign n23937 = n23934 | n23936 ;
  assign n23938 = x5 | n23937 ;
  assign n23939 = ~x5 & n23938 ;
  assign n23940 = ( ~n23937 & n23938 ) | ( ~n23937 & n23939 ) | ( n23938 & n23939 ) ;
  assign n23941 = n23616 & ~n23619 ;
  assign n23942 = n23618 & ~n23619 ;
  assign n23943 = n23941 | n23942 ;
  assign n23944 = n9245 & ~n20595 ;
  assign n23945 = n8680 & ~n20605 ;
  assign n23946 = n8681 & n20600 ;
  assign n23947 = n23945 | n23946 ;
  assign n23948 = n23944 | n23947 ;
  assign n23949 = n8685 | n23948 ;
  assign n23950 = ( ~n21554 & n23948 ) | ( ~n21554 & n23949 ) | ( n23948 & n23949 ) ;
  assign n23951 = ~x5 & n23950 ;
  assign n23952 = x5 | n23951 ;
  assign n23953 = ( ~n23950 & n23951 ) | ( ~n23950 & n23952 ) | ( n23951 & n23952 ) ;
  assign n23954 = n23611 & ~n23615 ;
  assign n23955 = n23614 & ~n23615 ;
  assign n23956 = n23954 | n23955 ;
  assign n23957 = n9245 & n20600 ;
  assign n23958 = n8680 & n20611 ;
  assign n23959 = n8681 & ~n20605 ;
  assign n23960 = n23958 | n23959 ;
  assign n23961 = n23957 | n23960 ;
  assign n23962 = n8685 | n23961 ;
  assign n23963 = ( ~n21432 & n23961 ) | ( ~n21432 & n23962 ) | ( n23961 & n23962 ) ;
  assign n23964 = ~x5 & n23963 ;
  assign n23965 = x5 | n23964 ;
  assign n23966 = ( ~n23963 & n23964 ) | ( ~n23963 & n23965 ) | ( n23964 & n23965 ) ;
  assign n23967 = n23607 | n23609 ;
  assign n23968 = ~n23610 & n23967 ;
  assign n23969 = n9245 & ~n20605 ;
  assign n23970 = n8680 & n20614 ;
  assign n23971 = n8681 & n20611 ;
  assign n23972 = n23970 | n23971 ;
  assign n23973 = n23969 | n23972 ;
  assign n23974 = n8685 | n23973 ;
  assign n23975 = ( ~n21275 & n23973 ) | ( ~n21275 & n23974 ) | ( n23973 & n23974 ) ;
  assign n23976 = ~x5 & n23975 ;
  assign n23977 = x5 | n23976 ;
  assign n23978 = ( ~n23975 & n23976 ) | ( ~n23975 & n23977 ) | ( n23976 & n23977 ) ;
  assign n23979 = n23968 & n23978 ;
  assign n23980 = n23533 | n23605 ;
  assign n23981 = ~n23606 & n23980 ;
  assign n23982 = n9245 & n20611 ;
  assign n23983 = n8680 & n20616 ;
  assign n23984 = n8681 & n20614 ;
  assign n23985 = n23983 | n23984 ;
  assign n23986 = n23982 | n23985 ;
  assign n23987 = n8685 | n23986 ;
  assign n23988 = ( n21293 & n23986 ) | ( n21293 & n23987 ) | ( n23986 & n23987 ) ;
  assign n23989 = x5 & n23988 ;
  assign n23990 = x5 & ~n23989 ;
  assign n23991 = ( n23988 & ~n23989 ) | ( n23988 & n23990 ) | ( ~n23989 & n23990 ) ;
  assign n23992 = n23981 & n23991 ;
  assign n23993 = n23601 | n23603 ;
  assign n23994 = ~n23604 & n23993 ;
  assign n23995 = n9245 & n20614 ;
  assign n23996 = n8680 & n20619 ;
  assign n23997 = n8681 | n23996 ;
  assign n23998 = ( n20616 & n23996 ) | ( n20616 & n23997 ) | ( n23996 & n23997 ) ;
  assign n23999 = n23995 | n23998 ;
  assign n24000 = n8685 | n23999 ;
  assign n24001 = ( n21302 & n23999 ) | ( n21302 & n24000 ) | ( n23999 & n24000 ) ;
  assign n24002 = x5 & n24001 ;
  assign n24003 = x5 & ~n24002 ;
  assign n24004 = ( n24001 & ~n24002 ) | ( n24001 & n24003 ) | ( ~n24002 & n24003 ) ;
  assign n24005 = n23994 & n24004 ;
  assign n24006 = n8680 & n20622 ;
  assign n24007 = n8681 | n24006 ;
  assign n24008 = ( n20619 & n24006 ) | ( n20619 & n24007 ) | ( n24006 & n24007 ) ;
  assign n24009 = n9245 | n24008 ;
  assign n24010 = ( n20616 & n24008 ) | ( n20616 & n24009 ) | ( n24008 & n24009 ) ;
  assign n24011 = n8685 | n24010 ;
  assign n24012 = ( n21190 & n24010 ) | ( n21190 & n24011 ) | ( n24010 & n24011 ) ;
  assign n24013 = ~x5 & n24012 ;
  assign n24014 = x5 & ~n24012 ;
  assign n24015 = n24013 | n24014 ;
  assign n24016 = n23561 | n23599 ;
  assign n24017 = ~n23600 & n24016 ;
  assign n24018 = n24015 & n24017 ;
  assign n24019 = n8680 & ~n20625 ;
  assign n24020 = n8681 | n24019 ;
  assign n24021 = ( n20622 & n24019 ) | ( n20622 & n24020 ) | ( n24019 & n24020 ) ;
  assign n24022 = n9245 | n24021 ;
  assign n24023 = ( n20619 & n24021 ) | ( n20619 & n24022 ) | ( n24021 & n24022 ) ;
  assign n24024 = n8685 | n24023 ;
  assign n24025 = ( ~n21056 & n24023 ) | ( ~n21056 & n24024 ) | ( n24023 & n24024 ) ;
  assign n24026 = ~x5 & n24025 ;
  assign n24027 = x5 | n24026 ;
  assign n24028 = ( ~n24025 & n24026 ) | ( ~n24025 & n24027 ) | ( n24026 & n24027 ) ;
  assign n24029 = n23587 & ~n23598 ;
  assign n24030 = ( n23597 & ~n23598 ) | ( n23597 & n24029 ) | ( ~n23598 & n24029 ) ;
  assign n24031 = n24028 & n24030 ;
  assign n24032 = n24028 | n24030 ;
  assign n24033 = ~n24031 & n24032 ;
  assign n24034 = n23571 | n23582 ;
  assign n24035 = ~n23585 & n24034 ;
  assign n24036 = n9245 & n20622 ;
  assign n24037 = n8680 & ~n20630 ;
  assign n24038 = n8681 & ~n20625 ;
  assign n24039 = n24037 | n24038 ;
  assign n24040 = n24036 | n24039 ;
  assign n24041 = n8685 | n24040 ;
  assign n24042 = ( n21114 & n24040 ) | ( n21114 & n24041 ) | ( n24040 & n24041 ) ;
  assign n24043 = x5 & n24042 ;
  assign n24044 = x5 | n24042 ;
  assign n24045 = ~n24043 & n24044 ;
  assign n24046 = n23562 | n23570 ;
  assign n24047 = ~n23571 & n24046 ;
  assign n24048 = n9245 & ~n20625 ;
  assign n24049 = n8680 & n20633 ;
  assign n24050 = n8681 & ~n20630 ;
  assign n24051 = n24049 | n24050 ;
  assign n24052 = n24048 | n24051 ;
  assign n24053 = n8685 | n24052 ;
  assign n24054 = ( ~n21129 & n24052 ) | ( ~n21129 & n24053 ) | ( n24052 & n24053 ) ;
  assign n24055 = ~x5 & n24054 ;
  assign n24056 = x5 | n24055 ;
  assign n24057 = ( ~n24054 & n24055 ) | ( ~n24054 & n24056 ) | ( n24055 & n24056 ) ;
  assign n24058 = n24047 & n24057 ;
  assign n24059 = n24047 | n24057 ;
  assign n24060 = ~n24058 & n24059 ;
  assign n24061 = n5502 & ~n20642 ;
  assign n24062 = ( x5 & n18451 ) | ( x5 & n20642 ) | ( n18451 & n20642 ) ;
  assign n24063 = n8685 & n21069 ;
  assign n24064 = n8681 & ~n20642 ;
  assign n24065 = n9245 & ~n20640 ;
  assign n24066 = n24064 | n24065 ;
  assign n24067 = n24063 | n24066 ;
  assign n24068 = x5 | n24067 ;
  assign n24069 = ~x5 & n24068 ;
  assign n24070 = ( ~n24067 & n24068 ) | ( ~n24067 & n24069 ) | ( n24068 & n24069 ) ;
  assign n24071 = n24062 & n24070 ;
  assign n24072 = n9245 & n20633 ;
  assign n24073 = n8680 & ~n20642 ;
  assign n24074 = n8681 & ~n20640 ;
  assign n24075 = n24073 | n24074 ;
  assign n24076 = n24072 | n24075 ;
  assign n24077 = n8685 & n21085 ;
  assign n24078 = n24076 | n24077 ;
  assign n24079 = ~x5 & n24078 ;
  assign n24080 = x5 | n24079 ;
  assign n24081 = ( ~n24078 & n24079 ) | ( ~n24078 & n24080 ) | ( n24079 & n24080 ) ;
  assign n24082 = n24071 & n24081 ;
  assign n24083 = n9245 & ~n20630 ;
  assign n24084 = n8680 & ~n20640 ;
  assign n24085 = n8681 & n20633 ;
  assign n24086 = n24084 | n24085 ;
  assign n24087 = n24083 | n24086 ;
  assign n24088 = n8685 | n24087 ;
  assign n24089 = ( n21099 & n24087 ) | ( n21099 & n24088 ) | ( n24087 & n24088 ) ;
  assign n24090 = x5 & n24089 ;
  assign n24091 = x5 | n24089 ;
  assign n24092 = ~n24090 & n24091 ;
  assign n24093 = ( n24061 & n24082 ) | ( n24061 & n24092 ) | ( n24082 & n24092 ) ;
  assign n24094 = n24060 & n24093 ;
  assign n24095 = n24058 | n24094 ;
  assign n24096 = ( n24035 & n24045 ) | ( n24035 & n24095 ) | ( n24045 & n24095 ) ;
  assign n24097 = n24033 & n24096 ;
  assign n24098 = n24031 | n24097 ;
  assign n24099 = n24015 | n24017 ;
  assign n24100 = ~n24018 & n24099 ;
  assign n24101 = n24098 & n24100 ;
  assign n24102 = n24018 | n24101 ;
  assign n24103 = n23994 & ~n24005 ;
  assign n24104 = n24004 & ~n24005 ;
  assign n24105 = n24103 | n24104 ;
  assign n24106 = n24102 & n24105 ;
  assign n24107 = n24005 | n24106 ;
  assign n24108 = n23991 & ~n23992 ;
  assign n24109 = ( n23981 & ~n23992 ) | ( n23981 & n24108 ) | ( ~n23992 & n24108 ) ;
  assign n24110 = n24107 & n24109 ;
  assign n24111 = n23968 | n23978 ;
  assign n24112 = ~n23979 & n24111 ;
  assign n24113 = ( n23992 & n24110 ) | ( n23992 & n24112 ) | ( n24110 & n24112 ) ;
  assign n24114 = n23979 | n24113 ;
  assign n24115 = ( n23956 & n23966 ) | ( n23956 & n24114 ) | ( n23966 & n24114 ) ;
  assign n24116 = ( n23943 & n23953 ) | ( n23943 & n24115 ) | ( n23953 & n24115 ) ;
  assign n24117 = ( n23929 & n23940 ) | ( n23929 & n24116 ) | ( n23940 & n24116 ) ;
  assign n24118 = ( n23916 & n23926 ) | ( n23916 & n24117 ) | ( n23926 & n24117 ) ;
  assign n24119 = ( n23904 & n23914 ) | ( n23904 & n24118 ) | ( n23914 & n24118 ) ;
  assign n24120 = n23902 & n24119 ;
  assign n24121 = n23900 | n24120 ;
  assign n24122 = ( n23407 & n23631 ) | ( n23407 & ~n23632 ) | ( n23631 & ~n23632 ) ;
  assign n24123 = ( n23417 & ~n23632 ) | ( n23417 & n24122 ) | ( ~n23632 & n24122 ) ;
  assign n24124 = ( n23887 & n24121 ) | ( n23887 & n24123 ) | ( n24121 & n24123 ) ;
  assign n24125 = ( n23395 & n23632 ) | ( n23395 & ~n23633 ) | ( n23632 & ~n23633 ) ;
  assign n24126 = ( n23405 & ~n23633 ) | ( n23405 & n24125 ) | ( ~n23633 & n24125 ) ;
  assign n24127 = ( n23876 & n24124 ) | ( n23876 & n24126 ) | ( n24124 & n24126 ) ;
  assign n24128 = n23866 & n24127 ;
  assign n24129 = n23864 | n24128 ;
  assign n24130 = n23839 & ~n23851 ;
  assign n24131 = ~n23839 & n23850 ;
  assign n24132 = ( n24129 & n24130 ) | ( n24129 & n24131 ) | ( n24130 & n24131 ) ;
  assign n24133 = n23851 | n24132 ;
  assign n24134 = n23824 & ~n23835 ;
  assign n24135 = ~n23824 & n23834 ;
  assign n24136 = ( n24133 & n24134 ) | ( n24133 & n24135 ) | ( n24134 & n24135 ) ;
  assign n24137 = ( n23835 & n23837 ) | ( n23835 & n24136 ) | ( n23837 & n24136 ) ;
  assign n24138 = n23822 | n24137 ;
  assign n24139 = ( n23798 & n23808 ) | ( n23798 & n24138 ) | ( n23808 & n24138 ) ;
  assign n24140 = ( n23785 & n23795 ) | ( n23785 & n24139 ) | ( n23795 & n24139 ) ;
  assign n24141 = ( n23771 & n23782 ) | ( n23771 & n24140 ) | ( n23782 & n24140 ) ;
  assign n24142 = ( n23758 & n23768 ) | ( n23758 & n24141 ) | ( n23768 & n24141 ) ;
  assign n24143 = n23756 & n24142 ;
  assign n24144 = n23754 | n24143 ;
  assign n24145 = ( ~n23665 & n23741 ) | ( ~n23665 & n24144 ) | ( n23741 & n24144 ) ;
  assign n24146 = ( ~n23721 & n23731 ) | ( ~n23721 & n24145 ) | ( n23731 & n24145 ) ;
  assign n24147 = ( n23717 & n23719 ) | ( n23717 & n24146 ) | ( n23719 & n24146 ) ;
  assign n24148 = ~n23703 & n24147 ;
  assign n24149 = n23701 | n24148 ;
  assign n24150 = n23685 & ~n24149 ;
  assign n24151 = ~n23685 & n24149 ;
  assign n24152 = n24150 | n24151 ;
  assign n24153 = n3744 & ~n12328 ;
  assign n24154 = n3639 & ~n12335 ;
  assign n24155 = n3727 & ~n12325 ;
  assign n24156 = n24154 | n24155 ;
  assign n24157 = n24153 | n24156 ;
  assign n24158 = n3636 | n24157 ;
  assign n24159 = ( ~n13544 & n24157 ) | ( ~n13544 & n24158 ) | ( n24157 & n24158 ) ;
  assign n24160 = n574 | n2722 ;
  assign n24161 = n342 & ~n24160 ;
  assign n24162 = n227 | n586 ;
  assign n24163 = n670 | n24162 ;
  assign n24164 = n665 | n24163 ;
  assign n24165 = n669 | n24164 ;
  assign n24166 = n55 | n24165 ;
  assign n24167 = n24161 & ~n24166 ;
  assign n24168 = n20958 | n24167 ;
  assign n24169 = n20958 & n24167 ;
  assign n24170 = n24168 & ~n24169 ;
  assign n24171 = n4481 | n4484 ;
  assign n24172 = n4479 | n24171 ;
  assign n24173 = n4487 | n24172 ;
  assign n24174 = ~n12314 & n24173 ;
  assign n24175 = ~x26 & n24174 ;
  assign n24176 = x26 | n24175 ;
  assign n24177 = ( ~n24174 & n24175 ) | ( ~n24174 & n24176 ) | ( n24175 & n24176 ) ;
  assign n24178 = n24170 & ~n24177 ;
  assign n24179 = n3628 | n3629 ;
  assign n24180 = n24164 | n24179 ;
  assign n24181 = n543 | n24180 ;
  assign n24182 = n669 | n24181 ;
  assign n24183 = ( n24168 & ~n24178 ) | ( n24168 & n24182 ) | ( ~n24178 & n24182 ) ;
  assign n24184 = ( n24168 & n24169 ) | ( n24168 & n24177 ) | ( n24169 & n24177 ) ;
  assign n24185 = n24182 & n24184 ;
  assign n24186 = n24183 & ~n24185 ;
  assign n24187 = n24159 & n24186 ;
  assign n24188 = n24186 & ~n24187 ;
  assign n24189 = ( n24159 & ~n24187 ) | ( n24159 & n24188 ) | ( ~n24187 & n24188 ) ;
  assign n24190 = n3636 & n13587 ;
  assign n24191 = ( n3636 & n13585 ) | ( n3636 & n24190 ) | ( n13585 & n24190 ) ;
  assign n24192 = n3074 | n3275 ;
  assign n24193 = n552 | n24192 ;
  assign n24194 = n3485 | n24193 ;
  assign n24195 = n3475 | n24194 ;
  assign n24196 = n371 | n1700 ;
  assign n24197 = n446 | n24196 ;
  assign n24198 = n24195 | n24197 ;
  assign n24199 = n3462 | n24198 ;
  assign n24200 = n528 | n670 ;
  assign n24201 = n451 | n24200 ;
  assign n24202 = ( n55 & ~n3413 ) | ( n55 & n24201 ) | ( ~n3413 & n24201 ) ;
  assign n24203 = n3413 | n24202 ;
  assign n24204 = n24199 | n24203 ;
  assign n24205 = n20958 | n24204 ;
  assign n24206 = n20958 & n24204 ;
  assign n24207 = n3744 & ~n12335 ;
  assign n24208 = n3639 & ~n12586 ;
  assign n24209 = n3727 & n12580 ;
  assign n24210 = n24208 | n24209 ;
  assign n24211 = n24207 | n24210 ;
  assign n24212 = ( n24205 & n24206 ) | ( n24205 & n24211 ) | ( n24206 & n24211 ) ;
  assign n24213 = ( n24191 & n24205 ) | ( n24191 & n24212 ) | ( n24205 & n24212 ) ;
  assign n24214 = ~n24170 & n24177 ;
  assign n24215 = n24178 | n24214 ;
  assign n24216 = n3744 & ~n12325 ;
  assign n24217 = n3639 & n12580 ;
  assign n24218 = n3727 & ~n12335 ;
  assign n24219 = n24217 | n24218 ;
  assign n24220 = n24216 | n24219 ;
  assign n24221 = n3636 | n24220 ;
  assign n24222 = ( ~n13720 & n24220 ) | ( ~n13720 & n24221 ) | ( n24220 & n24221 ) ;
  assign n24223 = ( ~n24213 & n24215 ) | ( ~n24213 & n24222 ) | ( n24215 & n24222 ) ;
  assign n24224 = ( n24213 & ~n24215 ) | ( n24213 & n24223 ) | ( ~n24215 & n24223 ) ;
  assign n24225 = n24189 | n24224 ;
  assign n24226 = n24189 & n24224 ;
  assign n24227 = n24225 & ~n24226 ;
  assign n24228 = n4045 & ~n12318 ;
  assign n24229 = n4043 & n12608 ;
  assign n24230 = n24228 | n24229 ;
  assign n24231 = n4048 & ~n12314 ;
  assign n24232 = n24230 | n24231 ;
  assign n24233 = n4051 | n24232 ;
  assign n24234 = ( ~n14302 & n24232 ) | ( ~n14302 & n24233 ) | ( n24232 & n24233 ) ;
  assign n24235 = ~x29 & n24234 ;
  assign n24236 = x29 | n24235 ;
  assign n24237 = ( ~n24234 & n24235 ) | ( ~n24234 & n24236 ) | ( n24235 & n24236 ) ;
  assign n24238 = n24227 & n24237 ;
  assign n24239 = n24227 | n24237 ;
  assign n24240 = ~n24238 & n24239 ;
  assign n24241 = ( ~n24222 & n24223 ) | ( ~n24222 & n24224 ) | ( n24223 & n24224 ) ;
  assign n24242 = n4048 & ~n12318 ;
  assign n24243 = n4043 & ~n12328 ;
  assign n24244 = n4045 & n12608 ;
  assign n24245 = n24243 | n24244 ;
  assign n24246 = n24242 | n24245 ;
  assign n24247 = n4051 | n24246 ;
  assign n24248 = ( n14320 & n24246 ) | ( n14320 & n24247 ) | ( n24246 & n24247 ) ;
  assign n24249 = x29 & n24248 ;
  assign n24250 = x29 & ~n24249 ;
  assign n24251 = ( n24248 & ~n24249 ) | ( n24248 & n24250 ) | ( ~n24249 & n24250 ) ;
  assign n24252 = ~n24241 & n24251 ;
  assign n24253 = n24241 & ~n24251 ;
  assign n24254 = n24252 | n24253 ;
  assign n24255 = n20959 | n20971 ;
  assign n24256 = n24205 & ~n24212 ;
  assign n24257 = ~n24191 & n24256 ;
  assign n24258 = n24255 & n24257 ;
  assign n24259 = n24205 & ~n24206 ;
  assign n24260 = n24191 & ~n24259 ;
  assign n24261 = ( n24211 & ~n24259 ) | ( n24211 & n24260 ) | ( ~n24259 & n24260 ) ;
  assign n24262 = ( n24255 & n24258 ) | ( n24255 & n24261 ) | ( n24258 & n24261 ) ;
  assign n24263 = n24255 | n24257 ;
  assign n24264 = n24261 | n24263 ;
  assign n24265 = ~n24262 & n24264 ;
  assign n24266 = n20975 | n20987 ;
  assign n24267 = n24265 & n24266 ;
  assign n24268 = n24262 | n24267 ;
  assign n24269 = ~n24254 & n24268 ;
  assign n24270 = n24252 | n24269 ;
  assign n24271 = n24240 & n24270 ;
  assign n24272 = n24240 | n24270 ;
  assign n24273 = ~n24271 & n24272 ;
  assign n24274 = n24254 & ~n24268 ;
  assign n24275 = n24269 | n24274 ;
  assign n24276 = ~n12314 & n24171 ;
  assign n24277 = ( ~n12318 & n24172 ) | ( ~n12318 & n24276 ) | ( n24172 & n24276 ) ;
  assign n24278 = n4487 & ~n17966 ;
  assign n24279 = n24277 | n24278 ;
  assign n24280 = x26 & ~n24279 ;
  assign n24281 = ~x26 & n24279 ;
  assign n24282 = n24280 | n24281 ;
  assign n24283 = n4051 & n13570 ;
  assign n24284 = ( n4051 & n13568 ) | ( n4051 & n24283 ) | ( n13568 & n24283 ) ;
  assign n24285 = n4043 & ~n12325 ;
  assign n24286 = n4045 & ~n12328 ;
  assign n24287 = n24285 | n24286 ;
  assign n24288 = n4048 & n12608 ;
  assign n24289 = n24287 | n24288 ;
  assign n24290 = n24284 | n24289 ;
  assign n24291 = ~x29 & n24290 ;
  assign n24292 = x29 & ~n24290 ;
  assign n24293 = n24291 | n24292 ;
  assign n24294 = n24282 & n24293 ;
  assign n24295 = n24265 | n24266 ;
  assign n24296 = ~n24267 & n24295 ;
  assign n24297 = n24282 | n24293 ;
  assign n24298 = ~n24294 & n24297 ;
  assign n24299 = n24296 & n24298 ;
  assign n24300 = n24294 | n24299 ;
  assign n24301 = ~n24275 & n24300 ;
  assign n24302 = n24275 & ~n24300 ;
  assign n24303 = n24301 | n24302 ;
  assign n24304 = n24296 | n24298 ;
  assign n24305 = ~n24299 & n24304 ;
  assign n24306 = n20990 & n24305 ;
  assign n24307 = n20990 | n24305 ;
  assign n24308 = ~n24306 & n24307 ;
  assign n24309 = n20994 | n20999 ;
  assign n24310 = n24308 & n24309 ;
  assign n24311 = n24306 | n24310 ;
  assign n24312 = ~n24303 & n24311 ;
  assign n24313 = n24301 | n24312 ;
  assign n24314 = n24273 & n24313 ;
  assign n24315 = n20994 | n21001 ;
  assign n24316 = n24308 & n24315 ;
  assign n24317 = n24306 | n24316 ;
  assign n24318 = ~n24303 & n24317 ;
  assign n24319 = n24301 | n24318 ;
  assign n24320 = n24273 & n24319 ;
  assign n24321 = ( n19561 & n24314 ) | ( n19561 & n24320 ) | ( n24314 & n24320 ) ;
  assign n24322 = ( n19561 & n24313 ) | ( n19561 & n24319 ) | ( n24313 & n24319 ) ;
  assign n24323 = n24273 | n24322 ;
  assign n24324 = ~n24321 & n24323 ;
  assign n24325 = n9798 & n24324 ;
  assign n24326 = ( n19561 & n24310 ) | ( n19561 & n24316 ) | ( n24310 & n24316 ) ;
  assign n24327 = ( n19561 & n24309 ) | ( n19561 & n24315 ) | ( n24309 & n24315 ) ;
  assign n24328 = n24308 | n24327 ;
  assign n24329 = ~n24326 & n24328 ;
  assign n24330 = n9782 & n24329 ;
  assign n24331 = ( n19561 & n24312 ) | ( n19561 & n24318 ) | ( n24312 & n24318 ) ;
  assign n24332 = ( n19561 & n24311 ) | ( n19561 & n24317 ) | ( n24311 & n24317 ) ;
  assign n24333 = n24303 & ~n24332 ;
  assign n24334 = n24331 | n24333 ;
  assign n24335 = n9783 & ~n24334 ;
  assign n24336 = n24330 | n24335 ;
  assign n24337 = n24325 | n24336 ;
  assign n24338 = ~n24324 & n24334 ;
  assign n24339 = n24324 & ~n24334 ;
  assign n24340 = ~n24329 & n24334 ;
  assign n24341 = n21005 & ~n24329 ;
  assign n24342 = n24340 | n24341 ;
  assign n24343 = n24338 | n24342 ;
  assign n24344 = n24339 | n24343 ;
  assign n24345 = ~n24339 & n24344 ;
  assign n24346 = n24329 & ~n24334 ;
  assign n24347 = ~n21005 & n24329 ;
  assign n24348 = n24346 | n24347 ;
  assign n24349 = ~n24338 & n24348 ;
  assign n24350 = ~n24339 & n24349 ;
  assign n24351 = n24339 | n24350 ;
  assign n24352 = ( n21013 & ~n24345 ) | ( n21013 & n24351 ) | ( ~n24345 & n24351 ) ;
  assign n24353 = n24338 | n24352 ;
  assign n24354 = ( n21013 & ~n24342 ) | ( n21013 & n24348 ) | ( ~n24342 & n24348 ) ;
  assign n24355 = ( n21013 & ~n24344 ) | ( n21013 & n24350 ) | ( ~n24344 & n24350 ) ;
  assign n24356 = n24354 & ~n24355 ;
  assign n24357 = n9787 & ~n24356 ;
  assign n24358 = n24353 & n24357 ;
  assign n24359 = ( n9787 & n24337 ) | ( n9787 & ~n24358 ) | ( n24337 & ~n24358 ) ;
  assign n24360 = x2 & n24359 ;
  assign n24361 = x2 & ~n24360 ;
  assign n24362 = ( n24359 & ~n24360 ) | ( n24359 & n24361 ) | ( ~n24360 & n24361 ) ;
  assign n24363 = ~n24152 & n24362 ;
  assign n24364 = n24152 & ~n24362 ;
  assign n24365 = n24363 | n24364 ;
  assign n24366 = n23703 & ~n24147 ;
  assign n24367 = n24148 | n24366 ;
  assign n24368 = n9798 & ~n24334 ;
  assign n24369 = n9782 & ~n21005 ;
  assign n24370 = n9783 & n24329 ;
  assign n24371 = n24369 | n24370 ;
  assign n24372 = n24368 | n24371 ;
  assign n24373 = n24340 | n24354 ;
  assign n24374 = ( ~n21013 & n24329 ) | ( ~n21013 & n24334 ) | ( n24329 & n24334 ) ;
  assign n24375 = ( ~n21005 & n24329 ) | ( ~n21005 & n24334 ) | ( n24329 & n24334 ) ;
  assign n24376 = ( n24346 & ~n24374 ) | ( n24346 & n24375 ) | ( ~n24374 & n24375 ) ;
  assign n24377 = n9787 & ~n24376 ;
  assign n24378 = n24373 & n24377 ;
  assign n24379 = ( n9787 & n24372 ) | ( n9787 & ~n24378 ) | ( n24372 & ~n24378 ) ;
  assign n24380 = x2 & n24379 ;
  assign n24381 = x2 & ~n24380 ;
  assign n24382 = ( n24379 & ~n24380 ) | ( n24379 & n24381 ) | ( ~n24380 & n24381 ) ;
  assign n24383 = ~n24367 & n24382 ;
  assign n24384 = ~n24365 & n24383 ;
  assign n24385 = n9798 & n24329 ;
  assign n24386 = n9782 & n20921 ;
  assign n24387 = n9783 & ~n21005 ;
  assign n24388 = n24386 | n24387 ;
  assign n24389 = n24385 | n24388 ;
  assign n24390 = n24341 | n24347 ;
  assign n24391 = n21013 | n24390 ;
  assign n24392 = n21013 & n24390 ;
  assign n24393 = n9787 & ~n24392 ;
  assign n24394 = n24391 & n24393 ;
  assign n24395 = ( n9787 & n24389 ) | ( n9787 & ~n24394 ) | ( n24389 & ~n24394 ) ;
  assign n24396 = x2 & n24395 ;
  assign n24397 = x2 & ~n24396 ;
  assign n24398 = ( n24395 & ~n24396 ) | ( n24395 & n24397 ) | ( ~n24396 & n24397 ) ;
  assign n24399 = n9798 & ~n21005 ;
  assign n24400 = n9782 & n20838 ;
  assign n24401 = n9783 & n20921 ;
  assign n24402 = n24400 | n24401 ;
  assign n24403 = n24399 | n24402 ;
  assign n24404 = n9787 | n24403 ;
  assign n24405 = ( ~n21015 & n24403 ) | ( ~n21015 & n24404 ) | ( n24403 & n24404 ) ;
  assign n24406 = ~x2 & n24405 ;
  assign n24407 = x2 | n24406 ;
  assign n24408 = ( ~n24405 & n24406 ) | ( ~n24405 & n24407 ) | ( n24406 & n24407 ) ;
  assign n24409 = n9798 & n20921 ;
  assign n24410 = n9782 & n20532 ;
  assign n24411 = n9783 & n20838 ;
  assign n24412 = n24410 | n24411 ;
  assign n24413 = n24409 | n24412 ;
  assign n24414 = n9787 & ~n23691 ;
  assign n24415 = ~n23695 & n24414 ;
  assign n24416 = ( n9787 & n24413 ) | ( n9787 & ~n24415 ) | ( n24413 & ~n24415 ) ;
  assign n24417 = ~x2 & n24416 ;
  assign n24418 = x2 | n24417 ;
  assign n24419 = ( ~n24416 & n24417 ) | ( ~n24416 & n24418 ) | ( n24417 & n24418 ) ;
  assign n24420 = n23756 | n24142 ;
  assign n24421 = ~n24143 & n24420 ;
  assign n24422 = ( n23758 & n24141 ) | ( n23758 & ~n24142 ) | ( n24141 & ~n24142 ) ;
  assign n24423 = ( n23768 & ~n24142 ) | ( n23768 & n24422 ) | ( ~n24142 & n24422 ) ;
  assign n24424 = n9798 & ~n20536 ;
  assign n24425 = n9782 & ~n20542 ;
  assign n24426 = n9783 & ~n20724 ;
  assign n24427 = n24425 | n24426 ;
  assign n24428 = n24424 | n24427 ;
  assign n24429 = n9787 & ~n23213 ;
  assign n24430 = n23217 & n24429 ;
  assign n24431 = ( n9787 & n24428 ) | ( n9787 & ~n24430 ) | ( n24428 & ~n24430 ) ;
  assign n24432 = x2 & n24431 ;
  assign n24433 = x2 & ~n24432 ;
  assign n24434 = ( n24431 & ~n24432 ) | ( n24431 & n24433 ) | ( ~n24432 & n24433 ) ;
  assign n24435 = n9798 & ~n20724 ;
  assign n24436 = n9782 & n20546 ;
  assign n24437 = n9783 & ~n20542 ;
  assign n24438 = n24436 | n24437 ;
  assign n24439 = n24435 | n24438 ;
  assign n24440 = n9787 | n24439 ;
  assign n24441 = ( n23229 & n24439 ) | ( n23229 & n24440 ) | ( n24439 & n24440 ) ;
  assign n24442 = x2 & n24441 ;
  assign n24443 = x2 & ~n24442 ;
  assign n24444 = ( n24441 & ~n24442 ) | ( n24441 & n24443 ) | ( ~n24442 & n24443 ) ;
  assign n24445 = n9798 & ~n20542 ;
  assign n24446 = n9782 & ~n20710 ;
  assign n24447 = n9783 & n20546 ;
  assign n24448 = n24446 | n24447 ;
  assign n24449 = n24445 | n24448 ;
  assign n24450 = n9787 | n24449 ;
  assign n24451 = ( ~n23042 & n24449 ) | ( ~n23042 & n24450 ) | ( n24449 & n24450 ) ;
  assign n24452 = ~x2 & n24451 ;
  assign n24453 = x2 | n24452 ;
  assign n24454 = ( ~n24451 & n24452 ) | ( ~n24451 & n24453 ) | ( n24452 & n24453 ) ;
  assign n24455 = n23835 | n23837 ;
  assign n24456 = n24136 | n24455 ;
  assign n24457 = ~n24137 & n24456 ;
  assign n24458 = ( ~n24133 & n24134 ) | ( ~n24133 & n24135 ) | ( n24134 & n24135 ) ;
  assign n24459 = n24133 | n24458 ;
  assign n24460 = ~n24136 & n24459 ;
  assign n24461 = n23866 | n24127 ;
  assign n24462 = ~n24128 & n24461 ;
  assign n24463 = n9798 & n20562 ;
  assign n24464 = n9782 & ~n20689 ;
  assign n24465 = n9783 & n20560 ;
  assign n24466 = n24464 | n24465 ;
  assign n24467 = n24463 | n24466 ;
  assign n24468 = n9787 | n24467 ;
  assign n24469 = ( ~n21044 & n24467 ) | ( ~n21044 & n24468 ) | ( n24467 & n24468 ) ;
  assign n24470 = ~x2 & n24469 ;
  assign n24471 = x2 | n24470 ;
  assign n24472 = ( ~n24469 & n24470 ) | ( ~n24469 & n24471 ) | ( n24470 & n24471 ) ;
  assign n24473 = n9798 & n20560 ;
  assign n24474 = n9782 & ~n20573 ;
  assign n24475 = n9783 & ~n20689 ;
  assign n24476 = n24474 | n24475 ;
  assign n24477 = n24473 | n24476 ;
  assign n24478 = n9787 & ~n22176 ;
  assign n24479 = ~n22173 & n24478 ;
  assign n24480 = ( n9787 & n24477 ) | ( n9787 & ~n24479 ) | ( n24477 & ~n24479 ) ;
  assign n24481 = ~x2 & n24480 ;
  assign n24482 = x2 | n24481 ;
  assign n24483 = ( ~n24480 & n24481 ) | ( ~n24480 & n24482 ) | ( n24481 & n24482 ) ;
  assign n24484 = n23902 | n24119 ;
  assign n24485 = ~n24120 & n24484 ;
  assign n24486 = n9787 & n21884 ;
  assign n24487 = ( n9787 & ~n21889 ) | ( n9787 & n24486 ) | ( ~n21889 & n24486 ) ;
  assign n24488 = n9798 & ~n20569 ;
  assign n24489 = n9782 & ~n20580 ;
  assign n24490 = n9783 & ~n20584 ;
  assign n24491 = n24489 | n24490 ;
  assign n24492 = n24488 | n24491 ;
  assign n24493 = n24487 | n24492 ;
  assign n24494 = x2 & n24493 ;
  assign n24495 = n9798 & ~n20584 ;
  assign n24496 = n9782 & n20588 ;
  assign n24497 = n9783 & ~n20580 ;
  assign n24498 = n24496 | n24497 ;
  assign n24499 = n24495 | n24498 ;
  assign n24500 = n9787 | n24499 ;
  assign n24501 = ( ~n21901 & n24499 ) | ( ~n21901 & n24500 ) | ( n24499 & n24500 ) ;
  assign n24502 = ~x2 & n24501 ;
  assign n24503 = x2 | n24502 ;
  assign n24504 = ( ~n24501 & n24502 ) | ( ~n24501 & n24503 ) | ( n24502 & n24503 ) ;
  assign n24505 = n9798 & ~n20580 ;
  assign n24506 = n9782 & ~n20591 ;
  assign n24507 = n9783 & n20588 ;
  assign n24508 = n24506 | n24507 ;
  assign n24509 = n24505 | n24508 ;
  assign n24510 = n9787 | n24509 ;
  assign n24511 = ( n21840 & n24509 ) | ( n21840 & n24510 ) | ( n24509 & n24510 ) ;
  assign n24512 = x2 & n24511 ;
  assign n24513 = x2 & ~n24512 ;
  assign n24514 = ( n24511 & ~n24512 ) | ( n24511 & n24513 ) | ( ~n24512 & n24513 ) ;
  assign n24515 = n9798 & n20588 ;
  assign n24516 = n9782 & ~n20595 ;
  assign n24517 = n9783 & ~n20591 ;
  assign n24518 = n24516 | n24517 ;
  assign n24519 = n24515 | n24518 ;
  assign n24520 = n9787 | n24519 ;
  assign n24521 = ( n21526 & n24519 ) | ( n21526 & n24520 ) | ( n24519 & n24520 ) ;
  assign n24522 = x2 & n24521 ;
  assign n24523 = x2 & ~n24522 ;
  assign n24524 = ( n24521 & ~n24522 ) | ( n24521 & n24523 ) | ( ~n24522 & n24523 ) ;
  assign n24525 = n23992 | n24112 ;
  assign n24526 = n24110 | n24525 ;
  assign n24527 = ~n24113 & n24526 ;
  assign n24528 = n24107 | n24109 ;
  assign n24529 = ~n24110 & n24528 ;
  assign n24530 = n24102 | n24105 ;
  assign n24531 = ~n24106 & n24530 ;
  assign n24532 = n24033 | n24096 ;
  assign n24533 = ~n24097 & n24532 ;
  assign n24534 = n9798 & n20614 ;
  assign n24535 = n9782 & n20619 ;
  assign n24536 = n9783 | n24535 ;
  assign n24537 = ( n20616 & n24535 ) | ( n20616 & n24536 ) | ( n24535 & n24536 ) ;
  assign n24538 = n24534 | n24537 ;
  assign n24539 = n9787 | n24538 ;
  assign n24540 = ( n21302 & n24538 ) | ( n21302 & n24539 ) | ( n24538 & n24539 ) ;
  assign n24541 = x2 & n24540 ;
  assign n24542 = x2 & ~n24541 ;
  assign n24543 = ( n24540 & ~n24541 ) | ( n24540 & n24542 ) | ( ~n24541 & n24542 ) ;
  assign n24544 = n24060 | n24093 ;
  assign n24545 = ~n24094 & n24544 ;
  assign n24546 = n24061 | n24082 ;
  assign n24547 = n24061 & n24082 ;
  assign n24548 = n24546 & ~n24547 ;
  assign n24549 = ~n24092 & n24548 ;
  assign n24550 = n9782 & ~n20625 ;
  assign n24551 = n9783 | n24550 ;
  assign n24552 = ( n20622 & n24550 ) | ( n20622 & n24551 ) | ( n24550 & n24551 ) ;
  assign n24553 = n9798 | n24552 ;
  assign n24554 = ( n20619 & n24552 ) | ( n20619 & n24553 ) | ( n24552 & n24553 ) ;
  assign n24555 = n9787 | n24554 ;
  assign n24556 = ( ~n21056 & n24554 ) | ( ~n21056 & n24555 ) | ( n24554 & n24555 ) ;
  assign n24557 = ~x2 & n24556 ;
  assign n24558 = x2 | n24557 ;
  assign n24559 = ( ~n24556 & n24557 ) | ( ~n24556 & n24558 ) | ( n24557 & n24558 ) ;
  assign n24560 = n8678 & ~n20642 ;
  assign n24561 = n10020 & n21069 ;
  assign n24562 = n10033 & ~n20642 ;
  assign n24563 = ( x2 & n10031 ) | ( x2 & n20640 ) | ( n10031 & n20640 ) ;
  assign n24564 = ~n24562 & n24563 ;
  assign n24565 = ~n24561 & n24564 ;
  assign n24566 = n9782 & ~n20642 ;
  assign n24567 = n9783 & ~n20640 ;
  assign n24568 = n24566 | n24567 ;
  assign n24569 = n9798 & n20633 ;
  assign n24570 = x2 & n24569 ;
  assign n24571 = ( x2 & n24568 ) | ( x2 & n24570 ) | ( n24568 & n24570 ) ;
  assign n24572 = n24565 & ~n24571 ;
  assign n24573 = x0 & ~n20642 ;
  assign n24574 = n10020 & n21085 ;
  assign n24575 = n24573 | n24574 ;
  assign n24576 = n24572 & ~n24575 ;
  assign n24577 = n9798 & ~n20630 ;
  assign n24578 = n9782 & ~n20640 ;
  assign n24579 = n9783 & n20633 ;
  assign n24580 = n24578 | n24579 ;
  assign n24581 = n24577 | n24580 ;
  assign n24582 = n9787 | n24581 ;
  assign n24583 = ( n21099 & n24581 ) | ( n21099 & n24582 ) | ( n24581 & n24582 ) ;
  assign n24584 = x2 & n24583 ;
  assign n24585 = x2 & ~n24584 ;
  assign n24586 = ( n24583 & ~n24584 ) | ( n24583 & n24585 ) | ( ~n24584 & n24585 ) ;
  assign n24587 = ( n24560 & n24576 ) | ( n24560 & n24586 ) | ( n24576 & n24586 ) ;
  assign n24588 = n9798 & ~n20625 ;
  assign n24589 = n9782 & n20633 ;
  assign n24590 = n9783 & ~n20630 ;
  assign n24591 = n24589 | n24590 ;
  assign n24592 = n24588 | n24591 ;
  assign n24593 = n9787 | n24592 ;
  assign n24594 = ( ~n21129 & n24592 ) | ( ~n21129 & n24593 ) | ( n24592 & n24593 ) ;
  assign n24595 = ~x2 & n24594 ;
  assign n24596 = x2 | n24595 ;
  assign n24597 = ( ~n24594 & n24595 ) | ( ~n24594 & n24596 ) | ( n24595 & n24596 ) ;
  assign n24598 = n24587 | n24597 ;
  assign n24599 = n24062 | n24070 ;
  assign n24600 = ~n24071 & n24599 ;
  assign n24601 = n24598 & n24600 ;
  assign n24602 = n24071 | n24081 ;
  assign n24603 = ~n24082 & n24602 ;
  assign n24604 = n24587 & n24597 ;
  assign n24605 = n24603 & n24604 ;
  assign n24606 = ( n24601 & n24603 ) | ( n24601 & n24605 ) | ( n24603 & n24605 ) ;
  assign n24607 = n24559 | n24606 ;
  assign n24608 = n9798 & n20622 ;
  assign n24609 = n9782 & ~n20630 ;
  assign n24610 = n9783 & ~n20625 ;
  assign n24611 = n24609 | n24610 ;
  assign n24612 = n24608 | n24611 ;
  assign n24613 = n9787 | n24612 ;
  assign n24614 = ( n21114 & n24612 ) | ( n21114 & n24613 ) | ( n24612 & n24613 ) ;
  assign n24615 = ~x2 & n24614 ;
  assign n24616 = n24603 | n24604 ;
  assign n24617 = n24601 | n24616 ;
  assign n24618 = ( ~n24614 & n24615 ) | ( ~n24614 & n24617 ) | ( n24615 & n24617 ) ;
  assign n24619 = ( x2 & n24615 ) | ( x2 & n24618 ) | ( n24615 & n24618 ) ;
  assign n24620 = n24607 | n24619 ;
  assign n24621 = ( n24092 & n24549 ) | ( n24092 & n24620 ) | ( n24549 & n24620 ) ;
  assign n24622 = ( ~n24548 & n24549 ) | ( ~n24548 & n24621 ) | ( n24549 & n24621 ) ;
  assign n24623 = n24559 & n24606 ;
  assign n24624 = ( n24559 & n24619 ) | ( n24559 & n24623 ) | ( n24619 & n24623 ) ;
  assign n24625 = n24545 & n24624 ;
  assign n24626 = ( n24545 & n24622 ) | ( n24545 & n24625 ) | ( n24622 & n24625 ) ;
  assign n24627 = n24543 & n24626 ;
  assign n24628 = n9782 & n20622 ;
  assign n24629 = n9783 | n24628 ;
  assign n24630 = ( n20619 & n24628 ) | ( n20619 & n24629 ) | ( n24628 & n24629 ) ;
  assign n24631 = n9798 | n24630 ;
  assign n24632 = ( n20616 & n24630 ) | ( n20616 & n24631 ) | ( n24630 & n24631 ) ;
  assign n24633 = n9787 | n24632 ;
  assign n24634 = ( n21190 & n24632 ) | ( n21190 & n24633 ) | ( n24632 & n24633 ) ;
  assign n24635 = ~x2 & n24634 ;
  assign n24636 = n24545 | n24624 ;
  assign n24637 = n24622 | n24636 ;
  assign n24638 = ( ~n24634 & n24635 ) | ( ~n24634 & n24637 ) | ( n24635 & n24637 ) ;
  assign n24639 = ( x2 & n24635 ) | ( x2 & n24638 ) | ( n24635 & n24638 ) ;
  assign n24640 = ( n24543 & n24627 ) | ( n24543 & n24639 ) | ( n24627 & n24639 ) ;
  assign n24641 = n9798 & n20611 ;
  assign n24642 = n9782 & n20616 ;
  assign n24643 = n9783 & n20614 ;
  assign n24644 = n24642 | n24643 ;
  assign n24645 = n24641 | n24644 ;
  assign n24646 = n9787 | n24645 ;
  assign n24647 = ( n21293 & n24645 ) | ( n21293 & n24646 ) | ( n24645 & n24646 ) ;
  assign n24648 = x2 & n24647 ;
  assign n24649 = x2 & ~n24648 ;
  assign n24650 = ( n24647 & ~n24648 ) | ( n24647 & n24649 ) | ( ~n24648 & n24649 ) ;
  assign n24651 = n24640 | n24650 ;
  assign n24652 = n24543 | n24626 ;
  assign n24653 = n24639 | n24652 ;
  assign n24654 = ( ~n24035 & n24045 ) | ( ~n24035 & n24095 ) | ( n24045 & n24095 ) ;
  assign n24655 = ( n24035 & ~n24045 ) | ( n24035 & n24095 ) | ( ~n24045 & n24095 ) ;
  assign n24656 = ( ~n24095 & n24654 ) | ( ~n24095 & n24655 ) | ( n24654 & n24655 ) ;
  assign n24657 = n24653 & n24656 ;
  assign n24658 = n24651 | n24657 ;
  assign n24659 = n24533 & n24658 ;
  assign n24660 = n9798 & ~n20605 ;
  assign n24661 = n9782 & n20614 ;
  assign n24662 = n9783 & n20611 ;
  assign n24663 = n24661 | n24662 ;
  assign n24664 = n24660 | n24663 ;
  assign n24665 = n9787 | n24664 ;
  assign n24666 = ( ~n21275 & n24664 ) | ( ~n21275 & n24665 ) | ( n24664 & n24665 ) ;
  assign n24667 = ~x2 & n24666 ;
  assign n24668 = x2 | n24667 ;
  assign n24669 = ( ~n24666 & n24667 ) | ( ~n24666 & n24668 ) | ( n24667 & n24668 ) ;
  assign n24670 = n24640 & n24650 ;
  assign n24671 = ( n24650 & n24657 ) | ( n24650 & n24670 ) | ( n24657 & n24670 ) ;
  assign n24672 = n24669 | n24671 ;
  assign n24673 = n24659 | n24672 ;
  assign n24674 = ( n24098 & n24100 ) | ( n24098 & n24673 ) | ( n24100 & n24673 ) ;
  assign n24675 = ~n24101 & n24674 ;
  assign n24676 = n24669 & n24671 ;
  assign n24677 = ( n24659 & n24669 ) | ( n24659 & n24676 ) | ( n24669 & n24676 ) ;
  assign n24678 = n24531 & n24677 ;
  assign n24679 = ( n24531 & n24675 ) | ( n24531 & n24678 ) | ( n24675 & n24678 ) ;
  assign n24680 = n24529 & n24679 ;
  assign n24681 = n9798 & n20600 ;
  assign n24682 = n9782 & n20611 ;
  assign n24683 = n9783 & ~n20605 ;
  assign n24684 = n24682 | n24683 ;
  assign n24685 = n24681 | n24684 ;
  assign n24686 = n9787 | n24685 ;
  assign n24687 = ( ~n21432 & n24685 ) | ( ~n21432 & n24686 ) | ( n24685 & n24686 ) ;
  assign n24688 = ~x2 & n24687 ;
  assign n24689 = n24531 | n24677 ;
  assign n24690 = n24675 | n24689 ;
  assign n24691 = ( ~n24687 & n24688 ) | ( ~n24687 & n24690 ) | ( n24688 & n24690 ) ;
  assign n24692 = ( x2 & n24688 ) | ( x2 & n24691 ) | ( n24688 & n24691 ) ;
  assign n24693 = ( n24529 & n24680 ) | ( n24529 & n24692 ) | ( n24680 & n24692 ) ;
  assign n24694 = n24527 & n24693 ;
  assign n24695 = n9798 & ~n20595 ;
  assign n24696 = n9782 & ~n20605 ;
  assign n24697 = n9783 & n20600 ;
  assign n24698 = n24696 | n24697 ;
  assign n24699 = n24695 | n24698 ;
  assign n24700 = n9787 | n24699 ;
  assign n24701 = ( ~n21554 & n24699 ) | ( ~n21554 & n24700 ) | ( n24699 & n24700 ) ;
  assign n24702 = ~x2 & n24701 ;
  assign n24703 = n24529 | n24679 ;
  assign n24704 = n24692 | n24703 ;
  assign n24705 = ( ~n24701 & n24702 ) | ( ~n24701 & n24704 ) | ( n24702 & n24704 ) ;
  assign n24706 = ( x2 & n24702 ) | ( x2 & n24705 ) | ( n24702 & n24705 ) ;
  assign n24707 = ( n24527 & n24694 ) | ( n24527 & n24706 ) | ( n24694 & n24706 ) ;
  assign n24708 = n24524 & n24707 ;
  assign n24709 = n9787 & n21539 ;
  assign n24710 = ( n9787 & n21543 ) | ( n9787 & n24709 ) | ( n21543 & n24709 ) ;
  assign n24711 = n9798 & ~n20591 ;
  assign n24712 = n9782 & n20600 ;
  assign n24713 = n9783 & ~n20595 ;
  assign n24714 = n24712 | n24713 ;
  assign n24715 = n24711 | n24714 ;
  assign n24716 = n24710 | n24715 ;
  assign n24717 = x2 & n24716 ;
  assign n24718 = n24527 | n24693 ;
  assign n24719 = n24706 | n24718 ;
  assign n24720 = ( x2 & n24716 ) | ( x2 & n24719 ) | ( n24716 & n24719 ) ;
  assign n24721 = ~n24717 & n24720 ;
  assign n24722 = ( n24524 & n24708 ) | ( n24524 & n24721 ) | ( n24708 & n24721 ) ;
  assign n24723 = n24514 & n24722 ;
  assign n24724 = n24524 | n24707 ;
  assign n24725 = n24721 | n24724 ;
  assign n24726 = ( ~n23956 & n23966 ) | ( ~n23956 & n24114 ) | ( n23966 & n24114 ) ;
  assign n24727 = ( n23956 & ~n23966 ) | ( n23956 & n24114 ) | ( ~n23966 & n24114 ) ;
  assign n24728 = ( ~n24114 & n24726 ) | ( ~n24114 & n24727 ) | ( n24726 & n24727 ) ;
  assign n24729 = n24725 & n24728 ;
  assign n24730 = ( n24514 & n24723 ) | ( n24514 & n24729 ) | ( n24723 & n24729 ) ;
  assign n24731 = n24504 & n24730 ;
  assign n24732 = n24514 | n24722 ;
  assign n24733 = n24729 | n24732 ;
  assign n24734 = ( ~n23943 & n23953 ) | ( ~n23943 & n24115 ) | ( n23953 & n24115 ) ;
  assign n24735 = ( n23943 & ~n23953 ) | ( n23943 & n24115 ) | ( ~n23953 & n24115 ) ;
  assign n24736 = ( ~n24115 & n24734 ) | ( ~n24115 & n24735 ) | ( n24734 & n24735 ) ;
  assign n24737 = n24733 & n24736 ;
  assign n24738 = ( n24504 & n24731 ) | ( n24504 & n24737 ) | ( n24731 & n24737 ) ;
  assign n24739 = ( n23916 & n24117 ) | ( n23916 & ~n24118 ) | ( n24117 & ~n24118 ) ;
  assign n24740 = ( n23926 & ~n24118 ) | ( n23926 & n24739 ) | ( ~n24118 & n24739 ) ;
  assign n24741 = n24738 | n24740 ;
  assign n24742 = n24504 | n24730 ;
  assign n24743 = n24737 | n24742 ;
  assign n24744 = ( ~n23929 & n23940 ) | ( ~n23929 & n24116 ) | ( n23940 & n24116 ) ;
  assign n24745 = ( n23929 & ~n23940 ) | ( n23929 & n24116 ) | ( ~n23940 & n24116 ) ;
  assign n24746 = ( ~n24116 & n24744 ) | ( ~n24116 & n24745 ) | ( n24744 & n24745 ) ;
  assign n24747 = n24743 & n24746 ;
  assign n24748 = n24741 | n24747 ;
  assign n24749 = ( x2 & n24493 ) | ( x2 & n24748 ) | ( n24493 & n24748 ) ;
  assign n24750 = ~n24494 & n24749 ;
  assign n24751 = ( n23904 & n24118 ) | ( n23904 & ~n24119 ) | ( n24118 & ~n24119 ) ;
  assign n24752 = ( n23914 & ~n24119 ) | ( n23914 & n24751 ) | ( ~n24119 & n24751 ) ;
  assign n24753 = n24738 & n24740 ;
  assign n24754 = ( n24740 & n24747 ) | ( n24740 & n24753 ) | ( n24747 & n24753 ) ;
  assign n24755 = n24752 & n24754 ;
  assign n24756 = ( n24750 & n24752 ) | ( n24750 & n24755 ) | ( n24752 & n24755 ) ;
  assign n24757 = n24485 & n24756 ;
  assign n24758 = n9798 & ~n20573 ;
  assign n24759 = n9782 & ~n20584 ;
  assign n24760 = n9783 & ~n20569 ;
  assign n24761 = n24759 | n24760 ;
  assign n24762 = n24758 | n24761 ;
  assign n24763 = n9787 | n24762 ;
  assign n24764 = ( ~n21860 & n24762 ) | ( ~n21860 & n24763 ) | ( n24762 & n24763 ) ;
  assign n24765 = ~x2 & n24764 ;
  assign n24766 = n24752 | n24754 ;
  assign n24767 = n24750 | n24766 ;
  assign n24768 = ( ~n24764 & n24765 ) | ( ~n24764 & n24767 ) | ( n24765 & n24767 ) ;
  assign n24769 = ( x2 & n24765 ) | ( x2 & n24768 ) | ( n24765 & n24768 ) ;
  assign n24770 = ( n24485 & n24757 ) | ( n24485 & n24769 ) | ( n24757 & n24769 ) ;
  assign n24771 = n24483 & n24770 ;
  assign n24772 = n9798 & ~n20689 ;
  assign n24773 = n9782 & ~n20569 ;
  assign n24774 = n9783 & ~n20573 ;
  assign n24775 = n24773 | n24774 ;
  assign n24776 = n24772 | n24775 ;
  assign n24777 = ( n9787 & ~n22192 ) | ( n9787 & n22193 ) | ( ~n22192 & n22193 ) ;
  assign n24778 = n24776 | n24777 ;
  assign n24779 = x2 & n24778 ;
  assign n24780 = n24485 | n24756 ;
  assign n24781 = n24769 | n24780 ;
  assign n24782 = ( x2 & n24778 ) | ( x2 & n24781 ) | ( n24778 & n24781 ) ;
  assign n24783 = ~n24779 & n24782 ;
  assign n24784 = ( n24483 & n24771 ) | ( n24483 & n24783 ) | ( n24771 & n24783 ) ;
  assign n24785 = n24472 & n24784 ;
  assign n24786 = n24483 | n24770 ;
  assign n24787 = n24783 | n24786 ;
  assign n24788 = ( n23887 & n24121 ) | ( n23887 & ~n24123 ) | ( n24121 & ~n24123 ) ;
  assign n24789 = ( ~n23887 & n24121 ) | ( ~n23887 & n24123 ) | ( n24121 & n24123 ) ;
  assign n24790 = ( ~n24121 & n24788 ) | ( ~n24121 & n24789 ) | ( n24788 & n24789 ) ;
  assign n24791 = n24787 & n24790 ;
  assign n24792 = ( n24472 & n24785 ) | ( n24472 & n24791 ) | ( n24785 & n24791 ) ;
  assign n24793 = n9798 & ~n20552 ;
  assign n24794 = n9782 & n20560 ;
  assign n24795 = n9783 & n20562 ;
  assign n24796 = n24794 | n24795 ;
  assign n24797 = n24793 | n24796 ;
  assign n24798 = n9787 & n22510 ;
  assign n24799 = ~n22512 & n24798 ;
  assign n24800 = ( n9787 & n24797 ) | ( n9787 & ~n24799 ) | ( n24797 & ~n24799 ) ;
  assign n24801 = x2 & n24800 ;
  assign n24802 = x2 & ~n24801 ;
  assign n24803 = ( n24800 & ~n24801 ) | ( n24800 & n24802 ) | ( ~n24801 & n24802 ) ;
  assign n24804 = n24792 | n24803 ;
  assign n24805 = n24472 | n24784 ;
  assign n24806 = n24791 | n24805 ;
  assign n24807 = ( n23876 & n24124 ) | ( n23876 & ~n24126 ) | ( n24124 & ~n24126 ) ;
  assign n24808 = ( ~n23876 & n24124 ) | ( ~n23876 & n24126 ) | ( n24124 & n24126 ) ;
  assign n24809 = ( ~n24124 & n24807 ) | ( ~n24124 & n24808 ) | ( n24807 & n24808 ) ;
  assign n24810 = n24806 & n24809 ;
  assign n24811 = n24804 | n24810 ;
  assign n24812 = n24462 & n24811 ;
  assign n24813 = ( ~n24129 & n24130 ) | ( ~n24129 & n24131 ) | ( n24130 & n24131 ) ;
  assign n24814 = n24129 | n24813 ;
  assign n24815 = ~n24132 & n24814 ;
  assign n24816 = n24792 & n24803 ;
  assign n24817 = ( n24803 & n24810 ) | ( n24803 & n24816 ) | ( n24810 & n24816 ) ;
  assign n24818 = n24815 & n24817 ;
  assign n24819 = ( n24812 & n24815 ) | ( n24812 & n24818 ) | ( n24815 & n24818 ) ;
  assign n24820 = n24460 & n24819 ;
  assign n24821 = n9798 & n20556 ;
  assign n24822 = n9782 & n20562 ;
  assign n24823 = n9783 & ~n20552 ;
  assign n24824 = n24822 | n24823 ;
  assign n24825 = n24821 | n24824 ;
  assign n24826 = n9787 | n24825 ;
  assign n24827 = ( ~n22655 & n24825 ) | ( ~n22655 & n24826 ) | ( n24825 & n24826 ) ;
  assign n24828 = ~x2 & n24827 ;
  assign n24829 = n24815 | n24817 ;
  assign n24830 = n24812 | n24829 ;
  assign n24831 = ( ~n24827 & n24828 ) | ( ~n24827 & n24830 ) | ( n24828 & n24830 ) ;
  assign n24832 = ( x2 & n24828 ) | ( x2 & n24831 ) | ( n24828 & n24831 ) ;
  assign n24833 = ( n24460 & n24820 ) | ( n24460 & n24832 ) | ( n24820 & n24832 ) ;
  assign n24834 = n24457 & n24833 ;
  assign n24835 = n9798 & ~n20710 ;
  assign n24836 = n9782 & ~n20552 ;
  assign n24837 = n9783 & n20556 ;
  assign n24838 = n24836 | n24837 ;
  assign n24839 = n24835 | n24838 ;
  assign n24840 = n9787 | n24839 ;
  assign n24841 = ( ~n22641 & n24839 ) | ( ~n22641 & n24840 ) | ( n24839 & n24840 ) ;
  assign n24842 = ~x2 & n24841 ;
  assign n24843 = n24460 | n24819 ;
  assign n24844 = n24832 | n24843 ;
  assign n24845 = ( ~n24841 & n24842 ) | ( ~n24841 & n24844 ) | ( n24842 & n24844 ) ;
  assign n24846 = ( x2 & n24842 ) | ( x2 & n24845 ) | ( n24842 & n24845 ) ;
  assign n24847 = ( n24457 & n24834 ) | ( n24457 & n24846 ) | ( n24834 & n24846 ) ;
  assign n24848 = n24454 & n24847 ;
  assign n24849 = n9787 & ~n21031 ;
  assign n24850 = ( n9787 & n21037 ) | ( n9787 & n24849 ) | ( n21037 & n24849 ) ;
  assign n24851 = n9798 & n20546 ;
  assign n24852 = n9782 & n20556 ;
  assign n24853 = n9783 & ~n20710 ;
  assign n24854 = n24852 | n24853 ;
  assign n24855 = n24851 | n24854 ;
  assign n24856 = n24850 | n24855 ;
  assign n24857 = x2 & n24856 ;
  assign n24858 = n24457 | n24833 ;
  assign n24859 = n24846 | n24858 ;
  assign n24860 = ( x2 & n24856 ) | ( x2 & n24859 ) | ( n24856 & n24859 ) ;
  assign n24861 = ~n24857 & n24860 ;
  assign n24862 = ( n24454 & n24848 ) | ( n24454 & n24861 ) | ( n24848 & n24861 ) ;
  assign n24863 = n24444 & n24862 ;
  assign n24864 = n24454 | n24847 ;
  assign n24865 = n24861 | n24864 ;
  assign n24866 = ( ~n23798 & n23808 ) | ( ~n23798 & n24138 ) | ( n23808 & n24138 ) ;
  assign n24867 = ( n23798 & ~n23808 ) | ( n23798 & n24138 ) | ( ~n23808 & n24138 ) ;
  assign n24868 = ( ~n24138 & n24866 ) | ( ~n24138 & n24867 ) | ( n24866 & n24867 ) ;
  assign n24869 = n24865 & n24868 ;
  assign n24870 = ( n24444 & n24863 ) | ( n24444 & n24869 ) | ( n24863 & n24869 ) ;
  assign n24871 = n24434 & n24870 ;
  assign n24872 = n24444 | n24862 ;
  assign n24873 = n24869 | n24872 ;
  assign n24874 = ( ~n23785 & n23795 ) | ( ~n23785 & n24139 ) | ( n23795 & n24139 ) ;
  assign n24875 = ( n23785 & ~n23795 ) | ( n23785 & n24139 ) | ( ~n23795 & n24139 ) ;
  assign n24876 = ( ~n24139 & n24874 ) | ( ~n24139 & n24875 ) | ( n24874 & n24875 ) ;
  assign n24877 = n24873 & n24876 ;
  assign n24878 = ( n24434 & n24871 ) | ( n24434 & n24877 ) | ( n24871 & n24877 ) ;
  assign n24879 = n24423 & n24878 ;
  assign n24880 = n24434 | n24870 ;
  assign n24881 = n24877 | n24880 ;
  assign n24882 = ( ~n23771 & n23782 ) | ( ~n23771 & n24140 ) | ( n23782 & n24140 ) ;
  assign n24883 = ( n23771 & ~n23782 ) | ( n23771 & n24140 ) | ( ~n23782 & n24140 ) ;
  assign n24884 = ( ~n24140 & n24882 ) | ( ~n24140 & n24883 ) | ( n24882 & n24883 ) ;
  assign n24885 = n24881 & n24884 ;
  assign n24886 = ( n24423 & n24879 ) | ( n24423 & n24885 ) | ( n24879 & n24885 ) ;
  assign n24887 = n24421 & n24886 ;
  assign n24888 = n9798 & n20532 ;
  assign n24889 = n9782 & ~n20724 ;
  assign n24890 = n9783 & ~n20536 ;
  assign n24891 = n24889 | n24890 ;
  assign n24892 = n24888 | n24891 ;
  assign n24893 = n9787 | n24892 ;
  assign n24894 = ( n23203 & n24892 ) | ( n23203 & n24893 ) | ( n24892 & n24893 ) ;
  assign n24895 = ~x2 & n24894 ;
  assign n24896 = n24423 | n24878 ;
  assign n24897 = n24885 | n24896 ;
  assign n24898 = ( ~n24894 & n24895 ) | ( ~n24894 & n24897 ) | ( n24895 & n24897 ) ;
  assign n24899 = ( x2 & n24895 ) | ( x2 & n24898 ) | ( n24895 & n24898 ) ;
  assign n24900 = ( n24421 & n24887 ) | ( n24421 & n24899 ) | ( n24887 & n24899 ) ;
  assign n24901 = n24419 & n24900 ;
  assign n24902 = n9798 & n20838 ;
  assign n24903 = n9782 & ~n20536 ;
  assign n24904 = n9783 & n20532 ;
  assign n24905 = n24903 | n24904 ;
  assign n24906 = n24902 | n24905 ;
  assign n24907 = n9787 | n24906 ;
  assign n24908 = ( ~n23712 & n24906 ) | ( ~n23712 & n24907 ) | ( n24906 & n24907 ) ;
  assign n24909 = ~x2 & n24908 ;
  assign n24910 = n24421 | n24886 ;
  assign n24911 = n24899 | n24910 ;
  assign n24912 = ( ~n24908 & n24909 ) | ( ~n24908 & n24911 ) | ( n24909 & n24911 ) ;
  assign n24913 = ( x2 & n24909 ) | ( x2 & n24912 ) | ( n24909 & n24912 ) ;
  assign n24914 = ( n24419 & n24901 ) | ( n24419 & n24913 ) | ( n24901 & n24913 ) ;
  assign n24915 = n24408 & n24914 ;
  assign n24916 = ~n23665 & n23741 ;
  assign n24917 = n23665 & ~n23741 ;
  assign n24918 = n24916 | n24917 ;
  assign n24919 = n24144 & ~n24918 ;
  assign n24920 = n24419 | n24900 ;
  assign n24921 = n24913 | n24920 ;
  assign n24922 = ( n24144 & ~n24918 ) | ( n24144 & n24921 ) | ( ~n24918 & n24921 ) ;
  assign n24923 = ~n24919 & n24922 ;
  assign n24924 = ( n24408 & n24915 ) | ( n24408 & n24923 ) | ( n24915 & n24923 ) ;
  assign n24925 = n24398 & n24924 ;
  assign n24926 = ~n23721 & n23731 ;
  assign n24927 = n23721 & ~n23731 ;
  assign n24928 = n24926 | n24927 ;
  assign n24929 = n24145 | n24928 ;
  assign n24930 = n24408 | n24914 ;
  assign n24931 = n24923 | n24930 ;
  assign n24932 = ( n24145 & ~n24929 ) | ( n24145 & n24931 ) | ( ~n24929 & n24931 ) ;
  assign n24933 = ( n24928 & ~n24929 ) | ( n24928 & n24932 ) | ( ~n24929 & n24932 ) ;
  assign n24934 = ( n24398 & n24925 ) | ( n24398 & n24933 ) | ( n24925 & n24933 ) ;
  assign n24935 = n24398 | n24924 ;
  assign n24936 = n24933 | n24935 ;
  assign n24937 = ( n23717 & ~n23719 ) | ( n23717 & n24146 ) | ( ~n23719 & n24146 ) ;
  assign n24938 = ( ~n23717 & n23719 ) | ( ~n23717 & n24146 ) | ( n23719 & n24146 ) ;
  assign n24939 = ( ~n24146 & n24937 ) | ( ~n24146 & n24938 ) | ( n24937 & n24938 ) ;
  assign n24940 = n24936 & n24939 ;
  assign n24941 = n24934 | n24940 ;
  assign n24942 = n24367 | n24383 ;
  assign n24943 = ( ~n24382 & n24383 ) | ( ~n24382 & n24942 ) | ( n24383 & n24942 ) ;
  assign n24944 = n24941 & ~n24943 ;
  assign n24945 = ( ~n24365 & n24384 ) | ( ~n24365 & n24944 ) | ( n24384 & n24944 ) ;
  assign n24946 = n24365 & ~n24383 ;
  assign n24947 = ~n24944 & n24946 ;
  assign n24948 = n24945 | n24947 ;
  assign n24949 = ~n24941 & n24943 ;
  assign n24950 = n24944 | n24949 ;
  assign n24951 = n24948 | n24950 ;
  assign n24952 = ~n24950 & n24951 ;
  assign n24953 = ( ~n24948 & n24951 ) | ( ~n24948 & n24952 ) | ( n24951 & n24952 ) ;
  assign n24954 = n9245 & n24329 ;
  assign n24955 = n8680 & n20921 ;
  assign n24956 = n8681 & ~n21005 ;
  assign n24957 = n24955 | n24956 ;
  assign n24958 = n24954 | n24957 ;
  assign n24959 = ( n8685 & ~n24391 ) | ( n8685 & n24392 ) | ( ~n24391 & n24392 ) ;
  assign n24960 = n24958 | n24959 ;
  assign n24961 = x5 | n24960 ;
  assign n24962 = ~x5 & n24961 ;
  assign n24963 = ( ~n24960 & n24961 ) | ( ~n24960 & n24962 ) | ( n24961 & n24962 ) ;
  assign n24964 = n23189 | n23193 ;
  assign n24965 = n7305 & ~n20724 ;
  assign n24966 = n7300 & n20546 ;
  assign n24967 = n7302 & ~n20542 ;
  assign n24968 = n24966 | n24967 ;
  assign n24969 = n24965 | n24968 ;
  assign n24970 = n7308 | n24969 ;
  assign n24971 = ( n23229 & n24969 ) | ( n23229 & n24970 ) | ( n24969 & n24970 ) ;
  assign n24972 = x11 & n24971 ;
  assign n24973 = x11 & ~n24972 ;
  assign n24974 = ( n24971 & ~n24972 ) | ( n24971 & n24973 ) | ( ~n24972 & n24973 ) ;
  assign n24975 = n23182 | n23185 ;
  assign n24976 = n7280 & ~n20710 ;
  assign n24977 = n5384 & ~n20552 ;
  assign n24978 = n7277 & n20556 ;
  assign n24979 = n24977 | n24978 ;
  assign n24980 = n24976 | n24979 ;
  assign n24981 = n39 | n24980 ;
  assign n24982 = ( ~n22641 & n24980 ) | ( ~n22641 & n24981 ) | ( n24980 & n24981 ) ;
  assign n24983 = ~x14 & n24982 ;
  assign n24984 = x14 | n24983 ;
  assign n24985 = ( ~n24982 & n24983 ) | ( ~n24982 & n24984 ) | ( n24983 & n24984 ) ;
  assign n24986 = n23176 | n23180 ;
  assign n24987 = n5083 & n20562 ;
  assign n24988 = n5069 & ~n20689 ;
  assign n24989 = n5070 & n20560 ;
  assign n24990 = n24988 | n24989 ;
  assign n24991 = n24987 | n24990 ;
  assign n24992 = n5074 | n24991 ;
  assign n24993 = ( ~n21044 & n24991 ) | ( ~n21044 & n24992 ) | ( n24991 & n24992 ) ;
  assign n24994 = ~x17 & n24993 ;
  assign n24995 = x17 | n24994 ;
  assign n24996 = ( ~n24993 & n24994 ) | ( ~n24993 & n24995 ) | ( n24994 & n24995 ) ;
  assign n24997 = n23169 | n23172 ;
  assign n24998 = n4781 & ~n20573 ;
  assign n24999 = n4776 & ~n20584 ;
  assign n25000 = n4778 & ~n20569 ;
  assign n25001 = n24999 | n25000 ;
  assign n25002 = n24998 | n25001 ;
  assign n25003 = n4784 | n25002 ;
  assign n25004 = ( ~n21860 & n25002 ) | ( ~n21860 & n25003 ) | ( n25002 & n25003 ) ;
  assign n25005 = ~x20 & n25004 ;
  assign n25006 = x20 | n25005 ;
  assign n25007 = ( ~n25004 & n25005 ) | ( ~n25004 & n25006 ) | ( n25005 & n25006 ) ;
  assign n25008 = n23163 | n23167 ;
  assign n25009 = n4551 & ~n20580 ;
  assign n25010 = n4546 & ~n20591 ;
  assign n25011 = n4548 & n20588 ;
  assign n25012 = n25010 | n25011 ;
  assign n25013 = n25009 | n25012 ;
  assign n25014 = n4554 | n25013 ;
  assign n25015 = ( n21840 & n25013 ) | ( n21840 & n25014 ) | ( n25013 & n25014 ) ;
  assign n25016 = x23 & n25015 ;
  assign n25017 = x23 & ~n25016 ;
  assign n25018 = ( n25015 & ~n25016 ) | ( n25015 & n25017 ) | ( ~n25016 & n25017 ) ;
  assign n25019 = n23156 | n23159 ;
  assign n25020 = n4484 & ~n20595 ;
  assign n25021 = n4479 & ~n20605 ;
  assign n25022 = n4481 & n20600 ;
  assign n25023 = n25021 | n25022 ;
  assign n25024 = n25020 | n25023 ;
  assign n25025 = n4487 | n25024 ;
  assign n25026 = ( ~n21554 & n25024 ) | ( ~n21554 & n25025 ) | ( n25024 & n25025 ) ;
  assign n25027 = ~x26 & n25026 ;
  assign n25028 = x26 | n25027 ;
  assign n25029 = ( ~n25026 & n25027 ) | ( ~n25026 & n25028 ) | ( n25027 & n25028 ) ;
  assign n25030 = n23150 | n23154 ;
  assign n25031 = n23142 | n23146 ;
  assign n25032 = n3744 & n20619 ;
  assign n25033 = n3727 & n20622 ;
  assign n25034 = n3639 & ~n20625 ;
  assign n25035 = n25033 | n25034 ;
  assign n25036 = n25032 | n25035 ;
  assign n25037 = n3636 | n25036 ;
  assign n25038 = ( ~n21056 & n25036 ) | ( ~n21056 & n25037 ) | ( n25036 & n25037 ) ;
  assign n25039 = n818 | n1575 ;
  assign n25040 = n1894 | n25039 ;
  assign n25041 = n5535 | n25040 ;
  assign n25042 = n5647 | n25041 ;
  assign n25043 = n12631 | n25042 ;
  assign n25044 = n971 | n25043 ;
  assign n25045 = n760 | n1613 ;
  assign n25046 = n430 | n25045 ;
  assign n25047 = n1522 | n25046 ;
  assign n25048 = n2361 | n25047 ;
  assign n25049 = n25044 | n25048 ;
  assign n25050 = n431 | n2943 ;
  assign n25051 = n409 | n25050 ;
  assign n25052 = n670 | n25051 ;
  assign n25053 = n226 & ~n25052 ;
  assign n25054 = ~n434 & n25053 ;
  assign n25055 = ~n157 & n25054 ;
  assign n25056 = ~n25049 & n25055 ;
  assign n25057 = n25038 & ~n25056 ;
  assign n25058 = n25038 & ~n25057 ;
  assign n25059 = n25038 | n25056 ;
  assign n25060 = ~n25058 & n25059 ;
  assign n25061 = n25031 & ~n25060 ;
  assign n25062 = n25031 & ~n25061 ;
  assign n25063 = n25060 | n25061 ;
  assign n25064 = ~n25062 & n25063 ;
  assign n25065 = n4048 & n20611 ;
  assign n25066 = n4043 & n20616 ;
  assign n25067 = n4045 & n20614 ;
  assign n25068 = n25066 | n25067 ;
  assign n25069 = n25065 | n25068 ;
  assign n25070 = n4051 | n25069 ;
  assign n25071 = ( n21293 & n25069 ) | ( n21293 & n25070 ) | ( n25069 & n25070 ) ;
  assign n25072 = x29 & n25071 ;
  assign n25073 = x29 & ~n25072 ;
  assign n25074 = ( n25071 & ~n25072 ) | ( n25071 & n25073 ) | ( ~n25072 & n25073 ) ;
  assign n25075 = ~n25064 & n25074 ;
  assign n25076 = n25064 & ~n25074 ;
  assign n25077 = n25075 | n25076 ;
  assign n25078 = n25030 & ~n25077 ;
  assign n25079 = ~n25030 & n25077 ;
  assign n25080 = n25078 | n25079 ;
  assign n25081 = n25029 & ~n25080 ;
  assign n25082 = n25080 | n25081 ;
  assign n25083 = ( ~n25029 & n25081 ) | ( ~n25029 & n25082 ) | ( n25081 & n25082 ) ;
  assign n25084 = n25019 & ~n25083 ;
  assign n25085 = n25019 & ~n25084 ;
  assign n25086 = n25083 | n25084 ;
  assign n25087 = ~n25085 & n25086 ;
  assign n25088 = n25018 & ~n25087 ;
  assign n25089 = n25087 | n25088 ;
  assign n25090 = ( ~n25018 & n25088 ) | ( ~n25018 & n25089 ) | ( n25088 & n25089 ) ;
  assign n25091 = ~n25008 & n25090 ;
  assign n25092 = n25008 & ~n25090 ;
  assign n25093 = n25091 | n25092 ;
  assign n25094 = n25007 & ~n25093 ;
  assign n25095 = n25093 | n25094 ;
  assign n25096 = ( ~n25007 & n25094 ) | ( ~n25007 & n25095 ) | ( n25094 & n25095 ) ;
  assign n25097 = n24997 & ~n25096 ;
  assign n25098 = n24997 & ~n25097 ;
  assign n25099 = n25096 | n25097 ;
  assign n25100 = ~n25098 & n25099 ;
  assign n25101 = n24996 & ~n25100 ;
  assign n25102 = n25100 | n25101 ;
  assign n25103 = ( ~n24996 & n25101 ) | ( ~n24996 & n25102 ) | ( n25101 & n25102 ) ;
  assign n25104 = ~n24986 & n25103 ;
  assign n25105 = n24986 & ~n25103 ;
  assign n25106 = n25104 | n25105 ;
  assign n25107 = n24985 & ~n25106 ;
  assign n25108 = n25106 | n25107 ;
  assign n25109 = ( ~n24985 & n25107 ) | ( ~n24985 & n25108 ) | ( n25107 & n25108 ) ;
  assign n25110 = n24975 & ~n25109 ;
  assign n25111 = n24975 & ~n25110 ;
  assign n25112 = n25109 | n25110 ;
  assign n25113 = ~n25111 & n25112 ;
  assign n25114 = n24974 & ~n25113 ;
  assign n25115 = n25113 | n25114 ;
  assign n25116 = ( ~n24974 & n25114 ) | ( ~n24974 & n25115 ) | ( n25114 & n25115 ) ;
  assign n25117 = ~n24964 & n25116 ;
  assign n25118 = n24964 & ~n25116 ;
  assign n25119 = n25117 | n25118 ;
  assign n25120 = n5503 & n20838 ;
  assign n25121 = n5512 & ~n20536 ;
  assign n25122 = n5508 & n20532 ;
  assign n25123 = n25121 | n25122 ;
  assign n25124 = n25120 | n25123 ;
  assign n25125 = n5515 | n25124 ;
  assign n25126 = ( ~n23712 & n25124 ) | ( ~n23712 & n25125 ) | ( n25124 & n25125 ) ;
  assign n25127 = ~x8 & n25126 ;
  assign n25128 = x8 | n25127 ;
  assign n25129 = ( ~n25126 & n25127 ) | ( ~n25126 & n25128 ) | ( n25127 & n25128 ) ;
  assign n25130 = ( n23681 & n25119 ) | ( n23681 & ~n25129 ) | ( n25119 & ~n25129 ) ;
  assign n25131 = ( ~n25119 & n25129 ) | ( ~n25119 & n25130 ) | ( n25129 & n25130 ) ;
  assign n25132 = ( ~n23681 & n25130 ) | ( ~n23681 & n25131 ) | ( n25130 & n25131 ) ;
  assign n25133 = n24963 & ~n25132 ;
  assign n25134 = ~n24963 & n25132 ;
  assign n25135 = n25133 | n25134 ;
  assign n25136 = n23683 | n24151 ;
  assign n25137 = n25135 & ~n25136 ;
  assign n25138 = ~n25135 & n25136 ;
  assign n25139 = n25137 | n25138 ;
  assign n25140 = n24157 & n24186 ;
  assign n25141 = n24183 & ~n25140 ;
  assign n25142 = ( ~n3636 & n24185 ) | ( ~n3636 & n25141 ) | ( n24185 & n25141 ) ;
  assign n25143 = ( n13544 & n25141 ) | ( n13544 & n25142 ) | ( n25141 & n25142 ) ;
  assign n25144 = n189 | n3633 ;
  assign n25145 = ~n24182 & n25144 ;
  assign n25146 = n24182 & ~n25144 ;
  assign n25147 = n25142 | n25146 ;
  assign n25148 = n25145 | n25147 ;
  assign n25149 = n25141 | n25146 ;
  assign n25150 = n25145 | n25149 ;
  assign n25151 = ( n13544 & n25148 ) | ( n13544 & n25150 ) | ( n25148 & n25150 ) ;
  assign n25152 = ~n25143 & n25151 ;
  assign n25153 = ~n25146 & n25151 ;
  assign n25154 = ~n25145 & n25153 ;
  assign n25155 = n25152 | n25154 ;
  assign n25156 = n4045 | n4048 ;
  assign n25157 = ~n12314 & n25156 ;
  assign n25158 = n4043 | n25157 ;
  assign n25159 = ( ~n12318 & n25157 ) | ( ~n12318 & n25158 ) | ( n25157 & n25158 ) ;
  assign n25160 = n4051 & ~n17966 ;
  assign n25161 = n25159 | n25160 ;
  assign n25162 = x29 & ~n25161 ;
  assign n25163 = ~x29 & n25161 ;
  assign n25164 = n25162 | n25163 ;
  assign n25165 = n3639 & ~n12325 ;
  assign n25166 = n3727 & ~n12328 ;
  assign n25167 = n25165 | n25166 ;
  assign n25168 = n3744 & n12608 ;
  assign n25169 = n25167 | n25168 ;
  assign n25170 = n3636 & n13570 ;
  assign n25171 = ( n3636 & n13568 ) | ( n3636 & n25170 ) | ( n13568 & n25170 ) ;
  assign n25172 = n25169 | n25171 ;
  assign n25173 = n25164 & n25172 ;
  assign n25174 = n25164 & ~n25173 ;
  assign n25175 = n25172 & ~n25173 ;
  assign n25176 = n25174 | n25175 ;
  assign n25177 = n25155 & ~n25176 ;
  assign n25178 = ~n25155 & n25176 ;
  assign n25179 = n25177 | n25178 ;
  assign n25180 = n24226 | n24238 ;
  assign n25181 = n25179 & n25180 ;
  assign n25182 = n25179 | n25180 ;
  assign n25183 = ~n25181 & n25182 ;
  assign n25184 = n24271 | n24321 ;
  assign n25185 = n25183 & n25184 ;
  assign n25186 = n25183 | n25184 ;
  assign n25187 = ~n25185 & n25186 ;
  assign n25188 = n24324 | n25187 ;
  assign n25189 = n24324 & n25187 ;
  assign n25190 = n25188 & ~n25189 ;
  assign n25191 = n24352 | n25190 ;
  assign n25192 = n24352 & n25190 ;
  assign n25193 = n25191 & ~n25192 ;
  assign n25194 = n9798 & n25187 ;
  assign n25195 = n9782 & ~n24334 ;
  assign n25196 = n9783 & n24324 ;
  assign n25197 = n25195 | n25196 ;
  assign n25198 = n25194 | n25197 ;
  assign n25199 = n9787 | n25198 ;
  assign n25200 = ( n25193 & n25198 ) | ( n25193 & n25199 ) | ( n25198 & n25199 ) ;
  assign n25201 = x2 & n25200 ;
  assign n25202 = x2 & ~n25201 ;
  assign n25203 = ( n25200 & ~n25201 ) | ( n25200 & n25202 ) | ( ~n25201 & n25202 ) ;
  assign n25204 = ~n25139 & n25203 ;
  assign n25205 = n25139 & ~n25203 ;
  assign n25206 = n25204 | n25205 ;
  assign n25207 = n24363 | n24384 ;
  assign n25208 = ( ~n24364 & n24944 ) | ( ~n24364 & n25207 ) | ( n24944 & n25207 ) ;
  assign n25209 = n25206 & ~n25208 ;
  assign n25210 = ~n25206 & n25208 ;
  assign n25211 = n25209 | n25210 ;
  assign n25212 = n24951 | n25211 ;
  assign n25213 = n24951 & n25211 ;
  assign n25214 = n25212 & ~n25213 ;
  assign n25215 = n9245 & ~n24334 ;
  assign n25216 = n8680 & ~n21005 ;
  assign n25217 = n8681 & n24329 ;
  assign n25218 = n25216 | n25217 ;
  assign n25219 = n25215 | n25218 ;
  assign n25220 = ( n8685 & ~n24373 ) | ( n8685 & n24376 ) | ( ~n24373 & n24376 ) ;
  assign n25221 = n25219 | n25220 ;
  assign n25222 = x5 | n25221 ;
  assign n25223 = ~x5 & n25222 ;
  assign n25224 = ( ~n25221 & n25222 ) | ( ~n25221 & n25223 ) | ( n25222 & n25223 ) ;
  assign n25225 = n5503 & n20921 ;
  assign n25226 = n5512 & n20532 ;
  assign n25227 = n5508 & n20838 ;
  assign n25228 = n25226 | n25227 ;
  assign n25229 = n25225 | n25228 ;
  assign n25230 = n5515 & ~n23691 ;
  assign n25231 = ~n23695 & n25230 ;
  assign n25232 = ( n5515 & n25229 ) | ( n5515 & ~n25231 ) | ( n25229 & ~n25231 ) ;
  assign n25233 = ~x8 & n25232 ;
  assign n25234 = x8 | n25233 ;
  assign n25235 = ( ~n25232 & n25233 ) | ( ~n25232 & n25234 ) | ( n25233 & n25234 ) ;
  assign n25236 = n25107 | n25110 ;
  assign n25237 = n25094 | n25097 ;
  assign n25238 = n25088 | n25092 ;
  assign n25239 = n4551 & ~n20584 ;
  assign n25240 = n4546 & n20588 ;
  assign n25241 = n4548 & ~n20580 ;
  assign n25242 = n25240 | n25241 ;
  assign n25243 = n25239 | n25242 ;
  assign n25244 = n4554 | n25243 ;
  assign n25245 = ( ~n21901 & n25243 ) | ( ~n21901 & n25244 ) | ( n25243 & n25244 ) ;
  assign n25246 = ~x23 & n25245 ;
  assign n25247 = x23 | n25246 ;
  assign n25248 = ( ~n25245 & n25246 ) | ( ~n25245 & n25247 ) | ( n25246 & n25247 ) ;
  assign n25249 = n4484 & ~n20591 ;
  assign n25250 = n4479 & n20600 ;
  assign n25251 = n4481 & ~n20595 ;
  assign n25252 = n25250 | n25251 ;
  assign n25253 = n25249 | n25252 ;
  assign n25254 = n4487 & ~n21539 ;
  assign n25255 = ~n21543 & n25254 ;
  assign n25256 = ( n4487 & n25253 ) | ( n4487 & ~n25255 ) | ( n25253 & ~n25255 ) ;
  assign n25257 = ~x26 & n25256 ;
  assign n25258 = x26 | n25257 ;
  assign n25259 = ( ~n25256 & n25257 ) | ( ~n25256 & n25258 ) | ( n25257 & n25258 ) ;
  assign n25260 = n25081 | n25084 ;
  assign n25261 = n25057 | n25061 ;
  assign n25262 = n3744 & n20616 ;
  assign n25263 = n3727 & n20619 ;
  assign n25264 = n3639 & n20622 ;
  assign n25265 = n25263 | n25264 ;
  assign n25266 = n25262 | n25265 ;
  assign n25267 = n3636 | n25266 ;
  assign n25268 = ( n21190 & n25266 ) | ( n21190 & n25267 ) | ( n25266 & n25267 ) ;
  assign n25269 = n435 | n12683 ;
  assign n25270 = n12992 | n25269 ;
  assign n25271 = n2315 | n5671 ;
  assign n25272 = n25270 | n25271 ;
  assign n25273 = n1222 | n25272 ;
  assign n25274 = n11389 | n25273 ;
  assign n25275 = n11385 | n25274 ;
  assign n25276 = n4858 | n25275 ;
  assign n25277 = n1560 | n25276 ;
  assign n25278 = n756 | n2807 ;
  assign n25279 = n1865 | n25278 ;
  assign n25280 = n352 | n25279 ;
  assign n25281 = n806 | n25280 ;
  assign n25282 = n260 | n25281 ;
  assign n25283 = n25277 | n25282 ;
  assign n25284 = n379 | n596 ;
  assign n25285 = n595 | n25284 ;
  assign n25286 = n164 | n25285 ;
  assign n25287 = n25283 | n25286 ;
  assign n25288 = n25268 & n25287 ;
  assign n25289 = n25268 & ~n25288 ;
  assign n25290 = ~n25268 & n25287 ;
  assign n25291 = n25289 | n25290 ;
  assign n25292 = n25261 & n25291 ;
  assign n25293 = n25261 & ~n25292 ;
  assign n25294 = n25291 & ~n25292 ;
  assign n25295 = n25293 | n25294 ;
  assign n25296 = n4048 & ~n20605 ;
  assign n25297 = n4043 & n20614 ;
  assign n25298 = n4045 & n20611 ;
  assign n25299 = n25297 | n25298 ;
  assign n25300 = n25296 | n25299 ;
  assign n25301 = n4051 | n25300 ;
  assign n25302 = ( ~n21275 & n25300 ) | ( ~n21275 & n25301 ) | ( n25300 & n25301 ) ;
  assign n25303 = ~x29 & n25302 ;
  assign n25304 = x29 | n25303 ;
  assign n25305 = ( ~n25302 & n25303 ) | ( ~n25302 & n25304 ) | ( n25303 & n25304 ) ;
  assign n25306 = n25295 & n25305 ;
  assign n25307 = n25295 | n25305 ;
  assign n25308 = ~n25306 & n25307 ;
  assign n25309 = n25075 | n25078 ;
  assign n25310 = n25308 & n25309 ;
  assign n25311 = n25308 | n25309 ;
  assign n25312 = ~n25310 & n25311 ;
  assign n25313 = ( n25259 & n25260 ) | ( n25259 & ~n25312 ) | ( n25260 & ~n25312 ) ;
  assign n25314 = ( ~n25260 & n25312 ) | ( ~n25260 & n25313 ) | ( n25312 & n25313 ) ;
  assign n25315 = ( ~n25259 & n25313 ) | ( ~n25259 & n25314 ) | ( n25313 & n25314 ) ;
  assign n25316 = n25248 & n25315 ;
  assign n25317 = n25248 | n25315 ;
  assign n25318 = ~n25316 & n25317 ;
  assign n25319 = n25238 | n25318 ;
  assign n25320 = n25238 & n25318 ;
  assign n25321 = n25319 & ~n25320 ;
  assign n25322 = n4781 & ~n20689 ;
  assign n25323 = n4776 & ~n20569 ;
  assign n25324 = n4778 & ~n20573 ;
  assign n25325 = n25323 | n25324 ;
  assign n25326 = n25322 | n25325 ;
  assign n25327 = n4784 & ~n22193 ;
  assign n25328 = n22192 & n25327 ;
  assign n25329 = ( n4784 & n25326 ) | ( n4784 & ~n25328 ) | ( n25326 & ~n25328 ) ;
  assign n25330 = x20 & n25329 ;
  assign n25331 = x20 & ~n25330 ;
  assign n25332 = ( n25329 & ~n25330 ) | ( n25329 & n25331 ) | ( ~n25330 & n25331 ) ;
  assign n25333 = n25321 & n25332 ;
  assign n25334 = n25321 & ~n25333 ;
  assign n25335 = ~n25321 & n25332 ;
  assign n25336 = n25334 | n25335 ;
  assign n25337 = n25237 & n25336 ;
  assign n25338 = n25237 & ~n25337 ;
  assign n25339 = n25336 & ~n25337 ;
  assign n25340 = n25338 | n25339 ;
  assign n25341 = n5083 & ~n20552 ;
  assign n25342 = n5069 & n20560 ;
  assign n25343 = n5070 & n20562 ;
  assign n25344 = n25342 | n25343 ;
  assign n25345 = n25341 | n25344 ;
  assign n25346 = n5074 & ~n22510 ;
  assign n25347 = ( n5074 & n22512 ) | ( n5074 & n25346 ) | ( n22512 & n25346 ) ;
  assign n25348 = n25345 | n25347 ;
  assign n25349 = x17 | n25348 ;
  assign n25350 = ~x17 & n25349 ;
  assign n25351 = ( ~n25348 & n25349 ) | ( ~n25348 & n25350 ) | ( n25349 & n25350 ) ;
  assign n25352 = n25340 & n25351 ;
  assign n25353 = n25340 & ~n25352 ;
  assign n25354 = ~n25340 & n25351 ;
  assign n25355 = n25353 | n25354 ;
  assign n25356 = n25101 | n25105 ;
  assign n25357 = n25355 | n25356 ;
  assign n25358 = n25355 & n25356 ;
  assign n25359 = n25357 & ~n25358 ;
  assign n25360 = n7280 & n20546 ;
  assign n25361 = n5384 & n20556 ;
  assign n25362 = n7277 & ~n20710 ;
  assign n25363 = n25361 | n25362 ;
  assign n25364 = n25360 | n25363 ;
  assign n25365 = n39 & n21031 ;
  assign n25366 = ~n21037 & n25365 ;
  assign n25367 = ( n39 & n25364 ) | ( n39 & ~n25366 ) | ( n25364 & ~n25366 ) ;
  assign n25368 = x14 & n25367 ;
  assign n25369 = x14 & ~n25368 ;
  assign n25370 = ( n25367 & ~n25368 ) | ( n25367 & n25369 ) | ( ~n25368 & n25369 ) ;
  assign n25371 = n25359 & n25370 ;
  assign n25372 = n25359 & ~n25371 ;
  assign n25373 = ~n25359 & n25370 ;
  assign n25374 = n25372 | n25373 ;
  assign n25375 = n25236 & n25374 ;
  assign n25376 = n25236 & ~n25375 ;
  assign n25377 = n25374 & ~n25375 ;
  assign n25378 = n25376 | n25377 ;
  assign n25379 = n7305 & ~n20536 ;
  assign n25380 = n7300 & ~n20542 ;
  assign n25381 = n7302 & ~n20724 ;
  assign n25382 = n25380 | n25381 ;
  assign n25383 = n25379 | n25382 ;
  assign n25384 = ( n7308 & n23213 ) | ( n7308 & ~n23217 ) | ( n23213 & ~n23217 ) ;
  assign n25385 = n25383 | n25384 ;
  assign n25386 = x11 | n25385 ;
  assign n25387 = ~x11 & n25386 ;
  assign n25388 = ( ~n25385 & n25386 ) | ( ~n25385 & n25387 ) | ( n25386 & n25387 ) ;
  assign n25389 = n25378 & n25388 ;
  assign n25390 = n25378 & ~n25389 ;
  assign n25391 = ~n25378 & n25388 ;
  assign n25392 = n25390 | n25391 ;
  assign n25393 = n25114 | n25118 ;
  assign n25394 = n25392 | n25393 ;
  assign n25395 = n25392 & n25393 ;
  assign n25396 = n25394 & ~n25395 ;
  assign n25397 = ( n25131 & n25235 ) | ( n25131 & n25396 ) | ( n25235 & n25396 ) ;
  assign n25398 = ( n25131 & n25396 ) | ( n25131 & ~n25397 ) | ( n25396 & ~n25397 ) ;
  assign n25399 = ( n25235 & ~n25397 ) | ( n25235 & n25398 ) | ( ~n25397 & n25398 ) ;
  assign n25400 = n25224 & n25399 ;
  assign n25401 = n25224 | n25399 ;
  assign n25402 = ~n25400 & n25401 ;
  assign n25403 = n25133 | n25138 ;
  assign n25404 = n25402 | n25403 ;
  assign n25405 = n25402 & n25403 ;
  assign n25406 = n25404 & ~n25405 ;
  assign n25407 = ( n25173 & n25176 ) | ( n25173 & ~n25178 ) | ( n25176 & ~n25178 ) ;
  assign n25408 = n3744 & ~n12318 ;
  assign n25409 = n3639 & ~n12328 ;
  assign n25410 = n3727 & n12608 ;
  assign n25411 = n25409 | n25410 ;
  assign n25412 = n25408 | n25411 ;
  assign n25413 = n3636 | n25412 ;
  assign n25414 = ( n14320 & n25412 ) | ( n14320 & n25413 ) | ( n25412 & n25413 ) ;
  assign n25415 = n12285 & n25144 ;
  assign n25416 = ( n12277 & n25144 ) | ( n12277 & n25415 ) | ( n25144 & n25415 ) ;
  assign n25417 = n12285 | n25144 ;
  assign n25418 = n12277 | n25417 ;
  assign n25419 = ~n25416 & n25418 ;
  assign n25420 = n4041 | n4045 ;
  assign n25421 = n4043 | n25420 ;
  assign n25422 = ~n12314 & n25421 ;
  assign n25423 = ~x29 & n25422 ;
  assign n25424 = x29 | n25423 ;
  assign n25425 = ( ~n25422 & n25423 ) | ( ~n25422 & n25424 ) | ( n25423 & n25424 ) ;
  assign n25426 = n25419 & ~n25425 ;
  assign n25427 = ~n25419 & n25425 ;
  assign n25428 = n25426 | n25427 ;
  assign n25429 = n25414 & ~n25428 ;
  assign n25430 = n25414 & ~n25429 ;
  assign n25431 = n25414 | n25428 ;
  assign n25432 = ( n25153 & ~n25430 ) | ( n25153 & n25431 ) | ( ~n25430 & n25431 ) ;
  assign n25433 = ( n25153 & n25431 ) | ( n25153 & ~n25432 ) | ( n25431 & ~n25432 ) ;
  assign n25434 = ( n25430 & n25432 ) | ( n25430 & ~n25433 ) | ( n25432 & ~n25433 ) ;
  assign n25435 = n25407 & n25434 ;
  assign n25436 = n25407 | n25434 ;
  assign n25437 = ~n25435 & n25436 ;
  assign n25438 = n25181 & n25437 ;
  assign n25439 = ( n25185 & n25437 ) | ( n25185 & n25438 ) | ( n25437 & n25438 ) ;
  assign n25440 = n25181 | n25437 ;
  assign n25441 = n25185 | n25440 ;
  assign n25442 = ~n25439 & n25441 ;
  assign n25443 = n9798 & n25442 ;
  assign n25444 = n9782 & n24324 ;
  assign n25445 = n9783 & n25187 ;
  assign n25446 = n25444 | n25445 ;
  assign n25447 = n25443 | n25446 ;
  assign n25448 = n9787 | n25447 ;
  assign n25449 = n25189 | n25192 ;
  assign n25450 = ( n25187 & ~n25442 ) | ( n25187 & n25449 ) | ( ~n25442 & n25449 ) ;
  assign n25451 = ( ~n25187 & n25442 ) | ( ~n25187 & n25450 ) | ( n25442 & n25450 ) ;
  assign n25452 = ( ~n25449 & n25450 ) | ( ~n25449 & n25451 ) | ( n25450 & n25451 ) ;
  assign n25453 = ( n25447 & n25448 ) | ( n25447 & n25452 ) | ( n25448 & n25452 ) ;
  assign n25454 = x2 & n25453 ;
  assign n25455 = x2 & ~n25454 ;
  assign n25456 = ( n25453 & ~n25454 ) | ( n25453 & n25455 ) | ( ~n25454 & n25455 ) ;
  assign n25457 = n25406 & n25456 ;
  assign n25458 = n25406 | n25456 ;
  assign n25459 = ~n25457 & n25458 ;
  assign n25460 = n25204 | n25210 ;
  assign n25461 = n25459 & n25460 ;
  assign n25462 = n25459 | n25460 ;
  assign n25463 = ~n25461 & n25462 ;
  assign n25464 = ~n25212 & n25463 ;
  assign n25465 = n25212 & ~n25463 ;
  assign n25466 = n25464 | n25465 ;
  assign n25467 = n5503 & ~n21005 ;
  assign n25468 = n5512 & n20838 ;
  assign n25469 = n5508 & n20921 ;
  assign n25470 = n25468 | n25469 ;
  assign n25471 = n25467 | n25470 ;
  assign n25472 = n5515 | n25471 ;
  assign n25473 = ( ~n21015 & n25471 ) | ( ~n21015 & n25472 ) | ( n25471 & n25472 ) ;
  assign n25474 = ~x8 & n25473 ;
  assign n25475 = x8 | n25474 ;
  assign n25476 = ( ~n25473 & n25474 ) | ( ~n25473 & n25475 ) | ( n25474 & n25475 ) ;
  assign n25477 = n25389 | n25395 ;
  assign n25478 = n7305 & n20532 ;
  assign n25479 = n7300 & ~n20724 ;
  assign n25480 = n7302 & ~n20536 ;
  assign n25481 = n25479 | n25480 ;
  assign n25482 = n25478 | n25481 ;
  assign n25483 = n7308 | n25482 ;
  assign n25484 = ( n23203 & n25482 ) | ( n23203 & n25483 ) | ( n25482 & n25483 ) ;
  assign n25485 = x11 & n25484 ;
  assign n25486 = x11 & ~n25485 ;
  assign n25487 = ( n25484 & ~n25485 ) | ( n25484 & n25486 ) | ( ~n25485 & n25486 ) ;
  assign n25488 = n25371 | n25375 ;
  assign n25489 = n7280 & ~n20542 ;
  assign n25490 = n5384 & ~n20710 ;
  assign n25491 = n7277 & n20546 ;
  assign n25492 = n25490 | n25491 ;
  assign n25493 = n25489 | n25492 ;
  assign n25494 = n39 | n25493 ;
  assign n25495 = ( ~n23042 & n25493 ) | ( ~n23042 & n25494 ) | ( n25493 & n25494 ) ;
  assign n25496 = ~x14 & n25495 ;
  assign n25497 = x14 | n25496 ;
  assign n25498 = ( ~n25495 & n25496 ) | ( ~n25495 & n25497 ) | ( n25496 & n25497 ) ;
  assign n25499 = n25352 | n25358 ;
  assign n25500 = n5083 & n20556 ;
  assign n25501 = n5069 & n20562 ;
  assign n25502 = n5070 & ~n20552 ;
  assign n25503 = n25501 | n25502 ;
  assign n25504 = n25500 | n25503 ;
  assign n25505 = n5074 | n25504 ;
  assign n25506 = ( ~n22655 & n25504 ) | ( ~n22655 & n25505 ) | ( n25504 & n25505 ) ;
  assign n25507 = ~x17 & n25506 ;
  assign n25508 = x17 | n25507 ;
  assign n25509 = ( ~n25506 & n25507 ) | ( ~n25506 & n25508 ) | ( n25507 & n25508 ) ;
  assign n25510 = n4781 & n20560 ;
  assign n25511 = n4776 & ~n20573 ;
  assign n25512 = n4778 & ~n20689 ;
  assign n25513 = n25511 | n25512 ;
  assign n25514 = n25510 | n25513 ;
  assign n25515 = n4784 & ~n22176 ;
  assign n25516 = ~n22173 & n25515 ;
  assign n25517 = ( n4784 & n25514 ) | ( n4784 & ~n25516 ) | ( n25514 & ~n25516 ) ;
  assign n25518 = ~x20 & n25517 ;
  assign n25519 = x20 | n25518 ;
  assign n25520 = ( ~n25517 & n25518 ) | ( ~n25517 & n25519 ) | ( n25518 & n25519 ) ;
  assign n25521 = n25333 | n25337 ;
  assign n25522 = ( n25259 & n25260 ) | ( n25259 & n25312 ) | ( n25260 & n25312 ) ;
  assign n25523 = n4484 & n20588 ;
  assign n25524 = n4479 & ~n20595 ;
  assign n25525 = n4481 & ~n20591 ;
  assign n25526 = n25524 | n25525 ;
  assign n25527 = n25523 | n25526 ;
  assign n25528 = n4487 | n25527 ;
  assign n25529 = ( n21526 & n25527 ) | ( n21526 & n25528 ) | ( n25527 & n25528 ) ;
  assign n25530 = x26 & n25529 ;
  assign n25531 = x26 & ~n25530 ;
  assign n25532 = ( n25529 & ~n25530 ) | ( n25529 & n25531 ) | ( ~n25530 & n25531 ) ;
  assign n25533 = n25288 | n25292 ;
  assign n25534 = n3744 & n20614 ;
  assign n25535 = n3727 & n20616 ;
  assign n25536 = n3639 & n20619 ;
  assign n25537 = n25535 | n25536 ;
  assign n25538 = n25534 | n25537 ;
  assign n25539 = n3636 | n25538 ;
  assign n25540 = ( n21302 & n25538 ) | ( n21302 & n25539 ) | ( n25538 & n25539 ) ;
  assign n25541 = n2118 | n5640 ;
  assign n25542 = n697 | n958 ;
  assign n25543 = n251 | n25542 ;
  assign n25544 = n1675 | n1689 ;
  assign n25545 = n25543 | n25544 ;
  assign n25546 = n2315 | n3844 ;
  assign n25547 = n25545 | n25546 ;
  assign n25548 = ( n5688 & n13807 ) | ( n5688 & n25547 ) | ( n13807 & n25547 ) ;
  assign n25549 = n5688 & ~n25548 ;
  assign n25550 = ~n25541 & n25549 ;
  assign n25551 = n732 | n2163 ;
  assign n25552 = n1336 | n25551 ;
  assign n25553 = n608 | n25552 ;
  assign n25554 = n100 | n25553 ;
  assign n25555 = n25550 & ~n25554 ;
  assign n25556 = n25540 & ~n25555 ;
  assign n25557 = n25540 & ~n25556 ;
  assign n25558 = n25540 | n25555 ;
  assign n25559 = ~n25557 & n25558 ;
  assign n25560 = n25533 & ~n25559 ;
  assign n25561 = n25533 & ~n25560 ;
  assign n25562 = n25559 | n25560 ;
  assign n25563 = ~n25561 & n25562 ;
  assign n25564 = n4048 & n20600 ;
  assign n25565 = n4043 & n20611 ;
  assign n25566 = n4045 & ~n20605 ;
  assign n25567 = n25565 | n25566 ;
  assign n25568 = n25564 | n25567 ;
  assign n25569 = n4051 | n25568 ;
  assign n25570 = ( ~n21432 & n25568 ) | ( ~n21432 & n25569 ) | ( n25568 & n25569 ) ;
  assign n25571 = ~x29 & n25570 ;
  assign n25572 = x29 | n25571 ;
  assign n25573 = ( ~n25570 & n25571 ) | ( ~n25570 & n25572 ) | ( n25571 & n25572 ) ;
  assign n25574 = ~n25563 & n25573 ;
  assign n25575 = n25563 & ~n25573 ;
  assign n25576 = n25574 | n25575 ;
  assign n25577 = n25306 | n25310 ;
  assign n25578 = ~n25576 & n25577 ;
  assign n25579 = n25576 & ~n25577 ;
  assign n25580 = n25578 | n25579 ;
  assign n25581 = n25532 & ~n25580 ;
  assign n25582 = n25580 | n25581 ;
  assign n25583 = ( ~n25532 & n25581 ) | ( ~n25532 & n25582 ) | ( n25581 & n25582 ) ;
  assign n25584 = n25522 & ~n25583 ;
  assign n25585 = n25522 & ~n25584 ;
  assign n25586 = n25522 | n25583 ;
  assign n25587 = ~n25585 & n25586 ;
  assign n25588 = n4551 & ~n20569 ;
  assign n25589 = n4546 & ~n20580 ;
  assign n25590 = n4548 & ~n20584 ;
  assign n25591 = n25589 | n25590 ;
  assign n25592 = n25588 | n25591 ;
  assign n25593 = n4554 & n21884 ;
  assign n25594 = ( n4554 & ~n21889 ) | ( n4554 & n25593 ) | ( ~n21889 & n25593 ) ;
  assign n25595 = n25592 | n25594 ;
  assign n25596 = x23 | n25595 ;
  assign n25597 = ~x23 & n25596 ;
  assign n25598 = ( ~n25595 & n25596 ) | ( ~n25595 & n25597 ) | ( n25596 & n25597 ) ;
  assign n25599 = ~n25587 & n25598 ;
  assign n25600 = n25587 & ~n25598 ;
  assign n25601 = n25599 | n25600 ;
  assign n25602 = n25316 | n25320 ;
  assign n25603 = n25601 & ~n25602 ;
  assign n25604 = ~n25601 & n25602 ;
  assign n25605 = n25603 | n25604 ;
  assign n25606 = ( n25520 & n25521 ) | ( n25520 & ~n25605 ) | ( n25521 & ~n25605 ) ;
  assign n25607 = ( ~n25521 & n25605 ) | ( ~n25521 & n25606 ) | ( n25605 & n25606 ) ;
  assign n25608 = ( ~n25520 & n25606 ) | ( ~n25520 & n25607 ) | ( n25606 & n25607 ) ;
  assign n25609 = n25509 & ~n25608 ;
  assign n25610 = ~n25509 & n25608 ;
  assign n25611 = n25609 | n25610 ;
  assign n25612 = ~n25499 & n25611 ;
  assign n25613 = n25499 & ~n25611 ;
  assign n25614 = n25612 | n25613 ;
  assign n25615 = n25498 & ~n25614 ;
  assign n25616 = n25614 | n25615 ;
  assign n25617 = ( ~n25498 & n25615 ) | ( ~n25498 & n25616 ) | ( n25615 & n25616 ) ;
  assign n25618 = n25488 & ~n25617 ;
  assign n25619 = n25488 & ~n25618 ;
  assign n25620 = n25617 | n25618 ;
  assign n25621 = ~n25619 & n25620 ;
  assign n25622 = n25487 & ~n25621 ;
  assign n25623 = n25621 | n25622 ;
  assign n25624 = ( ~n25487 & n25622 ) | ( ~n25487 & n25623 ) | ( n25622 & n25623 ) ;
  assign n25625 = ~n25477 & n25624 ;
  assign n25626 = n25477 & ~n25624 ;
  assign n25627 = n25625 | n25626 ;
  assign n25628 = n25476 & ~n25627 ;
  assign n25629 = n25627 | n25628 ;
  assign n25630 = ( ~n25476 & n25628 ) | ( ~n25476 & n25629 ) | ( n25628 & n25629 ) ;
  assign n25631 = n25397 & n25630 ;
  assign n25632 = n25397 | n25630 ;
  assign n25633 = ~n25631 & n25632 ;
  assign n25634 = n9245 & n24324 ;
  assign n25635 = n8680 & n24329 ;
  assign n25636 = n8681 & ~n24334 ;
  assign n25637 = n25635 | n25636 ;
  assign n25638 = n25634 | n25637 ;
  assign n25639 = n8685 & ~n24353 ;
  assign n25640 = ( n8685 & n24356 ) | ( n8685 & n25639 ) | ( n24356 & n25639 ) ;
  assign n25641 = n25638 | n25640 ;
  assign n25642 = x5 | n25641 ;
  assign n25643 = ~x5 & n25642 ;
  assign n25644 = ( ~n25641 & n25642 ) | ( ~n25641 & n25643 ) | ( n25642 & n25643 ) ;
  assign n25645 = ~n25633 & n25644 ;
  assign n25646 = n25633 & ~n25644 ;
  assign n25647 = n25645 | n25646 ;
  assign n25648 = n25400 | n25405 ;
  assign n25649 = n25647 & ~n25648 ;
  assign n25650 = ~n25647 & n25648 ;
  assign n25651 = n25649 | n25650 ;
  assign n25652 = ~n25429 & n25432 ;
  assign n25653 = n3727 & ~n12318 ;
  assign n25654 = n3639 & n12608 ;
  assign n25655 = n25653 | n25654 ;
  assign n25656 = n3744 & ~n12314 ;
  assign n25657 = n25655 | n25656 ;
  assign n25658 = n3636 | n25657 ;
  assign n25659 = ( ~n14302 & n25657 ) | ( ~n14302 & n25658 ) | ( n25657 & n25658 ) ;
  assign n25660 = ( n616 & n25416 ) | ( n616 & n25426 ) | ( n25416 & n25426 ) ;
  assign n25661 = ( n25416 & n25418 ) | ( n25416 & ~n25425 ) | ( n25418 & ~n25425 ) ;
  assign n25662 = n616 | n25661 ;
  assign n25663 = ~n25660 & n25662 ;
  assign n25664 = n25659 & n25663 ;
  assign n25665 = n25663 & ~n25664 ;
  assign n25666 = ( n25659 & ~n25664 ) | ( n25659 & n25665 ) | ( ~n25664 & n25665 ) ;
  assign n25667 = n25652 & ~n25666 ;
  assign n25668 = ~n25652 & n25666 ;
  assign n25669 = n25667 | n25668 ;
  assign n25670 = n25435 | n25438 ;
  assign n25671 = ~n25669 & n25670 ;
  assign n25672 = n25436 & ~n25669 ;
  assign n25673 = ( n25185 & n25671 ) | ( n25185 & n25672 ) | ( n25671 & n25672 ) ;
  assign n25674 = ( n25185 & n25436 ) | ( n25185 & n25670 ) | ( n25436 & n25670 ) ;
  assign n25675 = n25669 & ~n25674 ;
  assign n25676 = n25673 | n25675 ;
  assign n25677 = n9798 & ~n25676 ;
  assign n25678 = n9782 & n25187 ;
  assign n25679 = n9783 & n25442 ;
  assign n25680 = n25678 | n25679 ;
  assign n25681 = n25677 | n25680 ;
  assign n25682 = ~n25442 & n25676 ;
  assign n25683 = n25187 | n25442 ;
  assign n25684 = ~n25682 & n25683 ;
  assign n25685 = n25442 & ~n25676 ;
  assign n25686 = n25187 & n25442 ;
  assign n25687 = ~n25685 & n25686 ;
  assign n25688 = n25685 | n25687 ;
  assign n25689 = ( n25449 & n25684 ) | ( n25449 & n25688 ) | ( n25684 & n25688 ) ;
  assign n25690 = n25682 | n25689 ;
  assign n25691 = ( n25449 & n25683 ) | ( n25449 & n25686 ) | ( n25683 & n25686 ) ;
  assign n25692 = n25684 & ~n25685 ;
  assign n25693 = ( n25449 & n25687 ) | ( n25449 & n25692 ) | ( n25687 & n25692 ) ;
  assign n25694 = n25691 & ~n25693 ;
  assign n25695 = n9787 & ~n25694 ;
  assign n25696 = n25690 & n25695 ;
  assign n25697 = ( n9787 & n25681 ) | ( n9787 & ~n25696 ) | ( n25681 & ~n25696 ) ;
  assign n25698 = x2 & n25697 ;
  assign n25699 = x2 & ~n25698 ;
  assign n25700 = ( n25697 & ~n25698 ) | ( n25697 & n25699 ) | ( ~n25698 & n25699 ) ;
  assign n25701 = ~n25651 & n25700 ;
  assign n25702 = n25651 & ~n25700 ;
  assign n25703 = n25701 | n25702 ;
  assign n25704 = n25457 | n25461 ;
  assign n25705 = ~n25703 & n25704 ;
  assign n25706 = n25703 & ~n25704 ;
  assign n25707 = n25705 | n25706 ;
  assign n25708 = n25464 & ~n25707 ;
  assign n25709 = ~n25464 & n25707 ;
  assign n25710 = n25708 | n25709 ;
  assign n25711 = n25701 | n25705 ;
  assign n25712 = n25645 | n25650 ;
  assign n25713 = n9245 & n25187 ;
  assign n25714 = n8680 & ~n24334 ;
  assign n25715 = n8681 & n24324 ;
  assign n25716 = n25714 | n25715 ;
  assign n25717 = n25713 | n25716 ;
  assign n25718 = n8685 | n25717 ;
  assign n25719 = ( n25193 & n25717 ) | ( n25193 & n25718 ) | ( n25717 & n25718 ) ;
  assign n25720 = x5 & n25719 ;
  assign n25721 = x5 & ~n25720 ;
  assign n25722 = ( n25719 & ~n25720 ) | ( n25719 & n25721 ) | ( ~n25720 & n25721 ) ;
  assign n25897 = ( n25397 & n25476 ) | ( n25397 & n25633 ) | ( n25476 & n25633 ) ;
  assign n25723 = n5503 & n24329 ;
  assign n25724 = n5512 & n20921 ;
  assign n25725 = n5508 & ~n21005 ;
  assign n25726 = n25724 | n25725 ;
  assign n25727 = n25723 | n25726 ;
  assign n25728 = n5515 & n24391 ;
  assign n25729 = ~n24392 & n25728 ;
  assign n25730 = ( n5515 & n25727 ) | ( n5515 & ~n25729 ) | ( n25727 & ~n25729 ) ;
  assign n25731 = x8 & n25730 ;
  assign n25732 = x8 & ~n25731 ;
  assign n25733 = ( n25730 & ~n25731 ) | ( n25730 & n25732 ) | ( ~n25731 & n25732 ) ;
  assign n25734 = n7305 & n20838 ;
  assign n25735 = n7300 & ~n20536 ;
  assign n25736 = n7302 & n20532 ;
  assign n25737 = n25735 | n25736 ;
  assign n25738 = n25734 | n25737 ;
  assign n25739 = n7308 | n25738 ;
  assign n25740 = ( ~n23712 & n25738 ) | ( ~n23712 & n25739 ) | ( n25738 & n25739 ) ;
  assign n25741 = ~x11 & n25740 ;
  assign n25742 = x11 | n25741 ;
  assign n25743 = ( ~n25740 & n25741 ) | ( ~n25740 & n25742 ) | ( n25741 & n25742 ) ;
  assign n25744 = n7280 & ~n20724 ;
  assign n25745 = n5384 & n20546 ;
  assign n25746 = n7277 & ~n20542 ;
  assign n25747 = n25745 | n25746 ;
  assign n25748 = n25744 | n25747 ;
  assign n25749 = n39 | n25748 ;
  assign n25750 = ( n23229 & n25748 ) | ( n23229 & n25749 ) | ( n25748 & n25749 ) ;
  assign n25751 = x14 & n25750 ;
  assign n25752 = x14 & ~n25751 ;
  assign n25753 = ( n25750 & ~n25751 ) | ( n25750 & n25752 ) | ( ~n25751 & n25752 ) ;
  assign n25754 = n25615 | n25618 ;
  assign n25755 = n4781 & n20562 ;
  assign n25756 = n4776 & ~n20689 ;
  assign n25757 = n4778 & n20560 ;
  assign n25758 = n25756 | n25757 ;
  assign n25759 = n25755 | n25758 ;
  assign n25760 = n4784 | n25759 ;
  assign n25761 = ( ~n21044 & n25759 ) | ( ~n21044 & n25760 ) | ( n25759 & n25760 ) ;
  assign n25762 = ~x20 & n25761 ;
  assign n25763 = x20 | n25762 ;
  assign n25764 = ( ~n25761 & n25762 ) | ( ~n25761 & n25763 ) | ( n25762 & n25763 ) ;
  assign n25765 = n25581 | n25584 ;
  assign n25766 = n4484 & ~n20580 ;
  assign n25767 = n4479 & ~n20591 ;
  assign n25768 = n4481 & n20588 ;
  assign n25769 = n25767 | n25768 ;
  assign n25770 = n25766 | n25769 ;
  assign n25771 = n4487 | n25770 ;
  assign n25772 = ( n21840 & n25770 ) | ( n21840 & n25771 ) | ( n25770 & n25771 ) ;
  assign n25773 = x26 & n25772 ;
  assign n25774 = x26 & ~n25773 ;
  assign n25775 = ( n25772 & ~n25773 ) | ( n25772 & n25774 ) | ( ~n25773 & n25774 ) ;
  assign n25776 = n25556 | n25560 ;
  assign n25777 = n3744 & n20611 ;
  assign n25778 = n3727 & n20614 ;
  assign n25779 = n3639 & n20616 ;
  assign n25780 = n25778 | n25779 ;
  assign n25781 = n25777 | n25780 ;
  assign n25782 = n3636 | n25781 ;
  assign n25783 = ( n21293 & n25781 ) | ( n21293 & n25782 ) | ( n25781 & n25782 ) ;
  assign n25784 = n1353 | n2036 ;
  assign n25785 = n709 | n1457 ;
  assign n25786 = n25784 | n25785 ;
  assign n25787 = n82 | n3476 ;
  assign n25788 = n1657 | n25787 ;
  assign n25789 = ( ~n11341 & n25786 ) | ( ~n11341 & n25788 ) | ( n25786 & n25788 ) ;
  assign n25790 = n11341 | n25789 ;
  assign n25791 = n1886 & ~n25790 ;
  assign n25792 = ~n3968 & n25791 ;
  assign n25793 = n948 | n2037 ;
  assign n25794 = n25045 | n25793 ;
  assign n25795 = n301 | n529 ;
  assign n25796 = n319 | n25795 ;
  assign n25797 = n416 | n25796 ;
  assign n25798 = n25794 | n25797 ;
  assign n25799 = n190 | n379 ;
  assign n25800 = n601 | n25799 ;
  assign n25801 = n145 | n25800 ;
  assign n25802 = n25798 | n25801 ;
  assign n25803 = n1079 | n25802 ;
  assign n25804 = n421 | n25803 ;
  assign n25805 = n862 | n25804 ;
  assign n25806 = n409 | n25805 ;
  assign n25807 = n25792 & ~n25806 ;
  assign n25808 = n595 | n781 ;
  assign n25809 = n649 | n25808 ;
  assign n25810 = n25807 & ~n25809 ;
  assign n25811 = n25783 & ~n25810 ;
  assign n25812 = n25783 & ~n25811 ;
  assign n25813 = n25783 | n25810 ;
  assign n25814 = ~n25812 & n25813 ;
  assign n25815 = n25776 & ~n25814 ;
  assign n25816 = n25776 & ~n25815 ;
  assign n25817 = n25814 | n25815 ;
  assign n25818 = ~n25816 & n25817 ;
  assign n25819 = n4048 & ~n20595 ;
  assign n25820 = n4043 & ~n20605 ;
  assign n25821 = n4045 & n20600 ;
  assign n25822 = n25820 | n25821 ;
  assign n25823 = n25819 | n25822 ;
  assign n25824 = n4051 | n25823 ;
  assign n25825 = ( ~n21554 & n25823 ) | ( ~n21554 & n25824 ) | ( n25823 & n25824 ) ;
  assign n25826 = ~x29 & n25825 ;
  assign n25827 = x29 | n25826 ;
  assign n25828 = ( ~n25825 & n25826 ) | ( ~n25825 & n25827 ) | ( n25826 & n25827 ) ;
  assign n25829 = ~n25818 & n25828 ;
  assign n25830 = n25818 & ~n25828 ;
  assign n25831 = n25829 | n25830 ;
  assign n25832 = n25574 | n25578 ;
  assign n25833 = ~n25831 & n25832 ;
  assign n25834 = n25831 & ~n25832 ;
  assign n25835 = n25833 | n25834 ;
  assign n25836 = n25775 & ~n25835 ;
  assign n25837 = n25835 | n25836 ;
  assign n25838 = ( ~n25775 & n25836 ) | ( ~n25775 & n25837 ) | ( n25836 & n25837 ) ;
  assign n25839 = n25765 & ~n25838 ;
  assign n25840 = n25765 & ~n25839 ;
  assign n25841 = n25765 | n25838 ;
  assign n25842 = ~n25840 & n25841 ;
  assign n25843 = n4551 & ~n20573 ;
  assign n25844 = n4546 & ~n20584 ;
  assign n25845 = n4548 & ~n20569 ;
  assign n25846 = n25844 | n25845 ;
  assign n25847 = n25843 | n25846 ;
  assign n25848 = n4554 | n25847 ;
  assign n25849 = ( ~n21860 & n25847 ) | ( ~n21860 & n25848 ) | ( n25847 & n25848 ) ;
  assign n25850 = ~x23 & n25849 ;
  assign n25851 = x23 | n25850 ;
  assign n25852 = ( ~n25849 & n25850 ) | ( ~n25849 & n25851 ) | ( n25850 & n25851 ) ;
  assign n25853 = ~n25842 & n25852 ;
  assign n25854 = n25842 & ~n25852 ;
  assign n25855 = n25853 | n25854 ;
  assign n25856 = n25599 | n25604 ;
  assign n25857 = n25855 & ~n25856 ;
  assign n25858 = ~n25855 & n25856 ;
  assign n25859 = n25857 | n25858 ;
  assign n25860 = n25764 & ~n25859 ;
  assign n25861 = n25859 | n25860 ;
  assign n25862 = ( ~n25764 & n25860 ) | ( ~n25764 & n25861 ) | ( n25860 & n25861 ) ;
  assign n25863 = n25606 & ~n25862 ;
  assign n25864 = n25606 & ~n25863 ;
  assign n25865 = n25606 | n25862 ;
  assign n25866 = ~n25864 & n25865 ;
  assign n25867 = n5083 & ~n20710 ;
  assign n25868 = n5069 & ~n20552 ;
  assign n25869 = n5070 & n20556 ;
  assign n25870 = n25868 | n25869 ;
  assign n25871 = n25867 | n25870 ;
  assign n25872 = n5074 | n25871 ;
  assign n25873 = ( ~n22641 & n25871 ) | ( ~n22641 & n25872 ) | ( n25871 & n25872 ) ;
  assign n25874 = ~x17 & n25873 ;
  assign n25875 = x17 | n25874 ;
  assign n25876 = ( ~n25873 & n25874 ) | ( ~n25873 & n25875 ) | ( n25874 & n25875 ) ;
  assign n25877 = ~n25866 & n25876 ;
  assign n25878 = n25866 & ~n25876 ;
  assign n25879 = n25877 | n25878 ;
  assign n25880 = n25609 | n25613 ;
  assign n25881 = n25879 & ~n25880 ;
  assign n25882 = ~n25879 & n25880 ;
  assign n25883 = n25881 | n25882 ;
  assign n25884 = ( n25753 & n25754 ) | ( n25753 & ~n25883 ) | ( n25754 & ~n25883 ) ;
  assign n25885 = ( ~n25754 & n25883 ) | ( ~n25754 & n25884 ) | ( n25883 & n25884 ) ;
  assign n25886 = ( ~n25753 & n25884 ) | ( ~n25753 & n25885 ) | ( n25884 & n25885 ) ;
  assign n25887 = n25743 & ~n25886 ;
  assign n25888 = ~n25743 & n25886 ;
  assign n25889 = n25887 | n25888 ;
  assign n25890 = n25622 | n25626 ;
  assign n25891 = n25889 & ~n25890 ;
  assign n25892 = ~n25889 & n25890 ;
  assign n25893 = n25891 | n25892 ;
  assign n25894 = n25733 & ~n25893 ;
  assign n25895 = n25893 | n25894 ;
  assign n25896 = ( ~n25733 & n25894 ) | ( ~n25733 & n25895 ) | ( n25894 & n25895 ) ;
  assign n25898 = ~n25896 & n25897 ;
  assign n25899 = n25897 & ~n25898 ;
  assign n25900 = n25896 | n25898 ;
  assign n25901 = ~n25899 & n25900 ;
  assign n25902 = n25722 & ~n25901 ;
  assign n25903 = n25901 | n25902 ;
  assign n25904 = ( ~n25722 & n25902 ) | ( ~n25722 & n25903 ) | ( n25902 & n25903 ) ;
  assign n25905 = ~n25712 & n25904 ;
  assign n25906 = n25712 & ~n25904 ;
  assign n25907 = n25905 | n25906 ;
  assign n25908 = n3727 | n3744 ;
  assign n25909 = ~n12314 & n25908 ;
  assign n25910 = n3639 | n25909 ;
  assign n25911 = ( ~n12318 & n25909 ) | ( ~n12318 & n25910 ) | ( n25909 & n25910 ) ;
  assign n25912 = n3636 & ~n17966 ;
  assign n25913 = n25911 | n25912 ;
  assign n25914 = n616 & ~n25913 ;
  assign n25915 = ~n616 & n25913 ;
  assign n25916 = n25914 | n25915 ;
  assign n25917 = n25660 | n25664 ;
  assign n25918 = n25916 | n25917 ;
  assign n25919 = n25916 & n25917 ;
  assign n25920 = n25918 & ~n25919 ;
  assign n25921 = n25668 | n25671 ;
  assign n25922 = n25920 & n25921 ;
  assign n25923 = n25668 | n25672 ;
  assign n25924 = n25920 & n25923 ;
  assign n25925 = ( n25185 & n25922 ) | ( n25185 & n25924 ) | ( n25922 & n25924 ) ;
  assign n25926 = ( n25185 & n25921 ) | ( n25185 & n25923 ) | ( n25921 & n25923 ) ;
  assign n25927 = n25920 | n25926 ;
  assign n25928 = ~n25925 & n25927 ;
  assign n25929 = n25676 & ~n25928 ;
  assign n25930 = ~n25676 & n25928 ;
  assign n25931 = n25929 | n25930 ;
  assign n25932 = n25684 & ~n25931 ;
  assign n25933 = n25688 & ~n25931 ;
  assign n25934 = ( n25449 & n25932 ) | ( n25449 & n25933 ) | ( n25932 & n25933 ) ;
  assign n25935 = ~n25689 & n25931 ;
  assign n25936 = n25934 | n25935 ;
  assign n25937 = n9798 & n25928 ;
  assign n25938 = n9782 & n25442 ;
  assign n25939 = n9783 & ~n25676 ;
  assign n25940 = n25938 | n25939 ;
  assign n25941 = n25937 | n25940 ;
  assign n25942 = n9787 | n25941 ;
  assign n25943 = ( ~n25936 & n25941 ) | ( ~n25936 & n25942 ) | ( n25941 & n25942 ) ;
  assign n25944 = ~x2 & n25943 ;
  assign n25945 = x2 | n25944 ;
  assign n25946 = ( ~n25943 & n25944 ) | ( ~n25943 & n25945 ) | ( n25944 & n25945 ) ;
  assign n25947 = ~n25907 & n25946 ;
  assign n25948 = n25907 & ~n25946 ;
  assign n25949 = n25947 | n25948 ;
  assign n25950 = n25711 & ~n25949 ;
  assign n25951 = ~n25711 & n25949 ;
  assign n25952 = n25950 | n25951 ;
  assign n25953 = n25708 & ~n25952 ;
  assign n25954 = ~n25708 & n25952 ;
  assign n25955 = n25953 | n25954 ;
  assign n25956 = n25947 | n25950 ;
  assign n25957 = n25902 | n25906 ;
  assign n25958 = n9245 & n25442 ;
  assign n25959 = n8680 & n24324 ;
  assign n25960 = n8681 & n25187 ;
  assign n25961 = n25959 | n25960 ;
  assign n25962 = n25958 | n25961 ;
  assign n25963 = n8685 | n25962 ;
  assign n25964 = ( n25452 & n25962 ) | ( n25452 & n25963 ) | ( n25962 & n25963 ) ;
  assign n25965 = x5 & n25964 ;
  assign n25966 = x5 & ~n25965 ;
  assign n25967 = ( n25964 & ~n25965 ) | ( n25964 & n25966 ) | ( ~n25965 & n25966 ) ;
  assign n25968 = n25894 | n25898 ;
  assign n25969 = n5503 & ~n24334 ;
  assign n25970 = n5512 & ~n21005 ;
  assign n25971 = n5508 & n24329 ;
  assign n25972 = n25970 | n25971 ;
  assign n25973 = n25969 | n25972 ;
  assign n25974 = n5515 & ~n24376 ;
  assign n25975 = n24373 & n25974 ;
  assign n25976 = ( n5515 & n25973 ) | ( n5515 & ~n25975 ) | ( n25973 & ~n25975 ) ;
  assign n25977 = x8 & n25976 ;
  assign n25978 = x8 & ~n25977 ;
  assign n25979 = ( n25976 & ~n25977 ) | ( n25976 & n25978 ) | ( ~n25977 & n25978 ) ;
  assign n25980 = n25887 | n25892 ;
  assign n25981 = n7280 & ~n20536 ;
  assign n25982 = n5384 & ~n20542 ;
  assign n25983 = n7277 & ~n20724 ;
  assign n25984 = n25982 | n25983 ;
  assign n25985 = n25981 | n25984 ;
  assign n25986 = n39 & ~n23213 ;
  assign n25987 = n23217 & n25986 ;
  assign n25988 = ( n39 & n25985 ) | ( n39 & ~n25987 ) | ( n25985 & ~n25987 ) ;
  assign n25989 = x14 & n25988 ;
  assign n25990 = x14 & ~n25989 ;
  assign n25991 = ( n25988 & ~n25989 ) | ( n25988 & n25990 ) | ( ~n25989 & n25990 ) ;
  assign n25992 = n25860 | n25863 ;
  assign n25993 = n4781 & ~n20552 ;
  assign n25994 = n4776 & n20560 ;
  assign n25995 = n4778 & n20562 ;
  assign n25996 = n25994 | n25995 ;
  assign n25997 = n25993 | n25996 ;
  assign n25998 = n4784 & n22510 ;
  assign n25999 = ~n22512 & n25998 ;
  assign n26000 = ( n4784 & n25997 ) | ( n4784 & ~n25999 ) | ( n25997 & ~n25999 ) ;
  assign n26001 = x20 & n26000 ;
  assign n26002 = x20 & ~n26001 ;
  assign n26003 = ( n26000 & ~n26001 ) | ( n26000 & n26002 ) | ( ~n26001 & n26002 ) ;
  assign n26004 = n25853 | n25858 ;
  assign n26005 = n4551 & ~n20689 ;
  assign n26006 = n4546 & ~n20569 ;
  assign n26007 = n4548 & ~n20573 ;
  assign n26008 = n26006 | n26007 ;
  assign n26009 = n26005 | n26008 ;
  assign n26010 = ( n4554 & ~n22192 ) | ( n4554 & n22193 ) | ( ~n22192 & n22193 ) ;
  assign n26011 = n26009 | n26010 ;
  assign n26012 = x23 | n26011 ;
  assign n26013 = ~x23 & n26012 ;
  assign n26014 = ( ~n26011 & n26012 ) | ( ~n26011 & n26013 ) | ( n26012 & n26013 ) ;
  assign n26015 = n25836 | n25839 ;
  assign n26016 = n4484 & ~n20584 ;
  assign n26017 = n4479 & n20588 ;
  assign n26018 = n4481 & ~n20580 ;
  assign n26019 = n26017 | n26018 ;
  assign n26020 = n26016 | n26019 ;
  assign n26021 = n4487 | n26020 ;
  assign n26022 = ( ~n21901 & n26020 ) | ( ~n21901 & n26021 ) | ( n26020 & n26021 ) ;
  assign n26023 = ~x26 & n26022 ;
  assign n26024 = x26 | n26023 ;
  assign n26025 = ( ~n26022 & n26023 ) | ( ~n26022 & n26024 ) | ( n26023 & n26024 ) ;
  assign n26026 = n25829 | n25833 ;
  assign n26027 = n25811 | n25815 ;
  assign n26028 = n3744 & ~n20605 ;
  assign n26029 = n3727 & n20611 ;
  assign n26030 = n3639 & n20614 ;
  assign n26031 = n26029 | n26030 ;
  assign n26032 = n26028 | n26031 ;
  assign n26033 = n3636 | n26032 ;
  assign n26034 = ( ~n21275 & n26032 ) | ( ~n21275 & n26033 ) | ( n26032 & n26033 ) ;
  assign n26035 = n688 | n1200 ;
  assign n26036 = n736 | n26035 ;
  assign n26037 = n11181 | n26036 ;
  assign n26038 = ( n11139 & n14078 ) | ( n11139 & n26037 ) | ( n14078 & n26037 ) ;
  assign n26039 = n14078 & ~n26038 ;
  assign n26040 = ~n4417 & n26039 ;
  assign n26041 = n478 | n571 ;
  assign n26042 = n529 | n26041 ;
  assign n26043 = n428 | n26042 ;
  assign n26044 = n470 | n26043 ;
  assign n26045 = n55 | n26044 ;
  assign n26046 = n458 | n26045 ;
  assign n26047 = n441 | n26046 ;
  assign n26048 = n96 | n26047 ;
  assign n26049 = n26040 & ~n26048 ;
  assign n26050 = n122 | n126 ;
  assign n26051 = n646 | n26050 ;
  assign n26052 = n26049 & ~n26051 ;
  assign n26053 = n26034 & ~n26052 ;
  assign n26054 = n26034 & ~n26053 ;
  assign n26055 = n26034 | n26052 ;
  assign n26056 = ~n26054 & n26055 ;
  assign n26057 = n26027 & ~n26056 ;
  assign n26058 = ~n26027 & n26056 ;
  assign n26059 = n26057 | n26058 ;
  assign n26060 = n4048 & ~n20591 ;
  assign n26061 = n4043 & n20600 ;
  assign n26062 = n4045 & ~n20595 ;
  assign n26063 = n26061 | n26062 ;
  assign n26064 = n26060 | n26063 ;
  assign n26065 = n4051 & ~n21539 ;
  assign n26066 = ~n21543 & n26065 ;
  assign n26067 = ( n4051 & n26064 ) | ( n4051 & ~n26066 ) | ( n26064 & ~n26066 ) ;
  assign n26068 = ~x29 & n26067 ;
  assign n26069 = x29 | n26068 ;
  assign n26070 = ( ~n26067 & n26068 ) | ( ~n26067 & n26069 ) | ( n26068 & n26069 ) ;
  assign n26071 = ~n26059 & n26070 ;
  assign n26072 = n26059 & ~n26070 ;
  assign n26073 = n26071 | n26072 ;
  assign n26074 = n26026 & ~n26073 ;
  assign n26075 = ~n26026 & n26073 ;
  assign n26076 = n26074 | n26075 ;
  assign n26077 = n26025 & ~n26076 ;
  assign n26078 = n26076 | n26077 ;
  assign n26079 = ( ~n26025 & n26077 ) | ( ~n26025 & n26078 ) | ( n26077 & n26078 ) ;
  assign n26080 = n26015 & ~n26079 ;
  assign n26081 = n26015 & ~n26080 ;
  assign n26082 = n26079 | n26080 ;
  assign n26083 = ~n26081 & n26082 ;
  assign n26084 = n26014 & ~n26083 ;
  assign n26085 = n26083 | n26084 ;
  assign n26086 = ( ~n26014 & n26084 ) | ( ~n26014 & n26085 ) | ( n26084 & n26085 ) ;
  assign n26087 = ~n26004 & n26086 ;
  assign n26088 = n26004 & ~n26086 ;
  assign n26089 = n26087 | n26088 ;
  assign n26090 = n26003 & ~n26089 ;
  assign n26091 = n26089 | n26090 ;
  assign n26092 = ( ~n26003 & n26090 ) | ( ~n26003 & n26091 ) | ( n26090 & n26091 ) ;
  assign n26093 = n25992 & ~n26092 ;
  assign n26094 = n25992 & ~n26093 ;
  assign n26095 = n25992 | n26092 ;
  assign n26096 = ~n26094 & n26095 ;
  assign n26097 = n5083 & n20546 ;
  assign n26098 = n5069 & n20556 ;
  assign n26099 = n5070 & ~n20710 ;
  assign n26100 = n26098 | n26099 ;
  assign n26101 = n26097 | n26100 ;
  assign n26102 = n5074 & ~n21031 ;
  assign n26103 = ( n5074 & n21037 ) | ( n5074 & n26102 ) | ( n21037 & n26102 ) ;
  assign n26104 = n26101 | n26103 ;
  assign n26105 = x17 | n26104 ;
  assign n26106 = ~x17 & n26105 ;
  assign n26107 = ( ~n26104 & n26105 ) | ( ~n26104 & n26106 ) | ( n26105 & n26106 ) ;
  assign n26108 = ~n26096 & n26107 ;
  assign n26109 = n26096 & ~n26107 ;
  assign n26110 = n26108 | n26109 ;
  assign n26111 = n25877 | n25882 ;
  assign n26112 = n26110 & ~n26111 ;
  assign n26113 = ~n26110 & n26111 ;
  assign n26114 = n26112 | n26113 ;
  assign n26115 = n25991 & ~n26114 ;
  assign n26116 = n26114 | n26115 ;
  assign n26117 = ( ~n25991 & n26115 ) | ( ~n25991 & n26116 ) | ( n26115 & n26116 ) ;
  assign n26118 = n25884 & ~n26117 ;
  assign n26119 = n25884 & ~n26118 ;
  assign n26120 = n25884 | n26117 ;
  assign n26121 = ~n26119 & n26120 ;
  assign n26122 = n7305 & n20921 ;
  assign n26123 = n7300 & n20532 ;
  assign n26124 = n7302 & n20838 ;
  assign n26125 = n26123 | n26124 ;
  assign n26126 = n26122 | n26125 ;
  assign n26127 = ( n7308 & n23691 ) | ( n7308 & n23695 ) | ( n23691 & n23695 ) ;
  assign n26128 = n26126 | n26127 ;
  assign n26129 = x11 | n26128 ;
  assign n26130 = ~x11 & n26129 ;
  assign n26131 = ( ~n26128 & n26129 ) | ( ~n26128 & n26130 ) | ( n26129 & n26130 ) ;
  assign n26132 = ~n26121 & n26131 ;
  assign n26133 = n26121 & ~n26131 ;
  assign n26134 = n26132 | n26133 ;
  assign n26135 = ~n25980 & n26134 ;
  assign n26136 = n25980 & ~n26134 ;
  assign n26137 = n26135 | n26136 ;
  assign n26138 = n25979 & ~n26137 ;
  assign n26139 = n26137 | n26138 ;
  assign n26140 = ( ~n25979 & n26138 ) | ( ~n25979 & n26139 ) | ( n26138 & n26139 ) ;
  assign n26141 = n25968 & ~n26140 ;
  assign n26142 = n25968 & ~n26141 ;
  assign n26143 = n26140 | n26141 ;
  assign n26144 = ~n26142 & n26143 ;
  assign n26145 = n25967 & ~n26144 ;
  assign n26146 = n26144 | n26145 ;
  assign n26147 = ( ~n25967 & n26145 ) | ( ~n25967 & n26146 ) | ( n26145 & n26146 ) ;
  assign n26148 = ~n25957 & n26147 ;
  assign n26149 = n25957 & ~n26147 ;
  assign n26150 = n26148 | n26149 ;
  assign n26151 = x31 | n44 ;
  assign n26152 = ~n12314 & n26151 ;
  assign n26153 = n25919 | n25925 ;
  assign n26154 = ( n25914 & n26152 ) | ( n25914 & ~n26153 ) | ( n26152 & ~n26153 ) ;
  assign n26155 = ( ~n25914 & n26153 ) | ( ~n25914 & n26154 ) | ( n26153 & n26154 ) ;
  assign n26156 = ( ~n26152 & n26154 ) | ( ~n26152 & n26155 ) | ( n26154 & n26155 ) ;
  assign n26157 = n25928 & n26156 ;
  assign n26158 = n25928 | n26156 ;
  assign n26159 = ( n25930 & n25932 ) | ( n25930 & n26158 ) | ( n25932 & n26158 ) ;
  assign n26160 = ~n26157 & n26159 ;
  assign n26161 = ( n25930 & n25933 ) | ( n25930 & n26160 ) | ( n25933 & n26160 ) ;
  assign n26162 = ( n25449 & n26160 ) | ( n25449 & n26161 ) | ( n26160 & n26161 ) ;
  assign n26163 = n25930 | n25934 ;
  assign n26164 = ~n26162 & n26163 ;
  assign n26165 = n26157 | n26162 ;
  assign n26166 = n26158 & ~n26165 ;
  assign n26167 = n26164 | n26166 ;
  assign n26168 = n9798 & n26156 ;
  assign n26169 = n9782 & ~n25676 ;
  assign n26170 = n9783 & n25928 ;
  assign n26171 = n26169 | n26170 ;
  assign n26172 = n26168 | n26171 ;
  assign n26173 = n9787 | n26172 ;
  assign n26174 = ( n26167 & n26172 ) | ( n26167 & n26173 ) | ( n26172 & n26173 ) ;
  assign n26175 = x2 & n26174 ;
  assign n26176 = x2 & ~n26175 ;
  assign n26177 = ( n26174 & ~n26175 ) | ( n26174 & n26176 ) | ( ~n26175 & n26176 ) ;
  assign n26178 = ~n26150 & n26177 ;
  assign n26179 = n26150 & ~n26177 ;
  assign n26180 = n26178 | n26179 ;
  assign n26181 = n25956 & ~n26180 ;
  assign n26182 = ~n25956 & n26180 ;
  assign n26183 = n26181 | n26182 ;
  assign n26184 = n25953 & ~n26183 ;
  assign n26185 = ~n25953 & n26183 ;
  assign n26186 = n26184 | n26185 ;
  assign n26187 = n17962 & n26156 ;
  assign n26188 = n9782 & n25928 ;
  assign n26189 = n26187 | n26188 ;
  assign n26190 = n9787 | n26189 ;
  assign n26191 = ( n26165 & n26189 ) | ( n26165 & n26190 ) | ( n26189 & n26190 ) ;
  assign n26192 = x2 & n26191 ;
  assign n26193 = x2 & ~n26192 ;
  assign n26194 = ( n26191 & ~n26192 ) | ( n26191 & n26193 ) | ( ~n26192 & n26193 ) ;
  assign n26195 = n9245 & ~n25676 ;
  assign n26196 = n8680 & n25187 ;
  assign n26197 = n8681 & n25442 ;
  assign n26198 = n26196 | n26197 ;
  assign n26199 = n26195 | n26198 ;
  assign n26200 = n8685 & ~n25690 ;
  assign n26201 = ( n8685 & n25694 ) | ( n8685 & n26200 ) | ( n25694 & n26200 ) ;
  assign n26202 = n26199 | n26201 ;
  assign n26203 = x5 | n26202 ;
  assign n26204 = ~x5 & n26203 ;
  assign n26205 = ( ~n26202 & n26203 ) | ( ~n26202 & n26204 ) | ( n26203 & n26204 ) ;
  assign n26206 = n26132 | n26136 ;
  assign n26207 = n7305 & ~n21005 ;
  assign n26208 = n7300 & n20838 ;
  assign n26209 = n7302 & n20921 ;
  assign n26210 = n26208 | n26209 ;
  assign n26211 = n26207 | n26210 ;
  assign n26212 = n7308 | n26211 ;
  assign n26213 = ( ~n21015 & n26211 ) | ( ~n21015 & n26212 ) | ( n26211 & n26212 ) ;
  assign n26214 = ~x11 & n26213 ;
  assign n26215 = x11 | n26214 ;
  assign n26216 = ( ~n26213 & n26214 ) | ( ~n26213 & n26215 ) | ( n26214 & n26215 ) ;
  assign n26217 = n26108 | n26113 ;
  assign n26218 = n5083 & ~n20542 ;
  assign n26219 = n5069 & ~n20710 ;
  assign n26220 = n5070 & n20546 ;
  assign n26221 = n26219 | n26220 ;
  assign n26222 = n26218 | n26221 ;
  assign n26223 = n5074 | n26222 ;
  assign n26224 = ( ~n23042 & n26222 ) | ( ~n23042 & n26223 ) | ( n26222 & n26223 ) ;
  assign n26225 = ~x17 & n26224 ;
  assign n26226 = x17 | n26225 ;
  assign n26227 = ( ~n26224 & n26225 ) | ( ~n26224 & n26226 ) | ( n26225 & n26226 ) ;
  assign n26228 = n4551 & n20560 ;
  assign n26229 = n4546 & ~n20573 ;
  assign n26230 = n4548 & ~n20689 ;
  assign n26231 = n26229 | n26230 ;
  assign n26232 = n26228 | n26231 ;
  assign n26233 = ( n4554 & n22173 ) | ( n4554 & n22176 ) | ( n22173 & n22176 ) ;
  assign n26234 = n26232 | n26233 ;
  assign n26235 = x23 | n26234 ;
  assign n26236 = ~x23 & n26235 ;
  assign n26237 = ( ~n26234 & n26235 ) | ( ~n26234 & n26236 ) | ( n26235 & n26236 ) ;
  assign n26238 = n26053 | n26057 ;
  assign n26239 = n3744 & n20600 ;
  assign n26240 = n3727 & ~n20605 ;
  assign n26241 = n3639 & n20611 ;
  assign n26242 = n26240 | n26241 ;
  assign n26243 = n26239 | n26242 ;
  assign n26244 = n3636 | n26243 ;
  assign n26245 = ( ~n21432 & n26243 ) | ( ~n21432 & n26244 ) | ( n26243 & n26244 ) ;
  assign n26246 = n58 | n143 ;
  assign n26247 = n122 | n26246 ;
  assign n26248 = n1632 | n2169 ;
  assign n26249 = ( n242 & ~n2502 ) | ( n242 & n26248 ) | ( ~n2502 & n26248 ) ;
  assign n26250 = n2502 | n26249 ;
  assign n26251 = n26247 | n26250 ;
  assign n26252 = n843 | n3476 ;
  assign n26253 = n1921 | n25543 ;
  assign n26254 = n26252 | n26253 ;
  assign n26255 = n26251 | n26254 ;
  assign n26256 = n12688 | n26255 ;
  assign n26257 = n4088 | n26256 ;
  assign n26258 = n1261 | n13012 ;
  assign n26259 = n26257 | n26258 ;
  assign n26260 = n2361 | n3054 ;
  assign n26261 = n26259 | n26260 ;
  assign n26262 = n279 | n718 ;
  assign n26263 = n570 | n26262 ;
  assign n26264 = n226 & ~n26263 ;
  assign n26265 = ~n175 & n26264 ;
  assign n26266 = ~n110 & n26265 ;
  assign n26267 = ~n132 & n26266 ;
  assign n26268 = ~n145 & n26267 ;
  assign n26269 = ~n206 & n26268 ;
  assign n26270 = ~n26261 & n26269 ;
  assign n26271 = n26245 & ~n26270 ;
  assign n26272 = n26245 & ~n26271 ;
  assign n26273 = n26245 | n26270 ;
  assign n26274 = ~n26272 & n26273 ;
  assign n26275 = n26238 & ~n26274 ;
  assign n26276 = ~n26238 & n26274 ;
  assign n26277 = n26275 | n26276 ;
  assign n26278 = n4048 & n20588 ;
  assign n26279 = n4043 & ~n20595 ;
  assign n26280 = n4045 & ~n20591 ;
  assign n26281 = n26279 | n26280 ;
  assign n26282 = n26278 | n26281 ;
  assign n26283 = n4051 | n26282 ;
  assign n26284 = ( n21526 & n26282 ) | ( n21526 & n26283 ) | ( n26282 & n26283 ) ;
  assign n26285 = x29 & n26284 ;
  assign n26286 = x29 & ~n26285 ;
  assign n26287 = ( n26284 & ~n26285 ) | ( n26284 & n26286 ) | ( ~n26285 & n26286 ) ;
  assign n26288 = ~n26277 & n26287 ;
  assign n26289 = n26277 & ~n26287 ;
  assign n26290 = n26288 | n26289 ;
  assign n26291 = n26071 | n26074 ;
  assign n26292 = ~n26290 & n26291 ;
  assign n26293 = n26290 & ~n26291 ;
  assign n26294 = n26292 | n26293 ;
  assign n26295 = n4484 & ~n20569 ;
  assign n26296 = n4479 & ~n20580 ;
  assign n26297 = n4481 & ~n20584 ;
  assign n26298 = n26296 | n26297 ;
  assign n26299 = n26295 | n26298 ;
  assign n26300 = n4487 & ~n21884 ;
  assign n26301 = n21889 & n26300 ;
  assign n26302 = ( n4487 & n26299 ) | ( n4487 & ~n26301 ) | ( n26299 & ~n26301 ) ;
  assign n26303 = x26 & n26302 ;
  assign n26304 = x26 & ~n26303 ;
  assign n26305 = ( n26302 & ~n26303 ) | ( n26302 & n26304 ) | ( ~n26303 & n26304 ) ;
  assign n26306 = ~n26294 & n26305 ;
  assign n26307 = n26294 & ~n26305 ;
  assign n26308 = n26306 | n26307 ;
  assign n26309 = ~n26077 & n26308 ;
  assign n26310 = ~n26080 & n26309 ;
  assign n26311 = ( n26077 & n26080 ) | ( n26077 & ~n26308 ) | ( n26080 & ~n26308 ) ;
  assign n26312 = n26310 | n26311 ;
  assign n26313 = n26237 & ~n26312 ;
  assign n26314 = n26312 | n26313 ;
  assign n26315 = ( ~n26237 & n26313 ) | ( ~n26237 & n26314 ) | ( n26313 & n26314 ) ;
  assign n26316 = ~n26084 & n26315 ;
  assign n26317 = ~n26088 & n26316 ;
  assign n26318 = ( n26084 & n26088 ) | ( n26084 & ~n26315 ) | ( n26088 & ~n26315 ) ;
  assign n26319 = n26317 | n26318 ;
  assign n26320 = n4781 & n20556 ;
  assign n26321 = n4776 & n20562 ;
  assign n26322 = n4778 & ~n20552 ;
  assign n26323 = n26321 | n26322 ;
  assign n26324 = n26320 | n26323 ;
  assign n26325 = n4784 | n26324 ;
  assign n26326 = ( ~n22655 & n26324 ) | ( ~n22655 & n26325 ) | ( n26324 & n26325 ) ;
  assign n26327 = ~x20 & n26326 ;
  assign n26328 = x20 | n26327 ;
  assign n26329 = ( ~n26326 & n26327 ) | ( ~n26326 & n26328 ) | ( n26327 & n26328 ) ;
  assign n26330 = ~n26319 & n26329 ;
  assign n26331 = n26319 & ~n26329 ;
  assign n26332 = n26330 | n26331 ;
  assign n26333 = n26090 | n26093 ;
  assign n26334 = ~n26332 & n26333 ;
  assign n26335 = n26332 & ~n26333 ;
  assign n26336 = n26334 | n26335 ;
  assign n26337 = n26227 & ~n26336 ;
  assign n26338 = n26336 | n26337 ;
  assign n26339 = ( ~n26227 & n26337 ) | ( ~n26227 & n26338 ) | ( n26337 & n26338 ) ;
  assign n26340 = ~n26217 & n26339 ;
  assign n26341 = n26217 & ~n26339 ;
  assign n26342 = n26340 | n26341 ;
  assign n26343 = n7280 & n20532 ;
  assign n26344 = n5384 & ~n20724 ;
  assign n26345 = n7277 & ~n20536 ;
  assign n26346 = n26344 | n26345 ;
  assign n26347 = n26343 | n26346 ;
  assign n26348 = n39 | n26347 ;
  assign n26349 = ( n23203 & n26347 ) | ( n23203 & n26348 ) | ( n26347 & n26348 ) ;
  assign n26350 = x14 & n26349 ;
  assign n26351 = x14 & ~n26350 ;
  assign n26352 = ( n26349 & ~n26350 ) | ( n26349 & n26351 ) | ( ~n26350 & n26351 ) ;
  assign n26353 = ~n26342 & n26352 ;
  assign n26354 = n26342 & ~n26352 ;
  assign n26355 = n26353 | n26354 ;
  assign n26356 = n26115 | n26118 ;
  assign n26357 = ~n26355 & n26356 ;
  assign n26358 = n26355 & ~n26356 ;
  assign n26359 = n26357 | n26358 ;
  assign n26360 = n26216 & ~n26359 ;
  assign n26361 = n26359 | n26360 ;
  assign n26362 = ( ~n26216 & n26360 ) | ( ~n26216 & n26361 ) | ( n26360 & n26361 ) ;
  assign n26363 = ~n26206 & n26362 ;
  assign n26364 = n26206 & ~n26362 ;
  assign n26365 = n26363 | n26364 ;
  assign n26366 = n5503 & n24324 ;
  assign n26367 = n5512 & n24329 ;
  assign n26368 = n5508 & ~n24334 ;
  assign n26369 = n26367 | n26368 ;
  assign n26370 = n26366 | n26369 ;
  assign n26371 = n5515 & ~n24356 ;
  assign n26372 = n24353 & n26371 ;
  assign n26373 = ( n5515 & n26370 ) | ( n5515 & ~n26372 ) | ( n26370 & ~n26372 ) ;
  assign n26374 = x8 & n26373 ;
  assign n26375 = x8 & ~n26374 ;
  assign n26376 = ( n26373 & ~n26374 ) | ( n26373 & n26375 ) | ( ~n26374 & n26375 ) ;
  assign n26377 = ~n26365 & n26376 ;
  assign n26378 = n26365 & ~n26376 ;
  assign n26379 = n26377 | n26378 ;
  assign n26380 = ~n26138 & n26379 ;
  assign n26381 = ~n26141 & n26380 ;
  assign n26382 = ( n26138 & n26141 ) | ( n26138 & ~n26379 ) | ( n26141 & ~n26379 ) ;
  assign n26383 = n26381 | n26382 ;
  assign n26384 = n26205 & ~n26383 ;
  assign n26385 = n26383 | n26384 ;
  assign n26386 = ( ~n26205 & n26384 ) | ( ~n26205 & n26385 ) | ( n26384 & n26385 ) ;
  assign n26387 = n26194 & ~n26386 ;
  assign n26388 = ~n26194 & n26386 ;
  assign n26389 = n26387 | n26388 ;
  assign n26390 = n26145 | n26149 ;
  assign n26391 = n26389 & ~n26390 ;
  assign n26392 = ~n26389 & n26390 ;
  assign n26393 = n26391 | n26392 ;
  assign n26394 = ~n26178 & n26393 ;
  assign n26395 = ~n26181 & n26394 ;
  assign n26396 = ( n26178 & n26181 ) | ( n26178 & ~n26393 ) | ( n26181 & ~n26393 ) ;
  assign n26397 = n26395 | n26396 ;
  assign n26398 = n26184 & ~n26397 ;
  assign n26399 = ~n26184 & n26397 ;
  assign n26400 = n26398 | n26399 ;
  assign n26401 = n26306 | n26311 ;
  assign n26402 = n4484 & ~n20573 ;
  assign n26403 = n4479 & ~n20584 ;
  assign n26404 = n4481 & ~n20569 ;
  assign n26405 = n26403 | n26404 ;
  assign n26406 = n26402 | n26405 ;
  assign n26407 = n4487 | n26406 ;
  assign n26408 = ( ~n21860 & n26406 ) | ( ~n21860 & n26407 ) | ( n26406 & n26407 ) ;
  assign n26409 = ~x26 & n26408 ;
  assign n26410 = x26 | n26409 ;
  assign n26411 = ( ~n26408 & n26409 ) | ( ~n26408 & n26410 ) | ( n26409 & n26410 ) ;
  assign n26412 = n3744 & ~n20595 ;
  assign n26413 = n3639 & ~n20605 ;
  assign n26414 = n3727 & n20600 ;
  assign n26415 = n26413 | n26414 ;
  assign n26416 = n26412 | n26415 ;
  assign n26417 = n3636 | n26416 ;
  assign n26418 = ( ~n21554 & n26416 ) | ( ~n21554 & n26417 ) | ( n26416 & n26417 ) ;
  assign n26419 = n2015 | n2305 ;
  assign n26420 = n5690 | n19746 ;
  assign n26421 = n26419 | n26420 ;
  assign n26422 = n820 | n26421 ;
  assign n26423 = ~n555 & n19817 ;
  assign n26424 = ~n26422 & n26423 ;
  assign n26425 = ~n1784 & n26424 ;
  assign n26426 = ~n759 & n26425 ;
  assign n26427 = ~n3462 & n26426 ;
  assign n26428 = n362 | n2445 ;
  assign n26429 = n278 | n26428 ;
  assign n26430 = n26427 & ~n26429 ;
  assign n26431 = n55 | n13253 ;
  assign n26432 = n213 | n26431 ;
  assign n26433 = n457 | n26432 ;
  assign n26434 = n102 | n26433 ;
  assign n26435 = n26430 & ~n26434 ;
  assign n26436 = ( x2 & ~n12977 ) | ( x2 & n26156 ) | ( ~n12977 & n26156 ) ;
  assign n26437 = x2 & ~n26436 ;
  assign n26438 = ( n26156 & ~n26436 ) | ( n26156 & n26437 ) | ( ~n26436 & n26437 ) ;
  assign n26439 = ~n26435 & n26438 ;
  assign n26440 = n26435 & ~n26438 ;
  assign n26441 = n26439 | n26440 ;
  assign n26442 = n26418 & ~n26441 ;
  assign n26443 = n26418 & ~n26442 ;
  assign n26444 = n26441 | n26442 ;
  assign n26445 = ~n26443 & n26444 ;
  assign n26446 = n26271 | n26275 ;
  assign n26447 = n26445 & ~n26446 ;
  assign n26448 = ~n26445 & n26446 ;
  assign n26449 = n26447 | n26448 ;
  assign n26450 = n4048 & ~n20580 ;
  assign n26451 = n4043 & ~n20591 ;
  assign n26452 = n4045 & n20588 ;
  assign n26453 = n26451 | n26452 ;
  assign n26454 = n26450 | n26453 ;
  assign n26455 = n4051 | n26454 ;
  assign n26456 = ( n21840 & n26454 ) | ( n21840 & n26455 ) | ( n26454 & n26455 ) ;
  assign n26457 = x29 & n26456 ;
  assign n26458 = x29 & ~n26457 ;
  assign n26459 = ( n26456 & ~n26457 ) | ( n26456 & n26458 ) | ( ~n26457 & n26458 ) ;
  assign n26460 = ~n26449 & n26459 ;
  assign n26461 = n26449 & ~n26459 ;
  assign n26462 = n26460 | n26461 ;
  assign n26463 = n26288 | n26292 ;
  assign n26464 = ( n26411 & n26462 ) | ( n26411 & ~n26463 ) | ( n26462 & ~n26463 ) ;
  assign n26465 = ( ~n26462 & n26463 ) | ( ~n26462 & n26464 ) | ( n26463 & n26464 ) ;
  assign n26466 = ( ~n26411 & n26464 ) | ( ~n26411 & n26465 ) | ( n26464 & n26465 ) ;
  assign n26467 = ~n26401 & n26466 ;
  assign n26468 = n26401 & ~n26466 ;
  assign n26469 = n26467 | n26468 ;
  assign n26470 = n4551 & n20562 ;
  assign n26471 = n4546 & ~n20689 ;
  assign n26472 = n4548 & n20560 ;
  assign n26473 = n26471 | n26472 ;
  assign n26474 = n26470 | n26473 ;
  assign n26475 = n4554 | n26474 ;
  assign n26476 = ( ~n21044 & n26474 ) | ( ~n21044 & n26475 ) | ( n26474 & n26475 ) ;
  assign n26477 = ~x23 & n26476 ;
  assign n26478 = x23 | n26477 ;
  assign n26479 = ( ~n26476 & n26477 ) | ( ~n26476 & n26478 ) | ( n26477 & n26478 ) ;
  assign n26480 = n26469 & n26479 ;
  assign n26481 = ( n26401 & ~n26466 ) | ( n26401 & n26479 ) | ( ~n26466 & n26479 ) ;
  assign n26482 = n26467 | n26481 ;
  assign n26483 = ~n26480 & n26482 ;
  assign n26484 = n26313 | n26318 ;
  assign n26485 = n26483 & ~n26484 ;
  assign n26486 = ~n26483 & n26484 ;
  assign n26487 = n26485 | n26486 ;
  assign n26488 = n4781 & ~n20710 ;
  assign n26489 = n4776 & ~n20552 ;
  assign n26490 = n4778 & n20556 ;
  assign n26491 = n26489 | n26490 ;
  assign n26492 = n26488 | n26491 ;
  assign n26493 = n4784 | n26492 ;
  assign n26494 = ( ~n22641 & n26492 ) | ( ~n22641 & n26493 ) | ( n26492 & n26493 ) ;
  assign n26495 = ~x20 & n26494 ;
  assign n26496 = x20 | n26495 ;
  assign n26497 = ( ~n26494 & n26495 ) | ( ~n26494 & n26496 ) | ( n26495 & n26496 ) ;
  assign n26498 = n26487 & n26497 ;
  assign n26499 = ( ~n26483 & n26484 ) | ( ~n26483 & n26497 ) | ( n26484 & n26497 ) ;
  assign n26500 = n26485 | n26499 ;
  assign n26501 = ~n26498 & n26500 ;
  assign n26502 = n26330 | n26334 ;
  assign n26503 = n26501 & ~n26502 ;
  assign n26504 = ~n26501 & n26502 ;
  assign n26505 = n26503 | n26504 ;
  assign n26506 = n5083 & ~n20724 ;
  assign n26507 = n5069 & n20546 ;
  assign n26508 = n5070 & ~n20542 ;
  assign n26509 = n26507 | n26508 ;
  assign n26510 = n26506 | n26509 ;
  assign n26511 = n5074 | n26510 ;
  assign n26512 = ( n23229 & n26510 ) | ( n23229 & n26511 ) | ( n26510 & n26511 ) ;
  assign n26513 = x17 & n26512 ;
  assign n26514 = x17 & ~n26513 ;
  assign n26515 = ( n26512 & ~n26513 ) | ( n26512 & n26514 ) | ( ~n26513 & n26514 ) ;
  assign n26516 = n26505 & n26515 ;
  assign n26517 = ( ~n26501 & n26502 ) | ( ~n26501 & n26515 ) | ( n26502 & n26515 ) ;
  assign n26518 = n26503 | n26517 ;
  assign n26519 = ~n26516 & n26518 ;
  assign n26520 = n26337 | n26341 ;
  assign n26521 = n26519 & ~n26520 ;
  assign n26522 = ~n26519 & n26520 ;
  assign n26523 = n26521 | n26522 ;
  assign n26524 = n7280 & n20838 ;
  assign n26525 = n5384 & ~n20536 ;
  assign n26526 = n7277 & n20532 ;
  assign n26527 = n26525 | n26526 ;
  assign n26528 = n26524 | n26527 ;
  assign n26529 = n39 | n26528 ;
  assign n26530 = ( ~n23712 & n26528 ) | ( ~n23712 & n26529 ) | ( n26528 & n26529 ) ;
  assign n26531 = ~x14 & n26530 ;
  assign n26532 = x14 | n26531 ;
  assign n26533 = ( ~n26530 & n26531 ) | ( ~n26530 & n26532 ) | ( n26531 & n26532 ) ;
  assign n26534 = n26523 & n26533 ;
  assign n26535 = ( ~n26519 & n26520 ) | ( ~n26519 & n26533 ) | ( n26520 & n26533 ) ;
  assign n26536 = n26521 | n26535 ;
  assign n26537 = ~n26534 & n26536 ;
  assign n26538 = n26353 | n26357 ;
  assign n26539 = n26537 & ~n26538 ;
  assign n26540 = ~n26537 & n26538 ;
  assign n26541 = n26539 | n26540 ;
  assign n26542 = n7305 & n24329 ;
  assign n26543 = n7300 & n20921 ;
  assign n26544 = n7302 & ~n21005 ;
  assign n26545 = n26543 | n26544 ;
  assign n26546 = n26542 | n26545 ;
  assign n26547 = ( n7308 & ~n24391 ) | ( n7308 & n24392 ) | ( ~n24391 & n24392 ) ;
  assign n26548 = n26546 | n26547 ;
  assign n26549 = x11 | n26548 ;
  assign n26550 = ~x11 & n26549 ;
  assign n26551 = ( ~n26548 & n26549 ) | ( ~n26548 & n26550 ) | ( n26549 & n26550 ) ;
  assign n26552 = n26541 & n26551 ;
  assign n26553 = ( ~n26537 & n26538 ) | ( ~n26537 & n26551 ) | ( n26538 & n26551 ) ;
  assign n26554 = n26539 | n26553 ;
  assign n26555 = ~n26552 & n26554 ;
  assign n26556 = n26360 | n26364 ;
  assign n26557 = n26555 & ~n26556 ;
  assign n26558 = ~n26555 & n26556 ;
  assign n26559 = n26557 | n26558 ;
  assign n26560 = n5503 & n25187 ;
  assign n26561 = n5512 & ~n24334 ;
  assign n26562 = n5508 & n24324 ;
  assign n26563 = n26561 | n26562 ;
  assign n26564 = n26560 | n26563 ;
  assign n26565 = n5515 | n26564 ;
  assign n26566 = ( n25193 & n26564 ) | ( n25193 & n26565 ) | ( n26564 & n26565 ) ;
  assign n26567 = x8 & n26566 ;
  assign n26568 = x8 & ~n26567 ;
  assign n26569 = ( n26566 & ~n26567 ) | ( n26566 & n26568 ) | ( ~n26567 & n26568 ) ;
  assign n26570 = n26559 & n26569 ;
  assign n26571 = ( ~n26555 & n26556 ) | ( ~n26555 & n26569 ) | ( n26556 & n26569 ) ;
  assign n26572 = n26557 | n26571 ;
  assign n26573 = ~n26570 & n26572 ;
  assign n26574 = n26377 | n26382 ;
  assign n26575 = n26573 & ~n26574 ;
  assign n26576 = ~n26573 & n26574 ;
  assign n26577 = n26575 | n26576 ;
  assign n26578 = n9245 & n25928 ;
  assign n26579 = n8680 & n25442 ;
  assign n26580 = n8681 & ~n25676 ;
  assign n26581 = n26579 | n26580 ;
  assign n26582 = n26578 | n26581 ;
  assign n26583 = n8685 | n26582 ;
  assign n26584 = ( ~n25936 & n26582 ) | ( ~n25936 & n26583 ) | ( n26582 & n26583 ) ;
  assign n26585 = ~x5 & n26584 ;
  assign n26586 = x5 | n26585 ;
  assign n26587 = ( ~n26584 & n26585 ) | ( ~n26584 & n26586 ) | ( n26585 & n26586 ) ;
  assign n26588 = n26577 & n26587 ;
  assign n26589 = ( ~n26573 & n26574 ) | ( ~n26573 & n26587 ) | ( n26574 & n26587 ) ;
  assign n26590 = n26575 | n26589 ;
  assign n26591 = ~n26588 & n26590 ;
  assign n26592 = n26384 | n26387 ;
  assign n26593 = n26591 & ~n26592 ;
  assign n26594 = ~n26591 & n26592 ;
  assign n26595 = n26593 | n26594 ;
  assign n26596 = ~n26392 & n26595 ;
  assign n26597 = ~n26396 & n26596 ;
  assign n26598 = ( n26392 & n26396 ) | ( n26392 & ~n26595 ) | ( n26396 & ~n26595 ) ;
  assign n26599 = n26597 | n26598 ;
  assign n26600 = n26398 & ~n26599 ;
  assign n26601 = ~n26398 & n26599 ;
  assign n26602 = n26600 | n26601 ;
  assign n26603 = n26594 | n26598 ;
  assign n26604 = n9245 & n26156 ;
  assign n26605 = n8680 & ~n25676 ;
  assign n26606 = n8681 & n25928 ;
  assign n26607 = n26605 | n26606 ;
  assign n26608 = n26604 | n26607 ;
  assign n26609 = n8685 | n26608 ;
  assign n26610 = ( n26167 & n26608 ) | ( n26167 & n26609 ) | ( n26608 & n26609 ) ;
  assign n26611 = x5 & n26610 ;
  assign n26612 = x5 & ~n26611 ;
  assign n26613 = ( n26610 & ~n26611 ) | ( n26610 & n26612 ) | ( ~n26611 & n26612 ) ;
  assign n26614 = n5503 & n25442 ;
  assign n26615 = n5512 & n24324 ;
  assign n26616 = n5508 & n25187 ;
  assign n26617 = n26615 | n26616 ;
  assign n26618 = n26614 | n26617 ;
  assign n26619 = n5515 | n26618 ;
  assign n26620 = ( n25452 & n26618 ) | ( n25452 & n26619 ) | ( n26618 & n26619 ) ;
  assign n26621 = x8 & n26620 ;
  assign n26622 = x8 & ~n26621 ;
  assign n26623 = ( n26620 & ~n26621 ) | ( n26620 & n26622 ) | ( ~n26621 & n26622 ) ;
  assign n26624 = n7305 & ~n24334 ;
  assign n26625 = n7300 & ~n21005 ;
  assign n26626 = n7302 & n24329 ;
  assign n26627 = n26625 | n26626 ;
  assign n26628 = n26624 | n26627 ;
  assign n26629 = ( n7308 & ~n24373 ) | ( n7308 & n24376 ) | ( ~n24373 & n24376 ) ;
  assign n26630 = n26628 | n26629 ;
  assign n26631 = x11 | n26630 ;
  assign n26632 = ~x11 & n26631 ;
  assign n26633 = ( ~n26630 & n26631 ) | ( ~n26630 & n26632 ) | ( n26631 & n26632 ) ;
  assign n26634 = n7280 & n20921 ;
  assign n26635 = n5384 & n20532 ;
  assign n26636 = n7277 & n20838 ;
  assign n26637 = n26635 | n26636 ;
  assign n26638 = n26634 | n26637 ;
  assign n26639 = ( n39 & n23691 ) | ( n39 & n23695 ) | ( n23691 & n23695 ) ;
  assign n26640 = n26638 | n26639 ;
  assign n26641 = x14 | n26640 ;
  assign n26642 = ~x14 & n26641 ;
  assign n26643 = ( ~n26640 & n26641 ) | ( ~n26640 & n26642 ) | ( n26641 & n26642 ) ;
  assign n26644 = n5083 & ~n20536 ;
  assign n26645 = n5069 & ~n20542 ;
  assign n26646 = n5070 & ~n20724 ;
  assign n26647 = n26645 | n26646 ;
  assign n26648 = n26644 | n26647 ;
  assign n26649 = ( n5074 & n23213 ) | ( n5074 & ~n23217 ) | ( n23213 & ~n23217 ) ;
  assign n26650 = n26648 | n26649 ;
  assign n26651 = x17 | n26650 ;
  assign n26652 = ~x17 & n26651 ;
  assign n26653 = ( ~n26650 & n26651 ) | ( ~n26650 & n26652 ) | ( n26651 & n26652 ) ;
  assign n26654 = n4781 & n20546 ;
  assign n26655 = n4776 & n20556 ;
  assign n26656 = n4778 & ~n20710 ;
  assign n26657 = n26655 | n26656 ;
  assign n26658 = n26654 | n26657 ;
  assign n26659 = n4784 & ~n21031 ;
  assign n26660 = ( n4784 & n21037 ) | ( n4784 & n26659 ) | ( n21037 & n26659 ) ;
  assign n26661 = n26658 | n26660 ;
  assign n26662 = x20 | n26661 ;
  assign n26663 = ~x20 & n26662 ;
  assign n26664 = ( ~n26661 & n26662 ) | ( ~n26661 & n26663 ) | ( n26662 & n26663 ) ;
  assign n26665 = n302 | n1956 ;
  assign n26666 = n21475 | n26665 ;
  assign n26667 = n2315 | n26666 ;
  assign n26668 = n127 | n476 ;
  assign n26669 = n13931 | n26668 ;
  assign n26670 = n145 | n263 ;
  assign n26671 = n26669 | n26670 ;
  assign n26672 = n26667 | n26671 ;
  assign n26673 = n1492 | n26672 ;
  assign n26674 = n2623 | n26673 ;
  assign n26675 = n13984 | n26674 ;
  assign n26676 = ( n1253 & n1310 ) | ( n1253 & ~n2656 ) | ( n1310 & ~n2656 ) ;
  assign n26677 = n2656 | n26676 ;
  assign n26678 = n2089 | n26677 ;
  assign n26679 = n26675 | n26678 ;
  assign n26680 = n3204 | n4101 ;
  assign n26681 = n249 | n26680 ;
  assign n26682 = n57 | n26681 ;
  assign n26683 = n128 | n26682 ;
  assign n26684 = n207 | n26683 ;
  assign n26685 = n26679 | n26684 ;
  assign n26686 = n26438 & n26685 ;
  assign n26687 = n26438 | n26685 ;
  assign n26688 = ~n26686 & n26687 ;
  assign n26689 = ( n26439 & n26442 ) | ( n26439 & n26688 ) | ( n26442 & n26688 ) ;
  assign n26690 = n26688 & ~n26689 ;
  assign n26691 = ( n26439 & n26442 ) | ( n26439 & ~n26689 ) | ( n26442 & ~n26689 ) ;
  assign n26692 = n26690 | n26691 ;
  assign n26693 = n3744 & ~n20591 ;
  assign n26694 = n3639 & n20600 ;
  assign n26695 = n3727 & ~n20595 ;
  assign n26696 = n26694 | n26695 ;
  assign n26697 = n26693 | n26696 ;
  assign n26698 = n3636 & n21539 ;
  assign n26699 = ( n3636 & n21543 ) | ( n3636 & n26698 ) | ( n21543 & n26698 ) ;
  assign n26700 = n26697 | n26699 ;
  assign n26701 = n26692 & n26700 ;
  assign n26702 = n26692 & ~n26701 ;
  assign n26703 = ~n26692 & n26700 ;
  assign n26704 = n26702 | n26703 ;
  assign n26705 = n26448 | n26460 ;
  assign n26706 = n26704 | n26705 ;
  assign n26707 = n26704 & n26705 ;
  assign n26708 = n26706 & ~n26707 ;
  assign n26709 = n4048 & ~n20584 ;
  assign n26710 = n4043 & n20588 ;
  assign n26711 = n4045 & ~n20580 ;
  assign n26712 = n26710 | n26711 ;
  assign n26713 = n26709 | n26712 ;
  assign n26714 = n4051 | n26713 ;
  assign n26715 = ( ~n21901 & n26713 ) | ( ~n21901 & n26714 ) | ( n26713 & n26714 ) ;
  assign n26716 = ~x29 & n26715 ;
  assign n26717 = x29 | n26716 ;
  assign n26718 = ( ~n26715 & n26716 ) | ( ~n26715 & n26717 ) | ( n26716 & n26717 ) ;
  assign n26719 = n26708 & n26718 ;
  assign n26720 = n26708 & ~n26719 ;
  assign n26721 = ~n26708 & n26718 ;
  assign n26722 = n26720 | n26721 ;
  assign n26723 = n4484 & ~n20689 ;
  assign n26724 = n4479 & ~n20569 ;
  assign n26725 = n4481 & ~n20573 ;
  assign n26726 = n26724 | n26725 ;
  assign n26727 = n26723 | n26726 ;
  assign n26728 = ( n4487 & ~n22192 ) | ( n4487 & n22193 ) | ( ~n22192 & n22193 ) ;
  assign n26729 = n26727 | n26728 ;
  assign n26730 = x26 | n26729 ;
  assign n26731 = ~x26 & n26730 ;
  assign n26732 = ( ~n26729 & n26730 ) | ( ~n26729 & n26731 ) | ( n26730 & n26731 ) ;
  assign n26733 = n26722 & n26732 ;
  assign n26734 = n26722 | n26732 ;
  assign n26735 = ~n26733 & n26734 ;
  assign n26736 = n4551 & ~n20552 ;
  assign n26737 = n4546 & n20560 ;
  assign n26738 = n4548 & n20562 ;
  assign n26739 = n26737 | n26738 ;
  assign n26740 = n26736 | n26739 ;
  assign n26741 = n4554 & ~n22510 ;
  assign n26742 = ( n4554 & n22512 ) | ( n4554 & n26741 ) | ( n22512 & n26741 ) ;
  assign n26743 = n26740 | n26742 ;
  assign n26744 = x23 | n26743 ;
  assign n26745 = ~x23 & n26744 ;
  assign n26746 = ( ~n26743 & n26744 ) | ( ~n26743 & n26745 ) | ( n26744 & n26745 ) ;
  assign n26747 = ( n26465 & n26735 ) | ( n26465 & n26746 ) | ( n26735 & n26746 ) ;
  assign n26748 = ( n26735 & n26746 ) | ( n26735 & ~n26747 ) | ( n26746 & ~n26747 ) ;
  assign n26749 = ( n26465 & ~n26747 ) | ( n26465 & n26748 ) | ( ~n26747 & n26748 ) ;
  assign n26750 = ( n26481 & n26664 ) | ( n26481 & ~n26749 ) | ( n26664 & ~n26749 ) ;
  assign n26751 = ( ~n26481 & n26749 ) | ( ~n26481 & n26750 ) | ( n26749 & n26750 ) ;
  assign n26752 = ( ~n26664 & n26750 ) | ( ~n26664 & n26751 ) | ( n26750 & n26751 ) ;
  assign n26753 = ( n26499 & n26653 ) | ( n26499 & ~n26752 ) | ( n26653 & ~n26752 ) ;
  assign n26754 = ( ~n26499 & n26752 ) | ( ~n26499 & n26753 ) | ( n26752 & n26753 ) ;
  assign n26755 = ( ~n26653 & n26753 ) | ( ~n26653 & n26754 ) | ( n26753 & n26754 ) ;
  assign n26756 = ( n26517 & n26643 ) | ( n26517 & ~n26755 ) | ( n26643 & ~n26755 ) ;
  assign n26757 = ( ~n26517 & n26755 ) | ( ~n26517 & n26756 ) | ( n26755 & n26756 ) ;
  assign n26758 = ( ~n26643 & n26756 ) | ( ~n26643 & n26757 ) | ( n26756 & n26757 ) ;
  assign n26759 = ( n26535 & n26633 ) | ( n26535 & ~n26758 ) | ( n26633 & ~n26758 ) ;
  assign n26760 = ( ~n26535 & n26758 ) | ( ~n26535 & n26759 ) | ( n26758 & n26759 ) ;
  assign n26761 = ( ~n26633 & n26759 ) | ( ~n26633 & n26760 ) | ( n26759 & n26760 ) ;
  assign n26762 = ( n26553 & n26623 ) | ( n26553 & ~n26761 ) | ( n26623 & ~n26761 ) ;
  assign n26763 = ( ~n26553 & n26761 ) | ( ~n26553 & n26762 ) | ( n26761 & n26762 ) ;
  assign n26764 = ( ~n26623 & n26762 ) | ( ~n26623 & n26763 ) | ( n26762 & n26763 ) ;
  assign n26765 = ( n26571 & n26613 ) | ( n26571 & ~n26764 ) | ( n26613 & ~n26764 ) ;
  assign n26766 = ( ~n26571 & n26764 ) | ( ~n26571 & n26765 ) | ( n26764 & n26765 ) ;
  assign n26767 = ( ~n26613 & n26765 ) | ( ~n26613 & n26766 ) | ( n26765 & n26766 ) ;
  assign n26768 = ( n26589 & n26603 ) | ( n26589 & ~n26767 ) | ( n26603 & ~n26767 ) ;
  assign n26769 = ( ~n26589 & n26767 ) | ( ~n26589 & n26768 ) | ( n26767 & n26768 ) ;
  assign n26770 = ( ~n26603 & n26768 ) | ( ~n26603 & n26769 ) | ( n26768 & n26769 ) ;
  assign n26771 = n26600 & n26770 ;
  assign n26772 = n26600 | n26770 ;
  assign n26773 = ~n26771 & n26772 ;
  assign n26774 = n26589 | n26767 ;
  assign n26775 = ( n26571 & n26613 ) | ( n26571 & n26764 ) | ( n26613 & n26764 ) ;
  assign n26776 = n5503 & ~n25676 ;
  assign n26777 = n5512 & n25187 ;
  assign n26778 = n5508 & n25442 ;
  assign n26779 = n26777 | n26778 ;
  assign n26780 = n26776 | n26779 ;
  assign n26781 = n5515 & ~n25690 ;
  assign n26782 = ( n5515 & n25694 ) | ( n5515 & n26781 ) | ( n25694 & n26781 ) ;
  assign n26783 = n26780 | n26782 ;
  assign n26784 = x8 | n26783 ;
  assign n26785 = ~x8 & n26784 ;
  assign n26786 = ( ~n26783 & n26784 ) | ( ~n26783 & n26785 ) | ( n26784 & n26785 ) ;
  assign n26787 = ( n26535 & n26633 ) | ( n26535 & n26758 ) | ( n26633 & n26758 ) ;
  assign n26788 = n7305 & n24324 ;
  assign n26789 = n7300 & n24329 ;
  assign n26790 = n7302 & ~n24334 ;
  assign n26791 = n26789 | n26790 ;
  assign n26792 = n26788 | n26791 ;
  assign n26793 = n7308 & ~n24353 ;
  assign n26794 = ( n7308 & n24356 ) | ( n7308 & n26793 ) | ( n24356 & n26793 ) ;
  assign n26795 = n26792 | n26794 ;
  assign n26796 = x11 | n26795 ;
  assign n26797 = ~x11 & n26796 ;
  assign n26798 = ( ~n26795 & n26796 ) | ( ~n26795 & n26797 ) | ( n26796 & n26797 ) ;
  assign n26799 = ( n26517 & n26643 ) | ( n26517 & n26755 ) | ( n26643 & n26755 ) ;
  assign n26800 = n26719 | n26733 ;
  assign n26801 = n26701 | n26707 ;
  assign n26802 = n3744 & n20588 ;
  assign n26803 = n3639 & ~n20595 ;
  assign n26804 = n3727 & ~n20591 ;
  assign n26805 = n26803 | n26804 ;
  assign n26806 = n26802 | n26805 ;
  assign n26807 = n3636 | n26806 ;
  assign n26808 = ( n21526 & n26806 ) | ( n21526 & n26807 ) | ( n26806 & n26807 ) ;
  assign n26809 = n26686 | n26689 ;
  assign n26810 = n1336 | n2333 ;
  assign n26811 = n1284 | n26810 ;
  assign n26812 = n2001 | n26811 ;
  assign n26813 = n509 | n26812 ;
  assign n26814 = n1434 | n2612 ;
  assign n26815 = n2306 | n13191 ;
  assign n26816 = n26814 | n26815 ;
  assign n26817 = n11152 | n26816 ;
  assign n26818 = n4270 | n26817 ;
  assign n26819 = ( ~n1140 & n3344 ) | ( ~n1140 & n26818 ) | ( n3344 & n26818 ) ;
  assign n26820 = n1140 | n26819 ;
  assign n26821 = n26813 | n26820 ;
  assign n26822 = n373 | n639 ;
  assign n26823 = n498 | n26822 ;
  assign n26824 = n168 | n26823 ;
  assign n26825 = n26821 | n26824 ;
  assign n26826 = ( n26438 & n26809 ) | ( n26438 & ~n26825 ) | ( n26809 & ~n26825 ) ;
  assign n26827 = ( ~n26438 & n26825 ) | ( ~n26438 & n26826 ) | ( n26825 & n26826 ) ;
  assign n26828 = ( ~n26809 & n26826 ) | ( ~n26809 & n26827 ) | ( n26826 & n26827 ) ;
  assign n26829 = n26808 & n26828 ;
  assign n26830 = n26828 & ~n26829 ;
  assign n26831 = ( n26808 & ~n26829 ) | ( n26808 & n26830 ) | ( ~n26829 & n26830 ) ;
  assign n26832 = n26801 | n26831 ;
  assign n26833 = n26801 & n26831 ;
  assign n26834 = n26832 & ~n26833 ;
  assign n26835 = n4048 & ~n20569 ;
  assign n26836 = n4043 & ~n20580 ;
  assign n26837 = n4045 & ~n20584 ;
  assign n26838 = n26836 | n26837 ;
  assign n26839 = n26835 | n26838 ;
  assign n26840 = n4051 & n21884 ;
  assign n26841 = ( n4051 & ~n21889 ) | ( n4051 & n26840 ) | ( ~n21889 & n26840 ) ;
  assign n26842 = n26839 | n26841 ;
  assign n26843 = x29 | n26842 ;
  assign n26844 = ~x29 & n26843 ;
  assign n26845 = ( ~n26842 & n26843 ) | ( ~n26842 & n26844 ) | ( n26843 & n26844 ) ;
  assign n26846 = n26834 & n26845 ;
  assign n26847 = n26834 & ~n26846 ;
  assign n26848 = ~n26834 & n26845 ;
  assign n26849 = n26847 | n26848 ;
  assign n26850 = n4484 & n20560 ;
  assign n26851 = n4479 & ~n20573 ;
  assign n26852 = n4481 & ~n20689 ;
  assign n26853 = n26851 | n26852 ;
  assign n26854 = n26850 | n26853 ;
  assign n26855 = ( n4487 & n22173 ) | ( n4487 & n22176 ) | ( n22173 & n22176 ) ;
  assign n26856 = n26854 | n26855 ;
  assign n26857 = x26 | n26856 ;
  assign n26858 = ~x26 & n26857 ;
  assign n26859 = ( ~n26856 & n26857 ) | ( ~n26856 & n26858 ) | ( n26857 & n26858 ) ;
  assign n26860 = n26849 & n26859 ;
  assign n26861 = n26849 | n26859 ;
  assign n26862 = ~n26860 & n26861 ;
  assign n26863 = n26800 | n26862 ;
  assign n26864 = n4551 & n20556 ;
  assign n26865 = n4546 & n20562 ;
  assign n26866 = n4548 & ~n20552 ;
  assign n26867 = n26865 | n26866 ;
  assign n26868 = n26864 | n26867 ;
  assign n26869 = n4554 | n26868 ;
  assign n26870 = ( ~n22655 & n26868 ) | ( ~n22655 & n26869 ) | ( n26868 & n26869 ) ;
  assign n26871 = ~x23 & n26870 ;
  assign n26872 = x23 | n26871 ;
  assign n26873 = ( ~n26870 & n26871 ) | ( ~n26870 & n26872 ) | ( n26871 & n26872 ) ;
  assign n26874 = ( n26862 & ~n26863 ) | ( n26862 & n26873 ) | ( ~n26863 & n26873 ) ;
  assign n26875 = ( n26800 & ~n26863 ) | ( n26800 & n26874 ) | ( ~n26863 & n26874 ) ;
  assign n26876 = n26747 | n26875 ;
  assign n26877 = ( n26800 & n26862 ) | ( n26800 & n26873 ) | ( n26862 & n26873 ) ;
  assign n26878 = n26863 & ~n26877 ;
  assign n26879 = n26876 | n26878 ;
  assign n26880 = ( n26747 & n26875 ) | ( n26747 & n26878 ) | ( n26875 & n26878 ) ;
  assign n26881 = n26879 & ~n26880 ;
  assign n26882 = n4781 & ~n20542 ;
  assign n26883 = n4776 & ~n20710 ;
  assign n26884 = n4778 & n20546 ;
  assign n26885 = n26883 | n26884 ;
  assign n26886 = n26882 | n26885 ;
  assign n26887 = n4784 | n26886 ;
  assign n26888 = ( ~n23042 & n26886 ) | ( ~n23042 & n26887 ) | ( n26886 & n26887 ) ;
  assign n26889 = ~x20 & n26888 ;
  assign n26890 = x20 | n26889 ;
  assign n26891 = ( ~n26888 & n26889 ) | ( ~n26888 & n26890 ) | ( n26889 & n26890 ) ;
  assign n26892 = n26881 & n26891 ;
  assign n26893 = n26881 & ~n26892 ;
  assign n26894 = ( n26481 & n26664 ) | ( n26481 & n26749 ) | ( n26664 & n26749 ) ;
  assign n26895 = ~n26881 & n26891 ;
  assign n26896 = n26894 | n26895 ;
  assign n26897 = n26893 | n26896 ;
  assign n26898 = ( n26893 & n26894 ) | ( n26893 & n26895 ) | ( n26894 & n26895 ) ;
  assign n26899 = n26897 & ~n26898 ;
  assign n26900 = n5083 & n20532 ;
  assign n26901 = n5069 & ~n20724 ;
  assign n26902 = n5070 & ~n20536 ;
  assign n26903 = n26901 | n26902 ;
  assign n26904 = n26900 | n26903 ;
  assign n26905 = n5074 | n26904 ;
  assign n26906 = ( n23203 & n26904 ) | ( n23203 & n26905 ) | ( n26904 & n26905 ) ;
  assign n26907 = x17 & n26906 ;
  assign n26908 = x17 & ~n26907 ;
  assign n26909 = ( n26906 & ~n26907 ) | ( n26906 & n26908 ) | ( ~n26907 & n26908 ) ;
  assign n26910 = n26899 & n26909 ;
  assign n26911 = n26899 & ~n26910 ;
  assign n26912 = ( n26499 & n26653 ) | ( n26499 & n26752 ) | ( n26653 & n26752 ) ;
  assign n26913 = ~n26899 & n26909 ;
  assign n26914 = n26912 | n26913 ;
  assign n26915 = n26911 | n26914 ;
  assign n26916 = ( n26911 & n26912 ) | ( n26911 & n26913 ) | ( n26912 & n26913 ) ;
  assign n26917 = n26915 & ~n26916 ;
  assign n26918 = n7280 & ~n21005 ;
  assign n26919 = n5384 & n20838 ;
  assign n26920 = n7277 & n20921 ;
  assign n26921 = n26919 | n26920 ;
  assign n26922 = n26918 | n26921 ;
  assign n26923 = n39 | n26922 ;
  assign n26924 = ( ~n21015 & n26922 ) | ( ~n21015 & n26923 ) | ( n26922 & n26923 ) ;
  assign n26925 = ~x14 & n26924 ;
  assign n26926 = x14 | n26925 ;
  assign n26927 = ( ~n26924 & n26925 ) | ( ~n26924 & n26926 ) | ( n26925 & n26926 ) ;
  assign n26928 = n26917 & ~n26927 ;
  assign n26929 = n26927 | n26928 ;
  assign n26930 = ( ~n26917 & n26928 ) | ( ~n26917 & n26929 ) | ( n26928 & n26929 ) ;
  assign n26931 = ( n26798 & n26799 ) | ( n26798 & ~n26930 ) | ( n26799 & ~n26930 ) ;
  assign n26932 = ( ~n26799 & n26930 ) | ( ~n26799 & n26931 ) | ( n26930 & n26931 ) ;
  assign n26933 = ( ~n26798 & n26931 ) | ( ~n26798 & n26932 ) | ( n26931 & n26932 ) ;
  assign n26934 = ( n26786 & n26787 ) | ( n26786 & ~n26933 ) | ( n26787 & ~n26933 ) ;
  assign n26935 = ( ~n26787 & n26933 ) | ( ~n26787 & n26934 ) | ( n26933 & n26934 ) ;
  assign n26936 = ( ~n26786 & n26934 ) | ( ~n26786 & n26935 ) | ( n26934 & n26935 ) ;
  assign n26937 = ( n26553 & n26623 ) | ( n26553 & n26761 ) | ( n26623 & n26761 ) ;
  assign n26938 = n12982 & n26156 ;
  assign n26939 = n8680 & n25928 ;
  assign n26940 = n26938 | n26939 ;
  assign n26941 = n8685 | n26940 ;
  assign n26942 = ( n26165 & n26940 ) | ( n26165 & n26941 ) | ( n26940 & n26941 ) ;
  assign n26943 = x5 & n26942 ;
  assign n26944 = x5 & ~n26943 ;
  assign n26945 = ( n26942 & ~n26943 ) | ( n26942 & n26944 ) | ( ~n26943 & n26944 ) ;
  assign n26946 = ( n26936 & n26937 ) | ( n26936 & ~n26945 ) | ( n26937 & ~n26945 ) ;
  assign n26947 = ( ~n26937 & n26945 ) | ( ~n26937 & n26946 ) | ( n26945 & n26946 ) ;
  assign n26948 = ( ~n26936 & n26946 ) | ( ~n26936 & n26947 ) | ( n26946 & n26947 ) ;
  assign n26949 = n26775 | n26948 ;
  assign n26950 = n26775 & n26948 ;
  assign n26951 = n26949 & ~n26950 ;
  assign n26952 = n26774 & n26951 ;
  assign n26953 = n26589 & n26767 ;
  assign n26954 = n26951 & n26953 ;
  assign n26955 = ( n26603 & n26952 ) | ( n26603 & n26954 ) | ( n26952 & n26954 ) ;
  assign n26956 = ( n26589 & n26603 ) | ( n26589 & n26767 ) | ( n26603 & n26767 ) ;
  assign n26957 = n26951 | n26956 ;
  assign n26958 = ~n26955 & n26957 ;
  assign n26959 = n26771 & n26958 ;
  assign n26960 = n26771 | n26958 ;
  assign n26961 = ~n26959 & n26960 ;
  assign n26962 = ( n26786 & n26787 ) | ( n26786 & n26933 ) | ( n26787 & n26933 ) ;
  assign n26963 = n5503 & n25928 ;
  assign n26964 = n5512 & n25442 ;
  assign n26965 = n5508 & ~n25676 ;
  assign n26966 = n26964 | n26965 ;
  assign n26967 = n26963 | n26966 ;
  assign n26968 = n5515 | n26967 ;
  assign n26969 = ( ~n25936 & n26967 ) | ( ~n25936 & n26968 ) | ( n26967 & n26968 ) ;
  assign n26970 = ~x8 & n26969 ;
  assign n26971 = x8 | n26970 ;
  assign n26972 = ( ~n26969 & n26970 ) | ( ~n26969 & n26971 ) | ( n26970 & n26971 ) ;
  assign n26973 = n26962 & n26972 ;
  assign n26974 = n26962 & ~n26973 ;
  assign n26975 = ( n26915 & n26916 ) | ( n26915 & n26927 ) | ( n26916 & n26927 ) ;
  assign n26976 = n7280 & n24329 ;
  assign n26977 = n5384 & n20921 ;
  assign n26978 = n7277 & ~n21005 ;
  assign n26979 = n26977 | n26978 ;
  assign n26980 = n26976 | n26979 ;
  assign n26981 = ( n39 & ~n24391 ) | ( n39 & n24392 ) | ( ~n24391 & n24392 ) ;
  assign n26982 = n26980 | n26981 ;
  assign n26983 = x14 | n26982 ;
  assign n26984 = ~x14 & n26983 ;
  assign n26985 = ( ~n26982 & n26983 ) | ( ~n26982 & n26984 ) | ( n26983 & n26984 ) ;
  assign n26986 = n26975 & n26985 ;
  assign n26987 = n26975 & ~n26986 ;
  assign n26988 = n26846 | n26860 ;
  assign n26989 = n4484 & n20562 ;
  assign n26990 = n4479 & ~n20689 ;
  assign n26991 = n4481 & n20560 ;
  assign n26992 = n26990 | n26991 ;
  assign n26993 = n26989 | n26992 ;
  assign n26994 = n4487 | n26993 ;
  assign n26995 = ( ~n21044 & n26993 ) | ( ~n21044 & n26994 ) | ( n26993 & n26994 ) ;
  assign n26996 = ~x26 & n26995 ;
  assign n26997 = x26 | n26996 ;
  assign n26998 = ( ~n26995 & n26996 ) | ( ~n26995 & n26997 ) | ( n26996 & n26997 ) ;
  assign n26999 = n4048 & ~n20573 ;
  assign n27000 = n4043 & ~n20584 ;
  assign n27001 = n4045 & ~n20569 ;
  assign n27002 = n27000 | n27001 ;
  assign n27003 = n26999 | n27002 ;
  assign n27004 = n4051 | n27003 ;
  assign n27005 = ( ~n21860 & n27003 ) | ( ~n21860 & n27004 ) | ( n27003 & n27004 ) ;
  assign n27006 = ~x29 & n27005 ;
  assign n27007 = x29 | n27006 ;
  assign n27008 = ( ~n27005 & n27006 ) | ( ~n27005 & n27007 ) | ( n27006 & n27007 ) ;
  assign n27009 = n26829 | n26833 ;
  assign n27010 = n3744 & ~n20580 ;
  assign n27011 = n3639 & ~n20591 ;
  assign n27012 = n3727 & n20588 ;
  assign n27013 = n27011 | n27012 ;
  assign n27014 = n27010 | n27013 ;
  assign n27015 = n3636 | n27014 ;
  assign n27016 = ( n21840 & n27014 ) | ( n21840 & n27015 ) | ( n27014 & n27015 ) ;
  assign n27017 = ( n26438 & n26809 ) | ( n26438 & n26825 ) | ( n26809 & n26825 ) ;
  assign n27018 = n2824 | n3775 ;
  assign n27019 = n2816 | n27018 ;
  assign n27020 = n3149 | n4004 ;
  assign n27021 = n2967 | n27020 ;
  assign n27022 = n82 | n27021 ;
  assign n27023 = n19587 | n27022 ;
  assign n27024 = n11294 | n27023 ;
  assign n27025 = n27019 | n27024 ;
  assign n27026 = n2433 | n3375 ;
  assign n27027 = n66 | n27026 ;
  assign n27028 = n21226 | n27027 ;
  assign n27029 = n528 | n27028 ;
  assign n27030 = n505 | n27029 ;
  assign n27031 = n151 | n27030 ;
  assign n27032 = n27025 | n27031 ;
  assign n27033 = n146 | n27032 ;
  assign n27034 = n12984 & n26156 ;
  assign n27035 = ~x5 & n27034 ;
  assign n27036 = x5 | n27035 ;
  assign n27037 = ( ~n27034 & n27035 ) | ( ~n27034 & n27036 ) | ( n27035 & n27036 ) ;
  assign n27038 = ( n26438 & n27033 ) | ( n26438 & ~n27037 ) | ( n27033 & ~n27037 ) ;
  assign n27039 = ( ~n26438 & n27037 ) | ( ~n26438 & n27038 ) | ( n27037 & n27038 ) ;
  assign n27040 = ( ~n27033 & n27038 ) | ( ~n27033 & n27039 ) | ( n27038 & n27039 ) ;
  assign n27041 = ( n27016 & n27017 ) | ( n27016 & ~n27040 ) | ( n27017 & ~n27040 ) ;
  assign n27042 = ( ~n27017 & n27040 ) | ( ~n27017 & n27041 ) | ( n27040 & n27041 ) ;
  assign n27043 = ( ~n27016 & n27041 ) | ( ~n27016 & n27042 ) | ( n27041 & n27042 ) ;
  assign n27044 = ( n27008 & ~n27009 ) | ( n27008 & n27043 ) | ( ~n27009 & n27043 ) ;
  assign n27045 = ( n27009 & ~n27043 ) | ( n27009 & n27044 ) | ( ~n27043 & n27044 ) ;
  assign n27046 = ( ~n27008 & n27044 ) | ( ~n27008 & n27045 ) | ( n27044 & n27045 ) ;
  assign n27047 = n26998 & n27046 ;
  assign n27048 = n26998 | n27046 ;
  assign n27049 = ~n27047 & n27048 ;
  assign n27050 = n26988 | n27049 ;
  assign n27051 = n26988 & n27049 ;
  assign n27052 = n27050 & ~n27051 ;
  assign n27053 = n4551 & ~n20710 ;
  assign n27054 = n4546 & ~n20552 ;
  assign n27055 = n4548 & n20556 ;
  assign n27056 = n27054 | n27055 ;
  assign n27057 = n27053 | n27056 ;
  assign n27058 = n4554 | n27057 ;
  assign n27059 = ( ~n22641 & n27057 ) | ( ~n22641 & n27058 ) | ( n27057 & n27058 ) ;
  assign n27060 = ~x23 & n27059 ;
  assign n27061 = x23 | n27060 ;
  assign n27062 = ( ~n27059 & n27060 ) | ( ~n27059 & n27061 ) | ( n27060 & n27061 ) ;
  assign n27063 = n27052 & n27062 ;
  assign n27064 = n27052 & ~n27063 ;
  assign n27065 = ~n27052 & n27062 ;
  assign n27066 = n26877 | n27065 ;
  assign n27067 = n27064 | n27066 ;
  assign n27068 = ( n26877 & n27064 ) | ( n26877 & n27065 ) | ( n27064 & n27065 ) ;
  assign n27069 = n27067 & ~n27068 ;
  assign n27070 = n4781 & ~n20724 ;
  assign n27071 = n4776 & n20546 ;
  assign n27072 = n4778 & ~n20542 ;
  assign n27073 = n27071 | n27072 ;
  assign n27074 = n27070 | n27073 ;
  assign n27075 = n4784 | n27074 ;
  assign n27076 = ( n23229 & n27074 ) | ( n23229 & n27075 ) | ( n27074 & n27075 ) ;
  assign n27077 = x20 & n27076 ;
  assign n27078 = x20 & ~n27077 ;
  assign n27079 = ( n27076 & ~n27077 ) | ( n27076 & n27078 ) | ( ~n27077 & n27078 ) ;
  assign n27080 = n27069 & n27079 ;
  assign n27081 = n27069 & ~n27080 ;
  assign n27082 = ~n27069 & n27079 ;
  assign n27083 = n26880 | n26892 ;
  assign n27084 = n27082 | n27083 ;
  assign n27085 = n27081 | n27084 ;
  assign n27086 = ( n27081 & n27082 ) | ( n27081 & n27083 ) | ( n27082 & n27083 ) ;
  assign n27087 = n27085 & ~n27086 ;
  assign n27088 = n5083 & n20838 ;
  assign n27089 = n5069 & ~n20536 ;
  assign n27090 = n5070 & n20532 ;
  assign n27091 = n27089 | n27090 ;
  assign n27092 = n27088 | n27091 ;
  assign n27093 = n5074 | n27092 ;
  assign n27094 = ( ~n23712 & n27092 ) | ( ~n23712 & n27093 ) | ( n27092 & n27093 ) ;
  assign n27095 = ~x17 & n27094 ;
  assign n27096 = x17 | n27095 ;
  assign n27097 = ( ~n27094 & n27095 ) | ( ~n27094 & n27096 ) | ( n27095 & n27096 ) ;
  assign n27098 = n27087 & n27097 ;
  assign n27099 = n27087 & ~n27098 ;
  assign n27100 = ~n27087 & n27097 ;
  assign n27101 = n26898 | n26910 ;
  assign n27102 = n27100 | n27101 ;
  assign n27103 = n27099 | n27102 ;
  assign n27104 = ( n27099 & n27100 ) | ( n27099 & n27101 ) | ( n27100 & n27101 ) ;
  assign n27105 = n27103 & ~n27104 ;
  assign n27106 = ~n26975 & n26985 ;
  assign n27107 = n27105 | n27106 ;
  assign n27108 = n26987 | n27107 ;
  assign n27109 = ( n26987 & n27105 ) | ( n26987 & n27106 ) | ( n27105 & n27106 ) ;
  assign n27110 = n27108 & ~n27109 ;
  assign n27111 = n7305 & n25187 ;
  assign n27112 = n7300 & ~n24334 ;
  assign n27113 = n7302 & n24324 ;
  assign n27114 = n27112 | n27113 ;
  assign n27115 = n27111 | n27114 ;
  assign n27116 = n7308 | n27115 ;
  assign n27117 = ( n25193 & n27115 ) | ( n25193 & n27116 ) | ( n27115 & n27116 ) ;
  assign n27118 = x11 & n27117 ;
  assign n27119 = x11 & ~n27118 ;
  assign n27120 = ( n27117 & ~n27118 ) | ( n27117 & n27119 ) | ( ~n27118 & n27119 ) ;
  assign n27121 = n27110 & n27120 ;
  assign n27122 = n27110 & ~n27121 ;
  assign n27123 = ( n26798 & n26799 ) | ( n26798 & n26930 ) | ( n26799 & n26930 ) ;
  assign n27124 = ~n27110 & n27120 ;
  assign n27125 = n27123 | n27124 ;
  assign n27126 = n27122 | n27125 ;
  assign n27127 = ( n27122 & n27123 ) | ( n27122 & n27124 ) | ( n27123 & n27124 ) ;
  assign n27128 = n27126 & ~n27127 ;
  assign n27129 = ~n26962 & n26972 ;
  assign n27130 = n27128 | n27129 ;
  assign n27131 = n26974 | n27130 ;
  assign n27132 = ( n26974 & n27128 ) | ( n26974 & n27129 ) | ( n27128 & n27129 ) ;
  assign n27133 = n27131 & ~n27132 ;
  assign n27134 = ( n26936 & n26937 ) | ( n26936 & n26945 ) | ( n26937 & n26945 ) ;
  assign n27135 = n27133 & n27134 ;
  assign n27136 = n27133 | n27134 ;
  assign n27137 = ~n27135 & n27136 ;
  assign n27138 = n26950 | n26952 ;
  assign n27139 = n26950 | n26954 ;
  assign n27140 = ( n26603 & n27138 ) | ( n26603 & n27139 ) | ( n27138 & n27139 ) ;
  assign n27141 = n27137 | n27140 ;
  assign n27142 = n27137 & n27140 ;
  assign n27143 = n27141 & ~n27142 ;
  assign n27144 = n26959 | n27143 ;
  assign n27145 = n26958 & n27143 ;
  assign n27146 = n26771 & n27145 ;
  assign n27147 = n27144 & ~n27146 ;
  assign n27148 = n27135 | n27142 ;
  assign n27149 = n27121 | n27127 ;
  assign n27150 = n27098 | n27104 ;
  assign n27151 = n4781 & ~n20536 ;
  assign n27152 = n4776 & ~n20542 ;
  assign n27153 = n4778 & ~n20724 ;
  assign n27154 = n27152 | n27153 ;
  assign n27155 = n27151 | n27154 ;
  assign n27156 = ( n4784 & n23213 ) | ( n4784 & ~n23217 ) | ( n23213 & ~n23217 ) ;
  assign n27157 = n27155 | n27156 ;
  assign n27158 = x20 | n27157 ;
  assign n27159 = ~x20 & n27158 ;
  assign n27160 = ( ~n27157 & n27158 ) | ( ~n27157 & n27159 ) | ( n27158 & n27159 ) ;
  assign n27161 = n27063 | n27068 ;
  assign n27162 = n4551 & n20546 ;
  assign n27163 = n4546 & n20556 ;
  assign n27164 = n4548 & ~n20710 ;
  assign n27165 = n27163 | n27164 ;
  assign n27166 = n27162 | n27165 ;
  assign n27167 = n4554 & ~n21031 ;
  assign n27168 = ( n4554 & n21037 ) | ( n4554 & n27167 ) | ( n21037 & n27167 ) ;
  assign n27169 = n27166 | n27168 ;
  assign n27170 = x23 | n27169 ;
  assign n27171 = ~x23 & n27170 ;
  assign n27172 = ( ~n27169 & n27170 ) | ( ~n27169 & n27171 ) | ( n27170 & n27171 ) ;
  assign n27173 = n27047 | n27051 ;
  assign n27174 = n4484 & ~n20552 ;
  assign n27175 = n4479 & n20560 ;
  assign n27176 = n4481 & n20562 ;
  assign n27177 = n27175 | n27176 ;
  assign n27178 = n27174 | n27177 ;
  assign n27179 = n4487 & ~n22510 ;
  assign n27180 = ( n4487 & n22512 ) | ( n4487 & n27179 ) | ( n22512 & n27179 ) ;
  assign n27181 = n27178 | n27180 ;
  assign n27182 = x26 | n27181 ;
  assign n27183 = ~x26 & n27182 ;
  assign n27184 = ( ~n27181 & n27182 ) | ( ~n27181 & n27183 ) | ( n27182 & n27183 ) ;
  assign n27185 = ( n27008 & n27009 ) | ( n27008 & n27043 ) | ( n27009 & n27043 ) ;
  assign n27186 = n3744 & ~n20584 ;
  assign n27187 = n3639 & n20588 ;
  assign n27188 = n3727 & ~n20580 ;
  assign n27189 = n27187 | n27188 ;
  assign n27190 = n27186 | n27189 ;
  assign n27191 = n3636 | n27190 ;
  assign n27192 = ( ~n21901 & n27190 ) | ( ~n21901 & n27191 ) | ( n27190 & n27191 ) ;
  assign n27193 = n473 | n1469 ;
  assign n27194 = n5195 | n27193 ;
  assign n27195 = n1395 | n1513 ;
  assign n27196 = n27194 | n27195 ;
  assign n27197 = n1078 | n5701 ;
  assign n27198 = n27196 | n27197 ;
  assign n27199 = n856 | n1310 ;
  assign n27200 = n27198 | n27199 ;
  assign n27201 = n952 | n1692 ;
  assign n27202 = n4879 | n27201 ;
  assign n27203 = n5614 | n27202 ;
  assign n27204 = n432 | n1354 ;
  assign n27205 = n249 | n27204 ;
  assign n27206 = n269 | n27205 ;
  assign n27207 = n416 | n27206 ;
  assign n27208 = n27203 | n27207 ;
  assign n27209 = n27200 | n27208 ;
  assign n27210 = n2665 | n2930 ;
  assign n27211 = n1219 | n27210 ;
  assign n27212 = n27209 | n27211 ;
  assign n27213 = n3293 | n27212 ;
  assign n27214 = n959 | n995 ;
  assign n27215 = n2943 | n27214 ;
  assign n27216 = n373 | n27215 ;
  assign n27217 = n431 | n27216 ;
  assign n27218 = n253 | n27217 ;
  assign n27219 = n383 | n27218 ;
  assign n27220 = n190 | n27219 ;
  assign n27221 = n441 | n27220 ;
  assign n27222 = n27213 | n27221 ;
  assign n27223 = n224 | n27222 ;
  assign n27224 = ( n26438 & n27037 ) | ( n26438 & n27040 ) | ( n27037 & n27040 ) ;
  assign n27225 = n27223 | n27224 ;
  assign n27226 = n27223 & n27224 ;
  assign n27227 = n27225 & ~n27226 ;
  assign n27228 = n27192 & n27227 ;
  assign n27229 = n27227 & ~n27228 ;
  assign n27230 = ( n27192 & ~n27228 ) | ( n27192 & n27229 ) | ( ~n27228 & n27229 ) ;
  assign n27231 = ( n27016 & n27017 ) | ( n27016 & n27040 ) | ( n27017 & n27040 ) ;
  assign n27232 = n27230 | n27231 ;
  assign n27233 = n27230 & n27231 ;
  assign n27234 = n27232 & ~n27233 ;
  assign n27235 = n4048 & ~n20689 ;
  assign n27236 = n4043 & ~n20569 ;
  assign n27237 = n4045 & ~n20573 ;
  assign n27238 = n27236 | n27237 ;
  assign n27239 = n27235 | n27238 ;
  assign n27240 = n4051 & ~n22193 ;
  assign n27241 = n22192 & n27240 ;
  assign n27242 = ( n4051 & n27239 ) | ( n4051 & ~n27241 ) | ( n27239 & ~n27241 ) ;
  assign n27243 = x29 & n27242 ;
  assign n27244 = x29 & ~n27243 ;
  assign n27245 = ( n27242 & ~n27243 ) | ( n27242 & n27244 ) | ( ~n27243 & n27244 ) ;
  assign n27246 = n27234 & n27245 ;
  assign n27247 = n27234 | n27245 ;
  assign n27248 = ~n27246 & n27247 ;
  assign n27249 = ( n27184 & n27185 ) | ( n27184 & ~n27248 ) | ( n27185 & ~n27248 ) ;
  assign n27250 = ( ~n27185 & n27248 ) | ( ~n27185 & n27249 ) | ( n27248 & n27249 ) ;
  assign n27251 = ( ~n27184 & n27249 ) | ( ~n27184 & n27250 ) | ( n27249 & n27250 ) ;
  assign n27252 = ( n27172 & ~n27173 ) | ( n27172 & n27251 ) | ( ~n27173 & n27251 ) ;
  assign n27253 = ( n27173 & ~n27251 ) | ( n27173 & n27252 ) | ( ~n27251 & n27252 ) ;
  assign n27254 = ( ~n27172 & n27252 ) | ( ~n27172 & n27253 ) | ( n27252 & n27253 ) ;
  assign n27255 = ( n27160 & ~n27161 ) | ( n27160 & n27254 ) | ( ~n27161 & n27254 ) ;
  assign n27256 = ( n27161 & ~n27254 ) | ( n27161 & n27255 ) | ( ~n27254 & n27255 ) ;
  assign n27257 = ( ~n27160 & n27255 ) | ( ~n27160 & n27256 ) | ( n27255 & n27256 ) ;
  assign n27258 = n27080 | n27086 ;
  assign n27259 = n27257 | n27258 ;
  assign n27260 = n5083 & n20921 ;
  assign n27261 = n5069 & n20532 ;
  assign n27262 = n5070 & n20838 ;
  assign n27263 = n27261 | n27262 ;
  assign n27264 = n27260 | n27263 ;
  assign n27265 = ( n5074 & n23691 ) | ( n5074 & n23695 ) | ( n23691 & n23695 ) ;
  assign n27266 = n27264 | n27265 ;
  assign n27267 = x17 | n27266 ;
  assign n27268 = ~x17 & n27267 ;
  assign n27269 = ( ~n27266 & n27267 ) | ( ~n27266 & n27268 ) | ( n27267 & n27268 ) ;
  assign n27270 = ( n27258 & ~n27259 ) | ( n27258 & n27269 ) | ( ~n27259 & n27269 ) ;
  assign n27271 = ( n27257 & ~n27259 ) | ( n27257 & n27270 ) | ( ~n27259 & n27270 ) ;
  assign n27272 = n27150 | n27271 ;
  assign n27273 = ( n27257 & n27258 ) | ( n27257 & n27269 ) | ( n27258 & n27269 ) ;
  assign n27274 = n27259 & ~n27273 ;
  assign n27275 = n27272 | n27274 ;
  assign n27276 = ( n27150 & n27271 ) | ( n27150 & n27274 ) | ( n27271 & n27274 ) ;
  assign n27277 = n27275 & ~n27276 ;
  assign n27278 = n7280 & ~n24334 ;
  assign n27279 = n5384 & ~n21005 ;
  assign n27280 = n7277 & n24329 ;
  assign n27281 = n27279 | n27280 ;
  assign n27282 = n27278 | n27281 ;
  assign n27283 = ( n39 & ~n24373 ) | ( n39 & n24376 ) | ( ~n24373 & n24376 ) ;
  assign n27284 = n27282 | n27283 ;
  assign n27285 = x14 | n27284 ;
  assign n27286 = ~x14 & n27285 ;
  assign n27287 = ( ~n27284 & n27285 ) | ( ~n27284 & n27286 ) | ( n27285 & n27286 ) ;
  assign n27288 = n27277 & n27287 ;
  assign n27289 = n27277 & ~n27288 ;
  assign n27290 = ~n27277 & n27287 ;
  assign n27291 = n27289 | n27290 ;
  assign n27292 = n26986 | n27109 ;
  assign n27293 = n27291 & n27292 ;
  assign n27294 = n27291 | n27292 ;
  assign n27295 = ~n27293 & n27294 ;
  assign n27296 = n7305 & n25442 ;
  assign n27297 = n7300 & n24324 ;
  assign n27298 = n7302 & n25187 ;
  assign n27299 = n27297 | n27298 ;
  assign n27300 = n27296 | n27299 ;
  assign n27301 = n7308 | n27300 ;
  assign n27302 = ( n25452 & n27300 ) | ( n25452 & n27301 ) | ( n27300 & n27301 ) ;
  assign n27303 = x11 & n27302 ;
  assign n27304 = x11 & ~n27303 ;
  assign n27305 = ( n27302 & ~n27303 ) | ( n27302 & n27304 ) | ( ~n27303 & n27304 ) ;
  assign n27306 = ~n27295 & n27305 ;
  assign n27307 = n27149 | n27306 ;
  assign n27308 = n27295 & ~n27305 ;
  assign n27309 = n27307 | n27308 ;
  assign n27310 = ( n27149 & n27306 ) | ( n27149 & n27308 ) | ( n27306 & n27308 ) ;
  assign n27311 = n27309 & ~n27310 ;
  assign n27312 = n5503 & n26156 ;
  assign n27313 = n5512 & ~n25676 ;
  assign n27314 = n5508 & n25928 ;
  assign n27315 = n27313 | n27314 ;
  assign n27316 = n27312 | n27315 ;
  assign n27317 = n5515 | n27316 ;
  assign n27318 = ( n26167 & n27316 ) | ( n26167 & n27317 ) | ( n27316 & n27317 ) ;
  assign n27319 = x8 & n27318 ;
  assign n27320 = x8 & ~n27319 ;
  assign n27321 = ( n27318 & ~n27319 ) | ( n27318 & n27320 ) | ( ~n27319 & n27320 ) ;
  assign n27322 = n27311 & ~n27321 ;
  assign n27323 = n27321 | n27322 ;
  assign n27324 = ( ~n27311 & n27322 ) | ( ~n27311 & n27323 ) | ( n27322 & n27323 ) ;
  assign n27325 = n26973 | n27132 ;
  assign n27326 = ( n27148 & n27324 ) | ( n27148 & ~n27325 ) | ( n27324 & ~n27325 ) ;
  assign n27327 = ( ~n27324 & n27325 ) | ( ~n27324 & n27326 ) | ( n27325 & n27326 ) ;
  assign n27328 = ( ~n27148 & n27326 ) | ( ~n27148 & n27327 ) | ( n27326 & n27327 ) ;
  assign n27329 = n27146 & n27328 ;
  assign n27330 = n27146 & ~n27329 ;
  assign n27331 = ( n27328 & ~n27329 ) | ( n27328 & n27330 ) | ( ~n27329 & n27330 ) ;
  assign n27332 = n27324 & n27325 ;
  assign n27333 = ( n27160 & n27161 ) | ( n27160 & n27254 ) | ( n27161 & n27254 ) ;
  assign n27334 = ( n27172 & n27173 ) | ( n27172 & n27251 ) | ( n27173 & n27251 ) ;
  assign n27335 = n4484 & n20556 ;
  assign n27336 = n4479 & n20562 ;
  assign n27337 = n4481 & ~n20552 ;
  assign n27338 = n27336 | n27337 ;
  assign n27339 = n27335 | n27338 ;
  assign n27340 = n4487 | n27339 ;
  assign n27341 = ( ~n22655 & n27339 ) | ( ~n22655 & n27340 ) | ( n27339 & n27340 ) ;
  assign n27342 = ~x26 & n27341 ;
  assign n27343 = x26 | n27342 ;
  assign n27344 = ( ~n27341 & n27342 ) | ( ~n27341 & n27343 ) | ( n27342 & n27343 ) ;
  assign n27345 = n4048 & n20560 ;
  assign n27346 = n4043 & ~n20573 ;
  assign n27347 = n4045 & ~n20689 ;
  assign n27348 = n27346 | n27347 ;
  assign n27349 = n27345 | n27348 ;
  assign n27350 = ( n4051 & n22173 ) | ( n4051 & n22176 ) | ( n22173 & n22176 ) ;
  assign n27351 = n27349 | n27350 ;
  assign n27352 = x29 | n27351 ;
  assign n27353 = ~x29 & n27352 ;
  assign n27354 = ( ~n27351 & n27352 ) | ( ~n27351 & n27353 ) | ( n27352 & n27353 ) ;
  assign n27355 = n13357 | n19736 ;
  assign n27356 = n4138 | n27355 ;
  assign n27357 = n2332 | n10900 ;
  assign n27358 = n1287 | n27357 ;
  assign n27359 = n2362 | n3792 ;
  assign n27360 = n571 | n27359 ;
  assign n27361 = n27358 | n27360 ;
  assign n27362 = ~n1260 & n2322 ;
  assign n27363 = ~n27361 & n27362 ;
  assign n27364 = n299 | n655 ;
  assign n27365 = n125 | n27364 ;
  assign n27366 = n608 | n27365 ;
  assign n27367 = n595 | n27366 ;
  assign n27368 = n27363 & ~n27367 ;
  assign n27369 = ~n5805 & n27368 ;
  assign n27370 = ~n27356 & n27369 ;
  assign n27371 = n350 | n639 ;
  assign n27372 = n320 | n338 ;
  assign n27373 = n27371 | n27372 ;
  assign n27374 = n190 | n580 ;
  assign n27375 = n173 | n27374 ;
  assign n27376 = n27373 | n27375 ;
  assign n27377 = n94 | n661 ;
  assign n27378 = n27376 | n27377 ;
  assign n27379 = n11302 | n27378 ;
  assign n27380 = n11222 | n27379 ;
  assign n27381 = n531 | n27380 ;
  assign n27382 = n511 | n27381 ;
  assign n27383 = n327 | n27382 ;
  assign n27384 = n27370 & ~n27383 ;
  assign n27385 = n194 | n199 ;
  assign n27386 = n213 | n27385 ;
  assign n27387 = n181 | n27386 ;
  assign n27388 = n143 | n27387 ;
  assign n27389 = n27384 & ~n27388 ;
  assign n27390 = n27223 & n27389 ;
  assign n27391 = n27223 | n27389 ;
  assign n27392 = ~n27390 & n27391 ;
  assign n27393 = ( ~n27225 & n27228 ) | ( ~n27225 & n27392 ) | ( n27228 & n27392 ) ;
  assign n27394 = ( n27226 & n27229 ) | ( n27226 & ~n27392 ) | ( n27229 & ~n27392 ) ;
  assign n27395 = n27393 | n27394 ;
  assign n27396 = n3744 & ~n20569 ;
  assign n27397 = n3639 & ~n20580 ;
  assign n27398 = n3727 & ~n20584 ;
  assign n27399 = n27397 | n27398 ;
  assign n27400 = n27396 | n27399 ;
  assign n27401 = n3636 & n21884 ;
  assign n27402 = ( n3636 & ~n21889 ) | ( n3636 & n27401 ) | ( ~n21889 & n27401 ) ;
  assign n27403 = n27400 | n27402 ;
  assign n27404 = ~n27395 & n27403 ;
  assign n27405 = n27395 | n27404 ;
  assign n27406 = n27395 & n27403 ;
  assign n27407 = n27405 & ~n27406 ;
  assign n27408 = n27233 | n27246 ;
  assign n27409 = n27407 & ~n27408 ;
  assign n27410 = ~n27407 & n27408 ;
  assign n27411 = n27409 | n27410 ;
  assign n27412 = n27354 & ~n27411 ;
  assign n27413 = n27411 | n27412 ;
  assign n27414 = ( ~n27354 & n27412 ) | ( ~n27354 & n27413 ) | ( n27412 & n27413 ) ;
  assign n27415 = n27344 & ~n27414 ;
  assign n27416 = ~n27344 & n27414 ;
  assign n27417 = n27415 | n27416 ;
  assign n27418 = ( n27184 & n27185 ) | ( n27184 & n27248 ) | ( n27185 & n27248 ) ;
  assign n27419 = n27417 & ~n27418 ;
  assign n27420 = ~n27417 & n27418 ;
  assign n27421 = n27419 | n27420 ;
  assign n27422 = n4551 & ~n20542 ;
  assign n27423 = n4546 & ~n20710 ;
  assign n27424 = n4548 & n20546 ;
  assign n27425 = n27423 | n27424 ;
  assign n27426 = n27422 | n27425 ;
  assign n27427 = n4554 | n27426 ;
  assign n27428 = ( ~n23042 & n27426 ) | ( ~n23042 & n27427 ) | ( n27426 & n27427 ) ;
  assign n27429 = ~x23 & n27428 ;
  assign n27430 = x23 | n27429 ;
  assign n27431 = ( ~n27428 & n27429 ) | ( ~n27428 & n27430 ) | ( n27429 & n27430 ) ;
  assign n27432 = n27421 & n27431 ;
  assign n27433 = ( ~n27417 & n27418 ) | ( ~n27417 & n27431 ) | ( n27418 & n27431 ) ;
  assign n27434 = n27419 | n27433 ;
  assign n27435 = ~n27432 & n27434 ;
  assign n27436 = ~n27334 & n27435 ;
  assign n27437 = n27334 & ~n27435 ;
  assign n27438 = n27436 | n27437 ;
  assign n27439 = n4781 & n20532 ;
  assign n27440 = n4776 & ~n20724 ;
  assign n27441 = n4778 & ~n20536 ;
  assign n27442 = n27440 | n27441 ;
  assign n27443 = n27439 | n27442 ;
  assign n27444 = n4784 | n27443 ;
  assign n27445 = ( n23203 & n27443 ) | ( n23203 & n27444 ) | ( n27443 & n27444 ) ;
  assign n27446 = x20 & n27445 ;
  assign n27447 = x20 & ~n27446 ;
  assign n27448 = ( n27445 & ~n27446 ) | ( n27445 & n27447 ) | ( ~n27446 & n27447 ) ;
  assign n27449 = n27438 & n27448 ;
  assign n27450 = ( n27334 & ~n27435 ) | ( n27334 & n27448 ) | ( ~n27435 & n27448 ) ;
  assign n27451 = n27436 | n27450 ;
  assign n27452 = ~n27449 & n27451 ;
  assign n27453 = ~n27333 & n27452 ;
  assign n27454 = n27333 & ~n27452 ;
  assign n27455 = n27453 | n27454 ;
  assign n27456 = n5083 & ~n21005 ;
  assign n27457 = n5069 & n20838 ;
  assign n27458 = n5070 & n20921 ;
  assign n27459 = n27457 | n27458 ;
  assign n27460 = n27456 | n27459 ;
  assign n27461 = n5074 | n27460 ;
  assign n27462 = ( ~n21015 & n27460 ) | ( ~n21015 & n27461 ) | ( n27460 & n27461 ) ;
  assign n27463 = ~x17 & n27462 ;
  assign n27464 = x17 | n27463 ;
  assign n27465 = ( ~n27462 & n27463 ) | ( ~n27462 & n27464 ) | ( n27463 & n27464 ) ;
  assign n27466 = n27455 & n27465 ;
  assign n27467 = ( n27333 & ~n27452 ) | ( n27333 & n27465 ) | ( ~n27452 & n27465 ) ;
  assign n27468 = n27453 | n27467 ;
  assign n27469 = ~n27466 & n27468 ;
  assign n27470 = ~n27273 & n27469 ;
  assign n27471 = n27273 & ~n27469 ;
  assign n27472 = n27470 | n27471 ;
  assign n27473 = n7280 & n24324 ;
  assign n27474 = n5384 & n24329 ;
  assign n27475 = n7277 & ~n24334 ;
  assign n27476 = n27474 | n27475 ;
  assign n27477 = n27473 | n27476 ;
  assign n27478 = n39 & ~n24353 ;
  assign n27479 = ( n39 & n24356 ) | ( n39 & n27478 ) | ( n24356 & n27478 ) ;
  assign n27480 = n27477 | n27479 ;
  assign n27481 = x14 | n27480 ;
  assign n27482 = ~x14 & n27481 ;
  assign n27483 = ( ~n27480 & n27481 ) | ( ~n27480 & n27482 ) | ( n27481 & n27482 ) ;
  assign n27484 = n27472 & n27483 ;
  assign n27485 = n27276 | n27288 ;
  assign n27486 = n27484 | n27485 ;
  assign n27487 = ( n27273 & ~n27469 ) | ( n27273 & n27483 ) | ( ~n27469 & n27483 ) ;
  assign n27488 = n27470 | n27487 ;
  assign n27489 = ~n27486 & n27488 ;
  assign n27490 = ( n27484 & n27485 ) | ( n27484 & ~n27488 ) | ( n27485 & ~n27488 ) ;
  assign n27491 = n27489 | n27490 ;
  assign n27492 = n7305 & ~n25676 ;
  assign n27493 = n7300 & n25187 ;
  assign n27494 = n7302 & n25442 ;
  assign n27495 = n27493 | n27494 ;
  assign n27496 = n27492 | n27495 ;
  assign n27497 = n7308 & ~n25690 ;
  assign n27498 = ( n7308 & n25694 ) | ( n7308 & n27497 ) | ( n25694 & n27497 ) ;
  assign n27499 = n27496 | n27498 ;
  assign n27500 = x11 | n27499 ;
  assign n27501 = ~x11 & n27500 ;
  assign n27502 = ( ~n27499 & n27500 ) | ( ~n27499 & n27501 ) | ( n27500 & n27501 ) ;
  assign n27503 = n27491 | n27502 ;
  assign n27504 = ~n27502 & n27503 ;
  assign n27505 = ( ~n27491 & n27503 ) | ( ~n27491 & n27504 ) | ( n27503 & n27504 ) ;
  assign n27506 = n12701 & n26156 ;
  assign n27507 = n5512 & n25928 ;
  assign n27508 = n27506 | n27507 ;
  assign n27509 = n5515 | n27508 ;
  assign n27510 = ( n26165 & n27508 ) | ( n26165 & n27509 ) | ( n27508 & n27509 ) ;
  assign n27511 = x8 & n27510 ;
  assign n27512 = x8 & ~n27511 ;
  assign n27513 = ( n27510 & ~n27511 ) | ( n27510 & n27512 ) | ( ~n27511 & n27512 ) ;
  assign n27514 = ( n27293 & n27295 ) | ( n27293 & ~n27308 ) | ( n27295 & ~n27308 ) ;
  assign n27515 = n27513 & n27514 ;
  assign n27516 = n27513 | n27514 ;
  assign n27517 = ~n27515 & n27516 ;
  assign n27518 = ~n27505 & n27517 ;
  assign n27519 = n27505 | n27518 ;
  assign n27520 = n27517 & ~n27518 ;
  assign n27521 = n27519 & ~n27520 ;
  assign n27522 = ( n27309 & n27310 ) | ( n27309 & n27321 ) | ( n27310 & n27321 ) ;
  assign n27523 = n27521 & ~n27522 ;
  assign n27524 = ~n27521 & n27522 ;
  assign n27525 = n27523 | n27524 ;
  assign n27526 = n27332 & ~n27525 ;
  assign n27527 = n27324 & ~n27332 ;
  assign n27528 = ( n27325 & ~n27525 ) | ( n27325 & n27527 ) | ( ~n27525 & n27527 ) ;
  assign n27529 = ( n27148 & n27526 ) | ( n27148 & n27528 ) | ( n27526 & n27528 ) ;
  assign n27530 = ( n27148 & n27324 ) | ( n27148 & n27325 ) | ( n27324 & n27325 ) ;
  assign n27531 = n27525 & ~n27530 ;
  assign n27532 = n27529 | n27531 ;
  assign n27533 = ~n27329 & n27532 ;
  assign n27534 = ( n27329 & ~n27532 ) | ( n27329 & n27533 ) | ( ~n27532 & n27533 ) ;
  assign n27535 = n27533 | n27534 ;
  assign n27536 = n27515 | n27518 ;
  assign n27537 = ( n27486 & n27502 ) | ( n27486 & n27505 ) | ( n27502 & n27505 ) ;
  assign n27538 = n7305 & n25928 ;
  assign n27539 = n7300 & n25442 ;
  assign n27540 = n7302 & ~n25676 ;
  assign n27541 = n27539 | n27540 ;
  assign n27542 = n27538 | n27541 ;
  assign n27543 = n7308 | n27542 ;
  assign n27544 = ( ~n25936 & n27542 ) | ( ~n25936 & n27543 ) | ( n27542 & n27543 ) ;
  assign n27545 = ~x11 & n27544 ;
  assign n27546 = x11 | n27545 ;
  assign n27547 = ( ~n27544 & n27545 ) | ( ~n27544 & n27546 ) | ( n27545 & n27546 ) ;
  assign n27548 = n27537 & n27547 ;
  assign n27549 = n27537 & ~n27548 ;
  assign n27550 = n5083 & n24329 ;
  assign n27551 = n5069 & n20921 ;
  assign n27552 = n5070 & ~n21005 ;
  assign n27553 = n27551 | n27552 ;
  assign n27554 = n27550 | n27553 ;
  assign n27555 = ( n5074 & ~n24391 ) | ( n5074 & n24392 ) | ( ~n24391 & n24392 ) ;
  assign n27556 = n27554 | n27555 ;
  assign n27557 = x17 | n27556 ;
  assign n27558 = ~x17 & n27557 ;
  assign n27559 = ( ~n27556 & n27557 ) | ( ~n27556 & n27558 ) | ( n27557 & n27558 ) ;
  assign n27560 = n27467 & n27559 ;
  assign n27561 = n27467 & ~n27560 ;
  assign n27562 = n4781 & n20838 ;
  assign n27563 = n4776 & ~n20536 ;
  assign n27564 = n4778 & n20532 ;
  assign n27565 = n27563 | n27564 ;
  assign n27566 = n27562 | n27565 ;
  assign n27567 = n4784 | n27566 ;
  assign n27568 = ( ~n23712 & n27566 ) | ( ~n23712 & n27567 ) | ( n27566 & n27567 ) ;
  assign n27569 = ~x20 & n27568 ;
  assign n27570 = x20 | n27569 ;
  assign n27571 = ( ~n27568 & n27569 ) | ( ~n27568 & n27570 ) | ( n27569 & n27570 ) ;
  assign n27572 = n27412 | n27415 ;
  assign n27573 = n4484 & ~n20710 ;
  assign n27574 = n4479 & ~n20552 ;
  assign n27575 = n4481 & n20556 ;
  assign n27576 = n27574 | n27575 ;
  assign n27577 = n27573 | n27576 ;
  assign n27578 = n4487 | n27577 ;
  assign n27579 = ( ~n22641 & n27577 ) | ( ~n22641 & n27578 ) | ( n27577 & n27578 ) ;
  assign n27580 = ~x26 & n27579 ;
  assign n27581 = x26 | n27580 ;
  assign n27582 = ( ~n27579 & n27580 ) | ( ~n27579 & n27581 ) | ( n27580 & n27581 ) ;
  assign n27583 = n4048 & n20562 ;
  assign n27584 = n4043 & ~n20689 ;
  assign n27585 = n4045 & n20560 ;
  assign n27586 = n27584 | n27585 ;
  assign n27587 = n27583 | n27586 ;
  assign n27588 = n4051 | n27587 ;
  assign n27589 = ( ~n21044 & n27587 ) | ( ~n21044 & n27588 ) | ( n27587 & n27588 ) ;
  assign n27590 = ~x29 & n27589 ;
  assign n27591 = x29 | n27590 ;
  assign n27592 = ( ~n27589 & n27590 ) | ( ~n27589 & n27591 ) | ( n27590 & n27591 ) ;
  assign n27593 = n3744 & ~n20573 ;
  assign n27594 = n3639 & ~n20584 ;
  assign n27595 = n3727 & ~n20569 ;
  assign n27596 = n27594 | n27595 ;
  assign n27597 = n27593 | n27596 ;
  assign n27598 = n3636 | n27597 ;
  assign n27599 = ( ~n21860 & n27597 ) | ( ~n21860 & n27598 ) | ( n27597 & n27598 ) ;
  assign n27600 = n836 | n2967 ;
  assign n27601 = n2411 | n2891 ;
  assign n27602 = n27600 | n27601 ;
  assign n27603 = n19620 | n27602 ;
  assign n27604 = n1613 | n27603 ;
  assign n27605 = n1930 | n27604 ;
  assign n27606 = n1279 | n27605 ;
  assign n27607 = n2662 & ~n27606 ;
  assign n27608 = n944 | n2410 ;
  assign n27609 = n27607 & ~n27608 ;
  assign n27610 = n446 | n697 ;
  assign n27611 = n621 | n27610 ;
  assign n27612 = n212 | n27611 ;
  assign n27613 = n27609 & ~n27612 ;
  assign n27614 = ~n27223 & n27613 ;
  assign n27615 = n27223 & ~n27613 ;
  assign n27616 = n27614 | n27615 ;
  assign n27617 = n12703 & n26156 ;
  assign n27618 = ~x8 & n27617 ;
  assign n27619 = x8 | n27618 ;
  assign n27620 = ( ~n27617 & n27618 ) | ( ~n27617 & n27619 ) | ( n27618 & n27619 ) ;
  assign n27621 = n27616 | n27620 ;
  assign n27622 = n27616 & n27620 ;
  assign n27623 = n27621 & ~n27622 ;
  assign n27624 = n27391 & ~n27393 ;
  assign n27625 = ( n27599 & n27623 ) | ( n27599 & n27624 ) | ( n27623 & n27624 ) ;
  assign n27626 = ( n27623 & n27624 ) | ( n27623 & ~n27625 ) | ( n27624 & ~n27625 ) ;
  assign n27627 = ( n27599 & ~n27625 ) | ( n27599 & n27626 ) | ( ~n27625 & n27626 ) ;
  assign n27628 = n27592 & ~n27627 ;
  assign n27629 = ~n27592 & n27627 ;
  assign n27630 = n27628 | n27629 ;
  assign n27631 = n27404 | n27410 ;
  assign n27632 = n27630 & ~n27631 ;
  assign n27633 = ~n27630 & n27631 ;
  assign n27634 = n27632 | n27633 ;
  assign n27635 = n27582 & ~n27634 ;
  assign n27636 = n27634 | n27635 ;
  assign n27637 = ( ~n27582 & n27635 ) | ( ~n27582 & n27636 ) | ( n27635 & n27636 ) ;
  assign n27638 = ~n27572 & n27637 ;
  assign n27639 = n27572 & ~n27637 ;
  assign n27640 = n27638 | n27639 ;
  assign n27641 = n4551 & ~n20724 ;
  assign n27642 = n4546 & n20546 ;
  assign n27643 = n4548 & ~n20542 ;
  assign n27644 = n27642 | n27643 ;
  assign n27645 = n27641 | n27644 ;
  assign n27646 = n4554 | n27645 ;
  assign n27647 = ( n23229 & n27645 ) | ( n23229 & n27646 ) | ( n27645 & n27646 ) ;
  assign n27648 = x23 & n27647 ;
  assign n27649 = x23 & ~n27648 ;
  assign n27650 = ( n27647 & ~n27648 ) | ( n27647 & n27649 ) | ( ~n27648 & n27649 ) ;
  assign n27651 = ~n27640 & n27650 ;
  assign n27652 = n27640 | n27651 ;
  assign n27653 = n27640 & n27650 ;
  assign n27654 = n27433 | n27653 ;
  assign n27655 = n27652 & ~n27654 ;
  assign n27656 = ( n27433 & ~n27652 ) | ( n27433 & n27653 ) | ( ~n27652 & n27653 ) ;
  assign n27657 = n27655 | n27656 ;
  assign n27658 = n27571 & ~n27657 ;
  assign n27659 = n27657 | n27658 ;
  assign n27660 = ( ~n27571 & n27658 ) | ( ~n27571 & n27659 ) | ( n27658 & n27659 ) ;
  assign n27661 = ~n27450 & n27660 ;
  assign n27662 = n27450 & ~n27660 ;
  assign n27663 = n27661 | n27662 ;
  assign n27664 = ~n27467 & n27559 ;
  assign n27665 = n27663 & ~n27664 ;
  assign n27666 = ~n27561 & n27665 ;
  assign n27667 = ( n27561 & ~n27663 ) | ( n27561 & n27664 ) | ( ~n27663 & n27664 ) ;
  assign n27668 = n27666 | n27667 ;
  assign n27669 = n7280 & n25187 ;
  assign n27670 = n5384 & ~n24334 ;
  assign n27671 = n7277 & n24324 ;
  assign n27672 = n27670 | n27671 ;
  assign n27673 = n27669 | n27672 ;
  assign n27674 = n39 | n27673 ;
  assign n27675 = ( n25193 & n27673 ) | ( n25193 & n27674 ) | ( n27673 & n27674 ) ;
  assign n27676 = x14 & n27675 ;
  assign n27677 = x14 & ~n27676 ;
  assign n27678 = ( n27675 & ~n27676 ) | ( n27675 & n27677 ) | ( ~n27676 & n27677 ) ;
  assign n27679 = ~n27668 & n27678 ;
  assign n27680 = n27668 | n27679 ;
  assign n27681 = n27668 & n27678 ;
  assign n27682 = n27487 | n27681 ;
  assign n27683 = n27680 & ~n27682 ;
  assign n27684 = ( n27487 & ~n27680 ) | ( n27487 & n27681 ) | ( ~n27680 & n27681 ) ;
  assign n27685 = n27683 | n27684 ;
  assign n27686 = ~n27537 & n27547 ;
  assign n27687 = n27685 & ~n27686 ;
  assign n27688 = ~n27549 & n27687 ;
  assign n27689 = ( n27549 & ~n27685 ) | ( n27549 & n27686 ) | ( ~n27685 & n27686 ) ;
  assign n27690 = n27688 | n27689 ;
  assign n27691 = n27536 & ~n27690 ;
  assign n27692 = ~n27536 & n27690 ;
  assign n27693 = n27691 | n27692 ;
  assign n27694 = n27524 | n27528 ;
  assign n27695 = ~n27693 & n27694 ;
  assign n27696 = n27524 | n27526 ;
  assign n27697 = ~n27693 & n27696 ;
  assign n27698 = ( n27148 & n27695 ) | ( n27148 & n27697 ) | ( n27695 & n27697 ) ;
  assign n27699 = ( n27148 & n27694 ) | ( n27148 & n27696 ) | ( n27694 & n27696 ) ;
  assign n27700 = n27693 & ~n27699 ;
  assign n27701 = n27698 | n27700 ;
  assign n27702 = ~n27534 & n27701 ;
  assign n27703 = n27534 & ~n27701 ;
  assign n27704 = n27702 | n27703 ;
  assign n27705 = n27679 | n27684 ;
  assign n27706 = n27560 | n27667 ;
  assign n27707 = n27635 | n27639 ;
  assign n27708 = n4484 & n20546 ;
  assign n27709 = n4479 & n20556 ;
  assign n27710 = n4481 & ~n20710 ;
  assign n27711 = n27709 | n27710 ;
  assign n27712 = n27708 | n27711 ;
  assign n27713 = n4487 & ~n21031 ;
  assign n27714 = ( n4487 & n21037 ) | ( n4487 & n27713 ) | ( n21037 & n27713 ) ;
  assign n27715 = n27712 | n27714 ;
  assign n27716 = x26 | n27715 ;
  assign n27717 = ~x26 & n27716 ;
  assign n27718 = ( ~n27715 & n27716 ) | ( ~n27715 & n27717 ) | ( n27716 & n27717 ) ;
  assign n27719 = n3744 & ~n20689 ;
  assign n27720 = n3639 & ~n20569 ;
  assign n27721 = n3727 & ~n20573 ;
  assign n27722 = n27720 | n27721 ;
  assign n27723 = n27719 | n27722 ;
  assign n27724 = ( n3636 & ~n22192 ) | ( n3636 & n22193 ) | ( ~n22192 & n22193 ) ;
  assign n27725 = n27723 | n27724 ;
  assign n27726 = n428 | n2508 ;
  assign n27727 = n498 | n27726 ;
  assign n27728 = n383 | n27727 ;
  assign n27729 = n596 | n27728 ;
  assign n27730 = n444 | n27729 ;
  assign n27731 = n112 | n27730 ;
  assign n27732 = n661 | n27731 ;
  assign n27733 = n2802 | n2996 ;
  assign n27734 = n13889 | n27733 ;
  assign n27735 = n12867 | n27734 ;
  assign n27736 = n3873 | n3916 ;
  assign n27737 = n27735 | n27736 ;
  assign n27738 = ( n766 & n1673 ) | ( n766 & n27737 ) | ( n1673 & n27737 ) ;
  assign n27739 = n1673 & ~n27738 ;
  assign n27740 = ~n27732 & n27739 ;
  assign n27741 = ( n27615 & ~n27621 ) | ( n27615 & n27740 ) | ( ~n27621 & n27740 ) ;
  assign n27742 = ( n27614 & ~n27615 ) | ( n27614 & n27620 ) | ( ~n27615 & n27620 ) ;
  assign n27743 = ~n27740 & n27742 ;
  assign n27744 = n27741 | n27743 ;
  assign n27745 = n27725 | n27744 ;
  assign n27746 = ~n27744 & n27745 ;
  assign n27747 = ( ~n27725 & n27745 ) | ( ~n27725 & n27746 ) | ( n27745 & n27746 ) ;
  assign n27748 = ( n27599 & n27623 ) | ( n27599 & n27627 ) | ( n27623 & n27627 ) ;
  assign n27749 = n27747 & ~n27748 ;
  assign n27750 = ~n27747 & n27748 ;
  assign n27751 = n27749 | n27750 ;
  assign n27752 = n4048 & ~n20552 ;
  assign n27753 = n4043 & n20560 ;
  assign n27754 = n4045 & n20562 ;
  assign n27755 = n27753 | n27754 ;
  assign n27756 = n27752 | n27755 ;
  assign n27757 = n4051 & n22510 ;
  assign n27758 = ~n22512 & n27757 ;
  assign n27759 = ( n4051 & n27756 ) | ( n4051 & ~n27758 ) | ( n27756 & ~n27758 ) ;
  assign n27760 = x29 & n27759 ;
  assign n27761 = x29 & ~n27760 ;
  assign n27762 = ( n27759 & ~n27760 ) | ( n27759 & n27761 ) | ( ~n27760 & n27761 ) ;
  assign n27763 = ~n27751 & n27762 ;
  assign n27764 = n27751 & ~n27762 ;
  assign n27765 = n27763 | n27764 ;
  assign n27766 = n27628 | n27633 ;
  assign n27767 = ( n27718 & n27765 ) | ( n27718 & ~n27766 ) | ( n27765 & ~n27766 ) ;
  assign n27768 = ( ~n27765 & n27766 ) | ( ~n27765 & n27767 ) | ( n27766 & n27767 ) ;
  assign n27769 = ( ~n27718 & n27767 ) | ( ~n27718 & n27768 ) | ( n27767 & n27768 ) ;
  assign n27770 = ~n27707 & n27769 ;
  assign n27771 = n27707 & ~n27769 ;
  assign n27772 = n27770 | n27771 ;
  assign n27773 = n4551 & ~n20536 ;
  assign n27774 = n4546 & ~n20542 ;
  assign n27775 = n4548 & ~n20724 ;
  assign n27776 = n27774 | n27775 ;
  assign n27777 = n27773 | n27776 ;
  assign n27778 = ( n4554 & n23213 ) | ( n4554 & ~n23217 ) | ( n23213 & ~n23217 ) ;
  assign n27779 = n27777 | n27778 ;
  assign n27780 = x23 | n27779 ;
  assign n27781 = ~x23 & n27780 ;
  assign n27782 = ( ~n27779 & n27780 ) | ( ~n27779 & n27781 ) | ( n27780 & n27781 ) ;
  assign n27783 = n27772 & n27782 ;
  assign n27784 = ( n27707 & ~n27769 ) | ( n27707 & n27782 ) | ( ~n27769 & n27782 ) ;
  assign n27785 = n27770 | n27784 ;
  assign n27786 = ~n27783 & n27785 ;
  assign n27787 = n27651 | n27656 ;
  assign n27788 = n27786 & ~n27787 ;
  assign n27789 = ~n27786 & n27787 ;
  assign n27790 = n27788 | n27789 ;
  assign n27791 = n4781 & n20921 ;
  assign n27792 = n4776 & n20532 ;
  assign n27793 = n4778 & n20838 ;
  assign n27794 = n27792 | n27793 ;
  assign n27795 = n27791 | n27794 ;
  assign n27796 = ( n4784 & n23691 ) | ( n4784 & n23695 ) | ( n23691 & n23695 ) ;
  assign n27797 = n27795 | n27796 ;
  assign n27798 = x20 | n27797 ;
  assign n27799 = ~x20 & n27798 ;
  assign n27800 = ( ~n27797 & n27798 ) | ( ~n27797 & n27799 ) | ( n27798 & n27799 ) ;
  assign n27801 = n27790 & n27800 ;
  assign n27802 = ( ~n27786 & n27787 ) | ( ~n27786 & n27800 ) | ( n27787 & n27800 ) ;
  assign n27803 = n27788 | n27802 ;
  assign n27804 = ~n27801 & n27803 ;
  assign n27805 = n27658 | n27662 ;
  assign n27806 = n27804 & ~n27805 ;
  assign n27807 = ~n27804 & n27805 ;
  assign n27808 = n27806 | n27807 ;
  assign n27809 = n5083 & ~n24334 ;
  assign n27810 = n5069 & ~n21005 ;
  assign n27811 = n5070 & n24329 ;
  assign n27812 = n27810 | n27811 ;
  assign n27813 = n27809 | n27812 ;
  assign n27814 = ( n5074 & ~n24373 ) | ( n5074 & n24376 ) | ( ~n24373 & n24376 ) ;
  assign n27815 = n27813 | n27814 ;
  assign n27816 = x17 | n27815 ;
  assign n27817 = ~x17 & n27816 ;
  assign n27818 = ( ~n27815 & n27816 ) | ( ~n27815 & n27817 ) | ( n27816 & n27817 ) ;
  assign n27819 = n27808 & n27818 ;
  assign n27820 = ( ~n27804 & n27805 ) | ( ~n27804 & n27818 ) | ( n27805 & n27818 ) ;
  assign n27821 = n27806 | n27820 ;
  assign n27822 = ~n27819 & n27821 ;
  assign n27823 = n27706 & ~n27822 ;
  assign n27824 = n27706 & ~n27823 ;
  assign n27825 = n27706 | n27822 ;
  assign n27826 = ~n27824 & n27825 ;
  assign n27827 = n7280 & n25442 ;
  assign n27828 = n5384 & n24324 ;
  assign n27829 = n7277 & n25187 ;
  assign n27830 = n27828 | n27829 ;
  assign n27831 = n27827 | n27830 ;
  assign n27832 = n39 | n27831 ;
  assign n27833 = ( n25452 & n27831 ) | ( n25452 & n27832 ) | ( n27831 & n27832 ) ;
  assign n27834 = x14 & n27833 ;
  assign n27835 = x14 & ~n27834 ;
  assign n27836 = ( n27833 & ~n27834 ) | ( n27833 & n27835 ) | ( ~n27834 & n27835 ) ;
  assign n27837 = ~n27826 & n27836 ;
  assign n27838 = n27826 & ~n27836 ;
  assign n27839 = n27837 | n27838 ;
  assign n27840 = ~n27705 & n27839 ;
  assign n27841 = n27705 & ~n27839 ;
  assign n27842 = n27840 | n27841 ;
  assign n27843 = n7305 & n26156 ;
  assign n27844 = n7300 & ~n25676 ;
  assign n27845 = n7302 & n25928 ;
  assign n27846 = n27844 | n27845 ;
  assign n27847 = n27843 | n27846 ;
  assign n27848 = n7308 | n27847 ;
  assign n27849 = ( n26167 & n27847 ) | ( n26167 & n27848 ) | ( n27847 & n27848 ) ;
  assign n27850 = x11 & n27849 ;
  assign n27851 = x11 & ~n27850 ;
  assign n27852 = ( n27849 & ~n27850 ) | ( n27849 & n27851 ) | ( ~n27850 & n27851 ) ;
  assign n27853 = n27842 & n27852 ;
  assign n27854 = ( n27705 & ~n27839 ) | ( n27705 & n27852 ) | ( ~n27839 & n27852 ) ;
  assign n27855 = n27840 | n27854 ;
  assign n27856 = ~n27853 & n27855 ;
  assign n27857 = n27548 | n27689 ;
  assign n27858 = ~n27856 & n27857 ;
  assign n27859 = n27856 | n27858 ;
  assign n27860 = n27856 & n27857 ;
  assign n27861 = n27859 & ~n27860 ;
  assign n27862 = n27691 | n27695 ;
  assign n27863 = ~n27861 & n27862 ;
  assign n27864 = n27691 | n27697 ;
  assign n27865 = ~n27861 & n27864 ;
  assign n27866 = ( n27148 & n27863 ) | ( n27148 & n27865 ) | ( n27863 & n27865 ) ;
  assign n27867 = ( n27148 & n27862 ) | ( n27148 & n27864 ) | ( n27862 & n27864 ) ;
  assign n27868 = n27861 & ~n27867 ;
  assign n27869 = n27866 | n27868 ;
  assign n27870 = n27703 & n27869 ;
  assign n27871 = n27703 | n27869 ;
  assign n27872 = ~n27870 & n27871 ;
  assign n27873 = n12878 & n26156 ;
  assign n27874 = n7300 & n25928 ;
  assign n27875 = n27873 | n27874 ;
  assign n27876 = n7308 | n27875 ;
  assign n27877 = ( n26165 & n27875 ) | ( n26165 & n27876 ) | ( n27875 & n27876 ) ;
  assign n27878 = x11 & n27877 ;
  assign n27879 = x11 & ~n27878 ;
  assign n27880 = ( n27877 & ~n27878 ) | ( n27877 & n27879 ) | ( ~n27878 & n27879 ) ;
  assign n27881 = n27823 | n27880 ;
  assign n27882 = n27837 | n27881 ;
  assign n27883 = ( n27823 & n27837 ) | ( n27823 & n27880 ) | ( n27837 & n27880 ) ;
  assign n27884 = n27882 & ~n27883 ;
  assign n27885 = n7280 & ~n25676 ;
  assign n27886 = n5384 & n25187 ;
  assign n27887 = n7277 & n25442 ;
  assign n27888 = n27886 | n27887 ;
  assign n27889 = n27885 | n27888 ;
  assign n27890 = n39 & ~n25690 ;
  assign n27891 = ( n39 & n25694 ) | ( n39 & n27890 ) | ( n25694 & n27890 ) ;
  assign n27892 = n27889 | n27891 ;
  assign n27893 = x14 | n27892 ;
  assign n27894 = ~x14 & n27893 ;
  assign n27895 = ( ~n27892 & n27893 ) | ( ~n27892 & n27894 ) | ( n27893 & n27894 ) ;
  assign n27896 = n5083 & n24324 ;
  assign n27897 = n5069 & n24329 ;
  assign n27898 = n5070 & ~n24334 ;
  assign n27899 = n27897 | n27898 ;
  assign n27900 = n27896 | n27899 ;
  assign n27901 = n5074 & ~n24353 ;
  assign n27902 = ( n5074 & n24356 ) | ( n5074 & n27901 ) | ( n24356 & n27901 ) ;
  assign n27903 = n27900 | n27902 ;
  assign n27904 = x17 | n27903 ;
  assign n27905 = ~x17 & n27904 ;
  assign n27906 = ( ~n27903 & n27904 ) | ( ~n27903 & n27905 ) | ( n27904 & n27905 ) ;
  assign n27907 = n4781 & ~n21005 ;
  assign n27908 = n4776 & n20838 ;
  assign n27909 = n4778 & n20921 ;
  assign n27910 = n27908 | n27909 ;
  assign n27911 = n27907 | n27910 ;
  assign n27912 = n4784 | n27911 ;
  assign n27913 = ( ~n21015 & n27911 ) | ( ~n21015 & n27912 ) | ( n27911 & n27912 ) ;
  assign n27914 = ~x20 & n27913 ;
  assign n27915 = x20 | n27914 ;
  assign n27916 = ( ~n27913 & n27914 ) | ( ~n27913 & n27915 ) | ( n27914 & n27915 ) ;
  assign n27917 = n4551 & n20532 ;
  assign n27918 = n4546 & ~n20724 ;
  assign n27919 = n4548 & ~n20536 ;
  assign n27920 = n27918 | n27919 ;
  assign n27921 = n27917 | n27920 ;
  assign n27922 = n4554 | n27921 ;
  assign n27923 = ( n23203 & n27921 ) | ( n23203 & n27922 ) | ( n27921 & n27922 ) ;
  assign n27924 = x23 & n27923 ;
  assign n27925 = x23 & ~n27924 ;
  assign n27926 = ( n27923 & ~n27924 ) | ( n27923 & n27925 ) | ( ~n27924 & n27925 ) ;
  assign n27927 = n27750 | n27763 ;
  assign n27950 = ( n27725 & n27740 ) | ( n27725 & n27747 ) | ( n27740 & n27747 ) ;
  assign n27928 = n27200 | n27207 ;
  assign n27929 = n808 | n869 ;
  assign n27930 = n731 | n27929 ;
  assign n27931 = n27928 | n27930 ;
  assign n27932 = n752 | n2610 ;
  assign n27933 = n2684 | n27932 ;
  assign n27934 = n1271 | n1756 ;
  assign n27935 = n27933 | n27934 ;
  assign n27936 = n13223 | n27935 ;
  assign n27937 = ( ~n4417 & n19645 ) | ( ~n4417 & n27936 ) | ( n19645 & n27936 ) ;
  assign n27938 = n4417 | n27937 ;
  assign n27939 = n27931 | n27938 ;
  assign n27940 = n1115 | n1442 ;
  assign n27941 = n522 | n27940 ;
  assign n27942 = n326 | n27941 ;
  assign n27943 = n356 | n27942 ;
  assign n27944 = n602 | n27943 ;
  assign n27945 = n102 | n27944 ;
  assign n27946 = n27939 | n27945 ;
  assign n27947 = n27740 | n27946 ;
  assign n27948 = n27740 & n27946 ;
  assign n27949 = n27947 & ~n27948 ;
  assign n27951 = n27949 & n27950 ;
  assign n27952 = n27950 & ~n27951 ;
  assign n27953 = n27948 | n27951 ;
  assign n27954 = n27947 & ~n27953 ;
  assign n27955 = n27952 | n27954 ;
  assign n27956 = n3744 & n20560 ;
  assign n27957 = n3639 & ~n20573 ;
  assign n27958 = n3727 & ~n20689 ;
  assign n27959 = n27957 | n27958 ;
  assign n27960 = n27956 | n27959 ;
  assign n27961 = ( n3636 & n22173 ) | ( n3636 & n22176 ) | ( n22173 & n22176 ) ;
  assign n27962 = n27960 | n27961 ;
  assign n27963 = n27955 & n27962 ;
  assign n27964 = n27955 & ~n27963 ;
  assign n27965 = ~n27955 & n27962 ;
  assign n27966 = n4048 & n20556 ;
  assign n27967 = n4043 & n20562 ;
  assign n27968 = n4045 & ~n20552 ;
  assign n27969 = n27967 | n27968 ;
  assign n27970 = n27966 | n27969 ;
  assign n27971 = n4051 | n27970 ;
  assign n27972 = ( ~n22655 & n27970 ) | ( ~n22655 & n27971 ) | ( n27970 & n27971 ) ;
  assign n27973 = ~x29 & n27972 ;
  assign n27974 = x29 | n27973 ;
  assign n27975 = ( ~n27972 & n27973 ) | ( ~n27972 & n27974 ) | ( n27973 & n27974 ) ;
  assign n27976 = n27965 | n27975 ;
  assign n27977 = n27964 | n27976 ;
  assign n27978 = ( n27964 & n27965 ) | ( n27964 & n27975 ) | ( n27965 & n27975 ) ;
  assign n27979 = n27977 & ~n27978 ;
  assign n27980 = n4484 & ~n20542 ;
  assign n27981 = n4479 & ~n20710 ;
  assign n27982 = n4481 & n20546 ;
  assign n27983 = n27981 | n27982 ;
  assign n27984 = n27980 | n27983 ;
  assign n27985 = n4487 | n27984 ;
  assign n27986 = ( ~n23042 & n27984 ) | ( ~n23042 & n27985 ) | ( n27984 & n27985 ) ;
  assign n27987 = ~x26 & n27986 ;
  assign n27988 = x26 | n27987 ;
  assign n27989 = ( ~n27986 & n27987 ) | ( ~n27986 & n27988 ) | ( n27987 & n27988 ) ;
  assign n27990 = ( n27927 & n27979 ) | ( n27927 & n27989 ) | ( n27979 & n27989 ) ;
  assign n27991 = ( n27979 & n27989 ) | ( n27979 & ~n27990 ) | ( n27989 & ~n27990 ) ;
  assign n27992 = ( n27927 & ~n27990 ) | ( n27927 & n27991 ) | ( ~n27990 & n27991 ) ;
  assign n27993 = ( ~n27768 & n27926 ) | ( ~n27768 & n27992 ) | ( n27926 & n27992 ) ;
  assign n27994 = ( n27768 & ~n27992 ) | ( n27768 & n27993 ) | ( ~n27992 & n27993 ) ;
  assign n27995 = ( ~n27926 & n27993 ) | ( ~n27926 & n27994 ) | ( n27993 & n27994 ) ;
  assign n27996 = ( n27784 & n27916 ) | ( n27784 & ~n27995 ) | ( n27916 & ~n27995 ) ;
  assign n27997 = ( ~n27784 & n27995 ) | ( ~n27784 & n27996 ) | ( n27995 & n27996 ) ;
  assign n27998 = ( ~n27916 & n27996 ) | ( ~n27916 & n27997 ) | ( n27996 & n27997 ) ;
  assign n27999 = ( n27802 & n27906 ) | ( n27802 & ~n27998 ) | ( n27906 & ~n27998 ) ;
  assign n28000 = ( ~n27802 & n27998 ) | ( ~n27802 & n27999 ) | ( n27998 & n27999 ) ;
  assign n28001 = ( ~n27906 & n27999 ) | ( ~n27906 & n28000 ) | ( n27999 & n28000 ) ;
  assign n28002 = ( n27820 & n27895 ) | ( n27820 & ~n28001 ) | ( n27895 & ~n28001 ) ;
  assign n28003 = ( ~n27820 & n28001 ) | ( ~n27820 & n28002 ) | ( n28001 & n28002 ) ;
  assign n28004 = ( ~n27895 & n28002 ) | ( ~n27895 & n28003 ) | ( n28002 & n28003 ) ;
  assign n28005 = n27884 & ~n28004 ;
  assign n28006 = n28004 | n28005 ;
  assign n28007 = ( ~n27884 & n28005 ) | ( ~n27884 & n28006 ) | ( n28005 & n28006 ) ;
  assign n28008 = n27854 | n28007 ;
  assign n28009 = n27854 & n28007 ;
  assign n28010 = n28008 & ~n28009 ;
  assign n28011 = n27858 | n27863 ;
  assign n28012 = n28010 & n28011 ;
  assign n28013 = n27858 | n27865 ;
  assign n28014 = n28010 & n28013 ;
  assign n28015 = ( n27148 & n28012 ) | ( n27148 & n28014 ) | ( n28012 & n28014 ) ;
  assign n28016 = ( n27148 & n28011 ) | ( n27148 & n28013 ) | ( n28011 & n28013 ) ;
  assign n28017 = n28010 | n28016 ;
  assign n28018 = ~n28015 & n28017 ;
  assign n28019 = ( ~n27869 & n27871 ) | ( ~n27869 & n28018 ) | ( n27871 & n28018 ) ;
  assign n28020 = ( n27703 & n27869 ) | ( n27703 & ~n28018 ) | ( n27869 & ~n28018 ) ;
  assign n28021 = n27703 & ~n28020 ;
  assign n28022 = n28019 & ~n28021 ;
  assign n28023 = ( n27820 & n27895 ) | ( n27820 & n28001 ) | ( n27895 & n28001 ) ;
  assign n28024 = n7280 & n25928 ;
  assign n28025 = n5384 & n25442 ;
  assign n28026 = n7277 & ~n25676 ;
  assign n28027 = n28025 | n28026 ;
  assign n28028 = n28024 | n28027 ;
  assign n28029 = n39 | n28028 ;
  assign n28030 = ( ~n25936 & n28028 ) | ( ~n25936 & n28029 ) | ( n28028 & n28029 ) ;
  assign n28031 = ~x14 & n28030 ;
  assign n28032 = x14 | n28031 ;
  assign n28033 = ( ~n28030 & n28031 ) | ( ~n28030 & n28032 ) | ( n28031 & n28032 ) ;
  assign n28034 = n28023 & n28033 ;
  assign n28035 = n28023 & ~n28034 ;
  assign n28036 = ( n27784 & n27916 ) | ( n27784 & n27995 ) | ( n27916 & n27995 ) ;
  assign n28037 = n4781 & n24329 ;
  assign n28038 = n4776 & n20921 ;
  assign n28039 = n4778 & ~n21005 ;
  assign n28040 = n28038 | n28039 ;
  assign n28041 = n28037 | n28040 ;
  assign n28042 = ( n4784 & ~n24391 ) | ( n4784 & n24392 ) | ( ~n24391 & n24392 ) ;
  assign n28043 = n28041 | n28042 ;
  assign n28044 = x20 | n28043 ;
  assign n28045 = ~x20 & n28044 ;
  assign n28046 = ( ~n28043 & n28044 ) | ( ~n28043 & n28045 ) | ( n28044 & n28045 ) ;
  assign n28047 = n28036 & n28046 ;
  assign n28048 = n28036 & ~n28047 ;
  assign n28049 = n27963 | n27978 ;
  assign n28050 = n3744 & n20562 ;
  assign n28051 = n3639 & ~n20689 ;
  assign n28052 = n3727 & n20560 ;
  assign n28053 = n28051 | n28052 ;
  assign n28054 = n28050 | n28053 ;
  assign n28055 = n3636 | n28054 ;
  assign n28056 = ( ~n21044 & n28054 ) | ( ~n21044 & n28055 ) | ( n28054 & n28055 ) ;
  assign n28057 = n1188 | n4070 ;
  assign n28058 = n1974 | n28057 ;
  assign n28059 = n2689 | n28058 ;
  assign n28060 = n4094 | n28059 ;
  assign n28061 = n2919 & ~n28060 ;
  assign n28062 = n814 | n816 ;
  assign n28063 = n28061 & ~n28062 ;
  assign n28064 = n1963 | n2221 ;
  assign n28065 = n861 | n28064 ;
  assign n28066 = n1417 | n28065 ;
  assign n28067 = n3375 | n28066 ;
  assign n28068 = n28063 & ~n28067 ;
  assign n28069 = n428 | n648 ;
  assign n28070 = n327 | n28069 ;
  assign n28071 = n99 | n28070 ;
  assign n28072 = n207 | n28071 ;
  assign n28073 = n28068 & ~n28072 ;
  assign n28074 = n27740 & n28073 ;
  assign n28075 = n27740 | n28073 ;
  assign n28076 = ~n28074 & n28075 ;
  assign n28077 = n12880 & n26156 ;
  assign n28078 = ~x11 & n28077 ;
  assign n28079 = x11 | n28078 ;
  assign n28080 = ( ~n28077 & n28078 ) | ( ~n28077 & n28079 ) | ( n28078 & n28079 ) ;
  assign n28081 = n28076 & ~n28080 ;
  assign n28082 = ~n28076 & n28080 ;
  assign n28083 = n28081 | n28082 ;
  assign n28084 = n28056 & ~n28083 ;
  assign n28085 = n28056 & ~n28084 ;
  assign n28086 = n28056 | n28083 ;
  assign n28087 = ~n28085 & n28086 ;
  assign n28088 = n27953 & ~n28087 ;
  assign n28089 = n28087 | n28088 ;
  assign n28090 = n27953 & ~n28088 ;
  assign n28091 = n28089 & ~n28090 ;
  assign n28092 = n28049 & ~n28091 ;
  assign n28093 = ~n28049 & n28091 ;
  assign n28094 = n28092 | n28093 ;
  assign n28095 = n4048 & ~n20710 ;
  assign n28096 = n4043 & ~n20552 ;
  assign n28097 = n4045 & n20556 ;
  assign n28098 = n28096 | n28097 ;
  assign n28099 = n28095 | n28098 ;
  assign n28100 = n4051 | n28099 ;
  assign n28101 = ( ~n22641 & n28099 ) | ( ~n22641 & n28100 ) | ( n28099 & n28100 ) ;
  assign n28102 = ~x29 & n28101 ;
  assign n28103 = x29 | n28102 ;
  assign n28104 = ( ~n28101 & n28102 ) | ( ~n28101 & n28103 ) | ( n28102 & n28103 ) ;
  assign n28105 = n28094 & n28104 ;
  assign n28106 = n28094 | n28104 ;
  assign n28107 = ~n28105 & n28106 ;
  assign n28108 = n4484 & ~n20724 ;
  assign n28109 = n4479 & n20546 ;
  assign n28110 = n4481 & ~n20542 ;
  assign n28111 = n28109 | n28110 ;
  assign n28112 = n28108 | n28111 ;
  assign n28113 = n4487 | n28112 ;
  assign n28114 = ( n23229 & n28112 ) | ( n23229 & n28113 ) | ( n28112 & n28113 ) ;
  assign n28115 = x26 & n28114 ;
  assign n28116 = x26 & ~n28115 ;
  assign n28117 = ( n28114 & ~n28115 ) | ( n28114 & n28116 ) | ( ~n28115 & n28116 ) ;
  assign n28118 = ~n28107 & n28117 ;
  assign n28119 = n28107 & ~n28117 ;
  assign n28120 = n28118 | n28119 ;
  assign n28121 = ~n27990 & n28120 ;
  assign n28122 = n27990 & ~n28120 ;
  assign n28123 = n28121 | n28122 ;
  assign n28124 = n4551 & n20838 ;
  assign n28125 = n4546 & ~n20536 ;
  assign n28126 = n4548 & n20532 ;
  assign n28127 = n28125 | n28126 ;
  assign n28128 = n28124 | n28127 ;
  assign n28129 = n4554 | n28128 ;
  assign n28130 = ( ~n23712 & n28128 ) | ( ~n23712 & n28129 ) | ( n28128 & n28129 ) ;
  assign n28131 = ~x23 & n28130 ;
  assign n28132 = x23 | n28131 ;
  assign n28133 = ( ~n28130 & n28131 ) | ( ~n28130 & n28132 ) | ( n28131 & n28132 ) ;
  assign n28134 = ~n28123 & n28133 ;
  assign n28135 = n28123 | n28134 ;
  assign n28136 = ( n27768 & n27926 ) | ( n27768 & n27992 ) | ( n27926 & n27992 ) ;
  assign n28137 = n28123 & n28133 ;
  assign n28138 = n28136 | n28137 ;
  assign n28139 = n28135 & ~n28138 ;
  assign n28140 = ( ~n28135 & n28136 ) | ( ~n28135 & n28137 ) | ( n28136 & n28137 ) ;
  assign n28141 = n28139 | n28140 ;
  assign n28142 = ~n28036 & n28046 ;
  assign n28143 = n28141 & ~n28142 ;
  assign n28144 = ~n28048 & n28143 ;
  assign n28145 = ( n28048 & ~n28141 ) | ( n28048 & n28142 ) | ( ~n28141 & n28142 ) ;
  assign n28146 = n28144 | n28145 ;
  assign n28147 = n5083 & n25187 ;
  assign n28148 = n5069 & ~n24334 ;
  assign n28149 = n5070 & n24324 ;
  assign n28150 = n28148 | n28149 ;
  assign n28151 = n28147 | n28150 ;
  assign n28152 = n5074 | n28151 ;
  assign n28153 = ( n25193 & n28151 ) | ( n25193 & n28152 ) | ( n28151 & n28152 ) ;
  assign n28154 = x17 & n28153 ;
  assign n28155 = x17 & ~n28154 ;
  assign n28156 = ( n28153 & ~n28154 ) | ( n28153 & n28155 ) | ( ~n28154 & n28155 ) ;
  assign n28157 = ~n28146 & n28156 ;
  assign n28158 = n28146 | n28157 ;
  assign n28159 = ( n27802 & n27906 ) | ( n27802 & n27998 ) | ( n27906 & n27998 ) ;
  assign n28160 = n28146 & n28156 ;
  assign n28161 = n28159 | n28160 ;
  assign n28162 = n28158 & ~n28161 ;
  assign n28163 = ( ~n28158 & n28159 ) | ( ~n28158 & n28160 ) | ( n28159 & n28160 ) ;
  assign n28164 = n28162 | n28163 ;
  assign n28165 = ~n28023 & n28033 ;
  assign n28166 = n28164 & ~n28165 ;
  assign n28167 = ~n28035 & n28166 ;
  assign n28168 = ( n28035 & ~n28164 ) | ( n28035 & n28165 ) | ( ~n28164 & n28165 ) ;
  assign n28169 = n28167 | n28168 ;
  assign n28170 = ( n27882 & n27883 ) | ( n27882 & n28004 ) | ( n27883 & n28004 ) ;
  assign n28171 = ~n28169 & n28170 ;
  assign n28172 = n28169 & ~n28170 ;
  assign n28173 = n28171 | n28172 ;
  assign n28174 = n28009 | n28012 ;
  assign n28175 = ~n28173 & n28174 ;
  assign n28176 = n28009 | n28014 ;
  assign n28177 = ~n28173 & n28176 ;
  assign n28178 = ( n27148 & n28175 ) | ( n27148 & n28177 ) | ( n28175 & n28177 ) ;
  assign n28179 = ( n27148 & n28174 ) | ( n27148 & n28176 ) | ( n28174 & n28176 ) ;
  assign n28180 = n28173 & ~n28179 ;
  assign n28181 = n28178 | n28180 ;
  assign n28182 = ~n28021 & n28181 ;
  assign n28183 = n28021 & ~n28181 ;
  assign n28184 = n28182 | n28183 ;
  assign n28185 = n7280 & n26156 ;
  assign n28186 = n5384 & ~n25676 ;
  assign n28187 = n7277 & n25928 ;
  assign n28188 = n28186 | n28187 ;
  assign n28189 = n28185 | n28188 ;
  assign n28190 = n39 | n28189 ;
  assign n28191 = ( n26167 & n28189 ) | ( n26167 & n28190 ) | ( n28189 & n28190 ) ;
  assign n28192 = x14 & n28191 ;
  assign n28193 = x14 & ~n28192 ;
  assign n28194 = ( n28191 & ~n28192 ) | ( n28191 & n28193 ) | ( ~n28192 & n28193 ) ;
  assign n28195 = n28157 | n28163 ;
  assign n28196 = n4781 & ~n24334 ;
  assign n28197 = n4776 & ~n21005 ;
  assign n28198 = n4778 & n24329 ;
  assign n28199 = n28197 | n28198 ;
  assign n28200 = n28196 | n28199 ;
  assign n28201 = ( n4784 & ~n24373 ) | ( n4784 & n24376 ) | ( ~n24373 & n24376 ) ;
  assign n28202 = n28200 | n28201 ;
  assign n28203 = x20 | n28202 ;
  assign n28204 = ~x20 & n28203 ;
  assign n28205 = ( ~n28202 & n28203 ) | ( ~n28202 & n28204 ) | ( n28203 & n28204 ) ;
  assign n28206 = n28134 | n28140 ;
  assign n28207 = n4551 & n20921 ;
  assign n28208 = n4546 & n20532 ;
  assign n28209 = n4548 & n20838 ;
  assign n28210 = n28208 | n28209 ;
  assign n28211 = n28207 | n28210 ;
  assign n28212 = ( n4554 & n23691 ) | ( n4554 & n23695 ) | ( n23691 & n23695 ) ;
  assign n28213 = n28211 | n28212 ;
  assign n28214 = x23 | n28213 ;
  assign n28215 = ~x23 & n28214 ;
  assign n28216 = ( ~n28213 & n28214 ) | ( ~n28213 & n28215 ) | ( n28214 & n28215 ) ;
  assign n28217 = n28118 | n28122 ;
  assign n28218 = ( n28092 & ~n28094 ) | ( n28092 & n28106 ) | ( ~n28094 & n28106 ) ;
  assign n28219 = n28084 | n28088 ;
  assign n28220 = n3744 & ~n20552 ;
  assign n28221 = n3639 & n20560 ;
  assign n28222 = n3727 & n20562 ;
  assign n28223 = n28221 | n28222 ;
  assign n28224 = n28220 | n28223 ;
  assign n28225 = n3636 & ~n22510 ;
  assign n28226 = ( n3636 & n22512 ) | ( n3636 & n28225 ) | ( n22512 & n28225 ) ;
  assign n28227 = n28224 | n28226 ;
  assign n28228 = n1052 | n2060 ;
  assign n28229 = n2991 | n28228 ;
  assign n28230 = n474 | n28229 ;
  assign n28231 = n19923 | n28230 ;
  assign n28232 = n25802 | n28231 ;
  assign n28233 = n640 | n28232 ;
  assign n28234 = n20011 | n28233 ;
  assign n28235 = n13225 | n13228 ;
  assign n28236 = n26251 | n28235 ;
  assign n28237 = n28234 | n28236 ;
  assign n28238 = n1022 | n2341 ;
  assign n28239 = n478 | n28238 ;
  assign n28240 = n528 | n28239 ;
  assign n28241 = n520 | n28240 ;
  assign n28242 = ( ~n729 & n28237 ) | ( ~n729 & n28241 ) | ( n28237 & n28241 ) ;
  assign n28243 = n729 | n28242 ;
  assign n28244 = ( n28075 & ~n28081 ) | ( n28075 & n28243 ) | ( ~n28081 & n28243 ) ;
  assign n28245 = ( n28074 & n28075 ) | ( n28074 & n28080 ) | ( n28075 & n28080 ) ;
  assign n28246 = n28243 & n28245 ;
  assign n28247 = n28244 & ~n28246 ;
  assign n28248 = n28227 | n28247 ;
  assign n28249 = ~n28247 & n28248 ;
  assign n28250 = ( ~n28227 & n28248 ) | ( ~n28227 & n28249 ) | ( n28248 & n28249 ) ;
  assign n28251 = n28219 | n28250 ;
  assign n28252 = n28219 & n28250 ;
  assign n28253 = n28251 & ~n28252 ;
  assign n28254 = n4048 & n20546 ;
  assign n28255 = n4043 & n20556 ;
  assign n28256 = n4045 & ~n20710 ;
  assign n28257 = n28255 | n28256 ;
  assign n28258 = n28254 | n28257 ;
  assign n28259 = n4051 & n21031 ;
  assign n28260 = ~n21037 & n28259 ;
  assign n28261 = ( n4051 & n28258 ) | ( n4051 & ~n28260 ) | ( n28258 & ~n28260 ) ;
  assign n28262 = x29 & n28261 ;
  assign n28263 = x29 & ~n28262 ;
  assign n28264 = ( n28261 & ~n28262 ) | ( n28261 & n28263 ) | ( ~n28262 & n28263 ) ;
  assign n28265 = n28253 & n28264 ;
  assign n28266 = n28253 | n28264 ;
  assign n28267 = ~n28265 & n28266 ;
  assign n28268 = n4484 & ~n20536 ;
  assign n28269 = n4479 & ~n20542 ;
  assign n28270 = n4481 & ~n20724 ;
  assign n28271 = n28269 | n28270 ;
  assign n28272 = n28268 | n28271 ;
  assign n28273 = ( n4487 & n23213 ) | ( n4487 & ~n23217 ) | ( n23213 & ~n23217 ) ;
  assign n28274 = n28272 | n28273 ;
  assign n28275 = x26 | n28274 ;
  assign n28276 = ~x26 & n28275 ;
  assign n28277 = ( ~n28274 & n28275 ) | ( ~n28274 & n28276 ) | ( n28275 & n28276 ) ;
  assign n28278 = ( n28218 & n28267 ) | ( n28218 & n28277 ) | ( n28267 & n28277 ) ;
  assign n28279 = ( n28267 & n28277 ) | ( n28267 & ~n28278 ) | ( n28277 & ~n28278 ) ;
  assign n28280 = ( n28218 & ~n28278 ) | ( n28218 & n28279 ) | ( ~n28278 & n28279 ) ;
  assign n28281 = ( n28216 & ~n28217 ) | ( n28216 & n28280 ) | ( ~n28217 & n28280 ) ;
  assign n28282 = ( n28217 & ~n28280 ) | ( n28217 & n28281 ) | ( ~n28280 & n28281 ) ;
  assign n28283 = ( ~n28216 & n28281 ) | ( ~n28216 & n28282 ) | ( n28281 & n28282 ) ;
  assign n28284 = ( n28205 & ~n28206 ) | ( n28205 & n28283 ) | ( ~n28206 & n28283 ) ;
  assign n28285 = ( n28206 & ~n28283 ) | ( n28206 & n28284 ) | ( ~n28283 & n28284 ) ;
  assign n28286 = ( ~n28205 & n28284 ) | ( ~n28205 & n28285 ) | ( n28284 & n28285 ) ;
  assign n28287 = n28047 | n28145 ;
  assign n28288 = n28286 & n28287 ;
  assign n28289 = n28286 & ~n28288 ;
  assign n28290 = ~n28286 & n28287 ;
  assign n28291 = n28289 | n28290 ;
  assign n28292 = n5083 & n25442 ;
  assign n28293 = n5069 & n24324 ;
  assign n28294 = n5070 & n25187 ;
  assign n28295 = n28293 | n28294 ;
  assign n28296 = n28292 | n28295 ;
  assign n28297 = n5074 | n28296 ;
  assign n28298 = ( n25452 & n28296 ) | ( n25452 & n28297 ) | ( n28296 & n28297 ) ;
  assign n28299 = x17 & n28298 ;
  assign n28300 = x17 & ~n28299 ;
  assign n28301 = ( n28298 & ~n28299 ) | ( n28298 & n28300 ) | ( ~n28299 & n28300 ) ;
  assign n28302 = n28291 & n28301 ;
  assign n28303 = n28291 | n28301 ;
  assign n28304 = ~n28302 & n28303 ;
  assign n28305 = ( n28194 & n28195 ) | ( n28194 & ~n28304 ) | ( n28195 & ~n28304 ) ;
  assign n28306 = ( ~n28195 & n28304 ) | ( ~n28195 & n28305 ) | ( n28304 & n28305 ) ;
  assign n28307 = ( ~n28194 & n28305 ) | ( ~n28194 & n28306 ) | ( n28305 & n28306 ) ;
  assign n28308 = n28034 | n28168 ;
  assign n28309 = n28307 & n28308 ;
  assign n28310 = n28307 & ~n28309 ;
  assign n28311 = ~n28307 & n28308 ;
  assign n28312 = n28310 | n28311 ;
  assign n28313 = n28171 | n28178 ;
  assign n28314 = n28312 & n28313 ;
  assign n28315 = n28312 | n28313 ;
  assign n28316 = ~n28314 & n28315 ;
  assign n28317 = ~n28183 & n28316 ;
  assign n28318 = n28183 & ~n28316 ;
  assign n28319 = n28317 | n28318 ;
  assign n28320 = ( n28194 & n28195 ) | ( n28194 & n28304 ) | ( n28195 & n28304 ) ;
  assign n28321 = n12319 & n26156 ;
  assign n28322 = n5384 & n25928 ;
  assign n28323 = n28321 | n28322 ;
  assign n28324 = n39 | n28323 ;
  assign n28325 = ( n26165 & n28323 ) | ( n26165 & n28324 ) | ( n28323 & n28324 ) ;
  assign n28326 = x14 & n28325 ;
  assign n28327 = x14 & ~n28326 ;
  assign n28328 = ( n28325 & ~n28326 ) | ( n28325 & n28327 ) | ( ~n28326 & n28327 ) ;
  assign n28329 = n28288 | n28328 ;
  assign n28330 = n28302 | n28329 ;
  assign n28331 = ( n28288 & n28302 ) | ( n28288 & n28328 ) | ( n28302 & n28328 ) ;
  assign n28332 = n28330 & ~n28331 ;
  assign n28333 = ( n28205 & n28206 ) | ( n28205 & n28283 ) | ( n28206 & n28283 ) ;
  assign n28334 = ( n28216 & n28217 ) | ( n28216 & n28280 ) | ( n28217 & n28280 ) ;
  assign n28335 = n4484 & n20532 ;
  assign n28336 = n4479 & ~n20724 ;
  assign n28337 = n4481 & ~n20536 ;
  assign n28338 = n28336 | n28337 ;
  assign n28339 = n28335 | n28338 ;
  assign n28340 = n4487 | n28339 ;
  assign n28341 = ( n23203 & n28339 ) | ( n23203 & n28340 ) | ( n28339 & n28340 ) ;
  assign n28342 = x26 & n28341 ;
  assign n28343 = x26 & ~n28342 ;
  assign n28344 = ( n28341 & ~n28342 ) | ( n28341 & n28343 ) | ( ~n28342 & n28343 ) ;
  assign n28345 = n4048 & ~n20542 ;
  assign n28346 = n4043 & ~n20710 ;
  assign n28347 = n4045 & n20546 ;
  assign n28348 = n28346 | n28347 ;
  assign n28349 = n28345 | n28348 ;
  assign n28350 = n4051 | n28349 ;
  assign n28351 = ( ~n23042 & n28349 ) | ( ~n23042 & n28350 ) | ( n28349 & n28350 ) ;
  assign n28352 = ~x29 & n28351 ;
  assign n28353 = x29 | n28352 ;
  assign n28354 = ( ~n28351 & n28352 ) | ( ~n28351 & n28353 ) | ( n28352 & n28353 ) ;
  assign n28355 = n3744 & n20556 ;
  assign n28356 = n3639 & n20562 ;
  assign n28357 = n3727 & ~n20552 ;
  assign n28358 = n28356 | n28357 ;
  assign n28359 = n28355 | n28358 ;
  assign n28360 = n3636 | n28359 ;
  assign n28361 = ( ~n22655 & n28359 ) | ( ~n22655 & n28360 ) | ( n28359 & n28360 ) ;
  assign n28362 = ( n1203 & ~n1976 ) | ( n1203 & n5218 ) | ( ~n1976 & n5218 ) ;
  assign n28363 = n1976 | n28362 ;
  assign n28364 = n128 | n28363 ;
  assign n28365 = n10914 | n28364 ;
  assign n28366 = n3668 | n28365 ;
  assign n28367 = n11323 | n28366 ;
  assign n28368 = n2427 | n3565 ;
  assign n28369 = n4280 & ~n28368 ;
  assign n28370 = ~n28367 & n28369 ;
  assign n28371 = n281 | n514 ;
  assign n28372 = n520 | n28371 ;
  assign n28373 = n299 | n28372 ;
  assign n28374 = n269 | n28373 ;
  assign n28375 = n383 | n28374 ;
  assign n28376 = n197 | n28375 ;
  assign n28377 = n108 | n28376 ;
  assign n28378 = n218 | n28377 ;
  assign n28379 = n28370 & ~n28378 ;
  assign n28380 = n28243 & n28379 ;
  assign n28381 = n28243 | n28379 ;
  assign n28382 = n28360 & n28381 ;
  assign n28383 = ~n28380 & n28382 ;
  assign n28384 = n28359 & n28381 ;
  assign n28385 = ~n28380 & n28384 ;
  assign n28386 = ( ~n22655 & n28383 ) | ( ~n22655 & n28385 ) | ( n28383 & n28385 ) ;
  assign n28387 = n28361 & ~n28386 ;
  assign n28388 = ( n28226 & n28247 ) | ( n28226 & ~n28250 ) | ( n28247 & ~n28250 ) ;
  assign n28389 = n28244 & ~n28388 ;
  assign n28390 = n28381 & ~n28386 ;
  assign n28391 = ~n28380 & n28390 ;
  assign n28392 = ~n28389 & n28391 ;
  assign n28393 = ( n28387 & ~n28389 ) | ( n28387 & n28392 ) | ( ~n28389 & n28392 ) ;
  assign n28394 = n28389 & ~n28391 ;
  assign n28395 = ~n28387 & n28394 ;
  assign n28396 = n28393 | n28395 ;
  assign n28397 = n28252 | n28265 ;
  assign n28398 = n28396 & ~n28397 ;
  assign n28399 = ~n28396 & n28397 ;
  assign n28400 = n28398 | n28399 ;
  assign n28401 = n28354 & ~n28400 ;
  assign n28402 = n28400 | n28401 ;
  assign n28403 = ( ~n28354 & n28401 ) | ( ~n28354 & n28402 ) | ( n28401 & n28402 ) ;
  assign n28404 = n28344 & ~n28403 ;
  assign n28405 = ~n28344 & n28403 ;
  assign n28406 = n28404 | n28405 ;
  assign n28407 = ~n28278 & n28406 ;
  assign n28408 = n28278 & ~n28406 ;
  assign n28409 = n28407 | n28408 ;
  assign n28410 = n4551 & ~n21005 ;
  assign n28411 = n4546 & n20838 ;
  assign n28412 = n4548 & n20921 ;
  assign n28413 = n28411 | n28412 ;
  assign n28414 = n28410 | n28413 ;
  assign n28415 = n4554 | n28414 ;
  assign n28416 = ( ~n21015 & n28414 ) | ( ~n21015 & n28415 ) | ( n28414 & n28415 ) ;
  assign n28417 = ~x23 & n28416 ;
  assign n28418 = x23 | n28417 ;
  assign n28419 = ( ~n28416 & n28417 ) | ( ~n28416 & n28418 ) | ( n28417 & n28418 ) ;
  assign n28420 = n28409 & n28419 ;
  assign n28421 = ( n28278 & ~n28406 ) | ( n28278 & n28419 ) | ( ~n28406 & n28419 ) ;
  assign n28422 = n28407 | n28421 ;
  assign n28423 = ~n28420 & n28422 ;
  assign n28424 = ~n28334 & n28423 ;
  assign n28425 = n28334 & ~n28423 ;
  assign n28426 = n28424 | n28425 ;
  assign n28427 = n4781 & n24324 ;
  assign n28428 = n4776 & n24329 ;
  assign n28429 = n4778 & ~n24334 ;
  assign n28430 = n28428 | n28429 ;
  assign n28431 = n28427 | n28430 ;
  assign n28432 = n4784 & ~n24353 ;
  assign n28433 = ( n4784 & n24356 ) | ( n4784 & n28432 ) | ( n24356 & n28432 ) ;
  assign n28434 = n28431 | n28433 ;
  assign n28435 = x20 | n28434 ;
  assign n28436 = ~x20 & n28435 ;
  assign n28437 = ( ~n28434 & n28435 ) | ( ~n28434 & n28436 ) | ( n28435 & n28436 ) ;
  assign n28438 = n28426 & n28437 ;
  assign n28439 = ( n28334 & ~n28423 ) | ( n28334 & n28437 ) | ( ~n28423 & n28437 ) ;
  assign n28440 = n28424 | n28439 ;
  assign n28441 = ~n28438 & n28440 ;
  assign n28442 = ~n28333 & n28441 ;
  assign n28443 = n28333 & ~n28441 ;
  assign n28444 = n28442 | n28443 ;
  assign n28445 = n5083 & ~n25676 ;
  assign n28446 = n5069 & n25187 ;
  assign n28447 = n5070 & n25442 ;
  assign n28448 = n28446 | n28447 ;
  assign n28449 = n28445 | n28448 ;
  assign n28450 = n5074 & ~n25690 ;
  assign n28451 = ( n5074 & n25694 ) | ( n5074 & n28450 ) | ( n25694 & n28450 ) ;
  assign n28452 = n28449 | n28451 ;
  assign n28453 = x17 | n28452 ;
  assign n28454 = ~x17 & n28453 ;
  assign n28455 = ( ~n28452 & n28453 ) | ( ~n28452 & n28454 ) | ( n28453 & n28454 ) ;
  assign n28456 = n28444 & n28455 ;
  assign n28457 = ( n28333 & ~n28441 ) | ( n28333 & n28455 ) | ( ~n28441 & n28455 ) ;
  assign n28458 = n28442 | n28457 ;
  assign n28459 = ~n28456 & n28458 ;
  assign n28460 = n28332 & ~n28459 ;
  assign n28461 = n28459 | n28460 ;
  assign n28462 = ( ~n28332 & n28460 ) | ( ~n28332 & n28461 ) | ( n28460 & n28461 ) ;
  assign n28463 = ~n28320 & n28462 ;
  assign n28464 = n28320 & ~n28462 ;
  assign n28465 = n28463 | n28464 ;
  assign n28466 = n28309 & ~n28465 ;
  assign n28467 = ( n28314 & ~n28465 ) | ( n28314 & n28466 ) | ( ~n28465 & n28466 ) ;
  assign n28468 = ~n28309 & n28465 ;
  assign n28469 = ~n28314 & n28468 ;
  assign n28470 = n28467 | n28469 ;
  assign n28471 = ~n28181 & n28316 ;
  assign n28472 = n28021 & n28471 ;
  assign n28473 = n28470 & ~n28472 ;
  assign n28474 = ( ~n28470 & n28472 ) | ( ~n28470 & n28473 ) | ( n28472 & n28473 ) ;
  assign n28475 = n28473 | n28474 ;
  assign n28476 = n5083 & n25928 ;
  assign n28477 = n5069 & n25442 ;
  assign n28478 = n5070 & ~n25676 ;
  assign n28479 = n28477 | n28478 ;
  assign n28480 = n28476 | n28479 ;
  assign n28481 = n5074 | n28480 ;
  assign n28482 = ( ~n25936 & n28480 ) | ( ~n25936 & n28481 ) | ( n28480 & n28481 ) ;
  assign n28483 = ~x17 & n28482 ;
  assign n28484 = x17 | n28483 ;
  assign n28485 = ( ~n28482 & n28483 ) | ( ~n28482 & n28484 ) | ( n28483 & n28484 ) ;
  assign n28486 = n28457 & n28485 ;
  assign n28487 = n28457 & ~n28486 ;
  assign n28488 = n4551 & n24329 ;
  assign n28489 = n4546 & n20921 ;
  assign n28490 = n4548 & ~n21005 ;
  assign n28491 = n28489 | n28490 ;
  assign n28492 = n28488 | n28491 ;
  assign n28493 = ( n4554 & ~n24391 ) | ( n4554 & n24392 ) | ( ~n24391 & n24392 ) ;
  assign n28494 = n28492 | n28493 ;
  assign n28495 = x23 | n28494 ;
  assign n28496 = ~x23 & n28495 ;
  assign n28497 = ( ~n28494 & n28495 ) | ( ~n28494 & n28496 ) | ( n28495 & n28496 ) ;
  assign n28498 = n28421 & n28497 ;
  assign n28499 = n28421 & ~n28498 ;
  assign n28500 = n28401 | n28404 ;
  assign n28501 = n4484 & n20838 ;
  assign n28502 = n4479 & ~n20536 ;
  assign n28503 = n4481 & n20532 ;
  assign n28504 = n28502 | n28503 ;
  assign n28505 = n28501 | n28504 ;
  assign n28506 = n4487 | n28505 ;
  assign n28507 = ( ~n23712 & n28505 ) | ( ~n23712 & n28506 ) | ( n28505 & n28506 ) ;
  assign n28508 = ~x26 & n28507 ;
  assign n28509 = x26 | n28508 ;
  assign n28510 = ( ~n28507 & n28508 ) | ( ~n28507 & n28509 ) | ( n28508 & n28509 ) ;
  assign n28511 = n28393 | n28399 ;
  assign n28512 = n4048 & ~n20724 ;
  assign n28513 = n4043 & n20546 ;
  assign n28514 = n4045 & ~n20542 ;
  assign n28515 = n28513 | n28514 ;
  assign n28516 = n28512 | n28515 ;
  assign n28517 = n4051 | n28516 ;
  assign n28518 = ( n23229 & n28516 ) | ( n23229 & n28517 ) | ( n28516 & n28517 ) ;
  assign n28519 = x29 & n28518 ;
  assign n28520 = x29 & ~n28519 ;
  assign n28521 = ( n28518 & ~n28519 ) | ( n28518 & n28520 ) | ( ~n28519 & n28520 ) ;
  assign n28522 = n3744 & ~n20710 ;
  assign n28523 = n3639 & ~n20552 ;
  assign n28524 = n3727 & n20556 ;
  assign n28525 = n28523 | n28524 ;
  assign n28526 = n28522 | n28525 ;
  assign n28527 = n3636 | n28526 ;
  assign n28528 = ( ~n22641 & n28526 ) | ( ~n22641 & n28527 ) | ( n28526 & n28527 ) ;
  assign n28529 = n2578 | n11275 ;
  assign n28530 = n12762 | n28529 ;
  assign n28531 = n1737 | n28530 ;
  assign n28532 = n13615 | n28531 ;
  assign n28533 = n13612 | n28532 ;
  assign n28534 = n5670 & ~n28533 ;
  assign n28535 = ~n3096 & n28534 ;
  assign n28536 = ~n1454 & n28535 ;
  assign n28537 = n922 | n1352 ;
  assign n28538 = n383 | n28537 ;
  assign n28539 = n419 | n28538 ;
  assign n28540 = n610 | n28539 ;
  assign n28541 = n28536 & ~n28540 ;
  assign n28542 = ~n28243 & n28541 ;
  assign n28543 = n28243 & ~n28541 ;
  assign n28544 = n28542 | n28543 ;
  assign n28545 = n19606 & n26156 ;
  assign n28546 = ~x14 & n28545 ;
  assign n28547 = x14 | n28546 ;
  assign n28548 = ( ~n28545 & n28546 ) | ( ~n28545 & n28547 ) | ( n28546 & n28547 ) ;
  assign n28549 = n28544 | n28548 ;
  assign n28550 = n28544 & n28548 ;
  assign n28551 = n28549 & ~n28550 ;
  assign n28552 = ( n28390 & n28528 ) | ( n28390 & ~n28551 ) | ( n28528 & ~n28551 ) ;
  assign n28553 = ( ~n28390 & n28551 ) | ( ~n28390 & n28552 ) | ( n28551 & n28552 ) ;
  assign n28554 = ( ~n28528 & n28552 ) | ( ~n28528 & n28553 ) | ( n28552 & n28553 ) ;
  assign n28555 = n28521 & ~n28554 ;
  assign n28556 = n28554 | n28555 ;
  assign n28557 = ( ~n28521 & n28555 ) | ( ~n28521 & n28556 ) | ( n28555 & n28556 ) ;
  assign n28558 = ~n28511 & n28557 ;
  assign n28559 = n28511 & ~n28557 ;
  assign n28560 = n28558 | n28559 ;
  assign n28561 = n28510 & ~n28560 ;
  assign n28562 = n28560 | n28561 ;
  assign n28563 = ( ~n28510 & n28561 ) | ( ~n28510 & n28562 ) | ( n28561 & n28562 ) ;
  assign n28564 = ~n28500 & n28563 ;
  assign n28565 = n28500 & ~n28563 ;
  assign n28566 = n28564 | n28565 ;
  assign n28567 = ~n28421 & n28497 ;
  assign n28568 = n28566 & ~n28567 ;
  assign n28569 = ~n28499 & n28568 ;
  assign n28570 = ( n28499 & ~n28566 ) | ( n28499 & n28567 ) | ( ~n28566 & n28567 ) ;
  assign n28571 = n28569 | n28570 ;
  assign n28572 = n4781 & n25187 ;
  assign n28573 = n4776 & ~n24334 ;
  assign n28574 = n4778 & n24324 ;
  assign n28575 = n28573 | n28574 ;
  assign n28576 = n28572 | n28575 ;
  assign n28577 = n4784 | n28576 ;
  assign n28578 = ( n25193 & n28576 ) | ( n25193 & n28577 ) | ( n28576 & n28577 ) ;
  assign n28579 = x20 & n28578 ;
  assign n28580 = x20 & ~n28579 ;
  assign n28581 = ( n28578 & ~n28579 ) | ( n28578 & n28580 ) | ( ~n28579 & n28580 ) ;
  assign n28582 = ~n28571 & n28581 ;
  assign n28583 = n28571 | n28582 ;
  assign n28584 = n28571 & n28581 ;
  assign n28585 = n28439 | n28584 ;
  assign n28586 = n28583 & ~n28585 ;
  assign n28587 = ( n28439 & ~n28583 ) | ( n28439 & n28584 ) | ( ~n28583 & n28584 ) ;
  assign n28588 = n28586 | n28587 ;
  assign n28589 = ~n28457 & n28485 ;
  assign n28590 = n28588 & ~n28589 ;
  assign n28591 = ~n28487 & n28590 ;
  assign n28592 = ( n28487 & ~n28588 ) | ( n28487 & n28589 ) | ( ~n28588 & n28589 ) ;
  assign n28593 = n28591 | n28592 ;
  assign n28594 = n28331 | n28460 ;
  assign n28595 = ~n28593 & n28594 ;
  assign n28596 = n28593 & ~n28594 ;
  assign n28597 = n28595 | n28596 ;
  assign n28598 = n28464 | n28466 ;
  assign n28599 = ~n28597 & n28598 ;
  assign n28600 = n28463 | n28597 ;
  assign n28601 = ( n28314 & n28599 ) | ( n28314 & ~n28600 ) | ( n28599 & ~n28600 ) ;
  assign n28602 = ( n28314 & ~n28463 ) | ( n28314 & n28598 ) | ( ~n28463 & n28598 ) ;
  assign n28603 = n28597 & ~n28602 ;
  assign n28604 = n28601 | n28603 ;
  assign n28605 = ~n28474 & n28604 ;
  assign n28606 = ( n28474 & ~n28604 ) | ( n28474 & n28605 ) | ( ~n28604 & n28605 ) ;
  assign n28607 = n28605 | n28606 ;
  assign n28608 = n28582 | n28587 ;
  assign n28609 = n28498 | n28570 ;
  assign n28610 = n28561 | n28565 ;
  assign n28611 = n4484 & n20921 ;
  assign n28612 = n4479 & n20532 ;
  assign n28613 = n4481 & n20838 ;
  assign n28614 = n28612 | n28613 ;
  assign n28615 = n28611 | n28614 ;
  assign n28616 = ( n4487 & n23691 ) | ( n4487 & n23695 ) | ( n23691 & n23695 ) ;
  assign n28617 = n28615 | n28616 ;
  assign n28618 = x26 | n28617 ;
  assign n28619 = ~x26 & n28618 ;
  assign n28620 = ( ~n28617 & n28618 ) | ( ~n28617 & n28619 ) | ( n28618 & n28619 ) ;
  assign n28621 = n3744 & n20546 ;
  assign n28622 = n3639 & n20556 ;
  assign n28623 = n3727 & ~n20710 ;
  assign n28624 = n28622 | n28623 ;
  assign n28625 = n28621 | n28624 ;
  assign n28626 = n3636 & ~n21031 ;
  assign n28627 = ( n3636 & n21037 ) | ( n3636 & n28626 ) | ( n21037 & n28626 ) ;
  assign n28628 = n28625 | n28627 ;
  assign n28629 = n2199 | n2924 ;
  assign n28630 = n3551 | n28629 ;
  assign n28631 = n12646 | n28630 ;
  assign n28632 = n4955 | n28631 ;
  assign n28633 = n4110 | n28632 ;
  assign n28634 = n1852 | n3314 ;
  assign n28635 = n1337 | n28634 ;
  assign n28636 = n2219 | n28635 ;
  assign n28637 = n28633 | n28636 ;
  assign n28638 = ~n166 & n2662 ;
  assign n28639 = ~n28637 & n28638 ;
  assign n28640 = n629 | n2623 ;
  assign n28641 = n307 | n28640 ;
  assign n28642 = n96 | n28641 ;
  assign n28643 = n146 | n28642 ;
  assign n28644 = n28639 & ~n28643 ;
  assign n28645 = ( n28543 & ~n28549 ) | ( n28543 & n28644 ) | ( ~n28549 & n28644 ) ;
  assign n28646 = ( n28542 & ~n28543 ) | ( n28542 & n28548 ) | ( ~n28543 & n28548 ) ;
  assign n28647 = ~n28644 & n28646 ;
  assign n28648 = n28645 | n28647 ;
  assign n28649 = n28628 | n28648 ;
  assign n28650 = ~n28648 & n28649 ;
  assign n28651 = ( ~n28628 & n28649 ) | ( ~n28628 & n28650 ) | ( n28649 & n28650 ) ;
  assign n28652 = ~n28553 & n28651 ;
  assign n28653 = n28553 & ~n28651 ;
  assign n28654 = n28652 | n28653 ;
  assign n28655 = n4048 & ~n20536 ;
  assign n28656 = n4043 & ~n20542 ;
  assign n28657 = n4045 & ~n20724 ;
  assign n28658 = n28656 | n28657 ;
  assign n28659 = n28655 | n28658 ;
  assign n28660 = n4051 & ~n23213 ;
  assign n28661 = n23217 & n28660 ;
  assign n28662 = ( n4051 & n28659 ) | ( n4051 & ~n28661 ) | ( n28659 & ~n28661 ) ;
  assign n28663 = x29 & n28662 ;
  assign n28664 = x29 & ~n28663 ;
  assign n28665 = ( n28662 & ~n28663 ) | ( n28662 & n28664 ) | ( ~n28663 & n28664 ) ;
  assign n28666 = ~n28654 & n28665 ;
  assign n28667 = n28654 & ~n28665 ;
  assign n28668 = n28666 | n28667 ;
  assign n28669 = n28555 | n28559 ;
  assign n28670 = ( n28620 & n28668 ) | ( n28620 & ~n28669 ) | ( n28668 & ~n28669 ) ;
  assign n28671 = ( ~n28668 & n28669 ) | ( ~n28668 & n28670 ) | ( n28669 & n28670 ) ;
  assign n28672 = ( ~n28620 & n28670 ) | ( ~n28620 & n28671 ) | ( n28670 & n28671 ) ;
  assign n28673 = ~n28610 & n28672 ;
  assign n28674 = n28610 & ~n28672 ;
  assign n28675 = n28673 | n28674 ;
  assign n28676 = n4551 & ~n24334 ;
  assign n28677 = n4546 & ~n21005 ;
  assign n28678 = n4548 & n24329 ;
  assign n28679 = n28677 | n28678 ;
  assign n28680 = n28676 | n28679 ;
  assign n28681 = ( n4554 & ~n24373 ) | ( n4554 & n24376 ) | ( ~n24373 & n24376 ) ;
  assign n28682 = n28680 | n28681 ;
  assign n28683 = x23 | n28682 ;
  assign n28684 = ~x23 & n28683 ;
  assign n28685 = ( ~n28682 & n28683 ) | ( ~n28682 & n28684 ) | ( n28683 & n28684 ) ;
  assign n28686 = n28675 & n28685 ;
  assign n28687 = ( n28610 & ~n28672 ) | ( n28610 & n28685 ) | ( ~n28672 & n28685 ) ;
  assign n28688 = n28673 | n28687 ;
  assign n28689 = ~n28686 & n28688 ;
  assign n28690 = n28609 & ~n28689 ;
  assign n28691 = n28609 & ~n28690 ;
  assign n28692 = n28609 | n28689 ;
  assign n28693 = ~n28691 & n28692 ;
  assign n28694 = n4781 & n25442 ;
  assign n28695 = n4776 & n24324 ;
  assign n28696 = n4778 & n25187 ;
  assign n28697 = n28695 | n28696 ;
  assign n28698 = n28694 | n28697 ;
  assign n28699 = n4784 | n28698 ;
  assign n28700 = ( n25452 & n28698 ) | ( n25452 & n28699 ) | ( n28698 & n28699 ) ;
  assign n28701 = x20 & n28700 ;
  assign n28702 = x20 & ~n28701 ;
  assign n28703 = ( n28700 & ~n28701 ) | ( n28700 & n28702 ) | ( ~n28701 & n28702 ) ;
  assign n28704 = ~n28693 & n28703 ;
  assign n28705 = n28693 & ~n28703 ;
  assign n28706 = n28704 | n28705 ;
  assign n28707 = ~n28608 & n28706 ;
  assign n28708 = n28608 & ~n28706 ;
  assign n28709 = n28707 | n28708 ;
  assign n28710 = n5083 & n26156 ;
  assign n28711 = n5069 & ~n25676 ;
  assign n28712 = n5070 & n25928 ;
  assign n28713 = n28711 | n28712 ;
  assign n28714 = n28710 | n28713 ;
  assign n28715 = n5074 | n28714 ;
  assign n28716 = ( n26167 & n28714 ) | ( n26167 & n28715 ) | ( n28714 & n28715 ) ;
  assign n28717 = x17 & n28716 ;
  assign n28718 = x17 & ~n28717 ;
  assign n28719 = ( n28716 & ~n28717 ) | ( n28716 & n28718 ) | ( ~n28717 & n28718 ) ;
  assign n28720 = n28709 & n28719 ;
  assign n28721 = ( n28608 & ~n28706 ) | ( n28608 & n28719 ) | ( ~n28706 & n28719 ) ;
  assign n28722 = n28707 | n28721 ;
  assign n28723 = ~n28720 & n28722 ;
  assign n28724 = n28486 | n28592 ;
  assign n28725 = ~n28723 & n28724 ;
  assign n28726 = n28723 | n28725 ;
  assign n28727 = n28724 & ~n28725 ;
  assign n28728 = n28726 & ~n28727 ;
  assign n28729 = n28595 | n28599 ;
  assign n28730 = ~n28728 & n28729 ;
  assign n28731 = ~n28595 & n28600 ;
  assign n28732 = n28728 | n28731 ;
  assign n28733 = ( n28314 & n28730 ) | ( n28314 & ~n28732 ) | ( n28730 & ~n28732 ) ;
  assign n28734 = ( n28314 & n28729 ) | ( n28314 & ~n28731 ) | ( n28729 & ~n28731 ) ;
  assign n28735 = n28728 & ~n28734 ;
  assign n28736 = n28733 | n28735 ;
  assign n28737 = n28606 & ~n28736 ;
  assign n28738 = n28736 | n28737 ;
  assign n28739 = ( ~n28606 & n28737 ) | ( ~n28606 & n28738 ) | ( n28737 & n28738 ) ;
  assign n28740 = n19762 & n26156 ;
  assign n28741 = n5069 & n25928 ;
  assign n28742 = n28740 | n28741 ;
  assign n28743 = n5074 | n28742 ;
  assign n28744 = ( n26165 & n28742 ) | ( n26165 & n28743 ) | ( n28742 & n28743 ) ;
  assign n28745 = x17 & n28744 ;
  assign n28746 = x17 & ~n28745 ;
  assign n28747 = ( n28744 & ~n28745 ) | ( n28744 & n28746 ) | ( ~n28745 & n28746 ) ;
  assign n28748 = n28690 | n28747 ;
  assign n28749 = n28704 | n28748 ;
  assign n28750 = ( n28690 & n28704 ) | ( n28690 & n28747 ) | ( n28704 & n28747 ) ;
  assign n28751 = n28749 & ~n28750 ;
  assign n28752 = n4781 & ~n25676 ;
  assign n28753 = n4776 & n25187 ;
  assign n28754 = n4778 & n25442 ;
  assign n28755 = n28753 | n28754 ;
  assign n28756 = n28752 | n28755 ;
  assign n28757 = n4784 & ~n25690 ;
  assign n28758 = ( n4784 & n25694 ) | ( n4784 & n28757 ) | ( n25694 & n28757 ) ;
  assign n28759 = n28756 | n28758 ;
  assign n28760 = x20 | n28759 ;
  assign n28761 = ~x20 & n28760 ;
  assign n28762 = ( ~n28759 & n28760 ) | ( ~n28759 & n28761 ) | ( n28760 & n28761 ) ;
  assign n28763 = n4551 & n24324 ;
  assign n28764 = n4546 & n24329 ;
  assign n28765 = n4548 & ~n24334 ;
  assign n28766 = n28764 | n28765 ;
  assign n28767 = n28763 | n28766 ;
  assign n28768 = n4554 & ~n24353 ;
  assign n28769 = ( n4554 & n24356 ) | ( n4554 & n28768 ) | ( n24356 & n28768 ) ;
  assign n28770 = n28767 | n28769 ;
  assign n28771 = x23 | n28770 ;
  assign n28772 = ~x23 & n28771 ;
  assign n28773 = ( ~n28770 & n28771 ) | ( ~n28770 & n28772 ) | ( n28771 & n28772 ) ;
  assign n28774 = n28653 | n28666 ;
  assign n28775 = n28625 & ~n28648 ;
  assign n28776 = n28645 | n28775 ;
  assign n28777 = ( n28627 & ~n28647 ) | ( n28627 & n28776 ) | ( ~n28647 & n28776 ) ;
  assign n28778 = n1221 | n1889 ;
  assign n28779 = n428 | n626 ;
  assign n28780 = n1416 | n28779 ;
  assign n28781 = n28778 | n28780 ;
  assign n28782 = n952 | n28781 ;
  assign n28783 = n10934 | n28782 ;
  assign n28784 = n4324 | n28783 ;
  assign n28785 = n3171 | n28784 ;
  assign n28786 = n367 | n2385 ;
  assign n28787 = n3444 | n28786 ;
  assign n28788 = n2341 | n28787 ;
  assign n28789 = n484 | n28788 ;
  assign n28790 = n326 | n28789 ;
  assign n28791 = n191 | n28790 ;
  assign n28792 = n28785 | n28791 ;
  assign n28793 = n81 | n120 ;
  assign n28794 = n152 | n28793 ;
  assign n28795 = n28792 | n28794 ;
  assign n28796 = n28644 & n28795 ;
  assign n28797 = n28644 | n28795 ;
  assign n28798 = n28776 & n28797 ;
  assign n28799 = ~n28796 & n28798 ;
  assign n28800 = ~n28647 & n28797 ;
  assign n28801 = ~n28796 & n28800 ;
  assign n28802 = ( n28627 & n28799 ) | ( n28627 & n28801 ) | ( n28799 & n28801 ) ;
  assign n28803 = n28777 & ~n28802 ;
  assign n28804 = n28797 & ~n28802 ;
  assign n28805 = ~n28796 & n28804 ;
  assign n28806 = n28803 | n28805 ;
  assign n28807 = n3744 & ~n20542 ;
  assign n28808 = n3639 & ~n20710 ;
  assign n28809 = n3727 & n20546 ;
  assign n28810 = n28808 | n28809 ;
  assign n28811 = n28807 | n28810 ;
  assign n28812 = n3636 | n28811 ;
  assign n28813 = ( ~n23042 & n28811 ) | ( ~n23042 & n28812 ) | ( n28811 & n28812 ) ;
  assign n28814 = n28806 & n28813 ;
  assign n28815 = n28806 | n28813 ;
  assign n28816 = ~n28814 & n28815 ;
  assign n28817 = n4048 & n20532 ;
  assign n28818 = n4043 & ~n20724 ;
  assign n28819 = n4045 & ~n20536 ;
  assign n28820 = n28818 | n28819 ;
  assign n28821 = n28817 | n28820 ;
  assign n28822 = n4051 | n28821 ;
  assign n28823 = ( n23203 & n28821 ) | ( n23203 & n28822 ) | ( n28821 & n28822 ) ;
  assign n28824 = x29 & n28823 ;
  assign n28825 = x29 & ~n28824 ;
  assign n28826 = ( n28823 & ~n28824 ) | ( n28823 & n28825 ) | ( ~n28824 & n28825 ) ;
  assign n28827 = n28816 & n28826 ;
  assign n28828 = n28816 | n28826 ;
  assign n28829 = ~n28827 & n28828 ;
  assign n28830 = n4484 & ~n21005 ;
  assign n28831 = n4479 & n20838 ;
  assign n28832 = n4481 & n20921 ;
  assign n28833 = n28831 | n28832 ;
  assign n28834 = n28830 | n28833 ;
  assign n28835 = n4487 | n28834 ;
  assign n28836 = ( ~n21015 & n28834 ) | ( ~n21015 & n28835 ) | ( n28834 & n28835 ) ;
  assign n28837 = ~x26 & n28836 ;
  assign n28838 = x26 | n28837 ;
  assign n28839 = ( ~n28836 & n28837 ) | ( ~n28836 & n28838 ) | ( n28837 & n28838 ) ;
  assign n28840 = ( n28774 & n28829 ) | ( n28774 & n28839 ) | ( n28829 & n28839 ) ;
  assign n28841 = ( n28829 & n28839 ) | ( n28829 & ~n28840 ) | ( n28839 & ~n28840 ) ;
  assign n28842 = ( n28774 & ~n28840 ) | ( n28774 & n28841 ) | ( ~n28840 & n28841 ) ;
  assign n28843 = ( ~n28671 & n28773 ) | ( ~n28671 & n28842 ) | ( n28773 & n28842 ) ;
  assign n28844 = ( n28671 & ~n28842 ) | ( n28671 & n28843 ) | ( ~n28842 & n28843 ) ;
  assign n28845 = ( ~n28773 & n28843 ) | ( ~n28773 & n28844 ) | ( n28843 & n28844 ) ;
  assign n28846 = ( n28687 & n28762 ) | ( n28687 & ~n28845 ) | ( n28762 & ~n28845 ) ;
  assign n28847 = ( ~n28687 & n28845 ) | ( ~n28687 & n28846 ) | ( n28845 & n28846 ) ;
  assign n28848 = ( ~n28762 & n28846 ) | ( ~n28762 & n28847 ) | ( n28846 & n28847 ) ;
  assign n28849 = n28751 & ~n28848 ;
  assign n28850 = n28848 | n28849 ;
  assign n28851 = ( ~n28751 & n28849 ) | ( ~n28751 & n28850 ) | ( n28849 & n28850 ) ;
  assign n28852 = n28721 | n28851 ;
  assign n28853 = n28721 & n28851 ;
  assign n28854 = n28852 & ~n28853 ;
  assign n28855 = n28725 | n28730 ;
  assign n28856 = n28854 & n28855 ;
  assign n28857 = ~n28725 & n28732 ;
  assign n28858 = n28854 & ~n28857 ;
  assign n28859 = ( n28314 & n28856 ) | ( n28314 & n28858 ) | ( n28856 & n28858 ) ;
  assign n28860 = ( n28314 & n28855 ) | ( n28314 & ~n28857 ) | ( n28855 & ~n28857 ) ;
  assign n28861 = n28854 | n28860 ;
  assign n28862 = ~n28859 & n28861 ;
  assign n28863 = n28737 | n28862 ;
  assign n28864 = ~n28736 & n28862 ;
  assign n28865 = n28606 & n28864 ;
  assign n28866 = n28863 & ~n28865 ;
  assign n28867 = ( n28687 & n28762 ) | ( n28687 & n28845 ) | ( n28762 & n28845 ) ;
  assign n28868 = n4781 & n25928 ;
  assign n28869 = n4776 & n25442 ;
  assign n28870 = n4778 & ~n25676 ;
  assign n28871 = n28869 | n28870 ;
  assign n28872 = n28868 | n28871 ;
  assign n28873 = n4784 | n28872 ;
  assign n28874 = ( ~n25936 & n28872 ) | ( ~n25936 & n28873 ) | ( n28872 & n28873 ) ;
  assign n28875 = ~x20 & n28874 ;
  assign n28876 = x20 | n28875 ;
  assign n28877 = ( ~n28874 & n28875 ) | ( ~n28874 & n28876 ) | ( n28875 & n28876 ) ;
  assign n28878 = n28867 & n28877 ;
  assign n28879 = n28867 & ~n28878 ;
  assign n28880 = ( n28671 & n28773 ) | ( n28671 & n28842 ) | ( n28773 & n28842 ) ;
  assign n28881 = n4048 & n20838 ;
  assign n28882 = n4043 & ~n20536 ;
  assign n28883 = n4045 & n20532 ;
  assign n28884 = n28882 | n28883 ;
  assign n28885 = n28881 | n28884 ;
  assign n28886 = n4051 | n28885 ;
  assign n28887 = ( ~n23712 & n28885 ) | ( ~n23712 & n28886 ) | ( n28885 & n28886 ) ;
  assign n28888 = ~x29 & n28887 ;
  assign n28889 = x29 | n28888 ;
  assign n28890 = ( ~n28887 & n28888 ) | ( ~n28887 & n28889 ) | ( n28888 & n28889 ) ;
  assign n28891 = n3744 & ~n20724 ;
  assign n28892 = n3639 & n20546 ;
  assign n28893 = n3727 & ~n20542 ;
  assign n28894 = n28892 | n28893 ;
  assign n28895 = n28891 | n28894 ;
  assign n28896 = n3636 | n28895 ;
  assign n28897 = ( n23229 & n28895 ) | ( n23229 & n28896 ) | ( n28895 & n28896 ) ;
  assign n28898 = n1356 | n21774 ;
  assign n28899 = n2626 | n28898 ;
  assign n28900 = n3862 | n28899 ;
  assign n28901 = n11538 | n28900 ;
  assign n28902 = n1277 | n19837 ;
  assign n28903 = n3273 | n28902 ;
  assign n28904 = n3204 | n28903 ;
  assign n28905 = n432 | n28904 ;
  assign n28906 = n28901 | n28905 ;
  assign n28907 = n338 | n510 ;
  assign n28908 = n81 | n28907 ;
  assign n28909 = n157 | n28908 ;
  assign n28910 = n28906 | n28909 ;
  assign n28911 = n28795 | n28910 ;
  assign n28912 = n28795 & n28910 ;
  assign n28913 = n28911 & ~n28912 ;
  assign n28914 = n19764 & n26156 ;
  assign n28915 = ~x17 & n28914 ;
  assign n28916 = x17 | n28915 ;
  assign n28917 = ( ~n28914 & n28915 ) | ( ~n28914 & n28916 ) | ( n28915 & n28916 ) ;
  assign n28918 = n28913 & ~n28917 ;
  assign n28919 = ~n28913 & n28917 ;
  assign n28920 = n28918 | n28919 ;
  assign n28921 = n28897 & ~n28920 ;
  assign n28922 = n28897 & ~n28921 ;
  assign n28923 = n28897 | n28920 ;
  assign n28924 = ~n28922 & n28923 ;
  assign n28925 = n28804 | n28924 ;
  assign n28926 = n28804 & n28924 ;
  assign n28927 = n28925 & ~n28926 ;
  assign n28928 = n28814 | n28827 ;
  assign n28929 = n28927 & n28928 ;
  assign n28930 = n28928 & ~n28929 ;
  assign n28931 = ( n28927 & ~n28929 ) | ( n28927 & n28930 ) | ( ~n28929 & n28930 ) ;
  assign n28932 = n28890 & n28931 ;
  assign n28933 = n28890 | n28931 ;
  assign n28934 = ~n28932 & n28933 ;
  assign n28935 = n4484 & n24329 ;
  assign n28936 = n4479 & n20921 ;
  assign n28937 = n4481 & ~n21005 ;
  assign n28938 = n28936 | n28937 ;
  assign n28939 = n28935 | n28938 ;
  assign n28940 = ( n4487 & ~n24391 ) | ( n4487 & n24392 ) | ( ~n24391 & n24392 ) ;
  assign n28941 = n28939 | n28940 ;
  assign n28942 = x26 | n28941 ;
  assign n28943 = ~x26 & n28942 ;
  assign n28944 = ( ~n28941 & n28942 ) | ( ~n28941 & n28943 ) | ( n28942 & n28943 ) ;
  assign n28945 = ( ~n28840 & n28934 ) | ( ~n28840 & n28944 ) | ( n28934 & n28944 ) ;
  assign n28946 = ( n28840 & ~n28944 ) | ( n28840 & n28945 ) | ( ~n28944 & n28945 ) ;
  assign n28947 = ( ~n28934 & n28945 ) | ( ~n28934 & n28946 ) | ( n28945 & n28946 ) ;
  assign n28948 = n4551 & n25187 ;
  assign n28949 = n4546 & ~n24334 ;
  assign n28950 = n4548 & n24324 ;
  assign n28951 = n28949 | n28950 ;
  assign n28952 = n28948 | n28951 ;
  assign n28953 = n4554 | n28952 ;
  assign n28954 = ( n25193 & n28952 ) | ( n25193 & n28953 ) | ( n28952 & n28953 ) ;
  assign n28955 = x23 & n28954 ;
  assign n28956 = x23 & ~n28955 ;
  assign n28957 = ( n28954 & ~n28955 ) | ( n28954 & n28956 ) | ( ~n28955 & n28956 ) ;
  assign n28958 = n28947 & n28957 ;
  assign n28959 = n28947 | n28957 ;
  assign n28960 = ~n28958 & n28959 ;
  assign n28961 = n28880 | n28960 ;
  assign n28962 = n28880 & n28960 ;
  assign n28963 = n28961 & ~n28962 ;
  assign n28964 = ~n28867 & n28877 ;
  assign n28965 = n28963 | n28964 ;
  assign n28966 = n28879 | n28965 ;
  assign n28967 = ( n28879 & n28963 ) | ( n28879 & n28964 ) | ( n28963 & n28964 ) ;
  assign n28968 = n28966 & ~n28967 ;
  assign n28969 = ( n28749 & n28750 ) | ( n28749 & n28848 ) | ( n28750 & n28848 ) ;
  assign n28970 = n28968 & n28969 ;
  assign n28971 = n28968 | n28969 ;
  assign n28972 = ~n28970 & n28971 ;
  assign n28973 = n28853 | n28856 ;
  assign n28974 = n28972 & n28973 ;
  assign n28975 = n28853 | n28858 ;
  assign n28976 = n28972 & n28975 ;
  assign n28977 = ( n28314 & n28974 ) | ( n28314 & n28976 ) | ( n28974 & n28976 ) ;
  assign n28978 = ( n28314 & n28973 ) | ( n28314 & n28975 ) | ( n28973 & n28975 ) ;
  assign n28979 = n28972 | n28978 ;
  assign n28980 = ~n28977 & n28979 ;
  assign n28981 = n28865 | n28980 ;
  assign n28982 = n28864 & n28980 ;
  assign n28983 = n28606 & n28982 ;
  assign n28984 = n28981 & ~n28983 ;
  assign n28985 = n28958 | n28962 ;
  assign n28986 = ~n28921 & n28925 ;
  assign n28987 = n3744 & ~n20536 ;
  assign n28988 = n3639 & ~n20542 ;
  assign n28989 = n3727 & ~n20724 ;
  assign n28990 = n28988 | n28989 ;
  assign n28991 = n28987 | n28990 ;
  assign n28992 = ( n3636 & n23213 ) | ( n3636 & ~n23217 ) | ( n23213 & ~n23217 ) ;
  assign n28993 = n28991 | n28992 ;
  assign n28994 = n1164 | n12242 ;
  assign n28995 = n2548 | n28994 ;
  assign n28996 = n6006 | n28995 ;
  assign n28997 = n2584 | n28996 ;
  assign n28998 = n798 | n28997 ;
  assign n28999 = n6004 | n28998 ;
  assign n29000 = ~n1311 & n27368 ;
  assign n29001 = ~n28999 & n29000 ;
  assign n29002 = ( n834 & ~n2389 ) | ( n834 & n3856 ) | ( ~n2389 & n3856 ) ;
  assign n29003 = n2389 | n29002 ;
  assign n29004 = n505 | n29003 ;
  assign n29005 = n277 | n29004 ;
  assign n29006 = n381 | n29005 ;
  assign n29007 = n215 | n29006 ;
  assign n29008 = n29001 & ~n29007 ;
  assign n29009 = ( n28912 & n28918 ) | ( n28912 & n29008 ) | ( n28918 & n29008 ) ;
  assign n29010 = ( n28911 & n28912 ) | ( n28911 & ~n28917 ) | ( n28912 & ~n28917 ) ;
  assign n29011 = n29008 | n29010 ;
  assign n29012 = ~n29009 & n29011 ;
  assign n29013 = n28993 | n29012 ;
  assign n29014 = ~n29012 & n29013 ;
  assign n29015 = ( ~n28993 & n29013 ) | ( ~n28993 & n29014 ) | ( n29013 & n29014 ) ;
  assign n29016 = n28986 & ~n29015 ;
  assign n29017 = ~n28986 & n29015 ;
  assign n29018 = n29016 | n29017 ;
  assign n29019 = n4048 & n20921 ;
  assign n29020 = n4043 & n20532 ;
  assign n29021 = n4045 & n20838 ;
  assign n29022 = n29020 | n29021 ;
  assign n29023 = n29019 | n29022 ;
  assign n29024 = n4051 & ~n23691 ;
  assign n29025 = ~n23695 & n29024 ;
  assign n29026 = ( n4051 & n29023 ) | ( n4051 & ~n29025 ) | ( n29023 & ~n29025 ) ;
  assign n29027 = ~x29 & n29026 ;
  assign n29028 = x29 | n29027 ;
  assign n29029 = ( ~n29026 & n29027 ) | ( ~n29026 & n29028 ) | ( n29027 & n29028 ) ;
  assign n29030 = ~n29018 & n29029 ;
  assign n29031 = n29018 & ~n29029 ;
  assign n29032 = n29030 | n29031 ;
  assign n29033 = ~n28929 & n29032 ;
  assign n29034 = ~n28932 & n29033 ;
  assign n29035 = ( n28929 & n28932 ) | ( n28929 & ~n29032 ) | ( n28932 & ~n29032 ) ;
  assign n29036 = n29034 | n29035 ;
  assign n29037 = n4484 & ~n24334 ;
  assign n29038 = n4479 & ~n21005 ;
  assign n29039 = n4481 & n24329 ;
  assign n29040 = n29038 | n29039 ;
  assign n29041 = n29037 | n29040 ;
  assign n29042 = ( n4487 & ~n24373 ) | ( n4487 & n24376 ) | ( ~n24373 & n24376 ) ;
  assign n29043 = n29041 | n29042 ;
  assign n29044 = x26 | n29043 ;
  assign n29045 = ~x26 & n29044 ;
  assign n29046 = ( ~n29043 & n29044 ) | ( ~n29043 & n29045 ) | ( n29044 & n29045 ) ;
  assign n29047 = n29036 | n29046 ;
  assign n29048 = ~n29046 & n29047 ;
  assign n29049 = ( ~n29036 & n29047 ) | ( ~n29036 & n29048 ) | ( n29047 & n29048 ) ;
  assign n29050 = ( n28840 & n28934 ) | ( n28840 & n28944 ) | ( n28934 & n28944 ) ;
  assign n29051 = ~n29049 & n29050 ;
  assign n29052 = n29049 | n29051 ;
  assign n29053 = n29050 & ~n29051 ;
  assign n29054 = n29052 & ~n29053 ;
  assign n29055 = n4551 & n25442 ;
  assign n29056 = n4546 & n24324 ;
  assign n29057 = n4548 & n25187 ;
  assign n29058 = n29056 | n29057 ;
  assign n29059 = n29055 | n29058 ;
  assign n29060 = n4554 | n29059 ;
  assign n29061 = ( n25452 & n29059 ) | ( n25452 & n29060 ) | ( n29059 & n29060 ) ;
  assign n29062 = x23 & n29061 ;
  assign n29063 = x23 & ~n29062 ;
  assign n29064 = ( n29061 & ~n29062 ) | ( n29061 & n29063 ) | ( ~n29062 & n29063 ) ;
  assign n29065 = ( n28985 & n29054 ) | ( n28985 & ~n29064 ) | ( n29054 & ~n29064 ) ;
  assign n29066 = ( ~n29054 & n29064 ) | ( ~n29054 & n29065 ) | ( n29064 & n29065 ) ;
  assign n29067 = ( ~n28985 & n29065 ) | ( ~n28985 & n29066 ) | ( n29065 & n29066 ) ;
  assign n29068 = n4781 & n26156 ;
  assign n29069 = n4776 & ~n25676 ;
  assign n29070 = n4778 & n25928 ;
  assign n29071 = n29069 | n29070 ;
  assign n29072 = n29068 | n29071 ;
  assign n29073 = n4784 | n29072 ;
  assign n29074 = ( n26167 & n29072 ) | ( n26167 & n29073 ) | ( n29072 & n29073 ) ;
  assign n29075 = x20 & n29074 ;
  assign n29076 = x20 & ~n29075 ;
  assign n29077 = ( n29074 & ~n29075 ) | ( n29074 & n29076 ) | ( ~n29075 & n29076 ) ;
  assign n29078 = n29067 | n29077 ;
  assign n29079 = ~n29077 & n29078 ;
  assign n29080 = ( ~n29067 & n29078 ) | ( ~n29067 & n29079 ) | ( n29078 & n29079 ) ;
  assign n29081 = n28878 | n28967 ;
  assign n29082 = ~n29080 & n29081 ;
  assign n29083 = n29080 | n29082 ;
  assign n29084 = n29081 & ~n29082 ;
  assign n29085 = n29083 & ~n29084 ;
  assign n29086 = n28970 | n28974 ;
  assign n29087 = ~n29085 & n29086 ;
  assign n29088 = n28970 | n28976 ;
  assign n29089 = ~n29085 & n29088 ;
  assign n29090 = ( n28314 & n29087 ) | ( n28314 & n29089 ) | ( n29087 & n29089 ) ;
  assign n29091 = ( n28314 & n29086 ) | ( n28314 & n29088 ) | ( n29086 & n29088 ) ;
  assign n29092 = n29085 & ~n29091 ;
  assign n29093 = n29090 | n29092 ;
  assign n29094 = n28983 | n29093 ;
  assign n29095 = n28983 & n29093 ;
  assign n29096 = n29094 & ~n29095 ;
  assign n29097 = n4484 & n24324 ;
  assign n29098 = n4479 & n24329 ;
  assign n29099 = n4481 & ~n24334 ;
  assign n29100 = n29098 | n29099 ;
  assign n29101 = n29097 | n29100 ;
  assign n29102 = n4487 & ~n24353 ;
  assign n29103 = ( n4487 & n24356 ) | ( n4487 & n29102 ) | ( n24356 & n29102 ) ;
  assign n29104 = n29101 | n29103 ;
  assign n29105 = x26 | n29104 ;
  assign n29106 = ~x26 & n29105 ;
  assign n29107 = ( ~n29104 & n29105 ) | ( ~n29104 & n29106 ) | ( n29105 & n29106 ) ;
  assign n29108 = n4048 & ~n21005 ;
  assign n29109 = n4043 & n20838 ;
  assign n29110 = n4045 & n20921 ;
  assign n29111 = n29109 | n29110 ;
  assign n29112 = n29108 | n29111 ;
  assign n29113 = n4051 | n29112 ;
  assign n29114 = ( ~n21015 & n29112 ) | ( ~n21015 & n29113 ) | ( n29112 & n29113 ) ;
  assign n29115 = ~x29 & n29114 ;
  assign n29116 = x29 | n29115 ;
  assign n29117 = ( ~n29114 & n29115 ) | ( ~n29114 & n29116 ) | ( n29115 & n29116 ) ;
  assign n29118 = n3744 & n20532 ;
  assign n29119 = n3639 & ~n20724 ;
  assign n29120 = n3727 & ~n20536 ;
  assign n29121 = n29119 | n29120 ;
  assign n29122 = n29118 | n29121 ;
  assign n29123 = n3636 | n29122 ;
  assign n29124 = ( n23203 & n29122 ) | ( n23203 & n29123 ) | ( n29122 & n29123 ) ;
  assign n29125 = n19814 | n28780 ;
  assign n29126 = n4012 & ~n29125 ;
  assign n29127 = ~n11526 & n29126 ;
  assign n29128 = ~n5818 & n29127 ;
  assign n29129 = n869 | n2642 ;
  assign n29130 = n3224 | n29129 ;
  assign n29131 = n29128 & ~n29130 ;
  assign n29132 = n3293 | n26671 ;
  assign n29133 = n29131 & ~n29132 ;
  assign n29134 = n283 | n499 ;
  assign n29135 = n590 | n29134 ;
  assign n29136 = n139 | n29135 ;
  assign n29137 = n29133 & ~n29136 ;
  assign n29138 = ~n29008 & n29137 ;
  assign n29139 = n29008 & ~n29137 ;
  assign n29140 = n29123 & ~n29139 ;
  assign n29141 = ~n29138 & n29140 ;
  assign n29142 = n29122 & ~n29139 ;
  assign n29143 = ~n29138 & n29142 ;
  assign n29144 = ( n23203 & n29141 ) | ( n23203 & n29143 ) | ( n29141 & n29143 ) ;
  assign n29145 = n29124 & ~n29144 ;
  assign n29146 = ( n28992 & n29012 ) | ( n28992 & ~n29015 ) | ( n29012 & ~n29015 ) ;
  assign n29147 = n29009 | n29146 ;
  assign n29148 = n29139 | n29144 ;
  assign n29149 = n29138 | n29148 ;
  assign n29150 = n29147 & ~n29149 ;
  assign n29151 = ( n29145 & n29147 ) | ( n29145 & n29150 ) | ( n29147 & n29150 ) ;
  assign n29152 = ~n29147 & n29149 ;
  assign n29153 = ~n29145 & n29152 ;
  assign n29154 = n29151 | n29153 ;
  assign n29155 = n29017 | n29030 ;
  assign n29156 = n29154 & ~n29155 ;
  assign n29157 = ~n29154 & n29155 ;
  assign n29158 = n29156 | n29157 ;
  assign n29159 = n29117 & ~n29158 ;
  assign n29160 = n29158 | n29159 ;
  assign n29161 = ( ~n29117 & n29159 ) | ( ~n29117 & n29160 ) | ( n29159 & n29160 ) ;
  assign n29162 = n29107 & ~n29161 ;
  assign n29163 = ~n29107 & n29161 ;
  assign n29164 = n29162 | n29163 ;
  assign n29165 = ( n29035 & n29046 ) | ( n29035 & n29049 ) | ( n29046 & n29049 ) ;
  assign n29166 = n29164 & ~n29165 ;
  assign n29167 = ~n29164 & n29165 ;
  assign n29168 = n29166 | n29167 ;
  assign n29169 = n4551 & ~n25676 ;
  assign n29170 = n4546 & n25187 ;
  assign n29171 = n4548 & n25442 ;
  assign n29172 = n29170 | n29171 ;
  assign n29173 = n29169 | n29172 ;
  assign n29174 = n4554 & ~n25690 ;
  assign n29175 = ( n4554 & n25694 ) | ( n4554 & n29174 ) | ( n25694 & n29174 ) ;
  assign n29176 = n29173 | n29175 ;
  assign n29177 = x23 | n29176 ;
  assign n29178 = ~x23 & n29177 ;
  assign n29179 = ( ~n29176 & n29177 ) | ( ~n29176 & n29178 ) | ( n29177 & n29178 ) ;
  assign n29180 = n29168 & n29179 ;
  assign n29181 = ( ~n29164 & n29165 ) | ( ~n29164 & n29179 ) | ( n29165 & n29179 ) ;
  assign n29182 = n29166 | n29181 ;
  assign n29183 = ~n29180 & n29182 ;
  assign n29184 = n20032 & n26156 ;
  assign n29185 = n4776 & n25928 ;
  assign n29186 = n29184 | n29185 ;
  assign n29187 = n4784 | n29186 ;
  assign n29188 = ( n26165 & n29186 ) | ( n26165 & n29187 ) | ( n29186 & n29187 ) ;
  assign n29189 = x20 & n29188 ;
  assign n29190 = x20 & ~n29189 ;
  assign n29191 = ( n29188 & ~n29189 ) | ( n29188 & n29190 ) | ( ~n29189 & n29190 ) ;
  assign n29192 = ( ~n29049 & n29050 ) | ( ~n29049 & n29064 ) | ( n29050 & n29064 ) ;
  assign n29193 = n29191 & n29192 ;
  assign n29194 = n29191 | n29192 ;
  assign n29195 = ~n29193 & n29194 ;
  assign n29196 = ~n29183 & n29195 ;
  assign n29197 = n29183 | n29196 ;
  assign n29198 = n29195 & ~n29196 ;
  assign n29199 = n29197 & ~n29198 ;
  assign n29200 = ( n28985 & n29077 ) | ( n28985 & n29080 ) | ( n29077 & n29080 ) ;
  assign n29201 = n29199 & ~n29200 ;
  assign n29202 = ~n29199 & n29200 ;
  assign n29203 = n29201 | n29202 ;
  assign n29204 = n29082 | n29087 ;
  assign n29205 = ~n29203 & n29204 ;
  assign n29206 = n29082 | n29089 ;
  assign n29207 = ~n29203 & n29206 ;
  assign n29208 = ( n28314 & n29205 ) | ( n28314 & n29207 ) | ( n29205 & n29207 ) ;
  assign n29209 = ( n28314 & n29204 ) | ( n28314 & n29206 ) | ( n29204 & n29206 ) ;
  assign n29210 = n29203 & ~n29209 ;
  assign n29211 = n29208 | n29210 ;
  assign n29212 = ( n28983 & ~n29093 ) | ( n28983 & n29096 ) | ( ~n29093 & n29096 ) ;
  assign n29213 = ~n29211 & n29212 ;
  assign n29214 = n29211 & ~n29212 ;
  assign n29215 = n29213 | n29214 ;
  assign n29216 = n29193 | n29196 ;
  assign n29217 = n4551 & n25928 ;
  assign n29218 = n4546 & n25442 ;
  assign n29219 = n4548 & ~n25676 ;
  assign n29220 = n29218 | n29219 ;
  assign n29221 = n29217 | n29220 ;
  assign n29222 = n4554 | n29221 ;
  assign n29223 = ( ~n25936 & n29221 ) | ( ~n25936 & n29222 ) | ( n29221 & n29222 ) ;
  assign n29224 = ~x23 & n29223 ;
  assign n29225 = x23 | n29224 ;
  assign n29226 = ( ~n29223 & n29224 ) | ( ~n29223 & n29225 ) | ( n29224 & n29225 ) ;
  assign n29227 = n29181 & n29226 ;
  assign n29228 = n29181 & ~n29227 ;
  assign n29229 = n29159 | n29162 ;
  assign n29230 = n4484 & n25187 ;
  assign n29231 = n4479 & ~n24334 ;
  assign n29232 = n4481 & n24324 ;
  assign n29233 = n29231 | n29232 ;
  assign n29234 = n29230 | n29233 ;
  assign n29235 = n4487 | n29234 ;
  assign n29236 = ( n25193 & n29234 ) | ( n25193 & n29235 ) | ( n29234 & n29235 ) ;
  assign n29237 = x26 & n29236 ;
  assign n29238 = x26 & ~n29237 ;
  assign n29239 = ( n29236 & ~n29237 ) | ( n29236 & n29238 ) | ( ~n29237 & n29238 ) ;
  assign n29240 = n4048 & n24329 ;
  assign n29241 = n4043 & n20921 ;
  assign n29242 = n4045 & ~n21005 ;
  assign n29243 = n29241 | n29242 ;
  assign n29244 = n29240 | n29243 ;
  assign n29245 = ( n4051 & ~n24391 ) | ( n4051 & n24392 ) | ( ~n24391 & n24392 ) ;
  assign n29246 = n29244 | n29245 ;
  assign n29247 = x29 | n29246 ;
  assign n29248 = ~x29 & n29247 ;
  assign n29249 = ( ~n29246 & n29247 ) | ( ~n29246 & n29248 ) | ( n29247 & n29248 ) ;
  assign n29250 = n3744 & n20838 ;
  assign n29251 = n3639 & ~n20536 ;
  assign n29252 = n3727 & n20532 ;
  assign n29253 = n29251 | n29252 ;
  assign n29254 = n29250 | n29253 ;
  assign n29255 = n3636 | n29254 ;
  assign n29256 = ( ~n23712 & n29254 ) | ( ~n23712 & n29255 ) | ( n29254 & n29255 ) ;
  assign n29257 = n2733 | n3577 ;
  assign n29258 = n873 | n29257 ;
  assign n29259 = n12991 | n29258 ;
  assign n29260 = ( n3833 & n14065 ) | ( n3833 & ~n29259 ) | ( n14065 & ~n29259 ) ;
  assign n29261 = ~n3833 & n29260 ;
  assign n29262 = ~n3072 & n29261 ;
  assign n29263 = n216 | n1045 ;
  assign n29264 = n2385 | n29263 ;
  assign n29265 = n857 | n29264 ;
  assign n29266 = n759 | n29265 ;
  assign n29267 = n514 | n29266 ;
  assign n29268 = n335 | n29267 ;
  assign n29269 = n504 | n29268 ;
  assign n29270 = n29262 & ~n29269 ;
  assign n29271 = n592 | n610 ;
  assign n29272 = n92 | n29271 ;
  assign n29273 = n29270 & ~n29272 ;
  assign n29274 = n29008 & n29273 ;
  assign n29275 = n29008 | n29273 ;
  assign n29276 = ~n29274 & n29275 ;
  assign n29277 = n20034 & n26156 ;
  assign n29278 = ~x20 & n29277 ;
  assign n29279 = x20 | n29278 ;
  assign n29280 = ( ~n29277 & n29278 ) | ( ~n29277 & n29279 ) | ( n29278 & n29279 ) ;
  assign n29281 = n29276 & ~n29280 ;
  assign n29282 = ~n29276 & n29280 ;
  assign n29283 = n29281 | n29282 ;
  assign n29284 = ( n29148 & n29256 ) | ( n29148 & ~n29283 ) | ( n29256 & ~n29283 ) ;
  assign n29285 = ( ~n29148 & n29283 ) | ( ~n29148 & n29284 ) | ( n29283 & n29284 ) ;
  assign n29286 = ( ~n29256 & n29284 ) | ( ~n29256 & n29285 ) | ( n29284 & n29285 ) ;
  assign n29287 = ( n29151 & n29157 ) | ( n29151 & ~n29286 ) | ( n29157 & ~n29286 ) ;
  assign n29288 = ( n29151 & ~n29153 ) | ( n29151 & n29155 ) | ( ~n29153 & n29155 ) ;
  assign n29289 = n29286 & ~n29288 ;
  assign n29290 = n29287 | n29289 ;
  assign n29291 = n29249 & ~n29290 ;
  assign n29292 = n29290 | n29291 ;
  assign n29293 = ( ~n29249 & n29291 ) | ( ~n29249 & n29292 ) | ( n29291 & n29292 ) ;
  assign n29294 = n29239 & ~n29293 ;
  assign n29295 = ~n29239 & n29293 ;
  assign n29296 = n29294 | n29295 ;
  assign n29297 = ~n29229 & n29296 ;
  assign n29298 = n29229 & ~n29296 ;
  assign n29299 = n29297 | n29298 ;
  assign n29300 = ~n29181 & n29226 ;
  assign n29301 = n29299 & ~n29300 ;
  assign n29302 = ~n29228 & n29301 ;
  assign n29303 = ( n29228 & ~n29299 ) | ( n29228 & n29300 ) | ( ~n29299 & n29300 ) ;
  assign n29304 = n29302 | n29303 ;
  assign n29305 = n29216 & ~n29304 ;
  assign n29306 = ~n29216 & n29304 ;
  assign n29307 = n29305 | n29306 ;
  assign n29308 = n29202 | n29205 ;
  assign n29309 = ~n29307 & n29308 ;
  assign n29310 = n29202 | n29207 ;
  assign n29311 = ~n29307 & n29310 ;
  assign n29312 = ( n28314 & n29309 ) | ( n28314 & n29311 ) | ( n29309 & n29311 ) ;
  assign n29313 = ( n28314 & n29308 ) | ( n28314 & n29310 ) | ( n29308 & n29310 ) ;
  assign n29314 = n29307 & ~n29313 ;
  assign n29315 = n29312 | n29314 ;
  assign n29316 = ~n29213 & n29315 ;
  assign n29317 = n29211 | n29315 ;
  assign n29318 = n29212 & ~n29317 ;
  assign n29319 = n29316 | n29318 ;
  assign n29320 = n29227 | n29303 ;
  assign n29321 = n4551 & n26156 ;
  assign n29322 = n4546 & ~n25676 ;
  assign n29323 = n4548 & n25928 ;
  assign n29324 = n29322 | n29323 ;
  assign n29325 = n29321 | n29324 ;
  assign n29326 = n4554 | n29325 ;
  assign n29327 = ( n26167 & n29325 ) | ( n26167 & n29326 ) | ( n29325 & n29326 ) ;
  assign n29328 = x23 & n29327 ;
  assign n29329 = x23 & ~n29328 ;
  assign n29330 = ( n29327 & ~n29328 ) | ( n29327 & n29329 ) | ( ~n29328 & n29329 ) ;
  assign n29331 = n29294 | n29298 ;
  assign n29332 = n29287 | n29291 ;
  assign n29333 = n3744 & n20921 ;
  assign n29334 = n3639 & n20532 ;
  assign n29335 = n3727 & n20838 ;
  assign n29336 = n29334 | n29335 ;
  assign n29337 = n29333 | n29336 ;
  assign n29338 = ( n3636 & n23691 ) | ( n3636 & n23695 ) | ( n23691 & n23695 ) ;
  assign n29339 = n29337 | n29338 ;
  assign n29340 = n1654 | n11288 ;
  assign n29341 = n13976 | n29340 ;
  assign n29342 = n1682 | n3903 ;
  assign n29343 = n1576 | n29342 ;
  assign n29344 = n1605 | n29343 ;
  assign n29345 = n890 | n29344 ;
  assign n29346 = ( ~n11538 & n12657 ) | ( ~n11538 & n29345 ) | ( n12657 & n29345 ) ;
  assign n29347 = n11538 | n29346 ;
  assign n29348 = n29341 | n29347 ;
  assign n29349 = n431 | n1417 ;
  assign n29350 = n499 | n29349 ;
  assign n29351 = n198 | n29350 ;
  assign n29352 = n203 | n29351 ;
  assign n29353 = n646 | n29352 ;
  assign n29354 = n29348 | n29353 ;
  assign n29355 = ( n29275 & ~n29281 ) | ( n29275 & n29354 ) | ( ~n29281 & n29354 ) ;
  assign n29356 = ( n29274 & n29275 ) | ( n29274 & n29280 ) | ( n29275 & n29280 ) ;
  assign n29357 = n29354 & n29356 ;
  assign n29358 = n29355 & ~n29357 ;
  assign n29359 = n29339 | n29358 ;
  assign n29360 = ~n29358 & n29359 ;
  assign n29361 = ( ~n29339 & n29359 ) | ( ~n29339 & n29360 ) | ( n29359 & n29360 ) ;
  assign n29362 = n29284 | n29361 ;
  assign n29363 = n29284 & n29361 ;
  assign n29364 = n29362 & ~n29363 ;
  assign n29365 = n4048 & ~n24334 ;
  assign n29366 = n4043 & ~n21005 ;
  assign n29367 = n4045 & n24329 ;
  assign n29368 = n29366 | n29367 ;
  assign n29369 = n29365 | n29368 ;
  assign n29370 = n4051 & ~n24376 ;
  assign n29371 = n24373 & n29370 ;
  assign n29372 = ( n4051 & n29369 ) | ( n4051 & ~n29371 ) | ( n29369 & ~n29371 ) ;
  assign n29373 = x29 & n29372 ;
  assign n29374 = x29 & ~n29373 ;
  assign n29375 = ( n29372 & ~n29373 ) | ( n29372 & n29374 ) | ( ~n29373 & n29374 ) ;
  assign n29376 = n29364 & n29375 ;
  assign n29377 = n29364 | n29375 ;
  assign n29378 = ~n29376 & n29377 ;
  assign n29379 = n4484 & n25442 ;
  assign n29380 = n4479 & n24324 ;
  assign n29381 = n4481 & n25187 ;
  assign n29382 = n29380 | n29381 ;
  assign n29383 = n29379 | n29382 ;
  assign n29384 = n4487 | n29383 ;
  assign n29385 = ( n25452 & n29383 ) | ( n25452 & n29384 ) | ( n29383 & n29384 ) ;
  assign n29386 = x26 & n29385 ;
  assign n29387 = x26 & ~n29386 ;
  assign n29388 = ( n29385 & ~n29386 ) | ( n29385 & n29387 ) | ( ~n29386 & n29387 ) ;
  assign n29389 = ( n29332 & n29378 ) | ( n29332 & n29388 ) | ( n29378 & n29388 ) ;
  assign n29390 = ( n29378 & n29388 ) | ( n29378 & ~n29389 ) | ( n29388 & ~n29389 ) ;
  assign n29391 = ( n29332 & ~n29389 ) | ( n29332 & n29390 ) | ( ~n29389 & n29390 ) ;
  assign n29392 = ( n29330 & ~n29331 ) | ( n29330 & n29391 ) | ( ~n29331 & n29391 ) ;
  assign n29393 = ( n29331 & ~n29391 ) | ( n29331 & n29392 ) | ( ~n29391 & n29392 ) ;
  assign n29394 = ( ~n29330 & n29392 ) | ( ~n29330 & n29393 ) | ( n29392 & n29393 ) ;
  assign n29395 = n29320 & n29394 ;
  assign n29396 = n29320 & ~n29395 ;
  assign n29397 = ~n29320 & n29394 ;
  assign n29398 = n29396 | n29397 ;
  assign n29399 = n29305 | n29309 ;
  assign n29400 = n29398 & n29399 ;
  assign n29401 = n29305 | n29311 ;
  assign n29402 = n29398 & n29401 ;
  assign n29403 = ( n28314 & n29400 ) | ( n28314 & n29402 ) | ( n29400 & n29402 ) ;
  assign n29404 = ( n28314 & n29399 ) | ( n28314 & n29401 ) | ( n29399 & n29401 ) ;
  assign n29405 = n29398 | n29404 ;
  assign n29406 = ~n29403 & n29405 ;
  assign n29407 = n29318 & ~n29406 ;
  assign n29408 = ~n29318 & n29406 ;
  assign n29409 = n29407 | n29408 ;
  assign n29410 = ( n29330 & n29331 ) | ( n29330 & n29391 ) | ( n29331 & n29391 ) ;
  assign n29411 = n4484 & ~n25676 ;
  assign n29412 = n4479 & n25187 ;
  assign n29413 = n4481 & n25442 ;
  assign n29414 = n29412 | n29413 ;
  assign n29415 = n29411 | n29414 ;
  assign n29416 = n4487 & ~n25690 ;
  assign n29417 = ( n4487 & n25694 ) | ( n4487 & n29416 ) | ( n25694 & n29416 ) ;
  assign n29418 = n29415 | n29417 ;
  assign n29419 = x26 | n29418 ;
  assign n29420 = ~x26 & n29419 ;
  assign n29421 = ( ~n29418 & n29419 ) | ( ~n29418 & n29420 ) | ( n29419 & n29420 ) ;
  assign n29422 = n4048 & n24324 ;
  assign n29423 = n4043 & n24329 ;
  assign n29424 = n4045 & ~n24334 ;
  assign n29425 = n29423 | n29424 ;
  assign n29426 = n29422 | n29425 ;
  assign n29427 = n4051 & ~n24353 ;
  assign n29428 = ( n4051 & n24356 ) | ( n4051 & n29427 ) | ( n24356 & n29427 ) ;
  assign n29429 = n29426 | n29428 ;
  assign n29430 = x29 | n29429 ;
  assign n29431 = ~x29 & n29430 ;
  assign n29432 = ( ~n29429 & n29430 ) | ( ~n29429 & n29431 ) | ( n29430 & n29431 ) ;
  assign n29433 = ( ~n29337 & n29355 ) | ( ~n29337 & n29357 ) | ( n29355 & n29357 ) ;
  assign n29434 = ( ~n29338 & n29357 ) | ( ~n29338 & n29433 ) | ( n29357 & n29433 ) ;
  assign n29435 = n869 | n27378 ;
  assign n29436 = n1443 | n29435 ;
  assign n29437 = n1417 | n29436 ;
  assign n29438 = n127 | n29437 ;
  assign n29439 = n892 | n3152 ;
  assign n29440 = n12244 | n29439 ;
  assign n29441 = n13880 | n29440 ;
  assign n29442 = ( ~n4683 & n20952 ) | ( ~n4683 & n29441 ) | ( n20952 & n29441 ) ;
  assign n29443 = n4683 | n29442 ;
  assign n29444 = n29438 | n29443 ;
  assign n29445 = n21236 & ~n21242 ;
  assign n29446 = ~n280 & n29445 ;
  assign n29447 = ~n270 & n29446 ;
  assign n29448 = ~n29444 & n29447 ;
  assign n29449 = n193 | n417 ;
  assign n29450 = n29448 & ~n29449 ;
  assign n29451 = n29354 | n29450 ;
  assign n29452 = n29354 & n29450 ;
  assign n29453 = n29433 | n29452 ;
  assign n29454 = n29451 & ~n29453 ;
  assign n29455 = n29357 | n29452 ;
  assign n29456 = n29451 & ~n29455 ;
  assign n29457 = ( n29338 & n29454 ) | ( n29338 & n29456 ) | ( n29454 & n29456 ) ;
  assign n29458 = n29434 | n29457 ;
  assign n29459 = n29452 | n29457 ;
  assign n29460 = n29451 & ~n29459 ;
  assign n29461 = n29458 & ~n29460 ;
  assign n29462 = n3744 & ~n21005 ;
  assign n29463 = n3639 & n20838 ;
  assign n29464 = n3727 & n20921 ;
  assign n29465 = n29463 | n29464 ;
  assign n29466 = n29462 | n29465 ;
  assign n29467 = n3636 | n29466 ;
  assign n29468 = ( ~n21015 & n29466 ) | ( ~n21015 & n29467 ) | ( n29466 & n29467 ) ;
  assign n29469 = ~n29461 & n29468 ;
  assign n29470 = n29461 & ~n29468 ;
  assign n29471 = n29469 | n29470 ;
  assign n29472 = n29363 | n29376 ;
  assign n29473 = n29471 & ~n29472 ;
  assign n29474 = ~n29471 & n29472 ;
  assign n29475 = n29473 | n29474 ;
  assign n29476 = n29432 & ~n29475 ;
  assign n29477 = n29475 | n29476 ;
  assign n29478 = ( ~n29432 & n29476 ) | ( ~n29432 & n29477 ) | ( n29476 & n29477 ) ;
  assign n29479 = n29421 & ~n29478 ;
  assign n29480 = ~n29421 & n29478 ;
  assign n29481 = n29479 | n29480 ;
  assign n29482 = n20737 & n26156 ;
  assign n29483 = n4546 & n25928 ;
  assign n29484 = n29482 | n29483 ;
  assign n29485 = n4554 | n29484 ;
  assign n29486 = ( n26165 & n29484 ) | ( n26165 & n29485 ) | ( n29484 & n29485 ) ;
  assign n29487 = x23 & n29486 ;
  assign n29488 = x23 & ~n29487 ;
  assign n29489 = ( n29486 & ~n29487 ) | ( n29486 & n29488 ) | ( ~n29487 & n29488 ) ;
  assign n29490 = n29389 & n29489 ;
  assign n29491 = n29389 | n29489 ;
  assign n29492 = ~n29490 & n29491 ;
  assign n29493 = ~n29481 & n29492 ;
  assign n29494 = n29481 | n29493 ;
  assign n29495 = n29492 & ~n29493 ;
  assign n29496 = n29494 & ~n29495 ;
  assign n29497 = ~n29410 & n29496 ;
  assign n29498 = n29410 & ~n29496 ;
  assign n29499 = n29497 | n29498 ;
  assign n29500 = n29395 | n29400 ;
  assign n29501 = ~n29499 & n29500 ;
  assign n29502 = n29395 | n29402 ;
  assign n29503 = ~n29499 & n29502 ;
  assign n29504 = ( n28314 & n29501 ) | ( n28314 & n29503 ) | ( n29501 & n29503 ) ;
  assign n29505 = ( n28314 & n29500 ) | ( n28314 & n29502 ) | ( n29500 & n29502 ) ;
  assign n29506 = n29499 & ~n29505 ;
  assign n29507 = n29504 | n29506 ;
  assign n29508 = ~n29317 & n29406 ;
  assign n29509 = n29212 & n29508 ;
  assign n29510 = n29507 & ~n29509 ;
  assign n29511 = ~n29507 & n29508 ;
  assign n29512 = n29212 & n29511 ;
  assign n29513 = n29510 | n29512 ;
  assign n29514 = n29490 | n29493 ;
  assign n29515 = n4484 & n25928 ;
  assign n29516 = n4479 & n25442 ;
  assign n29517 = n4481 & ~n25676 ;
  assign n29518 = n29516 | n29517 ;
  assign n29519 = n29515 | n29518 ;
  assign n29520 = n4487 | n29519 ;
  assign n29521 = ( ~n25936 & n29519 ) | ( ~n25936 & n29520 ) | ( n29519 & n29520 ) ;
  assign n29522 = ~x26 & n29521 ;
  assign n29523 = x26 | n29522 ;
  assign n29524 = ( ~n29521 & n29522 ) | ( ~n29521 & n29523 ) | ( n29522 & n29523 ) ;
  assign n29525 = n29476 | n29479 ;
  assign n29526 = n644 | n657 ;
  assign n29527 = n3710 | n3866 ;
  assign n29528 = n115 | n29527 ;
  assign n29529 = n332 & ~n29528 ;
  assign n29530 = ~n29526 & n29529 ;
  assign n29531 = ~n3406 & n29530 ;
  assign n29532 = ( n348 & n960 ) | ( n348 & ~n13871 ) | ( n960 & ~n13871 ) ;
  assign n29533 = n13871 | n29532 ;
  assign n29534 = n429 | n29533 ;
  assign n29535 = n373 | n29534 ;
  assign n29536 = n351 | n29535 ;
  assign n29537 = n366 | n29536 ;
  assign n29538 = n591 | n29537 ;
  assign n29539 = n29531 & ~n29538 ;
  assign n29540 = ~n161 & n29539 ;
  assign n29541 = n29450 & n29540 ;
  assign n29542 = n29450 | n29540 ;
  assign n29543 = ~n29541 & n29542 ;
  assign n29544 = n20871 & n26156 ;
  assign n29545 = ~x23 & n29544 ;
  assign n29546 = x23 | n29545 ;
  assign n29547 = ( ~n29544 & n29545 ) | ( ~n29544 & n29546 ) | ( n29545 & n29546 ) ;
  assign n29548 = n29543 & ~n29547 ;
  assign n29549 = ~n29543 & n29547 ;
  assign n29550 = n29548 | n29549 ;
  assign n29551 = n29459 & ~n29550 ;
  assign n29552 = ~n29459 & n29550 ;
  assign n29553 = n29551 | n29552 ;
  assign n29554 = n3744 & n24329 ;
  assign n29555 = n3639 & n20921 ;
  assign n29556 = n3727 & ~n21005 ;
  assign n29557 = n29555 | n29556 ;
  assign n29558 = n29554 | n29557 ;
  assign n29559 = ( n3636 & ~n24391 ) | ( n3636 & n24392 ) | ( ~n24391 & n24392 ) ;
  assign n29560 = n29558 | n29559 ;
  assign n29561 = ~n29553 & n29560 ;
  assign n29562 = n29553 | n29561 ;
  assign n29563 = n29560 & ~n29561 ;
  assign n29564 = n29562 & ~n29563 ;
  assign n29565 = n29469 | n29474 ;
  assign n29566 = n29564 & ~n29565 ;
  assign n29567 = ~n29564 & n29565 ;
  assign n29568 = n29566 | n29567 ;
  assign n29569 = n4048 & n25187 ;
  assign n29570 = n4043 & ~n24334 ;
  assign n29571 = n4045 & n24324 ;
  assign n29572 = n29570 | n29571 ;
  assign n29573 = n29569 | n29572 ;
  assign n29574 = n4051 | n29573 ;
  assign n29575 = ( n25193 & n29573 ) | ( n25193 & n29574 ) | ( n29573 & n29574 ) ;
  assign n29576 = x29 & n29575 ;
  assign n29577 = x29 & ~n29576 ;
  assign n29578 = ( n29575 & ~n29576 ) | ( n29575 & n29577 ) | ( ~n29576 & n29577 ) ;
  assign n29579 = n29568 & n29578 ;
  assign n29580 = ( ~n29564 & n29565 ) | ( ~n29564 & n29578 ) | ( n29565 & n29578 ) ;
  assign n29581 = n29566 | n29580 ;
  assign n29582 = ~n29579 & n29581 ;
  assign n29583 = ( n29524 & ~n29525 ) | ( n29524 & n29582 ) | ( ~n29525 & n29582 ) ;
  assign n29584 = ( n29525 & ~n29582 ) | ( n29525 & n29583 ) | ( ~n29582 & n29583 ) ;
  assign n29585 = ( ~n29524 & n29583 ) | ( ~n29524 & n29584 ) | ( n29583 & n29584 ) ;
  assign n29586 = n29514 & ~n29585 ;
  assign n29587 = ~n29514 & n29585 ;
  assign n29588 = n29586 | n29587 ;
  assign n29589 = n29498 | n29501 ;
  assign n29590 = n29498 | n29503 ;
  assign n29591 = ( n28314 & n29589 ) | ( n28314 & n29590 ) | ( n29589 & n29590 ) ;
  assign n29592 = n29588 & ~n29591 ;
  assign n29593 = ~n29588 & n29591 ;
  assign n29594 = n29592 | n29593 ;
  assign n29595 = ~n29512 & n29594 ;
  assign n29596 = ( n29512 & ~n29594 ) | ( n29512 & n29595 ) | ( ~n29594 & n29595 ) ;
  assign n29597 = n29595 | n29596 ;
  assign n29598 = n29586 | n29593 ;
  assign n29599 = n4484 & n26156 ;
  assign n29600 = n4479 & ~n25676 ;
  assign n29601 = n4481 & n25928 ;
  assign n29602 = n29600 | n29601 ;
  assign n29603 = n29599 | n29602 ;
  assign n29604 = n4487 | n29603 ;
  assign n29605 = ( n26167 & n29603 ) | ( n26167 & n29604 ) | ( n29603 & n29604 ) ;
  assign n29606 = x26 & n29605 ;
  assign n29607 = x26 & ~n29606 ;
  assign n29608 = ( n29605 & ~n29606 ) | ( n29605 & n29607 ) | ( ~n29606 & n29607 ) ;
  assign n29609 = n29551 | n29561 ;
  assign n29610 = n3744 & ~n24334 ;
  assign n29611 = n3639 & ~n21005 ;
  assign n29612 = n3727 & n24329 ;
  assign n29613 = n29611 | n29612 ;
  assign n29614 = n29610 | n29613 ;
  assign n29615 = ( n3636 & ~n24373 ) | ( n3636 & n24376 ) | ( ~n24373 & n24376 ) ;
  assign n29616 = n29614 | n29615 ;
  assign n29617 = n1680 | n3532 ;
  assign n29618 = n12958 | n29617 ;
  assign n29619 = n5550 | n29618 ;
  assign n29620 = n24163 | n29619 ;
  assign n29621 = n665 | n29620 ;
  assign n29622 = n3418 | n29621 ;
  assign n29623 = n13877 | n29622 ;
  assign n29624 = n324 | n1337 ;
  assign n29625 = n130 | n29624 ;
  assign n29626 = n2922 | n29625 ;
  assign n29627 = n339 | n29626 ;
  assign n29628 = n3243 | n29627 ;
  assign n29629 = n29623 | n29628 ;
  assign n29630 = n199 | n335 ;
  assign n29631 = n203 | n29630 ;
  assign n29632 = n126 | n29631 ;
  assign n29633 = n29629 | n29632 ;
  assign n29634 = ( n29542 & ~n29548 ) | ( n29542 & n29633 ) | ( ~n29548 & n29633 ) ;
  assign n29635 = ( n29541 & n29542 ) | ( n29541 & n29547 ) | ( n29542 & n29547 ) ;
  assign n29636 = n29633 & n29635 ;
  assign n29637 = n29634 & ~n29636 ;
  assign n29638 = n29616 | n29637 ;
  assign n29639 = ~n29637 & n29638 ;
  assign n29640 = ( ~n29616 & n29638 ) | ( ~n29616 & n29639 ) | ( n29638 & n29639 ) ;
  assign n29641 = n29609 | n29640 ;
  assign n29642 = n29609 & n29640 ;
  assign n29643 = n29641 & ~n29642 ;
  assign n29644 = n4048 & n25442 ;
  assign n29645 = n4043 & n24324 ;
  assign n29646 = n4045 & n25187 ;
  assign n29647 = n29645 | n29646 ;
  assign n29648 = n29644 | n29647 ;
  assign n29649 = n4051 | n29648 ;
  assign n29650 = ( n25452 & n29648 ) | ( n25452 & n29649 ) | ( n29648 & n29649 ) ;
  assign n29651 = x29 & n29650 ;
  assign n29652 = x29 & ~n29651 ;
  assign n29653 = ( n29650 & ~n29651 ) | ( n29650 & n29652 ) | ( ~n29651 & n29652 ) ;
  assign n29654 = n29643 & n29653 ;
  assign n29655 = n29643 | n29653 ;
  assign n29656 = ~n29654 & n29655 ;
  assign n29657 = ( n29580 & n29608 ) | ( n29580 & ~n29656 ) | ( n29608 & ~n29656 ) ;
  assign n29658 = ( ~n29580 & n29656 ) | ( ~n29580 & n29657 ) | ( n29656 & n29657 ) ;
  assign n29659 = ( ~n29608 & n29657 ) | ( ~n29608 & n29658 ) | ( n29657 & n29658 ) ;
  assign n29660 = ( n29584 & n29598 ) | ( n29584 & ~n29659 ) | ( n29598 & ~n29659 ) ;
  assign n29661 = ( ~n29584 & n29659 ) | ( ~n29584 & n29660 ) | ( n29659 & n29660 ) ;
  assign n29662 = ( ~n29598 & n29660 ) | ( ~n29598 & n29661 ) | ( n29660 & n29661 ) ;
  assign n29663 = n29596 & n29662 ;
  assign n29664 = n29596 & ~n29663 ;
  assign n29665 = ( n29662 & ~n29663 ) | ( n29662 & n29664 ) | ( ~n29663 & n29664 ) ;
  assign n29666 = n29584 & n29659 ;
  assign n29667 = ( n29580 & n29608 ) | ( n29580 & n29656 ) | ( n29608 & n29656 ) ;
  assign n29668 = n24171 & n26156 ;
  assign n29669 = n4479 & n25928 ;
  assign n29670 = n29668 | n29669 ;
  assign n29671 = n4487 | n29670 ;
  assign n29672 = ( n26165 & n29670 ) | ( n26165 & n29671 ) | ( n29670 & n29671 ) ;
  assign n29673 = x26 & n29672 ;
  assign n29674 = x26 & ~n29673 ;
  assign n29675 = ( n29672 & ~n29673 ) | ( n29672 & n29674 ) | ( ~n29673 & n29674 ) ;
  assign n29676 = ( ~n29614 & n29634 ) | ( ~n29614 & n29636 ) | ( n29634 & n29636 ) ;
  assign n29677 = ( ~n29615 & n29636 ) | ( ~n29615 & n29676 ) | ( n29636 & n29676 ) ;
  assign n29678 = n289 | n12291 ;
  assign n29679 = n183 | n29678 ;
  assign n29680 = ~n119 & n616 ;
  assign n29681 = ~n29679 & n29680 ;
  assign n29682 = ( n553 & ~n24164 ) | ( n553 & n29681 ) | ( ~n24164 & n29681 ) ;
  assign n29683 = ~n553 & n29682 ;
  assign n29684 = n29633 & n29683 ;
  assign n29685 = n29633 | n29683 ;
  assign n29686 = ~n29676 & n29685 ;
  assign n29687 = ~n29684 & n29686 ;
  assign n29688 = ~n29636 & n29685 ;
  assign n29689 = ~n29684 & n29688 ;
  assign n29690 = ( n29615 & n29687 ) | ( n29615 & n29689 ) | ( n29687 & n29689 ) ;
  assign n29691 = n29677 | n29690 ;
  assign n29692 = n29685 & ~n29690 ;
  assign n29693 = ~n29684 & n29692 ;
  assign n29694 = n29691 & ~n29693 ;
  assign n29695 = n3744 & n24324 ;
  assign n29696 = n3639 & n24329 ;
  assign n29697 = n3727 & ~n24334 ;
  assign n29698 = n29696 | n29697 ;
  assign n29699 = n29695 | n29698 ;
  assign n29700 = n3636 & ~n24353 ;
  assign n29701 = ( n3636 & n24356 ) | ( n3636 & n29700 ) | ( n24356 & n29700 ) ;
  assign n29702 = n29699 | n29701 ;
  assign n29703 = ~n29694 & n29702 ;
  assign n29704 = n29694 & ~n29702 ;
  assign n29705 = n29703 | n29704 ;
  assign n29706 = n29642 | n29654 ;
  assign n29707 = n29705 & ~n29706 ;
  assign n29708 = ~n29705 & n29706 ;
  assign n29709 = n29707 | n29708 ;
  assign n29710 = n4051 & ~n25690 ;
  assign n29711 = ( n4051 & n25694 ) | ( n4051 & n29710 ) | ( n25694 & n29710 ) ;
  assign n29712 = n4048 & ~n25676 ;
  assign n29713 = n4043 & n25187 ;
  assign n29714 = n4045 & n25442 ;
  assign n29715 = n29713 | n29714 ;
  assign n29716 = n29712 | n29715 ;
  assign n29717 = n29711 | n29716 ;
  assign n29718 = ~x29 & n29717 ;
  assign n29719 = x29 & ~n29717 ;
  assign n29720 = n29718 | n29719 ;
  assign n29721 = ( n29675 & n29709 ) | ( n29675 & ~n29720 ) | ( n29709 & ~n29720 ) ;
  assign n29722 = n29675 & n29720 ;
  assign n29723 = n29675 | n29720 ;
  assign n29724 = ( ~n29709 & n29722 ) | ( ~n29709 & n29723 ) | ( n29722 & n29723 ) ;
  assign n29725 = ( ~n29675 & n29721 ) | ( ~n29675 & n29724 ) | ( n29721 & n29724 ) ;
  assign n29726 = n29667 & ~n29725 ;
  assign n29727 = ~n29667 & n29725 ;
  assign n29728 = n29726 | n29727 ;
  assign n29729 = n29666 & ~n29728 ;
  assign n29730 = n29584 & ~n29666 ;
  assign n29731 = ( n29659 & ~n29728 ) | ( n29659 & n29730 ) | ( ~n29728 & n29730 ) ;
  assign n29732 = ( n29598 & n29729 ) | ( n29598 & n29731 ) | ( n29729 & n29731 ) ;
  assign n29733 = ( n29584 & n29598 ) | ( n29584 & n29659 ) | ( n29598 & n29659 ) ;
  assign n29734 = n29728 & ~n29733 ;
  assign n29735 = n29732 | n29734 ;
  assign n29736 = ~n29663 & n29735 ;
  assign n29737 = n29662 & ~n29735 ;
  assign n29738 = n29596 & n29737 ;
  assign n29739 = n29736 | n29738 ;
  assign n29740 = n666 | n24179 ;
  assign n29741 = n189 | n29740 ;
  assign n29742 = ( x26 & ~n55 ) | ( x26 & n29741 ) | ( ~n55 & n29741 ) ;
  assign n29743 = ~x26 & n29742 ;
  assign n29744 = ( ~n29741 & n29742 ) | ( ~n29741 & n29743 ) | ( n29742 & n29743 ) ;
  assign n29745 = n24173 & n26156 ;
  assign n29746 = ( n29633 & n29744 ) | ( n29633 & n29745 ) | ( n29744 & n29745 ) ;
  assign n29747 = ( n29744 & n29745 ) | ( n29744 & ~n29746 ) | ( n29745 & ~n29746 ) ;
  assign n29748 = ( n29633 & ~n29746 ) | ( n29633 & n29747 ) | ( ~n29746 & n29747 ) ;
  assign n29749 = n3744 & n25187 ;
  assign n29750 = n3639 & ~n24334 ;
  assign n29751 = n3727 & n24324 ;
  assign n29752 = n29750 | n29751 ;
  assign n29753 = n29749 | n29752 ;
  assign n29754 = n3636 | n29753 ;
  assign n29755 = ( n25193 & n29753 ) | ( n25193 & n29754 ) | ( n29753 & n29754 ) ;
  assign n29756 = n4048 & n25928 ;
  assign n29757 = n4043 & n25442 ;
  assign n29758 = n4045 & ~n25676 ;
  assign n29759 = n29757 | n29758 ;
  assign n29760 = n29756 | n29759 ;
  assign n29761 = n4051 | n29760 ;
  assign n29762 = ( ~n25936 & n29760 ) | ( ~n25936 & n29761 ) | ( n29760 & n29761 ) ;
  assign n29763 = n29703 | n29708 ;
  assign n29764 = ( x29 & n29762 ) | ( x29 & ~n29763 ) | ( n29762 & ~n29763 ) ;
  assign n29765 = ( ~x29 & n29763 ) | ( ~x29 & n29764 ) | ( n29763 & n29764 ) ;
  assign n29766 = ( ~n29762 & n29764 ) | ( ~n29762 & n29765 ) | ( n29764 & n29765 ) ;
  assign n29767 = ( ~n29692 & n29755 ) | ( ~n29692 & n29766 ) | ( n29755 & n29766 ) ;
  assign n29768 = ( n29692 & ~n29766 ) | ( n29692 & n29767 ) | ( ~n29766 & n29767 ) ;
  assign n29769 = ( ~n29755 & n29767 ) | ( ~n29755 & n29768 ) | ( n29767 & n29768 ) ;
  assign n29770 = ( ~n29724 & n29748 ) | ( ~n29724 & n29769 ) | ( n29748 & n29769 ) ;
  assign n29771 = ( n29724 & ~n29769 ) | ( n29724 & n29770 ) | ( ~n29769 & n29770 ) ;
  assign n29772 = ( ~n29748 & n29770 ) | ( ~n29748 & n29771 ) | ( n29770 & n29771 ) ;
  assign n29773 = n29726 | n29732 ;
  assign n29774 = ( n29738 & n29772 ) | ( n29738 & ~n29773 ) | ( n29772 & ~n29773 ) ;
  assign n29775 = ( ~n29738 & n29773 ) | ( ~n29738 & n29774 ) | ( n29773 & n29774 ) ;
  assign n29776 = ( ~n29772 & n29774 ) | ( ~n29772 & n29775 ) | ( n29774 & n29775 ) ;
  assign y0 = n24953 ;
  assign y1 = n25214 ;
  assign y2 = ~n25466 ;
  assign y3 = ~n25710 ;
  assign y4 = ~n25955 ;
  assign y5 = ~n26186 ;
  assign y6 = ~n26400 ;
  assign y7 = ~n26602 ;
  assign y8 = n26773 ;
  assign y9 = n26961 ;
  assign y10 = n27147 ;
  assign y11 = n27331 ;
  assign y12 = ~n27535 ;
  assign y13 = ~n27704 ;
  assign y14 = ~n27872 ;
  assign y15 = n28022 ;
  assign y16 = ~n28184 ;
  assign y17 = n28319 ;
  assign y18 = ~n28475 ;
  assign y19 = ~n28607 ;
  assign y20 = ~n28739 ;
  assign y21 = n28866 ;
  assign y22 = n28984 ;
  assign y23 = ~n29096 ;
  assign y24 = ~n29215 ;
  assign y25 = ~n29319 ;
  assign y26 = n29409 ;
  assign y27 = ~n29513 ;
  assign y28 = ~n29597 ;
  assign y29 = n29665 ;
  assign y30 = ~n29739 ;
  assign y31 = n29776 ;
endmodule
